/*
rf_sqrt:
	jxor: 1822
	jspl: 7291
	jspl3: 4814
	jnot: 4227
	jand: 8708
	jor: 6453

Summary:
	jxor: 1822
	jspl: 7291
	jspl3: 4814
	jnot: 4227
	jand: 8708
	jor: 6453

The maximum logic level gap of any gate:
	rf_sqrt: 1
*/

module rf_sqrt(gclk, a, asqrt);
	input gclk;
	input [127:0] a;
	output [63:0] asqrt;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n199;
	wire n200;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n258;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n428;
	wire n429;
	wire n430;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n504;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n593;
	wire n594;
	wire n595;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n687;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n794;
	wire n795;
	wire n796;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n910;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1169;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1472;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1667;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1673;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1684;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1690;
	wire n1691;
	wire n1692;
	wire n1693;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1707;
	wire n1708;
	wire n1709;
	wire n1710;
	wire n1711;
	wire n1712;
	wire n1713;
	wire n1714;
	wire n1715;
	wire n1716;
	wire n1717;
	wire n1718;
	wire n1719;
	wire n1720;
	wire n1721;
	wire n1722;
	wire n1723;
	wire n1724;
	wire n1725;
	wire n1726;
	wire n1727;
	wire n1728;
	wire n1729;
	wire n1730;
	wire n1731;
	wire n1732;
	wire n1733;
	wire n1734;
	wire n1735;
	wire n1736;
	wire n1737;
	wire n1738;
	wire n1739;
	wire n1740;
	wire n1741;
	wire n1742;
	wire n1743;
	wire n1744;
	wire n1745;
	wire n1746;
	wire n1747;
	wire n1748;
	wire n1749;
	wire n1750;
	wire n1751;
	wire n1752;
	wire n1753;
	wire n1754;
	wire n1755;
	wire n1756;
	wire n1757;
	wire n1758;
	wire n1759;
	wire n1760;
	wire n1761;
	wire n1762;
	wire n1763;
	wire n1764;
	wire n1765;
	wire n1766;
	wire n1767;
	wire n1768;
	wire n1769;
	wire n1770;
	wire n1771;
	wire n1772;
	wire n1773;
	wire n1774;
	wire n1775;
	wire n1776;
	wire n1777;
	wire n1778;
	wire n1779;
	wire n1780;
	wire n1781;
	wire n1782;
	wire n1783;
	wire n1784;
	wire n1785;
	wire n1786;
	wire n1787;
	wire n1788;
	wire n1789;
	wire n1790;
	wire n1791;
	wire n1792;
	wire n1793;
	wire n1794;
	wire n1795;
	wire n1796;
	wire n1797;
	wire n1798;
	wire n1799;
	wire n1800;
	wire n1801;
	wire n1802;
	wire n1803;
	wire n1804;
	wire n1805;
	wire n1806;
	wire n1807;
	wire n1808;
	wire n1809;
	wire n1810;
	wire n1811;
	wire n1812;
	wire n1813;
	wire n1814;
	wire n1817;
	wire n1819;
	wire n1820;
	wire n1821;
	wire n1822;
	wire n1823;
	wire n1824;
	wire n1825;
	wire n1826;
	wire n1827;
	wire n1828;
	wire n1829;
	wire n1830;
	wire n1831;
	wire n1832;
	wire n1833;
	wire n1834;
	wire n1835;
	wire n1836;
	wire n1837;
	wire n1838;
	wire n1839;
	wire n1840;
	wire n1841;
	wire n1842;
	wire n1843;
	wire n1844;
	wire n1845;
	wire n1846;
	wire n1847;
	wire n1848;
	wire n1849;
	wire n1850;
	wire n1851;
	wire n1852;
	wire n1853;
	wire n1854;
	wire n1855;
	wire n1856;
	wire n1857;
	wire n1858;
	wire n1859;
	wire n1860;
	wire n1861;
	wire n1862;
	wire n1863;
	wire n1864;
	wire n1865;
	wire n1866;
	wire n1867;
	wire n1868;
	wire n1869;
	wire n1870;
	wire n1871;
	wire n1872;
	wire n1873;
	wire n1874;
	wire n1875;
	wire n1876;
	wire n1877;
	wire n1878;
	wire n1879;
	wire n1880;
	wire n1881;
	wire n1882;
	wire n1883;
	wire n1884;
	wire n1885;
	wire n1886;
	wire n1887;
	wire n1888;
	wire n1889;
	wire n1890;
	wire n1891;
	wire n1892;
	wire n1893;
	wire n1894;
	wire n1895;
	wire n1896;
	wire n1897;
	wire n1898;
	wire n1899;
	wire n1900;
	wire n1901;
	wire n1902;
	wire n1903;
	wire n1904;
	wire n1905;
	wire n1906;
	wire n1907;
	wire n1908;
	wire n1909;
	wire n1910;
	wire n1911;
	wire n1912;
	wire n1913;
	wire n1914;
	wire n1915;
	wire n1916;
	wire n1917;
	wire n1918;
	wire n1919;
	wire n1920;
	wire n1921;
	wire n1922;
	wire n1923;
	wire n1924;
	wire n1925;
	wire n1926;
	wire n1927;
	wire n1928;
	wire n1929;
	wire n1930;
	wire n1931;
	wire n1932;
	wire n1933;
	wire n1934;
	wire n1935;
	wire n1936;
	wire n1937;
	wire n1938;
	wire n1939;
	wire n1940;
	wire n1941;
	wire n1942;
	wire n1943;
	wire n1944;
	wire n1945;
	wire n1946;
	wire n1947;
	wire n1948;
	wire n1949;
	wire n1950;
	wire n1951;
	wire n1952;
	wire n1953;
	wire n1954;
	wire n1955;
	wire n1956;
	wire n1957;
	wire n1958;
	wire n1959;
	wire n1960;
	wire n1961;
	wire n1962;
	wire n1963;
	wire n1964;
	wire n1965;
	wire n1966;
	wire n1967;
	wire n1968;
	wire n1969;
	wire n1970;
	wire n1971;
	wire n1972;
	wire n1973;
	wire n1974;
	wire n1975;
	wire n1976;
	wire n1977;
	wire n1978;
	wire n1979;
	wire n1980;
	wire n1981;
	wire n1982;
	wire n1983;
	wire n1984;
	wire n1985;
	wire n1986;
	wire n1987;
	wire n1988;
	wire n1989;
	wire n1990;
	wire n1991;
	wire n1992;
	wire n1993;
	wire n1994;
	wire n1995;
	wire n1996;
	wire n1997;
	wire n1998;
	wire n1999;
	wire n2000;
	wire n2001;
	wire n2002;
	wire n2003;
	wire n2004;
	wire n2005;
	wire n2008;
	wire n2009;
	wire n2010;
	wire n2012;
	wire n2013;
	wire n2014;
	wire n2015;
	wire n2016;
	wire n2017;
	wire n2018;
	wire n2019;
	wire n2020;
	wire n2021;
	wire n2022;
	wire n2023;
	wire n2024;
	wire n2025;
	wire n2026;
	wire n2027;
	wire n2028;
	wire n2029;
	wire n2030;
	wire n2031;
	wire n2032;
	wire n2033;
	wire n2034;
	wire n2035;
	wire n2036;
	wire n2037;
	wire n2038;
	wire n2039;
	wire n2040;
	wire n2041;
	wire n2042;
	wire n2043;
	wire n2044;
	wire n2045;
	wire n2046;
	wire n2047;
	wire n2048;
	wire n2049;
	wire n2050;
	wire n2051;
	wire n2052;
	wire n2053;
	wire n2054;
	wire n2055;
	wire n2056;
	wire n2057;
	wire n2058;
	wire n2059;
	wire n2060;
	wire n2061;
	wire n2062;
	wire n2063;
	wire n2064;
	wire n2065;
	wire n2066;
	wire n2067;
	wire n2068;
	wire n2069;
	wire n2070;
	wire n2071;
	wire n2072;
	wire n2073;
	wire n2074;
	wire n2075;
	wire n2076;
	wire n2077;
	wire n2078;
	wire n2079;
	wire n2080;
	wire n2081;
	wire n2082;
	wire n2083;
	wire n2084;
	wire n2085;
	wire n2086;
	wire n2087;
	wire n2088;
	wire n2089;
	wire n2090;
	wire n2091;
	wire n2092;
	wire n2093;
	wire n2094;
	wire n2095;
	wire n2096;
	wire n2097;
	wire n2098;
	wire n2099;
	wire n2100;
	wire n2101;
	wire n2102;
	wire n2103;
	wire n2104;
	wire n2105;
	wire n2106;
	wire n2107;
	wire n2108;
	wire n2109;
	wire n2110;
	wire n2111;
	wire n2112;
	wire n2113;
	wire n2114;
	wire n2115;
	wire n2116;
	wire n2117;
	wire n2118;
	wire n2119;
	wire n2120;
	wire n2121;
	wire n2122;
	wire n2123;
	wire n2124;
	wire n2125;
	wire n2126;
	wire n2127;
	wire n2128;
	wire n2129;
	wire n2130;
	wire n2131;
	wire n2132;
	wire n2133;
	wire n2134;
	wire n2135;
	wire n2136;
	wire n2137;
	wire n2138;
	wire n2139;
	wire n2140;
	wire n2141;
	wire n2142;
	wire n2143;
	wire n2144;
	wire n2145;
	wire n2146;
	wire n2147;
	wire n2148;
	wire n2149;
	wire n2150;
	wire n2151;
	wire n2152;
	wire n2153;
	wire n2154;
	wire n2155;
	wire n2156;
	wire n2157;
	wire n2158;
	wire n2159;
	wire n2160;
	wire n2161;
	wire n2162;
	wire n2163;
	wire n2164;
	wire n2165;
	wire n2166;
	wire n2167;
	wire n2168;
	wire n2169;
	wire n2170;
	wire n2171;
	wire n2172;
	wire n2173;
	wire n2174;
	wire n2175;
	wire n2176;
	wire n2177;
	wire n2178;
	wire n2179;
	wire n2180;
	wire n2181;
	wire n2182;
	wire n2183;
	wire n2184;
	wire n2185;
	wire n2186;
	wire n2187;
	wire n2188;
	wire n2189;
	wire n2190;
	wire n2191;
	wire n2192;
	wire n2193;
	wire n2194;
	wire n2195;
	wire n2196;
	wire n2197;
	wire n2198;
	wire n2199;
	wire n2200;
	wire n2201;
	wire n2202;
	wire n2203;
	wire n2206;
	wire n2208;
	wire n2209;
	wire n2210;
	wire n2211;
	wire n2212;
	wire n2213;
	wire n2214;
	wire n2215;
	wire n2216;
	wire n2217;
	wire n2218;
	wire n2219;
	wire n2220;
	wire n2221;
	wire n2222;
	wire n2223;
	wire n2224;
	wire n2225;
	wire n2226;
	wire n2227;
	wire n2228;
	wire n2229;
	wire n2230;
	wire n2231;
	wire n2232;
	wire n2233;
	wire n2234;
	wire n2235;
	wire n2236;
	wire n2237;
	wire n2238;
	wire n2239;
	wire n2240;
	wire n2241;
	wire n2242;
	wire n2243;
	wire n2244;
	wire n2245;
	wire n2246;
	wire n2247;
	wire n2248;
	wire n2249;
	wire n2250;
	wire n2251;
	wire n2252;
	wire n2253;
	wire n2254;
	wire n2255;
	wire n2256;
	wire n2257;
	wire n2258;
	wire n2259;
	wire n2260;
	wire n2261;
	wire n2262;
	wire n2263;
	wire n2264;
	wire n2265;
	wire n2266;
	wire n2267;
	wire n2268;
	wire n2269;
	wire n2270;
	wire n2271;
	wire n2272;
	wire n2273;
	wire n2274;
	wire n2275;
	wire n2276;
	wire n2277;
	wire n2278;
	wire n2279;
	wire n2280;
	wire n2281;
	wire n2282;
	wire n2283;
	wire n2284;
	wire n2285;
	wire n2286;
	wire n2287;
	wire n2288;
	wire n2289;
	wire n2290;
	wire n2291;
	wire n2292;
	wire n2293;
	wire n2294;
	wire n2295;
	wire n2296;
	wire n2297;
	wire n2298;
	wire n2299;
	wire n2300;
	wire n2301;
	wire n2302;
	wire n2303;
	wire n2304;
	wire n2305;
	wire n2306;
	wire n2307;
	wire n2308;
	wire n2309;
	wire n2310;
	wire n2311;
	wire n2312;
	wire n2313;
	wire n2314;
	wire n2315;
	wire n2316;
	wire n2317;
	wire n2318;
	wire n2319;
	wire n2320;
	wire n2321;
	wire n2322;
	wire n2323;
	wire n2324;
	wire n2325;
	wire n2326;
	wire n2327;
	wire n2328;
	wire n2329;
	wire n2330;
	wire n2331;
	wire n2332;
	wire n2333;
	wire n2334;
	wire n2335;
	wire n2336;
	wire n2337;
	wire n2338;
	wire n2339;
	wire n2340;
	wire n2341;
	wire n2342;
	wire n2343;
	wire n2344;
	wire n2345;
	wire n2346;
	wire n2347;
	wire n2348;
	wire n2349;
	wire n2350;
	wire n2351;
	wire n2352;
	wire n2353;
	wire n2354;
	wire n2355;
	wire n2356;
	wire n2357;
	wire n2358;
	wire n2359;
	wire n2360;
	wire n2361;
	wire n2362;
	wire n2363;
	wire n2364;
	wire n2365;
	wire n2366;
	wire n2367;
	wire n2368;
	wire n2369;
	wire n2370;
	wire n2371;
	wire n2372;
	wire n2373;
	wire n2374;
	wire n2375;
	wire n2376;
	wire n2377;
	wire n2378;
	wire n2379;
	wire n2380;
	wire n2381;
	wire n2382;
	wire n2383;
	wire n2384;
	wire n2385;
	wire n2386;
	wire n2387;
	wire n2388;
	wire n2389;
	wire n2390;
	wire n2391;
	wire n2392;
	wire n2393;
	wire n2394;
	wire n2395;
	wire n2396;
	wire n2397;
	wire n2398;
	wire n2399;
	wire n2400;
	wire n2401;
	wire n2402;
	wire n2403;
	wire n2404;
	wire n2405;
	wire n2406;
	wire n2407;
	wire n2408;
	wire n2409;
	wire n2410;
	wire n2411;
	wire n2412;
	wire n2413;
	wire n2414;
	wire n2415;
	wire n2416;
	wire n2417;
	wire n2418;
	wire n2419;
	wire n2420;
	wire n2423;
	wire n2424;
	wire n2425;
	wire n2427;
	wire n2428;
	wire n2429;
	wire n2430;
	wire n2431;
	wire n2432;
	wire n2433;
	wire n2434;
	wire n2435;
	wire n2436;
	wire n2437;
	wire n2438;
	wire n2439;
	wire n2440;
	wire n2441;
	wire n2442;
	wire n2443;
	wire n2444;
	wire n2445;
	wire n2446;
	wire n2447;
	wire n2448;
	wire n2449;
	wire n2450;
	wire n2451;
	wire n2452;
	wire n2453;
	wire n2454;
	wire n2455;
	wire n2456;
	wire n2457;
	wire n2458;
	wire n2459;
	wire n2460;
	wire n2461;
	wire n2462;
	wire n2463;
	wire n2464;
	wire n2465;
	wire n2466;
	wire n2467;
	wire n2468;
	wire n2469;
	wire n2470;
	wire n2471;
	wire n2472;
	wire n2473;
	wire n2474;
	wire n2475;
	wire n2476;
	wire n2477;
	wire n2478;
	wire n2479;
	wire n2480;
	wire n2481;
	wire n2482;
	wire n2483;
	wire n2484;
	wire n2485;
	wire n2486;
	wire n2487;
	wire n2488;
	wire n2489;
	wire n2490;
	wire n2491;
	wire n2492;
	wire n2493;
	wire n2494;
	wire n2495;
	wire n2496;
	wire n2497;
	wire n2498;
	wire n2499;
	wire n2500;
	wire n2501;
	wire n2502;
	wire n2503;
	wire n2504;
	wire n2505;
	wire n2506;
	wire n2507;
	wire n2508;
	wire n2509;
	wire n2510;
	wire n2511;
	wire n2512;
	wire n2513;
	wire n2514;
	wire n2515;
	wire n2516;
	wire n2517;
	wire n2518;
	wire n2519;
	wire n2520;
	wire n2521;
	wire n2522;
	wire n2523;
	wire n2524;
	wire n2525;
	wire n2526;
	wire n2527;
	wire n2528;
	wire n2529;
	wire n2530;
	wire n2531;
	wire n2532;
	wire n2533;
	wire n2534;
	wire n2535;
	wire n2536;
	wire n2537;
	wire n2538;
	wire n2539;
	wire n2540;
	wire n2541;
	wire n2542;
	wire n2543;
	wire n2544;
	wire n2545;
	wire n2546;
	wire n2547;
	wire n2548;
	wire n2549;
	wire n2550;
	wire n2551;
	wire n2552;
	wire n2553;
	wire n2554;
	wire n2555;
	wire n2556;
	wire n2557;
	wire n2558;
	wire n2559;
	wire n2560;
	wire n2561;
	wire n2562;
	wire n2563;
	wire n2564;
	wire n2565;
	wire n2566;
	wire n2567;
	wire n2568;
	wire n2569;
	wire n2570;
	wire n2571;
	wire n2572;
	wire n2573;
	wire n2574;
	wire n2575;
	wire n2576;
	wire n2577;
	wire n2578;
	wire n2579;
	wire n2580;
	wire n2581;
	wire n2582;
	wire n2583;
	wire n2584;
	wire n2585;
	wire n2586;
	wire n2587;
	wire n2588;
	wire n2589;
	wire n2590;
	wire n2591;
	wire n2592;
	wire n2593;
	wire n2594;
	wire n2595;
	wire n2596;
	wire n2597;
	wire n2598;
	wire n2599;
	wire n2600;
	wire n2601;
	wire n2602;
	wire n2603;
	wire n2604;
	wire n2605;
	wire n2606;
	wire n2607;
	wire n2608;
	wire n2609;
	wire n2610;
	wire n2611;
	wire n2612;
	wire n2613;
	wire n2614;
	wire n2615;
	wire n2616;
	wire n2617;
	wire n2618;
	wire n2619;
	wire n2620;
	wire n2621;
	wire n2622;
	wire n2623;
	wire n2624;
	wire n2625;
	wire n2626;
	wire n2627;
	wire n2628;
	wire n2629;
	wire n2630;
	wire n2631;
	wire n2632;
	wire n2633;
	wire n2634;
	wire n2637;
	wire n2639;
	wire n2640;
	wire n2641;
	wire n2642;
	wire n2643;
	wire n2644;
	wire n2645;
	wire n2646;
	wire n2647;
	wire n2648;
	wire n2649;
	wire n2650;
	wire n2651;
	wire n2652;
	wire n2653;
	wire n2654;
	wire n2655;
	wire n2656;
	wire n2657;
	wire n2658;
	wire n2659;
	wire n2660;
	wire n2661;
	wire n2662;
	wire n2663;
	wire n2664;
	wire n2665;
	wire n2666;
	wire n2667;
	wire n2668;
	wire n2669;
	wire n2670;
	wire n2671;
	wire n2672;
	wire n2673;
	wire n2674;
	wire n2675;
	wire n2676;
	wire n2677;
	wire n2678;
	wire n2679;
	wire n2680;
	wire n2681;
	wire n2682;
	wire n2683;
	wire n2684;
	wire n2685;
	wire n2686;
	wire n2687;
	wire n2688;
	wire n2689;
	wire n2690;
	wire n2691;
	wire n2692;
	wire n2693;
	wire n2694;
	wire n2695;
	wire n2696;
	wire n2697;
	wire n2698;
	wire n2699;
	wire n2700;
	wire n2701;
	wire n2702;
	wire n2703;
	wire n2704;
	wire n2705;
	wire n2706;
	wire n2707;
	wire n2708;
	wire n2709;
	wire n2710;
	wire n2711;
	wire n2712;
	wire n2713;
	wire n2714;
	wire n2715;
	wire n2716;
	wire n2717;
	wire n2718;
	wire n2719;
	wire n2720;
	wire n2721;
	wire n2722;
	wire n2723;
	wire n2724;
	wire n2725;
	wire n2726;
	wire n2727;
	wire n2728;
	wire n2729;
	wire n2730;
	wire n2731;
	wire n2732;
	wire n2733;
	wire n2734;
	wire n2735;
	wire n2736;
	wire n2737;
	wire n2738;
	wire n2739;
	wire n2740;
	wire n2741;
	wire n2742;
	wire n2743;
	wire n2744;
	wire n2745;
	wire n2746;
	wire n2747;
	wire n2748;
	wire n2749;
	wire n2750;
	wire n2751;
	wire n2752;
	wire n2753;
	wire n2754;
	wire n2755;
	wire n2756;
	wire n2757;
	wire n2758;
	wire n2759;
	wire n2760;
	wire n2761;
	wire n2762;
	wire n2763;
	wire n2764;
	wire n2765;
	wire n2766;
	wire n2767;
	wire n2768;
	wire n2769;
	wire n2770;
	wire n2771;
	wire n2772;
	wire n2773;
	wire n2774;
	wire n2775;
	wire n2776;
	wire n2777;
	wire n2778;
	wire n2779;
	wire n2780;
	wire n2781;
	wire n2782;
	wire n2783;
	wire n2784;
	wire n2785;
	wire n2786;
	wire n2787;
	wire n2788;
	wire n2789;
	wire n2790;
	wire n2791;
	wire n2792;
	wire n2793;
	wire n2794;
	wire n2795;
	wire n2796;
	wire n2797;
	wire n2798;
	wire n2799;
	wire n2800;
	wire n2801;
	wire n2802;
	wire n2803;
	wire n2804;
	wire n2805;
	wire n2806;
	wire n2807;
	wire n2808;
	wire n2809;
	wire n2810;
	wire n2811;
	wire n2812;
	wire n2813;
	wire n2814;
	wire n2815;
	wire n2816;
	wire n2817;
	wire n2818;
	wire n2819;
	wire n2820;
	wire n2821;
	wire n2822;
	wire n2823;
	wire n2824;
	wire n2825;
	wire n2826;
	wire n2827;
	wire n2828;
	wire n2829;
	wire n2830;
	wire n2831;
	wire n2832;
	wire n2833;
	wire n2834;
	wire n2835;
	wire n2836;
	wire n2837;
	wire n2838;
	wire n2839;
	wire n2840;
	wire n2841;
	wire n2842;
	wire n2843;
	wire n2844;
	wire n2845;
	wire n2846;
	wire n2847;
	wire n2848;
	wire n2849;
	wire n2850;
	wire n2851;
	wire n2852;
	wire n2853;
	wire n2854;
	wire n2855;
	wire n2856;
	wire n2857;
	wire n2858;
	wire n2859;
	wire n2860;
	wire n2861;
	wire n2862;
	wire n2863;
	wire n2864;
	wire n2865;
	wire n2866;
	wire n2867;
	wire n2868;
	wire n2869;
	wire n2870;
	wire n2873;
	wire n2874;
	wire n2875;
	wire n2877;
	wire n2878;
	wire n2879;
	wire n2880;
	wire n2881;
	wire n2882;
	wire n2883;
	wire n2884;
	wire n2885;
	wire n2886;
	wire n2887;
	wire n2888;
	wire n2889;
	wire n2890;
	wire n2891;
	wire n2892;
	wire n2893;
	wire n2894;
	wire n2895;
	wire n2896;
	wire n2897;
	wire n2898;
	wire n2899;
	wire n2900;
	wire n2901;
	wire n2902;
	wire n2903;
	wire n2904;
	wire n2905;
	wire n2906;
	wire n2907;
	wire n2908;
	wire n2909;
	wire n2910;
	wire n2911;
	wire n2912;
	wire n2913;
	wire n2914;
	wire n2915;
	wire n2916;
	wire n2917;
	wire n2918;
	wire n2919;
	wire n2920;
	wire n2921;
	wire n2922;
	wire n2923;
	wire n2924;
	wire n2925;
	wire n2926;
	wire n2927;
	wire n2928;
	wire n2929;
	wire n2930;
	wire n2931;
	wire n2932;
	wire n2933;
	wire n2934;
	wire n2935;
	wire n2936;
	wire n2937;
	wire n2938;
	wire n2939;
	wire n2940;
	wire n2941;
	wire n2942;
	wire n2943;
	wire n2944;
	wire n2945;
	wire n2946;
	wire n2947;
	wire n2948;
	wire n2949;
	wire n2950;
	wire n2951;
	wire n2952;
	wire n2953;
	wire n2954;
	wire n2955;
	wire n2956;
	wire n2957;
	wire n2958;
	wire n2959;
	wire n2960;
	wire n2961;
	wire n2962;
	wire n2963;
	wire n2964;
	wire n2965;
	wire n2966;
	wire n2967;
	wire n2968;
	wire n2969;
	wire n2970;
	wire n2971;
	wire n2972;
	wire n2973;
	wire n2974;
	wire n2975;
	wire n2976;
	wire n2977;
	wire n2978;
	wire n2979;
	wire n2980;
	wire n2981;
	wire n2982;
	wire n2983;
	wire n2984;
	wire n2985;
	wire n2986;
	wire n2987;
	wire n2988;
	wire n2989;
	wire n2990;
	wire n2991;
	wire n2992;
	wire n2993;
	wire n2994;
	wire n2995;
	wire n2996;
	wire n2997;
	wire n2998;
	wire n2999;
	wire n3000;
	wire n3001;
	wire n3002;
	wire n3003;
	wire n3004;
	wire n3005;
	wire n3006;
	wire n3007;
	wire n3008;
	wire n3009;
	wire n3010;
	wire n3011;
	wire n3012;
	wire n3013;
	wire n3014;
	wire n3015;
	wire n3016;
	wire n3017;
	wire n3018;
	wire n3019;
	wire n3020;
	wire n3021;
	wire n3022;
	wire n3023;
	wire n3024;
	wire n3025;
	wire n3026;
	wire n3027;
	wire n3028;
	wire n3029;
	wire n3030;
	wire n3031;
	wire n3032;
	wire n3033;
	wire n3034;
	wire n3035;
	wire n3036;
	wire n3037;
	wire n3038;
	wire n3039;
	wire n3040;
	wire n3041;
	wire n3042;
	wire n3043;
	wire n3044;
	wire n3045;
	wire n3046;
	wire n3047;
	wire n3048;
	wire n3049;
	wire n3050;
	wire n3051;
	wire n3052;
	wire n3053;
	wire n3054;
	wire n3055;
	wire n3056;
	wire n3057;
	wire n3058;
	wire n3059;
	wire n3060;
	wire n3061;
	wire n3062;
	wire n3063;
	wire n3064;
	wire n3065;
	wire n3066;
	wire n3067;
	wire n3068;
	wire n3069;
	wire n3070;
	wire n3071;
	wire n3072;
	wire n3073;
	wire n3074;
	wire n3075;
	wire n3076;
	wire n3077;
	wire n3078;
	wire n3079;
	wire n3080;
	wire n3081;
	wire n3082;
	wire n3083;
	wire n3084;
	wire n3085;
	wire n3086;
	wire n3087;
	wire n3088;
	wire n3089;
	wire n3090;
	wire n3091;
	wire n3092;
	wire n3093;
	wire n3094;
	wire n3095;
	wire n3096;
	wire n3097;
	wire n3098;
	wire n3099;
	wire n3100;
	wire n3101;
	wire n3102;
	wire n3103;
	wire n3104;
	wire n3105;
	wire n3106;
	wire n3107;
	wire n3108;
	wire n3109;
	wire n3112;
	wire n3114;
	wire n3115;
	wire n3116;
	wire n3117;
	wire n3118;
	wire n3119;
	wire n3120;
	wire n3121;
	wire n3122;
	wire n3123;
	wire n3124;
	wire n3125;
	wire n3126;
	wire n3127;
	wire n3128;
	wire n3129;
	wire n3130;
	wire n3131;
	wire n3132;
	wire n3133;
	wire n3134;
	wire n3135;
	wire n3136;
	wire n3137;
	wire n3138;
	wire n3139;
	wire n3140;
	wire n3141;
	wire n3142;
	wire n3143;
	wire n3144;
	wire n3145;
	wire n3146;
	wire n3147;
	wire n3148;
	wire n3149;
	wire n3150;
	wire n3151;
	wire n3152;
	wire n3153;
	wire n3154;
	wire n3155;
	wire n3156;
	wire n3157;
	wire n3158;
	wire n3159;
	wire n3160;
	wire n3161;
	wire n3162;
	wire n3163;
	wire n3164;
	wire n3165;
	wire n3166;
	wire n3167;
	wire n3168;
	wire n3169;
	wire n3170;
	wire n3171;
	wire n3172;
	wire n3173;
	wire n3174;
	wire n3175;
	wire n3176;
	wire n3177;
	wire n3178;
	wire n3179;
	wire n3180;
	wire n3181;
	wire n3182;
	wire n3183;
	wire n3184;
	wire n3185;
	wire n3186;
	wire n3187;
	wire n3188;
	wire n3189;
	wire n3190;
	wire n3191;
	wire n3192;
	wire n3193;
	wire n3194;
	wire n3195;
	wire n3196;
	wire n3197;
	wire n3198;
	wire n3199;
	wire n3200;
	wire n3201;
	wire n3202;
	wire n3203;
	wire n3204;
	wire n3205;
	wire n3206;
	wire n3207;
	wire n3208;
	wire n3209;
	wire n3210;
	wire n3211;
	wire n3212;
	wire n3213;
	wire n3214;
	wire n3215;
	wire n3216;
	wire n3217;
	wire n3218;
	wire n3219;
	wire n3220;
	wire n3221;
	wire n3222;
	wire n3223;
	wire n3224;
	wire n3225;
	wire n3226;
	wire n3227;
	wire n3228;
	wire n3229;
	wire n3230;
	wire n3231;
	wire n3232;
	wire n3233;
	wire n3234;
	wire n3235;
	wire n3236;
	wire n3237;
	wire n3238;
	wire n3239;
	wire n3240;
	wire n3241;
	wire n3242;
	wire n3243;
	wire n3244;
	wire n3245;
	wire n3246;
	wire n3247;
	wire n3248;
	wire n3249;
	wire n3250;
	wire n3251;
	wire n3252;
	wire n3253;
	wire n3254;
	wire n3255;
	wire n3256;
	wire n3257;
	wire n3258;
	wire n3259;
	wire n3260;
	wire n3261;
	wire n3262;
	wire n3263;
	wire n3264;
	wire n3265;
	wire n3266;
	wire n3267;
	wire n3268;
	wire n3269;
	wire n3270;
	wire n3271;
	wire n3272;
	wire n3273;
	wire n3274;
	wire n3275;
	wire n3276;
	wire n3277;
	wire n3278;
	wire n3279;
	wire n3280;
	wire n3281;
	wire n3282;
	wire n3283;
	wire n3284;
	wire n3285;
	wire n3286;
	wire n3287;
	wire n3288;
	wire n3289;
	wire n3290;
	wire n3291;
	wire n3292;
	wire n3293;
	wire n3294;
	wire n3295;
	wire n3296;
	wire n3297;
	wire n3298;
	wire n3299;
	wire n3300;
	wire n3301;
	wire n3302;
	wire n3303;
	wire n3304;
	wire n3305;
	wire n3306;
	wire n3307;
	wire n3308;
	wire n3309;
	wire n3310;
	wire n3311;
	wire n3312;
	wire n3313;
	wire n3314;
	wire n3315;
	wire n3316;
	wire n3317;
	wire n3318;
	wire n3319;
	wire n3320;
	wire n3321;
	wire n3322;
	wire n3323;
	wire n3324;
	wire n3325;
	wire n3326;
	wire n3327;
	wire n3328;
	wire n3329;
	wire n3330;
	wire n3331;
	wire n3332;
	wire n3333;
	wire n3334;
	wire n3335;
	wire n3336;
	wire n3337;
	wire n3338;
	wire n3339;
	wire n3340;
	wire n3341;
	wire n3342;
	wire n3343;
	wire n3344;
	wire n3345;
	wire n3346;
	wire n3347;
	wire n3348;
	wire n3349;
	wire n3350;
	wire n3351;
	wire n3352;
	wire n3353;
	wire n3354;
	wire n3355;
	wire n3356;
	wire n3357;
	wire n3358;
	wire n3359;
	wire n3360;
	wire n3361;
	wire n3362;
	wire n3363;
	wire n3364;
	wire n3365;
	wire n3366;
	wire n3367;
	wire n3368;
	wire n3369;
	wire n3370;
	wire n3371;
	wire n3374;
	wire n3375;
	wire n3376;
	wire n3378;
	wire n3379;
	wire n3380;
	wire n3381;
	wire n3382;
	wire n3383;
	wire n3384;
	wire n3385;
	wire n3386;
	wire n3387;
	wire n3388;
	wire n3389;
	wire n3390;
	wire n3391;
	wire n3392;
	wire n3393;
	wire n3394;
	wire n3395;
	wire n3396;
	wire n3397;
	wire n3398;
	wire n3399;
	wire n3400;
	wire n3401;
	wire n3402;
	wire n3403;
	wire n3404;
	wire n3405;
	wire n3406;
	wire n3407;
	wire n3408;
	wire n3409;
	wire n3410;
	wire n3411;
	wire n3412;
	wire n3413;
	wire n3414;
	wire n3415;
	wire n3416;
	wire n3417;
	wire n3418;
	wire n3419;
	wire n3420;
	wire n3421;
	wire n3422;
	wire n3423;
	wire n3424;
	wire n3425;
	wire n3426;
	wire n3427;
	wire n3428;
	wire n3429;
	wire n3430;
	wire n3431;
	wire n3432;
	wire n3433;
	wire n3434;
	wire n3435;
	wire n3436;
	wire n3437;
	wire n3438;
	wire n3439;
	wire n3440;
	wire n3441;
	wire n3442;
	wire n3443;
	wire n3444;
	wire n3445;
	wire n3446;
	wire n3447;
	wire n3448;
	wire n3449;
	wire n3450;
	wire n3451;
	wire n3452;
	wire n3453;
	wire n3454;
	wire n3455;
	wire n3456;
	wire n3457;
	wire n3458;
	wire n3459;
	wire n3460;
	wire n3461;
	wire n3462;
	wire n3463;
	wire n3464;
	wire n3465;
	wire n3466;
	wire n3467;
	wire n3468;
	wire n3469;
	wire n3470;
	wire n3471;
	wire n3472;
	wire n3473;
	wire n3474;
	wire n3475;
	wire n3476;
	wire n3477;
	wire n3478;
	wire n3479;
	wire n3480;
	wire n3481;
	wire n3482;
	wire n3483;
	wire n3484;
	wire n3485;
	wire n3486;
	wire n3487;
	wire n3488;
	wire n3489;
	wire n3490;
	wire n3491;
	wire n3492;
	wire n3493;
	wire n3494;
	wire n3495;
	wire n3496;
	wire n3497;
	wire n3498;
	wire n3499;
	wire n3500;
	wire n3501;
	wire n3502;
	wire n3503;
	wire n3504;
	wire n3505;
	wire n3506;
	wire n3507;
	wire n3508;
	wire n3509;
	wire n3510;
	wire n3511;
	wire n3512;
	wire n3513;
	wire n3514;
	wire n3515;
	wire n3516;
	wire n3517;
	wire n3518;
	wire n3519;
	wire n3520;
	wire n3521;
	wire n3522;
	wire n3523;
	wire n3524;
	wire n3525;
	wire n3526;
	wire n3527;
	wire n3528;
	wire n3529;
	wire n3530;
	wire n3531;
	wire n3532;
	wire n3533;
	wire n3534;
	wire n3535;
	wire n3536;
	wire n3537;
	wire n3538;
	wire n3539;
	wire n3540;
	wire n3541;
	wire n3542;
	wire n3543;
	wire n3544;
	wire n3545;
	wire n3546;
	wire n3547;
	wire n3548;
	wire n3549;
	wire n3550;
	wire n3551;
	wire n3552;
	wire n3553;
	wire n3554;
	wire n3555;
	wire n3556;
	wire n3557;
	wire n3558;
	wire n3559;
	wire n3560;
	wire n3561;
	wire n3562;
	wire n3563;
	wire n3564;
	wire n3565;
	wire n3566;
	wire n3567;
	wire n3568;
	wire n3569;
	wire n3570;
	wire n3571;
	wire n3572;
	wire n3573;
	wire n3574;
	wire n3575;
	wire n3576;
	wire n3577;
	wire n3578;
	wire n3579;
	wire n3580;
	wire n3581;
	wire n3582;
	wire n3583;
	wire n3584;
	wire n3585;
	wire n3586;
	wire n3587;
	wire n3588;
	wire n3589;
	wire n3590;
	wire n3591;
	wire n3592;
	wire n3593;
	wire n3594;
	wire n3595;
	wire n3596;
	wire n3597;
	wire n3598;
	wire n3599;
	wire n3600;
	wire n3601;
	wire n3602;
	wire n3603;
	wire n3604;
	wire n3605;
	wire n3606;
	wire n3607;
	wire n3608;
	wire n3609;
	wire n3610;
	wire n3611;
	wire n3612;
	wire n3613;
	wire n3614;
	wire n3615;
	wire n3616;
	wire n3617;
	wire n3618;
	wire n3619;
	wire n3620;
	wire n3621;
	wire n3622;
	wire n3623;
	wire n3624;
	wire n3625;
	wire n3626;
	wire n3629;
	wire n3631;
	wire n3632;
	wire n3633;
	wire n3634;
	wire n3635;
	wire n3636;
	wire n3637;
	wire n3638;
	wire n3639;
	wire n3640;
	wire n3641;
	wire n3642;
	wire n3643;
	wire n3644;
	wire n3645;
	wire n3646;
	wire n3647;
	wire n3648;
	wire n3649;
	wire n3650;
	wire n3651;
	wire n3652;
	wire n3653;
	wire n3654;
	wire n3655;
	wire n3656;
	wire n3657;
	wire n3658;
	wire n3659;
	wire n3660;
	wire n3661;
	wire n3662;
	wire n3663;
	wire n3664;
	wire n3665;
	wire n3666;
	wire n3667;
	wire n3668;
	wire n3669;
	wire n3670;
	wire n3671;
	wire n3672;
	wire n3673;
	wire n3674;
	wire n3675;
	wire n3676;
	wire n3677;
	wire n3678;
	wire n3679;
	wire n3680;
	wire n3681;
	wire n3682;
	wire n3683;
	wire n3684;
	wire n3685;
	wire n3686;
	wire n3687;
	wire n3688;
	wire n3689;
	wire n3690;
	wire n3691;
	wire n3692;
	wire n3693;
	wire n3694;
	wire n3695;
	wire n3696;
	wire n3697;
	wire n3698;
	wire n3699;
	wire n3700;
	wire n3701;
	wire n3702;
	wire n3703;
	wire n3704;
	wire n3705;
	wire n3706;
	wire n3707;
	wire n3708;
	wire n3709;
	wire n3710;
	wire n3711;
	wire n3712;
	wire n3713;
	wire n3714;
	wire n3715;
	wire n3716;
	wire n3717;
	wire n3718;
	wire n3719;
	wire n3720;
	wire n3721;
	wire n3722;
	wire n3723;
	wire n3724;
	wire n3725;
	wire n3726;
	wire n3727;
	wire n3728;
	wire n3729;
	wire n3730;
	wire n3731;
	wire n3732;
	wire n3733;
	wire n3734;
	wire n3735;
	wire n3736;
	wire n3737;
	wire n3738;
	wire n3739;
	wire n3740;
	wire n3741;
	wire n3742;
	wire n3743;
	wire n3744;
	wire n3745;
	wire n3746;
	wire n3747;
	wire n3748;
	wire n3749;
	wire n3750;
	wire n3751;
	wire n3752;
	wire n3753;
	wire n3754;
	wire n3755;
	wire n3756;
	wire n3757;
	wire n3758;
	wire n3759;
	wire n3760;
	wire n3761;
	wire n3762;
	wire n3763;
	wire n3764;
	wire n3765;
	wire n3766;
	wire n3767;
	wire n3768;
	wire n3769;
	wire n3770;
	wire n3771;
	wire n3772;
	wire n3773;
	wire n3774;
	wire n3775;
	wire n3776;
	wire n3777;
	wire n3778;
	wire n3779;
	wire n3780;
	wire n3781;
	wire n3782;
	wire n3783;
	wire n3784;
	wire n3785;
	wire n3786;
	wire n3787;
	wire n3788;
	wire n3789;
	wire n3790;
	wire n3791;
	wire n3792;
	wire n3793;
	wire n3794;
	wire n3795;
	wire n3796;
	wire n3797;
	wire n3798;
	wire n3799;
	wire n3800;
	wire n3801;
	wire n3802;
	wire n3803;
	wire n3804;
	wire n3805;
	wire n3806;
	wire n3807;
	wire n3808;
	wire n3809;
	wire n3810;
	wire n3811;
	wire n3812;
	wire n3813;
	wire n3814;
	wire n3815;
	wire n3816;
	wire n3817;
	wire n3818;
	wire n3819;
	wire n3820;
	wire n3821;
	wire n3822;
	wire n3823;
	wire n3824;
	wire n3825;
	wire n3826;
	wire n3827;
	wire n3828;
	wire n3829;
	wire n3830;
	wire n3831;
	wire n3832;
	wire n3833;
	wire n3834;
	wire n3835;
	wire n3836;
	wire n3837;
	wire n3838;
	wire n3839;
	wire n3840;
	wire n3841;
	wire n3842;
	wire n3843;
	wire n3844;
	wire n3845;
	wire n3846;
	wire n3847;
	wire n3848;
	wire n3849;
	wire n3850;
	wire n3851;
	wire n3852;
	wire n3853;
	wire n3854;
	wire n3855;
	wire n3856;
	wire n3857;
	wire n3858;
	wire n3859;
	wire n3860;
	wire n3861;
	wire n3862;
	wire n3863;
	wire n3864;
	wire n3865;
	wire n3866;
	wire n3867;
	wire n3868;
	wire n3869;
	wire n3870;
	wire n3871;
	wire n3872;
	wire n3873;
	wire n3874;
	wire n3875;
	wire n3876;
	wire n3877;
	wire n3878;
	wire n3879;
	wire n3880;
	wire n3881;
	wire n3882;
	wire n3883;
	wire n3884;
	wire n3885;
	wire n3886;
	wire n3887;
	wire n3888;
	wire n3889;
	wire n3890;
	wire n3891;
	wire n3892;
	wire n3893;
	wire n3894;
	wire n3895;
	wire n3896;
	wire n3897;
	wire n3898;
	wire n3899;
	wire n3900;
	wire n3901;
	wire n3902;
	wire n3903;
	wire n3904;
	wire n3905;
	wire n3906;
	wire n3907;
	wire n3910;
	wire n3911;
	wire n3912;
	wire n3914;
	wire n3915;
	wire n3916;
	wire n3917;
	wire n3918;
	wire n3919;
	wire n3920;
	wire n3921;
	wire n3922;
	wire n3923;
	wire n3924;
	wire n3925;
	wire n3926;
	wire n3927;
	wire n3928;
	wire n3929;
	wire n3930;
	wire n3931;
	wire n3932;
	wire n3933;
	wire n3934;
	wire n3935;
	wire n3936;
	wire n3937;
	wire n3938;
	wire n3939;
	wire n3940;
	wire n3941;
	wire n3942;
	wire n3943;
	wire n3944;
	wire n3945;
	wire n3946;
	wire n3947;
	wire n3948;
	wire n3949;
	wire n3950;
	wire n3951;
	wire n3952;
	wire n3953;
	wire n3954;
	wire n3955;
	wire n3956;
	wire n3957;
	wire n3958;
	wire n3959;
	wire n3960;
	wire n3961;
	wire n3962;
	wire n3963;
	wire n3964;
	wire n3965;
	wire n3966;
	wire n3967;
	wire n3968;
	wire n3969;
	wire n3970;
	wire n3971;
	wire n3972;
	wire n3973;
	wire n3974;
	wire n3975;
	wire n3976;
	wire n3977;
	wire n3978;
	wire n3979;
	wire n3980;
	wire n3981;
	wire n3982;
	wire n3983;
	wire n3984;
	wire n3985;
	wire n3986;
	wire n3987;
	wire n3988;
	wire n3989;
	wire n3990;
	wire n3991;
	wire n3992;
	wire n3993;
	wire n3994;
	wire n3995;
	wire n3996;
	wire n3997;
	wire n3998;
	wire n3999;
	wire n4000;
	wire n4001;
	wire n4002;
	wire n4003;
	wire n4004;
	wire n4005;
	wire n4006;
	wire n4007;
	wire n4008;
	wire n4009;
	wire n4010;
	wire n4011;
	wire n4012;
	wire n4013;
	wire n4014;
	wire n4015;
	wire n4016;
	wire n4017;
	wire n4018;
	wire n4019;
	wire n4020;
	wire n4021;
	wire n4022;
	wire n4023;
	wire n4024;
	wire n4025;
	wire n4026;
	wire n4027;
	wire n4028;
	wire n4029;
	wire n4030;
	wire n4031;
	wire n4032;
	wire n4033;
	wire n4034;
	wire n4035;
	wire n4036;
	wire n4037;
	wire n4038;
	wire n4039;
	wire n4040;
	wire n4041;
	wire n4042;
	wire n4043;
	wire n4044;
	wire n4045;
	wire n4046;
	wire n4047;
	wire n4048;
	wire n4049;
	wire n4050;
	wire n4051;
	wire n4052;
	wire n4053;
	wire n4054;
	wire n4055;
	wire n4056;
	wire n4057;
	wire n4058;
	wire n4059;
	wire n4060;
	wire n4061;
	wire n4062;
	wire n4063;
	wire n4064;
	wire n4065;
	wire n4066;
	wire n4067;
	wire n4068;
	wire n4069;
	wire n4070;
	wire n4071;
	wire n4072;
	wire n4073;
	wire n4074;
	wire n4075;
	wire n4076;
	wire n4077;
	wire n4078;
	wire n4079;
	wire n4080;
	wire n4081;
	wire n4082;
	wire n4083;
	wire n4084;
	wire n4085;
	wire n4086;
	wire n4087;
	wire n4088;
	wire n4089;
	wire n4090;
	wire n4091;
	wire n4092;
	wire n4093;
	wire n4094;
	wire n4095;
	wire n4096;
	wire n4097;
	wire n4098;
	wire n4099;
	wire n4100;
	wire n4101;
	wire n4102;
	wire n4103;
	wire n4104;
	wire n4105;
	wire n4106;
	wire n4107;
	wire n4108;
	wire n4109;
	wire n4110;
	wire n4111;
	wire n4112;
	wire n4113;
	wire n4114;
	wire n4115;
	wire n4116;
	wire n4117;
	wire n4118;
	wire n4119;
	wire n4120;
	wire n4121;
	wire n4122;
	wire n4123;
	wire n4124;
	wire n4125;
	wire n4126;
	wire n4127;
	wire n4128;
	wire n4129;
	wire n4130;
	wire n4131;
	wire n4132;
	wire n4133;
	wire n4134;
	wire n4135;
	wire n4136;
	wire n4137;
	wire n4138;
	wire n4139;
	wire n4140;
	wire n4141;
	wire n4142;
	wire n4143;
	wire n4144;
	wire n4145;
	wire n4146;
	wire n4147;
	wire n4148;
	wire n4149;
	wire n4150;
	wire n4151;
	wire n4152;
	wire n4153;
	wire n4154;
	wire n4155;
	wire n4156;
	wire n4157;
	wire n4158;
	wire n4159;
	wire n4160;
	wire n4161;
	wire n4162;
	wire n4163;
	wire n4164;
	wire n4165;
	wire n4166;
	wire n4167;
	wire n4168;
	wire n4169;
	wire n4170;
	wire n4171;
	wire n4172;
	wire n4173;
	wire n4174;
	wire n4175;
	wire n4176;
	wire n4177;
	wire n4178;
	wire n4179;
	wire n4180;
	wire n4181;
	wire n4182;
	wire n4183;
	wire n4184;
	wire n4185;
	wire n4186;
	wire n4187;
	wire n4190;
	wire n4192;
	wire n4193;
	wire n4194;
	wire n4195;
	wire n4196;
	wire n4197;
	wire n4198;
	wire n4199;
	wire n4200;
	wire n4201;
	wire n4202;
	wire n4203;
	wire n4204;
	wire n4205;
	wire n4206;
	wire n4207;
	wire n4208;
	wire n4209;
	wire n4210;
	wire n4211;
	wire n4212;
	wire n4213;
	wire n4214;
	wire n4215;
	wire n4216;
	wire n4217;
	wire n4218;
	wire n4219;
	wire n4220;
	wire n4221;
	wire n4222;
	wire n4223;
	wire n4224;
	wire n4225;
	wire n4226;
	wire n4227;
	wire n4228;
	wire n4229;
	wire n4230;
	wire n4231;
	wire n4232;
	wire n4233;
	wire n4234;
	wire n4235;
	wire n4236;
	wire n4237;
	wire n4238;
	wire n4239;
	wire n4240;
	wire n4241;
	wire n4242;
	wire n4243;
	wire n4244;
	wire n4245;
	wire n4246;
	wire n4247;
	wire n4248;
	wire n4249;
	wire n4250;
	wire n4251;
	wire n4252;
	wire n4253;
	wire n4254;
	wire n4255;
	wire n4256;
	wire n4257;
	wire n4258;
	wire n4259;
	wire n4260;
	wire n4261;
	wire n4262;
	wire n4263;
	wire n4264;
	wire n4265;
	wire n4266;
	wire n4267;
	wire n4268;
	wire n4269;
	wire n4270;
	wire n4271;
	wire n4272;
	wire n4273;
	wire n4274;
	wire n4275;
	wire n4276;
	wire n4277;
	wire n4278;
	wire n4279;
	wire n4280;
	wire n4281;
	wire n4282;
	wire n4283;
	wire n4284;
	wire n4285;
	wire n4286;
	wire n4287;
	wire n4288;
	wire n4289;
	wire n4290;
	wire n4291;
	wire n4292;
	wire n4293;
	wire n4294;
	wire n4295;
	wire n4296;
	wire n4297;
	wire n4298;
	wire n4299;
	wire n4300;
	wire n4301;
	wire n4302;
	wire n4303;
	wire n4304;
	wire n4305;
	wire n4306;
	wire n4307;
	wire n4308;
	wire n4309;
	wire n4310;
	wire n4311;
	wire n4312;
	wire n4313;
	wire n4314;
	wire n4315;
	wire n4316;
	wire n4317;
	wire n4318;
	wire n4319;
	wire n4320;
	wire n4321;
	wire n4322;
	wire n4323;
	wire n4324;
	wire n4325;
	wire n4326;
	wire n4327;
	wire n4328;
	wire n4329;
	wire n4330;
	wire n4331;
	wire n4332;
	wire n4333;
	wire n4334;
	wire n4335;
	wire n4336;
	wire n4337;
	wire n4338;
	wire n4339;
	wire n4340;
	wire n4341;
	wire n4342;
	wire n4343;
	wire n4344;
	wire n4345;
	wire n4346;
	wire n4347;
	wire n4348;
	wire n4349;
	wire n4350;
	wire n4351;
	wire n4352;
	wire n4353;
	wire n4354;
	wire n4355;
	wire n4356;
	wire n4357;
	wire n4358;
	wire n4359;
	wire n4360;
	wire n4361;
	wire n4362;
	wire n4363;
	wire n4364;
	wire n4365;
	wire n4366;
	wire n4367;
	wire n4368;
	wire n4369;
	wire n4370;
	wire n4371;
	wire n4372;
	wire n4373;
	wire n4374;
	wire n4375;
	wire n4376;
	wire n4377;
	wire n4378;
	wire n4379;
	wire n4380;
	wire n4381;
	wire n4382;
	wire n4383;
	wire n4384;
	wire n4385;
	wire n4386;
	wire n4387;
	wire n4388;
	wire n4389;
	wire n4390;
	wire n4391;
	wire n4392;
	wire n4393;
	wire n4394;
	wire n4395;
	wire n4396;
	wire n4397;
	wire n4398;
	wire n4399;
	wire n4400;
	wire n4401;
	wire n4402;
	wire n4403;
	wire n4404;
	wire n4405;
	wire n4406;
	wire n4407;
	wire n4408;
	wire n4409;
	wire n4410;
	wire n4411;
	wire n4412;
	wire n4413;
	wire n4414;
	wire n4415;
	wire n4416;
	wire n4417;
	wire n4418;
	wire n4419;
	wire n4420;
	wire n4421;
	wire n4422;
	wire n4423;
	wire n4424;
	wire n4425;
	wire n4426;
	wire n4427;
	wire n4428;
	wire n4429;
	wire n4430;
	wire n4431;
	wire n4432;
	wire n4433;
	wire n4434;
	wire n4435;
	wire n4436;
	wire n4437;
	wire n4438;
	wire n4439;
	wire n4440;
	wire n4441;
	wire n4442;
	wire n4443;
	wire n4444;
	wire n4445;
	wire n4446;
	wire n4447;
	wire n4448;
	wire n4449;
	wire n4450;
	wire n4451;
	wire n4452;
	wire n4453;
	wire n4454;
	wire n4455;
	wire n4456;
	wire n4457;
	wire n4458;
	wire n4459;
	wire n4460;
	wire n4461;
	wire n4462;
	wire n4463;
	wire n4464;
	wire n4465;
	wire n4466;
	wire n4467;
	wire n4468;
	wire n4469;
	wire n4470;
	wire n4471;
	wire n4472;
	wire n4473;
	wire n4474;
	wire n4475;
	wire n4476;
	wire n4477;
	wire n4478;
	wire n4479;
	wire n4480;
	wire n4481;
	wire n4482;
	wire n4483;
	wire n4484;
	wire n4485;
	wire n4486;
	wire n4487;
	wire n4488;
	wire n4489;
	wire n4490;
	wire n4491;
	wire n4492;
	wire n4493;
	wire n4494;
	wire n4497;
	wire n4498;
	wire n4499;
	wire n4501;
	wire n4502;
	wire n4503;
	wire n4504;
	wire n4505;
	wire n4506;
	wire n4507;
	wire n4508;
	wire n4509;
	wire n4510;
	wire n4511;
	wire n4512;
	wire n4513;
	wire n4514;
	wire n4515;
	wire n4516;
	wire n4517;
	wire n4518;
	wire n4519;
	wire n4520;
	wire n4521;
	wire n4522;
	wire n4523;
	wire n4524;
	wire n4525;
	wire n4526;
	wire n4527;
	wire n4528;
	wire n4529;
	wire n4530;
	wire n4531;
	wire n4532;
	wire n4533;
	wire n4534;
	wire n4535;
	wire n4536;
	wire n4537;
	wire n4538;
	wire n4539;
	wire n4540;
	wire n4541;
	wire n4542;
	wire n4543;
	wire n4544;
	wire n4545;
	wire n4546;
	wire n4547;
	wire n4548;
	wire n4549;
	wire n4550;
	wire n4551;
	wire n4552;
	wire n4553;
	wire n4554;
	wire n4555;
	wire n4556;
	wire n4557;
	wire n4558;
	wire n4559;
	wire n4560;
	wire n4561;
	wire n4562;
	wire n4563;
	wire n4564;
	wire n4565;
	wire n4566;
	wire n4567;
	wire n4568;
	wire n4569;
	wire n4570;
	wire n4571;
	wire n4572;
	wire n4573;
	wire n4574;
	wire n4575;
	wire n4576;
	wire n4577;
	wire n4578;
	wire n4579;
	wire n4580;
	wire n4581;
	wire n4582;
	wire n4583;
	wire n4584;
	wire n4585;
	wire n4586;
	wire n4587;
	wire n4588;
	wire n4589;
	wire n4590;
	wire n4591;
	wire n4592;
	wire n4593;
	wire n4594;
	wire n4595;
	wire n4596;
	wire n4597;
	wire n4598;
	wire n4599;
	wire n4600;
	wire n4601;
	wire n4602;
	wire n4603;
	wire n4604;
	wire n4605;
	wire n4606;
	wire n4607;
	wire n4608;
	wire n4609;
	wire n4610;
	wire n4611;
	wire n4612;
	wire n4613;
	wire n4614;
	wire n4615;
	wire n4616;
	wire n4617;
	wire n4618;
	wire n4619;
	wire n4620;
	wire n4621;
	wire n4622;
	wire n4623;
	wire n4624;
	wire n4625;
	wire n4626;
	wire n4627;
	wire n4628;
	wire n4629;
	wire n4630;
	wire n4631;
	wire n4632;
	wire n4633;
	wire n4634;
	wire n4635;
	wire n4636;
	wire n4637;
	wire n4638;
	wire n4639;
	wire n4640;
	wire n4641;
	wire n4642;
	wire n4643;
	wire n4644;
	wire n4645;
	wire n4646;
	wire n4647;
	wire n4648;
	wire n4649;
	wire n4650;
	wire n4651;
	wire n4652;
	wire n4653;
	wire n4654;
	wire n4655;
	wire n4656;
	wire n4657;
	wire n4658;
	wire n4659;
	wire n4660;
	wire n4661;
	wire n4662;
	wire n4663;
	wire n4664;
	wire n4665;
	wire n4666;
	wire n4667;
	wire n4668;
	wire n4669;
	wire n4670;
	wire n4671;
	wire n4672;
	wire n4673;
	wire n4674;
	wire n4675;
	wire n4676;
	wire n4677;
	wire n4678;
	wire n4679;
	wire n4680;
	wire n4681;
	wire n4682;
	wire n4683;
	wire n4684;
	wire n4685;
	wire n4686;
	wire n4687;
	wire n4688;
	wire n4689;
	wire n4690;
	wire n4691;
	wire n4692;
	wire n4693;
	wire n4694;
	wire n4695;
	wire n4696;
	wire n4697;
	wire n4698;
	wire n4699;
	wire n4700;
	wire n4701;
	wire n4702;
	wire n4703;
	wire n4704;
	wire n4705;
	wire n4706;
	wire n4707;
	wire n4708;
	wire n4709;
	wire n4710;
	wire n4711;
	wire n4712;
	wire n4713;
	wire n4714;
	wire n4715;
	wire n4716;
	wire n4717;
	wire n4718;
	wire n4719;
	wire n4720;
	wire n4721;
	wire n4722;
	wire n4723;
	wire n4724;
	wire n4725;
	wire n4726;
	wire n4727;
	wire n4728;
	wire n4729;
	wire n4730;
	wire n4731;
	wire n4732;
	wire n4733;
	wire n4734;
	wire n4735;
	wire n4736;
	wire n4737;
	wire n4738;
	wire n4739;
	wire n4740;
	wire n4741;
	wire n4742;
	wire n4743;
	wire n4744;
	wire n4745;
	wire n4746;
	wire n4747;
	wire n4748;
	wire n4749;
	wire n4750;
	wire n4751;
	wire n4752;
	wire n4753;
	wire n4754;
	wire n4755;
	wire n4756;
	wire n4757;
	wire n4758;
	wire n4759;
	wire n4760;
	wire n4761;
	wire n4762;
	wire n4763;
	wire n4764;
	wire n4765;
	wire n4766;
	wire n4767;
	wire n4768;
	wire n4769;
	wire n4770;
	wire n4771;
	wire n4772;
	wire n4773;
	wire n4774;
	wire n4775;
	wire n4776;
	wire n4777;
	wire n4778;
	wire n4779;
	wire n4780;
	wire n4781;
	wire n4782;
	wire n4783;
	wire n4784;
	wire n4785;
	wire n4786;
	wire n4787;
	wire n4788;
	wire n4789;
	wire n4790;
	wire n4793;
	wire n4795;
	wire n4796;
	wire n4797;
	wire n4798;
	wire n4799;
	wire n4800;
	wire n4801;
	wire n4802;
	wire n4803;
	wire n4804;
	wire n4805;
	wire n4806;
	wire n4807;
	wire n4808;
	wire n4809;
	wire n4810;
	wire n4811;
	wire n4812;
	wire n4813;
	wire n4814;
	wire n4815;
	wire n4816;
	wire n4817;
	wire n4818;
	wire n4819;
	wire n4820;
	wire n4821;
	wire n4822;
	wire n4823;
	wire n4824;
	wire n4825;
	wire n4826;
	wire n4827;
	wire n4828;
	wire n4829;
	wire n4830;
	wire n4831;
	wire n4832;
	wire n4833;
	wire n4834;
	wire n4835;
	wire n4836;
	wire n4837;
	wire n4838;
	wire n4839;
	wire n4840;
	wire n4841;
	wire n4842;
	wire n4843;
	wire n4844;
	wire n4845;
	wire n4846;
	wire n4847;
	wire n4848;
	wire n4849;
	wire n4850;
	wire n4851;
	wire n4852;
	wire n4853;
	wire n4854;
	wire n4855;
	wire n4856;
	wire n4857;
	wire n4858;
	wire n4859;
	wire n4860;
	wire n4861;
	wire n4862;
	wire n4863;
	wire n4864;
	wire n4865;
	wire n4866;
	wire n4867;
	wire n4868;
	wire n4869;
	wire n4870;
	wire n4871;
	wire n4872;
	wire n4873;
	wire n4874;
	wire n4875;
	wire n4876;
	wire n4877;
	wire n4878;
	wire n4879;
	wire n4880;
	wire n4881;
	wire n4882;
	wire n4883;
	wire n4884;
	wire n4885;
	wire n4886;
	wire n4887;
	wire n4888;
	wire n4889;
	wire n4890;
	wire n4891;
	wire n4892;
	wire n4893;
	wire n4894;
	wire n4895;
	wire n4896;
	wire n4897;
	wire n4898;
	wire n4899;
	wire n4900;
	wire n4901;
	wire n4902;
	wire n4903;
	wire n4904;
	wire n4905;
	wire n4906;
	wire n4907;
	wire n4908;
	wire n4909;
	wire n4910;
	wire n4911;
	wire n4912;
	wire n4913;
	wire n4914;
	wire n4915;
	wire n4916;
	wire n4917;
	wire n4918;
	wire n4919;
	wire n4920;
	wire n4921;
	wire n4922;
	wire n4923;
	wire n4924;
	wire n4925;
	wire n4926;
	wire n4927;
	wire n4928;
	wire n4929;
	wire n4930;
	wire n4931;
	wire n4932;
	wire n4933;
	wire n4934;
	wire n4935;
	wire n4936;
	wire n4937;
	wire n4938;
	wire n4939;
	wire n4940;
	wire n4941;
	wire n4942;
	wire n4943;
	wire n4944;
	wire n4945;
	wire n4946;
	wire n4947;
	wire n4948;
	wire n4949;
	wire n4950;
	wire n4951;
	wire n4952;
	wire n4953;
	wire n4954;
	wire n4955;
	wire n4956;
	wire n4957;
	wire n4958;
	wire n4959;
	wire n4960;
	wire n4961;
	wire n4962;
	wire n4963;
	wire n4964;
	wire n4965;
	wire n4966;
	wire n4967;
	wire n4968;
	wire n4969;
	wire n4970;
	wire n4971;
	wire n4972;
	wire n4973;
	wire n4974;
	wire n4975;
	wire n4976;
	wire n4977;
	wire n4978;
	wire n4979;
	wire n4980;
	wire n4981;
	wire n4982;
	wire n4983;
	wire n4984;
	wire n4985;
	wire n4986;
	wire n4987;
	wire n4988;
	wire n4989;
	wire n4990;
	wire n4991;
	wire n4992;
	wire n4993;
	wire n4994;
	wire n4995;
	wire n4996;
	wire n4997;
	wire n4998;
	wire n4999;
	wire n5000;
	wire n5001;
	wire n5002;
	wire n5003;
	wire n5004;
	wire n5005;
	wire n5006;
	wire n5007;
	wire n5008;
	wire n5009;
	wire n5010;
	wire n5011;
	wire n5012;
	wire n5013;
	wire n5014;
	wire n5015;
	wire n5016;
	wire n5017;
	wire n5018;
	wire n5019;
	wire n5020;
	wire n5021;
	wire n5022;
	wire n5023;
	wire n5024;
	wire n5025;
	wire n5026;
	wire n5027;
	wire n5028;
	wire n5029;
	wire n5030;
	wire n5031;
	wire n5032;
	wire n5033;
	wire n5034;
	wire n5035;
	wire n5036;
	wire n5037;
	wire n5038;
	wire n5039;
	wire n5040;
	wire n5041;
	wire n5042;
	wire n5043;
	wire n5044;
	wire n5045;
	wire n5046;
	wire n5047;
	wire n5048;
	wire n5049;
	wire n5050;
	wire n5051;
	wire n5052;
	wire n5053;
	wire n5054;
	wire n5055;
	wire n5056;
	wire n5057;
	wire n5058;
	wire n5059;
	wire n5060;
	wire n5061;
	wire n5062;
	wire n5063;
	wire n5064;
	wire n5065;
	wire n5066;
	wire n5067;
	wire n5068;
	wire n5069;
	wire n5070;
	wire n5071;
	wire n5072;
	wire n5073;
	wire n5074;
	wire n5075;
	wire n5076;
	wire n5077;
	wire n5078;
	wire n5079;
	wire n5080;
	wire n5081;
	wire n5082;
	wire n5083;
	wire n5084;
	wire n5085;
	wire n5086;
	wire n5087;
	wire n5088;
	wire n5089;
	wire n5090;
	wire n5091;
	wire n5092;
	wire n5093;
	wire n5094;
	wire n5095;
	wire n5096;
	wire n5097;
	wire n5098;
	wire n5099;
	wire n5100;
	wire n5101;
	wire n5102;
	wire n5103;
	wire n5104;
	wire n5105;
	wire n5106;
	wire n5107;
	wire n5108;
	wire n5109;
	wire n5110;
	wire n5111;
	wire n5112;
	wire n5113;
	wire n5114;
	wire n5115;
	wire n5116;
	wire n5119;
	wire n5120;
	wire n5121;
	wire n5123;
	wire n5124;
	wire n5125;
	wire n5126;
	wire n5127;
	wire n5128;
	wire n5129;
	wire n5130;
	wire n5131;
	wire n5132;
	wire n5133;
	wire n5134;
	wire n5135;
	wire n5136;
	wire n5137;
	wire n5138;
	wire n5139;
	wire n5140;
	wire n5141;
	wire n5142;
	wire n5143;
	wire n5144;
	wire n5145;
	wire n5146;
	wire n5147;
	wire n5148;
	wire n5149;
	wire n5150;
	wire n5151;
	wire n5152;
	wire n5153;
	wire n5154;
	wire n5155;
	wire n5156;
	wire n5157;
	wire n5158;
	wire n5159;
	wire n5160;
	wire n5161;
	wire n5162;
	wire n5163;
	wire n5164;
	wire n5165;
	wire n5166;
	wire n5167;
	wire n5168;
	wire n5169;
	wire n5170;
	wire n5171;
	wire n5172;
	wire n5173;
	wire n5174;
	wire n5175;
	wire n5176;
	wire n5177;
	wire n5178;
	wire n5179;
	wire n5180;
	wire n5181;
	wire n5182;
	wire n5183;
	wire n5184;
	wire n5185;
	wire n5186;
	wire n5187;
	wire n5188;
	wire n5189;
	wire n5190;
	wire n5191;
	wire n5192;
	wire n5193;
	wire n5194;
	wire n5195;
	wire n5196;
	wire n5197;
	wire n5198;
	wire n5199;
	wire n5200;
	wire n5201;
	wire n5202;
	wire n5203;
	wire n5204;
	wire n5205;
	wire n5206;
	wire n5207;
	wire n5208;
	wire n5209;
	wire n5210;
	wire n5211;
	wire n5212;
	wire n5213;
	wire n5214;
	wire n5215;
	wire n5216;
	wire n5217;
	wire n5218;
	wire n5219;
	wire n5220;
	wire n5221;
	wire n5222;
	wire n5223;
	wire n5224;
	wire n5225;
	wire n5226;
	wire n5227;
	wire n5228;
	wire n5229;
	wire n5230;
	wire n5231;
	wire n5232;
	wire n5233;
	wire n5234;
	wire n5235;
	wire n5236;
	wire n5237;
	wire n5238;
	wire n5239;
	wire n5240;
	wire n5241;
	wire n5242;
	wire n5243;
	wire n5244;
	wire n5245;
	wire n5246;
	wire n5247;
	wire n5248;
	wire n5249;
	wire n5250;
	wire n5251;
	wire n5252;
	wire n5253;
	wire n5254;
	wire n5255;
	wire n5256;
	wire n5257;
	wire n5258;
	wire n5259;
	wire n5260;
	wire n5261;
	wire n5262;
	wire n5263;
	wire n5264;
	wire n5265;
	wire n5266;
	wire n5267;
	wire n5268;
	wire n5269;
	wire n5270;
	wire n5271;
	wire n5272;
	wire n5273;
	wire n5274;
	wire n5275;
	wire n5276;
	wire n5277;
	wire n5278;
	wire n5279;
	wire n5280;
	wire n5281;
	wire n5282;
	wire n5283;
	wire n5284;
	wire n5285;
	wire n5286;
	wire n5287;
	wire n5288;
	wire n5289;
	wire n5290;
	wire n5291;
	wire n5292;
	wire n5293;
	wire n5294;
	wire n5295;
	wire n5296;
	wire n5297;
	wire n5298;
	wire n5299;
	wire n5300;
	wire n5301;
	wire n5302;
	wire n5303;
	wire n5304;
	wire n5305;
	wire n5306;
	wire n5307;
	wire n5308;
	wire n5309;
	wire n5310;
	wire n5311;
	wire n5312;
	wire n5313;
	wire n5314;
	wire n5315;
	wire n5316;
	wire n5317;
	wire n5318;
	wire n5319;
	wire n5320;
	wire n5321;
	wire n5322;
	wire n5323;
	wire n5324;
	wire n5325;
	wire n5326;
	wire n5327;
	wire n5328;
	wire n5329;
	wire n5330;
	wire n5331;
	wire n5332;
	wire n5333;
	wire n5334;
	wire n5335;
	wire n5336;
	wire n5337;
	wire n5338;
	wire n5339;
	wire n5340;
	wire n5341;
	wire n5342;
	wire n5343;
	wire n5344;
	wire n5345;
	wire n5346;
	wire n5347;
	wire n5348;
	wire n5349;
	wire n5350;
	wire n5351;
	wire n5352;
	wire n5353;
	wire n5354;
	wire n5355;
	wire n5356;
	wire n5357;
	wire n5358;
	wire n5359;
	wire n5360;
	wire n5361;
	wire n5362;
	wire n5363;
	wire n5364;
	wire n5365;
	wire n5366;
	wire n5367;
	wire n5368;
	wire n5369;
	wire n5370;
	wire n5371;
	wire n5372;
	wire n5373;
	wire n5374;
	wire n5375;
	wire n5376;
	wire n5377;
	wire n5378;
	wire n5379;
	wire n5380;
	wire n5381;
	wire n5382;
	wire n5383;
	wire n5384;
	wire n5385;
	wire n5386;
	wire n5387;
	wire n5388;
	wire n5389;
	wire n5390;
	wire n5391;
	wire n5392;
	wire n5393;
	wire n5394;
	wire n5395;
	wire n5396;
	wire n5397;
	wire n5398;
	wire n5399;
	wire n5400;
	wire n5401;
	wire n5402;
	wire n5403;
	wire n5404;
	wire n5405;
	wire n5406;
	wire n5407;
	wire n5408;
	wire n5409;
	wire n5410;
	wire n5411;
	wire n5412;
	wire n5413;
	wire n5414;
	wire n5415;
	wire n5416;
	wire n5417;
	wire n5418;
	wire n5419;
	wire n5420;
	wire n5421;
	wire n5422;
	wire n5423;
	wire n5424;
	wire n5425;
	wire n5426;
	wire n5427;
	wire n5428;
	wire n5429;
	wire n5430;
	wire n5431;
	wire n5432;
	wire n5433;
	wire n5434;
	wire n5435;
	wire n5436;
	wire n5437;
	wire n5440;
	wire n5442;
	wire n5443;
	wire n5444;
	wire n5445;
	wire n5446;
	wire n5447;
	wire n5448;
	wire n5449;
	wire n5450;
	wire n5451;
	wire n5452;
	wire n5453;
	wire n5454;
	wire n5455;
	wire n5456;
	wire n5457;
	wire n5458;
	wire n5459;
	wire n5460;
	wire n5461;
	wire n5462;
	wire n5463;
	wire n5464;
	wire n5465;
	wire n5466;
	wire n5467;
	wire n5468;
	wire n5469;
	wire n5470;
	wire n5471;
	wire n5472;
	wire n5473;
	wire n5474;
	wire n5475;
	wire n5476;
	wire n5477;
	wire n5478;
	wire n5479;
	wire n5480;
	wire n5481;
	wire n5482;
	wire n5483;
	wire n5484;
	wire n5485;
	wire n5486;
	wire n5487;
	wire n5488;
	wire n5489;
	wire n5490;
	wire n5491;
	wire n5492;
	wire n5493;
	wire n5494;
	wire n5495;
	wire n5496;
	wire n5497;
	wire n5498;
	wire n5499;
	wire n5500;
	wire n5501;
	wire n5502;
	wire n5503;
	wire n5504;
	wire n5505;
	wire n5506;
	wire n5507;
	wire n5508;
	wire n5509;
	wire n5510;
	wire n5511;
	wire n5512;
	wire n5513;
	wire n5514;
	wire n5515;
	wire n5516;
	wire n5517;
	wire n5518;
	wire n5519;
	wire n5520;
	wire n5521;
	wire n5522;
	wire n5523;
	wire n5524;
	wire n5525;
	wire n5526;
	wire n5527;
	wire n5528;
	wire n5529;
	wire n5530;
	wire n5531;
	wire n5532;
	wire n5533;
	wire n5534;
	wire n5535;
	wire n5536;
	wire n5537;
	wire n5538;
	wire n5539;
	wire n5540;
	wire n5541;
	wire n5542;
	wire n5543;
	wire n5544;
	wire n5545;
	wire n5546;
	wire n5547;
	wire n5548;
	wire n5549;
	wire n5550;
	wire n5551;
	wire n5552;
	wire n5553;
	wire n5554;
	wire n5555;
	wire n5556;
	wire n5557;
	wire n5558;
	wire n5559;
	wire n5560;
	wire n5561;
	wire n5562;
	wire n5563;
	wire n5564;
	wire n5565;
	wire n5566;
	wire n5567;
	wire n5568;
	wire n5569;
	wire n5570;
	wire n5571;
	wire n5572;
	wire n5573;
	wire n5574;
	wire n5575;
	wire n5576;
	wire n5577;
	wire n5578;
	wire n5579;
	wire n5580;
	wire n5581;
	wire n5582;
	wire n5583;
	wire n5584;
	wire n5585;
	wire n5586;
	wire n5587;
	wire n5588;
	wire n5589;
	wire n5590;
	wire n5591;
	wire n5592;
	wire n5593;
	wire n5594;
	wire n5595;
	wire n5596;
	wire n5597;
	wire n5598;
	wire n5599;
	wire n5600;
	wire n5601;
	wire n5602;
	wire n5603;
	wire n5604;
	wire n5605;
	wire n5606;
	wire n5607;
	wire n5608;
	wire n5609;
	wire n5610;
	wire n5611;
	wire n5612;
	wire n5613;
	wire n5614;
	wire n5615;
	wire n5616;
	wire n5617;
	wire n5618;
	wire n5619;
	wire n5620;
	wire n5621;
	wire n5622;
	wire n5623;
	wire n5624;
	wire n5625;
	wire n5626;
	wire n5627;
	wire n5628;
	wire n5629;
	wire n5630;
	wire n5631;
	wire n5632;
	wire n5633;
	wire n5634;
	wire n5635;
	wire n5636;
	wire n5637;
	wire n5638;
	wire n5639;
	wire n5640;
	wire n5641;
	wire n5642;
	wire n5643;
	wire n5644;
	wire n5645;
	wire n5646;
	wire n5647;
	wire n5648;
	wire n5649;
	wire n5650;
	wire n5651;
	wire n5652;
	wire n5653;
	wire n5654;
	wire n5655;
	wire n5656;
	wire n5657;
	wire n5658;
	wire n5659;
	wire n5660;
	wire n5661;
	wire n5662;
	wire n5663;
	wire n5664;
	wire n5665;
	wire n5666;
	wire n5667;
	wire n5668;
	wire n5669;
	wire n5670;
	wire n5671;
	wire n5672;
	wire n5673;
	wire n5674;
	wire n5675;
	wire n5676;
	wire n5677;
	wire n5678;
	wire n5679;
	wire n5680;
	wire n5681;
	wire n5682;
	wire n5683;
	wire n5684;
	wire n5685;
	wire n5686;
	wire n5687;
	wire n5688;
	wire n5689;
	wire n5690;
	wire n5691;
	wire n5692;
	wire n5693;
	wire n5694;
	wire n5695;
	wire n5696;
	wire n5697;
	wire n5698;
	wire n5699;
	wire n5700;
	wire n5701;
	wire n5702;
	wire n5703;
	wire n5704;
	wire n5705;
	wire n5706;
	wire n5707;
	wire n5708;
	wire n5709;
	wire n5710;
	wire n5711;
	wire n5712;
	wire n5713;
	wire n5714;
	wire n5715;
	wire n5716;
	wire n5717;
	wire n5718;
	wire n5719;
	wire n5720;
	wire n5721;
	wire n5722;
	wire n5723;
	wire n5724;
	wire n5725;
	wire n5726;
	wire n5727;
	wire n5728;
	wire n5729;
	wire n5730;
	wire n5731;
	wire n5732;
	wire n5733;
	wire n5734;
	wire n5735;
	wire n5736;
	wire n5737;
	wire n5738;
	wire n5739;
	wire n5740;
	wire n5741;
	wire n5742;
	wire n5743;
	wire n5744;
	wire n5745;
	wire n5746;
	wire n5747;
	wire n5748;
	wire n5749;
	wire n5750;
	wire n5751;
	wire n5752;
	wire n5753;
	wire n5754;
	wire n5755;
	wire n5756;
	wire n5757;
	wire n5758;
	wire n5759;
	wire n5760;
	wire n5761;
	wire n5762;
	wire n5763;
	wire n5764;
	wire n5765;
	wire n5766;
	wire n5767;
	wire n5768;
	wire n5769;
	wire n5770;
	wire n5771;
	wire n5772;
	wire n5773;
	wire n5774;
	wire n5775;
	wire n5776;
	wire n5777;
	wire n5778;
	wire n5779;
	wire n5780;
	wire n5781;
	wire n5782;
	wire n5783;
	wire n5784;
	wire n5785;
	wire n5786;
	wire n5787;
	wire n5788;
	wire n5791;
	wire n5792;
	wire n5793;
	wire n5794;
	wire n5795;
	wire n5796;
	wire n5797;
	wire n5798;
	wire n5799;
	wire n5800;
	wire n5801;
	wire n5802;
	wire n5803;
	wire n5804;
	wire n5805;
	wire n5806;
	wire n5807;
	wire n5808;
	wire n5809;
	wire n5810;
	wire n5811;
	wire n5812;
	wire n5813;
	wire n5814;
	wire n5815;
	wire n5816;
	wire n5817;
	wire n5818;
	wire n5819;
	wire n5820;
	wire n5821;
	wire n5822;
	wire n5823;
	wire n5824;
	wire n5825;
	wire n5826;
	wire n5827;
	wire n5828;
	wire n5829;
	wire n5830;
	wire n5831;
	wire n5832;
	wire n5833;
	wire n5834;
	wire n5835;
	wire n5836;
	wire n5837;
	wire n5838;
	wire n5839;
	wire n5840;
	wire n5841;
	wire n5842;
	wire n5843;
	wire n5844;
	wire n5845;
	wire n5846;
	wire n5847;
	wire n5849;
	wire n5850;
	wire n5851;
	wire n5852;
	wire n5853;
	wire n5854;
	wire n5855;
	wire n5856;
	wire n5857;
	wire n5858;
	wire n5859;
	wire n5860;
	wire n5861;
	wire n5862;
	wire n5863;
	wire n5864;
	wire n5865;
	wire n5866;
	wire n5867;
	wire n5868;
	wire n5869;
	wire n5870;
	wire n5871;
	wire n5872;
	wire n5873;
	wire n5874;
	wire n5875;
	wire n5876;
	wire n5877;
	wire n5878;
	wire n5879;
	wire n5880;
	wire n5881;
	wire n5882;
	wire n5883;
	wire n5884;
	wire n5885;
	wire n5886;
	wire n5887;
	wire n5888;
	wire n5889;
	wire n5890;
	wire n5891;
	wire n5892;
	wire n5893;
	wire n5894;
	wire n5895;
	wire n5896;
	wire n5897;
	wire n5898;
	wire n5899;
	wire n5900;
	wire n5901;
	wire n5902;
	wire n5903;
	wire n5904;
	wire n5905;
	wire n5906;
	wire n5907;
	wire n5908;
	wire n5909;
	wire n5910;
	wire n5911;
	wire n5912;
	wire n5913;
	wire n5914;
	wire n5915;
	wire n5916;
	wire n5917;
	wire n5918;
	wire n5919;
	wire n5920;
	wire n5921;
	wire n5922;
	wire n5923;
	wire n5924;
	wire n5925;
	wire n5926;
	wire n5927;
	wire n5928;
	wire n5929;
	wire n5930;
	wire n5931;
	wire n5932;
	wire n5933;
	wire n5934;
	wire n5935;
	wire n5936;
	wire n5937;
	wire n5938;
	wire n5939;
	wire n5940;
	wire n5941;
	wire n5942;
	wire n5943;
	wire n5944;
	wire n5945;
	wire n5946;
	wire n5947;
	wire n5948;
	wire n5949;
	wire n5950;
	wire n5951;
	wire n5952;
	wire n5953;
	wire n5954;
	wire n5955;
	wire n5956;
	wire n5957;
	wire n5958;
	wire n5959;
	wire n5960;
	wire n5961;
	wire n5962;
	wire n5963;
	wire n5964;
	wire n5965;
	wire n5966;
	wire n5967;
	wire n5968;
	wire n5969;
	wire n5970;
	wire n5971;
	wire n5972;
	wire n5973;
	wire n5974;
	wire n5975;
	wire n5976;
	wire n5977;
	wire n5978;
	wire n5979;
	wire n5980;
	wire n5981;
	wire n5982;
	wire n5983;
	wire n5984;
	wire n5985;
	wire n5986;
	wire n5987;
	wire n5988;
	wire n5989;
	wire n5990;
	wire n5991;
	wire n5992;
	wire n5993;
	wire n5994;
	wire n5995;
	wire n5996;
	wire n5997;
	wire n5998;
	wire n5999;
	wire n6000;
	wire n6001;
	wire n6002;
	wire n6003;
	wire n6004;
	wire n6005;
	wire n6006;
	wire n6007;
	wire n6008;
	wire n6009;
	wire n6010;
	wire n6011;
	wire n6012;
	wire n6013;
	wire n6014;
	wire n6015;
	wire n6016;
	wire n6017;
	wire n6018;
	wire n6019;
	wire n6020;
	wire n6021;
	wire n6022;
	wire n6023;
	wire n6024;
	wire n6025;
	wire n6026;
	wire n6027;
	wire n6028;
	wire n6029;
	wire n6030;
	wire n6031;
	wire n6032;
	wire n6033;
	wire n6034;
	wire n6035;
	wire n6036;
	wire n6037;
	wire n6038;
	wire n6039;
	wire n6040;
	wire n6041;
	wire n6042;
	wire n6043;
	wire n6044;
	wire n6045;
	wire n6046;
	wire n6047;
	wire n6048;
	wire n6049;
	wire n6050;
	wire n6051;
	wire n6052;
	wire n6053;
	wire n6054;
	wire n6055;
	wire n6056;
	wire n6057;
	wire n6058;
	wire n6059;
	wire n6060;
	wire n6061;
	wire n6062;
	wire n6063;
	wire n6064;
	wire n6065;
	wire n6066;
	wire n6067;
	wire n6068;
	wire n6069;
	wire n6070;
	wire n6071;
	wire n6072;
	wire n6073;
	wire n6074;
	wire n6075;
	wire n6076;
	wire n6077;
	wire n6078;
	wire n6079;
	wire n6080;
	wire n6081;
	wire n6082;
	wire n6083;
	wire n6084;
	wire n6085;
	wire n6086;
	wire n6087;
	wire n6088;
	wire n6089;
	wire n6090;
	wire n6091;
	wire n6092;
	wire n6093;
	wire n6094;
	wire n6095;
	wire n6096;
	wire n6097;
	wire n6098;
	wire n6099;
	wire n6100;
	wire n6101;
	wire n6102;
	wire n6103;
	wire n6104;
	wire n6105;
	wire n6106;
	wire n6107;
	wire n6108;
	wire n6109;
	wire n6110;
	wire n6111;
	wire n6112;
	wire n6113;
	wire n6114;
	wire n6115;
	wire n6116;
	wire n6117;
	wire n6118;
	wire n6119;
	wire n6120;
	wire n6121;
	wire n6122;
	wire n6123;
	wire n6124;
	wire n6125;
	wire n6128;
	wire n6130;
	wire n6131;
	wire n6132;
	wire n6133;
	wire n6134;
	wire n6135;
	wire n6136;
	wire n6137;
	wire n6138;
	wire n6139;
	wire n6140;
	wire n6141;
	wire n6142;
	wire n6143;
	wire n6144;
	wire n6145;
	wire n6146;
	wire n6147;
	wire n6148;
	wire n6149;
	wire n6150;
	wire n6151;
	wire n6152;
	wire n6153;
	wire n6154;
	wire n6155;
	wire n6156;
	wire n6157;
	wire n6158;
	wire n6159;
	wire n6160;
	wire n6161;
	wire n6162;
	wire n6163;
	wire n6164;
	wire n6165;
	wire n6166;
	wire n6167;
	wire n6168;
	wire n6169;
	wire n6170;
	wire n6171;
	wire n6172;
	wire n6173;
	wire n6174;
	wire n6175;
	wire n6176;
	wire n6177;
	wire n6178;
	wire n6179;
	wire n6180;
	wire n6181;
	wire n6182;
	wire n6183;
	wire n6184;
	wire n6185;
	wire n6186;
	wire n6187;
	wire n6188;
	wire n6189;
	wire n6190;
	wire n6191;
	wire n6192;
	wire n6193;
	wire n6194;
	wire n6195;
	wire n6196;
	wire n6197;
	wire n6198;
	wire n6199;
	wire n6200;
	wire n6201;
	wire n6202;
	wire n6203;
	wire n6204;
	wire n6205;
	wire n6206;
	wire n6207;
	wire n6208;
	wire n6209;
	wire n6210;
	wire n6211;
	wire n6212;
	wire n6213;
	wire n6214;
	wire n6215;
	wire n6216;
	wire n6217;
	wire n6218;
	wire n6219;
	wire n6220;
	wire n6221;
	wire n6222;
	wire n6223;
	wire n6224;
	wire n6225;
	wire n6226;
	wire n6227;
	wire n6228;
	wire n6229;
	wire n6230;
	wire n6231;
	wire n6232;
	wire n6233;
	wire n6234;
	wire n6235;
	wire n6236;
	wire n6237;
	wire n6238;
	wire n6239;
	wire n6240;
	wire n6241;
	wire n6242;
	wire n6243;
	wire n6244;
	wire n6245;
	wire n6246;
	wire n6247;
	wire n6248;
	wire n6249;
	wire n6250;
	wire n6251;
	wire n6252;
	wire n6253;
	wire n6254;
	wire n6255;
	wire n6256;
	wire n6257;
	wire n6258;
	wire n6259;
	wire n6260;
	wire n6261;
	wire n6262;
	wire n6263;
	wire n6264;
	wire n6265;
	wire n6266;
	wire n6267;
	wire n6268;
	wire n6269;
	wire n6270;
	wire n6271;
	wire n6272;
	wire n6273;
	wire n6274;
	wire n6275;
	wire n6276;
	wire n6277;
	wire n6278;
	wire n6279;
	wire n6280;
	wire n6281;
	wire n6282;
	wire n6283;
	wire n6284;
	wire n6285;
	wire n6286;
	wire n6287;
	wire n6288;
	wire n6289;
	wire n6290;
	wire n6291;
	wire n6292;
	wire n6293;
	wire n6294;
	wire n6295;
	wire n6296;
	wire n6297;
	wire n6298;
	wire n6299;
	wire n6300;
	wire n6301;
	wire n6302;
	wire n6303;
	wire n6304;
	wire n6305;
	wire n6306;
	wire n6307;
	wire n6308;
	wire n6309;
	wire n6310;
	wire n6311;
	wire n6312;
	wire n6313;
	wire n6314;
	wire n6315;
	wire n6316;
	wire n6317;
	wire n6318;
	wire n6319;
	wire n6320;
	wire n6321;
	wire n6322;
	wire n6323;
	wire n6324;
	wire n6325;
	wire n6326;
	wire n6327;
	wire n6328;
	wire n6329;
	wire n6330;
	wire n6331;
	wire n6332;
	wire n6333;
	wire n6334;
	wire n6335;
	wire n6336;
	wire n6337;
	wire n6338;
	wire n6339;
	wire n6340;
	wire n6341;
	wire n6342;
	wire n6343;
	wire n6344;
	wire n6345;
	wire n6346;
	wire n6347;
	wire n6348;
	wire n6349;
	wire n6350;
	wire n6351;
	wire n6352;
	wire n6353;
	wire n6354;
	wire n6355;
	wire n6356;
	wire n6357;
	wire n6358;
	wire n6359;
	wire n6360;
	wire n6361;
	wire n6362;
	wire n6363;
	wire n6364;
	wire n6365;
	wire n6366;
	wire n6367;
	wire n6368;
	wire n6369;
	wire n6370;
	wire n6371;
	wire n6372;
	wire n6373;
	wire n6374;
	wire n6375;
	wire n6376;
	wire n6377;
	wire n6378;
	wire n6379;
	wire n6380;
	wire n6381;
	wire n6382;
	wire n6383;
	wire n6384;
	wire n6385;
	wire n6386;
	wire n6387;
	wire n6388;
	wire n6389;
	wire n6390;
	wire n6391;
	wire n6392;
	wire n6393;
	wire n6394;
	wire n6395;
	wire n6396;
	wire n6397;
	wire n6398;
	wire n6399;
	wire n6400;
	wire n6401;
	wire n6402;
	wire n6403;
	wire n6404;
	wire n6405;
	wire n6406;
	wire n6407;
	wire n6408;
	wire n6409;
	wire n6410;
	wire n6411;
	wire n6412;
	wire n6413;
	wire n6414;
	wire n6415;
	wire n6416;
	wire n6417;
	wire n6418;
	wire n6419;
	wire n6420;
	wire n6421;
	wire n6422;
	wire n6423;
	wire n6424;
	wire n6425;
	wire n6426;
	wire n6427;
	wire n6428;
	wire n6429;
	wire n6430;
	wire n6431;
	wire n6432;
	wire n6433;
	wire n6434;
	wire n6435;
	wire n6436;
	wire n6437;
	wire n6438;
	wire n6439;
	wire n6440;
	wire n6441;
	wire n6442;
	wire n6443;
	wire n6444;
	wire n6445;
	wire n6446;
	wire n6447;
	wire n6448;
	wire n6449;
	wire n6450;
	wire n6451;
	wire n6452;
	wire n6453;
	wire n6454;
	wire n6455;
	wire n6456;
	wire n6457;
	wire n6458;
	wire n6459;
	wire n6460;
	wire n6461;
	wire n6462;
	wire n6463;
	wire n6464;
	wire n6465;
	wire n6466;
	wire n6467;
	wire n6468;
	wire n6469;
	wire n6470;
	wire n6471;
	wire n6472;
	wire n6473;
	wire n6474;
	wire n6475;
	wire n6476;
	wire n6477;
	wire n6478;
	wire n6479;
	wire n6480;
	wire n6481;
	wire n6482;
	wire n6483;
	wire n6484;
	wire n6485;
	wire n6486;
	wire n6487;
	wire n6488;
	wire n6489;
	wire n6490;
	wire n6491;
	wire n6492;
	wire n6493;
	wire n6494;
	wire n6495;
	wire n6496;
	wire n6497;
	wire n6498;
	wire n6499;
	wire n6500;
	wire n6503;
	wire n6504;
	wire n6505;
	wire n6506;
	wire n6507;
	wire n6508;
	wire n6509;
	wire n6510;
	wire n6511;
	wire n6512;
	wire n6513;
	wire n6514;
	wire n6515;
	wire n6516;
	wire n6517;
	wire n6518;
	wire n6519;
	wire n6520;
	wire n6521;
	wire n6522;
	wire n6523;
	wire n6524;
	wire n6525;
	wire n6526;
	wire n6527;
	wire n6528;
	wire n6529;
	wire n6530;
	wire n6531;
	wire n6532;
	wire n6533;
	wire n6534;
	wire n6535;
	wire n6536;
	wire n6537;
	wire n6538;
	wire n6539;
	wire n6540;
	wire n6541;
	wire n6542;
	wire n6543;
	wire n6544;
	wire n6545;
	wire n6547;
	wire n6548;
	wire n6549;
	wire n6550;
	wire n6551;
	wire n6552;
	wire n6553;
	wire n6554;
	wire n6555;
	wire n6556;
	wire n6557;
	wire n6558;
	wire n6559;
	wire n6560;
	wire n6561;
	wire n6562;
	wire n6563;
	wire n6564;
	wire n6565;
	wire n6566;
	wire n6567;
	wire n6568;
	wire n6569;
	wire n6570;
	wire n6571;
	wire n6572;
	wire n6573;
	wire n6574;
	wire n6575;
	wire n6576;
	wire n6577;
	wire n6578;
	wire n6579;
	wire n6580;
	wire n6581;
	wire n6582;
	wire n6583;
	wire n6584;
	wire n6585;
	wire n6586;
	wire n6587;
	wire n6588;
	wire n6589;
	wire n6590;
	wire n6591;
	wire n6592;
	wire n6593;
	wire n6594;
	wire n6595;
	wire n6596;
	wire n6597;
	wire n6598;
	wire n6599;
	wire n6600;
	wire n6601;
	wire n6602;
	wire n6603;
	wire n6604;
	wire n6605;
	wire n6606;
	wire n6607;
	wire n6608;
	wire n6609;
	wire n6610;
	wire n6611;
	wire n6612;
	wire n6613;
	wire n6614;
	wire n6615;
	wire n6616;
	wire n6617;
	wire n6618;
	wire n6619;
	wire n6620;
	wire n6621;
	wire n6622;
	wire n6623;
	wire n6624;
	wire n6625;
	wire n6626;
	wire n6627;
	wire n6628;
	wire n6629;
	wire n6630;
	wire n6631;
	wire n6632;
	wire n6633;
	wire n6634;
	wire n6635;
	wire n6636;
	wire n6637;
	wire n6638;
	wire n6639;
	wire n6640;
	wire n6641;
	wire n6642;
	wire n6643;
	wire n6644;
	wire n6645;
	wire n6646;
	wire n6647;
	wire n6648;
	wire n6649;
	wire n6650;
	wire n6651;
	wire n6652;
	wire n6653;
	wire n6654;
	wire n6655;
	wire n6656;
	wire n6657;
	wire n6658;
	wire n6659;
	wire n6660;
	wire n6661;
	wire n6662;
	wire n6663;
	wire n6664;
	wire n6665;
	wire n6666;
	wire n6667;
	wire n6668;
	wire n6669;
	wire n6670;
	wire n6671;
	wire n6672;
	wire n6673;
	wire n6674;
	wire n6675;
	wire n6676;
	wire n6677;
	wire n6678;
	wire n6679;
	wire n6680;
	wire n6681;
	wire n6682;
	wire n6683;
	wire n6684;
	wire n6685;
	wire n6686;
	wire n6687;
	wire n6688;
	wire n6689;
	wire n6690;
	wire n6691;
	wire n6692;
	wire n6693;
	wire n6694;
	wire n6695;
	wire n6696;
	wire n6697;
	wire n6698;
	wire n6699;
	wire n6700;
	wire n6701;
	wire n6702;
	wire n6703;
	wire n6704;
	wire n6705;
	wire n6706;
	wire n6707;
	wire n6708;
	wire n6709;
	wire n6710;
	wire n6711;
	wire n6712;
	wire n6713;
	wire n6714;
	wire n6715;
	wire n6716;
	wire n6717;
	wire n6718;
	wire n6719;
	wire n6720;
	wire n6721;
	wire n6722;
	wire n6723;
	wire n6724;
	wire n6725;
	wire n6726;
	wire n6727;
	wire n6728;
	wire n6729;
	wire n6730;
	wire n6731;
	wire n6732;
	wire n6733;
	wire n6734;
	wire n6735;
	wire n6736;
	wire n6737;
	wire n6738;
	wire n6739;
	wire n6740;
	wire n6741;
	wire n6742;
	wire n6743;
	wire n6744;
	wire n6745;
	wire n6746;
	wire n6747;
	wire n6748;
	wire n6749;
	wire n6750;
	wire n6751;
	wire n6752;
	wire n6753;
	wire n6754;
	wire n6755;
	wire n6756;
	wire n6757;
	wire n6758;
	wire n6759;
	wire n6760;
	wire n6761;
	wire n6762;
	wire n6763;
	wire n6764;
	wire n6765;
	wire n6766;
	wire n6767;
	wire n6768;
	wire n6769;
	wire n6770;
	wire n6771;
	wire n6772;
	wire n6773;
	wire n6774;
	wire n6775;
	wire n6776;
	wire n6777;
	wire n6778;
	wire n6779;
	wire n6780;
	wire n6781;
	wire n6782;
	wire n6783;
	wire n6784;
	wire n6785;
	wire n6786;
	wire n6787;
	wire n6788;
	wire n6789;
	wire n6790;
	wire n6791;
	wire n6792;
	wire n6793;
	wire n6794;
	wire n6795;
	wire n6796;
	wire n6797;
	wire n6798;
	wire n6799;
	wire n6800;
	wire n6801;
	wire n6802;
	wire n6803;
	wire n6804;
	wire n6805;
	wire n6806;
	wire n6807;
	wire n6808;
	wire n6809;
	wire n6810;
	wire n6811;
	wire n6812;
	wire n6813;
	wire n6814;
	wire n6815;
	wire n6816;
	wire n6817;
	wire n6818;
	wire n6819;
	wire n6820;
	wire n6821;
	wire n6822;
	wire n6823;
	wire n6824;
	wire n6825;
	wire n6826;
	wire n6827;
	wire n6828;
	wire n6829;
	wire n6830;
	wire n6831;
	wire n6832;
	wire n6833;
	wire n6834;
	wire n6835;
	wire n6836;
	wire n6837;
	wire n6838;
	wire n6839;
	wire n6840;
	wire n6841;
	wire n6842;
	wire n6843;
	wire n6844;
	wire n6845;
	wire n6846;
	wire n6847;
	wire n6848;
	wire n6849;
	wire n6850;
	wire n6851;
	wire n6852;
	wire n6853;
	wire n6854;
	wire n6855;
	wire n6856;
	wire n6857;
	wire n6858;
	wire n6859;
	wire n6860;
	wire n6861;
	wire n6862;
	wire n6865;
	wire n6867;
	wire n6868;
	wire n6869;
	wire n6870;
	wire n6871;
	wire n6872;
	wire n6873;
	wire n6874;
	wire n6875;
	wire n6876;
	wire n6877;
	wire n6878;
	wire n6879;
	wire n6880;
	wire n6881;
	wire n6882;
	wire n6883;
	wire n6884;
	wire n6885;
	wire n6886;
	wire n6887;
	wire n6888;
	wire n6889;
	wire n6890;
	wire n6891;
	wire n6892;
	wire n6893;
	wire n6894;
	wire n6895;
	wire n6896;
	wire n6897;
	wire n6898;
	wire n6899;
	wire n6900;
	wire n6901;
	wire n6902;
	wire n6903;
	wire n6904;
	wire n6905;
	wire n6906;
	wire n6907;
	wire n6908;
	wire n6909;
	wire n6910;
	wire n6911;
	wire n6912;
	wire n6913;
	wire n6914;
	wire n6915;
	wire n6916;
	wire n6917;
	wire n6918;
	wire n6919;
	wire n6920;
	wire n6921;
	wire n6922;
	wire n6923;
	wire n6924;
	wire n6925;
	wire n6926;
	wire n6927;
	wire n6928;
	wire n6929;
	wire n6930;
	wire n6931;
	wire n6932;
	wire n6933;
	wire n6934;
	wire n6935;
	wire n6936;
	wire n6937;
	wire n6938;
	wire n6939;
	wire n6940;
	wire n6941;
	wire n6942;
	wire n6943;
	wire n6944;
	wire n6945;
	wire n6946;
	wire n6947;
	wire n6948;
	wire n6949;
	wire n6950;
	wire n6951;
	wire n6952;
	wire n6953;
	wire n6954;
	wire n6955;
	wire n6956;
	wire n6957;
	wire n6958;
	wire n6959;
	wire n6960;
	wire n6961;
	wire n6962;
	wire n6963;
	wire n6964;
	wire n6965;
	wire n6966;
	wire n6967;
	wire n6968;
	wire n6969;
	wire n6970;
	wire n6971;
	wire n6972;
	wire n6973;
	wire n6974;
	wire n6975;
	wire n6976;
	wire n6977;
	wire n6978;
	wire n6979;
	wire n6980;
	wire n6981;
	wire n6982;
	wire n6983;
	wire n6984;
	wire n6985;
	wire n6986;
	wire n6987;
	wire n6988;
	wire n6989;
	wire n6990;
	wire n6991;
	wire n6992;
	wire n6993;
	wire n6994;
	wire n6995;
	wire n6996;
	wire n6997;
	wire n6998;
	wire n6999;
	wire n7000;
	wire n7001;
	wire n7002;
	wire n7003;
	wire n7004;
	wire n7005;
	wire n7006;
	wire n7007;
	wire n7008;
	wire n7009;
	wire n7010;
	wire n7011;
	wire n7012;
	wire n7013;
	wire n7014;
	wire n7015;
	wire n7016;
	wire n7017;
	wire n7018;
	wire n7019;
	wire n7020;
	wire n7021;
	wire n7022;
	wire n7023;
	wire n7024;
	wire n7025;
	wire n7026;
	wire n7027;
	wire n7028;
	wire n7029;
	wire n7030;
	wire n7031;
	wire n7032;
	wire n7033;
	wire n7034;
	wire n7035;
	wire n7036;
	wire n7037;
	wire n7038;
	wire n7039;
	wire n7040;
	wire n7041;
	wire n7042;
	wire n7043;
	wire n7044;
	wire n7045;
	wire n7046;
	wire n7047;
	wire n7048;
	wire n7049;
	wire n7050;
	wire n7051;
	wire n7052;
	wire n7053;
	wire n7054;
	wire n7055;
	wire n7056;
	wire n7057;
	wire n7058;
	wire n7059;
	wire n7060;
	wire n7061;
	wire n7062;
	wire n7063;
	wire n7064;
	wire n7065;
	wire n7066;
	wire n7067;
	wire n7068;
	wire n7069;
	wire n7070;
	wire n7071;
	wire n7072;
	wire n7073;
	wire n7074;
	wire n7075;
	wire n7076;
	wire n7077;
	wire n7078;
	wire n7079;
	wire n7080;
	wire n7081;
	wire n7082;
	wire n7083;
	wire n7084;
	wire n7085;
	wire n7086;
	wire n7087;
	wire n7088;
	wire n7089;
	wire n7090;
	wire n7091;
	wire n7092;
	wire n7093;
	wire n7094;
	wire n7095;
	wire n7096;
	wire n7097;
	wire n7098;
	wire n7099;
	wire n7100;
	wire n7101;
	wire n7102;
	wire n7103;
	wire n7104;
	wire n7105;
	wire n7106;
	wire n7107;
	wire n7108;
	wire n7109;
	wire n7110;
	wire n7111;
	wire n7112;
	wire n7113;
	wire n7114;
	wire n7115;
	wire n7116;
	wire n7117;
	wire n7118;
	wire n7119;
	wire n7120;
	wire n7121;
	wire n7122;
	wire n7123;
	wire n7124;
	wire n7125;
	wire n7126;
	wire n7127;
	wire n7128;
	wire n7129;
	wire n7130;
	wire n7131;
	wire n7132;
	wire n7133;
	wire n7134;
	wire n7135;
	wire n7136;
	wire n7137;
	wire n7138;
	wire n7139;
	wire n7140;
	wire n7141;
	wire n7142;
	wire n7143;
	wire n7144;
	wire n7145;
	wire n7146;
	wire n7147;
	wire n7148;
	wire n7149;
	wire n7150;
	wire n7151;
	wire n7152;
	wire n7153;
	wire n7154;
	wire n7155;
	wire n7156;
	wire n7157;
	wire n7158;
	wire n7159;
	wire n7160;
	wire n7161;
	wire n7162;
	wire n7163;
	wire n7164;
	wire n7165;
	wire n7166;
	wire n7167;
	wire n7168;
	wire n7169;
	wire n7170;
	wire n7171;
	wire n7172;
	wire n7173;
	wire n7174;
	wire n7175;
	wire n7176;
	wire n7177;
	wire n7178;
	wire n7179;
	wire n7180;
	wire n7181;
	wire n7182;
	wire n7183;
	wire n7184;
	wire n7185;
	wire n7186;
	wire n7187;
	wire n7188;
	wire n7189;
	wire n7190;
	wire n7191;
	wire n7192;
	wire n7193;
	wire n7194;
	wire n7195;
	wire n7196;
	wire n7197;
	wire n7198;
	wire n7199;
	wire n7200;
	wire n7201;
	wire n7202;
	wire n7203;
	wire n7204;
	wire n7205;
	wire n7206;
	wire n7207;
	wire n7208;
	wire n7209;
	wire n7210;
	wire n7211;
	wire n7212;
	wire n7213;
	wire n7214;
	wire n7215;
	wire n7216;
	wire n7217;
	wire n7218;
	wire n7219;
	wire n7220;
	wire n7221;
	wire n7222;
	wire n7223;
	wire n7224;
	wire n7225;
	wire n7226;
	wire n7227;
	wire n7228;
	wire n7229;
	wire n7230;
	wire n7231;
	wire n7232;
	wire n7233;
	wire n7234;
	wire n7235;
	wire n7236;
	wire n7237;
	wire n7238;
	wire n7239;
	wire n7240;
	wire n7241;
	wire n7242;
	wire n7243;
	wire n7244;
	wire n7245;
	wire n7246;
	wire n7247;
	wire n7248;
	wire n7249;
	wire n7250;
	wire n7251;
	wire n7252;
	wire n7253;
	wire n7254;
	wire n7255;
	wire n7256;
	wire n7257;
	wire n7258;
	wire n7259;
	wire n7260;
	wire n7263;
	wire n7264;
	wire n7265;
	wire n7266;
	wire n7267;
	wire n7268;
	wire n7269;
	wire n7270;
	wire n7271;
	wire n7272;
	wire n7273;
	wire n7274;
	wire n7275;
	wire n7276;
	wire n7277;
	wire n7278;
	wire n7279;
	wire n7280;
	wire n7281;
	wire n7282;
	wire n7283;
	wire n7284;
	wire n7285;
	wire n7286;
	wire n7287;
	wire n7288;
	wire n7289;
	wire n7290;
	wire n7291;
	wire n7292;
	wire n7293;
	wire n7294;
	wire n7295;
	wire n7296;
	wire n7297;
	wire n7298;
	wire n7299;
	wire n7300;
	wire n7301;
	wire n7302;
	wire n7303;
	wire n7304;
	wire n7305;
	wire n7306;
	wire n7307;
	wire n7308;
	wire n7309;
	wire n7310;
	wire n7311;
	wire n7312;
	wire n7313;
	wire n7314;
	wire n7315;
	wire n7316;
	wire n7317;
	wire n7318;
	wire n7319;
	wire n7320;
	wire n7321;
	wire n7322;
	wire n7323;
	wire n7325;
	wire n7326;
	wire n7327;
	wire n7328;
	wire n7329;
	wire n7330;
	wire n7331;
	wire n7332;
	wire n7333;
	wire n7334;
	wire n7335;
	wire n7336;
	wire n7337;
	wire n7338;
	wire n7339;
	wire n7340;
	wire n7341;
	wire n7342;
	wire n7343;
	wire n7344;
	wire n7345;
	wire n7346;
	wire n7347;
	wire n7348;
	wire n7349;
	wire n7350;
	wire n7351;
	wire n7352;
	wire n7353;
	wire n7354;
	wire n7355;
	wire n7356;
	wire n7357;
	wire n7358;
	wire n7359;
	wire n7360;
	wire n7361;
	wire n7362;
	wire n7363;
	wire n7364;
	wire n7365;
	wire n7366;
	wire n7367;
	wire n7368;
	wire n7369;
	wire n7370;
	wire n7371;
	wire n7372;
	wire n7373;
	wire n7374;
	wire n7375;
	wire n7376;
	wire n7377;
	wire n7378;
	wire n7379;
	wire n7380;
	wire n7381;
	wire n7382;
	wire n7383;
	wire n7384;
	wire n7385;
	wire n7386;
	wire n7387;
	wire n7388;
	wire n7389;
	wire n7390;
	wire n7391;
	wire n7392;
	wire n7393;
	wire n7394;
	wire n7395;
	wire n7396;
	wire n7397;
	wire n7398;
	wire n7399;
	wire n7400;
	wire n7401;
	wire n7402;
	wire n7403;
	wire n7404;
	wire n7405;
	wire n7406;
	wire n7407;
	wire n7408;
	wire n7409;
	wire n7410;
	wire n7411;
	wire n7412;
	wire n7413;
	wire n7414;
	wire n7415;
	wire n7416;
	wire n7417;
	wire n7418;
	wire n7419;
	wire n7420;
	wire n7421;
	wire n7422;
	wire n7423;
	wire n7424;
	wire n7425;
	wire n7426;
	wire n7427;
	wire n7428;
	wire n7429;
	wire n7430;
	wire n7431;
	wire n7432;
	wire n7433;
	wire n7434;
	wire n7435;
	wire n7436;
	wire n7437;
	wire n7438;
	wire n7439;
	wire n7440;
	wire n7441;
	wire n7442;
	wire n7443;
	wire n7444;
	wire n7445;
	wire n7446;
	wire n7447;
	wire n7448;
	wire n7449;
	wire n7450;
	wire n7451;
	wire n7452;
	wire n7453;
	wire n7454;
	wire n7455;
	wire n7456;
	wire n7457;
	wire n7458;
	wire n7459;
	wire n7460;
	wire n7461;
	wire n7462;
	wire n7463;
	wire n7464;
	wire n7465;
	wire n7466;
	wire n7467;
	wire n7468;
	wire n7469;
	wire n7470;
	wire n7471;
	wire n7472;
	wire n7473;
	wire n7474;
	wire n7475;
	wire n7476;
	wire n7477;
	wire n7478;
	wire n7479;
	wire n7480;
	wire n7481;
	wire n7482;
	wire n7483;
	wire n7484;
	wire n7485;
	wire n7486;
	wire n7487;
	wire n7488;
	wire n7489;
	wire n7490;
	wire n7491;
	wire n7492;
	wire n7493;
	wire n7494;
	wire n7495;
	wire n7496;
	wire n7497;
	wire n7498;
	wire n7499;
	wire n7500;
	wire n7501;
	wire n7502;
	wire n7503;
	wire n7504;
	wire n7505;
	wire n7506;
	wire n7507;
	wire n7508;
	wire n7509;
	wire n7510;
	wire n7511;
	wire n7512;
	wire n7513;
	wire n7514;
	wire n7515;
	wire n7516;
	wire n7517;
	wire n7518;
	wire n7519;
	wire n7520;
	wire n7521;
	wire n7522;
	wire n7523;
	wire n7524;
	wire n7525;
	wire n7526;
	wire n7527;
	wire n7528;
	wire n7529;
	wire n7530;
	wire n7531;
	wire n7532;
	wire n7533;
	wire n7534;
	wire n7535;
	wire n7536;
	wire n7537;
	wire n7538;
	wire n7539;
	wire n7540;
	wire n7541;
	wire n7542;
	wire n7543;
	wire n7544;
	wire n7545;
	wire n7546;
	wire n7547;
	wire n7548;
	wire n7549;
	wire n7550;
	wire n7551;
	wire n7552;
	wire n7553;
	wire n7554;
	wire n7555;
	wire n7556;
	wire n7557;
	wire n7558;
	wire n7559;
	wire n7560;
	wire n7561;
	wire n7562;
	wire n7563;
	wire n7564;
	wire n7565;
	wire n7566;
	wire n7567;
	wire n7568;
	wire n7569;
	wire n7570;
	wire n7571;
	wire n7572;
	wire n7573;
	wire n7574;
	wire n7575;
	wire n7576;
	wire n7577;
	wire n7578;
	wire n7579;
	wire n7580;
	wire n7581;
	wire n7582;
	wire n7583;
	wire n7584;
	wire n7585;
	wire n7586;
	wire n7587;
	wire n7588;
	wire n7589;
	wire n7590;
	wire n7591;
	wire n7592;
	wire n7593;
	wire n7594;
	wire n7595;
	wire n7596;
	wire n7597;
	wire n7598;
	wire n7599;
	wire n7600;
	wire n7601;
	wire n7602;
	wire n7603;
	wire n7604;
	wire n7605;
	wire n7606;
	wire n7607;
	wire n7608;
	wire n7609;
	wire n7610;
	wire n7611;
	wire n7612;
	wire n7613;
	wire n7614;
	wire n7615;
	wire n7616;
	wire n7617;
	wire n7618;
	wire n7619;
	wire n7620;
	wire n7621;
	wire n7622;
	wire n7623;
	wire n7624;
	wire n7625;
	wire n7626;
	wire n7627;
	wire n7628;
	wire n7629;
	wire n7630;
	wire n7631;
	wire n7632;
	wire n7633;
	wire n7634;
	wire n7635;
	wire n7636;
	wire n7637;
	wire n7640;
	wire n7642;
	wire n7643;
	wire n7644;
	wire n7645;
	wire n7646;
	wire n7647;
	wire n7648;
	wire n7649;
	wire n7650;
	wire n7651;
	wire n7652;
	wire n7653;
	wire n7654;
	wire n7655;
	wire n7656;
	wire n7657;
	wire n7658;
	wire n7659;
	wire n7660;
	wire n7661;
	wire n7662;
	wire n7663;
	wire n7664;
	wire n7665;
	wire n7666;
	wire n7667;
	wire n7668;
	wire n7669;
	wire n7670;
	wire n7671;
	wire n7672;
	wire n7673;
	wire n7674;
	wire n7675;
	wire n7676;
	wire n7677;
	wire n7678;
	wire n7679;
	wire n7680;
	wire n7681;
	wire n7682;
	wire n7683;
	wire n7684;
	wire n7685;
	wire n7686;
	wire n7687;
	wire n7688;
	wire n7689;
	wire n7690;
	wire n7691;
	wire n7692;
	wire n7693;
	wire n7694;
	wire n7695;
	wire n7696;
	wire n7697;
	wire n7698;
	wire n7699;
	wire n7700;
	wire n7701;
	wire n7702;
	wire n7703;
	wire n7704;
	wire n7705;
	wire n7706;
	wire n7707;
	wire n7708;
	wire n7709;
	wire n7710;
	wire n7711;
	wire n7712;
	wire n7713;
	wire n7714;
	wire n7715;
	wire n7716;
	wire n7717;
	wire n7718;
	wire n7719;
	wire n7720;
	wire n7721;
	wire n7722;
	wire n7723;
	wire n7724;
	wire n7725;
	wire n7726;
	wire n7727;
	wire n7728;
	wire n7729;
	wire n7730;
	wire n7731;
	wire n7732;
	wire n7733;
	wire n7734;
	wire n7735;
	wire n7736;
	wire n7737;
	wire n7738;
	wire n7739;
	wire n7740;
	wire n7741;
	wire n7742;
	wire n7743;
	wire n7744;
	wire n7745;
	wire n7746;
	wire n7747;
	wire n7748;
	wire n7749;
	wire n7750;
	wire n7751;
	wire n7752;
	wire n7753;
	wire n7754;
	wire n7755;
	wire n7756;
	wire n7757;
	wire n7758;
	wire n7759;
	wire n7760;
	wire n7761;
	wire n7762;
	wire n7763;
	wire n7764;
	wire n7765;
	wire n7766;
	wire n7767;
	wire n7768;
	wire n7769;
	wire n7770;
	wire n7771;
	wire n7772;
	wire n7773;
	wire n7774;
	wire n7775;
	wire n7776;
	wire n7777;
	wire n7778;
	wire n7779;
	wire n7780;
	wire n7781;
	wire n7782;
	wire n7783;
	wire n7784;
	wire n7785;
	wire n7786;
	wire n7787;
	wire n7788;
	wire n7789;
	wire n7790;
	wire n7791;
	wire n7792;
	wire n7793;
	wire n7794;
	wire n7795;
	wire n7796;
	wire n7797;
	wire n7798;
	wire n7799;
	wire n7800;
	wire n7801;
	wire n7802;
	wire n7803;
	wire n7804;
	wire n7805;
	wire n7806;
	wire n7807;
	wire n7808;
	wire n7809;
	wire n7810;
	wire n7811;
	wire n7812;
	wire n7813;
	wire n7814;
	wire n7815;
	wire n7816;
	wire n7817;
	wire n7818;
	wire n7819;
	wire n7820;
	wire n7821;
	wire n7822;
	wire n7823;
	wire n7824;
	wire n7825;
	wire n7826;
	wire n7827;
	wire n7828;
	wire n7829;
	wire n7830;
	wire n7831;
	wire n7832;
	wire n7833;
	wire n7834;
	wire n7835;
	wire n7836;
	wire n7837;
	wire n7838;
	wire n7839;
	wire n7840;
	wire n7841;
	wire n7842;
	wire n7843;
	wire n7844;
	wire n7845;
	wire n7846;
	wire n7847;
	wire n7848;
	wire n7849;
	wire n7850;
	wire n7851;
	wire n7852;
	wire n7853;
	wire n7854;
	wire n7855;
	wire n7856;
	wire n7857;
	wire n7858;
	wire n7859;
	wire n7860;
	wire n7861;
	wire n7862;
	wire n7863;
	wire n7864;
	wire n7865;
	wire n7866;
	wire n7867;
	wire n7868;
	wire n7869;
	wire n7870;
	wire n7871;
	wire n7872;
	wire n7873;
	wire n7874;
	wire n7875;
	wire n7876;
	wire n7877;
	wire n7878;
	wire n7879;
	wire n7880;
	wire n7881;
	wire n7882;
	wire n7883;
	wire n7884;
	wire n7885;
	wire n7886;
	wire n7887;
	wire n7888;
	wire n7889;
	wire n7890;
	wire n7891;
	wire n7892;
	wire n7893;
	wire n7894;
	wire n7895;
	wire n7896;
	wire n7897;
	wire n7898;
	wire n7899;
	wire n7900;
	wire n7901;
	wire n7902;
	wire n7903;
	wire n7904;
	wire n7905;
	wire n7906;
	wire n7907;
	wire n7908;
	wire n7909;
	wire n7910;
	wire n7911;
	wire n7912;
	wire n7913;
	wire n7914;
	wire n7915;
	wire n7916;
	wire n7917;
	wire n7918;
	wire n7919;
	wire n7920;
	wire n7921;
	wire n7922;
	wire n7923;
	wire n7924;
	wire n7925;
	wire n7926;
	wire n7927;
	wire n7928;
	wire n7929;
	wire n7930;
	wire n7931;
	wire n7932;
	wire n7933;
	wire n7934;
	wire n7935;
	wire n7936;
	wire n7937;
	wire n7938;
	wire n7939;
	wire n7940;
	wire n7941;
	wire n7942;
	wire n7943;
	wire n7944;
	wire n7945;
	wire n7946;
	wire n7947;
	wire n7948;
	wire n7949;
	wire n7950;
	wire n7951;
	wire n7952;
	wire n7953;
	wire n7954;
	wire n7955;
	wire n7956;
	wire n7957;
	wire n7958;
	wire n7959;
	wire n7960;
	wire n7961;
	wire n7962;
	wire n7963;
	wire n7964;
	wire n7965;
	wire n7966;
	wire n7967;
	wire n7968;
	wire n7969;
	wire n7970;
	wire n7971;
	wire n7972;
	wire n7973;
	wire n7974;
	wire n7975;
	wire n7976;
	wire n7977;
	wire n7978;
	wire n7979;
	wire n7980;
	wire n7981;
	wire n7982;
	wire n7983;
	wire n7984;
	wire n7985;
	wire n7986;
	wire n7987;
	wire n7988;
	wire n7989;
	wire n7990;
	wire n7991;
	wire n7992;
	wire n7993;
	wire n7994;
	wire n7995;
	wire n7996;
	wire n7997;
	wire n7998;
	wire n7999;
	wire n8000;
	wire n8001;
	wire n8002;
	wire n8003;
	wire n8004;
	wire n8005;
	wire n8006;
	wire n8007;
	wire n8008;
	wire n8009;
	wire n8010;
	wire n8011;
	wire n8012;
	wire n8013;
	wire n8014;
	wire n8015;
	wire n8016;
	wire n8017;
	wire n8018;
	wire n8019;
	wire n8020;
	wire n8021;
	wire n8022;
	wire n8023;
	wire n8024;
	wire n8025;
	wire n8026;
	wire n8027;
	wire n8028;
	wire n8029;
	wire n8030;
	wire n8031;
	wire n8032;
	wire n8033;
	wire n8034;
	wire n8035;
	wire n8036;
	wire n8037;
	wire n8038;
	wire n8039;
	wire n8040;
	wire n8041;
	wire n8042;
	wire n8043;
	wire n8044;
	wire n8045;
	wire n8046;
	wire n8047;
	wire n8048;
	wire n8049;
	wire n8050;
	wire n8051;
	wire n8052;
	wire n8053;
	wire n8056;
	wire n8057;
	wire n8058;
	wire n8059;
	wire n8060;
	wire n8061;
	wire n8062;
	wire n8063;
	wire n8064;
	wire n8065;
	wire n8066;
	wire n8067;
	wire n8068;
	wire n8069;
	wire n8070;
	wire n8071;
	wire n8072;
	wire n8073;
	wire n8074;
	wire n8075;
	wire n8076;
	wire n8077;
	wire n8078;
	wire n8079;
	wire n8080;
	wire n8081;
	wire n8082;
	wire n8083;
	wire n8084;
	wire n8085;
	wire n8086;
	wire n8087;
	wire n8088;
	wire n8089;
	wire n8090;
	wire n8091;
	wire n8092;
	wire n8093;
	wire n8094;
	wire n8095;
	wire n8096;
	wire n8097;
	wire n8098;
	wire n8099;
	wire n8100;
	wire n8101;
	wire n8102;
	wire n8103;
	wire n8104;
	wire n8105;
	wire n8106;
	wire n8107;
	wire n8108;
	wire n8109;
	wire n8110;
	wire n8111;
	wire n8112;
	wire n8113;
	wire n8114;
	wire n8115;
	wire n8117;
	wire n8118;
	wire n8119;
	wire n8120;
	wire n8121;
	wire n8122;
	wire n8123;
	wire n8124;
	wire n8125;
	wire n8126;
	wire n8127;
	wire n8128;
	wire n8129;
	wire n8130;
	wire n8131;
	wire n8132;
	wire n8133;
	wire n8134;
	wire n8135;
	wire n8136;
	wire n8137;
	wire n8138;
	wire n8139;
	wire n8140;
	wire n8141;
	wire n8142;
	wire n8143;
	wire n8144;
	wire n8145;
	wire n8146;
	wire n8147;
	wire n8148;
	wire n8149;
	wire n8150;
	wire n8151;
	wire n8152;
	wire n8153;
	wire n8154;
	wire n8155;
	wire n8156;
	wire n8157;
	wire n8158;
	wire n8159;
	wire n8160;
	wire n8161;
	wire n8162;
	wire n8163;
	wire n8164;
	wire n8165;
	wire n8166;
	wire n8167;
	wire n8168;
	wire n8169;
	wire n8170;
	wire n8171;
	wire n8172;
	wire n8173;
	wire n8174;
	wire n8175;
	wire n8176;
	wire n8177;
	wire n8178;
	wire n8179;
	wire n8180;
	wire n8181;
	wire n8182;
	wire n8183;
	wire n8184;
	wire n8185;
	wire n8186;
	wire n8187;
	wire n8188;
	wire n8189;
	wire n8190;
	wire n8191;
	wire n8192;
	wire n8193;
	wire n8194;
	wire n8195;
	wire n8196;
	wire n8197;
	wire n8198;
	wire n8199;
	wire n8200;
	wire n8201;
	wire n8202;
	wire n8203;
	wire n8204;
	wire n8205;
	wire n8206;
	wire n8207;
	wire n8208;
	wire n8209;
	wire n8210;
	wire n8211;
	wire n8212;
	wire n8213;
	wire n8214;
	wire n8215;
	wire n8216;
	wire n8217;
	wire n8218;
	wire n8219;
	wire n8220;
	wire n8221;
	wire n8222;
	wire n8223;
	wire n8224;
	wire n8225;
	wire n8226;
	wire n8227;
	wire n8228;
	wire n8229;
	wire n8230;
	wire n8231;
	wire n8232;
	wire n8233;
	wire n8234;
	wire n8235;
	wire n8236;
	wire n8237;
	wire n8238;
	wire n8239;
	wire n8240;
	wire n8241;
	wire n8242;
	wire n8243;
	wire n8244;
	wire n8245;
	wire n8246;
	wire n8247;
	wire n8248;
	wire n8249;
	wire n8250;
	wire n8251;
	wire n8252;
	wire n8253;
	wire n8254;
	wire n8255;
	wire n8256;
	wire n8257;
	wire n8258;
	wire n8259;
	wire n8260;
	wire n8261;
	wire n8262;
	wire n8263;
	wire n8264;
	wire n8265;
	wire n8266;
	wire n8267;
	wire n8268;
	wire n8269;
	wire n8270;
	wire n8271;
	wire n8272;
	wire n8273;
	wire n8274;
	wire n8275;
	wire n8276;
	wire n8277;
	wire n8278;
	wire n8279;
	wire n8280;
	wire n8281;
	wire n8282;
	wire n8283;
	wire n8284;
	wire n8285;
	wire n8286;
	wire n8287;
	wire n8288;
	wire n8289;
	wire n8290;
	wire n8291;
	wire n8292;
	wire n8293;
	wire n8294;
	wire n8295;
	wire n8296;
	wire n8297;
	wire n8298;
	wire n8299;
	wire n8300;
	wire n8301;
	wire n8302;
	wire n8303;
	wire n8304;
	wire n8305;
	wire n8306;
	wire n8307;
	wire n8308;
	wire n8309;
	wire n8310;
	wire n8311;
	wire n8312;
	wire n8313;
	wire n8314;
	wire n8315;
	wire n8316;
	wire n8317;
	wire n8318;
	wire n8319;
	wire n8320;
	wire n8321;
	wire n8322;
	wire n8323;
	wire n8324;
	wire n8325;
	wire n8326;
	wire n8327;
	wire n8328;
	wire n8329;
	wire n8330;
	wire n8331;
	wire n8332;
	wire n8333;
	wire n8334;
	wire n8335;
	wire n8336;
	wire n8337;
	wire n8338;
	wire n8339;
	wire n8340;
	wire n8341;
	wire n8342;
	wire n8343;
	wire n8344;
	wire n8345;
	wire n8346;
	wire n8347;
	wire n8348;
	wire n8349;
	wire n8350;
	wire n8351;
	wire n8352;
	wire n8353;
	wire n8354;
	wire n8355;
	wire n8356;
	wire n8357;
	wire n8358;
	wire n8359;
	wire n8360;
	wire n8361;
	wire n8362;
	wire n8363;
	wire n8364;
	wire n8365;
	wire n8366;
	wire n8367;
	wire n8368;
	wire n8369;
	wire n8370;
	wire n8371;
	wire n8372;
	wire n8373;
	wire n8374;
	wire n8375;
	wire n8376;
	wire n8377;
	wire n8378;
	wire n8379;
	wire n8380;
	wire n8381;
	wire n8382;
	wire n8383;
	wire n8384;
	wire n8385;
	wire n8386;
	wire n8387;
	wire n8388;
	wire n8389;
	wire n8390;
	wire n8391;
	wire n8392;
	wire n8393;
	wire n8394;
	wire n8395;
	wire n8396;
	wire n8397;
	wire n8398;
	wire n8399;
	wire n8400;
	wire n8401;
	wire n8402;
	wire n8403;
	wire n8404;
	wire n8405;
	wire n8406;
	wire n8407;
	wire n8408;
	wire n8409;
	wire n8410;
	wire n8411;
	wire n8412;
	wire n8413;
	wire n8414;
	wire n8415;
	wire n8416;
	wire n8417;
	wire n8418;
	wire n8419;
	wire n8420;
	wire n8421;
	wire n8422;
	wire n8423;
	wire n8424;
	wire n8425;
	wire n8426;
	wire n8427;
	wire n8428;
	wire n8429;
	wire n8430;
	wire n8431;
	wire n8432;
	wire n8433;
	wire n8434;
	wire n8435;
	wire n8436;
	wire n8437;
	wire n8438;
	wire n8439;
	wire n8440;
	wire n8441;
	wire n8442;
	wire n8443;
	wire n8444;
	wire n8445;
	wire n8446;
	wire n8447;
	wire n8448;
	wire n8449;
	wire n8450;
	wire n8451;
	wire n8454;
	wire n8456;
	wire n8457;
	wire n8458;
	wire n8459;
	wire n8460;
	wire n8461;
	wire n8462;
	wire n8463;
	wire n8464;
	wire n8465;
	wire n8466;
	wire n8467;
	wire n8468;
	wire n8469;
	wire n8470;
	wire n8471;
	wire n8472;
	wire n8473;
	wire n8474;
	wire n8475;
	wire n8476;
	wire n8477;
	wire n8478;
	wire n8479;
	wire n8480;
	wire n8481;
	wire n8482;
	wire n8483;
	wire n8484;
	wire n8485;
	wire n8486;
	wire n8487;
	wire n8488;
	wire n8489;
	wire n8490;
	wire n8491;
	wire n8492;
	wire n8493;
	wire n8494;
	wire n8495;
	wire n8496;
	wire n8497;
	wire n8498;
	wire n8499;
	wire n8500;
	wire n8501;
	wire n8502;
	wire n8503;
	wire n8504;
	wire n8505;
	wire n8506;
	wire n8507;
	wire n8508;
	wire n8509;
	wire n8510;
	wire n8511;
	wire n8512;
	wire n8513;
	wire n8514;
	wire n8515;
	wire n8516;
	wire n8517;
	wire n8518;
	wire n8519;
	wire n8520;
	wire n8521;
	wire n8522;
	wire n8523;
	wire n8524;
	wire n8525;
	wire n8526;
	wire n8527;
	wire n8528;
	wire n8529;
	wire n8530;
	wire n8531;
	wire n8532;
	wire n8533;
	wire n8534;
	wire n8535;
	wire n8536;
	wire n8537;
	wire n8538;
	wire n8539;
	wire n8540;
	wire n8541;
	wire n8542;
	wire n8543;
	wire n8544;
	wire n8545;
	wire n8546;
	wire n8547;
	wire n8548;
	wire n8549;
	wire n8550;
	wire n8551;
	wire n8552;
	wire n8553;
	wire n8554;
	wire n8555;
	wire n8556;
	wire n8557;
	wire n8558;
	wire n8559;
	wire n8560;
	wire n8561;
	wire n8562;
	wire n8563;
	wire n8564;
	wire n8565;
	wire n8566;
	wire n8567;
	wire n8568;
	wire n8569;
	wire n8570;
	wire n8571;
	wire n8572;
	wire n8573;
	wire n8574;
	wire n8575;
	wire n8576;
	wire n8577;
	wire n8578;
	wire n8579;
	wire n8580;
	wire n8581;
	wire n8582;
	wire n8583;
	wire n8584;
	wire n8585;
	wire n8586;
	wire n8587;
	wire n8588;
	wire n8589;
	wire n8590;
	wire n8591;
	wire n8592;
	wire n8593;
	wire n8594;
	wire n8595;
	wire n8596;
	wire n8597;
	wire n8598;
	wire n8599;
	wire n8600;
	wire n8601;
	wire n8602;
	wire n8603;
	wire n8604;
	wire n8605;
	wire n8606;
	wire n8607;
	wire n8608;
	wire n8609;
	wire n8610;
	wire n8611;
	wire n8612;
	wire n8613;
	wire n8614;
	wire n8615;
	wire n8616;
	wire n8617;
	wire n8618;
	wire n8619;
	wire n8620;
	wire n8621;
	wire n8622;
	wire n8623;
	wire n8624;
	wire n8625;
	wire n8626;
	wire n8627;
	wire n8628;
	wire n8629;
	wire n8630;
	wire n8631;
	wire n8632;
	wire n8633;
	wire n8634;
	wire n8635;
	wire n8636;
	wire n8637;
	wire n8638;
	wire n8639;
	wire n8640;
	wire n8641;
	wire n8642;
	wire n8643;
	wire n8644;
	wire n8645;
	wire n8646;
	wire n8647;
	wire n8648;
	wire n8649;
	wire n8650;
	wire n8651;
	wire n8652;
	wire n8653;
	wire n8654;
	wire n8655;
	wire n8656;
	wire n8657;
	wire n8658;
	wire n8659;
	wire n8660;
	wire n8661;
	wire n8662;
	wire n8663;
	wire n8664;
	wire n8665;
	wire n8666;
	wire n8667;
	wire n8668;
	wire n8669;
	wire n8670;
	wire n8671;
	wire n8672;
	wire n8673;
	wire n8674;
	wire n8675;
	wire n8676;
	wire n8677;
	wire n8678;
	wire n8679;
	wire n8680;
	wire n8681;
	wire n8682;
	wire n8683;
	wire n8684;
	wire n8685;
	wire n8686;
	wire n8687;
	wire n8688;
	wire n8689;
	wire n8690;
	wire n8691;
	wire n8692;
	wire n8693;
	wire n8694;
	wire n8695;
	wire n8696;
	wire n8697;
	wire n8698;
	wire n8699;
	wire n8700;
	wire n8701;
	wire n8702;
	wire n8703;
	wire n8704;
	wire n8705;
	wire n8706;
	wire n8707;
	wire n8708;
	wire n8709;
	wire n8710;
	wire n8711;
	wire n8712;
	wire n8713;
	wire n8714;
	wire n8715;
	wire n8716;
	wire n8717;
	wire n8718;
	wire n8719;
	wire n8720;
	wire n8721;
	wire n8722;
	wire n8723;
	wire n8724;
	wire n8725;
	wire n8726;
	wire n8727;
	wire n8728;
	wire n8729;
	wire n8730;
	wire n8731;
	wire n8732;
	wire n8733;
	wire n8734;
	wire n8735;
	wire n8736;
	wire n8737;
	wire n8738;
	wire n8739;
	wire n8740;
	wire n8741;
	wire n8742;
	wire n8743;
	wire n8744;
	wire n8745;
	wire n8746;
	wire n8747;
	wire n8748;
	wire n8749;
	wire n8750;
	wire n8751;
	wire n8752;
	wire n8753;
	wire n8754;
	wire n8755;
	wire n8756;
	wire n8757;
	wire n8758;
	wire n8759;
	wire n8760;
	wire n8761;
	wire n8762;
	wire n8763;
	wire n8764;
	wire n8765;
	wire n8766;
	wire n8767;
	wire n8768;
	wire n8769;
	wire n8770;
	wire n8771;
	wire n8772;
	wire n8773;
	wire n8774;
	wire n8775;
	wire n8776;
	wire n8777;
	wire n8778;
	wire n8779;
	wire n8780;
	wire n8781;
	wire n8782;
	wire n8783;
	wire n8784;
	wire n8785;
	wire n8786;
	wire n8787;
	wire n8788;
	wire n8789;
	wire n8790;
	wire n8791;
	wire n8792;
	wire n8793;
	wire n8794;
	wire n8795;
	wire n8796;
	wire n8797;
	wire n8798;
	wire n8799;
	wire n8800;
	wire n8801;
	wire n8802;
	wire n8803;
	wire n8804;
	wire n8805;
	wire n8806;
	wire n8807;
	wire n8808;
	wire n8809;
	wire n8810;
	wire n8811;
	wire n8812;
	wire n8813;
	wire n8814;
	wire n8815;
	wire n8816;
	wire n8817;
	wire n8818;
	wire n8819;
	wire n8820;
	wire n8821;
	wire n8822;
	wire n8823;
	wire n8824;
	wire n8825;
	wire n8826;
	wire n8827;
	wire n8828;
	wire n8829;
	wire n8830;
	wire n8831;
	wire n8832;
	wire n8833;
	wire n8834;
	wire n8835;
	wire n8836;
	wire n8837;
	wire n8838;
	wire n8839;
	wire n8840;
	wire n8841;
	wire n8842;
	wire n8843;
	wire n8844;
	wire n8845;
	wire n8846;
	wire n8847;
	wire n8848;
	wire n8849;
	wire n8850;
	wire n8851;
	wire n8852;
	wire n8853;
	wire n8854;
	wire n8855;
	wire n8856;
	wire n8857;
	wire n8858;
	wire n8859;
	wire n8860;
	wire n8861;
	wire n8862;
	wire n8863;
	wire n8864;
	wire n8865;
	wire n8866;
	wire n8867;
	wire n8868;
	wire n8869;
	wire n8870;
	wire n8871;
	wire n8872;
	wire n8873;
	wire n8874;
	wire n8875;
	wire n8876;
	wire n8877;
	wire n8878;
	wire n8879;
	wire n8880;
	wire n8881;
	wire n8882;
	wire n8883;
	wire n8884;
	wire n8885;
	wire n8886;
	wire n8887;
	wire n8888;
	wire n8889;
	wire n8890;
	wire n8891;
	wire n8892;
	wire n8893;
	wire n8896;
	wire n8897;
	wire n8898;
	wire n8899;
	wire n8900;
	wire n8901;
	wire n8902;
	wire n8903;
	wire n8904;
	wire n8905;
	wire n8906;
	wire n8907;
	wire n8908;
	wire n8909;
	wire n8910;
	wire n8911;
	wire n8912;
	wire n8913;
	wire n8914;
	wire n8915;
	wire n8916;
	wire n8917;
	wire n8918;
	wire n8919;
	wire n8920;
	wire n8921;
	wire n8922;
	wire n8923;
	wire n8924;
	wire n8925;
	wire n8926;
	wire n8927;
	wire n8928;
	wire n8929;
	wire n8930;
	wire n8931;
	wire n8932;
	wire n8933;
	wire n8934;
	wire n8935;
	wire n8936;
	wire n8937;
	wire n8938;
	wire n8939;
	wire n8940;
	wire n8941;
	wire n8942;
	wire n8943;
	wire n8944;
	wire n8945;
	wire n8946;
	wire n8947;
	wire n8948;
	wire n8949;
	wire n8950;
	wire n8951;
	wire n8952;
	wire n8953;
	wire n8954;
	wire n8955;
	wire n8957;
	wire n8958;
	wire n8959;
	wire n8960;
	wire n8961;
	wire n8962;
	wire n8963;
	wire n8964;
	wire n8965;
	wire n8966;
	wire n8967;
	wire n8968;
	wire n8969;
	wire n8970;
	wire n8971;
	wire n8972;
	wire n8973;
	wire n8974;
	wire n8975;
	wire n8976;
	wire n8977;
	wire n8978;
	wire n8979;
	wire n8980;
	wire n8981;
	wire n8982;
	wire n8983;
	wire n8984;
	wire n8985;
	wire n8986;
	wire n8987;
	wire n8988;
	wire n8989;
	wire n8990;
	wire n8991;
	wire n8992;
	wire n8993;
	wire n8994;
	wire n8995;
	wire n8996;
	wire n8997;
	wire n8998;
	wire n8999;
	wire n9000;
	wire n9001;
	wire n9002;
	wire n9003;
	wire n9004;
	wire n9005;
	wire n9006;
	wire n9007;
	wire n9008;
	wire n9009;
	wire n9010;
	wire n9011;
	wire n9012;
	wire n9013;
	wire n9014;
	wire n9015;
	wire n9016;
	wire n9017;
	wire n9018;
	wire n9019;
	wire n9020;
	wire n9021;
	wire n9022;
	wire n9023;
	wire n9024;
	wire n9025;
	wire n9026;
	wire n9027;
	wire n9028;
	wire n9029;
	wire n9030;
	wire n9031;
	wire n9032;
	wire n9033;
	wire n9034;
	wire n9035;
	wire n9036;
	wire n9037;
	wire n9038;
	wire n9039;
	wire n9040;
	wire n9041;
	wire n9042;
	wire n9043;
	wire n9044;
	wire n9045;
	wire n9046;
	wire n9047;
	wire n9048;
	wire n9049;
	wire n9050;
	wire n9051;
	wire n9052;
	wire n9053;
	wire n9054;
	wire n9055;
	wire n9056;
	wire n9057;
	wire n9058;
	wire n9059;
	wire n9060;
	wire n9061;
	wire n9062;
	wire n9063;
	wire n9064;
	wire n9065;
	wire n9066;
	wire n9067;
	wire n9068;
	wire n9069;
	wire n9070;
	wire n9071;
	wire n9072;
	wire n9073;
	wire n9074;
	wire n9075;
	wire n9076;
	wire n9077;
	wire n9078;
	wire n9079;
	wire n9080;
	wire n9081;
	wire n9082;
	wire n9083;
	wire n9084;
	wire n9085;
	wire n9086;
	wire n9087;
	wire n9088;
	wire n9089;
	wire n9090;
	wire n9091;
	wire n9092;
	wire n9093;
	wire n9094;
	wire n9095;
	wire n9096;
	wire n9097;
	wire n9098;
	wire n9099;
	wire n9100;
	wire n9101;
	wire n9102;
	wire n9103;
	wire n9104;
	wire n9105;
	wire n9106;
	wire n9107;
	wire n9108;
	wire n9109;
	wire n9110;
	wire n9111;
	wire n9112;
	wire n9113;
	wire n9114;
	wire n9115;
	wire n9116;
	wire n9117;
	wire n9118;
	wire n9119;
	wire n9120;
	wire n9121;
	wire n9122;
	wire n9123;
	wire n9124;
	wire n9125;
	wire n9126;
	wire n9127;
	wire n9128;
	wire n9129;
	wire n9130;
	wire n9131;
	wire n9132;
	wire n9133;
	wire n9134;
	wire n9135;
	wire n9136;
	wire n9137;
	wire n9138;
	wire n9139;
	wire n9140;
	wire n9141;
	wire n9142;
	wire n9143;
	wire n9144;
	wire n9145;
	wire n9146;
	wire n9147;
	wire n9148;
	wire n9149;
	wire n9150;
	wire n9151;
	wire n9152;
	wire n9153;
	wire n9154;
	wire n9155;
	wire n9156;
	wire n9157;
	wire n9158;
	wire n9159;
	wire n9160;
	wire n9161;
	wire n9162;
	wire n9163;
	wire n9164;
	wire n9165;
	wire n9166;
	wire n9167;
	wire n9168;
	wire n9169;
	wire n9170;
	wire n9171;
	wire n9172;
	wire n9173;
	wire n9174;
	wire n9175;
	wire n9176;
	wire n9177;
	wire n9178;
	wire n9179;
	wire n9180;
	wire n9181;
	wire n9182;
	wire n9183;
	wire n9184;
	wire n9185;
	wire n9186;
	wire n9187;
	wire n9188;
	wire n9189;
	wire n9190;
	wire n9191;
	wire n9192;
	wire n9193;
	wire n9194;
	wire n9195;
	wire n9196;
	wire n9197;
	wire n9198;
	wire n9199;
	wire n9200;
	wire n9201;
	wire n9202;
	wire n9203;
	wire n9204;
	wire n9205;
	wire n9206;
	wire n9207;
	wire n9208;
	wire n9209;
	wire n9210;
	wire n9211;
	wire n9212;
	wire n9213;
	wire n9214;
	wire n9215;
	wire n9216;
	wire n9217;
	wire n9218;
	wire n9219;
	wire n9220;
	wire n9221;
	wire n9222;
	wire n9223;
	wire n9224;
	wire n9225;
	wire n9226;
	wire n9227;
	wire n9228;
	wire n9229;
	wire n9230;
	wire n9231;
	wire n9232;
	wire n9233;
	wire n9234;
	wire n9235;
	wire n9236;
	wire n9237;
	wire n9238;
	wire n9239;
	wire n9240;
	wire n9241;
	wire n9242;
	wire n9243;
	wire n9244;
	wire n9245;
	wire n9246;
	wire n9247;
	wire n9248;
	wire n9249;
	wire n9250;
	wire n9251;
	wire n9252;
	wire n9253;
	wire n9254;
	wire n9255;
	wire n9256;
	wire n9257;
	wire n9258;
	wire n9259;
	wire n9260;
	wire n9261;
	wire n9262;
	wire n9263;
	wire n9264;
	wire n9265;
	wire n9266;
	wire n9267;
	wire n9268;
	wire n9269;
	wire n9270;
	wire n9271;
	wire n9272;
	wire n9273;
	wire n9274;
	wire n9275;
	wire n9276;
	wire n9277;
	wire n9278;
	wire n9279;
	wire n9280;
	wire n9281;
	wire n9282;
	wire n9283;
	wire n9284;
	wire n9285;
	wire n9286;
	wire n9287;
	wire n9288;
	wire n9289;
	wire n9290;
	wire n9291;
	wire n9292;
	wire n9293;
	wire n9294;
	wire n9295;
	wire n9296;
	wire n9297;
	wire n9298;
	wire n9299;
	wire n9300;
	wire n9301;
	wire n9302;
	wire n9303;
	wire n9304;
	wire n9305;
	wire n9306;
	wire n9307;
	wire n9308;
	wire n9311;
	wire n9313;
	wire n9314;
	wire n9315;
	wire n9316;
	wire n9317;
	wire n9318;
	wire n9319;
	wire n9320;
	wire n9321;
	wire n9322;
	wire n9323;
	wire n9324;
	wire n9325;
	wire n9326;
	wire n9327;
	wire n9328;
	wire n9329;
	wire n9330;
	wire n9331;
	wire n9332;
	wire n9333;
	wire n9334;
	wire n9335;
	wire n9336;
	wire n9337;
	wire n9338;
	wire n9339;
	wire n9340;
	wire n9341;
	wire n9342;
	wire n9343;
	wire n9344;
	wire n9345;
	wire n9346;
	wire n9347;
	wire n9348;
	wire n9349;
	wire n9350;
	wire n9351;
	wire n9352;
	wire n9353;
	wire n9354;
	wire n9355;
	wire n9356;
	wire n9357;
	wire n9358;
	wire n9359;
	wire n9360;
	wire n9361;
	wire n9362;
	wire n9363;
	wire n9364;
	wire n9365;
	wire n9366;
	wire n9367;
	wire n9368;
	wire n9369;
	wire n9370;
	wire n9371;
	wire n9372;
	wire n9373;
	wire n9374;
	wire n9375;
	wire n9376;
	wire n9377;
	wire n9378;
	wire n9379;
	wire n9380;
	wire n9381;
	wire n9382;
	wire n9383;
	wire n9384;
	wire n9385;
	wire n9386;
	wire n9387;
	wire n9388;
	wire n9389;
	wire n9390;
	wire n9391;
	wire n9392;
	wire n9393;
	wire n9394;
	wire n9395;
	wire n9396;
	wire n9397;
	wire n9398;
	wire n9399;
	wire n9400;
	wire n9401;
	wire n9402;
	wire n9403;
	wire n9404;
	wire n9405;
	wire n9406;
	wire n9407;
	wire n9408;
	wire n9409;
	wire n9410;
	wire n9411;
	wire n9412;
	wire n9413;
	wire n9414;
	wire n9415;
	wire n9416;
	wire n9417;
	wire n9418;
	wire n9419;
	wire n9420;
	wire n9421;
	wire n9422;
	wire n9423;
	wire n9424;
	wire n9425;
	wire n9426;
	wire n9427;
	wire n9428;
	wire n9429;
	wire n9430;
	wire n9431;
	wire n9432;
	wire n9433;
	wire n9434;
	wire n9435;
	wire n9436;
	wire n9437;
	wire n9438;
	wire n9439;
	wire n9440;
	wire n9441;
	wire n9442;
	wire n9443;
	wire n9444;
	wire n9445;
	wire n9446;
	wire n9447;
	wire n9448;
	wire n9449;
	wire n9450;
	wire n9451;
	wire n9452;
	wire n9453;
	wire n9454;
	wire n9455;
	wire n9456;
	wire n9457;
	wire n9458;
	wire n9459;
	wire n9460;
	wire n9461;
	wire n9462;
	wire n9463;
	wire n9464;
	wire n9465;
	wire n9466;
	wire n9467;
	wire n9468;
	wire n9469;
	wire n9470;
	wire n9471;
	wire n9472;
	wire n9473;
	wire n9474;
	wire n9475;
	wire n9476;
	wire n9477;
	wire n9478;
	wire n9479;
	wire n9480;
	wire n9481;
	wire n9482;
	wire n9483;
	wire n9484;
	wire n9485;
	wire n9486;
	wire n9487;
	wire n9488;
	wire n9489;
	wire n9490;
	wire n9491;
	wire n9492;
	wire n9493;
	wire n9494;
	wire n9495;
	wire n9496;
	wire n9497;
	wire n9498;
	wire n9499;
	wire n9500;
	wire n9501;
	wire n9502;
	wire n9503;
	wire n9504;
	wire n9505;
	wire n9506;
	wire n9507;
	wire n9508;
	wire n9509;
	wire n9510;
	wire n9511;
	wire n9512;
	wire n9513;
	wire n9514;
	wire n9515;
	wire n9516;
	wire n9517;
	wire n9518;
	wire n9519;
	wire n9520;
	wire n9521;
	wire n9522;
	wire n9523;
	wire n9524;
	wire n9525;
	wire n9526;
	wire n9527;
	wire n9528;
	wire n9529;
	wire n9530;
	wire n9531;
	wire n9532;
	wire n9533;
	wire n9534;
	wire n9535;
	wire n9536;
	wire n9537;
	wire n9538;
	wire n9539;
	wire n9540;
	wire n9541;
	wire n9542;
	wire n9543;
	wire n9544;
	wire n9545;
	wire n9546;
	wire n9547;
	wire n9548;
	wire n9549;
	wire n9550;
	wire n9551;
	wire n9552;
	wire n9553;
	wire n9554;
	wire n9555;
	wire n9556;
	wire n9557;
	wire n9558;
	wire n9559;
	wire n9560;
	wire n9561;
	wire n9562;
	wire n9563;
	wire n9564;
	wire n9565;
	wire n9566;
	wire n9567;
	wire n9568;
	wire n9569;
	wire n9570;
	wire n9571;
	wire n9572;
	wire n9573;
	wire n9574;
	wire n9575;
	wire n9576;
	wire n9577;
	wire n9578;
	wire n9579;
	wire n9580;
	wire n9581;
	wire n9582;
	wire n9583;
	wire n9584;
	wire n9585;
	wire n9586;
	wire n9587;
	wire n9588;
	wire n9589;
	wire n9590;
	wire n9591;
	wire n9592;
	wire n9593;
	wire n9594;
	wire n9595;
	wire n9596;
	wire n9597;
	wire n9598;
	wire n9599;
	wire n9600;
	wire n9601;
	wire n9602;
	wire n9603;
	wire n9604;
	wire n9605;
	wire n9606;
	wire n9607;
	wire n9608;
	wire n9609;
	wire n9610;
	wire n9611;
	wire n9612;
	wire n9613;
	wire n9614;
	wire n9615;
	wire n9616;
	wire n9617;
	wire n9618;
	wire n9619;
	wire n9620;
	wire n9621;
	wire n9622;
	wire n9623;
	wire n9624;
	wire n9625;
	wire n9626;
	wire n9627;
	wire n9628;
	wire n9629;
	wire n9630;
	wire n9631;
	wire n9632;
	wire n9633;
	wire n9634;
	wire n9635;
	wire n9636;
	wire n9637;
	wire n9638;
	wire n9639;
	wire n9640;
	wire n9641;
	wire n9642;
	wire n9643;
	wire n9644;
	wire n9645;
	wire n9646;
	wire n9647;
	wire n9648;
	wire n9649;
	wire n9650;
	wire n9651;
	wire n9652;
	wire n9653;
	wire n9654;
	wire n9655;
	wire n9656;
	wire n9657;
	wire n9658;
	wire n9659;
	wire n9660;
	wire n9661;
	wire n9662;
	wire n9663;
	wire n9664;
	wire n9665;
	wire n9666;
	wire n9667;
	wire n9668;
	wire n9669;
	wire n9670;
	wire n9671;
	wire n9672;
	wire n9673;
	wire n9674;
	wire n9675;
	wire n9676;
	wire n9677;
	wire n9678;
	wire n9679;
	wire n9680;
	wire n9681;
	wire n9682;
	wire n9683;
	wire n9684;
	wire n9685;
	wire n9686;
	wire n9687;
	wire n9688;
	wire n9689;
	wire n9690;
	wire n9691;
	wire n9692;
	wire n9693;
	wire n9694;
	wire n9695;
	wire n9696;
	wire n9697;
	wire n9698;
	wire n9699;
	wire n9700;
	wire n9701;
	wire n9702;
	wire n9703;
	wire n9704;
	wire n9705;
	wire n9706;
	wire n9707;
	wire n9708;
	wire n9709;
	wire n9710;
	wire n9711;
	wire n9712;
	wire n9713;
	wire n9714;
	wire n9715;
	wire n9716;
	wire n9717;
	wire n9718;
	wire n9719;
	wire n9720;
	wire n9721;
	wire n9722;
	wire n9723;
	wire n9724;
	wire n9725;
	wire n9726;
	wire n9727;
	wire n9728;
	wire n9729;
	wire n9730;
	wire n9731;
	wire n9732;
	wire n9733;
	wire n9734;
	wire n9735;
	wire n9736;
	wire n9737;
	wire n9738;
	wire n9739;
	wire n9740;
	wire n9741;
	wire n9742;
	wire n9743;
	wire n9744;
	wire n9745;
	wire n9746;
	wire n9747;
	wire n9748;
	wire n9749;
	wire n9750;
	wire n9751;
	wire n9752;
	wire n9753;
	wire n9754;
	wire n9755;
	wire n9756;
	wire n9757;
	wire n9758;
	wire n9759;
	wire n9760;
	wire n9761;
	wire n9762;
	wire n9763;
	wire n9764;
	wire n9765;
	wire n9766;
	wire n9767;
	wire n9768;
	wire n9769;
	wire n9772;
	wire n9773;
	wire n9774;
	wire n9775;
	wire n9776;
	wire n9777;
	wire n9778;
	wire n9779;
	wire n9780;
	wire n9781;
	wire n9782;
	wire n9783;
	wire n9784;
	wire n9785;
	wire n9786;
	wire n9787;
	wire n9788;
	wire n9789;
	wire n9790;
	wire n9791;
	wire n9792;
	wire n9793;
	wire n9794;
	wire n9795;
	wire n9796;
	wire n9797;
	wire n9798;
	wire n9799;
	wire n9800;
	wire n9801;
	wire n9802;
	wire n9803;
	wire n9804;
	wire n9805;
	wire n9806;
	wire n9807;
	wire n9808;
	wire n9809;
	wire n9810;
	wire n9811;
	wire n9812;
	wire n9813;
	wire n9814;
	wire n9815;
	wire n9816;
	wire n9817;
	wire n9818;
	wire n9819;
	wire n9820;
	wire n9821;
	wire n9822;
	wire n9823;
	wire n9824;
	wire n9825;
	wire n9826;
	wire n9827;
	wire n9828;
	wire n9829;
	wire n9830;
	wire n9831;
	wire n9832;
	wire n9834;
	wire n9835;
	wire n9836;
	wire n9837;
	wire n9838;
	wire n9839;
	wire n9840;
	wire n9841;
	wire n9842;
	wire n9843;
	wire n9844;
	wire n9845;
	wire n9846;
	wire n9847;
	wire n9848;
	wire n9849;
	wire n9850;
	wire n9851;
	wire n9852;
	wire n9853;
	wire n9854;
	wire n9855;
	wire n9856;
	wire n9857;
	wire n9858;
	wire n9859;
	wire n9860;
	wire n9861;
	wire n9862;
	wire n9863;
	wire n9864;
	wire n9865;
	wire n9866;
	wire n9867;
	wire n9868;
	wire n9869;
	wire n9870;
	wire n9871;
	wire n9872;
	wire n9873;
	wire n9874;
	wire n9875;
	wire n9876;
	wire n9877;
	wire n9878;
	wire n9879;
	wire n9880;
	wire n9881;
	wire n9882;
	wire n9883;
	wire n9884;
	wire n9885;
	wire n9886;
	wire n9887;
	wire n9888;
	wire n9889;
	wire n9890;
	wire n9891;
	wire n9892;
	wire n9893;
	wire n9894;
	wire n9895;
	wire n9896;
	wire n9897;
	wire n9898;
	wire n9899;
	wire n9900;
	wire n9901;
	wire n9902;
	wire n9903;
	wire n9904;
	wire n9905;
	wire n9906;
	wire n9907;
	wire n9908;
	wire n9909;
	wire n9910;
	wire n9911;
	wire n9912;
	wire n9913;
	wire n9914;
	wire n9915;
	wire n9916;
	wire n9917;
	wire n9918;
	wire n9919;
	wire n9920;
	wire n9921;
	wire n9922;
	wire n9923;
	wire n9924;
	wire n9925;
	wire n9926;
	wire n9927;
	wire n9928;
	wire n9929;
	wire n9930;
	wire n9931;
	wire n9932;
	wire n9933;
	wire n9934;
	wire n9935;
	wire n9936;
	wire n9937;
	wire n9938;
	wire n9939;
	wire n9940;
	wire n9941;
	wire n9942;
	wire n9943;
	wire n9944;
	wire n9945;
	wire n9946;
	wire n9947;
	wire n9948;
	wire n9949;
	wire n9950;
	wire n9951;
	wire n9952;
	wire n9953;
	wire n9954;
	wire n9955;
	wire n9956;
	wire n9957;
	wire n9958;
	wire n9959;
	wire n9960;
	wire n9961;
	wire n9962;
	wire n9963;
	wire n9964;
	wire n9965;
	wire n9966;
	wire n9967;
	wire n9968;
	wire n9969;
	wire n9970;
	wire n9971;
	wire n9972;
	wire n9973;
	wire n9974;
	wire n9975;
	wire n9976;
	wire n9977;
	wire n9978;
	wire n9979;
	wire n9980;
	wire n9981;
	wire n9982;
	wire n9983;
	wire n9984;
	wire n9985;
	wire n9986;
	wire n9987;
	wire n9988;
	wire n9989;
	wire n9990;
	wire n9991;
	wire n9992;
	wire n9993;
	wire n9994;
	wire n9995;
	wire n9996;
	wire n9997;
	wire n9998;
	wire n9999;
	wire n10000;
	wire n10001;
	wire n10002;
	wire n10003;
	wire n10004;
	wire n10005;
	wire n10006;
	wire n10007;
	wire n10008;
	wire n10009;
	wire n10010;
	wire n10011;
	wire n10012;
	wire n10013;
	wire n10014;
	wire n10015;
	wire n10016;
	wire n10017;
	wire n10018;
	wire n10019;
	wire n10020;
	wire n10021;
	wire n10022;
	wire n10023;
	wire n10024;
	wire n10025;
	wire n10026;
	wire n10027;
	wire n10028;
	wire n10029;
	wire n10030;
	wire n10031;
	wire n10032;
	wire n10033;
	wire n10034;
	wire n10035;
	wire n10036;
	wire n10037;
	wire n10038;
	wire n10039;
	wire n10040;
	wire n10041;
	wire n10042;
	wire n10043;
	wire n10044;
	wire n10045;
	wire n10046;
	wire n10047;
	wire n10048;
	wire n10049;
	wire n10050;
	wire n10051;
	wire n10052;
	wire n10053;
	wire n10054;
	wire n10055;
	wire n10056;
	wire n10057;
	wire n10058;
	wire n10059;
	wire n10060;
	wire n10061;
	wire n10062;
	wire n10063;
	wire n10064;
	wire n10065;
	wire n10066;
	wire n10067;
	wire n10068;
	wire n10069;
	wire n10070;
	wire n10071;
	wire n10072;
	wire n10073;
	wire n10074;
	wire n10075;
	wire n10076;
	wire n10077;
	wire n10078;
	wire n10079;
	wire n10080;
	wire n10081;
	wire n10082;
	wire n10083;
	wire n10084;
	wire n10085;
	wire n10086;
	wire n10087;
	wire n10088;
	wire n10089;
	wire n10090;
	wire n10091;
	wire n10092;
	wire n10093;
	wire n10094;
	wire n10095;
	wire n10096;
	wire n10097;
	wire n10098;
	wire n10099;
	wire n10100;
	wire n10101;
	wire n10102;
	wire n10103;
	wire n10104;
	wire n10105;
	wire n10106;
	wire n10107;
	wire n10108;
	wire n10109;
	wire n10110;
	wire n10111;
	wire n10112;
	wire n10113;
	wire n10114;
	wire n10115;
	wire n10116;
	wire n10117;
	wire n10118;
	wire n10119;
	wire n10120;
	wire n10121;
	wire n10122;
	wire n10123;
	wire n10124;
	wire n10125;
	wire n10126;
	wire n10127;
	wire n10128;
	wire n10129;
	wire n10130;
	wire n10131;
	wire n10132;
	wire n10133;
	wire n10134;
	wire n10135;
	wire n10136;
	wire n10137;
	wire n10138;
	wire n10139;
	wire n10140;
	wire n10141;
	wire n10142;
	wire n10143;
	wire n10144;
	wire n10145;
	wire n10146;
	wire n10147;
	wire n10148;
	wire n10149;
	wire n10150;
	wire n10151;
	wire n10152;
	wire n10153;
	wire n10154;
	wire n10155;
	wire n10156;
	wire n10157;
	wire n10158;
	wire n10159;
	wire n10160;
	wire n10161;
	wire n10162;
	wire n10163;
	wire n10164;
	wire n10165;
	wire n10166;
	wire n10167;
	wire n10168;
	wire n10169;
	wire n10170;
	wire n10171;
	wire n10172;
	wire n10173;
	wire n10174;
	wire n10175;
	wire n10176;
	wire n10177;
	wire n10178;
	wire n10179;
	wire n10180;
	wire n10181;
	wire n10182;
	wire n10183;
	wire n10184;
	wire n10185;
	wire n10186;
	wire n10187;
	wire n10188;
	wire n10189;
	wire n10190;
	wire n10191;
	wire n10192;
	wire n10193;
	wire n10194;
	wire n10195;
	wire n10196;
	wire n10197;
	wire n10198;
	wire n10199;
	wire n10200;
	wire n10201;
	wire n10202;
	wire n10203;
	wire n10204;
	wire n10205;
	wire n10206;
	wire n10207;
	wire n10208;
	wire n10209;
	wire n10212;
	wire n10214;
	wire n10215;
	wire n10216;
	wire n10217;
	wire n10218;
	wire n10219;
	wire n10220;
	wire n10221;
	wire n10222;
	wire n10223;
	wire n10224;
	wire n10225;
	wire n10226;
	wire n10227;
	wire n10228;
	wire n10229;
	wire n10230;
	wire n10231;
	wire n10232;
	wire n10233;
	wire n10234;
	wire n10235;
	wire n10236;
	wire n10237;
	wire n10238;
	wire n10239;
	wire n10240;
	wire n10241;
	wire n10242;
	wire n10243;
	wire n10244;
	wire n10245;
	wire n10246;
	wire n10247;
	wire n10248;
	wire n10249;
	wire n10250;
	wire n10251;
	wire n10252;
	wire n10253;
	wire n10254;
	wire n10255;
	wire n10256;
	wire n10257;
	wire n10258;
	wire n10259;
	wire n10260;
	wire n10261;
	wire n10262;
	wire n10263;
	wire n10264;
	wire n10265;
	wire n10266;
	wire n10267;
	wire n10268;
	wire n10269;
	wire n10270;
	wire n10271;
	wire n10272;
	wire n10273;
	wire n10274;
	wire n10275;
	wire n10276;
	wire n10277;
	wire n10278;
	wire n10279;
	wire n10280;
	wire n10281;
	wire n10282;
	wire n10283;
	wire n10284;
	wire n10285;
	wire n10286;
	wire n10287;
	wire n10288;
	wire n10289;
	wire n10290;
	wire n10291;
	wire n10292;
	wire n10293;
	wire n10294;
	wire n10295;
	wire n10296;
	wire n10297;
	wire n10298;
	wire n10299;
	wire n10300;
	wire n10301;
	wire n10302;
	wire n10303;
	wire n10304;
	wire n10305;
	wire n10306;
	wire n10307;
	wire n10308;
	wire n10309;
	wire n10310;
	wire n10311;
	wire n10312;
	wire n10313;
	wire n10314;
	wire n10315;
	wire n10316;
	wire n10317;
	wire n10318;
	wire n10319;
	wire n10320;
	wire n10321;
	wire n10322;
	wire n10323;
	wire n10324;
	wire n10325;
	wire n10326;
	wire n10327;
	wire n10328;
	wire n10329;
	wire n10330;
	wire n10331;
	wire n10332;
	wire n10333;
	wire n10334;
	wire n10335;
	wire n10336;
	wire n10337;
	wire n10338;
	wire n10339;
	wire n10340;
	wire n10341;
	wire n10342;
	wire n10343;
	wire n10344;
	wire n10345;
	wire n10346;
	wire n10347;
	wire n10348;
	wire n10349;
	wire n10350;
	wire n10351;
	wire n10352;
	wire n10353;
	wire n10354;
	wire n10355;
	wire n10356;
	wire n10357;
	wire n10358;
	wire n10359;
	wire n10360;
	wire n10361;
	wire n10362;
	wire n10363;
	wire n10364;
	wire n10365;
	wire n10366;
	wire n10367;
	wire n10368;
	wire n10369;
	wire n10370;
	wire n10371;
	wire n10372;
	wire n10373;
	wire n10374;
	wire n10375;
	wire n10376;
	wire n10377;
	wire n10378;
	wire n10379;
	wire n10380;
	wire n10381;
	wire n10382;
	wire n10383;
	wire n10384;
	wire n10385;
	wire n10386;
	wire n10387;
	wire n10388;
	wire n10389;
	wire n10390;
	wire n10391;
	wire n10392;
	wire n10393;
	wire n10394;
	wire n10395;
	wire n10396;
	wire n10397;
	wire n10398;
	wire n10399;
	wire n10400;
	wire n10401;
	wire n10402;
	wire n10403;
	wire n10404;
	wire n10405;
	wire n10406;
	wire n10407;
	wire n10408;
	wire n10409;
	wire n10410;
	wire n10411;
	wire n10412;
	wire n10413;
	wire n10414;
	wire n10415;
	wire n10416;
	wire n10417;
	wire n10418;
	wire n10419;
	wire n10420;
	wire n10421;
	wire n10422;
	wire n10423;
	wire n10424;
	wire n10425;
	wire n10426;
	wire n10427;
	wire n10428;
	wire n10429;
	wire n10430;
	wire n10431;
	wire n10432;
	wire n10433;
	wire n10434;
	wire n10435;
	wire n10436;
	wire n10437;
	wire n10438;
	wire n10439;
	wire n10440;
	wire n10441;
	wire n10442;
	wire n10443;
	wire n10444;
	wire n10445;
	wire n10446;
	wire n10447;
	wire n10448;
	wire n10449;
	wire n10450;
	wire n10451;
	wire n10452;
	wire n10453;
	wire n10454;
	wire n10455;
	wire n10456;
	wire n10457;
	wire n10458;
	wire n10459;
	wire n10460;
	wire n10461;
	wire n10462;
	wire n10463;
	wire n10464;
	wire n10465;
	wire n10466;
	wire n10467;
	wire n10468;
	wire n10469;
	wire n10470;
	wire n10471;
	wire n10472;
	wire n10473;
	wire n10474;
	wire n10475;
	wire n10476;
	wire n10477;
	wire n10478;
	wire n10479;
	wire n10480;
	wire n10481;
	wire n10482;
	wire n10483;
	wire n10484;
	wire n10485;
	wire n10486;
	wire n10487;
	wire n10488;
	wire n10489;
	wire n10490;
	wire n10491;
	wire n10492;
	wire n10493;
	wire n10494;
	wire n10495;
	wire n10496;
	wire n10497;
	wire n10498;
	wire n10499;
	wire n10500;
	wire n10501;
	wire n10502;
	wire n10503;
	wire n10504;
	wire n10505;
	wire n10506;
	wire n10507;
	wire n10508;
	wire n10509;
	wire n10510;
	wire n10511;
	wire n10512;
	wire n10513;
	wire n10514;
	wire n10515;
	wire n10516;
	wire n10517;
	wire n10518;
	wire n10519;
	wire n10520;
	wire n10521;
	wire n10522;
	wire n10523;
	wire n10524;
	wire n10525;
	wire n10526;
	wire n10527;
	wire n10528;
	wire n10529;
	wire n10530;
	wire n10531;
	wire n10532;
	wire n10533;
	wire n10534;
	wire n10535;
	wire n10536;
	wire n10537;
	wire n10538;
	wire n10539;
	wire n10540;
	wire n10541;
	wire n10542;
	wire n10543;
	wire n10544;
	wire n10545;
	wire n10546;
	wire n10547;
	wire n10548;
	wire n10549;
	wire n10550;
	wire n10551;
	wire n10552;
	wire n10553;
	wire n10554;
	wire n10555;
	wire n10556;
	wire n10557;
	wire n10558;
	wire n10559;
	wire n10560;
	wire n10561;
	wire n10562;
	wire n10563;
	wire n10564;
	wire n10565;
	wire n10566;
	wire n10567;
	wire n10568;
	wire n10569;
	wire n10570;
	wire n10571;
	wire n10572;
	wire n10573;
	wire n10574;
	wire n10575;
	wire n10576;
	wire n10577;
	wire n10578;
	wire n10579;
	wire n10580;
	wire n10581;
	wire n10582;
	wire n10583;
	wire n10584;
	wire n10585;
	wire n10586;
	wire n10587;
	wire n10588;
	wire n10589;
	wire n10590;
	wire n10591;
	wire n10592;
	wire n10593;
	wire n10594;
	wire n10595;
	wire n10596;
	wire n10597;
	wire n10598;
	wire n10599;
	wire n10600;
	wire n10601;
	wire n10602;
	wire n10603;
	wire n10604;
	wire n10605;
	wire n10606;
	wire n10607;
	wire n10608;
	wire n10609;
	wire n10610;
	wire n10611;
	wire n10612;
	wire n10613;
	wire n10614;
	wire n10615;
	wire n10616;
	wire n10617;
	wire n10618;
	wire n10619;
	wire n10620;
	wire n10621;
	wire n10622;
	wire n10623;
	wire n10624;
	wire n10625;
	wire n10626;
	wire n10627;
	wire n10628;
	wire n10629;
	wire n10630;
	wire n10631;
	wire n10632;
	wire n10633;
	wire n10634;
	wire n10635;
	wire n10636;
	wire n10637;
	wire n10638;
	wire n10639;
	wire n10640;
	wire n10641;
	wire n10642;
	wire n10643;
	wire n10644;
	wire n10645;
	wire n10646;
	wire n10647;
	wire n10648;
	wire n10649;
	wire n10650;
	wire n10651;
	wire n10652;
	wire n10653;
	wire n10654;
	wire n10655;
	wire n10656;
	wire n10657;
	wire n10658;
	wire n10659;
	wire n10660;
	wire n10661;
	wire n10662;
	wire n10663;
	wire n10664;
	wire n10665;
	wire n10666;
	wire n10667;
	wire n10668;
	wire n10669;
	wire n10670;
	wire n10671;
	wire n10672;
	wire n10673;
	wire n10674;
	wire n10675;
	wire n10676;
	wire n10677;
	wire n10678;
	wire n10679;
	wire n10680;
	wire n10681;
	wire n10682;
	wire n10683;
	wire n10684;
	wire n10685;
	wire n10686;
	wire n10687;
	wire n10688;
	wire n10689;
	wire n10690;
	wire n10691;
	wire n10692;
	wire n10693;
	wire n10694;
	wire n10695;
	wire n10696;
	wire n10699;
	wire n10700;
	wire n10701;
	wire n10702;
	wire n10703;
	wire n10704;
	wire n10705;
	wire n10706;
	wire n10707;
	wire n10708;
	wire n10709;
	wire n10710;
	wire n10711;
	wire n10712;
	wire n10713;
	wire n10714;
	wire n10715;
	wire n10716;
	wire n10717;
	wire n10718;
	wire n10719;
	wire n10720;
	wire n10721;
	wire n10722;
	wire n10723;
	wire n10724;
	wire n10725;
	wire n10726;
	wire n10727;
	wire n10728;
	wire n10729;
	wire n10730;
	wire n10731;
	wire n10732;
	wire n10733;
	wire n10734;
	wire n10735;
	wire n10736;
	wire n10737;
	wire n10738;
	wire n10739;
	wire n10740;
	wire n10741;
	wire n10742;
	wire n10743;
	wire n10744;
	wire n10745;
	wire n10746;
	wire n10747;
	wire n10748;
	wire n10749;
	wire n10750;
	wire n10751;
	wire n10752;
	wire n10753;
	wire n10754;
	wire n10755;
	wire n10756;
	wire n10757;
	wire n10758;
	wire n10760;
	wire n10761;
	wire n10762;
	wire n10763;
	wire n10764;
	wire n10765;
	wire n10766;
	wire n10767;
	wire n10768;
	wire n10769;
	wire n10770;
	wire n10771;
	wire n10772;
	wire n10773;
	wire n10774;
	wire n10775;
	wire n10776;
	wire n10777;
	wire n10778;
	wire n10779;
	wire n10780;
	wire n10781;
	wire n10782;
	wire n10783;
	wire n10784;
	wire n10785;
	wire n10786;
	wire n10787;
	wire n10788;
	wire n10789;
	wire n10790;
	wire n10791;
	wire n10792;
	wire n10793;
	wire n10794;
	wire n10795;
	wire n10796;
	wire n10797;
	wire n10798;
	wire n10799;
	wire n10800;
	wire n10801;
	wire n10802;
	wire n10803;
	wire n10804;
	wire n10805;
	wire n10806;
	wire n10807;
	wire n10808;
	wire n10809;
	wire n10810;
	wire n10811;
	wire n10812;
	wire n10813;
	wire n10814;
	wire n10815;
	wire n10816;
	wire n10817;
	wire n10818;
	wire n10819;
	wire n10820;
	wire n10821;
	wire n10822;
	wire n10823;
	wire n10824;
	wire n10825;
	wire n10826;
	wire n10827;
	wire n10828;
	wire n10829;
	wire n10830;
	wire n10831;
	wire n10832;
	wire n10833;
	wire n10834;
	wire n10835;
	wire n10836;
	wire n10837;
	wire n10838;
	wire n10839;
	wire n10840;
	wire n10841;
	wire n10842;
	wire n10843;
	wire n10844;
	wire n10845;
	wire n10846;
	wire n10847;
	wire n10848;
	wire n10849;
	wire n10850;
	wire n10851;
	wire n10852;
	wire n10853;
	wire n10854;
	wire n10855;
	wire n10856;
	wire n10857;
	wire n10858;
	wire n10859;
	wire n10860;
	wire n10861;
	wire n10862;
	wire n10863;
	wire n10864;
	wire n10865;
	wire n10866;
	wire n10867;
	wire n10868;
	wire n10869;
	wire n10870;
	wire n10871;
	wire n10872;
	wire n10873;
	wire n10874;
	wire n10875;
	wire n10876;
	wire n10877;
	wire n10878;
	wire n10879;
	wire n10880;
	wire n10881;
	wire n10882;
	wire n10883;
	wire n10884;
	wire n10885;
	wire n10886;
	wire n10887;
	wire n10888;
	wire n10889;
	wire n10890;
	wire n10891;
	wire n10892;
	wire n10893;
	wire n10894;
	wire n10895;
	wire n10896;
	wire n10897;
	wire n10898;
	wire n10899;
	wire n10900;
	wire n10901;
	wire n10902;
	wire n10903;
	wire n10904;
	wire n10905;
	wire n10906;
	wire n10907;
	wire n10908;
	wire n10909;
	wire n10910;
	wire n10911;
	wire n10912;
	wire n10913;
	wire n10914;
	wire n10915;
	wire n10916;
	wire n10917;
	wire n10918;
	wire n10919;
	wire n10920;
	wire n10921;
	wire n10922;
	wire n10923;
	wire n10924;
	wire n10925;
	wire n10926;
	wire n10927;
	wire n10928;
	wire n10929;
	wire n10930;
	wire n10931;
	wire n10932;
	wire n10933;
	wire n10934;
	wire n10935;
	wire n10936;
	wire n10937;
	wire n10938;
	wire n10939;
	wire n10940;
	wire n10941;
	wire n10942;
	wire n10943;
	wire n10944;
	wire n10945;
	wire n10946;
	wire n10947;
	wire n10948;
	wire n10949;
	wire n10950;
	wire n10951;
	wire n10952;
	wire n10953;
	wire n10954;
	wire n10955;
	wire n10956;
	wire n10957;
	wire n10958;
	wire n10959;
	wire n10960;
	wire n10961;
	wire n10962;
	wire n10963;
	wire n10964;
	wire n10965;
	wire n10966;
	wire n10967;
	wire n10968;
	wire n10969;
	wire n10970;
	wire n10971;
	wire n10972;
	wire n10973;
	wire n10974;
	wire n10975;
	wire n10976;
	wire n10977;
	wire n10978;
	wire n10979;
	wire n10980;
	wire n10981;
	wire n10982;
	wire n10983;
	wire n10984;
	wire n10985;
	wire n10986;
	wire n10987;
	wire n10988;
	wire n10989;
	wire n10990;
	wire n10991;
	wire n10992;
	wire n10993;
	wire n10994;
	wire n10995;
	wire n10996;
	wire n10997;
	wire n10998;
	wire n10999;
	wire n11000;
	wire n11001;
	wire n11002;
	wire n11003;
	wire n11004;
	wire n11005;
	wire n11006;
	wire n11007;
	wire n11008;
	wire n11009;
	wire n11010;
	wire n11011;
	wire n11012;
	wire n11013;
	wire n11014;
	wire n11015;
	wire n11016;
	wire n11017;
	wire n11018;
	wire n11019;
	wire n11020;
	wire n11021;
	wire n11022;
	wire n11023;
	wire n11024;
	wire n11025;
	wire n11026;
	wire n11027;
	wire n11028;
	wire n11029;
	wire n11030;
	wire n11031;
	wire n11032;
	wire n11033;
	wire n11034;
	wire n11035;
	wire n11036;
	wire n11037;
	wire n11038;
	wire n11039;
	wire n11040;
	wire n11041;
	wire n11042;
	wire n11043;
	wire n11044;
	wire n11045;
	wire n11046;
	wire n11047;
	wire n11048;
	wire n11049;
	wire n11050;
	wire n11051;
	wire n11052;
	wire n11053;
	wire n11054;
	wire n11055;
	wire n11056;
	wire n11057;
	wire n11058;
	wire n11059;
	wire n11060;
	wire n11061;
	wire n11062;
	wire n11063;
	wire n11064;
	wire n11065;
	wire n11066;
	wire n11067;
	wire n11068;
	wire n11069;
	wire n11070;
	wire n11071;
	wire n11072;
	wire n11073;
	wire n11074;
	wire n11075;
	wire n11076;
	wire n11077;
	wire n11078;
	wire n11079;
	wire n11080;
	wire n11081;
	wire n11082;
	wire n11083;
	wire n11084;
	wire n11085;
	wire n11086;
	wire n11087;
	wire n11088;
	wire n11089;
	wire n11090;
	wire n11091;
	wire n11092;
	wire n11093;
	wire n11094;
	wire n11095;
	wire n11096;
	wire n11097;
	wire n11098;
	wire n11099;
	wire n11100;
	wire n11101;
	wire n11102;
	wire n11103;
	wire n11104;
	wire n11105;
	wire n11106;
	wire n11107;
	wire n11108;
	wire n11109;
	wire n11110;
	wire n11111;
	wire n11112;
	wire n11113;
	wire n11114;
	wire n11115;
	wire n11116;
	wire n11117;
	wire n11118;
	wire n11119;
	wire n11120;
	wire n11121;
	wire n11122;
	wire n11123;
	wire n11124;
	wire n11125;
	wire n11126;
	wire n11127;
	wire n11128;
	wire n11129;
	wire n11130;
	wire n11131;
	wire n11132;
	wire n11133;
	wire n11134;
	wire n11135;
	wire n11136;
	wire n11137;
	wire n11138;
	wire n11139;
	wire n11140;
	wire n11141;
	wire n11142;
	wire n11143;
	wire n11144;
	wire n11145;
	wire n11146;
	wire n11147;
	wire n11148;
	wire n11149;
	wire n11150;
	wire n11151;
	wire n11154;
	wire n11156;
	wire n11157;
	wire n11158;
	wire n11159;
	wire n11160;
	wire n11161;
	wire n11162;
	wire n11163;
	wire n11164;
	wire n11165;
	wire n11166;
	wire n11167;
	wire n11168;
	wire n11169;
	wire n11170;
	wire n11171;
	wire n11172;
	wire n11173;
	wire n11174;
	wire n11175;
	wire n11176;
	wire n11177;
	wire n11178;
	wire n11179;
	wire n11180;
	wire n11181;
	wire n11182;
	wire n11183;
	wire n11184;
	wire n11185;
	wire n11186;
	wire n11187;
	wire n11188;
	wire n11189;
	wire n11190;
	wire n11191;
	wire n11192;
	wire n11193;
	wire n11194;
	wire n11195;
	wire n11196;
	wire n11197;
	wire n11198;
	wire n11199;
	wire n11200;
	wire n11201;
	wire n11202;
	wire n11203;
	wire n11204;
	wire n11205;
	wire n11206;
	wire n11207;
	wire n11208;
	wire n11209;
	wire n11210;
	wire n11211;
	wire n11212;
	wire n11213;
	wire n11214;
	wire n11215;
	wire n11216;
	wire n11217;
	wire n11218;
	wire n11219;
	wire n11220;
	wire n11221;
	wire n11222;
	wire n11223;
	wire n11224;
	wire n11225;
	wire n11226;
	wire n11227;
	wire n11228;
	wire n11229;
	wire n11230;
	wire n11231;
	wire n11232;
	wire n11233;
	wire n11234;
	wire n11235;
	wire n11236;
	wire n11237;
	wire n11238;
	wire n11239;
	wire n11240;
	wire n11241;
	wire n11242;
	wire n11243;
	wire n11244;
	wire n11245;
	wire n11246;
	wire n11247;
	wire n11248;
	wire n11249;
	wire n11250;
	wire n11251;
	wire n11252;
	wire n11253;
	wire n11254;
	wire n11255;
	wire n11256;
	wire n11257;
	wire n11258;
	wire n11259;
	wire n11260;
	wire n11261;
	wire n11262;
	wire n11263;
	wire n11264;
	wire n11265;
	wire n11266;
	wire n11267;
	wire n11268;
	wire n11269;
	wire n11270;
	wire n11271;
	wire n11272;
	wire n11273;
	wire n11274;
	wire n11275;
	wire n11276;
	wire n11277;
	wire n11278;
	wire n11279;
	wire n11280;
	wire n11281;
	wire n11282;
	wire n11283;
	wire n11284;
	wire n11285;
	wire n11286;
	wire n11287;
	wire n11288;
	wire n11289;
	wire n11290;
	wire n11291;
	wire n11292;
	wire n11293;
	wire n11294;
	wire n11295;
	wire n11296;
	wire n11297;
	wire n11298;
	wire n11299;
	wire n11300;
	wire n11301;
	wire n11302;
	wire n11303;
	wire n11304;
	wire n11305;
	wire n11306;
	wire n11307;
	wire n11308;
	wire n11309;
	wire n11310;
	wire n11311;
	wire n11312;
	wire n11313;
	wire n11314;
	wire n11315;
	wire n11316;
	wire n11317;
	wire n11318;
	wire n11319;
	wire n11320;
	wire n11321;
	wire n11322;
	wire n11323;
	wire n11324;
	wire n11325;
	wire n11326;
	wire n11327;
	wire n11328;
	wire n11329;
	wire n11330;
	wire n11331;
	wire n11332;
	wire n11333;
	wire n11334;
	wire n11335;
	wire n11336;
	wire n11337;
	wire n11338;
	wire n11339;
	wire n11340;
	wire n11341;
	wire n11342;
	wire n11343;
	wire n11344;
	wire n11345;
	wire n11346;
	wire n11347;
	wire n11348;
	wire n11349;
	wire n11350;
	wire n11351;
	wire n11352;
	wire n11353;
	wire n11354;
	wire n11355;
	wire n11356;
	wire n11357;
	wire n11358;
	wire n11359;
	wire n11360;
	wire n11361;
	wire n11362;
	wire n11363;
	wire n11364;
	wire n11365;
	wire n11366;
	wire n11367;
	wire n11368;
	wire n11369;
	wire n11370;
	wire n11371;
	wire n11372;
	wire n11373;
	wire n11374;
	wire n11375;
	wire n11376;
	wire n11377;
	wire n11378;
	wire n11379;
	wire n11380;
	wire n11381;
	wire n11382;
	wire n11383;
	wire n11384;
	wire n11385;
	wire n11386;
	wire n11387;
	wire n11388;
	wire n11389;
	wire n11390;
	wire n11391;
	wire n11392;
	wire n11393;
	wire n11394;
	wire n11395;
	wire n11396;
	wire n11397;
	wire n11398;
	wire n11399;
	wire n11400;
	wire n11401;
	wire n11402;
	wire n11403;
	wire n11404;
	wire n11405;
	wire n11406;
	wire n11407;
	wire n11408;
	wire n11409;
	wire n11410;
	wire n11411;
	wire n11412;
	wire n11413;
	wire n11414;
	wire n11415;
	wire n11416;
	wire n11417;
	wire n11418;
	wire n11419;
	wire n11420;
	wire n11421;
	wire n11422;
	wire n11423;
	wire n11424;
	wire n11425;
	wire n11426;
	wire n11427;
	wire n11428;
	wire n11429;
	wire n11430;
	wire n11431;
	wire n11432;
	wire n11433;
	wire n11434;
	wire n11435;
	wire n11436;
	wire n11437;
	wire n11438;
	wire n11439;
	wire n11440;
	wire n11441;
	wire n11442;
	wire n11443;
	wire n11444;
	wire n11445;
	wire n11446;
	wire n11447;
	wire n11448;
	wire n11449;
	wire n11450;
	wire n11451;
	wire n11452;
	wire n11453;
	wire n11454;
	wire n11455;
	wire n11456;
	wire n11457;
	wire n11458;
	wire n11459;
	wire n11460;
	wire n11461;
	wire n11462;
	wire n11463;
	wire n11464;
	wire n11465;
	wire n11466;
	wire n11467;
	wire n11468;
	wire n11469;
	wire n11470;
	wire n11471;
	wire n11472;
	wire n11473;
	wire n11474;
	wire n11475;
	wire n11476;
	wire n11477;
	wire n11478;
	wire n11479;
	wire n11480;
	wire n11481;
	wire n11482;
	wire n11483;
	wire n11484;
	wire n11485;
	wire n11486;
	wire n11487;
	wire n11488;
	wire n11489;
	wire n11490;
	wire n11491;
	wire n11492;
	wire n11493;
	wire n11494;
	wire n11495;
	wire n11496;
	wire n11497;
	wire n11498;
	wire n11499;
	wire n11500;
	wire n11501;
	wire n11502;
	wire n11503;
	wire n11504;
	wire n11505;
	wire n11506;
	wire n11507;
	wire n11508;
	wire n11509;
	wire n11510;
	wire n11511;
	wire n11512;
	wire n11513;
	wire n11514;
	wire n11515;
	wire n11516;
	wire n11517;
	wire n11518;
	wire n11519;
	wire n11520;
	wire n11521;
	wire n11522;
	wire n11523;
	wire n11524;
	wire n11525;
	wire n11526;
	wire n11527;
	wire n11528;
	wire n11529;
	wire n11530;
	wire n11531;
	wire n11532;
	wire n11533;
	wire n11534;
	wire n11535;
	wire n11536;
	wire n11537;
	wire n11538;
	wire n11539;
	wire n11540;
	wire n11541;
	wire n11542;
	wire n11543;
	wire n11544;
	wire n11545;
	wire n11546;
	wire n11547;
	wire n11548;
	wire n11549;
	wire n11550;
	wire n11551;
	wire n11552;
	wire n11553;
	wire n11554;
	wire n11555;
	wire n11556;
	wire n11557;
	wire n11558;
	wire n11559;
	wire n11560;
	wire n11561;
	wire n11562;
	wire n11563;
	wire n11564;
	wire n11565;
	wire n11566;
	wire n11567;
	wire n11568;
	wire n11569;
	wire n11570;
	wire n11571;
	wire n11572;
	wire n11573;
	wire n11574;
	wire n11575;
	wire n11576;
	wire n11577;
	wire n11578;
	wire n11579;
	wire n11580;
	wire n11581;
	wire n11582;
	wire n11583;
	wire n11584;
	wire n11585;
	wire n11586;
	wire n11587;
	wire n11588;
	wire n11589;
	wire n11590;
	wire n11591;
	wire n11592;
	wire n11593;
	wire n11594;
	wire n11595;
	wire n11596;
	wire n11597;
	wire n11598;
	wire n11599;
	wire n11600;
	wire n11601;
	wire n11602;
	wire n11603;
	wire n11604;
	wire n11605;
	wire n11606;
	wire n11607;
	wire n11608;
	wire n11609;
	wire n11610;
	wire n11611;
	wire n11612;
	wire n11613;
	wire n11614;
	wire n11615;
	wire n11616;
	wire n11617;
	wire n11618;
	wire n11619;
	wire n11620;
	wire n11621;
	wire n11622;
	wire n11623;
	wire n11624;
	wire n11625;
	wire n11626;
	wire n11627;
	wire n11628;
	wire n11629;
	wire n11630;
	wire n11631;
	wire n11632;
	wire n11633;
	wire n11634;
	wire n11635;
	wire n11636;
	wire n11637;
	wire n11638;
	wire n11639;
	wire n11640;
	wire n11641;
	wire n11642;
	wire n11643;
	wire n11644;
	wire n11645;
	wire n11646;
	wire n11647;
	wire n11648;
	wire n11649;
	wire n11650;
	wire n11651;
	wire n11652;
	wire n11653;
	wire n11654;
	wire n11655;
	wire n11656;
	wire n11657;
	wire n11660;
	wire n11661;
	wire n11662;
	wire n11663;
	wire n11664;
	wire n11665;
	wire n11666;
	wire n11667;
	wire n11668;
	wire n11669;
	wire n11670;
	wire n11671;
	wire n11672;
	wire n11673;
	wire n11674;
	wire n11675;
	wire n11676;
	wire n11677;
	wire n11678;
	wire n11679;
	wire n11680;
	wire n11681;
	wire n11682;
	wire n11683;
	wire n11684;
	wire n11685;
	wire n11686;
	wire n11687;
	wire n11688;
	wire n11689;
	wire n11690;
	wire n11691;
	wire n11692;
	wire n11693;
	wire n11694;
	wire n11695;
	wire n11696;
	wire n11697;
	wire n11698;
	wire n11699;
	wire n11700;
	wire n11701;
	wire n11702;
	wire n11703;
	wire n11704;
	wire n11705;
	wire n11706;
	wire n11707;
	wire n11708;
	wire n11709;
	wire n11710;
	wire n11711;
	wire n11712;
	wire n11713;
	wire n11714;
	wire n11715;
	wire n11716;
	wire n11717;
	wire n11718;
	wire n11719;
	wire n11721;
	wire n11722;
	wire n11723;
	wire n11724;
	wire n11725;
	wire n11726;
	wire n11727;
	wire n11728;
	wire n11729;
	wire n11730;
	wire n11731;
	wire n11732;
	wire n11733;
	wire n11734;
	wire n11735;
	wire n11736;
	wire n11737;
	wire n11738;
	wire n11739;
	wire n11740;
	wire n11741;
	wire n11742;
	wire n11743;
	wire n11744;
	wire n11745;
	wire n11746;
	wire n11747;
	wire n11748;
	wire n11749;
	wire n11750;
	wire n11751;
	wire n11752;
	wire n11753;
	wire n11754;
	wire n11755;
	wire n11756;
	wire n11757;
	wire n11758;
	wire n11759;
	wire n11760;
	wire n11761;
	wire n11762;
	wire n11763;
	wire n11764;
	wire n11765;
	wire n11766;
	wire n11767;
	wire n11768;
	wire n11769;
	wire n11770;
	wire n11771;
	wire n11772;
	wire n11773;
	wire n11774;
	wire n11775;
	wire n11776;
	wire n11777;
	wire n11778;
	wire n11779;
	wire n11780;
	wire n11781;
	wire n11782;
	wire n11783;
	wire n11784;
	wire n11785;
	wire n11786;
	wire n11787;
	wire n11788;
	wire n11789;
	wire n11790;
	wire n11791;
	wire n11792;
	wire n11793;
	wire n11794;
	wire n11795;
	wire n11796;
	wire n11797;
	wire n11798;
	wire n11799;
	wire n11800;
	wire n11801;
	wire n11802;
	wire n11803;
	wire n11804;
	wire n11805;
	wire n11806;
	wire n11807;
	wire n11808;
	wire n11809;
	wire n11810;
	wire n11811;
	wire n11812;
	wire n11813;
	wire n11814;
	wire n11815;
	wire n11816;
	wire n11817;
	wire n11818;
	wire n11819;
	wire n11820;
	wire n11821;
	wire n11822;
	wire n11823;
	wire n11824;
	wire n11825;
	wire n11826;
	wire n11827;
	wire n11828;
	wire n11829;
	wire n11830;
	wire n11831;
	wire n11832;
	wire n11833;
	wire n11834;
	wire n11835;
	wire n11836;
	wire n11837;
	wire n11838;
	wire n11839;
	wire n11840;
	wire n11841;
	wire n11842;
	wire n11843;
	wire n11844;
	wire n11845;
	wire n11846;
	wire n11847;
	wire n11848;
	wire n11849;
	wire n11850;
	wire n11851;
	wire n11852;
	wire n11853;
	wire n11854;
	wire n11855;
	wire n11856;
	wire n11857;
	wire n11858;
	wire n11859;
	wire n11860;
	wire n11861;
	wire n11862;
	wire n11863;
	wire n11864;
	wire n11865;
	wire n11866;
	wire n11867;
	wire n11868;
	wire n11869;
	wire n11870;
	wire n11871;
	wire n11872;
	wire n11873;
	wire n11874;
	wire n11875;
	wire n11876;
	wire n11877;
	wire n11878;
	wire n11879;
	wire n11880;
	wire n11881;
	wire n11882;
	wire n11883;
	wire n11884;
	wire n11885;
	wire n11886;
	wire n11887;
	wire n11888;
	wire n11889;
	wire n11890;
	wire n11891;
	wire n11892;
	wire n11893;
	wire n11894;
	wire n11895;
	wire n11896;
	wire n11897;
	wire n11898;
	wire n11899;
	wire n11900;
	wire n11901;
	wire n11902;
	wire n11903;
	wire n11904;
	wire n11905;
	wire n11906;
	wire n11907;
	wire n11908;
	wire n11909;
	wire n11910;
	wire n11911;
	wire n11912;
	wire n11913;
	wire n11914;
	wire n11915;
	wire n11916;
	wire n11917;
	wire n11918;
	wire n11919;
	wire n11920;
	wire n11921;
	wire n11922;
	wire n11923;
	wire n11924;
	wire n11925;
	wire n11926;
	wire n11927;
	wire n11928;
	wire n11929;
	wire n11930;
	wire n11931;
	wire n11932;
	wire n11933;
	wire n11934;
	wire n11935;
	wire n11936;
	wire n11937;
	wire n11938;
	wire n11939;
	wire n11940;
	wire n11941;
	wire n11942;
	wire n11943;
	wire n11944;
	wire n11945;
	wire n11946;
	wire n11947;
	wire n11948;
	wire n11949;
	wire n11950;
	wire n11951;
	wire n11952;
	wire n11953;
	wire n11954;
	wire n11955;
	wire n11956;
	wire n11957;
	wire n11958;
	wire n11959;
	wire n11960;
	wire n11961;
	wire n11962;
	wire n11963;
	wire n11964;
	wire n11965;
	wire n11966;
	wire n11967;
	wire n11968;
	wire n11969;
	wire n11970;
	wire n11971;
	wire n11972;
	wire n11973;
	wire n11974;
	wire n11975;
	wire n11976;
	wire n11977;
	wire n11978;
	wire n11979;
	wire n11980;
	wire n11981;
	wire n11982;
	wire n11983;
	wire n11984;
	wire n11985;
	wire n11986;
	wire n11987;
	wire n11988;
	wire n11989;
	wire n11990;
	wire n11991;
	wire n11992;
	wire n11993;
	wire n11994;
	wire n11995;
	wire n11996;
	wire n11997;
	wire n11998;
	wire n11999;
	wire n12000;
	wire n12001;
	wire n12002;
	wire n12003;
	wire n12004;
	wire n12005;
	wire n12006;
	wire n12007;
	wire n12008;
	wire n12009;
	wire n12010;
	wire n12011;
	wire n12012;
	wire n12013;
	wire n12014;
	wire n12015;
	wire n12016;
	wire n12017;
	wire n12018;
	wire n12019;
	wire n12020;
	wire n12021;
	wire n12022;
	wire n12023;
	wire n12024;
	wire n12025;
	wire n12026;
	wire n12027;
	wire n12028;
	wire n12029;
	wire n12030;
	wire n12031;
	wire n12032;
	wire n12033;
	wire n12034;
	wire n12035;
	wire n12036;
	wire n12037;
	wire n12038;
	wire n12039;
	wire n12040;
	wire n12041;
	wire n12042;
	wire n12043;
	wire n12044;
	wire n12045;
	wire n12046;
	wire n12047;
	wire n12048;
	wire n12049;
	wire n12050;
	wire n12051;
	wire n12052;
	wire n12053;
	wire n12054;
	wire n12055;
	wire n12056;
	wire n12057;
	wire n12058;
	wire n12059;
	wire n12060;
	wire n12061;
	wire n12062;
	wire n12063;
	wire n12064;
	wire n12065;
	wire n12066;
	wire n12067;
	wire n12068;
	wire n12069;
	wire n12070;
	wire n12071;
	wire n12072;
	wire n12073;
	wire n12074;
	wire n12075;
	wire n12076;
	wire n12077;
	wire n12078;
	wire n12079;
	wire n12080;
	wire n12081;
	wire n12082;
	wire n12083;
	wire n12084;
	wire n12085;
	wire n12086;
	wire n12087;
	wire n12088;
	wire n12089;
	wire n12090;
	wire n12091;
	wire n12092;
	wire n12093;
	wire n12094;
	wire n12095;
	wire n12096;
	wire n12097;
	wire n12098;
	wire n12099;
	wire n12100;
	wire n12101;
	wire n12102;
	wire n12103;
	wire n12104;
	wire n12105;
	wire n12106;
	wire n12107;
	wire n12108;
	wire n12109;
	wire n12110;
	wire n12111;
	wire n12112;
	wire n12113;
	wire n12114;
	wire n12115;
	wire n12116;
	wire n12117;
	wire n12118;
	wire n12119;
	wire n12120;
	wire n12121;
	wire n12122;
	wire n12123;
	wire n12124;
	wire n12125;
	wire n12126;
	wire n12127;
	wire n12128;
	wire n12129;
	wire n12130;
	wire n12131;
	wire n12132;
	wire n12133;
	wire n12134;
	wire n12135;
	wire n12136;
	wire n12137;
	wire n12138;
	wire n12141;
	wire n12143;
	wire n12144;
	wire n12145;
	wire n12146;
	wire n12147;
	wire n12148;
	wire n12149;
	wire n12150;
	wire n12151;
	wire n12152;
	wire n12153;
	wire n12154;
	wire n12155;
	wire n12156;
	wire n12157;
	wire n12158;
	wire n12159;
	wire n12160;
	wire n12161;
	wire n12162;
	wire n12163;
	wire n12164;
	wire n12165;
	wire n12166;
	wire n12167;
	wire n12168;
	wire n12169;
	wire n12170;
	wire n12171;
	wire n12172;
	wire n12173;
	wire n12174;
	wire n12175;
	wire n12176;
	wire n12177;
	wire n12178;
	wire n12179;
	wire n12180;
	wire n12181;
	wire n12182;
	wire n12183;
	wire n12184;
	wire n12185;
	wire n12186;
	wire n12187;
	wire n12188;
	wire n12189;
	wire n12190;
	wire n12191;
	wire n12192;
	wire n12193;
	wire n12194;
	wire n12195;
	wire n12196;
	wire n12197;
	wire n12198;
	wire n12199;
	wire n12200;
	wire n12201;
	wire n12202;
	wire n12203;
	wire n12204;
	wire n12205;
	wire n12206;
	wire n12207;
	wire n12208;
	wire n12209;
	wire n12210;
	wire n12211;
	wire n12212;
	wire n12213;
	wire n12214;
	wire n12215;
	wire n12216;
	wire n12217;
	wire n12218;
	wire n12219;
	wire n12220;
	wire n12221;
	wire n12222;
	wire n12223;
	wire n12224;
	wire n12225;
	wire n12226;
	wire n12227;
	wire n12228;
	wire n12229;
	wire n12230;
	wire n12231;
	wire n12232;
	wire n12233;
	wire n12234;
	wire n12235;
	wire n12236;
	wire n12237;
	wire n12238;
	wire n12239;
	wire n12240;
	wire n12241;
	wire n12242;
	wire n12243;
	wire n12244;
	wire n12245;
	wire n12246;
	wire n12247;
	wire n12248;
	wire n12249;
	wire n12250;
	wire n12251;
	wire n12252;
	wire n12253;
	wire n12254;
	wire n12255;
	wire n12256;
	wire n12257;
	wire n12258;
	wire n12259;
	wire n12260;
	wire n12261;
	wire n12262;
	wire n12263;
	wire n12264;
	wire n12265;
	wire n12266;
	wire n12267;
	wire n12268;
	wire n12269;
	wire n12270;
	wire n12271;
	wire n12272;
	wire n12273;
	wire n12274;
	wire n12275;
	wire n12276;
	wire n12277;
	wire n12278;
	wire n12279;
	wire n12280;
	wire n12281;
	wire n12282;
	wire n12283;
	wire n12284;
	wire n12285;
	wire n12286;
	wire n12287;
	wire n12288;
	wire n12289;
	wire n12290;
	wire n12291;
	wire n12292;
	wire n12293;
	wire n12294;
	wire n12295;
	wire n12296;
	wire n12297;
	wire n12298;
	wire n12299;
	wire n12300;
	wire n12301;
	wire n12302;
	wire n12303;
	wire n12304;
	wire n12305;
	wire n12306;
	wire n12307;
	wire n12308;
	wire n12309;
	wire n12310;
	wire n12311;
	wire n12312;
	wire n12313;
	wire n12314;
	wire n12315;
	wire n12316;
	wire n12317;
	wire n12318;
	wire n12319;
	wire n12320;
	wire n12321;
	wire n12322;
	wire n12323;
	wire n12324;
	wire n12325;
	wire n12326;
	wire n12327;
	wire n12328;
	wire n12329;
	wire n12330;
	wire n12331;
	wire n12332;
	wire n12333;
	wire n12334;
	wire n12335;
	wire n12336;
	wire n12337;
	wire n12338;
	wire n12339;
	wire n12340;
	wire n12341;
	wire n12342;
	wire n12343;
	wire n12344;
	wire n12345;
	wire n12346;
	wire n12347;
	wire n12348;
	wire n12349;
	wire n12350;
	wire n12351;
	wire n12352;
	wire n12353;
	wire n12354;
	wire n12355;
	wire n12356;
	wire n12357;
	wire n12358;
	wire n12359;
	wire n12360;
	wire n12361;
	wire n12362;
	wire n12363;
	wire n12364;
	wire n12365;
	wire n12366;
	wire n12367;
	wire n12368;
	wire n12369;
	wire n12370;
	wire n12371;
	wire n12372;
	wire n12373;
	wire n12374;
	wire n12375;
	wire n12376;
	wire n12377;
	wire n12378;
	wire n12379;
	wire n12380;
	wire n12381;
	wire n12382;
	wire n12383;
	wire n12384;
	wire n12385;
	wire n12386;
	wire n12387;
	wire n12388;
	wire n12389;
	wire n12390;
	wire n12391;
	wire n12392;
	wire n12393;
	wire n12394;
	wire n12395;
	wire n12396;
	wire n12397;
	wire n12398;
	wire n12399;
	wire n12400;
	wire n12401;
	wire n12402;
	wire n12403;
	wire n12404;
	wire n12405;
	wire n12406;
	wire n12407;
	wire n12408;
	wire n12409;
	wire n12410;
	wire n12411;
	wire n12412;
	wire n12413;
	wire n12414;
	wire n12415;
	wire n12416;
	wire n12417;
	wire n12418;
	wire n12419;
	wire n12420;
	wire n12421;
	wire n12422;
	wire n12423;
	wire n12424;
	wire n12425;
	wire n12426;
	wire n12427;
	wire n12428;
	wire n12429;
	wire n12430;
	wire n12431;
	wire n12432;
	wire n12433;
	wire n12434;
	wire n12435;
	wire n12436;
	wire n12437;
	wire n12438;
	wire n12439;
	wire n12440;
	wire n12441;
	wire n12442;
	wire n12443;
	wire n12444;
	wire n12445;
	wire n12446;
	wire n12447;
	wire n12448;
	wire n12449;
	wire n12450;
	wire n12451;
	wire n12452;
	wire n12453;
	wire n12454;
	wire n12455;
	wire n12456;
	wire n12457;
	wire n12458;
	wire n12459;
	wire n12460;
	wire n12461;
	wire n12462;
	wire n12463;
	wire n12464;
	wire n12465;
	wire n12466;
	wire n12467;
	wire n12468;
	wire n12469;
	wire n12470;
	wire n12471;
	wire n12472;
	wire n12473;
	wire n12474;
	wire n12475;
	wire n12476;
	wire n12477;
	wire n12478;
	wire n12479;
	wire n12480;
	wire n12481;
	wire n12482;
	wire n12483;
	wire n12484;
	wire n12485;
	wire n12486;
	wire n12487;
	wire n12488;
	wire n12489;
	wire n12490;
	wire n12491;
	wire n12492;
	wire n12493;
	wire n12494;
	wire n12495;
	wire n12496;
	wire n12497;
	wire n12498;
	wire n12499;
	wire n12500;
	wire n12501;
	wire n12502;
	wire n12503;
	wire n12504;
	wire n12505;
	wire n12506;
	wire n12507;
	wire n12508;
	wire n12509;
	wire n12510;
	wire n12511;
	wire n12512;
	wire n12513;
	wire n12514;
	wire n12515;
	wire n12516;
	wire n12517;
	wire n12518;
	wire n12519;
	wire n12520;
	wire n12521;
	wire n12522;
	wire n12523;
	wire n12524;
	wire n12525;
	wire n12526;
	wire n12527;
	wire n12528;
	wire n12529;
	wire n12530;
	wire n12531;
	wire n12532;
	wire n12533;
	wire n12534;
	wire n12535;
	wire n12536;
	wire n12537;
	wire n12538;
	wire n12539;
	wire n12540;
	wire n12541;
	wire n12542;
	wire n12543;
	wire n12544;
	wire n12545;
	wire n12546;
	wire n12547;
	wire n12548;
	wire n12549;
	wire n12550;
	wire n12551;
	wire n12552;
	wire n12553;
	wire n12554;
	wire n12555;
	wire n12556;
	wire n12557;
	wire n12558;
	wire n12559;
	wire n12560;
	wire n12561;
	wire n12562;
	wire n12563;
	wire n12564;
	wire n12565;
	wire n12566;
	wire n12567;
	wire n12568;
	wire n12569;
	wire n12570;
	wire n12571;
	wire n12572;
	wire n12573;
	wire n12574;
	wire n12575;
	wire n12576;
	wire n12577;
	wire n12578;
	wire n12579;
	wire n12580;
	wire n12581;
	wire n12582;
	wire n12583;
	wire n12584;
	wire n12585;
	wire n12586;
	wire n12587;
	wire n12588;
	wire n12589;
	wire n12590;
	wire n12591;
	wire n12592;
	wire n12593;
	wire n12594;
	wire n12595;
	wire n12596;
	wire n12597;
	wire n12598;
	wire n12599;
	wire n12600;
	wire n12601;
	wire n12602;
	wire n12603;
	wire n12604;
	wire n12605;
	wire n12606;
	wire n12607;
	wire n12608;
	wire n12609;
	wire n12610;
	wire n12611;
	wire n12612;
	wire n12613;
	wire n12614;
	wire n12615;
	wire n12616;
	wire n12617;
	wire n12618;
	wire n12619;
	wire n12620;
	wire n12621;
	wire n12622;
	wire n12623;
	wire n12624;
	wire n12625;
	wire n12626;
	wire n12627;
	wire n12628;
	wire n12629;
	wire n12630;
	wire n12631;
	wire n12632;
	wire n12633;
	wire n12634;
	wire n12635;
	wire n12636;
	wire n12637;
	wire n12638;
	wire n12639;
	wire n12640;
	wire n12641;
	wire n12642;
	wire n12643;
	wire n12644;
	wire n12645;
	wire n12646;
	wire n12647;
	wire n12648;
	wire n12649;
	wire n12650;
	wire n12651;
	wire n12652;
	wire n12653;
	wire n12654;
	wire n12655;
	wire n12656;
	wire n12657;
	wire n12658;
	wire n12659;
	wire n12660;
	wire n12661;
	wire n12662;
	wire n12663;
	wire n12664;
	wire n12665;
	wire n12666;
	wire n12667;
	wire n12668;
	wire n12669;
	wire n12670;
	wire n12673;
	wire n12674;
	wire n12675;
	wire n12676;
	wire n12677;
	wire n12678;
	wire n12679;
	wire n12680;
	wire n12681;
	wire n12682;
	wire n12683;
	wire n12684;
	wire n12685;
	wire n12686;
	wire n12687;
	wire n12688;
	wire n12689;
	wire n12690;
	wire n12691;
	wire n12692;
	wire n12693;
	wire n12694;
	wire n12695;
	wire n12696;
	wire n12697;
	wire n12698;
	wire n12699;
	wire n12700;
	wire n12701;
	wire n12702;
	wire n12703;
	wire n12704;
	wire n12705;
	wire n12706;
	wire n12707;
	wire n12708;
	wire n12709;
	wire n12710;
	wire n12711;
	wire n12712;
	wire n12713;
	wire n12714;
	wire n12715;
	wire n12716;
	wire n12717;
	wire n12718;
	wire n12719;
	wire n12720;
	wire n12721;
	wire n12722;
	wire n12723;
	wire n12724;
	wire n12725;
	wire n12726;
	wire n12727;
	wire n12728;
	wire n12729;
	wire n12730;
	wire n12731;
	wire n12732;
	wire n12733;
	wire n12735;
	wire n12736;
	wire n12737;
	wire n12738;
	wire n12739;
	wire n12740;
	wire n12741;
	wire n12742;
	wire n12743;
	wire n12744;
	wire n12745;
	wire n12746;
	wire n12747;
	wire n12748;
	wire n12749;
	wire n12750;
	wire n12751;
	wire n12752;
	wire n12753;
	wire n12754;
	wire n12755;
	wire n12756;
	wire n12757;
	wire n12758;
	wire n12759;
	wire n12760;
	wire n12761;
	wire n12762;
	wire n12763;
	wire n12764;
	wire n12765;
	wire n12766;
	wire n12767;
	wire n12768;
	wire n12769;
	wire n12770;
	wire n12771;
	wire n12772;
	wire n12773;
	wire n12774;
	wire n12775;
	wire n12776;
	wire n12777;
	wire n12778;
	wire n12779;
	wire n12780;
	wire n12781;
	wire n12782;
	wire n12783;
	wire n12784;
	wire n12785;
	wire n12786;
	wire n12787;
	wire n12788;
	wire n12789;
	wire n12790;
	wire n12791;
	wire n12792;
	wire n12793;
	wire n12794;
	wire n12795;
	wire n12796;
	wire n12797;
	wire n12798;
	wire n12799;
	wire n12800;
	wire n12801;
	wire n12802;
	wire n12803;
	wire n12804;
	wire n12805;
	wire n12806;
	wire n12807;
	wire n12808;
	wire n12809;
	wire n12810;
	wire n12811;
	wire n12812;
	wire n12813;
	wire n12814;
	wire n12815;
	wire n12816;
	wire n12817;
	wire n12818;
	wire n12819;
	wire n12820;
	wire n12821;
	wire n12822;
	wire n12823;
	wire n12824;
	wire n12825;
	wire n12826;
	wire n12827;
	wire n12828;
	wire n12829;
	wire n12830;
	wire n12831;
	wire n12832;
	wire n12833;
	wire n12834;
	wire n12835;
	wire n12836;
	wire n12837;
	wire n12838;
	wire n12839;
	wire n12840;
	wire n12841;
	wire n12842;
	wire n12843;
	wire n12844;
	wire n12845;
	wire n12846;
	wire n12847;
	wire n12848;
	wire n12849;
	wire n12850;
	wire n12851;
	wire n12852;
	wire n12853;
	wire n12854;
	wire n12855;
	wire n12856;
	wire n12857;
	wire n12858;
	wire n12859;
	wire n12860;
	wire n12861;
	wire n12862;
	wire n12863;
	wire n12864;
	wire n12865;
	wire n12866;
	wire n12867;
	wire n12868;
	wire n12869;
	wire n12870;
	wire n12871;
	wire n12872;
	wire n12873;
	wire n12874;
	wire n12875;
	wire n12876;
	wire n12877;
	wire n12878;
	wire n12879;
	wire n12880;
	wire n12881;
	wire n12882;
	wire n12883;
	wire n12884;
	wire n12885;
	wire n12886;
	wire n12887;
	wire n12888;
	wire n12889;
	wire n12890;
	wire n12891;
	wire n12892;
	wire n12893;
	wire n12894;
	wire n12895;
	wire n12896;
	wire n12897;
	wire n12898;
	wire n12899;
	wire n12900;
	wire n12901;
	wire n12902;
	wire n12903;
	wire n12904;
	wire n12905;
	wire n12906;
	wire n12907;
	wire n12908;
	wire n12909;
	wire n12910;
	wire n12911;
	wire n12912;
	wire n12913;
	wire n12914;
	wire n12915;
	wire n12916;
	wire n12917;
	wire n12918;
	wire n12919;
	wire n12920;
	wire n12921;
	wire n12922;
	wire n12923;
	wire n12924;
	wire n12925;
	wire n12926;
	wire n12927;
	wire n12928;
	wire n12929;
	wire n12930;
	wire n12931;
	wire n12932;
	wire n12933;
	wire n12934;
	wire n12935;
	wire n12936;
	wire n12937;
	wire n12938;
	wire n12939;
	wire n12940;
	wire n12941;
	wire n12942;
	wire n12943;
	wire n12944;
	wire n12945;
	wire n12946;
	wire n12947;
	wire n12948;
	wire n12949;
	wire n12950;
	wire n12951;
	wire n12952;
	wire n12953;
	wire n12954;
	wire n12955;
	wire n12956;
	wire n12957;
	wire n12958;
	wire n12959;
	wire n12960;
	wire n12961;
	wire n12962;
	wire n12963;
	wire n12964;
	wire n12965;
	wire n12966;
	wire n12967;
	wire n12968;
	wire n12969;
	wire n12970;
	wire n12971;
	wire n12972;
	wire n12973;
	wire n12974;
	wire n12975;
	wire n12976;
	wire n12977;
	wire n12978;
	wire n12979;
	wire n12980;
	wire n12981;
	wire n12982;
	wire n12983;
	wire n12984;
	wire n12985;
	wire n12986;
	wire n12987;
	wire n12988;
	wire n12989;
	wire n12990;
	wire n12991;
	wire n12992;
	wire n12993;
	wire n12994;
	wire n12995;
	wire n12996;
	wire n12997;
	wire n12998;
	wire n12999;
	wire n13000;
	wire n13001;
	wire n13002;
	wire n13003;
	wire n13004;
	wire n13005;
	wire n13006;
	wire n13007;
	wire n13008;
	wire n13009;
	wire n13010;
	wire n13011;
	wire n13012;
	wire n13013;
	wire n13014;
	wire n13015;
	wire n13016;
	wire n13017;
	wire n13018;
	wire n13019;
	wire n13020;
	wire n13021;
	wire n13022;
	wire n13023;
	wire n13024;
	wire n13025;
	wire n13026;
	wire n13027;
	wire n13028;
	wire n13029;
	wire n13030;
	wire n13031;
	wire n13032;
	wire n13033;
	wire n13034;
	wire n13035;
	wire n13036;
	wire n13037;
	wire n13038;
	wire n13039;
	wire n13040;
	wire n13041;
	wire n13042;
	wire n13043;
	wire n13044;
	wire n13045;
	wire n13046;
	wire n13047;
	wire n13048;
	wire n13049;
	wire n13050;
	wire n13051;
	wire n13052;
	wire n13053;
	wire n13054;
	wire n13055;
	wire n13056;
	wire n13057;
	wire n13058;
	wire n13059;
	wire n13060;
	wire n13061;
	wire n13062;
	wire n13063;
	wire n13064;
	wire n13065;
	wire n13066;
	wire n13067;
	wire n13068;
	wire n13069;
	wire n13070;
	wire n13071;
	wire n13072;
	wire n13073;
	wire n13074;
	wire n13075;
	wire n13076;
	wire n13077;
	wire n13078;
	wire n13079;
	wire n13080;
	wire n13081;
	wire n13082;
	wire n13083;
	wire n13084;
	wire n13085;
	wire n13086;
	wire n13087;
	wire n13088;
	wire n13089;
	wire n13090;
	wire n13091;
	wire n13092;
	wire n13093;
	wire n13094;
	wire n13095;
	wire n13096;
	wire n13097;
	wire n13098;
	wire n13099;
	wire n13100;
	wire n13101;
	wire n13102;
	wire n13103;
	wire n13104;
	wire n13105;
	wire n13106;
	wire n13107;
	wire n13108;
	wire n13109;
	wire n13110;
	wire n13111;
	wire n13112;
	wire n13113;
	wire n13114;
	wire n13115;
	wire n13116;
	wire n13117;
	wire n13118;
	wire n13119;
	wire n13120;
	wire n13121;
	wire n13122;
	wire n13123;
	wire n13124;
	wire n13125;
	wire n13126;
	wire n13127;
	wire n13128;
	wire n13129;
	wire n13130;
	wire n13131;
	wire n13132;
	wire n13133;
	wire n13134;
	wire n13135;
	wire n13136;
	wire n13137;
	wire n13138;
	wire n13139;
	wire n13140;
	wire n13141;
	wire n13142;
	wire n13143;
	wire n13144;
	wire n13145;
	wire n13146;
	wire n13147;
	wire n13148;
	wire n13149;
	wire n13150;
	wire n13151;
	wire n13152;
	wire n13153;
	wire n13154;
	wire n13155;
	wire n13156;
	wire n13157;
	wire n13158;
	wire n13159;
	wire n13160;
	wire n13161;
	wire n13162;
	wire n13163;
	wire n13164;
	wire n13165;
	wire n13166;
	wire n13167;
	wire n13170;
	wire n13172;
	wire n13173;
	wire n13174;
	wire n13175;
	wire n13176;
	wire n13177;
	wire n13178;
	wire n13179;
	wire n13180;
	wire n13181;
	wire n13182;
	wire n13183;
	wire n13184;
	wire n13185;
	wire n13186;
	wire n13187;
	wire n13188;
	wire n13189;
	wire n13190;
	wire n13191;
	wire n13192;
	wire n13193;
	wire n13194;
	wire n13195;
	wire n13196;
	wire n13197;
	wire n13198;
	wire n13199;
	wire n13200;
	wire n13201;
	wire n13202;
	wire n13203;
	wire n13204;
	wire n13205;
	wire n13206;
	wire n13207;
	wire n13208;
	wire n13209;
	wire n13210;
	wire n13211;
	wire n13212;
	wire n13213;
	wire n13214;
	wire n13215;
	wire n13216;
	wire n13217;
	wire n13218;
	wire n13219;
	wire n13220;
	wire n13221;
	wire n13222;
	wire n13223;
	wire n13224;
	wire n13225;
	wire n13226;
	wire n13227;
	wire n13228;
	wire n13229;
	wire n13230;
	wire n13231;
	wire n13232;
	wire n13233;
	wire n13234;
	wire n13235;
	wire n13236;
	wire n13237;
	wire n13238;
	wire n13239;
	wire n13240;
	wire n13241;
	wire n13242;
	wire n13243;
	wire n13244;
	wire n13245;
	wire n13246;
	wire n13247;
	wire n13248;
	wire n13249;
	wire n13250;
	wire n13251;
	wire n13252;
	wire n13253;
	wire n13254;
	wire n13255;
	wire n13256;
	wire n13257;
	wire n13258;
	wire n13259;
	wire n13260;
	wire n13261;
	wire n13262;
	wire n13263;
	wire n13264;
	wire n13265;
	wire n13266;
	wire n13267;
	wire n13268;
	wire n13269;
	wire n13270;
	wire n13271;
	wire n13272;
	wire n13273;
	wire n13274;
	wire n13275;
	wire n13276;
	wire n13277;
	wire n13278;
	wire n13279;
	wire n13280;
	wire n13281;
	wire n13282;
	wire n13283;
	wire n13284;
	wire n13285;
	wire n13286;
	wire n13287;
	wire n13288;
	wire n13289;
	wire n13290;
	wire n13291;
	wire n13292;
	wire n13293;
	wire n13294;
	wire n13295;
	wire n13296;
	wire n13297;
	wire n13298;
	wire n13299;
	wire n13300;
	wire n13301;
	wire n13302;
	wire n13303;
	wire n13304;
	wire n13305;
	wire n13306;
	wire n13307;
	wire n13308;
	wire n13309;
	wire n13310;
	wire n13311;
	wire n13312;
	wire n13313;
	wire n13314;
	wire n13315;
	wire n13316;
	wire n13317;
	wire n13318;
	wire n13319;
	wire n13320;
	wire n13321;
	wire n13322;
	wire n13323;
	wire n13324;
	wire n13325;
	wire n13326;
	wire n13327;
	wire n13328;
	wire n13329;
	wire n13330;
	wire n13331;
	wire n13332;
	wire n13333;
	wire n13334;
	wire n13335;
	wire n13336;
	wire n13337;
	wire n13338;
	wire n13339;
	wire n13340;
	wire n13341;
	wire n13342;
	wire n13343;
	wire n13344;
	wire n13345;
	wire n13346;
	wire n13347;
	wire n13348;
	wire n13349;
	wire n13350;
	wire n13351;
	wire n13352;
	wire n13353;
	wire n13354;
	wire n13355;
	wire n13356;
	wire n13357;
	wire n13358;
	wire n13359;
	wire n13360;
	wire n13361;
	wire n13362;
	wire n13363;
	wire n13364;
	wire n13365;
	wire n13366;
	wire n13367;
	wire n13368;
	wire n13369;
	wire n13370;
	wire n13371;
	wire n13372;
	wire n13373;
	wire n13374;
	wire n13375;
	wire n13376;
	wire n13377;
	wire n13378;
	wire n13379;
	wire n13380;
	wire n13381;
	wire n13382;
	wire n13383;
	wire n13384;
	wire n13385;
	wire n13386;
	wire n13387;
	wire n13388;
	wire n13389;
	wire n13390;
	wire n13391;
	wire n13392;
	wire n13393;
	wire n13394;
	wire n13395;
	wire n13396;
	wire n13397;
	wire n13398;
	wire n13399;
	wire n13400;
	wire n13401;
	wire n13402;
	wire n13403;
	wire n13404;
	wire n13405;
	wire n13406;
	wire n13407;
	wire n13408;
	wire n13409;
	wire n13410;
	wire n13411;
	wire n13412;
	wire n13413;
	wire n13414;
	wire n13415;
	wire n13416;
	wire n13417;
	wire n13418;
	wire n13419;
	wire n13420;
	wire n13421;
	wire n13422;
	wire n13423;
	wire n13424;
	wire n13425;
	wire n13426;
	wire n13427;
	wire n13428;
	wire n13429;
	wire n13430;
	wire n13431;
	wire n13432;
	wire n13433;
	wire n13434;
	wire n13435;
	wire n13436;
	wire n13437;
	wire n13438;
	wire n13439;
	wire n13440;
	wire n13441;
	wire n13442;
	wire n13443;
	wire n13444;
	wire n13445;
	wire n13446;
	wire n13447;
	wire n13448;
	wire n13449;
	wire n13450;
	wire n13451;
	wire n13452;
	wire n13453;
	wire n13454;
	wire n13455;
	wire n13456;
	wire n13457;
	wire n13458;
	wire n13459;
	wire n13460;
	wire n13461;
	wire n13462;
	wire n13463;
	wire n13464;
	wire n13465;
	wire n13466;
	wire n13467;
	wire n13468;
	wire n13469;
	wire n13470;
	wire n13471;
	wire n13472;
	wire n13473;
	wire n13474;
	wire n13475;
	wire n13476;
	wire n13477;
	wire n13478;
	wire n13479;
	wire n13480;
	wire n13481;
	wire n13482;
	wire n13483;
	wire n13484;
	wire n13485;
	wire n13486;
	wire n13487;
	wire n13488;
	wire n13489;
	wire n13490;
	wire n13491;
	wire n13492;
	wire n13493;
	wire n13494;
	wire n13495;
	wire n13496;
	wire n13497;
	wire n13498;
	wire n13499;
	wire n13500;
	wire n13501;
	wire n13502;
	wire n13503;
	wire n13504;
	wire n13505;
	wire n13506;
	wire n13507;
	wire n13508;
	wire n13509;
	wire n13510;
	wire n13511;
	wire n13512;
	wire n13513;
	wire n13514;
	wire n13515;
	wire n13516;
	wire n13517;
	wire n13518;
	wire n13519;
	wire n13520;
	wire n13521;
	wire n13522;
	wire n13523;
	wire n13524;
	wire n13525;
	wire n13526;
	wire n13527;
	wire n13528;
	wire n13529;
	wire n13530;
	wire n13531;
	wire n13532;
	wire n13533;
	wire n13534;
	wire n13535;
	wire n13536;
	wire n13537;
	wire n13538;
	wire n13539;
	wire n13540;
	wire n13541;
	wire n13542;
	wire n13543;
	wire n13544;
	wire n13545;
	wire n13546;
	wire n13547;
	wire n13548;
	wire n13549;
	wire n13550;
	wire n13551;
	wire n13552;
	wire n13553;
	wire n13554;
	wire n13555;
	wire n13556;
	wire n13557;
	wire n13558;
	wire n13559;
	wire n13560;
	wire n13561;
	wire n13562;
	wire n13563;
	wire n13564;
	wire n13565;
	wire n13566;
	wire n13567;
	wire n13568;
	wire n13569;
	wire n13570;
	wire n13571;
	wire n13572;
	wire n13573;
	wire n13574;
	wire n13575;
	wire n13576;
	wire n13577;
	wire n13578;
	wire n13579;
	wire n13580;
	wire n13581;
	wire n13582;
	wire n13583;
	wire n13584;
	wire n13585;
	wire n13586;
	wire n13587;
	wire n13588;
	wire n13589;
	wire n13590;
	wire n13591;
	wire n13592;
	wire n13593;
	wire n13594;
	wire n13595;
	wire n13596;
	wire n13597;
	wire n13598;
	wire n13599;
	wire n13600;
	wire n13601;
	wire n13602;
	wire n13603;
	wire n13604;
	wire n13605;
	wire n13606;
	wire n13607;
	wire n13608;
	wire n13609;
	wire n13610;
	wire n13611;
	wire n13612;
	wire n13613;
	wire n13614;
	wire n13615;
	wire n13616;
	wire n13617;
	wire n13618;
	wire n13619;
	wire n13620;
	wire n13621;
	wire n13622;
	wire n13623;
	wire n13624;
	wire n13625;
	wire n13626;
	wire n13627;
	wire n13628;
	wire n13629;
	wire n13630;
	wire n13631;
	wire n13632;
	wire n13633;
	wire n13634;
	wire n13635;
	wire n13636;
	wire n13637;
	wire n13638;
	wire n13639;
	wire n13640;
	wire n13641;
	wire n13642;
	wire n13643;
	wire n13644;
	wire n13645;
	wire n13646;
	wire n13647;
	wire n13648;
	wire n13649;
	wire n13650;
	wire n13651;
	wire n13652;
	wire n13653;
	wire n13654;
	wire n13655;
	wire n13656;
	wire n13657;
	wire n13658;
	wire n13659;
	wire n13660;
	wire n13661;
	wire n13662;
	wire n13663;
	wire n13664;
	wire n13665;
	wire n13666;
	wire n13667;
	wire n13668;
	wire n13669;
	wire n13670;
	wire n13671;
	wire n13672;
	wire n13673;
	wire n13674;
	wire n13675;
	wire n13676;
	wire n13677;
	wire n13678;
	wire n13679;
	wire n13680;
	wire n13681;
	wire n13682;
	wire n13683;
	wire n13684;
	wire n13685;
	wire n13686;
	wire n13687;
	wire n13688;
	wire n13689;
	wire n13690;
	wire n13691;
	wire n13692;
	wire n13693;
	wire n13694;
	wire n13695;
	wire n13696;
	wire n13697;
	wire n13698;
	wire n13699;
	wire n13700;
	wire n13701;
	wire n13702;
	wire n13703;
	wire n13704;
	wire n13705;
	wire n13706;
	wire n13707;
	wire n13708;
	wire n13709;
	wire n13710;
	wire n13711;
	wire n13712;
	wire n13713;
	wire n13714;
	wire n13715;
	wire n13716;
	wire n13717;
	wire n13718;
	wire n13721;
	wire n13722;
	wire n13723;
	wire n13724;
	wire n13725;
	wire n13726;
	wire n13727;
	wire n13728;
	wire n13729;
	wire n13730;
	wire n13731;
	wire n13732;
	wire n13733;
	wire n13734;
	wire n13735;
	wire n13736;
	wire n13737;
	wire n13738;
	wire n13739;
	wire n13740;
	wire n13741;
	wire n13742;
	wire n13743;
	wire n13744;
	wire n13745;
	wire n13746;
	wire n13747;
	wire n13748;
	wire n13749;
	wire n13750;
	wire n13751;
	wire n13752;
	wire n13753;
	wire n13754;
	wire n13755;
	wire n13756;
	wire n13757;
	wire n13758;
	wire n13759;
	wire n13760;
	wire n13761;
	wire n13762;
	wire n13763;
	wire n13764;
	wire n13765;
	wire n13766;
	wire n13767;
	wire n13768;
	wire n13769;
	wire n13770;
	wire n13771;
	wire n13772;
	wire n13773;
	wire n13774;
	wire n13775;
	wire n13776;
	wire n13777;
	wire n13778;
	wire n13779;
	wire n13780;
	wire n13782;
	wire n13783;
	wire n13784;
	wire n13785;
	wire n13786;
	wire n13787;
	wire n13788;
	wire n13789;
	wire n13790;
	wire n13791;
	wire n13792;
	wire n13793;
	wire n13794;
	wire n13795;
	wire n13796;
	wire n13797;
	wire n13798;
	wire n13799;
	wire n13800;
	wire n13801;
	wire n13802;
	wire n13803;
	wire n13804;
	wire n13805;
	wire n13806;
	wire n13807;
	wire n13808;
	wire n13809;
	wire n13810;
	wire n13811;
	wire n13812;
	wire n13813;
	wire n13814;
	wire n13815;
	wire n13816;
	wire n13817;
	wire n13818;
	wire n13819;
	wire n13820;
	wire n13821;
	wire n13822;
	wire n13823;
	wire n13824;
	wire n13825;
	wire n13826;
	wire n13827;
	wire n13828;
	wire n13829;
	wire n13830;
	wire n13831;
	wire n13832;
	wire n13833;
	wire n13834;
	wire n13835;
	wire n13836;
	wire n13837;
	wire n13838;
	wire n13839;
	wire n13840;
	wire n13841;
	wire n13842;
	wire n13843;
	wire n13844;
	wire n13845;
	wire n13846;
	wire n13847;
	wire n13848;
	wire n13849;
	wire n13850;
	wire n13851;
	wire n13852;
	wire n13853;
	wire n13854;
	wire n13855;
	wire n13856;
	wire n13857;
	wire n13858;
	wire n13859;
	wire n13860;
	wire n13861;
	wire n13862;
	wire n13863;
	wire n13864;
	wire n13865;
	wire n13866;
	wire n13867;
	wire n13868;
	wire n13869;
	wire n13870;
	wire n13871;
	wire n13872;
	wire n13873;
	wire n13874;
	wire n13875;
	wire n13876;
	wire n13877;
	wire n13878;
	wire n13879;
	wire n13880;
	wire n13881;
	wire n13882;
	wire n13883;
	wire n13884;
	wire n13885;
	wire n13886;
	wire n13887;
	wire n13888;
	wire n13889;
	wire n13890;
	wire n13891;
	wire n13892;
	wire n13893;
	wire n13894;
	wire n13895;
	wire n13896;
	wire n13897;
	wire n13898;
	wire n13899;
	wire n13900;
	wire n13901;
	wire n13902;
	wire n13903;
	wire n13904;
	wire n13905;
	wire n13906;
	wire n13907;
	wire n13908;
	wire n13909;
	wire n13910;
	wire n13911;
	wire n13912;
	wire n13913;
	wire n13914;
	wire n13915;
	wire n13916;
	wire n13917;
	wire n13918;
	wire n13919;
	wire n13920;
	wire n13921;
	wire n13922;
	wire n13923;
	wire n13924;
	wire n13925;
	wire n13926;
	wire n13927;
	wire n13928;
	wire n13929;
	wire n13930;
	wire n13931;
	wire n13932;
	wire n13933;
	wire n13934;
	wire n13935;
	wire n13936;
	wire n13937;
	wire n13938;
	wire n13939;
	wire n13940;
	wire n13941;
	wire n13942;
	wire n13943;
	wire n13944;
	wire n13945;
	wire n13946;
	wire n13947;
	wire n13948;
	wire n13949;
	wire n13950;
	wire n13951;
	wire n13952;
	wire n13953;
	wire n13954;
	wire n13955;
	wire n13956;
	wire n13957;
	wire n13958;
	wire n13959;
	wire n13960;
	wire n13961;
	wire n13962;
	wire n13963;
	wire n13964;
	wire n13965;
	wire n13966;
	wire n13967;
	wire n13968;
	wire n13969;
	wire n13970;
	wire n13971;
	wire n13972;
	wire n13973;
	wire n13974;
	wire n13975;
	wire n13976;
	wire n13977;
	wire n13978;
	wire n13979;
	wire n13980;
	wire n13981;
	wire n13982;
	wire n13983;
	wire n13984;
	wire n13985;
	wire n13986;
	wire n13987;
	wire n13988;
	wire n13989;
	wire n13990;
	wire n13991;
	wire n13992;
	wire n13993;
	wire n13994;
	wire n13995;
	wire n13996;
	wire n13997;
	wire n13998;
	wire n13999;
	wire n14000;
	wire n14001;
	wire n14002;
	wire n14003;
	wire n14004;
	wire n14005;
	wire n14006;
	wire n14007;
	wire n14008;
	wire n14009;
	wire n14010;
	wire n14011;
	wire n14012;
	wire n14013;
	wire n14014;
	wire n14015;
	wire n14016;
	wire n14017;
	wire n14018;
	wire n14019;
	wire n14020;
	wire n14021;
	wire n14022;
	wire n14023;
	wire n14024;
	wire n14025;
	wire n14026;
	wire n14027;
	wire n14028;
	wire n14029;
	wire n14030;
	wire n14031;
	wire n14032;
	wire n14033;
	wire n14034;
	wire n14035;
	wire n14036;
	wire n14037;
	wire n14038;
	wire n14039;
	wire n14040;
	wire n14041;
	wire n14042;
	wire n14043;
	wire n14044;
	wire n14045;
	wire n14046;
	wire n14047;
	wire n14048;
	wire n14049;
	wire n14050;
	wire n14051;
	wire n14052;
	wire n14053;
	wire n14054;
	wire n14055;
	wire n14056;
	wire n14057;
	wire n14058;
	wire n14059;
	wire n14060;
	wire n14061;
	wire n14062;
	wire n14063;
	wire n14064;
	wire n14065;
	wire n14066;
	wire n14067;
	wire n14068;
	wire n14069;
	wire n14070;
	wire n14071;
	wire n14072;
	wire n14073;
	wire n14074;
	wire n14075;
	wire n14076;
	wire n14077;
	wire n14078;
	wire n14079;
	wire n14080;
	wire n14081;
	wire n14082;
	wire n14083;
	wire n14084;
	wire n14085;
	wire n14086;
	wire n14087;
	wire n14088;
	wire n14089;
	wire n14090;
	wire n14091;
	wire n14092;
	wire n14093;
	wire n14094;
	wire n14095;
	wire n14096;
	wire n14097;
	wire n14098;
	wire n14099;
	wire n14100;
	wire n14101;
	wire n14102;
	wire n14103;
	wire n14104;
	wire n14105;
	wire n14106;
	wire n14107;
	wire n14108;
	wire n14109;
	wire n14110;
	wire n14111;
	wire n14112;
	wire n14113;
	wire n14114;
	wire n14115;
	wire n14116;
	wire n14117;
	wire n14118;
	wire n14119;
	wire n14120;
	wire n14121;
	wire n14122;
	wire n14123;
	wire n14124;
	wire n14125;
	wire n14126;
	wire n14127;
	wire n14128;
	wire n14129;
	wire n14130;
	wire n14131;
	wire n14132;
	wire n14133;
	wire n14134;
	wire n14135;
	wire n14136;
	wire n14137;
	wire n14138;
	wire n14139;
	wire n14140;
	wire n14141;
	wire n14142;
	wire n14143;
	wire n14144;
	wire n14145;
	wire n14146;
	wire n14147;
	wire n14148;
	wire n14149;
	wire n14150;
	wire n14151;
	wire n14152;
	wire n14153;
	wire n14154;
	wire n14155;
	wire n14156;
	wire n14157;
	wire n14158;
	wire n14159;
	wire n14160;
	wire n14161;
	wire n14162;
	wire n14163;
	wire n14164;
	wire n14165;
	wire n14166;
	wire n14167;
	wire n14168;
	wire n14169;
	wire n14170;
	wire n14171;
	wire n14172;
	wire n14173;
	wire n14174;
	wire n14175;
	wire n14176;
	wire n14177;
	wire n14178;
	wire n14179;
	wire n14180;
	wire n14181;
	wire n14182;
	wire n14183;
	wire n14184;
	wire n14185;
	wire n14186;
	wire n14187;
	wire n14188;
	wire n14189;
	wire n14190;
	wire n14191;
	wire n14192;
	wire n14193;
	wire n14194;
	wire n14195;
	wire n14196;
	wire n14197;
	wire n14198;
	wire n14199;
	wire n14200;
	wire n14201;
	wire n14202;
	wire n14203;
	wire n14204;
	wire n14205;
	wire n14206;
	wire n14207;
	wire n14208;
	wire n14209;
	wire n14210;
	wire n14211;
	wire n14212;
	wire n14213;
	wire n14214;
	wire n14215;
	wire n14216;
	wire n14217;
	wire n14218;
	wire n14219;
	wire n14220;
	wire n14221;
	wire n14222;
	wire n14223;
	wire n14224;
	wire n14225;
	wire n14226;
	wire n14227;
	wire n14228;
	wire n14229;
	wire n14230;
	wire n14231;
	wire n14232;
	wire n14233;
	wire n14234;
	wire n14235;
	wire n14236;
	wire n14237;
	wire n14238;
	wire n14239;
	wire n14242;
	wire n14244;
	wire n14245;
	wire n14246;
	wire n14247;
	wire n14248;
	wire n14249;
	wire n14250;
	wire n14251;
	wire n14252;
	wire n14253;
	wire n14254;
	wire n14255;
	wire n14256;
	wire n14257;
	wire n14258;
	wire n14259;
	wire n14260;
	wire n14261;
	wire n14262;
	wire n14263;
	wire n14264;
	wire n14265;
	wire n14266;
	wire n14267;
	wire n14268;
	wire n14269;
	wire n14270;
	wire n14271;
	wire n14272;
	wire n14273;
	wire n14274;
	wire n14275;
	wire n14276;
	wire n14277;
	wire n14278;
	wire n14279;
	wire n14280;
	wire n14281;
	wire n14282;
	wire n14283;
	wire n14284;
	wire n14285;
	wire n14286;
	wire n14287;
	wire n14288;
	wire n14289;
	wire n14290;
	wire n14291;
	wire n14292;
	wire n14293;
	wire n14294;
	wire n14295;
	wire n14296;
	wire n14297;
	wire n14298;
	wire n14299;
	wire n14300;
	wire n14301;
	wire n14302;
	wire n14303;
	wire n14304;
	wire n14305;
	wire n14306;
	wire n14307;
	wire n14308;
	wire n14309;
	wire n14310;
	wire n14311;
	wire n14312;
	wire n14313;
	wire n14314;
	wire n14315;
	wire n14316;
	wire n14317;
	wire n14318;
	wire n14319;
	wire n14320;
	wire n14321;
	wire n14322;
	wire n14323;
	wire n14324;
	wire n14325;
	wire n14326;
	wire n14327;
	wire n14328;
	wire n14329;
	wire n14330;
	wire n14331;
	wire n14332;
	wire n14333;
	wire n14334;
	wire n14335;
	wire n14336;
	wire n14337;
	wire n14338;
	wire n14339;
	wire n14340;
	wire n14341;
	wire n14342;
	wire n14343;
	wire n14344;
	wire n14345;
	wire n14346;
	wire n14347;
	wire n14348;
	wire n14349;
	wire n14350;
	wire n14351;
	wire n14352;
	wire n14353;
	wire n14354;
	wire n14355;
	wire n14356;
	wire n14357;
	wire n14358;
	wire n14359;
	wire n14360;
	wire n14361;
	wire n14362;
	wire n14363;
	wire n14364;
	wire n14365;
	wire n14366;
	wire n14367;
	wire n14368;
	wire n14369;
	wire n14370;
	wire n14371;
	wire n14372;
	wire n14373;
	wire n14374;
	wire n14375;
	wire n14376;
	wire n14377;
	wire n14378;
	wire n14379;
	wire n14380;
	wire n14381;
	wire n14382;
	wire n14383;
	wire n14384;
	wire n14385;
	wire n14386;
	wire n14387;
	wire n14388;
	wire n14389;
	wire n14390;
	wire n14391;
	wire n14392;
	wire n14393;
	wire n14394;
	wire n14395;
	wire n14396;
	wire n14397;
	wire n14398;
	wire n14399;
	wire n14400;
	wire n14401;
	wire n14402;
	wire n14403;
	wire n14404;
	wire n14405;
	wire n14406;
	wire n14407;
	wire n14408;
	wire n14409;
	wire n14410;
	wire n14411;
	wire n14412;
	wire n14413;
	wire n14414;
	wire n14415;
	wire n14416;
	wire n14417;
	wire n14418;
	wire n14419;
	wire n14420;
	wire n14421;
	wire n14422;
	wire n14423;
	wire n14424;
	wire n14425;
	wire n14426;
	wire n14427;
	wire n14428;
	wire n14429;
	wire n14430;
	wire n14431;
	wire n14432;
	wire n14433;
	wire n14434;
	wire n14435;
	wire n14436;
	wire n14437;
	wire n14438;
	wire n14439;
	wire n14440;
	wire n14441;
	wire n14442;
	wire n14443;
	wire n14444;
	wire n14445;
	wire n14446;
	wire n14447;
	wire n14448;
	wire n14449;
	wire n14450;
	wire n14451;
	wire n14452;
	wire n14453;
	wire n14454;
	wire n14455;
	wire n14456;
	wire n14457;
	wire n14458;
	wire n14459;
	wire n14460;
	wire n14461;
	wire n14462;
	wire n14463;
	wire n14464;
	wire n14465;
	wire n14466;
	wire n14467;
	wire n14468;
	wire n14469;
	wire n14470;
	wire n14471;
	wire n14472;
	wire n14473;
	wire n14474;
	wire n14475;
	wire n14476;
	wire n14477;
	wire n14478;
	wire n14479;
	wire n14480;
	wire n14481;
	wire n14482;
	wire n14483;
	wire n14484;
	wire n14485;
	wire n14486;
	wire n14487;
	wire n14488;
	wire n14489;
	wire n14490;
	wire n14491;
	wire n14492;
	wire n14493;
	wire n14494;
	wire n14495;
	wire n14496;
	wire n14497;
	wire n14498;
	wire n14499;
	wire n14500;
	wire n14501;
	wire n14502;
	wire n14503;
	wire n14504;
	wire n14505;
	wire n14506;
	wire n14507;
	wire n14508;
	wire n14509;
	wire n14510;
	wire n14511;
	wire n14512;
	wire n14513;
	wire n14514;
	wire n14515;
	wire n14516;
	wire n14517;
	wire n14518;
	wire n14519;
	wire n14520;
	wire n14521;
	wire n14522;
	wire n14523;
	wire n14524;
	wire n14525;
	wire n14526;
	wire n14527;
	wire n14528;
	wire n14529;
	wire n14530;
	wire n14531;
	wire n14532;
	wire n14533;
	wire n14534;
	wire n14535;
	wire n14536;
	wire n14537;
	wire n14538;
	wire n14539;
	wire n14540;
	wire n14541;
	wire n14542;
	wire n14543;
	wire n14544;
	wire n14545;
	wire n14546;
	wire n14547;
	wire n14548;
	wire n14549;
	wire n14550;
	wire n14551;
	wire n14552;
	wire n14553;
	wire n14554;
	wire n14555;
	wire n14556;
	wire n14557;
	wire n14558;
	wire n14559;
	wire n14560;
	wire n14561;
	wire n14562;
	wire n14563;
	wire n14564;
	wire n14565;
	wire n14566;
	wire n14567;
	wire n14568;
	wire n14569;
	wire n14570;
	wire n14571;
	wire n14572;
	wire n14573;
	wire n14574;
	wire n14575;
	wire n14576;
	wire n14577;
	wire n14578;
	wire n14579;
	wire n14580;
	wire n14581;
	wire n14582;
	wire n14583;
	wire n14584;
	wire n14585;
	wire n14586;
	wire n14587;
	wire n14588;
	wire n14589;
	wire n14590;
	wire n14591;
	wire n14592;
	wire n14593;
	wire n14594;
	wire n14595;
	wire n14596;
	wire n14597;
	wire n14598;
	wire n14599;
	wire n14600;
	wire n14601;
	wire n14602;
	wire n14603;
	wire n14604;
	wire n14605;
	wire n14606;
	wire n14607;
	wire n14608;
	wire n14609;
	wire n14610;
	wire n14611;
	wire n14612;
	wire n14613;
	wire n14614;
	wire n14615;
	wire n14616;
	wire n14617;
	wire n14618;
	wire n14619;
	wire n14620;
	wire n14621;
	wire n14622;
	wire n14623;
	wire n14624;
	wire n14625;
	wire n14626;
	wire n14627;
	wire n14628;
	wire n14629;
	wire n14630;
	wire n14631;
	wire n14632;
	wire n14633;
	wire n14634;
	wire n14635;
	wire n14636;
	wire n14637;
	wire n14638;
	wire n14639;
	wire n14640;
	wire n14641;
	wire n14642;
	wire n14643;
	wire n14644;
	wire n14645;
	wire n14646;
	wire n14647;
	wire n14648;
	wire n14649;
	wire n14650;
	wire n14651;
	wire n14652;
	wire n14653;
	wire n14654;
	wire n14655;
	wire n14656;
	wire n14657;
	wire n14658;
	wire n14659;
	wire n14660;
	wire n14661;
	wire n14662;
	wire n14663;
	wire n14664;
	wire n14665;
	wire n14666;
	wire n14667;
	wire n14668;
	wire n14669;
	wire n14670;
	wire n14671;
	wire n14672;
	wire n14673;
	wire n14674;
	wire n14675;
	wire n14676;
	wire n14677;
	wire n14678;
	wire n14679;
	wire n14680;
	wire n14681;
	wire n14682;
	wire n14683;
	wire n14684;
	wire n14685;
	wire n14686;
	wire n14687;
	wire n14688;
	wire n14689;
	wire n14690;
	wire n14691;
	wire n14692;
	wire n14693;
	wire n14694;
	wire n14695;
	wire n14696;
	wire n14697;
	wire n14698;
	wire n14699;
	wire n14700;
	wire n14701;
	wire n14702;
	wire n14703;
	wire n14704;
	wire n14705;
	wire n14706;
	wire n14707;
	wire n14708;
	wire n14709;
	wire n14710;
	wire n14711;
	wire n14712;
	wire n14713;
	wire n14714;
	wire n14715;
	wire n14716;
	wire n14717;
	wire n14718;
	wire n14719;
	wire n14720;
	wire n14721;
	wire n14722;
	wire n14723;
	wire n14724;
	wire n14725;
	wire n14726;
	wire n14727;
	wire n14728;
	wire n14729;
	wire n14730;
	wire n14731;
	wire n14732;
	wire n14733;
	wire n14734;
	wire n14735;
	wire n14736;
	wire n14737;
	wire n14738;
	wire n14739;
	wire n14740;
	wire n14741;
	wire n14742;
	wire n14743;
	wire n14744;
	wire n14745;
	wire n14746;
	wire n14747;
	wire n14748;
	wire n14749;
	wire n14750;
	wire n14751;
	wire n14752;
	wire n14753;
	wire n14754;
	wire n14755;
	wire n14756;
	wire n14757;
	wire n14758;
	wire n14759;
	wire n14760;
	wire n14761;
	wire n14762;
	wire n14763;
	wire n14764;
	wire n14765;
	wire n14766;
	wire n14767;
	wire n14768;
	wire n14769;
	wire n14770;
	wire n14771;
	wire n14772;
	wire n14773;
	wire n14774;
	wire n14775;
	wire n14776;
	wire n14777;
	wire n14778;
	wire n14779;
	wire n14780;
	wire n14781;
	wire n14782;
	wire n14783;
	wire n14784;
	wire n14785;
	wire n14786;
	wire n14787;
	wire n14788;
	wire n14789;
	wire n14790;
	wire n14791;
	wire n14792;
	wire n14793;
	wire n14794;
	wire n14795;
	wire n14796;
	wire n14797;
	wire n14798;
	wire n14799;
	wire n14800;
	wire n14801;
	wire n14802;
	wire n14803;
	wire n14804;
	wire n14805;
	wire n14806;
	wire n14807;
	wire n14808;
	wire n14809;
	wire n14810;
	wire n14811;
	wire n14812;
	wire n14813;
	wire n14814;
	wire n14815;
	wire n14816;
	wire n14819;
	wire n14820;
	wire n14821;
	wire n14822;
	wire n14823;
	wire n14824;
	wire n14825;
	wire n14826;
	wire n14827;
	wire n14828;
	wire n14829;
	wire n14830;
	wire n14831;
	wire n14832;
	wire n14833;
	wire n14834;
	wire n14835;
	wire n14836;
	wire n14837;
	wire n14838;
	wire n14839;
	wire n14840;
	wire n14841;
	wire n14842;
	wire n14843;
	wire n14844;
	wire n14845;
	wire n14846;
	wire n14847;
	wire n14848;
	wire n14849;
	wire n14850;
	wire n14851;
	wire n14852;
	wire n14853;
	wire n14854;
	wire n14855;
	wire n14856;
	wire n14857;
	wire n14858;
	wire n14859;
	wire n14860;
	wire n14861;
	wire n14862;
	wire n14863;
	wire n14864;
	wire n14865;
	wire n14866;
	wire n14867;
	wire n14868;
	wire n14869;
	wire n14870;
	wire n14871;
	wire n14872;
	wire n14873;
	wire n14874;
	wire n14875;
	wire n14876;
	wire n14877;
	wire n14878;
	wire n14880;
	wire n14881;
	wire n14882;
	wire n14883;
	wire n14884;
	wire n14885;
	wire n14886;
	wire n14887;
	wire n14888;
	wire n14889;
	wire n14890;
	wire n14891;
	wire n14892;
	wire n14893;
	wire n14894;
	wire n14895;
	wire n14896;
	wire n14897;
	wire n14898;
	wire n14899;
	wire n14900;
	wire n14901;
	wire n14902;
	wire n14903;
	wire n14904;
	wire n14905;
	wire n14906;
	wire n14907;
	wire n14908;
	wire n14909;
	wire n14910;
	wire n14911;
	wire n14912;
	wire n14913;
	wire n14914;
	wire n14915;
	wire n14916;
	wire n14917;
	wire n14918;
	wire n14919;
	wire n14920;
	wire n14921;
	wire n14922;
	wire n14923;
	wire n14924;
	wire n14925;
	wire n14926;
	wire n14927;
	wire n14928;
	wire n14929;
	wire n14930;
	wire n14931;
	wire n14932;
	wire n14933;
	wire n14934;
	wire n14935;
	wire n14936;
	wire n14937;
	wire n14938;
	wire n14939;
	wire n14940;
	wire n14941;
	wire n14942;
	wire n14943;
	wire n14944;
	wire n14945;
	wire n14946;
	wire n14947;
	wire n14948;
	wire n14949;
	wire n14950;
	wire n14951;
	wire n14952;
	wire n14953;
	wire n14954;
	wire n14955;
	wire n14956;
	wire n14957;
	wire n14958;
	wire n14959;
	wire n14960;
	wire n14961;
	wire n14962;
	wire n14963;
	wire n14964;
	wire n14965;
	wire n14966;
	wire n14967;
	wire n14968;
	wire n14969;
	wire n14970;
	wire n14971;
	wire n14972;
	wire n14973;
	wire n14974;
	wire n14975;
	wire n14976;
	wire n14977;
	wire n14978;
	wire n14979;
	wire n14980;
	wire n14981;
	wire n14982;
	wire n14983;
	wire n14984;
	wire n14985;
	wire n14986;
	wire n14987;
	wire n14988;
	wire n14989;
	wire n14990;
	wire n14991;
	wire n14992;
	wire n14993;
	wire n14994;
	wire n14995;
	wire n14996;
	wire n14997;
	wire n14998;
	wire n14999;
	wire n15000;
	wire n15001;
	wire n15002;
	wire n15003;
	wire n15004;
	wire n15005;
	wire n15006;
	wire n15007;
	wire n15008;
	wire n15009;
	wire n15010;
	wire n15011;
	wire n15012;
	wire n15013;
	wire n15014;
	wire n15015;
	wire n15016;
	wire n15017;
	wire n15018;
	wire n15019;
	wire n15020;
	wire n15021;
	wire n15022;
	wire n15023;
	wire n15024;
	wire n15025;
	wire n15026;
	wire n15027;
	wire n15028;
	wire n15029;
	wire n15030;
	wire n15031;
	wire n15032;
	wire n15033;
	wire n15034;
	wire n15035;
	wire n15036;
	wire n15037;
	wire n15038;
	wire n15039;
	wire n15040;
	wire n15041;
	wire n15042;
	wire n15043;
	wire n15044;
	wire n15045;
	wire n15046;
	wire n15047;
	wire n15048;
	wire n15049;
	wire n15050;
	wire n15051;
	wire n15052;
	wire n15053;
	wire n15054;
	wire n15055;
	wire n15056;
	wire n15057;
	wire n15058;
	wire n15059;
	wire n15060;
	wire n15061;
	wire n15062;
	wire n15063;
	wire n15064;
	wire n15065;
	wire n15066;
	wire n15067;
	wire n15068;
	wire n15069;
	wire n15070;
	wire n15071;
	wire n15072;
	wire n15073;
	wire n15074;
	wire n15075;
	wire n15076;
	wire n15077;
	wire n15078;
	wire n15079;
	wire n15080;
	wire n15081;
	wire n15082;
	wire n15083;
	wire n15084;
	wire n15085;
	wire n15086;
	wire n15087;
	wire n15088;
	wire n15089;
	wire n15090;
	wire n15091;
	wire n15092;
	wire n15093;
	wire n15094;
	wire n15095;
	wire n15096;
	wire n15097;
	wire n15098;
	wire n15099;
	wire n15100;
	wire n15101;
	wire n15102;
	wire n15103;
	wire n15104;
	wire n15105;
	wire n15106;
	wire n15107;
	wire n15108;
	wire n15109;
	wire n15110;
	wire n15111;
	wire n15112;
	wire n15113;
	wire n15114;
	wire n15115;
	wire n15116;
	wire n15117;
	wire n15118;
	wire n15119;
	wire n15120;
	wire n15121;
	wire n15122;
	wire n15123;
	wire n15124;
	wire n15125;
	wire n15126;
	wire n15127;
	wire n15128;
	wire n15129;
	wire n15130;
	wire n15131;
	wire n15132;
	wire n15133;
	wire n15134;
	wire n15135;
	wire n15136;
	wire n15137;
	wire n15138;
	wire n15139;
	wire n15140;
	wire n15141;
	wire n15142;
	wire n15143;
	wire n15144;
	wire n15145;
	wire n15146;
	wire n15147;
	wire n15148;
	wire n15149;
	wire n15150;
	wire n15151;
	wire n15152;
	wire n15153;
	wire n15154;
	wire n15155;
	wire n15156;
	wire n15157;
	wire n15158;
	wire n15159;
	wire n15160;
	wire n15161;
	wire n15162;
	wire n15163;
	wire n15164;
	wire n15165;
	wire n15166;
	wire n15167;
	wire n15168;
	wire n15169;
	wire n15170;
	wire n15171;
	wire n15172;
	wire n15173;
	wire n15174;
	wire n15175;
	wire n15176;
	wire n15177;
	wire n15178;
	wire n15179;
	wire n15180;
	wire n15181;
	wire n15182;
	wire n15183;
	wire n15184;
	wire n15185;
	wire n15186;
	wire n15187;
	wire n15188;
	wire n15189;
	wire n15190;
	wire n15191;
	wire n15192;
	wire n15193;
	wire n15194;
	wire n15195;
	wire n15196;
	wire n15197;
	wire n15198;
	wire n15199;
	wire n15200;
	wire n15201;
	wire n15202;
	wire n15203;
	wire n15204;
	wire n15205;
	wire n15206;
	wire n15207;
	wire n15208;
	wire n15209;
	wire n15210;
	wire n15211;
	wire n15212;
	wire n15213;
	wire n15214;
	wire n15215;
	wire n15216;
	wire n15217;
	wire n15218;
	wire n15219;
	wire n15220;
	wire n15221;
	wire n15222;
	wire n15223;
	wire n15224;
	wire n15225;
	wire n15226;
	wire n15227;
	wire n15228;
	wire n15229;
	wire n15230;
	wire n15231;
	wire n15232;
	wire n15233;
	wire n15234;
	wire n15235;
	wire n15236;
	wire n15237;
	wire n15238;
	wire n15239;
	wire n15240;
	wire n15241;
	wire n15242;
	wire n15243;
	wire n15244;
	wire n15245;
	wire n15246;
	wire n15247;
	wire n15248;
	wire n15249;
	wire n15250;
	wire n15251;
	wire n15252;
	wire n15253;
	wire n15254;
	wire n15255;
	wire n15256;
	wire n15257;
	wire n15258;
	wire n15259;
	wire n15260;
	wire n15261;
	wire n15262;
	wire n15263;
	wire n15264;
	wire n15265;
	wire n15266;
	wire n15267;
	wire n15268;
	wire n15269;
	wire n15270;
	wire n15271;
	wire n15272;
	wire n15273;
	wire n15274;
	wire n15275;
	wire n15276;
	wire n15277;
	wire n15278;
	wire n15279;
	wire n15280;
	wire n15281;
	wire n15282;
	wire n15283;
	wire n15284;
	wire n15285;
	wire n15286;
	wire n15287;
	wire n15288;
	wire n15289;
	wire n15290;
	wire n15291;
	wire n15292;
	wire n15293;
	wire n15294;
	wire n15295;
	wire n15296;
	wire n15297;
	wire n15298;
	wire n15299;
	wire n15300;
	wire n15301;
	wire n15302;
	wire n15303;
	wire n15304;
	wire n15305;
	wire n15306;
	wire n15307;
	wire n15308;
	wire n15309;
	wire n15310;
	wire n15311;
	wire n15312;
	wire n15313;
	wire n15314;
	wire n15315;
	wire n15316;
	wire n15317;
	wire n15318;
	wire n15319;
	wire n15320;
	wire n15321;
	wire n15322;
	wire n15323;
	wire n15324;
	wire n15325;
	wire n15326;
	wire n15327;
	wire n15328;
	wire n15329;
	wire n15330;
	wire n15331;
	wire n15332;
	wire n15333;
	wire n15334;
	wire n15335;
	wire n15336;
	wire n15337;
	wire n15338;
	wire n15339;
	wire n15340;
	wire n15341;
	wire n15342;
	wire n15343;
	wire n15344;
	wire n15345;
	wire n15346;
	wire n15347;
	wire n15348;
	wire n15349;
	wire n15350;
	wire n15351;
	wire n15352;
	wire n15353;
	wire n15354;
	wire n15357;
	wire n15359;
	wire n15360;
	wire n15361;
	wire n15362;
	wire n15363;
	wire n15364;
	wire n15365;
	wire n15366;
	wire n15367;
	wire n15368;
	wire n15369;
	wire n15370;
	wire n15371;
	wire n15372;
	wire n15373;
	wire n15374;
	wire n15375;
	wire n15376;
	wire n15377;
	wire n15378;
	wire n15379;
	wire n15380;
	wire n15381;
	wire n15382;
	wire n15383;
	wire n15384;
	wire n15385;
	wire n15386;
	wire n15387;
	wire n15388;
	wire n15389;
	wire n15390;
	wire n15391;
	wire n15392;
	wire n15393;
	wire n15394;
	wire n15395;
	wire n15396;
	wire n15397;
	wire n15398;
	wire n15399;
	wire n15400;
	wire n15401;
	wire n15402;
	wire n15403;
	wire n15404;
	wire n15405;
	wire n15406;
	wire n15407;
	wire n15408;
	wire n15409;
	wire n15410;
	wire n15411;
	wire n15412;
	wire n15413;
	wire n15414;
	wire n15415;
	wire n15416;
	wire n15417;
	wire n15418;
	wire n15419;
	wire n15420;
	wire n15421;
	wire n15422;
	wire n15423;
	wire n15424;
	wire n15425;
	wire n15426;
	wire n15427;
	wire n15428;
	wire n15429;
	wire n15430;
	wire n15431;
	wire n15432;
	wire n15433;
	wire n15434;
	wire n15435;
	wire n15436;
	wire n15437;
	wire n15438;
	wire n15439;
	wire n15440;
	wire n15441;
	wire n15442;
	wire n15443;
	wire n15444;
	wire n15445;
	wire n15446;
	wire n15447;
	wire n15448;
	wire n15449;
	wire n15450;
	wire n15451;
	wire n15452;
	wire n15453;
	wire n15454;
	wire n15455;
	wire n15456;
	wire n15457;
	wire n15458;
	wire n15459;
	wire n15460;
	wire n15461;
	wire n15462;
	wire n15463;
	wire n15464;
	wire n15465;
	wire n15466;
	wire n15467;
	wire n15468;
	wire n15469;
	wire n15470;
	wire n15471;
	wire n15472;
	wire n15473;
	wire n15474;
	wire n15475;
	wire n15476;
	wire n15477;
	wire n15478;
	wire n15479;
	wire n15480;
	wire n15481;
	wire n15482;
	wire n15483;
	wire n15484;
	wire n15485;
	wire n15486;
	wire n15487;
	wire n15488;
	wire n15489;
	wire n15490;
	wire n15491;
	wire n15492;
	wire n15493;
	wire n15494;
	wire n15495;
	wire n15496;
	wire n15497;
	wire n15498;
	wire n15499;
	wire n15500;
	wire n15501;
	wire n15502;
	wire n15503;
	wire n15504;
	wire n15505;
	wire n15506;
	wire n15507;
	wire n15508;
	wire n15509;
	wire n15510;
	wire n15511;
	wire n15512;
	wire n15513;
	wire n15514;
	wire n15515;
	wire n15516;
	wire n15517;
	wire n15518;
	wire n15519;
	wire n15520;
	wire n15521;
	wire n15522;
	wire n15523;
	wire n15524;
	wire n15525;
	wire n15526;
	wire n15527;
	wire n15528;
	wire n15529;
	wire n15530;
	wire n15531;
	wire n15532;
	wire n15533;
	wire n15534;
	wire n15535;
	wire n15536;
	wire n15537;
	wire n15538;
	wire n15539;
	wire n15540;
	wire n15541;
	wire n15542;
	wire n15543;
	wire n15544;
	wire n15545;
	wire n15546;
	wire n15547;
	wire n15548;
	wire n15549;
	wire n15550;
	wire n15551;
	wire n15552;
	wire n15553;
	wire n15554;
	wire n15555;
	wire n15556;
	wire n15557;
	wire n15558;
	wire n15559;
	wire n15560;
	wire n15561;
	wire n15562;
	wire n15563;
	wire n15564;
	wire n15565;
	wire n15566;
	wire n15567;
	wire n15568;
	wire n15569;
	wire n15570;
	wire n15571;
	wire n15572;
	wire n15573;
	wire n15574;
	wire n15575;
	wire n15576;
	wire n15577;
	wire n15578;
	wire n15579;
	wire n15580;
	wire n15581;
	wire n15582;
	wire n15583;
	wire n15584;
	wire n15585;
	wire n15586;
	wire n15587;
	wire n15588;
	wire n15589;
	wire n15590;
	wire n15591;
	wire n15592;
	wire n15593;
	wire n15594;
	wire n15595;
	wire n15596;
	wire n15597;
	wire n15598;
	wire n15599;
	wire n15600;
	wire n15601;
	wire n15602;
	wire n15603;
	wire n15604;
	wire n15605;
	wire n15606;
	wire n15607;
	wire n15608;
	wire n15609;
	wire n15610;
	wire n15611;
	wire n15612;
	wire n15613;
	wire n15614;
	wire n15615;
	wire n15616;
	wire n15617;
	wire n15618;
	wire n15619;
	wire n15620;
	wire n15621;
	wire n15622;
	wire n15623;
	wire n15624;
	wire n15625;
	wire n15626;
	wire n15627;
	wire n15628;
	wire n15629;
	wire n15630;
	wire n15631;
	wire n15632;
	wire n15633;
	wire n15634;
	wire n15635;
	wire n15636;
	wire n15637;
	wire n15638;
	wire n15639;
	wire n15640;
	wire n15641;
	wire n15642;
	wire n15643;
	wire n15644;
	wire n15645;
	wire n15646;
	wire n15647;
	wire n15648;
	wire n15649;
	wire n15650;
	wire n15651;
	wire n15652;
	wire n15653;
	wire n15654;
	wire n15655;
	wire n15656;
	wire n15657;
	wire n15658;
	wire n15659;
	wire n15660;
	wire n15661;
	wire n15662;
	wire n15663;
	wire n15664;
	wire n15665;
	wire n15666;
	wire n15667;
	wire n15668;
	wire n15669;
	wire n15670;
	wire n15671;
	wire n15672;
	wire n15673;
	wire n15674;
	wire n15675;
	wire n15676;
	wire n15677;
	wire n15678;
	wire n15679;
	wire n15680;
	wire n15681;
	wire n15682;
	wire n15683;
	wire n15684;
	wire n15685;
	wire n15686;
	wire n15687;
	wire n15688;
	wire n15689;
	wire n15690;
	wire n15691;
	wire n15692;
	wire n15693;
	wire n15694;
	wire n15695;
	wire n15696;
	wire n15697;
	wire n15698;
	wire n15699;
	wire n15700;
	wire n15701;
	wire n15702;
	wire n15703;
	wire n15704;
	wire n15705;
	wire n15706;
	wire n15707;
	wire n15708;
	wire n15709;
	wire n15710;
	wire n15711;
	wire n15712;
	wire n15713;
	wire n15714;
	wire n15715;
	wire n15716;
	wire n15717;
	wire n15718;
	wire n15719;
	wire n15720;
	wire n15721;
	wire n15722;
	wire n15723;
	wire n15724;
	wire n15725;
	wire n15726;
	wire n15727;
	wire n15728;
	wire n15729;
	wire n15730;
	wire n15731;
	wire n15732;
	wire n15733;
	wire n15734;
	wire n15735;
	wire n15736;
	wire n15737;
	wire n15738;
	wire n15739;
	wire n15740;
	wire n15741;
	wire n15742;
	wire n15743;
	wire n15744;
	wire n15745;
	wire n15746;
	wire n15747;
	wire n15748;
	wire n15749;
	wire n15750;
	wire n15751;
	wire n15752;
	wire n15753;
	wire n15754;
	wire n15755;
	wire n15756;
	wire n15757;
	wire n15758;
	wire n15759;
	wire n15760;
	wire n15761;
	wire n15762;
	wire n15763;
	wire n15764;
	wire n15765;
	wire n15766;
	wire n15767;
	wire n15768;
	wire n15769;
	wire n15770;
	wire n15771;
	wire n15772;
	wire n15773;
	wire n15774;
	wire n15775;
	wire n15776;
	wire n15777;
	wire n15778;
	wire n15779;
	wire n15780;
	wire n15781;
	wire n15782;
	wire n15783;
	wire n15784;
	wire n15785;
	wire n15786;
	wire n15787;
	wire n15788;
	wire n15789;
	wire n15790;
	wire n15791;
	wire n15792;
	wire n15793;
	wire n15794;
	wire n15795;
	wire n15796;
	wire n15797;
	wire n15798;
	wire n15799;
	wire n15800;
	wire n15801;
	wire n15802;
	wire n15803;
	wire n15804;
	wire n15805;
	wire n15806;
	wire n15807;
	wire n15808;
	wire n15809;
	wire n15810;
	wire n15811;
	wire n15812;
	wire n15813;
	wire n15814;
	wire n15815;
	wire n15816;
	wire n15817;
	wire n15818;
	wire n15819;
	wire n15820;
	wire n15821;
	wire n15822;
	wire n15823;
	wire n15824;
	wire n15825;
	wire n15826;
	wire n15827;
	wire n15828;
	wire n15829;
	wire n15830;
	wire n15831;
	wire n15832;
	wire n15833;
	wire n15834;
	wire n15835;
	wire n15836;
	wire n15837;
	wire n15838;
	wire n15839;
	wire n15840;
	wire n15841;
	wire n15842;
	wire n15843;
	wire n15844;
	wire n15845;
	wire n15846;
	wire n15847;
	wire n15848;
	wire n15849;
	wire n15850;
	wire n15851;
	wire n15852;
	wire n15853;
	wire n15854;
	wire n15855;
	wire n15856;
	wire n15857;
	wire n15858;
	wire n15859;
	wire n15860;
	wire n15861;
	wire n15862;
	wire n15863;
	wire n15864;
	wire n15865;
	wire n15866;
	wire n15867;
	wire n15868;
	wire n15869;
	wire n15870;
	wire n15871;
	wire n15872;
	wire n15873;
	wire n15874;
	wire n15875;
	wire n15876;
	wire n15877;
	wire n15878;
	wire n15879;
	wire n15880;
	wire n15881;
	wire n15882;
	wire n15883;
	wire n15884;
	wire n15885;
	wire n15886;
	wire n15887;
	wire n15888;
	wire n15889;
	wire n15890;
	wire n15891;
	wire n15892;
	wire n15893;
	wire n15894;
	wire n15895;
	wire n15896;
	wire n15897;
	wire n15898;
	wire n15899;
	wire n15900;
	wire n15901;
	wire n15902;
	wire n15903;
	wire n15904;
	wire n15905;
	wire n15906;
	wire n15907;
	wire n15908;
	wire n15909;
	wire n15910;
	wire n15911;
	wire n15912;
	wire n15913;
	wire n15914;
	wire n15915;
	wire n15916;
	wire n15917;
	wire n15918;
	wire n15919;
	wire n15920;
	wire n15921;
	wire n15922;
	wire n15923;
	wire n15924;
	wire n15925;
	wire n15926;
	wire n15927;
	wire n15928;
	wire n15929;
	wire n15930;
	wire n15931;
	wire n15932;
	wire n15933;
	wire n15934;
	wire n15935;
	wire n15936;
	wire n15937;
	wire n15938;
	wire n15939;
	wire n15940;
	wire n15941;
	wire n15942;
	wire n15943;
	wire n15944;
	wire n15945;
	wire n15946;
	wire n15947;
	wire n15948;
	wire n15949;
	wire n15950;
	wire n15953;
	wire n15954;
	wire n15955;
	wire n15956;
	wire n15957;
	wire n15958;
	wire n15959;
	wire n15960;
	wire n15961;
	wire n15962;
	wire n15963;
	wire n15964;
	wire n15965;
	wire n15966;
	wire n15967;
	wire n15968;
	wire n15969;
	wire n15970;
	wire n15971;
	wire n15972;
	wire n15973;
	wire n15974;
	wire n15975;
	wire n15976;
	wire n15977;
	wire n15978;
	wire n15979;
	wire n15980;
	wire n15981;
	wire n15982;
	wire n15983;
	wire n15984;
	wire n15985;
	wire n15986;
	wire n15987;
	wire n15988;
	wire n15989;
	wire n15990;
	wire n15991;
	wire n15992;
	wire n15993;
	wire n15994;
	wire n15995;
	wire n15996;
	wire n15997;
	wire n15998;
	wire n15999;
	wire n16000;
	wire n16001;
	wire n16002;
	wire n16003;
	wire n16004;
	wire n16005;
	wire n16006;
	wire n16007;
	wire n16008;
	wire n16009;
	wire n16010;
	wire n16011;
	wire n16012;
	wire n16013;
	wire n16015;
	wire n16016;
	wire n16017;
	wire n16018;
	wire n16019;
	wire n16020;
	wire n16021;
	wire n16022;
	wire n16023;
	wire n16024;
	wire n16025;
	wire n16026;
	wire n16027;
	wire n16028;
	wire n16029;
	wire n16030;
	wire n16031;
	wire n16032;
	wire n16033;
	wire n16034;
	wire n16035;
	wire n16036;
	wire n16037;
	wire n16038;
	wire n16039;
	wire n16040;
	wire n16041;
	wire n16042;
	wire n16043;
	wire n16044;
	wire n16045;
	wire n16046;
	wire n16047;
	wire n16048;
	wire n16049;
	wire n16050;
	wire n16051;
	wire n16052;
	wire n16053;
	wire n16054;
	wire n16055;
	wire n16056;
	wire n16057;
	wire n16058;
	wire n16059;
	wire n16060;
	wire n16061;
	wire n16062;
	wire n16063;
	wire n16064;
	wire n16065;
	wire n16066;
	wire n16067;
	wire n16068;
	wire n16069;
	wire n16070;
	wire n16071;
	wire n16072;
	wire n16073;
	wire n16074;
	wire n16075;
	wire n16076;
	wire n16077;
	wire n16078;
	wire n16079;
	wire n16080;
	wire n16081;
	wire n16082;
	wire n16083;
	wire n16084;
	wire n16085;
	wire n16086;
	wire n16087;
	wire n16088;
	wire n16089;
	wire n16090;
	wire n16091;
	wire n16092;
	wire n16093;
	wire n16094;
	wire n16095;
	wire n16096;
	wire n16097;
	wire n16098;
	wire n16099;
	wire n16100;
	wire n16101;
	wire n16102;
	wire n16103;
	wire n16104;
	wire n16105;
	wire n16106;
	wire n16107;
	wire n16108;
	wire n16109;
	wire n16110;
	wire n16111;
	wire n16112;
	wire n16113;
	wire n16114;
	wire n16115;
	wire n16116;
	wire n16117;
	wire n16118;
	wire n16119;
	wire n16120;
	wire n16121;
	wire n16122;
	wire n16123;
	wire n16124;
	wire n16125;
	wire n16126;
	wire n16127;
	wire n16128;
	wire n16129;
	wire n16130;
	wire n16131;
	wire n16132;
	wire n16133;
	wire n16134;
	wire n16135;
	wire n16136;
	wire n16137;
	wire n16138;
	wire n16139;
	wire n16140;
	wire n16141;
	wire n16142;
	wire n16143;
	wire n16144;
	wire n16145;
	wire n16146;
	wire n16147;
	wire n16148;
	wire n16149;
	wire n16150;
	wire n16151;
	wire n16152;
	wire n16153;
	wire n16154;
	wire n16155;
	wire n16156;
	wire n16157;
	wire n16158;
	wire n16159;
	wire n16160;
	wire n16161;
	wire n16162;
	wire n16163;
	wire n16164;
	wire n16165;
	wire n16166;
	wire n16167;
	wire n16168;
	wire n16169;
	wire n16170;
	wire n16171;
	wire n16172;
	wire n16173;
	wire n16174;
	wire n16175;
	wire n16176;
	wire n16177;
	wire n16178;
	wire n16179;
	wire n16180;
	wire n16181;
	wire n16182;
	wire n16183;
	wire n16184;
	wire n16185;
	wire n16186;
	wire n16187;
	wire n16188;
	wire n16189;
	wire n16190;
	wire n16191;
	wire n16192;
	wire n16193;
	wire n16194;
	wire n16195;
	wire n16196;
	wire n16197;
	wire n16198;
	wire n16199;
	wire n16200;
	wire n16201;
	wire n16202;
	wire n16203;
	wire n16204;
	wire n16205;
	wire n16206;
	wire n16207;
	wire n16208;
	wire n16209;
	wire n16210;
	wire n16211;
	wire n16212;
	wire n16213;
	wire n16214;
	wire n16215;
	wire n16216;
	wire n16217;
	wire n16218;
	wire n16219;
	wire n16220;
	wire n16221;
	wire n16222;
	wire n16223;
	wire n16224;
	wire n16225;
	wire n16226;
	wire n16227;
	wire n16228;
	wire n16229;
	wire n16230;
	wire n16231;
	wire n16232;
	wire n16233;
	wire n16234;
	wire n16235;
	wire n16236;
	wire n16237;
	wire n16238;
	wire n16239;
	wire n16240;
	wire n16241;
	wire n16242;
	wire n16243;
	wire n16244;
	wire n16245;
	wire n16246;
	wire n16247;
	wire n16248;
	wire n16249;
	wire n16250;
	wire n16251;
	wire n16252;
	wire n16253;
	wire n16254;
	wire n16255;
	wire n16256;
	wire n16257;
	wire n16258;
	wire n16259;
	wire n16260;
	wire n16261;
	wire n16262;
	wire n16263;
	wire n16264;
	wire n16265;
	wire n16266;
	wire n16267;
	wire n16268;
	wire n16269;
	wire n16270;
	wire n16271;
	wire n16272;
	wire n16273;
	wire n16274;
	wire n16275;
	wire n16276;
	wire n16277;
	wire n16278;
	wire n16279;
	wire n16280;
	wire n16281;
	wire n16282;
	wire n16283;
	wire n16284;
	wire n16285;
	wire n16286;
	wire n16287;
	wire n16288;
	wire n16289;
	wire n16290;
	wire n16291;
	wire n16292;
	wire n16293;
	wire n16294;
	wire n16295;
	wire n16296;
	wire n16297;
	wire n16298;
	wire n16299;
	wire n16300;
	wire n16301;
	wire n16302;
	wire n16303;
	wire n16304;
	wire n16305;
	wire n16306;
	wire n16307;
	wire n16308;
	wire n16309;
	wire n16310;
	wire n16311;
	wire n16312;
	wire n16313;
	wire n16314;
	wire n16315;
	wire n16316;
	wire n16317;
	wire n16318;
	wire n16319;
	wire n16320;
	wire n16321;
	wire n16322;
	wire n16323;
	wire n16324;
	wire n16325;
	wire n16326;
	wire n16327;
	wire n16328;
	wire n16329;
	wire n16330;
	wire n16331;
	wire n16332;
	wire n16333;
	wire n16334;
	wire n16335;
	wire n16336;
	wire n16337;
	wire n16338;
	wire n16339;
	wire n16340;
	wire n16341;
	wire n16342;
	wire n16343;
	wire n16344;
	wire n16345;
	wire n16346;
	wire n16347;
	wire n16348;
	wire n16349;
	wire n16350;
	wire n16351;
	wire n16352;
	wire n16353;
	wire n16354;
	wire n16355;
	wire n16356;
	wire n16357;
	wire n16358;
	wire n16359;
	wire n16360;
	wire n16361;
	wire n16362;
	wire n16363;
	wire n16364;
	wire n16365;
	wire n16366;
	wire n16367;
	wire n16368;
	wire n16369;
	wire n16370;
	wire n16371;
	wire n16372;
	wire n16373;
	wire n16374;
	wire n16375;
	wire n16376;
	wire n16377;
	wire n16378;
	wire n16379;
	wire n16380;
	wire n16381;
	wire n16382;
	wire n16383;
	wire n16384;
	wire n16385;
	wire n16386;
	wire n16387;
	wire n16388;
	wire n16389;
	wire n16390;
	wire n16391;
	wire n16392;
	wire n16393;
	wire n16394;
	wire n16395;
	wire n16396;
	wire n16397;
	wire n16398;
	wire n16399;
	wire n16400;
	wire n16401;
	wire n16402;
	wire n16403;
	wire n16404;
	wire n16405;
	wire n16406;
	wire n16407;
	wire n16408;
	wire n16409;
	wire n16410;
	wire n16411;
	wire n16412;
	wire n16413;
	wire n16414;
	wire n16415;
	wire n16416;
	wire n16417;
	wire n16418;
	wire n16419;
	wire n16420;
	wire n16421;
	wire n16422;
	wire n16423;
	wire n16424;
	wire n16425;
	wire n16426;
	wire n16427;
	wire n16428;
	wire n16429;
	wire n16430;
	wire n16431;
	wire n16432;
	wire n16433;
	wire n16434;
	wire n16435;
	wire n16436;
	wire n16437;
	wire n16438;
	wire n16439;
	wire n16440;
	wire n16441;
	wire n16442;
	wire n16443;
	wire n16444;
	wire n16445;
	wire n16446;
	wire n16447;
	wire n16448;
	wire n16449;
	wire n16450;
	wire n16451;
	wire n16452;
	wire n16453;
	wire n16454;
	wire n16455;
	wire n16456;
	wire n16457;
	wire n16458;
	wire n16459;
	wire n16460;
	wire n16461;
	wire n16462;
	wire n16463;
	wire n16464;
	wire n16465;
	wire n16466;
	wire n16467;
	wire n16468;
	wire n16469;
	wire n16470;
	wire n16471;
	wire n16472;
	wire n16473;
	wire n16474;
	wire n16475;
	wire n16476;
	wire n16477;
	wire n16478;
	wire n16479;
	wire n16480;
	wire n16481;
	wire n16482;
	wire n16483;
	wire n16484;
	wire n16485;
	wire n16486;
	wire n16487;
	wire n16488;
	wire n16489;
	wire n16490;
	wire n16491;
	wire n16492;
	wire n16493;
	wire n16494;
	wire n16495;
	wire n16496;
	wire n16497;
	wire n16498;
	wire n16499;
	wire n16500;
	wire n16501;
	wire n16502;
	wire n16503;
	wire n16504;
	wire n16505;
	wire n16506;
	wire n16507;
	wire n16508;
	wire n16509;
	wire n16510;
	wire n16511;
	wire n16512;
	wire n16513;
	wire n16516;
	wire n16518;
	wire n16519;
	wire n16520;
	wire n16521;
	wire n16522;
	wire n16523;
	wire n16524;
	wire n16525;
	wire n16526;
	wire n16527;
	wire n16528;
	wire n16529;
	wire n16530;
	wire n16531;
	wire n16532;
	wire n16533;
	wire n16534;
	wire n16535;
	wire n16536;
	wire n16537;
	wire n16538;
	wire n16539;
	wire n16540;
	wire n16541;
	wire n16542;
	wire n16543;
	wire n16544;
	wire n16545;
	wire n16546;
	wire n16547;
	wire n16548;
	wire n16549;
	wire n16550;
	wire n16551;
	wire n16552;
	wire n16553;
	wire n16554;
	wire n16555;
	wire n16556;
	wire n16557;
	wire n16558;
	wire n16559;
	wire n16560;
	wire n16561;
	wire n16562;
	wire n16563;
	wire n16564;
	wire n16565;
	wire n16566;
	wire n16567;
	wire n16568;
	wire n16569;
	wire n16570;
	wire n16571;
	wire n16572;
	wire n16573;
	wire n16574;
	wire n16575;
	wire n16576;
	wire n16577;
	wire n16578;
	wire n16579;
	wire n16580;
	wire n16581;
	wire n16582;
	wire n16583;
	wire n16584;
	wire n16585;
	wire n16586;
	wire n16587;
	wire n16588;
	wire n16589;
	wire n16590;
	wire n16591;
	wire n16592;
	wire n16593;
	wire n16594;
	wire n16595;
	wire n16596;
	wire n16597;
	wire n16598;
	wire n16599;
	wire n16600;
	wire n16601;
	wire n16602;
	wire n16603;
	wire n16604;
	wire n16605;
	wire n16606;
	wire n16607;
	wire n16608;
	wire n16609;
	wire n16610;
	wire n16611;
	wire n16612;
	wire n16613;
	wire n16614;
	wire n16615;
	wire n16616;
	wire n16617;
	wire n16618;
	wire n16619;
	wire n16620;
	wire n16621;
	wire n16622;
	wire n16623;
	wire n16624;
	wire n16625;
	wire n16626;
	wire n16627;
	wire n16628;
	wire n16629;
	wire n16630;
	wire n16631;
	wire n16632;
	wire n16633;
	wire n16634;
	wire n16635;
	wire n16636;
	wire n16637;
	wire n16638;
	wire n16639;
	wire n16640;
	wire n16641;
	wire n16642;
	wire n16643;
	wire n16644;
	wire n16645;
	wire n16646;
	wire n16647;
	wire n16648;
	wire n16649;
	wire n16650;
	wire n16651;
	wire n16652;
	wire n16653;
	wire n16654;
	wire n16655;
	wire n16656;
	wire n16657;
	wire n16658;
	wire n16659;
	wire n16660;
	wire n16661;
	wire n16662;
	wire n16663;
	wire n16664;
	wire n16665;
	wire n16666;
	wire n16667;
	wire n16668;
	wire n16669;
	wire n16670;
	wire n16671;
	wire n16672;
	wire n16673;
	wire n16674;
	wire n16675;
	wire n16676;
	wire n16677;
	wire n16678;
	wire n16679;
	wire n16680;
	wire n16681;
	wire n16682;
	wire n16683;
	wire n16684;
	wire n16685;
	wire n16686;
	wire n16687;
	wire n16688;
	wire n16689;
	wire n16690;
	wire n16691;
	wire n16692;
	wire n16693;
	wire n16694;
	wire n16695;
	wire n16696;
	wire n16697;
	wire n16698;
	wire n16699;
	wire n16700;
	wire n16701;
	wire n16702;
	wire n16703;
	wire n16704;
	wire n16705;
	wire n16706;
	wire n16707;
	wire n16708;
	wire n16709;
	wire n16710;
	wire n16711;
	wire n16712;
	wire n16713;
	wire n16714;
	wire n16715;
	wire n16716;
	wire n16717;
	wire n16718;
	wire n16719;
	wire n16720;
	wire n16721;
	wire n16722;
	wire n16723;
	wire n16724;
	wire n16725;
	wire n16726;
	wire n16727;
	wire n16728;
	wire n16729;
	wire n16730;
	wire n16731;
	wire n16732;
	wire n16733;
	wire n16734;
	wire n16735;
	wire n16736;
	wire n16737;
	wire n16738;
	wire n16739;
	wire n16740;
	wire n16741;
	wire n16742;
	wire n16743;
	wire n16744;
	wire n16745;
	wire n16746;
	wire n16747;
	wire n16748;
	wire n16749;
	wire n16750;
	wire n16751;
	wire n16752;
	wire n16753;
	wire n16754;
	wire n16755;
	wire n16756;
	wire n16757;
	wire n16758;
	wire n16759;
	wire n16760;
	wire n16761;
	wire n16762;
	wire n16763;
	wire n16764;
	wire n16765;
	wire n16766;
	wire n16767;
	wire n16768;
	wire n16769;
	wire n16770;
	wire n16771;
	wire n16772;
	wire n16773;
	wire n16774;
	wire n16775;
	wire n16776;
	wire n16777;
	wire n16778;
	wire n16779;
	wire n16780;
	wire n16781;
	wire n16782;
	wire n16783;
	wire n16784;
	wire n16785;
	wire n16786;
	wire n16787;
	wire n16788;
	wire n16789;
	wire n16790;
	wire n16791;
	wire n16792;
	wire n16793;
	wire n16794;
	wire n16795;
	wire n16796;
	wire n16797;
	wire n16798;
	wire n16799;
	wire n16800;
	wire n16801;
	wire n16802;
	wire n16803;
	wire n16804;
	wire n16805;
	wire n16806;
	wire n16807;
	wire n16808;
	wire n16809;
	wire n16810;
	wire n16811;
	wire n16812;
	wire n16813;
	wire n16814;
	wire n16815;
	wire n16816;
	wire n16817;
	wire n16818;
	wire n16819;
	wire n16820;
	wire n16821;
	wire n16822;
	wire n16823;
	wire n16824;
	wire n16825;
	wire n16826;
	wire n16827;
	wire n16828;
	wire n16829;
	wire n16830;
	wire n16831;
	wire n16832;
	wire n16833;
	wire n16834;
	wire n16835;
	wire n16836;
	wire n16837;
	wire n16838;
	wire n16839;
	wire n16840;
	wire n16841;
	wire n16842;
	wire n16843;
	wire n16844;
	wire n16845;
	wire n16846;
	wire n16847;
	wire n16848;
	wire n16849;
	wire n16850;
	wire n16851;
	wire n16852;
	wire n16853;
	wire n16854;
	wire n16855;
	wire n16856;
	wire n16857;
	wire n16858;
	wire n16859;
	wire n16860;
	wire n16861;
	wire n16862;
	wire n16863;
	wire n16864;
	wire n16865;
	wire n16866;
	wire n16867;
	wire n16868;
	wire n16869;
	wire n16870;
	wire n16871;
	wire n16872;
	wire n16873;
	wire n16874;
	wire n16875;
	wire n16876;
	wire n16877;
	wire n16878;
	wire n16879;
	wire n16880;
	wire n16881;
	wire n16882;
	wire n16883;
	wire n16884;
	wire n16885;
	wire n16886;
	wire n16887;
	wire n16888;
	wire n16889;
	wire n16890;
	wire n16891;
	wire n16892;
	wire n16893;
	wire n16894;
	wire n16895;
	wire n16896;
	wire n16897;
	wire n16898;
	wire n16899;
	wire n16900;
	wire n16901;
	wire n16902;
	wire n16903;
	wire n16904;
	wire n16905;
	wire n16906;
	wire n16907;
	wire n16908;
	wire n16909;
	wire n16910;
	wire n16911;
	wire n16912;
	wire n16913;
	wire n16914;
	wire n16915;
	wire n16916;
	wire n16917;
	wire n16918;
	wire n16919;
	wire n16920;
	wire n16921;
	wire n16922;
	wire n16923;
	wire n16924;
	wire n16925;
	wire n16926;
	wire n16927;
	wire n16928;
	wire n16929;
	wire n16930;
	wire n16931;
	wire n16932;
	wire n16933;
	wire n16934;
	wire n16935;
	wire n16936;
	wire n16937;
	wire n16938;
	wire n16939;
	wire n16940;
	wire n16941;
	wire n16942;
	wire n16943;
	wire n16944;
	wire n16945;
	wire n16946;
	wire n16947;
	wire n16948;
	wire n16949;
	wire n16950;
	wire n16951;
	wire n16952;
	wire n16953;
	wire n16954;
	wire n16955;
	wire n16956;
	wire n16957;
	wire n16958;
	wire n16959;
	wire n16960;
	wire n16961;
	wire n16962;
	wire n16963;
	wire n16964;
	wire n16965;
	wire n16966;
	wire n16967;
	wire n16968;
	wire n16969;
	wire n16970;
	wire n16971;
	wire n16972;
	wire n16973;
	wire n16974;
	wire n16975;
	wire n16976;
	wire n16977;
	wire n16978;
	wire n16979;
	wire n16980;
	wire n16981;
	wire n16982;
	wire n16983;
	wire n16984;
	wire n16985;
	wire n16986;
	wire n16987;
	wire n16988;
	wire n16989;
	wire n16990;
	wire n16991;
	wire n16992;
	wire n16993;
	wire n16994;
	wire n16995;
	wire n16996;
	wire n16997;
	wire n16998;
	wire n16999;
	wire n17000;
	wire n17001;
	wire n17002;
	wire n17003;
	wire n17004;
	wire n17005;
	wire n17006;
	wire n17007;
	wire n17008;
	wire n17009;
	wire n17010;
	wire n17011;
	wire n17012;
	wire n17013;
	wire n17014;
	wire n17015;
	wire n17016;
	wire n17017;
	wire n17018;
	wire n17019;
	wire n17020;
	wire n17021;
	wire n17022;
	wire n17023;
	wire n17024;
	wire n17025;
	wire n17026;
	wire n17027;
	wire n17028;
	wire n17029;
	wire n17030;
	wire n17031;
	wire n17032;
	wire n17033;
	wire n17034;
	wire n17035;
	wire n17036;
	wire n17037;
	wire n17038;
	wire n17039;
	wire n17040;
	wire n17041;
	wire n17042;
	wire n17043;
	wire n17044;
	wire n17045;
	wire n17046;
	wire n17047;
	wire n17048;
	wire n17049;
	wire n17050;
	wire n17051;
	wire n17052;
	wire n17053;
	wire n17054;
	wire n17055;
	wire n17056;
	wire n17057;
	wire n17058;
	wire n17059;
	wire n17060;
	wire n17061;
	wire n17062;
	wire n17063;
	wire n17064;
	wire n17065;
	wire n17066;
	wire n17067;
	wire n17068;
	wire n17069;
	wire n17070;
	wire n17071;
	wire n17072;
	wire n17073;
	wire n17074;
	wire n17075;
	wire n17076;
	wire n17077;
	wire n17078;
	wire n17079;
	wire n17080;
	wire n17081;
	wire n17082;
	wire n17083;
	wire n17084;
	wire n17085;
	wire n17086;
	wire n17087;
	wire n17088;
	wire n17089;
	wire n17090;
	wire n17091;
	wire n17092;
	wire n17093;
	wire n17094;
	wire n17095;
	wire n17096;
	wire n17097;
	wire n17098;
	wire n17099;
	wire n17100;
	wire n17101;
	wire n17102;
	wire n17103;
	wire n17104;
	wire n17105;
	wire n17106;
	wire n17107;
	wire n17108;
	wire n17109;
	wire n17110;
	wire n17111;
	wire n17112;
	wire n17113;
	wire n17114;
	wire n17115;
	wire n17116;
	wire n17117;
	wire n17118;
	wire n17119;
	wire n17120;
	wire n17121;
	wire n17122;
	wire n17123;
	wire n17124;
	wire n17125;
	wire n17126;
	wire n17127;
	wire n17128;
	wire n17129;
	wire n17130;
	wire n17131;
	wire n17132;
	wire n17133;
	wire n17134;
	wire n17135;
	wire n17138;
	wire n17139;
	wire n17140;
	wire n17141;
	wire n17142;
	wire n17143;
	wire n17144;
	wire n17145;
	wire n17146;
	wire n17147;
	wire n17148;
	wire n17149;
	wire n17150;
	wire n17151;
	wire n17152;
	wire n17153;
	wire n17154;
	wire n17155;
	wire n17156;
	wire n17157;
	wire n17158;
	wire n17159;
	wire n17160;
	wire n17161;
	wire n17162;
	wire n17163;
	wire n17164;
	wire n17165;
	wire n17166;
	wire n17167;
	wire n17168;
	wire n17169;
	wire n17170;
	wire n17171;
	wire n17172;
	wire n17173;
	wire n17174;
	wire n17175;
	wire n17176;
	wire n17177;
	wire n17178;
	wire n17179;
	wire n17180;
	wire n17181;
	wire n17182;
	wire n17183;
	wire n17184;
	wire n17185;
	wire n17186;
	wire n17187;
	wire n17188;
	wire n17189;
	wire n17190;
	wire n17191;
	wire n17192;
	wire n17193;
	wire n17194;
	wire n17195;
	wire n17196;
	wire n17197;
	wire n17199;
	wire n17200;
	wire n17201;
	wire n17202;
	wire n17203;
	wire n17204;
	wire n17205;
	wire n17206;
	wire n17207;
	wire n17208;
	wire n17209;
	wire n17210;
	wire n17211;
	wire n17212;
	wire n17213;
	wire n17214;
	wire n17215;
	wire n17216;
	wire n17217;
	wire n17218;
	wire n17219;
	wire n17220;
	wire n17221;
	wire n17222;
	wire n17223;
	wire n17224;
	wire n17225;
	wire n17226;
	wire n17227;
	wire n17228;
	wire n17229;
	wire n17230;
	wire n17231;
	wire n17232;
	wire n17233;
	wire n17234;
	wire n17235;
	wire n17236;
	wire n17237;
	wire n17238;
	wire n17239;
	wire n17240;
	wire n17241;
	wire n17242;
	wire n17243;
	wire n17244;
	wire n17245;
	wire n17246;
	wire n17247;
	wire n17248;
	wire n17249;
	wire n17250;
	wire n17251;
	wire n17252;
	wire n17253;
	wire n17254;
	wire n17255;
	wire n17256;
	wire n17257;
	wire n17258;
	wire n17259;
	wire n17260;
	wire n17261;
	wire n17262;
	wire n17263;
	wire n17264;
	wire n17265;
	wire n17266;
	wire n17267;
	wire n17268;
	wire n17269;
	wire n17270;
	wire n17271;
	wire n17272;
	wire n17273;
	wire n17274;
	wire n17275;
	wire n17276;
	wire n17277;
	wire n17278;
	wire n17279;
	wire n17280;
	wire n17281;
	wire n17282;
	wire n17283;
	wire n17284;
	wire n17285;
	wire n17286;
	wire n17287;
	wire n17288;
	wire n17289;
	wire n17290;
	wire n17291;
	wire n17292;
	wire n17293;
	wire n17294;
	wire n17295;
	wire n17296;
	wire n17297;
	wire n17298;
	wire n17299;
	wire n17300;
	wire n17301;
	wire n17302;
	wire n17303;
	wire n17304;
	wire n17305;
	wire n17306;
	wire n17307;
	wire n17308;
	wire n17309;
	wire n17310;
	wire n17311;
	wire n17312;
	wire n17313;
	wire n17314;
	wire n17315;
	wire n17316;
	wire n17317;
	wire n17318;
	wire n17319;
	wire n17320;
	wire n17321;
	wire n17322;
	wire n17323;
	wire n17324;
	wire n17325;
	wire n17326;
	wire n17327;
	wire n17328;
	wire n17329;
	wire n17330;
	wire n17331;
	wire n17332;
	wire n17333;
	wire n17334;
	wire n17335;
	wire n17336;
	wire n17337;
	wire n17338;
	wire n17339;
	wire n17340;
	wire n17341;
	wire n17342;
	wire n17343;
	wire n17344;
	wire n17345;
	wire n17346;
	wire n17347;
	wire n17348;
	wire n17349;
	wire n17350;
	wire n17351;
	wire n17352;
	wire n17353;
	wire n17354;
	wire n17355;
	wire n17356;
	wire n17357;
	wire n17358;
	wire n17359;
	wire n17360;
	wire n17361;
	wire n17362;
	wire n17363;
	wire n17364;
	wire n17365;
	wire n17366;
	wire n17367;
	wire n17368;
	wire n17369;
	wire n17370;
	wire n17371;
	wire n17372;
	wire n17373;
	wire n17374;
	wire n17375;
	wire n17376;
	wire n17377;
	wire n17378;
	wire n17379;
	wire n17380;
	wire n17381;
	wire n17382;
	wire n17383;
	wire n17384;
	wire n17385;
	wire n17386;
	wire n17387;
	wire n17388;
	wire n17389;
	wire n17390;
	wire n17391;
	wire n17392;
	wire n17393;
	wire n17394;
	wire n17395;
	wire n17396;
	wire n17397;
	wire n17398;
	wire n17399;
	wire n17400;
	wire n17401;
	wire n17402;
	wire n17403;
	wire n17404;
	wire n17405;
	wire n17406;
	wire n17407;
	wire n17408;
	wire n17409;
	wire n17410;
	wire n17411;
	wire n17412;
	wire n17413;
	wire n17414;
	wire n17415;
	wire n17416;
	wire n17417;
	wire n17418;
	wire n17419;
	wire n17420;
	wire n17421;
	wire n17422;
	wire n17423;
	wire n17424;
	wire n17425;
	wire n17426;
	wire n17427;
	wire n17428;
	wire n17429;
	wire n17430;
	wire n17431;
	wire n17432;
	wire n17433;
	wire n17434;
	wire n17435;
	wire n17436;
	wire n17437;
	wire n17438;
	wire n17439;
	wire n17440;
	wire n17441;
	wire n17442;
	wire n17443;
	wire n17444;
	wire n17445;
	wire n17446;
	wire n17447;
	wire n17448;
	wire n17449;
	wire n17450;
	wire n17451;
	wire n17452;
	wire n17453;
	wire n17454;
	wire n17455;
	wire n17456;
	wire n17457;
	wire n17458;
	wire n17459;
	wire n17460;
	wire n17461;
	wire n17462;
	wire n17463;
	wire n17464;
	wire n17465;
	wire n17466;
	wire n17467;
	wire n17468;
	wire n17469;
	wire n17470;
	wire n17471;
	wire n17472;
	wire n17473;
	wire n17474;
	wire n17475;
	wire n17476;
	wire n17477;
	wire n17478;
	wire n17479;
	wire n17480;
	wire n17481;
	wire n17482;
	wire n17483;
	wire n17484;
	wire n17485;
	wire n17486;
	wire n17487;
	wire n17488;
	wire n17489;
	wire n17490;
	wire n17491;
	wire n17492;
	wire n17493;
	wire n17494;
	wire n17495;
	wire n17496;
	wire n17497;
	wire n17498;
	wire n17499;
	wire n17500;
	wire n17501;
	wire n17502;
	wire n17503;
	wire n17504;
	wire n17505;
	wire n17506;
	wire n17507;
	wire n17508;
	wire n17509;
	wire n17510;
	wire n17511;
	wire n17512;
	wire n17513;
	wire n17514;
	wire n17515;
	wire n17516;
	wire n17517;
	wire n17518;
	wire n17519;
	wire n17520;
	wire n17521;
	wire n17522;
	wire n17523;
	wire n17524;
	wire n17525;
	wire n17526;
	wire n17527;
	wire n17528;
	wire n17529;
	wire n17530;
	wire n17531;
	wire n17532;
	wire n17533;
	wire n17534;
	wire n17535;
	wire n17536;
	wire n17537;
	wire n17538;
	wire n17539;
	wire n17540;
	wire n17541;
	wire n17542;
	wire n17543;
	wire n17544;
	wire n17545;
	wire n17546;
	wire n17547;
	wire n17548;
	wire n17549;
	wire n17550;
	wire n17551;
	wire n17552;
	wire n17553;
	wire n17554;
	wire n17555;
	wire n17556;
	wire n17557;
	wire n17558;
	wire n17559;
	wire n17560;
	wire n17561;
	wire n17562;
	wire n17563;
	wire n17564;
	wire n17565;
	wire n17566;
	wire n17567;
	wire n17568;
	wire n17569;
	wire n17570;
	wire n17571;
	wire n17572;
	wire n17573;
	wire n17574;
	wire n17575;
	wire n17576;
	wire n17577;
	wire n17578;
	wire n17579;
	wire n17580;
	wire n17581;
	wire n17582;
	wire n17583;
	wire n17584;
	wire n17585;
	wire n17586;
	wire n17587;
	wire n17588;
	wire n17589;
	wire n17590;
	wire n17591;
	wire n17592;
	wire n17593;
	wire n17594;
	wire n17595;
	wire n17596;
	wire n17597;
	wire n17598;
	wire n17599;
	wire n17600;
	wire n17601;
	wire n17602;
	wire n17603;
	wire n17604;
	wire n17605;
	wire n17606;
	wire n17607;
	wire n17608;
	wire n17609;
	wire n17610;
	wire n17611;
	wire n17612;
	wire n17613;
	wire n17614;
	wire n17615;
	wire n17616;
	wire n17617;
	wire n17618;
	wire n17619;
	wire n17620;
	wire n17621;
	wire n17622;
	wire n17623;
	wire n17624;
	wire n17625;
	wire n17626;
	wire n17627;
	wire n17628;
	wire n17629;
	wire n17630;
	wire n17631;
	wire n17632;
	wire n17633;
	wire n17634;
	wire n17635;
	wire n17636;
	wire n17637;
	wire n17638;
	wire n17639;
	wire n17640;
	wire n17641;
	wire n17642;
	wire n17643;
	wire n17644;
	wire n17645;
	wire n17646;
	wire n17647;
	wire n17648;
	wire n17649;
	wire n17650;
	wire n17651;
	wire n17652;
	wire n17653;
	wire n17654;
	wire n17655;
	wire n17656;
	wire n17657;
	wire n17658;
	wire n17659;
	wire n17660;
	wire n17661;
	wire n17662;
	wire n17663;
	wire n17664;
	wire n17665;
	wire n17666;
	wire n17667;
	wire n17668;
	wire n17669;
	wire n17670;
	wire n17671;
	wire n17672;
	wire n17673;
	wire n17674;
	wire n17675;
	wire n17676;
	wire n17677;
	wire n17678;
	wire n17679;
	wire n17680;
	wire n17681;
	wire n17682;
	wire n17683;
	wire n17684;
	wire n17685;
	wire n17686;
	wire n17687;
	wire n17688;
	wire n17689;
	wire n17690;
	wire n17691;
	wire n17692;
	wire n17693;
	wire n17694;
	wire n17695;
	wire n17696;
	wire n17697;
	wire n17698;
	wire n17699;
	wire n17700;
	wire n17701;
	wire n17702;
	wire n17703;
	wire n17704;
	wire n17705;
	wire n17706;
	wire n17707;
	wire n17708;
	wire n17709;
	wire n17710;
	wire n17711;
	wire n17712;
	wire n17713;
	wire n17716;
	wire n17718;
	wire n17719;
	wire n17720;
	wire n17721;
	wire n17722;
	wire n17723;
	wire n17724;
	wire n17725;
	wire n17726;
	wire n17727;
	wire n17728;
	wire n17729;
	wire n17730;
	wire n17731;
	wire n17732;
	wire n17733;
	wire n17734;
	wire n17735;
	wire n17736;
	wire n17737;
	wire n17738;
	wire n17739;
	wire n17740;
	wire n17741;
	wire n17742;
	wire n17743;
	wire n17744;
	wire n17745;
	wire n17746;
	wire n17747;
	wire n17748;
	wire n17749;
	wire n17750;
	wire n17751;
	wire n17752;
	wire n17753;
	wire n17754;
	wire n17755;
	wire n17756;
	wire n17757;
	wire n17758;
	wire n17759;
	wire n17760;
	wire n17761;
	wire n17762;
	wire n17763;
	wire n17764;
	wire n17765;
	wire n17766;
	wire n17767;
	wire n17768;
	wire n17769;
	wire n17770;
	wire n17771;
	wire n17772;
	wire n17773;
	wire n17774;
	wire n17775;
	wire n17776;
	wire n17777;
	wire n17778;
	wire n17779;
	wire n17780;
	wire n17781;
	wire n17782;
	wire n17783;
	wire n17784;
	wire n17785;
	wire n17786;
	wire n17787;
	wire n17788;
	wire n17789;
	wire n17790;
	wire n17791;
	wire n17792;
	wire n17793;
	wire n17794;
	wire n17795;
	wire n17796;
	wire n17797;
	wire n17798;
	wire n17799;
	wire n17800;
	wire n17801;
	wire n17802;
	wire n17803;
	wire n17804;
	wire n17805;
	wire n17806;
	wire n17807;
	wire n17808;
	wire n17809;
	wire n17810;
	wire n17811;
	wire n17812;
	wire n17813;
	wire n17814;
	wire n17815;
	wire n17816;
	wire n17817;
	wire n17818;
	wire n17819;
	wire n17820;
	wire n17821;
	wire n17822;
	wire n17823;
	wire n17824;
	wire n17825;
	wire n17826;
	wire n17827;
	wire n17828;
	wire n17829;
	wire n17830;
	wire n17831;
	wire n17832;
	wire n17833;
	wire n17834;
	wire n17835;
	wire n17836;
	wire n17837;
	wire n17838;
	wire n17839;
	wire n17840;
	wire n17841;
	wire n17842;
	wire n17843;
	wire n17844;
	wire n17845;
	wire n17846;
	wire n17847;
	wire n17848;
	wire n17849;
	wire n17850;
	wire n17851;
	wire n17852;
	wire n17853;
	wire n17854;
	wire n17855;
	wire n17856;
	wire n17857;
	wire n17858;
	wire n17859;
	wire n17860;
	wire n17861;
	wire n17862;
	wire n17863;
	wire n17864;
	wire n17865;
	wire n17866;
	wire n17867;
	wire n17868;
	wire n17869;
	wire n17870;
	wire n17871;
	wire n17872;
	wire n17873;
	wire n17874;
	wire n17875;
	wire n17876;
	wire n17877;
	wire n17878;
	wire n17879;
	wire n17880;
	wire n17881;
	wire n17882;
	wire n17883;
	wire n17884;
	wire n17885;
	wire n17886;
	wire n17887;
	wire n17888;
	wire n17889;
	wire n17890;
	wire n17891;
	wire n17892;
	wire n17893;
	wire n17894;
	wire n17895;
	wire n17896;
	wire n17897;
	wire n17898;
	wire n17899;
	wire n17900;
	wire n17901;
	wire n17902;
	wire n17903;
	wire n17904;
	wire n17905;
	wire n17906;
	wire n17907;
	wire n17908;
	wire n17909;
	wire n17910;
	wire n17911;
	wire n17912;
	wire n17913;
	wire n17914;
	wire n17915;
	wire n17916;
	wire n17917;
	wire n17918;
	wire n17919;
	wire n17920;
	wire n17921;
	wire n17922;
	wire n17923;
	wire n17924;
	wire n17925;
	wire n17926;
	wire n17927;
	wire n17928;
	wire n17929;
	wire n17930;
	wire n17931;
	wire n17932;
	wire n17933;
	wire n17934;
	wire n17935;
	wire n17936;
	wire n17937;
	wire n17938;
	wire n17939;
	wire n17940;
	wire n17941;
	wire n17942;
	wire n17943;
	wire n17944;
	wire n17945;
	wire n17946;
	wire n17947;
	wire n17948;
	wire n17949;
	wire n17950;
	wire n17951;
	wire n17952;
	wire n17953;
	wire n17954;
	wire n17955;
	wire n17956;
	wire n17957;
	wire n17958;
	wire n17959;
	wire n17960;
	wire n17961;
	wire n17962;
	wire n17963;
	wire n17964;
	wire n17965;
	wire n17966;
	wire n17967;
	wire n17968;
	wire n17969;
	wire n17970;
	wire n17971;
	wire n17972;
	wire n17973;
	wire n17974;
	wire n17975;
	wire n17976;
	wire n17977;
	wire n17978;
	wire n17979;
	wire n17980;
	wire n17981;
	wire n17982;
	wire n17983;
	wire n17984;
	wire n17985;
	wire n17986;
	wire n17987;
	wire n17988;
	wire n17989;
	wire n17990;
	wire n17991;
	wire n17992;
	wire n17993;
	wire n17994;
	wire n17995;
	wire n17996;
	wire n17997;
	wire n17998;
	wire n17999;
	wire n18000;
	wire n18001;
	wire n18002;
	wire n18003;
	wire n18004;
	wire n18005;
	wire n18006;
	wire n18007;
	wire n18008;
	wire n18009;
	wire n18010;
	wire n18011;
	wire n18012;
	wire n18013;
	wire n18014;
	wire n18015;
	wire n18016;
	wire n18017;
	wire n18018;
	wire n18019;
	wire n18020;
	wire n18021;
	wire n18022;
	wire n18023;
	wire n18024;
	wire n18025;
	wire n18026;
	wire n18027;
	wire n18028;
	wire n18029;
	wire n18030;
	wire n18031;
	wire n18032;
	wire n18033;
	wire n18034;
	wire n18035;
	wire n18036;
	wire n18037;
	wire n18038;
	wire n18039;
	wire n18040;
	wire n18041;
	wire n18042;
	wire n18043;
	wire n18044;
	wire n18045;
	wire n18046;
	wire n18047;
	wire n18048;
	wire n18049;
	wire n18050;
	wire n18051;
	wire n18052;
	wire n18053;
	wire n18054;
	wire n18055;
	wire n18056;
	wire n18057;
	wire n18058;
	wire n18059;
	wire n18060;
	wire n18061;
	wire n18062;
	wire n18063;
	wire n18064;
	wire n18065;
	wire n18066;
	wire n18067;
	wire n18068;
	wire n18069;
	wire n18070;
	wire n18071;
	wire n18072;
	wire n18073;
	wire n18074;
	wire n18075;
	wire n18076;
	wire n18077;
	wire n18078;
	wire n18079;
	wire n18080;
	wire n18081;
	wire n18082;
	wire n18083;
	wire n18084;
	wire n18085;
	wire n18086;
	wire n18087;
	wire n18088;
	wire n18089;
	wire n18090;
	wire n18091;
	wire n18092;
	wire n18093;
	wire n18094;
	wire n18095;
	wire n18096;
	wire n18097;
	wire n18098;
	wire n18099;
	wire n18100;
	wire n18101;
	wire n18102;
	wire n18103;
	wire n18104;
	wire n18105;
	wire n18106;
	wire n18107;
	wire n18108;
	wire n18109;
	wire n18110;
	wire n18111;
	wire n18112;
	wire n18113;
	wire n18114;
	wire n18115;
	wire n18116;
	wire n18117;
	wire n18118;
	wire n18119;
	wire n18120;
	wire n18121;
	wire n18122;
	wire n18123;
	wire n18124;
	wire n18125;
	wire n18126;
	wire n18127;
	wire n18128;
	wire n18129;
	wire n18130;
	wire n18131;
	wire n18132;
	wire n18133;
	wire n18134;
	wire n18135;
	wire n18136;
	wire n18137;
	wire n18138;
	wire n18139;
	wire n18140;
	wire n18141;
	wire n18142;
	wire n18143;
	wire n18144;
	wire n18145;
	wire n18146;
	wire n18147;
	wire n18148;
	wire n18149;
	wire n18150;
	wire n18151;
	wire n18152;
	wire n18153;
	wire n18154;
	wire n18155;
	wire n18156;
	wire n18157;
	wire n18158;
	wire n18159;
	wire n18160;
	wire n18161;
	wire n18162;
	wire n18163;
	wire n18164;
	wire n18165;
	wire n18166;
	wire n18167;
	wire n18168;
	wire n18169;
	wire n18170;
	wire n18171;
	wire n18172;
	wire n18173;
	wire n18174;
	wire n18175;
	wire n18176;
	wire n18177;
	wire n18178;
	wire n18179;
	wire n18180;
	wire n18181;
	wire n18182;
	wire n18183;
	wire n18184;
	wire n18185;
	wire n18186;
	wire n18187;
	wire n18188;
	wire n18189;
	wire n18190;
	wire n18191;
	wire n18192;
	wire n18193;
	wire n18194;
	wire n18195;
	wire n18196;
	wire n18197;
	wire n18198;
	wire n18199;
	wire n18200;
	wire n18201;
	wire n18202;
	wire n18203;
	wire n18204;
	wire n18205;
	wire n18206;
	wire n18207;
	wire n18208;
	wire n18209;
	wire n18210;
	wire n18211;
	wire n18212;
	wire n18213;
	wire n18214;
	wire n18215;
	wire n18216;
	wire n18217;
	wire n18218;
	wire n18219;
	wire n18220;
	wire n18221;
	wire n18222;
	wire n18223;
	wire n18224;
	wire n18225;
	wire n18226;
	wire n18227;
	wire n18228;
	wire n18229;
	wire n18230;
	wire n18231;
	wire n18232;
	wire n18233;
	wire n18234;
	wire n18235;
	wire n18236;
	wire n18237;
	wire n18238;
	wire n18239;
	wire n18240;
	wire n18241;
	wire n18242;
	wire n18243;
	wire n18244;
	wire n18245;
	wire n18246;
	wire n18247;
	wire n18248;
	wire n18249;
	wire n18250;
	wire n18251;
	wire n18252;
	wire n18253;
	wire n18254;
	wire n18255;
	wire n18256;
	wire n18257;
	wire n18258;
	wire n18259;
	wire n18260;
	wire n18261;
	wire n18262;
	wire n18263;
	wire n18264;
	wire n18265;
	wire n18266;
	wire n18267;
	wire n18268;
	wire n18269;
	wire n18270;
	wire n18271;
	wire n18272;
	wire n18273;
	wire n18274;
	wire n18275;
	wire n18276;
	wire n18277;
	wire n18278;
	wire n18279;
	wire n18280;
	wire n18281;
	wire n18282;
	wire n18283;
	wire n18284;
	wire n18285;
	wire n18286;
	wire n18287;
	wire n18288;
	wire n18289;
	wire n18290;
	wire n18291;
	wire n18292;
	wire n18293;
	wire n18294;
	wire n18295;
	wire n18296;
	wire n18297;
	wire n18298;
	wire n18299;
	wire n18300;
	wire n18301;
	wire n18302;
	wire n18303;
	wire n18304;
	wire n18305;
	wire n18306;
	wire n18307;
	wire n18308;
	wire n18309;
	wire n18310;
	wire n18311;
	wire n18312;
	wire n18313;
	wire n18314;
	wire n18315;
	wire n18316;
	wire n18317;
	wire n18318;
	wire n18319;
	wire n18320;
	wire n18321;
	wire n18322;
	wire n18323;
	wire n18324;
	wire n18325;
	wire n18326;
	wire n18327;
	wire n18328;
	wire n18329;
	wire n18330;
	wire n18331;
	wire n18332;
	wire n18333;
	wire n18334;
	wire n18335;
	wire n18336;
	wire n18337;
	wire n18338;
	wire n18339;
	wire n18340;
	wire n18341;
	wire n18342;
	wire n18343;
	wire n18344;
	wire n18345;
	wire n18346;
	wire n18347;
	wire n18348;
	wire n18349;
	wire n18350;
	wire n18351;
	wire n18352;
	wire n18353;
	wire n18354;
	wire n18355;
	wire n18356;
	wire n18357;
	wire n18358;
	wire n18359;
	wire n18360;
	wire n18361;
	wire n18362;
	wire n18363;
	wire n18364;
	wire n18365;
	wire n18366;
	wire n18367;
	wire n18368;
	wire n18369;
	wire n18370;
	wire n18371;
	wire n18372;
	wire n18373;
	wire n18374;
	wire n18375;
	wire n18376;
	wire n18377;
	wire n18379;
	wire n18380;
	wire n18381;
	wire n18382;
	wire n18383;
	wire n18384;
	wire n18385;
	wire n18386;
	wire n18387;
	wire n18388;
	wire n18389;
	wire n18390;
	wire n18391;
	wire n18392;
	wire n18393;
	wire n18394;
	wire n18395;
	wire n18396;
	wire n18397;
	wire n18398;
	wire n18399;
	wire n18400;
	wire n18401;
	wire n18402;
	wire n18403;
	wire n18404;
	wire n18405;
	wire n18406;
	wire n18407;
	wire n18408;
	wire n18409;
	wire n18410;
	wire n18411;
	wire n18412;
	wire n18413;
	wire n18414;
	wire n18415;
	wire n18416;
	wire n18417;
	wire n18418;
	wire n18419;
	wire n18420;
	wire n18421;
	wire n18422;
	wire n18423;
	wire n18424;
	wire n18425;
	wire n18426;
	wire n18427;
	wire n18428;
	wire n18429;
	wire n18430;
	wire n18431;
	wire n18432;
	wire n18433;
	wire n18434;
	wire n18435;
	wire n18436;
	wire n18437;
	wire n18438;
	wire n18439;
	wire n18440;
	wire n18441;
	wire n18442;
	wire n18443;
	wire n18444;
	wire n18445;
	wire n18446;
	wire n18447;
	wire n18448;
	wire n18449;
	wire n18450;
	wire n18451;
	wire n18452;
	wire n18453;
	wire n18454;
	wire n18455;
	wire n18456;
	wire n18457;
	wire n18458;
	wire n18459;
	wire n18460;
	wire n18461;
	wire n18462;
	wire n18463;
	wire n18464;
	wire n18465;
	wire n18466;
	wire n18467;
	wire n18468;
	wire n18469;
	wire n18470;
	wire n18471;
	wire n18472;
	wire n18473;
	wire n18474;
	wire n18475;
	wire n18476;
	wire n18477;
	wire n18478;
	wire n18479;
	wire n18480;
	wire n18481;
	wire n18482;
	wire n18483;
	wire n18484;
	wire n18485;
	wire n18486;
	wire n18487;
	wire n18488;
	wire n18489;
	wire n18490;
	wire n18491;
	wire n18492;
	wire n18493;
	wire n18494;
	wire n18495;
	wire n18496;
	wire n18497;
	wire n18498;
	wire n18499;
	wire n18500;
	wire n18501;
	wire n18502;
	wire n18503;
	wire n18504;
	wire n18505;
	wire n18506;
	wire n18507;
	wire n18508;
	wire n18509;
	wire n18510;
	wire n18511;
	wire n18512;
	wire n18513;
	wire n18514;
	wire n18515;
	wire n18516;
	wire n18517;
	wire n18518;
	wire n18519;
	wire n18520;
	wire n18521;
	wire n18522;
	wire n18523;
	wire n18524;
	wire n18525;
	wire n18526;
	wire n18527;
	wire n18528;
	wire n18529;
	wire n18530;
	wire n18531;
	wire n18532;
	wire n18533;
	wire n18534;
	wire n18535;
	wire n18536;
	wire n18537;
	wire n18538;
	wire n18539;
	wire n18540;
	wire n18541;
	wire n18542;
	wire n18543;
	wire n18544;
	wire n18545;
	wire n18546;
	wire n18547;
	wire n18548;
	wire n18549;
	wire n18550;
	wire n18551;
	wire n18552;
	wire n18553;
	wire n18554;
	wire n18555;
	wire n18556;
	wire n18557;
	wire n18558;
	wire n18559;
	wire n18560;
	wire n18561;
	wire n18562;
	wire n18563;
	wire n18564;
	wire n18565;
	wire n18566;
	wire n18567;
	wire n18568;
	wire n18569;
	wire n18570;
	wire n18571;
	wire n18572;
	wire n18573;
	wire n18574;
	wire n18575;
	wire n18576;
	wire n18577;
	wire n18578;
	wire n18579;
	wire n18580;
	wire n18581;
	wire n18582;
	wire n18583;
	wire n18584;
	wire n18585;
	wire n18586;
	wire n18587;
	wire n18588;
	wire n18589;
	wire n18590;
	wire n18591;
	wire n18592;
	wire n18593;
	wire n18594;
	wire n18595;
	wire n18596;
	wire n18597;
	wire n18598;
	wire n18599;
	wire n18600;
	wire n18601;
	wire n18602;
	wire n18603;
	wire n18604;
	wire n18605;
	wire n18606;
	wire n18607;
	wire n18608;
	wire n18609;
	wire n18610;
	wire n18611;
	wire n18612;
	wire n18613;
	wire n18614;
	wire n18615;
	wire n18616;
	wire n18617;
	wire n18618;
	wire n18619;
	wire n18620;
	wire n18621;
	wire n18622;
	wire n18623;
	wire n18624;
	wire n18625;
	wire n18626;
	wire n18627;
	wire n18628;
	wire n18629;
	wire n18630;
	wire n18631;
	wire n18632;
	wire n18633;
	wire n18634;
	wire n18635;
	wire n18636;
	wire n18637;
	wire n18638;
	wire n18639;
	wire n18640;
	wire n18641;
	wire n18642;
	wire n18643;
	wire n18644;
	wire n18645;
	wire n18646;
	wire n18647;
	wire n18648;
	wire n18649;
	wire n18650;
	wire n18651;
	wire n18652;
	wire n18653;
	wire n18654;
	wire n18655;
	wire n18656;
	wire n18657;
	wire n18658;
	wire n18659;
	wire n18660;
	wire n18661;
	wire n18662;
	wire n18663;
	wire n18664;
	wire n18665;
	wire n18666;
	wire n18667;
	wire n18668;
	wire n18669;
	wire n18670;
	wire n18671;
	wire n18672;
	wire n18673;
	wire n18674;
	wire n18675;
	wire n18676;
	wire n18677;
	wire n18678;
	wire n18679;
	wire n18680;
	wire n18681;
	wire n18682;
	wire n18683;
	wire n18684;
	wire n18685;
	wire n18686;
	wire n18687;
	wire n18688;
	wire n18689;
	wire n18690;
	wire n18691;
	wire n18692;
	wire n18693;
	wire n18694;
	wire n18695;
	wire n18696;
	wire n18697;
	wire n18698;
	wire n18699;
	wire n18700;
	wire n18701;
	wire n18702;
	wire n18703;
	wire n18704;
	wire n18705;
	wire n18706;
	wire n18707;
	wire n18708;
	wire n18709;
	wire n18710;
	wire n18711;
	wire n18712;
	wire n18713;
	wire n18714;
	wire n18715;
	wire n18716;
	wire n18717;
	wire n18718;
	wire n18719;
	wire n18720;
	wire n18721;
	wire n18722;
	wire n18723;
	wire n18724;
	wire n18725;
	wire n18726;
	wire n18727;
	wire n18728;
	wire n18729;
	wire n18730;
	wire n18731;
	wire n18732;
	wire n18733;
	wire n18734;
	wire n18735;
	wire n18736;
	wire n18737;
	wire n18738;
	wire n18739;
	wire n18740;
	wire n18741;
	wire n18742;
	wire n18743;
	wire n18744;
	wire n18745;
	wire n18746;
	wire n18747;
	wire n18748;
	wire n18749;
	wire n18750;
	wire n18751;
	wire n18752;
	wire n18753;
	wire n18754;
	wire n18755;
	wire n18756;
	wire n18757;
	wire n18758;
	wire n18759;
	wire n18760;
	wire n18761;
	wire n18762;
	wire n18763;
	wire n18764;
	wire n18765;
	wire n18766;
	wire n18767;
	wire n18768;
	wire n18769;
	wire n18770;
	wire n18771;
	wire n18772;
	wire n18773;
	wire n18774;
	wire n18775;
	wire n18776;
	wire n18777;
	wire n18778;
	wire n18779;
	wire n18780;
	wire n18781;
	wire n18782;
	wire n18783;
	wire n18784;
	wire n18785;
	wire n18786;
	wire n18787;
	wire n18788;
	wire n18789;
	wire n18790;
	wire n18791;
	wire n18792;
	wire n18793;
	wire n18794;
	wire n18795;
	wire n18796;
	wire n18797;
	wire n18798;
	wire n18799;
	wire n18800;
	wire n18801;
	wire n18802;
	wire n18803;
	wire n18804;
	wire n18805;
	wire n18806;
	wire n18807;
	wire n18808;
	wire n18809;
	wire n18810;
	wire n18811;
	wire n18812;
	wire n18813;
	wire n18814;
	wire n18815;
	wire n18816;
	wire n18817;
	wire n18818;
	wire n18819;
	wire n18820;
	wire n18821;
	wire n18822;
	wire n18823;
	wire n18824;
	wire n18825;
	wire n18826;
	wire n18827;
	wire n18828;
	wire n18829;
	wire n18830;
	wire n18831;
	wire n18832;
	wire n18833;
	wire n18834;
	wire n18835;
	wire n18836;
	wire n18837;
	wire n18838;
	wire n18839;
	wire n18840;
	wire n18841;
	wire n18842;
	wire n18843;
	wire n18844;
	wire n18845;
	wire n18846;
	wire n18847;
	wire n18848;
	wire n18849;
	wire n18850;
	wire n18851;
	wire n18852;
	wire n18853;
	wire n18854;
	wire n18855;
	wire n18856;
	wire n18857;
	wire n18858;
	wire n18859;
	wire n18860;
	wire n18861;
	wire n18862;
	wire n18863;
	wire n18864;
	wire n18865;
	wire n18866;
	wire n18867;
	wire n18868;
	wire n18869;
	wire n18870;
	wire n18871;
	wire n18872;
	wire n18873;
	wire n18874;
	wire n18875;
	wire n18876;
	wire n18877;
	wire n18878;
	wire n18879;
	wire n18880;
	wire n18881;
	wire n18882;
	wire n18883;
	wire n18884;
	wire n18885;
	wire n18886;
	wire n18887;
	wire n18888;
	wire n18889;
	wire n18890;
	wire n18891;
	wire n18892;
	wire n18893;
	wire n18894;
	wire n18895;
	wire n18896;
	wire n18897;
	wire n18898;
	wire n18899;
	wire n18900;
	wire n18901;
	wire n18902;
	wire n18903;
	wire n18904;
	wire n18905;
	wire n18906;
	wire n18907;
	wire n18908;
	wire n18909;
	wire n18910;
	wire n18911;
	wire n18912;
	wire n18913;
	wire n18914;
	wire n18915;
	wire n18916;
	wire n18917;
	wire n18918;
	wire n18919;
	wire n18920;
	wire n18921;
	wire n18922;
	wire n18923;
	wire n18924;
	wire n18925;
	wire n18926;
	wire n18927;
	wire n18928;
	wire n18929;
	wire n18930;
	wire n18931;
	wire n18932;
	wire n18933;
	wire n18934;
	wire n18935;
	wire n18936;
	wire n18937;
	wire n18938;
	wire n18939;
	wire n18940;
	wire n18941;
	wire n18942;
	wire n18943;
	wire n18944;
	wire n18945;
	wire n18946;
	wire n18947;
	wire n18948;
	wire n18949;
	wire n18950;
	wire n18951;
	wire n18952;
	wire n18953;
	wire n18954;
	wire n18956;
	wire n18957;
	wire n18958;
	wire n18959;
	wire n18960;
	wire n18961;
	wire n18962;
	wire n18963;
	wire n18964;
	wire n18965;
	wire n18966;
	wire n18967;
	wire n18968;
	wire n18969;
	wire n18970;
	wire n18971;
	wire n18972;
	wire n18973;
	wire n18974;
	wire n18975;
	wire n18976;
	wire n18977;
	wire n18978;
	wire n18979;
	wire n18980;
	wire n18981;
	wire n18982;
	wire n18983;
	wire n18984;
	wire n18985;
	wire n18986;
	wire n18987;
	wire n18988;
	wire n18989;
	wire n18990;
	wire n18991;
	wire n18992;
	wire n18993;
	wire n18994;
	wire n18995;
	wire n18996;
	wire n18997;
	wire n18998;
	wire n18999;
	wire n19000;
	wire n19001;
	wire n19002;
	wire n19003;
	wire n19004;
	wire n19005;
	wire n19006;
	wire n19007;
	wire n19008;
	wire n19009;
	wire n19010;
	wire n19011;
	wire n19012;
	wire n19013;
	wire n19014;
	wire n19015;
	wire n19016;
	wire n19017;
	wire n19018;
	wire n19019;
	wire n19020;
	wire n19021;
	wire n19022;
	wire n19023;
	wire n19024;
	wire n19025;
	wire n19026;
	wire n19027;
	wire n19028;
	wire n19029;
	wire n19030;
	wire n19031;
	wire n19032;
	wire n19033;
	wire n19034;
	wire n19035;
	wire n19036;
	wire n19037;
	wire n19038;
	wire n19039;
	wire n19040;
	wire n19041;
	wire n19042;
	wire n19043;
	wire n19044;
	wire n19045;
	wire n19046;
	wire n19047;
	wire n19048;
	wire n19049;
	wire n19050;
	wire n19051;
	wire n19052;
	wire n19053;
	wire n19054;
	wire n19055;
	wire n19056;
	wire n19057;
	wire n19058;
	wire n19059;
	wire n19060;
	wire n19061;
	wire n19062;
	wire n19063;
	wire n19064;
	wire n19065;
	wire n19066;
	wire n19067;
	wire n19068;
	wire n19069;
	wire n19070;
	wire n19071;
	wire n19072;
	wire n19073;
	wire n19074;
	wire n19075;
	wire n19076;
	wire n19077;
	wire n19078;
	wire n19079;
	wire n19080;
	wire n19081;
	wire n19082;
	wire n19083;
	wire n19084;
	wire n19085;
	wire n19086;
	wire n19087;
	wire n19088;
	wire n19089;
	wire n19090;
	wire n19091;
	wire n19092;
	wire n19093;
	wire n19094;
	wire n19095;
	wire n19096;
	wire n19097;
	wire n19098;
	wire n19099;
	wire n19100;
	wire n19101;
	wire n19102;
	wire n19103;
	wire n19104;
	wire n19105;
	wire n19106;
	wire n19107;
	wire n19108;
	wire n19109;
	wire n19110;
	wire n19111;
	wire n19112;
	wire n19113;
	wire n19114;
	wire n19115;
	wire n19116;
	wire n19117;
	wire n19118;
	wire n19119;
	wire n19120;
	wire n19121;
	wire n19122;
	wire n19123;
	wire n19124;
	wire n19125;
	wire n19126;
	wire n19127;
	wire n19128;
	wire n19129;
	wire n19130;
	wire n19131;
	wire n19132;
	wire n19133;
	wire n19134;
	wire n19135;
	wire n19136;
	wire n19137;
	wire n19138;
	wire n19139;
	wire n19140;
	wire n19141;
	wire n19142;
	wire n19143;
	wire n19144;
	wire n19145;
	wire n19146;
	wire n19147;
	wire n19148;
	wire n19149;
	wire n19150;
	wire n19151;
	wire n19152;
	wire n19153;
	wire n19154;
	wire n19155;
	wire n19156;
	wire n19157;
	wire n19158;
	wire n19159;
	wire n19160;
	wire n19161;
	wire n19162;
	wire n19163;
	wire n19164;
	wire n19165;
	wire n19166;
	wire n19167;
	wire n19168;
	wire n19169;
	wire n19170;
	wire n19171;
	wire n19172;
	wire n19173;
	wire n19174;
	wire n19175;
	wire n19176;
	wire n19177;
	wire n19178;
	wire n19179;
	wire n19180;
	wire n19181;
	wire n19182;
	wire n19183;
	wire n19184;
	wire n19185;
	wire n19186;
	wire n19187;
	wire n19188;
	wire n19189;
	wire n19190;
	wire n19191;
	wire n19192;
	wire n19193;
	wire n19194;
	wire n19195;
	wire n19196;
	wire n19197;
	wire n19198;
	wire n19199;
	wire n19200;
	wire n19201;
	wire n19202;
	wire n19203;
	wire n19204;
	wire n19205;
	wire n19206;
	wire n19207;
	wire n19208;
	wire n19209;
	wire n19210;
	wire n19211;
	wire n19212;
	wire n19213;
	wire n19214;
	wire n19215;
	wire n19216;
	wire n19217;
	wire n19218;
	wire n19219;
	wire n19220;
	wire n19221;
	wire n19222;
	wire n19223;
	wire n19224;
	wire n19225;
	wire n19226;
	wire n19227;
	wire n19228;
	wire n19229;
	wire n19230;
	wire n19231;
	wire n19232;
	wire n19233;
	wire n19234;
	wire n19235;
	wire n19236;
	wire n19237;
	wire n19238;
	wire n19239;
	wire n19240;
	wire n19241;
	wire n19242;
	wire n19243;
	wire n19244;
	wire n19245;
	wire n19246;
	wire n19247;
	wire n19248;
	wire n19249;
	wire n19250;
	wire n19251;
	wire n19252;
	wire n19253;
	wire n19254;
	wire n19255;
	wire n19256;
	wire n19257;
	wire n19258;
	wire n19259;
	wire n19260;
	wire n19261;
	wire n19262;
	wire n19263;
	wire n19264;
	wire n19265;
	wire n19266;
	wire n19267;
	wire n19268;
	wire n19269;
	wire n19270;
	wire n19271;
	wire n19272;
	wire n19273;
	wire n19274;
	wire n19275;
	wire n19276;
	wire n19277;
	wire n19278;
	wire n19279;
	wire n19280;
	wire n19281;
	wire n19282;
	wire n19283;
	wire n19284;
	wire n19285;
	wire n19286;
	wire n19287;
	wire n19288;
	wire n19289;
	wire n19290;
	wire n19291;
	wire n19292;
	wire n19293;
	wire n19294;
	wire n19295;
	wire n19296;
	wire n19297;
	wire n19298;
	wire n19299;
	wire n19300;
	wire n19301;
	wire n19302;
	wire n19303;
	wire n19304;
	wire n19305;
	wire n19306;
	wire n19307;
	wire n19308;
	wire n19309;
	wire n19310;
	wire n19311;
	wire n19312;
	wire n19313;
	wire n19314;
	wire n19315;
	wire n19316;
	wire n19317;
	wire n19318;
	wire n19319;
	wire n19320;
	wire n19321;
	wire n19322;
	wire n19323;
	wire n19324;
	wire n19325;
	wire n19326;
	wire n19327;
	wire n19328;
	wire n19329;
	wire n19330;
	wire n19331;
	wire n19332;
	wire n19333;
	wire n19334;
	wire n19335;
	wire n19336;
	wire n19337;
	wire n19338;
	wire n19339;
	wire n19340;
	wire n19341;
	wire n19342;
	wire n19343;
	wire n19344;
	wire n19345;
	wire n19346;
	wire n19347;
	wire n19348;
	wire n19349;
	wire n19350;
	wire n19351;
	wire n19352;
	wire n19353;
	wire n19354;
	wire n19355;
	wire n19356;
	wire n19357;
	wire n19358;
	wire n19359;
	wire n19360;
	wire n19361;
	wire n19362;
	wire n19363;
	wire n19364;
	wire n19365;
	wire n19366;
	wire n19367;
	wire n19368;
	wire n19369;
	wire n19370;
	wire n19371;
	wire n19372;
	wire n19373;
	wire n19374;
	wire n19375;
	wire n19376;
	wire n19377;
	wire n19378;
	wire n19379;
	wire n19380;
	wire n19381;
	wire n19382;
	wire n19383;
	wire n19384;
	wire n19385;
	wire n19386;
	wire n19387;
	wire n19388;
	wire n19389;
	wire n19390;
	wire n19391;
	wire n19392;
	wire n19393;
	wire n19394;
	wire n19395;
	wire n19396;
	wire n19397;
	wire n19398;
	wire n19399;
	wire n19400;
	wire n19401;
	wire n19402;
	wire n19403;
	wire n19404;
	wire n19405;
	wire n19406;
	wire n19407;
	wire n19408;
	wire n19409;
	wire n19410;
	wire n19411;
	wire n19412;
	wire n19413;
	wire n19414;
	wire n19415;
	wire n19416;
	wire n19417;
	wire n19418;
	wire n19419;
	wire n19420;
	wire n19421;
	wire n19422;
	wire n19423;
	wire n19424;
	wire n19425;
	wire n19426;
	wire n19427;
	wire n19428;
	wire n19429;
	wire n19430;
	wire n19431;
	wire n19432;
	wire n19433;
	wire n19434;
	wire n19435;
	wire n19436;
	wire n19437;
	wire n19438;
	wire n19439;
	wire n19440;
	wire n19441;
	wire n19442;
	wire n19443;
	wire n19444;
	wire n19445;
	wire n19446;
	wire n19447;
	wire n19448;
	wire n19449;
	wire n19450;
	wire n19451;
	wire n19452;
	wire n19453;
	wire n19454;
	wire n19455;
	wire n19456;
	wire n19457;
	wire n19458;
	wire n19459;
	wire n19460;
	wire n19461;
	wire n19462;
	wire n19463;
	wire n19464;
	wire n19465;
	wire n19466;
	wire n19467;
	wire n19468;
	wire n19469;
	wire n19470;
	wire n19471;
	wire n19472;
	wire n19473;
	wire n19474;
	wire n19475;
	wire n19476;
	wire n19477;
	wire n19478;
	wire n19479;
	wire n19480;
	wire n19481;
	wire n19482;
	wire n19483;
	wire n19484;
	wire n19485;
	wire n19486;
	wire n19487;
	wire n19488;
	wire n19489;
	wire n19490;
	wire n19491;
	wire n19492;
	wire n19493;
	wire n19494;
	wire n19495;
	wire n19496;
	wire n19497;
	wire n19498;
	wire n19499;
	wire n19500;
	wire n19501;
	wire n19502;
	wire n19503;
	wire n19504;
	wire n19505;
	wire n19506;
	wire n19507;
	wire n19508;
	wire n19509;
	wire n19510;
	wire n19511;
	wire n19512;
	wire n19513;
	wire n19514;
	wire n19515;
	wire n19516;
	wire n19517;
	wire n19518;
	wire n19519;
	wire n19520;
	wire n19521;
	wire n19522;
	wire n19523;
	wire n19524;
	wire n19525;
	wire n19526;
	wire n19527;
	wire n19528;
	wire n19529;
	wire n19530;
	wire n19531;
	wire n19532;
	wire n19533;
	wire n19534;
	wire n19535;
	wire n19536;
	wire n19537;
	wire n19538;
	wire n19539;
	wire n19540;
	wire n19541;
	wire n19542;
	wire n19543;
	wire n19544;
	wire n19545;
	wire n19546;
	wire n19547;
	wire n19548;
	wire n19549;
	wire n19550;
	wire n19551;
	wire n19552;
	wire n19553;
	wire n19554;
	wire n19555;
	wire n19556;
	wire n19557;
	wire n19558;
	wire n19559;
	wire n19560;
	wire n19561;
	wire n19562;
	wire n19563;
	wire n19564;
	wire n19565;
	wire n19566;
	wire n19567;
	wire n19568;
	wire n19569;
	wire n19570;
	wire n19571;
	wire n19572;
	wire n19573;
	wire n19574;
	wire n19575;
	wire n19576;
	wire n19577;
	wire n19578;
	wire n19579;
	wire n19580;
	wire n19581;
	wire n19582;
	wire n19583;
	wire n19584;
	wire n19585;
	wire n19586;
	wire n19587;
	wire n19588;
	wire n19589;
	wire n19590;
	wire n19591;
	wire n19592;
	wire n19593;
	wire n19594;
	wire n19595;
	wire n19596;
	wire n19597;
	wire n19598;
	wire n19599;
	wire n19600;
	wire n19601;
	wire n19602;
	wire n19603;
	wire n19604;
	wire n19605;
	wire n19606;
	wire n19607;
	wire n19608;
	wire n19609;
	wire n19610;
	wire n19611;
	wire n19612;
	wire n19613;
	wire n19614;
	wire n19615;
	wire n19616;
	wire n19617;
	wire n19618;
	wire n19619;
	wire n19620;
	wire n19621;
	wire n19622;
	wire n19623;
	wire n19624;
	wire n19625;
	wire n19626;
	wire n19627;
	wire n19628;
	wire n19629;
	wire n19630;
	wire n19631;
	wire n19632;
	wire n19633;
	wire n19634;
	wire n19635;
	wire n19636;
	wire n19637;
	wire n19639;
	wire n19640;
	wire n19641;
	wire n19642;
	wire n19643;
	wire n19644;
	wire n19645;
	wire n19646;
	wire n19647;
	wire n19648;
	wire n19649;
	wire n19650;
	wire n19651;
	wire n19652;
	wire n19653;
	wire n19654;
	wire n19655;
	wire n19656;
	wire n19657;
	wire n19658;
	wire n19659;
	wire n19660;
	wire n19661;
	wire n19662;
	wire n19663;
	wire n19664;
	wire n19665;
	wire n19666;
	wire n19667;
	wire n19668;
	wire n19669;
	wire n19670;
	wire n19671;
	wire n19672;
	wire n19673;
	wire n19674;
	wire n19675;
	wire n19676;
	wire n19677;
	wire n19678;
	wire n19679;
	wire n19680;
	wire n19681;
	wire n19682;
	wire n19683;
	wire n19684;
	wire n19685;
	wire n19686;
	wire n19687;
	wire n19688;
	wire n19689;
	wire n19690;
	wire n19691;
	wire n19692;
	wire n19693;
	wire n19694;
	wire n19695;
	wire n19696;
	wire n19697;
	wire n19698;
	wire n19699;
	wire n19700;
	wire n19701;
	wire n19702;
	wire n19703;
	wire n19704;
	wire n19705;
	wire n19706;
	wire n19707;
	wire n19708;
	wire n19709;
	wire n19710;
	wire n19711;
	wire n19712;
	wire n19713;
	wire n19714;
	wire n19715;
	wire n19716;
	wire n19717;
	wire n19718;
	wire n19719;
	wire n19720;
	wire n19721;
	wire n19722;
	wire n19723;
	wire n19724;
	wire n19725;
	wire n19726;
	wire n19727;
	wire n19728;
	wire n19729;
	wire n19730;
	wire n19731;
	wire n19732;
	wire n19733;
	wire n19734;
	wire n19735;
	wire n19736;
	wire n19737;
	wire n19738;
	wire n19739;
	wire n19740;
	wire n19741;
	wire n19742;
	wire n19743;
	wire n19744;
	wire n19745;
	wire n19746;
	wire n19747;
	wire n19748;
	wire n19749;
	wire n19750;
	wire n19751;
	wire n19752;
	wire n19753;
	wire n19754;
	wire n19755;
	wire n19756;
	wire n19757;
	wire n19758;
	wire n19759;
	wire n19760;
	wire n19761;
	wire n19762;
	wire n19763;
	wire n19764;
	wire n19765;
	wire n19766;
	wire n19767;
	wire n19768;
	wire n19769;
	wire n19770;
	wire n19771;
	wire n19772;
	wire n19773;
	wire n19774;
	wire n19775;
	wire n19776;
	wire n19777;
	wire n19778;
	wire n19779;
	wire n19780;
	wire n19781;
	wire n19782;
	wire n19783;
	wire n19784;
	wire n19785;
	wire n19786;
	wire n19787;
	wire n19788;
	wire n19789;
	wire n19790;
	wire n19791;
	wire n19792;
	wire n19793;
	wire n19794;
	wire n19795;
	wire n19796;
	wire n19797;
	wire n19798;
	wire n19799;
	wire n19800;
	wire n19801;
	wire n19802;
	wire n19803;
	wire n19804;
	wire n19805;
	wire n19806;
	wire n19807;
	wire n19808;
	wire n19809;
	wire n19810;
	wire n19811;
	wire n19812;
	wire n19813;
	wire n19814;
	wire n19815;
	wire n19816;
	wire n19817;
	wire n19818;
	wire n19819;
	wire n19820;
	wire n19821;
	wire n19822;
	wire n19823;
	wire n19824;
	wire n19825;
	wire n19826;
	wire n19827;
	wire n19828;
	wire n19829;
	wire n19830;
	wire n19831;
	wire n19832;
	wire n19833;
	wire n19834;
	wire n19835;
	wire n19836;
	wire n19837;
	wire n19838;
	wire n19839;
	wire n19840;
	wire n19841;
	wire n19842;
	wire n19843;
	wire n19844;
	wire n19845;
	wire n19846;
	wire n19847;
	wire n19848;
	wire n19849;
	wire n19850;
	wire n19851;
	wire n19852;
	wire n19853;
	wire n19854;
	wire n19855;
	wire n19856;
	wire n19857;
	wire n19858;
	wire n19859;
	wire n19860;
	wire n19861;
	wire n19862;
	wire n19863;
	wire n19864;
	wire n19865;
	wire n19866;
	wire n19867;
	wire n19868;
	wire n19869;
	wire n19870;
	wire n19871;
	wire n19872;
	wire n19873;
	wire n19874;
	wire n19875;
	wire n19876;
	wire n19877;
	wire n19878;
	wire n19879;
	wire n19880;
	wire n19881;
	wire n19882;
	wire n19883;
	wire n19884;
	wire n19885;
	wire n19886;
	wire n19887;
	wire n19888;
	wire n19889;
	wire n19890;
	wire n19891;
	wire n19892;
	wire n19893;
	wire n19894;
	wire n19895;
	wire n19896;
	wire n19897;
	wire n19898;
	wire n19899;
	wire n19900;
	wire n19901;
	wire n19902;
	wire n19903;
	wire n19904;
	wire n19905;
	wire n19906;
	wire n19907;
	wire n19908;
	wire n19909;
	wire n19910;
	wire n19911;
	wire n19912;
	wire n19913;
	wire n19914;
	wire n19915;
	wire n19916;
	wire n19917;
	wire n19918;
	wire n19919;
	wire n19920;
	wire n19921;
	wire n19922;
	wire n19923;
	wire n19924;
	wire n19925;
	wire n19926;
	wire n19927;
	wire n19928;
	wire n19929;
	wire n19930;
	wire n19931;
	wire n19932;
	wire n19933;
	wire n19934;
	wire n19935;
	wire n19936;
	wire n19937;
	wire n19938;
	wire n19939;
	wire n19940;
	wire n19941;
	wire n19942;
	wire n19943;
	wire n19944;
	wire n19945;
	wire n19946;
	wire n19947;
	wire n19948;
	wire n19949;
	wire n19950;
	wire n19951;
	wire n19952;
	wire n19953;
	wire n19954;
	wire n19955;
	wire n19956;
	wire n19957;
	wire n19958;
	wire n19959;
	wire n19960;
	wire n19961;
	wire n19962;
	wire n19963;
	wire n19964;
	wire n19965;
	wire n19966;
	wire n19967;
	wire n19968;
	wire n19969;
	wire n19970;
	wire n19971;
	wire n19972;
	wire n19973;
	wire n19974;
	wire n19975;
	wire n19976;
	wire n19977;
	wire n19978;
	wire n19979;
	wire n19980;
	wire n19981;
	wire n19982;
	wire n19983;
	wire n19984;
	wire n19985;
	wire n19986;
	wire n19987;
	wire n19988;
	wire n19989;
	wire n19990;
	wire n19991;
	wire n19992;
	wire n19993;
	wire n19994;
	wire n19995;
	wire n19996;
	wire n19997;
	wire n19998;
	wire n19999;
	wire n20000;
	wire n20001;
	wire n20002;
	wire n20003;
	wire n20004;
	wire n20005;
	wire n20006;
	wire n20007;
	wire n20008;
	wire n20009;
	wire n20010;
	wire n20011;
	wire n20012;
	wire n20013;
	wire n20014;
	wire n20015;
	wire n20016;
	wire n20017;
	wire n20018;
	wire n20019;
	wire n20020;
	wire n20021;
	wire n20022;
	wire n20023;
	wire n20024;
	wire n20025;
	wire n20026;
	wire n20027;
	wire n20028;
	wire n20029;
	wire n20030;
	wire n20031;
	wire n20032;
	wire n20033;
	wire n20034;
	wire n20035;
	wire n20036;
	wire n20037;
	wire n20038;
	wire n20039;
	wire n20040;
	wire n20041;
	wire n20042;
	wire n20043;
	wire n20044;
	wire n20045;
	wire n20046;
	wire n20047;
	wire n20048;
	wire n20049;
	wire n20050;
	wire n20051;
	wire n20052;
	wire n20053;
	wire n20054;
	wire n20055;
	wire n20056;
	wire n20057;
	wire n20058;
	wire n20059;
	wire n20060;
	wire n20061;
	wire n20062;
	wire n20063;
	wire n20064;
	wire n20065;
	wire n20066;
	wire n20067;
	wire n20068;
	wire n20069;
	wire n20070;
	wire n20071;
	wire n20072;
	wire n20073;
	wire n20074;
	wire n20075;
	wire n20076;
	wire n20077;
	wire n20078;
	wire n20079;
	wire n20080;
	wire n20081;
	wire n20082;
	wire n20083;
	wire n20084;
	wire n20085;
	wire n20086;
	wire n20087;
	wire n20088;
	wire n20089;
	wire n20090;
	wire n20091;
	wire n20092;
	wire n20093;
	wire n20094;
	wire n20095;
	wire n20096;
	wire n20097;
	wire n20098;
	wire n20099;
	wire n20100;
	wire n20101;
	wire n20102;
	wire n20103;
	wire n20104;
	wire n20105;
	wire n20106;
	wire n20107;
	wire n20108;
	wire n20109;
	wire n20110;
	wire n20111;
	wire n20112;
	wire n20113;
	wire n20114;
	wire n20115;
	wire n20116;
	wire n20117;
	wire n20118;
	wire n20119;
	wire n20120;
	wire n20121;
	wire n20122;
	wire n20123;
	wire n20124;
	wire n20125;
	wire n20126;
	wire n20127;
	wire n20128;
	wire n20129;
	wire n20130;
	wire n20131;
	wire n20132;
	wire n20133;
	wire n20134;
	wire n20135;
	wire n20136;
	wire n20137;
	wire n20138;
	wire n20139;
	wire n20140;
	wire n20141;
	wire n20142;
	wire n20143;
	wire n20144;
	wire n20145;
	wire n20146;
	wire n20147;
	wire n20148;
	wire n20149;
	wire n20150;
	wire n20151;
	wire n20152;
	wire n20153;
	wire n20154;
	wire n20155;
	wire n20156;
	wire n20157;
	wire n20158;
	wire n20159;
	wire n20160;
	wire n20161;
	wire n20162;
	wire n20163;
	wire n20164;
	wire n20165;
	wire n20166;
	wire n20167;
	wire n20168;
	wire n20169;
	wire n20170;
	wire n20171;
	wire n20172;
	wire n20173;
	wire n20174;
	wire n20175;
	wire n20176;
	wire n20177;
	wire n20178;
	wire n20179;
	wire n20180;
	wire n20181;
	wire n20182;
	wire n20183;
	wire n20184;
	wire n20185;
	wire n20186;
	wire n20187;
	wire n20188;
	wire n20189;
	wire n20190;
	wire n20191;
	wire n20192;
	wire n20193;
	wire n20194;
	wire n20195;
	wire n20196;
	wire n20197;
	wire n20198;
	wire n20199;
	wire n20200;
	wire n20201;
	wire n20202;
	wire n20203;
	wire n20204;
	wire n20205;
	wire n20206;
	wire n20207;
	wire n20208;
	wire n20209;
	wire n20210;
	wire n20211;
	wire n20212;
	wire n20213;
	wire n20214;
	wire n20215;
	wire n20216;
	wire n20217;
	wire n20218;
	wire n20219;
	wire n20220;
	wire n20221;
	wire n20222;
	wire n20223;
	wire n20224;
	wire n20225;
	wire n20226;
	wire n20227;
	wire n20228;
	wire n20229;
	wire n20231;
	wire n20232;
	wire n20233;
	wire n20234;
	wire n20235;
	wire n20236;
	wire n20237;
	wire n20238;
	wire n20239;
	wire n20240;
	wire n20241;
	wire n20242;
	wire n20243;
	wire n20244;
	wire n20245;
	wire n20246;
	wire n20247;
	wire n20248;
	wire n20249;
	wire n20250;
	wire n20251;
	wire n20252;
	wire n20253;
	wire n20254;
	wire n20255;
	wire n20256;
	wire n20257;
	wire n20258;
	wire n20259;
	wire n20260;
	wire n20261;
	wire n20262;
	wire n20263;
	wire n20264;
	wire n20265;
	wire n20266;
	wire n20267;
	wire n20268;
	wire n20269;
	wire n20270;
	wire n20271;
	wire n20272;
	wire n20273;
	wire n20274;
	wire n20275;
	wire n20276;
	wire n20277;
	wire n20278;
	wire n20279;
	wire n20280;
	wire n20281;
	wire n20282;
	wire n20283;
	wire n20284;
	wire n20285;
	wire n20286;
	wire n20287;
	wire n20288;
	wire n20289;
	wire n20290;
	wire n20291;
	wire n20292;
	wire n20293;
	wire n20294;
	wire n20295;
	wire n20296;
	wire n20297;
	wire n20298;
	wire n20299;
	wire n20300;
	wire n20301;
	wire n20302;
	wire n20303;
	wire n20304;
	wire n20305;
	wire n20306;
	wire n20307;
	wire n20308;
	wire n20309;
	wire n20310;
	wire n20311;
	wire n20312;
	wire n20313;
	wire n20314;
	wire n20315;
	wire n20316;
	wire n20317;
	wire n20318;
	wire n20319;
	wire n20320;
	wire n20321;
	wire n20322;
	wire n20323;
	wire n20324;
	wire n20325;
	wire n20326;
	wire n20327;
	wire n20328;
	wire n20329;
	wire n20330;
	wire n20331;
	wire n20332;
	wire n20333;
	wire n20334;
	wire n20335;
	wire n20336;
	wire n20337;
	wire n20338;
	wire n20339;
	wire n20340;
	wire n20341;
	wire n20342;
	wire n20343;
	wire n20344;
	wire n20345;
	wire n20346;
	wire n20347;
	wire n20348;
	wire n20349;
	wire n20350;
	wire n20351;
	wire n20352;
	wire n20353;
	wire n20354;
	wire n20355;
	wire n20356;
	wire n20357;
	wire n20358;
	wire n20359;
	wire n20360;
	wire n20361;
	wire n20362;
	wire n20363;
	wire n20364;
	wire n20365;
	wire n20366;
	wire n20367;
	wire n20368;
	wire n20369;
	wire n20370;
	wire n20371;
	wire n20372;
	wire n20373;
	wire n20374;
	wire n20375;
	wire n20376;
	wire n20377;
	wire n20378;
	wire n20379;
	wire n20380;
	wire n20381;
	wire n20382;
	wire n20383;
	wire n20384;
	wire n20385;
	wire n20386;
	wire n20387;
	wire n20388;
	wire n20389;
	wire n20390;
	wire n20391;
	wire n20392;
	wire n20393;
	wire n20394;
	wire n20395;
	wire n20396;
	wire n20397;
	wire n20398;
	wire n20399;
	wire n20400;
	wire n20401;
	wire n20402;
	wire n20403;
	wire n20404;
	wire n20405;
	wire n20406;
	wire n20407;
	wire n20408;
	wire n20409;
	wire n20410;
	wire n20411;
	wire n20412;
	wire n20413;
	wire n20414;
	wire n20415;
	wire n20416;
	wire n20417;
	wire n20418;
	wire n20419;
	wire n20420;
	wire n20421;
	wire n20422;
	wire n20423;
	wire n20424;
	wire n20425;
	wire n20426;
	wire n20427;
	wire n20428;
	wire n20429;
	wire n20430;
	wire n20431;
	wire n20432;
	wire n20433;
	wire n20434;
	wire n20435;
	wire n20436;
	wire n20437;
	wire n20438;
	wire n20439;
	wire n20440;
	wire n20441;
	wire n20442;
	wire n20443;
	wire n20444;
	wire n20445;
	wire n20446;
	wire n20447;
	wire n20448;
	wire n20449;
	wire n20450;
	wire n20451;
	wire n20452;
	wire n20453;
	wire n20454;
	wire n20455;
	wire n20456;
	wire n20457;
	wire n20458;
	wire n20459;
	wire n20460;
	wire n20461;
	wire n20462;
	wire n20463;
	wire n20464;
	wire n20465;
	wire n20466;
	wire n20467;
	wire n20468;
	wire n20469;
	wire n20470;
	wire n20471;
	wire n20472;
	wire n20473;
	wire n20474;
	wire n20475;
	wire n20476;
	wire n20477;
	wire n20478;
	wire n20479;
	wire n20480;
	wire n20481;
	wire n20482;
	wire n20483;
	wire n20484;
	wire n20485;
	wire n20486;
	wire n20487;
	wire n20488;
	wire n20489;
	wire n20490;
	wire n20491;
	wire n20492;
	wire n20493;
	wire n20494;
	wire n20495;
	wire n20496;
	wire n20497;
	wire n20498;
	wire n20499;
	wire n20500;
	wire n20501;
	wire n20502;
	wire n20503;
	wire n20504;
	wire n20505;
	wire n20506;
	wire n20507;
	wire n20508;
	wire n20509;
	wire n20510;
	wire n20511;
	wire n20512;
	wire n20513;
	wire n20514;
	wire n20515;
	wire n20516;
	wire n20517;
	wire n20518;
	wire n20519;
	wire n20520;
	wire n20521;
	wire n20522;
	wire n20523;
	wire n20524;
	wire n20525;
	wire n20526;
	wire n20527;
	wire n20528;
	wire n20529;
	wire n20530;
	wire n20531;
	wire n20532;
	wire n20533;
	wire n20534;
	wire n20535;
	wire n20536;
	wire n20537;
	wire n20538;
	wire n20539;
	wire n20540;
	wire n20541;
	wire n20542;
	wire n20543;
	wire n20544;
	wire n20545;
	wire n20546;
	wire n20547;
	wire n20548;
	wire n20549;
	wire n20550;
	wire n20551;
	wire n20552;
	wire n20553;
	wire n20554;
	wire n20555;
	wire n20556;
	wire n20557;
	wire n20558;
	wire n20559;
	wire n20560;
	wire n20561;
	wire n20562;
	wire n20563;
	wire n20564;
	wire n20565;
	wire n20566;
	wire n20567;
	wire n20568;
	wire n20569;
	wire n20570;
	wire n20571;
	wire n20572;
	wire n20573;
	wire n20574;
	wire n20575;
	wire n20576;
	wire n20577;
	wire n20578;
	wire n20579;
	wire n20580;
	wire n20581;
	wire n20582;
	wire n20583;
	wire n20584;
	wire n20585;
	wire n20586;
	wire n20587;
	wire n20588;
	wire n20589;
	wire n20590;
	wire n20591;
	wire n20592;
	wire n20593;
	wire n20594;
	wire n20595;
	wire n20596;
	wire n20597;
	wire n20598;
	wire n20599;
	wire n20600;
	wire n20601;
	wire n20602;
	wire n20603;
	wire n20604;
	wire n20605;
	wire n20606;
	wire n20607;
	wire n20608;
	wire n20609;
	wire n20610;
	wire n20611;
	wire n20612;
	wire n20613;
	wire n20614;
	wire n20615;
	wire n20616;
	wire n20617;
	wire n20618;
	wire n20619;
	wire n20620;
	wire n20621;
	wire n20622;
	wire n20623;
	wire n20624;
	wire n20625;
	wire n20626;
	wire n20627;
	wire n20628;
	wire n20629;
	wire n20630;
	wire n20631;
	wire n20632;
	wire n20633;
	wire n20634;
	wire n20635;
	wire n20636;
	wire n20637;
	wire n20638;
	wire n20639;
	wire n20640;
	wire n20641;
	wire n20642;
	wire n20643;
	wire n20644;
	wire n20645;
	wire n20646;
	wire n20647;
	wire n20648;
	wire n20649;
	wire n20650;
	wire n20651;
	wire n20652;
	wire n20653;
	wire n20654;
	wire n20655;
	wire n20656;
	wire n20657;
	wire n20658;
	wire n20659;
	wire n20660;
	wire n20661;
	wire n20662;
	wire n20663;
	wire n20664;
	wire n20665;
	wire n20666;
	wire n20667;
	wire n20668;
	wire n20669;
	wire n20670;
	wire n20671;
	wire n20672;
	wire n20673;
	wire n20674;
	wire n20675;
	wire n20676;
	wire n20677;
	wire n20678;
	wire n20679;
	wire n20680;
	wire n20681;
	wire n20682;
	wire n20683;
	wire n20684;
	wire n20685;
	wire n20686;
	wire n20687;
	wire n20688;
	wire n20689;
	wire n20690;
	wire n20691;
	wire n20692;
	wire n20693;
	wire n20694;
	wire n20695;
	wire n20696;
	wire n20697;
	wire n20698;
	wire n20699;
	wire n20700;
	wire n20701;
	wire n20702;
	wire n20703;
	wire n20704;
	wire n20705;
	wire n20706;
	wire n20707;
	wire n20708;
	wire n20709;
	wire n20710;
	wire n20711;
	wire n20712;
	wire n20713;
	wire n20714;
	wire n20715;
	wire n20716;
	wire n20717;
	wire n20718;
	wire n20719;
	wire n20720;
	wire n20721;
	wire n20722;
	wire n20723;
	wire n20724;
	wire n20725;
	wire n20726;
	wire n20727;
	wire n20728;
	wire n20729;
	wire n20730;
	wire n20731;
	wire n20732;
	wire n20733;
	wire n20734;
	wire n20735;
	wire n20736;
	wire n20737;
	wire n20738;
	wire n20739;
	wire n20740;
	wire n20741;
	wire n20742;
	wire n20743;
	wire n20744;
	wire n20745;
	wire n20746;
	wire n20747;
	wire n20748;
	wire n20749;
	wire n20750;
	wire n20751;
	wire n20752;
	wire n20753;
	wire n20754;
	wire n20755;
	wire n20756;
	wire n20757;
	wire n20758;
	wire n20759;
	wire n20760;
	wire n20761;
	wire n20762;
	wire n20763;
	wire n20764;
	wire n20765;
	wire n20766;
	wire n20767;
	wire n20768;
	wire n20769;
	wire n20770;
	wire n20771;
	wire n20772;
	wire n20773;
	wire n20774;
	wire n20775;
	wire n20776;
	wire n20777;
	wire n20778;
	wire n20779;
	wire n20780;
	wire n20781;
	wire n20782;
	wire n20783;
	wire n20784;
	wire n20785;
	wire n20786;
	wire n20787;
	wire n20788;
	wire n20789;
	wire n20790;
	wire n20791;
	wire n20792;
	wire n20793;
	wire n20794;
	wire n20795;
	wire n20796;
	wire n20797;
	wire n20798;
	wire n20799;
	wire n20800;
	wire n20801;
	wire n20802;
	wire n20803;
	wire n20804;
	wire n20805;
	wire n20806;
	wire n20807;
	wire n20808;
	wire n20809;
	wire n20810;
	wire n20811;
	wire n20812;
	wire n20813;
	wire n20814;
	wire n20815;
	wire n20816;
	wire n20817;
	wire n20818;
	wire n20819;
	wire n20820;
	wire n20821;
	wire n20822;
	wire n20823;
	wire n20824;
	wire n20825;
	wire n20826;
	wire n20827;
	wire n20828;
	wire n20829;
	wire n20830;
	wire n20831;
	wire n20832;
	wire n20833;
	wire n20834;
	wire n20835;
	wire n20836;
	wire n20837;
	wire n20838;
	wire n20839;
	wire n20840;
	wire n20841;
	wire n20842;
	wire n20843;
	wire n20844;
	wire n20845;
	wire n20846;
	wire n20847;
	wire n20848;
	wire n20849;
	wire n20850;
	wire n20851;
	wire n20852;
	wire n20853;
	wire n20854;
	wire n20855;
	wire n20856;
	wire n20857;
	wire n20858;
	wire n20859;
	wire n20860;
	wire n20861;
	wire n20862;
	wire n20863;
	wire n20864;
	wire n20865;
	wire n20866;
	wire n20867;
	wire n20868;
	wire n20869;
	wire n20870;
	wire n20871;
	wire n20872;
	wire n20873;
	wire n20874;
	wire n20875;
	wire n20876;
	wire n20877;
	wire n20878;
	wire n20879;
	wire n20880;
	wire n20881;
	wire n20882;
	wire n20883;
	wire n20884;
	wire n20885;
	wire n20886;
	wire n20887;
	wire n20888;
	wire n20889;
	wire n20890;
	wire n20891;
	wire n20892;
	wire n20893;
	wire n20894;
	wire n20895;
	wire n20896;
	wire n20897;
	wire n20898;
	wire n20899;
	wire n20900;
	wire n20901;
	wire n20902;
	wire n20903;
	wire n20904;
	wire n20905;
	wire n20906;
	wire n20907;
	wire n20908;
	wire n20909;
	wire n20910;
	wire n20911;
	wire n20912;
	wire n20913;
	wire n20914;
	wire n20915;
	wire n20916;
	wire n20917;
	wire n20918;
	wire n20919;
	wire n20920;
	wire n20921;
	wire n20922;
	wire n20923;
	wire n20924;
	wire n20925;
	wire n20926;
	wire n20928;
	wire n20929;
	wire n20930;
	wire n20931;
	wire n20932;
	wire n20933;
	wire n20934;
	wire n20935;
	wire n20936;
	wire n20937;
	wire n20938;
	wire n20939;
	wire n20940;
	wire n20941;
	wire n20942;
	wire n20943;
	wire n20944;
	wire n20945;
	wire n20946;
	wire n20947;
	wire n20948;
	wire n20949;
	wire n20950;
	wire n20951;
	wire n20952;
	wire n20953;
	wire n20954;
	wire n20955;
	wire n20956;
	wire n20957;
	wire n20958;
	wire n20959;
	wire n20960;
	wire n20961;
	wire n20962;
	wire n20963;
	wire n20964;
	wire n20965;
	wire n20966;
	wire n20967;
	wire n20968;
	wire n20969;
	wire n20970;
	wire n20971;
	wire n20972;
	wire n20973;
	wire n20974;
	wire n20975;
	wire n20976;
	wire n20977;
	wire n20978;
	wire n20979;
	wire n20980;
	wire n20981;
	wire n20982;
	wire n20983;
	wire n20984;
	wire n20985;
	wire n20986;
	wire n20987;
	wire n20988;
	wire n20989;
	wire n20990;
	wire n20991;
	wire n20992;
	wire n20993;
	wire n20994;
	wire n20995;
	wire n20996;
	wire n20997;
	wire n20998;
	wire n20999;
	wire n21000;
	wire n21001;
	wire n21002;
	wire n21003;
	wire n21004;
	wire n21005;
	wire n21006;
	wire n21007;
	wire n21008;
	wire n21009;
	wire n21010;
	wire n21011;
	wire n21012;
	wire n21013;
	wire n21014;
	wire n21015;
	wire n21016;
	wire n21017;
	wire n21018;
	wire n21019;
	wire n21020;
	wire n21021;
	wire n21022;
	wire n21023;
	wire n21024;
	wire n21025;
	wire n21026;
	wire n21027;
	wire n21028;
	wire n21029;
	wire n21030;
	wire n21031;
	wire n21032;
	wire n21033;
	wire n21034;
	wire n21035;
	wire n21036;
	wire n21037;
	wire n21038;
	wire n21039;
	wire n21040;
	wire n21041;
	wire n21042;
	wire n21043;
	wire n21044;
	wire n21045;
	wire n21046;
	wire n21047;
	wire n21048;
	wire n21049;
	wire n21050;
	wire n21051;
	wire n21052;
	wire n21053;
	wire n21054;
	wire n21055;
	wire n21056;
	wire n21057;
	wire n21058;
	wire n21059;
	wire n21060;
	wire n21061;
	wire n21062;
	wire n21063;
	wire n21064;
	wire n21065;
	wire n21066;
	wire n21067;
	wire n21068;
	wire n21069;
	wire n21070;
	wire n21071;
	wire n21072;
	wire n21073;
	wire n21074;
	wire n21075;
	wire n21076;
	wire n21077;
	wire n21078;
	wire n21079;
	wire n21080;
	wire n21081;
	wire n21082;
	wire n21083;
	wire n21084;
	wire n21085;
	wire n21086;
	wire n21087;
	wire n21088;
	wire n21089;
	wire n21090;
	wire n21091;
	wire n21092;
	wire n21093;
	wire n21094;
	wire n21095;
	wire n21096;
	wire n21097;
	wire n21098;
	wire n21099;
	wire n21100;
	wire n21101;
	wire n21102;
	wire n21103;
	wire n21104;
	wire n21105;
	wire n21106;
	wire n21107;
	wire n21108;
	wire n21109;
	wire n21110;
	wire n21111;
	wire n21112;
	wire n21113;
	wire n21114;
	wire n21115;
	wire n21116;
	wire n21117;
	wire n21118;
	wire n21119;
	wire n21120;
	wire n21121;
	wire n21122;
	wire n21123;
	wire n21124;
	wire n21125;
	wire n21126;
	wire n21127;
	wire n21128;
	wire n21129;
	wire n21130;
	wire n21131;
	wire n21132;
	wire n21133;
	wire n21134;
	wire n21135;
	wire n21136;
	wire n21137;
	wire n21138;
	wire n21139;
	wire n21140;
	wire n21141;
	wire n21142;
	wire n21143;
	wire n21144;
	wire n21145;
	wire n21146;
	wire n21147;
	wire n21148;
	wire n21149;
	wire n21150;
	wire n21151;
	wire n21152;
	wire n21153;
	wire n21154;
	wire n21155;
	wire n21156;
	wire n21157;
	wire n21158;
	wire n21159;
	wire n21160;
	wire n21161;
	wire n21162;
	wire n21163;
	wire n21164;
	wire n21165;
	wire n21166;
	wire n21167;
	wire n21168;
	wire n21169;
	wire n21170;
	wire n21171;
	wire n21172;
	wire n21173;
	wire n21174;
	wire n21175;
	wire n21176;
	wire n21177;
	wire n21178;
	wire n21179;
	wire n21180;
	wire n21181;
	wire n21182;
	wire n21183;
	wire n21184;
	wire n21185;
	wire n21186;
	wire n21187;
	wire n21188;
	wire n21189;
	wire n21190;
	wire n21191;
	wire n21192;
	wire n21193;
	wire n21194;
	wire n21195;
	wire n21196;
	wire n21197;
	wire n21198;
	wire n21199;
	wire n21200;
	wire n21201;
	wire n21202;
	wire n21203;
	wire n21204;
	wire n21205;
	wire n21206;
	wire n21207;
	wire n21208;
	wire n21209;
	wire n21210;
	wire n21211;
	wire n21212;
	wire n21213;
	wire n21214;
	wire n21215;
	wire n21216;
	wire n21217;
	wire n21218;
	wire n21219;
	wire n21220;
	wire n21221;
	wire n21222;
	wire n21223;
	wire n21224;
	wire n21225;
	wire n21226;
	wire n21227;
	wire n21228;
	wire n21229;
	wire n21230;
	wire n21231;
	wire n21232;
	wire n21233;
	wire n21234;
	wire n21235;
	wire n21236;
	wire n21237;
	wire n21238;
	wire n21239;
	wire n21240;
	wire n21241;
	wire n21242;
	wire n21243;
	wire n21244;
	wire n21245;
	wire n21246;
	wire n21247;
	wire n21248;
	wire n21249;
	wire n21250;
	wire n21251;
	wire n21252;
	wire n21253;
	wire n21254;
	wire n21255;
	wire n21256;
	wire n21257;
	wire n21258;
	wire n21259;
	wire n21260;
	wire n21261;
	wire n21262;
	wire n21263;
	wire n21264;
	wire n21265;
	wire n21266;
	wire n21267;
	wire n21268;
	wire n21269;
	wire n21270;
	wire n21271;
	wire n21272;
	wire n21273;
	wire n21274;
	wire n21275;
	wire n21276;
	wire n21277;
	wire n21278;
	wire n21279;
	wire n21280;
	wire n21281;
	wire n21282;
	wire n21283;
	wire n21284;
	wire n21285;
	wire n21286;
	wire n21287;
	wire n21288;
	wire n21289;
	wire n21290;
	wire n21291;
	wire n21292;
	wire n21293;
	wire n21294;
	wire n21295;
	wire n21296;
	wire n21297;
	wire n21298;
	wire n21299;
	wire n21300;
	wire n21301;
	wire n21302;
	wire n21303;
	wire n21304;
	wire n21305;
	wire n21306;
	wire n21307;
	wire n21308;
	wire n21309;
	wire n21310;
	wire n21311;
	wire n21312;
	wire n21313;
	wire n21314;
	wire n21315;
	wire n21316;
	wire n21317;
	wire n21318;
	wire n21319;
	wire n21320;
	wire n21321;
	wire n21322;
	wire n21323;
	wire n21324;
	wire n21325;
	wire n21326;
	wire n21327;
	wire n21328;
	wire n21329;
	wire n21330;
	wire n21331;
	wire n21332;
	wire n21333;
	wire n21334;
	wire n21335;
	wire n21336;
	wire n21337;
	wire n21338;
	wire n21339;
	wire n21340;
	wire n21341;
	wire n21342;
	wire n21343;
	wire n21344;
	wire n21345;
	wire n21346;
	wire n21347;
	wire n21348;
	wire n21349;
	wire n21350;
	wire n21351;
	wire n21352;
	wire n21353;
	wire n21354;
	wire n21355;
	wire n21356;
	wire n21357;
	wire n21358;
	wire n21359;
	wire n21360;
	wire n21361;
	wire n21362;
	wire n21363;
	wire n21364;
	wire n21365;
	wire n21366;
	wire n21367;
	wire n21368;
	wire n21369;
	wire n21370;
	wire n21371;
	wire n21372;
	wire n21373;
	wire n21374;
	wire n21375;
	wire n21376;
	wire n21377;
	wire n21378;
	wire n21379;
	wire n21380;
	wire n21381;
	wire n21382;
	wire n21383;
	wire n21384;
	wire n21385;
	wire n21386;
	wire n21387;
	wire n21388;
	wire n21389;
	wire n21390;
	wire n21391;
	wire n21392;
	wire n21393;
	wire n21394;
	wire n21395;
	wire n21396;
	wire n21397;
	wire n21398;
	wire n21399;
	wire n21400;
	wire n21401;
	wire n21402;
	wire n21403;
	wire n21404;
	wire n21405;
	wire n21406;
	wire n21407;
	wire n21408;
	wire n21409;
	wire n21410;
	wire n21411;
	wire n21412;
	wire n21413;
	wire n21414;
	wire n21415;
	wire n21416;
	wire n21417;
	wire n21418;
	wire n21419;
	wire n21420;
	wire n21421;
	wire n21422;
	wire n21423;
	wire n21424;
	wire n21425;
	wire n21426;
	wire n21427;
	wire n21428;
	wire n21429;
	wire n21430;
	wire n21431;
	wire n21432;
	wire n21433;
	wire n21434;
	wire n21435;
	wire n21436;
	wire n21437;
	wire n21438;
	wire n21439;
	wire n21440;
	wire n21441;
	wire n21442;
	wire n21443;
	wire n21444;
	wire n21445;
	wire n21446;
	wire n21447;
	wire n21448;
	wire n21449;
	wire n21450;
	wire n21451;
	wire n21452;
	wire n21453;
	wire n21454;
	wire n21455;
	wire n21456;
	wire n21457;
	wire n21458;
	wire n21459;
	wire n21460;
	wire n21461;
	wire n21462;
	wire n21463;
	wire n21464;
	wire n21465;
	wire n21466;
	wire n21467;
	wire n21468;
	wire n21469;
	wire n21470;
	wire n21471;
	wire n21472;
	wire n21473;
	wire n21474;
	wire n21475;
	wire n21476;
	wire n21477;
	wire n21478;
	wire n21479;
	wire n21480;
	wire n21481;
	wire n21482;
	wire n21483;
	wire n21484;
	wire n21485;
	wire n21486;
	wire n21487;
	wire n21488;
	wire n21489;
	wire n21490;
	wire n21491;
	wire n21492;
	wire n21493;
	wire n21494;
	wire n21495;
	wire n21496;
	wire n21497;
	wire n21498;
	wire n21499;
	wire n21500;
	wire n21501;
	wire n21502;
	wire n21503;
	wire n21504;
	wire n21505;
	wire n21506;
	wire n21507;
	wire n21508;
	wire [2:0] w_a2_0;
	wire [1:0] w_a3_0;
	wire [1:0] w_a4_0;
	wire [1:0] w_a6_0;
	wire [1:0] w_a7_0;
	wire [1:0] w_a8_0;
	wire [1:0] w_a10_0;
	wire [1:0] w_a11_0;
	wire [1:0] w_a12_0;
	wire [1:0] w_a14_0;
	wire [1:0] w_a15_0;
	wire [1:0] w_a16_0;
	wire [1:0] w_a18_0;
	wire [1:0] w_a19_0;
	wire [1:0] w_a20_0;
	wire [1:0] w_a22_0;
	wire [1:0] w_a23_0;
	wire [1:0] w_a24_0;
	wire [1:0] w_a26_0;
	wire [1:0] w_a27_0;
	wire [1:0] w_a28_0;
	wire [1:0] w_a30_0;
	wire [1:0] w_a31_0;
	wire [1:0] w_a32_0;
	wire [1:0] w_a34_0;
	wire [1:0] w_a35_0;
	wire [1:0] w_a36_0;
	wire [1:0] w_a38_0;
	wire [1:0] w_a39_0;
	wire [1:0] w_a40_0;
	wire [1:0] w_a42_0;
	wire [1:0] w_a43_0;
	wire [1:0] w_a44_0;
	wire [1:0] w_a46_0;
	wire [1:0] w_a47_0;
	wire [1:0] w_a48_0;
	wire [1:0] w_a50_0;
	wire [1:0] w_a51_0;
	wire [1:0] w_a52_0;
	wire [1:0] w_a54_0;
	wire [1:0] w_a55_0;
	wire [1:0] w_a56_0;
	wire [1:0] w_a58_0;
	wire [1:0] w_a59_0;
	wire [1:0] w_a60_0;
	wire [1:0] w_a62_0;
	wire [1:0] w_a63_0;
	wire [1:0] w_a64_0;
	wire [1:0] w_a66_0;
	wire [1:0] w_a67_0;
	wire [1:0] w_a68_0;
	wire [1:0] w_a70_0;
	wire [1:0] w_a71_0;
	wire [1:0] w_a72_0;
	wire [1:0] w_a74_0;
	wire [1:0] w_a75_0;
	wire [1:0] w_a76_0;
	wire [1:0] w_a78_0;
	wire [1:0] w_a79_0;
	wire [1:0] w_a80_0;
	wire [1:0] w_a82_0;
	wire [1:0] w_a83_0;
	wire [1:0] w_a84_0;
	wire [1:0] w_a86_0;
	wire [1:0] w_a87_0;
	wire [1:0] w_a88_0;
	wire [1:0] w_a90_0;
	wire [1:0] w_a91_0;
	wire [1:0] w_a92_0;
	wire [1:0] w_a94_0;
	wire [1:0] w_a95_0;
	wire [1:0] w_a96_0;
	wire [1:0] w_a98_0;
	wire [1:0] w_a99_0;
	wire [1:0] w_a100_0;
	wire [1:0] w_a102_0;
	wire [1:0] w_a103_0;
	wire [1:0] w_a104_0;
	wire [1:0] w_a106_0;
	wire [1:0] w_a107_0;
	wire [1:0] w_a108_0;
	wire [1:0] w_a110_0;
	wire [1:0] w_a111_0;
	wire [1:0] w_a112_0;
	wire [1:0] w_a114_0;
	wire [1:0] w_a115_0;
	wire [1:0] w_a116_0;
	wire [1:0] w_a118_0;
	wire [1:0] w_a119_0;
	wire [1:0] w_a120_0;
	wire [1:0] w_a122_0;
	wire [1:0] w_a123_0;
	wire [2:0] w_a124_0;
	wire [1:0] w_a125_0;
	wire [2:0] w_a126_0;
	wire [1:0] w_a127_0;
	wire [2:0] w_asqrt1_0;
	wire [2:0] w_asqrt1_1;
	wire [2:0] w_asqrt1_2;
	wire [2:0] w_asqrt1_3;
	wire [2:0] w_asqrt1_4;
	wire [2:0] w_asqrt1_5;
	wire [2:0] w_asqrt1_6;
	wire [2:0] w_asqrt1_7;
	wire [2:0] w_asqrt1_8;
	wire [2:0] w_asqrt1_9;
	wire [2:0] w_asqrt1_10;
	wire [2:0] w_asqrt1_11;
	wire [2:0] w_asqrt1_12;
	wire [1:0] w_asqrt1_13;
	wire asqrt_fa_1;
	wire [2:0] w_asqrt2_0;
	wire [2:0] w_asqrt2_1;
	wire [2:0] w_asqrt2_2;
	wire [2:0] w_asqrt2_3;
	wire [2:0] w_asqrt2_4;
	wire [2:0] w_asqrt2_5;
	wire [2:0] w_asqrt2_6;
	wire [2:0] w_asqrt2_7;
	wire [2:0] w_asqrt2_8;
	wire [2:0] w_asqrt2_9;
	wire [2:0] w_asqrt2_10;
	wire [2:0] w_asqrt2_11;
	wire [2:0] w_asqrt2_12;
	wire [2:0] w_asqrt2_13;
	wire [2:0] w_asqrt2_14;
	wire [2:0] w_asqrt2_15;
	wire [2:0] w_asqrt2_16;
	wire [2:0] w_asqrt2_17;
	wire [2:0] w_asqrt2_18;
	wire [2:0] w_asqrt2_19;
	wire [2:0] w_asqrt2_20;
	wire [2:0] w_asqrt2_21;
	wire [2:0] w_asqrt2_22;
	wire [2:0] w_asqrt2_23;
	wire [2:0] w_asqrt2_24;
	wire [2:0] w_asqrt2_25;
	wire [2:0] w_asqrt2_26;
	wire [2:0] w_asqrt2_27;
	wire [2:0] w_asqrt2_28;
	wire [2:0] w_asqrt2_29;
	wire [2:0] w_asqrt2_30;
	wire w_asqrt2_31;
	wire asqrt_fa_2;
	wire [2:0] w_asqrt3_0;
	wire [2:0] w_asqrt3_1;
	wire [2:0] w_asqrt3_2;
	wire [2:0] w_asqrt3_3;
	wire [2:0] w_asqrt3_4;
	wire [2:0] w_asqrt3_5;
	wire [2:0] w_asqrt3_6;
	wire [2:0] w_asqrt3_7;
	wire [2:0] w_asqrt3_8;
	wire [2:0] w_asqrt3_9;
	wire [2:0] w_asqrt3_10;
	wire [2:0] w_asqrt3_11;
	wire [2:0] w_asqrt3_12;
	wire [2:0] w_asqrt3_13;
	wire [1:0] w_asqrt3_14;
	wire asqrt_fa_3;
	wire [2:0] w_asqrt4_0;
	wire [2:0] w_asqrt4_1;
	wire [2:0] w_asqrt4_2;
	wire [2:0] w_asqrt4_3;
	wire [2:0] w_asqrt4_4;
	wire [2:0] w_asqrt4_5;
	wire [2:0] w_asqrt4_6;
	wire [2:0] w_asqrt4_7;
	wire [2:0] w_asqrt4_8;
	wire [2:0] w_asqrt4_9;
	wire [2:0] w_asqrt4_10;
	wire [2:0] w_asqrt4_11;
	wire [2:0] w_asqrt4_12;
	wire [2:0] w_asqrt4_13;
	wire [2:0] w_asqrt4_14;
	wire [2:0] w_asqrt4_15;
	wire [2:0] w_asqrt4_16;
	wire [2:0] w_asqrt4_17;
	wire [2:0] w_asqrt4_18;
	wire [2:0] w_asqrt4_19;
	wire [2:0] w_asqrt4_20;
	wire [2:0] w_asqrt4_21;
	wire [2:0] w_asqrt4_22;
	wire [2:0] w_asqrt4_23;
	wire [2:0] w_asqrt4_24;
	wire [2:0] w_asqrt4_25;
	wire [2:0] w_asqrt4_26;
	wire [2:0] w_asqrt4_27;
	wire [2:0] w_asqrt4_28;
	wire [2:0] w_asqrt4_29;
	wire [2:0] w_asqrt4_30;
	wire w_asqrt4_31;
	wire asqrt_fa_4;
	wire [2:0] w_asqrt5_0;
	wire [2:0] w_asqrt5_1;
	wire [2:0] w_asqrt5_2;
	wire [2:0] w_asqrt5_3;
	wire [2:0] w_asqrt5_4;
	wire [2:0] w_asqrt5_5;
	wire [2:0] w_asqrt5_6;
	wire [2:0] w_asqrt5_7;
	wire [2:0] w_asqrt5_8;
	wire [2:0] w_asqrt5_9;
	wire [2:0] w_asqrt5_10;
	wire [2:0] w_asqrt5_11;
	wire [2:0] w_asqrt5_12;
	wire [2:0] w_asqrt5_13;
	wire [2:0] w_asqrt5_14;
	wire [1:0] w_asqrt5_15;
	wire asqrt_fa_5;
	wire [2:0] w_asqrt6_0;
	wire [2:0] w_asqrt6_1;
	wire [2:0] w_asqrt6_2;
	wire [2:0] w_asqrt6_3;
	wire [2:0] w_asqrt6_4;
	wire [2:0] w_asqrt6_5;
	wire [2:0] w_asqrt6_6;
	wire [2:0] w_asqrt6_7;
	wire [2:0] w_asqrt6_8;
	wire [2:0] w_asqrt6_9;
	wire [2:0] w_asqrt6_10;
	wire [2:0] w_asqrt6_11;
	wire [2:0] w_asqrt6_12;
	wire [2:0] w_asqrt6_13;
	wire [2:0] w_asqrt6_14;
	wire [2:0] w_asqrt6_15;
	wire [2:0] w_asqrt6_16;
	wire [2:0] w_asqrt6_17;
	wire [2:0] w_asqrt6_18;
	wire [2:0] w_asqrt6_19;
	wire [2:0] w_asqrt6_20;
	wire [2:0] w_asqrt6_21;
	wire [2:0] w_asqrt6_22;
	wire [2:0] w_asqrt6_23;
	wire [2:0] w_asqrt6_24;
	wire [2:0] w_asqrt6_25;
	wire [2:0] w_asqrt6_26;
	wire [2:0] w_asqrt6_27;
	wire [2:0] w_asqrt6_28;
	wire [2:0] w_asqrt6_29;
	wire [2:0] w_asqrt6_30;
	wire w_asqrt6_31;
	wire asqrt_fa_6;
	wire [2:0] w_asqrt7_0;
	wire [2:0] w_asqrt7_1;
	wire [2:0] w_asqrt7_2;
	wire [2:0] w_asqrt7_3;
	wire [2:0] w_asqrt7_4;
	wire [2:0] w_asqrt7_5;
	wire [2:0] w_asqrt7_6;
	wire [2:0] w_asqrt7_7;
	wire [2:0] w_asqrt7_8;
	wire [2:0] w_asqrt7_9;
	wire [2:0] w_asqrt7_10;
	wire [2:0] w_asqrt7_11;
	wire [2:0] w_asqrt7_12;
	wire [2:0] w_asqrt7_13;
	wire [2:0] w_asqrt7_14;
	wire w_asqrt7_15;
	wire asqrt_fa_7;
	wire [2:0] w_asqrt8_0;
	wire [2:0] w_asqrt8_1;
	wire [2:0] w_asqrt8_2;
	wire [2:0] w_asqrt8_3;
	wire [2:0] w_asqrt8_4;
	wire [2:0] w_asqrt8_5;
	wire [2:0] w_asqrt8_6;
	wire [2:0] w_asqrt8_7;
	wire [2:0] w_asqrt8_8;
	wire [2:0] w_asqrt8_9;
	wire [2:0] w_asqrt8_10;
	wire [2:0] w_asqrt8_11;
	wire [2:0] w_asqrt8_12;
	wire [2:0] w_asqrt8_13;
	wire [2:0] w_asqrt8_14;
	wire [2:0] w_asqrt8_15;
	wire [2:0] w_asqrt8_16;
	wire [2:0] w_asqrt8_17;
	wire [2:0] w_asqrt8_18;
	wire [2:0] w_asqrt8_19;
	wire [2:0] w_asqrt8_20;
	wire [2:0] w_asqrt8_21;
	wire [2:0] w_asqrt8_22;
	wire [2:0] w_asqrt8_23;
	wire [2:0] w_asqrt8_24;
	wire [2:0] w_asqrt8_25;
	wire [2:0] w_asqrt8_26;
	wire [2:0] w_asqrt8_27;
	wire [2:0] w_asqrt8_28;
	wire [2:0] w_asqrt8_29;
	wire [2:0] w_asqrt8_30;
	wire w_asqrt8_31;
	wire asqrt_fa_8;
	wire [2:0] w_asqrt9_0;
	wire [2:0] w_asqrt9_1;
	wire [2:0] w_asqrt9_2;
	wire [2:0] w_asqrt9_3;
	wire [2:0] w_asqrt9_4;
	wire [2:0] w_asqrt9_5;
	wire [2:0] w_asqrt9_6;
	wire [2:0] w_asqrt9_7;
	wire [2:0] w_asqrt9_8;
	wire [2:0] w_asqrt9_9;
	wire [2:0] w_asqrt9_10;
	wire [2:0] w_asqrt9_11;
	wire [2:0] w_asqrt9_12;
	wire [2:0] w_asqrt9_13;
	wire [2:0] w_asqrt9_14;
	wire [2:0] w_asqrt9_15;
	wire w_asqrt9_16;
	wire asqrt_fa_9;
	wire [2:0] w_asqrt10_0;
	wire [2:0] w_asqrt10_1;
	wire [2:0] w_asqrt10_2;
	wire [2:0] w_asqrt10_3;
	wire [2:0] w_asqrt10_4;
	wire [2:0] w_asqrt10_5;
	wire [2:0] w_asqrt10_6;
	wire [2:0] w_asqrt10_7;
	wire [2:0] w_asqrt10_8;
	wire [2:0] w_asqrt10_9;
	wire [2:0] w_asqrt10_10;
	wire [2:0] w_asqrt10_11;
	wire [2:0] w_asqrt10_12;
	wire [2:0] w_asqrt10_13;
	wire [2:0] w_asqrt10_14;
	wire [2:0] w_asqrt10_15;
	wire [2:0] w_asqrt10_16;
	wire [2:0] w_asqrt10_17;
	wire [2:0] w_asqrt10_18;
	wire [2:0] w_asqrt10_19;
	wire [2:0] w_asqrt10_20;
	wire [2:0] w_asqrt10_21;
	wire [2:0] w_asqrt10_22;
	wire [2:0] w_asqrt10_23;
	wire [2:0] w_asqrt10_24;
	wire [2:0] w_asqrt10_25;
	wire [2:0] w_asqrt10_26;
	wire [2:0] w_asqrt10_27;
	wire [2:0] w_asqrt10_28;
	wire [2:0] w_asqrt10_29;
	wire [2:0] w_asqrt10_30;
	wire w_asqrt10_31;
	wire asqrt_fa_10;
	wire [2:0] w_asqrt11_0;
	wire [2:0] w_asqrt11_1;
	wire [2:0] w_asqrt11_2;
	wire [2:0] w_asqrt11_3;
	wire [2:0] w_asqrt11_4;
	wire [2:0] w_asqrt11_5;
	wire [2:0] w_asqrt11_6;
	wire [2:0] w_asqrt11_7;
	wire [2:0] w_asqrt11_8;
	wire [2:0] w_asqrt11_9;
	wire [2:0] w_asqrt11_10;
	wire [2:0] w_asqrt11_11;
	wire [2:0] w_asqrt11_12;
	wire [2:0] w_asqrt11_13;
	wire [2:0] w_asqrt11_14;
	wire [2:0] w_asqrt11_15;
	wire w_asqrt11_16;
	wire asqrt_fa_11;
	wire [2:0] w_asqrt12_0;
	wire [2:0] w_asqrt12_1;
	wire [2:0] w_asqrt12_2;
	wire [2:0] w_asqrt12_3;
	wire [2:0] w_asqrt12_4;
	wire [2:0] w_asqrt12_5;
	wire [2:0] w_asqrt12_6;
	wire [2:0] w_asqrt12_7;
	wire [2:0] w_asqrt12_8;
	wire [2:0] w_asqrt12_9;
	wire [2:0] w_asqrt12_10;
	wire [2:0] w_asqrt12_11;
	wire [2:0] w_asqrt12_12;
	wire [2:0] w_asqrt12_13;
	wire [2:0] w_asqrt12_14;
	wire [2:0] w_asqrt12_15;
	wire [2:0] w_asqrt12_16;
	wire [2:0] w_asqrt12_17;
	wire [2:0] w_asqrt12_18;
	wire [2:0] w_asqrt12_19;
	wire [2:0] w_asqrt12_20;
	wire [2:0] w_asqrt12_21;
	wire [2:0] w_asqrt12_22;
	wire [2:0] w_asqrt12_23;
	wire [2:0] w_asqrt12_24;
	wire [2:0] w_asqrt12_25;
	wire [2:0] w_asqrt12_26;
	wire [2:0] w_asqrt12_27;
	wire [2:0] w_asqrt12_28;
	wire [2:0] w_asqrt12_29;
	wire [2:0] w_asqrt12_30;
	wire w_asqrt12_31;
	wire asqrt_fa_12;
	wire [2:0] w_asqrt13_0;
	wire [2:0] w_asqrt13_1;
	wire [2:0] w_asqrt13_2;
	wire [2:0] w_asqrt13_3;
	wire [2:0] w_asqrt13_4;
	wire [2:0] w_asqrt13_5;
	wire [2:0] w_asqrt13_6;
	wire [2:0] w_asqrt13_7;
	wire [2:0] w_asqrt13_8;
	wire [2:0] w_asqrt13_9;
	wire [2:0] w_asqrt13_10;
	wire [2:0] w_asqrt13_11;
	wire [2:0] w_asqrt13_12;
	wire [2:0] w_asqrt13_13;
	wire [2:0] w_asqrt13_14;
	wire [2:0] w_asqrt13_15;
	wire [2:0] w_asqrt13_16;
	wire w_asqrt13_17;
	wire asqrt_fa_13;
	wire [2:0] w_asqrt14_0;
	wire [2:0] w_asqrt14_1;
	wire [2:0] w_asqrt14_2;
	wire [2:0] w_asqrt14_3;
	wire [2:0] w_asqrt14_4;
	wire [2:0] w_asqrt14_5;
	wire [2:0] w_asqrt14_6;
	wire [2:0] w_asqrt14_7;
	wire [2:0] w_asqrt14_8;
	wire [2:0] w_asqrt14_9;
	wire [2:0] w_asqrt14_10;
	wire [2:0] w_asqrt14_11;
	wire [2:0] w_asqrt14_12;
	wire [2:0] w_asqrt14_13;
	wire [2:0] w_asqrt14_14;
	wire [2:0] w_asqrt14_15;
	wire [2:0] w_asqrt14_16;
	wire [2:0] w_asqrt14_17;
	wire [2:0] w_asqrt14_18;
	wire [2:0] w_asqrt14_19;
	wire [2:0] w_asqrt14_20;
	wire [2:0] w_asqrt14_21;
	wire [2:0] w_asqrt14_22;
	wire [2:0] w_asqrt14_23;
	wire [2:0] w_asqrt14_24;
	wire [2:0] w_asqrt14_25;
	wire [2:0] w_asqrt14_26;
	wire [2:0] w_asqrt14_27;
	wire [2:0] w_asqrt14_28;
	wire [2:0] w_asqrt14_29;
	wire [2:0] w_asqrt14_30;
	wire w_asqrt14_31;
	wire asqrt_fa_14;
	wire [2:0] w_asqrt15_0;
	wire [2:0] w_asqrt15_1;
	wire [2:0] w_asqrt15_2;
	wire [2:0] w_asqrt15_3;
	wire [2:0] w_asqrt15_4;
	wire [2:0] w_asqrt15_5;
	wire [2:0] w_asqrt15_6;
	wire [2:0] w_asqrt15_7;
	wire [2:0] w_asqrt15_8;
	wire [2:0] w_asqrt15_9;
	wire [2:0] w_asqrt15_10;
	wire [2:0] w_asqrt15_11;
	wire [2:0] w_asqrt15_12;
	wire [2:0] w_asqrt15_13;
	wire [2:0] w_asqrt15_14;
	wire [2:0] w_asqrt15_15;
	wire [2:0] w_asqrt15_16;
	wire w_asqrt15_17;
	wire asqrt_fa_15;
	wire [2:0] w_asqrt16_0;
	wire [2:0] w_asqrt16_1;
	wire [2:0] w_asqrt16_2;
	wire [2:0] w_asqrt16_3;
	wire [2:0] w_asqrt16_4;
	wire [2:0] w_asqrt16_5;
	wire [2:0] w_asqrt16_6;
	wire [2:0] w_asqrt16_7;
	wire [2:0] w_asqrt16_8;
	wire [2:0] w_asqrt16_9;
	wire [2:0] w_asqrt16_10;
	wire [2:0] w_asqrt16_11;
	wire [2:0] w_asqrt16_12;
	wire [2:0] w_asqrt16_13;
	wire [2:0] w_asqrt16_14;
	wire [2:0] w_asqrt16_15;
	wire [2:0] w_asqrt16_16;
	wire [2:0] w_asqrt16_17;
	wire [2:0] w_asqrt16_18;
	wire [2:0] w_asqrt16_19;
	wire [2:0] w_asqrt16_20;
	wire [2:0] w_asqrt16_21;
	wire [2:0] w_asqrt16_22;
	wire [2:0] w_asqrt16_23;
	wire [2:0] w_asqrt16_24;
	wire [2:0] w_asqrt16_25;
	wire [2:0] w_asqrt16_26;
	wire [2:0] w_asqrt16_27;
	wire [2:0] w_asqrt16_28;
	wire [2:0] w_asqrt16_29;
	wire [2:0] w_asqrt16_30;
	wire w_asqrt16_31;
	wire asqrt_fa_16;
	wire [2:0] w_asqrt17_0;
	wire [2:0] w_asqrt17_1;
	wire [2:0] w_asqrt17_2;
	wire [2:0] w_asqrt17_3;
	wire [2:0] w_asqrt17_4;
	wire [2:0] w_asqrt17_5;
	wire [2:0] w_asqrt17_6;
	wire [2:0] w_asqrt17_7;
	wire [2:0] w_asqrt17_8;
	wire [2:0] w_asqrt17_9;
	wire [2:0] w_asqrt17_10;
	wire [2:0] w_asqrt17_11;
	wire [2:0] w_asqrt17_12;
	wire [2:0] w_asqrt17_13;
	wire [2:0] w_asqrt17_14;
	wire [2:0] w_asqrt17_15;
	wire [2:0] w_asqrt17_16;
	wire [2:0] w_asqrt17_17;
	wire w_asqrt17_18;
	wire asqrt_fa_17;
	wire [2:0] w_asqrt18_0;
	wire [2:0] w_asqrt18_1;
	wire [2:0] w_asqrt18_2;
	wire [2:0] w_asqrt18_3;
	wire [2:0] w_asqrt18_4;
	wire [2:0] w_asqrt18_5;
	wire [2:0] w_asqrt18_6;
	wire [2:0] w_asqrt18_7;
	wire [2:0] w_asqrt18_8;
	wire [2:0] w_asqrt18_9;
	wire [2:0] w_asqrt18_10;
	wire [2:0] w_asqrt18_11;
	wire [2:0] w_asqrt18_12;
	wire [2:0] w_asqrt18_13;
	wire [2:0] w_asqrt18_14;
	wire [2:0] w_asqrt18_15;
	wire [2:0] w_asqrt18_16;
	wire [2:0] w_asqrt18_17;
	wire [2:0] w_asqrt18_18;
	wire [2:0] w_asqrt18_19;
	wire [2:0] w_asqrt18_20;
	wire [2:0] w_asqrt18_21;
	wire [2:0] w_asqrt18_22;
	wire [2:0] w_asqrt18_23;
	wire [2:0] w_asqrt18_24;
	wire [2:0] w_asqrt18_25;
	wire [2:0] w_asqrt18_26;
	wire [2:0] w_asqrt18_27;
	wire [2:0] w_asqrt18_28;
	wire [2:0] w_asqrt18_29;
	wire [2:0] w_asqrt18_30;
	wire w_asqrt18_31;
	wire asqrt_fa_18;
	wire [2:0] w_asqrt19_0;
	wire [2:0] w_asqrt19_1;
	wire [2:0] w_asqrt19_2;
	wire [2:0] w_asqrt19_3;
	wire [2:0] w_asqrt19_4;
	wire [2:0] w_asqrt19_5;
	wire [2:0] w_asqrt19_6;
	wire [2:0] w_asqrt19_7;
	wire [2:0] w_asqrt19_8;
	wire [2:0] w_asqrt19_9;
	wire [2:0] w_asqrt19_10;
	wire [2:0] w_asqrt19_11;
	wire [2:0] w_asqrt19_12;
	wire [2:0] w_asqrt19_13;
	wire [2:0] w_asqrt19_14;
	wire [2:0] w_asqrt19_15;
	wire [2:0] w_asqrt19_16;
	wire [2:0] w_asqrt19_17;
	wire w_asqrt19_18;
	wire asqrt_fa_19;
	wire [2:0] w_asqrt20_0;
	wire [2:0] w_asqrt20_1;
	wire [2:0] w_asqrt20_2;
	wire [2:0] w_asqrt20_3;
	wire [2:0] w_asqrt20_4;
	wire [2:0] w_asqrt20_5;
	wire [2:0] w_asqrt20_6;
	wire [2:0] w_asqrt20_7;
	wire [2:0] w_asqrt20_8;
	wire [2:0] w_asqrt20_9;
	wire [2:0] w_asqrt20_10;
	wire [2:0] w_asqrt20_11;
	wire [2:0] w_asqrt20_12;
	wire [2:0] w_asqrt20_13;
	wire [2:0] w_asqrt20_14;
	wire [2:0] w_asqrt20_15;
	wire [2:0] w_asqrt20_16;
	wire [2:0] w_asqrt20_17;
	wire [2:0] w_asqrt20_18;
	wire [2:0] w_asqrt20_19;
	wire [2:0] w_asqrt20_20;
	wire [2:0] w_asqrt20_21;
	wire [2:0] w_asqrt20_22;
	wire [2:0] w_asqrt20_23;
	wire [2:0] w_asqrt20_24;
	wire [2:0] w_asqrt20_25;
	wire [2:0] w_asqrt20_26;
	wire [2:0] w_asqrt20_27;
	wire [2:0] w_asqrt20_28;
	wire [2:0] w_asqrt20_29;
	wire [2:0] w_asqrt20_30;
	wire w_asqrt20_31;
	wire asqrt_fa_20;
	wire [2:0] w_asqrt21_0;
	wire [2:0] w_asqrt21_1;
	wire [2:0] w_asqrt21_2;
	wire [2:0] w_asqrt21_3;
	wire [2:0] w_asqrt21_4;
	wire [2:0] w_asqrt21_5;
	wire [2:0] w_asqrt21_6;
	wire [2:0] w_asqrt21_7;
	wire [2:0] w_asqrt21_8;
	wire [2:0] w_asqrt21_9;
	wire [2:0] w_asqrt21_10;
	wire [2:0] w_asqrt21_11;
	wire [2:0] w_asqrt21_12;
	wire [2:0] w_asqrt21_13;
	wire [2:0] w_asqrt21_14;
	wire [2:0] w_asqrt21_15;
	wire [2:0] w_asqrt21_16;
	wire [2:0] w_asqrt21_17;
	wire [2:0] w_asqrt21_18;
	wire w_asqrt21_19;
	wire asqrt_fa_21;
	wire [2:0] w_asqrt22_0;
	wire [2:0] w_asqrt22_1;
	wire [2:0] w_asqrt22_2;
	wire [2:0] w_asqrt22_3;
	wire [2:0] w_asqrt22_4;
	wire [2:0] w_asqrt22_5;
	wire [2:0] w_asqrt22_6;
	wire [2:0] w_asqrt22_7;
	wire [2:0] w_asqrt22_8;
	wire [2:0] w_asqrt22_9;
	wire [2:0] w_asqrt22_10;
	wire [2:0] w_asqrt22_11;
	wire [2:0] w_asqrt22_12;
	wire [2:0] w_asqrt22_13;
	wire [2:0] w_asqrt22_14;
	wire [2:0] w_asqrt22_15;
	wire [2:0] w_asqrt22_16;
	wire [2:0] w_asqrt22_17;
	wire [2:0] w_asqrt22_18;
	wire [2:0] w_asqrt22_19;
	wire [2:0] w_asqrt22_20;
	wire [2:0] w_asqrt22_21;
	wire [2:0] w_asqrt22_22;
	wire [2:0] w_asqrt22_23;
	wire [2:0] w_asqrt22_24;
	wire [2:0] w_asqrt22_25;
	wire [2:0] w_asqrt22_26;
	wire [2:0] w_asqrt22_27;
	wire [2:0] w_asqrt22_28;
	wire [2:0] w_asqrt22_29;
	wire [2:0] w_asqrt22_30;
	wire w_asqrt22_31;
	wire asqrt_fa_22;
	wire [2:0] w_asqrt23_0;
	wire [2:0] w_asqrt23_1;
	wire [2:0] w_asqrt23_2;
	wire [2:0] w_asqrt23_3;
	wire [2:0] w_asqrt23_4;
	wire [2:0] w_asqrt23_5;
	wire [2:0] w_asqrt23_6;
	wire [2:0] w_asqrt23_7;
	wire [2:0] w_asqrt23_8;
	wire [2:0] w_asqrt23_9;
	wire [2:0] w_asqrt23_10;
	wire [2:0] w_asqrt23_11;
	wire [2:0] w_asqrt23_12;
	wire [2:0] w_asqrt23_13;
	wire [2:0] w_asqrt23_14;
	wire [2:0] w_asqrt23_15;
	wire [2:0] w_asqrt23_16;
	wire [2:0] w_asqrt23_17;
	wire [2:0] w_asqrt23_18;
	wire w_asqrt23_19;
	wire asqrt_fa_23;
	wire [2:0] w_asqrt24_0;
	wire [2:0] w_asqrt24_1;
	wire [2:0] w_asqrt24_2;
	wire [2:0] w_asqrt24_3;
	wire [2:0] w_asqrt24_4;
	wire [2:0] w_asqrt24_5;
	wire [2:0] w_asqrt24_6;
	wire [2:0] w_asqrt24_7;
	wire [2:0] w_asqrt24_8;
	wire [2:0] w_asqrt24_9;
	wire [2:0] w_asqrt24_10;
	wire [2:0] w_asqrt24_11;
	wire [2:0] w_asqrt24_12;
	wire [2:0] w_asqrt24_13;
	wire [2:0] w_asqrt24_14;
	wire [2:0] w_asqrt24_15;
	wire [2:0] w_asqrt24_16;
	wire [2:0] w_asqrt24_17;
	wire [2:0] w_asqrt24_18;
	wire [2:0] w_asqrt24_19;
	wire [2:0] w_asqrt24_20;
	wire [2:0] w_asqrt24_21;
	wire [2:0] w_asqrt24_22;
	wire [2:0] w_asqrt24_23;
	wire [2:0] w_asqrt24_24;
	wire [2:0] w_asqrt24_25;
	wire [2:0] w_asqrt24_26;
	wire [2:0] w_asqrt24_27;
	wire [2:0] w_asqrt24_28;
	wire [2:0] w_asqrt24_29;
	wire [2:0] w_asqrt24_30;
	wire w_asqrt24_31;
	wire asqrt_fa_24;
	wire [2:0] w_asqrt25_0;
	wire [2:0] w_asqrt25_1;
	wire [2:0] w_asqrt25_2;
	wire [2:0] w_asqrt25_3;
	wire [2:0] w_asqrt25_4;
	wire [2:0] w_asqrt25_5;
	wire [2:0] w_asqrt25_6;
	wire [2:0] w_asqrt25_7;
	wire [2:0] w_asqrt25_8;
	wire [2:0] w_asqrt25_9;
	wire [2:0] w_asqrt25_10;
	wire [2:0] w_asqrt25_11;
	wire [2:0] w_asqrt25_12;
	wire [2:0] w_asqrt25_13;
	wire [2:0] w_asqrt25_14;
	wire [2:0] w_asqrt25_15;
	wire [2:0] w_asqrt25_16;
	wire [2:0] w_asqrt25_17;
	wire [2:0] w_asqrt25_18;
	wire [2:0] w_asqrt25_19;
	wire w_asqrt25_20;
	wire asqrt_fa_25;
	wire [2:0] w_asqrt26_0;
	wire [2:0] w_asqrt26_1;
	wire [2:0] w_asqrt26_2;
	wire [2:0] w_asqrt26_3;
	wire [2:0] w_asqrt26_4;
	wire [2:0] w_asqrt26_5;
	wire [2:0] w_asqrt26_6;
	wire [2:0] w_asqrt26_7;
	wire [2:0] w_asqrt26_8;
	wire [2:0] w_asqrt26_9;
	wire [2:0] w_asqrt26_10;
	wire [2:0] w_asqrt26_11;
	wire [2:0] w_asqrt26_12;
	wire [2:0] w_asqrt26_13;
	wire [2:0] w_asqrt26_14;
	wire [2:0] w_asqrt26_15;
	wire [2:0] w_asqrt26_16;
	wire [2:0] w_asqrt26_17;
	wire [2:0] w_asqrt26_18;
	wire [2:0] w_asqrt26_19;
	wire [2:0] w_asqrt26_20;
	wire [2:0] w_asqrt26_21;
	wire [2:0] w_asqrt26_22;
	wire [2:0] w_asqrt26_23;
	wire [2:0] w_asqrt26_24;
	wire [2:0] w_asqrt26_25;
	wire [2:0] w_asqrt26_26;
	wire [2:0] w_asqrt26_27;
	wire [2:0] w_asqrt26_28;
	wire [2:0] w_asqrt26_29;
	wire [2:0] w_asqrt26_30;
	wire w_asqrt26_31;
	wire asqrt_fa_26;
	wire [2:0] w_asqrt27_0;
	wire [2:0] w_asqrt27_1;
	wire [2:0] w_asqrt27_2;
	wire [2:0] w_asqrt27_3;
	wire [2:0] w_asqrt27_4;
	wire [2:0] w_asqrt27_5;
	wire [2:0] w_asqrt27_6;
	wire [2:0] w_asqrt27_7;
	wire [2:0] w_asqrt27_8;
	wire [2:0] w_asqrt27_9;
	wire [2:0] w_asqrt27_10;
	wire [2:0] w_asqrt27_11;
	wire [2:0] w_asqrt27_12;
	wire [2:0] w_asqrt27_13;
	wire [2:0] w_asqrt27_14;
	wire [2:0] w_asqrt27_15;
	wire [2:0] w_asqrt27_16;
	wire [2:0] w_asqrt27_17;
	wire [2:0] w_asqrt27_18;
	wire [2:0] w_asqrt27_19;
	wire [1:0] w_asqrt27_20;
	wire asqrt_fa_27;
	wire [2:0] w_asqrt28_0;
	wire [2:0] w_asqrt28_1;
	wire [2:0] w_asqrt28_2;
	wire [2:0] w_asqrt28_3;
	wire [2:0] w_asqrt28_4;
	wire [2:0] w_asqrt28_5;
	wire [2:0] w_asqrt28_6;
	wire [2:0] w_asqrt28_7;
	wire [2:0] w_asqrt28_8;
	wire [2:0] w_asqrt28_9;
	wire [2:0] w_asqrt28_10;
	wire [2:0] w_asqrt28_11;
	wire [2:0] w_asqrt28_12;
	wire [2:0] w_asqrt28_13;
	wire [2:0] w_asqrt28_14;
	wire [2:0] w_asqrt28_15;
	wire [2:0] w_asqrt28_16;
	wire [2:0] w_asqrt28_17;
	wire [2:0] w_asqrt28_18;
	wire [2:0] w_asqrt28_19;
	wire [2:0] w_asqrt28_20;
	wire [2:0] w_asqrt28_21;
	wire [2:0] w_asqrt28_22;
	wire [2:0] w_asqrt28_23;
	wire [2:0] w_asqrt28_24;
	wire [2:0] w_asqrt28_25;
	wire [2:0] w_asqrt28_26;
	wire [2:0] w_asqrt28_27;
	wire [2:0] w_asqrt28_28;
	wire [2:0] w_asqrt28_29;
	wire [2:0] w_asqrt28_30;
	wire w_asqrt28_31;
	wire asqrt_fa_28;
	wire [2:0] w_asqrt29_0;
	wire [2:0] w_asqrt29_1;
	wire [2:0] w_asqrt29_2;
	wire [2:0] w_asqrt29_3;
	wire [2:0] w_asqrt29_4;
	wire [2:0] w_asqrt29_5;
	wire [2:0] w_asqrt29_6;
	wire [2:0] w_asqrt29_7;
	wire [2:0] w_asqrt29_8;
	wire [2:0] w_asqrt29_9;
	wire [2:0] w_asqrt29_10;
	wire [2:0] w_asqrt29_11;
	wire [2:0] w_asqrt29_12;
	wire [2:0] w_asqrt29_13;
	wire [2:0] w_asqrt29_14;
	wire [2:0] w_asqrt29_15;
	wire [2:0] w_asqrt29_16;
	wire [2:0] w_asqrt29_17;
	wire [2:0] w_asqrt29_18;
	wire [2:0] w_asqrt29_19;
	wire [2:0] w_asqrt29_20;
	wire [1:0] w_asqrt29_21;
	wire asqrt_fa_29;
	wire [2:0] w_asqrt30_0;
	wire [2:0] w_asqrt30_1;
	wire [2:0] w_asqrt30_2;
	wire [2:0] w_asqrt30_3;
	wire [2:0] w_asqrt30_4;
	wire [2:0] w_asqrt30_5;
	wire [2:0] w_asqrt30_6;
	wire [2:0] w_asqrt30_7;
	wire [2:0] w_asqrt30_8;
	wire [2:0] w_asqrt30_9;
	wire [2:0] w_asqrt30_10;
	wire [2:0] w_asqrt30_11;
	wire [2:0] w_asqrt30_12;
	wire [2:0] w_asqrt30_13;
	wire [2:0] w_asqrt30_14;
	wire [2:0] w_asqrt30_15;
	wire [2:0] w_asqrt30_16;
	wire [2:0] w_asqrt30_17;
	wire [2:0] w_asqrt30_18;
	wire [2:0] w_asqrt30_19;
	wire [2:0] w_asqrt30_20;
	wire [2:0] w_asqrt30_21;
	wire [2:0] w_asqrt30_22;
	wire [2:0] w_asqrt30_23;
	wire [2:0] w_asqrt30_24;
	wire [2:0] w_asqrt30_25;
	wire [2:0] w_asqrt30_26;
	wire [2:0] w_asqrt30_27;
	wire [2:0] w_asqrt30_28;
	wire [2:0] w_asqrt30_29;
	wire [2:0] w_asqrt30_30;
	wire w_asqrt30_31;
	wire asqrt_fa_30;
	wire [2:0] w_asqrt31_0;
	wire [2:0] w_asqrt31_1;
	wire [2:0] w_asqrt31_2;
	wire [2:0] w_asqrt31_3;
	wire [2:0] w_asqrt31_4;
	wire [2:0] w_asqrt31_5;
	wire [2:0] w_asqrt31_6;
	wire [2:0] w_asqrt31_7;
	wire [2:0] w_asqrt31_8;
	wire [2:0] w_asqrt31_9;
	wire [2:0] w_asqrt31_10;
	wire [2:0] w_asqrt31_11;
	wire [2:0] w_asqrt31_12;
	wire [2:0] w_asqrt31_13;
	wire [2:0] w_asqrt31_14;
	wire [2:0] w_asqrt31_15;
	wire [2:0] w_asqrt31_16;
	wire [2:0] w_asqrt31_17;
	wire [2:0] w_asqrt31_18;
	wire [2:0] w_asqrt31_19;
	wire [2:0] w_asqrt31_20;
	wire [1:0] w_asqrt31_21;
	wire asqrt_fa_31;
	wire [2:0] w_asqrt32_0;
	wire [2:0] w_asqrt32_1;
	wire [2:0] w_asqrt32_2;
	wire [2:0] w_asqrt32_3;
	wire [2:0] w_asqrt32_4;
	wire [2:0] w_asqrt32_5;
	wire [2:0] w_asqrt32_6;
	wire [2:0] w_asqrt32_7;
	wire [2:0] w_asqrt32_8;
	wire [2:0] w_asqrt32_9;
	wire [2:0] w_asqrt32_10;
	wire [2:0] w_asqrt32_11;
	wire [2:0] w_asqrt32_12;
	wire [2:0] w_asqrt32_13;
	wire [2:0] w_asqrt32_14;
	wire [2:0] w_asqrt32_15;
	wire [2:0] w_asqrt32_16;
	wire [2:0] w_asqrt32_17;
	wire [2:0] w_asqrt32_18;
	wire [2:0] w_asqrt32_19;
	wire [2:0] w_asqrt32_20;
	wire [2:0] w_asqrt32_21;
	wire [2:0] w_asqrt32_22;
	wire [2:0] w_asqrt32_23;
	wire [2:0] w_asqrt32_24;
	wire [2:0] w_asqrt32_25;
	wire [2:0] w_asqrt32_26;
	wire [2:0] w_asqrt32_27;
	wire [2:0] w_asqrt32_28;
	wire [2:0] w_asqrt32_29;
	wire [2:0] w_asqrt32_30;
	wire w_asqrt32_31;
	wire asqrt_fa_32;
	wire [2:0] w_asqrt33_0;
	wire [2:0] w_asqrt33_1;
	wire [2:0] w_asqrt33_2;
	wire [2:0] w_asqrt33_3;
	wire [2:0] w_asqrt33_4;
	wire [2:0] w_asqrt33_5;
	wire [2:0] w_asqrt33_6;
	wire [2:0] w_asqrt33_7;
	wire [2:0] w_asqrt33_8;
	wire [2:0] w_asqrt33_9;
	wire [2:0] w_asqrt33_10;
	wire [2:0] w_asqrt33_11;
	wire [2:0] w_asqrt33_12;
	wire [2:0] w_asqrt33_13;
	wire [2:0] w_asqrt33_14;
	wire [2:0] w_asqrt33_15;
	wire [2:0] w_asqrt33_16;
	wire [2:0] w_asqrt33_17;
	wire [2:0] w_asqrt33_18;
	wire [2:0] w_asqrt33_19;
	wire [2:0] w_asqrt33_20;
	wire [2:0] w_asqrt33_21;
	wire [1:0] w_asqrt33_22;
	wire asqrt_fa_33;
	wire [2:0] w_asqrt34_0;
	wire [2:0] w_asqrt34_1;
	wire [2:0] w_asqrt34_2;
	wire [2:0] w_asqrt34_3;
	wire [2:0] w_asqrt34_4;
	wire [2:0] w_asqrt34_5;
	wire [2:0] w_asqrt34_6;
	wire [2:0] w_asqrt34_7;
	wire [2:0] w_asqrt34_8;
	wire [2:0] w_asqrt34_9;
	wire [2:0] w_asqrt34_10;
	wire [2:0] w_asqrt34_11;
	wire [2:0] w_asqrt34_12;
	wire [2:0] w_asqrt34_13;
	wire [2:0] w_asqrt34_14;
	wire [2:0] w_asqrt34_15;
	wire [2:0] w_asqrt34_16;
	wire [2:0] w_asqrt34_17;
	wire [2:0] w_asqrt34_18;
	wire [2:0] w_asqrt34_19;
	wire [2:0] w_asqrt34_20;
	wire [2:0] w_asqrt34_21;
	wire [2:0] w_asqrt34_22;
	wire [2:0] w_asqrt34_23;
	wire [2:0] w_asqrt34_24;
	wire [2:0] w_asqrt34_25;
	wire [2:0] w_asqrt34_26;
	wire [2:0] w_asqrt34_27;
	wire [2:0] w_asqrt34_28;
	wire [2:0] w_asqrt34_29;
	wire [2:0] w_asqrt34_30;
	wire w_asqrt34_31;
	wire asqrt_fa_34;
	wire [2:0] w_asqrt35_0;
	wire [2:0] w_asqrt35_1;
	wire [2:0] w_asqrt35_2;
	wire [2:0] w_asqrt35_3;
	wire [2:0] w_asqrt35_4;
	wire [2:0] w_asqrt35_5;
	wire [2:0] w_asqrt35_6;
	wire [2:0] w_asqrt35_7;
	wire [2:0] w_asqrt35_8;
	wire [2:0] w_asqrt35_9;
	wire [2:0] w_asqrt35_10;
	wire [2:0] w_asqrt35_11;
	wire [2:0] w_asqrt35_12;
	wire [2:0] w_asqrt35_13;
	wire [2:0] w_asqrt35_14;
	wire [2:0] w_asqrt35_15;
	wire [2:0] w_asqrt35_16;
	wire [2:0] w_asqrt35_17;
	wire [2:0] w_asqrt35_18;
	wire [2:0] w_asqrt35_19;
	wire [2:0] w_asqrt35_20;
	wire [2:0] w_asqrt35_21;
	wire [1:0] w_asqrt35_22;
	wire asqrt_fa_35;
	wire [2:0] w_asqrt36_0;
	wire [2:0] w_asqrt36_1;
	wire [2:0] w_asqrt36_2;
	wire [2:0] w_asqrt36_3;
	wire [2:0] w_asqrt36_4;
	wire [2:0] w_asqrt36_5;
	wire [2:0] w_asqrt36_6;
	wire [2:0] w_asqrt36_7;
	wire [2:0] w_asqrt36_8;
	wire [2:0] w_asqrt36_9;
	wire [2:0] w_asqrt36_10;
	wire [2:0] w_asqrt36_11;
	wire [2:0] w_asqrt36_12;
	wire [2:0] w_asqrt36_13;
	wire [2:0] w_asqrt36_14;
	wire [2:0] w_asqrt36_15;
	wire [2:0] w_asqrt36_16;
	wire [2:0] w_asqrt36_17;
	wire [2:0] w_asqrt36_18;
	wire [2:0] w_asqrt36_19;
	wire [2:0] w_asqrt36_20;
	wire [2:0] w_asqrt36_21;
	wire [2:0] w_asqrt36_22;
	wire [2:0] w_asqrt36_23;
	wire [2:0] w_asqrt36_24;
	wire [2:0] w_asqrt36_25;
	wire [2:0] w_asqrt36_26;
	wire [2:0] w_asqrt36_27;
	wire [2:0] w_asqrt36_28;
	wire [2:0] w_asqrt36_29;
	wire [2:0] w_asqrt36_30;
	wire w_asqrt36_31;
	wire asqrt_fa_36;
	wire [2:0] w_asqrt37_0;
	wire [2:0] w_asqrt37_1;
	wire [2:0] w_asqrt37_2;
	wire [2:0] w_asqrt37_3;
	wire [2:0] w_asqrt37_4;
	wire [2:0] w_asqrt37_5;
	wire [2:0] w_asqrt37_6;
	wire [2:0] w_asqrt37_7;
	wire [2:0] w_asqrt37_8;
	wire [2:0] w_asqrt37_9;
	wire [2:0] w_asqrt37_10;
	wire [2:0] w_asqrt37_11;
	wire [2:0] w_asqrt37_12;
	wire [2:0] w_asqrt37_13;
	wire [2:0] w_asqrt37_14;
	wire [2:0] w_asqrt37_15;
	wire [2:0] w_asqrt37_16;
	wire [2:0] w_asqrt37_17;
	wire [2:0] w_asqrt37_18;
	wire [2:0] w_asqrt37_19;
	wire [2:0] w_asqrt37_20;
	wire [2:0] w_asqrt37_21;
	wire [2:0] w_asqrt37_22;
	wire [1:0] w_asqrt37_23;
	wire asqrt_fa_37;
	wire [2:0] w_asqrt38_0;
	wire [2:0] w_asqrt38_1;
	wire [2:0] w_asqrt38_2;
	wire [2:0] w_asqrt38_3;
	wire [2:0] w_asqrt38_4;
	wire [2:0] w_asqrt38_5;
	wire [2:0] w_asqrt38_6;
	wire [2:0] w_asqrt38_7;
	wire [2:0] w_asqrt38_8;
	wire [2:0] w_asqrt38_9;
	wire [2:0] w_asqrt38_10;
	wire [2:0] w_asqrt38_11;
	wire [2:0] w_asqrt38_12;
	wire [2:0] w_asqrt38_13;
	wire [2:0] w_asqrt38_14;
	wire [2:0] w_asqrt38_15;
	wire [2:0] w_asqrt38_16;
	wire [2:0] w_asqrt38_17;
	wire [2:0] w_asqrt38_18;
	wire [2:0] w_asqrt38_19;
	wire [2:0] w_asqrt38_20;
	wire [2:0] w_asqrt38_21;
	wire [2:0] w_asqrt38_22;
	wire [2:0] w_asqrt38_23;
	wire [2:0] w_asqrt38_24;
	wire [2:0] w_asqrt38_25;
	wire [2:0] w_asqrt38_26;
	wire [2:0] w_asqrt38_27;
	wire [2:0] w_asqrt38_28;
	wire [2:0] w_asqrt38_29;
	wire [2:0] w_asqrt38_30;
	wire w_asqrt38_31;
	wire asqrt_fa_38;
	wire [2:0] w_asqrt39_0;
	wire [2:0] w_asqrt39_1;
	wire [2:0] w_asqrt39_2;
	wire [2:0] w_asqrt39_3;
	wire [2:0] w_asqrt39_4;
	wire [2:0] w_asqrt39_5;
	wire [2:0] w_asqrt39_6;
	wire [2:0] w_asqrt39_7;
	wire [2:0] w_asqrt39_8;
	wire [2:0] w_asqrt39_9;
	wire [2:0] w_asqrt39_10;
	wire [2:0] w_asqrt39_11;
	wire [2:0] w_asqrt39_12;
	wire [2:0] w_asqrt39_13;
	wire [2:0] w_asqrt39_14;
	wire [2:0] w_asqrt39_15;
	wire [2:0] w_asqrt39_16;
	wire [2:0] w_asqrt39_17;
	wire [2:0] w_asqrt39_18;
	wire [2:0] w_asqrt39_19;
	wire [2:0] w_asqrt39_20;
	wire [2:0] w_asqrt39_21;
	wire [2:0] w_asqrt39_22;
	wire [1:0] w_asqrt39_23;
	wire asqrt_fa_39;
	wire [2:0] w_asqrt40_0;
	wire [2:0] w_asqrt40_1;
	wire [2:0] w_asqrt40_2;
	wire [2:0] w_asqrt40_3;
	wire [2:0] w_asqrt40_4;
	wire [2:0] w_asqrt40_5;
	wire [2:0] w_asqrt40_6;
	wire [2:0] w_asqrt40_7;
	wire [2:0] w_asqrt40_8;
	wire [2:0] w_asqrt40_9;
	wire [2:0] w_asqrt40_10;
	wire [2:0] w_asqrt40_11;
	wire [2:0] w_asqrt40_12;
	wire [2:0] w_asqrt40_13;
	wire [2:0] w_asqrt40_14;
	wire [2:0] w_asqrt40_15;
	wire [2:0] w_asqrt40_16;
	wire [2:0] w_asqrt40_17;
	wire [2:0] w_asqrt40_18;
	wire [2:0] w_asqrt40_19;
	wire [2:0] w_asqrt40_20;
	wire [2:0] w_asqrt40_21;
	wire [2:0] w_asqrt40_22;
	wire [2:0] w_asqrt40_23;
	wire [2:0] w_asqrt40_24;
	wire [2:0] w_asqrt40_25;
	wire [2:0] w_asqrt40_26;
	wire [2:0] w_asqrt40_27;
	wire [2:0] w_asqrt40_28;
	wire [2:0] w_asqrt40_29;
	wire [2:0] w_asqrt40_30;
	wire w_asqrt40_31;
	wire asqrt_fa_40;
	wire [2:0] w_asqrt41_0;
	wire [2:0] w_asqrt41_1;
	wire [2:0] w_asqrt41_2;
	wire [2:0] w_asqrt41_3;
	wire [2:0] w_asqrt41_4;
	wire [2:0] w_asqrt41_5;
	wire [2:0] w_asqrt41_6;
	wire [2:0] w_asqrt41_7;
	wire [2:0] w_asqrt41_8;
	wire [2:0] w_asqrt41_9;
	wire [2:0] w_asqrt41_10;
	wire [2:0] w_asqrt41_11;
	wire [2:0] w_asqrt41_12;
	wire [2:0] w_asqrt41_13;
	wire [2:0] w_asqrt41_14;
	wire [2:0] w_asqrt41_15;
	wire [2:0] w_asqrt41_16;
	wire [2:0] w_asqrt41_17;
	wire [2:0] w_asqrt41_18;
	wire [2:0] w_asqrt41_19;
	wire [2:0] w_asqrt41_20;
	wire [2:0] w_asqrt41_21;
	wire [2:0] w_asqrt41_22;
	wire [2:0] w_asqrt41_23;
	wire [1:0] w_asqrt41_24;
	wire asqrt_fa_41;
	wire [2:0] w_asqrt42_0;
	wire [2:0] w_asqrt42_1;
	wire [2:0] w_asqrt42_2;
	wire [2:0] w_asqrt42_3;
	wire [2:0] w_asqrt42_4;
	wire [2:0] w_asqrt42_5;
	wire [2:0] w_asqrt42_6;
	wire [2:0] w_asqrt42_7;
	wire [2:0] w_asqrt42_8;
	wire [2:0] w_asqrt42_9;
	wire [2:0] w_asqrt42_10;
	wire [2:0] w_asqrt42_11;
	wire [2:0] w_asqrt42_12;
	wire [2:0] w_asqrt42_13;
	wire [2:0] w_asqrt42_14;
	wire [2:0] w_asqrt42_15;
	wire [2:0] w_asqrt42_16;
	wire [2:0] w_asqrt42_17;
	wire [2:0] w_asqrt42_18;
	wire [2:0] w_asqrt42_19;
	wire [2:0] w_asqrt42_20;
	wire [2:0] w_asqrt42_21;
	wire [2:0] w_asqrt42_22;
	wire [2:0] w_asqrt42_23;
	wire [2:0] w_asqrt42_24;
	wire [2:0] w_asqrt42_25;
	wire [2:0] w_asqrt42_26;
	wire [2:0] w_asqrt42_27;
	wire [2:0] w_asqrt42_28;
	wire [2:0] w_asqrt42_29;
	wire [2:0] w_asqrt42_30;
	wire w_asqrt42_31;
	wire asqrt_fa_42;
	wire [2:0] w_asqrt43_0;
	wire [2:0] w_asqrt43_1;
	wire [2:0] w_asqrt43_2;
	wire [2:0] w_asqrt43_3;
	wire [2:0] w_asqrt43_4;
	wire [2:0] w_asqrt43_5;
	wire [2:0] w_asqrt43_6;
	wire [2:0] w_asqrt43_7;
	wire [2:0] w_asqrt43_8;
	wire [2:0] w_asqrt43_9;
	wire [2:0] w_asqrt43_10;
	wire [2:0] w_asqrt43_11;
	wire [2:0] w_asqrt43_12;
	wire [2:0] w_asqrt43_13;
	wire [2:0] w_asqrt43_14;
	wire [2:0] w_asqrt43_15;
	wire [2:0] w_asqrt43_16;
	wire [2:0] w_asqrt43_17;
	wire [2:0] w_asqrt43_18;
	wire [2:0] w_asqrt43_19;
	wire [2:0] w_asqrt43_20;
	wire [2:0] w_asqrt43_21;
	wire [2:0] w_asqrt43_22;
	wire [2:0] w_asqrt43_23;
	wire [1:0] w_asqrt43_24;
	wire asqrt_fa_43;
	wire [2:0] w_asqrt44_0;
	wire [2:0] w_asqrt44_1;
	wire [2:0] w_asqrt44_2;
	wire [2:0] w_asqrt44_3;
	wire [2:0] w_asqrt44_4;
	wire [2:0] w_asqrt44_5;
	wire [2:0] w_asqrt44_6;
	wire [2:0] w_asqrt44_7;
	wire [2:0] w_asqrt44_8;
	wire [2:0] w_asqrt44_9;
	wire [2:0] w_asqrt44_10;
	wire [2:0] w_asqrt44_11;
	wire [2:0] w_asqrt44_12;
	wire [2:0] w_asqrt44_13;
	wire [2:0] w_asqrt44_14;
	wire [2:0] w_asqrt44_15;
	wire [2:0] w_asqrt44_16;
	wire [2:0] w_asqrt44_17;
	wire [2:0] w_asqrt44_18;
	wire [2:0] w_asqrt44_19;
	wire [2:0] w_asqrt44_20;
	wire [2:0] w_asqrt44_21;
	wire [2:0] w_asqrt44_22;
	wire [2:0] w_asqrt44_23;
	wire [2:0] w_asqrt44_24;
	wire [2:0] w_asqrt44_25;
	wire [2:0] w_asqrt44_26;
	wire [2:0] w_asqrt44_27;
	wire [2:0] w_asqrt44_28;
	wire [2:0] w_asqrt44_29;
	wire [2:0] w_asqrt44_30;
	wire w_asqrt44_31;
	wire asqrt_fa_44;
	wire [2:0] w_asqrt45_0;
	wire [2:0] w_asqrt45_1;
	wire [2:0] w_asqrt45_2;
	wire [2:0] w_asqrt45_3;
	wire [2:0] w_asqrt45_4;
	wire [2:0] w_asqrt45_5;
	wire [2:0] w_asqrt45_6;
	wire [2:0] w_asqrt45_7;
	wire [2:0] w_asqrt45_8;
	wire [2:0] w_asqrt45_9;
	wire [2:0] w_asqrt45_10;
	wire [2:0] w_asqrt45_11;
	wire [2:0] w_asqrt45_12;
	wire [2:0] w_asqrt45_13;
	wire [2:0] w_asqrt45_14;
	wire [2:0] w_asqrt45_15;
	wire [2:0] w_asqrt45_16;
	wire [2:0] w_asqrt45_17;
	wire [2:0] w_asqrt45_18;
	wire [2:0] w_asqrt45_19;
	wire [2:0] w_asqrt45_20;
	wire [2:0] w_asqrt45_21;
	wire [2:0] w_asqrt45_22;
	wire [2:0] w_asqrt45_23;
	wire [2:0] w_asqrt45_24;
	wire [1:0] w_asqrt45_25;
	wire asqrt_fa_45;
	wire [2:0] w_asqrt46_0;
	wire [2:0] w_asqrt46_1;
	wire [2:0] w_asqrt46_2;
	wire [2:0] w_asqrt46_3;
	wire [2:0] w_asqrt46_4;
	wire [2:0] w_asqrt46_5;
	wire [2:0] w_asqrt46_6;
	wire [2:0] w_asqrt46_7;
	wire [2:0] w_asqrt46_8;
	wire [2:0] w_asqrt46_9;
	wire [2:0] w_asqrt46_10;
	wire [2:0] w_asqrt46_11;
	wire [2:0] w_asqrt46_12;
	wire [2:0] w_asqrt46_13;
	wire [2:0] w_asqrt46_14;
	wire [2:0] w_asqrt46_15;
	wire [2:0] w_asqrt46_16;
	wire [2:0] w_asqrt46_17;
	wire [2:0] w_asqrt46_18;
	wire [2:0] w_asqrt46_19;
	wire [2:0] w_asqrt46_20;
	wire [2:0] w_asqrt46_21;
	wire [2:0] w_asqrt46_22;
	wire [2:0] w_asqrt46_23;
	wire [2:0] w_asqrt46_24;
	wire [2:0] w_asqrt46_25;
	wire [2:0] w_asqrt46_26;
	wire [2:0] w_asqrt46_27;
	wire [2:0] w_asqrt46_28;
	wire [2:0] w_asqrt46_29;
	wire [2:0] w_asqrt46_30;
	wire w_asqrt46_31;
	wire asqrt_fa_46;
	wire [2:0] w_asqrt47_0;
	wire [2:0] w_asqrt47_1;
	wire [2:0] w_asqrt47_2;
	wire [2:0] w_asqrt47_3;
	wire [2:0] w_asqrt47_4;
	wire [2:0] w_asqrt47_5;
	wire [2:0] w_asqrt47_6;
	wire [2:0] w_asqrt47_7;
	wire [2:0] w_asqrt47_8;
	wire [2:0] w_asqrt47_9;
	wire [2:0] w_asqrt47_10;
	wire [2:0] w_asqrt47_11;
	wire [2:0] w_asqrt47_12;
	wire [2:0] w_asqrt47_13;
	wire [2:0] w_asqrt47_14;
	wire [2:0] w_asqrt47_15;
	wire [2:0] w_asqrt47_16;
	wire [2:0] w_asqrt47_17;
	wire [2:0] w_asqrt47_18;
	wire [2:0] w_asqrt47_19;
	wire [2:0] w_asqrt47_20;
	wire [2:0] w_asqrt47_21;
	wire [2:0] w_asqrt47_22;
	wire [2:0] w_asqrt47_23;
	wire [2:0] w_asqrt47_24;
	wire [1:0] w_asqrt47_25;
	wire asqrt_fa_47;
	wire [2:0] w_asqrt48_0;
	wire [2:0] w_asqrt48_1;
	wire [2:0] w_asqrt48_2;
	wire [2:0] w_asqrt48_3;
	wire [2:0] w_asqrt48_4;
	wire [2:0] w_asqrt48_5;
	wire [2:0] w_asqrt48_6;
	wire [2:0] w_asqrt48_7;
	wire [2:0] w_asqrt48_8;
	wire [2:0] w_asqrt48_9;
	wire [2:0] w_asqrt48_10;
	wire [2:0] w_asqrt48_11;
	wire [2:0] w_asqrt48_12;
	wire [2:0] w_asqrt48_13;
	wire [2:0] w_asqrt48_14;
	wire [2:0] w_asqrt48_15;
	wire [2:0] w_asqrt48_16;
	wire [2:0] w_asqrt48_17;
	wire [2:0] w_asqrt48_18;
	wire [2:0] w_asqrt48_19;
	wire [2:0] w_asqrt48_20;
	wire [2:0] w_asqrt48_21;
	wire [2:0] w_asqrt48_22;
	wire [2:0] w_asqrt48_23;
	wire [2:0] w_asqrt48_24;
	wire [2:0] w_asqrt48_25;
	wire [2:0] w_asqrt48_26;
	wire [2:0] w_asqrt48_27;
	wire [2:0] w_asqrt48_28;
	wire [2:0] w_asqrt48_29;
	wire [2:0] w_asqrt48_30;
	wire w_asqrt48_31;
	wire asqrt_fa_48;
	wire [2:0] w_asqrt49_0;
	wire [2:0] w_asqrt49_1;
	wire [2:0] w_asqrt49_2;
	wire [2:0] w_asqrt49_3;
	wire [2:0] w_asqrt49_4;
	wire [2:0] w_asqrt49_5;
	wire [2:0] w_asqrt49_6;
	wire [2:0] w_asqrt49_7;
	wire [2:0] w_asqrt49_8;
	wire [2:0] w_asqrt49_9;
	wire [2:0] w_asqrt49_10;
	wire [2:0] w_asqrt49_11;
	wire [2:0] w_asqrt49_12;
	wire [2:0] w_asqrt49_13;
	wire [2:0] w_asqrt49_14;
	wire [2:0] w_asqrt49_15;
	wire [2:0] w_asqrt49_16;
	wire [2:0] w_asqrt49_17;
	wire [2:0] w_asqrt49_18;
	wire [2:0] w_asqrt49_19;
	wire [2:0] w_asqrt49_20;
	wire [2:0] w_asqrt49_21;
	wire [2:0] w_asqrt49_22;
	wire [2:0] w_asqrt49_23;
	wire [2:0] w_asqrt49_24;
	wire [2:0] w_asqrt49_25;
	wire [1:0] w_asqrt49_26;
	wire asqrt_fa_49;
	wire [2:0] w_asqrt50_0;
	wire [2:0] w_asqrt50_1;
	wire [2:0] w_asqrt50_2;
	wire [2:0] w_asqrt50_3;
	wire [2:0] w_asqrt50_4;
	wire [2:0] w_asqrt50_5;
	wire [2:0] w_asqrt50_6;
	wire [2:0] w_asqrt50_7;
	wire [2:0] w_asqrt50_8;
	wire [2:0] w_asqrt50_9;
	wire [2:0] w_asqrt50_10;
	wire [2:0] w_asqrt50_11;
	wire [2:0] w_asqrt50_12;
	wire [2:0] w_asqrt50_13;
	wire [2:0] w_asqrt50_14;
	wire [2:0] w_asqrt50_15;
	wire [2:0] w_asqrt50_16;
	wire [2:0] w_asqrt50_17;
	wire [2:0] w_asqrt50_18;
	wire [2:0] w_asqrt50_19;
	wire [2:0] w_asqrt50_20;
	wire [2:0] w_asqrt50_21;
	wire [2:0] w_asqrt50_22;
	wire [2:0] w_asqrt50_23;
	wire [2:0] w_asqrt50_24;
	wire [2:0] w_asqrt50_25;
	wire [2:0] w_asqrt50_26;
	wire [2:0] w_asqrt50_27;
	wire [2:0] w_asqrt50_28;
	wire [2:0] w_asqrt50_29;
	wire [2:0] w_asqrt50_30;
	wire w_asqrt50_31;
	wire asqrt_fa_50;
	wire [2:0] w_asqrt51_0;
	wire [2:0] w_asqrt51_1;
	wire [2:0] w_asqrt51_2;
	wire [2:0] w_asqrt51_3;
	wire [2:0] w_asqrt51_4;
	wire [2:0] w_asqrt51_5;
	wire [2:0] w_asqrt51_6;
	wire [2:0] w_asqrt51_7;
	wire [2:0] w_asqrt51_8;
	wire [2:0] w_asqrt51_9;
	wire [2:0] w_asqrt51_10;
	wire [2:0] w_asqrt51_11;
	wire [2:0] w_asqrt51_12;
	wire [2:0] w_asqrt51_13;
	wire [2:0] w_asqrt51_14;
	wire [2:0] w_asqrt51_15;
	wire [2:0] w_asqrt51_16;
	wire [2:0] w_asqrt51_17;
	wire [2:0] w_asqrt51_18;
	wire [2:0] w_asqrt51_19;
	wire [2:0] w_asqrt51_20;
	wire [2:0] w_asqrt51_21;
	wire [2:0] w_asqrt51_22;
	wire [2:0] w_asqrt51_23;
	wire [2:0] w_asqrt51_24;
	wire [2:0] w_asqrt51_25;
	wire [1:0] w_asqrt51_26;
	wire asqrt_fa_51;
	wire [2:0] w_asqrt52_0;
	wire [2:0] w_asqrt52_1;
	wire [2:0] w_asqrt52_2;
	wire [2:0] w_asqrt52_3;
	wire [2:0] w_asqrt52_4;
	wire [2:0] w_asqrt52_5;
	wire [2:0] w_asqrt52_6;
	wire [2:0] w_asqrt52_7;
	wire [2:0] w_asqrt52_8;
	wire [2:0] w_asqrt52_9;
	wire [2:0] w_asqrt52_10;
	wire [2:0] w_asqrt52_11;
	wire [2:0] w_asqrt52_12;
	wire [2:0] w_asqrt52_13;
	wire [2:0] w_asqrt52_14;
	wire [2:0] w_asqrt52_15;
	wire [2:0] w_asqrt52_16;
	wire [2:0] w_asqrt52_17;
	wire [2:0] w_asqrt52_18;
	wire [2:0] w_asqrt52_19;
	wire [2:0] w_asqrt52_20;
	wire [2:0] w_asqrt52_21;
	wire [2:0] w_asqrt52_22;
	wire [2:0] w_asqrt52_23;
	wire [2:0] w_asqrt52_24;
	wire [2:0] w_asqrt52_25;
	wire [2:0] w_asqrt52_26;
	wire [2:0] w_asqrt52_27;
	wire [2:0] w_asqrt52_28;
	wire [2:0] w_asqrt52_29;
	wire [2:0] w_asqrt52_30;
	wire w_asqrt52_31;
	wire asqrt_fa_52;
	wire [2:0] w_asqrt53_0;
	wire [2:0] w_asqrt53_1;
	wire [2:0] w_asqrt53_2;
	wire [2:0] w_asqrt53_3;
	wire [2:0] w_asqrt53_4;
	wire [2:0] w_asqrt53_5;
	wire [2:0] w_asqrt53_6;
	wire [2:0] w_asqrt53_7;
	wire [2:0] w_asqrt53_8;
	wire [2:0] w_asqrt53_9;
	wire [2:0] w_asqrt53_10;
	wire [2:0] w_asqrt53_11;
	wire [2:0] w_asqrt53_12;
	wire [2:0] w_asqrt53_13;
	wire [2:0] w_asqrt53_14;
	wire [2:0] w_asqrt53_15;
	wire [2:0] w_asqrt53_16;
	wire [2:0] w_asqrt53_17;
	wire [2:0] w_asqrt53_18;
	wire [2:0] w_asqrt53_19;
	wire [2:0] w_asqrt53_20;
	wire [2:0] w_asqrt53_21;
	wire [2:0] w_asqrt53_22;
	wire [2:0] w_asqrt53_23;
	wire [2:0] w_asqrt53_24;
	wire [2:0] w_asqrt53_25;
	wire [2:0] w_asqrt53_26;
	wire [1:0] w_asqrt53_27;
	wire asqrt_fa_53;
	wire [2:0] w_asqrt54_0;
	wire [2:0] w_asqrt54_1;
	wire [2:0] w_asqrt54_2;
	wire [2:0] w_asqrt54_3;
	wire [2:0] w_asqrt54_4;
	wire [2:0] w_asqrt54_5;
	wire [2:0] w_asqrt54_6;
	wire [2:0] w_asqrt54_7;
	wire [2:0] w_asqrt54_8;
	wire [2:0] w_asqrt54_9;
	wire [2:0] w_asqrt54_10;
	wire [2:0] w_asqrt54_11;
	wire [2:0] w_asqrt54_12;
	wire [2:0] w_asqrt54_13;
	wire [2:0] w_asqrt54_14;
	wire [2:0] w_asqrt54_15;
	wire [2:0] w_asqrt54_16;
	wire [2:0] w_asqrt54_17;
	wire [2:0] w_asqrt54_18;
	wire [2:0] w_asqrt54_19;
	wire [2:0] w_asqrt54_20;
	wire [2:0] w_asqrt54_21;
	wire [2:0] w_asqrt54_22;
	wire [2:0] w_asqrt54_23;
	wire [2:0] w_asqrt54_24;
	wire [2:0] w_asqrt54_25;
	wire [2:0] w_asqrt54_26;
	wire [2:0] w_asqrt54_27;
	wire [2:0] w_asqrt54_28;
	wire [2:0] w_asqrt54_29;
	wire [2:0] w_asqrt54_30;
	wire w_asqrt54_31;
	wire asqrt_fa_54;
	wire [2:0] w_asqrt55_0;
	wire [2:0] w_asqrt55_1;
	wire [2:0] w_asqrt55_2;
	wire [2:0] w_asqrt55_3;
	wire [2:0] w_asqrt55_4;
	wire [2:0] w_asqrt55_5;
	wire [2:0] w_asqrt55_6;
	wire [2:0] w_asqrt55_7;
	wire [2:0] w_asqrt55_8;
	wire [2:0] w_asqrt55_9;
	wire [2:0] w_asqrt55_10;
	wire [2:0] w_asqrt55_11;
	wire [2:0] w_asqrt55_12;
	wire [2:0] w_asqrt55_13;
	wire [2:0] w_asqrt55_14;
	wire [2:0] w_asqrt55_15;
	wire [2:0] w_asqrt55_16;
	wire [2:0] w_asqrt55_17;
	wire [2:0] w_asqrt55_18;
	wire [2:0] w_asqrt55_19;
	wire [2:0] w_asqrt55_20;
	wire [2:0] w_asqrt55_21;
	wire [2:0] w_asqrt55_22;
	wire [2:0] w_asqrt55_23;
	wire [2:0] w_asqrt55_24;
	wire [2:0] w_asqrt55_25;
	wire [2:0] w_asqrt55_26;
	wire [2:0] w_asqrt55_27;
	wire w_asqrt55_28;
	wire asqrt_fa_55;
	wire [2:0] w_asqrt56_0;
	wire [2:0] w_asqrt56_1;
	wire [2:0] w_asqrt56_2;
	wire [2:0] w_asqrt56_3;
	wire [2:0] w_asqrt56_4;
	wire [2:0] w_asqrt56_5;
	wire [2:0] w_asqrt56_6;
	wire [2:0] w_asqrt56_7;
	wire [2:0] w_asqrt56_8;
	wire [2:0] w_asqrt56_9;
	wire [2:0] w_asqrt56_10;
	wire [2:0] w_asqrt56_11;
	wire [2:0] w_asqrt56_12;
	wire [2:0] w_asqrt56_13;
	wire [2:0] w_asqrt56_14;
	wire [2:0] w_asqrt56_15;
	wire [2:0] w_asqrt56_16;
	wire [2:0] w_asqrt56_17;
	wire [2:0] w_asqrt56_18;
	wire [2:0] w_asqrt56_19;
	wire [2:0] w_asqrt56_20;
	wire [2:0] w_asqrt56_21;
	wire [2:0] w_asqrt56_22;
	wire [2:0] w_asqrt56_23;
	wire [2:0] w_asqrt56_24;
	wire [2:0] w_asqrt56_25;
	wire [2:0] w_asqrt56_26;
	wire [2:0] w_asqrt56_27;
	wire [2:0] w_asqrt56_28;
	wire [2:0] w_asqrt56_29;
	wire [2:0] w_asqrt56_30;
	wire w_asqrt56_31;
	wire asqrt_fa_56;
	wire [2:0] w_asqrt57_0;
	wire [2:0] w_asqrt57_1;
	wire [2:0] w_asqrt57_2;
	wire [2:0] w_asqrt57_3;
	wire [2:0] w_asqrt57_4;
	wire [2:0] w_asqrt57_5;
	wire [2:0] w_asqrt57_6;
	wire [2:0] w_asqrt57_7;
	wire [2:0] w_asqrt57_8;
	wire [2:0] w_asqrt57_9;
	wire [2:0] w_asqrt57_10;
	wire [2:0] w_asqrt57_11;
	wire [2:0] w_asqrt57_12;
	wire [2:0] w_asqrt57_13;
	wire [2:0] w_asqrt57_14;
	wire [2:0] w_asqrt57_15;
	wire [2:0] w_asqrt57_16;
	wire [2:0] w_asqrt57_17;
	wire [2:0] w_asqrt57_18;
	wire [2:0] w_asqrt57_19;
	wire [2:0] w_asqrt57_20;
	wire [2:0] w_asqrt57_21;
	wire [2:0] w_asqrt57_22;
	wire [2:0] w_asqrt57_23;
	wire [2:0] w_asqrt57_24;
	wire [2:0] w_asqrt57_25;
	wire [2:0] w_asqrt57_26;
	wire [2:0] w_asqrt57_27;
	wire [2:0] w_asqrt57_28;
	wire w_asqrt57_29;
	wire asqrt_fa_57;
	wire [2:0] w_asqrt58_0;
	wire [2:0] w_asqrt58_1;
	wire [2:0] w_asqrt58_2;
	wire [2:0] w_asqrt58_3;
	wire [2:0] w_asqrt58_4;
	wire [2:0] w_asqrt58_5;
	wire [2:0] w_asqrt58_6;
	wire [2:0] w_asqrt58_7;
	wire [2:0] w_asqrt58_8;
	wire [2:0] w_asqrt58_9;
	wire [2:0] w_asqrt58_10;
	wire [2:0] w_asqrt58_11;
	wire [2:0] w_asqrt58_12;
	wire [2:0] w_asqrt58_13;
	wire [2:0] w_asqrt58_14;
	wire [2:0] w_asqrt58_15;
	wire [2:0] w_asqrt58_16;
	wire [2:0] w_asqrt58_17;
	wire [2:0] w_asqrt58_18;
	wire [2:0] w_asqrt58_19;
	wire [2:0] w_asqrt58_20;
	wire [2:0] w_asqrt58_21;
	wire [2:0] w_asqrt58_22;
	wire [2:0] w_asqrt58_23;
	wire [2:0] w_asqrt58_24;
	wire [2:0] w_asqrt58_25;
	wire [2:0] w_asqrt58_26;
	wire [2:0] w_asqrt58_27;
	wire [2:0] w_asqrt58_28;
	wire [2:0] w_asqrt58_29;
	wire [2:0] w_asqrt58_30;
	wire w_asqrt58_31;
	wire asqrt_fa_58;
	wire [2:0] w_asqrt59_0;
	wire [2:0] w_asqrt59_1;
	wire [2:0] w_asqrt59_2;
	wire [2:0] w_asqrt59_3;
	wire [2:0] w_asqrt59_4;
	wire [2:0] w_asqrt59_5;
	wire [2:0] w_asqrt59_6;
	wire [2:0] w_asqrt59_7;
	wire [2:0] w_asqrt59_8;
	wire [2:0] w_asqrt59_9;
	wire [2:0] w_asqrt59_10;
	wire [2:0] w_asqrt59_11;
	wire [2:0] w_asqrt59_12;
	wire [2:0] w_asqrt59_13;
	wire [2:0] w_asqrt59_14;
	wire [2:0] w_asqrt59_15;
	wire [2:0] w_asqrt59_16;
	wire [2:0] w_asqrt59_17;
	wire [2:0] w_asqrt59_18;
	wire [2:0] w_asqrt59_19;
	wire [2:0] w_asqrt59_20;
	wire [2:0] w_asqrt59_21;
	wire [2:0] w_asqrt59_22;
	wire [2:0] w_asqrt59_23;
	wire [2:0] w_asqrt59_24;
	wire [2:0] w_asqrt59_25;
	wire [2:0] w_asqrt59_26;
	wire [2:0] w_asqrt59_27;
	wire [2:0] w_asqrt59_28;
	wire [2:0] w_asqrt59_29;
	wire [1:0] w_asqrt59_30;
	wire asqrt_fa_59;
	wire [2:0] w_asqrt60_0;
	wire [2:0] w_asqrt60_1;
	wire [2:0] w_asqrt60_2;
	wire [2:0] w_asqrt60_3;
	wire [2:0] w_asqrt60_4;
	wire [2:0] w_asqrt60_5;
	wire [2:0] w_asqrt60_6;
	wire [2:0] w_asqrt60_7;
	wire [2:0] w_asqrt60_8;
	wire [2:0] w_asqrt60_9;
	wire [2:0] w_asqrt60_10;
	wire [2:0] w_asqrt60_11;
	wire [2:0] w_asqrt60_12;
	wire [2:0] w_asqrt60_13;
	wire [2:0] w_asqrt60_14;
	wire [2:0] w_asqrt60_15;
	wire [2:0] w_asqrt60_16;
	wire [2:0] w_asqrt60_17;
	wire [2:0] w_asqrt60_18;
	wire [2:0] w_asqrt60_19;
	wire [2:0] w_asqrt60_20;
	wire [2:0] w_asqrt60_21;
	wire [2:0] w_asqrt60_22;
	wire [2:0] w_asqrt60_23;
	wire [2:0] w_asqrt60_24;
	wire [2:0] w_asqrt60_25;
	wire [2:0] w_asqrt60_26;
	wire [2:0] w_asqrt60_27;
	wire [2:0] w_asqrt60_28;
	wire [2:0] w_asqrt60_29;
	wire [1:0] w_asqrt60_30;
	wire asqrt_fa_60;
	wire [2:0] w_asqrt61_0;
	wire [2:0] w_asqrt61_1;
	wire [2:0] w_asqrt61_2;
	wire [2:0] w_asqrt61_3;
	wire [2:0] w_asqrt61_4;
	wire [2:0] w_asqrt61_5;
	wire [2:0] w_asqrt61_6;
	wire [2:0] w_asqrt61_7;
	wire [2:0] w_asqrt61_8;
	wire [2:0] w_asqrt61_9;
	wire [2:0] w_asqrt61_10;
	wire [2:0] w_asqrt61_11;
	wire [2:0] w_asqrt61_12;
	wire [2:0] w_asqrt61_13;
	wire [2:0] w_asqrt61_14;
	wire [2:0] w_asqrt61_15;
	wire [2:0] w_asqrt61_16;
	wire [2:0] w_asqrt61_17;
	wire [2:0] w_asqrt61_18;
	wire [2:0] w_asqrt61_19;
	wire [2:0] w_asqrt61_20;
	wire [2:0] w_asqrt61_21;
	wire [2:0] w_asqrt61_22;
	wire [2:0] w_asqrt61_23;
	wire [2:0] w_asqrt61_24;
	wire [2:0] w_asqrt61_25;
	wire [2:0] w_asqrt61_26;
	wire [2:0] w_asqrt61_27;
	wire [2:0] w_asqrt61_28;
	wire [2:0] w_asqrt61_29;
	wire [2:0] w_asqrt61_30;
	wire w_asqrt61_31;
	wire asqrt_fa_61;
	wire [2:0] w_asqrt62_0;
	wire [2:0] w_asqrt62_1;
	wire [2:0] w_asqrt62_2;
	wire [2:0] w_asqrt62_3;
	wire [2:0] w_asqrt62_4;
	wire [2:0] w_asqrt62_5;
	wire [2:0] w_asqrt62_6;
	wire [2:0] w_asqrt62_7;
	wire [2:0] w_asqrt62_8;
	wire [2:0] w_asqrt62_9;
	wire [2:0] w_asqrt62_10;
	wire [2:0] w_asqrt62_11;
	wire [2:0] w_asqrt62_12;
	wire [2:0] w_asqrt62_13;
	wire [2:0] w_asqrt62_14;
	wire [2:0] w_asqrt62_15;
	wire [2:0] w_asqrt62_16;
	wire [2:0] w_asqrt62_17;
	wire [2:0] w_asqrt62_18;
	wire [2:0] w_asqrt62_19;
	wire [2:0] w_asqrt62_20;
	wire [2:0] w_asqrt62_21;
	wire [2:0] w_asqrt62_22;
	wire [2:0] w_asqrt62_23;
	wire [2:0] w_asqrt62_24;
	wire [2:0] w_asqrt62_25;
	wire [2:0] w_asqrt62_26;
	wire [2:0] w_asqrt62_27;
	wire [2:0] w_asqrt62_28;
	wire [2:0] w_asqrt62_29;
	wire [2:0] w_asqrt62_30;
	wire w_asqrt62_31;
	wire asqrt_fa_62;
	wire [2:0] w_asqrt63_0;
	wire [2:0] w_asqrt63_1;
	wire [2:0] w_asqrt63_2;
	wire [2:0] w_asqrt63_3;
	wire [2:0] w_asqrt63_4;
	wire [2:0] w_asqrt63_5;
	wire [2:0] w_asqrt63_6;
	wire [2:0] w_asqrt63_7;
	wire [2:0] w_asqrt63_8;
	wire [2:0] w_asqrt63_9;
	wire [2:0] w_asqrt63_10;
	wire [2:0] w_asqrt63_11;
	wire [2:0] w_asqrt63_12;
	wire [2:0] w_asqrt63_13;
	wire [2:0] w_asqrt63_14;
	wire [2:0] w_asqrt63_15;
	wire [2:0] w_asqrt63_16;
	wire w_asqrt63_17;
	wire asqrt_fa_63;
	wire [1:0] w_n192_0;
	wire [1:0] w_n193_0;
	wire [2:0] w_n194_0;
	wire [2:0] w_n194_1;
	wire [2:0] w_n194_2;
	wire [2:0] w_n194_3;
	wire [2:0] w_n194_4;
	wire [2:0] w_n194_5;
	wire [2:0] w_n194_6;
	wire [2:0] w_n194_7;
	wire [2:0] w_n194_8;
	wire [2:0] w_n194_9;
	wire [2:0] w_n194_10;
	wire [2:0] w_n194_11;
	wire [2:0] w_n194_12;
	wire [2:0] w_n194_13;
	wire [2:0] w_n194_14;
	wire [2:0] w_n194_15;
	wire [2:0] w_n194_16;
	wire [2:0] w_n194_17;
	wire [2:0] w_n194_18;
	wire [2:0] w_n194_19;
	wire [2:0] w_n194_20;
	wire [2:0] w_n194_21;
	wire [2:0] w_n194_22;
	wire [2:0] w_n194_23;
	wire [2:0] w_n194_24;
	wire [2:0] w_n194_25;
	wire [2:0] w_n194_26;
	wire [2:0] w_n194_27;
	wire [2:0] w_n194_28;
	wire [2:0] w_n194_29;
	wire [2:0] w_n194_30;
	wire [2:0] w_n194_31;
	wire [2:0] w_n194_32;
	wire [2:0] w_n194_33;
	wire [2:0] w_n194_34;
	wire [2:0] w_n194_35;
	wire [2:0] w_n194_36;
	wire [2:0] w_n194_37;
	wire [2:0] w_n194_38;
	wire [2:0] w_n194_39;
	wire [2:0] w_n194_40;
	wire [2:0] w_n194_41;
	wire [2:0] w_n194_42;
	wire [2:0] w_n194_43;
	wire [1:0] w_n195_0;
	wire [1:0] w_n196_0;
	wire [1:0] w_n197_0;
	wire [2:0] w_n199_0;
	wire [2:0] w_n199_1;
	wire [2:0] w_n199_2;
	wire [2:0] w_n199_3;
	wire [2:0] w_n199_4;
	wire [2:0] w_n199_5;
	wire [2:0] w_n199_6;
	wire [2:0] w_n199_7;
	wire [2:0] w_n199_8;
	wire [2:0] w_n199_9;
	wire [2:0] w_n199_10;
	wire [2:0] w_n199_11;
	wire [2:0] w_n199_12;
	wire [2:0] w_n199_13;
	wire [2:0] w_n199_14;
	wire [2:0] w_n199_15;
	wire [2:0] w_n199_16;
	wire [2:0] w_n199_17;
	wire [2:0] w_n199_18;
	wire [2:0] w_n199_19;
	wire [2:0] w_n199_20;
	wire [2:0] w_n199_21;
	wire [2:0] w_n199_22;
	wire [2:0] w_n199_23;
	wire [2:0] w_n199_24;
	wire [2:0] w_n199_25;
	wire [2:0] w_n199_26;
	wire [2:0] w_n199_27;
	wire [2:0] w_n199_28;
	wire [2:0] w_n199_29;
	wire [2:0] w_n199_30;
	wire [2:0] w_n199_31;
	wire [2:0] w_n199_32;
	wire [2:0] w_n199_33;
	wire [2:0] w_n199_34;
	wire [2:0] w_n199_35;
	wire [2:0] w_n199_36;
	wire [2:0] w_n199_37;
	wire [2:0] w_n199_38;
	wire [2:0] w_n199_39;
	wire [2:0] w_n199_40;
	wire [2:0] w_n199_41;
	wire [2:0] w_n199_42;
	wire [2:0] w_n199_43;
	wire [2:0] w_n199_44;
	wire [2:0] w_n199_45;
	wire [1:0] w_n200_0;
	wire [2:0] w_n203_0;
	wire [1:0] w_n206_0;
	wire [2:0] w_n209_0;
	wire [2:0] w_n211_0;
	wire [1:0] w_n211_1;
	wire [1:0] w_n212_0;
	wire [2:0] w_n215_0;
	wire [2:0] w_n216_0;
	wire [1:0] w_n218_0;
	wire [1:0] w_n221_0;
	wire [2:0] w_n223_0;
	wire [2:0] w_n223_1;
	wire [2:0] w_n223_2;
	wire [2:0] w_n223_3;
	wire [2:0] w_n223_4;
	wire [2:0] w_n223_5;
	wire [2:0] w_n223_6;
	wire [2:0] w_n223_7;
	wire [2:0] w_n223_8;
	wire [2:0] w_n223_9;
	wire [2:0] w_n223_10;
	wire [2:0] w_n223_11;
	wire [2:0] w_n223_12;
	wire [2:0] w_n223_13;
	wire [2:0] w_n223_14;
	wire [2:0] w_n223_15;
	wire [2:0] w_n223_16;
	wire [2:0] w_n223_17;
	wire [2:0] w_n223_18;
	wire [2:0] w_n223_19;
	wire [2:0] w_n223_20;
	wire [2:0] w_n223_21;
	wire [2:0] w_n223_22;
	wire [2:0] w_n223_23;
	wire [2:0] w_n223_24;
	wire [2:0] w_n223_25;
	wire [2:0] w_n223_26;
	wire [2:0] w_n223_27;
	wire [2:0] w_n223_28;
	wire [2:0] w_n223_29;
	wire [2:0] w_n223_30;
	wire [2:0] w_n223_31;
	wire [2:0] w_n223_32;
	wire [2:0] w_n223_33;
	wire [2:0] w_n223_34;
	wire [2:0] w_n223_35;
	wire [2:0] w_n223_36;
	wire [2:0] w_n223_37;
	wire [2:0] w_n223_38;
	wire [2:0] w_n223_39;
	wire [1:0] w_n226_0;
	wire [2:0] w_n229_0;
	wire [2:0] w_n231_0;
	wire [1:0] w_n231_1;
	wire [2:0] w_n232_0;
	wire [2:0] w_n236_0;
	wire [1:0] w_n239_0;
	wire [1:0] w_n241_0;
	wire [2:0] w_n242_0;
	wire [1:0] w_n248_0;
	wire [1:0] w_n249_0;
	wire [1:0] w_n254_0;
	wire [2:0] w_n261_0;
	wire [1:0] w_n261_1;
	wire [1:0] w_n262_0;
	wire [2:0] w_n265_0;
	wire [1:0] w_n266_0;
	wire [1:0] w_n267_0;
	wire [1:0] w_n268_0;
	wire [1:0] w_n270_0;
	wire [1:0] w_n272_0;
	wire [1:0] w_n274_0;
	wire [2:0] w_n277_0;
	wire [1:0] w_n283_0;
	wire [2:0] w_n285_0;
	wire [1:0] w_n285_1;
	wire [2:0] w_n289_0;
	wire [1:0] w_n289_1;
	wire [2:0] w_n290_0;
	wire [2:0] w_n290_1;
	wire [2:0] w_n290_2;
	wire [2:0] w_n290_3;
	wire [2:0] w_n290_4;
	wire [2:0] w_n290_5;
	wire [2:0] w_n290_6;
	wire [2:0] w_n290_7;
	wire [2:0] w_n290_8;
	wire [2:0] w_n290_9;
	wire [2:0] w_n290_10;
	wire [2:0] w_n290_11;
	wire [2:0] w_n290_12;
	wire [2:0] w_n290_13;
	wire [2:0] w_n290_14;
	wire [2:0] w_n290_15;
	wire [2:0] w_n290_16;
	wire [2:0] w_n290_17;
	wire [2:0] w_n290_18;
	wire [2:0] w_n290_19;
	wire [2:0] w_n290_20;
	wire [2:0] w_n290_21;
	wire [2:0] w_n290_22;
	wire [2:0] w_n290_23;
	wire [2:0] w_n290_24;
	wire [2:0] w_n290_25;
	wire [2:0] w_n290_26;
	wire [2:0] w_n290_27;
	wire [2:0] w_n290_28;
	wire [2:0] w_n290_29;
	wire [2:0] w_n290_30;
	wire [2:0] w_n290_31;
	wire [2:0] w_n290_32;
	wire [2:0] w_n290_33;
	wire [2:0] w_n290_34;
	wire [2:0] w_n290_35;
	wire [2:0] w_n290_36;
	wire [2:0] w_n290_37;
	wire [2:0] w_n290_38;
	wire [1:0] w_n290_39;
	wire [1:0] w_n295_0;
	wire [2:0] w_n296_0;
	wire [1:0] w_n301_0;
	wire [2:0] w_n305_0;
	wire [2:0] w_n305_1;
	wire [2:0] w_n305_2;
	wire [2:0] w_n305_3;
	wire [2:0] w_n305_4;
	wire [2:0] w_n305_5;
	wire [2:0] w_n305_6;
	wire [2:0] w_n305_7;
	wire [2:0] w_n305_8;
	wire [2:0] w_n305_9;
	wire [2:0] w_n305_10;
	wire [2:0] w_n305_11;
	wire [2:0] w_n305_12;
	wire [2:0] w_n305_13;
	wire [2:0] w_n305_14;
	wire [2:0] w_n305_15;
	wire [2:0] w_n305_16;
	wire [2:0] w_n305_17;
	wire [2:0] w_n305_18;
	wire [2:0] w_n305_19;
	wire [2:0] w_n305_20;
	wire [2:0] w_n305_21;
	wire [2:0] w_n305_22;
	wire [2:0] w_n305_23;
	wire [2:0] w_n305_24;
	wire [2:0] w_n305_25;
	wire [2:0] w_n305_26;
	wire [2:0] w_n305_27;
	wire [2:0] w_n305_28;
	wire [2:0] w_n305_29;
	wire [2:0] w_n305_30;
	wire [2:0] w_n305_31;
	wire [2:0] w_n305_32;
	wire [2:0] w_n305_33;
	wire [2:0] w_n305_34;
	wire [2:0] w_n305_35;
	wire [2:0] w_n305_36;
	wire [2:0] w_n305_37;
	wire [2:0] w_n305_38;
	wire [2:0] w_n305_39;
	wire [2:0] w_n308_0;
	wire [1:0] w_n308_1;
	wire [2:0] w_n309_0;
	wire [2:0] w_n313_0;
	wire [1:0] w_n314_0;
	wire [1:0] w_n315_0;
	wire [1:0] w_n316_0;
	wire [1:0] w_n318_0;
	wire [1:0] w_n320_0;
	wire [1:0] w_n322_0;
	wire [1:0] w_n325_0;
	wire [1:0] w_n329_0;
	wire [2:0] w_n331_0;
	wire [1:0] w_n336_0;
	wire [2:0] w_n338_0;
	wire [2:0] w_n342_0;
	wire [1:0] w_n348_0;
	wire [2:0] w_n349_0;
	wire [1:0] w_n358_0;
	wire [2:0] w_n363_0;
	wire [1:0] w_n363_1;
	wire [1:0] w_n364_0;
	wire [2:0] w_n367_0;
	wire [1:0] w_n368_0;
	wire [1:0] w_n369_0;
	wire [1:0] w_n370_0;
	wire [1:0] w_n372_0;
	wire [1:0] w_n374_0;
	wire [1:0] w_n376_0;
	wire [1:0] w_n385_0;
	wire [2:0] w_n387_0;
	wire [1:0] w_n388_0;
	wire [1:0] w_n392_0;
	wire [1:0] w_n394_0;
	wire [1:0] w_n396_0;
	wire [1:0] w_n401_0;
	wire [1:0] w_n403_0;
	wire [1:0] w_n404_0;
	wire [2:0] w_n405_0;
	wire [2:0] w_n405_1;
	wire [1:0] w_n408_0;
	wire [2:0] w_n409_0;
	wire [1:0] w_n410_0;
	wire [1:0] w_n411_0;
	wire [1:0] w_n417_0;
	wire [2:0] w_n418_0;
	wire [1:0] w_n419_0;
	wire [1:0] w_n424_0;
	wire [2:0] w_n425_0;
	wire [2:0] w_n425_1;
	wire [2:0] w_n425_2;
	wire [2:0] w_n425_3;
	wire [2:0] w_n425_4;
	wire [2:0] w_n425_5;
	wire [2:0] w_n425_6;
	wire [2:0] w_n425_7;
	wire [2:0] w_n425_8;
	wire [2:0] w_n425_9;
	wire [2:0] w_n425_10;
	wire [2:0] w_n425_11;
	wire [2:0] w_n425_12;
	wire [2:0] w_n425_13;
	wire [2:0] w_n425_14;
	wire [2:0] w_n425_15;
	wire [2:0] w_n425_16;
	wire [2:0] w_n425_17;
	wire [2:0] w_n425_18;
	wire [2:0] w_n425_19;
	wire [2:0] w_n425_20;
	wire [2:0] w_n425_21;
	wire [2:0] w_n425_22;
	wire [2:0] w_n425_23;
	wire [2:0] w_n425_24;
	wire [2:0] w_n425_25;
	wire [2:0] w_n425_26;
	wire [2:0] w_n425_27;
	wire [2:0] w_n425_28;
	wire [2:0] w_n425_29;
	wire [2:0] w_n425_30;
	wire [2:0] w_n425_31;
	wire [2:0] w_n425_32;
	wire [2:0] w_n425_33;
	wire [2:0] w_n425_34;
	wire [2:0] w_n425_35;
	wire [2:0] w_n425_36;
	wire [2:0] w_n430_0;
	wire [2:0] w_n430_1;
	wire [2:0] w_n430_2;
	wire [2:0] w_n430_3;
	wire [2:0] w_n430_4;
	wire [2:0] w_n430_5;
	wire [2:0] w_n430_6;
	wire [2:0] w_n430_7;
	wire [2:0] w_n430_8;
	wire [2:0] w_n430_9;
	wire [2:0] w_n430_10;
	wire [2:0] w_n430_11;
	wire [2:0] w_n430_12;
	wire [2:0] w_n430_13;
	wire [2:0] w_n430_14;
	wire [2:0] w_n430_15;
	wire [2:0] w_n430_16;
	wire [2:0] w_n430_17;
	wire [2:0] w_n430_18;
	wire [2:0] w_n430_19;
	wire [2:0] w_n430_20;
	wire [2:0] w_n430_21;
	wire [2:0] w_n430_22;
	wire [2:0] w_n430_23;
	wire [2:0] w_n430_24;
	wire [2:0] w_n430_25;
	wire [2:0] w_n430_26;
	wire [2:0] w_n430_27;
	wire [2:0] w_n430_28;
	wire [2:0] w_n430_29;
	wire [2:0] w_n430_30;
	wire [2:0] w_n430_31;
	wire [2:0] w_n430_32;
	wire [2:0] w_n430_33;
	wire [2:0] w_n430_34;
	wire [2:0] w_n430_35;
	wire [2:0] w_n430_36;
	wire [2:0] w_n430_37;
	wire [2:0] w_n430_38;
	wire [2:0] w_n433_0;
	wire [1:0] w_n433_1;
	wire [2:0] w_n434_0;
	wire [2:0] w_n438_0;
	wire [1:0] w_n439_0;
	wire [1:0] w_n440_0;
	wire [1:0] w_n441_0;
	wire [1:0] w_n443_0;
	wire [1:0] w_n445_0;
	wire [1:0] w_n447_0;
	wire [1:0] w_n450_0;
	wire [1:0] w_n455_0;
	wire [2:0] w_n457_0;
	wire [1:0] w_n458_0;
	wire [1:0] w_n462_0;
	wire [1:0] w_n463_0;
	wire [1:0] w_n465_0;
	wire [1:0] w_n469_0;
	wire [1:0] w_n471_0;
	wire [1:0] w_n472_0;
	wire [2:0] w_n473_0;
	wire [1:0] w_n478_0;
	wire [2:0] w_n481_0;
	wire [1:0] w_n483_0;
	wire [2:0] w_n488_0;
	wire [1:0] w_n489_0;
	wire [1:0] w_n490_0;
	wire [1:0] w_n495_0;
	wire [2:0] w_n496_0;
	wire [1:0] w_n501_0;
	wire [2:0] w_n507_0;
	wire [1:0] w_n507_1;
	wire [1:0] w_n508_0;
	wire [2:0] w_n511_0;
	wire [1:0] w_n512_0;
	wire [1:0] w_n513_0;
	wire [1:0] w_n514_0;
	wire [1:0] w_n516_0;
	wire [1:0] w_n518_0;
	wire [1:0] w_n520_0;
	wire [1:0] w_n529_0;
	wire [2:0] w_n531_0;
	wire [1:0] w_n532_0;
	wire [1:0] w_n536_0;
	wire [1:0] w_n538_0;
	wire [1:0] w_n540_0;
	wire [1:0] w_n545_0;
	wire [1:0] w_n547_0;
	wire [1:0] w_n548_0;
	wire [2:0] w_n549_0;
	wire [1:0] w_n550_0;
	wire [1:0] w_n555_0;
	wire [1:0] w_n556_0;
	wire [1:0] w_n558_0;
	wire [1:0] w_n560_0;
	wire [1:0] w_n563_0;
	wire [1:0] w_n569_0;
	wire [2:0] w_n571_0;
	wire [2:0] w_n571_1;
	wire [2:0] w_n574_0;
	wire [1:0] w_n574_1;
	wire [2:0] w_n576_0;
	wire [1:0] w_n577_0;
	wire [1:0] w_n583_0;
	wire [1:0] w_n584_0;
	wire [1:0] w_n589_0;
	wire [2:0] w_n590_0;
	wire [2:0] w_n590_1;
	wire [2:0] w_n590_2;
	wire [2:0] w_n590_3;
	wire [2:0] w_n590_4;
	wire [2:0] w_n590_5;
	wire [2:0] w_n590_6;
	wire [2:0] w_n590_7;
	wire [2:0] w_n590_8;
	wire [2:0] w_n590_9;
	wire [2:0] w_n590_10;
	wire [2:0] w_n590_11;
	wire [2:0] w_n590_12;
	wire [2:0] w_n590_13;
	wire [2:0] w_n590_14;
	wire [2:0] w_n590_15;
	wire [2:0] w_n590_16;
	wire [2:0] w_n590_17;
	wire [2:0] w_n590_18;
	wire [2:0] w_n590_19;
	wire [2:0] w_n590_20;
	wire [2:0] w_n590_21;
	wire [2:0] w_n590_22;
	wire [2:0] w_n590_23;
	wire [2:0] w_n590_24;
	wire [2:0] w_n590_25;
	wire [2:0] w_n590_26;
	wire [2:0] w_n590_27;
	wire [2:0] w_n590_28;
	wire [2:0] w_n590_29;
	wire [2:0] w_n590_30;
	wire [2:0] w_n590_31;
	wire [2:0] w_n590_32;
	wire [2:0] w_n590_33;
	wire [2:0] w_n590_34;
	wire [2:0] w_n590_35;
	wire [2:0] w_n595_0;
	wire [2:0] w_n595_1;
	wire [2:0] w_n595_2;
	wire [2:0] w_n595_3;
	wire [2:0] w_n595_4;
	wire [2:0] w_n595_5;
	wire [2:0] w_n595_6;
	wire [2:0] w_n595_7;
	wire [2:0] w_n595_8;
	wire [2:0] w_n595_9;
	wire [2:0] w_n595_10;
	wire [2:0] w_n595_11;
	wire [2:0] w_n595_12;
	wire [2:0] w_n595_13;
	wire [2:0] w_n595_14;
	wire [2:0] w_n595_15;
	wire [2:0] w_n595_16;
	wire [2:0] w_n595_17;
	wire [2:0] w_n595_18;
	wire [2:0] w_n595_19;
	wire [2:0] w_n595_20;
	wire [2:0] w_n595_21;
	wire [2:0] w_n595_22;
	wire [2:0] w_n595_23;
	wire [2:0] w_n595_24;
	wire [2:0] w_n595_25;
	wire [2:0] w_n595_26;
	wire [2:0] w_n595_27;
	wire [2:0] w_n595_28;
	wire [2:0] w_n595_29;
	wire [2:0] w_n595_30;
	wire [2:0] w_n595_31;
	wire [2:0] w_n595_32;
	wire [2:0] w_n595_33;
	wire [2:0] w_n595_34;
	wire [2:0] w_n595_35;
	wire [2:0] w_n595_36;
	wire [2:0] w_n595_37;
	wire [2:0] w_n595_38;
	wire [2:0] w_n598_0;
	wire [1:0] w_n598_1;
	wire [2:0] w_n599_0;
	wire [2:0] w_n603_0;
	wire [1:0] w_n604_0;
	wire [1:0] w_n605_0;
	wire [1:0] w_n606_0;
	wire [1:0] w_n608_0;
	wire [1:0] w_n610_0;
	wire [1:0] w_n612_0;
	wire [1:0] w_n615_0;
	wire [1:0] w_n620_0;
	wire [2:0] w_n622_0;
	wire [1:0] w_n623_0;
	wire [1:0] w_n627_0;
	wire [1:0] w_n628_0;
	wire [1:0] w_n630_0;
	wire [1:0] w_n634_0;
	wire [1:0] w_n636_0;
	wire [1:0] w_n637_0;
	wire [2:0] w_n638_0;
	wire [1:0] w_n639_0;
	wire [1:0] w_n643_0;
	wire [1:0] w_n645_0;
	wire [1:0] w_n647_0;
	wire [1:0] w_n649_0;
	wire [1:0] w_n651_0;
	wire [1:0] w_n657_0;
	wire [2:0] w_n659_0;
	wire [1:0] w_n665_0;
	wire [2:0] w_n668_0;
	wire [2:0] w_n672_0;
	wire [1:0] w_n673_0;
	wire [1:0] w_n678_0;
	wire [2:0] w_n679_0;
	wire [1:0] w_n684_0;
	wire [2:0] w_n690_0;
	wire [1:0] w_n690_1;
	wire [1:0] w_n691_0;
	wire [2:0] w_n694_0;
	wire [1:0] w_n695_0;
	wire [1:0] w_n696_0;
	wire [1:0] w_n697_0;
	wire [1:0] w_n699_0;
	wire [1:0] w_n701_0;
	wire [1:0] w_n703_0;
	wire [1:0] w_n712_0;
	wire [2:0] w_n714_0;
	wire [1:0] w_n715_0;
	wire [1:0] w_n719_0;
	wire [1:0] w_n721_0;
	wire [1:0] w_n723_0;
	wire [1:0] w_n728_0;
	wire [1:0] w_n730_0;
	wire [1:0] w_n731_0;
	wire [2:0] w_n732_0;
	wire [1:0] w_n733_0;
	wire [1:0] w_n738_0;
	wire [1:0] w_n739_0;
	wire [1:0] w_n741_0;
	wire [1:0] w_n743_0;
	wire [1:0] w_n746_0;
	wire [1:0] w_n752_0;
	wire [2:0] w_n754_0;
	wire [1:0] w_n755_0;
	wire [1:0] w_n759_0;
	wire [1:0] w_n760_0;
	wire [1:0] w_n762_0;
	wire [1:0] w_n767_0;
	wire [1:0] w_n769_0;
	wire [1:0] w_n770_0;
	wire [2:0] w_n771_0;
	wire [2:0] w_n771_1;
	wire [2:0] w_n774_0;
	wire [1:0] w_n774_1;
	wire [2:0] w_n776_0;
	wire [1:0] w_n777_0;
	wire [1:0] w_n778_0;
	wire [1:0] w_n784_0;
	wire [1:0] w_n785_0;
	wire [1:0] w_n790_0;
	wire [2:0] w_n791_0;
	wire [2:0] w_n791_1;
	wire [2:0] w_n791_2;
	wire [2:0] w_n791_3;
	wire [2:0] w_n791_4;
	wire [2:0] w_n791_5;
	wire [2:0] w_n791_6;
	wire [2:0] w_n791_7;
	wire [2:0] w_n791_8;
	wire [2:0] w_n791_9;
	wire [2:0] w_n791_10;
	wire [2:0] w_n791_11;
	wire [2:0] w_n791_12;
	wire [2:0] w_n791_13;
	wire [2:0] w_n791_14;
	wire [2:0] w_n791_15;
	wire [2:0] w_n791_16;
	wire [2:0] w_n791_17;
	wire [2:0] w_n791_18;
	wire [2:0] w_n791_19;
	wire [2:0] w_n791_20;
	wire [2:0] w_n791_21;
	wire [2:0] w_n791_22;
	wire [2:0] w_n791_23;
	wire [2:0] w_n791_24;
	wire [2:0] w_n791_25;
	wire [2:0] w_n791_26;
	wire [2:0] w_n791_27;
	wire [2:0] w_n791_28;
	wire [2:0] w_n791_29;
	wire [2:0] w_n791_30;
	wire [2:0] w_n791_31;
	wire [2:0] w_n791_32;
	wire [2:0] w_n791_33;
	wire [1:0] w_n791_34;
	wire [2:0] w_n796_0;
	wire [2:0] w_n796_1;
	wire [2:0] w_n796_2;
	wire [2:0] w_n796_3;
	wire [2:0] w_n796_4;
	wire [2:0] w_n796_5;
	wire [2:0] w_n796_6;
	wire [2:0] w_n796_7;
	wire [2:0] w_n796_8;
	wire [2:0] w_n796_9;
	wire [2:0] w_n796_10;
	wire [2:0] w_n796_11;
	wire [2:0] w_n796_12;
	wire [2:0] w_n796_13;
	wire [2:0] w_n796_14;
	wire [2:0] w_n796_15;
	wire [2:0] w_n796_16;
	wire [2:0] w_n796_17;
	wire [2:0] w_n796_18;
	wire [2:0] w_n796_19;
	wire [2:0] w_n796_20;
	wire [2:0] w_n796_21;
	wire [2:0] w_n796_22;
	wire [2:0] w_n796_23;
	wire [2:0] w_n796_24;
	wire [2:0] w_n796_25;
	wire [2:0] w_n796_26;
	wire [2:0] w_n796_27;
	wire [2:0] w_n796_28;
	wire [2:0] w_n796_29;
	wire [2:0] w_n796_30;
	wire [2:0] w_n796_31;
	wire [2:0] w_n796_32;
	wire [2:0] w_n796_33;
	wire [2:0] w_n796_34;
	wire [2:0] w_n796_35;
	wire [2:0] w_n796_36;
	wire [2:0] w_n796_37;
	wire [2:0] w_n799_0;
	wire [1:0] w_n799_1;
	wire [2:0] w_n800_0;
	wire [2:0] w_n804_0;
	wire [1:0] w_n805_0;
	wire [1:0] w_n806_0;
	wire [1:0] w_n807_0;
	wire [1:0] w_n809_0;
	wire [1:0] w_n811_0;
	wire [1:0] w_n813_0;
	wire [1:0] w_n816_0;
	wire [1:0] w_n821_0;
	wire [2:0] w_n823_0;
	wire [1:0] w_n824_0;
	wire [1:0] w_n828_0;
	wire [1:0] w_n829_0;
	wire [1:0] w_n831_0;
	wire [1:0] w_n835_0;
	wire [1:0] w_n837_0;
	wire [1:0] w_n838_0;
	wire [2:0] w_n839_0;
	wire [1:0] w_n840_0;
	wire [1:0] w_n844_0;
	wire [1:0] w_n846_0;
	wire [1:0] w_n848_0;
	wire [1:0] w_n850_0;
	wire [1:0] w_n852_0;
	wire [1:0] w_n858_0;
	wire [2:0] w_n860_0;
	wire [1:0] w_n861_0;
	wire [1:0] w_n866_0;
	wire [1:0] w_n868_0;
	wire [1:0] w_n870_0;
	wire [1:0] w_n874_0;
	wire [1:0] w_n876_0;
	wire [1:0] w_n877_0;
	wire [2:0] w_n878_0;
	wire [1:0] w_n885_0;
	wire [2:0] w_n887_0;
	wire [1:0] w_n889_0;
	wire [2:0] w_n894_0;
	wire [1:0] w_n895_0;
	wire [1:0] w_n896_0;
	wire [1:0] w_n901_0;
	wire [2:0] w_n902_0;
	wire [1:0] w_n907_0;
	wire [2:0] w_n913_0;
	wire [1:0] w_n913_1;
	wire [1:0] w_n914_0;
	wire [2:0] w_n917_0;
	wire [1:0] w_n918_0;
	wire [1:0] w_n919_0;
	wire [1:0] w_n920_0;
	wire [1:0] w_n922_0;
	wire [1:0] w_n924_0;
	wire [1:0] w_n926_0;
	wire [1:0] w_n935_0;
	wire [2:0] w_n937_0;
	wire [1:0] w_n938_0;
	wire [1:0] w_n942_0;
	wire [1:0] w_n944_0;
	wire [1:0] w_n946_0;
	wire [1:0] w_n951_0;
	wire [1:0] w_n953_0;
	wire [1:0] w_n954_0;
	wire [2:0] w_n955_0;
	wire [1:0] w_n956_0;
	wire [1:0] w_n961_0;
	wire [1:0] w_n962_0;
	wire [1:0] w_n964_0;
	wire [1:0] w_n966_0;
	wire [1:0] w_n969_0;
	wire [1:0] w_n975_0;
	wire [2:0] w_n977_0;
	wire [1:0] w_n978_0;
	wire [1:0] w_n982_0;
	wire [1:0] w_n983_0;
	wire [1:0] w_n985_0;
	wire [1:0] w_n990_0;
	wire [1:0] w_n992_0;
	wire [1:0] w_n993_0;
	wire [2:0] w_n994_0;
	wire [1:0] w_n995_0;
	wire [1:0] w_n999_0;
	wire [1:0] w_n1000_0;
	wire [1:0] w_n1002_0;
	wire [1:0] w_n1004_0;
	wire [1:0] w_n1007_0;
	wire [1:0] w_n1013_0;
	wire [2:0] w_n1015_0;
	wire [2:0] w_n1015_1;
	wire [1:0] w_n1018_0;
	wire [2:0] w_n1019_0;
	wire [1:0] w_n1020_0;
	wire [1:0] w_n1026_0;
	wire [2:0] w_n1027_0;
	wire [1:0] w_n1028_0;
	wire [1:0] w_n1033_0;
	wire [2:0] w_n1034_0;
	wire [2:0] w_n1034_1;
	wire [2:0] w_n1034_2;
	wire [2:0] w_n1034_3;
	wire [2:0] w_n1034_4;
	wire [2:0] w_n1034_5;
	wire [2:0] w_n1034_6;
	wire [2:0] w_n1034_7;
	wire [2:0] w_n1034_8;
	wire [2:0] w_n1034_9;
	wire [2:0] w_n1034_10;
	wire [2:0] w_n1034_11;
	wire [2:0] w_n1034_12;
	wire [2:0] w_n1034_13;
	wire [2:0] w_n1034_14;
	wire [2:0] w_n1034_15;
	wire [2:0] w_n1034_16;
	wire [2:0] w_n1034_17;
	wire [2:0] w_n1034_18;
	wire [2:0] w_n1034_19;
	wire [2:0] w_n1034_20;
	wire [2:0] w_n1034_21;
	wire [2:0] w_n1034_22;
	wire [2:0] w_n1034_23;
	wire [2:0] w_n1034_24;
	wire [2:0] w_n1034_25;
	wire [2:0] w_n1034_26;
	wire [2:0] w_n1034_27;
	wire [2:0] w_n1034_28;
	wire [2:0] w_n1034_29;
	wire [2:0] w_n1034_30;
	wire [2:0] w_n1034_31;
	wire [2:0] w_n1034_32;
	wire [1:0] w_n1034_33;
	wire [2:0] w_n1039_0;
	wire [2:0] w_n1039_1;
	wire [2:0] w_n1039_2;
	wire [2:0] w_n1039_3;
	wire [2:0] w_n1039_4;
	wire [2:0] w_n1039_5;
	wire [2:0] w_n1039_6;
	wire [2:0] w_n1039_7;
	wire [2:0] w_n1039_8;
	wire [2:0] w_n1039_9;
	wire [2:0] w_n1039_10;
	wire [2:0] w_n1039_11;
	wire [2:0] w_n1039_12;
	wire [2:0] w_n1039_13;
	wire [2:0] w_n1039_14;
	wire [2:0] w_n1039_15;
	wire [2:0] w_n1039_16;
	wire [2:0] w_n1039_17;
	wire [2:0] w_n1039_18;
	wire [2:0] w_n1039_19;
	wire [2:0] w_n1039_20;
	wire [2:0] w_n1039_21;
	wire [2:0] w_n1039_22;
	wire [2:0] w_n1039_23;
	wire [2:0] w_n1039_24;
	wire [2:0] w_n1039_25;
	wire [2:0] w_n1039_26;
	wire [2:0] w_n1039_27;
	wire [2:0] w_n1039_28;
	wire [2:0] w_n1039_29;
	wire [2:0] w_n1039_30;
	wire [2:0] w_n1039_31;
	wire [2:0] w_n1039_32;
	wire [2:0] w_n1039_33;
	wire [2:0] w_n1039_34;
	wire [2:0] w_n1039_35;
	wire [2:0] w_n1039_36;
	wire [2:0] w_n1039_37;
	wire [2:0] w_n1042_0;
	wire [1:0] w_n1042_1;
	wire [2:0] w_n1043_0;
	wire [2:0] w_n1047_0;
	wire [1:0] w_n1048_0;
	wire [1:0] w_n1049_0;
	wire [1:0] w_n1050_0;
	wire [1:0] w_n1052_0;
	wire [1:0] w_n1054_0;
	wire [1:0] w_n1056_0;
	wire [1:0] w_n1059_0;
	wire [1:0] w_n1064_0;
	wire [2:0] w_n1066_0;
	wire [1:0] w_n1067_0;
	wire [1:0] w_n1071_0;
	wire [1:0] w_n1072_0;
	wire [1:0] w_n1074_0;
	wire [1:0] w_n1078_0;
	wire [1:0] w_n1080_0;
	wire [1:0] w_n1081_0;
	wire [2:0] w_n1082_0;
	wire [1:0] w_n1083_0;
	wire [1:0] w_n1087_0;
	wire [1:0] w_n1089_0;
	wire [1:0] w_n1091_0;
	wire [1:0] w_n1093_0;
	wire [1:0] w_n1095_0;
	wire [1:0] w_n1101_0;
	wire [2:0] w_n1103_0;
	wire [1:0] w_n1104_0;
	wire [1:0] w_n1109_0;
	wire [1:0] w_n1111_0;
	wire [1:0] w_n1113_0;
	wire [1:0] w_n1117_0;
	wire [1:0] w_n1119_0;
	wire [1:0] w_n1120_0;
	wire [2:0] w_n1121_0;
	wire [1:0] w_n1122_0;
	wire [1:0] w_n1128_0;
	wire [1:0] w_n1129_0;
	wire [1:0] w_n1131_0;
	wire [1:0] w_n1133_0;
	wire [1:0] w_n1135_0;
	wire [1:0] w_n1141_0;
	wire [2:0] w_n1143_0;
	wire [1:0] w_n1148_0;
	wire [2:0] w_n1150_0;
	wire [2:0] w_n1154_0;
	wire [1:0] w_n1155_0;
	wire [1:0] w_n1160_0;
	wire [2:0] w_n1161_0;
	wire [1:0] w_n1166_0;
	wire [2:0] w_n1172_0;
	wire [1:0] w_n1172_1;
	wire [1:0] w_n1173_0;
	wire [2:0] w_n1176_0;
	wire [1:0] w_n1177_0;
	wire [1:0] w_n1178_0;
	wire [1:0] w_n1179_0;
	wire [1:0] w_n1181_0;
	wire [1:0] w_n1183_0;
	wire [1:0] w_n1185_0;
	wire [1:0] w_n1194_0;
	wire [2:0] w_n1196_0;
	wire [1:0] w_n1197_0;
	wire [1:0] w_n1201_0;
	wire [1:0] w_n1203_0;
	wire [1:0] w_n1205_0;
	wire [1:0] w_n1210_0;
	wire [1:0] w_n1212_0;
	wire [1:0] w_n1213_0;
	wire [2:0] w_n1214_0;
	wire [1:0] w_n1215_0;
	wire [1:0] w_n1220_0;
	wire [1:0] w_n1221_0;
	wire [1:0] w_n1223_0;
	wire [1:0] w_n1225_0;
	wire [1:0] w_n1228_0;
	wire [1:0] w_n1234_0;
	wire [2:0] w_n1236_0;
	wire [1:0] w_n1237_0;
	wire [1:0] w_n1241_0;
	wire [1:0] w_n1242_0;
	wire [1:0] w_n1244_0;
	wire [1:0] w_n1249_0;
	wire [1:0] w_n1251_0;
	wire [1:0] w_n1252_0;
	wire [2:0] w_n1253_0;
	wire [1:0] w_n1254_0;
	wire [1:0] w_n1258_0;
	wire [1:0] w_n1259_0;
	wire [1:0] w_n1261_0;
	wire [1:0] w_n1263_0;
	wire [1:0] w_n1266_0;
	wire [1:0] w_n1272_0;
	wire [1:0] w_n1274_0;
	wire [2:0] w_n1275_0;
	wire [1:0] w_n1279_0;
	wire [1:0] w_n1280_0;
	wire [2:0] w_n1281_0;
	wire [1:0] w_n1283_0;
	wire [1:0] w_n1288_0;
	wire [1:0] w_n1290_0;
	wire [1:0] w_n1291_0;
	wire [2:0] w_n1292_0;
	wire [2:0] w_n1292_1;
	wire [1:0] w_n1295_0;
	wire [2:0] w_n1296_0;
	wire [1:0] w_n1297_0;
	wire [1:0] w_n1298_0;
	wire [1:0] w_n1304_0;
	wire [2:0] w_n1305_0;
	wire [1:0] w_n1306_0;
	wire [1:0] w_n1311_0;
	wire [2:0] w_n1312_0;
	wire [2:0] w_n1312_1;
	wire [2:0] w_n1312_2;
	wire [2:0] w_n1312_3;
	wire [2:0] w_n1312_4;
	wire [2:0] w_n1312_5;
	wire [2:0] w_n1312_6;
	wire [2:0] w_n1312_7;
	wire [2:0] w_n1312_8;
	wire [2:0] w_n1312_9;
	wire [2:0] w_n1312_10;
	wire [2:0] w_n1312_11;
	wire [2:0] w_n1312_12;
	wire [2:0] w_n1312_13;
	wire [2:0] w_n1312_14;
	wire [2:0] w_n1312_15;
	wire [2:0] w_n1312_16;
	wire [2:0] w_n1312_17;
	wire [2:0] w_n1312_18;
	wire [2:0] w_n1312_19;
	wire [2:0] w_n1312_20;
	wire [2:0] w_n1312_21;
	wire [2:0] w_n1312_22;
	wire [2:0] w_n1312_23;
	wire [2:0] w_n1312_24;
	wire [2:0] w_n1312_25;
	wire [2:0] w_n1312_26;
	wire [2:0] w_n1312_27;
	wire [2:0] w_n1312_28;
	wire [2:0] w_n1312_29;
	wire [2:0] w_n1312_30;
	wire [2:0] w_n1312_31;
	wire [2:0] w_n1317_0;
	wire [2:0] w_n1317_1;
	wire [2:0] w_n1317_2;
	wire [2:0] w_n1317_3;
	wire [2:0] w_n1317_4;
	wire [2:0] w_n1317_5;
	wire [2:0] w_n1317_6;
	wire [2:0] w_n1317_7;
	wire [2:0] w_n1317_8;
	wire [2:0] w_n1317_9;
	wire [2:0] w_n1317_10;
	wire [2:0] w_n1317_11;
	wire [2:0] w_n1317_12;
	wire [2:0] w_n1317_13;
	wire [2:0] w_n1317_14;
	wire [2:0] w_n1317_15;
	wire [2:0] w_n1317_16;
	wire [2:0] w_n1317_17;
	wire [2:0] w_n1317_18;
	wire [2:0] w_n1317_19;
	wire [2:0] w_n1317_20;
	wire [2:0] w_n1317_21;
	wire [2:0] w_n1317_22;
	wire [2:0] w_n1317_23;
	wire [2:0] w_n1317_24;
	wire [2:0] w_n1317_25;
	wire [2:0] w_n1317_26;
	wire [2:0] w_n1317_27;
	wire [2:0] w_n1317_28;
	wire [2:0] w_n1317_29;
	wire [2:0] w_n1317_30;
	wire [2:0] w_n1317_31;
	wire [2:0] w_n1317_32;
	wire [2:0] w_n1317_33;
	wire [2:0] w_n1317_34;
	wire [2:0] w_n1317_35;
	wire [1:0] w_n1317_36;
	wire [2:0] w_n1320_0;
	wire [1:0] w_n1320_1;
	wire [2:0] w_n1321_0;
	wire [2:0] w_n1325_0;
	wire [1:0] w_n1326_0;
	wire [1:0] w_n1327_0;
	wire [1:0] w_n1328_0;
	wire [1:0] w_n1330_0;
	wire [1:0] w_n1332_0;
	wire [1:0] w_n1334_0;
	wire [1:0] w_n1337_0;
	wire [1:0] w_n1342_0;
	wire [2:0] w_n1344_0;
	wire [1:0] w_n1345_0;
	wire [1:0] w_n1349_0;
	wire [1:0] w_n1350_0;
	wire [1:0] w_n1352_0;
	wire [1:0] w_n1356_0;
	wire [1:0] w_n1358_0;
	wire [1:0] w_n1359_0;
	wire [2:0] w_n1360_0;
	wire [1:0] w_n1361_0;
	wire [1:0] w_n1365_0;
	wire [1:0] w_n1367_0;
	wire [1:0] w_n1369_0;
	wire [1:0] w_n1371_0;
	wire [1:0] w_n1373_0;
	wire [1:0] w_n1379_0;
	wire [2:0] w_n1381_0;
	wire [1:0] w_n1382_0;
	wire [1:0] w_n1387_0;
	wire [1:0] w_n1389_0;
	wire [1:0] w_n1391_0;
	wire [1:0] w_n1395_0;
	wire [1:0] w_n1397_0;
	wire [1:0] w_n1398_0;
	wire [2:0] w_n1399_0;
	wire [1:0] w_n1400_0;
	wire [1:0] w_n1406_0;
	wire [1:0] w_n1407_0;
	wire [1:0] w_n1409_0;
	wire [1:0] w_n1411_0;
	wire [1:0] w_n1413_0;
	wire [1:0] w_n1419_0;
	wire [1:0] w_n1421_0;
	wire [2:0] w_n1422_0;
	wire [1:0] w_n1425_0;
	wire [1:0] w_n1426_0;
	wire [2:0] w_n1427_0;
	wire [1:0] w_n1429_0;
	wire [1:0] w_n1433_0;
	wire [1:0] w_n1435_0;
	wire [1:0] w_n1436_0;
	wire [2:0] w_n1437_0;
	wire [1:0] w_n1441_0;
	wire [1:0] w_n1447_0;
	wire [2:0] w_n1449_0;
	wire [1:0] w_n1451_0;
	wire [2:0] w_n1456_0;
	wire [1:0] w_n1457_0;
	wire [1:0] w_n1458_0;
	wire [1:0] w_n1463_0;
	wire [2:0] w_n1464_0;
	wire [1:0] w_n1469_0;
	wire [2:0] w_n1475_0;
	wire [1:0] w_n1475_1;
	wire [1:0] w_n1476_0;
	wire [2:0] w_n1479_0;
	wire [1:0] w_n1480_0;
	wire [1:0] w_n1481_0;
	wire [1:0] w_n1482_0;
	wire [1:0] w_n1484_0;
	wire [1:0] w_n1486_0;
	wire [1:0] w_n1488_0;
	wire [1:0] w_n1497_0;
	wire [2:0] w_n1499_0;
	wire [1:0] w_n1500_0;
	wire [1:0] w_n1504_0;
	wire [1:0] w_n1506_0;
	wire [1:0] w_n1508_0;
	wire [1:0] w_n1513_0;
	wire [1:0] w_n1515_0;
	wire [1:0] w_n1516_0;
	wire [2:0] w_n1517_0;
	wire [1:0] w_n1518_0;
	wire [1:0] w_n1523_0;
	wire [1:0] w_n1524_0;
	wire [1:0] w_n1526_0;
	wire [1:0] w_n1528_0;
	wire [1:0] w_n1531_0;
	wire [1:0] w_n1537_0;
	wire [2:0] w_n1539_0;
	wire [1:0] w_n1540_0;
	wire [1:0] w_n1544_0;
	wire [1:0] w_n1545_0;
	wire [1:0] w_n1547_0;
	wire [1:0] w_n1552_0;
	wire [1:0] w_n1554_0;
	wire [1:0] w_n1555_0;
	wire [2:0] w_n1556_0;
	wire [1:0] w_n1557_0;
	wire [1:0] w_n1561_0;
	wire [1:0] w_n1562_0;
	wire [1:0] w_n1564_0;
	wire [1:0] w_n1566_0;
	wire [1:0] w_n1569_0;
	wire [1:0] w_n1575_0;
	wire [1:0] w_n1577_0;
	wire [2:0] w_n1578_0;
	wire [1:0] w_n1582_0;
	wire [1:0] w_n1583_0;
	wire [2:0] w_n1584_0;
	wire [1:0] w_n1586_0;
	wire [1:0] w_n1591_0;
	wire [1:0] w_n1593_0;
	wire [1:0] w_n1594_0;
	wire [2:0] w_n1595_0;
	wire [1:0] w_n1596_0;
	wire [1:0] w_n1600_0;
	wire [1:0] w_n1606_0;
	wire [1:0] w_n1607_0;
	wire [1:0] w_n1609_0;
	wire [1:0] w_n1611_0;
	wire [1:0] w_n1614_0;
	wire [1:0] w_n1620_0;
	wire [2:0] w_n1622_0;
	wire [2:0] w_n1622_1;
	wire [1:0] w_n1625_0;
	wire [2:0] w_n1626_0;
	wire [1:0] w_n1627_0;
	wire [1:0] w_n1633_0;
	wire [2:0] w_n1634_0;
	wire [1:0] w_n1635_0;
	wire [1:0] w_n1640_0;
	wire [2:0] w_n1641_0;
	wire [2:0] w_n1641_1;
	wire [2:0] w_n1641_2;
	wire [2:0] w_n1641_3;
	wire [2:0] w_n1641_4;
	wire [2:0] w_n1641_5;
	wire [2:0] w_n1641_6;
	wire [2:0] w_n1641_7;
	wire [2:0] w_n1641_8;
	wire [2:0] w_n1641_9;
	wire [2:0] w_n1641_10;
	wire [2:0] w_n1641_11;
	wire [2:0] w_n1641_12;
	wire [2:0] w_n1641_13;
	wire [2:0] w_n1641_14;
	wire [2:0] w_n1641_15;
	wire [2:0] w_n1641_16;
	wire [2:0] w_n1641_17;
	wire [2:0] w_n1641_18;
	wire [2:0] w_n1641_19;
	wire [2:0] w_n1641_20;
	wire [2:0] w_n1641_21;
	wire [2:0] w_n1641_22;
	wire [2:0] w_n1641_23;
	wire [2:0] w_n1641_24;
	wire [2:0] w_n1641_25;
	wire [2:0] w_n1641_26;
	wire [2:0] w_n1641_27;
	wire [2:0] w_n1641_28;
	wire [2:0] w_n1641_29;
	wire [2:0] w_n1641_30;
	wire [2:0] w_n1646_0;
	wire [2:0] w_n1646_1;
	wire [2:0] w_n1646_2;
	wire [2:0] w_n1646_3;
	wire [2:0] w_n1646_4;
	wire [2:0] w_n1646_5;
	wire [2:0] w_n1646_6;
	wire [2:0] w_n1646_7;
	wire [2:0] w_n1646_8;
	wire [2:0] w_n1646_9;
	wire [2:0] w_n1646_10;
	wire [2:0] w_n1646_11;
	wire [2:0] w_n1646_12;
	wire [2:0] w_n1646_13;
	wire [2:0] w_n1646_14;
	wire [2:0] w_n1646_15;
	wire [2:0] w_n1646_16;
	wire [2:0] w_n1646_17;
	wire [2:0] w_n1646_18;
	wire [2:0] w_n1646_19;
	wire [2:0] w_n1646_20;
	wire [2:0] w_n1646_21;
	wire [2:0] w_n1646_22;
	wire [2:0] w_n1646_23;
	wire [2:0] w_n1646_24;
	wire [2:0] w_n1646_25;
	wire [2:0] w_n1646_26;
	wire [2:0] w_n1646_27;
	wire [2:0] w_n1646_28;
	wire [2:0] w_n1646_29;
	wire [2:0] w_n1646_30;
	wire [2:0] w_n1646_31;
	wire [2:0] w_n1646_32;
	wire [2:0] w_n1646_33;
	wire [2:0] w_n1646_34;
	wire [2:0] w_n1646_35;
	wire [1:0] w_n1646_36;
	wire [2:0] w_n1649_0;
	wire [1:0] w_n1649_1;
	wire [2:0] w_n1650_0;
	wire [2:0] w_n1654_0;
	wire [1:0] w_n1655_0;
	wire [1:0] w_n1656_0;
	wire [1:0] w_n1657_0;
	wire [1:0] w_n1659_0;
	wire [1:0] w_n1661_0;
	wire [1:0] w_n1663_0;
	wire [1:0] w_n1666_0;
	wire [1:0] w_n1671_0;
	wire [2:0] w_n1673_0;
	wire [1:0] w_n1674_0;
	wire [1:0] w_n1678_0;
	wire [1:0] w_n1679_0;
	wire [1:0] w_n1681_0;
	wire [1:0] w_n1685_0;
	wire [1:0] w_n1687_0;
	wire [1:0] w_n1688_0;
	wire [2:0] w_n1689_0;
	wire [1:0] w_n1690_0;
	wire [1:0] w_n1694_0;
	wire [1:0] w_n1696_0;
	wire [1:0] w_n1698_0;
	wire [1:0] w_n1700_0;
	wire [1:0] w_n1702_0;
	wire [1:0] w_n1708_0;
	wire [2:0] w_n1710_0;
	wire [1:0] w_n1711_0;
	wire [1:0] w_n1716_0;
	wire [1:0] w_n1718_0;
	wire [1:0] w_n1720_0;
	wire [1:0] w_n1724_0;
	wire [1:0] w_n1726_0;
	wire [1:0] w_n1727_0;
	wire [2:0] w_n1728_0;
	wire [1:0] w_n1729_0;
	wire [1:0] w_n1735_0;
	wire [1:0] w_n1736_0;
	wire [1:0] w_n1738_0;
	wire [1:0] w_n1740_0;
	wire [1:0] w_n1742_0;
	wire [1:0] w_n1748_0;
	wire [1:0] w_n1750_0;
	wire [2:0] w_n1751_0;
	wire [1:0] w_n1754_0;
	wire [1:0] w_n1755_0;
	wire [2:0] w_n1756_0;
	wire [1:0] w_n1758_0;
	wire [1:0] w_n1762_0;
	wire [1:0] w_n1764_0;
	wire [1:0] w_n1765_0;
	wire [2:0] w_n1766_0;
	wire [1:0] w_n1767_0;
	wire [1:0] w_n1770_0;
	wire [1:0] w_n1776_0;
	wire [1:0] w_n1777_0;
	wire [1:0] w_n1779_0;
	wire [1:0] w_n1781_0;
	wire [1:0] w_n1783_0;
	wire [1:0] w_n1789_0;
	wire [2:0] w_n1791_0;
	wire [1:0] w_n1796_0;
	wire [2:0] w_n1798_0;
	wire [2:0] w_n1802_0;
	wire [1:0] w_n1803_0;
	wire [1:0] w_n1808_0;
	wire [2:0] w_n1809_0;
	wire [1:0] w_n1814_0;
	wire [2:0] w_n1820_0;
	wire [1:0] w_n1820_1;
	wire [1:0] w_n1821_0;
	wire [2:0] w_n1824_0;
	wire [1:0] w_n1825_0;
	wire [1:0] w_n1826_0;
	wire [1:0] w_n1827_0;
	wire [1:0] w_n1829_0;
	wire [1:0] w_n1831_0;
	wire [1:0] w_n1833_0;
	wire [1:0] w_n1842_0;
	wire [2:0] w_n1844_0;
	wire [1:0] w_n1845_0;
	wire [1:0] w_n1849_0;
	wire [1:0] w_n1851_0;
	wire [1:0] w_n1853_0;
	wire [1:0] w_n1858_0;
	wire [1:0] w_n1860_0;
	wire [1:0] w_n1861_0;
	wire [2:0] w_n1862_0;
	wire [1:0] w_n1863_0;
	wire [1:0] w_n1868_0;
	wire [1:0] w_n1869_0;
	wire [1:0] w_n1871_0;
	wire [1:0] w_n1873_0;
	wire [1:0] w_n1876_0;
	wire [1:0] w_n1882_0;
	wire [2:0] w_n1884_0;
	wire [1:0] w_n1885_0;
	wire [1:0] w_n1889_0;
	wire [1:0] w_n1890_0;
	wire [1:0] w_n1892_0;
	wire [1:0] w_n1897_0;
	wire [1:0] w_n1899_0;
	wire [1:0] w_n1900_0;
	wire [2:0] w_n1901_0;
	wire [1:0] w_n1902_0;
	wire [1:0] w_n1906_0;
	wire [1:0] w_n1907_0;
	wire [1:0] w_n1909_0;
	wire [1:0] w_n1911_0;
	wire [1:0] w_n1914_0;
	wire [1:0] w_n1920_0;
	wire [1:0] w_n1922_0;
	wire [2:0] w_n1923_0;
	wire [1:0] w_n1927_0;
	wire [1:0] w_n1928_0;
	wire [2:0] w_n1929_0;
	wire [1:0] w_n1931_0;
	wire [1:0] w_n1936_0;
	wire [1:0] w_n1938_0;
	wire [1:0] w_n1939_0;
	wire [2:0] w_n1940_0;
	wire [1:0] w_n1941_0;
	wire [1:0] w_n1945_0;
	wire [1:0] w_n1951_0;
	wire [1:0] w_n1952_0;
	wire [1:0] w_n1954_0;
	wire [1:0] w_n1956_0;
	wire [1:0] w_n1959_0;
	wire [1:0] w_n1965_0;
	wire [1:0] w_n1967_0;
	wire [2:0] w_n1968_0;
	wire [1:0] w_n1972_0;
	wire [1:0] w_n1973_0;
	wire [2:0] w_n1974_0;
	wire [1:0] w_n1976_0;
	wire [1:0] w_n1981_0;
	wire [1:0] w_n1983_0;
	wire [1:0] w_n1984_0;
	wire [2:0] w_n1985_0;
	wire [2:0] w_n1985_1;
	wire [1:0] w_n1988_0;
	wire [2:0] w_n1989_0;
	wire [1:0] w_n1990_0;
	wire [1:0] w_n1991_0;
	wire [1:0] w_n1997_0;
	wire [2:0] w_n1998_0;
	wire [1:0] w_n1999_0;
	wire [1:0] w_n2004_0;
	wire [2:0] w_n2005_0;
	wire [2:0] w_n2005_1;
	wire [2:0] w_n2005_2;
	wire [2:0] w_n2005_3;
	wire [2:0] w_n2005_4;
	wire [2:0] w_n2005_5;
	wire [2:0] w_n2005_6;
	wire [2:0] w_n2005_7;
	wire [2:0] w_n2005_8;
	wire [2:0] w_n2005_9;
	wire [2:0] w_n2005_10;
	wire [2:0] w_n2005_11;
	wire [2:0] w_n2005_12;
	wire [2:0] w_n2005_13;
	wire [2:0] w_n2005_14;
	wire [2:0] w_n2005_15;
	wire [2:0] w_n2005_16;
	wire [2:0] w_n2005_17;
	wire [2:0] w_n2005_18;
	wire [2:0] w_n2005_19;
	wire [2:0] w_n2005_20;
	wire [2:0] w_n2005_21;
	wire [2:0] w_n2005_22;
	wire [2:0] w_n2005_23;
	wire [2:0] w_n2005_24;
	wire [2:0] w_n2005_25;
	wire [2:0] w_n2005_26;
	wire [2:0] w_n2005_27;
	wire [2:0] w_n2005_28;
	wire [1:0] w_n2005_29;
	wire [2:0] w_n2010_0;
	wire [2:0] w_n2010_1;
	wire [2:0] w_n2010_2;
	wire [2:0] w_n2010_3;
	wire [2:0] w_n2010_4;
	wire [2:0] w_n2010_5;
	wire [2:0] w_n2010_6;
	wire [2:0] w_n2010_7;
	wire [2:0] w_n2010_8;
	wire [2:0] w_n2010_9;
	wire [2:0] w_n2010_10;
	wire [2:0] w_n2010_11;
	wire [2:0] w_n2010_12;
	wire [2:0] w_n2010_13;
	wire [2:0] w_n2010_14;
	wire [2:0] w_n2010_15;
	wire [2:0] w_n2010_16;
	wire [2:0] w_n2010_17;
	wire [2:0] w_n2010_18;
	wire [2:0] w_n2010_19;
	wire [2:0] w_n2010_20;
	wire [2:0] w_n2010_21;
	wire [2:0] w_n2010_22;
	wire [2:0] w_n2010_23;
	wire [2:0] w_n2010_24;
	wire [2:0] w_n2010_25;
	wire [2:0] w_n2010_26;
	wire [2:0] w_n2010_27;
	wire [2:0] w_n2010_28;
	wire [2:0] w_n2010_29;
	wire [2:0] w_n2010_30;
	wire [2:0] w_n2010_31;
	wire [2:0] w_n2010_32;
	wire [2:0] w_n2010_33;
	wire [2:0] w_n2010_34;
	wire [2:0] w_n2013_0;
	wire [1:0] w_n2013_1;
	wire [2:0] w_n2014_0;
	wire [2:0] w_n2018_0;
	wire [1:0] w_n2019_0;
	wire [1:0] w_n2020_0;
	wire [1:0] w_n2021_0;
	wire [1:0] w_n2023_0;
	wire [1:0] w_n2025_0;
	wire [1:0] w_n2027_0;
	wire [1:0] w_n2030_0;
	wire [1:0] w_n2035_0;
	wire [2:0] w_n2037_0;
	wire [1:0] w_n2038_0;
	wire [1:0] w_n2042_0;
	wire [1:0] w_n2043_0;
	wire [1:0] w_n2045_0;
	wire [1:0] w_n2049_0;
	wire [1:0] w_n2051_0;
	wire [1:0] w_n2052_0;
	wire [2:0] w_n2053_0;
	wire [1:0] w_n2054_0;
	wire [1:0] w_n2058_0;
	wire [1:0] w_n2060_0;
	wire [1:0] w_n2062_0;
	wire [1:0] w_n2064_0;
	wire [1:0] w_n2066_0;
	wire [1:0] w_n2072_0;
	wire [2:0] w_n2074_0;
	wire [1:0] w_n2075_0;
	wire [1:0] w_n2080_0;
	wire [1:0] w_n2082_0;
	wire [1:0] w_n2084_0;
	wire [1:0] w_n2088_0;
	wire [1:0] w_n2090_0;
	wire [1:0] w_n2091_0;
	wire [2:0] w_n2092_0;
	wire [1:0] w_n2093_0;
	wire [1:0] w_n2099_0;
	wire [1:0] w_n2100_0;
	wire [1:0] w_n2102_0;
	wire [1:0] w_n2104_0;
	wire [1:0] w_n2106_0;
	wire [1:0] w_n2112_0;
	wire [1:0] w_n2114_0;
	wire [2:0] w_n2115_0;
	wire [1:0] w_n2118_0;
	wire [1:0] w_n2119_0;
	wire [2:0] w_n2120_0;
	wire [1:0] w_n2122_0;
	wire [1:0] w_n2126_0;
	wire [1:0] w_n2128_0;
	wire [1:0] w_n2129_0;
	wire [2:0] w_n2130_0;
	wire [1:0] w_n2131_0;
	wire [1:0] w_n2134_0;
	wire [1:0] w_n2140_0;
	wire [1:0] w_n2141_0;
	wire [1:0] w_n2143_0;
	wire [1:0] w_n2145_0;
	wire [1:0] w_n2147_0;
	wire [1:0] w_n2153_0;
	wire [1:0] w_n2155_0;
	wire [2:0] w_n2156_0;
	wire [1:0] w_n2159_0;
	wire [1:0] w_n2160_0;
	wire [2:0] w_n2161_0;
	wire [1:0] w_n2163_0;
	wire [1:0] w_n2167_0;
	wire [1:0] w_n2169_0;
	wire [1:0] w_n2170_0;
	wire [2:0] w_n2171_0;
	wire [1:0] w_n2175_0;
	wire [1:0] w_n2181_0;
	wire [2:0] w_n2183_0;
	wire [1:0] w_n2185_0;
	wire [2:0] w_n2190_0;
	wire [1:0] w_n2191_0;
	wire [1:0] w_n2192_0;
	wire [1:0] w_n2197_0;
	wire [2:0] w_n2198_0;
	wire [1:0] w_n2203_0;
	wire [2:0] w_n2209_0;
	wire [1:0] w_n2209_1;
	wire [1:0] w_n2210_0;
	wire [2:0] w_n2213_0;
	wire [1:0] w_n2214_0;
	wire [1:0] w_n2215_0;
	wire [1:0] w_n2216_0;
	wire [1:0] w_n2218_0;
	wire [1:0] w_n2220_0;
	wire [1:0] w_n2222_0;
	wire [1:0] w_n2231_0;
	wire [2:0] w_n2233_0;
	wire [1:0] w_n2234_0;
	wire [1:0] w_n2238_0;
	wire [1:0] w_n2240_0;
	wire [1:0] w_n2242_0;
	wire [1:0] w_n2247_0;
	wire [1:0] w_n2249_0;
	wire [1:0] w_n2250_0;
	wire [2:0] w_n2251_0;
	wire [1:0] w_n2252_0;
	wire [1:0] w_n2257_0;
	wire [1:0] w_n2258_0;
	wire [1:0] w_n2260_0;
	wire [1:0] w_n2262_0;
	wire [1:0] w_n2265_0;
	wire [1:0] w_n2271_0;
	wire [2:0] w_n2273_0;
	wire [1:0] w_n2274_0;
	wire [1:0] w_n2278_0;
	wire [1:0] w_n2279_0;
	wire [1:0] w_n2281_0;
	wire [1:0] w_n2286_0;
	wire [1:0] w_n2288_0;
	wire [1:0] w_n2289_0;
	wire [2:0] w_n2290_0;
	wire [1:0] w_n2291_0;
	wire [1:0] w_n2295_0;
	wire [1:0] w_n2296_0;
	wire [1:0] w_n2298_0;
	wire [1:0] w_n2300_0;
	wire [1:0] w_n2303_0;
	wire [1:0] w_n2309_0;
	wire [1:0] w_n2311_0;
	wire [2:0] w_n2312_0;
	wire [1:0] w_n2316_0;
	wire [1:0] w_n2317_0;
	wire [2:0] w_n2318_0;
	wire [1:0] w_n2320_0;
	wire [1:0] w_n2325_0;
	wire [1:0] w_n2327_0;
	wire [1:0] w_n2328_0;
	wire [2:0] w_n2329_0;
	wire [1:0] w_n2330_0;
	wire [1:0] w_n2334_0;
	wire [1:0] w_n2340_0;
	wire [1:0] w_n2341_0;
	wire [1:0] w_n2343_0;
	wire [1:0] w_n2345_0;
	wire [1:0] w_n2348_0;
	wire [1:0] w_n2354_0;
	wire [1:0] w_n2356_0;
	wire [2:0] w_n2357_0;
	wire [1:0] w_n2361_0;
	wire [1:0] w_n2362_0;
	wire [2:0] w_n2363_0;
	wire [1:0] w_n2365_0;
	wire [1:0] w_n2370_0;
	wire [1:0] w_n2372_0;
	wire [1:0] w_n2373_0;
	wire [2:0] w_n2374_0;
	wire [1:0] w_n2375_0;
	wire [1:0] w_n2379_0;
	wire [1:0] w_n2385_0;
	wire [1:0] w_n2386_0;
	wire [1:0] w_n2388_0;
	wire [1:0] w_n2390_0;
	wire [1:0] w_n2393_0;
	wire [1:0] w_n2399_0;
	wire [2:0] w_n2401_0;
	wire [2:0] w_n2401_1;
	wire [1:0] w_n2404_0;
	wire [2:0] w_n2405_0;
	wire [1:0] w_n2406_0;
	wire [1:0] w_n2412_0;
	wire [2:0] w_n2413_0;
	wire [1:0] w_n2414_0;
	wire [1:0] w_n2419_0;
	wire [2:0] w_n2420_0;
	wire [2:0] w_n2420_1;
	wire [2:0] w_n2420_2;
	wire [2:0] w_n2420_3;
	wire [2:0] w_n2420_4;
	wire [2:0] w_n2420_5;
	wire [2:0] w_n2420_6;
	wire [2:0] w_n2420_7;
	wire [2:0] w_n2420_8;
	wire [2:0] w_n2420_9;
	wire [2:0] w_n2420_10;
	wire [2:0] w_n2420_11;
	wire [2:0] w_n2420_12;
	wire [2:0] w_n2420_13;
	wire [2:0] w_n2420_14;
	wire [2:0] w_n2420_15;
	wire [2:0] w_n2420_16;
	wire [2:0] w_n2420_17;
	wire [2:0] w_n2420_18;
	wire [2:0] w_n2420_19;
	wire [2:0] w_n2420_20;
	wire [2:0] w_n2420_21;
	wire [2:0] w_n2420_22;
	wire [2:0] w_n2420_23;
	wire [2:0] w_n2420_24;
	wire [2:0] w_n2420_25;
	wire [2:0] w_n2420_26;
	wire [2:0] w_n2420_27;
	wire [1:0] w_n2420_28;
	wire [2:0] w_n2425_0;
	wire [2:0] w_n2425_1;
	wire [2:0] w_n2425_2;
	wire [2:0] w_n2425_3;
	wire [2:0] w_n2425_4;
	wire [2:0] w_n2425_5;
	wire [2:0] w_n2425_6;
	wire [2:0] w_n2425_7;
	wire [2:0] w_n2425_8;
	wire [2:0] w_n2425_9;
	wire [2:0] w_n2425_10;
	wire [2:0] w_n2425_11;
	wire [2:0] w_n2425_12;
	wire [2:0] w_n2425_13;
	wire [2:0] w_n2425_14;
	wire [2:0] w_n2425_15;
	wire [2:0] w_n2425_16;
	wire [2:0] w_n2425_17;
	wire [2:0] w_n2425_18;
	wire [2:0] w_n2425_19;
	wire [2:0] w_n2425_20;
	wire [2:0] w_n2425_21;
	wire [2:0] w_n2425_22;
	wire [2:0] w_n2425_23;
	wire [2:0] w_n2425_24;
	wire [2:0] w_n2425_25;
	wire [2:0] w_n2425_26;
	wire [2:0] w_n2425_27;
	wire [2:0] w_n2425_28;
	wire [2:0] w_n2425_29;
	wire [2:0] w_n2425_30;
	wire [2:0] w_n2425_31;
	wire [2:0] w_n2425_32;
	wire [2:0] w_n2425_33;
	wire [2:0] w_n2425_34;
	wire [2:0] w_n2428_0;
	wire [1:0] w_n2428_1;
	wire [2:0] w_n2429_0;
	wire [2:0] w_n2433_0;
	wire [1:0] w_n2434_0;
	wire [1:0] w_n2435_0;
	wire [1:0] w_n2436_0;
	wire [1:0] w_n2438_0;
	wire [1:0] w_n2440_0;
	wire [1:0] w_n2442_0;
	wire [1:0] w_n2445_0;
	wire [1:0] w_n2450_0;
	wire [2:0] w_n2452_0;
	wire [1:0] w_n2453_0;
	wire [1:0] w_n2457_0;
	wire [1:0] w_n2458_0;
	wire [1:0] w_n2460_0;
	wire [1:0] w_n2464_0;
	wire [1:0] w_n2466_0;
	wire [1:0] w_n2467_0;
	wire [2:0] w_n2468_0;
	wire [1:0] w_n2469_0;
	wire [1:0] w_n2473_0;
	wire [1:0] w_n2475_0;
	wire [1:0] w_n2477_0;
	wire [1:0] w_n2479_0;
	wire [1:0] w_n2481_0;
	wire [1:0] w_n2487_0;
	wire [2:0] w_n2489_0;
	wire [1:0] w_n2490_0;
	wire [1:0] w_n2495_0;
	wire [1:0] w_n2497_0;
	wire [1:0] w_n2499_0;
	wire [1:0] w_n2503_0;
	wire [1:0] w_n2505_0;
	wire [1:0] w_n2506_0;
	wire [2:0] w_n2507_0;
	wire [1:0] w_n2508_0;
	wire [1:0] w_n2514_0;
	wire [1:0] w_n2515_0;
	wire [1:0] w_n2517_0;
	wire [1:0] w_n2519_0;
	wire [1:0] w_n2521_0;
	wire [1:0] w_n2527_0;
	wire [1:0] w_n2529_0;
	wire [2:0] w_n2530_0;
	wire [1:0] w_n2533_0;
	wire [1:0] w_n2534_0;
	wire [2:0] w_n2535_0;
	wire [1:0] w_n2537_0;
	wire [1:0] w_n2541_0;
	wire [1:0] w_n2543_0;
	wire [1:0] w_n2544_0;
	wire [2:0] w_n2545_0;
	wire [1:0] w_n2546_0;
	wire [1:0] w_n2549_0;
	wire [1:0] w_n2555_0;
	wire [1:0] w_n2556_0;
	wire [1:0] w_n2558_0;
	wire [1:0] w_n2560_0;
	wire [1:0] w_n2562_0;
	wire [1:0] w_n2568_0;
	wire [1:0] w_n2570_0;
	wire [2:0] w_n2571_0;
	wire [1:0] w_n2574_0;
	wire [1:0] w_n2575_0;
	wire [2:0] w_n2576_0;
	wire [1:0] w_n2578_0;
	wire [1:0] w_n2582_0;
	wire [1:0] w_n2584_0;
	wire [1:0] w_n2585_0;
	wire [2:0] w_n2586_0;
	wire [1:0] w_n2587_0;
	wire [1:0] w_n2590_0;
	wire [1:0] w_n2596_0;
	wire [1:0] w_n2597_0;
	wire [1:0] w_n2599_0;
	wire [1:0] w_n2601_0;
	wire [1:0] w_n2603_0;
	wire [1:0] w_n2609_0;
	wire [2:0] w_n2611_0;
	wire [1:0] w_n2616_0;
	wire [2:0] w_n2618_0;
	wire [2:0] w_n2622_0;
	wire [1:0] w_n2623_0;
	wire [1:0] w_n2628_0;
	wire [2:0] w_n2629_0;
	wire [1:0] w_n2634_0;
	wire [2:0] w_n2640_0;
	wire [1:0] w_n2640_1;
	wire [1:0] w_n2641_0;
	wire [2:0] w_n2644_0;
	wire [1:0] w_n2645_0;
	wire [1:0] w_n2646_0;
	wire [1:0] w_n2647_0;
	wire [1:0] w_n2649_0;
	wire [1:0] w_n2651_0;
	wire [1:0] w_n2653_0;
	wire [1:0] w_n2662_0;
	wire [2:0] w_n2664_0;
	wire [1:0] w_n2665_0;
	wire [1:0] w_n2669_0;
	wire [1:0] w_n2671_0;
	wire [1:0] w_n2673_0;
	wire [1:0] w_n2678_0;
	wire [1:0] w_n2680_0;
	wire [1:0] w_n2681_0;
	wire [2:0] w_n2682_0;
	wire [1:0] w_n2683_0;
	wire [1:0] w_n2688_0;
	wire [1:0] w_n2689_0;
	wire [1:0] w_n2691_0;
	wire [1:0] w_n2693_0;
	wire [1:0] w_n2696_0;
	wire [1:0] w_n2702_0;
	wire [2:0] w_n2704_0;
	wire [1:0] w_n2705_0;
	wire [1:0] w_n2709_0;
	wire [1:0] w_n2710_0;
	wire [1:0] w_n2712_0;
	wire [1:0] w_n2717_0;
	wire [1:0] w_n2719_0;
	wire [1:0] w_n2720_0;
	wire [2:0] w_n2721_0;
	wire [1:0] w_n2722_0;
	wire [1:0] w_n2726_0;
	wire [1:0] w_n2727_0;
	wire [1:0] w_n2729_0;
	wire [1:0] w_n2731_0;
	wire [1:0] w_n2734_0;
	wire [1:0] w_n2740_0;
	wire [1:0] w_n2742_0;
	wire [2:0] w_n2743_0;
	wire [1:0] w_n2747_0;
	wire [1:0] w_n2748_0;
	wire [2:0] w_n2749_0;
	wire [1:0] w_n2751_0;
	wire [1:0] w_n2756_0;
	wire [1:0] w_n2758_0;
	wire [1:0] w_n2759_0;
	wire [2:0] w_n2760_0;
	wire [1:0] w_n2761_0;
	wire [1:0] w_n2765_0;
	wire [1:0] w_n2771_0;
	wire [1:0] w_n2772_0;
	wire [1:0] w_n2774_0;
	wire [1:0] w_n2776_0;
	wire [1:0] w_n2779_0;
	wire [1:0] w_n2785_0;
	wire [1:0] w_n2787_0;
	wire [2:0] w_n2788_0;
	wire [1:0] w_n2792_0;
	wire [1:0] w_n2793_0;
	wire [2:0] w_n2794_0;
	wire [1:0] w_n2796_0;
	wire [1:0] w_n2801_0;
	wire [1:0] w_n2803_0;
	wire [1:0] w_n2804_0;
	wire [2:0] w_n2805_0;
	wire [1:0] w_n2806_0;
	wire [1:0] w_n2810_0;
	wire [1:0] w_n2816_0;
	wire [1:0] w_n2817_0;
	wire [1:0] w_n2819_0;
	wire [1:0] w_n2821_0;
	wire [1:0] w_n2824_0;
	wire [1:0] w_n2830_0;
	wire [1:0] w_n2832_0;
	wire [2:0] w_n2833_0;
	wire [1:0] w_n2837_0;
	wire [1:0] w_n2838_0;
	wire [2:0] w_n2839_0;
	wire [1:0] w_n2841_0;
	wire [1:0] w_n2846_0;
	wire [1:0] w_n2848_0;
	wire [1:0] w_n2849_0;
	wire [2:0] w_n2850_0;
	wire [2:0] w_n2850_1;
	wire [1:0] w_n2853_0;
	wire [2:0] w_n2854_0;
	wire [1:0] w_n2855_0;
	wire [1:0] w_n2856_0;
	wire [1:0] w_n2862_0;
	wire [2:0] w_n2863_0;
	wire [1:0] w_n2864_0;
	wire [1:0] w_n2869_0;
	wire [2:0] w_n2870_0;
	wire [2:0] w_n2870_1;
	wire [2:0] w_n2870_2;
	wire [2:0] w_n2870_3;
	wire [2:0] w_n2870_4;
	wire [2:0] w_n2870_5;
	wire [2:0] w_n2870_6;
	wire [2:0] w_n2870_7;
	wire [2:0] w_n2870_8;
	wire [2:0] w_n2870_9;
	wire [2:0] w_n2870_10;
	wire [2:0] w_n2870_11;
	wire [2:0] w_n2870_12;
	wire [2:0] w_n2870_13;
	wire [2:0] w_n2870_14;
	wire [2:0] w_n2870_15;
	wire [2:0] w_n2870_16;
	wire [2:0] w_n2870_17;
	wire [2:0] w_n2870_18;
	wire [2:0] w_n2870_19;
	wire [2:0] w_n2870_20;
	wire [2:0] w_n2870_21;
	wire [2:0] w_n2870_22;
	wire [2:0] w_n2870_23;
	wire [2:0] w_n2870_24;
	wire [2:0] w_n2870_25;
	wire [2:0] w_n2870_26;
	wire [2:0] w_n2875_0;
	wire [2:0] w_n2875_1;
	wire [2:0] w_n2875_2;
	wire [2:0] w_n2875_3;
	wire [2:0] w_n2875_4;
	wire [2:0] w_n2875_5;
	wire [2:0] w_n2875_6;
	wire [2:0] w_n2875_7;
	wire [2:0] w_n2875_8;
	wire [2:0] w_n2875_9;
	wire [2:0] w_n2875_10;
	wire [2:0] w_n2875_11;
	wire [2:0] w_n2875_12;
	wire [2:0] w_n2875_13;
	wire [2:0] w_n2875_14;
	wire [2:0] w_n2875_15;
	wire [2:0] w_n2875_16;
	wire [2:0] w_n2875_17;
	wire [2:0] w_n2875_18;
	wire [2:0] w_n2875_19;
	wire [2:0] w_n2875_20;
	wire [2:0] w_n2875_21;
	wire [2:0] w_n2875_22;
	wire [2:0] w_n2875_23;
	wire [2:0] w_n2875_24;
	wire [2:0] w_n2875_25;
	wire [2:0] w_n2875_26;
	wire [2:0] w_n2875_27;
	wire [2:0] w_n2875_28;
	wire [2:0] w_n2875_29;
	wire [2:0] w_n2875_30;
	wire [2:0] w_n2875_31;
	wire [2:0] w_n2875_32;
	wire [1:0] w_n2875_33;
	wire [2:0] w_n2878_0;
	wire [1:0] w_n2878_1;
	wire [2:0] w_n2879_0;
	wire [2:0] w_n2883_0;
	wire [1:0] w_n2884_0;
	wire [1:0] w_n2885_0;
	wire [1:0] w_n2886_0;
	wire [1:0] w_n2888_0;
	wire [1:0] w_n2890_0;
	wire [1:0] w_n2892_0;
	wire [1:0] w_n2895_0;
	wire [1:0] w_n2900_0;
	wire [2:0] w_n2902_0;
	wire [1:0] w_n2903_0;
	wire [1:0] w_n2907_0;
	wire [1:0] w_n2908_0;
	wire [1:0] w_n2910_0;
	wire [1:0] w_n2914_0;
	wire [1:0] w_n2916_0;
	wire [1:0] w_n2917_0;
	wire [2:0] w_n2918_0;
	wire [1:0] w_n2919_0;
	wire [1:0] w_n2923_0;
	wire [1:0] w_n2925_0;
	wire [1:0] w_n2927_0;
	wire [1:0] w_n2929_0;
	wire [1:0] w_n2931_0;
	wire [1:0] w_n2937_0;
	wire [2:0] w_n2939_0;
	wire [1:0] w_n2940_0;
	wire [1:0] w_n2945_0;
	wire [1:0] w_n2947_0;
	wire [1:0] w_n2949_0;
	wire [1:0] w_n2953_0;
	wire [1:0] w_n2955_0;
	wire [1:0] w_n2956_0;
	wire [2:0] w_n2957_0;
	wire [1:0] w_n2958_0;
	wire [1:0] w_n2964_0;
	wire [1:0] w_n2965_0;
	wire [1:0] w_n2967_0;
	wire [1:0] w_n2969_0;
	wire [1:0] w_n2971_0;
	wire [1:0] w_n2977_0;
	wire [1:0] w_n2979_0;
	wire [2:0] w_n2980_0;
	wire [1:0] w_n2983_0;
	wire [1:0] w_n2984_0;
	wire [2:0] w_n2985_0;
	wire [1:0] w_n2987_0;
	wire [1:0] w_n2991_0;
	wire [1:0] w_n2993_0;
	wire [1:0] w_n2994_0;
	wire [2:0] w_n2995_0;
	wire [1:0] w_n2996_0;
	wire [1:0] w_n2999_0;
	wire [1:0] w_n3005_0;
	wire [1:0] w_n3006_0;
	wire [1:0] w_n3008_0;
	wire [1:0] w_n3010_0;
	wire [1:0] w_n3012_0;
	wire [1:0] w_n3018_0;
	wire [1:0] w_n3020_0;
	wire [2:0] w_n3021_0;
	wire [1:0] w_n3024_0;
	wire [1:0] w_n3025_0;
	wire [2:0] w_n3026_0;
	wire [1:0] w_n3028_0;
	wire [1:0] w_n3032_0;
	wire [1:0] w_n3034_0;
	wire [1:0] w_n3035_0;
	wire [2:0] w_n3036_0;
	wire [1:0] w_n3037_0;
	wire [1:0] w_n3040_0;
	wire [1:0] w_n3046_0;
	wire [1:0] w_n3047_0;
	wire [1:0] w_n3049_0;
	wire [1:0] w_n3051_0;
	wire [1:0] w_n3053_0;
	wire [1:0] w_n3059_0;
	wire [1:0] w_n3061_0;
	wire [2:0] w_n3062_0;
	wire [1:0] w_n3065_0;
	wire [1:0] w_n3066_0;
	wire [2:0] w_n3067_0;
	wire [1:0] w_n3069_0;
	wire [1:0] w_n3073_0;
	wire [1:0] w_n3075_0;
	wire [1:0] w_n3076_0;
	wire [2:0] w_n3077_0;
	wire [1:0] w_n3081_0;
	wire [1:0] w_n3087_0;
	wire [2:0] w_n3089_0;
	wire [1:0] w_n3091_0;
	wire [2:0] w_n3096_0;
	wire [1:0] w_n3097_0;
	wire [1:0] w_n3098_0;
	wire [1:0] w_n3103_0;
	wire [2:0] w_n3104_0;
	wire [1:0] w_n3109_0;
	wire [2:0] w_n3115_0;
	wire [1:0] w_n3115_1;
	wire [1:0] w_n3116_0;
	wire [2:0] w_n3119_0;
	wire [1:0] w_n3120_0;
	wire [1:0] w_n3121_0;
	wire [1:0] w_n3122_0;
	wire [1:0] w_n3124_0;
	wire [1:0] w_n3126_0;
	wire [1:0] w_n3128_0;
	wire [1:0] w_n3137_0;
	wire [2:0] w_n3139_0;
	wire [1:0] w_n3140_0;
	wire [1:0] w_n3144_0;
	wire [1:0] w_n3146_0;
	wire [1:0] w_n3148_0;
	wire [1:0] w_n3153_0;
	wire [1:0] w_n3155_0;
	wire [1:0] w_n3156_0;
	wire [2:0] w_n3157_0;
	wire [1:0] w_n3158_0;
	wire [1:0] w_n3163_0;
	wire [1:0] w_n3164_0;
	wire [1:0] w_n3166_0;
	wire [1:0] w_n3168_0;
	wire [1:0] w_n3171_0;
	wire [1:0] w_n3177_0;
	wire [2:0] w_n3179_0;
	wire [1:0] w_n3180_0;
	wire [1:0] w_n3184_0;
	wire [1:0] w_n3185_0;
	wire [1:0] w_n3187_0;
	wire [1:0] w_n3192_0;
	wire [1:0] w_n3194_0;
	wire [1:0] w_n3195_0;
	wire [2:0] w_n3196_0;
	wire [1:0] w_n3197_0;
	wire [1:0] w_n3201_0;
	wire [1:0] w_n3202_0;
	wire [1:0] w_n3204_0;
	wire [1:0] w_n3206_0;
	wire [1:0] w_n3209_0;
	wire [1:0] w_n3215_0;
	wire [1:0] w_n3217_0;
	wire [2:0] w_n3218_0;
	wire [1:0] w_n3222_0;
	wire [1:0] w_n3223_0;
	wire [2:0] w_n3224_0;
	wire [1:0] w_n3226_0;
	wire [1:0] w_n3231_0;
	wire [1:0] w_n3233_0;
	wire [1:0] w_n3234_0;
	wire [2:0] w_n3235_0;
	wire [1:0] w_n3236_0;
	wire [1:0] w_n3240_0;
	wire [1:0] w_n3246_0;
	wire [1:0] w_n3247_0;
	wire [1:0] w_n3249_0;
	wire [1:0] w_n3251_0;
	wire [1:0] w_n3254_0;
	wire [1:0] w_n3260_0;
	wire [1:0] w_n3262_0;
	wire [2:0] w_n3263_0;
	wire [1:0] w_n3267_0;
	wire [1:0] w_n3268_0;
	wire [2:0] w_n3269_0;
	wire [1:0] w_n3271_0;
	wire [1:0] w_n3276_0;
	wire [1:0] w_n3278_0;
	wire [1:0] w_n3279_0;
	wire [2:0] w_n3280_0;
	wire [1:0] w_n3281_0;
	wire [1:0] w_n3285_0;
	wire [1:0] w_n3291_0;
	wire [1:0] w_n3292_0;
	wire [1:0] w_n3294_0;
	wire [1:0] w_n3296_0;
	wire [1:0] w_n3299_0;
	wire [1:0] w_n3305_0;
	wire [1:0] w_n3307_0;
	wire [2:0] w_n3308_0;
	wire [1:0] w_n3312_0;
	wire [1:0] w_n3313_0;
	wire [2:0] w_n3314_0;
	wire [1:0] w_n3316_0;
	wire [1:0] w_n3321_0;
	wire [1:0] w_n3323_0;
	wire [1:0] w_n3324_0;
	wire [2:0] w_n3325_0;
	wire [1:0] w_n3326_0;
	wire [1:0] w_n3330_0;
	wire [1:0] w_n3336_0;
	wire [1:0] w_n3337_0;
	wire [1:0] w_n3339_0;
	wire [1:0] w_n3341_0;
	wire [1:0] w_n3344_0;
	wire [1:0] w_n3350_0;
	wire [2:0] w_n3352_0;
	wire [2:0] w_n3352_1;
	wire [1:0] w_n3355_0;
	wire [2:0] w_n3356_0;
	wire [1:0] w_n3357_0;
	wire [1:0] w_n3363_0;
	wire [2:0] w_n3364_0;
	wire [1:0] w_n3365_0;
	wire [1:0] w_n3370_0;
	wire [2:0] w_n3371_0;
	wire [2:0] w_n3371_1;
	wire [2:0] w_n3371_2;
	wire [2:0] w_n3371_3;
	wire [2:0] w_n3371_4;
	wire [2:0] w_n3371_5;
	wire [2:0] w_n3371_6;
	wire [2:0] w_n3371_7;
	wire [2:0] w_n3371_8;
	wire [2:0] w_n3371_9;
	wire [2:0] w_n3371_10;
	wire [2:0] w_n3371_11;
	wire [2:0] w_n3371_12;
	wire [2:0] w_n3371_13;
	wire [2:0] w_n3371_14;
	wire [2:0] w_n3371_15;
	wire [2:0] w_n3371_16;
	wire [2:0] w_n3371_17;
	wire [2:0] w_n3371_18;
	wire [2:0] w_n3371_19;
	wire [2:0] w_n3371_20;
	wire [2:0] w_n3371_21;
	wire [2:0] w_n3371_22;
	wire [2:0] w_n3371_23;
	wire [2:0] w_n3371_24;
	wire [2:0] w_n3371_25;
	wire [2:0] w_n3376_0;
	wire [2:0] w_n3376_1;
	wire [2:0] w_n3376_2;
	wire [2:0] w_n3376_3;
	wire [2:0] w_n3376_4;
	wire [2:0] w_n3376_5;
	wire [2:0] w_n3376_6;
	wire [2:0] w_n3376_7;
	wire [2:0] w_n3376_8;
	wire [2:0] w_n3376_9;
	wire [2:0] w_n3376_10;
	wire [2:0] w_n3376_11;
	wire [2:0] w_n3376_12;
	wire [2:0] w_n3376_13;
	wire [2:0] w_n3376_14;
	wire [2:0] w_n3376_15;
	wire [2:0] w_n3376_16;
	wire [2:0] w_n3376_17;
	wire [2:0] w_n3376_18;
	wire [2:0] w_n3376_19;
	wire [2:0] w_n3376_20;
	wire [2:0] w_n3376_21;
	wire [2:0] w_n3376_22;
	wire [2:0] w_n3376_23;
	wire [2:0] w_n3376_24;
	wire [2:0] w_n3376_25;
	wire [2:0] w_n3376_26;
	wire [2:0] w_n3376_27;
	wire [2:0] w_n3376_28;
	wire [2:0] w_n3376_29;
	wire [2:0] w_n3376_30;
	wire [2:0] w_n3376_31;
	wire [2:0] w_n3376_32;
	wire [1:0] w_n3376_33;
	wire [2:0] w_n3379_0;
	wire [1:0] w_n3379_1;
	wire [2:0] w_n3380_0;
	wire [2:0] w_n3384_0;
	wire [1:0] w_n3385_0;
	wire [1:0] w_n3386_0;
	wire [1:0] w_n3387_0;
	wire [1:0] w_n3389_0;
	wire [1:0] w_n3391_0;
	wire [1:0] w_n3393_0;
	wire [1:0] w_n3396_0;
	wire [1:0] w_n3401_0;
	wire [2:0] w_n3403_0;
	wire [1:0] w_n3404_0;
	wire [1:0] w_n3408_0;
	wire [1:0] w_n3409_0;
	wire [1:0] w_n3411_0;
	wire [1:0] w_n3415_0;
	wire [1:0] w_n3417_0;
	wire [1:0] w_n3418_0;
	wire [2:0] w_n3419_0;
	wire [1:0] w_n3420_0;
	wire [1:0] w_n3424_0;
	wire [1:0] w_n3426_0;
	wire [1:0] w_n3428_0;
	wire [1:0] w_n3430_0;
	wire [1:0] w_n3432_0;
	wire [1:0] w_n3438_0;
	wire [2:0] w_n3440_0;
	wire [1:0] w_n3441_0;
	wire [1:0] w_n3446_0;
	wire [1:0] w_n3448_0;
	wire [1:0] w_n3450_0;
	wire [1:0] w_n3454_0;
	wire [1:0] w_n3456_0;
	wire [1:0] w_n3457_0;
	wire [2:0] w_n3458_0;
	wire [1:0] w_n3459_0;
	wire [1:0] w_n3465_0;
	wire [1:0] w_n3466_0;
	wire [1:0] w_n3468_0;
	wire [1:0] w_n3470_0;
	wire [1:0] w_n3472_0;
	wire [1:0] w_n3478_0;
	wire [1:0] w_n3480_0;
	wire [2:0] w_n3481_0;
	wire [1:0] w_n3484_0;
	wire [1:0] w_n3485_0;
	wire [2:0] w_n3486_0;
	wire [1:0] w_n3488_0;
	wire [1:0] w_n3492_0;
	wire [1:0] w_n3494_0;
	wire [1:0] w_n3495_0;
	wire [2:0] w_n3496_0;
	wire [1:0] w_n3497_0;
	wire [1:0] w_n3500_0;
	wire [1:0] w_n3506_0;
	wire [1:0] w_n3507_0;
	wire [1:0] w_n3509_0;
	wire [1:0] w_n3511_0;
	wire [1:0] w_n3513_0;
	wire [1:0] w_n3519_0;
	wire [1:0] w_n3521_0;
	wire [2:0] w_n3522_0;
	wire [1:0] w_n3525_0;
	wire [1:0] w_n3526_0;
	wire [2:0] w_n3527_0;
	wire [1:0] w_n3529_0;
	wire [1:0] w_n3533_0;
	wire [1:0] w_n3535_0;
	wire [1:0] w_n3536_0;
	wire [2:0] w_n3537_0;
	wire [1:0] w_n3538_0;
	wire [1:0] w_n3541_0;
	wire [1:0] w_n3547_0;
	wire [1:0] w_n3548_0;
	wire [1:0] w_n3550_0;
	wire [1:0] w_n3552_0;
	wire [1:0] w_n3554_0;
	wire [1:0] w_n3560_0;
	wire [1:0] w_n3562_0;
	wire [2:0] w_n3563_0;
	wire [1:0] w_n3566_0;
	wire [1:0] w_n3567_0;
	wire [2:0] w_n3568_0;
	wire [1:0] w_n3570_0;
	wire [1:0] w_n3574_0;
	wire [1:0] w_n3576_0;
	wire [1:0] w_n3577_0;
	wire [2:0] w_n3578_0;
	wire [1:0] w_n3579_0;
	wire [1:0] w_n3582_0;
	wire [1:0] w_n3588_0;
	wire [1:0] w_n3589_0;
	wire [1:0] w_n3591_0;
	wire [1:0] w_n3593_0;
	wire [1:0] w_n3595_0;
	wire [1:0] w_n3601_0;
	wire [2:0] w_n3603_0;
	wire [1:0] w_n3608_0;
	wire [2:0] w_n3610_0;
	wire [2:0] w_n3614_0;
	wire [1:0] w_n3615_0;
	wire [1:0] w_n3620_0;
	wire [2:0] w_n3621_0;
	wire [1:0] w_n3626_0;
	wire [2:0] w_n3632_0;
	wire [1:0] w_n3632_1;
	wire [1:0] w_n3633_0;
	wire [2:0] w_n3636_0;
	wire [1:0] w_n3637_0;
	wire [1:0] w_n3638_0;
	wire [1:0] w_n3639_0;
	wire [1:0] w_n3641_0;
	wire [1:0] w_n3643_0;
	wire [1:0] w_n3645_0;
	wire [1:0] w_n3654_0;
	wire [2:0] w_n3656_0;
	wire [1:0] w_n3657_0;
	wire [1:0] w_n3661_0;
	wire [1:0] w_n3663_0;
	wire [1:0] w_n3665_0;
	wire [1:0] w_n3670_0;
	wire [1:0] w_n3672_0;
	wire [1:0] w_n3673_0;
	wire [2:0] w_n3674_0;
	wire [1:0] w_n3675_0;
	wire [1:0] w_n3680_0;
	wire [1:0] w_n3681_0;
	wire [1:0] w_n3683_0;
	wire [1:0] w_n3685_0;
	wire [1:0] w_n3688_0;
	wire [1:0] w_n3694_0;
	wire [2:0] w_n3696_0;
	wire [1:0] w_n3697_0;
	wire [1:0] w_n3701_0;
	wire [1:0] w_n3702_0;
	wire [1:0] w_n3704_0;
	wire [1:0] w_n3709_0;
	wire [1:0] w_n3711_0;
	wire [1:0] w_n3712_0;
	wire [2:0] w_n3713_0;
	wire [1:0] w_n3714_0;
	wire [1:0] w_n3718_0;
	wire [1:0] w_n3719_0;
	wire [1:0] w_n3721_0;
	wire [1:0] w_n3723_0;
	wire [1:0] w_n3726_0;
	wire [1:0] w_n3732_0;
	wire [1:0] w_n3734_0;
	wire [2:0] w_n3735_0;
	wire [1:0] w_n3739_0;
	wire [1:0] w_n3740_0;
	wire [2:0] w_n3741_0;
	wire [1:0] w_n3743_0;
	wire [1:0] w_n3748_0;
	wire [1:0] w_n3750_0;
	wire [1:0] w_n3751_0;
	wire [2:0] w_n3752_0;
	wire [1:0] w_n3753_0;
	wire [1:0] w_n3757_0;
	wire [1:0] w_n3763_0;
	wire [1:0] w_n3764_0;
	wire [1:0] w_n3766_0;
	wire [1:0] w_n3768_0;
	wire [1:0] w_n3771_0;
	wire [1:0] w_n3777_0;
	wire [1:0] w_n3779_0;
	wire [2:0] w_n3780_0;
	wire [1:0] w_n3784_0;
	wire [1:0] w_n3785_0;
	wire [2:0] w_n3786_0;
	wire [1:0] w_n3788_0;
	wire [1:0] w_n3793_0;
	wire [1:0] w_n3795_0;
	wire [1:0] w_n3796_0;
	wire [2:0] w_n3797_0;
	wire [1:0] w_n3798_0;
	wire [1:0] w_n3802_0;
	wire [1:0] w_n3808_0;
	wire [1:0] w_n3809_0;
	wire [1:0] w_n3811_0;
	wire [1:0] w_n3813_0;
	wire [1:0] w_n3816_0;
	wire [1:0] w_n3822_0;
	wire [1:0] w_n3824_0;
	wire [2:0] w_n3825_0;
	wire [1:0] w_n3829_0;
	wire [1:0] w_n3830_0;
	wire [2:0] w_n3831_0;
	wire [1:0] w_n3833_0;
	wire [1:0] w_n3838_0;
	wire [1:0] w_n3840_0;
	wire [1:0] w_n3841_0;
	wire [2:0] w_n3842_0;
	wire [1:0] w_n3843_0;
	wire [1:0] w_n3847_0;
	wire [1:0] w_n3853_0;
	wire [1:0] w_n3854_0;
	wire [1:0] w_n3856_0;
	wire [1:0] w_n3858_0;
	wire [1:0] w_n3861_0;
	wire [1:0] w_n3867_0;
	wire [1:0] w_n3869_0;
	wire [2:0] w_n3870_0;
	wire [1:0] w_n3874_0;
	wire [1:0] w_n3875_0;
	wire [2:0] w_n3876_0;
	wire [1:0] w_n3878_0;
	wire [1:0] w_n3883_0;
	wire [1:0] w_n3885_0;
	wire [1:0] w_n3886_0;
	wire [2:0] w_n3887_0;
	wire [2:0] w_n3887_1;
	wire [1:0] w_n3890_0;
	wire [2:0] w_n3891_0;
	wire [1:0] w_n3892_0;
	wire [1:0] w_n3893_0;
	wire [1:0] w_n3899_0;
	wire [2:0] w_n3900_0;
	wire [1:0] w_n3901_0;
	wire [1:0] w_n3906_0;
	wire [2:0] w_n3907_0;
	wire [2:0] w_n3907_1;
	wire [2:0] w_n3907_2;
	wire [2:0] w_n3907_3;
	wire [2:0] w_n3907_4;
	wire [2:0] w_n3907_5;
	wire [2:0] w_n3907_6;
	wire [2:0] w_n3907_7;
	wire [2:0] w_n3907_8;
	wire [2:0] w_n3907_9;
	wire [2:0] w_n3907_10;
	wire [2:0] w_n3907_11;
	wire [2:0] w_n3907_12;
	wire [2:0] w_n3907_13;
	wire [2:0] w_n3907_14;
	wire [2:0] w_n3907_15;
	wire [2:0] w_n3907_16;
	wire [2:0] w_n3907_17;
	wire [2:0] w_n3907_18;
	wire [2:0] w_n3907_19;
	wire [2:0] w_n3907_20;
	wire [2:0] w_n3907_21;
	wire [2:0] w_n3907_22;
	wire [2:0] w_n3907_23;
	wire [1:0] w_n3907_24;
	wire [2:0] w_n3912_0;
	wire [2:0] w_n3912_1;
	wire [2:0] w_n3912_2;
	wire [2:0] w_n3912_3;
	wire [2:0] w_n3912_4;
	wire [2:0] w_n3912_5;
	wire [2:0] w_n3912_6;
	wire [2:0] w_n3912_7;
	wire [2:0] w_n3912_8;
	wire [2:0] w_n3912_9;
	wire [2:0] w_n3912_10;
	wire [2:0] w_n3912_11;
	wire [2:0] w_n3912_12;
	wire [2:0] w_n3912_13;
	wire [2:0] w_n3912_14;
	wire [2:0] w_n3912_15;
	wire [2:0] w_n3912_16;
	wire [2:0] w_n3912_17;
	wire [2:0] w_n3912_18;
	wire [2:0] w_n3912_19;
	wire [2:0] w_n3912_20;
	wire [2:0] w_n3912_21;
	wire [2:0] w_n3912_22;
	wire [2:0] w_n3912_23;
	wire [2:0] w_n3912_24;
	wire [2:0] w_n3912_25;
	wire [2:0] w_n3912_26;
	wire [2:0] w_n3912_27;
	wire [2:0] w_n3912_28;
	wire [2:0] w_n3912_29;
	wire [2:0] w_n3912_30;
	wire [2:0] w_n3912_31;
	wire [2:0] w_n3915_0;
	wire [1:0] w_n3915_1;
	wire [2:0] w_n3916_0;
	wire [2:0] w_n3920_0;
	wire [1:0] w_n3921_0;
	wire [1:0] w_n3922_0;
	wire [1:0] w_n3923_0;
	wire [1:0] w_n3925_0;
	wire [1:0] w_n3927_0;
	wire [1:0] w_n3929_0;
	wire [1:0] w_n3932_0;
	wire [1:0] w_n3937_0;
	wire [2:0] w_n3939_0;
	wire [1:0] w_n3940_0;
	wire [1:0] w_n3944_0;
	wire [1:0] w_n3945_0;
	wire [1:0] w_n3947_0;
	wire [1:0] w_n3951_0;
	wire [1:0] w_n3953_0;
	wire [1:0] w_n3954_0;
	wire [2:0] w_n3955_0;
	wire [1:0] w_n3956_0;
	wire [1:0] w_n3960_0;
	wire [1:0] w_n3962_0;
	wire [1:0] w_n3964_0;
	wire [1:0] w_n3966_0;
	wire [1:0] w_n3968_0;
	wire [1:0] w_n3974_0;
	wire [2:0] w_n3976_0;
	wire [1:0] w_n3977_0;
	wire [1:0] w_n3982_0;
	wire [1:0] w_n3984_0;
	wire [1:0] w_n3986_0;
	wire [1:0] w_n3990_0;
	wire [1:0] w_n3992_0;
	wire [1:0] w_n3993_0;
	wire [2:0] w_n3994_0;
	wire [1:0] w_n3995_0;
	wire [1:0] w_n4001_0;
	wire [1:0] w_n4002_0;
	wire [1:0] w_n4004_0;
	wire [1:0] w_n4006_0;
	wire [1:0] w_n4008_0;
	wire [1:0] w_n4014_0;
	wire [1:0] w_n4016_0;
	wire [2:0] w_n4017_0;
	wire [1:0] w_n4020_0;
	wire [1:0] w_n4021_0;
	wire [2:0] w_n4022_0;
	wire [1:0] w_n4024_0;
	wire [1:0] w_n4028_0;
	wire [1:0] w_n4030_0;
	wire [1:0] w_n4031_0;
	wire [2:0] w_n4032_0;
	wire [1:0] w_n4033_0;
	wire [1:0] w_n4036_0;
	wire [1:0] w_n4042_0;
	wire [1:0] w_n4043_0;
	wire [1:0] w_n4045_0;
	wire [1:0] w_n4047_0;
	wire [1:0] w_n4049_0;
	wire [1:0] w_n4055_0;
	wire [1:0] w_n4057_0;
	wire [2:0] w_n4058_0;
	wire [1:0] w_n4061_0;
	wire [1:0] w_n4062_0;
	wire [2:0] w_n4063_0;
	wire [1:0] w_n4065_0;
	wire [1:0] w_n4069_0;
	wire [1:0] w_n4071_0;
	wire [1:0] w_n4072_0;
	wire [2:0] w_n4073_0;
	wire [1:0] w_n4074_0;
	wire [1:0] w_n4077_0;
	wire [1:0] w_n4083_0;
	wire [1:0] w_n4084_0;
	wire [1:0] w_n4086_0;
	wire [1:0] w_n4088_0;
	wire [1:0] w_n4090_0;
	wire [1:0] w_n4096_0;
	wire [1:0] w_n4098_0;
	wire [2:0] w_n4099_0;
	wire [1:0] w_n4102_0;
	wire [1:0] w_n4103_0;
	wire [2:0] w_n4104_0;
	wire [1:0] w_n4106_0;
	wire [1:0] w_n4110_0;
	wire [1:0] w_n4112_0;
	wire [1:0] w_n4113_0;
	wire [2:0] w_n4114_0;
	wire [1:0] w_n4115_0;
	wire [1:0] w_n4118_0;
	wire [1:0] w_n4124_0;
	wire [1:0] w_n4125_0;
	wire [1:0] w_n4127_0;
	wire [1:0] w_n4129_0;
	wire [1:0] w_n4131_0;
	wire [1:0] w_n4137_0;
	wire [1:0] w_n4139_0;
	wire [2:0] w_n4140_0;
	wire [1:0] w_n4143_0;
	wire [1:0] w_n4144_0;
	wire [2:0] w_n4145_0;
	wire [1:0] w_n4147_0;
	wire [1:0] w_n4151_0;
	wire [1:0] w_n4153_0;
	wire [1:0] w_n4154_0;
	wire [2:0] w_n4155_0;
	wire [1:0] w_n4159_0;
	wire [1:0] w_n4165_0;
	wire [2:0] w_n4167_0;
	wire [1:0] w_n4169_0;
	wire [2:0] w_n4174_0;
	wire [1:0] w_n4175_0;
	wire [1:0] w_n4176_0;
	wire [1:0] w_n4181_0;
	wire [2:0] w_n4182_0;
	wire [1:0] w_n4187_0;
	wire [2:0] w_n4193_0;
	wire [1:0] w_n4193_1;
	wire [1:0] w_n4194_0;
	wire [2:0] w_n4197_0;
	wire [1:0] w_n4198_0;
	wire [1:0] w_n4199_0;
	wire [1:0] w_n4200_0;
	wire [1:0] w_n4202_0;
	wire [1:0] w_n4204_0;
	wire [1:0] w_n4206_0;
	wire [1:0] w_n4215_0;
	wire [2:0] w_n4217_0;
	wire [1:0] w_n4218_0;
	wire [1:0] w_n4222_0;
	wire [1:0] w_n4224_0;
	wire [1:0] w_n4226_0;
	wire [1:0] w_n4231_0;
	wire [1:0] w_n4233_0;
	wire [1:0] w_n4234_0;
	wire [2:0] w_n4235_0;
	wire [1:0] w_n4236_0;
	wire [1:0] w_n4241_0;
	wire [1:0] w_n4242_0;
	wire [1:0] w_n4244_0;
	wire [1:0] w_n4246_0;
	wire [1:0] w_n4249_0;
	wire [1:0] w_n4255_0;
	wire [2:0] w_n4257_0;
	wire [1:0] w_n4258_0;
	wire [1:0] w_n4262_0;
	wire [1:0] w_n4263_0;
	wire [1:0] w_n4265_0;
	wire [1:0] w_n4270_0;
	wire [1:0] w_n4272_0;
	wire [1:0] w_n4273_0;
	wire [2:0] w_n4274_0;
	wire [1:0] w_n4275_0;
	wire [1:0] w_n4279_0;
	wire [1:0] w_n4280_0;
	wire [1:0] w_n4282_0;
	wire [1:0] w_n4284_0;
	wire [1:0] w_n4287_0;
	wire [1:0] w_n4293_0;
	wire [1:0] w_n4295_0;
	wire [2:0] w_n4296_0;
	wire [1:0] w_n4300_0;
	wire [1:0] w_n4301_0;
	wire [2:0] w_n4302_0;
	wire [1:0] w_n4304_0;
	wire [1:0] w_n4309_0;
	wire [1:0] w_n4311_0;
	wire [1:0] w_n4312_0;
	wire [2:0] w_n4313_0;
	wire [1:0] w_n4314_0;
	wire [1:0] w_n4318_0;
	wire [1:0] w_n4324_0;
	wire [1:0] w_n4325_0;
	wire [1:0] w_n4327_0;
	wire [1:0] w_n4329_0;
	wire [1:0] w_n4332_0;
	wire [1:0] w_n4338_0;
	wire [1:0] w_n4340_0;
	wire [2:0] w_n4341_0;
	wire [1:0] w_n4345_0;
	wire [1:0] w_n4346_0;
	wire [2:0] w_n4347_0;
	wire [1:0] w_n4349_0;
	wire [1:0] w_n4354_0;
	wire [1:0] w_n4356_0;
	wire [1:0] w_n4357_0;
	wire [2:0] w_n4358_0;
	wire [1:0] w_n4359_0;
	wire [1:0] w_n4363_0;
	wire [1:0] w_n4369_0;
	wire [1:0] w_n4370_0;
	wire [1:0] w_n4372_0;
	wire [1:0] w_n4374_0;
	wire [1:0] w_n4377_0;
	wire [1:0] w_n4383_0;
	wire [1:0] w_n4385_0;
	wire [2:0] w_n4386_0;
	wire [1:0] w_n4390_0;
	wire [1:0] w_n4391_0;
	wire [2:0] w_n4392_0;
	wire [1:0] w_n4394_0;
	wire [1:0] w_n4399_0;
	wire [1:0] w_n4401_0;
	wire [1:0] w_n4402_0;
	wire [2:0] w_n4403_0;
	wire [1:0] w_n4404_0;
	wire [1:0] w_n4408_0;
	wire [1:0] w_n4414_0;
	wire [1:0] w_n4415_0;
	wire [1:0] w_n4417_0;
	wire [1:0] w_n4419_0;
	wire [1:0] w_n4422_0;
	wire [1:0] w_n4428_0;
	wire [1:0] w_n4430_0;
	wire [2:0] w_n4431_0;
	wire [1:0] w_n4435_0;
	wire [1:0] w_n4436_0;
	wire [2:0] w_n4437_0;
	wire [1:0] w_n4439_0;
	wire [1:0] w_n4444_0;
	wire [1:0] w_n4446_0;
	wire [1:0] w_n4447_0;
	wire [2:0] w_n4448_0;
	wire [1:0] w_n4449_0;
	wire [1:0] w_n4453_0;
	wire [1:0] w_n4459_0;
	wire [1:0] w_n4460_0;
	wire [1:0] w_n4462_0;
	wire [1:0] w_n4464_0;
	wire [1:0] w_n4467_0;
	wire [1:0] w_n4473_0;
	wire [2:0] w_n4475_0;
	wire [2:0] w_n4475_1;
	wire [1:0] w_n4478_0;
	wire [2:0] w_n4479_0;
	wire [1:0] w_n4480_0;
	wire [1:0] w_n4486_0;
	wire [2:0] w_n4487_0;
	wire [1:0] w_n4488_0;
	wire [1:0] w_n4493_0;
	wire [2:0] w_n4494_0;
	wire [2:0] w_n4494_1;
	wire [2:0] w_n4494_2;
	wire [2:0] w_n4494_3;
	wire [2:0] w_n4494_4;
	wire [2:0] w_n4494_5;
	wire [2:0] w_n4494_6;
	wire [2:0] w_n4494_7;
	wire [2:0] w_n4494_8;
	wire [2:0] w_n4494_9;
	wire [2:0] w_n4494_10;
	wire [2:0] w_n4494_11;
	wire [2:0] w_n4494_12;
	wire [2:0] w_n4494_13;
	wire [2:0] w_n4494_14;
	wire [2:0] w_n4494_15;
	wire [2:0] w_n4494_16;
	wire [2:0] w_n4494_17;
	wire [2:0] w_n4494_18;
	wire [2:0] w_n4494_19;
	wire [2:0] w_n4494_20;
	wire [2:0] w_n4494_21;
	wire [2:0] w_n4494_22;
	wire [1:0] w_n4494_23;
	wire [2:0] w_n4499_0;
	wire [2:0] w_n4499_1;
	wire [2:0] w_n4499_2;
	wire [2:0] w_n4499_3;
	wire [2:0] w_n4499_4;
	wire [2:0] w_n4499_5;
	wire [2:0] w_n4499_6;
	wire [2:0] w_n4499_7;
	wire [2:0] w_n4499_8;
	wire [2:0] w_n4499_9;
	wire [2:0] w_n4499_10;
	wire [2:0] w_n4499_11;
	wire [2:0] w_n4499_12;
	wire [2:0] w_n4499_13;
	wire [2:0] w_n4499_14;
	wire [2:0] w_n4499_15;
	wire [2:0] w_n4499_16;
	wire [2:0] w_n4499_17;
	wire [2:0] w_n4499_18;
	wire [2:0] w_n4499_19;
	wire [2:0] w_n4499_20;
	wire [2:0] w_n4499_21;
	wire [2:0] w_n4499_22;
	wire [2:0] w_n4499_23;
	wire [2:0] w_n4499_24;
	wire [2:0] w_n4499_25;
	wire [2:0] w_n4499_26;
	wire [2:0] w_n4499_27;
	wire [2:0] w_n4499_28;
	wire [2:0] w_n4499_29;
	wire [2:0] w_n4499_30;
	wire [1:0] w_n4499_31;
	wire [2:0] w_n4502_0;
	wire [1:0] w_n4502_1;
	wire [2:0] w_n4503_0;
	wire [2:0] w_n4507_0;
	wire [1:0] w_n4508_0;
	wire [1:0] w_n4509_0;
	wire [1:0] w_n4510_0;
	wire [1:0] w_n4512_0;
	wire [1:0] w_n4514_0;
	wire [1:0] w_n4516_0;
	wire [1:0] w_n4519_0;
	wire [1:0] w_n4524_0;
	wire [2:0] w_n4526_0;
	wire [1:0] w_n4527_0;
	wire [1:0] w_n4531_0;
	wire [1:0] w_n4532_0;
	wire [1:0] w_n4534_0;
	wire [1:0] w_n4538_0;
	wire [1:0] w_n4540_0;
	wire [1:0] w_n4541_0;
	wire [2:0] w_n4542_0;
	wire [1:0] w_n4543_0;
	wire [1:0] w_n4547_0;
	wire [1:0] w_n4549_0;
	wire [1:0] w_n4551_0;
	wire [1:0] w_n4553_0;
	wire [1:0] w_n4555_0;
	wire [1:0] w_n4561_0;
	wire [2:0] w_n4563_0;
	wire [1:0] w_n4564_0;
	wire [1:0] w_n4569_0;
	wire [1:0] w_n4571_0;
	wire [1:0] w_n4573_0;
	wire [1:0] w_n4577_0;
	wire [1:0] w_n4579_0;
	wire [1:0] w_n4580_0;
	wire [2:0] w_n4581_0;
	wire [1:0] w_n4582_0;
	wire [1:0] w_n4588_0;
	wire [1:0] w_n4589_0;
	wire [1:0] w_n4591_0;
	wire [1:0] w_n4593_0;
	wire [1:0] w_n4595_0;
	wire [1:0] w_n4601_0;
	wire [1:0] w_n4603_0;
	wire [2:0] w_n4604_0;
	wire [1:0] w_n4607_0;
	wire [1:0] w_n4608_0;
	wire [2:0] w_n4609_0;
	wire [1:0] w_n4611_0;
	wire [1:0] w_n4615_0;
	wire [1:0] w_n4617_0;
	wire [1:0] w_n4618_0;
	wire [2:0] w_n4619_0;
	wire [1:0] w_n4620_0;
	wire [1:0] w_n4623_0;
	wire [1:0] w_n4629_0;
	wire [1:0] w_n4630_0;
	wire [1:0] w_n4632_0;
	wire [1:0] w_n4634_0;
	wire [1:0] w_n4636_0;
	wire [1:0] w_n4642_0;
	wire [1:0] w_n4644_0;
	wire [2:0] w_n4645_0;
	wire [1:0] w_n4648_0;
	wire [1:0] w_n4649_0;
	wire [2:0] w_n4650_0;
	wire [1:0] w_n4652_0;
	wire [1:0] w_n4656_0;
	wire [1:0] w_n4658_0;
	wire [1:0] w_n4659_0;
	wire [2:0] w_n4660_0;
	wire [1:0] w_n4661_0;
	wire [1:0] w_n4664_0;
	wire [1:0] w_n4670_0;
	wire [1:0] w_n4671_0;
	wire [1:0] w_n4673_0;
	wire [1:0] w_n4675_0;
	wire [1:0] w_n4677_0;
	wire [1:0] w_n4683_0;
	wire [1:0] w_n4685_0;
	wire [2:0] w_n4686_0;
	wire [1:0] w_n4689_0;
	wire [1:0] w_n4690_0;
	wire [2:0] w_n4691_0;
	wire [1:0] w_n4693_0;
	wire [1:0] w_n4697_0;
	wire [1:0] w_n4699_0;
	wire [1:0] w_n4700_0;
	wire [2:0] w_n4701_0;
	wire [1:0] w_n4702_0;
	wire [1:0] w_n4705_0;
	wire [1:0] w_n4711_0;
	wire [1:0] w_n4712_0;
	wire [1:0] w_n4714_0;
	wire [1:0] w_n4716_0;
	wire [1:0] w_n4718_0;
	wire [1:0] w_n4724_0;
	wire [1:0] w_n4726_0;
	wire [2:0] w_n4727_0;
	wire [1:0] w_n4730_0;
	wire [1:0] w_n4731_0;
	wire [2:0] w_n4732_0;
	wire [1:0] w_n4734_0;
	wire [1:0] w_n4738_0;
	wire [1:0] w_n4740_0;
	wire [1:0] w_n4741_0;
	wire [2:0] w_n4742_0;
	wire [1:0] w_n4743_0;
	wire [1:0] w_n4746_0;
	wire [1:0] w_n4752_0;
	wire [1:0] w_n4753_0;
	wire [1:0] w_n4755_0;
	wire [1:0] w_n4757_0;
	wire [1:0] w_n4759_0;
	wire [1:0] w_n4765_0;
	wire [2:0] w_n4767_0;
	wire [1:0] w_n4772_0;
	wire [2:0] w_n4774_0;
	wire [2:0] w_n4778_0;
	wire [1:0] w_n4779_0;
	wire [1:0] w_n4784_0;
	wire [2:0] w_n4785_0;
	wire [1:0] w_n4790_0;
	wire [2:0] w_n4796_0;
	wire [1:0] w_n4796_1;
	wire [1:0] w_n4797_0;
	wire [2:0] w_n4800_0;
	wire [1:0] w_n4801_0;
	wire [1:0] w_n4802_0;
	wire [1:0] w_n4803_0;
	wire [1:0] w_n4805_0;
	wire [1:0] w_n4807_0;
	wire [1:0] w_n4809_0;
	wire [1:0] w_n4818_0;
	wire [2:0] w_n4820_0;
	wire [1:0] w_n4821_0;
	wire [1:0] w_n4825_0;
	wire [1:0] w_n4827_0;
	wire [1:0] w_n4829_0;
	wire [1:0] w_n4834_0;
	wire [1:0] w_n4836_0;
	wire [1:0] w_n4837_0;
	wire [2:0] w_n4838_0;
	wire [1:0] w_n4839_0;
	wire [1:0] w_n4844_0;
	wire [1:0] w_n4845_0;
	wire [1:0] w_n4847_0;
	wire [1:0] w_n4849_0;
	wire [1:0] w_n4852_0;
	wire [1:0] w_n4858_0;
	wire [2:0] w_n4860_0;
	wire [1:0] w_n4861_0;
	wire [1:0] w_n4865_0;
	wire [1:0] w_n4866_0;
	wire [1:0] w_n4868_0;
	wire [1:0] w_n4873_0;
	wire [1:0] w_n4875_0;
	wire [1:0] w_n4876_0;
	wire [2:0] w_n4877_0;
	wire [1:0] w_n4878_0;
	wire [1:0] w_n4882_0;
	wire [1:0] w_n4883_0;
	wire [1:0] w_n4885_0;
	wire [1:0] w_n4887_0;
	wire [1:0] w_n4890_0;
	wire [1:0] w_n4896_0;
	wire [1:0] w_n4898_0;
	wire [2:0] w_n4899_0;
	wire [1:0] w_n4903_0;
	wire [1:0] w_n4904_0;
	wire [2:0] w_n4905_0;
	wire [1:0] w_n4907_0;
	wire [1:0] w_n4912_0;
	wire [1:0] w_n4914_0;
	wire [1:0] w_n4915_0;
	wire [2:0] w_n4916_0;
	wire [1:0] w_n4917_0;
	wire [1:0] w_n4921_0;
	wire [1:0] w_n4927_0;
	wire [1:0] w_n4928_0;
	wire [1:0] w_n4930_0;
	wire [1:0] w_n4932_0;
	wire [1:0] w_n4935_0;
	wire [1:0] w_n4941_0;
	wire [1:0] w_n4943_0;
	wire [2:0] w_n4944_0;
	wire [1:0] w_n4948_0;
	wire [1:0] w_n4949_0;
	wire [2:0] w_n4950_0;
	wire [1:0] w_n4952_0;
	wire [1:0] w_n4957_0;
	wire [1:0] w_n4959_0;
	wire [1:0] w_n4960_0;
	wire [2:0] w_n4961_0;
	wire [1:0] w_n4962_0;
	wire [1:0] w_n4966_0;
	wire [1:0] w_n4972_0;
	wire [1:0] w_n4973_0;
	wire [1:0] w_n4975_0;
	wire [1:0] w_n4977_0;
	wire [1:0] w_n4980_0;
	wire [1:0] w_n4986_0;
	wire [1:0] w_n4988_0;
	wire [2:0] w_n4989_0;
	wire [1:0] w_n4993_0;
	wire [1:0] w_n4994_0;
	wire [2:0] w_n4995_0;
	wire [1:0] w_n4997_0;
	wire [1:0] w_n5002_0;
	wire [1:0] w_n5004_0;
	wire [1:0] w_n5005_0;
	wire [2:0] w_n5006_0;
	wire [1:0] w_n5007_0;
	wire [1:0] w_n5011_0;
	wire [1:0] w_n5017_0;
	wire [1:0] w_n5018_0;
	wire [1:0] w_n5020_0;
	wire [1:0] w_n5022_0;
	wire [1:0] w_n5025_0;
	wire [1:0] w_n5031_0;
	wire [1:0] w_n5033_0;
	wire [2:0] w_n5034_0;
	wire [1:0] w_n5038_0;
	wire [1:0] w_n5039_0;
	wire [2:0] w_n5040_0;
	wire [1:0] w_n5042_0;
	wire [1:0] w_n5047_0;
	wire [1:0] w_n5049_0;
	wire [1:0] w_n5050_0;
	wire [2:0] w_n5051_0;
	wire [1:0] w_n5052_0;
	wire [1:0] w_n5056_0;
	wire [1:0] w_n5062_0;
	wire [1:0] w_n5063_0;
	wire [1:0] w_n5065_0;
	wire [1:0] w_n5067_0;
	wire [1:0] w_n5070_0;
	wire [1:0] w_n5076_0;
	wire [1:0] w_n5078_0;
	wire [2:0] w_n5079_0;
	wire [1:0] w_n5083_0;
	wire [1:0] w_n5084_0;
	wire [2:0] w_n5085_0;
	wire [1:0] w_n5087_0;
	wire [1:0] w_n5092_0;
	wire [1:0] w_n5094_0;
	wire [1:0] w_n5095_0;
	wire [2:0] w_n5096_0;
	wire [2:0] w_n5096_1;
	wire [1:0] w_n5099_0;
	wire [2:0] w_n5100_0;
	wire [1:0] w_n5101_0;
	wire [1:0] w_n5102_0;
	wire [1:0] w_n5108_0;
	wire [2:0] w_n5109_0;
	wire [1:0] w_n5110_0;
	wire [1:0] w_n5115_0;
	wire [2:0] w_n5116_0;
	wire [2:0] w_n5116_1;
	wire [2:0] w_n5116_2;
	wire [2:0] w_n5116_3;
	wire [2:0] w_n5116_4;
	wire [2:0] w_n5116_5;
	wire [2:0] w_n5116_6;
	wire [2:0] w_n5116_7;
	wire [2:0] w_n5116_8;
	wire [2:0] w_n5116_9;
	wire [2:0] w_n5116_10;
	wire [2:0] w_n5116_11;
	wire [2:0] w_n5116_12;
	wire [2:0] w_n5116_13;
	wire [2:0] w_n5116_14;
	wire [2:0] w_n5116_15;
	wire [2:0] w_n5116_16;
	wire [2:0] w_n5116_17;
	wire [2:0] w_n5116_18;
	wire [2:0] w_n5116_19;
	wire [2:0] w_n5116_20;
	wire [2:0] w_n5116_21;
	wire [2:0] w_n5121_0;
	wire [2:0] w_n5121_1;
	wire [2:0] w_n5121_2;
	wire [2:0] w_n5121_3;
	wire [2:0] w_n5121_4;
	wire [2:0] w_n5121_5;
	wire [2:0] w_n5121_6;
	wire [2:0] w_n5121_7;
	wire [2:0] w_n5121_8;
	wire [2:0] w_n5121_9;
	wire [2:0] w_n5121_10;
	wire [2:0] w_n5121_11;
	wire [2:0] w_n5121_12;
	wire [2:0] w_n5121_13;
	wire [2:0] w_n5121_14;
	wire [2:0] w_n5121_15;
	wire [2:0] w_n5121_16;
	wire [2:0] w_n5121_17;
	wire [2:0] w_n5121_18;
	wire [2:0] w_n5121_19;
	wire [2:0] w_n5121_20;
	wire [2:0] w_n5121_21;
	wire [2:0] w_n5121_22;
	wire [2:0] w_n5121_23;
	wire [2:0] w_n5121_24;
	wire [2:0] w_n5121_25;
	wire [2:0] w_n5121_26;
	wire [2:0] w_n5121_27;
	wire [2:0] w_n5121_28;
	wire [2:0] w_n5121_29;
	wire [2:0] w_n5124_0;
	wire [1:0] w_n5124_1;
	wire [2:0] w_n5125_0;
	wire [2:0] w_n5129_0;
	wire [1:0] w_n5130_0;
	wire [1:0] w_n5131_0;
	wire [1:0] w_n5132_0;
	wire [1:0] w_n5134_0;
	wire [1:0] w_n5136_0;
	wire [1:0] w_n5138_0;
	wire [1:0] w_n5141_0;
	wire [1:0] w_n5146_0;
	wire [2:0] w_n5148_0;
	wire [1:0] w_n5149_0;
	wire [1:0] w_n5153_0;
	wire [1:0] w_n5154_0;
	wire [1:0] w_n5156_0;
	wire [1:0] w_n5160_0;
	wire [1:0] w_n5162_0;
	wire [1:0] w_n5163_0;
	wire [2:0] w_n5164_0;
	wire [1:0] w_n5165_0;
	wire [1:0] w_n5169_0;
	wire [1:0] w_n5171_0;
	wire [1:0] w_n5173_0;
	wire [1:0] w_n5175_0;
	wire [1:0] w_n5177_0;
	wire [1:0] w_n5183_0;
	wire [2:0] w_n5185_0;
	wire [1:0] w_n5186_0;
	wire [1:0] w_n5191_0;
	wire [1:0] w_n5193_0;
	wire [1:0] w_n5195_0;
	wire [1:0] w_n5199_0;
	wire [1:0] w_n5201_0;
	wire [1:0] w_n5202_0;
	wire [2:0] w_n5203_0;
	wire [1:0] w_n5204_0;
	wire [1:0] w_n5210_0;
	wire [1:0] w_n5211_0;
	wire [1:0] w_n5213_0;
	wire [1:0] w_n5215_0;
	wire [1:0] w_n5217_0;
	wire [1:0] w_n5223_0;
	wire [1:0] w_n5225_0;
	wire [2:0] w_n5226_0;
	wire [1:0] w_n5229_0;
	wire [1:0] w_n5230_0;
	wire [2:0] w_n5231_0;
	wire [1:0] w_n5233_0;
	wire [1:0] w_n5237_0;
	wire [1:0] w_n5239_0;
	wire [1:0] w_n5240_0;
	wire [2:0] w_n5241_0;
	wire [1:0] w_n5242_0;
	wire [1:0] w_n5245_0;
	wire [1:0] w_n5251_0;
	wire [1:0] w_n5252_0;
	wire [1:0] w_n5254_0;
	wire [1:0] w_n5256_0;
	wire [1:0] w_n5258_0;
	wire [1:0] w_n5264_0;
	wire [1:0] w_n5266_0;
	wire [2:0] w_n5267_0;
	wire [1:0] w_n5270_0;
	wire [1:0] w_n5271_0;
	wire [2:0] w_n5272_0;
	wire [1:0] w_n5274_0;
	wire [1:0] w_n5278_0;
	wire [1:0] w_n5280_0;
	wire [1:0] w_n5281_0;
	wire [2:0] w_n5282_0;
	wire [1:0] w_n5283_0;
	wire [1:0] w_n5286_0;
	wire [1:0] w_n5292_0;
	wire [1:0] w_n5293_0;
	wire [1:0] w_n5295_0;
	wire [1:0] w_n5297_0;
	wire [1:0] w_n5299_0;
	wire [1:0] w_n5305_0;
	wire [1:0] w_n5307_0;
	wire [2:0] w_n5308_0;
	wire [1:0] w_n5311_0;
	wire [1:0] w_n5312_0;
	wire [2:0] w_n5313_0;
	wire [1:0] w_n5315_0;
	wire [1:0] w_n5319_0;
	wire [1:0] w_n5321_0;
	wire [1:0] w_n5322_0;
	wire [2:0] w_n5323_0;
	wire [1:0] w_n5324_0;
	wire [1:0] w_n5327_0;
	wire [1:0] w_n5333_0;
	wire [1:0] w_n5334_0;
	wire [1:0] w_n5336_0;
	wire [1:0] w_n5338_0;
	wire [1:0] w_n5340_0;
	wire [1:0] w_n5346_0;
	wire [1:0] w_n5348_0;
	wire [2:0] w_n5349_0;
	wire [1:0] w_n5352_0;
	wire [1:0] w_n5353_0;
	wire [2:0] w_n5354_0;
	wire [1:0] w_n5356_0;
	wire [1:0] w_n5360_0;
	wire [1:0] w_n5362_0;
	wire [1:0] w_n5363_0;
	wire [2:0] w_n5364_0;
	wire [1:0] w_n5365_0;
	wire [1:0] w_n5368_0;
	wire [1:0] w_n5374_0;
	wire [1:0] w_n5375_0;
	wire [1:0] w_n5377_0;
	wire [1:0] w_n5379_0;
	wire [1:0] w_n5381_0;
	wire [1:0] w_n5387_0;
	wire [1:0] w_n5389_0;
	wire [2:0] w_n5390_0;
	wire [1:0] w_n5393_0;
	wire [1:0] w_n5394_0;
	wire [2:0] w_n5395_0;
	wire [1:0] w_n5397_0;
	wire [1:0] w_n5401_0;
	wire [1:0] w_n5403_0;
	wire [1:0] w_n5404_0;
	wire [2:0] w_n5405_0;
	wire [1:0] w_n5409_0;
	wire [1:0] w_n5415_0;
	wire [2:0] w_n5417_0;
	wire [1:0] w_n5419_0;
	wire [2:0] w_n5424_0;
	wire [1:0] w_n5425_0;
	wire [1:0] w_n5426_0;
	wire [1:0] w_n5431_0;
	wire [2:0] w_n5432_0;
	wire [1:0] w_n5437_0;
	wire [2:0] w_n5443_0;
	wire [1:0] w_n5443_1;
	wire [2:0] w_n5446_0;
	wire [1:0] w_n5447_0;
	wire [1:0] w_n5448_0;
	wire [1:0] w_n5449_0;
	wire [1:0] w_n5451_0;
	wire [1:0] w_n5453_0;
	wire [1:0] w_n5455_0;
	wire [1:0] w_n5464_0;
	wire [2:0] w_n5466_0;
	wire [1:0] w_n5467_0;
	wire [1:0] w_n5471_0;
	wire [1:0] w_n5473_0;
	wire [1:0] w_n5475_0;
	wire [1:0] w_n5480_0;
	wire [1:0] w_n5482_0;
	wire [1:0] w_n5483_0;
	wire [2:0] w_n5484_0;
	wire [1:0] w_n5485_0;
	wire [1:0] w_n5490_0;
	wire [1:0] w_n5491_0;
	wire [1:0] w_n5493_0;
	wire [1:0] w_n5495_0;
	wire [1:0] w_n5498_0;
	wire [1:0] w_n5504_0;
	wire [2:0] w_n5506_0;
	wire [1:0] w_n5507_0;
	wire [1:0] w_n5511_0;
	wire [1:0] w_n5512_0;
	wire [1:0] w_n5514_0;
	wire [1:0] w_n5519_0;
	wire [1:0] w_n5521_0;
	wire [1:0] w_n5522_0;
	wire [2:0] w_n5523_0;
	wire [1:0] w_n5524_0;
	wire [1:0] w_n5528_0;
	wire [1:0] w_n5529_0;
	wire [1:0] w_n5531_0;
	wire [1:0] w_n5533_0;
	wire [1:0] w_n5536_0;
	wire [1:0] w_n5542_0;
	wire [1:0] w_n5544_0;
	wire [2:0] w_n5545_0;
	wire [1:0] w_n5549_0;
	wire [1:0] w_n5550_0;
	wire [2:0] w_n5551_0;
	wire [1:0] w_n5553_0;
	wire [1:0] w_n5558_0;
	wire [1:0] w_n5560_0;
	wire [1:0] w_n5561_0;
	wire [2:0] w_n5562_0;
	wire [1:0] w_n5563_0;
	wire [1:0] w_n5567_0;
	wire [1:0] w_n5573_0;
	wire [1:0] w_n5574_0;
	wire [1:0] w_n5576_0;
	wire [1:0] w_n5578_0;
	wire [1:0] w_n5581_0;
	wire [1:0] w_n5587_0;
	wire [1:0] w_n5589_0;
	wire [2:0] w_n5590_0;
	wire [1:0] w_n5594_0;
	wire [1:0] w_n5595_0;
	wire [2:0] w_n5596_0;
	wire [1:0] w_n5598_0;
	wire [1:0] w_n5603_0;
	wire [1:0] w_n5605_0;
	wire [1:0] w_n5606_0;
	wire [2:0] w_n5607_0;
	wire [1:0] w_n5608_0;
	wire [1:0] w_n5612_0;
	wire [1:0] w_n5618_0;
	wire [1:0] w_n5619_0;
	wire [1:0] w_n5621_0;
	wire [1:0] w_n5623_0;
	wire [1:0] w_n5626_0;
	wire [1:0] w_n5632_0;
	wire [1:0] w_n5634_0;
	wire [2:0] w_n5635_0;
	wire [1:0] w_n5639_0;
	wire [1:0] w_n5640_0;
	wire [2:0] w_n5641_0;
	wire [1:0] w_n5643_0;
	wire [1:0] w_n5648_0;
	wire [1:0] w_n5650_0;
	wire [1:0] w_n5651_0;
	wire [2:0] w_n5652_0;
	wire [1:0] w_n5653_0;
	wire [1:0] w_n5657_0;
	wire [1:0] w_n5663_0;
	wire [1:0] w_n5664_0;
	wire [1:0] w_n5666_0;
	wire [1:0] w_n5668_0;
	wire [1:0] w_n5671_0;
	wire [1:0] w_n5677_0;
	wire [1:0] w_n5679_0;
	wire [2:0] w_n5680_0;
	wire [1:0] w_n5684_0;
	wire [1:0] w_n5685_0;
	wire [2:0] w_n5686_0;
	wire [1:0] w_n5688_0;
	wire [1:0] w_n5693_0;
	wire [1:0] w_n5695_0;
	wire [1:0] w_n5696_0;
	wire [2:0] w_n5697_0;
	wire [1:0] w_n5698_0;
	wire [1:0] w_n5702_0;
	wire [1:0] w_n5708_0;
	wire [1:0] w_n5709_0;
	wire [1:0] w_n5711_0;
	wire [1:0] w_n5713_0;
	wire [1:0] w_n5716_0;
	wire [1:0] w_n5722_0;
	wire [1:0] w_n5724_0;
	wire [2:0] w_n5725_0;
	wire [1:0] w_n5729_0;
	wire [1:0] w_n5730_0;
	wire [2:0] w_n5731_0;
	wire [1:0] w_n5733_0;
	wire [1:0] w_n5738_0;
	wire [1:0] w_n5740_0;
	wire [1:0] w_n5741_0;
	wire [2:0] w_n5742_0;
	wire [1:0] w_n5743_0;
	wire [1:0] w_n5747_0;
	wire [1:0] w_n5753_0;
	wire [1:0] w_n5754_0;
	wire [1:0] w_n5756_0;
	wire [1:0] w_n5758_0;
	wire [1:0] w_n5761_0;
	wire [1:0] w_n5767_0;
	wire [2:0] w_n5769_0;
	wire [2:0] w_n5769_1;
	wire [1:0] w_n5772_0;
	wire [2:0] w_n5773_0;
	wire [1:0] w_n5774_0;
	wire [1:0] w_n5780_0;
	wire [2:0] w_n5781_0;
	wire [1:0] w_n5782_0;
	wire [1:0] w_n5787_0;
	wire [2:0] w_n5788_0;
	wire [2:0] w_n5788_1;
	wire [2:0] w_n5788_2;
	wire [2:0] w_n5788_3;
	wire [2:0] w_n5788_4;
	wire [2:0] w_n5788_5;
	wire [2:0] w_n5788_6;
	wire [2:0] w_n5788_7;
	wire [2:0] w_n5788_8;
	wire [2:0] w_n5788_9;
	wire [2:0] w_n5788_10;
	wire [2:0] w_n5788_11;
	wire [2:0] w_n5788_12;
	wire [2:0] w_n5788_13;
	wire [2:0] w_n5788_14;
	wire [2:0] w_n5788_15;
	wire [2:0] w_n5788_16;
	wire [2:0] w_n5788_17;
	wire [2:0] w_n5788_18;
	wire [2:0] w_n5788_19;
	wire [2:0] w_n5788_20;
	wire [2:0] w_n5793_0;
	wire [2:0] w_n5793_1;
	wire [2:0] w_n5793_2;
	wire [2:0] w_n5793_3;
	wire [2:0] w_n5793_4;
	wire [2:0] w_n5793_5;
	wire [2:0] w_n5793_6;
	wire [2:0] w_n5793_7;
	wire [2:0] w_n5793_8;
	wire [2:0] w_n5793_9;
	wire [2:0] w_n5793_10;
	wire [2:0] w_n5793_11;
	wire [2:0] w_n5793_12;
	wire [2:0] w_n5793_13;
	wire [2:0] w_n5793_14;
	wire [2:0] w_n5793_15;
	wire [2:0] w_n5793_16;
	wire [2:0] w_n5793_17;
	wire [2:0] w_n5793_18;
	wire [2:0] w_n5793_19;
	wire [2:0] w_n5793_20;
	wire [2:0] w_n5793_21;
	wire [2:0] w_n5793_22;
	wire [2:0] w_n5793_23;
	wire [2:0] w_n5793_24;
	wire [2:0] w_n5793_25;
	wire [2:0] w_n5793_26;
	wire [2:0] w_n5793_27;
	wire [2:0] w_n5793_28;
	wire [2:0] w_n5793_29;
	wire [1:0] w_n5794_0;
	wire [1:0] w_n5795_0;
	wire [2:0] w_n5797_0;
	wire [1:0] w_n5797_1;
	wire [2:0] w_n5798_0;
	wire [2:0] w_n5802_0;
	wire [1:0] w_n5803_0;
	wire [1:0] w_n5805_0;
	wire [1:0] w_n5807_0;
	wire [1:0] w_n5810_0;
	wire [1:0] w_n5815_0;
	wire [1:0] w_n5817_0;
	wire [1:0] w_n5818_0;
	wire [2:0] w_n5819_0;
	wire [1:0] w_n5820_0;
	wire [1:0] w_n5824_0;
	wire [1:0] w_n5825_0;
	wire [1:0] w_n5827_0;
	wire [1:0] w_n5831_0;
	wire [1:0] w_n5833_0;
	wire [1:0] w_n5834_0;
	wire [2:0] w_n5835_0;
	wire [1:0] w_n5836_0;
	wire [1:0] w_n5840_0;
	wire [1:0] w_n5842_0;
	wire [1:0] w_n5844_0;
	wire [1:0] w_n5846_0;
	wire [1:0] w_n5849_0;
	wire [1:0] w_n5855_0;
	wire [2:0] w_n5857_0;
	wire [1:0] w_n5858_0;
	wire [1:0] w_n5863_0;
	wire [1:0] w_n5865_0;
	wire [1:0] w_n5867_0;
	wire [1:0] w_n5871_0;
	wire [1:0] w_n5873_0;
	wire [1:0] w_n5874_0;
	wire [2:0] w_n5875_0;
	wire [1:0] w_n5876_0;
	wire [1:0] w_n5882_0;
	wire [1:0] w_n5883_0;
	wire [1:0] w_n5885_0;
	wire [1:0] w_n5887_0;
	wire [1:0] w_n5889_0;
	wire [1:0] w_n5895_0;
	wire [1:0] w_n5897_0;
	wire [2:0] w_n5898_0;
	wire [1:0] w_n5901_0;
	wire [1:0] w_n5902_0;
	wire [2:0] w_n5903_0;
	wire [1:0] w_n5905_0;
	wire [1:0] w_n5909_0;
	wire [1:0] w_n5911_0;
	wire [1:0] w_n5912_0;
	wire [2:0] w_n5913_0;
	wire [1:0] w_n5914_0;
	wire [1:0] w_n5917_0;
	wire [1:0] w_n5923_0;
	wire [1:0] w_n5924_0;
	wire [1:0] w_n5926_0;
	wire [1:0] w_n5928_0;
	wire [1:0] w_n5930_0;
	wire [1:0] w_n5936_0;
	wire [1:0] w_n5938_0;
	wire [2:0] w_n5939_0;
	wire [1:0] w_n5942_0;
	wire [1:0] w_n5943_0;
	wire [2:0] w_n5944_0;
	wire [1:0] w_n5946_0;
	wire [1:0] w_n5950_0;
	wire [1:0] w_n5952_0;
	wire [1:0] w_n5953_0;
	wire [2:0] w_n5954_0;
	wire [1:0] w_n5955_0;
	wire [1:0] w_n5958_0;
	wire [1:0] w_n5964_0;
	wire [1:0] w_n5965_0;
	wire [1:0] w_n5967_0;
	wire [1:0] w_n5969_0;
	wire [1:0] w_n5971_0;
	wire [1:0] w_n5977_0;
	wire [1:0] w_n5979_0;
	wire [2:0] w_n5980_0;
	wire [1:0] w_n5983_0;
	wire [1:0] w_n5984_0;
	wire [2:0] w_n5985_0;
	wire [1:0] w_n5987_0;
	wire [1:0] w_n5991_0;
	wire [1:0] w_n5993_0;
	wire [1:0] w_n5994_0;
	wire [2:0] w_n5995_0;
	wire [1:0] w_n5996_0;
	wire [1:0] w_n5999_0;
	wire [1:0] w_n6005_0;
	wire [1:0] w_n6006_0;
	wire [1:0] w_n6008_0;
	wire [1:0] w_n6010_0;
	wire [1:0] w_n6012_0;
	wire [1:0] w_n6018_0;
	wire [1:0] w_n6020_0;
	wire [2:0] w_n6021_0;
	wire [1:0] w_n6024_0;
	wire [1:0] w_n6025_0;
	wire [2:0] w_n6026_0;
	wire [1:0] w_n6028_0;
	wire [1:0] w_n6032_0;
	wire [1:0] w_n6034_0;
	wire [1:0] w_n6035_0;
	wire [2:0] w_n6036_0;
	wire [1:0] w_n6037_0;
	wire [1:0] w_n6040_0;
	wire [1:0] w_n6046_0;
	wire [1:0] w_n6047_0;
	wire [1:0] w_n6049_0;
	wire [1:0] w_n6051_0;
	wire [1:0] w_n6053_0;
	wire [1:0] w_n6059_0;
	wire [1:0] w_n6061_0;
	wire [2:0] w_n6062_0;
	wire [1:0] w_n6065_0;
	wire [1:0] w_n6066_0;
	wire [2:0] w_n6067_0;
	wire [1:0] w_n6069_0;
	wire [1:0] w_n6073_0;
	wire [1:0] w_n6075_0;
	wire [1:0] w_n6076_0;
	wire [2:0] w_n6077_0;
	wire [1:0] w_n6078_0;
	wire [1:0] w_n6081_0;
	wire [1:0] w_n6087_0;
	wire [1:0] w_n6088_0;
	wire [1:0] w_n6090_0;
	wire [1:0] w_n6092_0;
	wire [1:0] w_n6094_0;
	wire [1:0] w_n6100_0;
	wire [2:0] w_n6102_0;
	wire [1:0] w_n6107_0;
	wire [2:0] w_n6109_0;
	wire [2:0] w_n6113_0;
	wire [1:0] w_n6114_0;
	wire [1:0] w_n6119_0;
	wire [2:0] w_n6120_0;
	wire [1:0] w_n6125_0;
	wire [1:0] w_n6132_0;
	wire [2:0] w_n6134_0;
	wire [1:0] w_n6134_1;
	wire [1:0] w_n6135_0;
	wire [2:0] w_n6138_0;
	wire [1:0] w_n6139_0;
	wire [1:0] w_n6140_0;
	wire [1:0] w_n6141_0;
	wire [1:0] w_n6143_0;
	wire [1:0] w_n6145_0;
	wire [1:0] w_n6154_0;
	wire [1:0] w_n6156_0;
	wire [1:0] w_n6157_0;
	wire [2:0] w_n6158_0;
	wire [1:0] w_n6159_0;
	wire [1:0] w_n6162_0;
	wire [1:0] w_n6164_0;
	wire [1:0] w_n6166_0;
	wire [1:0] w_n6169_0;
	wire [1:0] w_n6175_0;
	wire [2:0] w_n6177_0;
	wire [1:0] w_n6178_0;
	wire [1:0] w_n6183_0;
	wire [1:0] w_n6184_0;
	wire [1:0] w_n6186_0;
	wire [1:0] w_n6188_0;
	wire [1:0] w_n6191_0;
	wire [1:0] w_n6197_0;
	wire [2:0] w_n6199_0;
	wire [1:0] w_n6200_0;
	wire [1:0] w_n6204_0;
	wire [1:0] w_n6205_0;
	wire [1:0] w_n6207_0;
	wire [1:0] w_n6212_0;
	wire [1:0] w_n6214_0;
	wire [1:0] w_n6215_0;
	wire [2:0] w_n6216_0;
	wire [1:0] w_n6217_0;
	wire [1:0] w_n6221_0;
	wire [1:0] w_n6222_0;
	wire [1:0] w_n6224_0;
	wire [1:0] w_n6226_0;
	wire [1:0] w_n6229_0;
	wire [1:0] w_n6235_0;
	wire [1:0] w_n6237_0;
	wire [2:0] w_n6238_0;
	wire [1:0] w_n6242_0;
	wire [1:0] w_n6243_0;
	wire [2:0] w_n6244_0;
	wire [1:0] w_n6246_0;
	wire [1:0] w_n6251_0;
	wire [1:0] w_n6253_0;
	wire [1:0] w_n6254_0;
	wire [2:0] w_n6255_0;
	wire [1:0] w_n6256_0;
	wire [1:0] w_n6260_0;
	wire [1:0] w_n6266_0;
	wire [1:0] w_n6267_0;
	wire [1:0] w_n6269_0;
	wire [1:0] w_n6271_0;
	wire [1:0] w_n6274_0;
	wire [1:0] w_n6280_0;
	wire [1:0] w_n6282_0;
	wire [2:0] w_n6283_0;
	wire [1:0] w_n6287_0;
	wire [1:0] w_n6288_0;
	wire [2:0] w_n6289_0;
	wire [1:0] w_n6291_0;
	wire [1:0] w_n6296_0;
	wire [1:0] w_n6298_0;
	wire [1:0] w_n6299_0;
	wire [2:0] w_n6300_0;
	wire [1:0] w_n6301_0;
	wire [1:0] w_n6305_0;
	wire [1:0] w_n6311_0;
	wire [1:0] w_n6312_0;
	wire [1:0] w_n6314_0;
	wire [1:0] w_n6316_0;
	wire [1:0] w_n6319_0;
	wire [1:0] w_n6325_0;
	wire [1:0] w_n6327_0;
	wire [2:0] w_n6328_0;
	wire [1:0] w_n6332_0;
	wire [1:0] w_n6333_0;
	wire [2:0] w_n6334_0;
	wire [1:0] w_n6336_0;
	wire [1:0] w_n6341_0;
	wire [1:0] w_n6343_0;
	wire [1:0] w_n6344_0;
	wire [2:0] w_n6345_0;
	wire [1:0] w_n6346_0;
	wire [1:0] w_n6350_0;
	wire [1:0] w_n6356_0;
	wire [1:0] w_n6357_0;
	wire [1:0] w_n6359_0;
	wire [1:0] w_n6361_0;
	wire [1:0] w_n6364_0;
	wire [1:0] w_n6370_0;
	wire [1:0] w_n6372_0;
	wire [2:0] w_n6373_0;
	wire [1:0] w_n6377_0;
	wire [1:0] w_n6378_0;
	wire [2:0] w_n6379_0;
	wire [1:0] w_n6381_0;
	wire [1:0] w_n6386_0;
	wire [1:0] w_n6388_0;
	wire [1:0] w_n6389_0;
	wire [2:0] w_n6390_0;
	wire [1:0] w_n6391_0;
	wire [1:0] w_n6395_0;
	wire [1:0] w_n6401_0;
	wire [1:0] w_n6402_0;
	wire [1:0] w_n6404_0;
	wire [1:0] w_n6406_0;
	wire [1:0] w_n6409_0;
	wire [1:0] w_n6415_0;
	wire [1:0] w_n6417_0;
	wire [2:0] w_n6418_0;
	wire [1:0] w_n6422_0;
	wire [1:0] w_n6423_0;
	wire [2:0] w_n6424_0;
	wire [1:0] w_n6426_0;
	wire [1:0] w_n6431_0;
	wire [1:0] w_n6433_0;
	wire [1:0] w_n6434_0;
	wire [2:0] w_n6435_0;
	wire [1:0] w_n6436_0;
	wire [1:0] w_n6440_0;
	wire [1:0] w_n6446_0;
	wire [1:0] w_n6447_0;
	wire [1:0] w_n6449_0;
	wire [1:0] w_n6451_0;
	wire [1:0] w_n6454_0;
	wire [1:0] w_n6460_0;
	wire [1:0] w_n6462_0;
	wire [2:0] w_n6463_0;
	wire [1:0] w_n6467_0;
	wire [1:0] w_n6468_0;
	wire [2:0] w_n6469_0;
	wire [1:0] w_n6471_0;
	wire [1:0] w_n6476_0;
	wire [1:0] w_n6478_0;
	wire [1:0] w_n6479_0;
	wire [2:0] w_n6480_0;
	wire [2:0] w_n6480_1;
	wire [1:0] w_n6483_0;
	wire [2:0] w_n6484_0;
	wire [1:0] w_n6485_0;
	wire [1:0] w_n6486_0;
	wire [1:0] w_n6492_0;
	wire [2:0] w_n6493_0;
	wire [1:0] w_n6494_0;
	wire [1:0] w_n6499_0;
	wire [2:0] w_n6500_0;
	wire [2:0] w_n6500_1;
	wire [2:0] w_n6500_2;
	wire [2:0] w_n6500_3;
	wire [2:0] w_n6500_4;
	wire [2:0] w_n6500_5;
	wire [2:0] w_n6500_6;
	wire [2:0] w_n6500_7;
	wire [2:0] w_n6500_8;
	wire [2:0] w_n6500_9;
	wire [2:0] w_n6500_10;
	wire [2:0] w_n6500_11;
	wire [2:0] w_n6500_12;
	wire [2:0] w_n6500_13;
	wire [2:0] w_n6500_14;
	wire [2:0] w_n6500_15;
	wire [2:0] w_n6500_16;
	wire [2:0] w_n6500_17;
	wire [2:0] w_n6500_18;
	wire [1:0] w_n6500_19;
	wire [2:0] w_n6505_0;
	wire [2:0] w_n6505_1;
	wire [2:0] w_n6505_2;
	wire [2:0] w_n6505_3;
	wire [2:0] w_n6505_4;
	wire [2:0] w_n6505_5;
	wire [2:0] w_n6505_6;
	wire [2:0] w_n6505_7;
	wire [2:0] w_n6505_8;
	wire [2:0] w_n6505_9;
	wire [2:0] w_n6505_10;
	wire [2:0] w_n6505_11;
	wire [2:0] w_n6505_12;
	wire [2:0] w_n6505_13;
	wire [2:0] w_n6505_14;
	wire [2:0] w_n6505_15;
	wire [2:0] w_n6505_16;
	wire [2:0] w_n6505_17;
	wire [2:0] w_n6505_18;
	wire [2:0] w_n6505_19;
	wire [2:0] w_n6505_20;
	wire [2:0] w_n6505_21;
	wire [2:0] w_n6505_22;
	wire [2:0] w_n6505_23;
	wire [2:0] w_n6505_24;
	wire [2:0] w_n6505_25;
	wire [2:0] w_n6505_26;
	wire [2:0] w_n6505_27;
	wire [1:0] w_n6505_28;
	wire [1:0] w_n6508_0;
	wire [2:0] w_n6510_0;
	wire [1:0] w_n6510_1;
	wire [2:0] w_n6511_0;
	wire [2:0] w_n6515_0;
	wire [1:0] w_n6516_0;
	wire [1:0] w_n6517_0;
	wire [1:0] w_n6518_0;
	wire [1:0] w_n6520_0;
	wire [1:0] w_n6522_0;
	wire [1:0] w_n6524_0;
	wire [1:0] w_n6527_0;
	wire [1:0] w_n6532_0;
	wire [2:0] w_n6534_0;
	wire [1:0] w_n6535_0;
	wire [1:0] w_n6539_0;
	wire [1:0] w_n6540_0;
	wire [1:0] w_n6542_0;
	wire [1:0] w_n6544_0;
	wire [1:0] w_n6547_0;
	wire [1:0] w_n6553_0;
	wire [2:0] w_n6555_0;
	wire [1:0] w_n6556_0;
	wire [1:0] w_n6559_0;
	wire [1:0] w_n6561_0;
	wire [1:0] w_n6565_0;
	wire [1:0] w_n6567_0;
	wire [1:0] w_n6568_0;
	wire [2:0] w_n6569_0;
	wire [1:0] w_n6570_0;
	wire [1:0] w_n6575_0;
	wire [1:0] w_n6577_0;
	wire [1:0] w_n6579_0;
	wire [1:0] w_n6583_0;
	wire [1:0] w_n6585_0;
	wire [1:0] w_n6586_0;
	wire [2:0] w_n6587_0;
	wire [1:0] w_n6588_0;
	wire [1:0] w_n6594_0;
	wire [1:0] w_n6595_0;
	wire [1:0] w_n6597_0;
	wire [1:0] w_n6599_0;
	wire [1:0] w_n6601_0;
	wire [1:0] w_n6607_0;
	wire [1:0] w_n6609_0;
	wire [2:0] w_n6610_0;
	wire [1:0] w_n6613_0;
	wire [1:0] w_n6614_0;
	wire [2:0] w_n6615_0;
	wire [1:0] w_n6617_0;
	wire [1:0] w_n6621_0;
	wire [1:0] w_n6623_0;
	wire [1:0] w_n6624_0;
	wire [2:0] w_n6625_0;
	wire [1:0] w_n6626_0;
	wire [1:0] w_n6629_0;
	wire [1:0] w_n6635_0;
	wire [1:0] w_n6636_0;
	wire [1:0] w_n6638_0;
	wire [1:0] w_n6640_0;
	wire [1:0] w_n6642_0;
	wire [1:0] w_n6648_0;
	wire [1:0] w_n6650_0;
	wire [2:0] w_n6651_0;
	wire [1:0] w_n6654_0;
	wire [1:0] w_n6655_0;
	wire [2:0] w_n6656_0;
	wire [1:0] w_n6658_0;
	wire [1:0] w_n6662_0;
	wire [1:0] w_n6664_0;
	wire [1:0] w_n6665_0;
	wire [2:0] w_n6666_0;
	wire [1:0] w_n6667_0;
	wire [1:0] w_n6670_0;
	wire [1:0] w_n6676_0;
	wire [1:0] w_n6677_0;
	wire [1:0] w_n6679_0;
	wire [1:0] w_n6681_0;
	wire [1:0] w_n6683_0;
	wire [1:0] w_n6689_0;
	wire [1:0] w_n6691_0;
	wire [2:0] w_n6692_0;
	wire [1:0] w_n6695_0;
	wire [1:0] w_n6696_0;
	wire [2:0] w_n6697_0;
	wire [1:0] w_n6699_0;
	wire [1:0] w_n6703_0;
	wire [1:0] w_n6705_0;
	wire [1:0] w_n6706_0;
	wire [2:0] w_n6707_0;
	wire [1:0] w_n6708_0;
	wire [1:0] w_n6711_0;
	wire [1:0] w_n6717_0;
	wire [1:0] w_n6718_0;
	wire [1:0] w_n6720_0;
	wire [1:0] w_n6722_0;
	wire [1:0] w_n6724_0;
	wire [1:0] w_n6730_0;
	wire [1:0] w_n6732_0;
	wire [2:0] w_n6733_0;
	wire [1:0] w_n6736_0;
	wire [1:0] w_n6737_0;
	wire [2:0] w_n6738_0;
	wire [1:0] w_n6740_0;
	wire [1:0] w_n6744_0;
	wire [1:0] w_n6746_0;
	wire [1:0] w_n6747_0;
	wire [2:0] w_n6748_0;
	wire [1:0] w_n6749_0;
	wire [1:0] w_n6752_0;
	wire [1:0] w_n6758_0;
	wire [1:0] w_n6759_0;
	wire [1:0] w_n6761_0;
	wire [1:0] w_n6763_0;
	wire [1:0] w_n6765_0;
	wire [1:0] w_n6771_0;
	wire [1:0] w_n6773_0;
	wire [2:0] w_n6774_0;
	wire [1:0] w_n6777_0;
	wire [1:0] w_n6778_0;
	wire [2:0] w_n6779_0;
	wire [1:0] w_n6781_0;
	wire [1:0] w_n6785_0;
	wire [1:0] w_n6787_0;
	wire [1:0] w_n6788_0;
	wire [2:0] w_n6789_0;
	wire [1:0] w_n6790_0;
	wire [1:0] w_n6793_0;
	wire [1:0] w_n6799_0;
	wire [1:0] w_n6800_0;
	wire [1:0] w_n6802_0;
	wire [1:0] w_n6804_0;
	wire [1:0] w_n6806_0;
	wire [1:0] w_n6812_0;
	wire [1:0] w_n6814_0;
	wire [2:0] w_n6815_0;
	wire [1:0] w_n6818_0;
	wire [1:0] w_n6819_0;
	wire [2:0] w_n6820_0;
	wire [1:0] w_n6822_0;
	wire [1:0] w_n6826_0;
	wire [1:0] w_n6828_0;
	wire [1:0] w_n6829_0;
	wire [2:0] w_n6830_0;
	wire [1:0] w_n6834_0;
	wire [1:0] w_n6840_0;
	wire [2:0] w_n6842_0;
	wire [1:0] w_n6844_0;
	wire [2:0] w_n6849_0;
	wire [1:0] w_n6850_0;
	wire [1:0] w_n6851_0;
	wire [1:0] w_n6856_0;
	wire [2:0] w_n6857_0;
	wire [1:0] w_n6862_0;
	wire [1:0] w_n6869_0;
	wire [2:0] w_n6872_0;
	wire [1:0] w_n6872_1;
	wire [1:0] w_n6873_0;
	wire [2:0] w_n6876_0;
	wire [1:0] w_n6877_0;
	wire [1:0] w_n6878_0;
	wire [1:0] w_n6879_0;
	wire [1:0] w_n6881_0;
	wire [1:0] w_n6883_0;
	wire [1:0] w_n6885_0;
	wire [1:0] w_n6894_0;
	wire [2:0] w_n6896_0;
	wire [1:0] w_n6897_0;
	wire [1:0] w_n6901_0;
	wire [1:0] w_n6903_0;
	wire [1:0] w_n6905_0;
	wire [1:0] w_n6910_0;
	wire [1:0] w_n6912_0;
	wire [1:0] w_n6913_0;
	wire [2:0] w_n6914_0;
	wire [1:0] w_n6915_0;
	wire [1:0] w_n6920_0;
	wire [1:0] w_n6921_0;
	wire [1:0] w_n6923_0;
	wire [1:0] w_n6928_0;
	wire [1:0] w_n6930_0;
	wire [1:0] w_n6931_0;
	wire [2:0] w_n6932_0;
	wire [1:0] w_n6933_0;
	wire [1:0] w_n6935_0;
	wire [1:0] w_n6937_0;
	wire [1:0] w_n6939_0;
	wire [1:0] w_n6942_0;
	wire [1:0] w_n6948_0;
	wire [2:0] w_n6950_0;
	wire [1:0] w_n6951_0;
	wire [1:0] w_n6955_0;
	wire [1:0] w_n6956_0;
	wire [1:0] w_n6958_0;
	wire [1:0] w_n6960_0;
	wire [1:0] w_n6963_0;
	wire [1:0] w_n6969_0;
	wire [1:0] w_n6971_0;
	wire [2:0] w_n6972_0;
	wire [1:0] w_n6976_0;
	wire [1:0] w_n6977_0;
	wire [2:0] w_n6978_0;
	wire [1:0] w_n6980_0;
	wire [1:0] w_n6985_0;
	wire [1:0] w_n6987_0;
	wire [1:0] w_n6988_0;
	wire [2:0] w_n6989_0;
	wire [1:0] w_n6990_0;
	wire [1:0] w_n6994_0;
	wire [1:0] w_n7000_0;
	wire [1:0] w_n7001_0;
	wire [1:0] w_n7003_0;
	wire [1:0] w_n7005_0;
	wire [1:0] w_n7008_0;
	wire [1:0] w_n7014_0;
	wire [1:0] w_n7016_0;
	wire [2:0] w_n7017_0;
	wire [1:0] w_n7021_0;
	wire [1:0] w_n7022_0;
	wire [2:0] w_n7023_0;
	wire [1:0] w_n7025_0;
	wire [1:0] w_n7030_0;
	wire [1:0] w_n7032_0;
	wire [1:0] w_n7033_0;
	wire [2:0] w_n7034_0;
	wire [1:0] w_n7035_0;
	wire [1:0] w_n7039_0;
	wire [1:0] w_n7045_0;
	wire [1:0] w_n7046_0;
	wire [1:0] w_n7048_0;
	wire [1:0] w_n7050_0;
	wire [1:0] w_n7053_0;
	wire [1:0] w_n7059_0;
	wire [1:0] w_n7061_0;
	wire [2:0] w_n7062_0;
	wire [1:0] w_n7066_0;
	wire [1:0] w_n7067_0;
	wire [2:0] w_n7068_0;
	wire [1:0] w_n7070_0;
	wire [1:0] w_n7075_0;
	wire [1:0] w_n7077_0;
	wire [1:0] w_n7078_0;
	wire [2:0] w_n7079_0;
	wire [1:0] w_n7080_0;
	wire [1:0] w_n7084_0;
	wire [1:0] w_n7090_0;
	wire [1:0] w_n7091_0;
	wire [1:0] w_n7093_0;
	wire [1:0] w_n7095_0;
	wire [1:0] w_n7098_0;
	wire [1:0] w_n7104_0;
	wire [1:0] w_n7106_0;
	wire [2:0] w_n7107_0;
	wire [1:0] w_n7111_0;
	wire [1:0] w_n7112_0;
	wire [2:0] w_n7113_0;
	wire [1:0] w_n7115_0;
	wire [1:0] w_n7120_0;
	wire [1:0] w_n7122_0;
	wire [1:0] w_n7123_0;
	wire [2:0] w_n7124_0;
	wire [1:0] w_n7125_0;
	wire [1:0] w_n7129_0;
	wire [1:0] w_n7135_0;
	wire [1:0] w_n7136_0;
	wire [1:0] w_n7138_0;
	wire [1:0] w_n7140_0;
	wire [1:0] w_n7143_0;
	wire [1:0] w_n7149_0;
	wire [1:0] w_n7151_0;
	wire [2:0] w_n7152_0;
	wire [1:0] w_n7156_0;
	wire [1:0] w_n7157_0;
	wire [2:0] w_n7158_0;
	wire [1:0] w_n7160_0;
	wire [1:0] w_n7165_0;
	wire [1:0] w_n7167_0;
	wire [1:0] w_n7168_0;
	wire [2:0] w_n7169_0;
	wire [1:0] w_n7170_0;
	wire [1:0] w_n7174_0;
	wire [1:0] w_n7180_0;
	wire [1:0] w_n7181_0;
	wire [1:0] w_n7183_0;
	wire [1:0] w_n7185_0;
	wire [1:0] w_n7188_0;
	wire [1:0] w_n7194_0;
	wire [1:0] w_n7196_0;
	wire [2:0] w_n7197_0;
	wire [1:0] w_n7201_0;
	wire [1:0] w_n7202_0;
	wire [2:0] w_n7203_0;
	wire [1:0] w_n7205_0;
	wire [1:0] w_n7210_0;
	wire [1:0] w_n7212_0;
	wire [1:0] w_n7213_0;
	wire [2:0] w_n7214_0;
	wire [1:0] w_n7215_0;
	wire [1:0] w_n7219_0;
	wire [1:0] w_n7225_0;
	wire [1:0] w_n7226_0;
	wire [1:0] w_n7228_0;
	wire [1:0] w_n7230_0;
	wire [1:0] w_n7233_0;
	wire [1:0] w_n7239_0;
	wire [2:0] w_n7241_0;
	wire [2:0] w_n7241_1;
	wire [1:0] w_n7244_0;
	wire [2:0] w_n7245_0;
	wire [1:0] w_n7246_0;
	wire [1:0] w_n7252_0;
	wire [2:0] w_n7253_0;
	wire [1:0] w_n7254_0;
	wire [1:0] w_n7259_0;
	wire [2:0] w_n7260_0;
	wire [2:0] w_n7260_1;
	wire [2:0] w_n7260_2;
	wire [2:0] w_n7260_3;
	wire [2:0] w_n7260_4;
	wire [2:0] w_n7260_5;
	wire [2:0] w_n7260_6;
	wire [2:0] w_n7260_7;
	wire [2:0] w_n7260_8;
	wire [2:0] w_n7260_9;
	wire [2:0] w_n7260_10;
	wire [2:0] w_n7260_11;
	wire [2:0] w_n7260_12;
	wire [2:0] w_n7260_13;
	wire [2:0] w_n7260_14;
	wire [2:0] w_n7260_15;
	wire [2:0] w_n7260_16;
	wire [2:0] w_n7260_17;
	wire [1:0] w_n7260_18;
	wire [2:0] w_n7265_0;
	wire [2:0] w_n7265_1;
	wire [2:0] w_n7265_2;
	wire [2:0] w_n7265_3;
	wire [2:0] w_n7265_4;
	wire [2:0] w_n7265_5;
	wire [2:0] w_n7265_6;
	wire [2:0] w_n7265_7;
	wire [2:0] w_n7265_8;
	wire [2:0] w_n7265_9;
	wire [2:0] w_n7265_10;
	wire [2:0] w_n7265_11;
	wire [2:0] w_n7265_12;
	wire [2:0] w_n7265_13;
	wire [2:0] w_n7265_14;
	wire [2:0] w_n7265_15;
	wire [2:0] w_n7265_16;
	wire [2:0] w_n7265_17;
	wire [2:0] w_n7265_18;
	wire [2:0] w_n7265_19;
	wire [2:0] w_n7265_20;
	wire [2:0] w_n7265_21;
	wire [2:0] w_n7265_22;
	wire [2:0] w_n7265_23;
	wire [2:0] w_n7265_24;
	wire [2:0] w_n7265_25;
	wire [2:0] w_n7265_26;
	wire [2:0] w_n7265_27;
	wire [1:0] w_n7265_28;
	wire [1:0] w_n7269_0;
	wire [2:0] w_n7271_0;
	wire [1:0] w_n7271_1;
	wire [2:0] w_n7272_0;
	wire [2:0] w_n7276_0;
	wire [1:0] w_n7277_0;
	wire [1:0] w_n7278_0;
	wire [1:0] w_n7279_0;
	wire [1:0] w_n7281_0;
	wire [1:0] w_n7283_0;
	wire [1:0] w_n7285_0;
	wire [1:0] w_n7288_0;
	wire [1:0] w_n7293_0;
	wire [2:0] w_n7295_0;
	wire [1:0] w_n7296_0;
	wire [1:0] w_n7300_0;
	wire [1:0] w_n7301_0;
	wire [1:0] w_n7303_0;
	wire [1:0] w_n7307_0;
	wire [1:0] w_n7309_0;
	wire [1:0] w_n7310_0;
	wire [2:0] w_n7311_0;
	wire [1:0] w_n7312_0;
	wire [1:0] w_n7316_0;
	wire [1:0] w_n7318_0;
	wire [1:0] w_n7320_0;
	wire [1:0] w_n7322_0;
	wire [1:0] w_n7325_0;
	wire [1:0] w_n7331_0;
	wire [2:0] w_n7333_0;
	wire [1:0] w_n7334_0;
	wire [1:0] w_n7339_0;
	wire [1:0] w_n7341_0;
	wire [1:0] w_n7343_0;
	wire [1:0] w_n7345_0;
	wire [1:0] w_n7347_0;
	wire [1:0] w_n7353_0;
	wire [2:0] w_n7355_0;
	wire [1:0] w_n7356_0;
	wire [1:0] w_n7358_0;
	wire [1:0] w_n7360_0;
	wire [1:0] w_n7364_0;
	wire [1:0] w_n7366_0;
	wire [1:0] w_n7367_0;
	wire [1:0] w_n7368_0;
	wire [2:0] w_n7369_0;
	wire [1:0] w_n7372_0;
	wire [1:0] w_n7373_0;
	wire [2:0] w_n7374_0;
	wire [1:0] w_n7376_0;
	wire [1:0] w_n7380_0;
	wire [1:0] w_n7382_0;
	wire [1:0] w_n7383_0;
	wire [2:0] w_n7384_0;
	wire [1:0] w_n7385_0;
	wire [1:0] w_n7388_0;
	wire [1:0] w_n7394_0;
	wire [1:0] w_n7395_0;
	wire [1:0] w_n7397_0;
	wire [1:0] w_n7399_0;
	wire [1:0] w_n7401_0;
	wire [1:0] w_n7407_0;
	wire [1:0] w_n7409_0;
	wire [2:0] w_n7410_0;
	wire [1:0] w_n7413_0;
	wire [1:0] w_n7414_0;
	wire [2:0] w_n7415_0;
	wire [1:0] w_n7417_0;
	wire [1:0] w_n7421_0;
	wire [1:0] w_n7423_0;
	wire [1:0] w_n7424_0;
	wire [2:0] w_n7425_0;
	wire [1:0] w_n7426_0;
	wire [1:0] w_n7429_0;
	wire [1:0] w_n7435_0;
	wire [1:0] w_n7436_0;
	wire [1:0] w_n7438_0;
	wire [1:0] w_n7440_0;
	wire [1:0] w_n7442_0;
	wire [1:0] w_n7448_0;
	wire [1:0] w_n7450_0;
	wire [2:0] w_n7451_0;
	wire [1:0] w_n7454_0;
	wire [1:0] w_n7455_0;
	wire [2:0] w_n7456_0;
	wire [1:0] w_n7458_0;
	wire [1:0] w_n7462_0;
	wire [1:0] w_n7464_0;
	wire [1:0] w_n7465_0;
	wire [2:0] w_n7466_0;
	wire [1:0] w_n7467_0;
	wire [1:0] w_n7470_0;
	wire [1:0] w_n7476_0;
	wire [1:0] w_n7477_0;
	wire [1:0] w_n7479_0;
	wire [1:0] w_n7481_0;
	wire [1:0] w_n7483_0;
	wire [1:0] w_n7489_0;
	wire [1:0] w_n7491_0;
	wire [2:0] w_n7492_0;
	wire [1:0] w_n7495_0;
	wire [1:0] w_n7496_0;
	wire [2:0] w_n7497_0;
	wire [1:0] w_n7499_0;
	wire [1:0] w_n7503_0;
	wire [1:0] w_n7505_0;
	wire [1:0] w_n7506_0;
	wire [2:0] w_n7507_0;
	wire [1:0] w_n7508_0;
	wire [1:0] w_n7511_0;
	wire [1:0] w_n7517_0;
	wire [1:0] w_n7518_0;
	wire [1:0] w_n7520_0;
	wire [1:0] w_n7522_0;
	wire [1:0] w_n7524_0;
	wire [1:0] w_n7530_0;
	wire [1:0] w_n7532_0;
	wire [2:0] w_n7533_0;
	wire [1:0] w_n7536_0;
	wire [1:0] w_n7537_0;
	wire [2:0] w_n7538_0;
	wire [1:0] w_n7540_0;
	wire [1:0] w_n7544_0;
	wire [1:0] w_n7546_0;
	wire [1:0] w_n7547_0;
	wire [2:0] w_n7548_0;
	wire [1:0] w_n7549_0;
	wire [1:0] w_n7552_0;
	wire [1:0] w_n7558_0;
	wire [1:0] w_n7559_0;
	wire [1:0] w_n7561_0;
	wire [1:0] w_n7563_0;
	wire [1:0] w_n7565_0;
	wire [1:0] w_n7571_0;
	wire [1:0] w_n7573_0;
	wire [2:0] w_n7574_0;
	wire [1:0] w_n7577_0;
	wire [1:0] w_n7578_0;
	wire [2:0] w_n7579_0;
	wire [1:0] w_n7581_0;
	wire [1:0] w_n7585_0;
	wire [1:0] w_n7587_0;
	wire [1:0] w_n7588_0;
	wire [2:0] w_n7589_0;
	wire [1:0] w_n7590_0;
	wire [1:0] w_n7593_0;
	wire [1:0] w_n7599_0;
	wire [1:0] w_n7600_0;
	wire [1:0] w_n7602_0;
	wire [1:0] w_n7604_0;
	wire [1:0] w_n7606_0;
	wire [1:0] w_n7612_0;
	wire [2:0] w_n7614_0;
	wire [1:0] w_n7619_0;
	wire [2:0] w_n7621_0;
	wire [2:0] w_n7625_0;
	wire [1:0] w_n7626_0;
	wire [1:0] w_n7631_0;
	wire [2:0] w_n7632_0;
	wire [1:0] w_n7637_0;
	wire [1:0] w_n7645_0;
	wire [2:0] w_n7647_0;
	wire [1:0] w_n7647_1;
	wire [1:0] w_n7648_0;
	wire [2:0] w_n7651_0;
	wire [1:0] w_n7652_0;
	wire [1:0] w_n7653_0;
	wire [1:0] w_n7654_0;
	wire [1:0] w_n7656_0;
	wire [1:0] w_n7658_0;
	wire [1:0] w_n7660_0;
	wire [1:0] w_n7669_0;
	wire [2:0] w_n7671_0;
	wire [1:0] w_n7672_0;
	wire [1:0] w_n7676_0;
	wire [1:0] w_n7678_0;
	wire [1:0] w_n7680_0;
	wire [1:0] w_n7685_0;
	wire [1:0] w_n7687_0;
	wire [1:0] w_n7688_0;
	wire [2:0] w_n7689_0;
	wire [1:0] w_n7690_0;
	wire [1:0] w_n7695_0;
	wire [1:0] w_n7696_0;
	wire [1:0] w_n7698_0;
	wire [1:0] w_n7700_0;
	wire [1:0] w_n7703_0;
	wire [1:0] w_n7709_0;
	wire [2:0] w_n7711_0;
	wire [1:0] w_n7712_0;
	wire [1:0] w_n7716_0;
	wire [1:0] w_n7717_0;
	wire [1:0] w_n7719_0;
	wire [1:0] w_n7724_0;
	wire [1:0] w_n7726_0;
	wire [1:0] w_n7727_0;
	wire [2:0] w_n7728_0;
	wire [1:0] w_n7729_0;
	wire [1:0] w_n7733_0;
	wire [1:0] w_n7734_0;
	wire [1:0] w_n7736_0;
	wire [1:0] w_n7741_0;
	wire [1:0] w_n7743_0;
	wire [1:0] w_n7744_0;
	wire [2:0] w_n7745_0;
	wire [1:0] w_n7746_0;
	wire [1:0] w_n7748_0;
	wire [1:0] w_n7750_0;
	wire [1:0] w_n7752_0;
	wire [1:0] w_n7755_0;
	wire [1:0] w_n7761_0;
	wire [2:0] w_n7763_0;
	wire [1:0] w_n7764_0;
	wire [1:0] w_n7768_0;
	wire [1:0] w_n7774_0;
	wire [1:0] w_n7775_0;
	wire [1:0] w_n7777_0;
	wire [1:0] w_n7779_0;
	wire [1:0] w_n7782_0;
	wire [1:0] w_n7788_0;
	wire [1:0] w_n7790_0;
	wire [2:0] w_n7791_0;
	wire [1:0] w_n7795_0;
	wire [1:0] w_n7796_0;
	wire [2:0] w_n7797_0;
	wire [1:0] w_n7799_0;
	wire [1:0] w_n7804_0;
	wire [1:0] w_n7806_0;
	wire [1:0] w_n7807_0;
	wire [2:0] w_n7808_0;
	wire [1:0] w_n7809_0;
	wire [1:0] w_n7813_0;
	wire [1:0] w_n7819_0;
	wire [1:0] w_n7820_0;
	wire [1:0] w_n7822_0;
	wire [1:0] w_n7824_0;
	wire [1:0] w_n7827_0;
	wire [1:0] w_n7833_0;
	wire [1:0] w_n7835_0;
	wire [2:0] w_n7836_0;
	wire [1:0] w_n7840_0;
	wire [1:0] w_n7841_0;
	wire [2:0] w_n7842_0;
	wire [1:0] w_n7844_0;
	wire [1:0] w_n7849_0;
	wire [1:0] w_n7851_0;
	wire [1:0] w_n7852_0;
	wire [2:0] w_n7853_0;
	wire [1:0] w_n7854_0;
	wire [1:0] w_n7858_0;
	wire [1:0] w_n7864_0;
	wire [1:0] w_n7865_0;
	wire [1:0] w_n7867_0;
	wire [1:0] w_n7869_0;
	wire [1:0] w_n7872_0;
	wire [1:0] w_n7878_0;
	wire [1:0] w_n7880_0;
	wire [2:0] w_n7881_0;
	wire [1:0] w_n7885_0;
	wire [1:0] w_n7886_0;
	wire [2:0] w_n7887_0;
	wire [1:0] w_n7889_0;
	wire [1:0] w_n7894_0;
	wire [1:0] w_n7896_0;
	wire [1:0] w_n7897_0;
	wire [2:0] w_n7898_0;
	wire [1:0] w_n7899_0;
	wire [1:0] w_n7903_0;
	wire [1:0] w_n7909_0;
	wire [1:0] w_n7910_0;
	wire [1:0] w_n7912_0;
	wire [1:0] w_n7914_0;
	wire [1:0] w_n7917_0;
	wire [1:0] w_n7923_0;
	wire [1:0] w_n7925_0;
	wire [2:0] w_n7926_0;
	wire [1:0] w_n7930_0;
	wire [1:0] w_n7931_0;
	wire [2:0] w_n7932_0;
	wire [1:0] w_n7934_0;
	wire [1:0] w_n7939_0;
	wire [1:0] w_n7941_0;
	wire [1:0] w_n7942_0;
	wire [2:0] w_n7943_0;
	wire [1:0] w_n7944_0;
	wire [1:0] w_n7948_0;
	wire [1:0] w_n7954_0;
	wire [1:0] w_n7955_0;
	wire [1:0] w_n7957_0;
	wire [1:0] w_n7959_0;
	wire [1:0] w_n7962_0;
	wire [1:0] w_n7968_0;
	wire [1:0] w_n7970_0;
	wire [2:0] w_n7971_0;
	wire [1:0] w_n7975_0;
	wire [1:0] w_n7976_0;
	wire [2:0] w_n7977_0;
	wire [1:0] w_n7979_0;
	wire [1:0] w_n7984_0;
	wire [1:0] w_n7986_0;
	wire [1:0] w_n7987_0;
	wire [2:0] w_n7988_0;
	wire [1:0] w_n7989_0;
	wire [1:0] w_n7993_0;
	wire [1:0] w_n7999_0;
	wire [1:0] w_n8000_0;
	wire [1:0] w_n8002_0;
	wire [1:0] w_n8004_0;
	wire [1:0] w_n8007_0;
	wire [1:0] w_n8013_0;
	wire [1:0] w_n8015_0;
	wire [2:0] w_n8016_0;
	wire [1:0] w_n8020_0;
	wire [1:0] w_n8021_0;
	wire [2:0] w_n8022_0;
	wire [1:0] w_n8024_0;
	wire [1:0] w_n8029_0;
	wire [1:0] w_n8031_0;
	wire [1:0] w_n8032_0;
	wire [2:0] w_n8033_0;
	wire [2:0] w_n8033_1;
	wire [1:0] w_n8036_0;
	wire [2:0] w_n8037_0;
	wire [1:0] w_n8038_0;
	wire [1:0] w_n8039_0;
	wire [1:0] w_n8045_0;
	wire [2:0] w_n8046_0;
	wire [1:0] w_n8047_0;
	wire [1:0] w_n8052_0;
	wire [2:0] w_n8053_0;
	wire [2:0] w_n8053_1;
	wire [2:0] w_n8053_2;
	wire [2:0] w_n8053_3;
	wire [2:0] w_n8053_4;
	wire [2:0] w_n8053_5;
	wire [2:0] w_n8053_6;
	wire [2:0] w_n8053_7;
	wire [2:0] w_n8053_8;
	wire [2:0] w_n8053_9;
	wire [2:0] w_n8053_10;
	wire [2:0] w_n8053_11;
	wire [2:0] w_n8053_12;
	wire [2:0] w_n8053_13;
	wire [2:0] w_n8053_14;
	wire [2:0] w_n8053_15;
	wire [2:0] w_n8053_16;
	wire [2:0] w_n8058_0;
	wire [2:0] w_n8058_1;
	wire [2:0] w_n8058_2;
	wire [2:0] w_n8058_3;
	wire [2:0] w_n8058_4;
	wire [2:0] w_n8058_5;
	wire [2:0] w_n8058_6;
	wire [2:0] w_n8058_7;
	wire [2:0] w_n8058_8;
	wire [2:0] w_n8058_9;
	wire [2:0] w_n8058_10;
	wire [2:0] w_n8058_11;
	wire [2:0] w_n8058_12;
	wire [2:0] w_n8058_13;
	wire [2:0] w_n8058_14;
	wire [2:0] w_n8058_15;
	wire [2:0] w_n8058_16;
	wire [2:0] w_n8058_17;
	wire [2:0] w_n8058_18;
	wire [2:0] w_n8058_19;
	wire [2:0] w_n8058_20;
	wire [2:0] w_n8058_21;
	wire [2:0] w_n8058_22;
	wire [2:0] w_n8058_23;
	wire [2:0] w_n8058_24;
	wire [2:0] w_n8058_25;
	wire [2:0] w_n8058_26;
	wire [1:0] w_n8058_27;
	wire [1:0] w_n8061_0;
	wire [2:0] w_n8063_0;
	wire [1:0] w_n8063_1;
	wire [2:0] w_n8064_0;
	wire [2:0] w_n8068_0;
	wire [1:0] w_n8069_0;
	wire [1:0] w_n8070_0;
	wire [1:0] w_n8071_0;
	wire [1:0] w_n8073_0;
	wire [1:0] w_n8075_0;
	wire [1:0] w_n8077_0;
	wire [1:0] w_n8080_0;
	wire [1:0] w_n8085_0;
	wire [2:0] w_n8087_0;
	wire [1:0] w_n8088_0;
	wire [1:0] w_n8092_0;
	wire [1:0] w_n8093_0;
	wire [1:0] w_n8095_0;
	wire [1:0] w_n8099_0;
	wire [1:0] w_n8101_0;
	wire [1:0] w_n8102_0;
	wire [2:0] w_n8103_0;
	wire [1:0] w_n8104_0;
	wire [1:0] w_n8108_0;
	wire [1:0] w_n8110_0;
	wire [1:0] w_n8112_0;
	wire [1:0] w_n8114_0;
	wire [1:0] w_n8117_0;
	wire [1:0] w_n8123_0;
	wire [2:0] w_n8125_0;
	wire [1:0] w_n8126_0;
	wire [1:0] w_n8131_0;
	wire [1:0] w_n8133_0;
	wire [1:0] w_n8135_0;
	wire [1:0] w_n8139_0;
	wire [1:0] w_n8141_0;
	wire [1:0] w_n8142_0;
	wire [2:0] w_n8143_0;
	wire [1:0] w_n8144_0;
	wire [1:0] w_n8150_0;
	wire [1:0] w_n8151_0;
	wire [1:0] w_n8153_0;
	wire [1:0] w_n8155_0;
	wire [1:0] w_n8157_0;
	wire [1:0] w_n8163_0;
	wire [1:0] w_n8165_0;
	wire [2:0] w_n8166_0;
	wire [1:0] w_n8169_0;
	wire [1:0] w_n8170_0;
	wire [2:0] w_n8171_0;
	wire [1:0] w_n8173_0;
	wire [1:0] w_n8175_0;
	wire [1:0] w_n8177_0;
	wire [1:0] w_n8183_0;
	wire [2:0] w_n8185_0;
	wire [1:0] w_n8186_0;
	wire [1:0] w_n8188_0;
	wire [1:0] w_n8190_0;
	wire [1:0] w_n8194_0;
	wire [1:0] w_n8196_0;
	wire [1:0] w_n8197_0;
	wire [1:0] w_n8198_0;
	wire [2:0] w_n8199_0;
	wire [1:0] w_n8202_0;
	wire [1:0] w_n8203_0;
	wire [2:0] w_n8204_0;
	wire [1:0] w_n8206_0;
	wire [1:0] w_n8210_0;
	wire [1:0] w_n8212_0;
	wire [1:0] w_n8213_0;
	wire [2:0] w_n8214_0;
	wire [1:0] w_n8215_0;
	wire [1:0] w_n8218_0;
	wire [1:0] w_n8224_0;
	wire [1:0] w_n8225_0;
	wire [1:0] w_n8227_0;
	wire [1:0] w_n8229_0;
	wire [1:0] w_n8231_0;
	wire [1:0] w_n8237_0;
	wire [1:0] w_n8239_0;
	wire [2:0] w_n8240_0;
	wire [1:0] w_n8243_0;
	wire [1:0] w_n8244_0;
	wire [2:0] w_n8245_0;
	wire [1:0] w_n8247_0;
	wire [1:0] w_n8251_0;
	wire [1:0] w_n8253_0;
	wire [1:0] w_n8254_0;
	wire [2:0] w_n8255_0;
	wire [1:0] w_n8256_0;
	wire [1:0] w_n8259_0;
	wire [1:0] w_n8265_0;
	wire [1:0] w_n8266_0;
	wire [1:0] w_n8268_0;
	wire [1:0] w_n8270_0;
	wire [1:0] w_n8272_0;
	wire [1:0] w_n8278_0;
	wire [1:0] w_n8280_0;
	wire [2:0] w_n8281_0;
	wire [1:0] w_n8284_0;
	wire [1:0] w_n8285_0;
	wire [2:0] w_n8286_0;
	wire [1:0] w_n8288_0;
	wire [1:0] w_n8292_0;
	wire [1:0] w_n8294_0;
	wire [1:0] w_n8295_0;
	wire [2:0] w_n8296_0;
	wire [1:0] w_n8297_0;
	wire [1:0] w_n8300_0;
	wire [1:0] w_n8306_0;
	wire [1:0] w_n8307_0;
	wire [1:0] w_n8309_0;
	wire [1:0] w_n8311_0;
	wire [1:0] w_n8313_0;
	wire [1:0] w_n8319_0;
	wire [1:0] w_n8321_0;
	wire [2:0] w_n8322_0;
	wire [1:0] w_n8325_0;
	wire [1:0] w_n8326_0;
	wire [2:0] w_n8327_0;
	wire [1:0] w_n8329_0;
	wire [1:0] w_n8333_0;
	wire [1:0] w_n8335_0;
	wire [1:0] w_n8336_0;
	wire [2:0] w_n8337_0;
	wire [1:0] w_n8338_0;
	wire [1:0] w_n8341_0;
	wire [1:0] w_n8347_0;
	wire [1:0] w_n8348_0;
	wire [1:0] w_n8350_0;
	wire [1:0] w_n8352_0;
	wire [1:0] w_n8354_0;
	wire [1:0] w_n8360_0;
	wire [1:0] w_n8362_0;
	wire [2:0] w_n8363_0;
	wire [1:0] w_n8366_0;
	wire [1:0] w_n8367_0;
	wire [2:0] w_n8368_0;
	wire [1:0] w_n8370_0;
	wire [1:0] w_n8374_0;
	wire [1:0] w_n8376_0;
	wire [1:0] w_n8377_0;
	wire [2:0] w_n8378_0;
	wire [1:0] w_n8379_0;
	wire [1:0] w_n8382_0;
	wire [1:0] w_n8388_0;
	wire [1:0] w_n8389_0;
	wire [1:0] w_n8391_0;
	wire [1:0] w_n8393_0;
	wire [1:0] w_n8395_0;
	wire [1:0] w_n8401_0;
	wire [1:0] w_n8403_0;
	wire [2:0] w_n8404_0;
	wire [1:0] w_n8407_0;
	wire [1:0] w_n8408_0;
	wire [2:0] w_n8409_0;
	wire [1:0] w_n8411_0;
	wire [1:0] w_n8415_0;
	wire [1:0] w_n8417_0;
	wire [1:0] w_n8418_0;
	wire [2:0] w_n8419_0;
	wire [1:0] w_n8423_0;
	wire [1:0] w_n8429_0;
	wire [2:0] w_n8431_0;
	wire [1:0] w_n8433_0;
	wire [2:0] w_n8438_0;
	wire [1:0] w_n8439_0;
	wire [1:0] w_n8440_0;
	wire [1:0] w_n8445_0;
	wire [2:0] w_n8446_0;
	wire [1:0] w_n8451_0;
	wire [1:0] w_n8458_0;
	wire [2:0] w_n8460_0;
	wire [1:0] w_n8460_1;
	wire [1:0] w_n8461_0;
	wire [2:0] w_n8464_0;
	wire [1:0] w_n8465_0;
	wire [1:0] w_n8466_0;
	wire [1:0] w_n8467_0;
	wire [1:0] w_n8469_0;
	wire [1:0] w_n8471_0;
	wire [1:0] w_n8473_0;
	wire [1:0] w_n8482_0;
	wire [2:0] w_n8484_0;
	wire [1:0] w_n8485_0;
	wire [1:0] w_n8489_0;
	wire [1:0] w_n8491_0;
	wire [1:0] w_n8493_0;
	wire [1:0] w_n8498_0;
	wire [1:0] w_n8500_0;
	wire [1:0] w_n8501_0;
	wire [2:0] w_n8502_0;
	wire [1:0] w_n8503_0;
	wire [1:0] w_n8508_0;
	wire [1:0] w_n8509_0;
	wire [1:0] w_n8511_0;
	wire [1:0] w_n8513_0;
	wire [1:0] w_n8516_0;
	wire [1:0] w_n8522_0;
	wire [2:0] w_n8524_0;
	wire [1:0] w_n8525_0;
	wire [1:0] w_n8529_0;
	wire [1:0] w_n8530_0;
	wire [1:0] w_n8532_0;
	wire [1:0] w_n8537_0;
	wire [1:0] w_n8539_0;
	wire [1:0] w_n8540_0;
	wire [2:0] w_n8541_0;
	wire [1:0] w_n8542_0;
	wire [1:0] w_n8546_0;
	wire [1:0] w_n8547_0;
	wire [1:0] w_n8549_0;
	wire [1:0] w_n8551_0;
	wire [1:0] w_n8554_0;
	wire [1:0] w_n8560_0;
	wire [1:0] w_n8562_0;
	wire [2:0] w_n8563_0;
	wire [1:0] w_n8567_0;
	wire [1:0] w_n8568_0;
	wire [2:0] w_n8569_0;
	wire [1:0] w_n8571_0;
	wire [1:0] w_n8576_0;
	wire [1:0] w_n8578_0;
	wire [1:0] w_n8579_0;
	wire [2:0] w_n8580_0;
	wire [1:0] w_n8581_0;
	wire [1:0] w_n8585_0;
	wire [1:0] w_n8591_0;
	wire [1:0] w_n8592_0;
	wire [1:0] w_n8594_0;
	wire [1:0] w_n8599_0;
	wire [1:0] w_n8601_0;
	wire [1:0] w_n8602_0;
	wire [2:0] w_n8603_0;
	wire [1:0] w_n8604_0;
	wire [1:0] w_n8607_0;
	wire [1:0] w_n8609_0;
	wire [1:0] w_n8611_0;
	wire [1:0] w_n8614_0;
	wire [1:0] w_n8620_0;
	wire [2:0] w_n8622_0;
	wire [1:0] w_n8623_0;
	wire [1:0] w_n8627_0;
	wire [1:0] w_n8633_0;
	wire [1:0] w_n8634_0;
	wire [1:0] w_n8636_0;
	wire [1:0] w_n8638_0;
	wire [1:0] w_n8641_0;
	wire [1:0] w_n8647_0;
	wire [1:0] w_n8649_0;
	wire [2:0] w_n8650_0;
	wire [1:0] w_n8654_0;
	wire [1:0] w_n8655_0;
	wire [2:0] w_n8656_0;
	wire [1:0] w_n8658_0;
	wire [1:0] w_n8663_0;
	wire [1:0] w_n8665_0;
	wire [1:0] w_n8666_0;
	wire [2:0] w_n8667_0;
	wire [1:0] w_n8668_0;
	wire [1:0] w_n8672_0;
	wire [1:0] w_n8678_0;
	wire [1:0] w_n8679_0;
	wire [1:0] w_n8681_0;
	wire [1:0] w_n8683_0;
	wire [1:0] w_n8686_0;
	wire [1:0] w_n8692_0;
	wire [1:0] w_n8694_0;
	wire [2:0] w_n8695_0;
	wire [1:0] w_n8699_0;
	wire [1:0] w_n8700_0;
	wire [2:0] w_n8701_0;
	wire [1:0] w_n8703_0;
	wire [1:0] w_n8708_0;
	wire [1:0] w_n8710_0;
	wire [1:0] w_n8711_0;
	wire [2:0] w_n8712_0;
	wire [1:0] w_n8713_0;
	wire [1:0] w_n8717_0;
	wire [1:0] w_n8723_0;
	wire [1:0] w_n8724_0;
	wire [1:0] w_n8726_0;
	wire [1:0] w_n8728_0;
	wire [1:0] w_n8731_0;
	wire [1:0] w_n8737_0;
	wire [1:0] w_n8739_0;
	wire [2:0] w_n8740_0;
	wire [1:0] w_n8744_0;
	wire [1:0] w_n8745_0;
	wire [2:0] w_n8746_0;
	wire [1:0] w_n8748_0;
	wire [1:0] w_n8753_0;
	wire [1:0] w_n8755_0;
	wire [1:0] w_n8756_0;
	wire [2:0] w_n8757_0;
	wire [1:0] w_n8758_0;
	wire [1:0] w_n8762_0;
	wire [1:0] w_n8768_0;
	wire [1:0] w_n8769_0;
	wire [1:0] w_n8771_0;
	wire [1:0] w_n8773_0;
	wire [1:0] w_n8776_0;
	wire [1:0] w_n8782_0;
	wire [1:0] w_n8784_0;
	wire [2:0] w_n8785_0;
	wire [1:0] w_n8789_0;
	wire [1:0] w_n8790_0;
	wire [2:0] w_n8791_0;
	wire [1:0] w_n8793_0;
	wire [1:0] w_n8798_0;
	wire [1:0] w_n8800_0;
	wire [1:0] w_n8801_0;
	wire [2:0] w_n8802_0;
	wire [1:0] w_n8803_0;
	wire [1:0] w_n8807_0;
	wire [1:0] w_n8813_0;
	wire [1:0] w_n8814_0;
	wire [1:0] w_n8816_0;
	wire [1:0] w_n8818_0;
	wire [1:0] w_n8821_0;
	wire [1:0] w_n8827_0;
	wire [1:0] w_n8829_0;
	wire [2:0] w_n8830_0;
	wire [1:0] w_n8834_0;
	wire [1:0] w_n8835_0;
	wire [2:0] w_n8836_0;
	wire [1:0] w_n8838_0;
	wire [1:0] w_n8843_0;
	wire [1:0] w_n8845_0;
	wire [1:0] w_n8846_0;
	wire [2:0] w_n8847_0;
	wire [1:0] w_n8848_0;
	wire [1:0] w_n8852_0;
	wire [1:0] w_n8858_0;
	wire [1:0] w_n8859_0;
	wire [1:0] w_n8861_0;
	wire [1:0] w_n8863_0;
	wire [1:0] w_n8866_0;
	wire [1:0] w_n8872_0;
	wire [2:0] w_n8874_0;
	wire [2:0] w_n8874_1;
	wire [1:0] w_n8877_0;
	wire [2:0] w_n8878_0;
	wire [1:0] w_n8879_0;
	wire [1:0] w_n8885_0;
	wire [2:0] w_n8886_0;
	wire [1:0] w_n8887_0;
	wire [1:0] w_n8892_0;
	wire [2:0] w_n8893_0;
	wire [2:0] w_n8893_1;
	wire [2:0] w_n8893_2;
	wire [2:0] w_n8893_3;
	wire [2:0] w_n8893_4;
	wire [2:0] w_n8893_5;
	wire [2:0] w_n8893_6;
	wire [2:0] w_n8893_7;
	wire [2:0] w_n8893_8;
	wire [2:0] w_n8893_9;
	wire [2:0] w_n8893_10;
	wire [2:0] w_n8893_11;
	wire [2:0] w_n8893_12;
	wire [2:0] w_n8893_13;
	wire [2:0] w_n8893_14;
	wire [2:0] w_n8893_15;
	wire [2:0] w_n8898_0;
	wire [2:0] w_n8898_1;
	wire [2:0] w_n8898_2;
	wire [2:0] w_n8898_3;
	wire [2:0] w_n8898_4;
	wire [2:0] w_n8898_5;
	wire [2:0] w_n8898_6;
	wire [2:0] w_n8898_7;
	wire [2:0] w_n8898_8;
	wire [2:0] w_n8898_9;
	wire [2:0] w_n8898_10;
	wire [2:0] w_n8898_11;
	wire [2:0] w_n8898_12;
	wire [2:0] w_n8898_13;
	wire [2:0] w_n8898_14;
	wire [2:0] w_n8898_15;
	wire [2:0] w_n8898_16;
	wire [2:0] w_n8898_17;
	wire [2:0] w_n8898_18;
	wire [2:0] w_n8898_19;
	wire [2:0] w_n8898_20;
	wire [2:0] w_n8898_21;
	wire [2:0] w_n8898_22;
	wire [2:0] w_n8898_23;
	wire [2:0] w_n8898_24;
	wire [2:0] w_n8898_25;
	wire [2:0] w_n8898_26;
	wire [1:0] w_n8898_27;
	wire [1:0] w_n8901_0;
	wire [2:0] w_n8903_0;
	wire [1:0] w_n8903_1;
	wire [2:0] w_n8904_0;
	wire [2:0] w_n8908_0;
	wire [1:0] w_n8909_0;
	wire [1:0] w_n8910_0;
	wire [1:0] w_n8911_0;
	wire [1:0] w_n8913_0;
	wire [1:0] w_n8915_0;
	wire [1:0] w_n8917_0;
	wire [1:0] w_n8920_0;
	wire [1:0] w_n8925_0;
	wire [2:0] w_n8927_0;
	wire [1:0] w_n8928_0;
	wire [1:0] w_n8932_0;
	wire [1:0] w_n8933_0;
	wire [1:0] w_n8935_0;
	wire [1:0] w_n8939_0;
	wire [1:0] w_n8941_0;
	wire [1:0] w_n8942_0;
	wire [2:0] w_n8943_0;
	wire [1:0] w_n8944_0;
	wire [1:0] w_n8948_0;
	wire [1:0] w_n8950_0;
	wire [1:0] w_n8952_0;
	wire [1:0] w_n8954_0;
	wire [1:0] w_n8957_0;
	wire [1:0] w_n8963_0;
	wire [2:0] w_n8965_0;
	wire [1:0] w_n8966_0;
	wire [1:0] w_n8971_0;
	wire [1:0] w_n8973_0;
	wire [1:0] w_n8975_0;
	wire [1:0] w_n8979_0;
	wire [1:0] w_n8981_0;
	wire [1:0] w_n8982_0;
	wire [2:0] w_n8983_0;
	wire [1:0] w_n8984_0;
	wire [1:0] w_n8990_0;
	wire [1:0] w_n8991_0;
	wire [1:0] w_n8993_0;
	wire [1:0] w_n8995_0;
	wire [1:0] w_n8997_0;
	wire [1:0] w_n9003_0;
	wire [1:0] w_n9005_0;
	wire [2:0] w_n9006_0;
	wire [1:0] w_n9009_0;
	wire [1:0] w_n9010_0;
	wire [2:0] w_n9011_0;
	wire [1:0] w_n9013_0;
	wire [1:0] w_n9017_0;
	wire [1:0] w_n9019_0;
	wire [1:0] w_n9020_0;
	wire [2:0] w_n9021_0;
	wire [1:0] w_n9022_0;
	wire [1:0] w_n9025_0;
	wire [1:0] w_n9031_0;
	wire [1:0] w_n9032_0;
	wire [1:0] w_n9034_0;
	wire [1:0] w_n9036_0;
	wire [1:0] w_n9038_0;
	wire [1:0] w_n9044_0;
	wire [1:0] w_n9046_0;
	wire [2:0] w_n9047_0;
	wire [1:0] w_n9050_0;
	wire [1:0] w_n9051_0;
	wire [2:0] w_n9052_0;
	wire [1:0] w_n9054_0;
	wire [1:0] w_n9056_0;
	wire [1:0] w_n9058_0;
	wire [1:0] w_n9064_0;
	wire [2:0] w_n9066_0;
	wire [1:0] w_n9067_0;
	wire [1:0] w_n9070_0;
	wire [1:0] w_n9072_0;
	wire [1:0] w_n9076_0;
	wire [1:0] w_n9078_0;
	wire [1:0] w_n9079_0;
	wire [1:0] w_n9080_0;
	wire [2:0] w_n9081_0;
	wire [1:0] w_n9084_0;
	wire [1:0] w_n9085_0;
	wire [2:0] w_n9086_0;
	wire [1:0] w_n9088_0;
	wire [1:0] w_n9092_0;
	wire [1:0] w_n9094_0;
	wire [1:0] w_n9095_0;
	wire [2:0] w_n9096_0;
	wire [1:0] w_n9097_0;
	wire [1:0] w_n9100_0;
	wire [1:0] w_n9106_0;
	wire [1:0] w_n9107_0;
	wire [1:0] w_n9109_0;
	wire [1:0] w_n9111_0;
	wire [1:0] w_n9113_0;
	wire [1:0] w_n9119_0;
	wire [1:0] w_n9121_0;
	wire [2:0] w_n9122_0;
	wire [1:0] w_n9125_0;
	wire [1:0] w_n9126_0;
	wire [2:0] w_n9127_0;
	wire [1:0] w_n9129_0;
	wire [1:0] w_n9133_0;
	wire [1:0] w_n9135_0;
	wire [1:0] w_n9136_0;
	wire [2:0] w_n9137_0;
	wire [1:0] w_n9138_0;
	wire [1:0] w_n9141_0;
	wire [1:0] w_n9147_0;
	wire [1:0] w_n9148_0;
	wire [1:0] w_n9150_0;
	wire [1:0] w_n9152_0;
	wire [1:0] w_n9154_0;
	wire [1:0] w_n9160_0;
	wire [1:0] w_n9162_0;
	wire [2:0] w_n9163_0;
	wire [1:0] w_n9166_0;
	wire [1:0] w_n9167_0;
	wire [2:0] w_n9168_0;
	wire [1:0] w_n9170_0;
	wire [1:0] w_n9174_0;
	wire [1:0] w_n9176_0;
	wire [1:0] w_n9177_0;
	wire [2:0] w_n9178_0;
	wire [1:0] w_n9179_0;
	wire [1:0] w_n9182_0;
	wire [1:0] w_n9188_0;
	wire [1:0] w_n9189_0;
	wire [1:0] w_n9191_0;
	wire [1:0] w_n9193_0;
	wire [1:0] w_n9195_0;
	wire [1:0] w_n9201_0;
	wire [1:0] w_n9203_0;
	wire [2:0] w_n9204_0;
	wire [1:0] w_n9207_0;
	wire [1:0] w_n9208_0;
	wire [2:0] w_n9209_0;
	wire [1:0] w_n9211_0;
	wire [1:0] w_n9215_0;
	wire [1:0] w_n9217_0;
	wire [1:0] w_n9218_0;
	wire [2:0] w_n9219_0;
	wire [1:0] w_n9220_0;
	wire [1:0] w_n9223_0;
	wire [1:0] w_n9229_0;
	wire [1:0] w_n9230_0;
	wire [1:0] w_n9232_0;
	wire [1:0] w_n9234_0;
	wire [1:0] w_n9236_0;
	wire [1:0] w_n9242_0;
	wire [1:0] w_n9244_0;
	wire [2:0] w_n9245_0;
	wire [1:0] w_n9248_0;
	wire [1:0] w_n9249_0;
	wire [2:0] w_n9250_0;
	wire [1:0] w_n9252_0;
	wire [1:0] w_n9256_0;
	wire [1:0] w_n9258_0;
	wire [1:0] w_n9259_0;
	wire [2:0] w_n9260_0;
	wire [1:0] w_n9261_0;
	wire [1:0] w_n9264_0;
	wire [1:0] w_n9270_0;
	wire [1:0] w_n9271_0;
	wire [1:0] w_n9273_0;
	wire [1:0] w_n9275_0;
	wire [1:0] w_n9277_0;
	wire [1:0] w_n9283_0;
	wire [2:0] w_n9285_0;
	wire [1:0] w_n9290_0;
	wire [2:0] w_n9292_0;
	wire [2:0] w_n9296_0;
	wire [1:0] w_n9297_0;
	wire [1:0] w_n9302_0;
	wire [2:0] w_n9303_0;
	wire [1:0] w_n9308_0;
	wire [1:0] w_n9315_0;
	wire [2:0] w_n9318_0;
	wire [1:0] w_n9318_1;
	wire [1:0] w_n9319_0;
	wire [2:0] w_n9322_0;
	wire [1:0] w_n9323_0;
	wire [1:0] w_n9324_0;
	wire [1:0] w_n9325_0;
	wire [1:0] w_n9327_0;
	wire [1:0] w_n9329_0;
	wire [1:0] w_n9331_0;
	wire [1:0] w_n9340_0;
	wire [2:0] w_n9342_0;
	wire [1:0] w_n9343_0;
	wire [1:0] w_n9347_0;
	wire [1:0] w_n9349_0;
	wire [1:0] w_n9351_0;
	wire [1:0] w_n9356_0;
	wire [1:0] w_n9358_0;
	wire [1:0] w_n9359_0;
	wire [2:0] w_n9360_0;
	wire [1:0] w_n9361_0;
	wire [1:0] w_n9366_0;
	wire [1:0] w_n9367_0;
	wire [1:0] w_n9369_0;
	wire [1:0] w_n9371_0;
	wire [1:0] w_n9374_0;
	wire [1:0] w_n9380_0;
	wire [2:0] w_n9382_0;
	wire [1:0] w_n9383_0;
	wire [1:0] w_n9387_0;
	wire [1:0] w_n9388_0;
	wire [1:0] w_n9390_0;
	wire [1:0] w_n9395_0;
	wire [1:0] w_n9397_0;
	wire [1:0] w_n9398_0;
	wire [2:0] w_n9399_0;
	wire [1:0] w_n9400_0;
	wire [1:0] w_n9404_0;
	wire [1:0] w_n9405_0;
	wire [1:0] w_n9407_0;
	wire [1:0] w_n9409_0;
	wire [1:0] w_n9412_0;
	wire [1:0] w_n9418_0;
	wire [1:0] w_n9420_0;
	wire [2:0] w_n9421_0;
	wire [1:0] w_n9425_0;
	wire [1:0] w_n9426_0;
	wire [2:0] w_n9427_0;
	wire [1:0] w_n9429_0;
	wire [1:0] w_n9434_0;
	wire [1:0] w_n9436_0;
	wire [1:0] w_n9437_0;
	wire [2:0] w_n9438_0;
	wire [1:0] w_n9439_0;
	wire [1:0] w_n9443_0;
	wire [1:0] w_n9449_0;
	wire [1:0] w_n9450_0;
	wire [1:0] w_n9452_0;
	wire [1:0] w_n9454_0;
	wire [1:0] w_n9457_0;
	wire [1:0] w_n9463_0;
	wire [1:0] w_n9465_0;
	wire [2:0] w_n9466_0;
	wire [1:0] w_n9470_0;
	wire [1:0] w_n9471_0;
	wire [2:0] w_n9472_0;
	wire [1:0] w_n9474_0;
	wire [1:0] w_n9479_0;
	wire [1:0] w_n9481_0;
	wire [1:0] w_n9482_0;
	wire [2:0] w_n9483_0;
	wire [1:0] w_n9484_0;
	wire [1:0] w_n9488_0;
	wire [1:0] w_n9494_0;
	wire [1:0] w_n9495_0;
	wire [1:0] w_n9497_0;
	wire [1:0] w_n9502_0;
	wire [1:0] w_n9504_0;
	wire [1:0] w_n9505_0;
	wire [2:0] w_n9506_0;
	wire [1:0] w_n9507_0;
	wire [1:0] w_n9509_0;
	wire [1:0] w_n9511_0;
	wire [1:0] w_n9513_0;
	wire [1:0] w_n9516_0;
	wire [1:0] w_n9522_0;
	wire [2:0] w_n9524_0;
	wire [1:0] w_n9525_0;
	wire [1:0] w_n9529_0;
	wire [1:0] w_n9535_0;
	wire [1:0] w_n9536_0;
	wire [1:0] w_n9538_0;
	wire [1:0] w_n9540_0;
	wire [1:0] w_n9543_0;
	wire [1:0] w_n9549_0;
	wire [1:0] w_n9551_0;
	wire [2:0] w_n9552_0;
	wire [1:0] w_n9556_0;
	wire [1:0] w_n9557_0;
	wire [2:0] w_n9558_0;
	wire [1:0] w_n9560_0;
	wire [1:0] w_n9565_0;
	wire [1:0] w_n9567_0;
	wire [1:0] w_n9568_0;
	wire [2:0] w_n9569_0;
	wire [1:0] w_n9570_0;
	wire [1:0] w_n9574_0;
	wire [1:0] w_n9580_0;
	wire [1:0] w_n9581_0;
	wire [1:0] w_n9583_0;
	wire [1:0] w_n9585_0;
	wire [1:0] w_n9588_0;
	wire [1:0] w_n9594_0;
	wire [1:0] w_n9596_0;
	wire [2:0] w_n9597_0;
	wire [1:0] w_n9601_0;
	wire [1:0] w_n9602_0;
	wire [2:0] w_n9603_0;
	wire [1:0] w_n9605_0;
	wire [1:0] w_n9610_0;
	wire [1:0] w_n9612_0;
	wire [1:0] w_n9613_0;
	wire [2:0] w_n9614_0;
	wire [1:0] w_n9615_0;
	wire [1:0] w_n9619_0;
	wire [1:0] w_n9625_0;
	wire [1:0] w_n9626_0;
	wire [1:0] w_n9628_0;
	wire [1:0] w_n9630_0;
	wire [1:0] w_n9633_0;
	wire [1:0] w_n9639_0;
	wire [1:0] w_n9641_0;
	wire [2:0] w_n9642_0;
	wire [1:0] w_n9646_0;
	wire [1:0] w_n9647_0;
	wire [2:0] w_n9648_0;
	wire [1:0] w_n9650_0;
	wire [1:0] w_n9655_0;
	wire [1:0] w_n9657_0;
	wire [1:0] w_n9658_0;
	wire [2:0] w_n9659_0;
	wire [1:0] w_n9660_0;
	wire [1:0] w_n9664_0;
	wire [1:0] w_n9670_0;
	wire [1:0] w_n9671_0;
	wire [1:0] w_n9673_0;
	wire [1:0] w_n9675_0;
	wire [1:0] w_n9678_0;
	wire [1:0] w_n9684_0;
	wire [1:0] w_n9686_0;
	wire [2:0] w_n9687_0;
	wire [1:0] w_n9691_0;
	wire [1:0] w_n9692_0;
	wire [2:0] w_n9693_0;
	wire [1:0] w_n9695_0;
	wire [1:0] w_n9700_0;
	wire [1:0] w_n9702_0;
	wire [1:0] w_n9703_0;
	wire [2:0] w_n9704_0;
	wire [1:0] w_n9705_0;
	wire [1:0] w_n9709_0;
	wire [1:0] w_n9715_0;
	wire [1:0] w_n9716_0;
	wire [1:0] w_n9718_0;
	wire [1:0] w_n9720_0;
	wire [1:0] w_n9723_0;
	wire [1:0] w_n9729_0;
	wire [1:0] w_n9731_0;
	wire [2:0] w_n9732_0;
	wire [1:0] w_n9736_0;
	wire [1:0] w_n9737_0;
	wire [2:0] w_n9738_0;
	wire [1:0] w_n9740_0;
	wire [1:0] w_n9745_0;
	wire [1:0] w_n9747_0;
	wire [1:0] w_n9748_0;
	wire [2:0] w_n9749_0;
	wire [2:0] w_n9749_1;
	wire [1:0] w_n9752_0;
	wire [2:0] w_n9753_0;
	wire [1:0] w_n9754_0;
	wire [1:0] w_n9755_0;
	wire [1:0] w_n9761_0;
	wire [2:0] w_n9762_0;
	wire [1:0] w_n9763_0;
	wire [1:0] w_n9768_0;
	wire [2:0] w_n9769_0;
	wire [2:0] w_n9769_1;
	wire [2:0] w_n9769_2;
	wire [2:0] w_n9769_3;
	wire [2:0] w_n9769_4;
	wire [2:0] w_n9769_5;
	wire [2:0] w_n9769_6;
	wire [2:0] w_n9769_7;
	wire [2:0] w_n9769_8;
	wire [2:0] w_n9769_9;
	wire [2:0] w_n9769_10;
	wire [2:0] w_n9769_11;
	wire [2:0] w_n9769_12;
	wire [2:0] w_n9769_13;
	wire [1:0] w_n9769_14;
	wire [2:0] w_n9774_0;
	wire [2:0] w_n9774_1;
	wire [2:0] w_n9774_2;
	wire [2:0] w_n9774_3;
	wire [2:0] w_n9774_4;
	wire [2:0] w_n9774_5;
	wire [2:0] w_n9774_6;
	wire [2:0] w_n9774_7;
	wire [2:0] w_n9774_8;
	wire [2:0] w_n9774_9;
	wire [2:0] w_n9774_10;
	wire [2:0] w_n9774_11;
	wire [2:0] w_n9774_12;
	wire [2:0] w_n9774_13;
	wire [2:0] w_n9774_14;
	wire [2:0] w_n9774_15;
	wire [2:0] w_n9774_16;
	wire [2:0] w_n9774_17;
	wire [2:0] w_n9774_18;
	wire [2:0] w_n9774_19;
	wire [2:0] w_n9774_20;
	wire [2:0] w_n9774_21;
	wire [2:0] w_n9774_22;
	wire [2:0] w_n9774_23;
	wire [2:0] w_n9774_24;
	wire [2:0] w_n9774_25;
	wire [1:0] w_n9778_0;
	wire [2:0] w_n9780_0;
	wire [1:0] w_n9780_1;
	wire [2:0] w_n9781_0;
	wire [2:0] w_n9785_0;
	wire [1:0] w_n9786_0;
	wire [1:0] w_n9787_0;
	wire [1:0] w_n9788_0;
	wire [1:0] w_n9790_0;
	wire [1:0] w_n9792_0;
	wire [1:0] w_n9794_0;
	wire [1:0] w_n9797_0;
	wire [1:0] w_n9802_0;
	wire [2:0] w_n9804_0;
	wire [1:0] w_n9805_0;
	wire [1:0] w_n9809_0;
	wire [1:0] w_n9810_0;
	wire [1:0] w_n9812_0;
	wire [1:0] w_n9816_0;
	wire [1:0] w_n9818_0;
	wire [1:0] w_n9819_0;
	wire [2:0] w_n9820_0;
	wire [1:0] w_n9821_0;
	wire [1:0] w_n9825_0;
	wire [1:0] w_n9827_0;
	wire [1:0] w_n9829_0;
	wire [1:0] w_n9831_0;
	wire [1:0] w_n9834_0;
	wire [1:0] w_n9840_0;
	wire [2:0] w_n9842_0;
	wire [1:0] w_n9843_0;
	wire [1:0] w_n9848_0;
	wire [1:0] w_n9850_0;
	wire [1:0] w_n9852_0;
	wire [1:0] w_n9856_0;
	wire [1:0] w_n9858_0;
	wire [1:0] w_n9859_0;
	wire [2:0] w_n9860_0;
	wire [1:0] w_n9861_0;
	wire [1:0] w_n9867_0;
	wire [1:0] w_n9868_0;
	wire [1:0] w_n9870_0;
	wire [1:0] w_n9872_0;
	wire [1:0] w_n9874_0;
	wire [1:0] w_n9880_0;
	wire [1:0] w_n9882_0;
	wire [2:0] w_n9883_0;
	wire [1:0] w_n9886_0;
	wire [1:0] w_n9887_0;
	wire [2:0] w_n9888_0;
	wire [1:0] w_n9890_0;
	wire [1:0] w_n9894_0;
	wire [1:0] w_n9896_0;
	wire [1:0] w_n9897_0;
	wire [2:0] w_n9898_0;
	wire [1:0] w_n9899_0;
	wire [1:0] w_n9902_0;
	wire [1:0] w_n9908_0;
	wire [1:0] w_n9909_0;
	wire [1:0] w_n9911_0;
	wire [1:0] w_n9913_0;
	wire [1:0] w_n9915_0;
	wire [1:0] w_n9921_0;
	wire [1:0] w_n9923_0;
	wire [2:0] w_n9924_0;
	wire [1:0] w_n9927_0;
	wire [1:0] w_n9928_0;
	wire [2:0] w_n9929_0;
	wire [1:0] w_n9931_0;
	wire [1:0] w_n9935_0;
	wire [1:0] w_n9937_0;
	wire [1:0] w_n9938_0;
	wire [2:0] w_n9939_0;
	wire [1:0] w_n9940_0;
	wire [1:0] w_n9943_0;
	wire [1:0] w_n9949_0;
	wire [1:0] w_n9950_0;
	wire [1:0] w_n9952_0;
	wire [1:0] w_n9954_0;
	wire [1:0] w_n9956_0;
	wire [1:0] w_n9962_0;
	wire [1:0] w_n9964_0;
	wire [2:0] w_n9965_0;
	wire [1:0] w_n9968_0;
	wire [1:0] w_n9969_0;
	wire [2:0] w_n9970_0;
	wire [1:0] w_n9972_0;
	wire [1:0] w_n9974_0;
	wire [1:0] w_n9976_0;
	wire [1:0] w_n9982_0;
	wire [2:0] w_n9984_0;
	wire [1:0] w_n9985_0;
	wire [1:0] w_n9987_0;
	wire [1:0] w_n9989_0;
	wire [1:0] w_n9993_0;
	wire [1:0] w_n9995_0;
	wire [1:0] w_n9996_0;
	wire [1:0] w_n9997_0;
	wire [2:0] w_n9998_0;
	wire [1:0] w_n10001_0;
	wire [1:0] w_n10002_0;
	wire [2:0] w_n10003_0;
	wire [1:0] w_n10005_0;
	wire [1:0] w_n10009_0;
	wire [1:0] w_n10011_0;
	wire [1:0] w_n10012_0;
	wire [2:0] w_n10013_0;
	wire [1:0] w_n10014_0;
	wire [1:0] w_n10017_0;
	wire [1:0] w_n10023_0;
	wire [1:0] w_n10024_0;
	wire [1:0] w_n10026_0;
	wire [1:0] w_n10028_0;
	wire [1:0] w_n10030_0;
	wire [1:0] w_n10036_0;
	wire [1:0] w_n10038_0;
	wire [2:0] w_n10039_0;
	wire [1:0] w_n10042_0;
	wire [1:0] w_n10043_0;
	wire [2:0] w_n10044_0;
	wire [1:0] w_n10046_0;
	wire [1:0] w_n10050_0;
	wire [1:0] w_n10052_0;
	wire [1:0] w_n10053_0;
	wire [2:0] w_n10054_0;
	wire [1:0] w_n10055_0;
	wire [1:0] w_n10058_0;
	wire [1:0] w_n10064_0;
	wire [1:0] w_n10065_0;
	wire [1:0] w_n10067_0;
	wire [1:0] w_n10069_0;
	wire [1:0] w_n10071_0;
	wire [1:0] w_n10077_0;
	wire [1:0] w_n10079_0;
	wire [2:0] w_n10080_0;
	wire [1:0] w_n10083_0;
	wire [1:0] w_n10084_0;
	wire [2:0] w_n10085_0;
	wire [1:0] w_n10087_0;
	wire [1:0] w_n10091_0;
	wire [1:0] w_n10093_0;
	wire [1:0] w_n10094_0;
	wire [2:0] w_n10095_0;
	wire [1:0] w_n10096_0;
	wire [1:0] w_n10099_0;
	wire [1:0] w_n10105_0;
	wire [1:0] w_n10106_0;
	wire [1:0] w_n10108_0;
	wire [1:0] w_n10110_0;
	wire [1:0] w_n10112_0;
	wire [1:0] w_n10118_0;
	wire [1:0] w_n10120_0;
	wire [2:0] w_n10121_0;
	wire [1:0] w_n10124_0;
	wire [1:0] w_n10125_0;
	wire [2:0] w_n10126_0;
	wire [1:0] w_n10128_0;
	wire [1:0] w_n10132_0;
	wire [1:0] w_n10134_0;
	wire [1:0] w_n10135_0;
	wire [2:0] w_n10136_0;
	wire [1:0] w_n10137_0;
	wire [1:0] w_n10140_0;
	wire [1:0] w_n10146_0;
	wire [1:0] w_n10147_0;
	wire [1:0] w_n10149_0;
	wire [1:0] w_n10151_0;
	wire [1:0] w_n10153_0;
	wire [1:0] w_n10159_0;
	wire [1:0] w_n10161_0;
	wire [2:0] w_n10162_0;
	wire [1:0] w_n10165_0;
	wire [1:0] w_n10166_0;
	wire [2:0] w_n10167_0;
	wire [1:0] w_n10169_0;
	wire [1:0] w_n10173_0;
	wire [1:0] w_n10175_0;
	wire [1:0] w_n10176_0;
	wire [2:0] w_n10177_0;
	wire [1:0] w_n10181_0;
	wire [1:0] w_n10187_0;
	wire [2:0] w_n10189_0;
	wire [1:0] w_n10191_0;
	wire [2:0] w_n10196_0;
	wire [1:0] w_n10197_0;
	wire [1:0] w_n10198_0;
	wire [1:0] w_n10203_0;
	wire [2:0] w_n10204_0;
	wire [1:0] w_n10209_0;
	wire [1:0] w_n10217_0;
	wire [2:0] w_n10219_0;
	wire [1:0] w_n10219_1;
	wire [1:0] w_n10220_0;
	wire [2:0] w_n10223_0;
	wire [1:0] w_n10224_0;
	wire [1:0] w_n10225_0;
	wire [1:0] w_n10226_0;
	wire [1:0] w_n10228_0;
	wire [1:0] w_n10230_0;
	wire [1:0] w_n10232_0;
	wire [1:0] w_n10241_0;
	wire [2:0] w_n10243_0;
	wire [1:0] w_n10244_0;
	wire [1:0] w_n10248_0;
	wire [1:0] w_n10250_0;
	wire [1:0] w_n10252_0;
	wire [1:0] w_n10257_0;
	wire [1:0] w_n10259_0;
	wire [1:0] w_n10260_0;
	wire [2:0] w_n10261_0;
	wire [1:0] w_n10262_0;
	wire [1:0] w_n10267_0;
	wire [1:0] w_n10268_0;
	wire [1:0] w_n10270_0;
	wire [1:0] w_n10272_0;
	wire [1:0] w_n10275_0;
	wire [1:0] w_n10281_0;
	wire [2:0] w_n10283_0;
	wire [1:0] w_n10284_0;
	wire [1:0] w_n10288_0;
	wire [1:0] w_n10289_0;
	wire [1:0] w_n10291_0;
	wire [1:0] w_n10296_0;
	wire [1:0] w_n10298_0;
	wire [1:0] w_n10299_0;
	wire [2:0] w_n10300_0;
	wire [1:0] w_n10301_0;
	wire [1:0] w_n10305_0;
	wire [1:0] w_n10306_0;
	wire [1:0] w_n10308_0;
	wire [1:0] w_n10310_0;
	wire [1:0] w_n10313_0;
	wire [1:0] w_n10319_0;
	wire [1:0] w_n10321_0;
	wire [2:0] w_n10322_0;
	wire [1:0] w_n10326_0;
	wire [1:0] w_n10327_0;
	wire [2:0] w_n10328_0;
	wire [1:0] w_n10330_0;
	wire [1:0] w_n10335_0;
	wire [1:0] w_n10337_0;
	wire [1:0] w_n10338_0;
	wire [2:0] w_n10339_0;
	wire [1:0] w_n10340_0;
	wire [1:0] w_n10344_0;
	wire [1:0] w_n10350_0;
	wire [1:0] w_n10351_0;
	wire [1:0] w_n10353_0;
	wire [1:0] w_n10355_0;
	wire [1:0] w_n10358_0;
	wire [1:0] w_n10364_0;
	wire [1:0] w_n10366_0;
	wire [2:0] w_n10367_0;
	wire [1:0] w_n10371_0;
	wire [1:0] w_n10372_0;
	wire [2:0] w_n10373_0;
	wire [1:0] w_n10375_0;
	wire [1:0] w_n10380_0;
	wire [1:0] w_n10382_0;
	wire [1:0] w_n10383_0;
	wire [2:0] w_n10384_0;
	wire [1:0] w_n10385_0;
	wire [1:0] w_n10389_0;
	wire [1:0] w_n10395_0;
	wire [1:0] w_n10396_0;
	wire [1:0] w_n10398_0;
	wire [1:0] w_n10400_0;
	wire [1:0] w_n10403_0;
	wire [1:0] w_n10409_0;
	wire [1:0] w_n10411_0;
	wire [2:0] w_n10412_0;
	wire [1:0] w_n10416_0;
	wire [1:0] w_n10417_0;
	wire [2:0] w_n10418_0;
	wire [1:0] w_n10420_0;
	wire [1:0] w_n10425_0;
	wire [1:0] w_n10427_0;
	wire [1:0] w_n10428_0;
	wire [2:0] w_n10429_0;
	wire [1:0] w_n10430_0;
	wire [1:0] w_n10434_0;
	wire [1:0] w_n10440_0;
	wire [1:0] w_n10441_0;
	wire [1:0] w_n10443_0;
	wire [1:0] w_n10448_0;
	wire [1:0] w_n10450_0;
	wire [1:0] w_n10451_0;
	wire [2:0] w_n10452_0;
	wire [1:0] w_n10453_0;
	wire [1:0] w_n10455_0;
	wire [1:0] w_n10457_0;
	wire [1:0] w_n10459_0;
	wire [1:0] w_n10462_0;
	wire [1:0] w_n10468_0;
	wire [2:0] w_n10470_0;
	wire [1:0] w_n10471_0;
	wire [1:0] w_n10475_0;
	wire [1:0] w_n10481_0;
	wire [1:0] w_n10482_0;
	wire [1:0] w_n10484_0;
	wire [1:0] w_n10486_0;
	wire [1:0] w_n10489_0;
	wire [1:0] w_n10495_0;
	wire [1:0] w_n10497_0;
	wire [2:0] w_n10498_0;
	wire [1:0] w_n10502_0;
	wire [1:0] w_n10503_0;
	wire [2:0] w_n10504_0;
	wire [1:0] w_n10506_0;
	wire [1:0] w_n10511_0;
	wire [1:0] w_n10513_0;
	wire [1:0] w_n10514_0;
	wire [2:0] w_n10515_0;
	wire [1:0] w_n10516_0;
	wire [1:0] w_n10520_0;
	wire [1:0] w_n10526_0;
	wire [1:0] w_n10527_0;
	wire [1:0] w_n10529_0;
	wire [1:0] w_n10531_0;
	wire [1:0] w_n10534_0;
	wire [1:0] w_n10540_0;
	wire [1:0] w_n10542_0;
	wire [2:0] w_n10543_0;
	wire [1:0] w_n10547_0;
	wire [1:0] w_n10548_0;
	wire [2:0] w_n10549_0;
	wire [1:0] w_n10551_0;
	wire [1:0] w_n10556_0;
	wire [1:0] w_n10558_0;
	wire [1:0] w_n10559_0;
	wire [2:0] w_n10560_0;
	wire [1:0] w_n10561_0;
	wire [1:0] w_n10565_0;
	wire [1:0] w_n10571_0;
	wire [1:0] w_n10572_0;
	wire [1:0] w_n10574_0;
	wire [1:0] w_n10576_0;
	wire [1:0] w_n10579_0;
	wire [1:0] w_n10585_0;
	wire [1:0] w_n10587_0;
	wire [2:0] w_n10588_0;
	wire [1:0] w_n10592_0;
	wire [1:0] w_n10593_0;
	wire [2:0] w_n10594_0;
	wire [1:0] w_n10596_0;
	wire [1:0] w_n10601_0;
	wire [1:0] w_n10603_0;
	wire [1:0] w_n10604_0;
	wire [2:0] w_n10605_0;
	wire [1:0] w_n10606_0;
	wire [1:0] w_n10610_0;
	wire [1:0] w_n10616_0;
	wire [1:0] w_n10617_0;
	wire [1:0] w_n10619_0;
	wire [1:0] w_n10621_0;
	wire [1:0] w_n10624_0;
	wire [1:0] w_n10630_0;
	wire [1:0] w_n10632_0;
	wire [2:0] w_n10633_0;
	wire [1:0] w_n10637_0;
	wire [1:0] w_n10638_0;
	wire [2:0] w_n10639_0;
	wire [1:0] w_n10641_0;
	wire [1:0] w_n10646_0;
	wire [1:0] w_n10648_0;
	wire [1:0] w_n10649_0;
	wire [2:0] w_n10650_0;
	wire [1:0] w_n10651_0;
	wire [1:0] w_n10655_0;
	wire [1:0] w_n10661_0;
	wire [1:0] w_n10662_0;
	wire [1:0] w_n10664_0;
	wire [1:0] w_n10666_0;
	wire [1:0] w_n10669_0;
	wire [1:0] w_n10675_0;
	wire [2:0] w_n10677_0;
	wire [2:0] w_n10677_1;
	wire [1:0] w_n10680_0;
	wire [2:0] w_n10681_0;
	wire [1:0] w_n10682_0;
	wire [1:0] w_n10688_0;
	wire [2:0] w_n10689_0;
	wire [1:0] w_n10690_0;
	wire [1:0] w_n10695_0;
	wire [2:0] w_n10696_0;
	wire [2:0] w_n10696_1;
	wire [2:0] w_n10696_2;
	wire [2:0] w_n10696_3;
	wire [2:0] w_n10696_4;
	wire [2:0] w_n10696_5;
	wire [2:0] w_n10696_6;
	wire [2:0] w_n10696_7;
	wire [2:0] w_n10696_8;
	wire [2:0] w_n10696_9;
	wire [2:0] w_n10696_10;
	wire [2:0] w_n10696_11;
	wire [2:0] w_n10696_12;
	wire [1:0] w_n10696_13;
	wire [2:0] w_n10701_0;
	wire [2:0] w_n10701_1;
	wire [2:0] w_n10701_2;
	wire [2:0] w_n10701_3;
	wire [2:0] w_n10701_4;
	wire [2:0] w_n10701_5;
	wire [2:0] w_n10701_6;
	wire [2:0] w_n10701_7;
	wire [2:0] w_n10701_8;
	wire [2:0] w_n10701_9;
	wire [2:0] w_n10701_10;
	wire [2:0] w_n10701_11;
	wire [2:0] w_n10701_12;
	wire [2:0] w_n10701_13;
	wire [2:0] w_n10701_14;
	wire [2:0] w_n10701_15;
	wire [2:0] w_n10701_16;
	wire [2:0] w_n10701_17;
	wire [2:0] w_n10701_18;
	wire [2:0] w_n10701_19;
	wire [2:0] w_n10701_20;
	wire [2:0] w_n10701_21;
	wire [2:0] w_n10701_22;
	wire [2:0] w_n10701_23;
	wire [2:0] w_n10701_24;
	wire [2:0] w_n10701_25;
	wire [1:0] w_n10704_0;
	wire [2:0] w_n10706_0;
	wire [1:0] w_n10706_1;
	wire [2:0] w_n10707_0;
	wire [2:0] w_n10711_0;
	wire [1:0] w_n10712_0;
	wire [1:0] w_n10713_0;
	wire [1:0] w_n10714_0;
	wire [1:0] w_n10716_0;
	wire [1:0] w_n10718_0;
	wire [1:0] w_n10720_0;
	wire [1:0] w_n10723_0;
	wire [1:0] w_n10728_0;
	wire [2:0] w_n10730_0;
	wire [1:0] w_n10731_0;
	wire [1:0] w_n10735_0;
	wire [1:0] w_n10736_0;
	wire [1:0] w_n10738_0;
	wire [1:0] w_n10742_0;
	wire [1:0] w_n10744_0;
	wire [1:0] w_n10745_0;
	wire [2:0] w_n10746_0;
	wire [1:0] w_n10747_0;
	wire [1:0] w_n10751_0;
	wire [1:0] w_n10753_0;
	wire [1:0] w_n10755_0;
	wire [1:0] w_n10757_0;
	wire [1:0] w_n10760_0;
	wire [1:0] w_n10766_0;
	wire [2:0] w_n10768_0;
	wire [1:0] w_n10769_0;
	wire [1:0] w_n10774_0;
	wire [1:0] w_n10776_0;
	wire [1:0] w_n10778_0;
	wire [1:0] w_n10782_0;
	wire [1:0] w_n10784_0;
	wire [1:0] w_n10785_0;
	wire [2:0] w_n10786_0;
	wire [1:0] w_n10787_0;
	wire [1:0] w_n10793_0;
	wire [1:0] w_n10794_0;
	wire [1:0] w_n10796_0;
	wire [1:0] w_n10798_0;
	wire [1:0] w_n10800_0;
	wire [1:0] w_n10806_0;
	wire [1:0] w_n10808_0;
	wire [2:0] w_n10809_0;
	wire [1:0] w_n10812_0;
	wire [1:0] w_n10813_0;
	wire [2:0] w_n10814_0;
	wire [1:0] w_n10816_0;
	wire [1:0] w_n10820_0;
	wire [1:0] w_n10822_0;
	wire [1:0] w_n10823_0;
	wire [2:0] w_n10824_0;
	wire [1:0] w_n10825_0;
	wire [1:0] w_n10828_0;
	wire [1:0] w_n10834_0;
	wire [1:0] w_n10835_0;
	wire [1:0] w_n10837_0;
	wire [1:0] w_n10839_0;
	wire [1:0] w_n10841_0;
	wire [1:0] w_n10847_0;
	wire [1:0] w_n10849_0;
	wire [2:0] w_n10850_0;
	wire [1:0] w_n10853_0;
	wire [1:0] w_n10854_0;
	wire [2:0] w_n10855_0;
	wire [1:0] w_n10857_0;
	wire [1:0] w_n10861_0;
	wire [1:0] w_n10863_0;
	wire [1:0] w_n10864_0;
	wire [2:0] w_n10865_0;
	wire [1:0] w_n10866_0;
	wire [1:0] w_n10869_0;
	wire [1:0] w_n10875_0;
	wire [1:0] w_n10876_0;
	wire [1:0] w_n10878_0;
	wire [1:0] w_n10880_0;
	wire [1:0] w_n10882_0;
	wire [1:0] w_n10888_0;
	wire [1:0] w_n10890_0;
	wire [2:0] w_n10891_0;
	wire [1:0] w_n10894_0;
	wire [1:0] w_n10895_0;
	wire [2:0] w_n10896_0;
	wire [1:0] w_n10898_0;
	wire [1:0] w_n10902_0;
	wire [1:0] w_n10904_0;
	wire [1:0] w_n10905_0;
	wire [2:0] w_n10906_0;
	wire [1:0] w_n10907_0;
	wire [1:0] w_n10910_0;
	wire [1:0] w_n10916_0;
	wire [1:0] w_n10917_0;
	wire [1:0] w_n10919_0;
	wire [1:0] w_n10921_0;
	wire [1:0] w_n10923_0;
	wire [1:0] w_n10929_0;
	wire [1:0] w_n10931_0;
	wire [2:0] w_n10932_0;
	wire [1:0] w_n10935_0;
	wire [1:0] w_n10936_0;
	wire [2:0] w_n10937_0;
	wire [1:0] w_n10939_0;
	wire [1:0] w_n10941_0;
	wire [1:0] w_n10943_0;
	wire [1:0] w_n10949_0;
	wire [2:0] w_n10951_0;
	wire [1:0] w_n10952_0;
	wire [1:0] w_n10954_0;
	wire [1:0] w_n10956_0;
	wire [1:0] w_n10960_0;
	wire [1:0] w_n10962_0;
	wire [1:0] w_n10963_0;
	wire [1:0] w_n10964_0;
	wire [2:0] w_n10965_0;
	wire [1:0] w_n10968_0;
	wire [1:0] w_n10969_0;
	wire [2:0] w_n10970_0;
	wire [1:0] w_n10972_0;
	wire [1:0] w_n10976_0;
	wire [1:0] w_n10978_0;
	wire [1:0] w_n10979_0;
	wire [2:0] w_n10980_0;
	wire [1:0] w_n10981_0;
	wire [1:0] w_n10984_0;
	wire [1:0] w_n10990_0;
	wire [1:0] w_n10991_0;
	wire [1:0] w_n10993_0;
	wire [1:0] w_n10995_0;
	wire [1:0] w_n10997_0;
	wire [1:0] w_n11003_0;
	wire [1:0] w_n11005_0;
	wire [2:0] w_n11006_0;
	wire [1:0] w_n11009_0;
	wire [1:0] w_n11010_0;
	wire [2:0] w_n11011_0;
	wire [1:0] w_n11013_0;
	wire [1:0] w_n11017_0;
	wire [1:0] w_n11019_0;
	wire [1:0] w_n11020_0;
	wire [2:0] w_n11021_0;
	wire [1:0] w_n11022_0;
	wire [1:0] w_n11025_0;
	wire [1:0] w_n11031_0;
	wire [1:0] w_n11032_0;
	wire [1:0] w_n11034_0;
	wire [1:0] w_n11036_0;
	wire [1:0] w_n11038_0;
	wire [1:0] w_n11044_0;
	wire [1:0] w_n11046_0;
	wire [2:0] w_n11047_0;
	wire [1:0] w_n11050_0;
	wire [1:0] w_n11051_0;
	wire [2:0] w_n11052_0;
	wire [1:0] w_n11054_0;
	wire [1:0] w_n11058_0;
	wire [1:0] w_n11060_0;
	wire [1:0] w_n11061_0;
	wire [2:0] w_n11062_0;
	wire [1:0] w_n11063_0;
	wire [1:0] w_n11066_0;
	wire [1:0] w_n11072_0;
	wire [1:0] w_n11073_0;
	wire [1:0] w_n11075_0;
	wire [1:0] w_n11077_0;
	wire [1:0] w_n11079_0;
	wire [1:0] w_n11085_0;
	wire [1:0] w_n11087_0;
	wire [2:0] w_n11088_0;
	wire [1:0] w_n11091_0;
	wire [1:0] w_n11092_0;
	wire [2:0] w_n11093_0;
	wire [1:0] w_n11095_0;
	wire [1:0] w_n11099_0;
	wire [1:0] w_n11101_0;
	wire [1:0] w_n11102_0;
	wire [2:0] w_n11103_0;
	wire [1:0] w_n11104_0;
	wire [1:0] w_n11107_0;
	wire [1:0] w_n11113_0;
	wire [1:0] w_n11114_0;
	wire [1:0] w_n11116_0;
	wire [1:0] w_n11118_0;
	wire [1:0] w_n11120_0;
	wire [1:0] w_n11126_0;
	wire [2:0] w_n11128_0;
	wire [1:0] w_n11133_0;
	wire [2:0] w_n11135_0;
	wire [2:0] w_n11139_0;
	wire [1:0] w_n11140_0;
	wire [1:0] w_n11145_0;
	wire [2:0] w_n11146_0;
	wire [1:0] w_n11151_0;
	wire [1:0] w_n11158_0;
	wire [2:0] w_n11160_0;
	wire [1:0] w_n11160_1;
	wire [1:0] w_n11161_0;
	wire [2:0] w_n11164_0;
	wire [1:0] w_n11165_0;
	wire [1:0] w_n11166_0;
	wire [1:0] w_n11167_0;
	wire [1:0] w_n11169_0;
	wire [1:0] w_n11171_0;
	wire [1:0] w_n11173_0;
	wire [1:0] w_n11182_0;
	wire [2:0] w_n11184_0;
	wire [1:0] w_n11185_0;
	wire [1:0] w_n11189_0;
	wire [1:0] w_n11191_0;
	wire [1:0] w_n11193_0;
	wire [1:0] w_n11198_0;
	wire [1:0] w_n11200_0;
	wire [1:0] w_n11201_0;
	wire [2:0] w_n11202_0;
	wire [1:0] w_n11203_0;
	wire [1:0] w_n11208_0;
	wire [1:0] w_n11209_0;
	wire [1:0] w_n11211_0;
	wire [1:0] w_n11213_0;
	wire [1:0] w_n11216_0;
	wire [1:0] w_n11222_0;
	wire [2:0] w_n11224_0;
	wire [1:0] w_n11225_0;
	wire [1:0] w_n11229_0;
	wire [1:0] w_n11230_0;
	wire [1:0] w_n11232_0;
	wire [1:0] w_n11237_0;
	wire [1:0] w_n11239_0;
	wire [1:0] w_n11240_0;
	wire [2:0] w_n11241_0;
	wire [1:0] w_n11242_0;
	wire [1:0] w_n11246_0;
	wire [1:0] w_n11247_0;
	wire [1:0] w_n11249_0;
	wire [1:0] w_n11251_0;
	wire [1:0] w_n11254_0;
	wire [1:0] w_n11260_0;
	wire [1:0] w_n11262_0;
	wire [2:0] w_n11263_0;
	wire [1:0] w_n11267_0;
	wire [1:0] w_n11268_0;
	wire [2:0] w_n11269_0;
	wire [1:0] w_n11271_0;
	wire [1:0] w_n11276_0;
	wire [1:0] w_n11278_0;
	wire [1:0] w_n11279_0;
	wire [2:0] w_n11280_0;
	wire [1:0] w_n11281_0;
	wire [1:0] w_n11285_0;
	wire [1:0] w_n11291_0;
	wire [1:0] w_n11292_0;
	wire [1:0] w_n11294_0;
	wire [1:0] w_n11296_0;
	wire [1:0] w_n11299_0;
	wire [1:0] w_n11305_0;
	wire [1:0] w_n11307_0;
	wire [2:0] w_n11308_0;
	wire [1:0] w_n11312_0;
	wire [1:0] w_n11313_0;
	wire [2:0] w_n11314_0;
	wire [1:0] w_n11316_0;
	wire [1:0] w_n11321_0;
	wire [1:0] w_n11323_0;
	wire [1:0] w_n11324_0;
	wire [2:0] w_n11325_0;
	wire [1:0] w_n11326_0;
	wire [1:0] w_n11330_0;
	wire [1:0] w_n11336_0;
	wire [1:0] w_n11337_0;
	wire [1:0] w_n11339_0;
	wire [1:0] w_n11341_0;
	wire [1:0] w_n11344_0;
	wire [1:0] w_n11350_0;
	wire [1:0] w_n11352_0;
	wire [2:0] w_n11353_0;
	wire [1:0] w_n11357_0;
	wire [1:0] w_n11358_0;
	wire [2:0] w_n11359_0;
	wire [1:0] w_n11361_0;
	wire [1:0] w_n11366_0;
	wire [1:0] w_n11368_0;
	wire [1:0] w_n11369_0;
	wire [2:0] w_n11370_0;
	wire [1:0] w_n11371_0;
	wire [1:0] w_n11375_0;
	wire [1:0] w_n11381_0;
	wire [1:0] w_n11382_0;
	wire [1:0] w_n11384_0;
	wire [1:0] w_n11386_0;
	wire [1:0] w_n11389_0;
	wire [1:0] w_n11395_0;
	wire [1:0] w_n11397_0;
	wire [2:0] w_n11398_0;
	wire [1:0] w_n11402_0;
	wire [1:0] w_n11403_0;
	wire [2:0] w_n11404_0;
	wire [1:0] w_n11406_0;
	wire [1:0] w_n11411_0;
	wire [1:0] w_n11413_0;
	wire [1:0] w_n11414_0;
	wire [2:0] w_n11415_0;
	wire [1:0] w_n11416_0;
	wire [1:0] w_n11420_0;
	wire [1:0] w_n11426_0;
	wire [1:0] w_n11427_0;
	wire [1:0] w_n11429_0;
	wire [1:0] w_n11434_0;
	wire [1:0] w_n11436_0;
	wire [1:0] w_n11437_0;
	wire [2:0] w_n11438_0;
	wire [1:0] w_n11439_0;
	wire [1:0] w_n11442_0;
	wire [1:0] w_n11444_0;
	wire [1:0] w_n11446_0;
	wire [1:0] w_n11449_0;
	wire [1:0] w_n11455_0;
	wire [2:0] w_n11457_0;
	wire [1:0] w_n11458_0;
	wire [1:0] w_n11462_0;
	wire [1:0] w_n11468_0;
	wire [1:0] w_n11469_0;
	wire [1:0] w_n11471_0;
	wire [1:0] w_n11473_0;
	wire [1:0] w_n11476_0;
	wire [1:0] w_n11482_0;
	wire [1:0] w_n11484_0;
	wire [2:0] w_n11485_0;
	wire [1:0] w_n11489_0;
	wire [1:0] w_n11490_0;
	wire [2:0] w_n11491_0;
	wire [1:0] w_n11493_0;
	wire [1:0] w_n11498_0;
	wire [1:0] w_n11500_0;
	wire [1:0] w_n11501_0;
	wire [2:0] w_n11502_0;
	wire [1:0] w_n11503_0;
	wire [1:0] w_n11507_0;
	wire [1:0] w_n11513_0;
	wire [1:0] w_n11514_0;
	wire [1:0] w_n11516_0;
	wire [1:0] w_n11518_0;
	wire [1:0] w_n11521_0;
	wire [1:0] w_n11527_0;
	wire [1:0] w_n11529_0;
	wire [2:0] w_n11530_0;
	wire [1:0] w_n11534_0;
	wire [1:0] w_n11535_0;
	wire [2:0] w_n11536_0;
	wire [1:0] w_n11538_0;
	wire [1:0] w_n11543_0;
	wire [1:0] w_n11545_0;
	wire [1:0] w_n11546_0;
	wire [2:0] w_n11547_0;
	wire [1:0] w_n11548_0;
	wire [1:0] w_n11552_0;
	wire [1:0] w_n11558_0;
	wire [1:0] w_n11559_0;
	wire [1:0] w_n11561_0;
	wire [1:0] w_n11563_0;
	wire [1:0] w_n11566_0;
	wire [1:0] w_n11572_0;
	wire [1:0] w_n11574_0;
	wire [2:0] w_n11575_0;
	wire [1:0] w_n11579_0;
	wire [1:0] w_n11580_0;
	wire [2:0] w_n11581_0;
	wire [1:0] w_n11583_0;
	wire [1:0] w_n11588_0;
	wire [1:0] w_n11590_0;
	wire [1:0] w_n11591_0;
	wire [2:0] w_n11592_0;
	wire [1:0] w_n11593_0;
	wire [1:0] w_n11597_0;
	wire [1:0] w_n11603_0;
	wire [1:0] w_n11604_0;
	wire [1:0] w_n11606_0;
	wire [1:0] w_n11608_0;
	wire [1:0] w_n11611_0;
	wire [1:0] w_n11617_0;
	wire [1:0] w_n11619_0;
	wire [2:0] w_n11620_0;
	wire [1:0] w_n11624_0;
	wire [1:0] w_n11625_0;
	wire [2:0] w_n11626_0;
	wire [1:0] w_n11628_0;
	wire [1:0] w_n11633_0;
	wire [1:0] w_n11635_0;
	wire [1:0] w_n11636_0;
	wire [2:0] w_n11637_0;
	wire [2:0] w_n11637_1;
	wire [1:0] w_n11640_0;
	wire [2:0] w_n11641_0;
	wire [1:0] w_n11642_0;
	wire [1:0] w_n11643_0;
	wire [1:0] w_n11649_0;
	wire [2:0] w_n11650_0;
	wire [1:0] w_n11651_0;
	wire [1:0] w_n11656_0;
	wire [2:0] w_n11657_0;
	wire [2:0] w_n11657_1;
	wire [2:0] w_n11657_2;
	wire [2:0] w_n11657_3;
	wire [2:0] w_n11657_4;
	wire [2:0] w_n11657_5;
	wire [2:0] w_n11657_6;
	wire [2:0] w_n11657_7;
	wire [2:0] w_n11657_8;
	wire [2:0] w_n11657_9;
	wire [2:0] w_n11657_10;
	wire [2:0] w_n11657_11;
	wire [2:0] w_n11662_0;
	wire [2:0] w_n11662_1;
	wire [2:0] w_n11662_2;
	wire [2:0] w_n11662_3;
	wire [2:0] w_n11662_4;
	wire [2:0] w_n11662_5;
	wire [2:0] w_n11662_6;
	wire [2:0] w_n11662_7;
	wire [2:0] w_n11662_8;
	wire [2:0] w_n11662_9;
	wire [2:0] w_n11662_10;
	wire [2:0] w_n11662_11;
	wire [2:0] w_n11662_12;
	wire [2:0] w_n11662_13;
	wire [2:0] w_n11662_14;
	wire [2:0] w_n11662_15;
	wire [2:0] w_n11662_16;
	wire [2:0] w_n11662_17;
	wire [2:0] w_n11662_18;
	wire [2:0] w_n11662_19;
	wire [2:0] w_n11662_20;
	wire [2:0] w_n11662_21;
	wire [2:0] w_n11662_22;
	wire [2:0] w_n11662_23;
	wire [1:0] w_n11662_24;
	wire [1:0] w_n11665_0;
	wire [2:0] w_n11667_0;
	wire [1:0] w_n11667_1;
	wire [2:0] w_n11668_0;
	wire [2:0] w_n11672_0;
	wire [1:0] w_n11673_0;
	wire [1:0] w_n11674_0;
	wire [1:0] w_n11675_0;
	wire [1:0] w_n11677_0;
	wire [1:0] w_n11679_0;
	wire [1:0] w_n11681_0;
	wire [1:0] w_n11684_0;
	wire [1:0] w_n11689_0;
	wire [2:0] w_n11691_0;
	wire [1:0] w_n11692_0;
	wire [1:0] w_n11696_0;
	wire [1:0] w_n11697_0;
	wire [1:0] w_n11699_0;
	wire [1:0] w_n11703_0;
	wire [1:0] w_n11705_0;
	wire [1:0] w_n11706_0;
	wire [2:0] w_n11707_0;
	wire [1:0] w_n11708_0;
	wire [1:0] w_n11712_0;
	wire [1:0] w_n11714_0;
	wire [1:0] w_n11716_0;
	wire [1:0] w_n11718_0;
	wire [1:0] w_n11721_0;
	wire [1:0] w_n11727_0;
	wire [2:0] w_n11729_0;
	wire [1:0] w_n11730_0;
	wire [1:0] w_n11735_0;
	wire [1:0] w_n11737_0;
	wire [1:0] w_n11739_0;
	wire [1:0] w_n11743_0;
	wire [1:0] w_n11745_0;
	wire [1:0] w_n11746_0;
	wire [2:0] w_n11747_0;
	wire [1:0] w_n11748_0;
	wire [1:0] w_n11754_0;
	wire [1:0] w_n11755_0;
	wire [1:0] w_n11757_0;
	wire [1:0] w_n11759_0;
	wire [1:0] w_n11761_0;
	wire [1:0] w_n11767_0;
	wire [1:0] w_n11769_0;
	wire [2:0] w_n11770_0;
	wire [1:0] w_n11773_0;
	wire [1:0] w_n11774_0;
	wire [2:0] w_n11775_0;
	wire [1:0] w_n11777_0;
	wire [1:0] w_n11781_0;
	wire [1:0] w_n11783_0;
	wire [1:0] w_n11784_0;
	wire [2:0] w_n11785_0;
	wire [1:0] w_n11786_0;
	wire [1:0] w_n11789_0;
	wire [1:0] w_n11795_0;
	wire [1:0] w_n11796_0;
	wire [1:0] w_n11798_0;
	wire [1:0] w_n11800_0;
	wire [1:0] w_n11802_0;
	wire [1:0] w_n11808_0;
	wire [1:0] w_n11810_0;
	wire [2:0] w_n11811_0;
	wire [1:0] w_n11814_0;
	wire [1:0] w_n11815_0;
	wire [2:0] w_n11816_0;
	wire [1:0] w_n11818_0;
	wire [1:0] w_n11822_0;
	wire [1:0] w_n11824_0;
	wire [1:0] w_n11825_0;
	wire [2:0] w_n11826_0;
	wire [1:0] w_n11827_0;
	wire [1:0] w_n11830_0;
	wire [1:0] w_n11836_0;
	wire [1:0] w_n11837_0;
	wire [1:0] w_n11839_0;
	wire [1:0] w_n11841_0;
	wire [1:0] w_n11843_0;
	wire [1:0] w_n11849_0;
	wire [1:0] w_n11851_0;
	wire [2:0] w_n11852_0;
	wire [1:0] w_n11855_0;
	wire [1:0] w_n11856_0;
	wire [2:0] w_n11857_0;
	wire [1:0] w_n11859_0;
	wire [1:0] w_n11863_0;
	wire [1:0] w_n11865_0;
	wire [1:0] w_n11866_0;
	wire [2:0] w_n11867_0;
	wire [1:0] w_n11868_0;
	wire [1:0] w_n11871_0;
	wire [1:0] w_n11877_0;
	wire [1:0] w_n11878_0;
	wire [1:0] w_n11880_0;
	wire [1:0] w_n11882_0;
	wire [1:0] w_n11884_0;
	wire [1:0] w_n11890_0;
	wire [1:0] w_n11892_0;
	wire [2:0] w_n11893_0;
	wire [1:0] w_n11896_0;
	wire [1:0] w_n11897_0;
	wire [2:0] w_n11898_0;
	wire [1:0] w_n11900_0;
	wire [1:0] w_n11904_0;
	wire [1:0] w_n11906_0;
	wire [1:0] w_n11907_0;
	wire [2:0] w_n11908_0;
	wire [1:0] w_n11909_0;
	wire [1:0] w_n11912_0;
	wire [1:0] w_n11918_0;
	wire [1:0] w_n11919_0;
	wire [1:0] w_n11921_0;
	wire [1:0] w_n11923_0;
	wire [1:0] w_n11925_0;
	wire [1:0] w_n11931_0;
	wire [1:0] w_n11933_0;
	wire [2:0] w_n11934_0;
	wire [1:0] w_n11937_0;
	wire [1:0] w_n11938_0;
	wire [2:0] w_n11939_0;
	wire [1:0] w_n11941_0;
	wire [1:0] w_n11943_0;
	wire [1:0] w_n11945_0;
	wire [1:0] w_n11951_0;
	wire [2:0] w_n11953_0;
	wire [1:0] w_n11954_0;
	wire [1:0] w_n11957_0;
	wire [1:0] w_n11959_0;
	wire [1:0] w_n11963_0;
	wire [1:0] w_n11965_0;
	wire [1:0] w_n11966_0;
	wire [1:0] w_n11967_0;
	wire [2:0] w_n11968_0;
	wire [1:0] w_n11971_0;
	wire [1:0] w_n11972_0;
	wire [2:0] w_n11973_0;
	wire [1:0] w_n11975_0;
	wire [1:0] w_n11979_0;
	wire [1:0] w_n11981_0;
	wire [1:0] w_n11982_0;
	wire [2:0] w_n11983_0;
	wire [1:0] w_n11984_0;
	wire [1:0] w_n11987_0;
	wire [1:0] w_n11993_0;
	wire [1:0] w_n11994_0;
	wire [1:0] w_n11996_0;
	wire [1:0] w_n11998_0;
	wire [1:0] w_n12000_0;
	wire [1:0] w_n12006_0;
	wire [1:0] w_n12008_0;
	wire [2:0] w_n12009_0;
	wire [1:0] w_n12012_0;
	wire [1:0] w_n12013_0;
	wire [2:0] w_n12014_0;
	wire [1:0] w_n12016_0;
	wire [1:0] w_n12020_0;
	wire [1:0] w_n12022_0;
	wire [1:0] w_n12023_0;
	wire [2:0] w_n12024_0;
	wire [1:0] w_n12025_0;
	wire [1:0] w_n12028_0;
	wire [1:0] w_n12034_0;
	wire [1:0] w_n12035_0;
	wire [1:0] w_n12037_0;
	wire [1:0] w_n12039_0;
	wire [1:0] w_n12041_0;
	wire [1:0] w_n12047_0;
	wire [1:0] w_n12049_0;
	wire [2:0] w_n12050_0;
	wire [1:0] w_n12053_0;
	wire [1:0] w_n12054_0;
	wire [2:0] w_n12055_0;
	wire [1:0] w_n12057_0;
	wire [1:0] w_n12061_0;
	wire [1:0] w_n12063_0;
	wire [1:0] w_n12064_0;
	wire [2:0] w_n12065_0;
	wire [1:0] w_n12066_0;
	wire [1:0] w_n12069_0;
	wire [1:0] w_n12075_0;
	wire [1:0] w_n12076_0;
	wire [1:0] w_n12078_0;
	wire [1:0] w_n12080_0;
	wire [1:0] w_n12082_0;
	wire [1:0] w_n12088_0;
	wire [1:0] w_n12090_0;
	wire [2:0] w_n12091_0;
	wire [1:0] w_n12094_0;
	wire [1:0] w_n12095_0;
	wire [2:0] w_n12096_0;
	wire [1:0] w_n12098_0;
	wire [1:0] w_n12102_0;
	wire [1:0] w_n12104_0;
	wire [1:0] w_n12105_0;
	wire [2:0] w_n12106_0;
	wire [1:0] w_n12110_0;
	wire [1:0] w_n12116_0;
	wire [2:0] w_n12118_0;
	wire [1:0] w_n12120_0;
	wire [2:0] w_n12125_0;
	wire [1:0] w_n12126_0;
	wire [1:0] w_n12127_0;
	wire [1:0] w_n12132_0;
	wire [2:0] w_n12133_0;
	wire [1:0] w_n12138_0;
	wire [1:0] w_n12145_0;
	wire [2:0] w_n12148_0;
	wire [1:0] w_n12148_1;
	wire [1:0] w_n12149_0;
	wire [2:0] w_n12152_0;
	wire [1:0] w_n12153_0;
	wire [1:0] w_n12154_0;
	wire [1:0] w_n12155_0;
	wire [1:0] w_n12157_0;
	wire [1:0] w_n12159_0;
	wire [1:0] w_n12161_0;
	wire [1:0] w_n12170_0;
	wire [2:0] w_n12172_0;
	wire [1:0] w_n12173_0;
	wire [1:0] w_n12177_0;
	wire [1:0] w_n12179_0;
	wire [1:0] w_n12181_0;
	wire [1:0] w_n12186_0;
	wire [1:0] w_n12188_0;
	wire [1:0] w_n12189_0;
	wire [2:0] w_n12190_0;
	wire [1:0] w_n12191_0;
	wire [1:0] w_n12196_0;
	wire [1:0] w_n12197_0;
	wire [1:0] w_n12199_0;
	wire [1:0] w_n12201_0;
	wire [1:0] w_n12204_0;
	wire [1:0] w_n12210_0;
	wire [2:0] w_n12212_0;
	wire [1:0] w_n12213_0;
	wire [1:0] w_n12217_0;
	wire [1:0] w_n12218_0;
	wire [1:0] w_n12220_0;
	wire [1:0] w_n12225_0;
	wire [1:0] w_n12227_0;
	wire [1:0] w_n12228_0;
	wire [2:0] w_n12229_0;
	wire [1:0] w_n12230_0;
	wire [1:0] w_n12234_0;
	wire [1:0] w_n12235_0;
	wire [1:0] w_n12237_0;
	wire [1:0] w_n12239_0;
	wire [1:0] w_n12242_0;
	wire [1:0] w_n12248_0;
	wire [1:0] w_n12250_0;
	wire [2:0] w_n12251_0;
	wire [1:0] w_n12255_0;
	wire [1:0] w_n12256_0;
	wire [2:0] w_n12257_0;
	wire [1:0] w_n12259_0;
	wire [1:0] w_n12264_0;
	wire [1:0] w_n12266_0;
	wire [1:0] w_n12267_0;
	wire [2:0] w_n12268_0;
	wire [1:0] w_n12269_0;
	wire [1:0] w_n12273_0;
	wire [1:0] w_n12279_0;
	wire [1:0] w_n12280_0;
	wire [1:0] w_n12282_0;
	wire [1:0] w_n12284_0;
	wire [1:0] w_n12287_0;
	wire [1:0] w_n12293_0;
	wire [1:0] w_n12295_0;
	wire [2:0] w_n12296_0;
	wire [1:0] w_n12300_0;
	wire [1:0] w_n12301_0;
	wire [2:0] w_n12302_0;
	wire [1:0] w_n12304_0;
	wire [1:0] w_n12309_0;
	wire [1:0] w_n12311_0;
	wire [1:0] w_n12312_0;
	wire [2:0] w_n12313_0;
	wire [1:0] w_n12314_0;
	wire [1:0] w_n12318_0;
	wire [1:0] w_n12324_0;
	wire [1:0] w_n12325_0;
	wire [1:0] w_n12327_0;
	wire [1:0] w_n12329_0;
	wire [1:0] w_n12332_0;
	wire [1:0] w_n12338_0;
	wire [1:0] w_n12340_0;
	wire [2:0] w_n12341_0;
	wire [1:0] w_n12345_0;
	wire [1:0] w_n12346_0;
	wire [2:0] w_n12347_0;
	wire [1:0] w_n12349_0;
	wire [1:0] w_n12354_0;
	wire [1:0] w_n12356_0;
	wire [1:0] w_n12357_0;
	wire [2:0] w_n12358_0;
	wire [1:0] w_n12359_0;
	wire [1:0] w_n12363_0;
	wire [1:0] w_n12369_0;
	wire [1:0] w_n12370_0;
	wire [1:0] w_n12372_0;
	wire [1:0] w_n12374_0;
	wire [1:0] w_n12377_0;
	wire [1:0] w_n12383_0;
	wire [1:0] w_n12385_0;
	wire [2:0] w_n12386_0;
	wire [1:0] w_n12390_0;
	wire [1:0] w_n12391_0;
	wire [2:0] w_n12392_0;
	wire [1:0] w_n12394_0;
	wire [1:0] w_n12399_0;
	wire [1:0] w_n12401_0;
	wire [1:0] w_n12402_0;
	wire [2:0] w_n12403_0;
	wire [1:0] w_n12404_0;
	wire [1:0] w_n12408_0;
	wire [1:0] w_n12414_0;
	wire [1:0] w_n12415_0;
	wire [1:0] w_n12417_0;
	wire [1:0] w_n12419_0;
	wire [1:0] w_n12422_0;
	wire [1:0] w_n12428_0;
	wire [1:0] w_n12430_0;
	wire [2:0] w_n12431_0;
	wire [1:0] w_n12435_0;
	wire [1:0] w_n12436_0;
	wire [2:0] w_n12437_0;
	wire [1:0] w_n12439_0;
	wire [1:0] w_n12444_0;
	wire [1:0] w_n12446_0;
	wire [1:0] w_n12447_0;
	wire [2:0] w_n12448_0;
	wire [1:0] w_n12449_0;
	wire [1:0] w_n12453_0;
	wire [1:0] w_n12459_0;
	wire [1:0] w_n12460_0;
	wire [1:0] w_n12462_0;
	wire [1:0] w_n12467_0;
	wire [1:0] w_n12469_0;
	wire [1:0] w_n12470_0;
	wire [2:0] w_n12471_0;
	wire [1:0] w_n12472_0;
	wire [1:0] w_n12474_0;
	wire [1:0] w_n12476_0;
	wire [1:0] w_n12478_0;
	wire [1:0] w_n12481_0;
	wire [1:0] w_n12487_0;
	wire [2:0] w_n12489_0;
	wire [1:0] w_n12490_0;
	wire [1:0] w_n12494_0;
	wire [1:0] w_n12500_0;
	wire [1:0] w_n12501_0;
	wire [1:0] w_n12503_0;
	wire [1:0] w_n12505_0;
	wire [1:0] w_n12508_0;
	wire [1:0] w_n12514_0;
	wire [1:0] w_n12516_0;
	wire [2:0] w_n12517_0;
	wire [1:0] w_n12521_0;
	wire [1:0] w_n12522_0;
	wire [2:0] w_n12523_0;
	wire [1:0] w_n12525_0;
	wire [1:0] w_n12530_0;
	wire [1:0] w_n12532_0;
	wire [1:0] w_n12533_0;
	wire [2:0] w_n12534_0;
	wire [1:0] w_n12535_0;
	wire [1:0] w_n12539_0;
	wire [1:0] w_n12545_0;
	wire [1:0] w_n12546_0;
	wire [1:0] w_n12548_0;
	wire [1:0] w_n12550_0;
	wire [1:0] w_n12553_0;
	wire [1:0] w_n12559_0;
	wire [1:0] w_n12561_0;
	wire [2:0] w_n12562_0;
	wire [1:0] w_n12566_0;
	wire [1:0] w_n12567_0;
	wire [2:0] w_n12568_0;
	wire [1:0] w_n12570_0;
	wire [1:0] w_n12575_0;
	wire [1:0] w_n12577_0;
	wire [1:0] w_n12578_0;
	wire [2:0] w_n12579_0;
	wire [1:0] w_n12580_0;
	wire [1:0] w_n12584_0;
	wire [1:0] w_n12590_0;
	wire [1:0] w_n12591_0;
	wire [1:0] w_n12593_0;
	wire [1:0] w_n12595_0;
	wire [1:0] w_n12598_0;
	wire [1:0] w_n12604_0;
	wire [1:0] w_n12606_0;
	wire [2:0] w_n12607_0;
	wire [1:0] w_n12611_0;
	wire [1:0] w_n12612_0;
	wire [2:0] w_n12613_0;
	wire [1:0] w_n12615_0;
	wire [1:0] w_n12620_0;
	wire [1:0] w_n12622_0;
	wire [1:0] w_n12623_0;
	wire [2:0] w_n12624_0;
	wire [1:0] w_n12625_0;
	wire [1:0] w_n12629_0;
	wire [1:0] w_n12635_0;
	wire [1:0] w_n12636_0;
	wire [1:0] w_n12638_0;
	wire [1:0] w_n12640_0;
	wire [1:0] w_n12643_0;
	wire [1:0] w_n12649_0;
	wire [2:0] w_n12651_0;
	wire [2:0] w_n12651_1;
	wire [1:0] w_n12654_0;
	wire [2:0] w_n12655_0;
	wire [1:0] w_n12656_0;
	wire [1:0] w_n12662_0;
	wire [2:0] w_n12663_0;
	wire [1:0] w_n12664_0;
	wire [1:0] w_n12669_0;
	wire [2:0] w_n12670_0;
	wire [2:0] w_n12670_1;
	wire [2:0] w_n12670_2;
	wire [2:0] w_n12670_3;
	wire [2:0] w_n12670_4;
	wire [2:0] w_n12670_5;
	wire [2:0] w_n12670_6;
	wire [2:0] w_n12670_7;
	wire [2:0] w_n12670_8;
	wire [2:0] w_n12670_9;
	wire [2:0] w_n12670_10;
	wire [2:0] w_n12675_0;
	wire [2:0] w_n12675_1;
	wire [2:0] w_n12675_2;
	wire [2:0] w_n12675_3;
	wire [2:0] w_n12675_4;
	wire [2:0] w_n12675_5;
	wire [2:0] w_n12675_6;
	wire [2:0] w_n12675_7;
	wire [2:0] w_n12675_8;
	wire [2:0] w_n12675_9;
	wire [2:0] w_n12675_10;
	wire [2:0] w_n12675_11;
	wire [2:0] w_n12675_12;
	wire [2:0] w_n12675_13;
	wire [2:0] w_n12675_14;
	wire [2:0] w_n12675_15;
	wire [2:0] w_n12675_16;
	wire [2:0] w_n12675_17;
	wire [2:0] w_n12675_18;
	wire [2:0] w_n12675_19;
	wire [2:0] w_n12675_20;
	wire [2:0] w_n12675_21;
	wire [2:0] w_n12675_22;
	wire [2:0] w_n12675_23;
	wire [1:0] w_n12675_24;
	wire [1:0] w_n12679_0;
	wire [2:0] w_n12681_0;
	wire [1:0] w_n12681_1;
	wire [2:0] w_n12682_0;
	wire [2:0] w_n12686_0;
	wire [1:0] w_n12687_0;
	wire [1:0] w_n12688_0;
	wire [1:0] w_n12689_0;
	wire [1:0] w_n12691_0;
	wire [1:0] w_n12693_0;
	wire [1:0] w_n12695_0;
	wire [1:0] w_n12698_0;
	wire [1:0] w_n12703_0;
	wire [2:0] w_n12705_0;
	wire [1:0] w_n12706_0;
	wire [1:0] w_n12710_0;
	wire [1:0] w_n12711_0;
	wire [1:0] w_n12713_0;
	wire [1:0] w_n12717_0;
	wire [1:0] w_n12719_0;
	wire [1:0] w_n12720_0;
	wire [2:0] w_n12721_0;
	wire [1:0] w_n12722_0;
	wire [1:0] w_n12726_0;
	wire [1:0] w_n12728_0;
	wire [1:0] w_n12730_0;
	wire [1:0] w_n12732_0;
	wire [1:0] w_n12735_0;
	wire [1:0] w_n12741_0;
	wire [2:0] w_n12743_0;
	wire [1:0] w_n12744_0;
	wire [1:0] w_n12749_0;
	wire [1:0] w_n12751_0;
	wire [1:0] w_n12753_0;
	wire [1:0] w_n12757_0;
	wire [1:0] w_n12759_0;
	wire [1:0] w_n12760_0;
	wire [2:0] w_n12761_0;
	wire [1:0] w_n12762_0;
	wire [1:0] w_n12768_0;
	wire [1:0] w_n12769_0;
	wire [1:0] w_n12771_0;
	wire [1:0] w_n12773_0;
	wire [1:0] w_n12775_0;
	wire [1:0] w_n12781_0;
	wire [1:0] w_n12783_0;
	wire [2:0] w_n12784_0;
	wire [1:0] w_n12787_0;
	wire [1:0] w_n12788_0;
	wire [2:0] w_n12789_0;
	wire [1:0] w_n12791_0;
	wire [1:0] w_n12795_0;
	wire [1:0] w_n12797_0;
	wire [1:0] w_n12798_0;
	wire [2:0] w_n12799_0;
	wire [1:0] w_n12800_0;
	wire [1:0] w_n12803_0;
	wire [1:0] w_n12809_0;
	wire [1:0] w_n12810_0;
	wire [1:0] w_n12812_0;
	wire [1:0] w_n12814_0;
	wire [1:0] w_n12816_0;
	wire [1:0] w_n12822_0;
	wire [1:0] w_n12824_0;
	wire [2:0] w_n12825_0;
	wire [1:0] w_n12828_0;
	wire [1:0] w_n12829_0;
	wire [2:0] w_n12830_0;
	wire [1:0] w_n12832_0;
	wire [1:0] w_n12836_0;
	wire [1:0] w_n12838_0;
	wire [1:0] w_n12839_0;
	wire [2:0] w_n12840_0;
	wire [1:0] w_n12841_0;
	wire [1:0] w_n12844_0;
	wire [1:0] w_n12850_0;
	wire [1:0] w_n12851_0;
	wire [1:0] w_n12853_0;
	wire [1:0] w_n12855_0;
	wire [1:0] w_n12857_0;
	wire [1:0] w_n12863_0;
	wire [1:0] w_n12865_0;
	wire [2:0] w_n12866_0;
	wire [1:0] w_n12869_0;
	wire [1:0] w_n12870_0;
	wire [2:0] w_n12871_0;
	wire [1:0] w_n12873_0;
	wire [1:0] w_n12877_0;
	wire [1:0] w_n12879_0;
	wire [1:0] w_n12880_0;
	wire [2:0] w_n12881_0;
	wire [1:0] w_n12882_0;
	wire [1:0] w_n12885_0;
	wire [1:0] w_n12891_0;
	wire [1:0] w_n12892_0;
	wire [1:0] w_n12894_0;
	wire [1:0] w_n12896_0;
	wire [1:0] w_n12898_0;
	wire [1:0] w_n12904_0;
	wire [1:0] w_n12906_0;
	wire [2:0] w_n12907_0;
	wire [1:0] w_n12910_0;
	wire [1:0] w_n12911_0;
	wire [2:0] w_n12912_0;
	wire [1:0] w_n12914_0;
	wire [1:0] w_n12918_0;
	wire [1:0] w_n12920_0;
	wire [1:0] w_n12921_0;
	wire [2:0] w_n12922_0;
	wire [1:0] w_n12923_0;
	wire [1:0] w_n12926_0;
	wire [1:0] w_n12932_0;
	wire [1:0] w_n12933_0;
	wire [1:0] w_n12935_0;
	wire [1:0] w_n12937_0;
	wire [1:0] w_n12939_0;
	wire [1:0] w_n12945_0;
	wire [1:0] w_n12947_0;
	wire [2:0] w_n12948_0;
	wire [1:0] w_n12951_0;
	wire [1:0] w_n12952_0;
	wire [2:0] w_n12953_0;
	wire [1:0] w_n12955_0;
	wire [1:0] w_n12959_0;
	wire [1:0] w_n12961_0;
	wire [1:0] w_n12962_0;
	wire [2:0] w_n12963_0;
	wire [1:0] w_n12964_0;
	wire [1:0] w_n12967_0;
	wire [1:0] w_n12973_0;
	wire [1:0] w_n12974_0;
	wire [1:0] w_n12976_0;
	wire [1:0] w_n12978_0;
	wire [1:0] w_n12980_0;
	wire [1:0] w_n12986_0;
	wire [1:0] w_n12988_0;
	wire [2:0] w_n12989_0;
	wire [1:0] w_n12992_0;
	wire [1:0] w_n12993_0;
	wire [2:0] w_n12994_0;
	wire [1:0] w_n12996_0;
	wire [1:0] w_n12998_0;
	wire [1:0] w_n13000_0;
	wire [1:0] w_n13006_0;
	wire [2:0] w_n13008_0;
	wire [1:0] w_n13009_0;
	wire [1:0] w_n13011_0;
	wire [1:0] w_n13013_0;
	wire [1:0] w_n13017_0;
	wire [1:0] w_n13019_0;
	wire [1:0] w_n13020_0;
	wire [1:0] w_n13021_0;
	wire [2:0] w_n13022_0;
	wire [1:0] w_n13025_0;
	wire [1:0] w_n13026_0;
	wire [2:0] w_n13027_0;
	wire [1:0] w_n13029_0;
	wire [1:0] w_n13033_0;
	wire [1:0] w_n13035_0;
	wire [1:0] w_n13036_0;
	wire [2:0] w_n13037_0;
	wire [1:0] w_n13038_0;
	wire [1:0] w_n13041_0;
	wire [1:0] w_n13047_0;
	wire [1:0] w_n13048_0;
	wire [1:0] w_n13050_0;
	wire [1:0] w_n13052_0;
	wire [1:0] w_n13054_0;
	wire [1:0] w_n13060_0;
	wire [1:0] w_n13062_0;
	wire [2:0] w_n13063_0;
	wire [1:0] w_n13066_0;
	wire [1:0] w_n13067_0;
	wire [2:0] w_n13068_0;
	wire [1:0] w_n13070_0;
	wire [1:0] w_n13074_0;
	wire [1:0] w_n13076_0;
	wire [1:0] w_n13077_0;
	wire [2:0] w_n13078_0;
	wire [1:0] w_n13079_0;
	wire [1:0] w_n13082_0;
	wire [1:0] w_n13088_0;
	wire [1:0] w_n13089_0;
	wire [1:0] w_n13091_0;
	wire [1:0] w_n13093_0;
	wire [1:0] w_n13095_0;
	wire [1:0] w_n13101_0;
	wire [1:0] w_n13103_0;
	wire [2:0] w_n13104_0;
	wire [1:0] w_n13107_0;
	wire [1:0] w_n13108_0;
	wire [2:0] w_n13109_0;
	wire [1:0] w_n13111_0;
	wire [1:0] w_n13115_0;
	wire [1:0] w_n13117_0;
	wire [1:0] w_n13118_0;
	wire [2:0] w_n13119_0;
	wire [1:0] w_n13120_0;
	wire [1:0] w_n13123_0;
	wire [1:0] w_n13129_0;
	wire [1:0] w_n13130_0;
	wire [1:0] w_n13132_0;
	wire [1:0] w_n13134_0;
	wire [1:0] w_n13136_0;
	wire [1:0] w_n13142_0;
	wire [2:0] w_n13144_0;
	wire [1:0] w_n13149_0;
	wire [2:0] w_n13151_0;
	wire [2:0] w_n13155_0;
	wire [1:0] w_n13156_0;
	wire [1:0] w_n13161_0;
	wire [2:0] w_n13162_0;
	wire [1:0] w_n13167_0;
	wire [1:0] w_n13175_0;
	wire [2:0] w_n13177_0;
	wire [1:0] w_n13177_1;
	wire [1:0] w_n13178_0;
	wire [2:0] w_n13181_0;
	wire [1:0] w_n13182_0;
	wire [1:0] w_n13183_0;
	wire [1:0] w_n13184_0;
	wire [1:0] w_n13186_0;
	wire [1:0] w_n13188_0;
	wire [1:0] w_n13190_0;
	wire [1:0] w_n13199_0;
	wire [2:0] w_n13201_0;
	wire [1:0] w_n13202_0;
	wire [1:0] w_n13206_0;
	wire [1:0] w_n13208_0;
	wire [1:0] w_n13210_0;
	wire [1:0] w_n13215_0;
	wire [1:0] w_n13217_0;
	wire [1:0] w_n13218_0;
	wire [2:0] w_n13219_0;
	wire [1:0] w_n13220_0;
	wire [1:0] w_n13225_0;
	wire [1:0] w_n13226_0;
	wire [1:0] w_n13228_0;
	wire [1:0] w_n13230_0;
	wire [1:0] w_n13233_0;
	wire [1:0] w_n13239_0;
	wire [2:0] w_n13241_0;
	wire [1:0] w_n13242_0;
	wire [1:0] w_n13246_0;
	wire [1:0] w_n13247_0;
	wire [1:0] w_n13249_0;
	wire [1:0] w_n13254_0;
	wire [1:0] w_n13256_0;
	wire [1:0] w_n13257_0;
	wire [2:0] w_n13258_0;
	wire [1:0] w_n13259_0;
	wire [1:0] w_n13263_0;
	wire [1:0] w_n13264_0;
	wire [1:0] w_n13266_0;
	wire [1:0] w_n13268_0;
	wire [1:0] w_n13271_0;
	wire [1:0] w_n13277_0;
	wire [1:0] w_n13279_0;
	wire [2:0] w_n13280_0;
	wire [1:0] w_n13284_0;
	wire [1:0] w_n13285_0;
	wire [2:0] w_n13286_0;
	wire [1:0] w_n13288_0;
	wire [1:0] w_n13293_0;
	wire [1:0] w_n13295_0;
	wire [1:0] w_n13296_0;
	wire [2:0] w_n13297_0;
	wire [1:0] w_n13298_0;
	wire [1:0] w_n13302_0;
	wire [1:0] w_n13308_0;
	wire [1:0] w_n13309_0;
	wire [1:0] w_n13311_0;
	wire [1:0] w_n13313_0;
	wire [1:0] w_n13316_0;
	wire [1:0] w_n13322_0;
	wire [1:0] w_n13324_0;
	wire [2:0] w_n13325_0;
	wire [1:0] w_n13329_0;
	wire [1:0] w_n13330_0;
	wire [2:0] w_n13331_0;
	wire [1:0] w_n13333_0;
	wire [1:0] w_n13338_0;
	wire [1:0] w_n13340_0;
	wire [1:0] w_n13341_0;
	wire [2:0] w_n13342_0;
	wire [1:0] w_n13343_0;
	wire [1:0] w_n13347_0;
	wire [1:0] w_n13353_0;
	wire [1:0] w_n13354_0;
	wire [1:0] w_n13356_0;
	wire [1:0] w_n13358_0;
	wire [1:0] w_n13361_0;
	wire [1:0] w_n13367_0;
	wire [1:0] w_n13369_0;
	wire [2:0] w_n13370_0;
	wire [1:0] w_n13374_0;
	wire [1:0] w_n13375_0;
	wire [2:0] w_n13376_0;
	wire [1:0] w_n13378_0;
	wire [1:0] w_n13383_0;
	wire [1:0] w_n13385_0;
	wire [1:0] w_n13386_0;
	wire [2:0] w_n13387_0;
	wire [1:0] w_n13388_0;
	wire [1:0] w_n13392_0;
	wire [1:0] w_n13398_0;
	wire [1:0] w_n13399_0;
	wire [1:0] w_n13401_0;
	wire [1:0] w_n13403_0;
	wire [1:0] w_n13406_0;
	wire [1:0] w_n13412_0;
	wire [1:0] w_n13414_0;
	wire [2:0] w_n13415_0;
	wire [1:0] w_n13419_0;
	wire [1:0] w_n13420_0;
	wire [2:0] w_n13421_0;
	wire [1:0] w_n13423_0;
	wire [1:0] w_n13428_0;
	wire [1:0] w_n13430_0;
	wire [1:0] w_n13431_0;
	wire [2:0] w_n13432_0;
	wire [1:0] w_n13433_0;
	wire [1:0] w_n13437_0;
	wire [1:0] w_n13443_0;
	wire [1:0] w_n13444_0;
	wire [1:0] w_n13446_0;
	wire [1:0] w_n13448_0;
	wire [1:0] w_n13451_0;
	wire [1:0] w_n13457_0;
	wire [1:0] w_n13459_0;
	wire [2:0] w_n13460_0;
	wire [1:0] w_n13464_0;
	wire [1:0] w_n13465_0;
	wire [2:0] w_n13466_0;
	wire [1:0] w_n13468_0;
	wire [1:0] w_n13473_0;
	wire [1:0] w_n13475_0;
	wire [1:0] w_n13476_0;
	wire [2:0] w_n13477_0;
	wire [1:0] w_n13478_0;
	wire [1:0] w_n13482_0;
	wire [1:0] w_n13488_0;
	wire [1:0] w_n13489_0;
	wire [1:0] w_n13491_0;
	wire [1:0] w_n13493_0;
	wire [1:0] w_n13496_0;
	wire [1:0] w_n13502_0;
	wire [1:0] w_n13504_0;
	wire [2:0] w_n13505_0;
	wire [1:0] w_n13509_0;
	wire [1:0] w_n13510_0;
	wire [2:0] w_n13511_0;
	wire [1:0] w_n13513_0;
	wire [1:0] w_n13518_0;
	wire [1:0] w_n13520_0;
	wire [1:0] w_n13521_0;
	wire [2:0] w_n13522_0;
	wire [1:0] w_n13523_0;
	wire [1:0] w_n13527_0;
	wire [1:0] w_n13533_0;
	wire [1:0] w_n13534_0;
	wire [1:0] w_n13536_0;
	wire [1:0] w_n13541_0;
	wire [1:0] w_n13543_0;
	wire [1:0] w_n13544_0;
	wire [2:0] w_n13545_0;
	wire [1:0] w_n13546_0;
	wire [1:0] w_n13548_0;
	wire [1:0] w_n13550_0;
	wire [1:0] w_n13552_0;
	wire [1:0] w_n13555_0;
	wire [1:0] w_n13561_0;
	wire [2:0] w_n13563_0;
	wire [1:0] w_n13564_0;
	wire [1:0] w_n13568_0;
	wire [1:0] w_n13574_0;
	wire [1:0] w_n13575_0;
	wire [1:0] w_n13577_0;
	wire [1:0] w_n13579_0;
	wire [1:0] w_n13582_0;
	wire [1:0] w_n13588_0;
	wire [1:0] w_n13590_0;
	wire [2:0] w_n13591_0;
	wire [1:0] w_n13595_0;
	wire [1:0] w_n13596_0;
	wire [2:0] w_n13597_0;
	wire [1:0] w_n13599_0;
	wire [1:0] w_n13604_0;
	wire [1:0] w_n13606_0;
	wire [1:0] w_n13607_0;
	wire [2:0] w_n13608_0;
	wire [1:0] w_n13609_0;
	wire [1:0] w_n13613_0;
	wire [1:0] w_n13619_0;
	wire [1:0] w_n13620_0;
	wire [1:0] w_n13622_0;
	wire [1:0] w_n13624_0;
	wire [1:0] w_n13627_0;
	wire [1:0] w_n13633_0;
	wire [1:0] w_n13635_0;
	wire [2:0] w_n13636_0;
	wire [1:0] w_n13640_0;
	wire [1:0] w_n13641_0;
	wire [2:0] w_n13642_0;
	wire [1:0] w_n13644_0;
	wire [1:0] w_n13649_0;
	wire [1:0] w_n13651_0;
	wire [1:0] w_n13652_0;
	wire [2:0] w_n13653_0;
	wire [1:0] w_n13654_0;
	wire [1:0] w_n13658_0;
	wire [1:0] w_n13664_0;
	wire [1:0] w_n13665_0;
	wire [1:0] w_n13667_0;
	wire [1:0] w_n13669_0;
	wire [1:0] w_n13672_0;
	wire [1:0] w_n13678_0;
	wire [1:0] w_n13680_0;
	wire [2:0] w_n13681_0;
	wire [1:0] w_n13685_0;
	wire [1:0] w_n13686_0;
	wire [2:0] w_n13687_0;
	wire [1:0] w_n13689_0;
	wire [1:0] w_n13694_0;
	wire [1:0] w_n13696_0;
	wire [1:0] w_n13697_0;
	wire [2:0] w_n13698_0;
	wire [2:0] w_n13698_1;
	wire [1:0] w_n13701_0;
	wire [2:0] w_n13702_0;
	wire [1:0] w_n13703_0;
	wire [1:0] w_n13704_0;
	wire [1:0] w_n13710_0;
	wire [2:0] w_n13711_0;
	wire [1:0] w_n13712_0;
	wire [1:0] w_n13717_0;
	wire [2:0] w_n13718_0;
	wire [2:0] w_n13718_1;
	wire [2:0] w_n13718_2;
	wire [2:0] w_n13718_3;
	wire [2:0] w_n13718_4;
	wire [2:0] w_n13718_5;
	wire [2:0] w_n13718_6;
	wire [2:0] w_n13718_7;
	wire [2:0] w_n13718_8;
	wire [1:0] w_n13718_9;
	wire [2:0] w_n13723_0;
	wire [2:0] w_n13723_1;
	wire [2:0] w_n13723_2;
	wire [2:0] w_n13723_3;
	wire [2:0] w_n13723_4;
	wire [2:0] w_n13723_5;
	wire [2:0] w_n13723_6;
	wire [2:0] w_n13723_7;
	wire [2:0] w_n13723_8;
	wire [2:0] w_n13723_9;
	wire [2:0] w_n13723_10;
	wire [2:0] w_n13723_11;
	wire [2:0] w_n13723_12;
	wire [2:0] w_n13723_13;
	wire [2:0] w_n13723_14;
	wire [2:0] w_n13723_15;
	wire [2:0] w_n13723_16;
	wire [2:0] w_n13723_17;
	wire [2:0] w_n13723_18;
	wire [2:0] w_n13723_19;
	wire [2:0] w_n13723_20;
	wire [2:0] w_n13723_21;
	wire [2:0] w_n13723_22;
	wire [1:0] w_n13726_0;
	wire [2:0] w_n13728_0;
	wire [1:0] w_n13728_1;
	wire [2:0] w_n13729_0;
	wire [2:0] w_n13733_0;
	wire [1:0] w_n13734_0;
	wire [1:0] w_n13735_0;
	wire [1:0] w_n13736_0;
	wire [1:0] w_n13738_0;
	wire [1:0] w_n13740_0;
	wire [1:0] w_n13742_0;
	wire [1:0] w_n13745_0;
	wire [1:0] w_n13750_0;
	wire [2:0] w_n13752_0;
	wire [1:0] w_n13753_0;
	wire [1:0] w_n13757_0;
	wire [1:0] w_n13758_0;
	wire [1:0] w_n13760_0;
	wire [1:0] w_n13764_0;
	wire [1:0] w_n13766_0;
	wire [1:0] w_n13767_0;
	wire [2:0] w_n13768_0;
	wire [1:0] w_n13769_0;
	wire [1:0] w_n13773_0;
	wire [1:0] w_n13775_0;
	wire [1:0] w_n13777_0;
	wire [1:0] w_n13779_0;
	wire [1:0] w_n13782_0;
	wire [1:0] w_n13788_0;
	wire [2:0] w_n13790_0;
	wire [1:0] w_n13791_0;
	wire [1:0] w_n13796_0;
	wire [1:0] w_n13798_0;
	wire [1:0] w_n13800_0;
	wire [1:0] w_n13804_0;
	wire [1:0] w_n13806_0;
	wire [1:0] w_n13807_0;
	wire [2:0] w_n13808_0;
	wire [1:0] w_n13809_0;
	wire [1:0] w_n13815_0;
	wire [1:0] w_n13816_0;
	wire [1:0] w_n13818_0;
	wire [1:0] w_n13820_0;
	wire [1:0] w_n13822_0;
	wire [1:0] w_n13828_0;
	wire [1:0] w_n13830_0;
	wire [2:0] w_n13831_0;
	wire [1:0] w_n13834_0;
	wire [1:0] w_n13835_0;
	wire [2:0] w_n13836_0;
	wire [1:0] w_n13838_0;
	wire [1:0] w_n13842_0;
	wire [1:0] w_n13844_0;
	wire [1:0] w_n13845_0;
	wire [2:0] w_n13846_0;
	wire [1:0] w_n13847_0;
	wire [1:0] w_n13850_0;
	wire [1:0] w_n13856_0;
	wire [1:0] w_n13857_0;
	wire [1:0] w_n13859_0;
	wire [1:0] w_n13861_0;
	wire [1:0] w_n13863_0;
	wire [1:0] w_n13869_0;
	wire [1:0] w_n13871_0;
	wire [2:0] w_n13872_0;
	wire [1:0] w_n13875_0;
	wire [1:0] w_n13876_0;
	wire [2:0] w_n13877_0;
	wire [1:0] w_n13879_0;
	wire [1:0] w_n13883_0;
	wire [1:0] w_n13885_0;
	wire [1:0] w_n13886_0;
	wire [2:0] w_n13887_0;
	wire [1:0] w_n13888_0;
	wire [1:0] w_n13891_0;
	wire [1:0] w_n13897_0;
	wire [1:0] w_n13898_0;
	wire [1:0] w_n13900_0;
	wire [1:0] w_n13902_0;
	wire [1:0] w_n13904_0;
	wire [1:0] w_n13910_0;
	wire [1:0] w_n13912_0;
	wire [2:0] w_n13913_0;
	wire [1:0] w_n13916_0;
	wire [1:0] w_n13917_0;
	wire [2:0] w_n13918_0;
	wire [1:0] w_n13920_0;
	wire [1:0] w_n13924_0;
	wire [1:0] w_n13926_0;
	wire [1:0] w_n13927_0;
	wire [2:0] w_n13928_0;
	wire [1:0] w_n13929_0;
	wire [1:0] w_n13932_0;
	wire [1:0] w_n13938_0;
	wire [1:0] w_n13939_0;
	wire [1:0] w_n13941_0;
	wire [1:0] w_n13943_0;
	wire [1:0] w_n13945_0;
	wire [1:0] w_n13951_0;
	wire [1:0] w_n13953_0;
	wire [2:0] w_n13954_0;
	wire [1:0] w_n13957_0;
	wire [1:0] w_n13958_0;
	wire [2:0] w_n13959_0;
	wire [1:0] w_n13961_0;
	wire [1:0] w_n13965_0;
	wire [1:0] w_n13967_0;
	wire [1:0] w_n13968_0;
	wire [2:0] w_n13969_0;
	wire [1:0] w_n13970_0;
	wire [1:0] w_n13973_0;
	wire [1:0] w_n13979_0;
	wire [1:0] w_n13980_0;
	wire [1:0] w_n13982_0;
	wire [1:0] w_n13984_0;
	wire [1:0] w_n13986_0;
	wire [1:0] w_n13992_0;
	wire [1:0] w_n13994_0;
	wire [2:0] w_n13995_0;
	wire [1:0] w_n13998_0;
	wire [1:0] w_n13999_0;
	wire [2:0] w_n14000_0;
	wire [1:0] w_n14002_0;
	wire [1:0] w_n14006_0;
	wire [1:0] w_n14008_0;
	wire [1:0] w_n14009_0;
	wire [2:0] w_n14010_0;
	wire [1:0] w_n14011_0;
	wire [1:0] w_n14014_0;
	wire [1:0] w_n14020_0;
	wire [1:0] w_n14021_0;
	wire [1:0] w_n14023_0;
	wire [1:0] w_n14025_0;
	wire [1:0] w_n14027_0;
	wire [1:0] w_n14033_0;
	wire [1:0] w_n14035_0;
	wire [2:0] w_n14036_0;
	wire [1:0] w_n14039_0;
	wire [1:0] w_n14040_0;
	wire [2:0] w_n14041_0;
	wire [1:0] w_n14043_0;
	wire [1:0] w_n14047_0;
	wire [1:0] w_n14049_0;
	wire [1:0] w_n14050_0;
	wire [2:0] w_n14051_0;
	wire [1:0] w_n14052_0;
	wire [1:0] w_n14055_0;
	wire [1:0] w_n14061_0;
	wire [1:0] w_n14062_0;
	wire [1:0] w_n14064_0;
	wire [1:0] w_n14066_0;
	wire [1:0] w_n14068_0;
	wire [1:0] w_n14074_0;
	wire [1:0] w_n14076_0;
	wire [2:0] w_n14077_0;
	wire [1:0] w_n14080_0;
	wire [1:0] w_n14081_0;
	wire [2:0] w_n14082_0;
	wire [1:0] w_n14084_0;
	wire [1:0] w_n14086_0;
	wire [1:0] w_n14088_0;
	wire [1:0] w_n14094_0;
	wire [2:0] w_n14096_0;
	wire [1:0] w_n14097_0;
	wire [1:0] w_n14099_0;
	wire [1:0] w_n14101_0;
	wire [1:0] w_n14105_0;
	wire [1:0] w_n14107_0;
	wire [1:0] w_n14108_0;
	wire [1:0] w_n14109_0;
	wire [2:0] w_n14110_0;
	wire [1:0] w_n14113_0;
	wire [1:0] w_n14114_0;
	wire [2:0] w_n14115_0;
	wire [1:0] w_n14117_0;
	wire [1:0] w_n14121_0;
	wire [1:0] w_n14123_0;
	wire [1:0] w_n14124_0;
	wire [2:0] w_n14125_0;
	wire [1:0] w_n14126_0;
	wire [1:0] w_n14129_0;
	wire [1:0] w_n14135_0;
	wire [1:0] w_n14136_0;
	wire [1:0] w_n14138_0;
	wire [1:0] w_n14140_0;
	wire [1:0] w_n14142_0;
	wire [1:0] w_n14148_0;
	wire [1:0] w_n14150_0;
	wire [2:0] w_n14151_0;
	wire [1:0] w_n14154_0;
	wire [1:0] w_n14155_0;
	wire [2:0] w_n14156_0;
	wire [1:0] w_n14158_0;
	wire [1:0] w_n14162_0;
	wire [1:0] w_n14164_0;
	wire [1:0] w_n14165_0;
	wire [2:0] w_n14166_0;
	wire [1:0] w_n14167_0;
	wire [1:0] w_n14170_0;
	wire [1:0] w_n14176_0;
	wire [1:0] w_n14177_0;
	wire [1:0] w_n14179_0;
	wire [1:0] w_n14181_0;
	wire [1:0] w_n14183_0;
	wire [1:0] w_n14189_0;
	wire [1:0] w_n14191_0;
	wire [2:0] w_n14192_0;
	wire [1:0] w_n14195_0;
	wire [1:0] w_n14196_0;
	wire [2:0] w_n14197_0;
	wire [1:0] w_n14199_0;
	wire [1:0] w_n14203_0;
	wire [1:0] w_n14205_0;
	wire [1:0] w_n14206_0;
	wire [2:0] w_n14207_0;
	wire [1:0] w_n14211_0;
	wire [1:0] w_n14217_0;
	wire [2:0] w_n14219_0;
	wire [1:0] w_n14221_0;
	wire [2:0] w_n14226_0;
	wire [1:0] w_n14227_0;
	wire [1:0] w_n14228_0;
	wire [1:0] w_n14233_0;
	wire [2:0] w_n14234_0;
	wire [1:0] w_n14239_0;
	wire [1:0] w_n14246_0;
	wire [2:0] w_n14248_0;
	wire [1:0] w_n14248_1;
	wire [1:0] w_n14249_0;
	wire [2:0] w_n14252_0;
	wire [1:0] w_n14253_0;
	wire [1:0] w_n14254_0;
	wire [1:0] w_n14255_0;
	wire [1:0] w_n14257_0;
	wire [1:0] w_n14259_0;
	wire [1:0] w_n14261_0;
	wire [1:0] w_n14270_0;
	wire [2:0] w_n14272_0;
	wire [1:0] w_n14273_0;
	wire [1:0] w_n14277_0;
	wire [1:0] w_n14279_0;
	wire [1:0] w_n14281_0;
	wire [1:0] w_n14286_0;
	wire [1:0] w_n14288_0;
	wire [1:0] w_n14289_0;
	wire [2:0] w_n14290_0;
	wire [1:0] w_n14291_0;
	wire [1:0] w_n14296_0;
	wire [1:0] w_n14297_0;
	wire [1:0] w_n14299_0;
	wire [1:0] w_n14301_0;
	wire [1:0] w_n14304_0;
	wire [1:0] w_n14310_0;
	wire [2:0] w_n14312_0;
	wire [1:0] w_n14313_0;
	wire [1:0] w_n14317_0;
	wire [1:0] w_n14318_0;
	wire [1:0] w_n14320_0;
	wire [1:0] w_n14325_0;
	wire [1:0] w_n14327_0;
	wire [1:0] w_n14328_0;
	wire [2:0] w_n14329_0;
	wire [1:0] w_n14330_0;
	wire [1:0] w_n14334_0;
	wire [1:0] w_n14335_0;
	wire [1:0] w_n14337_0;
	wire [1:0] w_n14339_0;
	wire [1:0] w_n14342_0;
	wire [1:0] w_n14348_0;
	wire [1:0] w_n14350_0;
	wire [2:0] w_n14351_0;
	wire [1:0] w_n14355_0;
	wire [1:0] w_n14356_0;
	wire [2:0] w_n14357_0;
	wire [1:0] w_n14359_0;
	wire [1:0] w_n14364_0;
	wire [1:0] w_n14366_0;
	wire [1:0] w_n14367_0;
	wire [2:0] w_n14368_0;
	wire [1:0] w_n14369_0;
	wire [1:0] w_n14373_0;
	wire [1:0] w_n14379_0;
	wire [1:0] w_n14380_0;
	wire [1:0] w_n14382_0;
	wire [1:0] w_n14384_0;
	wire [1:0] w_n14387_0;
	wire [1:0] w_n14393_0;
	wire [1:0] w_n14395_0;
	wire [2:0] w_n14396_0;
	wire [1:0] w_n14400_0;
	wire [1:0] w_n14401_0;
	wire [2:0] w_n14402_0;
	wire [1:0] w_n14404_0;
	wire [1:0] w_n14409_0;
	wire [1:0] w_n14411_0;
	wire [1:0] w_n14412_0;
	wire [2:0] w_n14413_0;
	wire [1:0] w_n14414_0;
	wire [1:0] w_n14418_0;
	wire [1:0] w_n14424_0;
	wire [1:0] w_n14425_0;
	wire [1:0] w_n14427_0;
	wire [1:0] w_n14429_0;
	wire [1:0] w_n14432_0;
	wire [1:0] w_n14438_0;
	wire [1:0] w_n14440_0;
	wire [2:0] w_n14441_0;
	wire [1:0] w_n14445_0;
	wire [1:0] w_n14446_0;
	wire [2:0] w_n14447_0;
	wire [1:0] w_n14449_0;
	wire [1:0] w_n14454_0;
	wire [1:0] w_n14456_0;
	wire [1:0] w_n14457_0;
	wire [2:0] w_n14458_0;
	wire [1:0] w_n14459_0;
	wire [1:0] w_n14463_0;
	wire [1:0] w_n14469_0;
	wire [1:0] w_n14470_0;
	wire [1:0] w_n14472_0;
	wire [1:0] w_n14474_0;
	wire [1:0] w_n14477_0;
	wire [1:0] w_n14483_0;
	wire [1:0] w_n14485_0;
	wire [2:0] w_n14486_0;
	wire [1:0] w_n14490_0;
	wire [1:0] w_n14491_0;
	wire [2:0] w_n14492_0;
	wire [1:0] w_n14494_0;
	wire [1:0] w_n14499_0;
	wire [1:0] w_n14501_0;
	wire [1:0] w_n14502_0;
	wire [2:0] w_n14503_0;
	wire [1:0] w_n14504_0;
	wire [1:0] w_n14508_0;
	wire [1:0] w_n14514_0;
	wire [1:0] w_n14515_0;
	wire [1:0] w_n14517_0;
	wire [1:0] w_n14519_0;
	wire [1:0] w_n14522_0;
	wire [1:0] w_n14528_0;
	wire [1:0] w_n14530_0;
	wire [2:0] w_n14531_0;
	wire [1:0] w_n14535_0;
	wire [1:0] w_n14536_0;
	wire [2:0] w_n14537_0;
	wire [1:0] w_n14539_0;
	wire [1:0] w_n14544_0;
	wire [1:0] w_n14546_0;
	wire [1:0] w_n14547_0;
	wire [2:0] w_n14548_0;
	wire [1:0] w_n14549_0;
	wire [1:0] w_n14553_0;
	wire [1:0] w_n14559_0;
	wire [1:0] w_n14560_0;
	wire [1:0] w_n14562_0;
	wire [1:0] w_n14564_0;
	wire [1:0] w_n14567_0;
	wire [1:0] w_n14573_0;
	wire [1:0] w_n14575_0;
	wire [2:0] w_n14576_0;
	wire [1:0] w_n14580_0;
	wire [1:0] w_n14581_0;
	wire [2:0] w_n14582_0;
	wire [1:0] w_n14584_0;
	wire [1:0] w_n14589_0;
	wire [1:0] w_n14591_0;
	wire [1:0] w_n14592_0;
	wire [2:0] w_n14593_0;
	wire [1:0] w_n14594_0;
	wire [1:0] w_n14598_0;
	wire [1:0] w_n14604_0;
	wire [1:0] w_n14605_0;
	wire [1:0] w_n14607_0;
	wire [1:0] w_n14609_0;
	wire [1:0] w_n14612_0;
	wire [1:0] w_n14618_0;
	wire [1:0] w_n14620_0;
	wire [2:0] w_n14621_0;
	wire [1:0] w_n14625_0;
	wire [1:0] w_n14626_0;
	wire [2:0] w_n14627_0;
	wire [1:0] w_n14629_0;
	wire [1:0] w_n14634_0;
	wire [1:0] w_n14636_0;
	wire [1:0] w_n14637_0;
	wire [2:0] w_n14638_0;
	wire [1:0] w_n14639_0;
	wire [1:0] w_n14643_0;
	wire [1:0] w_n14649_0;
	wire [1:0] w_n14650_0;
	wire [1:0] w_n14652_0;
	wire [1:0] w_n14657_0;
	wire [1:0] w_n14659_0;
	wire [1:0] w_n14660_0;
	wire [2:0] w_n14661_0;
	wire [1:0] w_n14662_0;
	wire [1:0] w_n14665_0;
	wire [1:0] w_n14667_0;
	wire [1:0] w_n14669_0;
	wire [1:0] w_n14672_0;
	wire [1:0] w_n14678_0;
	wire [2:0] w_n14680_0;
	wire [1:0] w_n14681_0;
	wire [1:0] w_n14685_0;
	wire [1:0] w_n14691_0;
	wire [1:0] w_n14692_0;
	wire [1:0] w_n14694_0;
	wire [1:0] w_n14696_0;
	wire [1:0] w_n14699_0;
	wire [1:0] w_n14705_0;
	wire [1:0] w_n14707_0;
	wire [2:0] w_n14708_0;
	wire [1:0] w_n14712_0;
	wire [1:0] w_n14713_0;
	wire [2:0] w_n14714_0;
	wire [1:0] w_n14716_0;
	wire [1:0] w_n14721_0;
	wire [1:0] w_n14723_0;
	wire [1:0] w_n14724_0;
	wire [2:0] w_n14725_0;
	wire [1:0] w_n14726_0;
	wire [1:0] w_n14730_0;
	wire [1:0] w_n14736_0;
	wire [1:0] w_n14737_0;
	wire [1:0] w_n14739_0;
	wire [1:0] w_n14741_0;
	wire [1:0] w_n14744_0;
	wire [1:0] w_n14750_0;
	wire [1:0] w_n14752_0;
	wire [2:0] w_n14753_0;
	wire [1:0] w_n14757_0;
	wire [1:0] w_n14758_0;
	wire [2:0] w_n14759_0;
	wire [1:0] w_n14761_0;
	wire [1:0] w_n14766_0;
	wire [1:0] w_n14768_0;
	wire [1:0] w_n14769_0;
	wire [2:0] w_n14770_0;
	wire [1:0] w_n14771_0;
	wire [1:0] w_n14775_0;
	wire [1:0] w_n14781_0;
	wire [1:0] w_n14782_0;
	wire [1:0] w_n14784_0;
	wire [1:0] w_n14786_0;
	wire [1:0] w_n14789_0;
	wire [1:0] w_n14795_0;
	wire [2:0] w_n14797_0;
	wire [2:0] w_n14797_1;
	wire [1:0] w_n14800_0;
	wire [2:0] w_n14801_0;
	wire [1:0] w_n14802_0;
	wire [1:0] w_n14808_0;
	wire [2:0] w_n14809_0;
	wire [1:0] w_n14810_0;
	wire [1:0] w_n14815_0;
	wire [2:0] w_n14816_0;
	wire [2:0] w_n14816_1;
	wire [2:0] w_n14816_2;
	wire [2:0] w_n14816_3;
	wire [2:0] w_n14816_4;
	wire [2:0] w_n14816_5;
	wire [2:0] w_n14816_6;
	wire [2:0] w_n14816_7;
	wire [1:0] w_n14816_8;
	wire [2:0] w_n14821_0;
	wire [2:0] w_n14821_1;
	wire [2:0] w_n14821_2;
	wire [2:0] w_n14821_3;
	wire [2:0] w_n14821_4;
	wire [2:0] w_n14821_5;
	wire [2:0] w_n14821_6;
	wire [2:0] w_n14821_7;
	wire [2:0] w_n14821_8;
	wire [2:0] w_n14821_9;
	wire [2:0] w_n14821_10;
	wire [2:0] w_n14821_11;
	wire [2:0] w_n14821_12;
	wire [2:0] w_n14821_13;
	wire [2:0] w_n14821_14;
	wire [2:0] w_n14821_15;
	wire [2:0] w_n14821_16;
	wire [2:0] w_n14821_17;
	wire [2:0] w_n14821_18;
	wire [2:0] w_n14821_19;
	wire [2:0] w_n14821_20;
	wire [2:0] w_n14821_21;
	wire [2:0] w_n14821_22;
	wire [1:0] w_n14824_0;
	wire [2:0] w_n14826_0;
	wire [1:0] w_n14826_1;
	wire [2:0] w_n14827_0;
	wire [2:0] w_n14831_0;
	wire [1:0] w_n14832_0;
	wire [1:0] w_n14833_0;
	wire [1:0] w_n14834_0;
	wire [1:0] w_n14836_0;
	wire [1:0] w_n14838_0;
	wire [1:0] w_n14840_0;
	wire [1:0] w_n14843_0;
	wire [1:0] w_n14848_0;
	wire [2:0] w_n14850_0;
	wire [1:0] w_n14851_0;
	wire [1:0] w_n14855_0;
	wire [1:0] w_n14856_0;
	wire [1:0] w_n14858_0;
	wire [1:0] w_n14862_0;
	wire [1:0] w_n14864_0;
	wire [1:0] w_n14865_0;
	wire [2:0] w_n14866_0;
	wire [1:0] w_n14867_0;
	wire [1:0] w_n14871_0;
	wire [1:0] w_n14873_0;
	wire [1:0] w_n14875_0;
	wire [1:0] w_n14877_0;
	wire [1:0] w_n14880_0;
	wire [1:0] w_n14886_0;
	wire [2:0] w_n14888_0;
	wire [1:0] w_n14889_0;
	wire [1:0] w_n14894_0;
	wire [1:0] w_n14896_0;
	wire [1:0] w_n14898_0;
	wire [1:0] w_n14902_0;
	wire [1:0] w_n14904_0;
	wire [1:0] w_n14905_0;
	wire [2:0] w_n14906_0;
	wire [1:0] w_n14907_0;
	wire [1:0] w_n14913_0;
	wire [1:0] w_n14914_0;
	wire [1:0] w_n14916_0;
	wire [1:0] w_n14918_0;
	wire [1:0] w_n14920_0;
	wire [1:0] w_n14926_0;
	wire [1:0] w_n14928_0;
	wire [2:0] w_n14929_0;
	wire [1:0] w_n14932_0;
	wire [1:0] w_n14933_0;
	wire [2:0] w_n14934_0;
	wire [1:0] w_n14936_0;
	wire [1:0] w_n14940_0;
	wire [1:0] w_n14942_0;
	wire [1:0] w_n14943_0;
	wire [2:0] w_n14944_0;
	wire [1:0] w_n14945_0;
	wire [1:0] w_n14948_0;
	wire [1:0] w_n14954_0;
	wire [1:0] w_n14955_0;
	wire [1:0] w_n14957_0;
	wire [1:0] w_n14959_0;
	wire [1:0] w_n14961_0;
	wire [1:0] w_n14967_0;
	wire [1:0] w_n14969_0;
	wire [2:0] w_n14970_0;
	wire [1:0] w_n14973_0;
	wire [1:0] w_n14974_0;
	wire [2:0] w_n14975_0;
	wire [1:0] w_n14977_0;
	wire [1:0] w_n14981_0;
	wire [1:0] w_n14983_0;
	wire [1:0] w_n14984_0;
	wire [2:0] w_n14985_0;
	wire [1:0] w_n14986_0;
	wire [1:0] w_n14989_0;
	wire [1:0] w_n14995_0;
	wire [1:0] w_n14996_0;
	wire [1:0] w_n14998_0;
	wire [1:0] w_n15000_0;
	wire [1:0] w_n15002_0;
	wire [1:0] w_n15008_0;
	wire [1:0] w_n15010_0;
	wire [2:0] w_n15011_0;
	wire [1:0] w_n15014_0;
	wire [1:0] w_n15015_0;
	wire [2:0] w_n15016_0;
	wire [1:0] w_n15018_0;
	wire [1:0] w_n15022_0;
	wire [1:0] w_n15024_0;
	wire [1:0] w_n15025_0;
	wire [2:0] w_n15026_0;
	wire [1:0] w_n15027_0;
	wire [1:0] w_n15030_0;
	wire [1:0] w_n15036_0;
	wire [1:0] w_n15037_0;
	wire [1:0] w_n15039_0;
	wire [1:0] w_n15041_0;
	wire [1:0] w_n15043_0;
	wire [1:0] w_n15049_0;
	wire [1:0] w_n15051_0;
	wire [2:0] w_n15052_0;
	wire [1:0] w_n15055_0;
	wire [1:0] w_n15056_0;
	wire [2:0] w_n15057_0;
	wire [1:0] w_n15059_0;
	wire [1:0] w_n15063_0;
	wire [1:0] w_n15065_0;
	wire [1:0] w_n15066_0;
	wire [2:0] w_n15067_0;
	wire [1:0] w_n15068_0;
	wire [1:0] w_n15071_0;
	wire [1:0] w_n15077_0;
	wire [1:0] w_n15078_0;
	wire [1:0] w_n15080_0;
	wire [1:0] w_n15082_0;
	wire [1:0] w_n15084_0;
	wire [1:0] w_n15090_0;
	wire [1:0] w_n15092_0;
	wire [2:0] w_n15093_0;
	wire [1:0] w_n15096_0;
	wire [1:0] w_n15097_0;
	wire [2:0] w_n15098_0;
	wire [1:0] w_n15100_0;
	wire [1:0] w_n15104_0;
	wire [1:0] w_n15106_0;
	wire [1:0] w_n15107_0;
	wire [2:0] w_n15108_0;
	wire [1:0] w_n15109_0;
	wire [1:0] w_n15112_0;
	wire [1:0] w_n15118_0;
	wire [1:0] w_n15119_0;
	wire [1:0] w_n15121_0;
	wire [1:0] w_n15123_0;
	wire [1:0] w_n15125_0;
	wire [1:0] w_n15131_0;
	wire [1:0] w_n15133_0;
	wire [2:0] w_n15134_0;
	wire [1:0] w_n15137_0;
	wire [1:0] w_n15138_0;
	wire [2:0] w_n15139_0;
	wire [1:0] w_n15141_0;
	wire [1:0] w_n15145_0;
	wire [1:0] w_n15147_0;
	wire [1:0] w_n15148_0;
	wire [2:0] w_n15149_0;
	wire [1:0] w_n15150_0;
	wire [1:0] w_n15153_0;
	wire [1:0] w_n15159_0;
	wire [1:0] w_n15160_0;
	wire [1:0] w_n15162_0;
	wire [1:0] w_n15164_0;
	wire [1:0] w_n15166_0;
	wire [1:0] w_n15172_0;
	wire [1:0] w_n15174_0;
	wire [2:0] w_n15175_0;
	wire [1:0] w_n15178_0;
	wire [1:0] w_n15179_0;
	wire [2:0] w_n15180_0;
	wire [1:0] w_n15182_0;
	wire [1:0] w_n15186_0;
	wire [1:0] w_n15188_0;
	wire [1:0] w_n15189_0;
	wire [2:0] w_n15190_0;
	wire [1:0] w_n15191_0;
	wire [1:0] w_n15194_0;
	wire [1:0] w_n15200_0;
	wire [1:0] w_n15201_0;
	wire [1:0] w_n15203_0;
	wire [1:0] w_n15205_0;
	wire [1:0] w_n15207_0;
	wire [1:0] w_n15213_0;
	wire [1:0] w_n15215_0;
	wire [2:0] w_n15216_0;
	wire [1:0] w_n15219_0;
	wire [1:0] w_n15220_0;
	wire [2:0] w_n15221_0;
	wire [1:0] w_n15223_0;
	wire [1:0] w_n15225_0;
	wire [1:0] w_n15227_0;
	wire [1:0] w_n15233_0;
	wire [2:0] w_n15235_0;
	wire [1:0] w_n15236_0;
	wire [1:0] w_n15239_0;
	wire [1:0] w_n15241_0;
	wire [1:0] w_n15245_0;
	wire [1:0] w_n15247_0;
	wire [1:0] w_n15248_0;
	wire [1:0] w_n15249_0;
	wire [2:0] w_n15250_0;
	wire [1:0] w_n15253_0;
	wire [1:0] w_n15254_0;
	wire [2:0] w_n15255_0;
	wire [1:0] w_n15257_0;
	wire [1:0] w_n15261_0;
	wire [1:0] w_n15263_0;
	wire [1:0] w_n15264_0;
	wire [2:0] w_n15265_0;
	wire [1:0] w_n15266_0;
	wire [1:0] w_n15269_0;
	wire [1:0] w_n15275_0;
	wire [1:0] w_n15276_0;
	wire [1:0] w_n15278_0;
	wire [1:0] w_n15280_0;
	wire [1:0] w_n15282_0;
	wire [1:0] w_n15288_0;
	wire [1:0] w_n15290_0;
	wire [2:0] w_n15291_0;
	wire [1:0] w_n15294_0;
	wire [1:0] w_n15295_0;
	wire [2:0] w_n15296_0;
	wire [1:0] w_n15298_0;
	wire [1:0] w_n15302_0;
	wire [1:0] w_n15304_0;
	wire [1:0] w_n15305_0;
	wire [2:0] w_n15306_0;
	wire [1:0] w_n15307_0;
	wire [1:0] w_n15310_0;
	wire [1:0] w_n15316_0;
	wire [1:0] w_n15317_0;
	wire [1:0] w_n15319_0;
	wire [1:0] w_n15321_0;
	wire [1:0] w_n15323_0;
	wire [1:0] w_n15329_0;
	wire [2:0] w_n15331_0;
	wire [1:0] w_n15336_0;
	wire [2:0] w_n15338_0;
	wire [2:0] w_n15342_0;
	wire [1:0] w_n15343_0;
	wire [1:0] w_n15348_0;
	wire [2:0] w_n15349_0;
	wire [1:0] w_n15354_0;
	wire [1:0] w_n15361_0;
	wire [2:0] w_n15364_0;
	wire [1:0] w_n15364_1;
	wire [1:0] w_n15365_0;
	wire [2:0] w_n15368_0;
	wire [1:0] w_n15369_0;
	wire [1:0] w_n15370_0;
	wire [1:0] w_n15371_0;
	wire [1:0] w_n15373_0;
	wire [1:0] w_n15375_0;
	wire [1:0] w_n15377_0;
	wire [1:0] w_n15386_0;
	wire [2:0] w_n15388_0;
	wire [1:0] w_n15389_0;
	wire [1:0] w_n15393_0;
	wire [1:0] w_n15395_0;
	wire [1:0] w_n15397_0;
	wire [1:0] w_n15402_0;
	wire [1:0] w_n15404_0;
	wire [1:0] w_n15405_0;
	wire [2:0] w_n15406_0;
	wire [1:0] w_n15407_0;
	wire [1:0] w_n15412_0;
	wire [1:0] w_n15413_0;
	wire [1:0] w_n15415_0;
	wire [1:0] w_n15417_0;
	wire [1:0] w_n15420_0;
	wire [1:0] w_n15426_0;
	wire [2:0] w_n15428_0;
	wire [1:0] w_n15429_0;
	wire [1:0] w_n15433_0;
	wire [1:0] w_n15434_0;
	wire [1:0] w_n15436_0;
	wire [1:0] w_n15441_0;
	wire [1:0] w_n15443_0;
	wire [1:0] w_n15444_0;
	wire [2:0] w_n15445_0;
	wire [1:0] w_n15446_0;
	wire [1:0] w_n15450_0;
	wire [1:0] w_n15451_0;
	wire [1:0] w_n15453_0;
	wire [1:0] w_n15455_0;
	wire [1:0] w_n15458_0;
	wire [1:0] w_n15464_0;
	wire [1:0] w_n15466_0;
	wire [2:0] w_n15467_0;
	wire [1:0] w_n15471_0;
	wire [1:0] w_n15472_0;
	wire [2:0] w_n15473_0;
	wire [1:0] w_n15475_0;
	wire [1:0] w_n15480_0;
	wire [1:0] w_n15482_0;
	wire [1:0] w_n15483_0;
	wire [2:0] w_n15484_0;
	wire [1:0] w_n15485_0;
	wire [1:0] w_n15489_0;
	wire [1:0] w_n15495_0;
	wire [1:0] w_n15496_0;
	wire [1:0] w_n15498_0;
	wire [1:0] w_n15500_0;
	wire [1:0] w_n15503_0;
	wire [1:0] w_n15509_0;
	wire [1:0] w_n15511_0;
	wire [2:0] w_n15512_0;
	wire [1:0] w_n15516_0;
	wire [1:0] w_n15517_0;
	wire [2:0] w_n15518_0;
	wire [1:0] w_n15520_0;
	wire [1:0] w_n15525_0;
	wire [1:0] w_n15527_0;
	wire [1:0] w_n15528_0;
	wire [2:0] w_n15529_0;
	wire [1:0] w_n15530_0;
	wire [1:0] w_n15534_0;
	wire [1:0] w_n15540_0;
	wire [1:0] w_n15541_0;
	wire [1:0] w_n15543_0;
	wire [1:0] w_n15545_0;
	wire [1:0] w_n15548_0;
	wire [1:0] w_n15554_0;
	wire [1:0] w_n15556_0;
	wire [2:0] w_n15557_0;
	wire [1:0] w_n15561_0;
	wire [1:0] w_n15562_0;
	wire [2:0] w_n15563_0;
	wire [1:0] w_n15565_0;
	wire [1:0] w_n15570_0;
	wire [1:0] w_n15572_0;
	wire [1:0] w_n15573_0;
	wire [2:0] w_n15574_0;
	wire [1:0] w_n15575_0;
	wire [1:0] w_n15579_0;
	wire [1:0] w_n15585_0;
	wire [1:0] w_n15586_0;
	wire [1:0] w_n15588_0;
	wire [1:0] w_n15590_0;
	wire [1:0] w_n15593_0;
	wire [1:0] w_n15599_0;
	wire [1:0] w_n15601_0;
	wire [2:0] w_n15602_0;
	wire [1:0] w_n15606_0;
	wire [1:0] w_n15607_0;
	wire [2:0] w_n15608_0;
	wire [1:0] w_n15610_0;
	wire [1:0] w_n15615_0;
	wire [1:0] w_n15617_0;
	wire [1:0] w_n15618_0;
	wire [2:0] w_n15619_0;
	wire [1:0] w_n15620_0;
	wire [1:0] w_n15624_0;
	wire [1:0] w_n15630_0;
	wire [1:0] w_n15631_0;
	wire [1:0] w_n15633_0;
	wire [1:0] w_n15635_0;
	wire [1:0] w_n15638_0;
	wire [1:0] w_n15644_0;
	wire [1:0] w_n15646_0;
	wire [2:0] w_n15647_0;
	wire [1:0] w_n15651_0;
	wire [1:0] w_n15652_0;
	wire [2:0] w_n15653_0;
	wire [1:0] w_n15655_0;
	wire [1:0] w_n15660_0;
	wire [1:0] w_n15662_0;
	wire [1:0] w_n15663_0;
	wire [2:0] w_n15664_0;
	wire [1:0] w_n15665_0;
	wire [1:0] w_n15669_0;
	wire [1:0] w_n15675_0;
	wire [1:0] w_n15676_0;
	wire [1:0] w_n15678_0;
	wire [1:0] w_n15680_0;
	wire [1:0] w_n15683_0;
	wire [1:0] w_n15689_0;
	wire [1:0] w_n15691_0;
	wire [2:0] w_n15692_0;
	wire [1:0] w_n15696_0;
	wire [1:0] w_n15697_0;
	wire [2:0] w_n15698_0;
	wire [1:0] w_n15700_0;
	wire [1:0] w_n15705_0;
	wire [1:0] w_n15707_0;
	wire [1:0] w_n15708_0;
	wire [2:0] w_n15709_0;
	wire [1:0] w_n15710_0;
	wire [1:0] w_n15714_0;
	wire [1:0] w_n15720_0;
	wire [1:0] w_n15721_0;
	wire [1:0] w_n15723_0;
	wire [1:0] w_n15725_0;
	wire [1:0] w_n15728_0;
	wire [1:0] w_n15734_0;
	wire [1:0] w_n15736_0;
	wire [2:0] w_n15737_0;
	wire [1:0] w_n15741_0;
	wire [1:0] w_n15742_0;
	wire [2:0] w_n15743_0;
	wire [1:0] w_n15745_0;
	wire [1:0] w_n15750_0;
	wire [1:0] w_n15752_0;
	wire [1:0] w_n15753_0;
	wire [2:0] w_n15754_0;
	wire [1:0] w_n15755_0;
	wire [1:0] w_n15759_0;
	wire [1:0] w_n15765_0;
	wire [1:0] w_n15766_0;
	wire [1:0] w_n15768_0;
	wire [1:0] w_n15770_0;
	wire [1:0] w_n15773_0;
	wire [1:0] w_n15779_0;
	wire [1:0] w_n15781_0;
	wire [2:0] w_n15782_0;
	wire [1:0] w_n15786_0;
	wire [1:0] w_n15787_0;
	wire [2:0] w_n15788_0;
	wire [1:0] w_n15790_0;
	wire [1:0] w_n15795_0;
	wire [1:0] w_n15797_0;
	wire [1:0] w_n15798_0;
	wire [2:0] w_n15799_0;
	wire [1:0] w_n15800_0;
	wire [1:0] w_n15804_0;
	wire [1:0] w_n15810_0;
	wire [1:0] w_n15811_0;
	wire [1:0] w_n15813_0;
	wire [1:0] w_n15818_0;
	wire [1:0] w_n15820_0;
	wire [1:0] w_n15821_0;
	wire [2:0] w_n15822_0;
	wire [1:0] w_n15823_0;
	wire [1:0] w_n15825_0;
	wire [1:0] w_n15827_0;
	wire [1:0] w_n15829_0;
	wire [1:0] w_n15832_0;
	wire [1:0] w_n15838_0;
	wire [2:0] w_n15840_0;
	wire [1:0] w_n15841_0;
	wire [1:0] w_n15845_0;
	wire [1:0] w_n15851_0;
	wire [1:0] w_n15852_0;
	wire [1:0] w_n15854_0;
	wire [1:0] w_n15856_0;
	wire [1:0] w_n15859_0;
	wire [1:0] w_n15865_0;
	wire [1:0] w_n15867_0;
	wire [2:0] w_n15868_0;
	wire [1:0] w_n15872_0;
	wire [1:0] w_n15873_0;
	wire [2:0] w_n15874_0;
	wire [1:0] w_n15876_0;
	wire [1:0] w_n15881_0;
	wire [1:0] w_n15883_0;
	wire [1:0] w_n15884_0;
	wire [2:0] w_n15885_0;
	wire [1:0] w_n15886_0;
	wire [1:0] w_n15890_0;
	wire [1:0] w_n15896_0;
	wire [1:0] w_n15897_0;
	wire [1:0] w_n15899_0;
	wire [1:0] w_n15901_0;
	wire [1:0] w_n15904_0;
	wire [1:0] w_n15910_0;
	wire [1:0] w_n15912_0;
	wire [2:0] w_n15913_0;
	wire [1:0] w_n15917_0;
	wire [1:0] w_n15918_0;
	wire [2:0] w_n15919_0;
	wire [1:0] w_n15921_0;
	wire [1:0] w_n15926_0;
	wire [1:0] w_n15928_0;
	wire [1:0] w_n15929_0;
	wire [2:0] w_n15930_0;
	wire [2:0] w_n15930_1;
	wire [1:0] w_n15933_0;
	wire [2:0] w_n15934_0;
	wire [1:0] w_n15935_0;
	wire [1:0] w_n15936_0;
	wire [1:0] w_n15942_0;
	wire [2:0] w_n15943_0;
	wire [1:0] w_n15944_0;
	wire [1:0] w_n15949_0;
	wire [2:0] w_n15950_0;
	wire [2:0] w_n15950_1;
	wire [2:0] w_n15950_2;
	wire [2:0] w_n15950_3;
	wire [2:0] w_n15950_4;
	wire [2:0] w_n15950_5;
	wire [2:0] w_n15950_6;
	wire [2:0] w_n15955_0;
	wire [2:0] w_n15955_1;
	wire [2:0] w_n15955_2;
	wire [2:0] w_n15955_3;
	wire [2:0] w_n15955_4;
	wire [2:0] w_n15955_5;
	wire [2:0] w_n15955_6;
	wire [2:0] w_n15955_7;
	wire [2:0] w_n15955_8;
	wire [2:0] w_n15955_9;
	wire [2:0] w_n15955_10;
	wire [2:0] w_n15955_11;
	wire [2:0] w_n15955_12;
	wire [2:0] w_n15955_13;
	wire [2:0] w_n15955_14;
	wire [2:0] w_n15955_15;
	wire [2:0] w_n15955_16;
	wire [2:0] w_n15955_17;
	wire [2:0] w_n15955_18;
	wire [2:0] w_n15955_19;
	wire [2:0] w_n15955_20;
	wire [1:0] w_n15955_21;
	wire [1:0] w_n15959_0;
	wire [2:0] w_n15961_0;
	wire [1:0] w_n15961_1;
	wire [2:0] w_n15962_0;
	wire [2:0] w_n15966_0;
	wire [1:0] w_n15967_0;
	wire [1:0] w_n15968_0;
	wire [1:0] w_n15969_0;
	wire [1:0] w_n15971_0;
	wire [1:0] w_n15973_0;
	wire [1:0] w_n15975_0;
	wire [1:0] w_n15978_0;
	wire [1:0] w_n15983_0;
	wire [2:0] w_n15985_0;
	wire [1:0] w_n15986_0;
	wire [1:0] w_n15990_0;
	wire [1:0] w_n15991_0;
	wire [1:0] w_n15993_0;
	wire [1:0] w_n15997_0;
	wire [1:0] w_n15999_0;
	wire [1:0] w_n16000_0;
	wire [2:0] w_n16001_0;
	wire [1:0] w_n16002_0;
	wire [1:0] w_n16006_0;
	wire [1:0] w_n16008_0;
	wire [1:0] w_n16010_0;
	wire [1:0] w_n16012_0;
	wire [1:0] w_n16015_0;
	wire [1:0] w_n16021_0;
	wire [2:0] w_n16023_0;
	wire [1:0] w_n16024_0;
	wire [1:0] w_n16029_0;
	wire [1:0] w_n16031_0;
	wire [1:0] w_n16033_0;
	wire [1:0] w_n16037_0;
	wire [1:0] w_n16039_0;
	wire [1:0] w_n16040_0;
	wire [2:0] w_n16041_0;
	wire [1:0] w_n16042_0;
	wire [1:0] w_n16048_0;
	wire [1:0] w_n16049_0;
	wire [1:0] w_n16051_0;
	wire [1:0] w_n16053_0;
	wire [1:0] w_n16055_0;
	wire [1:0] w_n16061_0;
	wire [1:0] w_n16063_0;
	wire [2:0] w_n16064_0;
	wire [1:0] w_n16067_0;
	wire [1:0] w_n16068_0;
	wire [2:0] w_n16069_0;
	wire [1:0] w_n16071_0;
	wire [1:0] w_n16075_0;
	wire [1:0] w_n16077_0;
	wire [1:0] w_n16078_0;
	wire [2:0] w_n16079_0;
	wire [1:0] w_n16080_0;
	wire [1:0] w_n16083_0;
	wire [1:0] w_n16089_0;
	wire [1:0] w_n16090_0;
	wire [1:0] w_n16092_0;
	wire [1:0] w_n16094_0;
	wire [1:0] w_n16096_0;
	wire [1:0] w_n16102_0;
	wire [1:0] w_n16104_0;
	wire [2:0] w_n16105_0;
	wire [1:0] w_n16108_0;
	wire [1:0] w_n16109_0;
	wire [2:0] w_n16110_0;
	wire [1:0] w_n16112_0;
	wire [1:0] w_n16116_0;
	wire [1:0] w_n16118_0;
	wire [1:0] w_n16119_0;
	wire [2:0] w_n16120_0;
	wire [1:0] w_n16121_0;
	wire [1:0] w_n16124_0;
	wire [1:0] w_n16130_0;
	wire [1:0] w_n16131_0;
	wire [1:0] w_n16133_0;
	wire [1:0] w_n16135_0;
	wire [1:0] w_n16137_0;
	wire [1:0] w_n16143_0;
	wire [1:0] w_n16145_0;
	wire [2:0] w_n16146_0;
	wire [1:0] w_n16149_0;
	wire [1:0] w_n16150_0;
	wire [2:0] w_n16151_0;
	wire [1:0] w_n16153_0;
	wire [1:0] w_n16157_0;
	wire [1:0] w_n16159_0;
	wire [1:0] w_n16160_0;
	wire [2:0] w_n16161_0;
	wire [1:0] w_n16162_0;
	wire [1:0] w_n16165_0;
	wire [1:0] w_n16171_0;
	wire [1:0] w_n16172_0;
	wire [1:0] w_n16174_0;
	wire [1:0] w_n16176_0;
	wire [1:0] w_n16178_0;
	wire [1:0] w_n16184_0;
	wire [1:0] w_n16186_0;
	wire [2:0] w_n16187_0;
	wire [1:0] w_n16190_0;
	wire [1:0] w_n16191_0;
	wire [2:0] w_n16192_0;
	wire [1:0] w_n16194_0;
	wire [1:0] w_n16198_0;
	wire [1:0] w_n16200_0;
	wire [1:0] w_n16201_0;
	wire [2:0] w_n16202_0;
	wire [1:0] w_n16203_0;
	wire [1:0] w_n16206_0;
	wire [1:0] w_n16212_0;
	wire [1:0] w_n16213_0;
	wire [1:0] w_n16215_0;
	wire [1:0] w_n16217_0;
	wire [1:0] w_n16219_0;
	wire [1:0] w_n16225_0;
	wire [1:0] w_n16227_0;
	wire [2:0] w_n16228_0;
	wire [1:0] w_n16231_0;
	wire [1:0] w_n16232_0;
	wire [2:0] w_n16233_0;
	wire [1:0] w_n16235_0;
	wire [1:0] w_n16239_0;
	wire [1:0] w_n16241_0;
	wire [1:0] w_n16242_0;
	wire [2:0] w_n16243_0;
	wire [1:0] w_n16244_0;
	wire [1:0] w_n16247_0;
	wire [1:0] w_n16253_0;
	wire [1:0] w_n16254_0;
	wire [1:0] w_n16256_0;
	wire [1:0] w_n16258_0;
	wire [1:0] w_n16260_0;
	wire [1:0] w_n16266_0;
	wire [1:0] w_n16268_0;
	wire [2:0] w_n16269_0;
	wire [1:0] w_n16272_0;
	wire [1:0] w_n16273_0;
	wire [2:0] w_n16274_0;
	wire [1:0] w_n16276_0;
	wire [1:0] w_n16280_0;
	wire [1:0] w_n16282_0;
	wire [1:0] w_n16283_0;
	wire [2:0] w_n16284_0;
	wire [1:0] w_n16285_0;
	wire [1:0] w_n16288_0;
	wire [1:0] w_n16294_0;
	wire [1:0] w_n16295_0;
	wire [1:0] w_n16297_0;
	wire [1:0] w_n16299_0;
	wire [1:0] w_n16301_0;
	wire [1:0] w_n16307_0;
	wire [1:0] w_n16309_0;
	wire [2:0] w_n16310_0;
	wire [1:0] w_n16313_0;
	wire [1:0] w_n16314_0;
	wire [2:0] w_n16315_0;
	wire [1:0] w_n16317_0;
	wire [1:0] w_n16321_0;
	wire [1:0] w_n16323_0;
	wire [1:0] w_n16324_0;
	wire [2:0] w_n16325_0;
	wire [1:0] w_n16326_0;
	wire [1:0] w_n16329_0;
	wire [1:0] w_n16335_0;
	wire [1:0] w_n16336_0;
	wire [1:0] w_n16338_0;
	wire [1:0] w_n16340_0;
	wire [1:0] w_n16342_0;
	wire [1:0] w_n16348_0;
	wire [1:0] w_n16350_0;
	wire [2:0] w_n16351_0;
	wire [1:0] w_n16354_0;
	wire [1:0] w_n16355_0;
	wire [2:0] w_n16356_0;
	wire [1:0] w_n16358_0;
	wire [1:0] w_n16362_0;
	wire [1:0] w_n16364_0;
	wire [1:0] w_n16365_0;
	wire [2:0] w_n16366_0;
	wire [1:0] w_n16367_0;
	wire [1:0] w_n16370_0;
	wire [1:0] w_n16376_0;
	wire [1:0] w_n16377_0;
	wire [1:0] w_n16379_0;
	wire [1:0] w_n16381_0;
	wire [1:0] w_n16383_0;
	wire [1:0] w_n16389_0;
	wire [1:0] w_n16391_0;
	wire [2:0] w_n16392_0;
	wire [1:0] w_n16395_0;
	wire [1:0] w_n16396_0;
	wire [2:0] w_n16397_0;
	wire [1:0] w_n16399_0;
	wire [1:0] w_n16401_0;
	wire [1:0] w_n16403_0;
	wire [1:0] w_n16409_0;
	wire [2:0] w_n16411_0;
	wire [1:0] w_n16412_0;
	wire [1:0] w_n16414_0;
	wire [1:0] w_n16416_0;
	wire [1:0] w_n16420_0;
	wire [1:0] w_n16422_0;
	wire [1:0] w_n16423_0;
	wire [1:0] w_n16424_0;
	wire [2:0] w_n16425_0;
	wire [1:0] w_n16428_0;
	wire [1:0] w_n16429_0;
	wire [2:0] w_n16430_0;
	wire [1:0] w_n16432_0;
	wire [1:0] w_n16436_0;
	wire [1:0] w_n16438_0;
	wire [1:0] w_n16439_0;
	wire [2:0] w_n16440_0;
	wire [1:0] w_n16441_0;
	wire [1:0] w_n16444_0;
	wire [1:0] w_n16450_0;
	wire [1:0] w_n16451_0;
	wire [1:0] w_n16453_0;
	wire [1:0] w_n16455_0;
	wire [1:0] w_n16457_0;
	wire [1:0] w_n16463_0;
	wire [1:0] w_n16465_0;
	wire [2:0] w_n16466_0;
	wire [1:0] w_n16469_0;
	wire [1:0] w_n16470_0;
	wire [2:0] w_n16471_0;
	wire [1:0] w_n16473_0;
	wire [1:0] w_n16477_0;
	wire [1:0] w_n16479_0;
	wire [1:0] w_n16480_0;
	wire [2:0] w_n16481_0;
	wire [1:0] w_n16485_0;
	wire [1:0] w_n16491_0;
	wire [2:0] w_n16493_0;
	wire [1:0] w_n16495_0;
	wire [2:0] w_n16500_0;
	wire [1:0] w_n16501_0;
	wire [1:0] w_n16502_0;
	wire [1:0] w_n16507_0;
	wire [2:0] w_n16508_0;
	wire [1:0] w_n16513_0;
	wire [1:0] w_n16521_0;
	wire [2:0] w_n16523_0;
	wire [1:0] w_n16523_1;
	wire [1:0] w_n16524_0;
	wire [2:0] w_n16527_0;
	wire [1:0] w_n16528_0;
	wire [1:0] w_n16529_0;
	wire [1:0] w_n16530_0;
	wire [1:0] w_n16532_0;
	wire [1:0] w_n16534_0;
	wire [1:0] w_n16536_0;
	wire [1:0] w_n16545_0;
	wire [2:0] w_n16547_0;
	wire [1:0] w_n16548_0;
	wire [1:0] w_n16552_0;
	wire [1:0] w_n16554_0;
	wire [1:0] w_n16556_0;
	wire [1:0] w_n16561_0;
	wire [1:0] w_n16563_0;
	wire [1:0] w_n16564_0;
	wire [2:0] w_n16565_0;
	wire [1:0] w_n16566_0;
	wire [1:0] w_n16571_0;
	wire [1:0] w_n16572_0;
	wire [1:0] w_n16574_0;
	wire [1:0] w_n16576_0;
	wire [1:0] w_n16579_0;
	wire [1:0] w_n16585_0;
	wire [2:0] w_n16587_0;
	wire [1:0] w_n16588_0;
	wire [1:0] w_n16592_0;
	wire [1:0] w_n16593_0;
	wire [1:0] w_n16595_0;
	wire [1:0] w_n16600_0;
	wire [1:0] w_n16602_0;
	wire [1:0] w_n16603_0;
	wire [2:0] w_n16604_0;
	wire [1:0] w_n16605_0;
	wire [1:0] w_n16609_0;
	wire [1:0] w_n16610_0;
	wire [1:0] w_n16612_0;
	wire [1:0] w_n16614_0;
	wire [1:0] w_n16617_0;
	wire [1:0] w_n16623_0;
	wire [1:0] w_n16625_0;
	wire [2:0] w_n16626_0;
	wire [1:0] w_n16630_0;
	wire [1:0] w_n16631_0;
	wire [2:0] w_n16632_0;
	wire [1:0] w_n16634_0;
	wire [1:0] w_n16639_0;
	wire [1:0] w_n16641_0;
	wire [1:0] w_n16642_0;
	wire [2:0] w_n16643_0;
	wire [1:0] w_n16644_0;
	wire [1:0] w_n16648_0;
	wire [1:0] w_n16654_0;
	wire [1:0] w_n16655_0;
	wire [1:0] w_n16657_0;
	wire [1:0] w_n16659_0;
	wire [1:0] w_n16662_0;
	wire [1:0] w_n16668_0;
	wire [1:0] w_n16670_0;
	wire [2:0] w_n16671_0;
	wire [1:0] w_n16675_0;
	wire [1:0] w_n16676_0;
	wire [2:0] w_n16677_0;
	wire [1:0] w_n16679_0;
	wire [1:0] w_n16684_0;
	wire [1:0] w_n16686_0;
	wire [1:0] w_n16687_0;
	wire [2:0] w_n16688_0;
	wire [1:0] w_n16689_0;
	wire [1:0] w_n16693_0;
	wire [1:0] w_n16699_0;
	wire [1:0] w_n16700_0;
	wire [1:0] w_n16702_0;
	wire [1:0] w_n16704_0;
	wire [1:0] w_n16707_0;
	wire [1:0] w_n16713_0;
	wire [1:0] w_n16715_0;
	wire [2:0] w_n16716_0;
	wire [1:0] w_n16720_0;
	wire [1:0] w_n16721_0;
	wire [2:0] w_n16722_0;
	wire [1:0] w_n16724_0;
	wire [1:0] w_n16729_0;
	wire [1:0] w_n16731_0;
	wire [1:0] w_n16732_0;
	wire [2:0] w_n16733_0;
	wire [1:0] w_n16734_0;
	wire [1:0] w_n16738_0;
	wire [1:0] w_n16744_0;
	wire [1:0] w_n16745_0;
	wire [1:0] w_n16747_0;
	wire [1:0] w_n16749_0;
	wire [1:0] w_n16752_0;
	wire [1:0] w_n16758_0;
	wire [1:0] w_n16760_0;
	wire [2:0] w_n16761_0;
	wire [1:0] w_n16765_0;
	wire [1:0] w_n16766_0;
	wire [2:0] w_n16767_0;
	wire [1:0] w_n16769_0;
	wire [1:0] w_n16774_0;
	wire [1:0] w_n16776_0;
	wire [1:0] w_n16777_0;
	wire [2:0] w_n16778_0;
	wire [1:0] w_n16779_0;
	wire [1:0] w_n16783_0;
	wire [1:0] w_n16789_0;
	wire [1:0] w_n16790_0;
	wire [1:0] w_n16792_0;
	wire [1:0] w_n16794_0;
	wire [1:0] w_n16797_0;
	wire [1:0] w_n16803_0;
	wire [1:0] w_n16805_0;
	wire [2:0] w_n16806_0;
	wire [1:0] w_n16810_0;
	wire [1:0] w_n16811_0;
	wire [2:0] w_n16812_0;
	wire [1:0] w_n16814_0;
	wire [1:0] w_n16819_0;
	wire [1:0] w_n16821_0;
	wire [1:0] w_n16822_0;
	wire [2:0] w_n16823_0;
	wire [1:0] w_n16824_0;
	wire [1:0] w_n16828_0;
	wire [1:0] w_n16834_0;
	wire [1:0] w_n16835_0;
	wire [1:0] w_n16837_0;
	wire [1:0] w_n16839_0;
	wire [1:0] w_n16842_0;
	wire [1:0] w_n16848_0;
	wire [1:0] w_n16850_0;
	wire [2:0] w_n16851_0;
	wire [1:0] w_n16855_0;
	wire [1:0] w_n16856_0;
	wire [2:0] w_n16857_0;
	wire [1:0] w_n16859_0;
	wire [1:0] w_n16864_0;
	wire [1:0] w_n16866_0;
	wire [1:0] w_n16867_0;
	wire [2:0] w_n16868_0;
	wire [1:0] w_n16869_0;
	wire [1:0] w_n16873_0;
	wire [1:0] w_n16879_0;
	wire [1:0] w_n16880_0;
	wire [1:0] w_n16882_0;
	wire [1:0] w_n16884_0;
	wire [1:0] w_n16887_0;
	wire [1:0] w_n16893_0;
	wire [1:0] w_n16895_0;
	wire [2:0] w_n16896_0;
	wire [1:0] w_n16900_0;
	wire [1:0] w_n16901_0;
	wire [2:0] w_n16902_0;
	wire [1:0] w_n16904_0;
	wire [1:0] w_n16909_0;
	wire [1:0] w_n16911_0;
	wire [1:0] w_n16912_0;
	wire [2:0] w_n16913_0;
	wire [1:0] w_n16914_0;
	wire [1:0] w_n16918_0;
	wire [1:0] w_n16924_0;
	wire [1:0] w_n16925_0;
	wire [1:0] w_n16927_0;
	wire [1:0] w_n16929_0;
	wire [1:0] w_n16932_0;
	wire [1:0] w_n16938_0;
	wire [1:0] w_n16940_0;
	wire [2:0] w_n16941_0;
	wire [1:0] w_n16945_0;
	wire [1:0] w_n16946_0;
	wire [2:0] w_n16947_0;
	wire [1:0] w_n16949_0;
	wire [1:0] w_n16954_0;
	wire [1:0] w_n16956_0;
	wire [1:0] w_n16957_0;
	wire [2:0] w_n16958_0;
	wire [1:0] w_n16959_0;
	wire [1:0] w_n16963_0;
	wire [1:0] w_n16969_0;
	wire [1:0] w_n16970_0;
	wire [1:0] w_n16972_0;
	wire [1:0] w_n16974_0;
	wire [1:0] w_n16977_0;
	wire [1:0] w_n16983_0;
	wire [1:0] w_n16985_0;
	wire [2:0] w_n16986_0;
	wire [1:0] w_n16990_0;
	wire [1:0] w_n16991_0;
	wire [2:0] w_n16992_0;
	wire [1:0] w_n16994_0;
	wire [1:0] w_n16999_0;
	wire [1:0] w_n17001_0;
	wire [1:0] w_n17002_0;
	wire [2:0] w_n17003_0;
	wire [1:0] w_n17004_0;
	wire [1:0] w_n17008_0;
	wire [1:0] w_n17014_0;
	wire [1:0] w_n17015_0;
	wire [1:0] w_n17017_0;
	wire [1:0] w_n17022_0;
	wire [1:0] w_n17024_0;
	wire [1:0] w_n17025_0;
	wire [2:0] w_n17026_0;
	wire [1:0] w_n17027_0;
	wire [1:0] w_n17029_0;
	wire [1:0] w_n17031_0;
	wire [1:0] w_n17033_0;
	wire [1:0] w_n17036_0;
	wire [1:0] w_n17042_0;
	wire [2:0] w_n17044_0;
	wire [1:0] w_n17045_0;
	wire [1:0] w_n17049_0;
	wire [1:0] w_n17055_0;
	wire [1:0] w_n17056_0;
	wire [1:0] w_n17058_0;
	wire [1:0] w_n17060_0;
	wire [1:0] w_n17063_0;
	wire [1:0] w_n17069_0;
	wire [1:0] w_n17071_0;
	wire [2:0] w_n17072_0;
	wire [1:0] w_n17076_0;
	wire [1:0] w_n17077_0;
	wire [2:0] w_n17078_0;
	wire [1:0] w_n17080_0;
	wire [1:0] w_n17085_0;
	wire [1:0] w_n17087_0;
	wire [1:0] w_n17088_0;
	wire [2:0] w_n17089_0;
	wire [1:0] w_n17090_0;
	wire [1:0] w_n17094_0;
	wire [1:0] w_n17100_0;
	wire [1:0] w_n17101_0;
	wire [1:0] w_n17103_0;
	wire [1:0] w_n17105_0;
	wire [1:0] w_n17108_0;
	wire [1:0] w_n17114_0;
	wire [2:0] w_n17116_0;
	wire [2:0] w_n17116_1;
	wire [1:0] w_n17119_0;
	wire [2:0] w_n17120_0;
	wire [1:0] w_n17121_0;
	wire [1:0] w_n17127_0;
	wire [2:0] w_n17128_0;
	wire [1:0] w_n17129_0;
	wire [1:0] w_n17134_0;
	wire [2:0] w_n17135_0;
	wire [2:0] w_n17135_1;
	wire [2:0] w_n17135_2;
	wire [2:0] w_n17135_3;
	wire [2:0] w_n17135_4;
	wire [1:0] w_n17135_5;
	wire [2:0] w_n17140_0;
	wire [2:0] w_n17140_1;
	wire [2:0] w_n17140_2;
	wire [2:0] w_n17140_3;
	wire [2:0] w_n17140_4;
	wire [2:0] w_n17140_5;
	wire [2:0] w_n17140_6;
	wire [2:0] w_n17140_7;
	wire [2:0] w_n17140_8;
	wire [2:0] w_n17140_9;
	wire [2:0] w_n17140_10;
	wire [2:0] w_n17140_11;
	wire [2:0] w_n17140_12;
	wire [2:0] w_n17140_13;
	wire [2:0] w_n17140_14;
	wire [2:0] w_n17140_15;
	wire [2:0] w_n17140_16;
	wire [2:0] w_n17140_17;
	wire [2:0] w_n17140_18;
	wire [2:0] w_n17140_19;
	wire [2:0] w_n17140_20;
	wire [1:0] w_n17143_0;
	wire [2:0] w_n17145_0;
	wire [1:0] w_n17145_1;
	wire [2:0] w_n17146_0;
	wire [2:0] w_n17150_0;
	wire [1:0] w_n17151_0;
	wire [1:0] w_n17152_0;
	wire [1:0] w_n17153_0;
	wire [1:0] w_n17155_0;
	wire [1:0] w_n17157_0;
	wire [1:0] w_n17159_0;
	wire [1:0] w_n17162_0;
	wire [1:0] w_n17167_0;
	wire [2:0] w_n17169_0;
	wire [1:0] w_n17170_0;
	wire [1:0] w_n17174_0;
	wire [1:0] w_n17175_0;
	wire [1:0] w_n17177_0;
	wire [1:0] w_n17181_0;
	wire [1:0] w_n17183_0;
	wire [1:0] w_n17184_0;
	wire [2:0] w_n17185_0;
	wire [1:0] w_n17186_0;
	wire [1:0] w_n17190_0;
	wire [1:0] w_n17192_0;
	wire [1:0] w_n17194_0;
	wire [1:0] w_n17196_0;
	wire [1:0] w_n17199_0;
	wire [1:0] w_n17205_0;
	wire [2:0] w_n17207_0;
	wire [1:0] w_n17208_0;
	wire [1:0] w_n17213_0;
	wire [1:0] w_n17215_0;
	wire [1:0] w_n17217_0;
	wire [1:0] w_n17221_0;
	wire [1:0] w_n17223_0;
	wire [1:0] w_n17224_0;
	wire [2:0] w_n17225_0;
	wire [1:0] w_n17226_0;
	wire [1:0] w_n17232_0;
	wire [1:0] w_n17233_0;
	wire [1:0] w_n17235_0;
	wire [1:0] w_n17237_0;
	wire [1:0] w_n17239_0;
	wire [1:0] w_n17245_0;
	wire [1:0] w_n17247_0;
	wire [2:0] w_n17248_0;
	wire [1:0] w_n17251_0;
	wire [1:0] w_n17252_0;
	wire [2:0] w_n17253_0;
	wire [1:0] w_n17255_0;
	wire [1:0] w_n17259_0;
	wire [1:0] w_n17261_0;
	wire [1:0] w_n17262_0;
	wire [2:0] w_n17263_0;
	wire [1:0] w_n17264_0;
	wire [1:0] w_n17267_0;
	wire [1:0] w_n17273_0;
	wire [1:0] w_n17274_0;
	wire [1:0] w_n17276_0;
	wire [1:0] w_n17278_0;
	wire [1:0] w_n17280_0;
	wire [1:0] w_n17286_0;
	wire [1:0] w_n17288_0;
	wire [2:0] w_n17289_0;
	wire [1:0] w_n17292_0;
	wire [1:0] w_n17293_0;
	wire [2:0] w_n17294_0;
	wire [1:0] w_n17296_0;
	wire [1:0] w_n17300_0;
	wire [1:0] w_n17302_0;
	wire [1:0] w_n17303_0;
	wire [2:0] w_n17304_0;
	wire [1:0] w_n17305_0;
	wire [1:0] w_n17308_0;
	wire [1:0] w_n17314_0;
	wire [1:0] w_n17315_0;
	wire [1:0] w_n17317_0;
	wire [1:0] w_n17319_0;
	wire [1:0] w_n17321_0;
	wire [1:0] w_n17327_0;
	wire [1:0] w_n17329_0;
	wire [2:0] w_n17330_0;
	wire [1:0] w_n17333_0;
	wire [1:0] w_n17334_0;
	wire [2:0] w_n17335_0;
	wire [1:0] w_n17337_0;
	wire [1:0] w_n17341_0;
	wire [1:0] w_n17343_0;
	wire [1:0] w_n17344_0;
	wire [2:0] w_n17345_0;
	wire [1:0] w_n17346_0;
	wire [1:0] w_n17349_0;
	wire [1:0] w_n17355_0;
	wire [1:0] w_n17356_0;
	wire [1:0] w_n17358_0;
	wire [1:0] w_n17360_0;
	wire [1:0] w_n17362_0;
	wire [1:0] w_n17368_0;
	wire [1:0] w_n17370_0;
	wire [2:0] w_n17371_0;
	wire [1:0] w_n17374_0;
	wire [1:0] w_n17375_0;
	wire [2:0] w_n17376_0;
	wire [1:0] w_n17378_0;
	wire [1:0] w_n17382_0;
	wire [1:0] w_n17384_0;
	wire [1:0] w_n17385_0;
	wire [2:0] w_n17386_0;
	wire [1:0] w_n17387_0;
	wire [1:0] w_n17390_0;
	wire [1:0] w_n17396_0;
	wire [1:0] w_n17397_0;
	wire [1:0] w_n17399_0;
	wire [1:0] w_n17401_0;
	wire [1:0] w_n17403_0;
	wire [1:0] w_n17409_0;
	wire [1:0] w_n17411_0;
	wire [2:0] w_n17412_0;
	wire [1:0] w_n17415_0;
	wire [1:0] w_n17416_0;
	wire [2:0] w_n17417_0;
	wire [1:0] w_n17419_0;
	wire [1:0] w_n17423_0;
	wire [1:0] w_n17425_0;
	wire [1:0] w_n17426_0;
	wire [2:0] w_n17427_0;
	wire [1:0] w_n17428_0;
	wire [1:0] w_n17431_0;
	wire [1:0] w_n17437_0;
	wire [1:0] w_n17438_0;
	wire [1:0] w_n17440_0;
	wire [1:0] w_n17442_0;
	wire [1:0] w_n17444_0;
	wire [1:0] w_n17450_0;
	wire [1:0] w_n17452_0;
	wire [2:0] w_n17453_0;
	wire [1:0] w_n17456_0;
	wire [1:0] w_n17457_0;
	wire [2:0] w_n17458_0;
	wire [1:0] w_n17460_0;
	wire [1:0] w_n17464_0;
	wire [1:0] w_n17466_0;
	wire [1:0] w_n17467_0;
	wire [2:0] w_n17468_0;
	wire [1:0] w_n17469_0;
	wire [1:0] w_n17472_0;
	wire [1:0] w_n17478_0;
	wire [1:0] w_n17479_0;
	wire [1:0] w_n17481_0;
	wire [1:0] w_n17483_0;
	wire [1:0] w_n17485_0;
	wire [1:0] w_n17491_0;
	wire [1:0] w_n17493_0;
	wire [2:0] w_n17494_0;
	wire [1:0] w_n17497_0;
	wire [1:0] w_n17498_0;
	wire [2:0] w_n17499_0;
	wire [1:0] w_n17501_0;
	wire [1:0] w_n17505_0;
	wire [1:0] w_n17507_0;
	wire [1:0] w_n17508_0;
	wire [2:0] w_n17509_0;
	wire [1:0] w_n17510_0;
	wire [1:0] w_n17513_0;
	wire [1:0] w_n17519_0;
	wire [1:0] w_n17520_0;
	wire [1:0] w_n17522_0;
	wire [1:0] w_n17524_0;
	wire [1:0] w_n17526_0;
	wire [1:0] w_n17532_0;
	wire [1:0] w_n17534_0;
	wire [2:0] w_n17535_0;
	wire [1:0] w_n17538_0;
	wire [1:0] w_n17539_0;
	wire [2:0] w_n17540_0;
	wire [1:0] w_n17542_0;
	wire [1:0] w_n17546_0;
	wire [1:0] w_n17548_0;
	wire [1:0] w_n17549_0;
	wire [2:0] w_n17550_0;
	wire [1:0] w_n17551_0;
	wire [1:0] w_n17554_0;
	wire [1:0] w_n17560_0;
	wire [1:0] w_n17561_0;
	wire [1:0] w_n17563_0;
	wire [1:0] w_n17565_0;
	wire [1:0] w_n17567_0;
	wire [1:0] w_n17573_0;
	wire [1:0] w_n17575_0;
	wire [2:0] w_n17576_0;
	wire [1:0] w_n17579_0;
	wire [1:0] w_n17580_0;
	wire [2:0] w_n17581_0;
	wire [1:0] w_n17583_0;
	wire [1:0] w_n17587_0;
	wire [1:0] w_n17589_0;
	wire [1:0] w_n17590_0;
	wire [2:0] w_n17591_0;
	wire [1:0] w_n17592_0;
	wire [1:0] w_n17595_0;
	wire [1:0] w_n17601_0;
	wire [1:0] w_n17602_0;
	wire [1:0] w_n17604_0;
	wire [1:0] w_n17606_0;
	wire [1:0] w_n17608_0;
	wire [1:0] w_n17614_0;
	wire [1:0] w_n17616_0;
	wire [2:0] w_n17617_0;
	wire [1:0] w_n17620_0;
	wire [1:0] w_n17621_0;
	wire [2:0] w_n17622_0;
	wire [1:0] w_n17624_0;
	wire [1:0] w_n17626_0;
	wire [1:0] w_n17628_0;
	wire [1:0] w_n17634_0;
	wire [2:0] w_n17636_0;
	wire [1:0] w_n17637_0;
	wire [1:0] w_n17639_0;
	wire [1:0] w_n17641_0;
	wire [1:0] w_n17645_0;
	wire [1:0] w_n17647_0;
	wire [1:0] w_n17648_0;
	wire [1:0] w_n17649_0;
	wire [2:0] w_n17650_0;
	wire [1:0] w_n17653_0;
	wire [1:0] w_n17654_0;
	wire [2:0] w_n17655_0;
	wire [1:0] w_n17657_0;
	wire [1:0] w_n17661_0;
	wire [1:0] w_n17663_0;
	wire [1:0] w_n17664_0;
	wire [2:0] w_n17665_0;
	wire [1:0] w_n17666_0;
	wire [1:0] w_n17669_0;
	wire [1:0] w_n17675_0;
	wire [1:0] w_n17676_0;
	wire [1:0] w_n17678_0;
	wire [1:0] w_n17680_0;
	wire [1:0] w_n17682_0;
	wire [1:0] w_n17688_0;
	wire [2:0] w_n17690_0;
	wire [1:0] w_n17695_0;
	wire [2:0] w_n17697_0;
	wire [2:0] w_n17701_0;
	wire [1:0] w_n17702_0;
	wire [1:0] w_n17707_0;
	wire [2:0] w_n17708_0;
	wire [1:0] w_n17713_0;
	wire [1:0] w_n17720_0;
	wire [2:0] w_n17722_0;
	wire [1:0] w_n17722_1;
	wire [1:0] w_n17723_0;
	wire [2:0] w_n17726_0;
	wire [1:0] w_n17727_0;
	wire [1:0] w_n17728_0;
	wire [1:0] w_n17729_0;
	wire [1:0] w_n17731_0;
	wire [1:0] w_n17733_0;
	wire [1:0] w_n17735_0;
	wire [1:0] w_n17744_0;
	wire [2:0] w_n17746_0;
	wire [1:0] w_n17747_0;
	wire [1:0] w_n17751_0;
	wire [1:0] w_n17753_0;
	wire [1:0] w_n17755_0;
	wire [1:0] w_n17760_0;
	wire [1:0] w_n17762_0;
	wire [1:0] w_n17763_0;
	wire [2:0] w_n17764_0;
	wire [1:0] w_n17765_0;
	wire [1:0] w_n17770_0;
	wire [1:0] w_n17771_0;
	wire [1:0] w_n17773_0;
	wire [1:0] w_n17775_0;
	wire [1:0] w_n17778_0;
	wire [1:0] w_n17784_0;
	wire [2:0] w_n17786_0;
	wire [1:0] w_n17787_0;
	wire [1:0] w_n17791_0;
	wire [1:0] w_n17792_0;
	wire [1:0] w_n17794_0;
	wire [1:0] w_n17799_0;
	wire [1:0] w_n17801_0;
	wire [1:0] w_n17802_0;
	wire [2:0] w_n17803_0;
	wire [1:0] w_n17804_0;
	wire [1:0] w_n17808_0;
	wire [1:0] w_n17809_0;
	wire [1:0] w_n17811_0;
	wire [1:0] w_n17813_0;
	wire [1:0] w_n17816_0;
	wire [1:0] w_n17822_0;
	wire [1:0] w_n17824_0;
	wire [2:0] w_n17825_0;
	wire [1:0] w_n17829_0;
	wire [1:0] w_n17830_0;
	wire [2:0] w_n17831_0;
	wire [1:0] w_n17833_0;
	wire [1:0] w_n17838_0;
	wire [1:0] w_n17840_0;
	wire [1:0] w_n17841_0;
	wire [2:0] w_n17842_0;
	wire [1:0] w_n17843_0;
	wire [1:0] w_n17847_0;
	wire [1:0] w_n17853_0;
	wire [1:0] w_n17854_0;
	wire [1:0] w_n17856_0;
	wire [1:0] w_n17858_0;
	wire [1:0] w_n17861_0;
	wire [1:0] w_n17867_0;
	wire [1:0] w_n17869_0;
	wire [2:0] w_n17870_0;
	wire [1:0] w_n17874_0;
	wire [1:0] w_n17875_0;
	wire [2:0] w_n17876_0;
	wire [1:0] w_n17878_0;
	wire [1:0] w_n17883_0;
	wire [1:0] w_n17885_0;
	wire [1:0] w_n17886_0;
	wire [2:0] w_n17887_0;
	wire [1:0] w_n17888_0;
	wire [1:0] w_n17892_0;
	wire [1:0] w_n17898_0;
	wire [1:0] w_n17899_0;
	wire [1:0] w_n17901_0;
	wire [1:0] w_n17903_0;
	wire [1:0] w_n17906_0;
	wire [1:0] w_n17912_0;
	wire [1:0] w_n17914_0;
	wire [2:0] w_n17915_0;
	wire [1:0] w_n17919_0;
	wire [1:0] w_n17920_0;
	wire [2:0] w_n17921_0;
	wire [1:0] w_n17923_0;
	wire [1:0] w_n17928_0;
	wire [1:0] w_n17930_0;
	wire [1:0] w_n17931_0;
	wire [2:0] w_n17932_0;
	wire [1:0] w_n17933_0;
	wire [1:0] w_n17937_0;
	wire [1:0] w_n17943_0;
	wire [1:0] w_n17944_0;
	wire [1:0] w_n17946_0;
	wire [1:0] w_n17948_0;
	wire [1:0] w_n17951_0;
	wire [1:0] w_n17957_0;
	wire [1:0] w_n17959_0;
	wire [2:0] w_n17960_0;
	wire [1:0] w_n17964_0;
	wire [1:0] w_n17965_0;
	wire [2:0] w_n17966_0;
	wire [1:0] w_n17968_0;
	wire [1:0] w_n17973_0;
	wire [1:0] w_n17975_0;
	wire [1:0] w_n17976_0;
	wire [2:0] w_n17977_0;
	wire [1:0] w_n17978_0;
	wire [1:0] w_n17982_0;
	wire [1:0] w_n17988_0;
	wire [1:0] w_n17989_0;
	wire [1:0] w_n17991_0;
	wire [1:0] w_n17993_0;
	wire [1:0] w_n17996_0;
	wire [1:0] w_n18002_0;
	wire [1:0] w_n18004_0;
	wire [2:0] w_n18005_0;
	wire [1:0] w_n18009_0;
	wire [1:0] w_n18010_0;
	wire [2:0] w_n18011_0;
	wire [1:0] w_n18013_0;
	wire [1:0] w_n18018_0;
	wire [1:0] w_n18020_0;
	wire [1:0] w_n18021_0;
	wire [2:0] w_n18022_0;
	wire [1:0] w_n18023_0;
	wire [1:0] w_n18027_0;
	wire [1:0] w_n18033_0;
	wire [1:0] w_n18034_0;
	wire [1:0] w_n18036_0;
	wire [1:0] w_n18038_0;
	wire [1:0] w_n18041_0;
	wire [1:0] w_n18047_0;
	wire [1:0] w_n18049_0;
	wire [2:0] w_n18050_0;
	wire [1:0] w_n18054_0;
	wire [1:0] w_n18055_0;
	wire [2:0] w_n18056_0;
	wire [1:0] w_n18058_0;
	wire [1:0] w_n18063_0;
	wire [1:0] w_n18065_0;
	wire [1:0] w_n18066_0;
	wire [2:0] w_n18067_0;
	wire [1:0] w_n18068_0;
	wire [1:0] w_n18072_0;
	wire [1:0] w_n18078_0;
	wire [1:0] w_n18079_0;
	wire [1:0] w_n18081_0;
	wire [1:0] w_n18083_0;
	wire [1:0] w_n18086_0;
	wire [1:0] w_n18092_0;
	wire [1:0] w_n18094_0;
	wire [2:0] w_n18095_0;
	wire [1:0] w_n18099_0;
	wire [1:0] w_n18100_0;
	wire [2:0] w_n18101_0;
	wire [1:0] w_n18103_0;
	wire [1:0] w_n18108_0;
	wire [1:0] w_n18110_0;
	wire [1:0] w_n18111_0;
	wire [2:0] w_n18112_0;
	wire [1:0] w_n18113_0;
	wire [1:0] w_n18117_0;
	wire [1:0] w_n18123_0;
	wire [1:0] w_n18124_0;
	wire [1:0] w_n18126_0;
	wire [1:0] w_n18128_0;
	wire [1:0] w_n18131_0;
	wire [1:0] w_n18137_0;
	wire [1:0] w_n18139_0;
	wire [2:0] w_n18140_0;
	wire [1:0] w_n18144_0;
	wire [1:0] w_n18145_0;
	wire [2:0] w_n18146_0;
	wire [1:0] w_n18148_0;
	wire [1:0] w_n18153_0;
	wire [1:0] w_n18155_0;
	wire [1:0] w_n18156_0;
	wire [2:0] w_n18157_0;
	wire [1:0] w_n18158_0;
	wire [1:0] w_n18162_0;
	wire [1:0] w_n18168_0;
	wire [1:0] w_n18169_0;
	wire [1:0] w_n18171_0;
	wire [1:0] w_n18173_0;
	wire [1:0] w_n18176_0;
	wire [1:0] w_n18182_0;
	wire [1:0] w_n18184_0;
	wire [2:0] w_n18185_0;
	wire [1:0] w_n18189_0;
	wire [1:0] w_n18190_0;
	wire [2:0] w_n18191_0;
	wire [1:0] w_n18193_0;
	wire [1:0] w_n18198_0;
	wire [1:0] w_n18200_0;
	wire [1:0] w_n18201_0;
	wire [2:0] w_n18202_0;
	wire [1:0] w_n18203_0;
	wire [1:0] w_n18207_0;
	wire [1:0] w_n18213_0;
	wire [1:0] w_n18214_0;
	wire [1:0] w_n18216_0;
	wire [1:0] w_n18218_0;
	wire [1:0] w_n18221_0;
	wire [1:0] w_n18227_0;
	wire [1:0] w_n18229_0;
	wire [2:0] w_n18230_0;
	wire [1:0] w_n18234_0;
	wire [1:0] w_n18235_0;
	wire [2:0] w_n18236_0;
	wire [1:0] w_n18238_0;
	wire [1:0] w_n18243_0;
	wire [1:0] w_n18245_0;
	wire [1:0] w_n18246_0;
	wire [2:0] w_n18247_0;
	wire [1:0] w_n18248_0;
	wire [1:0] w_n18252_0;
	wire [1:0] w_n18258_0;
	wire [1:0] w_n18259_0;
	wire [1:0] w_n18261_0;
	wire [1:0] w_n18266_0;
	wire [1:0] w_n18268_0;
	wire [1:0] w_n18269_0;
	wire [2:0] w_n18270_0;
	wire [1:0] w_n18271_0;
	wire [1:0] w_n18274_0;
	wire [1:0] w_n18276_0;
	wire [1:0] w_n18278_0;
	wire [1:0] w_n18281_0;
	wire [1:0] w_n18287_0;
	wire [2:0] w_n18289_0;
	wire [1:0] w_n18290_0;
	wire [1:0] w_n18294_0;
	wire [1:0] w_n18300_0;
	wire [1:0] w_n18301_0;
	wire [1:0] w_n18303_0;
	wire [1:0] w_n18305_0;
	wire [1:0] w_n18308_0;
	wire [1:0] w_n18314_0;
	wire [1:0] w_n18316_0;
	wire [2:0] w_n18317_0;
	wire [1:0] w_n18321_0;
	wire [1:0] w_n18322_0;
	wire [2:0] w_n18323_0;
	wire [1:0] w_n18325_0;
	wire [1:0] w_n18330_0;
	wire [1:0] w_n18332_0;
	wire [1:0] w_n18333_0;
	wire [2:0] w_n18334_0;
	wire [2:0] w_n18334_1;
	wire [1:0] w_n18337_0;
	wire [2:0] w_n18338_0;
	wire [1:0] w_n18339_0;
	wire [1:0] w_n18340_0;
	wire [2:0] w_n18347_0;
	wire [1:0] w_n18348_0;
	wire [2:0] w_n18356_0;
	wire [2:0] w_n18356_1;
	wire [2:0] w_n18356_2;
	wire [2:0] w_n18356_3;
	wire [2:0] w_n18356_4;
	wire [2:0] w_n18356_5;
	wire [2:0] w_n18356_6;
	wire [2:0] w_n18356_7;
	wire [2:0] w_n18356_8;
	wire [2:0] w_n18356_9;
	wire [2:0] w_n18356_10;
	wire [2:0] w_n18356_11;
	wire [2:0] w_n18356_12;
	wire [2:0] w_n18356_13;
	wire [2:0] w_n18356_14;
	wire [2:0] w_n18356_15;
	wire [2:0] w_n18356_16;
	wire [2:0] w_n18356_17;
	wire [2:0] w_n18356_18;
	wire [1:0] w_n18356_19;
	wire [1:0] w_n18359_0;
	wire [2:0] w_n18360_0;
	wire [2:0] w_n18360_1;
	wire [2:0] w_n18360_2;
	wire [2:0] w_n18360_3;
	wire [2:0] w_n18362_0;
	wire [1:0] w_n18362_1;
	wire [2:0] w_n18363_0;
	wire [2:0] w_n18367_0;
	wire [1:0] w_n18368_0;
	wire [1:0] w_n18369_0;
	wire [1:0] w_n18370_0;
	wire [1:0] w_n18372_0;
	wire [1:0] w_n18374_0;
	wire [1:0] w_n18376_0;
	wire [1:0] w_n18381_0;
	wire [2:0] w_n18383_0;
	wire [1:0] w_n18384_0;
	wire [1:0] w_n18388_0;
	wire [1:0] w_n18389_0;
	wire [1:0] w_n18391_0;
	wire [1:0] w_n18395_0;
	wire [1:0] w_n18397_0;
	wire [1:0] w_n18398_0;
	wire [2:0] w_n18399_0;
	wire [1:0] w_n18400_0;
	wire [1:0] w_n18404_0;
	wire [1:0] w_n18406_0;
	wire [1:0] w_n18408_0;
	wire [1:0] w_n18410_0;
	wire [1:0] w_n18412_0;
	wire [1:0] w_n18418_0;
	wire [2:0] w_n18420_0;
	wire [1:0] w_n18421_0;
	wire [1:0] w_n18426_0;
	wire [1:0] w_n18428_0;
	wire [1:0] w_n18430_0;
	wire [1:0] w_n18434_0;
	wire [1:0] w_n18436_0;
	wire [1:0] w_n18437_0;
	wire [2:0] w_n18438_0;
	wire [1:0] w_n18439_0;
	wire [1:0] w_n18445_0;
	wire [1:0] w_n18446_0;
	wire [1:0] w_n18448_0;
	wire [1:0] w_n18450_0;
	wire [1:0] w_n18452_0;
	wire [1:0] w_n18458_0;
	wire [1:0] w_n18460_0;
	wire [2:0] w_n18461_0;
	wire [1:0] w_n18464_0;
	wire [1:0] w_n18465_0;
	wire [2:0] w_n18466_0;
	wire [1:0] w_n18468_0;
	wire [1:0] w_n18472_0;
	wire [1:0] w_n18474_0;
	wire [1:0] w_n18475_0;
	wire [2:0] w_n18476_0;
	wire [1:0] w_n18477_0;
	wire [1:0] w_n18480_0;
	wire [1:0] w_n18486_0;
	wire [1:0] w_n18487_0;
	wire [1:0] w_n18489_0;
	wire [1:0] w_n18491_0;
	wire [1:0] w_n18493_0;
	wire [1:0] w_n18499_0;
	wire [1:0] w_n18501_0;
	wire [2:0] w_n18502_0;
	wire [1:0] w_n18505_0;
	wire [1:0] w_n18506_0;
	wire [2:0] w_n18507_0;
	wire [1:0] w_n18509_0;
	wire [1:0] w_n18513_0;
	wire [1:0] w_n18515_0;
	wire [1:0] w_n18516_0;
	wire [2:0] w_n18517_0;
	wire [1:0] w_n18518_0;
	wire [1:0] w_n18521_0;
	wire [1:0] w_n18527_0;
	wire [1:0] w_n18528_0;
	wire [1:0] w_n18530_0;
	wire [1:0] w_n18532_0;
	wire [1:0] w_n18534_0;
	wire [1:0] w_n18540_0;
	wire [1:0] w_n18542_0;
	wire [2:0] w_n18543_0;
	wire [1:0] w_n18546_0;
	wire [1:0] w_n18547_0;
	wire [2:0] w_n18548_0;
	wire [1:0] w_n18550_0;
	wire [1:0] w_n18554_0;
	wire [1:0] w_n18556_0;
	wire [1:0] w_n18557_0;
	wire [2:0] w_n18558_0;
	wire [1:0] w_n18559_0;
	wire [1:0] w_n18562_0;
	wire [1:0] w_n18568_0;
	wire [1:0] w_n18569_0;
	wire [1:0] w_n18571_0;
	wire [1:0] w_n18573_0;
	wire [1:0] w_n18575_0;
	wire [1:0] w_n18581_0;
	wire [1:0] w_n18583_0;
	wire [2:0] w_n18584_0;
	wire [1:0] w_n18587_0;
	wire [1:0] w_n18588_0;
	wire [2:0] w_n18589_0;
	wire [1:0] w_n18591_0;
	wire [1:0] w_n18595_0;
	wire [1:0] w_n18597_0;
	wire [1:0] w_n18598_0;
	wire [2:0] w_n18599_0;
	wire [1:0] w_n18600_0;
	wire [1:0] w_n18603_0;
	wire [1:0] w_n18609_0;
	wire [1:0] w_n18610_0;
	wire [1:0] w_n18612_0;
	wire [1:0] w_n18614_0;
	wire [1:0] w_n18616_0;
	wire [1:0] w_n18622_0;
	wire [1:0] w_n18624_0;
	wire [2:0] w_n18625_0;
	wire [1:0] w_n18628_0;
	wire [1:0] w_n18629_0;
	wire [2:0] w_n18630_0;
	wire [1:0] w_n18632_0;
	wire [1:0] w_n18636_0;
	wire [1:0] w_n18638_0;
	wire [1:0] w_n18639_0;
	wire [2:0] w_n18640_0;
	wire [1:0] w_n18641_0;
	wire [1:0] w_n18644_0;
	wire [1:0] w_n18650_0;
	wire [1:0] w_n18651_0;
	wire [1:0] w_n18653_0;
	wire [1:0] w_n18655_0;
	wire [1:0] w_n18657_0;
	wire [1:0] w_n18663_0;
	wire [1:0] w_n18665_0;
	wire [2:0] w_n18666_0;
	wire [1:0] w_n18669_0;
	wire [1:0] w_n18670_0;
	wire [2:0] w_n18671_0;
	wire [1:0] w_n18673_0;
	wire [1:0] w_n18677_0;
	wire [1:0] w_n18679_0;
	wire [1:0] w_n18680_0;
	wire [2:0] w_n18681_0;
	wire [1:0] w_n18682_0;
	wire [1:0] w_n18685_0;
	wire [1:0] w_n18691_0;
	wire [1:0] w_n18692_0;
	wire [1:0] w_n18694_0;
	wire [1:0] w_n18696_0;
	wire [1:0] w_n18698_0;
	wire [1:0] w_n18704_0;
	wire [1:0] w_n18706_0;
	wire [2:0] w_n18707_0;
	wire [1:0] w_n18710_0;
	wire [1:0] w_n18711_0;
	wire [2:0] w_n18712_0;
	wire [1:0] w_n18714_0;
	wire [1:0] w_n18718_0;
	wire [1:0] w_n18720_0;
	wire [1:0] w_n18721_0;
	wire [2:0] w_n18722_0;
	wire [1:0] w_n18723_0;
	wire [1:0] w_n18726_0;
	wire [1:0] w_n18732_0;
	wire [1:0] w_n18733_0;
	wire [1:0] w_n18735_0;
	wire [1:0] w_n18737_0;
	wire [1:0] w_n18739_0;
	wire [1:0] w_n18745_0;
	wire [1:0] w_n18747_0;
	wire [2:0] w_n18748_0;
	wire [1:0] w_n18751_0;
	wire [1:0] w_n18752_0;
	wire [2:0] w_n18753_0;
	wire [1:0] w_n18755_0;
	wire [1:0] w_n18759_0;
	wire [1:0] w_n18761_0;
	wire [1:0] w_n18762_0;
	wire [2:0] w_n18763_0;
	wire [1:0] w_n18764_0;
	wire [1:0] w_n18767_0;
	wire [1:0] w_n18773_0;
	wire [1:0] w_n18774_0;
	wire [1:0] w_n18776_0;
	wire [1:0] w_n18778_0;
	wire [1:0] w_n18780_0;
	wire [1:0] w_n18786_0;
	wire [1:0] w_n18788_0;
	wire [2:0] w_n18789_0;
	wire [1:0] w_n18792_0;
	wire [1:0] w_n18793_0;
	wire [2:0] w_n18794_0;
	wire [1:0] w_n18796_0;
	wire [1:0] w_n18800_0;
	wire [1:0] w_n18802_0;
	wire [1:0] w_n18803_0;
	wire [2:0] w_n18804_0;
	wire [1:0] w_n18805_0;
	wire [1:0] w_n18808_0;
	wire [1:0] w_n18814_0;
	wire [1:0] w_n18815_0;
	wire [1:0] w_n18817_0;
	wire [1:0] w_n18819_0;
	wire [1:0] w_n18821_0;
	wire [1:0] w_n18827_0;
	wire [1:0] w_n18829_0;
	wire [2:0] w_n18830_0;
	wire [1:0] w_n18833_0;
	wire [1:0] w_n18834_0;
	wire [2:0] w_n18835_0;
	wire [1:0] w_n18837_0;
	wire [1:0] w_n18841_0;
	wire [1:0] w_n18843_0;
	wire [1:0] w_n18844_0;
	wire [2:0] w_n18845_0;
	wire [1:0] w_n18846_0;
	wire [1:0] w_n18849_0;
	wire [1:0] w_n18855_0;
	wire [1:0] w_n18856_0;
	wire [1:0] w_n18858_0;
	wire [1:0] w_n18860_0;
	wire [1:0] w_n18862_0;
	wire [1:0] w_n18868_0;
	wire [1:0] w_n18870_0;
	wire [2:0] w_n18871_0;
	wire [1:0] w_n18874_0;
	wire [1:0] w_n18875_0;
	wire [2:0] w_n18876_0;
	wire [1:0] w_n18878_0;
	wire [1:0] w_n18880_0;
	wire [1:0] w_n18882_0;
	wire [1:0] w_n18888_0;
	wire [2:0] w_n18890_0;
	wire [1:0] w_n18891_0;
	wire [1:0] w_n18894_0;
	wire [1:0] w_n18896_0;
	wire [1:0] w_n18900_0;
	wire [1:0] w_n18902_0;
	wire [1:0] w_n18903_0;
	wire [1:0] w_n18904_0;
	wire [2:0] w_n18905_0;
	wire [1:0] w_n18908_0;
	wire [1:0] w_n18909_0;
	wire [2:0] w_n18910_0;
	wire [1:0] w_n18912_0;
	wire [1:0] w_n18916_0;
	wire [1:0] w_n18918_0;
	wire [1:0] w_n18919_0;
	wire [2:0] w_n18920_0;
	wire [1:0] w_n18924_0;
	wire [1:0] w_n18930_0;
	wire [2:0] w_n18932_0;
	wire [1:0] w_n18934_0;
	wire [2:0] w_n18939_0;
	wire [1:0] w_n18940_0;
	wire [1:0] w_n18942_0;
	wire [1:0] w_n18948_0;
	wire [1:0] w_n18958_0;
	wire [2:0] w_n18961_0;
	wire [1:0] w_n18961_1;
	wire [1:0] w_n18962_0;
	wire [2:0] w_n18965_0;
	wire [1:0] w_n18966_0;
	wire [1:0] w_n18967_0;
	wire [1:0] w_n18968_0;
	wire [1:0] w_n18970_0;
	wire [1:0] w_n18972_0;
	wire [1:0] w_n18974_0;
	wire [2:0] w_n18976_0;
	wire [2:0] w_n18976_1;
	wire [2:0] w_n18976_2;
	wire [1:0] w_n18979_0;
	wire [2:0] w_n18981_0;
	wire [1:0] w_n18982_0;
	wire [1:0] w_n18986_0;
	wire [1:0] w_n18988_0;
	wire [1:0] w_n18990_0;
	wire [1:0] w_n18995_0;
	wire [1:0] w_n18997_0;
	wire [1:0] w_n18998_0;
	wire [2:0] w_n18999_0;
	wire [1:0] w_n19000_0;
	wire [1:0] w_n19005_0;
	wire [1:0] w_n19006_0;
	wire [1:0] w_n19008_0;
	wire [1:0] w_n19010_0;
	wire [1:0] w_n19013_0;
	wire [1:0] w_n19019_0;
	wire [2:0] w_n19021_0;
	wire [1:0] w_n19022_0;
	wire [1:0] w_n19026_0;
	wire [1:0] w_n19027_0;
	wire [1:0] w_n19029_0;
	wire [1:0] w_n19034_0;
	wire [1:0] w_n19036_0;
	wire [1:0] w_n19037_0;
	wire [2:0] w_n19038_0;
	wire [1:0] w_n19039_0;
	wire [1:0] w_n19043_0;
	wire [1:0] w_n19044_0;
	wire [1:0] w_n19046_0;
	wire [1:0] w_n19048_0;
	wire [1:0] w_n19051_0;
	wire [1:0] w_n19057_0;
	wire [1:0] w_n19059_0;
	wire [2:0] w_n19060_0;
	wire [1:0] w_n19064_0;
	wire [1:0] w_n19065_0;
	wire [2:0] w_n19066_0;
	wire [1:0] w_n19068_0;
	wire [1:0] w_n19073_0;
	wire [1:0] w_n19075_0;
	wire [1:0] w_n19076_0;
	wire [2:0] w_n19077_0;
	wire [1:0] w_n19078_0;
	wire [1:0] w_n19082_0;
	wire [1:0] w_n19088_0;
	wire [1:0] w_n19089_0;
	wire [1:0] w_n19091_0;
	wire [1:0] w_n19093_0;
	wire [1:0] w_n19096_0;
	wire [1:0] w_n19102_0;
	wire [1:0] w_n19104_0;
	wire [2:0] w_n19105_0;
	wire [1:0] w_n19109_0;
	wire [1:0] w_n19110_0;
	wire [2:0] w_n19111_0;
	wire [1:0] w_n19113_0;
	wire [1:0] w_n19118_0;
	wire [1:0] w_n19120_0;
	wire [1:0] w_n19121_0;
	wire [2:0] w_n19122_0;
	wire [1:0] w_n19123_0;
	wire [1:0] w_n19127_0;
	wire [1:0] w_n19133_0;
	wire [1:0] w_n19134_0;
	wire [1:0] w_n19136_0;
	wire [1:0] w_n19138_0;
	wire [1:0] w_n19141_0;
	wire [1:0] w_n19147_0;
	wire [1:0] w_n19149_0;
	wire [2:0] w_n19150_0;
	wire [1:0] w_n19154_0;
	wire [1:0] w_n19155_0;
	wire [2:0] w_n19156_0;
	wire [1:0] w_n19158_0;
	wire [1:0] w_n19163_0;
	wire [1:0] w_n19165_0;
	wire [1:0] w_n19166_0;
	wire [2:0] w_n19167_0;
	wire [1:0] w_n19168_0;
	wire [1:0] w_n19172_0;
	wire [1:0] w_n19178_0;
	wire [1:0] w_n19179_0;
	wire [1:0] w_n19181_0;
	wire [1:0] w_n19183_0;
	wire [1:0] w_n19186_0;
	wire [1:0] w_n19192_0;
	wire [1:0] w_n19194_0;
	wire [2:0] w_n19195_0;
	wire [1:0] w_n19199_0;
	wire [1:0] w_n19200_0;
	wire [2:0] w_n19201_0;
	wire [1:0] w_n19203_0;
	wire [1:0] w_n19208_0;
	wire [1:0] w_n19210_0;
	wire [1:0] w_n19211_0;
	wire [2:0] w_n19212_0;
	wire [1:0] w_n19213_0;
	wire [1:0] w_n19217_0;
	wire [1:0] w_n19223_0;
	wire [1:0] w_n19224_0;
	wire [1:0] w_n19226_0;
	wire [1:0] w_n19228_0;
	wire [1:0] w_n19231_0;
	wire [1:0] w_n19237_0;
	wire [1:0] w_n19239_0;
	wire [2:0] w_n19240_0;
	wire [1:0] w_n19244_0;
	wire [1:0] w_n19245_0;
	wire [2:0] w_n19246_0;
	wire [1:0] w_n19248_0;
	wire [1:0] w_n19253_0;
	wire [1:0] w_n19255_0;
	wire [1:0] w_n19256_0;
	wire [2:0] w_n19257_0;
	wire [1:0] w_n19258_0;
	wire [1:0] w_n19262_0;
	wire [1:0] w_n19268_0;
	wire [1:0] w_n19269_0;
	wire [1:0] w_n19271_0;
	wire [1:0] w_n19273_0;
	wire [1:0] w_n19276_0;
	wire [1:0] w_n19282_0;
	wire [1:0] w_n19284_0;
	wire [2:0] w_n19285_0;
	wire [1:0] w_n19289_0;
	wire [1:0] w_n19290_0;
	wire [2:0] w_n19291_0;
	wire [1:0] w_n19293_0;
	wire [1:0] w_n19298_0;
	wire [1:0] w_n19300_0;
	wire [1:0] w_n19301_0;
	wire [2:0] w_n19302_0;
	wire [1:0] w_n19303_0;
	wire [1:0] w_n19307_0;
	wire [1:0] w_n19313_0;
	wire [1:0] w_n19314_0;
	wire [1:0] w_n19316_0;
	wire [1:0] w_n19318_0;
	wire [1:0] w_n19321_0;
	wire [1:0] w_n19327_0;
	wire [1:0] w_n19329_0;
	wire [2:0] w_n19330_0;
	wire [1:0] w_n19334_0;
	wire [1:0] w_n19335_0;
	wire [2:0] w_n19336_0;
	wire [1:0] w_n19338_0;
	wire [1:0] w_n19343_0;
	wire [1:0] w_n19345_0;
	wire [1:0] w_n19346_0;
	wire [2:0] w_n19347_0;
	wire [1:0] w_n19348_0;
	wire [1:0] w_n19352_0;
	wire [1:0] w_n19358_0;
	wire [1:0] w_n19359_0;
	wire [1:0] w_n19361_0;
	wire [1:0] w_n19363_0;
	wire [1:0] w_n19366_0;
	wire [1:0] w_n19372_0;
	wire [1:0] w_n19374_0;
	wire [2:0] w_n19375_0;
	wire [1:0] w_n19379_0;
	wire [1:0] w_n19380_0;
	wire [2:0] w_n19381_0;
	wire [1:0] w_n19383_0;
	wire [1:0] w_n19388_0;
	wire [1:0] w_n19390_0;
	wire [1:0] w_n19391_0;
	wire [2:0] w_n19392_0;
	wire [1:0] w_n19393_0;
	wire [1:0] w_n19397_0;
	wire [1:0] w_n19403_0;
	wire [1:0] w_n19404_0;
	wire [1:0] w_n19406_0;
	wire [1:0] w_n19408_0;
	wire [1:0] w_n19411_0;
	wire [1:0] w_n19417_0;
	wire [1:0] w_n19419_0;
	wire [2:0] w_n19420_0;
	wire [1:0] w_n19424_0;
	wire [1:0] w_n19425_0;
	wire [2:0] w_n19426_0;
	wire [1:0] w_n19428_0;
	wire [1:0] w_n19433_0;
	wire [1:0] w_n19435_0;
	wire [1:0] w_n19436_0;
	wire [2:0] w_n19437_0;
	wire [1:0] w_n19438_0;
	wire [1:0] w_n19442_0;
	wire [1:0] w_n19448_0;
	wire [1:0] w_n19449_0;
	wire [1:0] w_n19451_0;
	wire [1:0] w_n19453_0;
	wire [1:0] w_n19456_0;
	wire [1:0] w_n19462_0;
	wire [1:0] w_n19464_0;
	wire [2:0] w_n19465_0;
	wire [1:0] w_n19469_0;
	wire [1:0] w_n19470_0;
	wire [2:0] w_n19471_0;
	wire [1:0] w_n19473_0;
	wire [1:0] w_n19478_0;
	wire [1:0] w_n19480_0;
	wire [1:0] w_n19481_0;
	wire [2:0] w_n19482_0;
	wire [1:0] w_n19483_0;
	wire [1:0] w_n19487_0;
	wire [1:0] w_n19493_0;
	wire [1:0] w_n19494_0;
	wire [1:0] w_n19496_0;
	wire [1:0] w_n19498_0;
	wire [1:0] w_n19501_0;
	wire [1:0] w_n19507_0;
	wire [1:0] w_n19509_0;
	wire [2:0] w_n19510_0;
	wire [1:0] w_n19514_0;
	wire [1:0] w_n19515_0;
	wire [2:0] w_n19516_0;
	wire [1:0] w_n19518_0;
	wire [1:0] w_n19523_0;
	wire [1:0] w_n19525_0;
	wire [1:0] w_n19526_0;
	wire [2:0] w_n19527_0;
	wire [1:0] w_n19528_0;
	wire [1:0] w_n19532_0;
	wire [1:0] w_n19538_0;
	wire [1:0] w_n19539_0;
	wire [1:0] w_n19541_0;
	wire [1:0] w_n19546_0;
	wire [1:0] w_n19548_0;
	wire [1:0] w_n19549_0;
	wire [2:0] w_n19550_0;
	wire [1:0] w_n19551_0;
	wire [1:0] w_n19553_0;
	wire [1:0] w_n19555_0;
	wire [1:0] w_n19557_0;
	wire [1:0] w_n19560_0;
	wire [1:0] w_n19566_0;
	wire [2:0] w_n19568_0;
	wire [1:0] w_n19569_0;
	wire [1:0] w_n19573_0;
	wire [1:0] w_n19579_0;
	wire [1:0] w_n19580_0;
	wire [1:0] w_n19582_0;
	wire [1:0] w_n19584_0;
	wire [1:0] w_n19587_0;
	wire [1:0] w_n19593_0;
	wire [2:0] w_n19595_0;
	wire [2:0] w_n19595_1;
	wire [1:0] w_n19598_0;
	wire [2:0] w_n19599_0;
	wire [1:0] w_n19600_0;
	wire [2:0] w_n19607_0;
	wire [1:0] w_n19608_0;
	wire [2:0] w_n19616_0;
	wire [2:0] w_n19616_1;
	wire [2:0] w_n19616_2;
	wire [2:0] w_n19616_3;
	wire [2:0] w_n19616_4;
	wire [2:0] w_n19616_5;
	wire [2:0] w_n19616_6;
	wire [2:0] w_n19616_7;
	wire [2:0] w_n19616_8;
	wire [2:0] w_n19616_9;
	wire [2:0] w_n19616_10;
	wire [2:0] w_n19616_11;
	wire [2:0] w_n19616_12;
	wire [2:0] w_n19616_13;
	wire [2:0] w_n19616_14;
	wire [2:0] w_n19616_15;
	wire [2:0] w_n19616_16;
	wire [2:0] w_n19616_17;
	wire [2:0] w_n19616_18;
	wire [1:0] w_n19620_0;
	wire [2:0] w_n19622_0;
	wire [1:0] w_n19622_1;
	wire [2:0] w_n19623_0;
	wire [2:0] w_n19627_0;
	wire [1:0] w_n19628_0;
	wire [1:0] w_n19629_0;
	wire [1:0] w_n19630_0;
	wire [1:0] w_n19632_0;
	wire [1:0] w_n19634_0;
	wire [1:0] w_n19636_0;
	wire [1:0] w_n19641_0;
	wire [2:0] w_n19643_0;
	wire [1:0] w_n19644_0;
	wire [1:0] w_n19648_0;
	wire [1:0] w_n19649_0;
	wire [1:0] w_n19651_0;
	wire [1:0] w_n19655_0;
	wire [1:0] w_n19657_0;
	wire [1:0] w_n19658_0;
	wire [2:0] w_n19659_0;
	wire [1:0] w_n19660_0;
	wire [1:0] w_n19664_0;
	wire [1:0] w_n19666_0;
	wire [1:0] w_n19668_0;
	wire [1:0] w_n19670_0;
	wire [1:0] w_n19672_0;
	wire [1:0] w_n19678_0;
	wire [2:0] w_n19680_0;
	wire [1:0] w_n19681_0;
	wire [1:0] w_n19686_0;
	wire [1:0] w_n19688_0;
	wire [1:0] w_n19690_0;
	wire [1:0] w_n19694_0;
	wire [1:0] w_n19696_0;
	wire [1:0] w_n19697_0;
	wire [2:0] w_n19698_0;
	wire [1:0] w_n19699_0;
	wire [1:0] w_n19705_0;
	wire [1:0] w_n19706_0;
	wire [1:0] w_n19708_0;
	wire [1:0] w_n19710_0;
	wire [1:0] w_n19712_0;
	wire [1:0] w_n19718_0;
	wire [1:0] w_n19720_0;
	wire [2:0] w_n19721_0;
	wire [1:0] w_n19724_0;
	wire [1:0] w_n19725_0;
	wire [2:0] w_n19726_0;
	wire [1:0] w_n19728_0;
	wire [1:0] w_n19732_0;
	wire [1:0] w_n19734_0;
	wire [1:0] w_n19735_0;
	wire [2:0] w_n19736_0;
	wire [1:0] w_n19737_0;
	wire [1:0] w_n19740_0;
	wire [1:0] w_n19746_0;
	wire [1:0] w_n19747_0;
	wire [1:0] w_n19749_0;
	wire [1:0] w_n19751_0;
	wire [1:0] w_n19753_0;
	wire [1:0] w_n19759_0;
	wire [1:0] w_n19761_0;
	wire [2:0] w_n19762_0;
	wire [1:0] w_n19765_0;
	wire [1:0] w_n19766_0;
	wire [2:0] w_n19767_0;
	wire [1:0] w_n19769_0;
	wire [1:0] w_n19773_0;
	wire [1:0] w_n19775_0;
	wire [1:0] w_n19776_0;
	wire [2:0] w_n19777_0;
	wire [1:0] w_n19778_0;
	wire [1:0] w_n19781_0;
	wire [1:0] w_n19787_0;
	wire [1:0] w_n19788_0;
	wire [1:0] w_n19790_0;
	wire [1:0] w_n19792_0;
	wire [1:0] w_n19794_0;
	wire [1:0] w_n19800_0;
	wire [1:0] w_n19802_0;
	wire [2:0] w_n19803_0;
	wire [1:0] w_n19806_0;
	wire [1:0] w_n19807_0;
	wire [2:0] w_n19808_0;
	wire [1:0] w_n19810_0;
	wire [1:0] w_n19814_0;
	wire [1:0] w_n19816_0;
	wire [1:0] w_n19817_0;
	wire [2:0] w_n19818_0;
	wire [1:0] w_n19819_0;
	wire [1:0] w_n19822_0;
	wire [1:0] w_n19828_0;
	wire [1:0] w_n19829_0;
	wire [1:0] w_n19831_0;
	wire [1:0] w_n19833_0;
	wire [1:0] w_n19835_0;
	wire [1:0] w_n19841_0;
	wire [1:0] w_n19843_0;
	wire [2:0] w_n19844_0;
	wire [1:0] w_n19847_0;
	wire [1:0] w_n19848_0;
	wire [2:0] w_n19849_0;
	wire [1:0] w_n19851_0;
	wire [1:0] w_n19855_0;
	wire [1:0] w_n19857_0;
	wire [1:0] w_n19858_0;
	wire [2:0] w_n19859_0;
	wire [1:0] w_n19860_0;
	wire [1:0] w_n19863_0;
	wire [1:0] w_n19869_0;
	wire [1:0] w_n19870_0;
	wire [1:0] w_n19872_0;
	wire [1:0] w_n19874_0;
	wire [1:0] w_n19876_0;
	wire [1:0] w_n19882_0;
	wire [1:0] w_n19884_0;
	wire [2:0] w_n19885_0;
	wire [1:0] w_n19888_0;
	wire [1:0] w_n19889_0;
	wire [2:0] w_n19890_0;
	wire [1:0] w_n19892_0;
	wire [1:0] w_n19896_0;
	wire [1:0] w_n19898_0;
	wire [1:0] w_n19899_0;
	wire [2:0] w_n19900_0;
	wire [1:0] w_n19901_0;
	wire [1:0] w_n19904_0;
	wire [1:0] w_n19910_0;
	wire [1:0] w_n19911_0;
	wire [1:0] w_n19913_0;
	wire [1:0] w_n19915_0;
	wire [1:0] w_n19917_0;
	wire [1:0] w_n19923_0;
	wire [1:0] w_n19925_0;
	wire [2:0] w_n19926_0;
	wire [1:0] w_n19929_0;
	wire [1:0] w_n19930_0;
	wire [2:0] w_n19931_0;
	wire [1:0] w_n19933_0;
	wire [1:0] w_n19937_0;
	wire [1:0] w_n19939_0;
	wire [1:0] w_n19940_0;
	wire [2:0] w_n19941_0;
	wire [1:0] w_n19942_0;
	wire [1:0] w_n19945_0;
	wire [1:0] w_n19951_0;
	wire [1:0] w_n19952_0;
	wire [1:0] w_n19954_0;
	wire [1:0] w_n19956_0;
	wire [1:0] w_n19958_0;
	wire [1:0] w_n19964_0;
	wire [1:0] w_n19966_0;
	wire [2:0] w_n19967_0;
	wire [1:0] w_n19970_0;
	wire [1:0] w_n19971_0;
	wire [2:0] w_n19972_0;
	wire [1:0] w_n19974_0;
	wire [1:0] w_n19978_0;
	wire [1:0] w_n19980_0;
	wire [1:0] w_n19981_0;
	wire [2:0] w_n19982_0;
	wire [1:0] w_n19983_0;
	wire [1:0] w_n19986_0;
	wire [1:0] w_n19992_0;
	wire [1:0] w_n19993_0;
	wire [1:0] w_n19995_0;
	wire [1:0] w_n19997_0;
	wire [1:0] w_n19999_0;
	wire [1:0] w_n20005_0;
	wire [1:0] w_n20007_0;
	wire [2:0] w_n20008_0;
	wire [1:0] w_n20011_0;
	wire [1:0] w_n20012_0;
	wire [2:0] w_n20013_0;
	wire [1:0] w_n20015_0;
	wire [1:0] w_n20019_0;
	wire [1:0] w_n20021_0;
	wire [1:0] w_n20022_0;
	wire [2:0] w_n20023_0;
	wire [1:0] w_n20024_0;
	wire [1:0] w_n20027_0;
	wire [1:0] w_n20033_0;
	wire [1:0] w_n20034_0;
	wire [1:0] w_n20036_0;
	wire [1:0] w_n20038_0;
	wire [1:0] w_n20040_0;
	wire [1:0] w_n20046_0;
	wire [1:0] w_n20048_0;
	wire [2:0] w_n20049_0;
	wire [1:0] w_n20052_0;
	wire [1:0] w_n20053_0;
	wire [2:0] w_n20054_0;
	wire [1:0] w_n20056_0;
	wire [1:0] w_n20060_0;
	wire [1:0] w_n20062_0;
	wire [1:0] w_n20063_0;
	wire [2:0] w_n20064_0;
	wire [1:0] w_n20065_0;
	wire [1:0] w_n20068_0;
	wire [1:0] w_n20074_0;
	wire [1:0] w_n20075_0;
	wire [1:0] w_n20077_0;
	wire [1:0] w_n20079_0;
	wire [1:0] w_n20081_0;
	wire [1:0] w_n20087_0;
	wire [1:0] w_n20089_0;
	wire [2:0] w_n20090_0;
	wire [1:0] w_n20093_0;
	wire [1:0] w_n20094_0;
	wire [2:0] w_n20095_0;
	wire [1:0] w_n20097_0;
	wire [1:0] w_n20101_0;
	wire [1:0] w_n20103_0;
	wire [1:0] w_n20104_0;
	wire [2:0] w_n20105_0;
	wire [1:0] w_n20106_0;
	wire [1:0] w_n20109_0;
	wire [1:0] w_n20115_0;
	wire [1:0] w_n20116_0;
	wire [1:0] w_n20118_0;
	wire [1:0] w_n20120_0;
	wire [1:0] w_n20122_0;
	wire [1:0] w_n20128_0;
	wire [1:0] w_n20130_0;
	wire [2:0] w_n20131_0;
	wire [1:0] w_n20134_0;
	wire [1:0] w_n20135_0;
	wire [2:0] w_n20136_0;
	wire [1:0] w_n20138_0;
	wire [1:0] w_n20142_0;
	wire [1:0] w_n20144_0;
	wire [1:0] w_n20145_0;
	wire [2:0] w_n20146_0;
	wire [1:0] w_n20147_0;
	wire [1:0] w_n20150_0;
	wire [1:0] w_n20156_0;
	wire [1:0] w_n20157_0;
	wire [1:0] w_n20159_0;
	wire [1:0] w_n20161_0;
	wire [1:0] w_n20163_0;
	wire [1:0] w_n20169_0;
	wire [1:0] w_n20171_0;
	wire [2:0] w_n20172_0;
	wire [1:0] w_n20175_0;
	wire [1:0] w_n20176_0;
	wire [2:0] w_n20177_0;
	wire [1:0] w_n20179_0;
	wire [1:0] w_n20181_0;
	wire [1:0] w_n20183_0;
	wire [1:0] w_n20189_0;
	wire [2:0] w_n20191_0;
	wire [1:0] w_n20192_0;
	wire [1:0] w_n20194_0;
	wire [1:0] w_n20196_0;
	wire [1:0] w_n20200_0;
	wire [1:0] w_n20202_0;
	wire [1:0] w_n20203_0;
	wire [2:0] w_n20204_0;
	wire [1:0] w_n20209_0;
	wire [2:0] w_n20211_0;
	wire [2:0] w_n20215_0;
	wire [1:0] w_n20217_0;
	wire [1:0] w_n20223_0;
	wire [1:0] w_n20234_0;
	wire [1:0] w_n20236_0;
	wire [1:0] w_n20237_0;
	wire [2:0] w_n20240_0;
	wire [1:0] w_n20241_0;
	wire [1:0] w_n20242_0;
	wire [1:0] w_n20243_0;
	wire [1:0] w_n20245_0;
	wire [1:0] w_n20247_0;
	wire [1:0] w_n20249_0;
	wire [2:0] w_n20251_0;
	wire [1:0] w_n20251_1;
	wire [1:0] w_n20254_0;
	wire [2:0] w_n20256_0;
	wire [1:0] w_n20257_0;
	wire [1:0] w_n20262_0;
	wire [1:0] w_n20263_0;
	wire [1:0] w_n20265_0;
	wire [1:0] w_n20269_0;
	wire [1:0] w_n20272_0;
	wire [1:0] w_n20273_0;
	wire [2:0] w_n20274_0;
	wire [1:0] w_n20275_0;
	wire [1:0] w_n20280_0;
	wire [1:0] w_n20281_0;
	wire [1:0] w_n20283_0;
	wire [1:0] w_n20285_0;
	wire [1:0] w_n20288_0;
	wire [1:0] w_n20294_0;
	wire [2:0] w_n20296_0;
	wire [1:0] w_n20297_0;
	wire [1:0] w_n20301_0;
	wire [1:0] w_n20302_0;
	wire [1:0] w_n20304_0;
	wire [1:0] w_n20308_0;
	wire [1:0] w_n20311_0;
	wire [1:0] w_n20312_0;
	wire [2:0] w_n20313_0;
	wire [1:0] w_n20314_0;
	wire [1:0] w_n20318_0;
	wire [1:0] w_n20319_0;
	wire [1:0] w_n20321_0;
	wire [1:0] w_n20323_0;
	wire [1:0] w_n20326_0;
	wire [1:0] w_n20332_0;
	wire [1:0] w_n20334_0;
	wire [2:0] w_n20335_0;
	wire [1:0] w_n20338_0;
	wire [1:0] w_n20340_0;
	wire [2:0] w_n20341_0;
	wire [1:0] w_n20343_0;
	wire [1:0] w_n20347_0;
	wire [1:0] w_n20350_0;
	wire [1:0] w_n20351_0;
	wire [2:0] w_n20352_0;
	wire [1:0] w_n20353_0;
	wire [1:0] w_n20357_0;
	wire [1:0] w_n20363_0;
	wire [1:0] w_n20364_0;
	wire [1:0] w_n20366_0;
	wire [1:0] w_n20368_0;
	wire [1:0] w_n20371_0;
	wire [1:0] w_n20377_0;
	wire [1:0] w_n20379_0;
	wire [2:0] w_n20380_0;
	wire [1:0] w_n20383_0;
	wire [1:0] w_n20385_0;
	wire [2:0] w_n20386_0;
	wire [1:0] w_n20388_0;
	wire [1:0] w_n20392_0;
	wire [1:0] w_n20395_0;
	wire [1:0] w_n20396_0;
	wire [2:0] w_n20397_0;
	wire [1:0] w_n20398_0;
	wire [1:0] w_n20402_0;
	wire [1:0] w_n20408_0;
	wire [1:0] w_n20409_0;
	wire [1:0] w_n20411_0;
	wire [1:0] w_n20413_0;
	wire [1:0] w_n20416_0;
	wire [1:0] w_n20422_0;
	wire [1:0] w_n20424_0;
	wire [2:0] w_n20425_0;
	wire [1:0] w_n20428_0;
	wire [1:0] w_n20430_0;
	wire [2:0] w_n20431_0;
	wire [1:0] w_n20433_0;
	wire [1:0] w_n20437_0;
	wire [1:0] w_n20440_0;
	wire [1:0] w_n20441_0;
	wire [2:0] w_n20442_0;
	wire [1:0] w_n20443_0;
	wire [1:0] w_n20447_0;
	wire [1:0] w_n20453_0;
	wire [1:0] w_n20454_0;
	wire [1:0] w_n20456_0;
	wire [1:0] w_n20458_0;
	wire [1:0] w_n20461_0;
	wire [1:0] w_n20467_0;
	wire [1:0] w_n20469_0;
	wire [2:0] w_n20470_0;
	wire [1:0] w_n20473_0;
	wire [1:0] w_n20475_0;
	wire [2:0] w_n20476_0;
	wire [1:0] w_n20478_0;
	wire [1:0] w_n20482_0;
	wire [1:0] w_n20485_0;
	wire [1:0] w_n20486_0;
	wire [2:0] w_n20487_0;
	wire [1:0] w_n20488_0;
	wire [1:0] w_n20492_0;
	wire [1:0] w_n20498_0;
	wire [1:0] w_n20499_0;
	wire [1:0] w_n20501_0;
	wire [1:0] w_n20503_0;
	wire [1:0] w_n20506_0;
	wire [1:0] w_n20512_0;
	wire [1:0] w_n20514_0;
	wire [2:0] w_n20515_0;
	wire [1:0] w_n20518_0;
	wire [1:0] w_n20520_0;
	wire [2:0] w_n20521_0;
	wire [1:0] w_n20523_0;
	wire [1:0] w_n20527_0;
	wire [1:0] w_n20530_0;
	wire [1:0] w_n20531_0;
	wire [2:0] w_n20532_0;
	wire [1:0] w_n20533_0;
	wire [1:0] w_n20537_0;
	wire [1:0] w_n20543_0;
	wire [1:0] w_n20544_0;
	wire [1:0] w_n20546_0;
	wire [1:0] w_n20548_0;
	wire [1:0] w_n20551_0;
	wire [1:0] w_n20557_0;
	wire [1:0] w_n20559_0;
	wire [2:0] w_n20560_0;
	wire [1:0] w_n20563_0;
	wire [1:0] w_n20565_0;
	wire [2:0] w_n20566_0;
	wire [1:0] w_n20568_0;
	wire [1:0] w_n20572_0;
	wire [1:0] w_n20575_0;
	wire [1:0] w_n20576_0;
	wire [2:0] w_n20577_0;
	wire [1:0] w_n20578_0;
	wire [1:0] w_n20582_0;
	wire [1:0] w_n20588_0;
	wire [1:0] w_n20589_0;
	wire [1:0] w_n20591_0;
	wire [1:0] w_n20593_0;
	wire [1:0] w_n20596_0;
	wire [1:0] w_n20602_0;
	wire [1:0] w_n20604_0;
	wire [2:0] w_n20605_0;
	wire [1:0] w_n20608_0;
	wire [1:0] w_n20610_0;
	wire [2:0] w_n20611_0;
	wire [1:0] w_n20613_0;
	wire [1:0] w_n20617_0;
	wire [1:0] w_n20620_0;
	wire [1:0] w_n20621_0;
	wire [2:0] w_n20622_0;
	wire [1:0] w_n20623_0;
	wire [1:0] w_n20627_0;
	wire [1:0] w_n20633_0;
	wire [1:0] w_n20634_0;
	wire [1:0] w_n20636_0;
	wire [1:0] w_n20638_0;
	wire [1:0] w_n20641_0;
	wire [1:0] w_n20647_0;
	wire [1:0] w_n20649_0;
	wire [2:0] w_n20650_0;
	wire [1:0] w_n20653_0;
	wire [1:0] w_n20655_0;
	wire [2:0] w_n20656_0;
	wire [1:0] w_n20658_0;
	wire [1:0] w_n20662_0;
	wire [1:0] w_n20665_0;
	wire [1:0] w_n20666_0;
	wire [2:0] w_n20667_0;
	wire [1:0] w_n20668_0;
	wire [1:0] w_n20672_0;
	wire [1:0] w_n20678_0;
	wire [1:0] w_n20679_0;
	wire [1:0] w_n20681_0;
	wire [1:0] w_n20683_0;
	wire [1:0] w_n20686_0;
	wire [1:0] w_n20692_0;
	wire [1:0] w_n20694_0;
	wire [2:0] w_n20695_0;
	wire [1:0] w_n20698_0;
	wire [1:0] w_n20700_0;
	wire [2:0] w_n20701_0;
	wire [1:0] w_n20703_0;
	wire [1:0] w_n20707_0;
	wire [1:0] w_n20710_0;
	wire [1:0] w_n20711_0;
	wire [2:0] w_n20712_0;
	wire [1:0] w_n20713_0;
	wire [1:0] w_n20717_0;
	wire [1:0] w_n20723_0;
	wire [1:0] w_n20724_0;
	wire [1:0] w_n20726_0;
	wire [1:0] w_n20728_0;
	wire [1:0] w_n20731_0;
	wire [1:0] w_n20737_0;
	wire [1:0] w_n20739_0;
	wire [2:0] w_n20740_0;
	wire [1:0] w_n20743_0;
	wire [1:0] w_n20745_0;
	wire [2:0] w_n20746_0;
	wire [1:0] w_n20748_0;
	wire [1:0] w_n20752_0;
	wire [1:0] w_n20755_0;
	wire [1:0] w_n20756_0;
	wire [2:0] w_n20757_0;
	wire [1:0] w_n20758_0;
	wire [1:0] w_n20762_0;
	wire [1:0] w_n20768_0;
	wire [1:0] w_n20769_0;
	wire [1:0] w_n20771_0;
	wire [1:0] w_n20773_0;
	wire [1:0] w_n20776_0;
	wire [1:0] w_n20782_0;
	wire [1:0] w_n20784_0;
	wire [2:0] w_n20785_0;
	wire [1:0] w_n20788_0;
	wire [1:0] w_n20790_0;
	wire [2:0] w_n20791_0;
	wire [1:0] w_n20793_0;
	wire [1:0] w_n20797_0;
	wire [1:0] w_n20800_0;
	wire [1:0] w_n20801_0;
	wire [2:0] w_n20802_0;
	wire [1:0] w_n20803_0;
	wire [1:0] w_n20807_0;
	wire [1:0] w_n20813_0;
	wire [1:0] w_n20814_0;
	wire [1:0] w_n20816_0;
	wire [1:0] w_n20818_0;
	wire [1:0] w_n20821_0;
	wire [1:0] w_n20827_0;
	wire [1:0] w_n20829_0;
	wire [2:0] w_n20830_0;
	wire [1:0] w_n20833_0;
	wire [1:0] w_n20835_0;
	wire [2:0] w_n20836_0;
	wire [1:0] w_n20838_0;
	wire [1:0] w_n20842_0;
	wire [1:0] w_n20845_0;
	wire [1:0] w_n20846_0;
	wire [2:0] w_n20847_0;
	wire [1:0] w_n20848_0;
	wire [1:0] w_n20852_0;
	wire [1:0] w_n20858_0;
	wire [1:0] w_n20859_0;
	wire [1:0] w_n20861_0;
	wire [1:0] w_n20865_0;
	wire [1:0] w_n20868_0;
	wire [1:0] w_n20869_0;
	wire [2:0] w_n20870_0;
	wire [1:0] w_n20871_0;
	wire [1:0] w_n20873_0;
	wire [1:0] w_n20875_0;
	wire [1:0] w_n20877_0;
	wire [1:0] w_n20880_0;
	wire [1:0] w_n20886_0;
	wire [2:0] w_n20888_0;
	wire [2:0] w_n20888_1;
	wire [2:0] w_n20891_0;
	wire [2:0] w_n20892_0;
	wire [1:0] w_n20893_0;
	wire [1:0] w_n20894_0;
	wire [1:0] w_n20901_0;
	wire [1:0] w_n20902_0;
	wire [2:0] w_n20910_0;
	wire [2:0] w_n20910_1;
	wire [2:0] w_n20910_2;
	wire [2:0] w_n20910_3;
	wire [2:0] w_n20910_4;
	wire [2:0] w_n20910_5;
	wire [2:0] w_n20910_6;
	wire [2:0] w_n20910_7;
	wire [2:0] w_n20910_8;
	wire [2:0] w_n20910_9;
	wire [2:0] w_n20910_10;
	wire [2:0] w_n20910_11;
	wire [2:0] w_n20910_12;
	wire [2:0] w_n20910_13;
	wire [2:0] w_n20910_14;
	wire [2:0] w_n20910_15;
	wire [2:0] w_n20910_16;
	wire [2:0] w_n20910_17;
	wire [1:0] w_n20913_0;
	wire [1:0] w_n20918_0;
	wire [1:0] w_n20921_0;
	wire [1:0] w_n20924_0;
	wire [1:0] w_n20934_0;
	wire [1:0] w_n20942_0;
	wire [1:0] w_n20950_0;
	wire [1:0] w_n20955_0;
	wire [1:0] w_n20960_0;
	wire [1:0] w_n20967_0;
	wire [1:0] w_n20975_0;
	wire [1:0] w_n20982_0;
	wire [1:0] w_n20989_0;
	wire [1:0] w_n20994_0;
	wire [1:0] w_n21001_0;
	wire [1:0] w_n21009_0;
	wire [1:0] w_n21016_0;
	wire [1:0] w_n21021_0;
	wire [1:0] w_n21028_0;
	wire [1:0] w_n21033_0;
	wire [1:0] w_n21040_0;
	wire [1:0] w_n21048_0;
	wire [1:0] w_n21055_0;
	wire [1:0] w_n21060_0;
	wire [1:0] w_n21067_0;
	wire [1:0] w_n21072_0;
	wire [1:0] w_n21079_0;
	wire [1:0] w_n21087_0;
	wire [1:0] w_n21094_0;
	wire [1:0] w_n21099_0;
	wire [1:0] w_n21106_0;
	wire [1:0] w_n21111_0;
	wire [1:0] w_n21118_0;
	wire [1:0] w_n21126_0;
	wire [1:0] w_n21133_0;
	wire [1:0] w_n21138_0;
	wire [1:0] w_n21145_0;
	wire [1:0] w_n21150_0;
	wire [1:0] w_n21157_0;
	wire [1:0] w_n21165_0;
	wire [1:0] w_n21172_0;
	wire [1:0] w_n21177_0;
	wire [1:0] w_n21184_0;
	wire [1:0] w_n21189_0;
	wire [1:0] w_n21196_0;
	wire [1:0] w_n21204_0;
	wire [1:0] w_n21211_0;
	wire [1:0] w_n21216_0;
	wire [1:0] w_n21223_0;
	wire [1:0] w_n21228_0;
	wire [1:0] w_n21235_0;
	wire [1:0] w_n21243_0;
	wire [1:0] w_n21250_0;
	wire [1:0] w_n21255_0;
	wire [1:0] w_n21262_0;
	wire [1:0] w_n21267_0;
	wire [1:0] w_n21274_0;
	wire [1:0] w_n21282_0;
	wire [1:0] w_n21289_0;
	wire [1:0] w_n21294_0;
	wire [1:0] w_n21301_0;
	wire [1:0] w_n21306_0;
	wire [1:0] w_n21313_0;
	wire [1:0] w_n21321_0;
	wire [1:0] w_n21328_0;
	wire [1:0] w_n21333_0;
	wire [1:0] w_n21340_0;
	wire [1:0] w_n21345_0;
	wire [1:0] w_n21352_0;
	wire [1:0] w_n21360_0;
	wire [1:0] w_n21367_0;
	wire [1:0] w_n21372_0;
	wire [1:0] w_n21379_0;
	wire [1:0] w_n21384_0;
	wire [1:0] w_n21391_0;
	wire [1:0] w_n21399_0;
	wire [1:0] w_n21406_0;
	wire [1:0] w_n21411_0;
	wire [1:0] w_n21418_0;
	wire [1:0] w_n21423_0;
	wire [1:0] w_n21430_0;
	wire [1:0] w_n21438_0;
	wire [1:0] w_n21445_0;
	wire [1:0] w_n21450_0;
	wire [1:0] w_n21457_0;
	wire [1:0] w_n21462_0;
	wire [1:0] w_n21469_0;
	wire [1:0] w_n21476_0;
	wire [1:0] w_n21481_0;
	wire [1:0] w_n21490_0;
	wire [1:0] w_n21494_0;
	wire [1:0] w_n21496_0;
	jnot g00000(.din(w_a126_0[2]),.dout(n192),.clk(gclk));
	jnot g00001(.din(w_a127_0[1]),.dout(n193),.clk(gclk));
	jand g00002(.dina(w_n193_0[1]),.dinb(w_n192_0[1]),.dout(n194),.clk(gclk));
	jand g00003(.dina(w_a127_0[0]),.dinb(w_a126_0[1]),.dout(n195),.clk(gclk));
	jor g00004(.dina(w_a125_0[1]),.dinb(w_a124_0[2]),.dout(n196),.clk(gclk));
	jand g00005(.dina(w_n196_0[1]),.dinb(w_n192_0[0]),.dout(n197),.clk(gclk));
	jor g00006(.dina(w_n197_0[1]),.dinb(w_n195_0[1]),.dout(asqrt_fa_63),.clk(gclk));
	jnot g00007(.din(w_asqrt62_31),.dout(n199),.clk(gclk));
	jnot g00008(.din(w_a63_0[1]),.dout(n200),.clk(gclk));
	jnot g00009(.din(w_n194_43[2]),.dout(asqrt[63]),.clk(gclk));
	jnot g00010(.din(w_a125_0[0]),.dout(n202),.clk(gclk));
	jnot g00011(.din(w_a124_0[1]),.dout(n203),.clk(gclk));
	jand g00012(.dina(w_asqrt62_30[2]),.dinb(w_n203_0[2]),.dout(n204),.clk(gclk));
	jor g00013(.dina(n204),.dinb(n202),.dout(n205),.clk(gclk));
	jnot g00014(.din(w_n196_0[0]),.dout(n206),.clk(gclk));
	jand g00015(.dina(w_n206_0[1]),.dinb(w_n195_0[0]),.dout(n207),.clk(gclk));
	jnot g00016(.din(n207),.dout(n208),.clk(gclk));
	jand g00017(.dina(n208),.dinb(n205),.dout(n209),.clk(gclk));
	jand g00018(.dina(w_asqrt62_30[1]),.dinb(w_a124_0[0]),.dout(n210),.clk(gclk));
	jnot g00019(.din(w_a122_0[1]),.dout(n211),.clk(gclk));
	jnot g00020(.din(w_a123_0[1]),.dout(n212),.clk(gclk));
	jand g00021(.dina(w_n203_0[1]),.dinb(w_n212_0[1]),.dout(n213),.clk(gclk));
	jand g00022(.dina(n213),.dinb(w_n211_1[1]),.dout(n214),.clk(gclk));
	jor g00023(.dina(n214),.dinb(n210),.dout(n215),.clk(gclk));
	jand g00024(.dina(w_n215_0[2]),.dinb(w_n209_0[2]),.dout(n216),.clk(gclk));
	jor g00025(.dina(w_n216_0[2]),.dinb(w_asqrt63_17),.dout(n217),.clk(gclk));
	jor g00026(.dina(w_n215_0[1]),.dinb(w_n209_0[1]),.dout(n218),.clk(gclk));
	jand g00027(.dina(w_n206_0[0]),.dinb(w_a126_0[0]),.dout(n219),.clk(gclk));
	jor g00028(.dina(w_n197_0[0]),.dinb(w_n193_0[0]),.dout(n220),.clk(gclk));
	jor g00029(.dina(n220),.dinb(n219),.dout(n221),.clk(gclk));
	jand g00030(.dina(w_n221_0[1]),.dinb(w_n218_0[1]),.dout(n222),.clk(gclk));
	jand g00031(.dina(n222),.dinb(n217),.dout(n223),.clk(gclk));
	jnot g00032(.din(w_n223_39[2]),.dout(asqrt_fa_62),.clk(gclk));
	jor g00033(.dina(w_asqrt61_31),.dinb(w_n199_45[2]),.dout(n225),.clk(gclk));
	jor g00034(.dina(w_n223_39[1]),.dinb(w_a122_0[0]),.dout(n226),.clk(gclk));
	jor g00035(.dina(w_n226_0[1]),.dinb(w_a123_0[0]),.dout(n227),.clk(gclk));
	jand g00036(.dina(n227),.dinb(n225),.dout(n228),.clk(gclk));
	jxor g00037(.dina(n228),.dinb(w_n203_0[0]),.dout(n229),.clk(gclk));
	jor g00038(.dina(w_n223_39[0]),.dinb(w_n211_1[0]),.dout(n230),.clk(gclk));
	jnot g00039(.din(w_a120_0[1]),.dout(n231),.clk(gclk));
	jnot g00040(.din(a[121]),.dout(n232),.clk(gclk));
	jand g00041(.dina(w_n211_0[2]),.dinb(w_n232_0[2]),.dout(n233),.clk(gclk));
	jand g00042(.dina(n233),.dinb(w_n231_1[1]),.dout(n234),.clk(gclk));
	jnot g00043(.din(n234),.dout(n235),.clk(gclk));
	jand g00044(.dina(n235),.dinb(n230),.dout(n236),.clk(gclk));
	jor g00045(.dina(w_n236_0[2]),.dinb(w_n199_45[1]),.dout(n237),.clk(gclk));
	jand g00046(.dina(w_n236_0[1]),.dinb(w_n199_45[0]),.dout(n238),.clk(gclk));
	jxor g00047(.dina(w_n226_0[0]),.dinb(w_n212_0[0]),.dout(n239),.clk(gclk));
	jor g00048(.dina(w_n239_0[1]),.dinb(n238),.dout(n240),.clk(gclk));
	jand g00049(.dina(n240),.dinb(n237),.dout(n241),.clk(gclk));
	jor g00050(.dina(w_n241_0[1]),.dinb(w_n229_0[2]),.dout(n242),.clk(gclk));
	jnot g00051(.din(w_n218_0[0]),.dout(n243),.clk(gclk));
	jnot g00052(.din(w_n221_0[0]),.dout(n244),.clk(gclk));
	jand g00053(.dina(n244),.dinb(w_n216_0[1]),.dout(n245),.clk(gclk));
	jor g00054(.dina(n245),.dinb(n243),.dout(n246),.clk(gclk));
	jor g00055(.dina(n246),.dinb(w_n242_0[2]),.dout(n247),.clk(gclk));
	jand g00056(.dina(n247),.dinb(w_n194_43[1]),.dout(n248),.clk(gclk));
	jand g00057(.dina(w_n241_0[0]),.dinb(w_n229_0[1]),.dout(n249),.clk(gclk));
	jand g00058(.dina(w_asqrt61_30[2]),.dinb(w_n209_0[0]),.dout(n250),.clk(gclk));
	jor g00059(.dina(n250),.dinb(w_n215_0[0]),.dout(n251),.clk(gclk));
	jnot g00060(.din(w_n216_0[0]),.dout(n252),.clk(gclk));
	jand g00061(.dina(n252),.dinb(w_asqrt63_16[2]),.dout(n253),.clk(gclk));
	jand g00062(.dina(n253),.dinb(n251),.dout(n254),.clk(gclk));
	jor g00063(.dina(w_n254_0[1]),.dinb(w_n249_0[1]),.dout(n258),.clk(gclk));
	jor g00064(.dina(n258),.dinb(w_n248_0[1]),.dout(asqrt_fa_61),.clk(gclk));
	jand g00065(.dina(w_asqrt60_30[1]),.dinb(w_a120_0[0]),.dout(n260),.clk(gclk));
	jnot g00066(.din(w_a118_0[1]),.dout(n261),.clk(gclk));
	jnot g00067(.din(w_a119_0[1]),.dout(n262),.clk(gclk));
	jand g00068(.dina(w_n231_1[0]),.dinb(w_n262_0[1]),.dout(n263),.clk(gclk));
	jand g00069(.dina(n263),.dinb(w_n261_1[1]),.dout(n264),.clk(gclk));
	jor g00070(.dina(n264),.dinb(n260),.dout(n265),.clk(gclk));
	jand g00071(.dina(w_n265_0[2]),.dinb(w_asqrt61_30[1]),.dout(n266),.clk(gclk));
	jand g00072(.dina(w_asqrt60_30[0]),.dinb(w_n231_0[2]),.dout(n267),.clk(gclk));
	jxor g00073(.dina(w_n267_0[1]),.dinb(w_n232_0[1]),.dout(n268),.clk(gclk));
	jor g00074(.dina(w_n265_0[1]),.dinb(w_asqrt61_30[0]),.dout(n269),.clk(gclk));
	jand g00075(.dina(n269),.dinb(w_n268_0[1]),.dout(n270),.clk(gclk));
	jor g00076(.dina(w_n270_0[1]),.dinb(w_n266_0[1]),.dout(n271),.clk(gclk));
	jand g00077(.dina(n271),.dinb(w_asqrt62_30[0]),.dout(n272),.clk(gclk));
	jor g00078(.dina(w_n266_0[0]),.dinb(w_asqrt62_29[2]),.dout(n273),.clk(gclk));
	jor g00079(.dina(n273),.dinb(w_n270_0[0]),.dout(n274),.clk(gclk));
	jand g00080(.dina(w_n267_0[0]),.dinb(w_n232_0[0]),.dout(n275),.clk(gclk));
	jnot g00081(.din(w_n248_0[0]),.dout(n276),.clk(gclk));
	jnot g00082(.din(w_n249_0[0]),.dout(n277),.clk(gclk));
	jnot g00083(.din(w_n254_0[0]),.dout(n278),.clk(gclk));
	jand g00084(.dina(n278),.dinb(w_asqrt61_29[2]),.dout(n279),.clk(gclk));
	jand g00085(.dina(n279),.dinb(w_n277_0[2]),.dout(n280),.clk(gclk));
	jand g00086(.dina(n280),.dinb(n276),.dout(n281),.clk(gclk));
	jor g00087(.dina(n281),.dinb(n275),.dout(n282),.clk(gclk));
	jxor g00088(.dina(n282),.dinb(w_n211_0[1]),.dout(n283),.clk(gclk));
	jand g00089(.dina(w_n283_0[1]),.dinb(w_n274_0[1]),.dout(n284),.clk(gclk));
	jor g00090(.dina(n284),.dinb(w_n272_0[1]),.dout(n285),.clk(gclk));
	jnot g00091(.din(w_n239_0[0]),.dout(n286),.clk(gclk));
	jxor g00092(.dina(w_n236_0[0]),.dinb(w_n199_44[2]),.dout(n287),.clk(gclk));
	jand g00093(.dina(n287),.dinb(w_asqrt60_29[2]),.dout(n288),.clk(gclk));
	jxor g00094(.dina(n288),.dinb(n286),.dout(n289),.clk(gclk));
	jnot g00095(.din(w_asqrt60_29[1]),.dout(n290),.clk(gclk));
	jor g00096(.dina(w_n290_39[1]),.dinb(w_n242_0[1]),.dout(n291),.clk(gclk));
	jand g00097(.dina(n291),.dinb(w_n277_0[1]),.dout(n292),.clk(gclk));
	jand g00098(.dina(n292),.dinb(w_n289_1[1]),.dout(n293),.clk(gclk));
	jand g00099(.dina(n293),.dinb(w_n285_1[1]),.dout(n294),.clk(gclk));
	jor g00100(.dina(n294),.dinb(w_asqrt63_16[1]),.dout(n295),.clk(gclk));
	jor g00101(.dina(w_n289_1[0]),.dinb(w_n285_1[0]),.dout(n296),.clk(gclk));
	jnot g00102(.din(w_n229_0[0]),.dout(n297),.clk(gclk));
	jand g00103(.dina(w_n290_39[0]),.dinb(n297),.dout(n298),.clk(gclk));
	jand g00104(.dina(w_n277_0[0]),.dinb(w_asqrt63_16[0]),.dout(n299),.clk(gclk));
	jand g00105(.dina(n299),.dinb(w_n242_0[0]),.dout(n300),.clk(gclk));
	jor g00106(.dina(n300),.dinb(w_n290_38[2]),.dout(n301),.clk(gclk));
	jnot g00107(.din(w_n301_0[1]),.dout(n302),.clk(gclk));
	jor g00108(.dina(n302),.dinb(n298),.dout(n303),.clk(gclk));
	jand g00109(.dina(n303),.dinb(w_n296_0[2]),.dout(n304),.clk(gclk));
	jand g00110(.dina(n304),.dinb(w_n295_0[1]),.dout(n305),.clk(gclk));
	jnot g00111(.din(w_n305_39[2]),.dout(asqrt_fa_60),.clk(gclk));
	jor g00112(.dina(w_n305_39[1]),.dinb(w_n261_1[0]),.dout(n307),.clk(gclk));
	jnot g00113(.din(w_a116_0[1]),.dout(n308),.clk(gclk));
	jnot g00114(.din(a[117]),.dout(n309),.clk(gclk));
	jand g00115(.dina(w_n261_0[2]),.dinb(w_n309_0[2]),.dout(n310),.clk(gclk));
	jand g00116(.dina(n310),.dinb(w_n308_1[1]),.dout(n311),.clk(gclk));
	jnot g00117(.din(n311),.dout(n312),.clk(gclk));
	jand g00118(.dina(n312),.dinb(n307),.dout(n313),.clk(gclk));
	jor g00119(.dina(w_n313_0[2]),.dinb(w_n290_38[1]),.dout(n314),.clk(gclk));
	jor g00120(.dina(w_n305_39[0]),.dinb(w_a118_0[0]),.dout(n315),.clk(gclk));
	jxor g00121(.dina(w_n315_0[1]),.dinb(w_n262_0[0]),.dout(n316),.clk(gclk));
	jand g00122(.dina(w_n313_0[1]),.dinb(w_n290_38[0]),.dout(n317),.clk(gclk));
	jor g00123(.dina(n317),.dinb(w_n316_0[1]),.dout(n318),.clk(gclk));
	jand g00124(.dina(w_n318_0[1]),.dinb(w_n314_0[1]),.dout(n319),.clk(gclk));
	jor g00125(.dina(n319),.dinb(w_n223_38[2]),.dout(n320),.clk(gclk));
	jand g00126(.dina(w_n314_0[0]),.dinb(w_n223_38[1]),.dout(n321),.clk(gclk));
	jand g00127(.dina(n321),.dinb(w_n318_0[0]),.dout(n322),.clk(gclk));
	jor g00128(.dina(w_n315_0[0]),.dinb(w_a119_0[0]),.dout(n323),.clk(gclk));
	jnot g00129(.din(w_n295_0[0]),.dout(n324),.clk(gclk));
	jnot g00130(.din(w_n296_0[1]),.dout(n325),.clk(gclk));
	jor g00131(.dina(w_n301_0[0]),.dinb(w_n325_0[1]),.dout(n326),.clk(gclk));
	jor g00132(.dina(n326),.dinb(n324),.dout(n327),.clk(gclk));
	jand g00133(.dina(n327),.dinb(n323),.dout(n328),.clk(gclk));
	jxor g00134(.dina(n328),.dinb(w_n231_0[1]),.dout(n329),.clk(gclk));
	jor g00135(.dina(w_n329_0[1]),.dinb(w_n322_0[1]),.dout(n330),.clk(gclk));
	jand g00136(.dina(n330),.dinb(w_n320_0[1]),.dout(n331),.clk(gclk));
	jor g00137(.dina(w_n331_0[2]),.dinb(w_n199_44[1]),.dout(n332),.clk(gclk));
	jand g00138(.dina(w_n331_0[1]),.dinb(w_n199_44[0]),.dout(n333),.clk(gclk));
	jxor g00139(.dina(w_n265_0[0]),.dinb(w_n223_38[0]),.dout(n334),.clk(gclk));
	jor g00140(.dina(n334),.dinb(w_n305_38[2]),.dout(n335),.clk(gclk));
	jxor g00141(.dina(n335),.dinb(w_n268_0[0]),.dout(n336),.clk(gclk));
	jor g00142(.dina(w_n336_0[1]),.dinb(n333),.dout(n337),.clk(gclk));
	jand g00143(.dina(n337),.dinb(n332),.dout(n338),.clk(gclk));
	jnot g00144(.din(w_n274_0[0]),.dout(n339),.clk(gclk));
	jor g00145(.dina(n339),.dinb(w_n272_0[0]),.dout(n340),.clk(gclk));
	jor g00146(.dina(n340),.dinb(w_n305_38[1]),.dout(n341),.clk(gclk));
	jxor g00147(.dina(n341),.dinb(w_n283_0[0]),.dout(n342),.clk(gclk));
	jand g00148(.dina(w_n289_0[2]),.dinb(w_n285_0[2]),.dout(n343),.clk(gclk));
	jand g00149(.dina(n343),.dinb(w_asqrt59_30[1]),.dout(n344),.clk(gclk));
	jor g00150(.dina(n344),.dinb(w_n325_0[0]),.dout(n345),.clk(gclk));
	jor g00151(.dina(n345),.dinb(w_n342_0[2]),.dout(n346),.clk(gclk));
	jor g00152(.dina(n346),.dinb(w_n338_0[2]),.dout(n347),.clk(gclk));
	jand g00153(.dina(n347),.dinb(w_n194_43[0]),.dout(n348),.clk(gclk));
	jand g00154(.dina(w_n342_0[1]),.dinb(w_n338_0[1]),.dout(n349),.clk(gclk));
	jnot g00155(.din(w_n289_0[1]),.dout(n350),.clk(gclk));
	jnot g00156(.din(w_n285_0[1]),.dout(n351),.clk(gclk));
	jand g00157(.dina(w_asqrt59_30[0]),.dinb(n351),.dout(n352),.clk(gclk));
	jor g00158(.dina(n352),.dinb(n350),.dout(n353),.clk(gclk));
	jnot g00159(.din(n353),.dout(n354),.clk(gclk));
	jand g00160(.dina(w_n296_0[0]),.dinb(w_asqrt63_15[2]),.dout(n355),.clk(gclk));
	jnot g00161(.din(n355),.dout(n356),.clk(gclk));
	jand g00162(.dina(n356),.dinb(w_asqrt59_29[2]),.dout(n357),.clk(gclk));
	jor g00163(.dina(n357),.dinb(n354),.dout(n358),.clk(gclk));
	jnot g00164(.din(w_n358_0[1]),.dout(n359),.clk(gclk));
	jor g00165(.dina(n359),.dinb(w_n349_0[2]),.dout(n360),.clk(gclk));
	jor g00166(.dina(n360),.dinb(w_n348_0[1]),.dout(asqrt_fa_59),.clk(gclk));
	jand g00167(.dina(w_asqrt58_31),.dinb(w_a116_0[0]),.dout(n362),.clk(gclk));
	jnot g00168(.din(w_a114_0[1]),.dout(n363),.clk(gclk));
	jnot g00169(.din(w_a115_0[1]),.dout(n364),.clk(gclk));
	jand g00170(.dina(w_n308_1[0]),.dinb(w_n364_0[1]),.dout(n365),.clk(gclk));
	jand g00171(.dina(n365),.dinb(w_n363_1[1]),.dout(n366),.clk(gclk));
	jor g00172(.dina(n366),.dinb(n362),.dout(n367),.clk(gclk));
	jand g00173(.dina(w_n367_0[2]),.dinb(w_asqrt59_29[1]),.dout(n368),.clk(gclk));
	jand g00174(.dina(w_asqrt58_30[2]),.dinb(w_n308_0[2]),.dout(n369),.clk(gclk));
	jxor g00175(.dina(w_n369_0[1]),.dinb(w_n309_0[1]),.dout(n370),.clk(gclk));
	jor g00176(.dina(w_n367_0[1]),.dinb(w_asqrt59_29[0]),.dout(n371),.clk(gclk));
	jand g00177(.dina(n371),.dinb(w_n370_0[1]),.dout(n372),.clk(gclk));
	jor g00178(.dina(w_n372_0[1]),.dinb(w_n368_0[1]),.dout(n373),.clk(gclk));
	jand g00179(.dina(n373),.dinb(w_asqrt60_29[0]),.dout(n374),.clk(gclk));
	jor g00180(.dina(w_n368_0[0]),.dinb(w_asqrt60_28[2]),.dout(n375),.clk(gclk));
	jor g00181(.dina(n375),.dinb(w_n372_0[0]),.dout(n376),.clk(gclk));
	jand g00182(.dina(w_n369_0[0]),.dinb(w_n309_0[0]),.dout(n377),.clk(gclk));
	jnot g00183(.din(w_n348_0[0]),.dout(n378),.clk(gclk));
	jnot g00184(.din(w_n349_0[1]),.dout(n379),.clk(gclk));
	jand g00185(.dina(w_n358_0[0]),.dinb(w_asqrt59_28[2]),.dout(n381),.clk(gclk));
	jand g00186(.dina(n381),.dinb(n379),.dout(n382),.clk(gclk));
	jand g00187(.dina(n382),.dinb(n378),.dout(n383),.clk(gclk));
	jor g00188(.dina(n383),.dinb(n377),.dout(n384),.clk(gclk));
	jxor g00189(.dina(n384),.dinb(w_n261_0[1]),.dout(n385),.clk(gclk));
	jand g00190(.dina(w_n385_0[1]),.dinb(w_n376_0[1]),.dout(n386),.clk(gclk));
	jor g00191(.dina(n386),.dinb(w_n374_0[1]),.dout(n387),.clk(gclk));
	jand g00192(.dina(w_n387_0[2]),.dinb(w_asqrt61_29[1]),.dout(n388),.clk(gclk));
	jor g00193(.dina(w_n387_0[1]),.dinb(w_asqrt61_29[0]),.dout(n389),.clk(gclk));
	jxor g00194(.dina(w_n313_0[0]),.dinb(w_n290_37[2]),.dout(n390),.clk(gclk));
	jand g00195(.dina(n390),.dinb(w_asqrt58_30[1]),.dout(n391),.clk(gclk));
	jxor g00196(.dina(n391),.dinb(w_n316_0[0]),.dout(n392),.clk(gclk));
	jnot g00197(.din(w_n392_0[1]),.dout(n393),.clk(gclk));
	jand g00198(.dina(n393),.dinb(n389),.dout(n394),.clk(gclk));
	jor g00199(.dina(w_n394_0[1]),.dinb(w_n388_0[1]),.dout(n395),.clk(gclk));
	jand g00200(.dina(n395),.dinb(w_asqrt62_29[1]),.dout(n396),.clk(gclk));
	jnot g00201(.din(w_n322_0[0]),.dout(n397),.clk(gclk));
	jand g00202(.dina(n397),.dinb(w_n320_0[0]),.dout(n398),.clk(gclk));
	jand g00203(.dina(n398),.dinb(w_asqrt58_30[0]),.dout(n399),.clk(gclk));
	jxor g00204(.dina(n399),.dinb(w_n329_0[0]),.dout(n400),.clk(gclk));
	jnot g00205(.din(n400),.dout(n401),.clk(gclk));
	jor g00206(.dina(w_n388_0[0]),.dinb(w_asqrt62_29[0]),.dout(n402),.clk(gclk));
	jor g00207(.dina(n402),.dinb(w_n394_0[0]),.dout(n403),.clk(gclk));
	jand g00208(.dina(w_n403_0[1]),.dinb(w_n401_0[1]),.dout(n404),.clk(gclk));
	jor g00209(.dina(w_n404_0[1]),.dinb(w_n396_0[1]),.dout(n405),.clk(gclk));
	jxor g00210(.dina(w_n331_0[0]),.dinb(w_n199_43[2]),.dout(n406),.clk(gclk));
	jand g00211(.dina(n406),.dinb(w_asqrt58_29[2]),.dout(n407),.clk(gclk));
	jxor g00212(.dina(n407),.dinb(w_n336_0[0]),.dout(n408),.clk(gclk));
	jnot g00213(.din(w_n338_0[0]),.dout(n409),.clk(gclk));
	jnot g00214(.din(w_n342_0[0]),.dout(n410),.clk(gclk));
	jand g00215(.dina(w_asqrt58_29[1]),.dinb(w_n410_0[1]),.dout(n411),.clk(gclk));
	jand g00216(.dina(w_n411_0[1]),.dinb(w_n409_0[2]),.dout(n412),.clk(gclk));
	jor g00217(.dina(n412),.dinb(w_n349_0[0]),.dout(n413),.clk(gclk));
	jor g00218(.dina(n413),.dinb(w_n408_0[1]),.dout(n414),.clk(gclk));
	jnot g00219(.din(n414),.dout(n415),.clk(gclk));
	jand g00220(.dina(n415),.dinb(w_n405_1[2]),.dout(n416),.clk(gclk));
	jor g00221(.dina(n416),.dinb(w_asqrt63_15[1]),.dout(n417),.clk(gclk));
	jnot g00222(.din(w_n408_0[0]),.dout(n418),.clk(gclk));
	jor g00223(.dina(w_n418_0[2]),.dinb(w_n405_1[1]),.dout(n419),.clk(gclk));
	jor g00224(.dina(w_n411_0[0]),.dinb(w_n409_0[1]),.dout(n420),.clk(gclk));
	jand g00225(.dina(w_n410_0[0]),.dinb(w_n409_0[0]),.dout(n421),.clk(gclk));
	jor g00226(.dina(n421),.dinb(w_n194_42[2]),.dout(n422),.clk(gclk));
	jnot g00227(.din(n422),.dout(n423),.clk(gclk));
	jand g00228(.dina(n423),.dinb(n420),.dout(n424),.clk(gclk));
	jnot g00229(.din(w_asqrt58_29[0]),.dout(n425),.clk(gclk));
	jnot g00230(.din(w_n424_0[1]),.dout(n428),.clk(gclk));
	jand g00231(.dina(n428),.dinb(w_n419_0[1]),.dout(n429),.clk(gclk));
	jand g00232(.dina(n429),.dinb(w_n417_0[1]),.dout(n430),.clk(gclk));
	jnot g00233(.din(w_n430_38[2]),.dout(asqrt_fa_58),.clk(gclk));
	jor g00234(.dina(w_n430_38[1]),.dinb(w_n363_1[0]),.dout(n432),.clk(gclk));
	jnot g00235(.din(w_a112_0[1]),.dout(n433),.clk(gclk));
	jnot g00236(.din(a[113]),.dout(n434),.clk(gclk));
	jand g00237(.dina(w_n363_0[2]),.dinb(w_n434_0[2]),.dout(n435),.clk(gclk));
	jand g00238(.dina(n435),.dinb(w_n433_1[1]),.dout(n436),.clk(gclk));
	jnot g00239(.din(n436),.dout(n437),.clk(gclk));
	jand g00240(.dina(n437),.dinb(n432),.dout(n438),.clk(gclk));
	jor g00241(.dina(w_n438_0[2]),.dinb(w_n425_36[2]),.dout(n439),.clk(gclk));
	jor g00242(.dina(w_n430_38[0]),.dinb(w_a114_0[0]),.dout(n440),.clk(gclk));
	jxor g00243(.dina(w_n440_0[1]),.dinb(w_n364_0[0]),.dout(n441),.clk(gclk));
	jand g00244(.dina(w_n438_0[1]),.dinb(w_n425_36[1]),.dout(n442),.clk(gclk));
	jor g00245(.dina(n442),.dinb(w_n441_0[1]),.dout(n443),.clk(gclk));
	jand g00246(.dina(w_n443_0[1]),.dinb(w_n439_0[1]),.dout(n444),.clk(gclk));
	jor g00247(.dina(n444),.dinb(w_n305_38[0]),.dout(n445),.clk(gclk));
	jand g00248(.dina(w_n439_0[0]),.dinb(w_n305_37[2]),.dout(n446),.clk(gclk));
	jand g00249(.dina(n446),.dinb(w_n443_0[0]),.dout(n447),.clk(gclk));
	jor g00250(.dina(w_n440_0[0]),.dinb(w_a115_0[0]),.dout(n448),.clk(gclk));
	jnot g00251(.din(w_n417_0[0]),.dout(n449),.clk(gclk));
	jnot g00252(.din(w_n419_0[0]),.dout(n450),.clk(gclk));
	jor g00253(.dina(w_n424_0[0]),.dinb(w_n425_36[0]),.dout(n451),.clk(gclk));
	jor g00254(.dina(n451),.dinb(w_n450_0[1]),.dout(n452),.clk(gclk));
	jor g00255(.dina(n452),.dinb(n449),.dout(n453),.clk(gclk));
	jand g00256(.dina(n453),.dinb(n448),.dout(n454),.clk(gclk));
	jxor g00257(.dina(n454),.dinb(w_n308_0[1]),.dout(n455),.clk(gclk));
	jor g00258(.dina(w_n455_0[1]),.dinb(w_n447_0[1]),.dout(n456),.clk(gclk));
	jand g00259(.dina(n456),.dinb(w_n445_0[1]),.dout(n457),.clk(gclk));
	jor g00260(.dina(w_n457_0[2]),.dinb(w_n290_37[1]),.dout(n458),.clk(gclk));
	jand g00261(.dina(w_n457_0[1]),.dinb(w_n290_37[0]),.dout(n459),.clk(gclk));
	jxor g00262(.dina(w_n367_0[0]),.dinb(w_n305_37[1]),.dout(n460),.clk(gclk));
	jor g00263(.dina(n460),.dinb(w_n430_37[2]),.dout(n461),.clk(gclk));
	jxor g00264(.dina(n461),.dinb(w_n370_0[0]),.dout(n462),.clk(gclk));
	jor g00265(.dina(w_n462_0[1]),.dinb(n459),.dout(n463),.clk(gclk));
	jand g00266(.dina(w_n463_0[1]),.dinb(w_n458_0[1]),.dout(n464),.clk(gclk));
	jor g00267(.dina(n464),.dinb(w_n223_37[2]),.dout(n465),.clk(gclk));
	jnot g00268(.din(w_n376_0[0]),.dout(n466),.clk(gclk));
	jor g00269(.dina(n466),.dinb(w_n374_0[0]),.dout(n467),.clk(gclk));
	jor g00270(.dina(n467),.dinb(w_n430_37[1]),.dout(n468),.clk(gclk));
	jxor g00271(.dina(n468),.dinb(w_n385_0[0]),.dout(n469),.clk(gclk));
	jand g00272(.dina(w_n458_0[0]),.dinb(w_n223_37[1]),.dout(n470),.clk(gclk));
	jand g00273(.dina(n470),.dinb(w_n463_0[0]),.dout(n471),.clk(gclk));
	jor g00274(.dina(w_n471_0[1]),.dinb(w_n469_0[1]),.dout(n472),.clk(gclk));
	jand g00275(.dina(w_n472_0[1]),.dinb(w_n465_0[1]),.dout(n473),.clk(gclk));
	jor g00276(.dina(w_n473_0[2]),.dinb(w_n199_43[1]),.dout(n474),.clk(gclk));
	jand g00277(.dina(w_n473_0[1]),.dinb(w_n199_43[0]),.dout(n475),.clk(gclk));
	jxor g00278(.dina(w_n387_0[0]),.dinb(w_n223_37[0]),.dout(n476),.clk(gclk));
	jor g00279(.dina(n476),.dinb(w_n430_37[0]),.dout(n477),.clk(gclk));
	jxor g00280(.dina(n477),.dinb(w_n392_0[0]),.dout(n478),.clk(gclk));
	jnot g00281(.din(w_n478_0[1]),.dout(n479),.clk(gclk));
	jor g00282(.dina(n479),.dinb(n475),.dout(n480),.clk(gclk));
	jand g00283(.dina(n480),.dinb(n474),.dout(n481),.clk(gclk));
	jnot g00284(.din(w_n396_0[0]),.dout(n482),.clk(gclk));
	jand g00285(.dina(w_asqrt57_29),.dinb(n482),.dout(n483),.clk(gclk));
	jand g00286(.dina(w_n483_0[1]),.dinb(w_n403_0[0]),.dout(n484),.clk(gclk));
	jor g00287(.dina(n484),.dinb(w_n401_0[0]),.dout(n485),.clk(gclk));
	jand g00288(.dina(w_n483_0[0]),.dinb(w_n404_0[0]),.dout(n486),.clk(gclk));
	jnot g00289(.din(n486),.dout(n487),.clk(gclk));
	jand g00290(.dina(n487),.dinb(n485),.dout(n488),.clk(gclk));
	jnot g00291(.din(w_n488_0[2]),.dout(n489),.clk(gclk));
	jand g00292(.dina(w_asqrt57_28[2]),.dinb(w_n418_0[1]),.dout(n490),.clk(gclk));
	jand g00293(.dina(w_n490_0[1]),.dinb(w_n405_1[0]),.dout(n491),.clk(gclk));
	jor g00294(.dina(n491),.dinb(w_n450_0[0]),.dout(n492),.clk(gclk));
	jor g00295(.dina(n492),.dinb(w_n489_0[1]),.dout(n493),.clk(gclk));
	jor g00296(.dina(n493),.dinb(w_n481_0[2]),.dout(n494),.clk(gclk));
	jand g00297(.dina(n494),.dinb(w_n194_42[1]),.dout(n495),.clk(gclk));
	jand g00298(.dina(w_n489_0[0]),.dinb(w_n481_0[1]),.dout(n496),.clk(gclk));
	jor g00299(.dina(w_n490_0[0]),.dinb(w_n405_0[2]),.dout(n497),.clk(gclk));
	jand g00300(.dina(w_n418_0[0]),.dinb(w_n405_0[1]),.dout(n498),.clk(gclk));
	jor g00301(.dina(n498),.dinb(w_n194_42[0]),.dout(n499),.clk(gclk));
	jnot g00302(.din(n499),.dout(n500),.clk(gclk));
	jand g00303(.dina(n500),.dinb(n497),.dout(n501),.clk(gclk));
	jor g00304(.dina(w_n501_0[1]),.dinb(w_n496_0[2]),.dout(n504),.clk(gclk));
	jor g00305(.dina(n504),.dinb(w_n495_0[1]),.dout(asqrt_fa_57),.clk(gclk));
	jand g00306(.dina(w_asqrt56_31),.dinb(w_a112_0[0]),.dout(n506),.clk(gclk));
	jnot g00307(.din(w_a110_0[1]),.dout(n507),.clk(gclk));
	jnot g00308(.din(w_a111_0[1]),.dout(n508),.clk(gclk));
	jand g00309(.dina(w_n433_1[0]),.dinb(w_n508_0[1]),.dout(n509),.clk(gclk));
	jand g00310(.dina(n509),.dinb(w_n507_1[1]),.dout(n510),.clk(gclk));
	jor g00311(.dina(n510),.dinb(n506),.dout(n511),.clk(gclk));
	jand g00312(.dina(w_n511_0[2]),.dinb(w_asqrt57_28[1]),.dout(n512),.clk(gclk));
	jand g00313(.dina(w_asqrt56_30[2]),.dinb(w_n433_0[2]),.dout(n513),.clk(gclk));
	jxor g00314(.dina(w_n513_0[1]),.dinb(w_n434_0[1]),.dout(n514),.clk(gclk));
	jor g00315(.dina(w_n511_0[1]),.dinb(w_asqrt57_28[0]),.dout(n515),.clk(gclk));
	jand g00316(.dina(n515),.dinb(w_n514_0[1]),.dout(n516),.clk(gclk));
	jor g00317(.dina(w_n516_0[1]),.dinb(w_n512_0[1]),.dout(n517),.clk(gclk));
	jand g00318(.dina(n517),.dinb(w_asqrt58_28[2]),.dout(n518),.clk(gclk));
	jor g00319(.dina(w_n512_0[0]),.dinb(w_asqrt58_28[1]),.dout(n519),.clk(gclk));
	jor g00320(.dina(n519),.dinb(w_n516_0[0]),.dout(n520),.clk(gclk));
	jand g00321(.dina(w_n513_0[0]),.dinb(w_n434_0[0]),.dout(n521),.clk(gclk));
	jnot g00322(.din(w_n495_0[0]),.dout(n522),.clk(gclk));
	jnot g00323(.din(w_n496_0[1]),.dout(n523),.clk(gclk));
	jnot g00324(.din(w_n501_0[0]),.dout(n524),.clk(gclk));
	jand g00325(.dina(n524),.dinb(w_asqrt57_27[2]),.dout(n525),.clk(gclk));
	jand g00326(.dina(n525),.dinb(n523),.dout(n526),.clk(gclk));
	jand g00327(.dina(n526),.dinb(n522),.dout(n527),.clk(gclk));
	jor g00328(.dina(n527),.dinb(n521),.dout(n528),.clk(gclk));
	jxor g00329(.dina(n528),.dinb(w_n363_0[1]),.dout(n529),.clk(gclk));
	jand g00330(.dina(w_n529_0[1]),.dinb(w_n520_0[1]),.dout(n530),.clk(gclk));
	jor g00331(.dina(n530),.dinb(w_n518_0[1]),.dout(n531),.clk(gclk));
	jand g00332(.dina(w_n531_0[2]),.dinb(w_asqrt59_28[1]),.dout(n532),.clk(gclk));
	jor g00333(.dina(w_n531_0[1]),.dinb(w_asqrt59_28[0]),.dout(n533),.clk(gclk));
	jxor g00334(.dina(w_n438_0[0]),.dinb(w_n425_35[2]),.dout(n534),.clk(gclk));
	jand g00335(.dina(n534),.dinb(w_asqrt56_30[1]),.dout(n535),.clk(gclk));
	jxor g00336(.dina(n535),.dinb(w_n441_0[0]),.dout(n536),.clk(gclk));
	jnot g00337(.din(w_n536_0[1]),.dout(n537),.clk(gclk));
	jand g00338(.dina(n537),.dinb(n533),.dout(n538),.clk(gclk));
	jor g00339(.dina(w_n538_0[1]),.dinb(w_n532_0[1]),.dout(n539),.clk(gclk));
	jand g00340(.dina(n539),.dinb(w_asqrt60_28[1]),.dout(n540),.clk(gclk));
	jnot g00341(.din(w_n447_0[0]),.dout(n541),.clk(gclk));
	jand g00342(.dina(n541),.dinb(w_n445_0[0]),.dout(n542),.clk(gclk));
	jand g00343(.dina(n542),.dinb(w_asqrt56_30[0]),.dout(n543),.clk(gclk));
	jxor g00344(.dina(n543),.dinb(w_n455_0[0]),.dout(n544),.clk(gclk));
	jnot g00345(.din(n544),.dout(n545),.clk(gclk));
	jor g00346(.dina(w_n532_0[0]),.dinb(w_asqrt60_28[0]),.dout(n546),.clk(gclk));
	jor g00347(.dina(n546),.dinb(w_n538_0[0]),.dout(n547),.clk(gclk));
	jand g00348(.dina(w_n547_0[1]),.dinb(w_n545_0[1]),.dout(n548),.clk(gclk));
	jor g00349(.dina(w_n548_0[1]),.dinb(w_n540_0[1]),.dout(n549),.clk(gclk));
	jand g00350(.dina(w_n549_0[2]),.dinb(w_asqrt61_28[2]),.dout(n550),.clk(gclk));
	jor g00351(.dina(w_n549_0[1]),.dinb(w_asqrt61_28[1]),.dout(n551),.clk(gclk));
	jnot g00352(.din(w_n462_0[0]),.dout(n552),.clk(gclk));
	jxor g00353(.dina(w_n457_0[0]),.dinb(w_n290_36[2]),.dout(n553),.clk(gclk));
	jand g00354(.dina(n553),.dinb(w_asqrt56_29[2]),.dout(n554),.clk(gclk));
	jxor g00355(.dina(n554),.dinb(n552),.dout(n555),.clk(gclk));
	jand g00356(.dina(w_n555_0[1]),.dinb(n551),.dout(n556),.clk(gclk));
	jor g00357(.dina(w_n556_0[1]),.dinb(w_n550_0[1]),.dout(n557),.clk(gclk));
	jand g00358(.dina(n557),.dinb(w_asqrt62_28[2]),.dout(n558),.clk(gclk));
	jor g00359(.dina(w_n550_0[0]),.dinb(w_asqrt62_28[1]),.dout(n559),.clk(gclk));
	jor g00360(.dina(n559),.dinb(w_n556_0[0]),.dout(n560),.clk(gclk));
	jnot g00361(.din(w_n469_0[0]),.dout(n561),.clk(gclk));
	jnot g00362(.din(w_n471_0[0]),.dout(n562),.clk(gclk));
	jand g00363(.dina(w_asqrt56_29[1]),.dinb(w_n465_0[0]),.dout(n563),.clk(gclk));
	jand g00364(.dina(w_n563_0[1]),.dinb(n562),.dout(n564),.clk(gclk));
	jor g00365(.dina(n564),.dinb(n561),.dout(n565),.clk(gclk));
	jnot g00366(.din(w_n472_0[0]),.dout(n566),.clk(gclk));
	jand g00367(.dina(w_n563_0[0]),.dinb(n566),.dout(n567),.clk(gclk));
	jnot g00368(.din(n567),.dout(n568),.clk(gclk));
	jand g00369(.dina(n568),.dinb(n565),.dout(n569),.clk(gclk));
	jand g00370(.dina(w_n569_0[1]),.dinb(w_n560_0[1]),.dout(n570),.clk(gclk));
	jor g00371(.dina(n570),.dinb(w_n558_0[1]),.dout(n571),.clk(gclk));
	jxor g00372(.dina(w_n473_0[0]),.dinb(w_n199_42[2]),.dout(n572),.clk(gclk));
	jand g00373(.dina(n572),.dinb(w_asqrt56_29[0]),.dout(n573),.clk(gclk));
	jxor g00374(.dina(n573),.dinb(w_n478_0[0]),.dout(n574),.clk(gclk));
	jnot g00375(.din(w_n574_1[1]),.dout(n575),.clk(gclk));
	jnot g00376(.din(w_n481_0[0]),.dout(n576),.clk(gclk));
	jand g00377(.dina(w_asqrt56_28[2]),.dinb(w_n488_0[1]),.dout(n577),.clk(gclk));
	jand g00378(.dina(w_n577_0[1]),.dinb(w_n576_0[2]),.dout(n578),.clk(gclk));
	jor g00379(.dina(n578),.dinb(w_n496_0[0]),.dout(n579),.clk(gclk));
	jor g00380(.dina(n579),.dinb(n575),.dout(n580),.clk(gclk));
	jnot g00381(.din(n580),.dout(n581),.clk(gclk));
	jand g00382(.dina(n581),.dinb(w_n571_1[2]),.dout(n582),.clk(gclk));
	jor g00383(.dina(n582),.dinb(w_asqrt63_15[0]),.dout(n583),.clk(gclk));
	jor g00384(.dina(w_n574_1[0]),.dinb(w_n571_1[1]),.dout(n584),.clk(gclk));
	jor g00385(.dina(w_n577_0[0]),.dinb(w_n576_0[1]),.dout(n585),.clk(gclk));
	jand g00386(.dina(w_n488_0[0]),.dinb(w_n576_0[0]),.dout(n586),.clk(gclk));
	jor g00387(.dina(n586),.dinb(w_n194_41[2]),.dout(n587),.clk(gclk));
	jnot g00388(.din(n587),.dout(n588),.clk(gclk));
	jand g00389(.dina(n588),.dinb(n585),.dout(n589),.clk(gclk));
	jnot g00390(.din(w_asqrt56_28[1]),.dout(n590),.clk(gclk));
	jnot g00391(.din(w_n589_0[1]),.dout(n593),.clk(gclk));
	jand g00392(.dina(n593),.dinb(w_n584_0[1]),.dout(n594),.clk(gclk));
	jand g00393(.dina(n594),.dinb(w_n583_0[1]),.dout(n595),.clk(gclk));
	jnot g00394(.din(w_n595_38[2]),.dout(asqrt_fa_56),.clk(gclk));
	jor g00395(.dina(w_n595_38[1]),.dinb(w_n507_1[0]),.dout(n597),.clk(gclk));
	jnot g00396(.din(w_a108_0[1]),.dout(n598),.clk(gclk));
	jnot g00397(.din(a[109]),.dout(n599),.clk(gclk));
	jand g00398(.dina(w_n507_0[2]),.dinb(w_n599_0[2]),.dout(n600),.clk(gclk));
	jand g00399(.dina(n600),.dinb(w_n598_1[1]),.dout(n601),.clk(gclk));
	jnot g00400(.din(n601),.dout(n602),.clk(gclk));
	jand g00401(.dina(n602),.dinb(n597),.dout(n603),.clk(gclk));
	jor g00402(.dina(w_n603_0[2]),.dinb(w_n590_35[2]),.dout(n604),.clk(gclk));
	jor g00403(.dina(w_n595_38[0]),.dinb(w_a110_0[0]),.dout(n605),.clk(gclk));
	jxor g00404(.dina(w_n605_0[1]),.dinb(w_n508_0[0]),.dout(n606),.clk(gclk));
	jand g00405(.dina(w_n603_0[1]),.dinb(w_n590_35[1]),.dout(n607),.clk(gclk));
	jor g00406(.dina(n607),.dinb(w_n606_0[1]),.dout(n608),.clk(gclk));
	jand g00407(.dina(w_n608_0[1]),.dinb(w_n604_0[1]),.dout(n609),.clk(gclk));
	jor g00408(.dina(n609),.dinb(w_n430_36[2]),.dout(n610),.clk(gclk));
	jand g00409(.dina(w_n604_0[0]),.dinb(w_n430_36[1]),.dout(n611),.clk(gclk));
	jand g00410(.dina(n611),.dinb(w_n608_0[0]),.dout(n612),.clk(gclk));
	jor g00411(.dina(w_n605_0[0]),.dinb(w_a111_0[0]),.dout(n613),.clk(gclk));
	jnot g00412(.din(w_n583_0[0]),.dout(n614),.clk(gclk));
	jnot g00413(.din(w_n584_0[0]),.dout(n615),.clk(gclk));
	jor g00414(.dina(w_n589_0[0]),.dinb(w_n590_35[0]),.dout(n616),.clk(gclk));
	jor g00415(.dina(n616),.dinb(w_n615_0[1]),.dout(n617),.clk(gclk));
	jor g00416(.dina(n617),.dinb(n614),.dout(n618),.clk(gclk));
	jand g00417(.dina(n618),.dinb(n613),.dout(n619),.clk(gclk));
	jxor g00418(.dina(n619),.dinb(w_n433_0[1]),.dout(n620),.clk(gclk));
	jor g00419(.dina(w_n620_0[1]),.dinb(w_n612_0[1]),.dout(n621),.clk(gclk));
	jand g00420(.dina(n621),.dinb(w_n610_0[1]),.dout(n622),.clk(gclk));
	jor g00421(.dina(w_n622_0[2]),.dinb(w_n425_35[1]),.dout(n623),.clk(gclk));
	jand g00422(.dina(w_n622_0[1]),.dinb(w_n425_35[0]),.dout(n624),.clk(gclk));
	jxor g00423(.dina(w_n511_0[0]),.dinb(w_n430_36[0]),.dout(n625),.clk(gclk));
	jor g00424(.dina(n625),.dinb(w_n595_37[2]),.dout(n626),.clk(gclk));
	jxor g00425(.dina(n626),.dinb(w_n514_0[0]),.dout(n627),.clk(gclk));
	jor g00426(.dina(w_n627_0[1]),.dinb(n624),.dout(n628),.clk(gclk));
	jand g00427(.dina(w_n628_0[1]),.dinb(w_n623_0[1]),.dout(n629),.clk(gclk));
	jor g00428(.dina(n629),.dinb(w_n305_37[0]),.dout(n630),.clk(gclk));
	jnot g00429(.din(w_n520_0[0]),.dout(n631),.clk(gclk));
	jor g00430(.dina(n631),.dinb(w_n518_0[0]),.dout(n632),.clk(gclk));
	jor g00431(.dina(n632),.dinb(w_n595_37[1]),.dout(n633),.clk(gclk));
	jxor g00432(.dina(n633),.dinb(w_n529_0[0]),.dout(n634),.clk(gclk));
	jand g00433(.dina(w_n623_0[0]),.dinb(w_n305_36[2]),.dout(n635),.clk(gclk));
	jand g00434(.dina(n635),.dinb(w_n628_0[0]),.dout(n636),.clk(gclk));
	jor g00435(.dina(w_n636_0[1]),.dinb(w_n634_0[1]),.dout(n637),.clk(gclk));
	jand g00436(.dina(w_n637_0[1]),.dinb(w_n630_0[1]),.dout(n638),.clk(gclk));
	jor g00437(.dina(w_n638_0[2]),.dinb(w_n290_36[1]),.dout(n639),.clk(gclk));
	jand g00438(.dina(w_n638_0[1]),.dinb(w_n290_36[0]),.dout(n640),.clk(gclk));
	jxor g00439(.dina(w_n531_0[0]),.dinb(w_n305_36[1]),.dout(n641),.clk(gclk));
	jor g00440(.dina(n641),.dinb(w_n595_37[0]),.dout(n642),.clk(gclk));
	jxor g00441(.dina(n642),.dinb(w_n536_0[0]),.dout(n643),.clk(gclk));
	jnot g00442(.din(w_n643_0[1]),.dout(n644),.clk(gclk));
	jor g00443(.dina(n644),.dinb(n640),.dout(n645),.clk(gclk));
	jand g00444(.dina(w_n645_0[1]),.dinb(w_n639_0[1]),.dout(n646),.clk(gclk));
	jor g00445(.dina(n646),.dinb(w_n223_36[2]),.dout(n647),.clk(gclk));
	jand g00446(.dina(w_n639_0[0]),.dinb(w_n223_36[1]),.dout(n648),.clk(gclk));
	jand g00447(.dina(n648),.dinb(w_n645_0[0]),.dout(n649),.clk(gclk));
	jnot g00448(.din(w_n540_0[0]),.dout(n650),.clk(gclk));
	jand g00449(.dina(w_asqrt55_28),.dinb(n650),.dout(n651),.clk(gclk));
	jand g00450(.dina(w_n651_0[1]),.dinb(w_n547_0[0]),.dout(n652),.clk(gclk));
	jor g00451(.dina(n652),.dinb(w_n545_0[0]),.dout(n653),.clk(gclk));
	jand g00452(.dina(w_n651_0[0]),.dinb(w_n548_0[0]),.dout(n654),.clk(gclk));
	jnot g00453(.din(n654),.dout(n655),.clk(gclk));
	jand g00454(.dina(n655),.dinb(n653),.dout(n656),.clk(gclk));
	jnot g00455(.din(n656),.dout(n657),.clk(gclk));
	jor g00456(.dina(w_n657_0[1]),.dinb(w_n649_0[1]),.dout(n658),.clk(gclk));
	jand g00457(.dina(n658),.dinb(w_n647_0[1]),.dout(n659),.clk(gclk));
	jor g00458(.dina(w_n659_0[2]),.dinb(w_n199_42[1]),.dout(n660),.clk(gclk));
	jand g00459(.dina(w_n659_0[1]),.dinb(w_n199_42[0]),.dout(n661),.clk(gclk));
	jnot g00460(.din(w_n555_0[0]),.dout(n662),.clk(gclk));
	jxor g00461(.dina(w_n549_0[0]),.dinb(w_n223_36[0]),.dout(n663),.clk(gclk));
	jor g00462(.dina(n663),.dinb(w_n595_36[2]),.dout(n664),.clk(gclk));
	jxor g00463(.dina(n664),.dinb(n662),.dout(n665),.clk(gclk));
	jnot g00464(.din(w_n665_0[1]),.dout(n666),.clk(gclk));
	jor g00465(.dina(n666),.dinb(n661),.dout(n667),.clk(gclk));
	jand g00466(.dina(n667),.dinb(n660),.dout(n668),.clk(gclk));
	jnot g00467(.din(w_n560_0[0]),.dout(n669),.clk(gclk));
	jor g00468(.dina(n669),.dinb(w_n558_0[0]),.dout(n670),.clk(gclk));
	jor g00469(.dina(n670),.dinb(w_n595_36[1]),.dout(n671),.clk(gclk));
	jxor g00470(.dina(n671),.dinb(w_n569_0[0]),.dout(n672),.clk(gclk));
	jand g00471(.dina(w_asqrt55_27[2]),.dinb(w_n574_0[2]),.dout(n673),.clk(gclk));
	jand g00472(.dina(w_n673_0[1]),.dinb(w_n571_1[0]),.dout(n674),.clk(gclk));
	jor g00473(.dina(n674),.dinb(w_n615_0[0]),.dout(n675),.clk(gclk));
	jor g00474(.dina(n675),.dinb(w_n672_0[2]),.dout(n676),.clk(gclk));
	jor g00475(.dina(n676),.dinb(w_n668_0[2]),.dout(n677),.clk(gclk));
	jand g00476(.dina(n677),.dinb(w_n194_41[1]),.dout(n678),.clk(gclk));
	jand g00477(.dina(w_n672_0[1]),.dinb(w_n668_0[1]),.dout(n679),.clk(gclk));
	jor g00478(.dina(w_n673_0[0]),.dinb(w_n571_0[2]),.dout(n680),.clk(gclk));
	jand g00479(.dina(w_n574_0[1]),.dinb(w_n571_0[1]),.dout(n681),.clk(gclk));
	jor g00480(.dina(n681),.dinb(w_n194_41[0]),.dout(n682),.clk(gclk));
	jnot g00481(.din(n682),.dout(n683),.clk(gclk));
	jand g00482(.dina(n683),.dinb(n680),.dout(n684),.clk(gclk));
	jor g00483(.dina(w_n684_0[1]),.dinb(w_n679_0[2]),.dout(n687),.clk(gclk));
	jor g00484(.dina(n687),.dinb(w_n678_0[1]),.dout(asqrt_fa_55),.clk(gclk));
	jand g00485(.dina(w_asqrt54_31),.dinb(w_a108_0[0]),.dout(n689),.clk(gclk));
	jnot g00486(.din(w_a106_0[1]),.dout(n690),.clk(gclk));
	jnot g00487(.din(w_a107_0[1]),.dout(n691),.clk(gclk));
	jand g00488(.dina(w_n598_1[0]),.dinb(w_n691_0[1]),.dout(n692),.clk(gclk));
	jand g00489(.dina(n692),.dinb(w_n690_1[1]),.dout(n693),.clk(gclk));
	jor g00490(.dina(n693),.dinb(n689),.dout(n694),.clk(gclk));
	jand g00491(.dina(w_n694_0[2]),.dinb(w_asqrt55_27[1]),.dout(n695),.clk(gclk));
	jand g00492(.dina(w_asqrt54_30[2]),.dinb(w_n598_0[2]),.dout(n696),.clk(gclk));
	jxor g00493(.dina(w_n696_0[1]),.dinb(w_n599_0[1]),.dout(n697),.clk(gclk));
	jor g00494(.dina(w_n694_0[1]),.dinb(w_asqrt55_27[0]),.dout(n698),.clk(gclk));
	jand g00495(.dina(n698),.dinb(w_n697_0[1]),.dout(n699),.clk(gclk));
	jor g00496(.dina(w_n699_0[1]),.dinb(w_n695_0[1]),.dout(n700),.clk(gclk));
	jand g00497(.dina(n700),.dinb(w_asqrt56_28[0]),.dout(n701),.clk(gclk));
	jor g00498(.dina(w_n695_0[0]),.dinb(w_asqrt56_27[2]),.dout(n702),.clk(gclk));
	jor g00499(.dina(n702),.dinb(w_n699_0[0]),.dout(n703),.clk(gclk));
	jand g00500(.dina(w_n696_0[0]),.dinb(w_n599_0[0]),.dout(n704),.clk(gclk));
	jnot g00501(.din(w_n678_0[0]),.dout(n705),.clk(gclk));
	jnot g00502(.din(w_n679_0[1]),.dout(n706),.clk(gclk));
	jnot g00503(.din(w_n684_0[0]),.dout(n707),.clk(gclk));
	jand g00504(.dina(n707),.dinb(w_asqrt55_26[2]),.dout(n708),.clk(gclk));
	jand g00505(.dina(n708),.dinb(n706),.dout(n709),.clk(gclk));
	jand g00506(.dina(n709),.dinb(n705),.dout(n710),.clk(gclk));
	jor g00507(.dina(n710),.dinb(n704),.dout(n711),.clk(gclk));
	jxor g00508(.dina(n711),.dinb(w_n507_0[1]),.dout(n712),.clk(gclk));
	jand g00509(.dina(w_n712_0[1]),.dinb(w_n703_0[1]),.dout(n713),.clk(gclk));
	jor g00510(.dina(n713),.dinb(w_n701_0[1]),.dout(n714),.clk(gclk));
	jand g00511(.dina(w_n714_0[2]),.dinb(w_asqrt57_27[1]),.dout(n715),.clk(gclk));
	jor g00512(.dina(w_n714_0[1]),.dinb(w_asqrt57_27[0]),.dout(n716),.clk(gclk));
	jxor g00513(.dina(w_n603_0[0]),.dinb(w_n590_34[2]),.dout(n717),.clk(gclk));
	jand g00514(.dina(n717),.dinb(w_asqrt54_30[1]),.dout(n718),.clk(gclk));
	jxor g00515(.dina(n718),.dinb(w_n606_0[0]),.dout(n719),.clk(gclk));
	jnot g00516(.din(w_n719_0[1]),.dout(n720),.clk(gclk));
	jand g00517(.dina(n720),.dinb(n716),.dout(n721),.clk(gclk));
	jor g00518(.dina(w_n721_0[1]),.dinb(w_n715_0[1]),.dout(n722),.clk(gclk));
	jand g00519(.dina(n722),.dinb(w_asqrt58_28[0]),.dout(n723),.clk(gclk));
	jnot g00520(.din(w_n612_0[0]),.dout(n724),.clk(gclk));
	jand g00521(.dina(n724),.dinb(w_n610_0[0]),.dout(n725),.clk(gclk));
	jand g00522(.dina(n725),.dinb(w_asqrt54_30[0]),.dout(n726),.clk(gclk));
	jxor g00523(.dina(n726),.dinb(w_n620_0[0]),.dout(n727),.clk(gclk));
	jnot g00524(.din(n727),.dout(n728),.clk(gclk));
	jor g00525(.dina(w_n715_0[0]),.dinb(w_asqrt58_27[2]),.dout(n729),.clk(gclk));
	jor g00526(.dina(n729),.dinb(w_n721_0[0]),.dout(n730),.clk(gclk));
	jand g00527(.dina(w_n730_0[1]),.dinb(w_n728_0[1]),.dout(n731),.clk(gclk));
	jor g00528(.dina(w_n731_0[1]),.dinb(w_n723_0[1]),.dout(n732),.clk(gclk));
	jand g00529(.dina(w_n732_0[2]),.dinb(w_asqrt59_27[2]),.dout(n733),.clk(gclk));
	jor g00530(.dina(w_n732_0[1]),.dinb(w_asqrt59_27[1]),.dout(n734),.clk(gclk));
	jnot g00531(.din(w_n627_0[0]),.dout(n735),.clk(gclk));
	jxor g00532(.dina(w_n622_0[0]),.dinb(w_n425_34[2]),.dout(n736),.clk(gclk));
	jand g00533(.dina(n736),.dinb(w_asqrt54_29[2]),.dout(n737),.clk(gclk));
	jxor g00534(.dina(n737),.dinb(n735),.dout(n738),.clk(gclk));
	jand g00535(.dina(w_n738_0[1]),.dinb(n734),.dout(n739),.clk(gclk));
	jor g00536(.dina(w_n739_0[1]),.dinb(w_n733_0[1]),.dout(n740),.clk(gclk));
	jand g00537(.dina(n740),.dinb(w_asqrt60_27[2]),.dout(n741),.clk(gclk));
	jor g00538(.dina(w_n733_0[0]),.dinb(w_asqrt60_27[1]),.dout(n742),.clk(gclk));
	jor g00539(.dina(n742),.dinb(w_n739_0[0]),.dout(n743),.clk(gclk));
	jnot g00540(.din(w_n634_0[0]),.dout(n744),.clk(gclk));
	jnot g00541(.din(w_n636_0[0]),.dout(n745),.clk(gclk));
	jand g00542(.dina(w_asqrt54_29[1]),.dinb(w_n630_0[0]),.dout(n746),.clk(gclk));
	jand g00543(.dina(w_n746_0[1]),.dinb(n745),.dout(n747),.clk(gclk));
	jor g00544(.dina(n747),.dinb(n744),.dout(n748),.clk(gclk));
	jnot g00545(.din(w_n637_0[0]),.dout(n749),.clk(gclk));
	jand g00546(.dina(w_n746_0[0]),.dinb(n749),.dout(n750),.clk(gclk));
	jnot g00547(.din(n750),.dout(n751),.clk(gclk));
	jand g00548(.dina(n751),.dinb(n748),.dout(n752),.clk(gclk));
	jand g00549(.dina(w_n752_0[1]),.dinb(w_n743_0[1]),.dout(n753),.clk(gclk));
	jor g00550(.dina(n753),.dinb(w_n741_0[1]),.dout(n754),.clk(gclk));
	jand g00551(.dina(w_n754_0[2]),.dinb(w_asqrt61_28[0]),.dout(n755),.clk(gclk));
	jor g00552(.dina(w_n754_0[1]),.dinb(w_asqrt61_27[2]),.dout(n756),.clk(gclk));
	jxor g00553(.dina(w_n638_0[0]),.dinb(w_n290_35[2]),.dout(n757),.clk(gclk));
	jand g00554(.dina(n757),.dinb(w_asqrt54_29[0]),.dout(n758),.clk(gclk));
	jxor g00555(.dina(n758),.dinb(w_n643_0[0]),.dout(n759),.clk(gclk));
	jand g00556(.dina(w_n759_0[1]),.dinb(n756),.dout(n760),.clk(gclk));
	jor g00557(.dina(w_n760_0[1]),.dinb(w_n755_0[1]),.dout(n761),.clk(gclk));
	jand g00558(.dina(n761),.dinb(w_asqrt62_28[0]),.dout(n762),.clk(gclk));
	jnot g00559(.din(w_n649_0[0]),.dout(n763),.clk(gclk));
	jand g00560(.dina(n763),.dinb(w_n647_0[0]),.dout(n764),.clk(gclk));
	jand g00561(.dina(n764),.dinb(w_asqrt54_28[2]),.dout(n765),.clk(gclk));
	jxor g00562(.dina(n765),.dinb(w_n657_0[0]),.dout(n766),.clk(gclk));
	jnot g00563(.din(n766),.dout(n767),.clk(gclk));
	jor g00564(.dina(w_n755_0[0]),.dinb(w_asqrt62_27[2]),.dout(n768),.clk(gclk));
	jor g00565(.dina(n768),.dinb(w_n760_0[0]),.dout(n769),.clk(gclk));
	jand g00566(.dina(w_n769_0[1]),.dinb(w_n767_0[1]),.dout(n770),.clk(gclk));
	jor g00567(.dina(w_n770_0[1]),.dinb(w_n762_0[1]),.dout(n771),.clk(gclk));
	jxor g00568(.dina(w_n659_0[0]),.dinb(w_n199_41[2]),.dout(n772),.clk(gclk));
	jand g00569(.dina(n772),.dinb(w_asqrt54_28[1]),.dout(n773),.clk(gclk));
	jxor g00570(.dina(n773),.dinb(w_n665_0[0]),.dout(n774),.clk(gclk));
	jnot g00571(.din(w_n774_1[1]),.dout(n775),.clk(gclk));
	jnot g00572(.din(w_n668_0[0]),.dout(n776),.clk(gclk));
	jnot g00573(.din(w_n672_0[0]),.dout(n777),.clk(gclk));
	jand g00574(.dina(w_asqrt54_28[0]),.dinb(w_n777_0[1]),.dout(n778),.clk(gclk));
	jand g00575(.dina(w_n778_0[1]),.dinb(w_n776_0[2]),.dout(n779),.clk(gclk));
	jor g00576(.dina(n779),.dinb(w_n679_0[0]),.dout(n780),.clk(gclk));
	jor g00577(.dina(n780),.dinb(n775),.dout(n781),.clk(gclk));
	jnot g00578(.din(n781),.dout(n782),.clk(gclk));
	jand g00579(.dina(n782),.dinb(w_n771_1[2]),.dout(n783),.clk(gclk));
	jor g00580(.dina(n783),.dinb(w_asqrt63_14[2]),.dout(n784),.clk(gclk));
	jor g00581(.dina(w_n774_1[0]),.dinb(w_n771_1[1]),.dout(n785),.clk(gclk));
	jor g00582(.dina(w_n778_0[0]),.dinb(w_n776_0[1]),.dout(n786),.clk(gclk));
	jand g00583(.dina(w_n777_0[0]),.dinb(w_n776_0[0]),.dout(n787),.clk(gclk));
	jor g00584(.dina(n787),.dinb(w_n194_40[2]),.dout(n788),.clk(gclk));
	jnot g00585(.din(n788),.dout(n789),.clk(gclk));
	jand g00586(.dina(n789),.dinb(n786),.dout(n790),.clk(gclk));
	jnot g00587(.din(w_asqrt54_27[2]),.dout(n791),.clk(gclk));
	jnot g00588(.din(w_n790_0[1]),.dout(n794),.clk(gclk));
	jand g00589(.dina(n794),.dinb(w_n785_0[1]),.dout(n795),.clk(gclk));
	jand g00590(.dina(n795),.dinb(w_n784_0[1]),.dout(n796),.clk(gclk));
	jnot g00591(.din(w_n796_37[2]),.dout(asqrt_fa_54),.clk(gclk));
	jor g00592(.dina(w_n796_37[1]),.dinb(w_n690_1[0]),.dout(n798),.clk(gclk));
	jnot g00593(.din(w_a104_0[1]),.dout(n799),.clk(gclk));
	jnot g00594(.din(a[105]),.dout(n800),.clk(gclk));
	jand g00595(.dina(w_n690_0[2]),.dinb(w_n800_0[2]),.dout(n801),.clk(gclk));
	jand g00596(.dina(n801),.dinb(w_n799_1[1]),.dout(n802),.clk(gclk));
	jnot g00597(.din(n802),.dout(n803),.clk(gclk));
	jand g00598(.dina(n803),.dinb(n798),.dout(n804),.clk(gclk));
	jor g00599(.dina(w_n804_0[2]),.dinb(w_n791_34[1]),.dout(n805),.clk(gclk));
	jor g00600(.dina(w_n796_37[0]),.dinb(w_a106_0[0]),.dout(n806),.clk(gclk));
	jxor g00601(.dina(w_n806_0[1]),.dinb(w_n691_0[0]),.dout(n807),.clk(gclk));
	jand g00602(.dina(w_n804_0[1]),.dinb(w_n791_34[0]),.dout(n808),.clk(gclk));
	jor g00603(.dina(n808),.dinb(w_n807_0[1]),.dout(n809),.clk(gclk));
	jand g00604(.dina(w_n809_0[1]),.dinb(w_n805_0[1]),.dout(n810),.clk(gclk));
	jor g00605(.dina(n810),.dinb(w_n595_36[0]),.dout(n811),.clk(gclk));
	jand g00606(.dina(w_n805_0[0]),.dinb(w_n595_35[2]),.dout(n812),.clk(gclk));
	jand g00607(.dina(n812),.dinb(w_n809_0[0]),.dout(n813),.clk(gclk));
	jor g00608(.dina(w_n806_0[0]),.dinb(w_a107_0[0]),.dout(n814),.clk(gclk));
	jnot g00609(.din(w_n784_0[0]),.dout(n815),.clk(gclk));
	jnot g00610(.din(w_n785_0[0]),.dout(n816),.clk(gclk));
	jor g00611(.dina(w_n790_0[0]),.dinb(w_n791_33[2]),.dout(n817),.clk(gclk));
	jor g00612(.dina(n817),.dinb(w_n816_0[1]),.dout(n818),.clk(gclk));
	jor g00613(.dina(n818),.dinb(n815),.dout(n819),.clk(gclk));
	jand g00614(.dina(n819),.dinb(n814),.dout(n820),.clk(gclk));
	jxor g00615(.dina(n820),.dinb(w_n598_0[1]),.dout(n821),.clk(gclk));
	jor g00616(.dina(w_n821_0[1]),.dinb(w_n813_0[1]),.dout(n822),.clk(gclk));
	jand g00617(.dina(n822),.dinb(w_n811_0[1]),.dout(n823),.clk(gclk));
	jor g00618(.dina(w_n823_0[2]),.dinb(w_n590_34[1]),.dout(n824),.clk(gclk));
	jand g00619(.dina(w_n823_0[1]),.dinb(w_n590_34[0]),.dout(n825),.clk(gclk));
	jxor g00620(.dina(w_n694_0[0]),.dinb(w_n595_35[1]),.dout(n826),.clk(gclk));
	jor g00621(.dina(n826),.dinb(w_n796_36[2]),.dout(n827),.clk(gclk));
	jxor g00622(.dina(n827),.dinb(w_n697_0[0]),.dout(n828),.clk(gclk));
	jor g00623(.dina(w_n828_0[1]),.dinb(n825),.dout(n829),.clk(gclk));
	jand g00624(.dina(w_n829_0[1]),.dinb(w_n824_0[1]),.dout(n830),.clk(gclk));
	jor g00625(.dina(n830),.dinb(w_n430_35[2]),.dout(n831),.clk(gclk));
	jnot g00626(.din(w_n703_0[0]),.dout(n832),.clk(gclk));
	jor g00627(.dina(n832),.dinb(w_n701_0[0]),.dout(n833),.clk(gclk));
	jor g00628(.dina(n833),.dinb(w_n796_36[1]),.dout(n834),.clk(gclk));
	jxor g00629(.dina(n834),.dinb(w_n712_0[0]),.dout(n835),.clk(gclk));
	jand g00630(.dina(w_n824_0[0]),.dinb(w_n430_35[1]),.dout(n836),.clk(gclk));
	jand g00631(.dina(n836),.dinb(w_n829_0[0]),.dout(n837),.clk(gclk));
	jor g00632(.dina(w_n837_0[1]),.dinb(w_n835_0[1]),.dout(n838),.clk(gclk));
	jand g00633(.dina(w_n838_0[1]),.dinb(w_n831_0[1]),.dout(n839),.clk(gclk));
	jor g00634(.dina(w_n839_0[2]),.dinb(w_n425_34[1]),.dout(n840),.clk(gclk));
	jand g00635(.dina(w_n839_0[1]),.dinb(w_n425_34[0]),.dout(n841),.clk(gclk));
	jxor g00636(.dina(w_n714_0[0]),.dinb(w_n430_35[0]),.dout(n842),.clk(gclk));
	jor g00637(.dina(n842),.dinb(w_n796_36[0]),.dout(n843),.clk(gclk));
	jxor g00638(.dina(n843),.dinb(w_n719_0[0]),.dout(n844),.clk(gclk));
	jnot g00639(.din(w_n844_0[1]),.dout(n845),.clk(gclk));
	jor g00640(.dina(n845),.dinb(n841),.dout(n846),.clk(gclk));
	jand g00641(.dina(w_n846_0[1]),.dinb(w_n840_0[1]),.dout(n847),.clk(gclk));
	jor g00642(.dina(n847),.dinb(w_n305_36[0]),.dout(n848),.clk(gclk));
	jand g00643(.dina(w_n840_0[0]),.dinb(w_n305_35[2]),.dout(n849),.clk(gclk));
	jand g00644(.dina(n849),.dinb(w_n846_0[0]),.dout(n850),.clk(gclk));
	jnot g00645(.din(w_n723_0[0]),.dout(n851),.clk(gclk));
	jand g00646(.dina(w_asqrt53_27[1]),.dinb(n851),.dout(n852),.clk(gclk));
	jand g00647(.dina(w_n852_0[1]),.dinb(w_n730_0[0]),.dout(n853),.clk(gclk));
	jor g00648(.dina(n853),.dinb(w_n728_0[0]),.dout(n854),.clk(gclk));
	jand g00649(.dina(w_n852_0[0]),.dinb(w_n731_0[0]),.dout(n855),.clk(gclk));
	jnot g00650(.din(n855),.dout(n856),.clk(gclk));
	jand g00651(.dina(n856),.dinb(n854),.dout(n857),.clk(gclk));
	jnot g00652(.din(n857),.dout(n858),.clk(gclk));
	jor g00653(.dina(w_n858_0[1]),.dinb(w_n850_0[1]),.dout(n859),.clk(gclk));
	jand g00654(.dina(n859),.dinb(w_n848_0[1]),.dout(n860),.clk(gclk));
	jor g00655(.dina(w_n860_0[2]),.dinb(w_n290_35[1]),.dout(n861),.clk(gclk));
	jand g00656(.dina(w_n860_0[1]),.dinb(w_n290_35[0]),.dout(n862),.clk(gclk));
	jnot g00657(.din(w_n738_0[0]),.dout(n863),.clk(gclk));
	jxor g00658(.dina(w_n732_0[0]),.dinb(w_n305_35[1]),.dout(n864),.clk(gclk));
	jor g00659(.dina(n864),.dinb(w_n796_35[2]),.dout(n865),.clk(gclk));
	jxor g00660(.dina(n865),.dinb(n863),.dout(n866),.clk(gclk));
	jnot g00661(.din(w_n866_0[1]),.dout(n867),.clk(gclk));
	jor g00662(.dina(n867),.dinb(n862),.dout(n868),.clk(gclk));
	jand g00663(.dina(w_n868_0[1]),.dinb(w_n861_0[1]),.dout(n869),.clk(gclk));
	jor g00664(.dina(n869),.dinb(w_n223_35[2]),.dout(n870),.clk(gclk));
	jnot g00665(.din(w_n743_0[0]),.dout(n871),.clk(gclk));
	jor g00666(.dina(n871),.dinb(w_n741_0[0]),.dout(n872),.clk(gclk));
	jor g00667(.dina(n872),.dinb(w_n796_35[1]),.dout(n873),.clk(gclk));
	jxor g00668(.dina(n873),.dinb(w_n752_0[0]),.dout(n874),.clk(gclk));
	jand g00669(.dina(w_n861_0[0]),.dinb(w_n223_35[1]),.dout(n875),.clk(gclk));
	jand g00670(.dina(n875),.dinb(w_n868_0[0]),.dout(n876),.clk(gclk));
	jor g00671(.dina(w_n876_0[1]),.dinb(w_n874_0[1]),.dout(n877),.clk(gclk));
	jand g00672(.dina(w_n877_0[1]),.dinb(w_n870_0[1]),.dout(n878),.clk(gclk));
	jor g00673(.dina(w_n878_0[2]),.dinb(w_n199_41[1]),.dout(n879),.clk(gclk));
	jand g00674(.dina(w_n878_0[1]),.dinb(w_n199_41[0]),.dout(n880),.clk(gclk));
	jnot g00675(.din(w_n759_0[0]),.dout(n881),.clk(gclk));
	jxor g00676(.dina(w_n754_0[0]),.dinb(w_n223_35[0]),.dout(n882),.clk(gclk));
	jor g00677(.dina(n882),.dinb(w_n796_35[0]),.dout(n883),.clk(gclk));
	jxor g00678(.dina(n883),.dinb(n881),.dout(n884),.clk(gclk));
	jnot g00679(.din(n884),.dout(n885),.clk(gclk));
	jor g00680(.dina(w_n885_0[1]),.dinb(n880),.dout(n886),.clk(gclk));
	jand g00681(.dina(n886),.dinb(n879),.dout(n887),.clk(gclk));
	jnot g00682(.din(w_n762_0[0]),.dout(n888),.clk(gclk));
	jand g00683(.dina(w_asqrt53_27[0]),.dinb(n888),.dout(n889),.clk(gclk));
	jand g00684(.dina(w_n889_0[1]),.dinb(w_n769_0[0]),.dout(n890),.clk(gclk));
	jor g00685(.dina(n890),.dinb(w_n767_0[0]),.dout(n891),.clk(gclk));
	jand g00686(.dina(w_n889_0[0]),.dinb(w_n770_0[0]),.dout(n892),.clk(gclk));
	jnot g00687(.din(n892),.dout(n893),.clk(gclk));
	jand g00688(.dina(n893),.dinb(n891),.dout(n894),.clk(gclk));
	jnot g00689(.din(w_n894_0[2]),.dout(n895),.clk(gclk));
	jand g00690(.dina(w_asqrt53_26[2]),.dinb(w_n774_0[2]),.dout(n896),.clk(gclk));
	jand g00691(.dina(w_n896_0[1]),.dinb(w_n771_1[0]),.dout(n897),.clk(gclk));
	jor g00692(.dina(n897),.dinb(w_n816_0[0]),.dout(n898),.clk(gclk));
	jor g00693(.dina(n898),.dinb(w_n895_0[1]),.dout(n899),.clk(gclk));
	jor g00694(.dina(n899),.dinb(w_n887_0[2]),.dout(n900),.clk(gclk));
	jand g00695(.dina(n900),.dinb(w_n194_40[1]),.dout(n901),.clk(gclk));
	jand g00696(.dina(w_n895_0[0]),.dinb(w_n887_0[1]),.dout(n902),.clk(gclk));
	jor g00697(.dina(w_n896_0[0]),.dinb(w_n771_0[2]),.dout(n903),.clk(gclk));
	jand g00698(.dina(w_n774_0[1]),.dinb(w_n771_0[1]),.dout(n904),.clk(gclk));
	jor g00699(.dina(n904),.dinb(w_n194_40[0]),.dout(n905),.clk(gclk));
	jnot g00700(.din(n905),.dout(n906),.clk(gclk));
	jand g00701(.dina(n906),.dinb(n903),.dout(n907),.clk(gclk));
	jor g00702(.dina(w_n907_0[1]),.dinb(w_n902_0[2]),.dout(n910),.clk(gclk));
	jor g00703(.dina(n910),.dinb(w_n901_0[1]),.dout(asqrt_fa_53),.clk(gclk));
	jand g00704(.dina(w_asqrt52_31),.dinb(w_a104_0[0]),.dout(n912),.clk(gclk));
	jnot g00705(.din(w_a102_0[1]),.dout(n913),.clk(gclk));
	jnot g00706(.din(w_a103_0[1]),.dout(n914),.clk(gclk));
	jand g00707(.dina(w_n799_1[0]),.dinb(w_n914_0[1]),.dout(n915),.clk(gclk));
	jand g00708(.dina(n915),.dinb(w_n913_1[1]),.dout(n916),.clk(gclk));
	jor g00709(.dina(n916),.dinb(n912),.dout(n917),.clk(gclk));
	jand g00710(.dina(w_n917_0[2]),.dinb(w_asqrt53_26[1]),.dout(n918),.clk(gclk));
	jand g00711(.dina(w_asqrt52_30[2]),.dinb(w_n799_0[2]),.dout(n919),.clk(gclk));
	jxor g00712(.dina(w_n919_0[1]),.dinb(w_n800_0[1]),.dout(n920),.clk(gclk));
	jor g00713(.dina(w_n917_0[1]),.dinb(w_asqrt53_26[0]),.dout(n921),.clk(gclk));
	jand g00714(.dina(n921),.dinb(w_n920_0[1]),.dout(n922),.clk(gclk));
	jor g00715(.dina(w_n922_0[1]),.dinb(w_n918_0[1]),.dout(n923),.clk(gclk));
	jand g00716(.dina(n923),.dinb(w_asqrt54_27[1]),.dout(n924),.clk(gclk));
	jor g00717(.dina(w_n918_0[0]),.dinb(w_asqrt54_27[0]),.dout(n925),.clk(gclk));
	jor g00718(.dina(n925),.dinb(w_n922_0[0]),.dout(n926),.clk(gclk));
	jand g00719(.dina(w_n919_0[0]),.dinb(w_n800_0[0]),.dout(n927),.clk(gclk));
	jnot g00720(.din(w_n901_0[0]),.dout(n928),.clk(gclk));
	jnot g00721(.din(w_n902_0[1]),.dout(n929),.clk(gclk));
	jnot g00722(.din(w_n907_0[0]),.dout(n930),.clk(gclk));
	jand g00723(.dina(n930),.dinb(w_asqrt53_25[2]),.dout(n931),.clk(gclk));
	jand g00724(.dina(n931),.dinb(n929),.dout(n932),.clk(gclk));
	jand g00725(.dina(n932),.dinb(n928),.dout(n933),.clk(gclk));
	jor g00726(.dina(n933),.dinb(n927),.dout(n934),.clk(gclk));
	jxor g00727(.dina(n934),.dinb(w_n690_0[1]),.dout(n935),.clk(gclk));
	jand g00728(.dina(w_n935_0[1]),.dinb(w_n926_0[1]),.dout(n936),.clk(gclk));
	jor g00729(.dina(n936),.dinb(w_n924_0[1]),.dout(n937),.clk(gclk));
	jand g00730(.dina(w_n937_0[2]),.dinb(w_asqrt55_26[1]),.dout(n938),.clk(gclk));
	jor g00731(.dina(w_n937_0[1]),.dinb(w_asqrt55_26[0]),.dout(n939),.clk(gclk));
	jxor g00732(.dina(w_n804_0[0]),.dinb(w_n791_33[1]),.dout(n940),.clk(gclk));
	jand g00733(.dina(n940),.dinb(w_asqrt52_30[1]),.dout(n941),.clk(gclk));
	jxor g00734(.dina(n941),.dinb(w_n807_0[0]),.dout(n942),.clk(gclk));
	jnot g00735(.din(w_n942_0[1]),.dout(n943),.clk(gclk));
	jand g00736(.dina(n943),.dinb(n939),.dout(n944),.clk(gclk));
	jor g00737(.dina(w_n944_0[1]),.dinb(w_n938_0[1]),.dout(n945),.clk(gclk));
	jand g00738(.dina(n945),.dinb(w_asqrt56_27[1]),.dout(n946),.clk(gclk));
	jnot g00739(.din(w_n813_0[0]),.dout(n947),.clk(gclk));
	jand g00740(.dina(n947),.dinb(w_n811_0[0]),.dout(n948),.clk(gclk));
	jand g00741(.dina(n948),.dinb(w_asqrt52_30[0]),.dout(n949),.clk(gclk));
	jxor g00742(.dina(n949),.dinb(w_n821_0[0]),.dout(n950),.clk(gclk));
	jnot g00743(.din(n950),.dout(n951),.clk(gclk));
	jor g00744(.dina(w_n938_0[0]),.dinb(w_asqrt56_27[0]),.dout(n952),.clk(gclk));
	jor g00745(.dina(n952),.dinb(w_n944_0[0]),.dout(n953),.clk(gclk));
	jand g00746(.dina(w_n953_0[1]),.dinb(w_n951_0[1]),.dout(n954),.clk(gclk));
	jor g00747(.dina(w_n954_0[1]),.dinb(w_n946_0[1]),.dout(n955),.clk(gclk));
	jand g00748(.dina(w_n955_0[2]),.dinb(w_asqrt57_26[2]),.dout(n956),.clk(gclk));
	jor g00749(.dina(w_n955_0[1]),.dinb(w_asqrt57_26[1]),.dout(n957),.clk(gclk));
	jnot g00750(.din(w_n828_0[0]),.dout(n958),.clk(gclk));
	jxor g00751(.dina(w_n823_0[0]),.dinb(w_n590_33[2]),.dout(n959),.clk(gclk));
	jand g00752(.dina(n959),.dinb(w_asqrt52_29[2]),.dout(n960),.clk(gclk));
	jxor g00753(.dina(n960),.dinb(n958),.dout(n961),.clk(gclk));
	jand g00754(.dina(w_n961_0[1]),.dinb(n957),.dout(n962),.clk(gclk));
	jor g00755(.dina(w_n962_0[1]),.dinb(w_n956_0[1]),.dout(n963),.clk(gclk));
	jand g00756(.dina(n963),.dinb(w_asqrt58_27[1]),.dout(n964),.clk(gclk));
	jor g00757(.dina(w_n956_0[0]),.dinb(w_asqrt58_27[0]),.dout(n965),.clk(gclk));
	jor g00758(.dina(n965),.dinb(w_n962_0[0]),.dout(n966),.clk(gclk));
	jnot g00759(.din(w_n835_0[0]),.dout(n967),.clk(gclk));
	jnot g00760(.din(w_n837_0[0]),.dout(n968),.clk(gclk));
	jand g00761(.dina(w_asqrt52_29[1]),.dinb(w_n831_0[0]),.dout(n969),.clk(gclk));
	jand g00762(.dina(w_n969_0[1]),.dinb(n968),.dout(n970),.clk(gclk));
	jor g00763(.dina(n970),.dinb(n967),.dout(n971),.clk(gclk));
	jnot g00764(.din(w_n838_0[0]),.dout(n972),.clk(gclk));
	jand g00765(.dina(w_n969_0[0]),.dinb(n972),.dout(n973),.clk(gclk));
	jnot g00766(.din(n973),.dout(n974),.clk(gclk));
	jand g00767(.dina(n974),.dinb(n971),.dout(n975),.clk(gclk));
	jand g00768(.dina(w_n975_0[1]),.dinb(w_n966_0[1]),.dout(n976),.clk(gclk));
	jor g00769(.dina(n976),.dinb(w_n964_0[1]),.dout(n977),.clk(gclk));
	jand g00770(.dina(w_n977_0[2]),.dinb(w_asqrt59_27[0]),.dout(n978),.clk(gclk));
	jor g00771(.dina(w_n977_0[1]),.dinb(w_asqrt59_26[2]),.dout(n979),.clk(gclk));
	jxor g00772(.dina(w_n839_0[0]),.dinb(w_n425_33[2]),.dout(n980),.clk(gclk));
	jand g00773(.dina(n980),.dinb(w_asqrt52_29[0]),.dout(n981),.clk(gclk));
	jxor g00774(.dina(n981),.dinb(w_n844_0[0]),.dout(n982),.clk(gclk));
	jand g00775(.dina(w_n982_0[1]),.dinb(n979),.dout(n983),.clk(gclk));
	jor g00776(.dina(w_n983_0[1]),.dinb(w_n978_0[1]),.dout(n984),.clk(gclk));
	jand g00777(.dina(n984),.dinb(w_asqrt60_27[0]),.dout(n985),.clk(gclk));
	jnot g00778(.din(w_n850_0[0]),.dout(n986),.clk(gclk));
	jand g00779(.dina(n986),.dinb(w_n848_0[0]),.dout(n987),.clk(gclk));
	jand g00780(.dina(n987),.dinb(w_asqrt52_28[2]),.dout(n988),.clk(gclk));
	jxor g00781(.dina(n988),.dinb(w_n858_0[0]),.dout(n989),.clk(gclk));
	jnot g00782(.din(n989),.dout(n990),.clk(gclk));
	jor g00783(.dina(w_n978_0[0]),.dinb(w_asqrt60_26[2]),.dout(n991),.clk(gclk));
	jor g00784(.dina(n991),.dinb(w_n983_0[0]),.dout(n992),.clk(gclk));
	jand g00785(.dina(w_n992_0[1]),.dinb(w_n990_0[1]),.dout(n993),.clk(gclk));
	jor g00786(.dina(w_n993_0[1]),.dinb(w_n985_0[1]),.dout(n994),.clk(gclk));
	jand g00787(.dina(w_n994_0[2]),.dinb(w_asqrt61_27[1]),.dout(n995),.clk(gclk));
	jor g00788(.dina(w_n994_0[1]),.dinb(w_asqrt61_27[0]),.dout(n996),.clk(gclk));
	jxor g00789(.dina(w_n860_0[0]),.dinb(w_n290_34[2]),.dout(n997),.clk(gclk));
	jand g00790(.dina(n997),.dinb(w_asqrt52_28[1]),.dout(n998),.clk(gclk));
	jxor g00791(.dina(n998),.dinb(w_n866_0[0]),.dout(n999),.clk(gclk));
	jand g00792(.dina(w_n999_0[1]),.dinb(n996),.dout(n1000),.clk(gclk));
	jor g00793(.dina(w_n1000_0[1]),.dinb(w_n995_0[1]),.dout(n1001),.clk(gclk));
	jand g00794(.dina(n1001),.dinb(w_asqrt62_27[1]),.dout(n1002),.clk(gclk));
	jor g00795(.dina(w_n995_0[0]),.dinb(w_asqrt62_27[0]),.dout(n1003),.clk(gclk));
	jor g00796(.dina(n1003),.dinb(w_n1000_0[0]),.dout(n1004),.clk(gclk));
	jnot g00797(.din(w_n874_0[0]),.dout(n1005),.clk(gclk));
	jnot g00798(.din(w_n876_0[0]),.dout(n1006),.clk(gclk));
	jand g00799(.dina(w_asqrt52_28[0]),.dinb(w_n870_0[0]),.dout(n1007),.clk(gclk));
	jand g00800(.dina(w_n1007_0[1]),.dinb(n1006),.dout(n1008),.clk(gclk));
	jor g00801(.dina(n1008),.dinb(n1005),.dout(n1009),.clk(gclk));
	jnot g00802(.din(w_n877_0[0]),.dout(n1010),.clk(gclk));
	jand g00803(.dina(w_n1007_0[0]),.dinb(n1010),.dout(n1011),.clk(gclk));
	jnot g00804(.din(n1011),.dout(n1012),.clk(gclk));
	jand g00805(.dina(n1012),.dinb(n1009),.dout(n1013),.clk(gclk));
	jand g00806(.dina(w_n1013_0[1]),.dinb(w_n1004_0[1]),.dout(n1014),.clk(gclk));
	jor g00807(.dina(n1014),.dinb(w_n1002_0[1]),.dout(n1015),.clk(gclk));
	jxor g00808(.dina(w_n878_0[0]),.dinb(w_n199_40[2]),.dout(n1016),.clk(gclk));
	jand g00809(.dina(n1016),.dinb(w_asqrt52_27[2]),.dout(n1017),.clk(gclk));
	jxor g00810(.dina(n1017),.dinb(w_n885_0[0]),.dout(n1018),.clk(gclk));
	jnot g00811(.din(w_n887_0[0]),.dout(n1019),.clk(gclk));
	jand g00812(.dina(w_asqrt52_27[1]),.dinb(w_n894_0[1]),.dout(n1020),.clk(gclk));
	jand g00813(.dina(w_n1020_0[1]),.dinb(w_n1019_0[2]),.dout(n1021),.clk(gclk));
	jor g00814(.dina(n1021),.dinb(w_n902_0[0]),.dout(n1022),.clk(gclk));
	jor g00815(.dina(n1022),.dinb(w_n1018_0[1]),.dout(n1023),.clk(gclk));
	jnot g00816(.din(n1023),.dout(n1024),.clk(gclk));
	jand g00817(.dina(n1024),.dinb(w_n1015_1[2]),.dout(n1025),.clk(gclk));
	jor g00818(.dina(n1025),.dinb(w_asqrt63_14[1]),.dout(n1026),.clk(gclk));
	jnot g00819(.din(w_n1018_0[0]),.dout(n1027),.clk(gclk));
	jor g00820(.dina(w_n1027_0[2]),.dinb(w_n1015_1[1]),.dout(n1028),.clk(gclk));
	jor g00821(.dina(w_n1020_0[0]),.dinb(w_n1019_0[1]),.dout(n1029),.clk(gclk));
	jand g00822(.dina(w_n894_0[0]),.dinb(w_n1019_0[0]),.dout(n1030),.clk(gclk));
	jor g00823(.dina(n1030),.dinb(w_n194_39[2]),.dout(n1031),.clk(gclk));
	jnot g00824(.din(n1031),.dout(n1032),.clk(gclk));
	jand g00825(.dina(n1032),.dinb(n1029),.dout(n1033),.clk(gclk));
	jnot g00826(.din(w_asqrt52_27[0]),.dout(n1034),.clk(gclk));
	jnot g00827(.din(w_n1033_0[1]),.dout(n1037),.clk(gclk));
	jand g00828(.dina(n1037),.dinb(w_n1028_0[1]),.dout(n1038),.clk(gclk));
	jand g00829(.dina(n1038),.dinb(w_n1026_0[1]),.dout(n1039),.clk(gclk));
	jnot g00830(.din(w_n1039_37[2]),.dout(asqrt_fa_52),.clk(gclk));
	jor g00831(.dina(w_n1039_37[1]),.dinb(w_n913_1[0]),.dout(n1041),.clk(gclk));
	jnot g00832(.din(w_a100_0[1]),.dout(n1042),.clk(gclk));
	jnot g00833(.din(a[101]),.dout(n1043),.clk(gclk));
	jand g00834(.dina(w_n913_0[2]),.dinb(w_n1043_0[2]),.dout(n1044),.clk(gclk));
	jand g00835(.dina(n1044),.dinb(w_n1042_1[1]),.dout(n1045),.clk(gclk));
	jnot g00836(.din(n1045),.dout(n1046),.clk(gclk));
	jand g00837(.dina(n1046),.dinb(n1041),.dout(n1047),.clk(gclk));
	jor g00838(.dina(w_n1047_0[2]),.dinb(w_n1034_33[1]),.dout(n1048),.clk(gclk));
	jor g00839(.dina(w_n1039_37[0]),.dinb(w_a102_0[0]),.dout(n1049),.clk(gclk));
	jxor g00840(.dina(w_n1049_0[1]),.dinb(w_n914_0[0]),.dout(n1050),.clk(gclk));
	jand g00841(.dina(w_n1047_0[1]),.dinb(w_n1034_33[0]),.dout(n1051),.clk(gclk));
	jor g00842(.dina(n1051),.dinb(w_n1050_0[1]),.dout(n1052),.clk(gclk));
	jand g00843(.dina(w_n1052_0[1]),.dinb(w_n1048_0[1]),.dout(n1053),.clk(gclk));
	jor g00844(.dina(n1053),.dinb(w_n796_34[2]),.dout(n1054),.clk(gclk));
	jand g00845(.dina(w_n1048_0[0]),.dinb(w_n796_34[1]),.dout(n1055),.clk(gclk));
	jand g00846(.dina(n1055),.dinb(w_n1052_0[0]),.dout(n1056),.clk(gclk));
	jor g00847(.dina(w_n1049_0[0]),.dinb(w_a103_0[0]),.dout(n1057),.clk(gclk));
	jnot g00848(.din(w_n1026_0[0]),.dout(n1058),.clk(gclk));
	jnot g00849(.din(w_n1028_0[0]),.dout(n1059),.clk(gclk));
	jor g00850(.dina(w_n1033_0[0]),.dinb(w_n1034_32[2]),.dout(n1060),.clk(gclk));
	jor g00851(.dina(n1060),.dinb(w_n1059_0[1]),.dout(n1061),.clk(gclk));
	jor g00852(.dina(n1061),.dinb(n1058),.dout(n1062),.clk(gclk));
	jand g00853(.dina(n1062),.dinb(n1057),.dout(n1063),.clk(gclk));
	jxor g00854(.dina(n1063),.dinb(w_n799_0[1]),.dout(n1064),.clk(gclk));
	jor g00855(.dina(w_n1064_0[1]),.dinb(w_n1056_0[1]),.dout(n1065),.clk(gclk));
	jand g00856(.dina(n1065),.dinb(w_n1054_0[1]),.dout(n1066),.clk(gclk));
	jor g00857(.dina(w_n1066_0[2]),.dinb(w_n791_33[0]),.dout(n1067),.clk(gclk));
	jand g00858(.dina(w_n1066_0[1]),.dinb(w_n791_32[2]),.dout(n1068),.clk(gclk));
	jxor g00859(.dina(w_n917_0[0]),.dinb(w_n796_34[0]),.dout(n1069),.clk(gclk));
	jor g00860(.dina(n1069),.dinb(w_n1039_36[2]),.dout(n1070),.clk(gclk));
	jxor g00861(.dina(n1070),.dinb(w_n920_0[0]),.dout(n1071),.clk(gclk));
	jor g00862(.dina(w_n1071_0[1]),.dinb(n1068),.dout(n1072),.clk(gclk));
	jand g00863(.dina(w_n1072_0[1]),.dinb(w_n1067_0[1]),.dout(n1073),.clk(gclk));
	jor g00864(.dina(n1073),.dinb(w_n595_35[0]),.dout(n1074),.clk(gclk));
	jnot g00865(.din(w_n926_0[0]),.dout(n1075),.clk(gclk));
	jor g00866(.dina(n1075),.dinb(w_n924_0[0]),.dout(n1076),.clk(gclk));
	jor g00867(.dina(n1076),.dinb(w_n1039_36[1]),.dout(n1077),.clk(gclk));
	jxor g00868(.dina(n1077),.dinb(w_n935_0[0]),.dout(n1078),.clk(gclk));
	jand g00869(.dina(w_n1067_0[0]),.dinb(w_n595_34[2]),.dout(n1079),.clk(gclk));
	jand g00870(.dina(n1079),.dinb(w_n1072_0[0]),.dout(n1080),.clk(gclk));
	jor g00871(.dina(w_n1080_0[1]),.dinb(w_n1078_0[1]),.dout(n1081),.clk(gclk));
	jand g00872(.dina(w_n1081_0[1]),.dinb(w_n1074_0[1]),.dout(n1082),.clk(gclk));
	jor g00873(.dina(w_n1082_0[2]),.dinb(w_n590_33[1]),.dout(n1083),.clk(gclk));
	jand g00874(.dina(w_n1082_0[1]),.dinb(w_n590_33[0]),.dout(n1084),.clk(gclk));
	jxor g00875(.dina(w_n937_0[0]),.dinb(w_n595_34[1]),.dout(n1085),.clk(gclk));
	jor g00876(.dina(n1085),.dinb(w_n1039_36[0]),.dout(n1086),.clk(gclk));
	jxor g00877(.dina(n1086),.dinb(w_n942_0[0]),.dout(n1087),.clk(gclk));
	jnot g00878(.din(w_n1087_0[1]),.dout(n1088),.clk(gclk));
	jor g00879(.dina(n1088),.dinb(n1084),.dout(n1089),.clk(gclk));
	jand g00880(.dina(w_n1089_0[1]),.dinb(w_n1083_0[1]),.dout(n1090),.clk(gclk));
	jor g00881(.dina(n1090),.dinb(w_n430_34[2]),.dout(n1091),.clk(gclk));
	jand g00882(.dina(w_n1083_0[0]),.dinb(w_n430_34[1]),.dout(n1092),.clk(gclk));
	jand g00883(.dina(n1092),.dinb(w_n1089_0[0]),.dout(n1093),.clk(gclk));
	jnot g00884(.din(w_n946_0[0]),.dout(n1094),.clk(gclk));
	jand g00885(.dina(w_asqrt51_26[1]),.dinb(n1094),.dout(n1095),.clk(gclk));
	jand g00886(.dina(w_n1095_0[1]),.dinb(w_n953_0[0]),.dout(n1096),.clk(gclk));
	jor g00887(.dina(n1096),.dinb(w_n951_0[0]),.dout(n1097),.clk(gclk));
	jand g00888(.dina(w_n1095_0[0]),.dinb(w_n954_0[0]),.dout(n1098),.clk(gclk));
	jnot g00889(.din(n1098),.dout(n1099),.clk(gclk));
	jand g00890(.dina(n1099),.dinb(n1097),.dout(n1100),.clk(gclk));
	jnot g00891(.din(n1100),.dout(n1101),.clk(gclk));
	jor g00892(.dina(w_n1101_0[1]),.dinb(w_n1093_0[1]),.dout(n1102),.clk(gclk));
	jand g00893(.dina(n1102),.dinb(w_n1091_0[1]),.dout(n1103),.clk(gclk));
	jor g00894(.dina(w_n1103_0[2]),.dinb(w_n425_33[1]),.dout(n1104),.clk(gclk));
	jand g00895(.dina(w_n1103_0[1]),.dinb(w_n425_33[0]),.dout(n1105),.clk(gclk));
	jnot g00896(.din(w_n961_0[0]),.dout(n1106),.clk(gclk));
	jxor g00897(.dina(w_n955_0[0]),.dinb(w_n430_34[0]),.dout(n1107),.clk(gclk));
	jor g00898(.dina(n1107),.dinb(w_n1039_35[2]),.dout(n1108),.clk(gclk));
	jxor g00899(.dina(n1108),.dinb(n1106),.dout(n1109),.clk(gclk));
	jnot g00900(.din(w_n1109_0[1]),.dout(n1110),.clk(gclk));
	jor g00901(.dina(n1110),.dinb(n1105),.dout(n1111),.clk(gclk));
	jand g00902(.dina(w_n1111_0[1]),.dinb(w_n1104_0[1]),.dout(n1112),.clk(gclk));
	jor g00903(.dina(n1112),.dinb(w_n305_35[0]),.dout(n1113),.clk(gclk));
	jnot g00904(.din(w_n966_0[0]),.dout(n1114),.clk(gclk));
	jor g00905(.dina(n1114),.dinb(w_n964_0[0]),.dout(n1115),.clk(gclk));
	jor g00906(.dina(n1115),.dinb(w_n1039_35[1]),.dout(n1116),.clk(gclk));
	jxor g00907(.dina(n1116),.dinb(w_n975_0[0]),.dout(n1117),.clk(gclk));
	jand g00908(.dina(w_n1104_0[0]),.dinb(w_n305_34[2]),.dout(n1118),.clk(gclk));
	jand g00909(.dina(n1118),.dinb(w_n1111_0[0]),.dout(n1119),.clk(gclk));
	jor g00910(.dina(w_n1119_0[1]),.dinb(w_n1117_0[1]),.dout(n1120),.clk(gclk));
	jand g00911(.dina(w_n1120_0[1]),.dinb(w_n1113_0[1]),.dout(n1121),.clk(gclk));
	jor g00912(.dina(w_n1121_0[2]),.dinb(w_n290_34[1]),.dout(n1122),.clk(gclk));
	jand g00913(.dina(w_n1121_0[1]),.dinb(w_n290_34[0]),.dout(n1123),.clk(gclk));
	jnot g00914(.din(w_n982_0[0]),.dout(n1124),.clk(gclk));
	jxor g00915(.dina(w_n977_0[0]),.dinb(w_n305_34[1]),.dout(n1125),.clk(gclk));
	jor g00916(.dina(n1125),.dinb(w_n1039_35[0]),.dout(n1126),.clk(gclk));
	jxor g00917(.dina(n1126),.dinb(n1124),.dout(n1127),.clk(gclk));
	jnot g00918(.din(n1127),.dout(n1128),.clk(gclk));
	jor g00919(.dina(w_n1128_0[1]),.dinb(n1123),.dout(n1129),.clk(gclk));
	jand g00920(.dina(w_n1129_0[1]),.dinb(w_n1122_0[1]),.dout(n1130),.clk(gclk));
	jor g00921(.dina(n1130),.dinb(w_n223_34[2]),.dout(n1131),.clk(gclk));
	jand g00922(.dina(w_n1122_0[0]),.dinb(w_n223_34[1]),.dout(n1132),.clk(gclk));
	jand g00923(.dina(n1132),.dinb(w_n1129_0[0]),.dout(n1133),.clk(gclk));
	jnot g00924(.din(w_n985_0[0]),.dout(n1134),.clk(gclk));
	jand g00925(.dina(w_asqrt51_26[0]),.dinb(n1134),.dout(n1135),.clk(gclk));
	jand g00926(.dina(w_n1135_0[1]),.dinb(w_n992_0[0]),.dout(n1136),.clk(gclk));
	jor g00927(.dina(n1136),.dinb(w_n990_0[0]),.dout(n1137),.clk(gclk));
	jand g00928(.dina(w_n1135_0[0]),.dinb(w_n993_0[0]),.dout(n1138),.clk(gclk));
	jnot g00929(.din(n1138),.dout(n1139),.clk(gclk));
	jand g00930(.dina(n1139),.dinb(n1137),.dout(n1140),.clk(gclk));
	jnot g00931(.din(n1140),.dout(n1141),.clk(gclk));
	jor g00932(.dina(w_n1141_0[1]),.dinb(w_n1133_0[1]),.dout(n1142),.clk(gclk));
	jand g00933(.dina(n1142),.dinb(w_n1131_0[1]),.dout(n1143),.clk(gclk));
	jor g00934(.dina(w_n1143_0[2]),.dinb(w_n199_40[1]),.dout(n1144),.clk(gclk));
	jand g00935(.dina(w_n1143_0[1]),.dinb(w_n199_40[0]),.dout(n1145),.clk(gclk));
	jxor g00936(.dina(w_n994_0[0]),.dinb(w_n223_34[0]),.dout(n1146),.clk(gclk));
	jor g00937(.dina(n1146),.dinb(w_n1039_34[2]),.dout(n1147),.clk(gclk));
	jxor g00938(.dina(n1147),.dinb(w_n999_0[0]),.dout(n1148),.clk(gclk));
	jor g00939(.dina(w_n1148_0[1]),.dinb(n1145),.dout(n1149),.clk(gclk));
	jand g00940(.dina(n1149),.dinb(n1144),.dout(n1150),.clk(gclk));
	jnot g00941(.din(w_n1004_0[0]),.dout(n1151),.clk(gclk));
	jor g00942(.dina(n1151),.dinb(w_n1002_0[0]),.dout(n1152),.clk(gclk));
	jor g00943(.dina(n1152),.dinb(w_n1039_34[1]),.dout(n1153),.clk(gclk));
	jxor g00944(.dina(n1153),.dinb(w_n1013_0[0]),.dout(n1154),.clk(gclk));
	jand g00945(.dina(w_asqrt51_25[2]),.dinb(w_n1027_0[1]),.dout(n1155),.clk(gclk));
	jand g00946(.dina(w_n1155_0[1]),.dinb(w_n1015_1[0]),.dout(n1156),.clk(gclk));
	jor g00947(.dina(n1156),.dinb(w_n1059_0[0]),.dout(n1157),.clk(gclk));
	jor g00948(.dina(n1157),.dinb(w_n1154_0[2]),.dout(n1158),.clk(gclk));
	jor g00949(.dina(n1158),.dinb(w_n1150_0[2]),.dout(n1159),.clk(gclk));
	jand g00950(.dina(n1159),.dinb(w_n194_39[1]),.dout(n1160),.clk(gclk));
	jand g00951(.dina(w_n1154_0[1]),.dinb(w_n1150_0[1]),.dout(n1161),.clk(gclk));
	jor g00952(.dina(w_n1155_0[0]),.dinb(w_n1015_0[2]),.dout(n1162),.clk(gclk));
	jand g00953(.dina(w_n1027_0[0]),.dinb(w_n1015_0[1]),.dout(n1163),.clk(gclk));
	jor g00954(.dina(n1163),.dinb(w_n194_39[0]),.dout(n1164),.clk(gclk));
	jnot g00955(.din(n1164),.dout(n1165),.clk(gclk));
	jand g00956(.dina(n1165),.dinb(n1162),.dout(n1166),.clk(gclk));
	jor g00957(.dina(w_n1166_0[1]),.dinb(w_n1161_0[2]),.dout(n1169),.clk(gclk));
	jor g00958(.dina(n1169),.dinb(w_n1160_0[1]),.dout(asqrt_fa_51),.clk(gclk));
	jand g00959(.dina(w_asqrt50_31),.dinb(w_a100_0[0]),.dout(n1171),.clk(gclk));
	jnot g00960(.din(w_a98_0[1]),.dout(n1172),.clk(gclk));
	jnot g00961(.din(w_a99_0[1]),.dout(n1173),.clk(gclk));
	jand g00962(.dina(w_n1042_1[0]),.dinb(w_n1173_0[1]),.dout(n1174),.clk(gclk));
	jand g00963(.dina(n1174),.dinb(w_n1172_1[1]),.dout(n1175),.clk(gclk));
	jor g00964(.dina(n1175),.dinb(n1171),.dout(n1176),.clk(gclk));
	jand g00965(.dina(w_n1176_0[2]),.dinb(w_asqrt51_25[1]),.dout(n1177),.clk(gclk));
	jand g00966(.dina(w_asqrt50_30[2]),.dinb(w_n1042_0[2]),.dout(n1178),.clk(gclk));
	jxor g00967(.dina(w_n1178_0[1]),.dinb(w_n1043_0[1]),.dout(n1179),.clk(gclk));
	jor g00968(.dina(w_n1176_0[1]),.dinb(w_asqrt51_25[0]),.dout(n1180),.clk(gclk));
	jand g00969(.dina(n1180),.dinb(w_n1179_0[1]),.dout(n1181),.clk(gclk));
	jor g00970(.dina(w_n1181_0[1]),.dinb(w_n1177_0[1]),.dout(n1182),.clk(gclk));
	jand g00971(.dina(n1182),.dinb(w_asqrt52_26[2]),.dout(n1183),.clk(gclk));
	jor g00972(.dina(w_n1177_0[0]),.dinb(w_asqrt52_26[1]),.dout(n1184),.clk(gclk));
	jor g00973(.dina(n1184),.dinb(w_n1181_0[0]),.dout(n1185),.clk(gclk));
	jand g00974(.dina(w_n1178_0[0]),.dinb(w_n1043_0[0]),.dout(n1186),.clk(gclk));
	jnot g00975(.din(w_n1160_0[0]),.dout(n1187),.clk(gclk));
	jnot g00976(.din(w_n1161_0[1]),.dout(n1188),.clk(gclk));
	jnot g00977(.din(w_n1166_0[0]),.dout(n1189),.clk(gclk));
	jand g00978(.dina(n1189),.dinb(w_asqrt51_24[2]),.dout(n1190),.clk(gclk));
	jand g00979(.dina(n1190),.dinb(n1188),.dout(n1191),.clk(gclk));
	jand g00980(.dina(n1191),.dinb(n1187),.dout(n1192),.clk(gclk));
	jor g00981(.dina(n1192),.dinb(n1186),.dout(n1193),.clk(gclk));
	jxor g00982(.dina(n1193),.dinb(w_n913_0[1]),.dout(n1194),.clk(gclk));
	jand g00983(.dina(w_n1194_0[1]),.dinb(w_n1185_0[1]),.dout(n1195),.clk(gclk));
	jor g00984(.dina(n1195),.dinb(w_n1183_0[1]),.dout(n1196),.clk(gclk));
	jand g00985(.dina(w_n1196_0[2]),.dinb(w_asqrt53_25[1]),.dout(n1197),.clk(gclk));
	jor g00986(.dina(w_n1196_0[1]),.dinb(w_asqrt53_25[0]),.dout(n1198),.clk(gclk));
	jxor g00987(.dina(w_n1047_0[0]),.dinb(w_n1034_32[1]),.dout(n1199),.clk(gclk));
	jand g00988(.dina(n1199),.dinb(w_asqrt50_30[1]),.dout(n1200),.clk(gclk));
	jxor g00989(.dina(n1200),.dinb(w_n1050_0[0]),.dout(n1201),.clk(gclk));
	jnot g00990(.din(w_n1201_0[1]),.dout(n1202),.clk(gclk));
	jand g00991(.dina(n1202),.dinb(n1198),.dout(n1203),.clk(gclk));
	jor g00992(.dina(w_n1203_0[1]),.dinb(w_n1197_0[1]),.dout(n1204),.clk(gclk));
	jand g00993(.dina(n1204),.dinb(w_asqrt54_26[2]),.dout(n1205),.clk(gclk));
	jnot g00994(.din(w_n1056_0[0]),.dout(n1206),.clk(gclk));
	jand g00995(.dina(n1206),.dinb(w_n1054_0[0]),.dout(n1207),.clk(gclk));
	jand g00996(.dina(n1207),.dinb(w_asqrt50_30[0]),.dout(n1208),.clk(gclk));
	jxor g00997(.dina(n1208),.dinb(w_n1064_0[0]),.dout(n1209),.clk(gclk));
	jnot g00998(.din(n1209),.dout(n1210),.clk(gclk));
	jor g00999(.dina(w_n1197_0[0]),.dinb(w_asqrt54_26[1]),.dout(n1211),.clk(gclk));
	jor g01000(.dina(n1211),.dinb(w_n1203_0[0]),.dout(n1212),.clk(gclk));
	jand g01001(.dina(w_n1212_0[1]),.dinb(w_n1210_0[1]),.dout(n1213),.clk(gclk));
	jor g01002(.dina(w_n1213_0[1]),.dinb(w_n1205_0[1]),.dout(n1214),.clk(gclk));
	jand g01003(.dina(w_n1214_0[2]),.dinb(w_asqrt55_25[2]),.dout(n1215),.clk(gclk));
	jor g01004(.dina(w_n1214_0[1]),.dinb(w_asqrt55_25[1]),.dout(n1216),.clk(gclk));
	jnot g01005(.din(w_n1071_0[0]),.dout(n1217),.clk(gclk));
	jxor g01006(.dina(w_n1066_0[0]),.dinb(w_n791_32[1]),.dout(n1218),.clk(gclk));
	jand g01007(.dina(n1218),.dinb(w_asqrt50_29[2]),.dout(n1219),.clk(gclk));
	jxor g01008(.dina(n1219),.dinb(n1217),.dout(n1220),.clk(gclk));
	jand g01009(.dina(w_n1220_0[1]),.dinb(n1216),.dout(n1221),.clk(gclk));
	jor g01010(.dina(w_n1221_0[1]),.dinb(w_n1215_0[1]),.dout(n1222),.clk(gclk));
	jand g01011(.dina(n1222),.dinb(w_asqrt56_26[2]),.dout(n1223),.clk(gclk));
	jor g01012(.dina(w_n1215_0[0]),.dinb(w_asqrt56_26[1]),.dout(n1224),.clk(gclk));
	jor g01013(.dina(n1224),.dinb(w_n1221_0[0]),.dout(n1225),.clk(gclk));
	jnot g01014(.din(w_n1078_0[0]),.dout(n1226),.clk(gclk));
	jnot g01015(.din(w_n1080_0[0]),.dout(n1227),.clk(gclk));
	jand g01016(.dina(w_asqrt50_29[1]),.dinb(w_n1074_0[0]),.dout(n1228),.clk(gclk));
	jand g01017(.dina(w_n1228_0[1]),.dinb(n1227),.dout(n1229),.clk(gclk));
	jor g01018(.dina(n1229),.dinb(n1226),.dout(n1230),.clk(gclk));
	jnot g01019(.din(w_n1081_0[0]),.dout(n1231),.clk(gclk));
	jand g01020(.dina(w_n1228_0[0]),.dinb(n1231),.dout(n1232),.clk(gclk));
	jnot g01021(.din(n1232),.dout(n1233),.clk(gclk));
	jand g01022(.dina(n1233),.dinb(n1230),.dout(n1234),.clk(gclk));
	jand g01023(.dina(w_n1234_0[1]),.dinb(w_n1225_0[1]),.dout(n1235),.clk(gclk));
	jor g01024(.dina(n1235),.dinb(w_n1223_0[1]),.dout(n1236),.clk(gclk));
	jand g01025(.dina(w_n1236_0[2]),.dinb(w_asqrt57_26[0]),.dout(n1237),.clk(gclk));
	jor g01026(.dina(w_n1236_0[1]),.dinb(w_asqrt57_25[2]),.dout(n1238),.clk(gclk));
	jxor g01027(.dina(w_n1082_0[0]),.dinb(w_n590_32[2]),.dout(n1239),.clk(gclk));
	jand g01028(.dina(n1239),.dinb(w_asqrt50_29[0]),.dout(n1240),.clk(gclk));
	jxor g01029(.dina(n1240),.dinb(w_n1087_0[0]),.dout(n1241),.clk(gclk));
	jand g01030(.dina(w_n1241_0[1]),.dinb(n1238),.dout(n1242),.clk(gclk));
	jor g01031(.dina(w_n1242_0[1]),.dinb(w_n1237_0[1]),.dout(n1243),.clk(gclk));
	jand g01032(.dina(n1243),.dinb(w_asqrt58_26[2]),.dout(n1244),.clk(gclk));
	jnot g01033(.din(w_n1093_0[0]),.dout(n1245),.clk(gclk));
	jand g01034(.dina(n1245),.dinb(w_n1091_0[0]),.dout(n1246),.clk(gclk));
	jand g01035(.dina(n1246),.dinb(w_asqrt50_28[2]),.dout(n1247),.clk(gclk));
	jxor g01036(.dina(n1247),.dinb(w_n1101_0[0]),.dout(n1248),.clk(gclk));
	jnot g01037(.din(n1248),.dout(n1249),.clk(gclk));
	jor g01038(.dina(w_n1237_0[0]),.dinb(w_asqrt58_26[1]),.dout(n1250),.clk(gclk));
	jor g01039(.dina(n1250),.dinb(w_n1242_0[0]),.dout(n1251),.clk(gclk));
	jand g01040(.dina(w_n1251_0[1]),.dinb(w_n1249_0[1]),.dout(n1252),.clk(gclk));
	jor g01041(.dina(w_n1252_0[1]),.dinb(w_n1244_0[1]),.dout(n1253),.clk(gclk));
	jand g01042(.dina(w_n1253_0[2]),.dinb(w_asqrt59_26[1]),.dout(n1254),.clk(gclk));
	jor g01043(.dina(w_n1253_0[1]),.dinb(w_asqrt59_26[0]),.dout(n1255),.clk(gclk));
	jxor g01044(.dina(w_n1103_0[0]),.dinb(w_n425_32[2]),.dout(n1256),.clk(gclk));
	jand g01045(.dina(n1256),.dinb(w_asqrt50_28[1]),.dout(n1257),.clk(gclk));
	jxor g01046(.dina(n1257),.dinb(w_n1109_0[0]),.dout(n1258),.clk(gclk));
	jand g01047(.dina(w_n1258_0[1]),.dinb(n1255),.dout(n1259),.clk(gclk));
	jor g01048(.dina(w_n1259_0[1]),.dinb(w_n1254_0[1]),.dout(n1260),.clk(gclk));
	jand g01049(.dina(n1260),.dinb(w_asqrt60_26[1]),.dout(n1261),.clk(gclk));
	jor g01050(.dina(w_n1254_0[0]),.dinb(w_asqrt60_26[0]),.dout(n1262),.clk(gclk));
	jor g01051(.dina(n1262),.dinb(w_n1259_0[0]),.dout(n1263),.clk(gclk));
	jnot g01052(.din(w_n1117_0[0]),.dout(n1264),.clk(gclk));
	jnot g01053(.din(w_n1119_0[0]),.dout(n1265),.clk(gclk));
	jand g01054(.dina(w_asqrt50_28[0]),.dinb(w_n1113_0[0]),.dout(n1266),.clk(gclk));
	jand g01055(.dina(w_n1266_0[1]),.dinb(n1265),.dout(n1267),.clk(gclk));
	jor g01056(.dina(n1267),.dinb(n1264),.dout(n1268),.clk(gclk));
	jnot g01057(.din(w_n1120_0[0]),.dout(n1269),.clk(gclk));
	jand g01058(.dina(w_n1266_0[0]),.dinb(n1269),.dout(n1270),.clk(gclk));
	jnot g01059(.din(n1270),.dout(n1271),.clk(gclk));
	jand g01060(.dina(n1271),.dinb(n1268),.dout(n1272),.clk(gclk));
	jand g01061(.dina(w_n1272_0[1]),.dinb(w_n1263_0[1]),.dout(n1273),.clk(gclk));
	jor g01062(.dina(n1273),.dinb(w_n1261_0[1]),.dout(n1274),.clk(gclk));
	jand g01063(.dina(w_n1274_0[1]),.dinb(w_asqrt61_26[2]),.dout(n1275),.clk(gclk));
	jxor g01064(.dina(w_n1121_0[0]),.dinb(w_n290_33[2]),.dout(n1276),.clk(gclk));
	jand g01065(.dina(n1276),.dinb(w_asqrt50_27[2]),.dout(n1277),.clk(gclk));
	jxor g01066(.dina(n1277),.dinb(w_n1128_0[0]),.dout(n1278),.clk(gclk));
	jnot g01067(.din(n1278),.dout(n1279),.clk(gclk));
	jor g01068(.dina(w_n1274_0[0]),.dinb(w_asqrt61_26[1]),.dout(n1280),.clk(gclk));
	jand g01069(.dina(w_n1280_0[1]),.dinb(w_n1279_0[1]),.dout(n1281),.clk(gclk));
	jor g01070(.dina(w_n1281_0[2]),.dinb(w_n1275_0[2]),.dout(n1282),.clk(gclk));
	jand g01071(.dina(n1282),.dinb(w_asqrt62_26[2]),.dout(n1283),.clk(gclk));
	jnot g01072(.din(w_n1133_0[0]),.dout(n1284),.clk(gclk));
	jand g01073(.dina(n1284),.dinb(w_n1131_0[0]),.dout(n1285),.clk(gclk));
	jand g01074(.dina(n1285),.dinb(w_asqrt50_27[1]),.dout(n1286),.clk(gclk));
	jxor g01075(.dina(n1286),.dinb(w_n1141_0[0]),.dout(n1287),.clk(gclk));
	jnot g01076(.din(n1287),.dout(n1288),.clk(gclk));
	jor g01077(.dina(w_n1275_0[1]),.dinb(w_asqrt62_26[1]),.dout(n1289),.clk(gclk));
	jor g01078(.dina(n1289),.dinb(w_n1281_0[1]),.dout(n1290),.clk(gclk));
	jand g01079(.dina(w_n1290_0[1]),.dinb(w_n1288_0[1]),.dout(n1291),.clk(gclk));
	jor g01080(.dina(w_n1291_0[1]),.dinb(w_n1283_0[1]),.dout(n1292),.clk(gclk));
	jxor g01081(.dina(w_n1143_0[0]),.dinb(w_n199_39[2]),.dout(n1293),.clk(gclk));
	jand g01082(.dina(n1293),.dinb(w_asqrt50_27[0]),.dout(n1294),.clk(gclk));
	jxor g01083(.dina(n1294),.dinb(w_n1148_0[0]),.dout(n1295),.clk(gclk));
	jnot g01084(.din(w_n1150_0[0]),.dout(n1296),.clk(gclk));
	jnot g01085(.din(w_n1154_0[0]),.dout(n1297),.clk(gclk));
	jand g01086(.dina(w_asqrt50_26[2]),.dinb(w_n1297_0[1]),.dout(n1298),.clk(gclk));
	jand g01087(.dina(w_n1298_0[1]),.dinb(w_n1296_0[2]),.dout(n1299),.clk(gclk));
	jor g01088(.dina(n1299),.dinb(w_n1161_0[0]),.dout(n1300),.clk(gclk));
	jor g01089(.dina(n1300),.dinb(w_n1295_0[1]),.dout(n1301),.clk(gclk));
	jnot g01090(.din(n1301),.dout(n1302),.clk(gclk));
	jand g01091(.dina(n1302),.dinb(w_n1292_1[2]),.dout(n1303),.clk(gclk));
	jor g01092(.dina(n1303),.dinb(w_asqrt63_14[0]),.dout(n1304),.clk(gclk));
	jnot g01093(.din(w_n1295_0[0]),.dout(n1305),.clk(gclk));
	jor g01094(.dina(w_n1305_0[2]),.dinb(w_n1292_1[1]),.dout(n1306),.clk(gclk));
	jor g01095(.dina(w_n1298_0[0]),.dinb(w_n1296_0[1]),.dout(n1307),.clk(gclk));
	jand g01096(.dina(w_n1297_0[0]),.dinb(w_n1296_0[0]),.dout(n1308),.clk(gclk));
	jor g01097(.dina(n1308),.dinb(w_n194_38[2]),.dout(n1309),.clk(gclk));
	jnot g01098(.din(n1309),.dout(n1310),.clk(gclk));
	jand g01099(.dina(n1310),.dinb(n1307),.dout(n1311),.clk(gclk));
	jnot g01100(.din(w_asqrt50_26[1]),.dout(n1312),.clk(gclk));
	jnot g01101(.din(w_n1311_0[1]),.dout(n1315),.clk(gclk));
	jand g01102(.dina(n1315),.dinb(w_n1306_0[1]),.dout(n1316),.clk(gclk));
	jand g01103(.dina(n1316),.dinb(w_n1304_0[1]),.dout(n1317),.clk(gclk));
	jnot g01104(.din(w_n1317_36[1]),.dout(asqrt_fa_50),.clk(gclk));
	jor g01105(.dina(w_n1317_36[0]),.dinb(w_n1172_1[0]),.dout(n1319),.clk(gclk));
	jnot g01106(.din(w_a96_0[1]),.dout(n1320),.clk(gclk));
	jnot g01107(.din(a[97]),.dout(n1321),.clk(gclk));
	jand g01108(.dina(w_n1172_0[2]),.dinb(w_n1321_0[2]),.dout(n1322),.clk(gclk));
	jand g01109(.dina(n1322),.dinb(w_n1320_1[1]),.dout(n1323),.clk(gclk));
	jnot g01110(.din(n1323),.dout(n1324),.clk(gclk));
	jand g01111(.dina(n1324),.dinb(n1319),.dout(n1325),.clk(gclk));
	jor g01112(.dina(w_n1325_0[2]),.dinb(w_n1312_31[2]),.dout(n1326),.clk(gclk));
	jor g01113(.dina(w_n1317_35[2]),.dinb(w_a98_0[0]),.dout(n1327),.clk(gclk));
	jxor g01114(.dina(w_n1327_0[1]),.dinb(w_n1173_0[0]),.dout(n1328),.clk(gclk));
	jand g01115(.dina(w_n1325_0[1]),.dinb(w_n1312_31[1]),.dout(n1329),.clk(gclk));
	jor g01116(.dina(n1329),.dinb(w_n1328_0[1]),.dout(n1330),.clk(gclk));
	jand g01117(.dina(w_n1330_0[1]),.dinb(w_n1326_0[1]),.dout(n1331),.clk(gclk));
	jor g01118(.dina(n1331),.dinb(w_n1039_34[0]),.dout(n1332),.clk(gclk));
	jand g01119(.dina(w_n1326_0[0]),.dinb(w_n1039_33[2]),.dout(n1333),.clk(gclk));
	jand g01120(.dina(n1333),.dinb(w_n1330_0[0]),.dout(n1334),.clk(gclk));
	jor g01121(.dina(w_n1327_0[0]),.dinb(w_a99_0[0]),.dout(n1335),.clk(gclk));
	jnot g01122(.din(w_n1304_0[0]),.dout(n1336),.clk(gclk));
	jnot g01123(.din(w_n1306_0[0]),.dout(n1337),.clk(gclk));
	jor g01124(.dina(w_n1311_0[0]),.dinb(w_n1312_31[0]),.dout(n1338),.clk(gclk));
	jor g01125(.dina(n1338),.dinb(w_n1337_0[1]),.dout(n1339),.clk(gclk));
	jor g01126(.dina(n1339),.dinb(n1336),.dout(n1340),.clk(gclk));
	jand g01127(.dina(n1340),.dinb(n1335),.dout(n1341),.clk(gclk));
	jxor g01128(.dina(n1341),.dinb(w_n1042_0[1]),.dout(n1342),.clk(gclk));
	jor g01129(.dina(w_n1342_0[1]),.dinb(w_n1334_0[1]),.dout(n1343),.clk(gclk));
	jand g01130(.dina(n1343),.dinb(w_n1332_0[1]),.dout(n1344),.clk(gclk));
	jor g01131(.dina(w_n1344_0[2]),.dinb(w_n1034_32[0]),.dout(n1345),.clk(gclk));
	jand g01132(.dina(w_n1344_0[1]),.dinb(w_n1034_31[2]),.dout(n1346),.clk(gclk));
	jxor g01133(.dina(w_n1176_0[0]),.dinb(w_n1039_33[1]),.dout(n1347),.clk(gclk));
	jor g01134(.dina(n1347),.dinb(w_n1317_35[1]),.dout(n1348),.clk(gclk));
	jxor g01135(.dina(n1348),.dinb(w_n1179_0[0]),.dout(n1349),.clk(gclk));
	jor g01136(.dina(w_n1349_0[1]),.dinb(n1346),.dout(n1350),.clk(gclk));
	jand g01137(.dina(w_n1350_0[1]),.dinb(w_n1345_0[1]),.dout(n1351),.clk(gclk));
	jor g01138(.dina(n1351),.dinb(w_n796_33[2]),.dout(n1352),.clk(gclk));
	jnot g01139(.din(w_n1185_0[0]),.dout(n1353),.clk(gclk));
	jor g01140(.dina(n1353),.dinb(w_n1183_0[0]),.dout(n1354),.clk(gclk));
	jor g01141(.dina(n1354),.dinb(w_n1317_35[0]),.dout(n1355),.clk(gclk));
	jxor g01142(.dina(n1355),.dinb(w_n1194_0[0]),.dout(n1356),.clk(gclk));
	jand g01143(.dina(w_n1345_0[0]),.dinb(w_n796_33[1]),.dout(n1357),.clk(gclk));
	jand g01144(.dina(n1357),.dinb(w_n1350_0[0]),.dout(n1358),.clk(gclk));
	jor g01145(.dina(w_n1358_0[1]),.dinb(w_n1356_0[1]),.dout(n1359),.clk(gclk));
	jand g01146(.dina(w_n1359_0[1]),.dinb(w_n1352_0[1]),.dout(n1360),.clk(gclk));
	jor g01147(.dina(w_n1360_0[2]),.dinb(w_n791_32[0]),.dout(n1361),.clk(gclk));
	jand g01148(.dina(w_n1360_0[1]),.dinb(w_n791_31[2]),.dout(n1362),.clk(gclk));
	jxor g01149(.dina(w_n1196_0[0]),.dinb(w_n796_33[0]),.dout(n1363),.clk(gclk));
	jor g01150(.dina(n1363),.dinb(w_n1317_34[2]),.dout(n1364),.clk(gclk));
	jxor g01151(.dina(n1364),.dinb(w_n1201_0[0]),.dout(n1365),.clk(gclk));
	jnot g01152(.din(w_n1365_0[1]),.dout(n1366),.clk(gclk));
	jor g01153(.dina(n1366),.dinb(n1362),.dout(n1367),.clk(gclk));
	jand g01154(.dina(w_n1367_0[1]),.dinb(w_n1361_0[1]),.dout(n1368),.clk(gclk));
	jor g01155(.dina(n1368),.dinb(w_n595_34[0]),.dout(n1369),.clk(gclk));
	jand g01156(.dina(w_n1361_0[0]),.dinb(w_n595_33[2]),.dout(n1370),.clk(gclk));
	jand g01157(.dina(n1370),.dinb(w_n1367_0[0]),.dout(n1371),.clk(gclk));
	jnot g01158(.din(w_n1205_0[0]),.dout(n1372),.clk(gclk));
	jand g01159(.dina(w_asqrt49_26[1]),.dinb(n1372),.dout(n1373),.clk(gclk));
	jand g01160(.dina(w_n1373_0[1]),.dinb(w_n1212_0[0]),.dout(n1374),.clk(gclk));
	jor g01161(.dina(n1374),.dinb(w_n1210_0[0]),.dout(n1375),.clk(gclk));
	jand g01162(.dina(w_n1373_0[0]),.dinb(w_n1213_0[0]),.dout(n1376),.clk(gclk));
	jnot g01163(.din(n1376),.dout(n1377),.clk(gclk));
	jand g01164(.dina(n1377),.dinb(n1375),.dout(n1378),.clk(gclk));
	jnot g01165(.din(n1378),.dout(n1379),.clk(gclk));
	jor g01166(.dina(w_n1379_0[1]),.dinb(w_n1371_0[1]),.dout(n1380),.clk(gclk));
	jand g01167(.dina(n1380),.dinb(w_n1369_0[1]),.dout(n1381),.clk(gclk));
	jor g01168(.dina(w_n1381_0[2]),.dinb(w_n590_32[1]),.dout(n1382),.clk(gclk));
	jand g01169(.dina(w_n1381_0[1]),.dinb(w_n590_32[0]),.dout(n1383),.clk(gclk));
	jnot g01170(.din(w_n1220_0[0]),.dout(n1384),.clk(gclk));
	jxor g01171(.dina(w_n1214_0[0]),.dinb(w_n595_33[1]),.dout(n1385),.clk(gclk));
	jor g01172(.dina(n1385),.dinb(w_n1317_34[1]),.dout(n1386),.clk(gclk));
	jxor g01173(.dina(n1386),.dinb(n1384),.dout(n1387),.clk(gclk));
	jnot g01174(.din(w_n1387_0[1]),.dout(n1388),.clk(gclk));
	jor g01175(.dina(n1388),.dinb(n1383),.dout(n1389),.clk(gclk));
	jand g01176(.dina(w_n1389_0[1]),.dinb(w_n1382_0[1]),.dout(n1390),.clk(gclk));
	jor g01177(.dina(n1390),.dinb(w_n430_33[2]),.dout(n1391),.clk(gclk));
	jnot g01178(.din(w_n1225_0[0]),.dout(n1392),.clk(gclk));
	jor g01179(.dina(n1392),.dinb(w_n1223_0[0]),.dout(n1393),.clk(gclk));
	jor g01180(.dina(n1393),.dinb(w_n1317_34[0]),.dout(n1394),.clk(gclk));
	jxor g01181(.dina(n1394),.dinb(w_n1234_0[0]),.dout(n1395),.clk(gclk));
	jand g01182(.dina(w_n1382_0[0]),.dinb(w_n430_33[1]),.dout(n1396),.clk(gclk));
	jand g01183(.dina(n1396),.dinb(w_n1389_0[0]),.dout(n1397),.clk(gclk));
	jor g01184(.dina(w_n1397_0[1]),.dinb(w_n1395_0[1]),.dout(n1398),.clk(gclk));
	jand g01185(.dina(w_n1398_0[1]),.dinb(w_n1391_0[1]),.dout(n1399),.clk(gclk));
	jor g01186(.dina(w_n1399_0[2]),.dinb(w_n425_32[1]),.dout(n1400),.clk(gclk));
	jand g01187(.dina(w_n1399_0[1]),.dinb(w_n425_32[0]),.dout(n1401),.clk(gclk));
	jnot g01188(.din(w_n1241_0[0]),.dout(n1402),.clk(gclk));
	jxor g01189(.dina(w_n1236_0[0]),.dinb(w_n430_33[0]),.dout(n1403),.clk(gclk));
	jor g01190(.dina(n1403),.dinb(w_n1317_33[2]),.dout(n1404),.clk(gclk));
	jxor g01191(.dina(n1404),.dinb(n1402),.dout(n1405),.clk(gclk));
	jnot g01192(.din(n1405),.dout(n1406),.clk(gclk));
	jor g01193(.dina(w_n1406_0[1]),.dinb(n1401),.dout(n1407),.clk(gclk));
	jand g01194(.dina(w_n1407_0[1]),.dinb(w_n1400_0[1]),.dout(n1408),.clk(gclk));
	jor g01195(.dina(n1408),.dinb(w_n305_34[0]),.dout(n1409),.clk(gclk));
	jand g01196(.dina(w_n1400_0[0]),.dinb(w_n305_33[2]),.dout(n1410),.clk(gclk));
	jand g01197(.dina(n1410),.dinb(w_n1407_0[0]),.dout(n1411),.clk(gclk));
	jnot g01198(.din(w_n1244_0[0]),.dout(n1412),.clk(gclk));
	jand g01199(.dina(w_asqrt49_26[0]),.dinb(n1412),.dout(n1413),.clk(gclk));
	jand g01200(.dina(w_n1413_0[1]),.dinb(w_n1251_0[0]),.dout(n1414),.clk(gclk));
	jor g01201(.dina(n1414),.dinb(w_n1249_0[0]),.dout(n1415),.clk(gclk));
	jand g01202(.dina(w_n1413_0[0]),.dinb(w_n1252_0[0]),.dout(n1416),.clk(gclk));
	jnot g01203(.din(n1416),.dout(n1417),.clk(gclk));
	jand g01204(.dina(n1417),.dinb(n1415),.dout(n1418),.clk(gclk));
	jnot g01205(.din(n1418),.dout(n1419),.clk(gclk));
	jor g01206(.dina(w_n1419_0[1]),.dinb(w_n1411_0[1]),.dout(n1420),.clk(gclk));
	jand g01207(.dina(n1420),.dinb(w_n1409_0[1]),.dout(n1421),.clk(gclk));
	jor g01208(.dina(w_n1421_0[1]),.dinb(w_n290_33[1]),.dout(n1422),.clk(gclk));
	jxor g01209(.dina(w_n1253_0[0]),.dinb(w_n305_33[1]),.dout(n1423),.clk(gclk));
	jor g01210(.dina(n1423),.dinb(w_n1317_33[1]),.dout(n1424),.clk(gclk));
	jxor g01211(.dina(n1424),.dinb(w_n1258_0[0]),.dout(n1425),.clk(gclk));
	jand g01212(.dina(w_n1421_0[0]),.dinb(w_n290_33[0]),.dout(n1426),.clk(gclk));
	jor g01213(.dina(w_n1426_0[1]),.dinb(w_n1425_0[1]),.dout(n1427),.clk(gclk));
	jand g01214(.dina(w_n1427_0[2]),.dinb(w_n1422_0[2]),.dout(n1428),.clk(gclk));
	jor g01215(.dina(n1428),.dinb(w_n223_33[2]),.dout(n1429),.clk(gclk));
	jnot g01216(.din(w_n1263_0[0]),.dout(n1430),.clk(gclk));
	jor g01217(.dina(n1430),.dinb(w_n1261_0[0]),.dout(n1431),.clk(gclk));
	jor g01218(.dina(n1431),.dinb(w_n1317_33[0]),.dout(n1432),.clk(gclk));
	jxor g01219(.dina(n1432),.dinb(w_n1272_0[0]),.dout(n1433),.clk(gclk));
	jand g01220(.dina(w_n1422_0[1]),.dinb(w_n223_33[1]),.dout(n1434),.clk(gclk));
	jand g01221(.dina(n1434),.dinb(w_n1427_0[1]),.dout(n1435),.clk(gclk));
	jor g01222(.dina(w_n1435_0[1]),.dinb(w_n1433_0[1]),.dout(n1436),.clk(gclk));
	jand g01223(.dina(w_n1436_0[1]),.dinb(w_n1429_0[1]),.dout(n1437),.clk(gclk));
	jor g01224(.dina(w_n1437_0[2]),.dinb(w_n199_39[1]),.dout(n1438),.clk(gclk));
	jand g01225(.dina(w_n1437_0[1]),.dinb(w_n199_39[0]),.dout(n1439),.clk(gclk));
	jnot g01226(.din(w_n1275_0[0]),.dout(n1440),.clk(gclk));
	jand g01227(.dina(w_asqrt49_25[2]),.dinb(n1440),.dout(n1441),.clk(gclk));
	jand g01228(.dina(w_n1441_0[1]),.dinb(w_n1280_0[0]),.dout(n1442),.clk(gclk));
	jor g01229(.dina(n1442),.dinb(w_n1279_0[0]),.dout(n1443),.clk(gclk));
	jand g01230(.dina(w_n1441_0[0]),.dinb(w_n1281_0[0]),.dout(n1444),.clk(gclk));
	jnot g01231(.din(n1444),.dout(n1445),.clk(gclk));
	jand g01232(.dina(n1445),.dinb(n1443),.dout(n1446),.clk(gclk));
	jnot g01233(.din(n1446),.dout(n1447),.clk(gclk));
	jor g01234(.dina(w_n1447_0[1]),.dinb(n1439),.dout(n1448),.clk(gclk));
	jand g01235(.dina(n1448),.dinb(n1438),.dout(n1449),.clk(gclk));
	jnot g01236(.din(w_n1283_0[0]),.dout(n1450),.clk(gclk));
	jand g01237(.dina(w_asqrt49_25[1]),.dinb(n1450),.dout(n1451),.clk(gclk));
	jand g01238(.dina(w_n1451_0[1]),.dinb(w_n1290_0[0]),.dout(n1452),.clk(gclk));
	jor g01239(.dina(n1452),.dinb(w_n1288_0[0]),.dout(n1453),.clk(gclk));
	jand g01240(.dina(w_n1451_0[0]),.dinb(w_n1291_0[0]),.dout(n1454),.clk(gclk));
	jnot g01241(.din(n1454),.dout(n1455),.clk(gclk));
	jand g01242(.dina(n1455),.dinb(n1453),.dout(n1456),.clk(gclk));
	jnot g01243(.din(w_n1456_0[2]),.dout(n1457),.clk(gclk));
	jand g01244(.dina(w_asqrt49_25[0]),.dinb(w_n1305_0[1]),.dout(n1458),.clk(gclk));
	jand g01245(.dina(w_n1458_0[1]),.dinb(w_n1292_1[0]),.dout(n1459),.clk(gclk));
	jor g01246(.dina(n1459),.dinb(w_n1337_0[0]),.dout(n1460),.clk(gclk));
	jor g01247(.dina(n1460),.dinb(w_n1457_0[1]),.dout(n1461),.clk(gclk));
	jor g01248(.dina(n1461),.dinb(w_n1449_0[2]),.dout(n1462),.clk(gclk));
	jand g01249(.dina(n1462),.dinb(w_n194_38[1]),.dout(n1463),.clk(gclk));
	jand g01250(.dina(w_n1457_0[0]),.dinb(w_n1449_0[1]),.dout(n1464),.clk(gclk));
	jor g01251(.dina(w_n1458_0[0]),.dinb(w_n1292_0[2]),.dout(n1465),.clk(gclk));
	jand g01252(.dina(w_n1305_0[0]),.dinb(w_n1292_0[1]),.dout(n1466),.clk(gclk));
	jor g01253(.dina(n1466),.dinb(w_n194_38[0]),.dout(n1467),.clk(gclk));
	jnot g01254(.din(n1467),.dout(n1468),.clk(gclk));
	jand g01255(.dina(n1468),.dinb(n1465),.dout(n1469),.clk(gclk));
	jor g01256(.dina(w_n1469_0[1]),.dinb(w_n1464_0[2]),.dout(n1472),.clk(gclk));
	jor g01257(.dina(n1472),.dinb(w_n1463_0[1]),.dout(asqrt_fa_49),.clk(gclk));
	jand g01258(.dina(w_asqrt48_31),.dinb(w_a96_0[0]),.dout(n1474),.clk(gclk));
	jnot g01259(.din(w_a94_0[1]),.dout(n1475),.clk(gclk));
	jnot g01260(.din(w_a95_0[1]),.dout(n1476),.clk(gclk));
	jand g01261(.dina(w_n1320_1[0]),.dinb(w_n1476_0[1]),.dout(n1477),.clk(gclk));
	jand g01262(.dina(n1477),.dinb(w_n1475_1[1]),.dout(n1478),.clk(gclk));
	jor g01263(.dina(n1478),.dinb(n1474),.dout(n1479),.clk(gclk));
	jand g01264(.dina(w_n1479_0[2]),.dinb(w_asqrt49_24[2]),.dout(n1480),.clk(gclk));
	jand g01265(.dina(w_asqrt48_30[2]),.dinb(w_n1320_0[2]),.dout(n1481),.clk(gclk));
	jxor g01266(.dina(w_n1481_0[1]),.dinb(w_n1321_0[1]),.dout(n1482),.clk(gclk));
	jor g01267(.dina(w_n1479_0[1]),.dinb(w_asqrt49_24[1]),.dout(n1483),.clk(gclk));
	jand g01268(.dina(n1483),.dinb(w_n1482_0[1]),.dout(n1484),.clk(gclk));
	jor g01269(.dina(w_n1484_0[1]),.dinb(w_n1480_0[1]),.dout(n1485),.clk(gclk));
	jand g01270(.dina(n1485),.dinb(w_asqrt50_26[0]),.dout(n1486),.clk(gclk));
	jor g01271(.dina(w_n1480_0[0]),.dinb(w_asqrt50_25[2]),.dout(n1487),.clk(gclk));
	jor g01272(.dina(n1487),.dinb(w_n1484_0[0]),.dout(n1488),.clk(gclk));
	jand g01273(.dina(w_n1481_0[0]),.dinb(w_n1321_0[0]),.dout(n1489),.clk(gclk));
	jnot g01274(.din(w_n1463_0[0]),.dout(n1490),.clk(gclk));
	jnot g01275(.din(w_n1464_0[1]),.dout(n1491),.clk(gclk));
	jnot g01276(.din(w_n1469_0[0]),.dout(n1492),.clk(gclk));
	jand g01277(.dina(n1492),.dinb(w_asqrt49_24[0]),.dout(n1493),.clk(gclk));
	jand g01278(.dina(n1493),.dinb(n1491),.dout(n1494),.clk(gclk));
	jand g01279(.dina(n1494),.dinb(n1490),.dout(n1495),.clk(gclk));
	jor g01280(.dina(n1495),.dinb(n1489),.dout(n1496),.clk(gclk));
	jxor g01281(.dina(n1496),.dinb(w_n1172_0[1]),.dout(n1497),.clk(gclk));
	jand g01282(.dina(w_n1497_0[1]),.dinb(w_n1488_0[1]),.dout(n1498),.clk(gclk));
	jor g01283(.dina(n1498),.dinb(w_n1486_0[1]),.dout(n1499),.clk(gclk));
	jand g01284(.dina(w_n1499_0[2]),.dinb(w_asqrt51_24[1]),.dout(n1500),.clk(gclk));
	jor g01285(.dina(w_n1499_0[1]),.dinb(w_asqrt51_24[0]),.dout(n1501),.clk(gclk));
	jxor g01286(.dina(w_n1325_0[0]),.dinb(w_n1312_30[2]),.dout(n1502),.clk(gclk));
	jand g01287(.dina(n1502),.dinb(w_asqrt48_30[1]),.dout(n1503),.clk(gclk));
	jxor g01288(.dina(n1503),.dinb(w_n1328_0[0]),.dout(n1504),.clk(gclk));
	jnot g01289(.din(w_n1504_0[1]),.dout(n1505),.clk(gclk));
	jand g01290(.dina(n1505),.dinb(n1501),.dout(n1506),.clk(gclk));
	jor g01291(.dina(w_n1506_0[1]),.dinb(w_n1500_0[1]),.dout(n1507),.clk(gclk));
	jand g01292(.dina(n1507),.dinb(w_asqrt52_26[0]),.dout(n1508),.clk(gclk));
	jnot g01293(.din(w_n1334_0[0]),.dout(n1509),.clk(gclk));
	jand g01294(.dina(n1509),.dinb(w_n1332_0[0]),.dout(n1510),.clk(gclk));
	jand g01295(.dina(n1510),.dinb(w_asqrt48_30[0]),.dout(n1511),.clk(gclk));
	jxor g01296(.dina(n1511),.dinb(w_n1342_0[0]),.dout(n1512),.clk(gclk));
	jnot g01297(.din(n1512),.dout(n1513),.clk(gclk));
	jor g01298(.dina(w_n1500_0[0]),.dinb(w_asqrt52_25[2]),.dout(n1514),.clk(gclk));
	jor g01299(.dina(n1514),.dinb(w_n1506_0[0]),.dout(n1515),.clk(gclk));
	jand g01300(.dina(w_n1515_0[1]),.dinb(w_n1513_0[1]),.dout(n1516),.clk(gclk));
	jor g01301(.dina(w_n1516_0[1]),.dinb(w_n1508_0[1]),.dout(n1517),.clk(gclk));
	jand g01302(.dina(w_n1517_0[2]),.dinb(w_asqrt53_24[2]),.dout(n1518),.clk(gclk));
	jor g01303(.dina(w_n1517_0[1]),.dinb(w_asqrt53_24[1]),.dout(n1519),.clk(gclk));
	jnot g01304(.din(w_n1349_0[0]),.dout(n1520),.clk(gclk));
	jxor g01305(.dina(w_n1344_0[0]),.dinb(w_n1034_31[1]),.dout(n1521),.clk(gclk));
	jand g01306(.dina(n1521),.dinb(w_asqrt48_29[2]),.dout(n1522),.clk(gclk));
	jxor g01307(.dina(n1522),.dinb(n1520),.dout(n1523),.clk(gclk));
	jand g01308(.dina(w_n1523_0[1]),.dinb(n1519),.dout(n1524),.clk(gclk));
	jor g01309(.dina(w_n1524_0[1]),.dinb(w_n1518_0[1]),.dout(n1525),.clk(gclk));
	jand g01310(.dina(n1525),.dinb(w_asqrt54_26[0]),.dout(n1526),.clk(gclk));
	jor g01311(.dina(w_n1518_0[0]),.dinb(w_asqrt54_25[2]),.dout(n1527),.clk(gclk));
	jor g01312(.dina(n1527),.dinb(w_n1524_0[0]),.dout(n1528),.clk(gclk));
	jnot g01313(.din(w_n1356_0[0]),.dout(n1529),.clk(gclk));
	jnot g01314(.din(w_n1358_0[0]),.dout(n1530),.clk(gclk));
	jand g01315(.dina(w_asqrt48_29[1]),.dinb(w_n1352_0[0]),.dout(n1531),.clk(gclk));
	jand g01316(.dina(w_n1531_0[1]),.dinb(n1530),.dout(n1532),.clk(gclk));
	jor g01317(.dina(n1532),.dinb(n1529),.dout(n1533),.clk(gclk));
	jnot g01318(.din(w_n1359_0[0]),.dout(n1534),.clk(gclk));
	jand g01319(.dina(w_n1531_0[0]),.dinb(n1534),.dout(n1535),.clk(gclk));
	jnot g01320(.din(n1535),.dout(n1536),.clk(gclk));
	jand g01321(.dina(n1536),.dinb(n1533),.dout(n1537),.clk(gclk));
	jand g01322(.dina(w_n1537_0[1]),.dinb(w_n1528_0[1]),.dout(n1538),.clk(gclk));
	jor g01323(.dina(n1538),.dinb(w_n1526_0[1]),.dout(n1539),.clk(gclk));
	jand g01324(.dina(w_n1539_0[2]),.dinb(w_asqrt55_25[0]),.dout(n1540),.clk(gclk));
	jor g01325(.dina(w_n1539_0[1]),.dinb(w_asqrt55_24[2]),.dout(n1541),.clk(gclk));
	jxor g01326(.dina(w_n1360_0[0]),.dinb(w_n791_31[1]),.dout(n1542),.clk(gclk));
	jand g01327(.dina(n1542),.dinb(w_asqrt48_29[0]),.dout(n1543),.clk(gclk));
	jxor g01328(.dina(n1543),.dinb(w_n1365_0[0]),.dout(n1544),.clk(gclk));
	jand g01329(.dina(w_n1544_0[1]),.dinb(n1541),.dout(n1545),.clk(gclk));
	jor g01330(.dina(w_n1545_0[1]),.dinb(w_n1540_0[1]),.dout(n1546),.clk(gclk));
	jand g01331(.dina(n1546),.dinb(w_asqrt56_26[0]),.dout(n1547),.clk(gclk));
	jnot g01332(.din(w_n1371_0[0]),.dout(n1548),.clk(gclk));
	jand g01333(.dina(n1548),.dinb(w_n1369_0[0]),.dout(n1549),.clk(gclk));
	jand g01334(.dina(n1549),.dinb(w_asqrt48_28[2]),.dout(n1550),.clk(gclk));
	jxor g01335(.dina(n1550),.dinb(w_n1379_0[0]),.dout(n1551),.clk(gclk));
	jnot g01336(.din(n1551),.dout(n1552),.clk(gclk));
	jor g01337(.dina(w_n1540_0[0]),.dinb(w_asqrt56_25[2]),.dout(n1553),.clk(gclk));
	jor g01338(.dina(n1553),.dinb(w_n1545_0[0]),.dout(n1554),.clk(gclk));
	jand g01339(.dina(w_n1554_0[1]),.dinb(w_n1552_0[1]),.dout(n1555),.clk(gclk));
	jor g01340(.dina(w_n1555_0[1]),.dinb(w_n1547_0[1]),.dout(n1556),.clk(gclk));
	jand g01341(.dina(w_n1556_0[2]),.dinb(w_asqrt57_25[1]),.dout(n1557),.clk(gclk));
	jor g01342(.dina(w_n1556_0[1]),.dinb(w_asqrt57_25[0]),.dout(n1558),.clk(gclk));
	jxor g01343(.dina(w_n1381_0[0]),.dinb(w_n590_31[2]),.dout(n1559),.clk(gclk));
	jand g01344(.dina(n1559),.dinb(w_asqrt48_28[1]),.dout(n1560),.clk(gclk));
	jxor g01345(.dina(n1560),.dinb(w_n1387_0[0]),.dout(n1561),.clk(gclk));
	jand g01346(.dina(w_n1561_0[1]),.dinb(n1558),.dout(n1562),.clk(gclk));
	jor g01347(.dina(w_n1562_0[1]),.dinb(w_n1557_0[1]),.dout(n1563),.clk(gclk));
	jand g01348(.dina(n1563),.dinb(w_asqrt58_26[0]),.dout(n1564),.clk(gclk));
	jor g01349(.dina(w_n1557_0[0]),.dinb(w_asqrt58_25[2]),.dout(n1565),.clk(gclk));
	jor g01350(.dina(n1565),.dinb(w_n1562_0[0]),.dout(n1566),.clk(gclk));
	jnot g01351(.din(w_n1395_0[0]),.dout(n1567),.clk(gclk));
	jnot g01352(.din(w_n1397_0[0]),.dout(n1568),.clk(gclk));
	jand g01353(.dina(w_asqrt48_28[0]),.dinb(w_n1391_0[0]),.dout(n1569),.clk(gclk));
	jand g01354(.dina(w_n1569_0[1]),.dinb(n1568),.dout(n1570),.clk(gclk));
	jor g01355(.dina(n1570),.dinb(n1567),.dout(n1571),.clk(gclk));
	jnot g01356(.din(w_n1398_0[0]),.dout(n1572),.clk(gclk));
	jand g01357(.dina(w_n1569_0[0]),.dinb(n1572),.dout(n1573),.clk(gclk));
	jnot g01358(.din(n1573),.dout(n1574),.clk(gclk));
	jand g01359(.dina(n1574),.dinb(n1571),.dout(n1575),.clk(gclk));
	jand g01360(.dina(w_n1575_0[1]),.dinb(w_n1566_0[1]),.dout(n1576),.clk(gclk));
	jor g01361(.dina(n1576),.dinb(w_n1564_0[1]),.dout(n1577),.clk(gclk));
	jand g01362(.dina(w_n1577_0[1]),.dinb(w_asqrt59_25[2]),.dout(n1578),.clk(gclk));
	jxor g01363(.dina(w_n1399_0[0]),.dinb(w_n425_31[2]),.dout(n1579),.clk(gclk));
	jand g01364(.dina(n1579),.dinb(w_asqrt48_27[2]),.dout(n1580),.clk(gclk));
	jxor g01365(.dina(n1580),.dinb(w_n1406_0[0]),.dout(n1581),.clk(gclk));
	jnot g01366(.din(n1581),.dout(n1582),.clk(gclk));
	jor g01367(.dina(w_n1577_0[0]),.dinb(w_asqrt59_25[1]),.dout(n1583),.clk(gclk));
	jand g01368(.dina(w_n1583_0[1]),.dinb(w_n1582_0[1]),.dout(n1584),.clk(gclk));
	jor g01369(.dina(w_n1584_0[2]),.dinb(w_n1578_0[2]),.dout(n1585),.clk(gclk));
	jand g01370(.dina(n1585),.dinb(w_asqrt60_25[2]),.dout(n1586),.clk(gclk));
	jnot g01371(.din(w_n1411_0[0]),.dout(n1587),.clk(gclk));
	jand g01372(.dina(n1587),.dinb(w_n1409_0[0]),.dout(n1588),.clk(gclk));
	jand g01373(.dina(n1588),.dinb(w_asqrt48_27[1]),.dout(n1589),.clk(gclk));
	jxor g01374(.dina(n1589),.dinb(w_n1419_0[0]),.dout(n1590),.clk(gclk));
	jnot g01375(.din(n1590),.dout(n1591),.clk(gclk));
	jor g01376(.dina(w_n1578_0[1]),.dinb(w_asqrt60_25[1]),.dout(n1592),.clk(gclk));
	jor g01377(.dina(n1592),.dinb(w_n1584_0[1]),.dout(n1593),.clk(gclk));
	jand g01378(.dina(w_n1593_0[1]),.dinb(w_n1591_0[1]),.dout(n1594),.clk(gclk));
	jor g01379(.dina(w_n1594_0[1]),.dinb(w_n1586_0[1]),.dout(n1595),.clk(gclk));
	jand g01380(.dina(w_n1595_0[2]),.dinb(w_asqrt61_26[0]),.dout(n1596),.clk(gclk));
	jor g01381(.dina(w_n1595_0[1]),.dinb(w_asqrt61_25[2]),.dout(n1597),.clk(gclk));
	jnot g01382(.din(w_n1425_0[0]),.dout(n1598),.clk(gclk));
	jnot g01383(.din(w_n1426_0[0]),.dout(n1599),.clk(gclk));
	jand g01384(.dina(w_asqrt48_27[0]),.dinb(w_n1422_0[0]),.dout(n1600),.clk(gclk));
	jand g01385(.dina(w_n1600_0[1]),.dinb(n1599),.dout(n1601),.clk(gclk));
	jor g01386(.dina(n1601),.dinb(n1598),.dout(n1602),.clk(gclk));
	jnot g01387(.din(w_n1427_0[0]),.dout(n1603),.clk(gclk));
	jand g01388(.dina(w_n1600_0[0]),.dinb(n1603),.dout(n1604),.clk(gclk));
	jnot g01389(.din(n1604),.dout(n1605),.clk(gclk));
	jand g01390(.dina(n1605),.dinb(n1602),.dout(n1606),.clk(gclk));
	jand g01391(.dina(w_n1606_0[1]),.dinb(n1597),.dout(n1607),.clk(gclk));
	jor g01392(.dina(w_n1607_0[1]),.dinb(w_n1596_0[1]),.dout(n1608),.clk(gclk));
	jand g01393(.dina(n1608),.dinb(w_asqrt62_26[0]),.dout(n1609),.clk(gclk));
	jor g01394(.dina(w_n1596_0[0]),.dinb(w_asqrt62_25[2]),.dout(n1610),.clk(gclk));
	jor g01395(.dina(n1610),.dinb(w_n1607_0[0]),.dout(n1611),.clk(gclk));
	jnot g01396(.din(w_n1433_0[0]),.dout(n1612),.clk(gclk));
	jnot g01397(.din(w_n1435_0[0]),.dout(n1613),.clk(gclk));
	jand g01398(.dina(w_asqrt48_26[2]),.dinb(w_n1429_0[0]),.dout(n1614),.clk(gclk));
	jand g01399(.dina(w_n1614_0[1]),.dinb(n1613),.dout(n1615),.clk(gclk));
	jor g01400(.dina(n1615),.dinb(n1612),.dout(n1616),.clk(gclk));
	jnot g01401(.din(w_n1436_0[0]),.dout(n1617),.clk(gclk));
	jand g01402(.dina(w_n1614_0[0]),.dinb(n1617),.dout(n1618),.clk(gclk));
	jnot g01403(.din(n1618),.dout(n1619),.clk(gclk));
	jand g01404(.dina(n1619),.dinb(n1616),.dout(n1620),.clk(gclk));
	jand g01405(.dina(w_n1620_0[1]),.dinb(w_n1611_0[1]),.dout(n1621),.clk(gclk));
	jor g01406(.dina(n1621),.dinb(w_n1609_0[1]),.dout(n1622),.clk(gclk));
	jxor g01407(.dina(w_n1437_0[0]),.dinb(w_n199_38[2]),.dout(n1623),.clk(gclk));
	jand g01408(.dina(n1623),.dinb(w_asqrt48_26[1]),.dout(n1624),.clk(gclk));
	jxor g01409(.dina(n1624),.dinb(w_n1447_0[0]),.dout(n1625),.clk(gclk));
	jnot g01410(.din(w_n1449_0[0]),.dout(n1626),.clk(gclk));
	jand g01411(.dina(w_asqrt48_26[0]),.dinb(w_n1456_0[1]),.dout(n1627),.clk(gclk));
	jand g01412(.dina(w_n1627_0[1]),.dinb(w_n1626_0[2]),.dout(n1628),.clk(gclk));
	jor g01413(.dina(n1628),.dinb(w_n1464_0[0]),.dout(n1629),.clk(gclk));
	jor g01414(.dina(n1629),.dinb(w_n1625_0[1]),.dout(n1630),.clk(gclk));
	jnot g01415(.din(n1630),.dout(n1631),.clk(gclk));
	jand g01416(.dina(n1631),.dinb(w_n1622_1[2]),.dout(n1632),.clk(gclk));
	jor g01417(.dina(n1632),.dinb(w_asqrt63_13[2]),.dout(n1633),.clk(gclk));
	jnot g01418(.din(w_n1625_0[0]),.dout(n1634),.clk(gclk));
	jor g01419(.dina(w_n1634_0[2]),.dinb(w_n1622_1[1]),.dout(n1635),.clk(gclk));
	jor g01420(.dina(w_n1627_0[0]),.dinb(w_n1626_0[1]),.dout(n1636),.clk(gclk));
	jand g01421(.dina(w_n1456_0[0]),.dinb(w_n1626_0[0]),.dout(n1637),.clk(gclk));
	jor g01422(.dina(n1637),.dinb(w_n194_37[2]),.dout(n1638),.clk(gclk));
	jnot g01423(.din(n1638),.dout(n1639),.clk(gclk));
	jand g01424(.dina(n1639),.dinb(n1636),.dout(n1640),.clk(gclk));
	jnot g01425(.din(w_asqrt48_25[2]),.dout(n1641),.clk(gclk));
	jnot g01426(.din(w_n1640_0[1]),.dout(n1644),.clk(gclk));
	jand g01427(.dina(n1644),.dinb(w_n1635_0[1]),.dout(n1645),.clk(gclk));
	jand g01428(.dina(n1645),.dinb(w_n1633_0[1]),.dout(n1646),.clk(gclk));
	jnot g01429(.din(w_n1646_36[1]),.dout(asqrt_fa_48),.clk(gclk));
	jor g01430(.dina(w_n1646_36[0]),.dinb(w_n1475_1[0]),.dout(n1648),.clk(gclk));
	jnot g01431(.din(w_a92_0[1]),.dout(n1649),.clk(gclk));
	jnot g01432(.din(a[93]),.dout(n1650),.clk(gclk));
	jand g01433(.dina(w_n1475_0[2]),.dinb(w_n1650_0[2]),.dout(n1651),.clk(gclk));
	jand g01434(.dina(n1651),.dinb(w_n1649_1[1]),.dout(n1652),.clk(gclk));
	jnot g01435(.din(n1652),.dout(n1653),.clk(gclk));
	jand g01436(.dina(n1653),.dinb(n1648),.dout(n1654),.clk(gclk));
	jor g01437(.dina(w_n1654_0[2]),.dinb(w_n1641_30[2]),.dout(n1655),.clk(gclk));
	jor g01438(.dina(w_n1646_35[2]),.dinb(w_a94_0[0]),.dout(n1656),.clk(gclk));
	jxor g01439(.dina(w_n1656_0[1]),.dinb(w_n1476_0[0]),.dout(n1657),.clk(gclk));
	jand g01440(.dina(w_n1654_0[1]),.dinb(w_n1641_30[1]),.dout(n1658),.clk(gclk));
	jor g01441(.dina(n1658),.dinb(w_n1657_0[1]),.dout(n1659),.clk(gclk));
	jand g01442(.dina(w_n1659_0[1]),.dinb(w_n1655_0[1]),.dout(n1660),.clk(gclk));
	jor g01443(.dina(n1660),.dinb(w_n1317_32[2]),.dout(n1661),.clk(gclk));
	jand g01444(.dina(w_n1655_0[0]),.dinb(w_n1317_32[1]),.dout(n1662),.clk(gclk));
	jand g01445(.dina(n1662),.dinb(w_n1659_0[0]),.dout(n1663),.clk(gclk));
	jor g01446(.dina(w_n1656_0[0]),.dinb(w_a95_0[0]),.dout(n1664),.clk(gclk));
	jnot g01447(.din(w_n1633_0[0]),.dout(n1665),.clk(gclk));
	jnot g01448(.din(w_n1635_0[0]),.dout(n1666),.clk(gclk));
	jor g01449(.dina(w_n1640_0[0]),.dinb(w_n1641_30[0]),.dout(n1667),.clk(gclk));
	jor g01450(.dina(n1667),.dinb(w_n1666_0[1]),.dout(n1668),.clk(gclk));
	jor g01451(.dina(n1668),.dinb(n1665),.dout(n1669),.clk(gclk));
	jand g01452(.dina(n1669),.dinb(n1664),.dout(n1670),.clk(gclk));
	jxor g01453(.dina(n1670),.dinb(w_n1320_0[1]),.dout(n1671),.clk(gclk));
	jor g01454(.dina(w_n1671_0[1]),.dinb(w_n1663_0[1]),.dout(n1672),.clk(gclk));
	jand g01455(.dina(n1672),.dinb(w_n1661_0[1]),.dout(n1673),.clk(gclk));
	jor g01456(.dina(w_n1673_0[2]),.dinb(w_n1312_30[1]),.dout(n1674),.clk(gclk));
	jand g01457(.dina(w_n1673_0[1]),.dinb(w_n1312_30[0]),.dout(n1675),.clk(gclk));
	jxor g01458(.dina(w_n1479_0[0]),.dinb(w_n1317_32[0]),.dout(n1676),.clk(gclk));
	jor g01459(.dina(n1676),.dinb(w_n1646_35[1]),.dout(n1677),.clk(gclk));
	jxor g01460(.dina(n1677),.dinb(w_n1482_0[0]),.dout(n1678),.clk(gclk));
	jor g01461(.dina(w_n1678_0[1]),.dinb(n1675),.dout(n1679),.clk(gclk));
	jand g01462(.dina(w_n1679_0[1]),.dinb(w_n1674_0[1]),.dout(n1680),.clk(gclk));
	jor g01463(.dina(n1680),.dinb(w_n1039_33[0]),.dout(n1681),.clk(gclk));
	jnot g01464(.din(w_n1488_0[0]),.dout(n1682),.clk(gclk));
	jor g01465(.dina(n1682),.dinb(w_n1486_0[0]),.dout(n1683),.clk(gclk));
	jor g01466(.dina(n1683),.dinb(w_n1646_35[0]),.dout(n1684),.clk(gclk));
	jxor g01467(.dina(n1684),.dinb(w_n1497_0[0]),.dout(n1685),.clk(gclk));
	jand g01468(.dina(w_n1674_0[0]),.dinb(w_n1039_32[2]),.dout(n1686),.clk(gclk));
	jand g01469(.dina(n1686),.dinb(w_n1679_0[0]),.dout(n1687),.clk(gclk));
	jor g01470(.dina(w_n1687_0[1]),.dinb(w_n1685_0[1]),.dout(n1688),.clk(gclk));
	jand g01471(.dina(w_n1688_0[1]),.dinb(w_n1681_0[1]),.dout(n1689),.clk(gclk));
	jor g01472(.dina(w_n1689_0[2]),.dinb(w_n1034_31[0]),.dout(n1690),.clk(gclk));
	jand g01473(.dina(w_n1689_0[1]),.dinb(w_n1034_30[2]),.dout(n1691),.clk(gclk));
	jxor g01474(.dina(w_n1499_0[0]),.dinb(w_n1039_32[1]),.dout(n1692),.clk(gclk));
	jor g01475(.dina(n1692),.dinb(w_n1646_34[2]),.dout(n1693),.clk(gclk));
	jxor g01476(.dina(n1693),.dinb(w_n1504_0[0]),.dout(n1694),.clk(gclk));
	jnot g01477(.din(w_n1694_0[1]),.dout(n1695),.clk(gclk));
	jor g01478(.dina(n1695),.dinb(n1691),.dout(n1696),.clk(gclk));
	jand g01479(.dina(w_n1696_0[1]),.dinb(w_n1690_0[1]),.dout(n1697),.clk(gclk));
	jor g01480(.dina(n1697),.dinb(w_n796_32[2]),.dout(n1698),.clk(gclk));
	jand g01481(.dina(w_n1690_0[0]),.dinb(w_n796_32[1]),.dout(n1699),.clk(gclk));
	jand g01482(.dina(n1699),.dinb(w_n1696_0[0]),.dout(n1700),.clk(gclk));
	jnot g01483(.din(w_n1508_0[0]),.dout(n1701),.clk(gclk));
	jand g01484(.dina(w_asqrt47_25[1]),.dinb(n1701),.dout(n1702),.clk(gclk));
	jand g01485(.dina(w_n1702_0[1]),.dinb(w_n1515_0[0]),.dout(n1703),.clk(gclk));
	jor g01486(.dina(n1703),.dinb(w_n1513_0[0]),.dout(n1704),.clk(gclk));
	jand g01487(.dina(w_n1702_0[0]),.dinb(w_n1516_0[0]),.dout(n1705),.clk(gclk));
	jnot g01488(.din(n1705),.dout(n1706),.clk(gclk));
	jand g01489(.dina(n1706),.dinb(n1704),.dout(n1707),.clk(gclk));
	jnot g01490(.din(n1707),.dout(n1708),.clk(gclk));
	jor g01491(.dina(w_n1708_0[1]),.dinb(w_n1700_0[1]),.dout(n1709),.clk(gclk));
	jand g01492(.dina(n1709),.dinb(w_n1698_0[1]),.dout(n1710),.clk(gclk));
	jor g01493(.dina(w_n1710_0[2]),.dinb(w_n791_31[0]),.dout(n1711),.clk(gclk));
	jand g01494(.dina(w_n1710_0[1]),.dinb(w_n791_30[2]),.dout(n1712),.clk(gclk));
	jnot g01495(.din(w_n1523_0[0]),.dout(n1713),.clk(gclk));
	jxor g01496(.dina(w_n1517_0[0]),.dinb(w_n796_32[0]),.dout(n1714),.clk(gclk));
	jor g01497(.dina(n1714),.dinb(w_n1646_34[1]),.dout(n1715),.clk(gclk));
	jxor g01498(.dina(n1715),.dinb(n1713),.dout(n1716),.clk(gclk));
	jnot g01499(.din(w_n1716_0[1]),.dout(n1717),.clk(gclk));
	jor g01500(.dina(n1717),.dinb(n1712),.dout(n1718),.clk(gclk));
	jand g01501(.dina(w_n1718_0[1]),.dinb(w_n1711_0[1]),.dout(n1719),.clk(gclk));
	jor g01502(.dina(n1719),.dinb(w_n595_33[0]),.dout(n1720),.clk(gclk));
	jnot g01503(.din(w_n1528_0[0]),.dout(n1721),.clk(gclk));
	jor g01504(.dina(n1721),.dinb(w_n1526_0[0]),.dout(n1722),.clk(gclk));
	jor g01505(.dina(n1722),.dinb(w_n1646_34[0]),.dout(n1723),.clk(gclk));
	jxor g01506(.dina(n1723),.dinb(w_n1537_0[0]),.dout(n1724),.clk(gclk));
	jand g01507(.dina(w_n1711_0[0]),.dinb(w_n595_32[2]),.dout(n1725),.clk(gclk));
	jand g01508(.dina(n1725),.dinb(w_n1718_0[0]),.dout(n1726),.clk(gclk));
	jor g01509(.dina(w_n1726_0[1]),.dinb(w_n1724_0[1]),.dout(n1727),.clk(gclk));
	jand g01510(.dina(w_n1727_0[1]),.dinb(w_n1720_0[1]),.dout(n1728),.clk(gclk));
	jor g01511(.dina(w_n1728_0[2]),.dinb(w_n590_31[1]),.dout(n1729),.clk(gclk));
	jand g01512(.dina(w_n1728_0[1]),.dinb(w_n590_31[0]),.dout(n1730),.clk(gclk));
	jnot g01513(.din(w_n1544_0[0]),.dout(n1731),.clk(gclk));
	jxor g01514(.dina(w_n1539_0[0]),.dinb(w_n595_32[1]),.dout(n1732),.clk(gclk));
	jor g01515(.dina(n1732),.dinb(w_n1646_33[2]),.dout(n1733),.clk(gclk));
	jxor g01516(.dina(n1733),.dinb(n1731),.dout(n1734),.clk(gclk));
	jnot g01517(.din(n1734),.dout(n1735),.clk(gclk));
	jor g01518(.dina(w_n1735_0[1]),.dinb(n1730),.dout(n1736),.clk(gclk));
	jand g01519(.dina(w_n1736_0[1]),.dinb(w_n1729_0[1]),.dout(n1737),.clk(gclk));
	jor g01520(.dina(n1737),.dinb(w_n430_32[2]),.dout(n1738),.clk(gclk));
	jand g01521(.dina(w_n1729_0[0]),.dinb(w_n430_32[1]),.dout(n1739),.clk(gclk));
	jand g01522(.dina(n1739),.dinb(w_n1736_0[0]),.dout(n1740),.clk(gclk));
	jnot g01523(.din(w_n1547_0[0]),.dout(n1741),.clk(gclk));
	jand g01524(.dina(w_asqrt47_25[0]),.dinb(n1741),.dout(n1742),.clk(gclk));
	jand g01525(.dina(w_n1742_0[1]),.dinb(w_n1554_0[0]),.dout(n1743),.clk(gclk));
	jor g01526(.dina(n1743),.dinb(w_n1552_0[0]),.dout(n1744),.clk(gclk));
	jand g01527(.dina(w_n1742_0[0]),.dinb(w_n1555_0[0]),.dout(n1745),.clk(gclk));
	jnot g01528(.din(n1745),.dout(n1746),.clk(gclk));
	jand g01529(.dina(n1746),.dinb(n1744),.dout(n1747),.clk(gclk));
	jnot g01530(.din(n1747),.dout(n1748),.clk(gclk));
	jor g01531(.dina(w_n1748_0[1]),.dinb(w_n1740_0[1]),.dout(n1749),.clk(gclk));
	jand g01532(.dina(n1749),.dinb(w_n1738_0[1]),.dout(n1750),.clk(gclk));
	jor g01533(.dina(w_n1750_0[1]),.dinb(w_n425_31[1]),.dout(n1751),.clk(gclk));
	jxor g01534(.dina(w_n1556_0[0]),.dinb(w_n430_32[0]),.dout(n1752),.clk(gclk));
	jor g01535(.dina(n1752),.dinb(w_n1646_33[1]),.dout(n1753),.clk(gclk));
	jxor g01536(.dina(n1753),.dinb(w_n1561_0[0]),.dout(n1754),.clk(gclk));
	jand g01537(.dina(w_n1750_0[0]),.dinb(w_n425_31[0]),.dout(n1755),.clk(gclk));
	jor g01538(.dina(w_n1755_0[1]),.dinb(w_n1754_0[1]),.dout(n1756),.clk(gclk));
	jand g01539(.dina(w_n1756_0[2]),.dinb(w_n1751_0[2]),.dout(n1757),.clk(gclk));
	jor g01540(.dina(n1757),.dinb(w_n305_33[0]),.dout(n1758),.clk(gclk));
	jnot g01541(.din(w_n1566_0[0]),.dout(n1759),.clk(gclk));
	jor g01542(.dina(n1759),.dinb(w_n1564_0[0]),.dout(n1760),.clk(gclk));
	jor g01543(.dina(n1760),.dinb(w_n1646_33[0]),.dout(n1761),.clk(gclk));
	jxor g01544(.dina(n1761),.dinb(w_n1575_0[0]),.dout(n1762),.clk(gclk));
	jand g01545(.dina(w_n1751_0[1]),.dinb(w_n305_32[2]),.dout(n1763),.clk(gclk));
	jand g01546(.dina(n1763),.dinb(w_n1756_0[1]),.dout(n1764),.clk(gclk));
	jor g01547(.dina(w_n1764_0[1]),.dinb(w_n1762_0[1]),.dout(n1765),.clk(gclk));
	jand g01548(.dina(w_n1765_0[1]),.dinb(w_n1758_0[1]),.dout(n1766),.clk(gclk));
	jor g01549(.dina(w_n1766_0[2]),.dinb(w_n290_32[2]),.dout(n1767),.clk(gclk));
	jand g01550(.dina(w_n1766_0[1]),.dinb(w_n290_32[1]),.dout(n1768),.clk(gclk));
	jnot g01551(.din(w_n1578_0[0]),.dout(n1769),.clk(gclk));
	jand g01552(.dina(w_asqrt47_24[2]),.dinb(n1769),.dout(n1770),.clk(gclk));
	jand g01553(.dina(w_n1770_0[1]),.dinb(w_n1583_0[0]),.dout(n1771),.clk(gclk));
	jor g01554(.dina(n1771),.dinb(w_n1582_0[0]),.dout(n1772),.clk(gclk));
	jand g01555(.dina(w_n1770_0[0]),.dinb(w_n1584_0[0]),.dout(n1773),.clk(gclk));
	jnot g01556(.din(n1773),.dout(n1774),.clk(gclk));
	jand g01557(.dina(n1774),.dinb(n1772),.dout(n1775),.clk(gclk));
	jnot g01558(.din(n1775),.dout(n1776),.clk(gclk));
	jor g01559(.dina(w_n1776_0[1]),.dinb(n1768),.dout(n1777),.clk(gclk));
	jand g01560(.dina(w_n1777_0[1]),.dinb(w_n1767_0[1]),.dout(n1778),.clk(gclk));
	jor g01561(.dina(n1778),.dinb(w_n223_33[0]),.dout(n1779),.clk(gclk));
	jand g01562(.dina(w_n1767_0[0]),.dinb(w_n223_32[2]),.dout(n1780),.clk(gclk));
	jand g01563(.dina(n1780),.dinb(w_n1777_0[0]),.dout(n1781),.clk(gclk));
	jnot g01564(.din(w_n1586_0[0]),.dout(n1782),.clk(gclk));
	jand g01565(.dina(w_asqrt47_24[1]),.dinb(n1782),.dout(n1783),.clk(gclk));
	jand g01566(.dina(w_n1783_0[1]),.dinb(w_n1593_0[0]),.dout(n1784),.clk(gclk));
	jor g01567(.dina(n1784),.dinb(w_n1591_0[0]),.dout(n1785),.clk(gclk));
	jand g01568(.dina(w_n1783_0[0]),.dinb(w_n1594_0[0]),.dout(n1786),.clk(gclk));
	jnot g01569(.din(n1786),.dout(n1787),.clk(gclk));
	jand g01570(.dina(n1787),.dinb(n1785),.dout(n1788),.clk(gclk));
	jnot g01571(.din(n1788),.dout(n1789),.clk(gclk));
	jor g01572(.dina(w_n1789_0[1]),.dinb(w_n1781_0[1]),.dout(n1790),.clk(gclk));
	jand g01573(.dina(n1790),.dinb(w_n1779_0[1]),.dout(n1791),.clk(gclk));
	jor g01574(.dina(w_n1791_0[2]),.dinb(w_n199_38[1]),.dout(n1792),.clk(gclk));
	jand g01575(.dina(w_n1791_0[1]),.dinb(w_n199_38[0]),.dout(n1793),.clk(gclk));
	jxor g01576(.dina(w_n1595_0[0]),.dinb(w_n223_32[1]),.dout(n1794),.clk(gclk));
	jor g01577(.dina(n1794),.dinb(w_n1646_32[2]),.dout(n1795),.clk(gclk));
	jxor g01578(.dina(n1795),.dinb(w_n1606_0[0]),.dout(n1796),.clk(gclk));
	jor g01579(.dina(w_n1796_0[1]),.dinb(n1793),.dout(n1797),.clk(gclk));
	jand g01580(.dina(n1797),.dinb(n1792),.dout(n1798),.clk(gclk));
	jnot g01581(.din(w_n1611_0[0]),.dout(n1799),.clk(gclk));
	jor g01582(.dina(n1799),.dinb(w_n1609_0[0]),.dout(n1800),.clk(gclk));
	jor g01583(.dina(n1800),.dinb(w_n1646_32[1]),.dout(n1801),.clk(gclk));
	jxor g01584(.dina(n1801),.dinb(w_n1620_0[0]),.dout(n1802),.clk(gclk));
	jand g01585(.dina(w_asqrt47_24[0]),.dinb(w_n1634_0[1]),.dout(n1803),.clk(gclk));
	jand g01586(.dina(w_n1803_0[1]),.dinb(w_n1622_1[0]),.dout(n1804),.clk(gclk));
	jor g01587(.dina(n1804),.dinb(w_n1666_0[0]),.dout(n1805),.clk(gclk));
	jor g01588(.dina(n1805),.dinb(w_n1802_0[2]),.dout(n1806),.clk(gclk));
	jor g01589(.dina(n1806),.dinb(w_n1798_0[2]),.dout(n1807),.clk(gclk));
	jand g01590(.dina(n1807),.dinb(w_n194_37[1]),.dout(n1808),.clk(gclk));
	jand g01591(.dina(w_n1802_0[1]),.dinb(w_n1798_0[1]),.dout(n1809),.clk(gclk));
	jor g01592(.dina(w_n1803_0[0]),.dinb(w_n1622_0[2]),.dout(n1810),.clk(gclk));
	jand g01593(.dina(w_n1634_0[0]),.dinb(w_n1622_0[1]),.dout(n1811),.clk(gclk));
	jor g01594(.dina(n1811),.dinb(w_n194_37[0]),.dout(n1812),.clk(gclk));
	jnot g01595(.din(n1812),.dout(n1813),.clk(gclk));
	jand g01596(.dina(n1813),.dinb(n1810),.dout(n1814),.clk(gclk));
	jor g01597(.dina(w_n1814_0[1]),.dinb(w_n1809_0[2]),.dout(n1817),.clk(gclk));
	jor g01598(.dina(n1817),.dinb(w_n1808_0[1]),.dout(asqrt_fa_47),.clk(gclk));
	jand g01599(.dina(w_asqrt46_31),.dinb(w_a92_0[0]),.dout(n1819),.clk(gclk));
	jnot g01600(.din(w_a90_0[1]),.dout(n1820),.clk(gclk));
	jnot g01601(.din(w_a91_0[1]),.dout(n1821),.clk(gclk));
	jand g01602(.dina(w_n1649_1[0]),.dinb(w_n1821_0[1]),.dout(n1822),.clk(gclk));
	jand g01603(.dina(n1822),.dinb(w_n1820_1[1]),.dout(n1823),.clk(gclk));
	jor g01604(.dina(n1823),.dinb(n1819),.dout(n1824),.clk(gclk));
	jand g01605(.dina(w_n1824_0[2]),.dinb(w_asqrt47_23[2]),.dout(n1825),.clk(gclk));
	jand g01606(.dina(w_asqrt46_30[2]),.dinb(w_n1649_0[2]),.dout(n1826),.clk(gclk));
	jxor g01607(.dina(w_n1826_0[1]),.dinb(w_n1650_0[1]),.dout(n1827),.clk(gclk));
	jor g01608(.dina(w_n1824_0[1]),.dinb(w_asqrt47_23[1]),.dout(n1828),.clk(gclk));
	jand g01609(.dina(n1828),.dinb(w_n1827_0[1]),.dout(n1829),.clk(gclk));
	jor g01610(.dina(w_n1829_0[1]),.dinb(w_n1825_0[1]),.dout(n1830),.clk(gclk));
	jand g01611(.dina(n1830),.dinb(w_asqrt48_25[1]),.dout(n1831),.clk(gclk));
	jor g01612(.dina(w_n1825_0[0]),.dinb(w_asqrt48_25[0]),.dout(n1832),.clk(gclk));
	jor g01613(.dina(n1832),.dinb(w_n1829_0[0]),.dout(n1833),.clk(gclk));
	jand g01614(.dina(w_n1826_0[0]),.dinb(w_n1650_0[0]),.dout(n1834),.clk(gclk));
	jnot g01615(.din(w_n1808_0[0]),.dout(n1835),.clk(gclk));
	jnot g01616(.din(w_n1809_0[1]),.dout(n1836),.clk(gclk));
	jnot g01617(.din(w_n1814_0[0]),.dout(n1837),.clk(gclk));
	jand g01618(.dina(n1837),.dinb(w_asqrt47_23[0]),.dout(n1838),.clk(gclk));
	jand g01619(.dina(n1838),.dinb(n1836),.dout(n1839),.clk(gclk));
	jand g01620(.dina(n1839),.dinb(n1835),.dout(n1840),.clk(gclk));
	jor g01621(.dina(n1840),.dinb(n1834),.dout(n1841),.clk(gclk));
	jxor g01622(.dina(n1841),.dinb(w_n1475_0[1]),.dout(n1842),.clk(gclk));
	jand g01623(.dina(w_n1842_0[1]),.dinb(w_n1833_0[1]),.dout(n1843),.clk(gclk));
	jor g01624(.dina(n1843),.dinb(w_n1831_0[1]),.dout(n1844),.clk(gclk));
	jand g01625(.dina(w_n1844_0[2]),.dinb(w_asqrt49_23[2]),.dout(n1845),.clk(gclk));
	jor g01626(.dina(w_n1844_0[1]),.dinb(w_asqrt49_23[1]),.dout(n1846),.clk(gclk));
	jxor g01627(.dina(w_n1654_0[0]),.dinb(w_n1641_29[2]),.dout(n1847),.clk(gclk));
	jand g01628(.dina(n1847),.dinb(w_asqrt46_30[1]),.dout(n1848),.clk(gclk));
	jxor g01629(.dina(n1848),.dinb(w_n1657_0[0]),.dout(n1849),.clk(gclk));
	jnot g01630(.din(w_n1849_0[1]),.dout(n1850),.clk(gclk));
	jand g01631(.dina(n1850),.dinb(n1846),.dout(n1851),.clk(gclk));
	jor g01632(.dina(w_n1851_0[1]),.dinb(w_n1845_0[1]),.dout(n1852),.clk(gclk));
	jand g01633(.dina(n1852),.dinb(w_asqrt50_25[1]),.dout(n1853),.clk(gclk));
	jnot g01634(.din(w_n1663_0[0]),.dout(n1854),.clk(gclk));
	jand g01635(.dina(n1854),.dinb(w_n1661_0[0]),.dout(n1855),.clk(gclk));
	jand g01636(.dina(n1855),.dinb(w_asqrt46_30[0]),.dout(n1856),.clk(gclk));
	jxor g01637(.dina(n1856),.dinb(w_n1671_0[0]),.dout(n1857),.clk(gclk));
	jnot g01638(.din(n1857),.dout(n1858),.clk(gclk));
	jor g01639(.dina(w_n1845_0[0]),.dinb(w_asqrt50_25[0]),.dout(n1859),.clk(gclk));
	jor g01640(.dina(n1859),.dinb(w_n1851_0[0]),.dout(n1860),.clk(gclk));
	jand g01641(.dina(w_n1860_0[1]),.dinb(w_n1858_0[1]),.dout(n1861),.clk(gclk));
	jor g01642(.dina(w_n1861_0[1]),.dinb(w_n1853_0[1]),.dout(n1862),.clk(gclk));
	jand g01643(.dina(w_n1862_0[2]),.dinb(w_asqrt51_23[2]),.dout(n1863),.clk(gclk));
	jor g01644(.dina(w_n1862_0[1]),.dinb(w_asqrt51_23[1]),.dout(n1864),.clk(gclk));
	jnot g01645(.din(w_n1678_0[0]),.dout(n1865),.clk(gclk));
	jxor g01646(.dina(w_n1673_0[0]),.dinb(w_n1312_29[2]),.dout(n1866),.clk(gclk));
	jand g01647(.dina(n1866),.dinb(w_asqrt46_29[2]),.dout(n1867),.clk(gclk));
	jxor g01648(.dina(n1867),.dinb(n1865),.dout(n1868),.clk(gclk));
	jand g01649(.dina(w_n1868_0[1]),.dinb(n1864),.dout(n1869),.clk(gclk));
	jor g01650(.dina(w_n1869_0[1]),.dinb(w_n1863_0[1]),.dout(n1870),.clk(gclk));
	jand g01651(.dina(n1870),.dinb(w_asqrt52_25[1]),.dout(n1871),.clk(gclk));
	jor g01652(.dina(w_n1863_0[0]),.dinb(w_asqrt52_25[0]),.dout(n1872),.clk(gclk));
	jor g01653(.dina(n1872),.dinb(w_n1869_0[0]),.dout(n1873),.clk(gclk));
	jnot g01654(.din(w_n1685_0[0]),.dout(n1874),.clk(gclk));
	jnot g01655(.din(w_n1687_0[0]),.dout(n1875),.clk(gclk));
	jand g01656(.dina(w_asqrt46_29[1]),.dinb(w_n1681_0[0]),.dout(n1876),.clk(gclk));
	jand g01657(.dina(w_n1876_0[1]),.dinb(n1875),.dout(n1877),.clk(gclk));
	jor g01658(.dina(n1877),.dinb(n1874),.dout(n1878),.clk(gclk));
	jnot g01659(.din(w_n1688_0[0]),.dout(n1879),.clk(gclk));
	jand g01660(.dina(w_n1876_0[0]),.dinb(n1879),.dout(n1880),.clk(gclk));
	jnot g01661(.din(n1880),.dout(n1881),.clk(gclk));
	jand g01662(.dina(n1881),.dinb(n1878),.dout(n1882),.clk(gclk));
	jand g01663(.dina(w_n1882_0[1]),.dinb(w_n1873_0[1]),.dout(n1883),.clk(gclk));
	jor g01664(.dina(n1883),.dinb(w_n1871_0[1]),.dout(n1884),.clk(gclk));
	jand g01665(.dina(w_n1884_0[2]),.dinb(w_asqrt53_24[0]),.dout(n1885),.clk(gclk));
	jor g01666(.dina(w_n1884_0[1]),.dinb(w_asqrt53_23[2]),.dout(n1886),.clk(gclk));
	jxor g01667(.dina(w_n1689_0[0]),.dinb(w_n1034_30[1]),.dout(n1887),.clk(gclk));
	jand g01668(.dina(n1887),.dinb(w_asqrt46_29[0]),.dout(n1888),.clk(gclk));
	jxor g01669(.dina(n1888),.dinb(w_n1694_0[0]),.dout(n1889),.clk(gclk));
	jand g01670(.dina(w_n1889_0[1]),.dinb(n1886),.dout(n1890),.clk(gclk));
	jor g01671(.dina(w_n1890_0[1]),.dinb(w_n1885_0[1]),.dout(n1891),.clk(gclk));
	jand g01672(.dina(n1891),.dinb(w_asqrt54_25[1]),.dout(n1892),.clk(gclk));
	jnot g01673(.din(w_n1700_0[0]),.dout(n1893),.clk(gclk));
	jand g01674(.dina(n1893),.dinb(w_n1698_0[0]),.dout(n1894),.clk(gclk));
	jand g01675(.dina(n1894),.dinb(w_asqrt46_28[2]),.dout(n1895),.clk(gclk));
	jxor g01676(.dina(n1895),.dinb(w_n1708_0[0]),.dout(n1896),.clk(gclk));
	jnot g01677(.din(n1896),.dout(n1897),.clk(gclk));
	jor g01678(.dina(w_n1885_0[0]),.dinb(w_asqrt54_25[0]),.dout(n1898),.clk(gclk));
	jor g01679(.dina(n1898),.dinb(w_n1890_0[0]),.dout(n1899),.clk(gclk));
	jand g01680(.dina(w_n1899_0[1]),.dinb(w_n1897_0[1]),.dout(n1900),.clk(gclk));
	jor g01681(.dina(w_n1900_0[1]),.dinb(w_n1892_0[1]),.dout(n1901),.clk(gclk));
	jand g01682(.dina(w_n1901_0[2]),.dinb(w_asqrt55_24[1]),.dout(n1902),.clk(gclk));
	jor g01683(.dina(w_n1901_0[1]),.dinb(w_asqrt55_24[0]),.dout(n1903),.clk(gclk));
	jxor g01684(.dina(w_n1710_0[0]),.dinb(w_n791_30[1]),.dout(n1904),.clk(gclk));
	jand g01685(.dina(n1904),.dinb(w_asqrt46_28[1]),.dout(n1905),.clk(gclk));
	jxor g01686(.dina(n1905),.dinb(w_n1716_0[0]),.dout(n1906),.clk(gclk));
	jand g01687(.dina(w_n1906_0[1]),.dinb(n1903),.dout(n1907),.clk(gclk));
	jor g01688(.dina(w_n1907_0[1]),.dinb(w_n1902_0[1]),.dout(n1908),.clk(gclk));
	jand g01689(.dina(n1908),.dinb(w_asqrt56_25[1]),.dout(n1909),.clk(gclk));
	jor g01690(.dina(w_n1902_0[0]),.dinb(w_asqrt56_25[0]),.dout(n1910),.clk(gclk));
	jor g01691(.dina(n1910),.dinb(w_n1907_0[0]),.dout(n1911),.clk(gclk));
	jnot g01692(.din(w_n1724_0[0]),.dout(n1912),.clk(gclk));
	jnot g01693(.din(w_n1726_0[0]),.dout(n1913),.clk(gclk));
	jand g01694(.dina(w_asqrt46_28[0]),.dinb(w_n1720_0[0]),.dout(n1914),.clk(gclk));
	jand g01695(.dina(w_n1914_0[1]),.dinb(n1913),.dout(n1915),.clk(gclk));
	jor g01696(.dina(n1915),.dinb(n1912),.dout(n1916),.clk(gclk));
	jnot g01697(.din(w_n1727_0[0]),.dout(n1917),.clk(gclk));
	jand g01698(.dina(w_n1914_0[0]),.dinb(n1917),.dout(n1918),.clk(gclk));
	jnot g01699(.din(n1918),.dout(n1919),.clk(gclk));
	jand g01700(.dina(n1919),.dinb(n1916),.dout(n1920),.clk(gclk));
	jand g01701(.dina(w_n1920_0[1]),.dinb(w_n1911_0[1]),.dout(n1921),.clk(gclk));
	jor g01702(.dina(n1921),.dinb(w_n1909_0[1]),.dout(n1922),.clk(gclk));
	jand g01703(.dina(w_n1922_0[1]),.dinb(w_asqrt57_24[2]),.dout(n1923),.clk(gclk));
	jxor g01704(.dina(w_n1728_0[0]),.dinb(w_n590_30[2]),.dout(n1924),.clk(gclk));
	jand g01705(.dina(n1924),.dinb(w_asqrt46_27[2]),.dout(n1925),.clk(gclk));
	jxor g01706(.dina(n1925),.dinb(w_n1735_0[0]),.dout(n1926),.clk(gclk));
	jnot g01707(.din(n1926),.dout(n1927),.clk(gclk));
	jor g01708(.dina(w_n1922_0[0]),.dinb(w_asqrt57_24[1]),.dout(n1928),.clk(gclk));
	jand g01709(.dina(w_n1928_0[1]),.dinb(w_n1927_0[1]),.dout(n1929),.clk(gclk));
	jor g01710(.dina(w_n1929_0[2]),.dinb(w_n1923_0[2]),.dout(n1930),.clk(gclk));
	jand g01711(.dina(n1930),.dinb(w_asqrt58_25[1]),.dout(n1931),.clk(gclk));
	jnot g01712(.din(w_n1740_0[0]),.dout(n1932),.clk(gclk));
	jand g01713(.dina(n1932),.dinb(w_n1738_0[0]),.dout(n1933),.clk(gclk));
	jand g01714(.dina(n1933),.dinb(w_asqrt46_27[1]),.dout(n1934),.clk(gclk));
	jxor g01715(.dina(n1934),.dinb(w_n1748_0[0]),.dout(n1935),.clk(gclk));
	jnot g01716(.din(n1935),.dout(n1936),.clk(gclk));
	jor g01717(.dina(w_n1923_0[1]),.dinb(w_asqrt58_25[0]),.dout(n1937),.clk(gclk));
	jor g01718(.dina(n1937),.dinb(w_n1929_0[1]),.dout(n1938),.clk(gclk));
	jand g01719(.dina(w_n1938_0[1]),.dinb(w_n1936_0[1]),.dout(n1939),.clk(gclk));
	jor g01720(.dina(w_n1939_0[1]),.dinb(w_n1931_0[1]),.dout(n1940),.clk(gclk));
	jand g01721(.dina(w_n1940_0[2]),.dinb(w_asqrt59_25[0]),.dout(n1941),.clk(gclk));
	jor g01722(.dina(w_n1940_0[1]),.dinb(w_asqrt59_24[2]),.dout(n1942),.clk(gclk));
	jnot g01723(.din(w_n1754_0[0]),.dout(n1943),.clk(gclk));
	jnot g01724(.din(w_n1755_0[0]),.dout(n1944),.clk(gclk));
	jand g01725(.dina(w_asqrt46_27[0]),.dinb(w_n1751_0[0]),.dout(n1945),.clk(gclk));
	jand g01726(.dina(w_n1945_0[1]),.dinb(n1944),.dout(n1946),.clk(gclk));
	jor g01727(.dina(n1946),.dinb(n1943),.dout(n1947),.clk(gclk));
	jnot g01728(.din(w_n1756_0[0]),.dout(n1948),.clk(gclk));
	jand g01729(.dina(w_n1945_0[0]),.dinb(n1948),.dout(n1949),.clk(gclk));
	jnot g01730(.din(n1949),.dout(n1950),.clk(gclk));
	jand g01731(.dina(n1950),.dinb(n1947),.dout(n1951),.clk(gclk));
	jand g01732(.dina(w_n1951_0[1]),.dinb(n1942),.dout(n1952),.clk(gclk));
	jor g01733(.dina(w_n1952_0[1]),.dinb(w_n1941_0[1]),.dout(n1953),.clk(gclk));
	jand g01734(.dina(n1953),.dinb(w_asqrt60_25[0]),.dout(n1954),.clk(gclk));
	jor g01735(.dina(w_n1941_0[0]),.dinb(w_asqrt60_24[2]),.dout(n1955),.clk(gclk));
	jor g01736(.dina(n1955),.dinb(w_n1952_0[0]),.dout(n1956),.clk(gclk));
	jnot g01737(.din(w_n1762_0[0]),.dout(n1957),.clk(gclk));
	jnot g01738(.din(w_n1764_0[0]),.dout(n1958),.clk(gclk));
	jand g01739(.dina(w_asqrt46_26[2]),.dinb(w_n1758_0[0]),.dout(n1959),.clk(gclk));
	jand g01740(.dina(w_n1959_0[1]),.dinb(n1958),.dout(n1960),.clk(gclk));
	jor g01741(.dina(n1960),.dinb(n1957),.dout(n1961),.clk(gclk));
	jnot g01742(.din(w_n1765_0[0]),.dout(n1962),.clk(gclk));
	jand g01743(.dina(w_n1959_0[0]),.dinb(n1962),.dout(n1963),.clk(gclk));
	jnot g01744(.din(n1963),.dout(n1964),.clk(gclk));
	jand g01745(.dina(n1964),.dinb(n1961),.dout(n1965),.clk(gclk));
	jand g01746(.dina(w_n1965_0[1]),.dinb(w_n1956_0[1]),.dout(n1966),.clk(gclk));
	jor g01747(.dina(n1966),.dinb(w_n1954_0[1]),.dout(n1967),.clk(gclk));
	jand g01748(.dina(w_n1967_0[1]),.dinb(w_asqrt61_25[1]),.dout(n1968),.clk(gclk));
	jxor g01749(.dina(w_n1766_0[0]),.dinb(w_n290_32[0]),.dout(n1969),.clk(gclk));
	jand g01750(.dina(n1969),.dinb(w_asqrt46_26[1]),.dout(n1970),.clk(gclk));
	jxor g01751(.dina(n1970),.dinb(w_n1776_0[0]),.dout(n1971),.clk(gclk));
	jnot g01752(.din(n1971),.dout(n1972),.clk(gclk));
	jor g01753(.dina(w_n1967_0[0]),.dinb(w_asqrt61_25[0]),.dout(n1973),.clk(gclk));
	jand g01754(.dina(w_n1973_0[1]),.dinb(w_n1972_0[1]),.dout(n1974),.clk(gclk));
	jor g01755(.dina(w_n1974_0[2]),.dinb(w_n1968_0[2]),.dout(n1975),.clk(gclk));
	jand g01756(.dina(n1975),.dinb(w_asqrt62_25[1]),.dout(n1976),.clk(gclk));
	jnot g01757(.din(w_n1781_0[0]),.dout(n1977),.clk(gclk));
	jand g01758(.dina(n1977),.dinb(w_n1779_0[0]),.dout(n1978),.clk(gclk));
	jand g01759(.dina(n1978),.dinb(w_asqrt46_26[0]),.dout(n1979),.clk(gclk));
	jxor g01760(.dina(n1979),.dinb(w_n1789_0[0]),.dout(n1980),.clk(gclk));
	jnot g01761(.din(n1980),.dout(n1981),.clk(gclk));
	jor g01762(.dina(w_n1968_0[1]),.dinb(w_asqrt62_25[0]),.dout(n1982),.clk(gclk));
	jor g01763(.dina(n1982),.dinb(w_n1974_0[1]),.dout(n1983),.clk(gclk));
	jand g01764(.dina(w_n1983_0[1]),.dinb(w_n1981_0[1]),.dout(n1984),.clk(gclk));
	jor g01765(.dina(w_n1984_0[1]),.dinb(w_n1976_0[1]),.dout(n1985),.clk(gclk));
	jxor g01766(.dina(w_n1791_0[0]),.dinb(w_n199_37[2]),.dout(n1986),.clk(gclk));
	jand g01767(.dina(n1986),.dinb(w_asqrt46_25[2]),.dout(n1987),.clk(gclk));
	jxor g01768(.dina(n1987),.dinb(w_n1796_0[0]),.dout(n1988),.clk(gclk));
	jnot g01769(.din(w_n1798_0[0]),.dout(n1989),.clk(gclk));
	jnot g01770(.din(w_n1802_0[0]),.dout(n1990),.clk(gclk));
	jand g01771(.dina(w_asqrt46_25[1]),.dinb(w_n1990_0[1]),.dout(n1991),.clk(gclk));
	jand g01772(.dina(w_n1991_0[1]),.dinb(w_n1989_0[2]),.dout(n1992),.clk(gclk));
	jor g01773(.dina(n1992),.dinb(w_n1809_0[0]),.dout(n1993),.clk(gclk));
	jor g01774(.dina(n1993),.dinb(w_n1988_0[1]),.dout(n1994),.clk(gclk));
	jnot g01775(.din(n1994),.dout(n1995),.clk(gclk));
	jand g01776(.dina(n1995),.dinb(w_n1985_1[2]),.dout(n1996),.clk(gclk));
	jor g01777(.dina(n1996),.dinb(w_asqrt63_13[1]),.dout(n1997),.clk(gclk));
	jnot g01778(.din(w_n1988_0[0]),.dout(n1998),.clk(gclk));
	jor g01779(.dina(w_n1998_0[2]),.dinb(w_n1985_1[1]),.dout(n1999),.clk(gclk));
	jor g01780(.dina(w_n1991_0[0]),.dinb(w_n1989_0[1]),.dout(n2000),.clk(gclk));
	jand g01781(.dina(w_n1990_0[0]),.dinb(w_n1989_0[0]),.dout(n2001),.clk(gclk));
	jor g01782(.dina(n2001),.dinb(w_n194_36[2]),.dout(n2002),.clk(gclk));
	jnot g01783(.din(n2002),.dout(n2003),.clk(gclk));
	jand g01784(.dina(n2003),.dinb(n2000),.dout(n2004),.clk(gclk));
	jnot g01785(.din(w_asqrt46_25[0]),.dout(n2005),.clk(gclk));
	jnot g01786(.din(w_n2004_0[1]),.dout(n2008),.clk(gclk));
	jand g01787(.dina(n2008),.dinb(w_n1999_0[1]),.dout(n2009),.clk(gclk));
	jand g01788(.dina(n2009),.dinb(w_n1997_0[1]),.dout(n2010),.clk(gclk));
	jnot g01789(.din(w_n2010_34[2]),.dout(asqrt_fa_46),.clk(gclk));
	jor g01790(.dina(w_n2010_34[1]),.dinb(w_n1820_1[0]),.dout(n2012),.clk(gclk));
	jnot g01791(.din(w_a88_0[1]),.dout(n2013),.clk(gclk));
	jnot g01792(.din(a[89]),.dout(n2014),.clk(gclk));
	jand g01793(.dina(w_n1820_0[2]),.dinb(w_n2014_0[2]),.dout(n2015),.clk(gclk));
	jand g01794(.dina(n2015),.dinb(w_n2013_1[1]),.dout(n2016),.clk(gclk));
	jnot g01795(.din(n2016),.dout(n2017),.clk(gclk));
	jand g01796(.dina(n2017),.dinb(n2012),.dout(n2018),.clk(gclk));
	jor g01797(.dina(w_n2018_0[2]),.dinb(w_n2005_29[1]),.dout(n2019),.clk(gclk));
	jor g01798(.dina(w_n2010_34[0]),.dinb(w_a90_0[0]),.dout(n2020),.clk(gclk));
	jxor g01799(.dina(w_n2020_0[1]),.dinb(w_n1821_0[0]),.dout(n2021),.clk(gclk));
	jand g01800(.dina(w_n2018_0[1]),.dinb(w_n2005_29[0]),.dout(n2022),.clk(gclk));
	jor g01801(.dina(n2022),.dinb(w_n2021_0[1]),.dout(n2023),.clk(gclk));
	jand g01802(.dina(w_n2023_0[1]),.dinb(w_n2019_0[1]),.dout(n2024),.clk(gclk));
	jor g01803(.dina(n2024),.dinb(w_n1646_32[0]),.dout(n2025),.clk(gclk));
	jand g01804(.dina(w_n2019_0[0]),.dinb(w_n1646_31[2]),.dout(n2026),.clk(gclk));
	jand g01805(.dina(n2026),.dinb(w_n2023_0[0]),.dout(n2027),.clk(gclk));
	jor g01806(.dina(w_n2020_0[0]),.dinb(w_a91_0[0]),.dout(n2028),.clk(gclk));
	jnot g01807(.din(w_n1997_0[0]),.dout(n2029),.clk(gclk));
	jnot g01808(.din(w_n1999_0[0]),.dout(n2030),.clk(gclk));
	jor g01809(.dina(w_n2004_0[0]),.dinb(w_n2005_28[2]),.dout(n2031),.clk(gclk));
	jor g01810(.dina(n2031),.dinb(w_n2030_0[1]),.dout(n2032),.clk(gclk));
	jor g01811(.dina(n2032),.dinb(n2029),.dout(n2033),.clk(gclk));
	jand g01812(.dina(n2033),.dinb(n2028),.dout(n2034),.clk(gclk));
	jxor g01813(.dina(n2034),.dinb(w_n1649_0[1]),.dout(n2035),.clk(gclk));
	jor g01814(.dina(w_n2035_0[1]),.dinb(w_n2027_0[1]),.dout(n2036),.clk(gclk));
	jand g01815(.dina(n2036),.dinb(w_n2025_0[1]),.dout(n2037),.clk(gclk));
	jor g01816(.dina(w_n2037_0[2]),.dinb(w_n1641_29[1]),.dout(n2038),.clk(gclk));
	jand g01817(.dina(w_n2037_0[1]),.dinb(w_n1641_29[0]),.dout(n2039),.clk(gclk));
	jxor g01818(.dina(w_n1824_0[0]),.dinb(w_n1646_31[1]),.dout(n2040),.clk(gclk));
	jor g01819(.dina(n2040),.dinb(w_n2010_33[2]),.dout(n2041),.clk(gclk));
	jxor g01820(.dina(n2041),.dinb(w_n1827_0[0]),.dout(n2042),.clk(gclk));
	jor g01821(.dina(w_n2042_0[1]),.dinb(n2039),.dout(n2043),.clk(gclk));
	jand g01822(.dina(w_n2043_0[1]),.dinb(w_n2038_0[1]),.dout(n2044),.clk(gclk));
	jor g01823(.dina(n2044),.dinb(w_n1317_31[2]),.dout(n2045),.clk(gclk));
	jnot g01824(.din(w_n1833_0[0]),.dout(n2046),.clk(gclk));
	jor g01825(.dina(n2046),.dinb(w_n1831_0[0]),.dout(n2047),.clk(gclk));
	jor g01826(.dina(n2047),.dinb(w_n2010_33[1]),.dout(n2048),.clk(gclk));
	jxor g01827(.dina(n2048),.dinb(w_n1842_0[0]),.dout(n2049),.clk(gclk));
	jand g01828(.dina(w_n2038_0[0]),.dinb(w_n1317_31[1]),.dout(n2050),.clk(gclk));
	jand g01829(.dina(n2050),.dinb(w_n2043_0[0]),.dout(n2051),.clk(gclk));
	jor g01830(.dina(w_n2051_0[1]),.dinb(w_n2049_0[1]),.dout(n2052),.clk(gclk));
	jand g01831(.dina(w_n2052_0[1]),.dinb(w_n2045_0[1]),.dout(n2053),.clk(gclk));
	jor g01832(.dina(w_n2053_0[2]),.dinb(w_n1312_29[1]),.dout(n2054),.clk(gclk));
	jand g01833(.dina(w_n2053_0[1]),.dinb(w_n1312_29[0]),.dout(n2055),.clk(gclk));
	jxor g01834(.dina(w_n1844_0[0]),.dinb(w_n1317_31[0]),.dout(n2056),.clk(gclk));
	jor g01835(.dina(n2056),.dinb(w_n2010_33[0]),.dout(n2057),.clk(gclk));
	jxor g01836(.dina(n2057),.dinb(w_n1849_0[0]),.dout(n2058),.clk(gclk));
	jnot g01837(.din(w_n2058_0[1]),.dout(n2059),.clk(gclk));
	jor g01838(.dina(n2059),.dinb(n2055),.dout(n2060),.clk(gclk));
	jand g01839(.dina(w_n2060_0[1]),.dinb(w_n2054_0[1]),.dout(n2061),.clk(gclk));
	jor g01840(.dina(n2061),.dinb(w_n1039_32[0]),.dout(n2062),.clk(gclk));
	jand g01841(.dina(w_n2054_0[0]),.dinb(w_n1039_31[2]),.dout(n2063),.clk(gclk));
	jand g01842(.dina(n2063),.dinb(w_n2060_0[0]),.dout(n2064),.clk(gclk));
	jnot g01843(.din(w_n1853_0[0]),.dout(n2065),.clk(gclk));
	jand g01844(.dina(w_asqrt45_25[1]),.dinb(n2065),.dout(n2066),.clk(gclk));
	jand g01845(.dina(w_n2066_0[1]),.dinb(w_n1860_0[0]),.dout(n2067),.clk(gclk));
	jor g01846(.dina(n2067),.dinb(w_n1858_0[0]),.dout(n2068),.clk(gclk));
	jand g01847(.dina(w_n2066_0[0]),.dinb(w_n1861_0[0]),.dout(n2069),.clk(gclk));
	jnot g01848(.din(n2069),.dout(n2070),.clk(gclk));
	jand g01849(.dina(n2070),.dinb(n2068),.dout(n2071),.clk(gclk));
	jnot g01850(.din(n2071),.dout(n2072),.clk(gclk));
	jor g01851(.dina(w_n2072_0[1]),.dinb(w_n2064_0[1]),.dout(n2073),.clk(gclk));
	jand g01852(.dina(n2073),.dinb(w_n2062_0[1]),.dout(n2074),.clk(gclk));
	jor g01853(.dina(w_n2074_0[2]),.dinb(w_n1034_30[0]),.dout(n2075),.clk(gclk));
	jand g01854(.dina(w_n2074_0[1]),.dinb(w_n1034_29[2]),.dout(n2076),.clk(gclk));
	jnot g01855(.din(w_n1868_0[0]),.dout(n2077),.clk(gclk));
	jxor g01856(.dina(w_n1862_0[0]),.dinb(w_n1039_31[1]),.dout(n2078),.clk(gclk));
	jor g01857(.dina(n2078),.dinb(w_n2010_32[2]),.dout(n2079),.clk(gclk));
	jxor g01858(.dina(n2079),.dinb(n2077),.dout(n2080),.clk(gclk));
	jnot g01859(.din(w_n2080_0[1]),.dout(n2081),.clk(gclk));
	jor g01860(.dina(n2081),.dinb(n2076),.dout(n2082),.clk(gclk));
	jand g01861(.dina(w_n2082_0[1]),.dinb(w_n2075_0[1]),.dout(n2083),.clk(gclk));
	jor g01862(.dina(n2083),.dinb(w_n796_31[2]),.dout(n2084),.clk(gclk));
	jnot g01863(.din(w_n1873_0[0]),.dout(n2085),.clk(gclk));
	jor g01864(.dina(n2085),.dinb(w_n1871_0[0]),.dout(n2086),.clk(gclk));
	jor g01865(.dina(n2086),.dinb(w_n2010_32[1]),.dout(n2087),.clk(gclk));
	jxor g01866(.dina(n2087),.dinb(w_n1882_0[0]),.dout(n2088),.clk(gclk));
	jand g01867(.dina(w_n2075_0[0]),.dinb(w_n796_31[1]),.dout(n2089),.clk(gclk));
	jand g01868(.dina(n2089),.dinb(w_n2082_0[0]),.dout(n2090),.clk(gclk));
	jor g01869(.dina(w_n2090_0[1]),.dinb(w_n2088_0[1]),.dout(n2091),.clk(gclk));
	jand g01870(.dina(w_n2091_0[1]),.dinb(w_n2084_0[1]),.dout(n2092),.clk(gclk));
	jor g01871(.dina(w_n2092_0[2]),.dinb(w_n791_30[0]),.dout(n2093),.clk(gclk));
	jand g01872(.dina(w_n2092_0[1]),.dinb(w_n791_29[2]),.dout(n2094),.clk(gclk));
	jnot g01873(.din(w_n1889_0[0]),.dout(n2095),.clk(gclk));
	jxor g01874(.dina(w_n1884_0[0]),.dinb(w_n796_31[0]),.dout(n2096),.clk(gclk));
	jor g01875(.dina(n2096),.dinb(w_n2010_32[0]),.dout(n2097),.clk(gclk));
	jxor g01876(.dina(n2097),.dinb(n2095),.dout(n2098),.clk(gclk));
	jnot g01877(.din(n2098),.dout(n2099),.clk(gclk));
	jor g01878(.dina(w_n2099_0[1]),.dinb(n2094),.dout(n2100),.clk(gclk));
	jand g01879(.dina(w_n2100_0[1]),.dinb(w_n2093_0[1]),.dout(n2101),.clk(gclk));
	jor g01880(.dina(n2101),.dinb(w_n595_32[0]),.dout(n2102),.clk(gclk));
	jand g01881(.dina(w_n2093_0[0]),.dinb(w_n595_31[2]),.dout(n2103),.clk(gclk));
	jand g01882(.dina(n2103),.dinb(w_n2100_0[0]),.dout(n2104),.clk(gclk));
	jnot g01883(.din(w_n1892_0[0]),.dout(n2105),.clk(gclk));
	jand g01884(.dina(w_asqrt45_25[0]),.dinb(n2105),.dout(n2106),.clk(gclk));
	jand g01885(.dina(w_n2106_0[1]),.dinb(w_n1899_0[0]),.dout(n2107),.clk(gclk));
	jor g01886(.dina(n2107),.dinb(w_n1897_0[0]),.dout(n2108),.clk(gclk));
	jand g01887(.dina(w_n2106_0[0]),.dinb(w_n1900_0[0]),.dout(n2109),.clk(gclk));
	jnot g01888(.din(n2109),.dout(n2110),.clk(gclk));
	jand g01889(.dina(n2110),.dinb(n2108),.dout(n2111),.clk(gclk));
	jnot g01890(.din(n2111),.dout(n2112),.clk(gclk));
	jor g01891(.dina(w_n2112_0[1]),.dinb(w_n2104_0[1]),.dout(n2113),.clk(gclk));
	jand g01892(.dina(n2113),.dinb(w_n2102_0[1]),.dout(n2114),.clk(gclk));
	jor g01893(.dina(w_n2114_0[1]),.dinb(w_n590_30[1]),.dout(n2115),.clk(gclk));
	jxor g01894(.dina(w_n1901_0[0]),.dinb(w_n595_31[1]),.dout(n2116),.clk(gclk));
	jor g01895(.dina(n2116),.dinb(w_n2010_31[2]),.dout(n2117),.clk(gclk));
	jxor g01896(.dina(n2117),.dinb(w_n1906_0[0]),.dout(n2118),.clk(gclk));
	jand g01897(.dina(w_n2114_0[0]),.dinb(w_n590_30[0]),.dout(n2119),.clk(gclk));
	jor g01898(.dina(w_n2119_0[1]),.dinb(w_n2118_0[1]),.dout(n2120),.clk(gclk));
	jand g01899(.dina(w_n2120_0[2]),.dinb(w_n2115_0[2]),.dout(n2121),.clk(gclk));
	jor g01900(.dina(n2121),.dinb(w_n430_31[2]),.dout(n2122),.clk(gclk));
	jnot g01901(.din(w_n1911_0[0]),.dout(n2123),.clk(gclk));
	jor g01902(.dina(n2123),.dinb(w_n1909_0[0]),.dout(n2124),.clk(gclk));
	jor g01903(.dina(n2124),.dinb(w_n2010_31[1]),.dout(n2125),.clk(gclk));
	jxor g01904(.dina(n2125),.dinb(w_n1920_0[0]),.dout(n2126),.clk(gclk));
	jand g01905(.dina(w_n2115_0[1]),.dinb(w_n430_31[1]),.dout(n2127),.clk(gclk));
	jand g01906(.dina(n2127),.dinb(w_n2120_0[1]),.dout(n2128),.clk(gclk));
	jor g01907(.dina(w_n2128_0[1]),.dinb(w_n2126_0[1]),.dout(n2129),.clk(gclk));
	jand g01908(.dina(w_n2129_0[1]),.dinb(w_n2122_0[1]),.dout(n2130),.clk(gclk));
	jor g01909(.dina(w_n2130_0[2]),.dinb(w_n425_30[2]),.dout(n2131),.clk(gclk));
	jand g01910(.dina(w_n2130_0[1]),.dinb(w_n425_30[1]),.dout(n2132),.clk(gclk));
	jnot g01911(.din(w_n1923_0[0]),.dout(n2133),.clk(gclk));
	jand g01912(.dina(w_asqrt45_24[2]),.dinb(n2133),.dout(n2134),.clk(gclk));
	jand g01913(.dina(w_n2134_0[1]),.dinb(w_n1928_0[0]),.dout(n2135),.clk(gclk));
	jor g01914(.dina(n2135),.dinb(w_n1927_0[0]),.dout(n2136),.clk(gclk));
	jand g01915(.dina(w_n2134_0[0]),.dinb(w_n1929_0[0]),.dout(n2137),.clk(gclk));
	jnot g01916(.din(n2137),.dout(n2138),.clk(gclk));
	jand g01917(.dina(n2138),.dinb(n2136),.dout(n2139),.clk(gclk));
	jnot g01918(.din(n2139),.dout(n2140),.clk(gclk));
	jor g01919(.dina(w_n2140_0[1]),.dinb(n2132),.dout(n2141),.clk(gclk));
	jand g01920(.dina(w_n2141_0[1]),.dinb(w_n2131_0[1]),.dout(n2142),.clk(gclk));
	jor g01921(.dina(n2142),.dinb(w_n305_32[1]),.dout(n2143),.clk(gclk));
	jand g01922(.dina(w_n2131_0[0]),.dinb(w_n305_32[0]),.dout(n2144),.clk(gclk));
	jand g01923(.dina(n2144),.dinb(w_n2141_0[0]),.dout(n2145),.clk(gclk));
	jnot g01924(.din(w_n1931_0[0]),.dout(n2146),.clk(gclk));
	jand g01925(.dina(w_asqrt45_24[1]),.dinb(n2146),.dout(n2147),.clk(gclk));
	jand g01926(.dina(w_n2147_0[1]),.dinb(w_n1938_0[0]),.dout(n2148),.clk(gclk));
	jor g01927(.dina(n2148),.dinb(w_n1936_0[0]),.dout(n2149),.clk(gclk));
	jand g01928(.dina(w_n2147_0[0]),.dinb(w_n1939_0[0]),.dout(n2150),.clk(gclk));
	jnot g01929(.din(n2150),.dout(n2151),.clk(gclk));
	jand g01930(.dina(n2151),.dinb(n2149),.dout(n2152),.clk(gclk));
	jnot g01931(.din(n2152),.dout(n2153),.clk(gclk));
	jor g01932(.dina(w_n2153_0[1]),.dinb(w_n2145_0[1]),.dout(n2154),.clk(gclk));
	jand g01933(.dina(n2154),.dinb(w_n2143_0[1]),.dout(n2155),.clk(gclk));
	jor g01934(.dina(w_n2155_0[1]),.dinb(w_n290_31[2]),.dout(n2156),.clk(gclk));
	jxor g01935(.dina(w_n1940_0[0]),.dinb(w_n305_31[2]),.dout(n2157),.clk(gclk));
	jor g01936(.dina(n2157),.dinb(w_n2010_31[0]),.dout(n2158),.clk(gclk));
	jxor g01937(.dina(n2158),.dinb(w_n1951_0[0]),.dout(n2159),.clk(gclk));
	jand g01938(.dina(w_n2155_0[0]),.dinb(w_n290_31[1]),.dout(n2160),.clk(gclk));
	jor g01939(.dina(w_n2160_0[1]),.dinb(w_n2159_0[1]),.dout(n2161),.clk(gclk));
	jand g01940(.dina(w_n2161_0[2]),.dinb(w_n2156_0[2]),.dout(n2162),.clk(gclk));
	jor g01941(.dina(n2162),.dinb(w_n223_32[0]),.dout(n2163),.clk(gclk));
	jnot g01942(.din(w_n1956_0[0]),.dout(n2164),.clk(gclk));
	jor g01943(.dina(n2164),.dinb(w_n1954_0[0]),.dout(n2165),.clk(gclk));
	jor g01944(.dina(n2165),.dinb(w_n2010_30[2]),.dout(n2166),.clk(gclk));
	jxor g01945(.dina(n2166),.dinb(w_n1965_0[0]),.dout(n2167),.clk(gclk));
	jand g01946(.dina(w_n2156_0[1]),.dinb(w_n223_31[2]),.dout(n2168),.clk(gclk));
	jand g01947(.dina(n2168),.dinb(w_n2161_0[1]),.dout(n2169),.clk(gclk));
	jor g01948(.dina(w_n2169_0[1]),.dinb(w_n2167_0[1]),.dout(n2170),.clk(gclk));
	jand g01949(.dina(w_n2170_0[1]),.dinb(w_n2163_0[1]),.dout(n2171),.clk(gclk));
	jor g01950(.dina(w_n2171_0[2]),.dinb(w_n199_37[1]),.dout(n2172),.clk(gclk));
	jand g01951(.dina(w_n2171_0[1]),.dinb(w_n199_37[0]),.dout(n2173),.clk(gclk));
	jnot g01952(.din(w_n1968_0[0]),.dout(n2174),.clk(gclk));
	jand g01953(.dina(w_asqrt45_24[0]),.dinb(n2174),.dout(n2175),.clk(gclk));
	jand g01954(.dina(w_n2175_0[1]),.dinb(w_n1973_0[0]),.dout(n2176),.clk(gclk));
	jor g01955(.dina(n2176),.dinb(w_n1972_0[0]),.dout(n2177),.clk(gclk));
	jand g01956(.dina(w_n2175_0[0]),.dinb(w_n1974_0[0]),.dout(n2178),.clk(gclk));
	jnot g01957(.din(n2178),.dout(n2179),.clk(gclk));
	jand g01958(.dina(n2179),.dinb(n2177),.dout(n2180),.clk(gclk));
	jnot g01959(.din(n2180),.dout(n2181),.clk(gclk));
	jor g01960(.dina(w_n2181_0[1]),.dinb(n2173),.dout(n2182),.clk(gclk));
	jand g01961(.dina(n2182),.dinb(n2172),.dout(n2183),.clk(gclk));
	jnot g01962(.din(w_n1976_0[0]),.dout(n2184),.clk(gclk));
	jand g01963(.dina(w_asqrt45_23[2]),.dinb(n2184),.dout(n2185),.clk(gclk));
	jand g01964(.dina(w_n2185_0[1]),.dinb(w_n1983_0[0]),.dout(n2186),.clk(gclk));
	jor g01965(.dina(n2186),.dinb(w_n1981_0[0]),.dout(n2187),.clk(gclk));
	jand g01966(.dina(w_n2185_0[0]),.dinb(w_n1984_0[0]),.dout(n2188),.clk(gclk));
	jnot g01967(.din(n2188),.dout(n2189),.clk(gclk));
	jand g01968(.dina(n2189),.dinb(n2187),.dout(n2190),.clk(gclk));
	jnot g01969(.din(w_n2190_0[2]),.dout(n2191),.clk(gclk));
	jand g01970(.dina(w_asqrt45_23[1]),.dinb(w_n1998_0[1]),.dout(n2192),.clk(gclk));
	jand g01971(.dina(w_n2192_0[1]),.dinb(w_n1985_1[0]),.dout(n2193),.clk(gclk));
	jor g01972(.dina(n2193),.dinb(w_n2030_0[0]),.dout(n2194),.clk(gclk));
	jor g01973(.dina(n2194),.dinb(w_n2191_0[1]),.dout(n2195),.clk(gclk));
	jor g01974(.dina(n2195),.dinb(w_n2183_0[2]),.dout(n2196),.clk(gclk));
	jand g01975(.dina(n2196),.dinb(w_n194_36[1]),.dout(n2197),.clk(gclk));
	jand g01976(.dina(w_n2191_0[0]),.dinb(w_n2183_0[1]),.dout(n2198),.clk(gclk));
	jor g01977(.dina(w_n2192_0[0]),.dinb(w_n1985_0[2]),.dout(n2199),.clk(gclk));
	jand g01978(.dina(w_n1998_0[0]),.dinb(w_n1985_0[1]),.dout(n2200),.clk(gclk));
	jor g01979(.dina(n2200),.dinb(w_n194_36[0]),.dout(n2201),.clk(gclk));
	jnot g01980(.din(n2201),.dout(n2202),.clk(gclk));
	jand g01981(.dina(n2202),.dinb(n2199),.dout(n2203),.clk(gclk));
	jor g01982(.dina(w_n2203_0[1]),.dinb(w_n2198_0[2]),.dout(n2206),.clk(gclk));
	jor g01983(.dina(n2206),.dinb(w_n2197_0[1]),.dout(asqrt_fa_45),.clk(gclk));
	jand g01984(.dina(w_asqrt44_31),.dinb(w_a88_0[0]),.dout(n2208),.clk(gclk));
	jnot g01985(.din(w_a86_0[1]),.dout(n2209),.clk(gclk));
	jnot g01986(.din(w_a87_0[1]),.dout(n2210),.clk(gclk));
	jand g01987(.dina(w_n2013_1[0]),.dinb(w_n2210_0[1]),.dout(n2211),.clk(gclk));
	jand g01988(.dina(n2211),.dinb(w_n2209_1[1]),.dout(n2212),.clk(gclk));
	jor g01989(.dina(n2212),.dinb(n2208),.dout(n2213),.clk(gclk));
	jand g01990(.dina(w_n2213_0[2]),.dinb(w_asqrt45_23[0]),.dout(n2214),.clk(gclk));
	jand g01991(.dina(w_asqrt44_30[2]),.dinb(w_n2013_0[2]),.dout(n2215),.clk(gclk));
	jxor g01992(.dina(w_n2215_0[1]),.dinb(w_n2014_0[1]),.dout(n2216),.clk(gclk));
	jor g01993(.dina(w_n2213_0[1]),.dinb(w_asqrt45_22[2]),.dout(n2217),.clk(gclk));
	jand g01994(.dina(n2217),.dinb(w_n2216_0[1]),.dout(n2218),.clk(gclk));
	jor g01995(.dina(w_n2218_0[1]),.dinb(w_n2214_0[1]),.dout(n2219),.clk(gclk));
	jand g01996(.dina(n2219),.dinb(w_asqrt46_24[2]),.dout(n2220),.clk(gclk));
	jor g01997(.dina(w_n2214_0[0]),.dinb(w_asqrt46_24[1]),.dout(n2221),.clk(gclk));
	jor g01998(.dina(n2221),.dinb(w_n2218_0[0]),.dout(n2222),.clk(gclk));
	jand g01999(.dina(w_n2215_0[0]),.dinb(w_n2014_0[0]),.dout(n2223),.clk(gclk));
	jnot g02000(.din(w_n2197_0[0]),.dout(n2224),.clk(gclk));
	jnot g02001(.din(w_n2198_0[1]),.dout(n2225),.clk(gclk));
	jnot g02002(.din(w_n2203_0[0]),.dout(n2226),.clk(gclk));
	jand g02003(.dina(n2226),.dinb(w_asqrt45_22[1]),.dout(n2227),.clk(gclk));
	jand g02004(.dina(n2227),.dinb(n2225),.dout(n2228),.clk(gclk));
	jand g02005(.dina(n2228),.dinb(n2224),.dout(n2229),.clk(gclk));
	jor g02006(.dina(n2229),.dinb(n2223),.dout(n2230),.clk(gclk));
	jxor g02007(.dina(n2230),.dinb(w_n1820_0[1]),.dout(n2231),.clk(gclk));
	jand g02008(.dina(w_n2231_0[1]),.dinb(w_n2222_0[1]),.dout(n2232),.clk(gclk));
	jor g02009(.dina(n2232),.dinb(w_n2220_0[1]),.dout(n2233),.clk(gclk));
	jand g02010(.dina(w_n2233_0[2]),.dinb(w_asqrt47_22[2]),.dout(n2234),.clk(gclk));
	jor g02011(.dina(w_n2233_0[1]),.dinb(w_asqrt47_22[1]),.dout(n2235),.clk(gclk));
	jxor g02012(.dina(w_n2018_0[0]),.dinb(w_n2005_28[1]),.dout(n2236),.clk(gclk));
	jand g02013(.dina(n2236),.dinb(w_asqrt44_30[1]),.dout(n2237),.clk(gclk));
	jxor g02014(.dina(n2237),.dinb(w_n2021_0[0]),.dout(n2238),.clk(gclk));
	jnot g02015(.din(w_n2238_0[1]),.dout(n2239),.clk(gclk));
	jand g02016(.dina(n2239),.dinb(n2235),.dout(n2240),.clk(gclk));
	jor g02017(.dina(w_n2240_0[1]),.dinb(w_n2234_0[1]),.dout(n2241),.clk(gclk));
	jand g02018(.dina(n2241),.dinb(w_asqrt48_24[2]),.dout(n2242),.clk(gclk));
	jnot g02019(.din(w_n2027_0[0]),.dout(n2243),.clk(gclk));
	jand g02020(.dina(n2243),.dinb(w_n2025_0[0]),.dout(n2244),.clk(gclk));
	jand g02021(.dina(n2244),.dinb(w_asqrt44_30[0]),.dout(n2245),.clk(gclk));
	jxor g02022(.dina(n2245),.dinb(w_n2035_0[0]),.dout(n2246),.clk(gclk));
	jnot g02023(.din(n2246),.dout(n2247),.clk(gclk));
	jor g02024(.dina(w_n2234_0[0]),.dinb(w_asqrt48_24[1]),.dout(n2248),.clk(gclk));
	jor g02025(.dina(n2248),.dinb(w_n2240_0[0]),.dout(n2249),.clk(gclk));
	jand g02026(.dina(w_n2249_0[1]),.dinb(w_n2247_0[1]),.dout(n2250),.clk(gclk));
	jor g02027(.dina(w_n2250_0[1]),.dinb(w_n2242_0[1]),.dout(n2251),.clk(gclk));
	jand g02028(.dina(w_n2251_0[2]),.dinb(w_asqrt49_23[0]),.dout(n2252),.clk(gclk));
	jor g02029(.dina(w_n2251_0[1]),.dinb(w_asqrt49_22[2]),.dout(n2253),.clk(gclk));
	jnot g02030(.din(w_n2042_0[0]),.dout(n2254),.clk(gclk));
	jxor g02031(.dina(w_n2037_0[0]),.dinb(w_n1641_28[2]),.dout(n2255),.clk(gclk));
	jand g02032(.dina(n2255),.dinb(w_asqrt44_29[2]),.dout(n2256),.clk(gclk));
	jxor g02033(.dina(n2256),.dinb(n2254),.dout(n2257),.clk(gclk));
	jand g02034(.dina(w_n2257_0[1]),.dinb(n2253),.dout(n2258),.clk(gclk));
	jor g02035(.dina(w_n2258_0[1]),.dinb(w_n2252_0[1]),.dout(n2259),.clk(gclk));
	jand g02036(.dina(n2259),.dinb(w_asqrt50_24[2]),.dout(n2260),.clk(gclk));
	jor g02037(.dina(w_n2252_0[0]),.dinb(w_asqrt50_24[1]),.dout(n2261),.clk(gclk));
	jor g02038(.dina(n2261),.dinb(w_n2258_0[0]),.dout(n2262),.clk(gclk));
	jnot g02039(.din(w_n2049_0[0]),.dout(n2263),.clk(gclk));
	jnot g02040(.din(w_n2051_0[0]),.dout(n2264),.clk(gclk));
	jand g02041(.dina(w_asqrt44_29[1]),.dinb(w_n2045_0[0]),.dout(n2265),.clk(gclk));
	jand g02042(.dina(w_n2265_0[1]),.dinb(n2264),.dout(n2266),.clk(gclk));
	jor g02043(.dina(n2266),.dinb(n2263),.dout(n2267),.clk(gclk));
	jnot g02044(.din(w_n2052_0[0]),.dout(n2268),.clk(gclk));
	jand g02045(.dina(w_n2265_0[0]),.dinb(n2268),.dout(n2269),.clk(gclk));
	jnot g02046(.din(n2269),.dout(n2270),.clk(gclk));
	jand g02047(.dina(n2270),.dinb(n2267),.dout(n2271),.clk(gclk));
	jand g02048(.dina(w_n2271_0[1]),.dinb(w_n2262_0[1]),.dout(n2272),.clk(gclk));
	jor g02049(.dina(n2272),.dinb(w_n2260_0[1]),.dout(n2273),.clk(gclk));
	jand g02050(.dina(w_n2273_0[2]),.dinb(w_asqrt51_23[0]),.dout(n2274),.clk(gclk));
	jor g02051(.dina(w_n2273_0[1]),.dinb(w_asqrt51_22[2]),.dout(n2275),.clk(gclk));
	jxor g02052(.dina(w_n2053_0[0]),.dinb(w_n1312_28[2]),.dout(n2276),.clk(gclk));
	jand g02053(.dina(n2276),.dinb(w_asqrt44_29[0]),.dout(n2277),.clk(gclk));
	jxor g02054(.dina(n2277),.dinb(w_n2058_0[0]),.dout(n2278),.clk(gclk));
	jand g02055(.dina(w_n2278_0[1]),.dinb(n2275),.dout(n2279),.clk(gclk));
	jor g02056(.dina(w_n2279_0[1]),.dinb(w_n2274_0[1]),.dout(n2280),.clk(gclk));
	jand g02057(.dina(n2280),.dinb(w_asqrt52_24[2]),.dout(n2281),.clk(gclk));
	jnot g02058(.din(w_n2064_0[0]),.dout(n2282),.clk(gclk));
	jand g02059(.dina(n2282),.dinb(w_n2062_0[0]),.dout(n2283),.clk(gclk));
	jand g02060(.dina(n2283),.dinb(w_asqrt44_28[2]),.dout(n2284),.clk(gclk));
	jxor g02061(.dina(n2284),.dinb(w_n2072_0[0]),.dout(n2285),.clk(gclk));
	jnot g02062(.din(n2285),.dout(n2286),.clk(gclk));
	jor g02063(.dina(w_n2274_0[0]),.dinb(w_asqrt52_24[1]),.dout(n2287),.clk(gclk));
	jor g02064(.dina(n2287),.dinb(w_n2279_0[0]),.dout(n2288),.clk(gclk));
	jand g02065(.dina(w_n2288_0[1]),.dinb(w_n2286_0[1]),.dout(n2289),.clk(gclk));
	jor g02066(.dina(w_n2289_0[1]),.dinb(w_n2281_0[1]),.dout(n2290),.clk(gclk));
	jand g02067(.dina(w_n2290_0[2]),.dinb(w_asqrt53_23[1]),.dout(n2291),.clk(gclk));
	jor g02068(.dina(w_n2290_0[1]),.dinb(w_asqrt53_23[0]),.dout(n2292),.clk(gclk));
	jxor g02069(.dina(w_n2074_0[0]),.dinb(w_n1034_29[1]),.dout(n2293),.clk(gclk));
	jand g02070(.dina(n2293),.dinb(w_asqrt44_28[1]),.dout(n2294),.clk(gclk));
	jxor g02071(.dina(n2294),.dinb(w_n2080_0[0]),.dout(n2295),.clk(gclk));
	jand g02072(.dina(w_n2295_0[1]),.dinb(n2292),.dout(n2296),.clk(gclk));
	jor g02073(.dina(w_n2296_0[1]),.dinb(w_n2291_0[1]),.dout(n2297),.clk(gclk));
	jand g02074(.dina(n2297),.dinb(w_asqrt54_24[2]),.dout(n2298),.clk(gclk));
	jor g02075(.dina(w_n2291_0[0]),.dinb(w_asqrt54_24[1]),.dout(n2299),.clk(gclk));
	jor g02076(.dina(n2299),.dinb(w_n2296_0[0]),.dout(n2300),.clk(gclk));
	jnot g02077(.din(w_n2088_0[0]),.dout(n2301),.clk(gclk));
	jnot g02078(.din(w_n2090_0[0]),.dout(n2302),.clk(gclk));
	jand g02079(.dina(w_asqrt44_28[0]),.dinb(w_n2084_0[0]),.dout(n2303),.clk(gclk));
	jand g02080(.dina(w_n2303_0[1]),.dinb(n2302),.dout(n2304),.clk(gclk));
	jor g02081(.dina(n2304),.dinb(n2301),.dout(n2305),.clk(gclk));
	jnot g02082(.din(w_n2091_0[0]),.dout(n2306),.clk(gclk));
	jand g02083(.dina(w_n2303_0[0]),.dinb(n2306),.dout(n2307),.clk(gclk));
	jnot g02084(.din(n2307),.dout(n2308),.clk(gclk));
	jand g02085(.dina(n2308),.dinb(n2305),.dout(n2309),.clk(gclk));
	jand g02086(.dina(w_n2309_0[1]),.dinb(w_n2300_0[1]),.dout(n2310),.clk(gclk));
	jor g02087(.dina(n2310),.dinb(w_n2298_0[1]),.dout(n2311),.clk(gclk));
	jand g02088(.dina(w_n2311_0[1]),.dinb(w_asqrt55_23[2]),.dout(n2312),.clk(gclk));
	jxor g02089(.dina(w_n2092_0[0]),.dinb(w_n791_29[1]),.dout(n2313),.clk(gclk));
	jand g02090(.dina(n2313),.dinb(w_asqrt44_27[2]),.dout(n2314),.clk(gclk));
	jxor g02091(.dina(n2314),.dinb(w_n2099_0[0]),.dout(n2315),.clk(gclk));
	jnot g02092(.din(n2315),.dout(n2316),.clk(gclk));
	jor g02093(.dina(w_n2311_0[0]),.dinb(w_asqrt55_23[1]),.dout(n2317),.clk(gclk));
	jand g02094(.dina(w_n2317_0[1]),.dinb(w_n2316_0[1]),.dout(n2318),.clk(gclk));
	jor g02095(.dina(w_n2318_0[2]),.dinb(w_n2312_0[2]),.dout(n2319),.clk(gclk));
	jand g02096(.dina(n2319),.dinb(w_asqrt56_24[2]),.dout(n2320),.clk(gclk));
	jnot g02097(.din(w_n2104_0[0]),.dout(n2321),.clk(gclk));
	jand g02098(.dina(n2321),.dinb(w_n2102_0[0]),.dout(n2322),.clk(gclk));
	jand g02099(.dina(n2322),.dinb(w_asqrt44_27[1]),.dout(n2323),.clk(gclk));
	jxor g02100(.dina(n2323),.dinb(w_n2112_0[0]),.dout(n2324),.clk(gclk));
	jnot g02101(.din(n2324),.dout(n2325),.clk(gclk));
	jor g02102(.dina(w_n2312_0[1]),.dinb(w_asqrt56_24[1]),.dout(n2326),.clk(gclk));
	jor g02103(.dina(n2326),.dinb(w_n2318_0[1]),.dout(n2327),.clk(gclk));
	jand g02104(.dina(w_n2327_0[1]),.dinb(w_n2325_0[1]),.dout(n2328),.clk(gclk));
	jor g02105(.dina(w_n2328_0[1]),.dinb(w_n2320_0[1]),.dout(n2329),.clk(gclk));
	jand g02106(.dina(w_n2329_0[2]),.dinb(w_asqrt57_24[0]),.dout(n2330),.clk(gclk));
	jor g02107(.dina(w_n2329_0[1]),.dinb(w_asqrt57_23[2]),.dout(n2331),.clk(gclk));
	jnot g02108(.din(w_n2118_0[0]),.dout(n2332),.clk(gclk));
	jnot g02109(.din(w_n2119_0[0]),.dout(n2333),.clk(gclk));
	jand g02110(.dina(w_asqrt44_27[0]),.dinb(w_n2115_0[0]),.dout(n2334),.clk(gclk));
	jand g02111(.dina(w_n2334_0[1]),.dinb(n2333),.dout(n2335),.clk(gclk));
	jor g02112(.dina(n2335),.dinb(n2332),.dout(n2336),.clk(gclk));
	jnot g02113(.din(w_n2120_0[0]),.dout(n2337),.clk(gclk));
	jand g02114(.dina(w_n2334_0[0]),.dinb(n2337),.dout(n2338),.clk(gclk));
	jnot g02115(.din(n2338),.dout(n2339),.clk(gclk));
	jand g02116(.dina(n2339),.dinb(n2336),.dout(n2340),.clk(gclk));
	jand g02117(.dina(w_n2340_0[1]),.dinb(n2331),.dout(n2341),.clk(gclk));
	jor g02118(.dina(w_n2341_0[1]),.dinb(w_n2330_0[1]),.dout(n2342),.clk(gclk));
	jand g02119(.dina(n2342),.dinb(w_asqrt58_24[2]),.dout(n2343),.clk(gclk));
	jor g02120(.dina(w_n2330_0[0]),.dinb(w_asqrt58_24[1]),.dout(n2344),.clk(gclk));
	jor g02121(.dina(n2344),.dinb(w_n2341_0[0]),.dout(n2345),.clk(gclk));
	jnot g02122(.din(w_n2126_0[0]),.dout(n2346),.clk(gclk));
	jnot g02123(.din(w_n2128_0[0]),.dout(n2347),.clk(gclk));
	jand g02124(.dina(w_asqrt44_26[2]),.dinb(w_n2122_0[0]),.dout(n2348),.clk(gclk));
	jand g02125(.dina(w_n2348_0[1]),.dinb(n2347),.dout(n2349),.clk(gclk));
	jor g02126(.dina(n2349),.dinb(n2346),.dout(n2350),.clk(gclk));
	jnot g02127(.din(w_n2129_0[0]),.dout(n2351),.clk(gclk));
	jand g02128(.dina(w_n2348_0[0]),.dinb(n2351),.dout(n2352),.clk(gclk));
	jnot g02129(.din(n2352),.dout(n2353),.clk(gclk));
	jand g02130(.dina(n2353),.dinb(n2350),.dout(n2354),.clk(gclk));
	jand g02131(.dina(w_n2354_0[1]),.dinb(w_n2345_0[1]),.dout(n2355),.clk(gclk));
	jor g02132(.dina(n2355),.dinb(w_n2343_0[1]),.dout(n2356),.clk(gclk));
	jand g02133(.dina(w_n2356_0[1]),.dinb(w_asqrt59_24[1]),.dout(n2357),.clk(gclk));
	jxor g02134(.dina(w_n2130_0[0]),.dinb(w_n425_30[0]),.dout(n2358),.clk(gclk));
	jand g02135(.dina(n2358),.dinb(w_asqrt44_26[1]),.dout(n2359),.clk(gclk));
	jxor g02136(.dina(n2359),.dinb(w_n2140_0[0]),.dout(n2360),.clk(gclk));
	jnot g02137(.din(n2360),.dout(n2361),.clk(gclk));
	jor g02138(.dina(w_n2356_0[0]),.dinb(w_asqrt59_24[0]),.dout(n2362),.clk(gclk));
	jand g02139(.dina(w_n2362_0[1]),.dinb(w_n2361_0[1]),.dout(n2363),.clk(gclk));
	jor g02140(.dina(w_n2363_0[2]),.dinb(w_n2357_0[2]),.dout(n2364),.clk(gclk));
	jand g02141(.dina(n2364),.dinb(w_asqrt60_24[1]),.dout(n2365),.clk(gclk));
	jnot g02142(.din(w_n2145_0[0]),.dout(n2366),.clk(gclk));
	jand g02143(.dina(n2366),.dinb(w_n2143_0[0]),.dout(n2367),.clk(gclk));
	jand g02144(.dina(n2367),.dinb(w_asqrt44_26[0]),.dout(n2368),.clk(gclk));
	jxor g02145(.dina(n2368),.dinb(w_n2153_0[0]),.dout(n2369),.clk(gclk));
	jnot g02146(.din(n2369),.dout(n2370),.clk(gclk));
	jor g02147(.dina(w_n2357_0[1]),.dinb(w_asqrt60_24[0]),.dout(n2371),.clk(gclk));
	jor g02148(.dina(n2371),.dinb(w_n2363_0[1]),.dout(n2372),.clk(gclk));
	jand g02149(.dina(w_n2372_0[1]),.dinb(w_n2370_0[1]),.dout(n2373),.clk(gclk));
	jor g02150(.dina(w_n2373_0[1]),.dinb(w_n2365_0[1]),.dout(n2374),.clk(gclk));
	jand g02151(.dina(w_n2374_0[2]),.dinb(w_asqrt61_24[2]),.dout(n2375),.clk(gclk));
	jor g02152(.dina(w_n2374_0[1]),.dinb(w_asqrt61_24[1]),.dout(n2376),.clk(gclk));
	jnot g02153(.din(w_n2159_0[0]),.dout(n2377),.clk(gclk));
	jnot g02154(.din(w_n2160_0[0]),.dout(n2378),.clk(gclk));
	jand g02155(.dina(w_asqrt44_25[2]),.dinb(w_n2156_0[0]),.dout(n2379),.clk(gclk));
	jand g02156(.dina(w_n2379_0[1]),.dinb(n2378),.dout(n2380),.clk(gclk));
	jor g02157(.dina(n2380),.dinb(n2377),.dout(n2381),.clk(gclk));
	jnot g02158(.din(w_n2161_0[0]),.dout(n2382),.clk(gclk));
	jand g02159(.dina(w_n2379_0[0]),.dinb(n2382),.dout(n2383),.clk(gclk));
	jnot g02160(.din(n2383),.dout(n2384),.clk(gclk));
	jand g02161(.dina(n2384),.dinb(n2381),.dout(n2385),.clk(gclk));
	jand g02162(.dina(w_n2385_0[1]),.dinb(n2376),.dout(n2386),.clk(gclk));
	jor g02163(.dina(w_n2386_0[1]),.dinb(w_n2375_0[1]),.dout(n2387),.clk(gclk));
	jand g02164(.dina(n2387),.dinb(w_asqrt62_24[2]),.dout(n2388),.clk(gclk));
	jor g02165(.dina(w_n2375_0[0]),.dinb(w_asqrt62_24[1]),.dout(n2389),.clk(gclk));
	jor g02166(.dina(n2389),.dinb(w_n2386_0[0]),.dout(n2390),.clk(gclk));
	jnot g02167(.din(w_n2167_0[0]),.dout(n2391),.clk(gclk));
	jnot g02168(.din(w_n2169_0[0]),.dout(n2392),.clk(gclk));
	jand g02169(.dina(w_asqrt44_25[1]),.dinb(w_n2163_0[0]),.dout(n2393),.clk(gclk));
	jand g02170(.dina(w_n2393_0[1]),.dinb(n2392),.dout(n2394),.clk(gclk));
	jor g02171(.dina(n2394),.dinb(n2391),.dout(n2395),.clk(gclk));
	jnot g02172(.din(w_n2170_0[0]),.dout(n2396),.clk(gclk));
	jand g02173(.dina(w_n2393_0[0]),.dinb(n2396),.dout(n2397),.clk(gclk));
	jnot g02174(.din(n2397),.dout(n2398),.clk(gclk));
	jand g02175(.dina(n2398),.dinb(n2395),.dout(n2399),.clk(gclk));
	jand g02176(.dina(w_n2399_0[1]),.dinb(w_n2390_0[1]),.dout(n2400),.clk(gclk));
	jor g02177(.dina(n2400),.dinb(w_n2388_0[1]),.dout(n2401),.clk(gclk));
	jxor g02178(.dina(w_n2171_0[0]),.dinb(w_n199_36[2]),.dout(n2402),.clk(gclk));
	jand g02179(.dina(n2402),.dinb(w_asqrt44_25[0]),.dout(n2403),.clk(gclk));
	jxor g02180(.dina(n2403),.dinb(w_n2181_0[0]),.dout(n2404),.clk(gclk));
	jnot g02181(.din(w_n2183_0[0]),.dout(n2405),.clk(gclk));
	jand g02182(.dina(w_asqrt44_24[2]),.dinb(w_n2190_0[1]),.dout(n2406),.clk(gclk));
	jand g02183(.dina(w_n2406_0[1]),.dinb(w_n2405_0[2]),.dout(n2407),.clk(gclk));
	jor g02184(.dina(n2407),.dinb(w_n2198_0[0]),.dout(n2408),.clk(gclk));
	jor g02185(.dina(n2408),.dinb(w_n2404_0[1]),.dout(n2409),.clk(gclk));
	jnot g02186(.din(n2409),.dout(n2410),.clk(gclk));
	jand g02187(.dina(n2410),.dinb(w_n2401_1[2]),.dout(n2411),.clk(gclk));
	jor g02188(.dina(n2411),.dinb(w_asqrt63_13[0]),.dout(n2412),.clk(gclk));
	jnot g02189(.din(w_n2404_0[0]),.dout(n2413),.clk(gclk));
	jor g02190(.dina(w_n2413_0[2]),.dinb(w_n2401_1[1]),.dout(n2414),.clk(gclk));
	jor g02191(.dina(w_n2406_0[0]),.dinb(w_n2405_0[1]),.dout(n2415),.clk(gclk));
	jand g02192(.dina(w_n2190_0[0]),.dinb(w_n2405_0[0]),.dout(n2416),.clk(gclk));
	jor g02193(.dina(n2416),.dinb(w_n194_35[2]),.dout(n2417),.clk(gclk));
	jnot g02194(.din(n2417),.dout(n2418),.clk(gclk));
	jand g02195(.dina(n2418),.dinb(n2415),.dout(n2419),.clk(gclk));
	jnot g02196(.din(w_asqrt44_24[1]),.dout(n2420),.clk(gclk));
	jnot g02197(.din(w_n2419_0[1]),.dout(n2423),.clk(gclk));
	jand g02198(.dina(n2423),.dinb(w_n2414_0[1]),.dout(n2424),.clk(gclk));
	jand g02199(.dina(n2424),.dinb(w_n2412_0[1]),.dout(n2425),.clk(gclk));
	jnot g02200(.din(w_n2425_34[2]),.dout(asqrt_fa_44),.clk(gclk));
	jor g02201(.dina(w_n2425_34[1]),.dinb(w_n2209_1[0]),.dout(n2427),.clk(gclk));
	jnot g02202(.din(w_a84_0[1]),.dout(n2428),.clk(gclk));
	jnot g02203(.din(a[85]),.dout(n2429),.clk(gclk));
	jand g02204(.dina(w_n2209_0[2]),.dinb(w_n2429_0[2]),.dout(n2430),.clk(gclk));
	jand g02205(.dina(n2430),.dinb(w_n2428_1[1]),.dout(n2431),.clk(gclk));
	jnot g02206(.din(n2431),.dout(n2432),.clk(gclk));
	jand g02207(.dina(n2432),.dinb(n2427),.dout(n2433),.clk(gclk));
	jor g02208(.dina(w_n2433_0[2]),.dinb(w_n2420_28[1]),.dout(n2434),.clk(gclk));
	jor g02209(.dina(w_n2425_34[0]),.dinb(w_a86_0[0]),.dout(n2435),.clk(gclk));
	jxor g02210(.dina(w_n2435_0[1]),.dinb(w_n2210_0[0]),.dout(n2436),.clk(gclk));
	jand g02211(.dina(w_n2433_0[1]),.dinb(w_n2420_28[0]),.dout(n2437),.clk(gclk));
	jor g02212(.dina(n2437),.dinb(w_n2436_0[1]),.dout(n2438),.clk(gclk));
	jand g02213(.dina(w_n2438_0[1]),.dinb(w_n2434_0[1]),.dout(n2439),.clk(gclk));
	jor g02214(.dina(n2439),.dinb(w_n2010_30[1]),.dout(n2440),.clk(gclk));
	jand g02215(.dina(w_n2434_0[0]),.dinb(w_n2010_30[0]),.dout(n2441),.clk(gclk));
	jand g02216(.dina(n2441),.dinb(w_n2438_0[0]),.dout(n2442),.clk(gclk));
	jor g02217(.dina(w_n2435_0[0]),.dinb(w_a87_0[0]),.dout(n2443),.clk(gclk));
	jnot g02218(.din(w_n2412_0[0]),.dout(n2444),.clk(gclk));
	jnot g02219(.din(w_n2414_0[0]),.dout(n2445),.clk(gclk));
	jor g02220(.dina(w_n2419_0[0]),.dinb(w_n2420_27[2]),.dout(n2446),.clk(gclk));
	jor g02221(.dina(n2446),.dinb(w_n2445_0[1]),.dout(n2447),.clk(gclk));
	jor g02222(.dina(n2447),.dinb(n2444),.dout(n2448),.clk(gclk));
	jand g02223(.dina(n2448),.dinb(n2443),.dout(n2449),.clk(gclk));
	jxor g02224(.dina(n2449),.dinb(w_n2013_0[1]),.dout(n2450),.clk(gclk));
	jor g02225(.dina(w_n2450_0[1]),.dinb(w_n2442_0[1]),.dout(n2451),.clk(gclk));
	jand g02226(.dina(n2451),.dinb(w_n2440_0[1]),.dout(n2452),.clk(gclk));
	jor g02227(.dina(w_n2452_0[2]),.dinb(w_n2005_28[0]),.dout(n2453),.clk(gclk));
	jand g02228(.dina(w_n2452_0[1]),.dinb(w_n2005_27[2]),.dout(n2454),.clk(gclk));
	jxor g02229(.dina(w_n2213_0[0]),.dinb(w_n2010_29[2]),.dout(n2455),.clk(gclk));
	jor g02230(.dina(n2455),.dinb(w_n2425_33[2]),.dout(n2456),.clk(gclk));
	jxor g02231(.dina(n2456),.dinb(w_n2216_0[0]),.dout(n2457),.clk(gclk));
	jor g02232(.dina(w_n2457_0[1]),.dinb(n2454),.dout(n2458),.clk(gclk));
	jand g02233(.dina(w_n2458_0[1]),.dinb(w_n2453_0[1]),.dout(n2459),.clk(gclk));
	jor g02234(.dina(n2459),.dinb(w_n1646_31[0]),.dout(n2460),.clk(gclk));
	jnot g02235(.din(w_n2222_0[0]),.dout(n2461),.clk(gclk));
	jor g02236(.dina(n2461),.dinb(w_n2220_0[0]),.dout(n2462),.clk(gclk));
	jor g02237(.dina(n2462),.dinb(w_n2425_33[1]),.dout(n2463),.clk(gclk));
	jxor g02238(.dina(n2463),.dinb(w_n2231_0[0]),.dout(n2464),.clk(gclk));
	jand g02239(.dina(w_n2453_0[0]),.dinb(w_n1646_30[2]),.dout(n2465),.clk(gclk));
	jand g02240(.dina(n2465),.dinb(w_n2458_0[0]),.dout(n2466),.clk(gclk));
	jor g02241(.dina(w_n2466_0[1]),.dinb(w_n2464_0[1]),.dout(n2467),.clk(gclk));
	jand g02242(.dina(w_n2467_0[1]),.dinb(w_n2460_0[1]),.dout(n2468),.clk(gclk));
	jor g02243(.dina(w_n2468_0[2]),.dinb(w_n1641_28[1]),.dout(n2469),.clk(gclk));
	jand g02244(.dina(w_n2468_0[1]),.dinb(w_n1641_28[0]),.dout(n2470),.clk(gclk));
	jxor g02245(.dina(w_n2233_0[0]),.dinb(w_n1646_30[1]),.dout(n2471),.clk(gclk));
	jor g02246(.dina(n2471),.dinb(w_n2425_33[0]),.dout(n2472),.clk(gclk));
	jxor g02247(.dina(n2472),.dinb(w_n2238_0[0]),.dout(n2473),.clk(gclk));
	jnot g02248(.din(w_n2473_0[1]),.dout(n2474),.clk(gclk));
	jor g02249(.dina(n2474),.dinb(n2470),.dout(n2475),.clk(gclk));
	jand g02250(.dina(w_n2475_0[1]),.dinb(w_n2469_0[1]),.dout(n2476),.clk(gclk));
	jor g02251(.dina(n2476),.dinb(w_n1317_30[2]),.dout(n2477),.clk(gclk));
	jand g02252(.dina(w_n2469_0[0]),.dinb(w_n1317_30[1]),.dout(n2478),.clk(gclk));
	jand g02253(.dina(n2478),.dinb(w_n2475_0[0]),.dout(n2479),.clk(gclk));
	jnot g02254(.din(w_n2242_0[0]),.dout(n2480),.clk(gclk));
	jand g02255(.dina(w_asqrt43_24[1]),.dinb(n2480),.dout(n2481),.clk(gclk));
	jand g02256(.dina(w_n2481_0[1]),.dinb(w_n2249_0[0]),.dout(n2482),.clk(gclk));
	jor g02257(.dina(n2482),.dinb(w_n2247_0[0]),.dout(n2483),.clk(gclk));
	jand g02258(.dina(w_n2481_0[0]),.dinb(w_n2250_0[0]),.dout(n2484),.clk(gclk));
	jnot g02259(.din(n2484),.dout(n2485),.clk(gclk));
	jand g02260(.dina(n2485),.dinb(n2483),.dout(n2486),.clk(gclk));
	jnot g02261(.din(n2486),.dout(n2487),.clk(gclk));
	jor g02262(.dina(w_n2487_0[1]),.dinb(w_n2479_0[1]),.dout(n2488),.clk(gclk));
	jand g02263(.dina(n2488),.dinb(w_n2477_0[1]),.dout(n2489),.clk(gclk));
	jor g02264(.dina(w_n2489_0[2]),.dinb(w_n1312_28[1]),.dout(n2490),.clk(gclk));
	jand g02265(.dina(w_n2489_0[1]),.dinb(w_n1312_28[0]),.dout(n2491),.clk(gclk));
	jnot g02266(.din(w_n2257_0[0]),.dout(n2492),.clk(gclk));
	jxor g02267(.dina(w_n2251_0[0]),.dinb(w_n1317_30[0]),.dout(n2493),.clk(gclk));
	jor g02268(.dina(n2493),.dinb(w_n2425_32[2]),.dout(n2494),.clk(gclk));
	jxor g02269(.dina(n2494),.dinb(n2492),.dout(n2495),.clk(gclk));
	jnot g02270(.din(w_n2495_0[1]),.dout(n2496),.clk(gclk));
	jor g02271(.dina(n2496),.dinb(n2491),.dout(n2497),.clk(gclk));
	jand g02272(.dina(w_n2497_0[1]),.dinb(w_n2490_0[1]),.dout(n2498),.clk(gclk));
	jor g02273(.dina(n2498),.dinb(w_n1039_31[0]),.dout(n2499),.clk(gclk));
	jnot g02274(.din(w_n2262_0[0]),.dout(n2500),.clk(gclk));
	jor g02275(.dina(n2500),.dinb(w_n2260_0[0]),.dout(n2501),.clk(gclk));
	jor g02276(.dina(n2501),.dinb(w_n2425_32[1]),.dout(n2502),.clk(gclk));
	jxor g02277(.dina(n2502),.dinb(w_n2271_0[0]),.dout(n2503),.clk(gclk));
	jand g02278(.dina(w_n2490_0[0]),.dinb(w_n1039_30[2]),.dout(n2504),.clk(gclk));
	jand g02279(.dina(n2504),.dinb(w_n2497_0[0]),.dout(n2505),.clk(gclk));
	jor g02280(.dina(w_n2505_0[1]),.dinb(w_n2503_0[1]),.dout(n2506),.clk(gclk));
	jand g02281(.dina(w_n2506_0[1]),.dinb(w_n2499_0[1]),.dout(n2507),.clk(gclk));
	jor g02282(.dina(w_n2507_0[2]),.dinb(w_n1034_29[0]),.dout(n2508),.clk(gclk));
	jand g02283(.dina(w_n2507_0[1]),.dinb(w_n1034_28[2]),.dout(n2509),.clk(gclk));
	jnot g02284(.din(w_n2278_0[0]),.dout(n2510),.clk(gclk));
	jxor g02285(.dina(w_n2273_0[0]),.dinb(w_n1039_30[1]),.dout(n2511),.clk(gclk));
	jor g02286(.dina(n2511),.dinb(w_n2425_32[0]),.dout(n2512),.clk(gclk));
	jxor g02287(.dina(n2512),.dinb(n2510),.dout(n2513),.clk(gclk));
	jnot g02288(.din(n2513),.dout(n2514),.clk(gclk));
	jor g02289(.dina(w_n2514_0[1]),.dinb(n2509),.dout(n2515),.clk(gclk));
	jand g02290(.dina(w_n2515_0[1]),.dinb(w_n2508_0[1]),.dout(n2516),.clk(gclk));
	jor g02291(.dina(n2516),.dinb(w_n796_30[2]),.dout(n2517),.clk(gclk));
	jand g02292(.dina(w_n2508_0[0]),.dinb(w_n796_30[1]),.dout(n2518),.clk(gclk));
	jand g02293(.dina(n2518),.dinb(w_n2515_0[0]),.dout(n2519),.clk(gclk));
	jnot g02294(.din(w_n2281_0[0]),.dout(n2520),.clk(gclk));
	jand g02295(.dina(w_asqrt43_24[0]),.dinb(n2520),.dout(n2521),.clk(gclk));
	jand g02296(.dina(w_n2521_0[1]),.dinb(w_n2288_0[0]),.dout(n2522),.clk(gclk));
	jor g02297(.dina(n2522),.dinb(w_n2286_0[0]),.dout(n2523),.clk(gclk));
	jand g02298(.dina(w_n2521_0[0]),.dinb(w_n2289_0[0]),.dout(n2524),.clk(gclk));
	jnot g02299(.din(n2524),.dout(n2525),.clk(gclk));
	jand g02300(.dina(n2525),.dinb(n2523),.dout(n2526),.clk(gclk));
	jnot g02301(.din(n2526),.dout(n2527),.clk(gclk));
	jor g02302(.dina(w_n2527_0[1]),.dinb(w_n2519_0[1]),.dout(n2528),.clk(gclk));
	jand g02303(.dina(n2528),.dinb(w_n2517_0[1]),.dout(n2529),.clk(gclk));
	jor g02304(.dina(w_n2529_0[1]),.dinb(w_n791_29[0]),.dout(n2530),.clk(gclk));
	jxor g02305(.dina(w_n2290_0[0]),.dinb(w_n796_30[0]),.dout(n2531),.clk(gclk));
	jor g02306(.dina(n2531),.dinb(w_n2425_31[2]),.dout(n2532),.clk(gclk));
	jxor g02307(.dina(n2532),.dinb(w_n2295_0[0]),.dout(n2533),.clk(gclk));
	jand g02308(.dina(w_n2529_0[0]),.dinb(w_n791_28[2]),.dout(n2534),.clk(gclk));
	jor g02309(.dina(w_n2534_0[1]),.dinb(w_n2533_0[1]),.dout(n2535),.clk(gclk));
	jand g02310(.dina(w_n2535_0[2]),.dinb(w_n2530_0[2]),.dout(n2536),.clk(gclk));
	jor g02311(.dina(n2536),.dinb(w_n595_31[0]),.dout(n2537),.clk(gclk));
	jnot g02312(.din(w_n2300_0[0]),.dout(n2538),.clk(gclk));
	jor g02313(.dina(n2538),.dinb(w_n2298_0[0]),.dout(n2539),.clk(gclk));
	jor g02314(.dina(n2539),.dinb(w_n2425_31[1]),.dout(n2540),.clk(gclk));
	jxor g02315(.dina(n2540),.dinb(w_n2309_0[0]),.dout(n2541),.clk(gclk));
	jand g02316(.dina(w_n2530_0[1]),.dinb(w_n595_30[2]),.dout(n2542),.clk(gclk));
	jand g02317(.dina(n2542),.dinb(w_n2535_0[1]),.dout(n2543),.clk(gclk));
	jor g02318(.dina(w_n2543_0[1]),.dinb(w_n2541_0[1]),.dout(n2544),.clk(gclk));
	jand g02319(.dina(w_n2544_0[1]),.dinb(w_n2537_0[1]),.dout(n2545),.clk(gclk));
	jor g02320(.dina(w_n2545_0[2]),.dinb(w_n590_29[2]),.dout(n2546),.clk(gclk));
	jand g02321(.dina(w_n2545_0[1]),.dinb(w_n590_29[1]),.dout(n2547),.clk(gclk));
	jnot g02322(.din(w_n2312_0[0]),.dout(n2548),.clk(gclk));
	jand g02323(.dina(w_asqrt43_23[2]),.dinb(n2548),.dout(n2549),.clk(gclk));
	jand g02324(.dina(w_n2549_0[1]),.dinb(w_n2317_0[0]),.dout(n2550),.clk(gclk));
	jor g02325(.dina(n2550),.dinb(w_n2316_0[0]),.dout(n2551),.clk(gclk));
	jand g02326(.dina(w_n2549_0[0]),.dinb(w_n2318_0[0]),.dout(n2552),.clk(gclk));
	jnot g02327(.din(n2552),.dout(n2553),.clk(gclk));
	jand g02328(.dina(n2553),.dinb(n2551),.dout(n2554),.clk(gclk));
	jnot g02329(.din(n2554),.dout(n2555),.clk(gclk));
	jor g02330(.dina(w_n2555_0[1]),.dinb(n2547),.dout(n2556),.clk(gclk));
	jand g02331(.dina(w_n2556_0[1]),.dinb(w_n2546_0[1]),.dout(n2557),.clk(gclk));
	jor g02332(.dina(n2557),.dinb(w_n430_31[0]),.dout(n2558),.clk(gclk));
	jand g02333(.dina(w_n2546_0[0]),.dinb(w_n430_30[2]),.dout(n2559),.clk(gclk));
	jand g02334(.dina(n2559),.dinb(w_n2556_0[0]),.dout(n2560),.clk(gclk));
	jnot g02335(.din(w_n2320_0[0]),.dout(n2561),.clk(gclk));
	jand g02336(.dina(w_asqrt43_23[1]),.dinb(n2561),.dout(n2562),.clk(gclk));
	jand g02337(.dina(w_n2562_0[1]),.dinb(w_n2327_0[0]),.dout(n2563),.clk(gclk));
	jor g02338(.dina(n2563),.dinb(w_n2325_0[0]),.dout(n2564),.clk(gclk));
	jand g02339(.dina(w_n2562_0[0]),.dinb(w_n2328_0[0]),.dout(n2565),.clk(gclk));
	jnot g02340(.din(n2565),.dout(n2566),.clk(gclk));
	jand g02341(.dina(n2566),.dinb(n2564),.dout(n2567),.clk(gclk));
	jnot g02342(.din(n2567),.dout(n2568),.clk(gclk));
	jor g02343(.dina(w_n2568_0[1]),.dinb(w_n2560_0[1]),.dout(n2569),.clk(gclk));
	jand g02344(.dina(n2569),.dinb(w_n2558_0[1]),.dout(n2570),.clk(gclk));
	jor g02345(.dina(w_n2570_0[1]),.dinb(w_n425_29[2]),.dout(n2571),.clk(gclk));
	jxor g02346(.dina(w_n2329_0[0]),.dinb(w_n430_30[1]),.dout(n2572),.clk(gclk));
	jor g02347(.dina(n2572),.dinb(w_n2425_31[0]),.dout(n2573),.clk(gclk));
	jxor g02348(.dina(n2573),.dinb(w_n2340_0[0]),.dout(n2574),.clk(gclk));
	jand g02349(.dina(w_n2570_0[0]),.dinb(w_n425_29[1]),.dout(n2575),.clk(gclk));
	jor g02350(.dina(w_n2575_0[1]),.dinb(w_n2574_0[1]),.dout(n2576),.clk(gclk));
	jand g02351(.dina(w_n2576_0[2]),.dinb(w_n2571_0[2]),.dout(n2577),.clk(gclk));
	jor g02352(.dina(n2577),.dinb(w_n305_31[1]),.dout(n2578),.clk(gclk));
	jnot g02353(.din(w_n2345_0[0]),.dout(n2579),.clk(gclk));
	jor g02354(.dina(n2579),.dinb(w_n2343_0[0]),.dout(n2580),.clk(gclk));
	jor g02355(.dina(n2580),.dinb(w_n2425_30[2]),.dout(n2581),.clk(gclk));
	jxor g02356(.dina(n2581),.dinb(w_n2354_0[0]),.dout(n2582),.clk(gclk));
	jand g02357(.dina(w_n2571_0[1]),.dinb(w_n305_31[0]),.dout(n2583),.clk(gclk));
	jand g02358(.dina(n2583),.dinb(w_n2576_0[1]),.dout(n2584),.clk(gclk));
	jor g02359(.dina(w_n2584_0[1]),.dinb(w_n2582_0[1]),.dout(n2585),.clk(gclk));
	jand g02360(.dina(w_n2585_0[1]),.dinb(w_n2578_0[1]),.dout(n2586),.clk(gclk));
	jor g02361(.dina(w_n2586_0[2]),.dinb(w_n290_31[0]),.dout(n2587),.clk(gclk));
	jand g02362(.dina(w_n2586_0[1]),.dinb(w_n290_30[2]),.dout(n2588),.clk(gclk));
	jnot g02363(.din(w_n2357_0[0]),.dout(n2589),.clk(gclk));
	jand g02364(.dina(w_asqrt43_23[0]),.dinb(n2589),.dout(n2590),.clk(gclk));
	jand g02365(.dina(w_n2590_0[1]),.dinb(w_n2362_0[0]),.dout(n2591),.clk(gclk));
	jor g02366(.dina(n2591),.dinb(w_n2361_0[0]),.dout(n2592),.clk(gclk));
	jand g02367(.dina(w_n2590_0[0]),.dinb(w_n2363_0[0]),.dout(n2593),.clk(gclk));
	jnot g02368(.din(n2593),.dout(n2594),.clk(gclk));
	jand g02369(.dina(n2594),.dinb(n2592),.dout(n2595),.clk(gclk));
	jnot g02370(.din(n2595),.dout(n2596),.clk(gclk));
	jor g02371(.dina(w_n2596_0[1]),.dinb(n2588),.dout(n2597),.clk(gclk));
	jand g02372(.dina(w_n2597_0[1]),.dinb(w_n2587_0[1]),.dout(n2598),.clk(gclk));
	jor g02373(.dina(n2598),.dinb(w_n223_31[1]),.dout(n2599),.clk(gclk));
	jand g02374(.dina(w_n2587_0[0]),.dinb(w_n223_31[0]),.dout(n2600),.clk(gclk));
	jand g02375(.dina(n2600),.dinb(w_n2597_0[0]),.dout(n2601),.clk(gclk));
	jnot g02376(.din(w_n2365_0[0]),.dout(n2602),.clk(gclk));
	jand g02377(.dina(w_asqrt43_22[2]),.dinb(n2602),.dout(n2603),.clk(gclk));
	jand g02378(.dina(w_n2603_0[1]),.dinb(w_n2372_0[0]),.dout(n2604),.clk(gclk));
	jor g02379(.dina(n2604),.dinb(w_n2370_0[0]),.dout(n2605),.clk(gclk));
	jand g02380(.dina(w_n2603_0[0]),.dinb(w_n2373_0[0]),.dout(n2606),.clk(gclk));
	jnot g02381(.din(n2606),.dout(n2607),.clk(gclk));
	jand g02382(.dina(n2607),.dinb(n2605),.dout(n2608),.clk(gclk));
	jnot g02383(.din(n2608),.dout(n2609),.clk(gclk));
	jor g02384(.dina(w_n2609_0[1]),.dinb(w_n2601_0[1]),.dout(n2610),.clk(gclk));
	jand g02385(.dina(n2610),.dinb(w_n2599_0[1]),.dout(n2611),.clk(gclk));
	jor g02386(.dina(w_n2611_0[2]),.dinb(w_n199_36[1]),.dout(n2612),.clk(gclk));
	jand g02387(.dina(w_n2611_0[1]),.dinb(w_n199_36[0]),.dout(n2613),.clk(gclk));
	jxor g02388(.dina(w_n2374_0[0]),.dinb(w_n223_30[2]),.dout(n2614),.clk(gclk));
	jor g02389(.dina(n2614),.dinb(w_n2425_30[1]),.dout(n2615),.clk(gclk));
	jxor g02390(.dina(n2615),.dinb(w_n2385_0[0]),.dout(n2616),.clk(gclk));
	jor g02391(.dina(w_n2616_0[1]),.dinb(n2613),.dout(n2617),.clk(gclk));
	jand g02392(.dina(n2617),.dinb(n2612),.dout(n2618),.clk(gclk));
	jnot g02393(.din(w_n2390_0[0]),.dout(n2619),.clk(gclk));
	jor g02394(.dina(n2619),.dinb(w_n2388_0[0]),.dout(n2620),.clk(gclk));
	jor g02395(.dina(n2620),.dinb(w_n2425_30[0]),.dout(n2621),.clk(gclk));
	jxor g02396(.dina(n2621),.dinb(w_n2399_0[0]),.dout(n2622),.clk(gclk));
	jand g02397(.dina(w_asqrt43_22[1]),.dinb(w_n2413_0[1]),.dout(n2623),.clk(gclk));
	jand g02398(.dina(w_n2623_0[1]),.dinb(w_n2401_1[0]),.dout(n2624),.clk(gclk));
	jor g02399(.dina(n2624),.dinb(w_n2445_0[0]),.dout(n2625),.clk(gclk));
	jor g02400(.dina(n2625),.dinb(w_n2622_0[2]),.dout(n2626),.clk(gclk));
	jor g02401(.dina(n2626),.dinb(w_n2618_0[2]),.dout(n2627),.clk(gclk));
	jand g02402(.dina(n2627),.dinb(w_n194_35[1]),.dout(n2628),.clk(gclk));
	jand g02403(.dina(w_n2622_0[1]),.dinb(w_n2618_0[1]),.dout(n2629),.clk(gclk));
	jor g02404(.dina(w_n2623_0[0]),.dinb(w_n2401_0[2]),.dout(n2630),.clk(gclk));
	jand g02405(.dina(w_n2413_0[0]),.dinb(w_n2401_0[1]),.dout(n2631),.clk(gclk));
	jor g02406(.dina(n2631),.dinb(w_n194_35[0]),.dout(n2632),.clk(gclk));
	jnot g02407(.din(n2632),.dout(n2633),.clk(gclk));
	jand g02408(.dina(n2633),.dinb(n2630),.dout(n2634),.clk(gclk));
	jor g02409(.dina(w_n2634_0[1]),.dinb(w_n2629_0[2]),.dout(n2637),.clk(gclk));
	jor g02410(.dina(n2637),.dinb(w_n2628_0[1]),.dout(asqrt_fa_43),.clk(gclk));
	jand g02411(.dina(w_asqrt42_31),.dinb(w_a84_0[0]),.dout(n2639),.clk(gclk));
	jnot g02412(.din(w_a82_0[1]),.dout(n2640),.clk(gclk));
	jnot g02413(.din(w_a83_0[1]),.dout(n2641),.clk(gclk));
	jand g02414(.dina(w_n2428_1[0]),.dinb(w_n2641_0[1]),.dout(n2642),.clk(gclk));
	jand g02415(.dina(n2642),.dinb(w_n2640_1[1]),.dout(n2643),.clk(gclk));
	jor g02416(.dina(n2643),.dinb(n2639),.dout(n2644),.clk(gclk));
	jand g02417(.dina(w_n2644_0[2]),.dinb(w_asqrt43_22[0]),.dout(n2645),.clk(gclk));
	jand g02418(.dina(w_asqrt42_30[2]),.dinb(w_n2428_0[2]),.dout(n2646),.clk(gclk));
	jxor g02419(.dina(w_n2646_0[1]),.dinb(w_n2429_0[1]),.dout(n2647),.clk(gclk));
	jor g02420(.dina(w_n2644_0[1]),.dinb(w_asqrt43_21[2]),.dout(n2648),.clk(gclk));
	jand g02421(.dina(n2648),.dinb(w_n2647_0[1]),.dout(n2649),.clk(gclk));
	jor g02422(.dina(w_n2649_0[1]),.dinb(w_n2645_0[1]),.dout(n2650),.clk(gclk));
	jand g02423(.dina(n2650),.dinb(w_asqrt44_24[0]),.dout(n2651),.clk(gclk));
	jor g02424(.dina(w_n2645_0[0]),.dinb(w_asqrt44_23[2]),.dout(n2652),.clk(gclk));
	jor g02425(.dina(n2652),.dinb(w_n2649_0[0]),.dout(n2653),.clk(gclk));
	jand g02426(.dina(w_n2646_0[0]),.dinb(w_n2429_0[0]),.dout(n2654),.clk(gclk));
	jnot g02427(.din(w_n2628_0[0]),.dout(n2655),.clk(gclk));
	jnot g02428(.din(w_n2629_0[1]),.dout(n2656),.clk(gclk));
	jnot g02429(.din(w_n2634_0[0]),.dout(n2657),.clk(gclk));
	jand g02430(.dina(n2657),.dinb(w_asqrt43_21[1]),.dout(n2658),.clk(gclk));
	jand g02431(.dina(n2658),.dinb(n2656),.dout(n2659),.clk(gclk));
	jand g02432(.dina(n2659),.dinb(n2655),.dout(n2660),.clk(gclk));
	jor g02433(.dina(n2660),.dinb(n2654),.dout(n2661),.clk(gclk));
	jxor g02434(.dina(n2661),.dinb(w_n2209_0[1]),.dout(n2662),.clk(gclk));
	jand g02435(.dina(w_n2662_0[1]),.dinb(w_n2653_0[1]),.dout(n2663),.clk(gclk));
	jor g02436(.dina(n2663),.dinb(w_n2651_0[1]),.dout(n2664),.clk(gclk));
	jand g02437(.dina(w_n2664_0[2]),.dinb(w_asqrt45_22[0]),.dout(n2665),.clk(gclk));
	jor g02438(.dina(w_n2664_0[1]),.dinb(w_asqrt45_21[2]),.dout(n2666),.clk(gclk));
	jxor g02439(.dina(w_n2433_0[0]),.dinb(w_n2420_27[1]),.dout(n2667),.clk(gclk));
	jand g02440(.dina(n2667),.dinb(w_asqrt42_30[1]),.dout(n2668),.clk(gclk));
	jxor g02441(.dina(n2668),.dinb(w_n2436_0[0]),.dout(n2669),.clk(gclk));
	jnot g02442(.din(w_n2669_0[1]),.dout(n2670),.clk(gclk));
	jand g02443(.dina(n2670),.dinb(n2666),.dout(n2671),.clk(gclk));
	jor g02444(.dina(w_n2671_0[1]),.dinb(w_n2665_0[1]),.dout(n2672),.clk(gclk));
	jand g02445(.dina(n2672),.dinb(w_asqrt46_24[0]),.dout(n2673),.clk(gclk));
	jnot g02446(.din(w_n2442_0[0]),.dout(n2674),.clk(gclk));
	jand g02447(.dina(n2674),.dinb(w_n2440_0[0]),.dout(n2675),.clk(gclk));
	jand g02448(.dina(n2675),.dinb(w_asqrt42_30[0]),.dout(n2676),.clk(gclk));
	jxor g02449(.dina(n2676),.dinb(w_n2450_0[0]),.dout(n2677),.clk(gclk));
	jnot g02450(.din(n2677),.dout(n2678),.clk(gclk));
	jor g02451(.dina(w_n2665_0[0]),.dinb(w_asqrt46_23[2]),.dout(n2679),.clk(gclk));
	jor g02452(.dina(n2679),.dinb(w_n2671_0[0]),.dout(n2680),.clk(gclk));
	jand g02453(.dina(w_n2680_0[1]),.dinb(w_n2678_0[1]),.dout(n2681),.clk(gclk));
	jor g02454(.dina(w_n2681_0[1]),.dinb(w_n2673_0[1]),.dout(n2682),.clk(gclk));
	jand g02455(.dina(w_n2682_0[2]),.dinb(w_asqrt47_22[0]),.dout(n2683),.clk(gclk));
	jor g02456(.dina(w_n2682_0[1]),.dinb(w_asqrt47_21[2]),.dout(n2684),.clk(gclk));
	jnot g02457(.din(w_n2457_0[0]),.dout(n2685),.clk(gclk));
	jxor g02458(.dina(w_n2452_0[0]),.dinb(w_n2005_27[1]),.dout(n2686),.clk(gclk));
	jand g02459(.dina(n2686),.dinb(w_asqrt42_29[2]),.dout(n2687),.clk(gclk));
	jxor g02460(.dina(n2687),.dinb(n2685),.dout(n2688),.clk(gclk));
	jand g02461(.dina(w_n2688_0[1]),.dinb(n2684),.dout(n2689),.clk(gclk));
	jor g02462(.dina(w_n2689_0[1]),.dinb(w_n2683_0[1]),.dout(n2690),.clk(gclk));
	jand g02463(.dina(n2690),.dinb(w_asqrt48_24[0]),.dout(n2691),.clk(gclk));
	jor g02464(.dina(w_n2683_0[0]),.dinb(w_asqrt48_23[2]),.dout(n2692),.clk(gclk));
	jor g02465(.dina(n2692),.dinb(w_n2689_0[0]),.dout(n2693),.clk(gclk));
	jnot g02466(.din(w_n2464_0[0]),.dout(n2694),.clk(gclk));
	jnot g02467(.din(w_n2466_0[0]),.dout(n2695),.clk(gclk));
	jand g02468(.dina(w_asqrt42_29[1]),.dinb(w_n2460_0[0]),.dout(n2696),.clk(gclk));
	jand g02469(.dina(w_n2696_0[1]),.dinb(n2695),.dout(n2697),.clk(gclk));
	jor g02470(.dina(n2697),.dinb(n2694),.dout(n2698),.clk(gclk));
	jnot g02471(.din(w_n2467_0[0]),.dout(n2699),.clk(gclk));
	jand g02472(.dina(w_n2696_0[0]),.dinb(n2699),.dout(n2700),.clk(gclk));
	jnot g02473(.din(n2700),.dout(n2701),.clk(gclk));
	jand g02474(.dina(n2701),.dinb(n2698),.dout(n2702),.clk(gclk));
	jand g02475(.dina(w_n2702_0[1]),.dinb(w_n2693_0[1]),.dout(n2703),.clk(gclk));
	jor g02476(.dina(n2703),.dinb(w_n2691_0[1]),.dout(n2704),.clk(gclk));
	jand g02477(.dina(w_n2704_0[2]),.dinb(w_asqrt49_22[1]),.dout(n2705),.clk(gclk));
	jor g02478(.dina(w_n2704_0[1]),.dinb(w_asqrt49_22[0]),.dout(n2706),.clk(gclk));
	jxor g02479(.dina(w_n2468_0[0]),.dinb(w_n1641_27[2]),.dout(n2707),.clk(gclk));
	jand g02480(.dina(n2707),.dinb(w_asqrt42_29[0]),.dout(n2708),.clk(gclk));
	jxor g02481(.dina(n2708),.dinb(w_n2473_0[0]),.dout(n2709),.clk(gclk));
	jand g02482(.dina(w_n2709_0[1]),.dinb(n2706),.dout(n2710),.clk(gclk));
	jor g02483(.dina(w_n2710_0[1]),.dinb(w_n2705_0[1]),.dout(n2711),.clk(gclk));
	jand g02484(.dina(n2711),.dinb(w_asqrt50_24[0]),.dout(n2712),.clk(gclk));
	jnot g02485(.din(w_n2479_0[0]),.dout(n2713),.clk(gclk));
	jand g02486(.dina(n2713),.dinb(w_n2477_0[0]),.dout(n2714),.clk(gclk));
	jand g02487(.dina(n2714),.dinb(w_asqrt42_28[2]),.dout(n2715),.clk(gclk));
	jxor g02488(.dina(n2715),.dinb(w_n2487_0[0]),.dout(n2716),.clk(gclk));
	jnot g02489(.din(n2716),.dout(n2717),.clk(gclk));
	jor g02490(.dina(w_n2705_0[0]),.dinb(w_asqrt50_23[2]),.dout(n2718),.clk(gclk));
	jor g02491(.dina(n2718),.dinb(w_n2710_0[0]),.dout(n2719),.clk(gclk));
	jand g02492(.dina(w_n2719_0[1]),.dinb(w_n2717_0[1]),.dout(n2720),.clk(gclk));
	jor g02493(.dina(w_n2720_0[1]),.dinb(w_n2712_0[1]),.dout(n2721),.clk(gclk));
	jand g02494(.dina(w_n2721_0[2]),.dinb(w_asqrt51_22[1]),.dout(n2722),.clk(gclk));
	jor g02495(.dina(w_n2721_0[1]),.dinb(w_asqrt51_22[0]),.dout(n2723),.clk(gclk));
	jxor g02496(.dina(w_n2489_0[0]),.dinb(w_n1312_27[2]),.dout(n2724),.clk(gclk));
	jand g02497(.dina(n2724),.dinb(w_asqrt42_28[1]),.dout(n2725),.clk(gclk));
	jxor g02498(.dina(n2725),.dinb(w_n2495_0[0]),.dout(n2726),.clk(gclk));
	jand g02499(.dina(w_n2726_0[1]),.dinb(n2723),.dout(n2727),.clk(gclk));
	jor g02500(.dina(w_n2727_0[1]),.dinb(w_n2722_0[1]),.dout(n2728),.clk(gclk));
	jand g02501(.dina(n2728),.dinb(w_asqrt52_24[0]),.dout(n2729),.clk(gclk));
	jor g02502(.dina(w_n2722_0[0]),.dinb(w_asqrt52_23[2]),.dout(n2730),.clk(gclk));
	jor g02503(.dina(n2730),.dinb(w_n2727_0[0]),.dout(n2731),.clk(gclk));
	jnot g02504(.din(w_n2503_0[0]),.dout(n2732),.clk(gclk));
	jnot g02505(.din(w_n2505_0[0]),.dout(n2733),.clk(gclk));
	jand g02506(.dina(w_asqrt42_28[0]),.dinb(w_n2499_0[0]),.dout(n2734),.clk(gclk));
	jand g02507(.dina(w_n2734_0[1]),.dinb(n2733),.dout(n2735),.clk(gclk));
	jor g02508(.dina(n2735),.dinb(n2732),.dout(n2736),.clk(gclk));
	jnot g02509(.din(w_n2506_0[0]),.dout(n2737),.clk(gclk));
	jand g02510(.dina(w_n2734_0[0]),.dinb(n2737),.dout(n2738),.clk(gclk));
	jnot g02511(.din(n2738),.dout(n2739),.clk(gclk));
	jand g02512(.dina(n2739),.dinb(n2736),.dout(n2740),.clk(gclk));
	jand g02513(.dina(w_n2740_0[1]),.dinb(w_n2731_0[1]),.dout(n2741),.clk(gclk));
	jor g02514(.dina(n2741),.dinb(w_n2729_0[1]),.dout(n2742),.clk(gclk));
	jand g02515(.dina(w_n2742_0[1]),.dinb(w_asqrt53_22[2]),.dout(n2743),.clk(gclk));
	jxor g02516(.dina(w_n2507_0[0]),.dinb(w_n1034_28[1]),.dout(n2744),.clk(gclk));
	jand g02517(.dina(n2744),.dinb(w_asqrt42_27[2]),.dout(n2745),.clk(gclk));
	jxor g02518(.dina(n2745),.dinb(w_n2514_0[0]),.dout(n2746),.clk(gclk));
	jnot g02519(.din(n2746),.dout(n2747),.clk(gclk));
	jor g02520(.dina(w_n2742_0[0]),.dinb(w_asqrt53_22[1]),.dout(n2748),.clk(gclk));
	jand g02521(.dina(w_n2748_0[1]),.dinb(w_n2747_0[1]),.dout(n2749),.clk(gclk));
	jor g02522(.dina(w_n2749_0[2]),.dinb(w_n2743_0[2]),.dout(n2750),.clk(gclk));
	jand g02523(.dina(n2750),.dinb(w_asqrt54_24[0]),.dout(n2751),.clk(gclk));
	jnot g02524(.din(w_n2519_0[0]),.dout(n2752),.clk(gclk));
	jand g02525(.dina(n2752),.dinb(w_n2517_0[0]),.dout(n2753),.clk(gclk));
	jand g02526(.dina(n2753),.dinb(w_asqrt42_27[1]),.dout(n2754),.clk(gclk));
	jxor g02527(.dina(n2754),.dinb(w_n2527_0[0]),.dout(n2755),.clk(gclk));
	jnot g02528(.din(n2755),.dout(n2756),.clk(gclk));
	jor g02529(.dina(w_n2743_0[1]),.dinb(w_asqrt54_23[2]),.dout(n2757),.clk(gclk));
	jor g02530(.dina(n2757),.dinb(w_n2749_0[1]),.dout(n2758),.clk(gclk));
	jand g02531(.dina(w_n2758_0[1]),.dinb(w_n2756_0[1]),.dout(n2759),.clk(gclk));
	jor g02532(.dina(w_n2759_0[1]),.dinb(w_n2751_0[1]),.dout(n2760),.clk(gclk));
	jand g02533(.dina(w_n2760_0[2]),.dinb(w_asqrt55_23[0]),.dout(n2761),.clk(gclk));
	jor g02534(.dina(w_n2760_0[1]),.dinb(w_asqrt55_22[2]),.dout(n2762),.clk(gclk));
	jnot g02535(.din(w_n2533_0[0]),.dout(n2763),.clk(gclk));
	jnot g02536(.din(w_n2534_0[0]),.dout(n2764),.clk(gclk));
	jand g02537(.dina(w_asqrt42_27[0]),.dinb(w_n2530_0[0]),.dout(n2765),.clk(gclk));
	jand g02538(.dina(w_n2765_0[1]),.dinb(n2764),.dout(n2766),.clk(gclk));
	jor g02539(.dina(n2766),.dinb(n2763),.dout(n2767),.clk(gclk));
	jnot g02540(.din(w_n2535_0[0]),.dout(n2768),.clk(gclk));
	jand g02541(.dina(w_n2765_0[0]),.dinb(n2768),.dout(n2769),.clk(gclk));
	jnot g02542(.din(n2769),.dout(n2770),.clk(gclk));
	jand g02543(.dina(n2770),.dinb(n2767),.dout(n2771),.clk(gclk));
	jand g02544(.dina(w_n2771_0[1]),.dinb(n2762),.dout(n2772),.clk(gclk));
	jor g02545(.dina(w_n2772_0[1]),.dinb(w_n2761_0[1]),.dout(n2773),.clk(gclk));
	jand g02546(.dina(n2773),.dinb(w_asqrt56_24[0]),.dout(n2774),.clk(gclk));
	jor g02547(.dina(w_n2761_0[0]),.dinb(w_asqrt56_23[2]),.dout(n2775),.clk(gclk));
	jor g02548(.dina(n2775),.dinb(w_n2772_0[0]),.dout(n2776),.clk(gclk));
	jnot g02549(.din(w_n2541_0[0]),.dout(n2777),.clk(gclk));
	jnot g02550(.din(w_n2543_0[0]),.dout(n2778),.clk(gclk));
	jand g02551(.dina(w_asqrt42_26[2]),.dinb(w_n2537_0[0]),.dout(n2779),.clk(gclk));
	jand g02552(.dina(w_n2779_0[1]),.dinb(n2778),.dout(n2780),.clk(gclk));
	jor g02553(.dina(n2780),.dinb(n2777),.dout(n2781),.clk(gclk));
	jnot g02554(.din(w_n2544_0[0]),.dout(n2782),.clk(gclk));
	jand g02555(.dina(w_n2779_0[0]),.dinb(n2782),.dout(n2783),.clk(gclk));
	jnot g02556(.din(n2783),.dout(n2784),.clk(gclk));
	jand g02557(.dina(n2784),.dinb(n2781),.dout(n2785),.clk(gclk));
	jand g02558(.dina(w_n2785_0[1]),.dinb(w_n2776_0[1]),.dout(n2786),.clk(gclk));
	jor g02559(.dina(n2786),.dinb(w_n2774_0[1]),.dout(n2787),.clk(gclk));
	jand g02560(.dina(w_n2787_0[1]),.dinb(w_asqrt57_23[1]),.dout(n2788),.clk(gclk));
	jxor g02561(.dina(w_n2545_0[0]),.dinb(w_n590_29[0]),.dout(n2789),.clk(gclk));
	jand g02562(.dina(n2789),.dinb(w_asqrt42_26[1]),.dout(n2790),.clk(gclk));
	jxor g02563(.dina(n2790),.dinb(w_n2555_0[0]),.dout(n2791),.clk(gclk));
	jnot g02564(.din(n2791),.dout(n2792),.clk(gclk));
	jor g02565(.dina(w_n2787_0[0]),.dinb(w_asqrt57_23[0]),.dout(n2793),.clk(gclk));
	jand g02566(.dina(w_n2793_0[1]),.dinb(w_n2792_0[1]),.dout(n2794),.clk(gclk));
	jor g02567(.dina(w_n2794_0[2]),.dinb(w_n2788_0[2]),.dout(n2795),.clk(gclk));
	jand g02568(.dina(n2795),.dinb(w_asqrt58_24[0]),.dout(n2796),.clk(gclk));
	jnot g02569(.din(w_n2560_0[0]),.dout(n2797),.clk(gclk));
	jand g02570(.dina(n2797),.dinb(w_n2558_0[0]),.dout(n2798),.clk(gclk));
	jand g02571(.dina(n2798),.dinb(w_asqrt42_26[0]),.dout(n2799),.clk(gclk));
	jxor g02572(.dina(n2799),.dinb(w_n2568_0[0]),.dout(n2800),.clk(gclk));
	jnot g02573(.din(n2800),.dout(n2801),.clk(gclk));
	jor g02574(.dina(w_n2788_0[1]),.dinb(w_asqrt58_23[2]),.dout(n2802),.clk(gclk));
	jor g02575(.dina(n2802),.dinb(w_n2794_0[1]),.dout(n2803),.clk(gclk));
	jand g02576(.dina(w_n2803_0[1]),.dinb(w_n2801_0[1]),.dout(n2804),.clk(gclk));
	jor g02577(.dina(w_n2804_0[1]),.dinb(w_n2796_0[1]),.dout(n2805),.clk(gclk));
	jand g02578(.dina(w_n2805_0[2]),.dinb(w_asqrt59_23[2]),.dout(n2806),.clk(gclk));
	jor g02579(.dina(w_n2805_0[1]),.dinb(w_asqrt59_23[1]),.dout(n2807),.clk(gclk));
	jnot g02580(.din(w_n2574_0[0]),.dout(n2808),.clk(gclk));
	jnot g02581(.din(w_n2575_0[0]),.dout(n2809),.clk(gclk));
	jand g02582(.dina(w_asqrt42_25[2]),.dinb(w_n2571_0[0]),.dout(n2810),.clk(gclk));
	jand g02583(.dina(w_n2810_0[1]),.dinb(n2809),.dout(n2811),.clk(gclk));
	jor g02584(.dina(n2811),.dinb(n2808),.dout(n2812),.clk(gclk));
	jnot g02585(.din(w_n2576_0[0]),.dout(n2813),.clk(gclk));
	jand g02586(.dina(w_n2810_0[0]),.dinb(n2813),.dout(n2814),.clk(gclk));
	jnot g02587(.din(n2814),.dout(n2815),.clk(gclk));
	jand g02588(.dina(n2815),.dinb(n2812),.dout(n2816),.clk(gclk));
	jand g02589(.dina(w_n2816_0[1]),.dinb(n2807),.dout(n2817),.clk(gclk));
	jor g02590(.dina(w_n2817_0[1]),.dinb(w_n2806_0[1]),.dout(n2818),.clk(gclk));
	jand g02591(.dina(n2818),.dinb(w_asqrt60_23[2]),.dout(n2819),.clk(gclk));
	jor g02592(.dina(w_n2806_0[0]),.dinb(w_asqrt60_23[1]),.dout(n2820),.clk(gclk));
	jor g02593(.dina(n2820),.dinb(w_n2817_0[0]),.dout(n2821),.clk(gclk));
	jnot g02594(.din(w_n2582_0[0]),.dout(n2822),.clk(gclk));
	jnot g02595(.din(w_n2584_0[0]),.dout(n2823),.clk(gclk));
	jand g02596(.dina(w_asqrt42_25[1]),.dinb(w_n2578_0[0]),.dout(n2824),.clk(gclk));
	jand g02597(.dina(w_n2824_0[1]),.dinb(n2823),.dout(n2825),.clk(gclk));
	jor g02598(.dina(n2825),.dinb(n2822),.dout(n2826),.clk(gclk));
	jnot g02599(.din(w_n2585_0[0]),.dout(n2827),.clk(gclk));
	jand g02600(.dina(w_n2824_0[0]),.dinb(n2827),.dout(n2828),.clk(gclk));
	jnot g02601(.din(n2828),.dout(n2829),.clk(gclk));
	jand g02602(.dina(n2829),.dinb(n2826),.dout(n2830),.clk(gclk));
	jand g02603(.dina(w_n2830_0[1]),.dinb(w_n2821_0[1]),.dout(n2831),.clk(gclk));
	jor g02604(.dina(n2831),.dinb(w_n2819_0[1]),.dout(n2832),.clk(gclk));
	jand g02605(.dina(w_n2832_0[1]),.dinb(w_asqrt61_24[0]),.dout(n2833),.clk(gclk));
	jxor g02606(.dina(w_n2586_0[0]),.dinb(w_n290_30[1]),.dout(n2834),.clk(gclk));
	jand g02607(.dina(n2834),.dinb(w_asqrt42_25[0]),.dout(n2835),.clk(gclk));
	jxor g02608(.dina(n2835),.dinb(w_n2596_0[0]),.dout(n2836),.clk(gclk));
	jnot g02609(.din(n2836),.dout(n2837),.clk(gclk));
	jor g02610(.dina(w_n2832_0[0]),.dinb(w_asqrt61_23[2]),.dout(n2838),.clk(gclk));
	jand g02611(.dina(w_n2838_0[1]),.dinb(w_n2837_0[1]),.dout(n2839),.clk(gclk));
	jor g02612(.dina(w_n2839_0[2]),.dinb(w_n2833_0[2]),.dout(n2840),.clk(gclk));
	jand g02613(.dina(n2840),.dinb(w_asqrt62_24[0]),.dout(n2841),.clk(gclk));
	jnot g02614(.din(w_n2601_0[0]),.dout(n2842),.clk(gclk));
	jand g02615(.dina(n2842),.dinb(w_n2599_0[0]),.dout(n2843),.clk(gclk));
	jand g02616(.dina(n2843),.dinb(w_asqrt42_24[2]),.dout(n2844),.clk(gclk));
	jxor g02617(.dina(n2844),.dinb(w_n2609_0[0]),.dout(n2845),.clk(gclk));
	jnot g02618(.din(n2845),.dout(n2846),.clk(gclk));
	jor g02619(.dina(w_n2833_0[1]),.dinb(w_asqrt62_23[2]),.dout(n2847),.clk(gclk));
	jor g02620(.dina(n2847),.dinb(w_n2839_0[1]),.dout(n2848),.clk(gclk));
	jand g02621(.dina(w_n2848_0[1]),.dinb(w_n2846_0[1]),.dout(n2849),.clk(gclk));
	jor g02622(.dina(w_n2849_0[1]),.dinb(w_n2841_0[1]),.dout(n2850),.clk(gclk));
	jxor g02623(.dina(w_n2611_0[0]),.dinb(w_n199_35[2]),.dout(n2851),.clk(gclk));
	jand g02624(.dina(n2851),.dinb(w_asqrt42_24[1]),.dout(n2852),.clk(gclk));
	jxor g02625(.dina(n2852),.dinb(w_n2616_0[0]),.dout(n2853),.clk(gclk));
	jnot g02626(.din(w_n2618_0[0]),.dout(n2854),.clk(gclk));
	jnot g02627(.din(w_n2622_0[0]),.dout(n2855),.clk(gclk));
	jand g02628(.dina(w_asqrt42_24[0]),.dinb(w_n2855_0[1]),.dout(n2856),.clk(gclk));
	jand g02629(.dina(w_n2856_0[1]),.dinb(w_n2854_0[2]),.dout(n2857),.clk(gclk));
	jor g02630(.dina(n2857),.dinb(w_n2629_0[0]),.dout(n2858),.clk(gclk));
	jor g02631(.dina(n2858),.dinb(w_n2853_0[1]),.dout(n2859),.clk(gclk));
	jnot g02632(.din(n2859),.dout(n2860),.clk(gclk));
	jand g02633(.dina(n2860),.dinb(w_n2850_1[2]),.dout(n2861),.clk(gclk));
	jor g02634(.dina(n2861),.dinb(w_asqrt63_12[2]),.dout(n2862),.clk(gclk));
	jnot g02635(.din(w_n2853_0[0]),.dout(n2863),.clk(gclk));
	jor g02636(.dina(w_n2863_0[2]),.dinb(w_n2850_1[1]),.dout(n2864),.clk(gclk));
	jor g02637(.dina(w_n2856_0[0]),.dinb(w_n2854_0[1]),.dout(n2865),.clk(gclk));
	jand g02638(.dina(w_n2855_0[0]),.dinb(w_n2854_0[0]),.dout(n2866),.clk(gclk));
	jor g02639(.dina(n2866),.dinb(w_n194_34[2]),.dout(n2867),.clk(gclk));
	jnot g02640(.din(n2867),.dout(n2868),.clk(gclk));
	jand g02641(.dina(n2868),.dinb(n2865),.dout(n2869),.clk(gclk));
	jnot g02642(.din(w_asqrt42_23[2]),.dout(n2870),.clk(gclk));
	jnot g02643(.din(w_n2869_0[1]),.dout(n2873),.clk(gclk));
	jand g02644(.dina(n2873),.dinb(w_n2864_0[1]),.dout(n2874),.clk(gclk));
	jand g02645(.dina(n2874),.dinb(w_n2862_0[1]),.dout(n2875),.clk(gclk));
	jnot g02646(.din(w_n2875_33[1]),.dout(asqrt_fa_42),.clk(gclk));
	jor g02647(.dina(w_n2875_33[0]),.dinb(w_n2640_1[0]),.dout(n2877),.clk(gclk));
	jnot g02648(.din(w_a80_0[1]),.dout(n2878),.clk(gclk));
	jnot g02649(.din(a[81]),.dout(n2879),.clk(gclk));
	jand g02650(.dina(w_n2640_0[2]),.dinb(w_n2879_0[2]),.dout(n2880),.clk(gclk));
	jand g02651(.dina(n2880),.dinb(w_n2878_1[1]),.dout(n2881),.clk(gclk));
	jnot g02652(.din(n2881),.dout(n2882),.clk(gclk));
	jand g02653(.dina(n2882),.dinb(n2877),.dout(n2883),.clk(gclk));
	jor g02654(.dina(w_n2883_0[2]),.dinb(w_n2870_26[2]),.dout(n2884),.clk(gclk));
	jor g02655(.dina(w_n2875_32[2]),.dinb(w_a82_0[0]),.dout(n2885),.clk(gclk));
	jxor g02656(.dina(w_n2885_0[1]),.dinb(w_n2641_0[0]),.dout(n2886),.clk(gclk));
	jand g02657(.dina(w_n2883_0[1]),.dinb(w_n2870_26[1]),.dout(n2887),.clk(gclk));
	jor g02658(.dina(n2887),.dinb(w_n2886_0[1]),.dout(n2888),.clk(gclk));
	jand g02659(.dina(w_n2888_0[1]),.dinb(w_n2884_0[1]),.dout(n2889),.clk(gclk));
	jor g02660(.dina(n2889),.dinb(w_n2425_29[2]),.dout(n2890),.clk(gclk));
	jand g02661(.dina(w_n2884_0[0]),.dinb(w_n2425_29[1]),.dout(n2891),.clk(gclk));
	jand g02662(.dina(n2891),.dinb(w_n2888_0[0]),.dout(n2892),.clk(gclk));
	jor g02663(.dina(w_n2885_0[0]),.dinb(w_a83_0[0]),.dout(n2893),.clk(gclk));
	jnot g02664(.din(w_n2862_0[0]),.dout(n2894),.clk(gclk));
	jnot g02665(.din(w_n2864_0[0]),.dout(n2895),.clk(gclk));
	jor g02666(.dina(w_n2869_0[0]),.dinb(w_n2870_26[0]),.dout(n2896),.clk(gclk));
	jor g02667(.dina(n2896),.dinb(w_n2895_0[1]),.dout(n2897),.clk(gclk));
	jor g02668(.dina(n2897),.dinb(n2894),.dout(n2898),.clk(gclk));
	jand g02669(.dina(n2898),.dinb(n2893),.dout(n2899),.clk(gclk));
	jxor g02670(.dina(n2899),.dinb(w_n2428_0[1]),.dout(n2900),.clk(gclk));
	jor g02671(.dina(w_n2900_0[1]),.dinb(w_n2892_0[1]),.dout(n2901),.clk(gclk));
	jand g02672(.dina(n2901),.dinb(w_n2890_0[1]),.dout(n2902),.clk(gclk));
	jor g02673(.dina(w_n2902_0[2]),.dinb(w_n2420_27[0]),.dout(n2903),.clk(gclk));
	jand g02674(.dina(w_n2902_0[1]),.dinb(w_n2420_26[2]),.dout(n2904),.clk(gclk));
	jxor g02675(.dina(w_n2644_0[0]),.dinb(w_n2425_29[0]),.dout(n2905),.clk(gclk));
	jor g02676(.dina(n2905),.dinb(w_n2875_32[1]),.dout(n2906),.clk(gclk));
	jxor g02677(.dina(n2906),.dinb(w_n2647_0[0]),.dout(n2907),.clk(gclk));
	jor g02678(.dina(w_n2907_0[1]),.dinb(n2904),.dout(n2908),.clk(gclk));
	jand g02679(.dina(w_n2908_0[1]),.dinb(w_n2903_0[1]),.dout(n2909),.clk(gclk));
	jor g02680(.dina(n2909),.dinb(w_n2010_29[1]),.dout(n2910),.clk(gclk));
	jnot g02681(.din(w_n2653_0[0]),.dout(n2911),.clk(gclk));
	jor g02682(.dina(n2911),.dinb(w_n2651_0[0]),.dout(n2912),.clk(gclk));
	jor g02683(.dina(n2912),.dinb(w_n2875_32[0]),.dout(n2913),.clk(gclk));
	jxor g02684(.dina(n2913),.dinb(w_n2662_0[0]),.dout(n2914),.clk(gclk));
	jand g02685(.dina(w_n2903_0[0]),.dinb(w_n2010_29[0]),.dout(n2915),.clk(gclk));
	jand g02686(.dina(n2915),.dinb(w_n2908_0[0]),.dout(n2916),.clk(gclk));
	jor g02687(.dina(w_n2916_0[1]),.dinb(w_n2914_0[1]),.dout(n2917),.clk(gclk));
	jand g02688(.dina(w_n2917_0[1]),.dinb(w_n2910_0[1]),.dout(n2918),.clk(gclk));
	jor g02689(.dina(w_n2918_0[2]),.dinb(w_n2005_27[0]),.dout(n2919),.clk(gclk));
	jand g02690(.dina(w_n2918_0[1]),.dinb(w_n2005_26[2]),.dout(n2920),.clk(gclk));
	jxor g02691(.dina(w_n2664_0[0]),.dinb(w_n2010_28[2]),.dout(n2921),.clk(gclk));
	jor g02692(.dina(n2921),.dinb(w_n2875_31[2]),.dout(n2922),.clk(gclk));
	jxor g02693(.dina(n2922),.dinb(w_n2669_0[0]),.dout(n2923),.clk(gclk));
	jnot g02694(.din(w_n2923_0[1]),.dout(n2924),.clk(gclk));
	jor g02695(.dina(n2924),.dinb(n2920),.dout(n2925),.clk(gclk));
	jand g02696(.dina(w_n2925_0[1]),.dinb(w_n2919_0[1]),.dout(n2926),.clk(gclk));
	jor g02697(.dina(n2926),.dinb(w_n1646_30[0]),.dout(n2927),.clk(gclk));
	jand g02698(.dina(w_n2919_0[0]),.dinb(w_n1646_29[2]),.dout(n2928),.clk(gclk));
	jand g02699(.dina(n2928),.dinb(w_n2925_0[0]),.dout(n2929),.clk(gclk));
	jnot g02700(.din(w_n2673_0[0]),.dout(n2930),.clk(gclk));
	jand g02701(.dina(w_asqrt41_24[1]),.dinb(n2930),.dout(n2931),.clk(gclk));
	jand g02702(.dina(w_n2931_0[1]),.dinb(w_n2680_0[0]),.dout(n2932),.clk(gclk));
	jor g02703(.dina(n2932),.dinb(w_n2678_0[0]),.dout(n2933),.clk(gclk));
	jand g02704(.dina(w_n2931_0[0]),.dinb(w_n2681_0[0]),.dout(n2934),.clk(gclk));
	jnot g02705(.din(n2934),.dout(n2935),.clk(gclk));
	jand g02706(.dina(n2935),.dinb(n2933),.dout(n2936),.clk(gclk));
	jnot g02707(.din(n2936),.dout(n2937),.clk(gclk));
	jor g02708(.dina(w_n2937_0[1]),.dinb(w_n2929_0[1]),.dout(n2938),.clk(gclk));
	jand g02709(.dina(n2938),.dinb(w_n2927_0[1]),.dout(n2939),.clk(gclk));
	jor g02710(.dina(w_n2939_0[2]),.dinb(w_n1641_27[1]),.dout(n2940),.clk(gclk));
	jand g02711(.dina(w_n2939_0[1]),.dinb(w_n1641_27[0]),.dout(n2941),.clk(gclk));
	jnot g02712(.din(w_n2688_0[0]),.dout(n2942),.clk(gclk));
	jxor g02713(.dina(w_n2682_0[0]),.dinb(w_n1646_29[1]),.dout(n2943),.clk(gclk));
	jor g02714(.dina(n2943),.dinb(w_n2875_31[1]),.dout(n2944),.clk(gclk));
	jxor g02715(.dina(n2944),.dinb(n2942),.dout(n2945),.clk(gclk));
	jnot g02716(.din(w_n2945_0[1]),.dout(n2946),.clk(gclk));
	jor g02717(.dina(n2946),.dinb(n2941),.dout(n2947),.clk(gclk));
	jand g02718(.dina(w_n2947_0[1]),.dinb(w_n2940_0[1]),.dout(n2948),.clk(gclk));
	jor g02719(.dina(n2948),.dinb(w_n1317_29[2]),.dout(n2949),.clk(gclk));
	jnot g02720(.din(w_n2693_0[0]),.dout(n2950),.clk(gclk));
	jor g02721(.dina(n2950),.dinb(w_n2691_0[0]),.dout(n2951),.clk(gclk));
	jor g02722(.dina(n2951),.dinb(w_n2875_31[0]),.dout(n2952),.clk(gclk));
	jxor g02723(.dina(n2952),.dinb(w_n2702_0[0]),.dout(n2953),.clk(gclk));
	jand g02724(.dina(w_n2940_0[0]),.dinb(w_n1317_29[1]),.dout(n2954),.clk(gclk));
	jand g02725(.dina(n2954),.dinb(w_n2947_0[0]),.dout(n2955),.clk(gclk));
	jor g02726(.dina(w_n2955_0[1]),.dinb(w_n2953_0[1]),.dout(n2956),.clk(gclk));
	jand g02727(.dina(w_n2956_0[1]),.dinb(w_n2949_0[1]),.dout(n2957),.clk(gclk));
	jor g02728(.dina(w_n2957_0[2]),.dinb(w_n1312_27[1]),.dout(n2958),.clk(gclk));
	jand g02729(.dina(w_n2957_0[1]),.dinb(w_n1312_27[0]),.dout(n2959),.clk(gclk));
	jnot g02730(.din(w_n2709_0[0]),.dout(n2960),.clk(gclk));
	jxor g02731(.dina(w_n2704_0[0]),.dinb(w_n1317_29[0]),.dout(n2961),.clk(gclk));
	jor g02732(.dina(n2961),.dinb(w_n2875_30[2]),.dout(n2962),.clk(gclk));
	jxor g02733(.dina(n2962),.dinb(n2960),.dout(n2963),.clk(gclk));
	jnot g02734(.din(n2963),.dout(n2964),.clk(gclk));
	jor g02735(.dina(w_n2964_0[1]),.dinb(n2959),.dout(n2965),.clk(gclk));
	jand g02736(.dina(w_n2965_0[1]),.dinb(w_n2958_0[1]),.dout(n2966),.clk(gclk));
	jor g02737(.dina(n2966),.dinb(w_n1039_30[0]),.dout(n2967),.clk(gclk));
	jand g02738(.dina(w_n2958_0[0]),.dinb(w_n1039_29[2]),.dout(n2968),.clk(gclk));
	jand g02739(.dina(n2968),.dinb(w_n2965_0[0]),.dout(n2969),.clk(gclk));
	jnot g02740(.din(w_n2712_0[0]),.dout(n2970),.clk(gclk));
	jand g02741(.dina(w_asqrt41_24[0]),.dinb(n2970),.dout(n2971),.clk(gclk));
	jand g02742(.dina(w_n2971_0[1]),.dinb(w_n2719_0[0]),.dout(n2972),.clk(gclk));
	jor g02743(.dina(n2972),.dinb(w_n2717_0[0]),.dout(n2973),.clk(gclk));
	jand g02744(.dina(w_n2971_0[0]),.dinb(w_n2720_0[0]),.dout(n2974),.clk(gclk));
	jnot g02745(.din(n2974),.dout(n2975),.clk(gclk));
	jand g02746(.dina(n2975),.dinb(n2973),.dout(n2976),.clk(gclk));
	jnot g02747(.din(n2976),.dout(n2977),.clk(gclk));
	jor g02748(.dina(w_n2977_0[1]),.dinb(w_n2969_0[1]),.dout(n2978),.clk(gclk));
	jand g02749(.dina(n2978),.dinb(w_n2967_0[1]),.dout(n2979),.clk(gclk));
	jor g02750(.dina(w_n2979_0[1]),.dinb(w_n1034_28[0]),.dout(n2980),.clk(gclk));
	jxor g02751(.dina(w_n2721_0[0]),.dinb(w_n1039_29[1]),.dout(n2981),.clk(gclk));
	jor g02752(.dina(n2981),.dinb(w_n2875_30[1]),.dout(n2982),.clk(gclk));
	jxor g02753(.dina(n2982),.dinb(w_n2726_0[0]),.dout(n2983),.clk(gclk));
	jand g02754(.dina(w_n2979_0[0]),.dinb(w_n1034_27[2]),.dout(n2984),.clk(gclk));
	jor g02755(.dina(w_n2984_0[1]),.dinb(w_n2983_0[1]),.dout(n2985),.clk(gclk));
	jand g02756(.dina(w_n2985_0[2]),.dinb(w_n2980_0[2]),.dout(n2986),.clk(gclk));
	jor g02757(.dina(n2986),.dinb(w_n796_29[2]),.dout(n2987),.clk(gclk));
	jnot g02758(.din(w_n2731_0[0]),.dout(n2988),.clk(gclk));
	jor g02759(.dina(n2988),.dinb(w_n2729_0[0]),.dout(n2989),.clk(gclk));
	jor g02760(.dina(n2989),.dinb(w_n2875_30[0]),.dout(n2990),.clk(gclk));
	jxor g02761(.dina(n2990),.dinb(w_n2740_0[0]),.dout(n2991),.clk(gclk));
	jand g02762(.dina(w_n2980_0[1]),.dinb(w_n796_29[1]),.dout(n2992),.clk(gclk));
	jand g02763(.dina(n2992),.dinb(w_n2985_0[1]),.dout(n2993),.clk(gclk));
	jor g02764(.dina(w_n2993_0[1]),.dinb(w_n2991_0[1]),.dout(n2994),.clk(gclk));
	jand g02765(.dina(w_n2994_0[1]),.dinb(w_n2987_0[1]),.dout(n2995),.clk(gclk));
	jor g02766(.dina(w_n2995_0[2]),.dinb(w_n791_28[1]),.dout(n2996),.clk(gclk));
	jand g02767(.dina(w_n2995_0[1]),.dinb(w_n791_28[0]),.dout(n2997),.clk(gclk));
	jnot g02768(.din(w_n2743_0[0]),.dout(n2998),.clk(gclk));
	jand g02769(.dina(w_asqrt41_23[2]),.dinb(n2998),.dout(n2999),.clk(gclk));
	jand g02770(.dina(w_n2999_0[1]),.dinb(w_n2748_0[0]),.dout(n3000),.clk(gclk));
	jor g02771(.dina(n3000),.dinb(w_n2747_0[0]),.dout(n3001),.clk(gclk));
	jand g02772(.dina(w_n2999_0[0]),.dinb(w_n2749_0[0]),.dout(n3002),.clk(gclk));
	jnot g02773(.din(n3002),.dout(n3003),.clk(gclk));
	jand g02774(.dina(n3003),.dinb(n3001),.dout(n3004),.clk(gclk));
	jnot g02775(.din(n3004),.dout(n3005),.clk(gclk));
	jor g02776(.dina(w_n3005_0[1]),.dinb(n2997),.dout(n3006),.clk(gclk));
	jand g02777(.dina(w_n3006_0[1]),.dinb(w_n2996_0[1]),.dout(n3007),.clk(gclk));
	jor g02778(.dina(n3007),.dinb(w_n595_30[1]),.dout(n3008),.clk(gclk));
	jand g02779(.dina(w_n2996_0[0]),.dinb(w_n595_30[0]),.dout(n3009),.clk(gclk));
	jand g02780(.dina(n3009),.dinb(w_n3006_0[0]),.dout(n3010),.clk(gclk));
	jnot g02781(.din(w_n2751_0[0]),.dout(n3011),.clk(gclk));
	jand g02782(.dina(w_asqrt41_23[1]),.dinb(n3011),.dout(n3012),.clk(gclk));
	jand g02783(.dina(w_n3012_0[1]),.dinb(w_n2758_0[0]),.dout(n3013),.clk(gclk));
	jor g02784(.dina(n3013),.dinb(w_n2756_0[0]),.dout(n3014),.clk(gclk));
	jand g02785(.dina(w_n3012_0[0]),.dinb(w_n2759_0[0]),.dout(n3015),.clk(gclk));
	jnot g02786(.din(n3015),.dout(n3016),.clk(gclk));
	jand g02787(.dina(n3016),.dinb(n3014),.dout(n3017),.clk(gclk));
	jnot g02788(.din(n3017),.dout(n3018),.clk(gclk));
	jor g02789(.dina(w_n3018_0[1]),.dinb(w_n3010_0[1]),.dout(n3019),.clk(gclk));
	jand g02790(.dina(n3019),.dinb(w_n3008_0[1]),.dout(n3020),.clk(gclk));
	jor g02791(.dina(w_n3020_0[1]),.dinb(w_n590_28[2]),.dout(n3021),.clk(gclk));
	jxor g02792(.dina(w_n2760_0[0]),.dinb(w_n595_29[2]),.dout(n3022),.clk(gclk));
	jor g02793(.dina(n3022),.dinb(w_n2875_29[2]),.dout(n3023),.clk(gclk));
	jxor g02794(.dina(n3023),.dinb(w_n2771_0[0]),.dout(n3024),.clk(gclk));
	jand g02795(.dina(w_n3020_0[0]),.dinb(w_n590_28[1]),.dout(n3025),.clk(gclk));
	jor g02796(.dina(w_n3025_0[1]),.dinb(w_n3024_0[1]),.dout(n3026),.clk(gclk));
	jand g02797(.dina(w_n3026_0[2]),.dinb(w_n3021_0[2]),.dout(n3027),.clk(gclk));
	jor g02798(.dina(n3027),.dinb(w_n430_30[0]),.dout(n3028),.clk(gclk));
	jnot g02799(.din(w_n2776_0[0]),.dout(n3029),.clk(gclk));
	jor g02800(.dina(n3029),.dinb(w_n2774_0[0]),.dout(n3030),.clk(gclk));
	jor g02801(.dina(n3030),.dinb(w_n2875_29[1]),.dout(n3031),.clk(gclk));
	jxor g02802(.dina(n3031),.dinb(w_n2785_0[0]),.dout(n3032),.clk(gclk));
	jand g02803(.dina(w_n3021_0[1]),.dinb(w_n430_29[2]),.dout(n3033),.clk(gclk));
	jand g02804(.dina(n3033),.dinb(w_n3026_0[1]),.dout(n3034),.clk(gclk));
	jor g02805(.dina(w_n3034_0[1]),.dinb(w_n3032_0[1]),.dout(n3035),.clk(gclk));
	jand g02806(.dina(w_n3035_0[1]),.dinb(w_n3028_0[1]),.dout(n3036),.clk(gclk));
	jor g02807(.dina(w_n3036_0[2]),.dinb(w_n425_29[0]),.dout(n3037),.clk(gclk));
	jand g02808(.dina(w_n3036_0[1]),.dinb(w_n425_28[2]),.dout(n3038),.clk(gclk));
	jnot g02809(.din(w_n2788_0[0]),.dout(n3039),.clk(gclk));
	jand g02810(.dina(w_asqrt41_23[0]),.dinb(n3039),.dout(n3040),.clk(gclk));
	jand g02811(.dina(w_n3040_0[1]),.dinb(w_n2793_0[0]),.dout(n3041),.clk(gclk));
	jor g02812(.dina(n3041),.dinb(w_n2792_0[0]),.dout(n3042),.clk(gclk));
	jand g02813(.dina(w_n3040_0[0]),.dinb(w_n2794_0[0]),.dout(n3043),.clk(gclk));
	jnot g02814(.din(n3043),.dout(n3044),.clk(gclk));
	jand g02815(.dina(n3044),.dinb(n3042),.dout(n3045),.clk(gclk));
	jnot g02816(.din(n3045),.dout(n3046),.clk(gclk));
	jor g02817(.dina(w_n3046_0[1]),.dinb(n3038),.dout(n3047),.clk(gclk));
	jand g02818(.dina(w_n3047_0[1]),.dinb(w_n3037_0[1]),.dout(n3048),.clk(gclk));
	jor g02819(.dina(n3048),.dinb(w_n305_30[2]),.dout(n3049),.clk(gclk));
	jand g02820(.dina(w_n3037_0[0]),.dinb(w_n305_30[1]),.dout(n3050),.clk(gclk));
	jand g02821(.dina(n3050),.dinb(w_n3047_0[0]),.dout(n3051),.clk(gclk));
	jnot g02822(.din(w_n2796_0[0]),.dout(n3052),.clk(gclk));
	jand g02823(.dina(w_asqrt41_22[2]),.dinb(n3052),.dout(n3053),.clk(gclk));
	jand g02824(.dina(w_n3053_0[1]),.dinb(w_n2803_0[0]),.dout(n3054),.clk(gclk));
	jor g02825(.dina(n3054),.dinb(w_n2801_0[0]),.dout(n3055),.clk(gclk));
	jand g02826(.dina(w_n3053_0[0]),.dinb(w_n2804_0[0]),.dout(n3056),.clk(gclk));
	jnot g02827(.din(n3056),.dout(n3057),.clk(gclk));
	jand g02828(.dina(n3057),.dinb(n3055),.dout(n3058),.clk(gclk));
	jnot g02829(.din(n3058),.dout(n3059),.clk(gclk));
	jor g02830(.dina(w_n3059_0[1]),.dinb(w_n3051_0[1]),.dout(n3060),.clk(gclk));
	jand g02831(.dina(n3060),.dinb(w_n3049_0[1]),.dout(n3061),.clk(gclk));
	jor g02832(.dina(w_n3061_0[1]),.dinb(w_n290_30[0]),.dout(n3062),.clk(gclk));
	jxor g02833(.dina(w_n2805_0[0]),.dinb(w_n305_30[0]),.dout(n3063),.clk(gclk));
	jor g02834(.dina(n3063),.dinb(w_n2875_29[0]),.dout(n3064),.clk(gclk));
	jxor g02835(.dina(n3064),.dinb(w_n2816_0[0]),.dout(n3065),.clk(gclk));
	jand g02836(.dina(w_n3061_0[0]),.dinb(w_n290_29[2]),.dout(n3066),.clk(gclk));
	jor g02837(.dina(w_n3066_0[1]),.dinb(w_n3065_0[1]),.dout(n3067),.clk(gclk));
	jand g02838(.dina(w_n3067_0[2]),.dinb(w_n3062_0[2]),.dout(n3068),.clk(gclk));
	jor g02839(.dina(n3068),.dinb(w_n223_30[1]),.dout(n3069),.clk(gclk));
	jnot g02840(.din(w_n2821_0[0]),.dout(n3070),.clk(gclk));
	jor g02841(.dina(n3070),.dinb(w_n2819_0[0]),.dout(n3071),.clk(gclk));
	jor g02842(.dina(n3071),.dinb(w_n2875_28[2]),.dout(n3072),.clk(gclk));
	jxor g02843(.dina(n3072),.dinb(w_n2830_0[0]),.dout(n3073),.clk(gclk));
	jand g02844(.dina(w_n3062_0[1]),.dinb(w_n223_30[0]),.dout(n3074),.clk(gclk));
	jand g02845(.dina(n3074),.dinb(w_n3067_0[1]),.dout(n3075),.clk(gclk));
	jor g02846(.dina(w_n3075_0[1]),.dinb(w_n3073_0[1]),.dout(n3076),.clk(gclk));
	jand g02847(.dina(w_n3076_0[1]),.dinb(w_n3069_0[1]),.dout(n3077),.clk(gclk));
	jor g02848(.dina(w_n3077_0[2]),.dinb(w_n199_35[1]),.dout(n3078),.clk(gclk));
	jand g02849(.dina(w_n3077_0[1]),.dinb(w_n199_35[0]),.dout(n3079),.clk(gclk));
	jnot g02850(.din(w_n2833_0[0]),.dout(n3080),.clk(gclk));
	jand g02851(.dina(w_asqrt41_22[1]),.dinb(n3080),.dout(n3081),.clk(gclk));
	jand g02852(.dina(w_n3081_0[1]),.dinb(w_n2838_0[0]),.dout(n3082),.clk(gclk));
	jor g02853(.dina(n3082),.dinb(w_n2837_0[0]),.dout(n3083),.clk(gclk));
	jand g02854(.dina(w_n3081_0[0]),.dinb(w_n2839_0[0]),.dout(n3084),.clk(gclk));
	jnot g02855(.din(n3084),.dout(n3085),.clk(gclk));
	jand g02856(.dina(n3085),.dinb(n3083),.dout(n3086),.clk(gclk));
	jnot g02857(.din(n3086),.dout(n3087),.clk(gclk));
	jor g02858(.dina(w_n3087_0[1]),.dinb(n3079),.dout(n3088),.clk(gclk));
	jand g02859(.dina(n3088),.dinb(n3078),.dout(n3089),.clk(gclk));
	jnot g02860(.din(w_n2841_0[0]),.dout(n3090),.clk(gclk));
	jand g02861(.dina(w_asqrt41_22[0]),.dinb(n3090),.dout(n3091),.clk(gclk));
	jand g02862(.dina(w_n3091_0[1]),.dinb(w_n2848_0[0]),.dout(n3092),.clk(gclk));
	jor g02863(.dina(n3092),.dinb(w_n2846_0[0]),.dout(n3093),.clk(gclk));
	jand g02864(.dina(w_n3091_0[0]),.dinb(w_n2849_0[0]),.dout(n3094),.clk(gclk));
	jnot g02865(.din(n3094),.dout(n3095),.clk(gclk));
	jand g02866(.dina(n3095),.dinb(n3093),.dout(n3096),.clk(gclk));
	jnot g02867(.din(w_n3096_0[2]),.dout(n3097),.clk(gclk));
	jand g02868(.dina(w_asqrt41_21[2]),.dinb(w_n2863_0[1]),.dout(n3098),.clk(gclk));
	jand g02869(.dina(w_n3098_0[1]),.dinb(w_n2850_1[0]),.dout(n3099),.clk(gclk));
	jor g02870(.dina(n3099),.dinb(w_n2895_0[0]),.dout(n3100),.clk(gclk));
	jor g02871(.dina(n3100),.dinb(w_n3097_0[1]),.dout(n3101),.clk(gclk));
	jor g02872(.dina(n3101),.dinb(w_n3089_0[2]),.dout(n3102),.clk(gclk));
	jand g02873(.dina(n3102),.dinb(w_n194_34[1]),.dout(n3103),.clk(gclk));
	jand g02874(.dina(w_n3097_0[0]),.dinb(w_n3089_0[1]),.dout(n3104),.clk(gclk));
	jor g02875(.dina(w_n3098_0[0]),.dinb(w_n2850_0[2]),.dout(n3105),.clk(gclk));
	jand g02876(.dina(w_n2863_0[0]),.dinb(w_n2850_0[1]),.dout(n3106),.clk(gclk));
	jor g02877(.dina(n3106),.dinb(w_n194_34[0]),.dout(n3107),.clk(gclk));
	jnot g02878(.din(n3107),.dout(n3108),.clk(gclk));
	jand g02879(.dina(n3108),.dinb(n3105),.dout(n3109),.clk(gclk));
	jor g02880(.dina(w_n3109_0[1]),.dinb(w_n3104_0[2]),.dout(n3112),.clk(gclk));
	jor g02881(.dina(n3112),.dinb(w_n3103_0[1]),.dout(asqrt_fa_41),.clk(gclk));
	jand g02882(.dina(w_asqrt40_31),.dinb(w_a80_0[0]),.dout(n3114),.clk(gclk));
	jnot g02883(.din(w_a78_0[1]),.dout(n3115),.clk(gclk));
	jnot g02884(.din(w_a79_0[1]),.dout(n3116),.clk(gclk));
	jand g02885(.dina(w_n2878_1[0]),.dinb(w_n3116_0[1]),.dout(n3117),.clk(gclk));
	jand g02886(.dina(n3117),.dinb(w_n3115_1[1]),.dout(n3118),.clk(gclk));
	jor g02887(.dina(n3118),.dinb(n3114),.dout(n3119),.clk(gclk));
	jand g02888(.dina(w_n3119_0[2]),.dinb(w_asqrt41_21[1]),.dout(n3120),.clk(gclk));
	jand g02889(.dina(w_asqrt40_30[2]),.dinb(w_n2878_0[2]),.dout(n3121),.clk(gclk));
	jxor g02890(.dina(w_n3121_0[1]),.dinb(w_n2879_0[1]),.dout(n3122),.clk(gclk));
	jor g02891(.dina(w_n3119_0[1]),.dinb(w_asqrt41_21[0]),.dout(n3123),.clk(gclk));
	jand g02892(.dina(n3123),.dinb(w_n3122_0[1]),.dout(n3124),.clk(gclk));
	jor g02893(.dina(w_n3124_0[1]),.dinb(w_n3120_0[1]),.dout(n3125),.clk(gclk));
	jand g02894(.dina(n3125),.dinb(w_asqrt42_23[1]),.dout(n3126),.clk(gclk));
	jor g02895(.dina(w_n3120_0[0]),.dinb(w_asqrt42_23[0]),.dout(n3127),.clk(gclk));
	jor g02896(.dina(n3127),.dinb(w_n3124_0[0]),.dout(n3128),.clk(gclk));
	jand g02897(.dina(w_n3121_0[0]),.dinb(w_n2879_0[0]),.dout(n3129),.clk(gclk));
	jnot g02898(.din(w_n3103_0[0]),.dout(n3130),.clk(gclk));
	jnot g02899(.din(w_n3104_0[1]),.dout(n3131),.clk(gclk));
	jnot g02900(.din(w_n3109_0[0]),.dout(n3132),.clk(gclk));
	jand g02901(.dina(n3132),.dinb(w_asqrt41_20[2]),.dout(n3133),.clk(gclk));
	jand g02902(.dina(n3133),.dinb(n3131),.dout(n3134),.clk(gclk));
	jand g02903(.dina(n3134),.dinb(n3130),.dout(n3135),.clk(gclk));
	jor g02904(.dina(n3135),.dinb(n3129),.dout(n3136),.clk(gclk));
	jxor g02905(.dina(n3136),.dinb(w_n2640_0[1]),.dout(n3137),.clk(gclk));
	jand g02906(.dina(w_n3137_0[1]),.dinb(w_n3128_0[1]),.dout(n3138),.clk(gclk));
	jor g02907(.dina(n3138),.dinb(w_n3126_0[1]),.dout(n3139),.clk(gclk));
	jand g02908(.dina(w_n3139_0[2]),.dinb(w_asqrt43_21[0]),.dout(n3140),.clk(gclk));
	jor g02909(.dina(w_n3139_0[1]),.dinb(w_asqrt43_20[2]),.dout(n3141),.clk(gclk));
	jxor g02910(.dina(w_n2883_0[0]),.dinb(w_n2870_25[2]),.dout(n3142),.clk(gclk));
	jand g02911(.dina(n3142),.dinb(w_asqrt40_30[1]),.dout(n3143),.clk(gclk));
	jxor g02912(.dina(n3143),.dinb(w_n2886_0[0]),.dout(n3144),.clk(gclk));
	jnot g02913(.din(w_n3144_0[1]),.dout(n3145),.clk(gclk));
	jand g02914(.dina(n3145),.dinb(n3141),.dout(n3146),.clk(gclk));
	jor g02915(.dina(w_n3146_0[1]),.dinb(w_n3140_0[1]),.dout(n3147),.clk(gclk));
	jand g02916(.dina(n3147),.dinb(w_asqrt44_23[1]),.dout(n3148),.clk(gclk));
	jnot g02917(.din(w_n2892_0[0]),.dout(n3149),.clk(gclk));
	jand g02918(.dina(n3149),.dinb(w_n2890_0[0]),.dout(n3150),.clk(gclk));
	jand g02919(.dina(n3150),.dinb(w_asqrt40_30[0]),.dout(n3151),.clk(gclk));
	jxor g02920(.dina(n3151),.dinb(w_n2900_0[0]),.dout(n3152),.clk(gclk));
	jnot g02921(.din(n3152),.dout(n3153),.clk(gclk));
	jor g02922(.dina(w_n3140_0[0]),.dinb(w_asqrt44_23[0]),.dout(n3154),.clk(gclk));
	jor g02923(.dina(n3154),.dinb(w_n3146_0[0]),.dout(n3155),.clk(gclk));
	jand g02924(.dina(w_n3155_0[1]),.dinb(w_n3153_0[1]),.dout(n3156),.clk(gclk));
	jor g02925(.dina(w_n3156_0[1]),.dinb(w_n3148_0[1]),.dout(n3157),.clk(gclk));
	jand g02926(.dina(w_n3157_0[2]),.dinb(w_asqrt45_21[1]),.dout(n3158),.clk(gclk));
	jor g02927(.dina(w_n3157_0[1]),.dinb(w_asqrt45_21[0]),.dout(n3159),.clk(gclk));
	jnot g02928(.din(w_n2907_0[0]),.dout(n3160),.clk(gclk));
	jxor g02929(.dina(w_n2902_0[0]),.dinb(w_n2420_26[1]),.dout(n3161),.clk(gclk));
	jand g02930(.dina(n3161),.dinb(w_asqrt40_29[2]),.dout(n3162),.clk(gclk));
	jxor g02931(.dina(n3162),.dinb(n3160),.dout(n3163),.clk(gclk));
	jand g02932(.dina(w_n3163_0[1]),.dinb(n3159),.dout(n3164),.clk(gclk));
	jor g02933(.dina(w_n3164_0[1]),.dinb(w_n3158_0[1]),.dout(n3165),.clk(gclk));
	jand g02934(.dina(n3165),.dinb(w_asqrt46_23[1]),.dout(n3166),.clk(gclk));
	jor g02935(.dina(w_n3158_0[0]),.dinb(w_asqrt46_23[0]),.dout(n3167),.clk(gclk));
	jor g02936(.dina(n3167),.dinb(w_n3164_0[0]),.dout(n3168),.clk(gclk));
	jnot g02937(.din(w_n2914_0[0]),.dout(n3169),.clk(gclk));
	jnot g02938(.din(w_n2916_0[0]),.dout(n3170),.clk(gclk));
	jand g02939(.dina(w_asqrt40_29[1]),.dinb(w_n2910_0[0]),.dout(n3171),.clk(gclk));
	jand g02940(.dina(w_n3171_0[1]),.dinb(n3170),.dout(n3172),.clk(gclk));
	jor g02941(.dina(n3172),.dinb(n3169),.dout(n3173),.clk(gclk));
	jnot g02942(.din(w_n2917_0[0]),.dout(n3174),.clk(gclk));
	jand g02943(.dina(w_n3171_0[0]),.dinb(n3174),.dout(n3175),.clk(gclk));
	jnot g02944(.din(n3175),.dout(n3176),.clk(gclk));
	jand g02945(.dina(n3176),.dinb(n3173),.dout(n3177),.clk(gclk));
	jand g02946(.dina(w_n3177_0[1]),.dinb(w_n3168_0[1]),.dout(n3178),.clk(gclk));
	jor g02947(.dina(n3178),.dinb(w_n3166_0[1]),.dout(n3179),.clk(gclk));
	jand g02948(.dina(w_n3179_0[2]),.dinb(w_asqrt47_21[1]),.dout(n3180),.clk(gclk));
	jor g02949(.dina(w_n3179_0[1]),.dinb(w_asqrt47_21[0]),.dout(n3181),.clk(gclk));
	jxor g02950(.dina(w_n2918_0[0]),.dinb(w_n2005_26[1]),.dout(n3182),.clk(gclk));
	jand g02951(.dina(n3182),.dinb(w_asqrt40_29[0]),.dout(n3183),.clk(gclk));
	jxor g02952(.dina(n3183),.dinb(w_n2923_0[0]),.dout(n3184),.clk(gclk));
	jand g02953(.dina(w_n3184_0[1]),.dinb(n3181),.dout(n3185),.clk(gclk));
	jor g02954(.dina(w_n3185_0[1]),.dinb(w_n3180_0[1]),.dout(n3186),.clk(gclk));
	jand g02955(.dina(n3186),.dinb(w_asqrt48_23[1]),.dout(n3187),.clk(gclk));
	jnot g02956(.din(w_n2929_0[0]),.dout(n3188),.clk(gclk));
	jand g02957(.dina(n3188),.dinb(w_n2927_0[0]),.dout(n3189),.clk(gclk));
	jand g02958(.dina(n3189),.dinb(w_asqrt40_28[2]),.dout(n3190),.clk(gclk));
	jxor g02959(.dina(n3190),.dinb(w_n2937_0[0]),.dout(n3191),.clk(gclk));
	jnot g02960(.din(n3191),.dout(n3192),.clk(gclk));
	jor g02961(.dina(w_n3180_0[0]),.dinb(w_asqrt48_23[0]),.dout(n3193),.clk(gclk));
	jor g02962(.dina(n3193),.dinb(w_n3185_0[0]),.dout(n3194),.clk(gclk));
	jand g02963(.dina(w_n3194_0[1]),.dinb(w_n3192_0[1]),.dout(n3195),.clk(gclk));
	jor g02964(.dina(w_n3195_0[1]),.dinb(w_n3187_0[1]),.dout(n3196),.clk(gclk));
	jand g02965(.dina(w_n3196_0[2]),.dinb(w_asqrt49_21[2]),.dout(n3197),.clk(gclk));
	jor g02966(.dina(w_n3196_0[1]),.dinb(w_asqrt49_21[1]),.dout(n3198),.clk(gclk));
	jxor g02967(.dina(w_n2939_0[0]),.dinb(w_n1641_26[2]),.dout(n3199),.clk(gclk));
	jand g02968(.dina(n3199),.dinb(w_asqrt40_28[1]),.dout(n3200),.clk(gclk));
	jxor g02969(.dina(n3200),.dinb(w_n2945_0[0]),.dout(n3201),.clk(gclk));
	jand g02970(.dina(w_n3201_0[1]),.dinb(n3198),.dout(n3202),.clk(gclk));
	jor g02971(.dina(w_n3202_0[1]),.dinb(w_n3197_0[1]),.dout(n3203),.clk(gclk));
	jand g02972(.dina(n3203),.dinb(w_asqrt50_23[1]),.dout(n3204),.clk(gclk));
	jor g02973(.dina(w_n3197_0[0]),.dinb(w_asqrt50_23[0]),.dout(n3205),.clk(gclk));
	jor g02974(.dina(n3205),.dinb(w_n3202_0[0]),.dout(n3206),.clk(gclk));
	jnot g02975(.din(w_n2953_0[0]),.dout(n3207),.clk(gclk));
	jnot g02976(.din(w_n2955_0[0]),.dout(n3208),.clk(gclk));
	jand g02977(.dina(w_asqrt40_28[0]),.dinb(w_n2949_0[0]),.dout(n3209),.clk(gclk));
	jand g02978(.dina(w_n3209_0[1]),.dinb(n3208),.dout(n3210),.clk(gclk));
	jor g02979(.dina(n3210),.dinb(n3207),.dout(n3211),.clk(gclk));
	jnot g02980(.din(w_n2956_0[0]),.dout(n3212),.clk(gclk));
	jand g02981(.dina(w_n3209_0[0]),.dinb(n3212),.dout(n3213),.clk(gclk));
	jnot g02982(.din(n3213),.dout(n3214),.clk(gclk));
	jand g02983(.dina(n3214),.dinb(n3211),.dout(n3215),.clk(gclk));
	jand g02984(.dina(w_n3215_0[1]),.dinb(w_n3206_0[1]),.dout(n3216),.clk(gclk));
	jor g02985(.dina(n3216),.dinb(w_n3204_0[1]),.dout(n3217),.clk(gclk));
	jand g02986(.dina(w_n3217_0[1]),.dinb(w_asqrt51_21[2]),.dout(n3218),.clk(gclk));
	jxor g02987(.dina(w_n2957_0[0]),.dinb(w_n1312_26[2]),.dout(n3219),.clk(gclk));
	jand g02988(.dina(n3219),.dinb(w_asqrt40_27[2]),.dout(n3220),.clk(gclk));
	jxor g02989(.dina(n3220),.dinb(w_n2964_0[0]),.dout(n3221),.clk(gclk));
	jnot g02990(.din(n3221),.dout(n3222),.clk(gclk));
	jor g02991(.dina(w_n3217_0[0]),.dinb(w_asqrt51_21[1]),.dout(n3223),.clk(gclk));
	jand g02992(.dina(w_n3223_0[1]),.dinb(w_n3222_0[1]),.dout(n3224),.clk(gclk));
	jor g02993(.dina(w_n3224_0[2]),.dinb(w_n3218_0[2]),.dout(n3225),.clk(gclk));
	jand g02994(.dina(n3225),.dinb(w_asqrt52_23[1]),.dout(n3226),.clk(gclk));
	jnot g02995(.din(w_n2969_0[0]),.dout(n3227),.clk(gclk));
	jand g02996(.dina(n3227),.dinb(w_n2967_0[0]),.dout(n3228),.clk(gclk));
	jand g02997(.dina(n3228),.dinb(w_asqrt40_27[1]),.dout(n3229),.clk(gclk));
	jxor g02998(.dina(n3229),.dinb(w_n2977_0[0]),.dout(n3230),.clk(gclk));
	jnot g02999(.din(n3230),.dout(n3231),.clk(gclk));
	jor g03000(.dina(w_n3218_0[1]),.dinb(w_asqrt52_23[0]),.dout(n3232),.clk(gclk));
	jor g03001(.dina(n3232),.dinb(w_n3224_0[1]),.dout(n3233),.clk(gclk));
	jand g03002(.dina(w_n3233_0[1]),.dinb(w_n3231_0[1]),.dout(n3234),.clk(gclk));
	jor g03003(.dina(w_n3234_0[1]),.dinb(w_n3226_0[1]),.dout(n3235),.clk(gclk));
	jand g03004(.dina(w_n3235_0[2]),.dinb(w_asqrt53_22[0]),.dout(n3236),.clk(gclk));
	jor g03005(.dina(w_n3235_0[1]),.dinb(w_asqrt53_21[2]),.dout(n3237),.clk(gclk));
	jnot g03006(.din(w_n2983_0[0]),.dout(n3238),.clk(gclk));
	jnot g03007(.din(w_n2984_0[0]),.dout(n3239),.clk(gclk));
	jand g03008(.dina(w_asqrt40_27[0]),.dinb(w_n2980_0[0]),.dout(n3240),.clk(gclk));
	jand g03009(.dina(w_n3240_0[1]),.dinb(n3239),.dout(n3241),.clk(gclk));
	jor g03010(.dina(n3241),.dinb(n3238),.dout(n3242),.clk(gclk));
	jnot g03011(.din(w_n2985_0[0]),.dout(n3243),.clk(gclk));
	jand g03012(.dina(w_n3240_0[0]),.dinb(n3243),.dout(n3244),.clk(gclk));
	jnot g03013(.din(n3244),.dout(n3245),.clk(gclk));
	jand g03014(.dina(n3245),.dinb(n3242),.dout(n3246),.clk(gclk));
	jand g03015(.dina(w_n3246_0[1]),.dinb(n3237),.dout(n3247),.clk(gclk));
	jor g03016(.dina(w_n3247_0[1]),.dinb(w_n3236_0[1]),.dout(n3248),.clk(gclk));
	jand g03017(.dina(n3248),.dinb(w_asqrt54_23[1]),.dout(n3249),.clk(gclk));
	jor g03018(.dina(w_n3236_0[0]),.dinb(w_asqrt54_23[0]),.dout(n3250),.clk(gclk));
	jor g03019(.dina(n3250),.dinb(w_n3247_0[0]),.dout(n3251),.clk(gclk));
	jnot g03020(.din(w_n2991_0[0]),.dout(n3252),.clk(gclk));
	jnot g03021(.din(w_n2993_0[0]),.dout(n3253),.clk(gclk));
	jand g03022(.dina(w_asqrt40_26[2]),.dinb(w_n2987_0[0]),.dout(n3254),.clk(gclk));
	jand g03023(.dina(w_n3254_0[1]),.dinb(n3253),.dout(n3255),.clk(gclk));
	jor g03024(.dina(n3255),.dinb(n3252),.dout(n3256),.clk(gclk));
	jnot g03025(.din(w_n2994_0[0]),.dout(n3257),.clk(gclk));
	jand g03026(.dina(w_n3254_0[0]),.dinb(n3257),.dout(n3258),.clk(gclk));
	jnot g03027(.din(n3258),.dout(n3259),.clk(gclk));
	jand g03028(.dina(n3259),.dinb(n3256),.dout(n3260),.clk(gclk));
	jand g03029(.dina(w_n3260_0[1]),.dinb(w_n3251_0[1]),.dout(n3261),.clk(gclk));
	jor g03030(.dina(n3261),.dinb(w_n3249_0[1]),.dout(n3262),.clk(gclk));
	jand g03031(.dina(w_n3262_0[1]),.dinb(w_asqrt55_22[1]),.dout(n3263),.clk(gclk));
	jxor g03032(.dina(w_n2995_0[0]),.dinb(w_n791_27[2]),.dout(n3264),.clk(gclk));
	jand g03033(.dina(n3264),.dinb(w_asqrt40_26[1]),.dout(n3265),.clk(gclk));
	jxor g03034(.dina(n3265),.dinb(w_n3005_0[0]),.dout(n3266),.clk(gclk));
	jnot g03035(.din(n3266),.dout(n3267),.clk(gclk));
	jor g03036(.dina(w_n3262_0[0]),.dinb(w_asqrt55_22[0]),.dout(n3268),.clk(gclk));
	jand g03037(.dina(w_n3268_0[1]),.dinb(w_n3267_0[1]),.dout(n3269),.clk(gclk));
	jor g03038(.dina(w_n3269_0[2]),.dinb(w_n3263_0[2]),.dout(n3270),.clk(gclk));
	jand g03039(.dina(n3270),.dinb(w_asqrt56_23[1]),.dout(n3271),.clk(gclk));
	jnot g03040(.din(w_n3010_0[0]),.dout(n3272),.clk(gclk));
	jand g03041(.dina(n3272),.dinb(w_n3008_0[0]),.dout(n3273),.clk(gclk));
	jand g03042(.dina(n3273),.dinb(w_asqrt40_26[0]),.dout(n3274),.clk(gclk));
	jxor g03043(.dina(n3274),.dinb(w_n3018_0[0]),.dout(n3275),.clk(gclk));
	jnot g03044(.din(n3275),.dout(n3276),.clk(gclk));
	jor g03045(.dina(w_n3263_0[1]),.dinb(w_asqrt56_23[0]),.dout(n3277),.clk(gclk));
	jor g03046(.dina(n3277),.dinb(w_n3269_0[1]),.dout(n3278),.clk(gclk));
	jand g03047(.dina(w_n3278_0[1]),.dinb(w_n3276_0[1]),.dout(n3279),.clk(gclk));
	jor g03048(.dina(w_n3279_0[1]),.dinb(w_n3271_0[1]),.dout(n3280),.clk(gclk));
	jand g03049(.dina(w_n3280_0[2]),.dinb(w_asqrt57_22[2]),.dout(n3281),.clk(gclk));
	jor g03050(.dina(w_n3280_0[1]),.dinb(w_asqrt57_22[1]),.dout(n3282),.clk(gclk));
	jnot g03051(.din(w_n3024_0[0]),.dout(n3283),.clk(gclk));
	jnot g03052(.din(w_n3025_0[0]),.dout(n3284),.clk(gclk));
	jand g03053(.dina(w_asqrt40_25[2]),.dinb(w_n3021_0[0]),.dout(n3285),.clk(gclk));
	jand g03054(.dina(w_n3285_0[1]),.dinb(n3284),.dout(n3286),.clk(gclk));
	jor g03055(.dina(n3286),.dinb(n3283),.dout(n3287),.clk(gclk));
	jnot g03056(.din(w_n3026_0[0]),.dout(n3288),.clk(gclk));
	jand g03057(.dina(w_n3285_0[0]),.dinb(n3288),.dout(n3289),.clk(gclk));
	jnot g03058(.din(n3289),.dout(n3290),.clk(gclk));
	jand g03059(.dina(n3290),.dinb(n3287),.dout(n3291),.clk(gclk));
	jand g03060(.dina(w_n3291_0[1]),.dinb(n3282),.dout(n3292),.clk(gclk));
	jor g03061(.dina(w_n3292_0[1]),.dinb(w_n3281_0[1]),.dout(n3293),.clk(gclk));
	jand g03062(.dina(n3293),.dinb(w_asqrt58_23[1]),.dout(n3294),.clk(gclk));
	jor g03063(.dina(w_n3281_0[0]),.dinb(w_asqrt58_23[0]),.dout(n3295),.clk(gclk));
	jor g03064(.dina(n3295),.dinb(w_n3292_0[0]),.dout(n3296),.clk(gclk));
	jnot g03065(.din(w_n3032_0[0]),.dout(n3297),.clk(gclk));
	jnot g03066(.din(w_n3034_0[0]),.dout(n3298),.clk(gclk));
	jand g03067(.dina(w_asqrt40_25[1]),.dinb(w_n3028_0[0]),.dout(n3299),.clk(gclk));
	jand g03068(.dina(w_n3299_0[1]),.dinb(n3298),.dout(n3300),.clk(gclk));
	jor g03069(.dina(n3300),.dinb(n3297),.dout(n3301),.clk(gclk));
	jnot g03070(.din(w_n3035_0[0]),.dout(n3302),.clk(gclk));
	jand g03071(.dina(w_n3299_0[0]),.dinb(n3302),.dout(n3303),.clk(gclk));
	jnot g03072(.din(n3303),.dout(n3304),.clk(gclk));
	jand g03073(.dina(n3304),.dinb(n3301),.dout(n3305),.clk(gclk));
	jand g03074(.dina(w_n3305_0[1]),.dinb(w_n3296_0[1]),.dout(n3306),.clk(gclk));
	jor g03075(.dina(n3306),.dinb(w_n3294_0[1]),.dout(n3307),.clk(gclk));
	jand g03076(.dina(w_n3307_0[1]),.dinb(w_asqrt59_23[0]),.dout(n3308),.clk(gclk));
	jxor g03077(.dina(w_n3036_0[0]),.dinb(w_n425_28[1]),.dout(n3309),.clk(gclk));
	jand g03078(.dina(n3309),.dinb(w_asqrt40_25[0]),.dout(n3310),.clk(gclk));
	jxor g03079(.dina(n3310),.dinb(w_n3046_0[0]),.dout(n3311),.clk(gclk));
	jnot g03080(.din(n3311),.dout(n3312),.clk(gclk));
	jor g03081(.dina(w_n3307_0[0]),.dinb(w_asqrt59_22[2]),.dout(n3313),.clk(gclk));
	jand g03082(.dina(w_n3313_0[1]),.dinb(w_n3312_0[1]),.dout(n3314),.clk(gclk));
	jor g03083(.dina(w_n3314_0[2]),.dinb(w_n3308_0[2]),.dout(n3315),.clk(gclk));
	jand g03084(.dina(n3315),.dinb(w_asqrt60_23[0]),.dout(n3316),.clk(gclk));
	jnot g03085(.din(w_n3051_0[0]),.dout(n3317),.clk(gclk));
	jand g03086(.dina(n3317),.dinb(w_n3049_0[0]),.dout(n3318),.clk(gclk));
	jand g03087(.dina(n3318),.dinb(w_asqrt40_24[2]),.dout(n3319),.clk(gclk));
	jxor g03088(.dina(n3319),.dinb(w_n3059_0[0]),.dout(n3320),.clk(gclk));
	jnot g03089(.din(n3320),.dout(n3321),.clk(gclk));
	jor g03090(.dina(w_n3308_0[1]),.dinb(w_asqrt60_22[2]),.dout(n3322),.clk(gclk));
	jor g03091(.dina(n3322),.dinb(w_n3314_0[1]),.dout(n3323),.clk(gclk));
	jand g03092(.dina(w_n3323_0[1]),.dinb(w_n3321_0[1]),.dout(n3324),.clk(gclk));
	jor g03093(.dina(w_n3324_0[1]),.dinb(w_n3316_0[1]),.dout(n3325),.clk(gclk));
	jand g03094(.dina(w_n3325_0[2]),.dinb(w_asqrt61_23[1]),.dout(n3326),.clk(gclk));
	jor g03095(.dina(w_n3325_0[1]),.dinb(w_asqrt61_23[0]),.dout(n3327),.clk(gclk));
	jnot g03096(.din(w_n3065_0[0]),.dout(n3328),.clk(gclk));
	jnot g03097(.din(w_n3066_0[0]),.dout(n3329),.clk(gclk));
	jand g03098(.dina(w_asqrt40_24[1]),.dinb(w_n3062_0[0]),.dout(n3330),.clk(gclk));
	jand g03099(.dina(w_n3330_0[1]),.dinb(n3329),.dout(n3331),.clk(gclk));
	jor g03100(.dina(n3331),.dinb(n3328),.dout(n3332),.clk(gclk));
	jnot g03101(.din(w_n3067_0[0]),.dout(n3333),.clk(gclk));
	jand g03102(.dina(w_n3330_0[0]),.dinb(n3333),.dout(n3334),.clk(gclk));
	jnot g03103(.din(n3334),.dout(n3335),.clk(gclk));
	jand g03104(.dina(n3335),.dinb(n3332),.dout(n3336),.clk(gclk));
	jand g03105(.dina(w_n3336_0[1]),.dinb(n3327),.dout(n3337),.clk(gclk));
	jor g03106(.dina(w_n3337_0[1]),.dinb(w_n3326_0[1]),.dout(n3338),.clk(gclk));
	jand g03107(.dina(n3338),.dinb(w_asqrt62_23[1]),.dout(n3339),.clk(gclk));
	jor g03108(.dina(w_n3326_0[0]),.dinb(w_asqrt62_23[0]),.dout(n3340),.clk(gclk));
	jor g03109(.dina(n3340),.dinb(w_n3337_0[0]),.dout(n3341),.clk(gclk));
	jnot g03110(.din(w_n3073_0[0]),.dout(n3342),.clk(gclk));
	jnot g03111(.din(w_n3075_0[0]),.dout(n3343),.clk(gclk));
	jand g03112(.dina(w_asqrt40_24[0]),.dinb(w_n3069_0[0]),.dout(n3344),.clk(gclk));
	jand g03113(.dina(w_n3344_0[1]),.dinb(n3343),.dout(n3345),.clk(gclk));
	jor g03114(.dina(n3345),.dinb(n3342),.dout(n3346),.clk(gclk));
	jnot g03115(.din(w_n3076_0[0]),.dout(n3347),.clk(gclk));
	jand g03116(.dina(w_n3344_0[0]),.dinb(n3347),.dout(n3348),.clk(gclk));
	jnot g03117(.din(n3348),.dout(n3349),.clk(gclk));
	jand g03118(.dina(n3349),.dinb(n3346),.dout(n3350),.clk(gclk));
	jand g03119(.dina(w_n3350_0[1]),.dinb(w_n3341_0[1]),.dout(n3351),.clk(gclk));
	jor g03120(.dina(n3351),.dinb(w_n3339_0[1]),.dout(n3352),.clk(gclk));
	jxor g03121(.dina(w_n3077_0[0]),.dinb(w_n199_34[2]),.dout(n3353),.clk(gclk));
	jand g03122(.dina(n3353),.dinb(w_asqrt40_23[2]),.dout(n3354),.clk(gclk));
	jxor g03123(.dina(n3354),.dinb(w_n3087_0[0]),.dout(n3355),.clk(gclk));
	jnot g03124(.din(w_n3089_0[0]),.dout(n3356),.clk(gclk));
	jand g03125(.dina(w_asqrt40_23[1]),.dinb(w_n3096_0[1]),.dout(n3357),.clk(gclk));
	jand g03126(.dina(w_n3357_0[1]),.dinb(w_n3356_0[2]),.dout(n3358),.clk(gclk));
	jor g03127(.dina(n3358),.dinb(w_n3104_0[0]),.dout(n3359),.clk(gclk));
	jor g03128(.dina(n3359),.dinb(w_n3355_0[1]),.dout(n3360),.clk(gclk));
	jnot g03129(.din(n3360),.dout(n3361),.clk(gclk));
	jand g03130(.dina(n3361),.dinb(w_n3352_1[2]),.dout(n3362),.clk(gclk));
	jor g03131(.dina(n3362),.dinb(w_asqrt63_12[1]),.dout(n3363),.clk(gclk));
	jnot g03132(.din(w_n3355_0[0]),.dout(n3364),.clk(gclk));
	jor g03133(.dina(w_n3364_0[2]),.dinb(w_n3352_1[1]),.dout(n3365),.clk(gclk));
	jor g03134(.dina(w_n3357_0[0]),.dinb(w_n3356_0[1]),.dout(n3366),.clk(gclk));
	jand g03135(.dina(w_n3096_0[0]),.dinb(w_n3356_0[0]),.dout(n3367),.clk(gclk));
	jor g03136(.dina(n3367),.dinb(w_n194_33[2]),.dout(n3368),.clk(gclk));
	jnot g03137(.din(n3368),.dout(n3369),.clk(gclk));
	jand g03138(.dina(n3369),.dinb(n3366),.dout(n3370),.clk(gclk));
	jnot g03139(.din(w_asqrt40_23[0]),.dout(n3371),.clk(gclk));
	jnot g03140(.din(w_n3370_0[1]),.dout(n3374),.clk(gclk));
	jand g03141(.dina(n3374),.dinb(w_n3365_0[1]),.dout(n3375),.clk(gclk));
	jand g03142(.dina(n3375),.dinb(w_n3363_0[1]),.dout(n3376),.clk(gclk));
	jnot g03143(.din(w_n3376_33[1]),.dout(asqrt_fa_40),.clk(gclk));
	jor g03144(.dina(w_n3376_33[0]),.dinb(w_n3115_1[0]),.dout(n3378),.clk(gclk));
	jnot g03145(.din(w_a76_0[1]),.dout(n3379),.clk(gclk));
	jnot g03146(.din(a[77]),.dout(n3380),.clk(gclk));
	jand g03147(.dina(w_n3115_0[2]),.dinb(w_n3380_0[2]),.dout(n3381),.clk(gclk));
	jand g03148(.dina(n3381),.dinb(w_n3379_1[1]),.dout(n3382),.clk(gclk));
	jnot g03149(.din(n3382),.dout(n3383),.clk(gclk));
	jand g03150(.dina(n3383),.dinb(n3378),.dout(n3384),.clk(gclk));
	jor g03151(.dina(w_n3384_0[2]),.dinb(w_n3371_25[2]),.dout(n3385),.clk(gclk));
	jor g03152(.dina(w_n3376_32[2]),.dinb(w_a78_0[0]),.dout(n3386),.clk(gclk));
	jxor g03153(.dina(w_n3386_0[1]),.dinb(w_n3116_0[0]),.dout(n3387),.clk(gclk));
	jand g03154(.dina(w_n3384_0[1]),.dinb(w_n3371_25[1]),.dout(n3388),.clk(gclk));
	jor g03155(.dina(n3388),.dinb(w_n3387_0[1]),.dout(n3389),.clk(gclk));
	jand g03156(.dina(w_n3389_0[1]),.dinb(w_n3385_0[1]),.dout(n3390),.clk(gclk));
	jor g03157(.dina(n3390),.dinb(w_n2875_28[1]),.dout(n3391),.clk(gclk));
	jand g03158(.dina(w_n3385_0[0]),.dinb(w_n2875_28[0]),.dout(n3392),.clk(gclk));
	jand g03159(.dina(n3392),.dinb(w_n3389_0[0]),.dout(n3393),.clk(gclk));
	jor g03160(.dina(w_n3386_0[0]),.dinb(w_a79_0[0]),.dout(n3394),.clk(gclk));
	jnot g03161(.din(w_n3363_0[0]),.dout(n3395),.clk(gclk));
	jnot g03162(.din(w_n3365_0[0]),.dout(n3396),.clk(gclk));
	jor g03163(.dina(w_n3370_0[0]),.dinb(w_n3371_25[0]),.dout(n3397),.clk(gclk));
	jor g03164(.dina(n3397),.dinb(w_n3396_0[1]),.dout(n3398),.clk(gclk));
	jor g03165(.dina(n3398),.dinb(n3395),.dout(n3399),.clk(gclk));
	jand g03166(.dina(n3399),.dinb(n3394),.dout(n3400),.clk(gclk));
	jxor g03167(.dina(n3400),.dinb(w_n2878_0[1]),.dout(n3401),.clk(gclk));
	jor g03168(.dina(w_n3401_0[1]),.dinb(w_n3393_0[1]),.dout(n3402),.clk(gclk));
	jand g03169(.dina(n3402),.dinb(w_n3391_0[1]),.dout(n3403),.clk(gclk));
	jor g03170(.dina(w_n3403_0[2]),.dinb(w_n2870_25[1]),.dout(n3404),.clk(gclk));
	jand g03171(.dina(w_n3403_0[1]),.dinb(w_n2870_25[0]),.dout(n3405),.clk(gclk));
	jxor g03172(.dina(w_n3119_0[0]),.dinb(w_n2875_27[2]),.dout(n3406),.clk(gclk));
	jor g03173(.dina(n3406),.dinb(w_n3376_32[1]),.dout(n3407),.clk(gclk));
	jxor g03174(.dina(n3407),.dinb(w_n3122_0[0]),.dout(n3408),.clk(gclk));
	jor g03175(.dina(w_n3408_0[1]),.dinb(n3405),.dout(n3409),.clk(gclk));
	jand g03176(.dina(w_n3409_0[1]),.dinb(w_n3404_0[1]),.dout(n3410),.clk(gclk));
	jor g03177(.dina(n3410),.dinb(w_n2425_28[2]),.dout(n3411),.clk(gclk));
	jnot g03178(.din(w_n3128_0[0]),.dout(n3412),.clk(gclk));
	jor g03179(.dina(n3412),.dinb(w_n3126_0[0]),.dout(n3413),.clk(gclk));
	jor g03180(.dina(n3413),.dinb(w_n3376_32[0]),.dout(n3414),.clk(gclk));
	jxor g03181(.dina(n3414),.dinb(w_n3137_0[0]),.dout(n3415),.clk(gclk));
	jand g03182(.dina(w_n3404_0[0]),.dinb(w_n2425_28[1]),.dout(n3416),.clk(gclk));
	jand g03183(.dina(n3416),.dinb(w_n3409_0[0]),.dout(n3417),.clk(gclk));
	jor g03184(.dina(w_n3417_0[1]),.dinb(w_n3415_0[1]),.dout(n3418),.clk(gclk));
	jand g03185(.dina(w_n3418_0[1]),.dinb(w_n3411_0[1]),.dout(n3419),.clk(gclk));
	jor g03186(.dina(w_n3419_0[2]),.dinb(w_n2420_26[0]),.dout(n3420),.clk(gclk));
	jand g03187(.dina(w_n3419_0[1]),.dinb(w_n2420_25[2]),.dout(n3421),.clk(gclk));
	jxor g03188(.dina(w_n3139_0[0]),.dinb(w_n2425_28[0]),.dout(n3422),.clk(gclk));
	jor g03189(.dina(n3422),.dinb(w_n3376_31[2]),.dout(n3423),.clk(gclk));
	jxor g03190(.dina(n3423),.dinb(w_n3144_0[0]),.dout(n3424),.clk(gclk));
	jnot g03191(.din(w_n3424_0[1]),.dout(n3425),.clk(gclk));
	jor g03192(.dina(n3425),.dinb(n3421),.dout(n3426),.clk(gclk));
	jand g03193(.dina(w_n3426_0[1]),.dinb(w_n3420_0[1]),.dout(n3427),.clk(gclk));
	jor g03194(.dina(n3427),.dinb(w_n2010_28[1]),.dout(n3428),.clk(gclk));
	jand g03195(.dina(w_n3420_0[0]),.dinb(w_n2010_28[0]),.dout(n3429),.clk(gclk));
	jand g03196(.dina(n3429),.dinb(w_n3426_0[0]),.dout(n3430),.clk(gclk));
	jnot g03197(.din(w_n3148_0[0]),.dout(n3431),.clk(gclk));
	jand g03198(.dina(w_asqrt39_23[1]),.dinb(n3431),.dout(n3432),.clk(gclk));
	jand g03199(.dina(w_n3432_0[1]),.dinb(w_n3155_0[0]),.dout(n3433),.clk(gclk));
	jor g03200(.dina(n3433),.dinb(w_n3153_0[0]),.dout(n3434),.clk(gclk));
	jand g03201(.dina(w_n3432_0[0]),.dinb(w_n3156_0[0]),.dout(n3435),.clk(gclk));
	jnot g03202(.din(n3435),.dout(n3436),.clk(gclk));
	jand g03203(.dina(n3436),.dinb(n3434),.dout(n3437),.clk(gclk));
	jnot g03204(.din(n3437),.dout(n3438),.clk(gclk));
	jor g03205(.dina(w_n3438_0[1]),.dinb(w_n3430_0[1]),.dout(n3439),.clk(gclk));
	jand g03206(.dina(n3439),.dinb(w_n3428_0[1]),.dout(n3440),.clk(gclk));
	jor g03207(.dina(w_n3440_0[2]),.dinb(w_n2005_26[0]),.dout(n3441),.clk(gclk));
	jand g03208(.dina(w_n3440_0[1]),.dinb(w_n2005_25[2]),.dout(n3442),.clk(gclk));
	jnot g03209(.din(w_n3163_0[0]),.dout(n3443),.clk(gclk));
	jxor g03210(.dina(w_n3157_0[0]),.dinb(w_n2010_27[2]),.dout(n3444),.clk(gclk));
	jor g03211(.dina(n3444),.dinb(w_n3376_31[1]),.dout(n3445),.clk(gclk));
	jxor g03212(.dina(n3445),.dinb(n3443),.dout(n3446),.clk(gclk));
	jnot g03213(.din(w_n3446_0[1]),.dout(n3447),.clk(gclk));
	jor g03214(.dina(n3447),.dinb(n3442),.dout(n3448),.clk(gclk));
	jand g03215(.dina(w_n3448_0[1]),.dinb(w_n3441_0[1]),.dout(n3449),.clk(gclk));
	jor g03216(.dina(n3449),.dinb(w_n1646_29[0]),.dout(n3450),.clk(gclk));
	jnot g03217(.din(w_n3168_0[0]),.dout(n3451),.clk(gclk));
	jor g03218(.dina(n3451),.dinb(w_n3166_0[0]),.dout(n3452),.clk(gclk));
	jor g03219(.dina(n3452),.dinb(w_n3376_31[0]),.dout(n3453),.clk(gclk));
	jxor g03220(.dina(n3453),.dinb(w_n3177_0[0]),.dout(n3454),.clk(gclk));
	jand g03221(.dina(w_n3441_0[0]),.dinb(w_n1646_28[2]),.dout(n3455),.clk(gclk));
	jand g03222(.dina(n3455),.dinb(w_n3448_0[0]),.dout(n3456),.clk(gclk));
	jor g03223(.dina(w_n3456_0[1]),.dinb(w_n3454_0[1]),.dout(n3457),.clk(gclk));
	jand g03224(.dina(w_n3457_0[1]),.dinb(w_n3450_0[1]),.dout(n3458),.clk(gclk));
	jor g03225(.dina(w_n3458_0[2]),.dinb(w_n1641_26[1]),.dout(n3459),.clk(gclk));
	jand g03226(.dina(w_n3458_0[1]),.dinb(w_n1641_26[0]),.dout(n3460),.clk(gclk));
	jnot g03227(.din(w_n3184_0[0]),.dout(n3461),.clk(gclk));
	jxor g03228(.dina(w_n3179_0[0]),.dinb(w_n1646_28[1]),.dout(n3462),.clk(gclk));
	jor g03229(.dina(n3462),.dinb(w_n3376_30[2]),.dout(n3463),.clk(gclk));
	jxor g03230(.dina(n3463),.dinb(n3461),.dout(n3464),.clk(gclk));
	jnot g03231(.din(n3464),.dout(n3465),.clk(gclk));
	jor g03232(.dina(w_n3465_0[1]),.dinb(n3460),.dout(n3466),.clk(gclk));
	jand g03233(.dina(w_n3466_0[1]),.dinb(w_n3459_0[1]),.dout(n3467),.clk(gclk));
	jor g03234(.dina(n3467),.dinb(w_n1317_28[2]),.dout(n3468),.clk(gclk));
	jand g03235(.dina(w_n3459_0[0]),.dinb(w_n1317_28[1]),.dout(n3469),.clk(gclk));
	jand g03236(.dina(n3469),.dinb(w_n3466_0[0]),.dout(n3470),.clk(gclk));
	jnot g03237(.din(w_n3187_0[0]),.dout(n3471),.clk(gclk));
	jand g03238(.dina(w_asqrt39_23[0]),.dinb(n3471),.dout(n3472),.clk(gclk));
	jand g03239(.dina(w_n3472_0[1]),.dinb(w_n3194_0[0]),.dout(n3473),.clk(gclk));
	jor g03240(.dina(n3473),.dinb(w_n3192_0[0]),.dout(n3474),.clk(gclk));
	jand g03241(.dina(w_n3472_0[0]),.dinb(w_n3195_0[0]),.dout(n3475),.clk(gclk));
	jnot g03242(.din(n3475),.dout(n3476),.clk(gclk));
	jand g03243(.dina(n3476),.dinb(n3474),.dout(n3477),.clk(gclk));
	jnot g03244(.din(n3477),.dout(n3478),.clk(gclk));
	jor g03245(.dina(w_n3478_0[1]),.dinb(w_n3470_0[1]),.dout(n3479),.clk(gclk));
	jand g03246(.dina(n3479),.dinb(w_n3468_0[1]),.dout(n3480),.clk(gclk));
	jor g03247(.dina(w_n3480_0[1]),.dinb(w_n1312_26[1]),.dout(n3481),.clk(gclk));
	jxor g03248(.dina(w_n3196_0[0]),.dinb(w_n1317_28[0]),.dout(n3482),.clk(gclk));
	jor g03249(.dina(n3482),.dinb(w_n3376_30[1]),.dout(n3483),.clk(gclk));
	jxor g03250(.dina(n3483),.dinb(w_n3201_0[0]),.dout(n3484),.clk(gclk));
	jand g03251(.dina(w_n3480_0[0]),.dinb(w_n1312_26[0]),.dout(n3485),.clk(gclk));
	jor g03252(.dina(w_n3485_0[1]),.dinb(w_n3484_0[1]),.dout(n3486),.clk(gclk));
	jand g03253(.dina(w_n3486_0[2]),.dinb(w_n3481_0[2]),.dout(n3487),.clk(gclk));
	jor g03254(.dina(n3487),.dinb(w_n1039_29[0]),.dout(n3488),.clk(gclk));
	jnot g03255(.din(w_n3206_0[0]),.dout(n3489),.clk(gclk));
	jor g03256(.dina(n3489),.dinb(w_n3204_0[0]),.dout(n3490),.clk(gclk));
	jor g03257(.dina(n3490),.dinb(w_n3376_30[0]),.dout(n3491),.clk(gclk));
	jxor g03258(.dina(n3491),.dinb(w_n3215_0[0]),.dout(n3492),.clk(gclk));
	jand g03259(.dina(w_n3481_0[1]),.dinb(w_n1039_28[2]),.dout(n3493),.clk(gclk));
	jand g03260(.dina(n3493),.dinb(w_n3486_0[1]),.dout(n3494),.clk(gclk));
	jor g03261(.dina(w_n3494_0[1]),.dinb(w_n3492_0[1]),.dout(n3495),.clk(gclk));
	jand g03262(.dina(w_n3495_0[1]),.dinb(w_n3488_0[1]),.dout(n3496),.clk(gclk));
	jor g03263(.dina(w_n3496_0[2]),.dinb(w_n1034_27[1]),.dout(n3497),.clk(gclk));
	jand g03264(.dina(w_n3496_0[1]),.dinb(w_n1034_27[0]),.dout(n3498),.clk(gclk));
	jnot g03265(.din(w_n3218_0[0]),.dout(n3499),.clk(gclk));
	jand g03266(.dina(w_asqrt39_22[2]),.dinb(n3499),.dout(n3500),.clk(gclk));
	jand g03267(.dina(w_n3500_0[1]),.dinb(w_n3223_0[0]),.dout(n3501),.clk(gclk));
	jor g03268(.dina(n3501),.dinb(w_n3222_0[0]),.dout(n3502),.clk(gclk));
	jand g03269(.dina(w_n3500_0[0]),.dinb(w_n3224_0[0]),.dout(n3503),.clk(gclk));
	jnot g03270(.din(n3503),.dout(n3504),.clk(gclk));
	jand g03271(.dina(n3504),.dinb(n3502),.dout(n3505),.clk(gclk));
	jnot g03272(.din(n3505),.dout(n3506),.clk(gclk));
	jor g03273(.dina(w_n3506_0[1]),.dinb(n3498),.dout(n3507),.clk(gclk));
	jand g03274(.dina(w_n3507_0[1]),.dinb(w_n3497_0[1]),.dout(n3508),.clk(gclk));
	jor g03275(.dina(n3508),.dinb(w_n796_29[0]),.dout(n3509),.clk(gclk));
	jand g03276(.dina(w_n3497_0[0]),.dinb(w_n796_28[2]),.dout(n3510),.clk(gclk));
	jand g03277(.dina(n3510),.dinb(w_n3507_0[0]),.dout(n3511),.clk(gclk));
	jnot g03278(.din(w_n3226_0[0]),.dout(n3512),.clk(gclk));
	jand g03279(.dina(w_asqrt39_22[1]),.dinb(n3512),.dout(n3513),.clk(gclk));
	jand g03280(.dina(w_n3513_0[1]),.dinb(w_n3233_0[0]),.dout(n3514),.clk(gclk));
	jor g03281(.dina(n3514),.dinb(w_n3231_0[0]),.dout(n3515),.clk(gclk));
	jand g03282(.dina(w_n3513_0[0]),.dinb(w_n3234_0[0]),.dout(n3516),.clk(gclk));
	jnot g03283(.din(n3516),.dout(n3517),.clk(gclk));
	jand g03284(.dina(n3517),.dinb(n3515),.dout(n3518),.clk(gclk));
	jnot g03285(.din(n3518),.dout(n3519),.clk(gclk));
	jor g03286(.dina(w_n3519_0[1]),.dinb(w_n3511_0[1]),.dout(n3520),.clk(gclk));
	jand g03287(.dina(n3520),.dinb(w_n3509_0[1]),.dout(n3521),.clk(gclk));
	jor g03288(.dina(w_n3521_0[1]),.dinb(w_n791_27[1]),.dout(n3522),.clk(gclk));
	jxor g03289(.dina(w_n3235_0[0]),.dinb(w_n796_28[1]),.dout(n3523),.clk(gclk));
	jor g03290(.dina(n3523),.dinb(w_n3376_29[2]),.dout(n3524),.clk(gclk));
	jxor g03291(.dina(n3524),.dinb(w_n3246_0[0]),.dout(n3525),.clk(gclk));
	jand g03292(.dina(w_n3521_0[0]),.dinb(w_n791_27[0]),.dout(n3526),.clk(gclk));
	jor g03293(.dina(w_n3526_0[1]),.dinb(w_n3525_0[1]),.dout(n3527),.clk(gclk));
	jand g03294(.dina(w_n3527_0[2]),.dinb(w_n3522_0[2]),.dout(n3528),.clk(gclk));
	jor g03295(.dina(n3528),.dinb(w_n595_29[1]),.dout(n3529),.clk(gclk));
	jnot g03296(.din(w_n3251_0[0]),.dout(n3530),.clk(gclk));
	jor g03297(.dina(n3530),.dinb(w_n3249_0[0]),.dout(n3531),.clk(gclk));
	jor g03298(.dina(n3531),.dinb(w_n3376_29[1]),.dout(n3532),.clk(gclk));
	jxor g03299(.dina(n3532),.dinb(w_n3260_0[0]),.dout(n3533),.clk(gclk));
	jand g03300(.dina(w_n3522_0[1]),.dinb(w_n595_29[0]),.dout(n3534),.clk(gclk));
	jand g03301(.dina(n3534),.dinb(w_n3527_0[1]),.dout(n3535),.clk(gclk));
	jor g03302(.dina(w_n3535_0[1]),.dinb(w_n3533_0[1]),.dout(n3536),.clk(gclk));
	jand g03303(.dina(w_n3536_0[1]),.dinb(w_n3529_0[1]),.dout(n3537),.clk(gclk));
	jor g03304(.dina(w_n3537_0[2]),.dinb(w_n590_28[0]),.dout(n3538),.clk(gclk));
	jand g03305(.dina(w_n3537_0[1]),.dinb(w_n590_27[2]),.dout(n3539),.clk(gclk));
	jnot g03306(.din(w_n3263_0[0]),.dout(n3540),.clk(gclk));
	jand g03307(.dina(w_asqrt39_22[0]),.dinb(n3540),.dout(n3541),.clk(gclk));
	jand g03308(.dina(w_n3541_0[1]),.dinb(w_n3268_0[0]),.dout(n3542),.clk(gclk));
	jor g03309(.dina(n3542),.dinb(w_n3267_0[0]),.dout(n3543),.clk(gclk));
	jand g03310(.dina(w_n3541_0[0]),.dinb(w_n3269_0[0]),.dout(n3544),.clk(gclk));
	jnot g03311(.din(n3544),.dout(n3545),.clk(gclk));
	jand g03312(.dina(n3545),.dinb(n3543),.dout(n3546),.clk(gclk));
	jnot g03313(.din(n3546),.dout(n3547),.clk(gclk));
	jor g03314(.dina(w_n3547_0[1]),.dinb(n3539),.dout(n3548),.clk(gclk));
	jand g03315(.dina(w_n3548_0[1]),.dinb(w_n3538_0[1]),.dout(n3549),.clk(gclk));
	jor g03316(.dina(n3549),.dinb(w_n430_29[1]),.dout(n3550),.clk(gclk));
	jand g03317(.dina(w_n3538_0[0]),.dinb(w_n430_29[0]),.dout(n3551),.clk(gclk));
	jand g03318(.dina(n3551),.dinb(w_n3548_0[0]),.dout(n3552),.clk(gclk));
	jnot g03319(.din(w_n3271_0[0]),.dout(n3553),.clk(gclk));
	jand g03320(.dina(w_asqrt39_21[2]),.dinb(n3553),.dout(n3554),.clk(gclk));
	jand g03321(.dina(w_n3554_0[1]),.dinb(w_n3278_0[0]),.dout(n3555),.clk(gclk));
	jor g03322(.dina(n3555),.dinb(w_n3276_0[0]),.dout(n3556),.clk(gclk));
	jand g03323(.dina(w_n3554_0[0]),.dinb(w_n3279_0[0]),.dout(n3557),.clk(gclk));
	jnot g03324(.din(n3557),.dout(n3558),.clk(gclk));
	jand g03325(.dina(n3558),.dinb(n3556),.dout(n3559),.clk(gclk));
	jnot g03326(.din(n3559),.dout(n3560),.clk(gclk));
	jor g03327(.dina(w_n3560_0[1]),.dinb(w_n3552_0[1]),.dout(n3561),.clk(gclk));
	jand g03328(.dina(n3561),.dinb(w_n3550_0[1]),.dout(n3562),.clk(gclk));
	jor g03329(.dina(w_n3562_0[1]),.dinb(w_n425_28[0]),.dout(n3563),.clk(gclk));
	jxor g03330(.dina(w_n3280_0[0]),.dinb(w_n430_28[2]),.dout(n3564),.clk(gclk));
	jor g03331(.dina(n3564),.dinb(w_n3376_29[0]),.dout(n3565),.clk(gclk));
	jxor g03332(.dina(n3565),.dinb(w_n3291_0[0]),.dout(n3566),.clk(gclk));
	jand g03333(.dina(w_n3562_0[0]),.dinb(w_n425_27[2]),.dout(n3567),.clk(gclk));
	jor g03334(.dina(w_n3567_0[1]),.dinb(w_n3566_0[1]),.dout(n3568),.clk(gclk));
	jand g03335(.dina(w_n3568_0[2]),.dinb(w_n3563_0[2]),.dout(n3569),.clk(gclk));
	jor g03336(.dina(n3569),.dinb(w_n305_29[2]),.dout(n3570),.clk(gclk));
	jnot g03337(.din(w_n3296_0[0]),.dout(n3571),.clk(gclk));
	jor g03338(.dina(n3571),.dinb(w_n3294_0[0]),.dout(n3572),.clk(gclk));
	jor g03339(.dina(n3572),.dinb(w_n3376_28[2]),.dout(n3573),.clk(gclk));
	jxor g03340(.dina(n3573),.dinb(w_n3305_0[0]),.dout(n3574),.clk(gclk));
	jand g03341(.dina(w_n3563_0[1]),.dinb(w_n305_29[1]),.dout(n3575),.clk(gclk));
	jand g03342(.dina(n3575),.dinb(w_n3568_0[1]),.dout(n3576),.clk(gclk));
	jor g03343(.dina(w_n3576_0[1]),.dinb(w_n3574_0[1]),.dout(n3577),.clk(gclk));
	jand g03344(.dina(w_n3577_0[1]),.dinb(w_n3570_0[1]),.dout(n3578),.clk(gclk));
	jor g03345(.dina(w_n3578_0[2]),.dinb(w_n290_29[1]),.dout(n3579),.clk(gclk));
	jand g03346(.dina(w_n3578_0[1]),.dinb(w_n290_29[0]),.dout(n3580),.clk(gclk));
	jnot g03347(.din(w_n3308_0[0]),.dout(n3581),.clk(gclk));
	jand g03348(.dina(w_asqrt39_21[1]),.dinb(n3581),.dout(n3582),.clk(gclk));
	jand g03349(.dina(w_n3582_0[1]),.dinb(w_n3313_0[0]),.dout(n3583),.clk(gclk));
	jor g03350(.dina(n3583),.dinb(w_n3312_0[0]),.dout(n3584),.clk(gclk));
	jand g03351(.dina(w_n3582_0[0]),.dinb(w_n3314_0[0]),.dout(n3585),.clk(gclk));
	jnot g03352(.din(n3585),.dout(n3586),.clk(gclk));
	jand g03353(.dina(n3586),.dinb(n3584),.dout(n3587),.clk(gclk));
	jnot g03354(.din(n3587),.dout(n3588),.clk(gclk));
	jor g03355(.dina(w_n3588_0[1]),.dinb(n3580),.dout(n3589),.clk(gclk));
	jand g03356(.dina(w_n3589_0[1]),.dinb(w_n3579_0[1]),.dout(n3590),.clk(gclk));
	jor g03357(.dina(n3590),.dinb(w_n223_29[2]),.dout(n3591),.clk(gclk));
	jand g03358(.dina(w_n3579_0[0]),.dinb(w_n223_29[1]),.dout(n3592),.clk(gclk));
	jand g03359(.dina(n3592),.dinb(w_n3589_0[0]),.dout(n3593),.clk(gclk));
	jnot g03360(.din(w_n3316_0[0]),.dout(n3594),.clk(gclk));
	jand g03361(.dina(w_asqrt39_21[0]),.dinb(n3594),.dout(n3595),.clk(gclk));
	jand g03362(.dina(w_n3595_0[1]),.dinb(w_n3323_0[0]),.dout(n3596),.clk(gclk));
	jor g03363(.dina(n3596),.dinb(w_n3321_0[0]),.dout(n3597),.clk(gclk));
	jand g03364(.dina(w_n3595_0[0]),.dinb(w_n3324_0[0]),.dout(n3598),.clk(gclk));
	jnot g03365(.din(n3598),.dout(n3599),.clk(gclk));
	jand g03366(.dina(n3599),.dinb(n3597),.dout(n3600),.clk(gclk));
	jnot g03367(.din(n3600),.dout(n3601),.clk(gclk));
	jor g03368(.dina(w_n3601_0[1]),.dinb(w_n3593_0[1]),.dout(n3602),.clk(gclk));
	jand g03369(.dina(n3602),.dinb(w_n3591_0[1]),.dout(n3603),.clk(gclk));
	jor g03370(.dina(w_n3603_0[2]),.dinb(w_n199_34[1]),.dout(n3604),.clk(gclk));
	jand g03371(.dina(w_n3603_0[1]),.dinb(w_n199_34[0]),.dout(n3605),.clk(gclk));
	jxor g03372(.dina(w_n3325_0[0]),.dinb(w_n223_29[0]),.dout(n3606),.clk(gclk));
	jor g03373(.dina(n3606),.dinb(w_n3376_28[1]),.dout(n3607),.clk(gclk));
	jxor g03374(.dina(n3607),.dinb(w_n3336_0[0]),.dout(n3608),.clk(gclk));
	jor g03375(.dina(w_n3608_0[1]),.dinb(n3605),.dout(n3609),.clk(gclk));
	jand g03376(.dina(n3609),.dinb(n3604),.dout(n3610),.clk(gclk));
	jnot g03377(.din(w_n3341_0[0]),.dout(n3611),.clk(gclk));
	jor g03378(.dina(n3611),.dinb(w_n3339_0[0]),.dout(n3612),.clk(gclk));
	jor g03379(.dina(n3612),.dinb(w_n3376_28[0]),.dout(n3613),.clk(gclk));
	jxor g03380(.dina(n3613),.dinb(w_n3350_0[0]),.dout(n3614),.clk(gclk));
	jand g03381(.dina(w_asqrt39_20[2]),.dinb(w_n3364_0[1]),.dout(n3615),.clk(gclk));
	jand g03382(.dina(w_n3615_0[1]),.dinb(w_n3352_1[0]),.dout(n3616),.clk(gclk));
	jor g03383(.dina(n3616),.dinb(w_n3396_0[0]),.dout(n3617),.clk(gclk));
	jor g03384(.dina(n3617),.dinb(w_n3614_0[2]),.dout(n3618),.clk(gclk));
	jor g03385(.dina(n3618),.dinb(w_n3610_0[2]),.dout(n3619),.clk(gclk));
	jand g03386(.dina(n3619),.dinb(w_n194_33[1]),.dout(n3620),.clk(gclk));
	jand g03387(.dina(w_n3614_0[1]),.dinb(w_n3610_0[1]),.dout(n3621),.clk(gclk));
	jor g03388(.dina(w_n3615_0[0]),.dinb(w_n3352_0[2]),.dout(n3622),.clk(gclk));
	jand g03389(.dina(w_n3364_0[0]),.dinb(w_n3352_0[1]),.dout(n3623),.clk(gclk));
	jor g03390(.dina(n3623),.dinb(w_n194_33[0]),.dout(n3624),.clk(gclk));
	jnot g03391(.din(n3624),.dout(n3625),.clk(gclk));
	jand g03392(.dina(n3625),.dinb(n3622),.dout(n3626),.clk(gclk));
	jor g03393(.dina(w_n3626_0[1]),.dinb(w_n3621_0[2]),.dout(n3629),.clk(gclk));
	jor g03394(.dina(n3629),.dinb(w_n3620_0[1]),.dout(asqrt_fa_39),.clk(gclk));
	jand g03395(.dina(w_asqrt38_31),.dinb(w_a76_0[0]),.dout(n3631),.clk(gclk));
	jnot g03396(.din(w_a74_0[1]),.dout(n3632),.clk(gclk));
	jnot g03397(.din(w_a75_0[1]),.dout(n3633),.clk(gclk));
	jand g03398(.dina(w_n3379_1[0]),.dinb(w_n3633_0[1]),.dout(n3634),.clk(gclk));
	jand g03399(.dina(n3634),.dinb(w_n3632_1[1]),.dout(n3635),.clk(gclk));
	jor g03400(.dina(n3635),.dinb(n3631),.dout(n3636),.clk(gclk));
	jand g03401(.dina(w_n3636_0[2]),.dinb(w_asqrt39_20[1]),.dout(n3637),.clk(gclk));
	jand g03402(.dina(w_asqrt38_30[2]),.dinb(w_n3379_0[2]),.dout(n3638),.clk(gclk));
	jxor g03403(.dina(w_n3638_0[1]),.dinb(w_n3380_0[1]),.dout(n3639),.clk(gclk));
	jor g03404(.dina(w_n3636_0[1]),.dinb(w_asqrt39_20[0]),.dout(n3640),.clk(gclk));
	jand g03405(.dina(n3640),.dinb(w_n3639_0[1]),.dout(n3641),.clk(gclk));
	jor g03406(.dina(w_n3641_0[1]),.dinb(w_n3637_0[1]),.dout(n3642),.clk(gclk));
	jand g03407(.dina(n3642),.dinb(w_asqrt40_22[2]),.dout(n3643),.clk(gclk));
	jor g03408(.dina(w_n3637_0[0]),.dinb(w_asqrt40_22[1]),.dout(n3644),.clk(gclk));
	jor g03409(.dina(n3644),.dinb(w_n3641_0[0]),.dout(n3645),.clk(gclk));
	jand g03410(.dina(w_n3638_0[0]),.dinb(w_n3380_0[0]),.dout(n3646),.clk(gclk));
	jnot g03411(.din(w_n3620_0[0]),.dout(n3647),.clk(gclk));
	jnot g03412(.din(w_n3621_0[1]),.dout(n3648),.clk(gclk));
	jnot g03413(.din(w_n3626_0[0]),.dout(n3649),.clk(gclk));
	jand g03414(.dina(n3649),.dinb(w_asqrt39_19[2]),.dout(n3650),.clk(gclk));
	jand g03415(.dina(n3650),.dinb(n3648),.dout(n3651),.clk(gclk));
	jand g03416(.dina(n3651),.dinb(n3647),.dout(n3652),.clk(gclk));
	jor g03417(.dina(n3652),.dinb(n3646),.dout(n3653),.clk(gclk));
	jxor g03418(.dina(n3653),.dinb(w_n3115_0[1]),.dout(n3654),.clk(gclk));
	jand g03419(.dina(w_n3654_0[1]),.dinb(w_n3645_0[1]),.dout(n3655),.clk(gclk));
	jor g03420(.dina(n3655),.dinb(w_n3643_0[1]),.dout(n3656),.clk(gclk));
	jand g03421(.dina(w_n3656_0[2]),.dinb(w_asqrt41_20[1]),.dout(n3657),.clk(gclk));
	jor g03422(.dina(w_n3656_0[1]),.dinb(w_asqrt41_20[0]),.dout(n3658),.clk(gclk));
	jxor g03423(.dina(w_n3384_0[0]),.dinb(w_n3371_24[2]),.dout(n3659),.clk(gclk));
	jand g03424(.dina(n3659),.dinb(w_asqrt38_30[1]),.dout(n3660),.clk(gclk));
	jxor g03425(.dina(n3660),.dinb(w_n3387_0[0]),.dout(n3661),.clk(gclk));
	jnot g03426(.din(w_n3661_0[1]),.dout(n3662),.clk(gclk));
	jand g03427(.dina(n3662),.dinb(n3658),.dout(n3663),.clk(gclk));
	jor g03428(.dina(w_n3663_0[1]),.dinb(w_n3657_0[1]),.dout(n3664),.clk(gclk));
	jand g03429(.dina(n3664),.dinb(w_asqrt42_22[2]),.dout(n3665),.clk(gclk));
	jnot g03430(.din(w_n3393_0[0]),.dout(n3666),.clk(gclk));
	jand g03431(.dina(n3666),.dinb(w_n3391_0[0]),.dout(n3667),.clk(gclk));
	jand g03432(.dina(n3667),.dinb(w_asqrt38_30[0]),.dout(n3668),.clk(gclk));
	jxor g03433(.dina(n3668),.dinb(w_n3401_0[0]),.dout(n3669),.clk(gclk));
	jnot g03434(.din(n3669),.dout(n3670),.clk(gclk));
	jor g03435(.dina(w_n3657_0[0]),.dinb(w_asqrt42_22[1]),.dout(n3671),.clk(gclk));
	jor g03436(.dina(n3671),.dinb(w_n3663_0[0]),.dout(n3672),.clk(gclk));
	jand g03437(.dina(w_n3672_0[1]),.dinb(w_n3670_0[1]),.dout(n3673),.clk(gclk));
	jor g03438(.dina(w_n3673_0[1]),.dinb(w_n3665_0[1]),.dout(n3674),.clk(gclk));
	jand g03439(.dina(w_n3674_0[2]),.dinb(w_asqrt43_20[1]),.dout(n3675),.clk(gclk));
	jor g03440(.dina(w_n3674_0[1]),.dinb(w_asqrt43_20[0]),.dout(n3676),.clk(gclk));
	jnot g03441(.din(w_n3408_0[0]),.dout(n3677),.clk(gclk));
	jxor g03442(.dina(w_n3403_0[0]),.dinb(w_n2870_24[2]),.dout(n3678),.clk(gclk));
	jand g03443(.dina(n3678),.dinb(w_asqrt38_29[2]),.dout(n3679),.clk(gclk));
	jxor g03444(.dina(n3679),.dinb(n3677),.dout(n3680),.clk(gclk));
	jand g03445(.dina(w_n3680_0[1]),.dinb(n3676),.dout(n3681),.clk(gclk));
	jor g03446(.dina(w_n3681_0[1]),.dinb(w_n3675_0[1]),.dout(n3682),.clk(gclk));
	jand g03447(.dina(n3682),.dinb(w_asqrt44_22[2]),.dout(n3683),.clk(gclk));
	jor g03448(.dina(w_n3675_0[0]),.dinb(w_asqrt44_22[1]),.dout(n3684),.clk(gclk));
	jor g03449(.dina(n3684),.dinb(w_n3681_0[0]),.dout(n3685),.clk(gclk));
	jnot g03450(.din(w_n3415_0[0]),.dout(n3686),.clk(gclk));
	jnot g03451(.din(w_n3417_0[0]),.dout(n3687),.clk(gclk));
	jand g03452(.dina(w_asqrt38_29[1]),.dinb(w_n3411_0[0]),.dout(n3688),.clk(gclk));
	jand g03453(.dina(w_n3688_0[1]),.dinb(n3687),.dout(n3689),.clk(gclk));
	jor g03454(.dina(n3689),.dinb(n3686),.dout(n3690),.clk(gclk));
	jnot g03455(.din(w_n3418_0[0]),.dout(n3691),.clk(gclk));
	jand g03456(.dina(w_n3688_0[0]),.dinb(n3691),.dout(n3692),.clk(gclk));
	jnot g03457(.din(n3692),.dout(n3693),.clk(gclk));
	jand g03458(.dina(n3693),.dinb(n3690),.dout(n3694),.clk(gclk));
	jand g03459(.dina(w_n3694_0[1]),.dinb(w_n3685_0[1]),.dout(n3695),.clk(gclk));
	jor g03460(.dina(n3695),.dinb(w_n3683_0[1]),.dout(n3696),.clk(gclk));
	jand g03461(.dina(w_n3696_0[2]),.dinb(w_asqrt45_20[2]),.dout(n3697),.clk(gclk));
	jor g03462(.dina(w_n3696_0[1]),.dinb(w_asqrt45_20[1]),.dout(n3698),.clk(gclk));
	jxor g03463(.dina(w_n3419_0[0]),.dinb(w_n2420_25[1]),.dout(n3699),.clk(gclk));
	jand g03464(.dina(n3699),.dinb(w_asqrt38_29[0]),.dout(n3700),.clk(gclk));
	jxor g03465(.dina(n3700),.dinb(w_n3424_0[0]),.dout(n3701),.clk(gclk));
	jand g03466(.dina(w_n3701_0[1]),.dinb(n3698),.dout(n3702),.clk(gclk));
	jor g03467(.dina(w_n3702_0[1]),.dinb(w_n3697_0[1]),.dout(n3703),.clk(gclk));
	jand g03468(.dina(n3703),.dinb(w_asqrt46_22[2]),.dout(n3704),.clk(gclk));
	jnot g03469(.din(w_n3430_0[0]),.dout(n3705),.clk(gclk));
	jand g03470(.dina(n3705),.dinb(w_n3428_0[0]),.dout(n3706),.clk(gclk));
	jand g03471(.dina(n3706),.dinb(w_asqrt38_28[2]),.dout(n3707),.clk(gclk));
	jxor g03472(.dina(n3707),.dinb(w_n3438_0[0]),.dout(n3708),.clk(gclk));
	jnot g03473(.din(n3708),.dout(n3709),.clk(gclk));
	jor g03474(.dina(w_n3697_0[0]),.dinb(w_asqrt46_22[1]),.dout(n3710),.clk(gclk));
	jor g03475(.dina(n3710),.dinb(w_n3702_0[0]),.dout(n3711),.clk(gclk));
	jand g03476(.dina(w_n3711_0[1]),.dinb(w_n3709_0[1]),.dout(n3712),.clk(gclk));
	jor g03477(.dina(w_n3712_0[1]),.dinb(w_n3704_0[1]),.dout(n3713),.clk(gclk));
	jand g03478(.dina(w_n3713_0[2]),.dinb(w_asqrt47_20[2]),.dout(n3714),.clk(gclk));
	jor g03479(.dina(w_n3713_0[1]),.dinb(w_asqrt47_20[1]),.dout(n3715),.clk(gclk));
	jxor g03480(.dina(w_n3440_0[0]),.dinb(w_n2005_25[1]),.dout(n3716),.clk(gclk));
	jand g03481(.dina(n3716),.dinb(w_asqrt38_28[1]),.dout(n3717),.clk(gclk));
	jxor g03482(.dina(n3717),.dinb(w_n3446_0[0]),.dout(n3718),.clk(gclk));
	jand g03483(.dina(w_n3718_0[1]),.dinb(n3715),.dout(n3719),.clk(gclk));
	jor g03484(.dina(w_n3719_0[1]),.dinb(w_n3714_0[1]),.dout(n3720),.clk(gclk));
	jand g03485(.dina(n3720),.dinb(w_asqrt48_22[2]),.dout(n3721),.clk(gclk));
	jor g03486(.dina(w_n3714_0[0]),.dinb(w_asqrt48_22[1]),.dout(n3722),.clk(gclk));
	jor g03487(.dina(n3722),.dinb(w_n3719_0[0]),.dout(n3723),.clk(gclk));
	jnot g03488(.din(w_n3454_0[0]),.dout(n3724),.clk(gclk));
	jnot g03489(.din(w_n3456_0[0]),.dout(n3725),.clk(gclk));
	jand g03490(.dina(w_asqrt38_28[0]),.dinb(w_n3450_0[0]),.dout(n3726),.clk(gclk));
	jand g03491(.dina(w_n3726_0[1]),.dinb(n3725),.dout(n3727),.clk(gclk));
	jor g03492(.dina(n3727),.dinb(n3724),.dout(n3728),.clk(gclk));
	jnot g03493(.din(w_n3457_0[0]),.dout(n3729),.clk(gclk));
	jand g03494(.dina(w_n3726_0[0]),.dinb(n3729),.dout(n3730),.clk(gclk));
	jnot g03495(.din(n3730),.dout(n3731),.clk(gclk));
	jand g03496(.dina(n3731),.dinb(n3728),.dout(n3732),.clk(gclk));
	jand g03497(.dina(w_n3732_0[1]),.dinb(w_n3723_0[1]),.dout(n3733),.clk(gclk));
	jor g03498(.dina(n3733),.dinb(w_n3721_0[1]),.dout(n3734),.clk(gclk));
	jand g03499(.dina(w_n3734_0[1]),.dinb(w_asqrt49_21[0]),.dout(n3735),.clk(gclk));
	jxor g03500(.dina(w_n3458_0[0]),.dinb(w_n1641_25[2]),.dout(n3736),.clk(gclk));
	jand g03501(.dina(n3736),.dinb(w_asqrt38_27[2]),.dout(n3737),.clk(gclk));
	jxor g03502(.dina(n3737),.dinb(w_n3465_0[0]),.dout(n3738),.clk(gclk));
	jnot g03503(.din(n3738),.dout(n3739),.clk(gclk));
	jor g03504(.dina(w_n3734_0[0]),.dinb(w_asqrt49_20[2]),.dout(n3740),.clk(gclk));
	jand g03505(.dina(w_n3740_0[1]),.dinb(w_n3739_0[1]),.dout(n3741),.clk(gclk));
	jor g03506(.dina(w_n3741_0[2]),.dinb(w_n3735_0[2]),.dout(n3742),.clk(gclk));
	jand g03507(.dina(n3742),.dinb(w_asqrt50_22[2]),.dout(n3743),.clk(gclk));
	jnot g03508(.din(w_n3470_0[0]),.dout(n3744),.clk(gclk));
	jand g03509(.dina(n3744),.dinb(w_n3468_0[0]),.dout(n3745),.clk(gclk));
	jand g03510(.dina(n3745),.dinb(w_asqrt38_27[1]),.dout(n3746),.clk(gclk));
	jxor g03511(.dina(n3746),.dinb(w_n3478_0[0]),.dout(n3747),.clk(gclk));
	jnot g03512(.din(n3747),.dout(n3748),.clk(gclk));
	jor g03513(.dina(w_n3735_0[1]),.dinb(w_asqrt50_22[1]),.dout(n3749),.clk(gclk));
	jor g03514(.dina(n3749),.dinb(w_n3741_0[1]),.dout(n3750),.clk(gclk));
	jand g03515(.dina(w_n3750_0[1]),.dinb(w_n3748_0[1]),.dout(n3751),.clk(gclk));
	jor g03516(.dina(w_n3751_0[1]),.dinb(w_n3743_0[1]),.dout(n3752),.clk(gclk));
	jand g03517(.dina(w_n3752_0[2]),.dinb(w_asqrt51_21[0]),.dout(n3753),.clk(gclk));
	jor g03518(.dina(w_n3752_0[1]),.dinb(w_asqrt51_20[2]),.dout(n3754),.clk(gclk));
	jnot g03519(.din(w_n3484_0[0]),.dout(n3755),.clk(gclk));
	jnot g03520(.din(w_n3485_0[0]),.dout(n3756),.clk(gclk));
	jand g03521(.dina(w_asqrt38_27[0]),.dinb(w_n3481_0[0]),.dout(n3757),.clk(gclk));
	jand g03522(.dina(w_n3757_0[1]),.dinb(n3756),.dout(n3758),.clk(gclk));
	jor g03523(.dina(n3758),.dinb(n3755),.dout(n3759),.clk(gclk));
	jnot g03524(.din(w_n3486_0[0]),.dout(n3760),.clk(gclk));
	jand g03525(.dina(w_n3757_0[0]),.dinb(n3760),.dout(n3761),.clk(gclk));
	jnot g03526(.din(n3761),.dout(n3762),.clk(gclk));
	jand g03527(.dina(n3762),.dinb(n3759),.dout(n3763),.clk(gclk));
	jand g03528(.dina(w_n3763_0[1]),.dinb(n3754),.dout(n3764),.clk(gclk));
	jor g03529(.dina(w_n3764_0[1]),.dinb(w_n3753_0[1]),.dout(n3765),.clk(gclk));
	jand g03530(.dina(n3765),.dinb(w_asqrt52_22[2]),.dout(n3766),.clk(gclk));
	jor g03531(.dina(w_n3753_0[0]),.dinb(w_asqrt52_22[1]),.dout(n3767),.clk(gclk));
	jor g03532(.dina(n3767),.dinb(w_n3764_0[0]),.dout(n3768),.clk(gclk));
	jnot g03533(.din(w_n3492_0[0]),.dout(n3769),.clk(gclk));
	jnot g03534(.din(w_n3494_0[0]),.dout(n3770),.clk(gclk));
	jand g03535(.dina(w_asqrt38_26[2]),.dinb(w_n3488_0[0]),.dout(n3771),.clk(gclk));
	jand g03536(.dina(w_n3771_0[1]),.dinb(n3770),.dout(n3772),.clk(gclk));
	jor g03537(.dina(n3772),.dinb(n3769),.dout(n3773),.clk(gclk));
	jnot g03538(.din(w_n3495_0[0]),.dout(n3774),.clk(gclk));
	jand g03539(.dina(w_n3771_0[0]),.dinb(n3774),.dout(n3775),.clk(gclk));
	jnot g03540(.din(n3775),.dout(n3776),.clk(gclk));
	jand g03541(.dina(n3776),.dinb(n3773),.dout(n3777),.clk(gclk));
	jand g03542(.dina(w_n3777_0[1]),.dinb(w_n3768_0[1]),.dout(n3778),.clk(gclk));
	jor g03543(.dina(n3778),.dinb(w_n3766_0[1]),.dout(n3779),.clk(gclk));
	jand g03544(.dina(w_n3779_0[1]),.dinb(w_asqrt53_21[1]),.dout(n3780),.clk(gclk));
	jxor g03545(.dina(w_n3496_0[0]),.dinb(w_n1034_26[2]),.dout(n3781),.clk(gclk));
	jand g03546(.dina(n3781),.dinb(w_asqrt38_26[1]),.dout(n3782),.clk(gclk));
	jxor g03547(.dina(n3782),.dinb(w_n3506_0[0]),.dout(n3783),.clk(gclk));
	jnot g03548(.din(n3783),.dout(n3784),.clk(gclk));
	jor g03549(.dina(w_n3779_0[0]),.dinb(w_asqrt53_21[0]),.dout(n3785),.clk(gclk));
	jand g03550(.dina(w_n3785_0[1]),.dinb(w_n3784_0[1]),.dout(n3786),.clk(gclk));
	jor g03551(.dina(w_n3786_0[2]),.dinb(w_n3780_0[2]),.dout(n3787),.clk(gclk));
	jand g03552(.dina(n3787),.dinb(w_asqrt54_22[2]),.dout(n3788),.clk(gclk));
	jnot g03553(.din(w_n3511_0[0]),.dout(n3789),.clk(gclk));
	jand g03554(.dina(n3789),.dinb(w_n3509_0[0]),.dout(n3790),.clk(gclk));
	jand g03555(.dina(n3790),.dinb(w_asqrt38_26[0]),.dout(n3791),.clk(gclk));
	jxor g03556(.dina(n3791),.dinb(w_n3519_0[0]),.dout(n3792),.clk(gclk));
	jnot g03557(.din(n3792),.dout(n3793),.clk(gclk));
	jor g03558(.dina(w_n3780_0[1]),.dinb(w_asqrt54_22[1]),.dout(n3794),.clk(gclk));
	jor g03559(.dina(n3794),.dinb(w_n3786_0[1]),.dout(n3795),.clk(gclk));
	jand g03560(.dina(w_n3795_0[1]),.dinb(w_n3793_0[1]),.dout(n3796),.clk(gclk));
	jor g03561(.dina(w_n3796_0[1]),.dinb(w_n3788_0[1]),.dout(n3797),.clk(gclk));
	jand g03562(.dina(w_n3797_0[2]),.dinb(w_asqrt55_21[2]),.dout(n3798),.clk(gclk));
	jor g03563(.dina(w_n3797_0[1]),.dinb(w_asqrt55_21[1]),.dout(n3799),.clk(gclk));
	jnot g03564(.din(w_n3525_0[0]),.dout(n3800),.clk(gclk));
	jnot g03565(.din(w_n3526_0[0]),.dout(n3801),.clk(gclk));
	jand g03566(.dina(w_asqrt38_25[2]),.dinb(w_n3522_0[0]),.dout(n3802),.clk(gclk));
	jand g03567(.dina(w_n3802_0[1]),.dinb(n3801),.dout(n3803),.clk(gclk));
	jor g03568(.dina(n3803),.dinb(n3800),.dout(n3804),.clk(gclk));
	jnot g03569(.din(w_n3527_0[0]),.dout(n3805),.clk(gclk));
	jand g03570(.dina(w_n3802_0[0]),.dinb(n3805),.dout(n3806),.clk(gclk));
	jnot g03571(.din(n3806),.dout(n3807),.clk(gclk));
	jand g03572(.dina(n3807),.dinb(n3804),.dout(n3808),.clk(gclk));
	jand g03573(.dina(w_n3808_0[1]),.dinb(n3799),.dout(n3809),.clk(gclk));
	jor g03574(.dina(w_n3809_0[1]),.dinb(w_n3798_0[1]),.dout(n3810),.clk(gclk));
	jand g03575(.dina(n3810),.dinb(w_asqrt56_22[2]),.dout(n3811),.clk(gclk));
	jor g03576(.dina(w_n3798_0[0]),.dinb(w_asqrt56_22[1]),.dout(n3812),.clk(gclk));
	jor g03577(.dina(n3812),.dinb(w_n3809_0[0]),.dout(n3813),.clk(gclk));
	jnot g03578(.din(w_n3533_0[0]),.dout(n3814),.clk(gclk));
	jnot g03579(.din(w_n3535_0[0]),.dout(n3815),.clk(gclk));
	jand g03580(.dina(w_asqrt38_25[1]),.dinb(w_n3529_0[0]),.dout(n3816),.clk(gclk));
	jand g03581(.dina(w_n3816_0[1]),.dinb(n3815),.dout(n3817),.clk(gclk));
	jor g03582(.dina(n3817),.dinb(n3814),.dout(n3818),.clk(gclk));
	jnot g03583(.din(w_n3536_0[0]),.dout(n3819),.clk(gclk));
	jand g03584(.dina(w_n3816_0[0]),.dinb(n3819),.dout(n3820),.clk(gclk));
	jnot g03585(.din(n3820),.dout(n3821),.clk(gclk));
	jand g03586(.dina(n3821),.dinb(n3818),.dout(n3822),.clk(gclk));
	jand g03587(.dina(w_n3822_0[1]),.dinb(w_n3813_0[1]),.dout(n3823),.clk(gclk));
	jor g03588(.dina(n3823),.dinb(w_n3811_0[1]),.dout(n3824),.clk(gclk));
	jand g03589(.dina(w_n3824_0[1]),.dinb(w_asqrt57_22[0]),.dout(n3825),.clk(gclk));
	jxor g03590(.dina(w_n3537_0[0]),.dinb(w_n590_27[1]),.dout(n3826),.clk(gclk));
	jand g03591(.dina(n3826),.dinb(w_asqrt38_25[0]),.dout(n3827),.clk(gclk));
	jxor g03592(.dina(n3827),.dinb(w_n3547_0[0]),.dout(n3828),.clk(gclk));
	jnot g03593(.din(n3828),.dout(n3829),.clk(gclk));
	jor g03594(.dina(w_n3824_0[0]),.dinb(w_asqrt57_21[2]),.dout(n3830),.clk(gclk));
	jand g03595(.dina(w_n3830_0[1]),.dinb(w_n3829_0[1]),.dout(n3831),.clk(gclk));
	jor g03596(.dina(w_n3831_0[2]),.dinb(w_n3825_0[2]),.dout(n3832),.clk(gclk));
	jand g03597(.dina(n3832),.dinb(w_asqrt58_22[2]),.dout(n3833),.clk(gclk));
	jnot g03598(.din(w_n3552_0[0]),.dout(n3834),.clk(gclk));
	jand g03599(.dina(n3834),.dinb(w_n3550_0[0]),.dout(n3835),.clk(gclk));
	jand g03600(.dina(n3835),.dinb(w_asqrt38_24[2]),.dout(n3836),.clk(gclk));
	jxor g03601(.dina(n3836),.dinb(w_n3560_0[0]),.dout(n3837),.clk(gclk));
	jnot g03602(.din(n3837),.dout(n3838),.clk(gclk));
	jor g03603(.dina(w_n3825_0[1]),.dinb(w_asqrt58_22[1]),.dout(n3839),.clk(gclk));
	jor g03604(.dina(n3839),.dinb(w_n3831_0[1]),.dout(n3840),.clk(gclk));
	jand g03605(.dina(w_n3840_0[1]),.dinb(w_n3838_0[1]),.dout(n3841),.clk(gclk));
	jor g03606(.dina(w_n3841_0[1]),.dinb(w_n3833_0[1]),.dout(n3842),.clk(gclk));
	jand g03607(.dina(w_n3842_0[2]),.dinb(w_asqrt59_22[1]),.dout(n3843),.clk(gclk));
	jor g03608(.dina(w_n3842_0[1]),.dinb(w_asqrt59_22[0]),.dout(n3844),.clk(gclk));
	jnot g03609(.din(w_n3566_0[0]),.dout(n3845),.clk(gclk));
	jnot g03610(.din(w_n3567_0[0]),.dout(n3846),.clk(gclk));
	jand g03611(.dina(w_asqrt38_24[1]),.dinb(w_n3563_0[0]),.dout(n3847),.clk(gclk));
	jand g03612(.dina(w_n3847_0[1]),.dinb(n3846),.dout(n3848),.clk(gclk));
	jor g03613(.dina(n3848),.dinb(n3845),.dout(n3849),.clk(gclk));
	jnot g03614(.din(w_n3568_0[0]),.dout(n3850),.clk(gclk));
	jand g03615(.dina(w_n3847_0[0]),.dinb(n3850),.dout(n3851),.clk(gclk));
	jnot g03616(.din(n3851),.dout(n3852),.clk(gclk));
	jand g03617(.dina(n3852),.dinb(n3849),.dout(n3853),.clk(gclk));
	jand g03618(.dina(w_n3853_0[1]),.dinb(n3844),.dout(n3854),.clk(gclk));
	jor g03619(.dina(w_n3854_0[1]),.dinb(w_n3843_0[1]),.dout(n3855),.clk(gclk));
	jand g03620(.dina(n3855),.dinb(w_asqrt60_22[1]),.dout(n3856),.clk(gclk));
	jor g03621(.dina(w_n3843_0[0]),.dinb(w_asqrt60_22[0]),.dout(n3857),.clk(gclk));
	jor g03622(.dina(n3857),.dinb(w_n3854_0[0]),.dout(n3858),.clk(gclk));
	jnot g03623(.din(w_n3574_0[0]),.dout(n3859),.clk(gclk));
	jnot g03624(.din(w_n3576_0[0]),.dout(n3860),.clk(gclk));
	jand g03625(.dina(w_asqrt38_24[0]),.dinb(w_n3570_0[0]),.dout(n3861),.clk(gclk));
	jand g03626(.dina(w_n3861_0[1]),.dinb(n3860),.dout(n3862),.clk(gclk));
	jor g03627(.dina(n3862),.dinb(n3859),.dout(n3863),.clk(gclk));
	jnot g03628(.din(w_n3577_0[0]),.dout(n3864),.clk(gclk));
	jand g03629(.dina(w_n3861_0[0]),.dinb(n3864),.dout(n3865),.clk(gclk));
	jnot g03630(.din(n3865),.dout(n3866),.clk(gclk));
	jand g03631(.dina(n3866),.dinb(n3863),.dout(n3867),.clk(gclk));
	jand g03632(.dina(w_n3867_0[1]),.dinb(w_n3858_0[1]),.dout(n3868),.clk(gclk));
	jor g03633(.dina(n3868),.dinb(w_n3856_0[1]),.dout(n3869),.clk(gclk));
	jand g03634(.dina(w_n3869_0[1]),.dinb(w_asqrt61_22[2]),.dout(n3870),.clk(gclk));
	jxor g03635(.dina(w_n3578_0[0]),.dinb(w_n290_28[2]),.dout(n3871),.clk(gclk));
	jand g03636(.dina(n3871),.dinb(w_asqrt38_23[2]),.dout(n3872),.clk(gclk));
	jxor g03637(.dina(n3872),.dinb(w_n3588_0[0]),.dout(n3873),.clk(gclk));
	jnot g03638(.din(n3873),.dout(n3874),.clk(gclk));
	jor g03639(.dina(w_n3869_0[0]),.dinb(w_asqrt61_22[1]),.dout(n3875),.clk(gclk));
	jand g03640(.dina(w_n3875_0[1]),.dinb(w_n3874_0[1]),.dout(n3876),.clk(gclk));
	jor g03641(.dina(w_n3876_0[2]),.dinb(w_n3870_0[2]),.dout(n3877),.clk(gclk));
	jand g03642(.dina(n3877),.dinb(w_asqrt62_22[2]),.dout(n3878),.clk(gclk));
	jnot g03643(.din(w_n3593_0[0]),.dout(n3879),.clk(gclk));
	jand g03644(.dina(n3879),.dinb(w_n3591_0[0]),.dout(n3880),.clk(gclk));
	jand g03645(.dina(n3880),.dinb(w_asqrt38_23[1]),.dout(n3881),.clk(gclk));
	jxor g03646(.dina(n3881),.dinb(w_n3601_0[0]),.dout(n3882),.clk(gclk));
	jnot g03647(.din(n3882),.dout(n3883),.clk(gclk));
	jor g03648(.dina(w_n3870_0[1]),.dinb(w_asqrt62_22[1]),.dout(n3884),.clk(gclk));
	jor g03649(.dina(n3884),.dinb(w_n3876_0[1]),.dout(n3885),.clk(gclk));
	jand g03650(.dina(w_n3885_0[1]),.dinb(w_n3883_0[1]),.dout(n3886),.clk(gclk));
	jor g03651(.dina(w_n3886_0[1]),.dinb(w_n3878_0[1]),.dout(n3887),.clk(gclk));
	jxor g03652(.dina(w_n3603_0[0]),.dinb(w_n199_33[2]),.dout(n3888),.clk(gclk));
	jand g03653(.dina(n3888),.dinb(w_asqrt38_23[0]),.dout(n3889),.clk(gclk));
	jxor g03654(.dina(n3889),.dinb(w_n3608_0[0]),.dout(n3890),.clk(gclk));
	jnot g03655(.din(w_n3610_0[0]),.dout(n3891),.clk(gclk));
	jnot g03656(.din(w_n3614_0[0]),.dout(n3892),.clk(gclk));
	jand g03657(.dina(w_asqrt38_22[2]),.dinb(w_n3892_0[1]),.dout(n3893),.clk(gclk));
	jand g03658(.dina(w_n3893_0[1]),.dinb(w_n3891_0[2]),.dout(n3894),.clk(gclk));
	jor g03659(.dina(n3894),.dinb(w_n3621_0[0]),.dout(n3895),.clk(gclk));
	jor g03660(.dina(n3895),.dinb(w_n3890_0[1]),.dout(n3896),.clk(gclk));
	jnot g03661(.din(n3896),.dout(n3897),.clk(gclk));
	jand g03662(.dina(n3897),.dinb(w_n3887_1[2]),.dout(n3898),.clk(gclk));
	jor g03663(.dina(n3898),.dinb(w_asqrt63_12[0]),.dout(n3899),.clk(gclk));
	jnot g03664(.din(w_n3890_0[0]),.dout(n3900),.clk(gclk));
	jor g03665(.dina(w_n3900_0[2]),.dinb(w_n3887_1[1]),.dout(n3901),.clk(gclk));
	jor g03666(.dina(w_n3893_0[0]),.dinb(w_n3891_0[1]),.dout(n3902),.clk(gclk));
	jand g03667(.dina(w_n3892_0[0]),.dinb(w_n3891_0[0]),.dout(n3903),.clk(gclk));
	jor g03668(.dina(n3903),.dinb(w_n194_32[2]),.dout(n3904),.clk(gclk));
	jnot g03669(.din(n3904),.dout(n3905),.clk(gclk));
	jand g03670(.dina(n3905),.dinb(n3902),.dout(n3906),.clk(gclk));
	jnot g03671(.din(w_asqrt38_22[1]),.dout(n3907),.clk(gclk));
	jnot g03672(.din(w_n3906_0[1]),.dout(n3910),.clk(gclk));
	jand g03673(.dina(n3910),.dinb(w_n3901_0[1]),.dout(n3911),.clk(gclk));
	jand g03674(.dina(n3911),.dinb(w_n3899_0[1]),.dout(n3912),.clk(gclk));
	jnot g03675(.din(w_n3912_31[2]),.dout(asqrt_fa_38),.clk(gclk));
	jor g03676(.dina(w_n3912_31[1]),.dinb(w_n3632_1[0]),.dout(n3914),.clk(gclk));
	jnot g03677(.din(w_a72_0[1]),.dout(n3915),.clk(gclk));
	jnot g03678(.din(a[73]),.dout(n3916),.clk(gclk));
	jand g03679(.dina(w_n3632_0[2]),.dinb(w_n3916_0[2]),.dout(n3917),.clk(gclk));
	jand g03680(.dina(n3917),.dinb(w_n3915_1[1]),.dout(n3918),.clk(gclk));
	jnot g03681(.din(n3918),.dout(n3919),.clk(gclk));
	jand g03682(.dina(n3919),.dinb(n3914),.dout(n3920),.clk(gclk));
	jor g03683(.dina(w_n3920_0[2]),.dinb(w_n3907_24[1]),.dout(n3921),.clk(gclk));
	jor g03684(.dina(w_n3912_31[0]),.dinb(w_a74_0[0]),.dout(n3922),.clk(gclk));
	jxor g03685(.dina(w_n3922_0[1]),.dinb(w_n3633_0[0]),.dout(n3923),.clk(gclk));
	jand g03686(.dina(w_n3920_0[1]),.dinb(w_n3907_24[0]),.dout(n3924),.clk(gclk));
	jor g03687(.dina(n3924),.dinb(w_n3923_0[1]),.dout(n3925),.clk(gclk));
	jand g03688(.dina(w_n3925_0[1]),.dinb(w_n3921_0[1]),.dout(n3926),.clk(gclk));
	jor g03689(.dina(n3926),.dinb(w_n3376_27[2]),.dout(n3927),.clk(gclk));
	jand g03690(.dina(w_n3921_0[0]),.dinb(w_n3376_27[1]),.dout(n3928),.clk(gclk));
	jand g03691(.dina(n3928),.dinb(w_n3925_0[0]),.dout(n3929),.clk(gclk));
	jor g03692(.dina(w_n3922_0[0]),.dinb(w_a75_0[0]),.dout(n3930),.clk(gclk));
	jnot g03693(.din(w_n3899_0[0]),.dout(n3931),.clk(gclk));
	jnot g03694(.din(w_n3901_0[0]),.dout(n3932),.clk(gclk));
	jor g03695(.dina(w_n3906_0[0]),.dinb(w_n3907_23[2]),.dout(n3933),.clk(gclk));
	jor g03696(.dina(n3933),.dinb(w_n3932_0[1]),.dout(n3934),.clk(gclk));
	jor g03697(.dina(n3934),.dinb(n3931),.dout(n3935),.clk(gclk));
	jand g03698(.dina(n3935),.dinb(n3930),.dout(n3936),.clk(gclk));
	jxor g03699(.dina(n3936),.dinb(w_n3379_0[1]),.dout(n3937),.clk(gclk));
	jor g03700(.dina(w_n3937_0[1]),.dinb(w_n3929_0[1]),.dout(n3938),.clk(gclk));
	jand g03701(.dina(n3938),.dinb(w_n3927_0[1]),.dout(n3939),.clk(gclk));
	jor g03702(.dina(w_n3939_0[2]),.dinb(w_n3371_24[1]),.dout(n3940),.clk(gclk));
	jand g03703(.dina(w_n3939_0[1]),.dinb(w_n3371_24[0]),.dout(n3941),.clk(gclk));
	jxor g03704(.dina(w_n3636_0[0]),.dinb(w_n3376_27[0]),.dout(n3942),.clk(gclk));
	jor g03705(.dina(n3942),.dinb(w_n3912_30[2]),.dout(n3943),.clk(gclk));
	jxor g03706(.dina(n3943),.dinb(w_n3639_0[0]),.dout(n3944),.clk(gclk));
	jor g03707(.dina(w_n3944_0[1]),.dinb(n3941),.dout(n3945),.clk(gclk));
	jand g03708(.dina(w_n3945_0[1]),.dinb(w_n3940_0[1]),.dout(n3946),.clk(gclk));
	jor g03709(.dina(n3946),.dinb(w_n2875_27[1]),.dout(n3947),.clk(gclk));
	jnot g03710(.din(w_n3645_0[0]),.dout(n3948),.clk(gclk));
	jor g03711(.dina(n3948),.dinb(w_n3643_0[0]),.dout(n3949),.clk(gclk));
	jor g03712(.dina(n3949),.dinb(w_n3912_30[1]),.dout(n3950),.clk(gclk));
	jxor g03713(.dina(n3950),.dinb(w_n3654_0[0]),.dout(n3951),.clk(gclk));
	jand g03714(.dina(w_n3940_0[0]),.dinb(w_n2875_27[0]),.dout(n3952),.clk(gclk));
	jand g03715(.dina(n3952),.dinb(w_n3945_0[0]),.dout(n3953),.clk(gclk));
	jor g03716(.dina(w_n3953_0[1]),.dinb(w_n3951_0[1]),.dout(n3954),.clk(gclk));
	jand g03717(.dina(w_n3954_0[1]),.dinb(w_n3947_0[1]),.dout(n3955),.clk(gclk));
	jor g03718(.dina(w_n3955_0[2]),.dinb(w_n2870_24[1]),.dout(n3956),.clk(gclk));
	jand g03719(.dina(w_n3955_0[1]),.dinb(w_n2870_24[0]),.dout(n3957),.clk(gclk));
	jxor g03720(.dina(w_n3656_0[0]),.dinb(w_n2875_26[2]),.dout(n3958),.clk(gclk));
	jor g03721(.dina(n3958),.dinb(w_n3912_30[0]),.dout(n3959),.clk(gclk));
	jxor g03722(.dina(n3959),.dinb(w_n3661_0[0]),.dout(n3960),.clk(gclk));
	jnot g03723(.din(w_n3960_0[1]),.dout(n3961),.clk(gclk));
	jor g03724(.dina(n3961),.dinb(n3957),.dout(n3962),.clk(gclk));
	jand g03725(.dina(w_n3962_0[1]),.dinb(w_n3956_0[1]),.dout(n3963),.clk(gclk));
	jor g03726(.dina(n3963),.dinb(w_n2425_27[2]),.dout(n3964),.clk(gclk));
	jand g03727(.dina(w_n3956_0[0]),.dinb(w_n2425_27[1]),.dout(n3965),.clk(gclk));
	jand g03728(.dina(n3965),.dinb(w_n3962_0[0]),.dout(n3966),.clk(gclk));
	jnot g03729(.din(w_n3665_0[0]),.dout(n3967),.clk(gclk));
	jand g03730(.dina(w_asqrt37_23[1]),.dinb(n3967),.dout(n3968),.clk(gclk));
	jand g03731(.dina(w_n3968_0[1]),.dinb(w_n3672_0[0]),.dout(n3969),.clk(gclk));
	jor g03732(.dina(n3969),.dinb(w_n3670_0[0]),.dout(n3970),.clk(gclk));
	jand g03733(.dina(w_n3968_0[0]),.dinb(w_n3673_0[0]),.dout(n3971),.clk(gclk));
	jnot g03734(.din(n3971),.dout(n3972),.clk(gclk));
	jand g03735(.dina(n3972),.dinb(n3970),.dout(n3973),.clk(gclk));
	jnot g03736(.din(n3973),.dout(n3974),.clk(gclk));
	jor g03737(.dina(w_n3974_0[1]),.dinb(w_n3966_0[1]),.dout(n3975),.clk(gclk));
	jand g03738(.dina(n3975),.dinb(w_n3964_0[1]),.dout(n3976),.clk(gclk));
	jor g03739(.dina(w_n3976_0[2]),.dinb(w_n2420_25[0]),.dout(n3977),.clk(gclk));
	jand g03740(.dina(w_n3976_0[1]),.dinb(w_n2420_24[2]),.dout(n3978),.clk(gclk));
	jnot g03741(.din(w_n3680_0[0]),.dout(n3979),.clk(gclk));
	jxor g03742(.dina(w_n3674_0[0]),.dinb(w_n2425_27[0]),.dout(n3980),.clk(gclk));
	jor g03743(.dina(n3980),.dinb(w_n3912_29[2]),.dout(n3981),.clk(gclk));
	jxor g03744(.dina(n3981),.dinb(n3979),.dout(n3982),.clk(gclk));
	jnot g03745(.din(w_n3982_0[1]),.dout(n3983),.clk(gclk));
	jor g03746(.dina(n3983),.dinb(n3978),.dout(n3984),.clk(gclk));
	jand g03747(.dina(w_n3984_0[1]),.dinb(w_n3977_0[1]),.dout(n3985),.clk(gclk));
	jor g03748(.dina(n3985),.dinb(w_n2010_27[1]),.dout(n3986),.clk(gclk));
	jnot g03749(.din(w_n3685_0[0]),.dout(n3987),.clk(gclk));
	jor g03750(.dina(n3987),.dinb(w_n3683_0[0]),.dout(n3988),.clk(gclk));
	jor g03751(.dina(n3988),.dinb(w_n3912_29[1]),.dout(n3989),.clk(gclk));
	jxor g03752(.dina(n3989),.dinb(w_n3694_0[0]),.dout(n3990),.clk(gclk));
	jand g03753(.dina(w_n3977_0[0]),.dinb(w_n2010_27[0]),.dout(n3991),.clk(gclk));
	jand g03754(.dina(n3991),.dinb(w_n3984_0[0]),.dout(n3992),.clk(gclk));
	jor g03755(.dina(w_n3992_0[1]),.dinb(w_n3990_0[1]),.dout(n3993),.clk(gclk));
	jand g03756(.dina(w_n3993_0[1]),.dinb(w_n3986_0[1]),.dout(n3994),.clk(gclk));
	jor g03757(.dina(w_n3994_0[2]),.dinb(w_n2005_25[0]),.dout(n3995),.clk(gclk));
	jand g03758(.dina(w_n3994_0[1]),.dinb(w_n2005_24[2]),.dout(n3996),.clk(gclk));
	jnot g03759(.din(w_n3701_0[0]),.dout(n3997),.clk(gclk));
	jxor g03760(.dina(w_n3696_0[0]),.dinb(w_n2010_26[2]),.dout(n3998),.clk(gclk));
	jor g03761(.dina(n3998),.dinb(w_n3912_29[0]),.dout(n3999),.clk(gclk));
	jxor g03762(.dina(n3999),.dinb(n3997),.dout(n4000),.clk(gclk));
	jnot g03763(.din(n4000),.dout(n4001),.clk(gclk));
	jor g03764(.dina(w_n4001_0[1]),.dinb(n3996),.dout(n4002),.clk(gclk));
	jand g03765(.dina(w_n4002_0[1]),.dinb(w_n3995_0[1]),.dout(n4003),.clk(gclk));
	jor g03766(.dina(n4003),.dinb(w_n1646_28[0]),.dout(n4004),.clk(gclk));
	jand g03767(.dina(w_n3995_0[0]),.dinb(w_n1646_27[2]),.dout(n4005),.clk(gclk));
	jand g03768(.dina(n4005),.dinb(w_n4002_0[0]),.dout(n4006),.clk(gclk));
	jnot g03769(.din(w_n3704_0[0]),.dout(n4007),.clk(gclk));
	jand g03770(.dina(w_asqrt37_23[0]),.dinb(n4007),.dout(n4008),.clk(gclk));
	jand g03771(.dina(w_n4008_0[1]),.dinb(w_n3711_0[0]),.dout(n4009),.clk(gclk));
	jor g03772(.dina(n4009),.dinb(w_n3709_0[0]),.dout(n4010),.clk(gclk));
	jand g03773(.dina(w_n4008_0[0]),.dinb(w_n3712_0[0]),.dout(n4011),.clk(gclk));
	jnot g03774(.din(n4011),.dout(n4012),.clk(gclk));
	jand g03775(.dina(n4012),.dinb(n4010),.dout(n4013),.clk(gclk));
	jnot g03776(.din(n4013),.dout(n4014),.clk(gclk));
	jor g03777(.dina(w_n4014_0[1]),.dinb(w_n4006_0[1]),.dout(n4015),.clk(gclk));
	jand g03778(.dina(n4015),.dinb(w_n4004_0[1]),.dout(n4016),.clk(gclk));
	jor g03779(.dina(w_n4016_0[1]),.dinb(w_n1641_25[1]),.dout(n4017),.clk(gclk));
	jxor g03780(.dina(w_n3713_0[0]),.dinb(w_n1646_27[1]),.dout(n4018),.clk(gclk));
	jor g03781(.dina(n4018),.dinb(w_n3912_28[2]),.dout(n4019),.clk(gclk));
	jxor g03782(.dina(n4019),.dinb(w_n3718_0[0]),.dout(n4020),.clk(gclk));
	jand g03783(.dina(w_n4016_0[0]),.dinb(w_n1641_25[0]),.dout(n4021),.clk(gclk));
	jor g03784(.dina(w_n4021_0[1]),.dinb(w_n4020_0[1]),.dout(n4022),.clk(gclk));
	jand g03785(.dina(w_n4022_0[2]),.dinb(w_n4017_0[2]),.dout(n4023),.clk(gclk));
	jor g03786(.dina(n4023),.dinb(w_n1317_27[2]),.dout(n4024),.clk(gclk));
	jnot g03787(.din(w_n3723_0[0]),.dout(n4025),.clk(gclk));
	jor g03788(.dina(n4025),.dinb(w_n3721_0[0]),.dout(n4026),.clk(gclk));
	jor g03789(.dina(n4026),.dinb(w_n3912_28[1]),.dout(n4027),.clk(gclk));
	jxor g03790(.dina(n4027),.dinb(w_n3732_0[0]),.dout(n4028),.clk(gclk));
	jand g03791(.dina(w_n4017_0[1]),.dinb(w_n1317_27[1]),.dout(n4029),.clk(gclk));
	jand g03792(.dina(n4029),.dinb(w_n4022_0[1]),.dout(n4030),.clk(gclk));
	jor g03793(.dina(w_n4030_0[1]),.dinb(w_n4028_0[1]),.dout(n4031),.clk(gclk));
	jand g03794(.dina(w_n4031_0[1]),.dinb(w_n4024_0[1]),.dout(n4032),.clk(gclk));
	jor g03795(.dina(w_n4032_0[2]),.dinb(w_n1312_25[2]),.dout(n4033),.clk(gclk));
	jand g03796(.dina(w_n4032_0[1]),.dinb(w_n1312_25[1]),.dout(n4034),.clk(gclk));
	jnot g03797(.din(w_n3735_0[0]),.dout(n4035),.clk(gclk));
	jand g03798(.dina(w_asqrt37_22[2]),.dinb(n4035),.dout(n4036),.clk(gclk));
	jand g03799(.dina(w_n4036_0[1]),.dinb(w_n3740_0[0]),.dout(n4037),.clk(gclk));
	jor g03800(.dina(n4037),.dinb(w_n3739_0[0]),.dout(n4038),.clk(gclk));
	jand g03801(.dina(w_n4036_0[0]),.dinb(w_n3741_0[0]),.dout(n4039),.clk(gclk));
	jnot g03802(.din(n4039),.dout(n4040),.clk(gclk));
	jand g03803(.dina(n4040),.dinb(n4038),.dout(n4041),.clk(gclk));
	jnot g03804(.din(n4041),.dout(n4042),.clk(gclk));
	jor g03805(.dina(w_n4042_0[1]),.dinb(n4034),.dout(n4043),.clk(gclk));
	jand g03806(.dina(w_n4043_0[1]),.dinb(w_n4033_0[1]),.dout(n4044),.clk(gclk));
	jor g03807(.dina(n4044),.dinb(w_n1039_28[1]),.dout(n4045),.clk(gclk));
	jand g03808(.dina(w_n4033_0[0]),.dinb(w_n1039_28[0]),.dout(n4046),.clk(gclk));
	jand g03809(.dina(n4046),.dinb(w_n4043_0[0]),.dout(n4047),.clk(gclk));
	jnot g03810(.din(w_n3743_0[0]),.dout(n4048),.clk(gclk));
	jand g03811(.dina(w_asqrt37_22[1]),.dinb(n4048),.dout(n4049),.clk(gclk));
	jand g03812(.dina(w_n4049_0[1]),.dinb(w_n3750_0[0]),.dout(n4050),.clk(gclk));
	jor g03813(.dina(n4050),.dinb(w_n3748_0[0]),.dout(n4051),.clk(gclk));
	jand g03814(.dina(w_n4049_0[0]),.dinb(w_n3751_0[0]),.dout(n4052),.clk(gclk));
	jnot g03815(.din(n4052),.dout(n4053),.clk(gclk));
	jand g03816(.dina(n4053),.dinb(n4051),.dout(n4054),.clk(gclk));
	jnot g03817(.din(n4054),.dout(n4055),.clk(gclk));
	jor g03818(.dina(w_n4055_0[1]),.dinb(w_n4047_0[1]),.dout(n4056),.clk(gclk));
	jand g03819(.dina(n4056),.dinb(w_n4045_0[1]),.dout(n4057),.clk(gclk));
	jor g03820(.dina(w_n4057_0[1]),.dinb(w_n1034_26[1]),.dout(n4058),.clk(gclk));
	jxor g03821(.dina(w_n3752_0[0]),.dinb(w_n1039_27[2]),.dout(n4059),.clk(gclk));
	jor g03822(.dina(n4059),.dinb(w_n3912_28[0]),.dout(n4060),.clk(gclk));
	jxor g03823(.dina(n4060),.dinb(w_n3763_0[0]),.dout(n4061),.clk(gclk));
	jand g03824(.dina(w_n4057_0[0]),.dinb(w_n1034_26[0]),.dout(n4062),.clk(gclk));
	jor g03825(.dina(w_n4062_0[1]),.dinb(w_n4061_0[1]),.dout(n4063),.clk(gclk));
	jand g03826(.dina(w_n4063_0[2]),.dinb(w_n4058_0[2]),.dout(n4064),.clk(gclk));
	jor g03827(.dina(n4064),.dinb(w_n796_28[0]),.dout(n4065),.clk(gclk));
	jnot g03828(.din(w_n3768_0[0]),.dout(n4066),.clk(gclk));
	jor g03829(.dina(n4066),.dinb(w_n3766_0[0]),.dout(n4067),.clk(gclk));
	jor g03830(.dina(n4067),.dinb(w_n3912_27[2]),.dout(n4068),.clk(gclk));
	jxor g03831(.dina(n4068),.dinb(w_n3777_0[0]),.dout(n4069),.clk(gclk));
	jand g03832(.dina(w_n4058_0[1]),.dinb(w_n796_27[2]),.dout(n4070),.clk(gclk));
	jand g03833(.dina(n4070),.dinb(w_n4063_0[1]),.dout(n4071),.clk(gclk));
	jor g03834(.dina(w_n4071_0[1]),.dinb(w_n4069_0[1]),.dout(n4072),.clk(gclk));
	jand g03835(.dina(w_n4072_0[1]),.dinb(w_n4065_0[1]),.dout(n4073),.clk(gclk));
	jor g03836(.dina(w_n4073_0[2]),.dinb(w_n791_26[2]),.dout(n4074),.clk(gclk));
	jand g03837(.dina(w_n4073_0[1]),.dinb(w_n791_26[1]),.dout(n4075),.clk(gclk));
	jnot g03838(.din(w_n3780_0[0]),.dout(n4076),.clk(gclk));
	jand g03839(.dina(w_asqrt37_22[0]),.dinb(n4076),.dout(n4077),.clk(gclk));
	jand g03840(.dina(w_n4077_0[1]),.dinb(w_n3785_0[0]),.dout(n4078),.clk(gclk));
	jor g03841(.dina(n4078),.dinb(w_n3784_0[0]),.dout(n4079),.clk(gclk));
	jand g03842(.dina(w_n4077_0[0]),.dinb(w_n3786_0[0]),.dout(n4080),.clk(gclk));
	jnot g03843(.din(n4080),.dout(n4081),.clk(gclk));
	jand g03844(.dina(n4081),.dinb(n4079),.dout(n4082),.clk(gclk));
	jnot g03845(.din(n4082),.dout(n4083),.clk(gclk));
	jor g03846(.dina(w_n4083_0[1]),.dinb(n4075),.dout(n4084),.clk(gclk));
	jand g03847(.dina(w_n4084_0[1]),.dinb(w_n4074_0[1]),.dout(n4085),.clk(gclk));
	jor g03848(.dina(n4085),.dinb(w_n595_28[2]),.dout(n4086),.clk(gclk));
	jand g03849(.dina(w_n4074_0[0]),.dinb(w_n595_28[1]),.dout(n4087),.clk(gclk));
	jand g03850(.dina(n4087),.dinb(w_n4084_0[0]),.dout(n4088),.clk(gclk));
	jnot g03851(.din(w_n3788_0[0]),.dout(n4089),.clk(gclk));
	jand g03852(.dina(w_asqrt37_21[2]),.dinb(n4089),.dout(n4090),.clk(gclk));
	jand g03853(.dina(w_n4090_0[1]),.dinb(w_n3795_0[0]),.dout(n4091),.clk(gclk));
	jor g03854(.dina(n4091),.dinb(w_n3793_0[0]),.dout(n4092),.clk(gclk));
	jand g03855(.dina(w_n4090_0[0]),.dinb(w_n3796_0[0]),.dout(n4093),.clk(gclk));
	jnot g03856(.din(n4093),.dout(n4094),.clk(gclk));
	jand g03857(.dina(n4094),.dinb(n4092),.dout(n4095),.clk(gclk));
	jnot g03858(.din(n4095),.dout(n4096),.clk(gclk));
	jor g03859(.dina(w_n4096_0[1]),.dinb(w_n4088_0[1]),.dout(n4097),.clk(gclk));
	jand g03860(.dina(n4097),.dinb(w_n4086_0[1]),.dout(n4098),.clk(gclk));
	jor g03861(.dina(w_n4098_0[1]),.dinb(w_n590_27[0]),.dout(n4099),.clk(gclk));
	jxor g03862(.dina(w_n3797_0[0]),.dinb(w_n595_28[0]),.dout(n4100),.clk(gclk));
	jor g03863(.dina(n4100),.dinb(w_n3912_27[1]),.dout(n4101),.clk(gclk));
	jxor g03864(.dina(n4101),.dinb(w_n3808_0[0]),.dout(n4102),.clk(gclk));
	jand g03865(.dina(w_n4098_0[0]),.dinb(w_n590_26[2]),.dout(n4103),.clk(gclk));
	jor g03866(.dina(w_n4103_0[1]),.dinb(w_n4102_0[1]),.dout(n4104),.clk(gclk));
	jand g03867(.dina(w_n4104_0[2]),.dinb(w_n4099_0[2]),.dout(n4105),.clk(gclk));
	jor g03868(.dina(n4105),.dinb(w_n430_28[1]),.dout(n4106),.clk(gclk));
	jnot g03869(.din(w_n3813_0[0]),.dout(n4107),.clk(gclk));
	jor g03870(.dina(n4107),.dinb(w_n3811_0[0]),.dout(n4108),.clk(gclk));
	jor g03871(.dina(n4108),.dinb(w_n3912_27[0]),.dout(n4109),.clk(gclk));
	jxor g03872(.dina(n4109),.dinb(w_n3822_0[0]),.dout(n4110),.clk(gclk));
	jand g03873(.dina(w_n4099_0[1]),.dinb(w_n430_28[0]),.dout(n4111),.clk(gclk));
	jand g03874(.dina(n4111),.dinb(w_n4104_0[1]),.dout(n4112),.clk(gclk));
	jor g03875(.dina(w_n4112_0[1]),.dinb(w_n4110_0[1]),.dout(n4113),.clk(gclk));
	jand g03876(.dina(w_n4113_0[1]),.dinb(w_n4106_0[1]),.dout(n4114),.clk(gclk));
	jor g03877(.dina(w_n4114_0[2]),.dinb(w_n425_27[1]),.dout(n4115),.clk(gclk));
	jand g03878(.dina(w_n4114_0[1]),.dinb(w_n425_27[0]),.dout(n4116),.clk(gclk));
	jnot g03879(.din(w_n3825_0[0]),.dout(n4117),.clk(gclk));
	jand g03880(.dina(w_asqrt37_21[1]),.dinb(n4117),.dout(n4118),.clk(gclk));
	jand g03881(.dina(w_n4118_0[1]),.dinb(w_n3830_0[0]),.dout(n4119),.clk(gclk));
	jor g03882(.dina(n4119),.dinb(w_n3829_0[0]),.dout(n4120),.clk(gclk));
	jand g03883(.dina(w_n4118_0[0]),.dinb(w_n3831_0[0]),.dout(n4121),.clk(gclk));
	jnot g03884(.din(n4121),.dout(n4122),.clk(gclk));
	jand g03885(.dina(n4122),.dinb(n4120),.dout(n4123),.clk(gclk));
	jnot g03886(.din(n4123),.dout(n4124),.clk(gclk));
	jor g03887(.dina(w_n4124_0[1]),.dinb(n4116),.dout(n4125),.clk(gclk));
	jand g03888(.dina(w_n4125_0[1]),.dinb(w_n4115_0[1]),.dout(n4126),.clk(gclk));
	jor g03889(.dina(n4126),.dinb(w_n305_29[0]),.dout(n4127),.clk(gclk));
	jand g03890(.dina(w_n4115_0[0]),.dinb(w_n305_28[2]),.dout(n4128),.clk(gclk));
	jand g03891(.dina(n4128),.dinb(w_n4125_0[0]),.dout(n4129),.clk(gclk));
	jnot g03892(.din(w_n3833_0[0]),.dout(n4130),.clk(gclk));
	jand g03893(.dina(w_asqrt37_21[0]),.dinb(n4130),.dout(n4131),.clk(gclk));
	jand g03894(.dina(w_n4131_0[1]),.dinb(w_n3840_0[0]),.dout(n4132),.clk(gclk));
	jor g03895(.dina(n4132),.dinb(w_n3838_0[0]),.dout(n4133),.clk(gclk));
	jand g03896(.dina(w_n4131_0[0]),.dinb(w_n3841_0[0]),.dout(n4134),.clk(gclk));
	jnot g03897(.din(n4134),.dout(n4135),.clk(gclk));
	jand g03898(.dina(n4135),.dinb(n4133),.dout(n4136),.clk(gclk));
	jnot g03899(.din(n4136),.dout(n4137),.clk(gclk));
	jor g03900(.dina(w_n4137_0[1]),.dinb(w_n4129_0[1]),.dout(n4138),.clk(gclk));
	jand g03901(.dina(n4138),.dinb(w_n4127_0[1]),.dout(n4139),.clk(gclk));
	jor g03902(.dina(w_n4139_0[1]),.dinb(w_n290_28[1]),.dout(n4140),.clk(gclk));
	jxor g03903(.dina(w_n3842_0[0]),.dinb(w_n305_28[1]),.dout(n4141),.clk(gclk));
	jor g03904(.dina(n4141),.dinb(w_n3912_26[2]),.dout(n4142),.clk(gclk));
	jxor g03905(.dina(n4142),.dinb(w_n3853_0[0]),.dout(n4143),.clk(gclk));
	jand g03906(.dina(w_n4139_0[0]),.dinb(w_n290_28[0]),.dout(n4144),.clk(gclk));
	jor g03907(.dina(w_n4144_0[1]),.dinb(w_n4143_0[1]),.dout(n4145),.clk(gclk));
	jand g03908(.dina(w_n4145_0[2]),.dinb(w_n4140_0[2]),.dout(n4146),.clk(gclk));
	jor g03909(.dina(n4146),.dinb(w_n223_28[2]),.dout(n4147),.clk(gclk));
	jnot g03910(.din(w_n3858_0[0]),.dout(n4148),.clk(gclk));
	jor g03911(.dina(n4148),.dinb(w_n3856_0[0]),.dout(n4149),.clk(gclk));
	jor g03912(.dina(n4149),.dinb(w_n3912_26[1]),.dout(n4150),.clk(gclk));
	jxor g03913(.dina(n4150),.dinb(w_n3867_0[0]),.dout(n4151),.clk(gclk));
	jand g03914(.dina(w_n4140_0[1]),.dinb(w_n223_28[1]),.dout(n4152),.clk(gclk));
	jand g03915(.dina(n4152),.dinb(w_n4145_0[1]),.dout(n4153),.clk(gclk));
	jor g03916(.dina(w_n4153_0[1]),.dinb(w_n4151_0[1]),.dout(n4154),.clk(gclk));
	jand g03917(.dina(w_n4154_0[1]),.dinb(w_n4147_0[1]),.dout(n4155),.clk(gclk));
	jor g03918(.dina(w_n4155_0[2]),.dinb(w_n199_33[1]),.dout(n4156),.clk(gclk));
	jand g03919(.dina(w_n4155_0[1]),.dinb(w_n199_33[0]),.dout(n4157),.clk(gclk));
	jnot g03920(.din(w_n3870_0[0]),.dout(n4158),.clk(gclk));
	jand g03921(.dina(w_asqrt37_20[2]),.dinb(n4158),.dout(n4159),.clk(gclk));
	jand g03922(.dina(w_n4159_0[1]),.dinb(w_n3875_0[0]),.dout(n4160),.clk(gclk));
	jor g03923(.dina(n4160),.dinb(w_n3874_0[0]),.dout(n4161),.clk(gclk));
	jand g03924(.dina(w_n4159_0[0]),.dinb(w_n3876_0[0]),.dout(n4162),.clk(gclk));
	jnot g03925(.din(n4162),.dout(n4163),.clk(gclk));
	jand g03926(.dina(n4163),.dinb(n4161),.dout(n4164),.clk(gclk));
	jnot g03927(.din(n4164),.dout(n4165),.clk(gclk));
	jor g03928(.dina(w_n4165_0[1]),.dinb(n4157),.dout(n4166),.clk(gclk));
	jand g03929(.dina(n4166),.dinb(n4156),.dout(n4167),.clk(gclk));
	jnot g03930(.din(w_n3878_0[0]),.dout(n4168),.clk(gclk));
	jand g03931(.dina(w_asqrt37_20[1]),.dinb(n4168),.dout(n4169),.clk(gclk));
	jand g03932(.dina(w_n4169_0[1]),.dinb(w_n3885_0[0]),.dout(n4170),.clk(gclk));
	jor g03933(.dina(n4170),.dinb(w_n3883_0[0]),.dout(n4171),.clk(gclk));
	jand g03934(.dina(w_n4169_0[0]),.dinb(w_n3886_0[0]),.dout(n4172),.clk(gclk));
	jnot g03935(.din(n4172),.dout(n4173),.clk(gclk));
	jand g03936(.dina(n4173),.dinb(n4171),.dout(n4174),.clk(gclk));
	jnot g03937(.din(w_n4174_0[2]),.dout(n4175),.clk(gclk));
	jand g03938(.dina(w_asqrt37_20[0]),.dinb(w_n3900_0[1]),.dout(n4176),.clk(gclk));
	jand g03939(.dina(w_n4176_0[1]),.dinb(w_n3887_1[0]),.dout(n4177),.clk(gclk));
	jor g03940(.dina(n4177),.dinb(w_n3932_0[0]),.dout(n4178),.clk(gclk));
	jor g03941(.dina(n4178),.dinb(w_n4175_0[1]),.dout(n4179),.clk(gclk));
	jor g03942(.dina(n4179),.dinb(w_n4167_0[2]),.dout(n4180),.clk(gclk));
	jand g03943(.dina(n4180),.dinb(w_n194_32[1]),.dout(n4181),.clk(gclk));
	jand g03944(.dina(w_n4175_0[0]),.dinb(w_n4167_0[1]),.dout(n4182),.clk(gclk));
	jor g03945(.dina(w_n4176_0[0]),.dinb(w_n3887_0[2]),.dout(n4183),.clk(gclk));
	jand g03946(.dina(w_n3900_0[0]),.dinb(w_n3887_0[1]),.dout(n4184),.clk(gclk));
	jor g03947(.dina(n4184),.dinb(w_n194_32[0]),.dout(n4185),.clk(gclk));
	jnot g03948(.din(n4185),.dout(n4186),.clk(gclk));
	jand g03949(.dina(n4186),.dinb(n4183),.dout(n4187),.clk(gclk));
	jor g03950(.dina(w_n4187_0[1]),.dinb(w_n4182_0[2]),.dout(n4190),.clk(gclk));
	jor g03951(.dina(n4190),.dinb(w_n4181_0[1]),.dout(asqrt_fa_37),.clk(gclk));
	jand g03952(.dina(w_asqrt36_31),.dinb(w_a72_0[0]),.dout(n4192),.clk(gclk));
	jnot g03953(.din(w_a70_0[1]),.dout(n4193),.clk(gclk));
	jnot g03954(.din(w_a71_0[1]),.dout(n4194),.clk(gclk));
	jand g03955(.dina(w_n3915_1[0]),.dinb(w_n4194_0[1]),.dout(n4195),.clk(gclk));
	jand g03956(.dina(n4195),.dinb(w_n4193_1[1]),.dout(n4196),.clk(gclk));
	jor g03957(.dina(n4196),.dinb(n4192),.dout(n4197),.clk(gclk));
	jand g03958(.dina(w_n4197_0[2]),.dinb(w_asqrt37_19[2]),.dout(n4198),.clk(gclk));
	jand g03959(.dina(w_asqrt36_30[2]),.dinb(w_n3915_0[2]),.dout(n4199),.clk(gclk));
	jxor g03960(.dina(w_n4199_0[1]),.dinb(w_n3916_0[1]),.dout(n4200),.clk(gclk));
	jor g03961(.dina(w_n4197_0[1]),.dinb(w_asqrt37_19[1]),.dout(n4201),.clk(gclk));
	jand g03962(.dina(n4201),.dinb(w_n4200_0[1]),.dout(n4202),.clk(gclk));
	jor g03963(.dina(w_n4202_0[1]),.dinb(w_n4198_0[1]),.dout(n4203),.clk(gclk));
	jand g03964(.dina(n4203),.dinb(w_asqrt38_22[0]),.dout(n4204),.clk(gclk));
	jor g03965(.dina(w_n4198_0[0]),.dinb(w_asqrt38_21[2]),.dout(n4205),.clk(gclk));
	jor g03966(.dina(n4205),.dinb(w_n4202_0[0]),.dout(n4206),.clk(gclk));
	jand g03967(.dina(w_n4199_0[0]),.dinb(w_n3916_0[0]),.dout(n4207),.clk(gclk));
	jnot g03968(.din(w_n4181_0[0]),.dout(n4208),.clk(gclk));
	jnot g03969(.din(w_n4182_0[1]),.dout(n4209),.clk(gclk));
	jnot g03970(.din(w_n4187_0[0]),.dout(n4210),.clk(gclk));
	jand g03971(.dina(n4210),.dinb(w_asqrt37_19[0]),.dout(n4211),.clk(gclk));
	jand g03972(.dina(n4211),.dinb(n4209),.dout(n4212),.clk(gclk));
	jand g03973(.dina(n4212),.dinb(n4208),.dout(n4213),.clk(gclk));
	jor g03974(.dina(n4213),.dinb(n4207),.dout(n4214),.clk(gclk));
	jxor g03975(.dina(n4214),.dinb(w_n3632_0[1]),.dout(n4215),.clk(gclk));
	jand g03976(.dina(w_n4215_0[1]),.dinb(w_n4206_0[1]),.dout(n4216),.clk(gclk));
	jor g03977(.dina(n4216),.dinb(w_n4204_0[1]),.dout(n4217),.clk(gclk));
	jand g03978(.dina(w_n4217_0[2]),.dinb(w_asqrt39_19[1]),.dout(n4218),.clk(gclk));
	jor g03979(.dina(w_n4217_0[1]),.dinb(w_asqrt39_19[0]),.dout(n4219),.clk(gclk));
	jxor g03980(.dina(w_n3920_0[0]),.dinb(w_n3907_23[1]),.dout(n4220),.clk(gclk));
	jand g03981(.dina(n4220),.dinb(w_asqrt36_30[1]),.dout(n4221),.clk(gclk));
	jxor g03982(.dina(n4221),.dinb(w_n3923_0[0]),.dout(n4222),.clk(gclk));
	jnot g03983(.din(w_n4222_0[1]),.dout(n4223),.clk(gclk));
	jand g03984(.dina(n4223),.dinb(n4219),.dout(n4224),.clk(gclk));
	jor g03985(.dina(w_n4224_0[1]),.dinb(w_n4218_0[1]),.dout(n4225),.clk(gclk));
	jand g03986(.dina(n4225),.dinb(w_asqrt40_22[0]),.dout(n4226),.clk(gclk));
	jnot g03987(.din(w_n3929_0[0]),.dout(n4227),.clk(gclk));
	jand g03988(.dina(n4227),.dinb(w_n3927_0[0]),.dout(n4228),.clk(gclk));
	jand g03989(.dina(n4228),.dinb(w_asqrt36_30[0]),.dout(n4229),.clk(gclk));
	jxor g03990(.dina(n4229),.dinb(w_n3937_0[0]),.dout(n4230),.clk(gclk));
	jnot g03991(.din(n4230),.dout(n4231),.clk(gclk));
	jor g03992(.dina(w_n4218_0[0]),.dinb(w_asqrt40_21[2]),.dout(n4232),.clk(gclk));
	jor g03993(.dina(n4232),.dinb(w_n4224_0[0]),.dout(n4233),.clk(gclk));
	jand g03994(.dina(w_n4233_0[1]),.dinb(w_n4231_0[1]),.dout(n4234),.clk(gclk));
	jor g03995(.dina(w_n4234_0[1]),.dinb(w_n4226_0[1]),.dout(n4235),.clk(gclk));
	jand g03996(.dina(w_n4235_0[2]),.dinb(w_asqrt41_19[2]),.dout(n4236),.clk(gclk));
	jor g03997(.dina(w_n4235_0[1]),.dinb(w_asqrt41_19[1]),.dout(n4237),.clk(gclk));
	jnot g03998(.din(w_n3944_0[0]),.dout(n4238),.clk(gclk));
	jxor g03999(.dina(w_n3939_0[0]),.dinb(w_n3371_23[2]),.dout(n4239),.clk(gclk));
	jand g04000(.dina(n4239),.dinb(w_asqrt36_29[2]),.dout(n4240),.clk(gclk));
	jxor g04001(.dina(n4240),.dinb(n4238),.dout(n4241),.clk(gclk));
	jand g04002(.dina(w_n4241_0[1]),.dinb(n4237),.dout(n4242),.clk(gclk));
	jor g04003(.dina(w_n4242_0[1]),.dinb(w_n4236_0[1]),.dout(n4243),.clk(gclk));
	jand g04004(.dina(n4243),.dinb(w_asqrt42_22[0]),.dout(n4244),.clk(gclk));
	jor g04005(.dina(w_n4236_0[0]),.dinb(w_asqrt42_21[2]),.dout(n4245),.clk(gclk));
	jor g04006(.dina(n4245),.dinb(w_n4242_0[0]),.dout(n4246),.clk(gclk));
	jnot g04007(.din(w_n3951_0[0]),.dout(n4247),.clk(gclk));
	jnot g04008(.din(w_n3953_0[0]),.dout(n4248),.clk(gclk));
	jand g04009(.dina(w_asqrt36_29[1]),.dinb(w_n3947_0[0]),.dout(n4249),.clk(gclk));
	jand g04010(.dina(w_n4249_0[1]),.dinb(n4248),.dout(n4250),.clk(gclk));
	jor g04011(.dina(n4250),.dinb(n4247),.dout(n4251),.clk(gclk));
	jnot g04012(.din(w_n3954_0[0]),.dout(n4252),.clk(gclk));
	jand g04013(.dina(w_n4249_0[0]),.dinb(n4252),.dout(n4253),.clk(gclk));
	jnot g04014(.din(n4253),.dout(n4254),.clk(gclk));
	jand g04015(.dina(n4254),.dinb(n4251),.dout(n4255),.clk(gclk));
	jand g04016(.dina(w_n4255_0[1]),.dinb(w_n4246_0[1]),.dout(n4256),.clk(gclk));
	jor g04017(.dina(n4256),.dinb(w_n4244_0[1]),.dout(n4257),.clk(gclk));
	jand g04018(.dina(w_n4257_0[2]),.dinb(w_asqrt43_19[2]),.dout(n4258),.clk(gclk));
	jor g04019(.dina(w_n4257_0[1]),.dinb(w_asqrt43_19[1]),.dout(n4259),.clk(gclk));
	jxor g04020(.dina(w_n3955_0[0]),.dinb(w_n2870_23[2]),.dout(n4260),.clk(gclk));
	jand g04021(.dina(n4260),.dinb(w_asqrt36_29[0]),.dout(n4261),.clk(gclk));
	jxor g04022(.dina(n4261),.dinb(w_n3960_0[0]),.dout(n4262),.clk(gclk));
	jand g04023(.dina(w_n4262_0[1]),.dinb(n4259),.dout(n4263),.clk(gclk));
	jor g04024(.dina(w_n4263_0[1]),.dinb(w_n4258_0[1]),.dout(n4264),.clk(gclk));
	jand g04025(.dina(n4264),.dinb(w_asqrt44_22[0]),.dout(n4265),.clk(gclk));
	jnot g04026(.din(w_n3966_0[0]),.dout(n4266),.clk(gclk));
	jand g04027(.dina(n4266),.dinb(w_n3964_0[0]),.dout(n4267),.clk(gclk));
	jand g04028(.dina(n4267),.dinb(w_asqrt36_28[2]),.dout(n4268),.clk(gclk));
	jxor g04029(.dina(n4268),.dinb(w_n3974_0[0]),.dout(n4269),.clk(gclk));
	jnot g04030(.din(n4269),.dout(n4270),.clk(gclk));
	jor g04031(.dina(w_n4258_0[0]),.dinb(w_asqrt44_21[2]),.dout(n4271),.clk(gclk));
	jor g04032(.dina(n4271),.dinb(w_n4263_0[0]),.dout(n4272),.clk(gclk));
	jand g04033(.dina(w_n4272_0[1]),.dinb(w_n4270_0[1]),.dout(n4273),.clk(gclk));
	jor g04034(.dina(w_n4273_0[1]),.dinb(w_n4265_0[1]),.dout(n4274),.clk(gclk));
	jand g04035(.dina(w_n4274_0[2]),.dinb(w_asqrt45_20[0]),.dout(n4275),.clk(gclk));
	jor g04036(.dina(w_n4274_0[1]),.dinb(w_asqrt45_19[2]),.dout(n4276),.clk(gclk));
	jxor g04037(.dina(w_n3976_0[0]),.dinb(w_n2420_24[1]),.dout(n4277),.clk(gclk));
	jand g04038(.dina(n4277),.dinb(w_asqrt36_28[1]),.dout(n4278),.clk(gclk));
	jxor g04039(.dina(n4278),.dinb(w_n3982_0[0]),.dout(n4279),.clk(gclk));
	jand g04040(.dina(w_n4279_0[1]),.dinb(n4276),.dout(n4280),.clk(gclk));
	jor g04041(.dina(w_n4280_0[1]),.dinb(w_n4275_0[1]),.dout(n4281),.clk(gclk));
	jand g04042(.dina(n4281),.dinb(w_asqrt46_22[0]),.dout(n4282),.clk(gclk));
	jor g04043(.dina(w_n4275_0[0]),.dinb(w_asqrt46_21[2]),.dout(n4283),.clk(gclk));
	jor g04044(.dina(n4283),.dinb(w_n4280_0[0]),.dout(n4284),.clk(gclk));
	jnot g04045(.din(w_n3990_0[0]),.dout(n4285),.clk(gclk));
	jnot g04046(.din(w_n3992_0[0]),.dout(n4286),.clk(gclk));
	jand g04047(.dina(w_asqrt36_28[0]),.dinb(w_n3986_0[0]),.dout(n4287),.clk(gclk));
	jand g04048(.dina(w_n4287_0[1]),.dinb(n4286),.dout(n4288),.clk(gclk));
	jor g04049(.dina(n4288),.dinb(n4285),.dout(n4289),.clk(gclk));
	jnot g04050(.din(w_n3993_0[0]),.dout(n4290),.clk(gclk));
	jand g04051(.dina(w_n4287_0[0]),.dinb(n4290),.dout(n4291),.clk(gclk));
	jnot g04052(.din(n4291),.dout(n4292),.clk(gclk));
	jand g04053(.dina(n4292),.dinb(n4289),.dout(n4293),.clk(gclk));
	jand g04054(.dina(w_n4293_0[1]),.dinb(w_n4284_0[1]),.dout(n4294),.clk(gclk));
	jor g04055(.dina(n4294),.dinb(w_n4282_0[1]),.dout(n4295),.clk(gclk));
	jand g04056(.dina(w_n4295_0[1]),.dinb(w_asqrt47_20[0]),.dout(n4296),.clk(gclk));
	jxor g04057(.dina(w_n3994_0[0]),.dinb(w_n2005_24[1]),.dout(n4297),.clk(gclk));
	jand g04058(.dina(n4297),.dinb(w_asqrt36_27[2]),.dout(n4298),.clk(gclk));
	jxor g04059(.dina(n4298),.dinb(w_n4001_0[0]),.dout(n4299),.clk(gclk));
	jnot g04060(.din(n4299),.dout(n4300),.clk(gclk));
	jor g04061(.dina(w_n4295_0[0]),.dinb(w_asqrt47_19[2]),.dout(n4301),.clk(gclk));
	jand g04062(.dina(w_n4301_0[1]),.dinb(w_n4300_0[1]),.dout(n4302),.clk(gclk));
	jor g04063(.dina(w_n4302_0[2]),.dinb(w_n4296_0[2]),.dout(n4303),.clk(gclk));
	jand g04064(.dina(n4303),.dinb(w_asqrt48_22[0]),.dout(n4304),.clk(gclk));
	jnot g04065(.din(w_n4006_0[0]),.dout(n4305),.clk(gclk));
	jand g04066(.dina(n4305),.dinb(w_n4004_0[0]),.dout(n4306),.clk(gclk));
	jand g04067(.dina(n4306),.dinb(w_asqrt36_27[1]),.dout(n4307),.clk(gclk));
	jxor g04068(.dina(n4307),.dinb(w_n4014_0[0]),.dout(n4308),.clk(gclk));
	jnot g04069(.din(n4308),.dout(n4309),.clk(gclk));
	jor g04070(.dina(w_n4296_0[1]),.dinb(w_asqrt48_21[2]),.dout(n4310),.clk(gclk));
	jor g04071(.dina(n4310),.dinb(w_n4302_0[1]),.dout(n4311),.clk(gclk));
	jand g04072(.dina(w_n4311_0[1]),.dinb(w_n4309_0[1]),.dout(n4312),.clk(gclk));
	jor g04073(.dina(w_n4312_0[1]),.dinb(w_n4304_0[1]),.dout(n4313),.clk(gclk));
	jand g04074(.dina(w_n4313_0[2]),.dinb(w_asqrt49_20[1]),.dout(n4314),.clk(gclk));
	jor g04075(.dina(w_n4313_0[1]),.dinb(w_asqrt49_20[0]),.dout(n4315),.clk(gclk));
	jnot g04076(.din(w_n4020_0[0]),.dout(n4316),.clk(gclk));
	jnot g04077(.din(w_n4021_0[0]),.dout(n4317),.clk(gclk));
	jand g04078(.dina(w_asqrt36_27[0]),.dinb(w_n4017_0[0]),.dout(n4318),.clk(gclk));
	jand g04079(.dina(w_n4318_0[1]),.dinb(n4317),.dout(n4319),.clk(gclk));
	jor g04080(.dina(n4319),.dinb(n4316),.dout(n4320),.clk(gclk));
	jnot g04081(.din(w_n4022_0[0]),.dout(n4321),.clk(gclk));
	jand g04082(.dina(w_n4318_0[0]),.dinb(n4321),.dout(n4322),.clk(gclk));
	jnot g04083(.din(n4322),.dout(n4323),.clk(gclk));
	jand g04084(.dina(n4323),.dinb(n4320),.dout(n4324),.clk(gclk));
	jand g04085(.dina(w_n4324_0[1]),.dinb(n4315),.dout(n4325),.clk(gclk));
	jor g04086(.dina(w_n4325_0[1]),.dinb(w_n4314_0[1]),.dout(n4326),.clk(gclk));
	jand g04087(.dina(n4326),.dinb(w_asqrt50_22[0]),.dout(n4327),.clk(gclk));
	jor g04088(.dina(w_n4314_0[0]),.dinb(w_asqrt50_21[2]),.dout(n4328),.clk(gclk));
	jor g04089(.dina(n4328),.dinb(w_n4325_0[0]),.dout(n4329),.clk(gclk));
	jnot g04090(.din(w_n4028_0[0]),.dout(n4330),.clk(gclk));
	jnot g04091(.din(w_n4030_0[0]),.dout(n4331),.clk(gclk));
	jand g04092(.dina(w_asqrt36_26[2]),.dinb(w_n4024_0[0]),.dout(n4332),.clk(gclk));
	jand g04093(.dina(w_n4332_0[1]),.dinb(n4331),.dout(n4333),.clk(gclk));
	jor g04094(.dina(n4333),.dinb(n4330),.dout(n4334),.clk(gclk));
	jnot g04095(.din(w_n4031_0[0]),.dout(n4335),.clk(gclk));
	jand g04096(.dina(w_n4332_0[0]),.dinb(n4335),.dout(n4336),.clk(gclk));
	jnot g04097(.din(n4336),.dout(n4337),.clk(gclk));
	jand g04098(.dina(n4337),.dinb(n4334),.dout(n4338),.clk(gclk));
	jand g04099(.dina(w_n4338_0[1]),.dinb(w_n4329_0[1]),.dout(n4339),.clk(gclk));
	jor g04100(.dina(n4339),.dinb(w_n4327_0[1]),.dout(n4340),.clk(gclk));
	jand g04101(.dina(w_n4340_0[1]),.dinb(w_asqrt51_20[1]),.dout(n4341),.clk(gclk));
	jxor g04102(.dina(w_n4032_0[0]),.dinb(w_n1312_25[0]),.dout(n4342),.clk(gclk));
	jand g04103(.dina(n4342),.dinb(w_asqrt36_26[1]),.dout(n4343),.clk(gclk));
	jxor g04104(.dina(n4343),.dinb(w_n4042_0[0]),.dout(n4344),.clk(gclk));
	jnot g04105(.din(n4344),.dout(n4345),.clk(gclk));
	jor g04106(.dina(w_n4340_0[0]),.dinb(w_asqrt51_20[0]),.dout(n4346),.clk(gclk));
	jand g04107(.dina(w_n4346_0[1]),.dinb(w_n4345_0[1]),.dout(n4347),.clk(gclk));
	jor g04108(.dina(w_n4347_0[2]),.dinb(w_n4341_0[2]),.dout(n4348),.clk(gclk));
	jand g04109(.dina(n4348),.dinb(w_asqrt52_22[0]),.dout(n4349),.clk(gclk));
	jnot g04110(.din(w_n4047_0[0]),.dout(n4350),.clk(gclk));
	jand g04111(.dina(n4350),.dinb(w_n4045_0[0]),.dout(n4351),.clk(gclk));
	jand g04112(.dina(n4351),.dinb(w_asqrt36_26[0]),.dout(n4352),.clk(gclk));
	jxor g04113(.dina(n4352),.dinb(w_n4055_0[0]),.dout(n4353),.clk(gclk));
	jnot g04114(.din(n4353),.dout(n4354),.clk(gclk));
	jor g04115(.dina(w_n4341_0[1]),.dinb(w_asqrt52_21[2]),.dout(n4355),.clk(gclk));
	jor g04116(.dina(n4355),.dinb(w_n4347_0[1]),.dout(n4356),.clk(gclk));
	jand g04117(.dina(w_n4356_0[1]),.dinb(w_n4354_0[1]),.dout(n4357),.clk(gclk));
	jor g04118(.dina(w_n4357_0[1]),.dinb(w_n4349_0[1]),.dout(n4358),.clk(gclk));
	jand g04119(.dina(w_n4358_0[2]),.dinb(w_asqrt53_20[2]),.dout(n4359),.clk(gclk));
	jor g04120(.dina(w_n4358_0[1]),.dinb(w_asqrt53_20[1]),.dout(n4360),.clk(gclk));
	jnot g04121(.din(w_n4061_0[0]),.dout(n4361),.clk(gclk));
	jnot g04122(.din(w_n4062_0[0]),.dout(n4362),.clk(gclk));
	jand g04123(.dina(w_asqrt36_25[2]),.dinb(w_n4058_0[0]),.dout(n4363),.clk(gclk));
	jand g04124(.dina(w_n4363_0[1]),.dinb(n4362),.dout(n4364),.clk(gclk));
	jor g04125(.dina(n4364),.dinb(n4361),.dout(n4365),.clk(gclk));
	jnot g04126(.din(w_n4063_0[0]),.dout(n4366),.clk(gclk));
	jand g04127(.dina(w_n4363_0[0]),.dinb(n4366),.dout(n4367),.clk(gclk));
	jnot g04128(.din(n4367),.dout(n4368),.clk(gclk));
	jand g04129(.dina(n4368),.dinb(n4365),.dout(n4369),.clk(gclk));
	jand g04130(.dina(w_n4369_0[1]),.dinb(n4360),.dout(n4370),.clk(gclk));
	jor g04131(.dina(w_n4370_0[1]),.dinb(w_n4359_0[1]),.dout(n4371),.clk(gclk));
	jand g04132(.dina(n4371),.dinb(w_asqrt54_22[0]),.dout(n4372),.clk(gclk));
	jor g04133(.dina(w_n4359_0[0]),.dinb(w_asqrt54_21[2]),.dout(n4373),.clk(gclk));
	jor g04134(.dina(n4373),.dinb(w_n4370_0[0]),.dout(n4374),.clk(gclk));
	jnot g04135(.din(w_n4069_0[0]),.dout(n4375),.clk(gclk));
	jnot g04136(.din(w_n4071_0[0]),.dout(n4376),.clk(gclk));
	jand g04137(.dina(w_asqrt36_25[1]),.dinb(w_n4065_0[0]),.dout(n4377),.clk(gclk));
	jand g04138(.dina(w_n4377_0[1]),.dinb(n4376),.dout(n4378),.clk(gclk));
	jor g04139(.dina(n4378),.dinb(n4375),.dout(n4379),.clk(gclk));
	jnot g04140(.din(w_n4072_0[0]),.dout(n4380),.clk(gclk));
	jand g04141(.dina(w_n4377_0[0]),.dinb(n4380),.dout(n4381),.clk(gclk));
	jnot g04142(.din(n4381),.dout(n4382),.clk(gclk));
	jand g04143(.dina(n4382),.dinb(n4379),.dout(n4383),.clk(gclk));
	jand g04144(.dina(w_n4383_0[1]),.dinb(w_n4374_0[1]),.dout(n4384),.clk(gclk));
	jor g04145(.dina(n4384),.dinb(w_n4372_0[1]),.dout(n4385),.clk(gclk));
	jand g04146(.dina(w_n4385_0[1]),.dinb(w_asqrt55_21[0]),.dout(n4386),.clk(gclk));
	jxor g04147(.dina(w_n4073_0[0]),.dinb(w_n791_26[0]),.dout(n4387),.clk(gclk));
	jand g04148(.dina(n4387),.dinb(w_asqrt36_25[0]),.dout(n4388),.clk(gclk));
	jxor g04149(.dina(n4388),.dinb(w_n4083_0[0]),.dout(n4389),.clk(gclk));
	jnot g04150(.din(n4389),.dout(n4390),.clk(gclk));
	jor g04151(.dina(w_n4385_0[0]),.dinb(w_asqrt55_20[2]),.dout(n4391),.clk(gclk));
	jand g04152(.dina(w_n4391_0[1]),.dinb(w_n4390_0[1]),.dout(n4392),.clk(gclk));
	jor g04153(.dina(w_n4392_0[2]),.dinb(w_n4386_0[2]),.dout(n4393),.clk(gclk));
	jand g04154(.dina(n4393),.dinb(w_asqrt56_22[0]),.dout(n4394),.clk(gclk));
	jnot g04155(.din(w_n4088_0[0]),.dout(n4395),.clk(gclk));
	jand g04156(.dina(n4395),.dinb(w_n4086_0[0]),.dout(n4396),.clk(gclk));
	jand g04157(.dina(n4396),.dinb(w_asqrt36_24[2]),.dout(n4397),.clk(gclk));
	jxor g04158(.dina(n4397),.dinb(w_n4096_0[0]),.dout(n4398),.clk(gclk));
	jnot g04159(.din(n4398),.dout(n4399),.clk(gclk));
	jor g04160(.dina(w_n4386_0[1]),.dinb(w_asqrt56_21[2]),.dout(n4400),.clk(gclk));
	jor g04161(.dina(n4400),.dinb(w_n4392_0[1]),.dout(n4401),.clk(gclk));
	jand g04162(.dina(w_n4401_0[1]),.dinb(w_n4399_0[1]),.dout(n4402),.clk(gclk));
	jor g04163(.dina(w_n4402_0[1]),.dinb(w_n4394_0[1]),.dout(n4403),.clk(gclk));
	jand g04164(.dina(w_n4403_0[2]),.dinb(w_asqrt57_21[1]),.dout(n4404),.clk(gclk));
	jor g04165(.dina(w_n4403_0[1]),.dinb(w_asqrt57_21[0]),.dout(n4405),.clk(gclk));
	jnot g04166(.din(w_n4102_0[0]),.dout(n4406),.clk(gclk));
	jnot g04167(.din(w_n4103_0[0]),.dout(n4407),.clk(gclk));
	jand g04168(.dina(w_asqrt36_24[1]),.dinb(w_n4099_0[0]),.dout(n4408),.clk(gclk));
	jand g04169(.dina(w_n4408_0[1]),.dinb(n4407),.dout(n4409),.clk(gclk));
	jor g04170(.dina(n4409),.dinb(n4406),.dout(n4410),.clk(gclk));
	jnot g04171(.din(w_n4104_0[0]),.dout(n4411),.clk(gclk));
	jand g04172(.dina(w_n4408_0[0]),.dinb(n4411),.dout(n4412),.clk(gclk));
	jnot g04173(.din(n4412),.dout(n4413),.clk(gclk));
	jand g04174(.dina(n4413),.dinb(n4410),.dout(n4414),.clk(gclk));
	jand g04175(.dina(w_n4414_0[1]),.dinb(n4405),.dout(n4415),.clk(gclk));
	jor g04176(.dina(w_n4415_0[1]),.dinb(w_n4404_0[1]),.dout(n4416),.clk(gclk));
	jand g04177(.dina(n4416),.dinb(w_asqrt58_22[0]),.dout(n4417),.clk(gclk));
	jor g04178(.dina(w_n4404_0[0]),.dinb(w_asqrt58_21[2]),.dout(n4418),.clk(gclk));
	jor g04179(.dina(n4418),.dinb(w_n4415_0[0]),.dout(n4419),.clk(gclk));
	jnot g04180(.din(w_n4110_0[0]),.dout(n4420),.clk(gclk));
	jnot g04181(.din(w_n4112_0[0]),.dout(n4421),.clk(gclk));
	jand g04182(.dina(w_asqrt36_24[0]),.dinb(w_n4106_0[0]),.dout(n4422),.clk(gclk));
	jand g04183(.dina(w_n4422_0[1]),.dinb(n4421),.dout(n4423),.clk(gclk));
	jor g04184(.dina(n4423),.dinb(n4420),.dout(n4424),.clk(gclk));
	jnot g04185(.din(w_n4113_0[0]),.dout(n4425),.clk(gclk));
	jand g04186(.dina(w_n4422_0[0]),.dinb(n4425),.dout(n4426),.clk(gclk));
	jnot g04187(.din(n4426),.dout(n4427),.clk(gclk));
	jand g04188(.dina(n4427),.dinb(n4424),.dout(n4428),.clk(gclk));
	jand g04189(.dina(w_n4428_0[1]),.dinb(w_n4419_0[1]),.dout(n4429),.clk(gclk));
	jor g04190(.dina(n4429),.dinb(w_n4417_0[1]),.dout(n4430),.clk(gclk));
	jand g04191(.dina(w_n4430_0[1]),.dinb(w_asqrt59_21[2]),.dout(n4431),.clk(gclk));
	jxor g04192(.dina(w_n4114_0[0]),.dinb(w_n425_26[2]),.dout(n4432),.clk(gclk));
	jand g04193(.dina(n4432),.dinb(w_asqrt36_23[2]),.dout(n4433),.clk(gclk));
	jxor g04194(.dina(n4433),.dinb(w_n4124_0[0]),.dout(n4434),.clk(gclk));
	jnot g04195(.din(n4434),.dout(n4435),.clk(gclk));
	jor g04196(.dina(w_n4430_0[0]),.dinb(w_asqrt59_21[1]),.dout(n4436),.clk(gclk));
	jand g04197(.dina(w_n4436_0[1]),.dinb(w_n4435_0[1]),.dout(n4437),.clk(gclk));
	jor g04198(.dina(w_n4437_0[2]),.dinb(w_n4431_0[2]),.dout(n4438),.clk(gclk));
	jand g04199(.dina(n4438),.dinb(w_asqrt60_21[2]),.dout(n4439),.clk(gclk));
	jnot g04200(.din(w_n4129_0[0]),.dout(n4440),.clk(gclk));
	jand g04201(.dina(n4440),.dinb(w_n4127_0[0]),.dout(n4441),.clk(gclk));
	jand g04202(.dina(n4441),.dinb(w_asqrt36_23[1]),.dout(n4442),.clk(gclk));
	jxor g04203(.dina(n4442),.dinb(w_n4137_0[0]),.dout(n4443),.clk(gclk));
	jnot g04204(.din(n4443),.dout(n4444),.clk(gclk));
	jor g04205(.dina(w_n4431_0[1]),.dinb(w_asqrt60_21[1]),.dout(n4445),.clk(gclk));
	jor g04206(.dina(n4445),.dinb(w_n4437_0[1]),.dout(n4446),.clk(gclk));
	jand g04207(.dina(w_n4446_0[1]),.dinb(w_n4444_0[1]),.dout(n4447),.clk(gclk));
	jor g04208(.dina(w_n4447_0[1]),.dinb(w_n4439_0[1]),.dout(n4448),.clk(gclk));
	jand g04209(.dina(w_n4448_0[2]),.dinb(w_asqrt61_22[0]),.dout(n4449),.clk(gclk));
	jor g04210(.dina(w_n4448_0[1]),.dinb(w_asqrt61_21[2]),.dout(n4450),.clk(gclk));
	jnot g04211(.din(w_n4143_0[0]),.dout(n4451),.clk(gclk));
	jnot g04212(.din(w_n4144_0[0]),.dout(n4452),.clk(gclk));
	jand g04213(.dina(w_asqrt36_23[0]),.dinb(w_n4140_0[0]),.dout(n4453),.clk(gclk));
	jand g04214(.dina(w_n4453_0[1]),.dinb(n4452),.dout(n4454),.clk(gclk));
	jor g04215(.dina(n4454),.dinb(n4451),.dout(n4455),.clk(gclk));
	jnot g04216(.din(w_n4145_0[0]),.dout(n4456),.clk(gclk));
	jand g04217(.dina(w_n4453_0[0]),.dinb(n4456),.dout(n4457),.clk(gclk));
	jnot g04218(.din(n4457),.dout(n4458),.clk(gclk));
	jand g04219(.dina(n4458),.dinb(n4455),.dout(n4459),.clk(gclk));
	jand g04220(.dina(w_n4459_0[1]),.dinb(n4450),.dout(n4460),.clk(gclk));
	jor g04221(.dina(w_n4460_0[1]),.dinb(w_n4449_0[1]),.dout(n4461),.clk(gclk));
	jand g04222(.dina(n4461),.dinb(w_asqrt62_22[0]),.dout(n4462),.clk(gclk));
	jor g04223(.dina(w_n4449_0[0]),.dinb(w_asqrt62_21[2]),.dout(n4463),.clk(gclk));
	jor g04224(.dina(n4463),.dinb(w_n4460_0[0]),.dout(n4464),.clk(gclk));
	jnot g04225(.din(w_n4151_0[0]),.dout(n4465),.clk(gclk));
	jnot g04226(.din(w_n4153_0[0]),.dout(n4466),.clk(gclk));
	jand g04227(.dina(w_asqrt36_22[2]),.dinb(w_n4147_0[0]),.dout(n4467),.clk(gclk));
	jand g04228(.dina(w_n4467_0[1]),.dinb(n4466),.dout(n4468),.clk(gclk));
	jor g04229(.dina(n4468),.dinb(n4465),.dout(n4469),.clk(gclk));
	jnot g04230(.din(w_n4154_0[0]),.dout(n4470),.clk(gclk));
	jand g04231(.dina(w_n4467_0[0]),.dinb(n4470),.dout(n4471),.clk(gclk));
	jnot g04232(.din(n4471),.dout(n4472),.clk(gclk));
	jand g04233(.dina(n4472),.dinb(n4469),.dout(n4473),.clk(gclk));
	jand g04234(.dina(w_n4473_0[1]),.dinb(w_n4464_0[1]),.dout(n4474),.clk(gclk));
	jor g04235(.dina(n4474),.dinb(w_n4462_0[1]),.dout(n4475),.clk(gclk));
	jxor g04236(.dina(w_n4155_0[0]),.dinb(w_n199_32[2]),.dout(n4476),.clk(gclk));
	jand g04237(.dina(n4476),.dinb(w_asqrt36_22[1]),.dout(n4477),.clk(gclk));
	jxor g04238(.dina(n4477),.dinb(w_n4165_0[0]),.dout(n4478),.clk(gclk));
	jnot g04239(.din(w_n4167_0[0]),.dout(n4479),.clk(gclk));
	jand g04240(.dina(w_asqrt36_22[0]),.dinb(w_n4174_0[1]),.dout(n4480),.clk(gclk));
	jand g04241(.dina(w_n4480_0[1]),.dinb(w_n4479_0[2]),.dout(n4481),.clk(gclk));
	jor g04242(.dina(n4481),.dinb(w_n4182_0[0]),.dout(n4482),.clk(gclk));
	jor g04243(.dina(n4482),.dinb(w_n4478_0[1]),.dout(n4483),.clk(gclk));
	jnot g04244(.din(n4483),.dout(n4484),.clk(gclk));
	jand g04245(.dina(n4484),.dinb(w_n4475_1[2]),.dout(n4485),.clk(gclk));
	jor g04246(.dina(n4485),.dinb(w_asqrt63_11[2]),.dout(n4486),.clk(gclk));
	jnot g04247(.din(w_n4478_0[0]),.dout(n4487),.clk(gclk));
	jor g04248(.dina(w_n4487_0[2]),.dinb(w_n4475_1[1]),.dout(n4488),.clk(gclk));
	jor g04249(.dina(w_n4480_0[0]),.dinb(w_n4479_0[1]),.dout(n4489),.clk(gclk));
	jand g04250(.dina(w_n4174_0[0]),.dinb(w_n4479_0[0]),.dout(n4490),.clk(gclk));
	jor g04251(.dina(n4490),.dinb(w_n194_31[2]),.dout(n4491),.clk(gclk));
	jnot g04252(.din(n4491),.dout(n4492),.clk(gclk));
	jand g04253(.dina(n4492),.dinb(n4489),.dout(n4493),.clk(gclk));
	jnot g04254(.din(w_asqrt36_21[2]),.dout(n4494),.clk(gclk));
	jnot g04255(.din(w_n4493_0[1]),.dout(n4497),.clk(gclk));
	jand g04256(.dina(n4497),.dinb(w_n4488_0[1]),.dout(n4498),.clk(gclk));
	jand g04257(.dina(n4498),.dinb(w_n4486_0[1]),.dout(n4499),.clk(gclk));
	jnot g04258(.din(w_n4499_31[1]),.dout(asqrt_fa_36),.clk(gclk));
	jor g04259(.dina(w_n4499_31[0]),.dinb(w_n4193_1[0]),.dout(n4501),.clk(gclk));
	jnot g04260(.din(w_a68_0[1]),.dout(n4502),.clk(gclk));
	jnot g04261(.din(a[69]),.dout(n4503),.clk(gclk));
	jand g04262(.dina(w_n4193_0[2]),.dinb(w_n4503_0[2]),.dout(n4504),.clk(gclk));
	jand g04263(.dina(n4504),.dinb(w_n4502_1[1]),.dout(n4505),.clk(gclk));
	jnot g04264(.din(n4505),.dout(n4506),.clk(gclk));
	jand g04265(.dina(n4506),.dinb(n4501),.dout(n4507),.clk(gclk));
	jor g04266(.dina(w_n4507_0[2]),.dinb(w_n4494_23[1]),.dout(n4508),.clk(gclk));
	jor g04267(.dina(w_n4499_30[2]),.dinb(w_a70_0[0]),.dout(n4509),.clk(gclk));
	jxor g04268(.dina(w_n4509_0[1]),.dinb(w_n4194_0[0]),.dout(n4510),.clk(gclk));
	jand g04269(.dina(w_n4507_0[1]),.dinb(w_n4494_23[0]),.dout(n4511),.clk(gclk));
	jor g04270(.dina(n4511),.dinb(w_n4510_0[1]),.dout(n4512),.clk(gclk));
	jand g04271(.dina(w_n4512_0[1]),.dinb(w_n4508_0[1]),.dout(n4513),.clk(gclk));
	jor g04272(.dina(n4513),.dinb(w_n3912_26[0]),.dout(n4514),.clk(gclk));
	jand g04273(.dina(w_n4508_0[0]),.dinb(w_n3912_25[2]),.dout(n4515),.clk(gclk));
	jand g04274(.dina(n4515),.dinb(w_n4512_0[0]),.dout(n4516),.clk(gclk));
	jor g04275(.dina(w_n4509_0[0]),.dinb(w_a71_0[0]),.dout(n4517),.clk(gclk));
	jnot g04276(.din(w_n4486_0[0]),.dout(n4518),.clk(gclk));
	jnot g04277(.din(w_n4488_0[0]),.dout(n4519),.clk(gclk));
	jor g04278(.dina(w_n4493_0[0]),.dinb(w_n4494_22[2]),.dout(n4520),.clk(gclk));
	jor g04279(.dina(n4520),.dinb(w_n4519_0[1]),.dout(n4521),.clk(gclk));
	jor g04280(.dina(n4521),.dinb(n4518),.dout(n4522),.clk(gclk));
	jand g04281(.dina(n4522),.dinb(n4517),.dout(n4523),.clk(gclk));
	jxor g04282(.dina(n4523),.dinb(w_n3915_0[1]),.dout(n4524),.clk(gclk));
	jor g04283(.dina(w_n4524_0[1]),.dinb(w_n4516_0[1]),.dout(n4525),.clk(gclk));
	jand g04284(.dina(n4525),.dinb(w_n4514_0[1]),.dout(n4526),.clk(gclk));
	jor g04285(.dina(w_n4526_0[2]),.dinb(w_n3907_23[0]),.dout(n4527),.clk(gclk));
	jand g04286(.dina(w_n4526_0[1]),.dinb(w_n3907_22[2]),.dout(n4528),.clk(gclk));
	jxor g04287(.dina(w_n4197_0[0]),.dinb(w_n3912_25[1]),.dout(n4529),.clk(gclk));
	jor g04288(.dina(n4529),.dinb(w_n4499_30[1]),.dout(n4530),.clk(gclk));
	jxor g04289(.dina(n4530),.dinb(w_n4200_0[0]),.dout(n4531),.clk(gclk));
	jor g04290(.dina(w_n4531_0[1]),.dinb(n4528),.dout(n4532),.clk(gclk));
	jand g04291(.dina(w_n4532_0[1]),.dinb(w_n4527_0[1]),.dout(n4533),.clk(gclk));
	jor g04292(.dina(n4533),.dinb(w_n3376_26[2]),.dout(n4534),.clk(gclk));
	jnot g04293(.din(w_n4206_0[0]),.dout(n4535),.clk(gclk));
	jor g04294(.dina(n4535),.dinb(w_n4204_0[0]),.dout(n4536),.clk(gclk));
	jor g04295(.dina(n4536),.dinb(w_n4499_30[0]),.dout(n4537),.clk(gclk));
	jxor g04296(.dina(n4537),.dinb(w_n4215_0[0]),.dout(n4538),.clk(gclk));
	jand g04297(.dina(w_n4527_0[0]),.dinb(w_n3376_26[1]),.dout(n4539),.clk(gclk));
	jand g04298(.dina(n4539),.dinb(w_n4532_0[0]),.dout(n4540),.clk(gclk));
	jor g04299(.dina(w_n4540_0[1]),.dinb(w_n4538_0[1]),.dout(n4541),.clk(gclk));
	jand g04300(.dina(w_n4541_0[1]),.dinb(w_n4534_0[1]),.dout(n4542),.clk(gclk));
	jor g04301(.dina(w_n4542_0[2]),.dinb(w_n3371_23[1]),.dout(n4543),.clk(gclk));
	jand g04302(.dina(w_n4542_0[1]),.dinb(w_n3371_23[0]),.dout(n4544),.clk(gclk));
	jxor g04303(.dina(w_n4217_0[0]),.dinb(w_n3376_26[0]),.dout(n4545),.clk(gclk));
	jor g04304(.dina(n4545),.dinb(w_n4499_29[2]),.dout(n4546),.clk(gclk));
	jxor g04305(.dina(n4546),.dinb(w_n4222_0[0]),.dout(n4547),.clk(gclk));
	jnot g04306(.din(w_n4547_0[1]),.dout(n4548),.clk(gclk));
	jor g04307(.dina(n4548),.dinb(n4544),.dout(n4549),.clk(gclk));
	jand g04308(.dina(w_n4549_0[1]),.dinb(w_n4543_0[1]),.dout(n4550),.clk(gclk));
	jor g04309(.dina(n4550),.dinb(w_n2875_26[1]),.dout(n4551),.clk(gclk));
	jand g04310(.dina(w_n4543_0[0]),.dinb(w_n2875_26[0]),.dout(n4552),.clk(gclk));
	jand g04311(.dina(n4552),.dinb(w_n4549_0[0]),.dout(n4553),.clk(gclk));
	jnot g04312(.din(w_n4226_0[0]),.dout(n4554),.clk(gclk));
	jand g04313(.dina(w_asqrt35_22[1]),.dinb(n4554),.dout(n4555),.clk(gclk));
	jand g04314(.dina(w_n4555_0[1]),.dinb(w_n4233_0[0]),.dout(n4556),.clk(gclk));
	jor g04315(.dina(n4556),.dinb(w_n4231_0[0]),.dout(n4557),.clk(gclk));
	jand g04316(.dina(w_n4555_0[0]),.dinb(w_n4234_0[0]),.dout(n4558),.clk(gclk));
	jnot g04317(.din(n4558),.dout(n4559),.clk(gclk));
	jand g04318(.dina(n4559),.dinb(n4557),.dout(n4560),.clk(gclk));
	jnot g04319(.din(n4560),.dout(n4561),.clk(gclk));
	jor g04320(.dina(w_n4561_0[1]),.dinb(w_n4553_0[1]),.dout(n4562),.clk(gclk));
	jand g04321(.dina(n4562),.dinb(w_n4551_0[1]),.dout(n4563),.clk(gclk));
	jor g04322(.dina(w_n4563_0[2]),.dinb(w_n2870_23[1]),.dout(n4564),.clk(gclk));
	jand g04323(.dina(w_n4563_0[1]),.dinb(w_n2870_23[0]),.dout(n4565),.clk(gclk));
	jnot g04324(.din(w_n4241_0[0]),.dout(n4566),.clk(gclk));
	jxor g04325(.dina(w_n4235_0[0]),.dinb(w_n2875_25[2]),.dout(n4567),.clk(gclk));
	jor g04326(.dina(n4567),.dinb(w_n4499_29[1]),.dout(n4568),.clk(gclk));
	jxor g04327(.dina(n4568),.dinb(n4566),.dout(n4569),.clk(gclk));
	jnot g04328(.din(w_n4569_0[1]),.dout(n4570),.clk(gclk));
	jor g04329(.dina(n4570),.dinb(n4565),.dout(n4571),.clk(gclk));
	jand g04330(.dina(w_n4571_0[1]),.dinb(w_n4564_0[1]),.dout(n4572),.clk(gclk));
	jor g04331(.dina(n4572),.dinb(w_n2425_26[2]),.dout(n4573),.clk(gclk));
	jnot g04332(.din(w_n4246_0[0]),.dout(n4574),.clk(gclk));
	jor g04333(.dina(n4574),.dinb(w_n4244_0[0]),.dout(n4575),.clk(gclk));
	jor g04334(.dina(n4575),.dinb(w_n4499_29[0]),.dout(n4576),.clk(gclk));
	jxor g04335(.dina(n4576),.dinb(w_n4255_0[0]),.dout(n4577),.clk(gclk));
	jand g04336(.dina(w_n4564_0[0]),.dinb(w_n2425_26[1]),.dout(n4578),.clk(gclk));
	jand g04337(.dina(n4578),.dinb(w_n4571_0[0]),.dout(n4579),.clk(gclk));
	jor g04338(.dina(w_n4579_0[1]),.dinb(w_n4577_0[1]),.dout(n4580),.clk(gclk));
	jand g04339(.dina(w_n4580_0[1]),.dinb(w_n4573_0[1]),.dout(n4581),.clk(gclk));
	jor g04340(.dina(w_n4581_0[2]),.dinb(w_n2420_24[0]),.dout(n4582),.clk(gclk));
	jand g04341(.dina(w_n4581_0[1]),.dinb(w_n2420_23[2]),.dout(n4583),.clk(gclk));
	jnot g04342(.din(w_n4262_0[0]),.dout(n4584),.clk(gclk));
	jxor g04343(.dina(w_n4257_0[0]),.dinb(w_n2425_26[0]),.dout(n4585),.clk(gclk));
	jor g04344(.dina(n4585),.dinb(w_n4499_28[2]),.dout(n4586),.clk(gclk));
	jxor g04345(.dina(n4586),.dinb(n4584),.dout(n4587),.clk(gclk));
	jnot g04346(.din(n4587),.dout(n4588),.clk(gclk));
	jor g04347(.dina(w_n4588_0[1]),.dinb(n4583),.dout(n4589),.clk(gclk));
	jand g04348(.dina(w_n4589_0[1]),.dinb(w_n4582_0[1]),.dout(n4590),.clk(gclk));
	jor g04349(.dina(n4590),.dinb(w_n2010_26[1]),.dout(n4591),.clk(gclk));
	jand g04350(.dina(w_n4582_0[0]),.dinb(w_n2010_26[0]),.dout(n4592),.clk(gclk));
	jand g04351(.dina(n4592),.dinb(w_n4589_0[0]),.dout(n4593),.clk(gclk));
	jnot g04352(.din(w_n4265_0[0]),.dout(n4594),.clk(gclk));
	jand g04353(.dina(w_asqrt35_22[0]),.dinb(n4594),.dout(n4595),.clk(gclk));
	jand g04354(.dina(w_n4595_0[1]),.dinb(w_n4272_0[0]),.dout(n4596),.clk(gclk));
	jor g04355(.dina(n4596),.dinb(w_n4270_0[0]),.dout(n4597),.clk(gclk));
	jand g04356(.dina(w_n4595_0[0]),.dinb(w_n4273_0[0]),.dout(n4598),.clk(gclk));
	jnot g04357(.din(n4598),.dout(n4599),.clk(gclk));
	jand g04358(.dina(n4599),.dinb(n4597),.dout(n4600),.clk(gclk));
	jnot g04359(.din(n4600),.dout(n4601),.clk(gclk));
	jor g04360(.dina(w_n4601_0[1]),.dinb(w_n4593_0[1]),.dout(n4602),.clk(gclk));
	jand g04361(.dina(n4602),.dinb(w_n4591_0[1]),.dout(n4603),.clk(gclk));
	jor g04362(.dina(w_n4603_0[1]),.dinb(w_n2005_24[0]),.dout(n4604),.clk(gclk));
	jxor g04363(.dina(w_n4274_0[0]),.dinb(w_n2010_25[2]),.dout(n4605),.clk(gclk));
	jor g04364(.dina(n4605),.dinb(w_n4499_28[1]),.dout(n4606),.clk(gclk));
	jxor g04365(.dina(n4606),.dinb(w_n4279_0[0]),.dout(n4607),.clk(gclk));
	jand g04366(.dina(w_n4603_0[0]),.dinb(w_n2005_23[2]),.dout(n4608),.clk(gclk));
	jor g04367(.dina(w_n4608_0[1]),.dinb(w_n4607_0[1]),.dout(n4609),.clk(gclk));
	jand g04368(.dina(w_n4609_0[2]),.dinb(w_n4604_0[2]),.dout(n4610),.clk(gclk));
	jor g04369(.dina(n4610),.dinb(w_n1646_27[0]),.dout(n4611),.clk(gclk));
	jnot g04370(.din(w_n4284_0[0]),.dout(n4612),.clk(gclk));
	jor g04371(.dina(n4612),.dinb(w_n4282_0[0]),.dout(n4613),.clk(gclk));
	jor g04372(.dina(n4613),.dinb(w_n4499_28[0]),.dout(n4614),.clk(gclk));
	jxor g04373(.dina(n4614),.dinb(w_n4293_0[0]),.dout(n4615),.clk(gclk));
	jand g04374(.dina(w_n4604_0[1]),.dinb(w_n1646_26[2]),.dout(n4616),.clk(gclk));
	jand g04375(.dina(n4616),.dinb(w_n4609_0[1]),.dout(n4617),.clk(gclk));
	jor g04376(.dina(w_n4617_0[1]),.dinb(w_n4615_0[1]),.dout(n4618),.clk(gclk));
	jand g04377(.dina(w_n4618_0[1]),.dinb(w_n4611_0[1]),.dout(n4619),.clk(gclk));
	jor g04378(.dina(w_n4619_0[2]),.dinb(w_n1641_24[2]),.dout(n4620),.clk(gclk));
	jand g04379(.dina(w_n4619_0[1]),.dinb(w_n1641_24[1]),.dout(n4621),.clk(gclk));
	jnot g04380(.din(w_n4296_0[0]),.dout(n4622),.clk(gclk));
	jand g04381(.dina(w_asqrt35_21[2]),.dinb(n4622),.dout(n4623),.clk(gclk));
	jand g04382(.dina(w_n4623_0[1]),.dinb(w_n4301_0[0]),.dout(n4624),.clk(gclk));
	jor g04383(.dina(n4624),.dinb(w_n4300_0[0]),.dout(n4625),.clk(gclk));
	jand g04384(.dina(w_n4623_0[0]),.dinb(w_n4302_0[0]),.dout(n4626),.clk(gclk));
	jnot g04385(.din(n4626),.dout(n4627),.clk(gclk));
	jand g04386(.dina(n4627),.dinb(n4625),.dout(n4628),.clk(gclk));
	jnot g04387(.din(n4628),.dout(n4629),.clk(gclk));
	jor g04388(.dina(w_n4629_0[1]),.dinb(n4621),.dout(n4630),.clk(gclk));
	jand g04389(.dina(w_n4630_0[1]),.dinb(w_n4620_0[1]),.dout(n4631),.clk(gclk));
	jor g04390(.dina(n4631),.dinb(w_n1317_27[0]),.dout(n4632),.clk(gclk));
	jand g04391(.dina(w_n4620_0[0]),.dinb(w_n1317_26[2]),.dout(n4633),.clk(gclk));
	jand g04392(.dina(n4633),.dinb(w_n4630_0[0]),.dout(n4634),.clk(gclk));
	jnot g04393(.din(w_n4304_0[0]),.dout(n4635),.clk(gclk));
	jand g04394(.dina(w_asqrt35_21[1]),.dinb(n4635),.dout(n4636),.clk(gclk));
	jand g04395(.dina(w_n4636_0[1]),.dinb(w_n4311_0[0]),.dout(n4637),.clk(gclk));
	jor g04396(.dina(n4637),.dinb(w_n4309_0[0]),.dout(n4638),.clk(gclk));
	jand g04397(.dina(w_n4636_0[0]),.dinb(w_n4312_0[0]),.dout(n4639),.clk(gclk));
	jnot g04398(.din(n4639),.dout(n4640),.clk(gclk));
	jand g04399(.dina(n4640),.dinb(n4638),.dout(n4641),.clk(gclk));
	jnot g04400(.din(n4641),.dout(n4642),.clk(gclk));
	jor g04401(.dina(w_n4642_0[1]),.dinb(w_n4634_0[1]),.dout(n4643),.clk(gclk));
	jand g04402(.dina(n4643),.dinb(w_n4632_0[1]),.dout(n4644),.clk(gclk));
	jor g04403(.dina(w_n4644_0[1]),.dinb(w_n1312_24[2]),.dout(n4645),.clk(gclk));
	jxor g04404(.dina(w_n4313_0[0]),.dinb(w_n1317_26[1]),.dout(n4646),.clk(gclk));
	jor g04405(.dina(n4646),.dinb(w_n4499_27[2]),.dout(n4647),.clk(gclk));
	jxor g04406(.dina(n4647),.dinb(w_n4324_0[0]),.dout(n4648),.clk(gclk));
	jand g04407(.dina(w_n4644_0[0]),.dinb(w_n1312_24[1]),.dout(n4649),.clk(gclk));
	jor g04408(.dina(w_n4649_0[1]),.dinb(w_n4648_0[1]),.dout(n4650),.clk(gclk));
	jand g04409(.dina(w_n4650_0[2]),.dinb(w_n4645_0[2]),.dout(n4651),.clk(gclk));
	jor g04410(.dina(n4651),.dinb(w_n1039_27[1]),.dout(n4652),.clk(gclk));
	jnot g04411(.din(w_n4329_0[0]),.dout(n4653),.clk(gclk));
	jor g04412(.dina(n4653),.dinb(w_n4327_0[0]),.dout(n4654),.clk(gclk));
	jor g04413(.dina(n4654),.dinb(w_n4499_27[1]),.dout(n4655),.clk(gclk));
	jxor g04414(.dina(n4655),.dinb(w_n4338_0[0]),.dout(n4656),.clk(gclk));
	jand g04415(.dina(w_n4645_0[1]),.dinb(w_n1039_27[0]),.dout(n4657),.clk(gclk));
	jand g04416(.dina(n4657),.dinb(w_n4650_0[1]),.dout(n4658),.clk(gclk));
	jor g04417(.dina(w_n4658_0[1]),.dinb(w_n4656_0[1]),.dout(n4659),.clk(gclk));
	jand g04418(.dina(w_n4659_0[1]),.dinb(w_n4652_0[1]),.dout(n4660),.clk(gclk));
	jor g04419(.dina(w_n4660_0[2]),.dinb(w_n1034_25[2]),.dout(n4661),.clk(gclk));
	jand g04420(.dina(w_n4660_0[1]),.dinb(w_n1034_25[1]),.dout(n4662),.clk(gclk));
	jnot g04421(.din(w_n4341_0[0]),.dout(n4663),.clk(gclk));
	jand g04422(.dina(w_asqrt35_21[0]),.dinb(n4663),.dout(n4664),.clk(gclk));
	jand g04423(.dina(w_n4664_0[1]),.dinb(w_n4346_0[0]),.dout(n4665),.clk(gclk));
	jor g04424(.dina(n4665),.dinb(w_n4345_0[0]),.dout(n4666),.clk(gclk));
	jand g04425(.dina(w_n4664_0[0]),.dinb(w_n4347_0[0]),.dout(n4667),.clk(gclk));
	jnot g04426(.din(n4667),.dout(n4668),.clk(gclk));
	jand g04427(.dina(n4668),.dinb(n4666),.dout(n4669),.clk(gclk));
	jnot g04428(.din(n4669),.dout(n4670),.clk(gclk));
	jor g04429(.dina(w_n4670_0[1]),.dinb(n4662),.dout(n4671),.clk(gclk));
	jand g04430(.dina(w_n4671_0[1]),.dinb(w_n4661_0[1]),.dout(n4672),.clk(gclk));
	jor g04431(.dina(n4672),.dinb(w_n796_27[1]),.dout(n4673),.clk(gclk));
	jand g04432(.dina(w_n4661_0[0]),.dinb(w_n796_27[0]),.dout(n4674),.clk(gclk));
	jand g04433(.dina(n4674),.dinb(w_n4671_0[0]),.dout(n4675),.clk(gclk));
	jnot g04434(.din(w_n4349_0[0]),.dout(n4676),.clk(gclk));
	jand g04435(.dina(w_asqrt35_20[2]),.dinb(n4676),.dout(n4677),.clk(gclk));
	jand g04436(.dina(w_n4677_0[1]),.dinb(w_n4356_0[0]),.dout(n4678),.clk(gclk));
	jor g04437(.dina(n4678),.dinb(w_n4354_0[0]),.dout(n4679),.clk(gclk));
	jand g04438(.dina(w_n4677_0[0]),.dinb(w_n4357_0[0]),.dout(n4680),.clk(gclk));
	jnot g04439(.din(n4680),.dout(n4681),.clk(gclk));
	jand g04440(.dina(n4681),.dinb(n4679),.dout(n4682),.clk(gclk));
	jnot g04441(.din(n4682),.dout(n4683),.clk(gclk));
	jor g04442(.dina(w_n4683_0[1]),.dinb(w_n4675_0[1]),.dout(n4684),.clk(gclk));
	jand g04443(.dina(n4684),.dinb(w_n4673_0[1]),.dout(n4685),.clk(gclk));
	jor g04444(.dina(w_n4685_0[1]),.dinb(w_n791_25[2]),.dout(n4686),.clk(gclk));
	jxor g04445(.dina(w_n4358_0[0]),.dinb(w_n796_26[2]),.dout(n4687),.clk(gclk));
	jor g04446(.dina(n4687),.dinb(w_n4499_27[0]),.dout(n4688),.clk(gclk));
	jxor g04447(.dina(n4688),.dinb(w_n4369_0[0]),.dout(n4689),.clk(gclk));
	jand g04448(.dina(w_n4685_0[0]),.dinb(w_n791_25[1]),.dout(n4690),.clk(gclk));
	jor g04449(.dina(w_n4690_0[1]),.dinb(w_n4689_0[1]),.dout(n4691),.clk(gclk));
	jand g04450(.dina(w_n4691_0[2]),.dinb(w_n4686_0[2]),.dout(n4692),.clk(gclk));
	jor g04451(.dina(n4692),.dinb(w_n595_27[2]),.dout(n4693),.clk(gclk));
	jnot g04452(.din(w_n4374_0[0]),.dout(n4694),.clk(gclk));
	jor g04453(.dina(n4694),.dinb(w_n4372_0[0]),.dout(n4695),.clk(gclk));
	jor g04454(.dina(n4695),.dinb(w_n4499_26[2]),.dout(n4696),.clk(gclk));
	jxor g04455(.dina(n4696),.dinb(w_n4383_0[0]),.dout(n4697),.clk(gclk));
	jand g04456(.dina(w_n4686_0[1]),.dinb(w_n595_27[1]),.dout(n4698),.clk(gclk));
	jand g04457(.dina(n4698),.dinb(w_n4691_0[1]),.dout(n4699),.clk(gclk));
	jor g04458(.dina(w_n4699_0[1]),.dinb(w_n4697_0[1]),.dout(n4700),.clk(gclk));
	jand g04459(.dina(w_n4700_0[1]),.dinb(w_n4693_0[1]),.dout(n4701),.clk(gclk));
	jor g04460(.dina(w_n4701_0[2]),.dinb(w_n590_26[1]),.dout(n4702),.clk(gclk));
	jand g04461(.dina(w_n4701_0[1]),.dinb(w_n590_26[0]),.dout(n4703),.clk(gclk));
	jnot g04462(.din(w_n4386_0[0]),.dout(n4704),.clk(gclk));
	jand g04463(.dina(w_asqrt35_20[1]),.dinb(n4704),.dout(n4705),.clk(gclk));
	jand g04464(.dina(w_n4705_0[1]),.dinb(w_n4391_0[0]),.dout(n4706),.clk(gclk));
	jor g04465(.dina(n4706),.dinb(w_n4390_0[0]),.dout(n4707),.clk(gclk));
	jand g04466(.dina(w_n4705_0[0]),.dinb(w_n4392_0[0]),.dout(n4708),.clk(gclk));
	jnot g04467(.din(n4708),.dout(n4709),.clk(gclk));
	jand g04468(.dina(n4709),.dinb(n4707),.dout(n4710),.clk(gclk));
	jnot g04469(.din(n4710),.dout(n4711),.clk(gclk));
	jor g04470(.dina(w_n4711_0[1]),.dinb(n4703),.dout(n4712),.clk(gclk));
	jand g04471(.dina(w_n4712_0[1]),.dinb(w_n4702_0[1]),.dout(n4713),.clk(gclk));
	jor g04472(.dina(n4713),.dinb(w_n430_27[2]),.dout(n4714),.clk(gclk));
	jand g04473(.dina(w_n4702_0[0]),.dinb(w_n430_27[1]),.dout(n4715),.clk(gclk));
	jand g04474(.dina(n4715),.dinb(w_n4712_0[0]),.dout(n4716),.clk(gclk));
	jnot g04475(.din(w_n4394_0[0]),.dout(n4717),.clk(gclk));
	jand g04476(.dina(w_asqrt35_20[0]),.dinb(n4717),.dout(n4718),.clk(gclk));
	jand g04477(.dina(w_n4718_0[1]),.dinb(w_n4401_0[0]),.dout(n4719),.clk(gclk));
	jor g04478(.dina(n4719),.dinb(w_n4399_0[0]),.dout(n4720),.clk(gclk));
	jand g04479(.dina(w_n4718_0[0]),.dinb(w_n4402_0[0]),.dout(n4721),.clk(gclk));
	jnot g04480(.din(n4721),.dout(n4722),.clk(gclk));
	jand g04481(.dina(n4722),.dinb(n4720),.dout(n4723),.clk(gclk));
	jnot g04482(.din(n4723),.dout(n4724),.clk(gclk));
	jor g04483(.dina(w_n4724_0[1]),.dinb(w_n4716_0[1]),.dout(n4725),.clk(gclk));
	jand g04484(.dina(n4725),.dinb(w_n4714_0[1]),.dout(n4726),.clk(gclk));
	jor g04485(.dina(w_n4726_0[1]),.dinb(w_n425_26[1]),.dout(n4727),.clk(gclk));
	jxor g04486(.dina(w_n4403_0[0]),.dinb(w_n430_27[0]),.dout(n4728),.clk(gclk));
	jor g04487(.dina(n4728),.dinb(w_n4499_26[1]),.dout(n4729),.clk(gclk));
	jxor g04488(.dina(n4729),.dinb(w_n4414_0[0]),.dout(n4730),.clk(gclk));
	jand g04489(.dina(w_n4726_0[0]),.dinb(w_n425_26[0]),.dout(n4731),.clk(gclk));
	jor g04490(.dina(w_n4731_0[1]),.dinb(w_n4730_0[1]),.dout(n4732),.clk(gclk));
	jand g04491(.dina(w_n4732_0[2]),.dinb(w_n4727_0[2]),.dout(n4733),.clk(gclk));
	jor g04492(.dina(n4733),.dinb(w_n305_28[0]),.dout(n4734),.clk(gclk));
	jnot g04493(.din(w_n4419_0[0]),.dout(n4735),.clk(gclk));
	jor g04494(.dina(n4735),.dinb(w_n4417_0[0]),.dout(n4736),.clk(gclk));
	jor g04495(.dina(n4736),.dinb(w_n4499_26[0]),.dout(n4737),.clk(gclk));
	jxor g04496(.dina(n4737),.dinb(w_n4428_0[0]),.dout(n4738),.clk(gclk));
	jand g04497(.dina(w_n4727_0[1]),.dinb(w_n305_27[2]),.dout(n4739),.clk(gclk));
	jand g04498(.dina(n4739),.dinb(w_n4732_0[1]),.dout(n4740),.clk(gclk));
	jor g04499(.dina(w_n4740_0[1]),.dinb(w_n4738_0[1]),.dout(n4741),.clk(gclk));
	jand g04500(.dina(w_n4741_0[1]),.dinb(w_n4734_0[1]),.dout(n4742),.clk(gclk));
	jor g04501(.dina(w_n4742_0[2]),.dinb(w_n290_27[2]),.dout(n4743),.clk(gclk));
	jand g04502(.dina(w_n4742_0[1]),.dinb(w_n290_27[1]),.dout(n4744),.clk(gclk));
	jnot g04503(.din(w_n4431_0[0]),.dout(n4745),.clk(gclk));
	jand g04504(.dina(w_asqrt35_19[2]),.dinb(n4745),.dout(n4746),.clk(gclk));
	jand g04505(.dina(w_n4746_0[1]),.dinb(w_n4436_0[0]),.dout(n4747),.clk(gclk));
	jor g04506(.dina(n4747),.dinb(w_n4435_0[0]),.dout(n4748),.clk(gclk));
	jand g04507(.dina(w_n4746_0[0]),.dinb(w_n4437_0[0]),.dout(n4749),.clk(gclk));
	jnot g04508(.din(n4749),.dout(n4750),.clk(gclk));
	jand g04509(.dina(n4750),.dinb(n4748),.dout(n4751),.clk(gclk));
	jnot g04510(.din(n4751),.dout(n4752),.clk(gclk));
	jor g04511(.dina(w_n4752_0[1]),.dinb(n4744),.dout(n4753),.clk(gclk));
	jand g04512(.dina(w_n4753_0[1]),.dinb(w_n4743_0[1]),.dout(n4754),.clk(gclk));
	jor g04513(.dina(n4754),.dinb(w_n223_28[0]),.dout(n4755),.clk(gclk));
	jand g04514(.dina(w_n4743_0[0]),.dinb(w_n223_27[2]),.dout(n4756),.clk(gclk));
	jand g04515(.dina(n4756),.dinb(w_n4753_0[0]),.dout(n4757),.clk(gclk));
	jnot g04516(.din(w_n4439_0[0]),.dout(n4758),.clk(gclk));
	jand g04517(.dina(w_asqrt35_19[1]),.dinb(n4758),.dout(n4759),.clk(gclk));
	jand g04518(.dina(w_n4759_0[1]),.dinb(w_n4446_0[0]),.dout(n4760),.clk(gclk));
	jor g04519(.dina(n4760),.dinb(w_n4444_0[0]),.dout(n4761),.clk(gclk));
	jand g04520(.dina(w_n4759_0[0]),.dinb(w_n4447_0[0]),.dout(n4762),.clk(gclk));
	jnot g04521(.din(n4762),.dout(n4763),.clk(gclk));
	jand g04522(.dina(n4763),.dinb(n4761),.dout(n4764),.clk(gclk));
	jnot g04523(.din(n4764),.dout(n4765),.clk(gclk));
	jor g04524(.dina(w_n4765_0[1]),.dinb(w_n4757_0[1]),.dout(n4766),.clk(gclk));
	jand g04525(.dina(n4766),.dinb(w_n4755_0[1]),.dout(n4767),.clk(gclk));
	jor g04526(.dina(w_n4767_0[2]),.dinb(w_n199_32[1]),.dout(n4768),.clk(gclk));
	jand g04527(.dina(w_n4767_0[1]),.dinb(w_n199_32[0]),.dout(n4769),.clk(gclk));
	jxor g04528(.dina(w_n4448_0[0]),.dinb(w_n223_27[1]),.dout(n4770),.clk(gclk));
	jor g04529(.dina(n4770),.dinb(w_n4499_25[2]),.dout(n4771),.clk(gclk));
	jxor g04530(.dina(n4771),.dinb(w_n4459_0[0]),.dout(n4772),.clk(gclk));
	jor g04531(.dina(w_n4772_0[1]),.dinb(n4769),.dout(n4773),.clk(gclk));
	jand g04532(.dina(n4773),.dinb(n4768),.dout(n4774),.clk(gclk));
	jnot g04533(.din(w_n4464_0[0]),.dout(n4775),.clk(gclk));
	jor g04534(.dina(n4775),.dinb(w_n4462_0[0]),.dout(n4776),.clk(gclk));
	jor g04535(.dina(n4776),.dinb(w_n4499_25[1]),.dout(n4777),.clk(gclk));
	jxor g04536(.dina(n4777),.dinb(w_n4473_0[0]),.dout(n4778),.clk(gclk));
	jand g04537(.dina(w_asqrt35_19[0]),.dinb(w_n4487_0[1]),.dout(n4779),.clk(gclk));
	jand g04538(.dina(w_n4779_0[1]),.dinb(w_n4475_1[0]),.dout(n4780),.clk(gclk));
	jor g04539(.dina(n4780),.dinb(w_n4519_0[0]),.dout(n4781),.clk(gclk));
	jor g04540(.dina(n4781),.dinb(w_n4778_0[2]),.dout(n4782),.clk(gclk));
	jor g04541(.dina(n4782),.dinb(w_n4774_0[2]),.dout(n4783),.clk(gclk));
	jand g04542(.dina(n4783),.dinb(w_n194_31[1]),.dout(n4784),.clk(gclk));
	jand g04543(.dina(w_n4778_0[1]),.dinb(w_n4774_0[1]),.dout(n4785),.clk(gclk));
	jor g04544(.dina(w_n4779_0[0]),.dinb(w_n4475_0[2]),.dout(n4786),.clk(gclk));
	jand g04545(.dina(w_n4487_0[0]),.dinb(w_n4475_0[1]),.dout(n4787),.clk(gclk));
	jor g04546(.dina(n4787),.dinb(w_n194_31[0]),.dout(n4788),.clk(gclk));
	jnot g04547(.din(n4788),.dout(n4789),.clk(gclk));
	jand g04548(.dina(n4789),.dinb(n4786),.dout(n4790),.clk(gclk));
	jor g04549(.dina(w_n4790_0[1]),.dinb(w_n4785_0[2]),.dout(n4793),.clk(gclk));
	jor g04550(.dina(n4793),.dinb(w_n4784_0[1]),.dout(asqrt_fa_35),.clk(gclk));
	jand g04551(.dina(w_asqrt34_31),.dinb(w_a68_0[0]),.dout(n4795),.clk(gclk));
	jnot g04552(.din(w_a66_0[1]),.dout(n4796),.clk(gclk));
	jnot g04553(.din(w_a67_0[1]),.dout(n4797),.clk(gclk));
	jand g04554(.dina(w_n4502_1[0]),.dinb(w_n4797_0[1]),.dout(n4798),.clk(gclk));
	jand g04555(.dina(n4798),.dinb(w_n4796_1[1]),.dout(n4799),.clk(gclk));
	jor g04556(.dina(n4799),.dinb(n4795),.dout(n4800),.clk(gclk));
	jand g04557(.dina(w_n4800_0[2]),.dinb(w_asqrt35_18[2]),.dout(n4801),.clk(gclk));
	jand g04558(.dina(w_asqrt34_30[2]),.dinb(w_n4502_0[2]),.dout(n4802),.clk(gclk));
	jxor g04559(.dina(w_n4802_0[1]),.dinb(w_n4503_0[1]),.dout(n4803),.clk(gclk));
	jor g04560(.dina(w_n4800_0[1]),.dinb(w_asqrt35_18[1]),.dout(n4804),.clk(gclk));
	jand g04561(.dina(n4804),.dinb(w_n4803_0[1]),.dout(n4805),.clk(gclk));
	jor g04562(.dina(w_n4805_0[1]),.dinb(w_n4801_0[1]),.dout(n4806),.clk(gclk));
	jand g04563(.dina(n4806),.dinb(w_asqrt36_21[1]),.dout(n4807),.clk(gclk));
	jor g04564(.dina(w_n4801_0[0]),.dinb(w_asqrt36_21[0]),.dout(n4808),.clk(gclk));
	jor g04565(.dina(n4808),.dinb(w_n4805_0[0]),.dout(n4809),.clk(gclk));
	jand g04566(.dina(w_n4802_0[0]),.dinb(w_n4503_0[0]),.dout(n4810),.clk(gclk));
	jnot g04567(.din(w_n4784_0[0]),.dout(n4811),.clk(gclk));
	jnot g04568(.din(w_n4785_0[1]),.dout(n4812),.clk(gclk));
	jnot g04569(.din(w_n4790_0[0]),.dout(n4813),.clk(gclk));
	jand g04570(.dina(n4813),.dinb(w_asqrt35_18[0]),.dout(n4814),.clk(gclk));
	jand g04571(.dina(n4814),.dinb(n4812),.dout(n4815),.clk(gclk));
	jand g04572(.dina(n4815),.dinb(n4811),.dout(n4816),.clk(gclk));
	jor g04573(.dina(n4816),.dinb(n4810),.dout(n4817),.clk(gclk));
	jxor g04574(.dina(n4817),.dinb(w_n4193_0[1]),.dout(n4818),.clk(gclk));
	jand g04575(.dina(w_n4818_0[1]),.dinb(w_n4809_0[1]),.dout(n4819),.clk(gclk));
	jor g04576(.dina(n4819),.dinb(w_n4807_0[1]),.dout(n4820),.clk(gclk));
	jand g04577(.dina(w_n4820_0[2]),.dinb(w_asqrt37_18[2]),.dout(n4821),.clk(gclk));
	jor g04578(.dina(w_n4820_0[1]),.dinb(w_asqrt37_18[1]),.dout(n4822),.clk(gclk));
	jxor g04579(.dina(w_n4507_0[0]),.dinb(w_n4494_22[1]),.dout(n4823),.clk(gclk));
	jand g04580(.dina(n4823),.dinb(w_asqrt34_30[1]),.dout(n4824),.clk(gclk));
	jxor g04581(.dina(n4824),.dinb(w_n4510_0[0]),.dout(n4825),.clk(gclk));
	jnot g04582(.din(w_n4825_0[1]),.dout(n4826),.clk(gclk));
	jand g04583(.dina(n4826),.dinb(n4822),.dout(n4827),.clk(gclk));
	jor g04584(.dina(w_n4827_0[1]),.dinb(w_n4821_0[1]),.dout(n4828),.clk(gclk));
	jand g04585(.dina(n4828),.dinb(w_asqrt38_21[1]),.dout(n4829),.clk(gclk));
	jnot g04586(.din(w_n4516_0[0]),.dout(n4830),.clk(gclk));
	jand g04587(.dina(n4830),.dinb(w_n4514_0[0]),.dout(n4831),.clk(gclk));
	jand g04588(.dina(n4831),.dinb(w_asqrt34_30[0]),.dout(n4832),.clk(gclk));
	jxor g04589(.dina(n4832),.dinb(w_n4524_0[0]),.dout(n4833),.clk(gclk));
	jnot g04590(.din(n4833),.dout(n4834),.clk(gclk));
	jor g04591(.dina(w_n4821_0[0]),.dinb(w_asqrt38_21[0]),.dout(n4835),.clk(gclk));
	jor g04592(.dina(n4835),.dinb(w_n4827_0[0]),.dout(n4836),.clk(gclk));
	jand g04593(.dina(w_n4836_0[1]),.dinb(w_n4834_0[1]),.dout(n4837),.clk(gclk));
	jor g04594(.dina(w_n4837_0[1]),.dinb(w_n4829_0[1]),.dout(n4838),.clk(gclk));
	jand g04595(.dina(w_n4838_0[2]),.dinb(w_asqrt39_18[2]),.dout(n4839),.clk(gclk));
	jor g04596(.dina(w_n4838_0[1]),.dinb(w_asqrt39_18[1]),.dout(n4840),.clk(gclk));
	jnot g04597(.din(w_n4531_0[0]),.dout(n4841),.clk(gclk));
	jxor g04598(.dina(w_n4526_0[0]),.dinb(w_n3907_22[1]),.dout(n4842),.clk(gclk));
	jand g04599(.dina(n4842),.dinb(w_asqrt34_29[2]),.dout(n4843),.clk(gclk));
	jxor g04600(.dina(n4843),.dinb(n4841),.dout(n4844),.clk(gclk));
	jand g04601(.dina(w_n4844_0[1]),.dinb(n4840),.dout(n4845),.clk(gclk));
	jor g04602(.dina(w_n4845_0[1]),.dinb(w_n4839_0[1]),.dout(n4846),.clk(gclk));
	jand g04603(.dina(n4846),.dinb(w_asqrt40_21[1]),.dout(n4847),.clk(gclk));
	jor g04604(.dina(w_n4839_0[0]),.dinb(w_asqrt40_21[0]),.dout(n4848),.clk(gclk));
	jor g04605(.dina(n4848),.dinb(w_n4845_0[0]),.dout(n4849),.clk(gclk));
	jnot g04606(.din(w_n4538_0[0]),.dout(n4850),.clk(gclk));
	jnot g04607(.din(w_n4540_0[0]),.dout(n4851),.clk(gclk));
	jand g04608(.dina(w_asqrt34_29[1]),.dinb(w_n4534_0[0]),.dout(n4852),.clk(gclk));
	jand g04609(.dina(w_n4852_0[1]),.dinb(n4851),.dout(n4853),.clk(gclk));
	jor g04610(.dina(n4853),.dinb(n4850),.dout(n4854),.clk(gclk));
	jnot g04611(.din(w_n4541_0[0]),.dout(n4855),.clk(gclk));
	jand g04612(.dina(w_n4852_0[0]),.dinb(n4855),.dout(n4856),.clk(gclk));
	jnot g04613(.din(n4856),.dout(n4857),.clk(gclk));
	jand g04614(.dina(n4857),.dinb(n4854),.dout(n4858),.clk(gclk));
	jand g04615(.dina(w_n4858_0[1]),.dinb(w_n4849_0[1]),.dout(n4859),.clk(gclk));
	jor g04616(.dina(n4859),.dinb(w_n4847_0[1]),.dout(n4860),.clk(gclk));
	jand g04617(.dina(w_n4860_0[2]),.dinb(w_asqrt41_19[0]),.dout(n4861),.clk(gclk));
	jor g04618(.dina(w_n4860_0[1]),.dinb(w_asqrt41_18[2]),.dout(n4862),.clk(gclk));
	jxor g04619(.dina(w_n4542_0[0]),.dinb(w_n3371_22[2]),.dout(n4863),.clk(gclk));
	jand g04620(.dina(n4863),.dinb(w_asqrt34_29[0]),.dout(n4864),.clk(gclk));
	jxor g04621(.dina(n4864),.dinb(w_n4547_0[0]),.dout(n4865),.clk(gclk));
	jand g04622(.dina(w_n4865_0[1]),.dinb(n4862),.dout(n4866),.clk(gclk));
	jor g04623(.dina(w_n4866_0[1]),.dinb(w_n4861_0[1]),.dout(n4867),.clk(gclk));
	jand g04624(.dina(n4867),.dinb(w_asqrt42_21[1]),.dout(n4868),.clk(gclk));
	jnot g04625(.din(w_n4553_0[0]),.dout(n4869),.clk(gclk));
	jand g04626(.dina(n4869),.dinb(w_n4551_0[0]),.dout(n4870),.clk(gclk));
	jand g04627(.dina(n4870),.dinb(w_asqrt34_28[2]),.dout(n4871),.clk(gclk));
	jxor g04628(.dina(n4871),.dinb(w_n4561_0[0]),.dout(n4872),.clk(gclk));
	jnot g04629(.din(n4872),.dout(n4873),.clk(gclk));
	jor g04630(.dina(w_n4861_0[0]),.dinb(w_asqrt42_21[0]),.dout(n4874),.clk(gclk));
	jor g04631(.dina(n4874),.dinb(w_n4866_0[0]),.dout(n4875),.clk(gclk));
	jand g04632(.dina(w_n4875_0[1]),.dinb(w_n4873_0[1]),.dout(n4876),.clk(gclk));
	jor g04633(.dina(w_n4876_0[1]),.dinb(w_n4868_0[1]),.dout(n4877),.clk(gclk));
	jand g04634(.dina(w_n4877_0[2]),.dinb(w_asqrt43_19[0]),.dout(n4878),.clk(gclk));
	jor g04635(.dina(w_n4877_0[1]),.dinb(w_asqrt43_18[2]),.dout(n4879),.clk(gclk));
	jxor g04636(.dina(w_n4563_0[0]),.dinb(w_n2870_22[2]),.dout(n4880),.clk(gclk));
	jand g04637(.dina(n4880),.dinb(w_asqrt34_28[1]),.dout(n4881),.clk(gclk));
	jxor g04638(.dina(n4881),.dinb(w_n4569_0[0]),.dout(n4882),.clk(gclk));
	jand g04639(.dina(w_n4882_0[1]),.dinb(n4879),.dout(n4883),.clk(gclk));
	jor g04640(.dina(w_n4883_0[1]),.dinb(w_n4878_0[1]),.dout(n4884),.clk(gclk));
	jand g04641(.dina(n4884),.dinb(w_asqrt44_21[1]),.dout(n4885),.clk(gclk));
	jor g04642(.dina(w_n4878_0[0]),.dinb(w_asqrt44_21[0]),.dout(n4886),.clk(gclk));
	jor g04643(.dina(n4886),.dinb(w_n4883_0[0]),.dout(n4887),.clk(gclk));
	jnot g04644(.din(w_n4577_0[0]),.dout(n4888),.clk(gclk));
	jnot g04645(.din(w_n4579_0[0]),.dout(n4889),.clk(gclk));
	jand g04646(.dina(w_asqrt34_28[0]),.dinb(w_n4573_0[0]),.dout(n4890),.clk(gclk));
	jand g04647(.dina(w_n4890_0[1]),.dinb(n4889),.dout(n4891),.clk(gclk));
	jor g04648(.dina(n4891),.dinb(n4888),.dout(n4892),.clk(gclk));
	jnot g04649(.din(w_n4580_0[0]),.dout(n4893),.clk(gclk));
	jand g04650(.dina(w_n4890_0[0]),.dinb(n4893),.dout(n4894),.clk(gclk));
	jnot g04651(.din(n4894),.dout(n4895),.clk(gclk));
	jand g04652(.dina(n4895),.dinb(n4892),.dout(n4896),.clk(gclk));
	jand g04653(.dina(w_n4896_0[1]),.dinb(w_n4887_0[1]),.dout(n4897),.clk(gclk));
	jor g04654(.dina(n4897),.dinb(w_n4885_0[1]),.dout(n4898),.clk(gclk));
	jand g04655(.dina(w_n4898_0[1]),.dinb(w_asqrt45_19[1]),.dout(n4899),.clk(gclk));
	jxor g04656(.dina(w_n4581_0[0]),.dinb(w_n2420_23[1]),.dout(n4900),.clk(gclk));
	jand g04657(.dina(n4900),.dinb(w_asqrt34_27[2]),.dout(n4901),.clk(gclk));
	jxor g04658(.dina(n4901),.dinb(w_n4588_0[0]),.dout(n4902),.clk(gclk));
	jnot g04659(.din(n4902),.dout(n4903),.clk(gclk));
	jor g04660(.dina(w_n4898_0[0]),.dinb(w_asqrt45_19[0]),.dout(n4904),.clk(gclk));
	jand g04661(.dina(w_n4904_0[1]),.dinb(w_n4903_0[1]),.dout(n4905),.clk(gclk));
	jor g04662(.dina(w_n4905_0[2]),.dinb(w_n4899_0[2]),.dout(n4906),.clk(gclk));
	jand g04663(.dina(n4906),.dinb(w_asqrt46_21[1]),.dout(n4907),.clk(gclk));
	jnot g04664(.din(w_n4593_0[0]),.dout(n4908),.clk(gclk));
	jand g04665(.dina(n4908),.dinb(w_n4591_0[0]),.dout(n4909),.clk(gclk));
	jand g04666(.dina(n4909),.dinb(w_asqrt34_27[1]),.dout(n4910),.clk(gclk));
	jxor g04667(.dina(n4910),.dinb(w_n4601_0[0]),.dout(n4911),.clk(gclk));
	jnot g04668(.din(n4911),.dout(n4912),.clk(gclk));
	jor g04669(.dina(w_n4899_0[1]),.dinb(w_asqrt46_21[0]),.dout(n4913),.clk(gclk));
	jor g04670(.dina(n4913),.dinb(w_n4905_0[1]),.dout(n4914),.clk(gclk));
	jand g04671(.dina(w_n4914_0[1]),.dinb(w_n4912_0[1]),.dout(n4915),.clk(gclk));
	jor g04672(.dina(w_n4915_0[1]),.dinb(w_n4907_0[1]),.dout(n4916),.clk(gclk));
	jand g04673(.dina(w_n4916_0[2]),.dinb(w_asqrt47_19[1]),.dout(n4917),.clk(gclk));
	jor g04674(.dina(w_n4916_0[1]),.dinb(w_asqrt47_19[0]),.dout(n4918),.clk(gclk));
	jnot g04675(.din(w_n4607_0[0]),.dout(n4919),.clk(gclk));
	jnot g04676(.din(w_n4608_0[0]),.dout(n4920),.clk(gclk));
	jand g04677(.dina(w_asqrt34_27[0]),.dinb(w_n4604_0[0]),.dout(n4921),.clk(gclk));
	jand g04678(.dina(w_n4921_0[1]),.dinb(n4920),.dout(n4922),.clk(gclk));
	jor g04679(.dina(n4922),.dinb(n4919),.dout(n4923),.clk(gclk));
	jnot g04680(.din(w_n4609_0[0]),.dout(n4924),.clk(gclk));
	jand g04681(.dina(w_n4921_0[0]),.dinb(n4924),.dout(n4925),.clk(gclk));
	jnot g04682(.din(n4925),.dout(n4926),.clk(gclk));
	jand g04683(.dina(n4926),.dinb(n4923),.dout(n4927),.clk(gclk));
	jand g04684(.dina(w_n4927_0[1]),.dinb(n4918),.dout(n4928),.clk(gclk));
	jor g04685(.dina(w_n4928_0[1]),.dinb(w_n4917_0[1]),.dout(n4929),.clk(gclk));
	jand g04686(.dina(n4929),.dinb(w_asqrt48_21[1]),.dout(n4930),.clk(gclk));
	jor g04687(.dina(w_n4917_0[0]),.dinb(w_asqrt48_21[0]),.dout(n4931),.clk(gclk));
	jor g04688(.dina(n4931),.dinb(w_n4928_0[0]),.dout(n4932),.clk(gclk));
	jnot g04689(.din(w_n4615_0[0]),.dout(n4933),.clk(gclk));
	jnot g04690(.din(w_n4617_0[0]),.dout(n4934),.clk(gclk));
	jand g04691(.dina(w_asqrt34_26[2]),.dinb(w_n4611_0[0]),.dout(n4935),.clk(gclk));
	jand g04692(.dina(w_n4935_0[1]),.dinb(n4934),.dout(n4936),.clk(gclk));
	jor g04693(.dina(n4936),.dinb(n4933),.dout(n4937),.clk(gclk));
	jnot g04694(.din(w_n4618_0[0]),.dout(n4938),.clk(gclk));
	jand g04695(.dina(w_n4935_0[0]),.dinb(n4938),.dout(n4939),.clk(gclk));
	jnot g04696(.din(n4939),.dout(n4940),.clk(gclk));
	jand g04697(.dina(n4940),.dinb(n4937),.dout(n4941),.clk(gclk));
	jand g04698(.dina(w_n4941_0[1]),.dinb(w_n4932_0[1]),.dout(n4942),.clk(gclk));
	jor g04699(.dina(n4942),.dinb(w_n4930_0[1]),.dout(n4943),.clk(gclk));
	jand g04700(.dina(w_n4943_0[1]),.dinb(w_asqrt49_19[2]),.dout(n4944),.clk(gclk));
	jxor g04701(.dina(w_n4619_0[0]),.dinb(w_n1641_24[0]),.dout(n4945),.clk(gclk));
	jand g04702(.dina(n4945),.dinb(w_asqrt34_26[1]),.dout(n4946),.clk(gclk));
	jxor g04703(.dina(n4946),.dinb(w_n4629_0[0]),.dout(n4947),.clk(gclk));
	jnot g04704(.din(n4947),.dout(n4948),.clk(gclk));
	jor g04705(.dina(w_n4943_0[0]),.dinb(w_asqrt49_19[1]),.dout(n4949),.clk(gclk));
	jand g04706(.dina(w_n4949_0[1]),.dinb(w_n4948_0[1]),.dout(n4950),.clk(gclk));
	jor g04707(.dina(w_n4950_0[2]),.dinb(w_n4944_0[2]),.dout(n4951),.clk(gclk));
	jand g04708(.dina(n4951),.dinb(w_asqrt50_21[1]),.dout(n4952),.clk(gclk));
	jnot g04709(.din(w_n4634_0[0]),.dout(n4953),.clk(gclk));
	jand g04710(.dina(n4953),.dinb(w_n4632_0[0]),.dout(n4954),.clk(gclk));
	jand g04711(.dina(n4954),.dinb(w_asqrt34_26[0]),.dout(n4955),.clk(gclk));
	jxor g04712(.dina(n4955),.dinb(w_n4642_0[0]),.dout(n4956),.clk(gclk));
	jnot g04713(.din(n4956),.dout(n4957),.clk(gclk));
	jor g04714(.dina(w_n4944_0[1]),.dinb(w_asqrt50_21[0]),.dout(n4958),.clk(gclk));
	jor g04715(.dina(n4958),.dinb(w_n4950_0[1]),.dout(n4959),.clk(gclk));
	jand g04716(.dina(w_n4959_0[1]),.dinb(w_n4957_0[1]),.dout(n4960),.clk(gclk));
	jor g04717(.dina(w_n4960_0[1]),.dinb(w_n4952_0[1]),.dout(n4961),.clk(gclk));
	jand g04718(.dina(w_n4961_0[2]),.dinb(w_asqrt51_19[2]),.dout(n4962),.clk(gclk));
	jor g04719(.dina(w_n4961_0[1]),.dinb(w_asqrt51_19[1]),.dout(n4963),.clk(gclk));
	jnot g04720(.din(w_n4648_0[0]),.dout(n4964),.clk(gclk));
	jnot g04721(.din(w_n4649_0[0]),.dout(n4965),.clk(gclk));
	jand g04722(.dina(w_asqrt34_25[2]),.dinb(w_n4645_0[0]),.dout(n4966),.clk(gclk));
	jand g04723(.dina(w_n4966_0[1]),.dinb(n4965),.dout(n4967),.clk(gclk));
	jor g04724(.dina(n4967),.dinb(n4964),.dout(n4968),.clk(gclk));
	jnot g04725(.din(w_n4650_0[0]),.dout(n4969),.clk(gclk));
	jand g04726(.dina(w_n4966_0[0]),.dinb(n4969),.dout(n4970),.clk(gclk));
	jnot g04727(.din(n4970),.dout(n4971),.clk(gclk));
	jand g04728(.dina(n4971),.dinb(n4968),.dout(n4972),.clk(gclk));
	jand g04729(.dina(w_n4972_0[1]),.dinb(n4963),.dout(n4973),.clk(gclk));
	jor g04730(.dina(w_n4973_0[1]),.dinb(w_n4962_0[1]),.dout(n4974),.clk(gclk));
	jand g04731(.dina(n4974),.dinb(w_asqrt52_21[1]),.dout(n4975),.clk(gclk));
	jor g04732(.dina(w_n4962_0[0]),.dinb(w_asqrt52_21[0]),.dout(n4976),.clk(gclk));
	jor g04733(.dina(n4976),.dinb(w_n4973_0[0]),.dout(n4977),.clk(gclk));
	jnot g04734(.din(w_n4656_0[0]),.dout(n4978),.clk(gclk));
	jnot g04735(.din(w_n4658_0[0]),.dout(n4979),.clk(gclk));
	jand g04736(.dina(w_asqrt34_25[1]),.dinb(w_n4652_0[0]),.dout(n4980),.clk(gclk));
	jand g04737(.dina(w_n4980_0[1]),.dinb(n4979),.dout(n4981),.clk(gclk));
	jor g04738(.dina(n4981),.dinb(n4978),.dout(n4982),.clk(gclk));
	jnot g04739(.din(w_n4659_0[0]),.dout(n4983),.clk(gclk));
	jand g04740(.dina(w_n4980_0[0]),.dinb(n4983),.dout(n4984),.clk(gclk));
	jnot g04741(.din(n4984),.dout(n4985),.clk(gclk));
	jand g04742(.dina(n4985),.dinb(n4982),.dout(n4986),.clk(gclk));
	jand g04743(.dina(w_n4986_0[1]),.dinb(w_n4977_0[1]),.dout(n4987),.clk(gclk));
	jor g04744(.dina(n4987),.dinb(w_n4975_0[1]),.dout(n4988),.clk(gclk));
	jand g04745(.dina(w_n4988_0[1]),.dinb(w_asqrt53_20[0]),.dout(n4989),.clk(gclk));
	jxor g04746(.dina(w_n4660_0[0]),.dinb(w_n1034_25[0]),.dout(n4990),.clk(gclk));
	jand g04747(.dina(n4990),.dinb(w_asqrt34_25[0]),.dout(n4991),.clk(gclk));
	jxor g04748(.dina(n4991),.dinb(w_n4670_0[0]),.dout(n4992),.clk(gclk));
	jnot g04749(.din(n4992),.dout(n4993),.clk(gclk));
	jor g04750(.dina(w_n4988_0[0]),.dinb(w_asqrt53_19[2]),.dout(n4994),.clk(gclk));
	jand g04751(.dina(w_n4994_0[1]),.dinb(w_n4993_0[1]),.dout(n4995),.clk(gclk));
	jor g04752(.dina(w_n4995_0[2]),.dinb(w_n4989_0[2]),.dout(n4996),.clk(gclk));
	jand g04753(.dina(n4996),.dinb(w_asqrt54_21[1]),.dout(n4997),.clk(gclk));
	jnot g04754(.din(w_n4675_0[0]),.dout(n4998),.clk(gclk));
	jand g04755(.dina(n4998),.dinb(w_n4673_0[0]),.dout(n4999),.clk(gclk));
	jand g04756(.dina(n4999),.dinb(w_asqrt34_24[2]),.dout(n5000),.clk(gclk));
	jxor g04757(.dina(n5000),.dinb(w_n4683_0[0]),.dout(n5001),.clk(gclk));
	jnot g04758(.din(n5001),.dout(n5002),.clk(gclk));
	jor g04759(.dina(w_n4989_0[1]),.dinb(w_asqrt54_21[0]),.dout(n5003),.clk(gclk));
	jor g04760(.dina(n5003),.dinb(w_n4995_0[1]),.dout(n5004),.clk(gclk));
	jand g04761(.dina(w_n5004_0[1]),.dinb(w_n5002_0[1]),.dout(n5005),.clk(gclk));
	jor g04762(.dina(w_n5005_0[1]),.dinb(w_n4997_0[1]),.dout(n5006),.clk(gclk));
	jand g04763(.dina(w_n5006_0[2]),.dinb(w_asqrt55_20[1]),.dout(n5007),.clk(gclk));
	jor g04764(.dina(w_n5006_0[1]),.dinb(w_asqrt55_20[0]),.dout(n5008),.clk(gclk));
	jnot g04765(.din(w_n4689_0[0]),.dout(n5009),.clk(gclk));
	jnot g04766(.din(w_n4690_0[0]),.dout(n5010),.clk(gclk));
	jand g04767(.dina(w_asqrt34_24[1]),.dinb(w_n4686_0[0]),.dout(n5011),.clk(gclk));
	jand g04768(.dina(w_n5011_0[1]),.dinb(n5010),.dout(n5012),.clk(gclk));
	jor g04769(.dina(n5012),.dinb(n5009),.dout(n5013),.clk(gclk));
	jnot g04770(.din(w_n4691_0[0]),.dout(n5014),.clk(gclk));
	jand g04771(.dina(w_n5011_0[0]),.dinb(n5014),.dout(n5015),.clk(gclk));
	jnot g04772(.din(n5015),.dout(n5016),.clk(gclk));
	jand g04773(.dina(n5016),.dinb(n5013),.dout(n5017),.clk(gclk));
	jand g04774(.dina(w_n5017_0[1]),.dinb(n5008),.dout(n5018),.clk(gclk));
	jor g04775(.dina(w_n5018_0[1]),.dinb(w_n5007_0[1]),.dout(n5019),.clk(gclk));
	jand g04776(.dina(n5019),.dinb(w_asqrt56_21[1]),.dout(n5020),.clk(gclk));
	jor g04777(.dina(w_n5007_0[0]),.dinb(w_asqrt56_21[0]),.dout(n5021),.clk(gclk));
	jor g04778(.dina(n5021),.dinb(w_n5018_0[0]),.dout(n5022),.clk(gclk));
	jnot g04779(.din(w_n4697_0[0]),.dout(n5023),.clk(gclk));
	jnot g04780(.din(w_n4699_0[0]),.dout(n5024),.clk(gclk));
	jand g04781(.dina(w_asqrt34_24[0]),.dinb(w_n4693_0[0]),.dout(n5025),.clk(gclk));
	jand g04782(.dina(w_n5025_0[1]),.dinb(n5024),.dout(n5026),.clk(gclk));
	jor g04783(.dina(n5026),.dinb(n5023),.dout(n5027),.clk(gclk));
	jnot g04784(.din(w_n4700_0[0]),.dout(n5028),.clk(gclk));
	jand g04785(.dina(w_n5025_0[0]),.dinb(n5028),.dout(n5029),.clk(gclk));
	jnot g04786(.din(n5029),.dout(n5030),.clk(gclk));
	jand g04787(.dina(n5030),.dinb(n5027),.dout(n5031),.clk(gclk));
	jand g04788(.dina(w_n5031_0[1]),.dinb(w_n5022_0[1]),.dout(n5032),.clk(gclk));
	jor g04789(.dina(n5032),.dinb(w_n5020_0[1]),.dout(n5033),.clk(gclk));
	jand g04790(.dina(w_n5033_0[1]),.dinb(w_asqrt57_20[2]),.dout(n5034),.clk(gclk));
	jxor g04791(.dina(w_n4701_0[0]),.dinb(w_n590_25[2]),.dout(n5035),.clk(gclk));
	jand g04792(.dina(n5035),.dinb(w_asqrt34_23[2]),.dout(n5036),.clk(gclk));
	jxor g04793(.dina(n5036),.dinb(w_n4711_0[0]),.dout(n5037),.clk(gclk));
	jnot g04794(.din(n5037),.dout(n5038),.clk(gclk));
	jor g04795(.dina(w_n5033_0[0]),.dinb(w_asqrt57_20[1]),.dout(n5039),.clk(gclk));
	jand g04796(.dina(w_n5039_0[1]),.dinb(w_n5038_0[1]),.dout(n5040),.clk(gclk));
	jor g04797(.dina(w_n5040_0[2]),.dinb(w_n5034_0[2]),.dout(n5041),.clk(gclk));
	jand g04798(.dina(n5041),.dinb(w_asqrt58_21[1]),.dout(n5042),.clk(gclk));
	jnot g04799(.din(w_n4716_0[0]),.dout(n5043),.clk(gclk));
	jand g04800(.dina(n5043),.dinb(w_n4714_0[0]),.dout(n5044),.clk(gclk));
	jand g04801(.dina(n5044),.dinb(w_asqrt34_23[1]),.dout(n5045),.clk(gclk));
	jxor g04802(.dina(n5045),.dinb(w_n4724_0[0]),.dout(n5046),.clk(gclk));
	jnot g04803(.din(n5046),.dout(n5047),.clk(gclk));
	jor g04804(.dina(w_n5034_0[1]),.dinb(w_asqrt58_21[0]),.dout(n5048),.clk(gclk));
	jor g04805(.dina(n5048),.dinb(w_n5040_0[1]),.dout(n5049),.clk(gclk));
	jand g04806(.dina(w_n5049_0[1]),.dinb(w_n5047_0[1]),.dout(n5050),.clk(gclk));
	jor g04807(.dina(w_n5050_0[1]),.dinb(w_n5042_0[1]),.dout(n5051),.clk(gclk));
	jand g04808(.dina(w_n5051_0[2]),.dinb(w_asqrt59_21[0]),.dout(n5052),.clk(gclk));
	jor g04809(.dina(w_n5051_0[1]),.dinb(w_asqrt59_20[2]),.dout(n5053),.clk(gclk));
	jnot g04810(.din(w_n4730_0[0]),.dout(n5054),.clk(gclk));
	jnot g04811(.din(w_n4731_0[0]),.dout(n5055),.clk(gclk));
	jand g04812(.dina(w_asqrt34_23[0]),.dinb(w_n4727_0[0]),.dout(n5056),.clk(gclk));
	jand g04813(.dina(w_n5056_0[1]),.dinb(n5055),.dout(n5057),.clk(gclk));
	jor g04814(.dina(n5057),.dinb(n5054),.dout(n5058),.clk(gclk));
	jnot g04815(.din(w_n4732_0[0]),.dout(n5059),.clk(gclk));
	jand g04816(.dina(w_n5056_0[0]),.dinb(n5059),.dout(n5060),.clk(gclk));
	jnot g04817(.din(n5060),.dout(n5061),.clk(gclk));
	jand g04818(.dina(n5061),.dinb(n5058),.dout(n5062),.clk(gclk));
	jand g04819(.dina(w_n5062_0[1]),.dinb(n5053),.dout(n5063),.clk(gclk));
	jor g04820(.dina(w_n5063_0[1]),.dinb(w_n5052_0[1]),.dout(n5064),.clk(gclk));
	jand g04821(.dina(n5064),.dinb(w_asqrt60_21[0]),.dout(n5065),.clk(gclk));
	jor g04822(.dina(w_n5052_0[0]),.dinb(w_asqrt60_20[2]),.dout(n5066),.clk(gclk));
	jor g04823(.dina(n5066),.dinb(w_n5063_0[0]),.dout(n5067),.clk(gclk));
	jnot g04824(.din(w_n4738_0[0]),.dout(n5068),.clk(gclk));
	jnot g04825(.din(w_n4740_0[0]),.dout(n5069),.clk(gclk));
	jand g04826(.dina(w_asqrt34_22[2]),.dinb(w_n4734_0[0]),.dout(n5070),.clk(gclk));
	jand g04827(.dina(w_n5070_0[1]),.dinb(n5069),.dout(n5071),.clk(gclk));
	jor g04828(.dina(n5071),.dinb(n5068),.dout(n5072),.clk(gclk));
	jnot g04829(.din(w_n4741_0[0]),.dout(n5073),.clk(gclk));
	jand g04830(.dina(w_n5070_0[0]),.dinb(n5073),.dout(n5074),.clk(gclk));
	jnot g04831(.din(n5074),.dout(n5075),.clk(gclk));
	jand g04832(.dina(n5075),.dinb(n5072),.dout(n5076),.clk(gclk));
	jand g04833(.dina(w_n5076_0[1]),.dinb(w_n5067_0[1]),.dout(n5077),.clk(gclk));
	jor g04834(.dina(n5077),.dinb(w_n5065_0[1]),.dout(n5078),.clk(gclk));
	jand g04835(.dina(w_n5078_0[1]),.dinb(w_asqrt61_21[1]),.dout(n5079),.clk(gclk));
	jxor g04836(.dina(w_n4742_0[0]),.dinb(w_n290_27[0]),.dout(n5080),.clk(gclk));
	jand g04837(.dina(n5080),.dinb(w_asqrt34_22[1]),.dout(n5081),.clk(gclk));
	jxor g04838(.dina(n5081),.dinb(w_n4752_0[0]),.dout(n5082),.clk(gclk));
	jnot g04839(.din(n5082),.dout(n5083),.clk(gclk));
	jor g04840(.dina(w_n5078_0[0]),.dinb(w_asqrt61_21[0]),.dout(n5084),.clk(gclk));
	jand g04841(.dina(w_n5084_0[1]),.dinb(w_n5083_0[1]),.dout(n5085),.clk(gclk));
	jor g04842(.dina(w_n5085_0[2]),.dinb(w_n5079_0[2]),.dout(n5086),.clk(gclk));
	jand g04843(.dina(n5086),.dinb(w_asqrt62_21[1]),.dout(n5087),.clk(gclk));
	jnot g04844(.din(w_n4757_0[0]),.dout(n5088),.clk(gclk));
	jand g04845(.dina(n5088),.dinb(w_n4755_0[0]),.dout(n5089),.clk(gclk));
	jand g04846(.dina(n5089),.dinb(w_asqrt34_22[0]),.dout(n5090),.clk(gclk));
	jxor g04847(.dina(n5090),.dinb(w_n4765_0[0]),.dout(n5091),.clk(gclk));
	jnot g04848(.din(n5091),.dout(n5092),.clk(gclk));
	jor g04849(.dina(w_n5079_0[1]),.dinb(w_asqrt62_21[0]),.dout(n5093),.clk(gclk));
	jor g04850(.dina(n5093),.dinb(w_n5085_0[1]),.dout(n5094),.clk(gclk));
	jand g04851(.dina(w_n5094_0[1]),.dinb(w_n5092_0[1]),.dout(n5095),.clk(gclk));
	jor g04852(.dina(w_n5095_0[1]),.dinb(w_n5087_0[1]),.dout(n5096),.clk(gclk));
	jxor g04853(.dina(w_n4767_0[0]),.dinb(w_n199_31[2]),.dout(n5097),.clk(gclk));
	jand g04854(.dina(n5097),.dinb(w_asqrt34_21[2]),.dout(n5098),.clk(gclk));
	jxor g04855(.dina(n5098),.dinb(w_n4772_0[0]),.dout(n5099),.clk(gclk));
	jnot g04856(.din(w_n4774_0[0]),.dout(n5100),.clk(gclk));
	jnot g04857(.din(w_n4778_0[0]),.dout(n5101),.clk(gclk));
	jand g04858(.dina(w_asqrt34_21[1]),.dinb(w_n5101_0[1]),.dout(n5102),.clk(gclk));
	jand g04859(.dina(w_n5102_0[1]),.dinb(w_n5100_0[2]),.dout(n5103),.clk(gclk));
	jor g04860(.dina(n5103),.dinb(w_n4785_0[0]),.dout(n5104),.clk(gclk));
	jor g04861(.dina(n5104),.dinb(w_n5099_0[1]),.dout(n5105),.clk(gclk));
	jnot g04862(.din(n5105),.dout(n5106),.clk(gclk));
	jand g04863(.dina(n5106),.dinb(w_n5096_1[2]),.dout(n5107),.clk(gclk));
	jor g04864(.dina(n5107),.dinb(w_asqrt63_11[1]),.dout(n5108),.clk(gclk));
	jnot g04865(.din(w_n5099_0[0]),.dout(n5109),.clk(gclk));
	jor g04866(.dina(w_n5109_0[2]),.dinb(w_n5096_1[1]),.dout(n5110),.clk(gclk));
	jor g04867(.dina(w_n5102_0[0]),.dinb(w_n5100_0[1]),.dout(n5111),.clk(gclk));
	jand g04868(.dina(w_n5101_0[0]),.dinb(w_n5100_0[0]),.dout(n5112),.clk(gclk));
	jor g04869(.dina(n5112),.dinb(w_n194_30[2]),.dout(n5113),.clk(gclk));
	jnot g04870(.din(n5113),.dout(n5114),.clk(gclk));
	jand g04871(.dina(n5114),.dinb(n5111),.dout(n5115),.clk(gclk));
	jnot g04872(.din(w_asqrt34_21[0]),.dout(n5116),.clk(gclk));
	jnot g04873(.din(w_n5115_0[1]),.dout(n5119),.clk(gclk));
	jand g04874(.dina(n5119),.dinb(w_n5110_0[1]),.dout(n5120),.clk(gclk));
	jand g04875(.dina(n5120),.dinb(w_n5108_0[1]),.dout(n5121),.clk(gclk));
	jnot g04876(.din(w_n5121_29[2]),.dout(asqrt_fa_34),.clk(gclk));
	jor g04877(.dina(w_n5121_29[1]),.dinb(w_n4796_1[0]),.dout(n5123),.clk(gclk));
	jnot g04878(.din(w_a64_0[1]),.dout(n5124),.clk(gclk));
	jnot g04879(.din(a[65]),.dout(n5125),.clk(gclk));
	jand g04880(.dina(w_n4796_0[2]),.dinb(w_n5125_0[2]),.dout(n5126),.clk(gclk));
	jand g04881(.dina(n5126),.dinb(w_n5124_1[1]),.dout(n5127),.clk(gclk));
	jnot g04882(.din(n5127),.dout(n5128),.clk(gclk));
	jand g04883(.dina(n5128),.dinb(n5123),.dout(n5129),.clk(gclk));
	jor g04884(.dina(w_n5129_0[2]),.dinb(w_n5116_21[2]),.dout(n5130),.clk(gclk));
	jor g04885(.dina(w_n5121_29[0]),.dinb(w_a66_0[0]),.dout(n5131),.clk(gclk));
	jxor g04886(.dina(w_n5131_0[1]),.dinb(w_n4797_0[0]),.dout(n5132),.clk(gclk));
	jand g04887(.dina(w_n5129_0[1]),.dinb(w_n5116_21[1]),.dout(n5133),.clk(gclk));
	jor g04888(.dina(n5133),.dinb(w_n5132_0[1]),.dout(n5134),.clk(gclk));
	jand g04889(.dina(w_n5134_0[1]),.dinb(w_n5130_0[1]),.dout(n5135),.clk(gclk));
	jor g04890(.dina(n5135),.dinb(w_n4499_25[0]),.dout(n5136),.clk(gclk));
	jand g04891(.dina(w_n5130_0[0]),.dinb(w_n4499_24[2]),.dout(n5137),.clk(gclk));
	jand g04892(.dina(n5137),.dinb(w_n5134_0[0]),.dout(n5138),.clk(gclk));
	jor g04893(.dina(w_n5131_0[0]),.dinb(w_a67_0[0]),.dout(n5139),.clk(gclk));
	jnot g04894(.din(w_n5108_0[0]),.dout(n5140),.clk(gclk));
	jnot g04895(.din(w_n5110_0[0]),.dout(n5141),.clk(gclk));
	jor g04896(.dina(w_n5115_0[0]),.dinb(w_n5116_21[0]),.dout(n5142),.clk(gclk));
	jor g04897(.dina(n5142),.dinb(w_n5141_0[1]),.dout(n5143),.clk(gclk));
	jor g04898(.dina(n5143),.dinb(n5140),.dout(n5144),.clk(gclk));
	jand g04899(.dina(n5144),.dinb(n5139),.dout(n5145),.clk(gclk));
	jxor g04900(.dina(n5145),.dinb(w_n4502_0[1]),.dout(n5146),.clk(gclk));
	jor g04901(.dina(w_n5146_0[1]),.dinb(w_n5138_0[1]),.dout(n5147),.clk(gclk));
	jand g04902(.dina(n5147),.dinb(w_n5136_0[1]),.dout(n5148),.clk(gclk));
	jor g04903(.dina(w_n5148_0[2]),.dinb(w_n4494_22[0]),.dout(n5149),.clk(gclk));
	jand g04904(.dina(w_n5148_0[1]),.dinb(w_n4494_21[2]),.dout(n5150),.clk(gclk));
	jxor g04905(.dina(w_n4800_0[0]),.dinb(w_n4499_24[1]),.dout(n5151),.clk(gclk));
	jor g04906(.dina(n5151),.dinb(w_n5121_28[2]),.dout(n5152),.clk(gclk));
	jxor g04907(.dina(n5152),.dinb(w_n4803_0[0]),.dout(n5153),.clk(gclk));
	jor g04908(.dina(w_n5153_0[1]),.dinb(n5150),.dout(n5154),.clk(gclk));
	jand g04909(.dina(w_n5154_0[1]),.dinb(w_n5149_0[1]),.dout(n5155),.clk(gclk));
	jor g04910(.dina(n5155),.dinb(w_n3912_25[0]),.dout(n5156),.clk(gclk));
	jnot g04911(.din(w_n4809_0[0]),.dout(n5157),.clk(gclk));
	jor g04912(.dina(n5157),.dinb(w_n4807_0[0]),.dout(n5158),.clk(gclk));
	jor g04913(.dina(n5158),.dinb(w_n5121_28[1]),.dout(n5159),.clk(gclk));
	jxor g04914(.dina(n5159),.dinb(w_n4818_0[0]),.dout(n5160),.clk(gclk));
	jand g04915(.dina(w_n5149_0[0]),.dinb(w_n3912_24[2]),.dout(n5161),.clk(gclk));
	jand g04916(.dina(n5161),.dinb(w_n5154_0[0]),.dout(n5162),.clk(gclk));
	jor g04917(.dina(w_n5162_0[1]),.dinb(w_n5160_0[1]),.dout(n5163),.clk(gclk));
	jand g04918(.dina(w_n5163_0[1]),.dinb(w_n5156_0[1]),.dout(n5164),.clk(gclk));
	jor g04919(.dina(w_n5164_0[2]),.dinb(w_n3907_22[0]),.dout(n5165),.clk(gclk));
	jand g04920(.dina(w_n5164_0[1]),.dinb(w_n3907_21[2]),.dout(n5166),.clk(gclk));
	jxor g04921(.dina(w_n4820_0[0]),.dinb(w_n3912_24[1]),.dout(n5167),.clk(gclk));
	jor g04922(.dina(n5167),.dinb(w_n5121_28[0]),.dout(n5168),.clk(gclk));
	jxor g04923(.dina(n5168),.dinb(w_n4825_0[0]),.dout(n5169),.clk(gclk));
	jnot g04924(.din(w_n5169_0[1]),.dout(n5170),.clk(gclk));
	jor g04925(.dina(n5170),.dinb(n5166),.dout(n5171),.clk(gclk));
	jand g04926(.dina(w_n5171_0[1]),.dinb(w_n5165_0[1]),.dout(n5172),.clk(gclk));
	jor g04927(.dina(n5172),.dinb(w_n3376_25[2]),.dout(n5173),.clk(gclk));
	jand g04928(.dina(w_n5165_0[0]),.dinb(w_n3376_25[1]),.dout(n5174),.clk(gclk));
	jand g04929(.dina(n5174),.dinb(w_n5171_0[0]),.dout(n5175),.clk(gclk));
	jnot g04930(.din(w_n4829_0[0]),.dout(n5176),.clk(gclk));
	jand g04931(.dina(w_asqrt33_22[1]),.dinb(n5176),.dout(n5177),.clk(gclk));
	jand g04932(.dina(w_n5177_0[1]),.dinb(w_n4836_0[0]),.dout(n5178),.clk(gclk));
	jor g04933(.dina(n5178),.dinb(w_n4834_0[0]),.dout(n5179),.clk(gclk));
	jand g04934(.dina(w_n5177_0[0]),.dinb(w_n4837_0[0]),.dout(n5180),.clk(gclk));
	jnot g04935(.din(n5180),.dout(n5181),.clk(gclk));
	jand g04936(.dina(n5181),.dinb(n5179),.dout(n5182),.clk(gclk));
	jnot g04937(.din(n5182),.dout(n5183),.clk(gclk));
	jor g04938(.dina(w_n5183_0[1]),.dinb(w_n5175_0[1]),.dout(n5184),.clk(gclk));
	jand g04939(.dina(n5184),.dinb(w_n5173_0[1]),.dout(n5185),.clk(gclk));
	jor g04940(.dina(w_n5185_0[2]),.dinb(w_n3371_22[1]),.dout(n5186),.clk(gclk));
	jand g04941(.dina(w_n5185_0[1]),.dinb(w_n3371_22[0]),.dout(n5187),.clk(gclk));
	jnot g04942(.din(w_n4844_0[0]),.dout(n5188),.clk(gclk));
	jxor g04943(.dina(w_n4838_0[0]),.dinb(w_n3376_25[0]),.dout(n5189),.clk(gclk));
	jor g04944(.dina(n5189),.dinb(w_n5121_27[2]),.dout(n5190),.clk(gclk));
	jxor g04945(.dina(n5190),.dinb(n5188),.dout(n5191),.clk(gclk));
	jnot g04946(.din(w_n5191_0[1]),.dout(n5192),.clk(gclk));
	jor g04947(.dina(n5192),.dinb(n5187),.dout(n5193),.clk(gclk));
	jand g04948(.dina(w_n5193_0[1]),.dinb(w_n5186_0[1]),.dout(n5194),.clk(gclk));
	jor g04949(.dina(n5194),.dinb(w_n2875_25[1]),.dout(n5195),.clk(gclk));
	jnot g04950(.din(w_n4849_0[0]),.dout(n5196),.clk(gclk));
	jor g04951(.dina(n5196),.dinb(w_n4847_0[0]),.dout(n5197),.clk(gclk));
	jor g04952(.dina(n5197),.dinb(w_n5121_27[1]),.dout(n5198),.clk(gclk));
	jxor g04953(.dina(n5198),.dinb(w_n4858_0[0]),.dout(n5199),.clk(gclk));
	jand g04954(.dina(w_n5186_0[0]),.dinb(w_n2875_25[0]),.dout(n5200),.clk(gclk));
	jand g04955(.dina(n5200),.dinb(w_n5193_0[0]),.dout(n5201),.clk(gclk));
	jor g04956(.dina(w_n5201_0[1]),.dinb(w_n5199_0[1]),.dout(n5202),.clk(gclk));
	jand g04957(.dina(w_n5202_0[1]),.dinb(w_n5195_0[1]),.dout(n5203),.clk(gclk));
	jor g04958(.dina(w_n5203_0[2]),.dinb(w_n2870_22[1]),.dout(n5204),.clk(gclk));
	jand g04959(.dina(w_n5203_0[1]),.dinb(w_n2870_22[0]),.dout(n5205),.clk(gclk));
	jnot g04960(.din(w_n4865_0[0]),.dout(n5206),.clk(gclk));
	jxor g04961(.dina(w_n4860_0[0]),.dinb(w_n2875_24[2]),.dout(n5207),.clk(gclk));
	jor g04962(.dina(n5207),.dinb(w_n5121_27[0]),.dout(n5208),.clk(gclk));
	jxor g04963(.dina(n5208),.dinb(n5206),.dout(n5209),.clk(gclk));
	jnot g04964(.din(n5209),.dout(n5210),.clk(gclk));
	jor g04965(.dina(w_n5210_0[1]),.dinb(n5205),.dout(n5211),.clk(gclk));
	jand g04966(.dina(w_n5211_0[1]),.dinb(w_n5204_0[1]),.dout(n5212),.clk(gclk));
	jor g04967(.dina(n5212),.dinb(w_n2425_25[2]),.dout(n5213),.clk(gclk));
	jand g04968(.dina(w_n5204_0[0]),.dinb(w_n2425_25[1]),.dout(n5214),.clk(gclk));
	jand g04969(.dina(n5214),.dinb(w_n5211_0[0]),.dout(n5215),.clk(gclk));
	jnot g04970(.din(w_n4868_0[0]),.dout(n5216),.clk(gclk));
	jand g04971(.dina(w_asqrt33_22[0]),.dinb(n5216),.dout(n5217),.clk(gclk));
	jand g04972(.dina(w_n5217_0[1]),.dinb(w_n4875_0[0]),.dout(n5218),.clk(gclk));
	jor g04973(.dina(n5218),.dinb(w_n4873_0[0]),.dout(n5219),.clk(gclk));
	jand g04974(.dina(w_n5217_0[0]),.dinb(w_n4876_0[0]),.dout(n5220),.clk(gclk));
	jnot g04975(.din(n5220),.dout(n5221),.clk(gclk));
	jand g04976(.dina(n5221),.dinb(n5219),.dout(n5222),.clk(gclk));
	jnot g04977(.din(n5222),.dout(n5223),.clk(gclk));
	jor g04978(.dina(w_n5223_0[1]),.dinb(w_n5215_0[1]),.dout(n5224),.clk(gclk));
	jand g04979(.dina(n5224),.dinb(w_n5213_0[1]),.dout(n5225),.clk(gclk));
	jor g04980(.dina(w_n5225_0[1]),.dinb(w_n2420_23[0]),.dout(n5226),.clk(gclk));
	jxor g04981(.dina(w_n4877_0[0]),.dinb(w_n2425_25[0]),.dout(n5227),.clk(gclk));
	jor g04982(.dina(n5227),.dinb(w_n5121_26[2]),.dout(n5228),.clk(gclk));
	jxor g04983(.dina(n5228),.dinb(w_n4882_0[0]),.dout(n5229),.clk(gclk));
	jand g04984(.dina(w_n5225_0[0]),.dinb(w_n2420_22[2]),.dout(n5230),.clk(gclk));
	jor g04985(.dina(w_n5230_0[1]),.dinb(w_n5229_0[1]),.dout(n5231),.clk(gclk));
	jand g04986(.dina(w_n5231_0[2]),.dinb(w_n5226_0[2]),.dout(n5232),.clk(gclk));
	jor g04987(.dina(n5232),.dinb(w_n2010_25[1]),.dout(n5233),.clk(gclk));
	jnot g04988(.din(w_n4887_0[0]),.dout(n5234),.clk(gclk));
	jor g04989(.dina(n5234),.dinb(w_n4885_0[0]),.dout(n5235),.clk(gclk));
	jor g04990(.dina(n5235),.dinb(w_n5121_26[1]),.dout(n5236),.clk(gclk));
	jxor g04991(.dina(n5236),.dinb(w_n4896_0[0]),.dout(n5237),.clk(gclk));
	jand g04992(.dina(w_n5226_0[1]),.dinb(w_n2010_25[0]),.dout(n5238),.clk(gclk));
	jand g04993(.dina(n5238),.dinb(w_n5231_0[1]),.dout(n5239),.clk(gclk));
	jor g04994(.dina(w_n5239_0[1]),.dinb(w_n5237_0[1]),.dout(n5240),.clk(gclk));
	jand g04995(.dina(w_n5240_0[1]),.dinb(w_n5233_0[1]),.dout(n5241),.clk(gclk));
	jor g04996(.dina(w_n5241_0[2]),.dinb(w_n2005_23[1]),.dout(n5242),.clk(gclk));
	jand g04997(.dina(w_n5241_0[1]),.dinb(w_n2005_23[0]),.dout(n5243),.clk(gclk));
	jnot g04998(.din(w_n4899_0[0]),.dout(n5244),.clk(gclk));
	jand g04999(.dina(w_asqrt33_21[2]),.dinb(n5244),.dout(n5245),.clk(gclk));
	jand g05000(.dina(w_n5245_0[1]),.dinb(w_n4904_0[0]),.dout(n5246),.clk(gclk));
	jor g05001(.dina(n5246),.dinb(w_n4903_0[0]),.dout(n5247),.clk(gclk));
	jand g05002(.dina(w_n5245_0[0]),.dinb(w_n4905_0[0]),.dout(n5248),.clk(gclk));
	jnot g05003(.din(n5248),.dout(n5249),.clk(gclk));
	jand g05004(.dina(n5249),.dinb(n5247),.dout(n5250),.clk(gclk));
	jnot g05005(.din(n5250),.dout(n5251),.clk(gclk));
	jor g05006(.dina(w_n5251_0[1]),.dinb(n5243),.dout(n5252),.clk(gclk));
	jand g05007(.dina(w_n5252_0[1]),.dinb(w_n5242_0[1]),.dout(n5253),.clk(gclk));
	jor g05008(.dina(n5253),.dinb(w_n1646_26[1]),.dout(n5254),.clk(gclk));
	jand g05009(.dina(w_n5242_0[0]),.dinb(w_n1646_26[0]),.dout(n5255),.clk(gclk));
	jand g05010(.dina(n5255),.dinb(w_n5252_0[0]),.dout(n5256),.clk(gclk));
	jnot g05011(.din(w_n4907_0[0]),.dout(n5257),.clk(gclk));
	jand g05012(.dina(w_asqrt33_21[1]),.dinb(n5257),.dout(n5258),.clk(gclk));
	jand g05013(.dina(w_n5258_0[1]),.dinb(w_n4914_0[0]),.dout(n5259),.clk(gclk));
	jor g05014(.dina(n5259),.dinb(w_n4912_0[0]),.dout(n5260),.clk(gclk));
	jand g05015(.dina(w_n5258_0[0]),.dinb(w_n4915_0[0]),.dout(n5261),.clk(gclk));
	jnot g05016(.din(n5261),.dout(n5262),.clk(gclk));
	jand g05017(.dina(n5262),.dinb(n5260),.dout(n5263),.clk(gclk));
	jnot g05018(.din(n5263),.dout(n5264),.clk(gclk));
	jor g05019(.dina(w_n5264_0[1]),.dinb(w_n5256_0[1]),.dout(n5265),.clk(gclk));
	jand g05020(.dina(n5265),.dinb(w_n5254_0[1]),.dout(n5266),.clk(gclk));
	jor g05021(.dina(w_n5266_0[1]),.dinb(w_n1641_23[2]),.dout(n5267),.clk(gclk));
	jxor g05022(.dina(w_n4916_0[0]),.dinb(w_n1646_25[2]),.dout(n5268),.clk(gclk));
	jor g05023(.dina(n5268),.dinb(w_n5121_26[0]),.dout(n5269),.clk(gclk));
	jxor g05024(.dina(n5269),.dinb(w_n4927_0[0]),.dout(n5270),.clk(gclk));
	jand g05025(.dina(w_n5266_0[0]),.dinb(w_n1641_23[1]),.dout(n5271),.clk(gclk));
	jor g05026(.dina(w_n5271_0[1]),.dinb(w_n5270_0[1]),.dout(n5272),.clk(gclk));
	jand g05027(.dina(w_n5272_0[2]),.dinb(w_n5267_0[2]),.dout(n5273),.clk(gclk));
	jor g05028(.dina(n5273),.dinb(w_n1317_26[0]),.dout(n5274),.clk(gclk));
	jnot g05029(.din(w_n4932_0[0]),.dout(n5275),.clk(gclk));
	jor g05030(.dina(n5275),.dinb(w_n4930_0[0]),.dout(n5276),.clk(gclk));
	jor g05031(.dina(n5276),.dinb(w_n5121_25[2]),.dout(n5277),.clk(gclk));
	jxor g05032(.dina(n5277),.dinb(w_n4941_0[0]),.dout(n5278),.clk(gclk));
	jand g05033(.dina(w_n5267_0[1]),.dinb(w_n1317_25[2]),.dout(n5279),.clk(gclk));
	jand g05034(.dina(n5279),.dinb(w_n5272_0[1]),.dout(n5280),.clk(gclk));
	jor g05035(.dina(w_n5280_0[1]),.dinb(w_n5278_0[1]),.dout(n5281),.clk(gclk));
	jand g05036(.dina(w_n5281_0[1]),.dinb(w_n5274_0[1]),.dout(n5282),.clk(gclk));
	jor g05037(.dina(w_n5282_0[2]),.dinb(w_n1312_24[0]),.dout(n5283),.clk(gclk));
	jand g05038(.dina(w_n5282_0[1]),.dinb(w_n1312_23[2]),.dout(n5284),.clk(gclk));
	jnot g05039(.din(w_n4944_0[0]),.dout(n5285),.clk(gclk));
	jand g05040(.dina(w_asqrt33_21[0]),.dinb(n5285),.dout(n5286),.clk(gclk));
	jand g05041(.dina(w_n5286_0[1]),.dinb(w_n4949_0[0]),.dout(n5287),.clk(gclk));
	jor g05042(.dina(n5287),.dinb(w_n4948_0[0]),.dout(n5288),.clk(gclk));
	jand g05043(.dina(w_n5286_0[0]),.dinb(w_n4950_0[0]),.dout(n5289),.clk(gclk));
	jnot g05044(.din(n5289),.dout(n5290),.clk(gclk));
	jand g05045(.dina(n5290),.dinb(n5288),.dout(n5291),.clk(gclk));
	jnot g05046(.din(n5291),.dout(n5292),.clk(gclk));
	jor g05047(.dina(w_n5292_0[1]),.dinb(n5284),.dout(n5293),.clk(gclk));
	jand g05048(.dina(w_n5293_0[1]),.dinb(w_n5283_0[1]),.dout(n5294),.clk(gclk));
	jor g05049(.dina(n5294),.dinb(w_n1039_26[2]),.dout(n5295),.clk(gclk));
	jand g05050(.dina(w_n5283_0[0]),.dinb(w_n1039_26[1]),.dout(n5296),.clk(gclk));
	jand g05051(.dina(n5296),.dinb(w_n5293_0[0]),.dout(n5297),.clk(gclk));
	jnot g05052(.din(w_n4952_0[0]),.dout(n5298),.clk(gclk));
	jand g05053(.dina(w_asqrt33_20[2]),.dinb(n5298),.dout(n5299),.clk(gclk));
	jand g05054(.dina(w_n5299_0[1]),.dinb(w_n4959_0[0]),.dout(n5300),.clk(gclk));
	jor g05055(.dina(n5300),.dinb(w_n4957_0[0]),.dout(n5301),.clk(gclk));
	jand g05056(.dina(w_n5299_0[0]),.dinb(w_n4960_0[0]),.dout(n5302),.clk(gclk));
	jnot g05057(.din(n5302),.dout(n5303),.clk(gclk));
	jand g05058(.dina(n5303),.dinb(n5301),.dout(n5304),.clk(gclk));
	jnot g05059(.din(n5304),.dout(n5305),.clk(gclk));
	jor g05060(.dina(w_n5305_0[1]),.dinb(w_n5297_0[1]),.dout(n5306),.clk(gclk));
	jand g05061(.dina(n5306),.dinb(w_n5295_0[1]),.dout(n5307),.clk(gclk));
	jor g05062(.dina(w_n5307_0[1]),.dinb(w_n1034_24[2]),.dout(n5308),.clk(gclk));
	jxor g05063(.dina(w_n4961_0[0]),.dinb(w_n1039_26[0]),.dout(n5309),.clk(gclk));
	jor g05064(.dina(n5309),.dinb(w_n5121_25[1]),.dout(n5310),.clk(gclk));
	jxor g05065(.dina(n5310),.dinb(w_n4972_0[0]),.dout(n5311),.clk(gclk));
	jand g05066(.dina(w_n5307_0[0]),.dinb(w_n1034_24[1]),.dout(n5312),.clk(gclk));
	jor g05067(.dina(w_n5312_0[1]),.dinb(w_n5311_0[1]),.dout(n5313),.clk(gclk));
	jand g05068(.dina(w_n5313_0[2]),.dinb(w_n5308_0[2]),.dout(n5314),.clk(gclk));
	jor g05069(.dina(n5314),.dinb(w_n796_26[1]),.dout(n5315),.clk(gclk));
	jnot g05070(.din(w_n4977_0[0]),.dout(n5316),.clk(gclk));
	jor g05071(.dina(n5316),.dinb(w_n4975_0[0]),.dout(n5317),.clk(gclk));
	jor g05072(.dina(n5317),.dinb(w_n5121_25[0]),.dout(n5318),.clk(gclk));
	jxor g05073(.dina(n5318),.dinb(w_n4986_0[0]),.dout(n5319),.clk(gclk));
	jand g05074(.dina(w_n5308_0[1]),.dinb(w_n796_26[0]),.dout(n5320),.clk(gclk));
	jand g05075(.dina(n5320),.dinb(w_n5313_0[1]),.dout(n5321),.clk(gclk));
	jor g05076(.dina(w_n5321_0[1]),.dinb(w_n5319_0[1]),.dout(n5322),.clk(gclk));
	jand g05077(.dina(w_n5322_0[1]),.dinb(w_n5315_0[1]),.dout(n5323),.clk(gclk));
	jor g05078(.dina(w_n5323_0[2]),.dinb(w_n791_25[0]),.dout(n5324),.clk(gclk));
	jand g05079(.dina(w_n5323_0[1]),.dinb(w_n791_24[2]),.dout(n5325),.clk(gclk));
	jnot g05080(.din(w_n4989_0[0]),.dout(n5326),.clk(gclk));
	jand g05081(.dina(w_asqrt33_20[1]),.dinb(n5326),.dout(n5327),.clk(gclk));
	jand g05082(.dina(w_n5327_0[1]),.dinb(w_n4994_0[0]),.dout(n5328),.clk(gclk));
	jor g05083(.dina(n5328),.dinb(w_n4993_0[0]),.dout(n5329),.clk(gclk));
	jand g05084(.dina(w_n5327_0[0]),.dinb(w_n4995_0[0]),.dout(n5330),.clk(gclk));
	jnot g05085(.din(n5330),.dout(n5331),.clk(gclk));
	jand g05086(.dina(n5331),.dinb(n5329),.dout(n5332),.clk(gclk));
	jnot g05087(.din(n5332),.dout(n5333),.clk(gclk));
	jor g05088(.dina(w_n5333_0[1]),.dinb(n5325),.dout(n5334),.clk(gclk));
	jand g05089(.dina(w_n5334_0[1]),.dinb(w_n5324_0[1]),.dout(n5335),.clk(gclk));
	jor g05090(.dina(n5335),.dinb(w_n595_27[0]),.dout(n5336),.clk(gclk));
	jand g05091(.dina(w_n5324_0[0]),.dinb(w_n595_26[2]),.dout(n5337),.clk(gclk));
	jand g05092(.dina(n5337),.dinb(w_n5334_0[0]),.dout(n5338),.clk(gclk));
	jnot g05093(.din(w_n4997_0[0]),.dout(n5339),.clk(gclk));
	jand g05094(.dina(w_asqrt33_20[0]),.dinb(n5339),.dout(n5340),.clk(gclk));
	jand g05095(.dina(w_n5340_0[1]),.dinb(w_n5004_0[0]),.dout(n5341),.clk(gclk));
	jor g05096(.dina(n5341),.dinb(w_n5002_0[0]),.dout(n5342),.clk(gclk));
	jand g05097(.dina(w_n5340_0[0]),.dinb(w_n5005_0[0]),.dout(n5343),.clk(gclk));
	jnot g05098(.din(n5343),.dout(n5344),.clk(gclk));
	jand g05099(.dina(n5344),.dinb(n5342),.dout(n5345),.clk(gclk));
	jnot g05100(.din(n5345),.dout(n5346),.clk(gclk));
	jor g05101(.dina(w_n5346_0[1]),.dinb(w_n5338_0[1]),.dout(n5347),.clk(gclk));
	jand g05102(.dina(n5347),.dinb(w_n5336_0[1]),.dout(n5348),.clk(gclk));
	jor g05103(.dina(w_n5348_0[1]),.dinb(w_n590_25[1]),.dout(n5349),.clk(gclk));
	jxor g05104(.dina(w_n5006_0[0]),.dinb(w_n595_26[1]),.dout(n5350),.clk(gclk));
	jor g05105(.dina(n5350),.dinb(w_n5121_24[2]),.dout(n5351),.clk(gclk));
	jxor g05106(.dina(n5351),.dinb(w_n5017_0[0]),.dout(n5352),.clk(gclk));
	jand g05107(.dina(w_n5348_0[0]),.dinb(w_n590_25[0]),.dout(n5353),.clk(gclk));
	jor g05108(.dina(w_n5353_0[1]),.dinb(w_n5352_0[1]),.dout(n5354),.clk(gclk));
	jand g05109(.dina(w_n5354_0[2]),.dinb(w_n5349_0[2]),.dout(n5355),.clk(gclk));
	jor g05110(.dina(n5355),.dinb(w_n430_26[2]),.dout(n5356),.clk(gclk));
	jnot g05111(.din(w_n5022_0[0]),.dout(n5357),.clk(gclk));
	jor g05112(.dina(n5357),.dinb(w_n5020_0[0]),.dout(n5358),.clk(gclk));
	jor g05113(.dina(n5358),.dinb(w_n5121_24[1]),.dout(n5359),.clk(gclk));
	jxor g05114(.dina(n5359),.dinb(w_n5031_0[0]),.dout(n5360),.clk(gclk));
	jand g05115(.dina(w_n5349_0[1]),.dinb(w_n430_26[1]),.dout(n5361),.clk(gclk));
	jand g05116(.dina(n5361),.dinb(w_n5354_0[1]),.dout(n5362),.clk(gclk));
	jor g05117(.dina(w_n5362_0[1]),.dinb(w_n5360_0[1]),.dout(n5363),.clk(gclk));
	jand g05118(.dina(w_n5363_0[1]),.dinb(w_n5356_0[1]),.dout(n5364),.clk(gclk));
	jor g05119(.dina(w_n5364_0[2]),.dinb(w_n425_25[2]),.dout(n5365),.clk(gclk));
	jand g05120(.dina(w_n5364_0[1]),.dinb(w_n425_25[1]),.dout(n5366),.clk(gclk));
	jnot g05121(.din(w_n5034_0[0]),.dout(n5367),.clk(gclk));
	jand g05122(.dina(w_asqrt33_19[2]),.dinb(n5367),.dout(n5368),.clk(gclk));
	jand g05123(.dina(w_n5368_0[1]),.dinb(w_n5039_0[0]),.dout(n5369),.clk(gclk));
	jor g05124(.dina(n5369),.dinb(w_n5038_0[0]),.dout(n5370),.clk(gclk));
	jand g05125(.dina(w_n5368_0[0]),.dinb(w_n5040_0[0]),.dout(n5371),.clk(gclk));
	jnot g05126(.din(n5371),.dout(n5372),.clk(gclk));
	jand g05127(.dina(n5372),.dinb(n5370),.dout(n5373),.clk(gclk));
	jnot g05128(.din(n5373),.dout(n5374),.clk(gclk));
	jor g05129(.dina(w_n5374_0[1]),.dinb(n5366),.dout(n5375),.clk(gclk));
	jand g05130(.dina(w_n5375_0[1]),.dinb(w_n5365_0[1]),.dout(n5376),.clk(gclk));
	jor g05131(.dina(n5376),.dinb(w_n305_27[1]),.dout(n5377),.clk(gclk));
	jand g05132(.dina(w_n5365_0[0]),.dinb(w_n305_27[0]),.dout(n5378),.clk(gclk));
	jand g05133(.dina(n5378),.dinb(w_n5375_0[0]),.dout(n5379),.clk(gclk));
	jnot g05134(.din(w_n5042_0[0]),.dout(n5380),.clk(gclk));
	jand g05135(.dina(w_asqrt33_19[1]),.dinb(n5380),.dout(n5381),.clk(gclk));
	jand g05136(.dina(w_n5381_0[1]),.dinb(w_n5049_0[0]),.dout(n5382),.clk(gclk));
	jor g05137(.dina(n5382),.dinb(w_n5047_0[0]),.dout(n5383),.clk(gclk));
	jand g05138(.dina(w_n5381_0[0]),.dinb(w_n5050_0[0]),.dout(n5384),.clk(gclk));
	jnot g05139(.din(n5384),.dout(n5385),.clk(gclk));
	jand g05140(.dina(n5385),.dinb(n5383),.dout(n5386),.clk(gclk));
	jnot g05141(.din(n5386),.dout(n5387),.clk(gclk));
	jor g05142(.dina(w_n5387_0[1]),.dinb(w_n5379_0[1]),.dout(n5388),.clk(gclk));
	jand g05143(.dina(n5388),.dinb(w_n5377_0[1]),.dout(n5389),.clk(gclk));
	jor g05144(.dina(w_n5389_0[1]),.dinb(w_n290_26[2]),.dout(n5390),.clk(gclk));
	jxor g05145(.dina(w_n5051_0[0]),.dinb(w_n305_26[2]),.dout(n5391),.clk(gclk));
	jor g05146(.dina(n5391),.dinb(w_n5121_24[0]),.dout(n5392),.clk(gclk));
	jxor g05147(.dina(n5392),.dinb(w_n5062_0[0]),.dout(n5393),.clk(gclk));
	jand g05148(.dina(w_n5389_0[0]),.dinb(w_n290_26[1]),.dout(n5394),.clk(gclk));
	jor g05149(.dina(w_n5394_0[1]),.dinb(w_n5393_0[1]),.dout(n5395),.clk(gclk));
	jand g05150(.dina(w_n5395_0[2]),.dinb(w_n5390_0[2]),.dout(n5396),.clk(gclk));
	jor g05151(.dina(n5396),.dinb(w_n223_27[0]),.dout(n5397),.clk(gclk));
	jnot g05152(.din(w_n5067_0[0]),.dout(n5398),.clk(gclk));
	jor g05153(.dina(n5398),.dinb(w_n5065_0[0]),.dout(n5399),.clk(gclk));
	jor g05154(.dina(n5399),.dinb(w_n5121_23[2]),.dout(n5400),.clk(gclk));
	jxor g05155(.dina(n5400),.dinb(w_n5076_0[0]),.dout(n5401),.clk(gclk));
	jand g05156(.dina(w_n5390_0[1]),.dinb(w_n223_26[2]),.dout(n5402),.clk(gclk));
	jand g05157(.dina(n5402),.dinb(w_n5395_0[1]),.dout(n5403),.clk(gclk));
	jor g05158(.dina(w_n5403_0[1]),.dinb(w_n5401_0[1]),.dout(n5404),.clk(gclk));
	jand g05159(.dina(w_n5404_0[1]),.dinb(w_n5397_0[1]),.dout(n5405),.clk(gclk));
	jor g05160(.dina(w_n5405_0[2]),.dinb(w_n199_31[1]),.dout(n5406),.clk(gclk));
	jand g05161(.dina(w_n5405_0[1]),.dinb(w_n199_31[0]),.dout(n5407),.clk(gclk));
	jnot g05162(.din(w_n5079_0[0]),.dout(n5408),.clk(gclk));
	jand g05163(.dina(w_asqrt33_19[0]),.dinb(n5408),.dout(n5409),.clk(gclk));
	jand g05164(.dina(w_n5409_0[1]),.dinb(w_n5084_0[0]),.dout(n5410),.clk(gclk));
	jor g05165(.dina(n5410),.dinb(w_n5083_0[0]),.dout(n5411),.clk(gclk));
	jand g05166(.dina(w_n5409_0[0]),.dinb(w_n5085_0[0]),.dout(n5412),.clk(gclk));
	jnot g05167(.din(n5412),.dout(n5413),.clk(gclk));
	jand g05168(.dina(n5413),.dinb(n5411),.dout(n5414),.clk(gclk));
	jnot g05169(.din(n5414),.dout(n5415),.clk(gclk));
	jor g05170(.dina(w_n5415_0[1]),.dinb(n5407),.dout(n5416),.clk(gclk));
	jand g05171(.dina(n5416),.dinb(n5406),.dout(n5417),.clk(gclk));
	jnot g05172(.din(w_n5087_0[0]),.dout(n5418),.clk(gclk));
	jand g05173(.dina(w_asqrt33_18[2]),.dinb(n5418),.dout(n5419),.clk(gclk));
	jand g05174(.dina(w_n5419_0[1]),.dinb(w_n5094_0[0]),.dout(n5420),.clk(gclk));
	jor g05175(.dina(n5420),.dinb(w_n5092_0[0]),.dout(n5421),.clk(gclk));
	jand g05176(.dina(w_n5419_0[0]),.dinb(w_n5095_0[0]),.dout(n5422),.clk(gclk));
	jnot g05177(.din(n5422),.dout(n5423),.clk(gclk));
	jand g05178(.dina(n5423),.dinb(n5421),.dout(n5424),.clk(gclk));
	jnot g05179(.din(w_n5424_0[2]),.dout(n5425),.clk(gclk));
	jand g05180(.dina(w_asqrt33_18[1]),.dinb(w_n5109_0[1]),.dout(n5426),.clk(gclk));
	jand g05181(.dina(w_n5426_0[1]),.dinb(w_n5096_1[0]),.dout(n5427),.clk(gclk));
	jor g05182(.dina(n5427),.dinb(w_n5141_0[0]),.dout(n5428),.clk(gclk));
	jor g05183(.dina(n5428),.dinb(w_n5425_0[1]),.dout(n5429),.clk(gclk));
	jor g05184(.dina(n5429),.dinb(w_n5417_0[2]),.dout(n5430),.clk(gclk));
	jand g05185(.dina(n5430),.dinb(w_n194_30[1]),.dout(n5431),.clk(gclk));
	jand g05186(.dina(w_n5425_0[0]),.dinb(w_n5417_0[1]),.dout(n5432),.clk(gclk));
	jor g05187(.dina(w_n5426_0[0]),.dinb(w_n5096_0[2]),.dout(n5433),.clk(gclk));
	jand g05188(.dina(w_n5109_0[0]),.dinb(w_n5096_0[1]),.dout(n5434),.clk(gclk));
	jor g05189(.dina(n5434),.dinb(w_n194_30[0]),.dout(n5435),.clk(gclk));
	jnot g05190(.din(n5435),.dout(n5436),.clk(gclk));
	jand g05191(.dina(n5436),.dinb(n5433),.dout(n5437),.clk(gclk));
	jor g05192(.dina(w_n5437_0[1]),.dinb(w_n5432_0[2]),.dout(n5440),.clk(gclk));
	jor g05193(.dina(n5440),.dinb(w_n5431_0[1]),.dout(asqrt_fa_33),.clk(gclk));
	jand g05194(.dina(w_asqrt32_31),.dinb(w_a64_0[0]),.dout(n5442),.clk(gclk));
	jnot g05195(.din(w_a62_0[1]),.dout(n5443),.clk(gclk));
	jand g05196(.dina(w_n5124_1[0]),.dinb(w_n200_0[1]),.dout(n5444),.clk(gclk));
	jand g05197(.dina(n5444),.dinb(w_n5443_1[1]),.dout(n5445),.clk(gclk));
	jor g05198(.dina(n5445),.dinb(n5442),.dout(n5446),.clk(gclk));
	jand g05199(.dina(w_n5446_0[2]),.dinb(w_asqrt33_18[0]),.dout(n5447),.clk(gclk));
	jand g05200(.dina(w_asqrt32_30[2]),.dinb(w_n5124_0[2]),.dout(n5448),.clk(gclk));
	jxor g05201(.dina(w_n5448_0[1]),.dinb(w_n5125_0[1]),.dout(n5449),.clk(gclk));
	jor g05202(.dina(w_n5446_0[1]),.dinb(w_asqrt33_17[2]),.dout(n5450),.clk(gclk));
	jand g05203(.dina(n5450),.dinb(w_n5449_0[1]),.dout(n5451),.clk(gclk));
	jor g05204(.dina(w_n5451_0[1]),.dinb(w_n5447_0[1]),.dout(n5452),.clk(gclk));
	jand g05205(.dina(n5452),.dinb(w_asqrt34_20[2]),.dout(n5453),.clk(gclk));
	jor g05206(.dina(w_n5447_0[0]),.dinb(w_asqrt34_20[1]),.dout(n5454),.clk(gclk));
	jor g05207(.dina(n5454),.dinb(w_n5451_0[0]),.dout(n5455),.clk(gclk));
	jand g05208(.dina(w_n5448_0[0]),.dinb(w_n5125_0[0]),.dout(n5456),.clk(gclk));
	jnot g05209(.din(w_n5431_0[0]),.dout(n5457),.clk(gclk));
	jnot g05210(.din(w_n5432_0[1]),.dout(n5458),.clk(gclk));
	jnot g05211(.din(w_n5437_0[0]),.dout(n5459),.clk(gclk));
	jand g05212(.dina(n5459),.dinb(w_asqrt33_17[1]),.dout(n5460),.clk(gclk));
	jand g05213(.dina(n5460),.dinb(n5458),.dout(n5461),.clk(gclk));
	jand g05214(.dina(n5461),.dinb(n5457),.dout(n5462),.clk(gclk));
	jor g05215(.dina(n5462),.dinb(n5456),.dout(n5463),.clk(gclk));
	jxor g05216(.dina(n5463),.dinb(w_n4796_0[1]),.dout(n5464),.clk(gclk));
	jand g05217(.dina(w_n5464_0[1]),.dinb(w_n5455_0[1]),.dout(n5465),.clk(gclk));
	jor g05218(.dina(n5465),.dinb(w_n5453_0[1]),.dout(n5466),.clk(gclk));
	jand g05219(.dina(w_n5466_0[2]),.dinb(w_asqrt35_17[2]),.dout(n5467),.clk(gclk));
	jor g05220(.dina(w_n5466_0[1]),.dinb(w_asqrt35_17[1]),.dout(n5468),.clk(gclk));
	jxor g05221(.dina(w_n5129_0[0]),.dinb(w_n5116_20[2]),.dout(n5469),.clk(gclk));
	jand g05222(.dina(n5469),.dinb(w_asqrt32_30[1]),.dout(n5470),.clk(gclk));
	jxor g05223(.dina(n5470),.dinb(w_n5132_0[0]),.dout(n5471),.clk(gclk));
	jnot g05224(.din(w_n5471_0[1]),.dout(n5472),.clk(gclk));
	jand g05225(.dina(n5472),.dinb(n5468),.dout(n5473),.clk(gclk));
	jor g05226(.dina(w_n5473_0[1]),.dinb(w_n5467_0[1]),.dout(n5474),.clk(gclk));
	jand g05227(.dina(n5474),.dinb(w_asqrt36_20[2]),.dout(n5475),.clk(gclk));
	jnot g05228(.din(w_n5138_0[0]),.dout(n5476),.clk(gclk));
	jand g05229(.dina(n5476),.dinb(w_n5136_0[0]),.dout(n5477),.clk(gclk));
	jand g05230(.dina(n5477),.dinb(w_asqrt32_30[0]),.dout(n5478),.clk(gclk));
	jxor g05231(.dina(n5478),.dinb(w_n5146_0[0]),.dout(n5479),.clk(gclk));
	jnot g05232(.din(n5479),.dout(n5480),.clk(gclk));
	jor g05233(.dina(w_n5467_0[0]),.dinb(w_asqrt36_20[1]),.dout(n5481),.clk(gclk));
	jor g05234(.dina(n5481),.dinb(w_n5473_0[0]),.dout(n5482),.clk(gclk));
	jand g05235(.dina(w_n5482_0[1]),.dinb(w_n5480_0[1]),.dout(n5483),.clk(gclk));
	jor g05236(.dina(w_n5483_0[1]),.dinb(w_n5475_0[1]),.dout(n5484),.clk(gclk));
	jand g05237(.dina(w_n5484_0[2]),.dinb(w_asqrt37_18[0]),.dout(n5485),.clk(gclk));
	jor g05238(.dina(w_n5484_0[1]),.dinb(w_asqrt37_17[2]),.dout(n5486),.clk(gclk));
	jnot g05239(.din(w_n5153_0[0]),.dout(n5487),.clk(gclk));
	jxor g05240(.dina(w_n5148_0[0]),.dinb(w_n4494_21[1]),.dout(n5488),.clk(gclk));
	jand g05241(.dina(n5488),.dinb(w_asqrt32_29[2]),.dout(n5489),.clk(gclk));
	jxor g05242(.dina(n5489),.dinb(n5487),.dout(n5490),.clk(gclk));
	jand g05243(.dina(w_n5490_0[1]),.dinb(n5486),.dout(n5491),.clk(gclk));
	jor g05244(.dina(w_n5491_0[1]),.dinb(w_n5485_0[1]),.dout(n5492),.clk(gclk));
	jand g05245(.dina(n5492),.dinb(w_asqrt38_20[2]),.dout(n5493),.clk(gclk));
	jor g05246(.dina(w_n5485_0[0]),.dinb(w_asqrt38_20[1]),.dout(n5494),.clk(gclk));
	jor g05247(.dina(n5494),.dinb(w_n5491_0[0]),.dout(n5495),.clk(gclk));
	jnot g05248(.din(w_n5160_0[0]),.dout(n5496),.clk(gclk));
	jnot g05249(.din(w_n5162_0[0]),.dout(n5497),.clk(gclk));
	jand g05250(.dina(w_asqrt32_29[1]),.dinb(w_n5156_0[0]),.dout(n5498),.clk(gclk));
	jand g05251(.dina(w_n5498_0[1]),.dinb(n5497),.dout(n5499),.clk(gclk));
	jor g05252(.dina(n5499),.dinb(n5496),.dout(n5500),.clk(gclk));
	jnot g05253(.din(w_n5163_0[0]),.dout(n5501),.clk(gclk));
	jand g05254(.dina(w_n5498_0[0]),.dinb(n5501),.dout(n5502),.clk(gclk));
	jnot g05255(.din(n5502),.dout(n5503),.clk(gclk));
	jand g05256(.dina(n5503),.dinb(n5500),.dout(n5504),.clk(gclk));
	jand g05257(.dina(w_n5504_0[1]),.dinb(w_n5495_0[1]),.dout(n5505),.clk(gclk));
	jor g05258(.dina(n5505),.dinb(w_n5493_0[1]),.dout(n5506),.clk(gclk));
	jand g05259(.dina(w_n5506_0[2]),.dinb(w_asqrt39_18[0]),.dout(n5507),.clk(gclk));
	jor g05260(.dina(w_n5506_0[1]),.dinb(w_asqrt39_17[2]),.dout(n5508),.clk(gclk));
	jxor g05261(.dina(w_n5164_0[0]),.dinb(w_n3907_21[1]),.dout(n5509),.clk(gclk));
	jand g05262(.dina(n5509),.dinb(w_asqrt32_29[0]),.dout(n5510),.clk(gclk));
	jxor g05263(.dina(n5510),.dinb(w_n5169_0[0]),.dout(n5511),.clk(gclk));
	jand g05264(.dina(w_n5511_0[1]),.dinb(n5508),.dout(n5512),.clk(gclk));
	jor g05265(.dina(w_n5512_0[1]),.dinb(w_n5507_0[1]),.dout(n5513),.clk(gclk));
	jand g05266(.dina(n5513),.dinb(w_asqrt40_20[2]),.dout(n5514),.clk(gclk));
	jnot g05267(.din(w_n5175_0[0]),.dout(n5515),.clk(gclk));
	jand g05268(.dina(n5515),.dinb(w_n5173_0[0]),.dout(n5516),.clk(gclk));
	jand g05269(.dina(n5516),.dinb(w_asqrt32_28[2]),.dout(n5517),.clk(gclk));
	jxor g05270(.dina(n5517),.dinb(w_n5183_0[0]),.dout(n5518),.clk(gclk));
	jnot g05271(.din(n5518),.dout(n5519),.clk(gclk));
	jor g05272(.dina(w_n5507_0[0]),.dinb(w_asqrt40_20[1]),.dout(n5520),.clk(gclk));
	jor g05273(.dina(n5520),.dinb(w_n5512_0[0]),.dout(n5521),.clk(gclk));
	jand g05274(.dina(w_n5521_0[1]),.dinb(w_n5519_0[1]),.dout(n5522),.clk(gclk));
	jor g05275(.dina(w_n5522_0[1]),.dinb(w_n5514_0[1]),.dout(n5523),.clk(gclk));
	jand g05276(.dina(w_n5523_0[2]),.dinb(w_asqrt41_18[1]),.dout(n5524),.clk(gclk));
	jor g05277(.dina(w_n5523_0[1]),.dinb(w_asqrt41_18[0]),.dout(n5525),.clk(gclk));
	jxor g05278(.dina(w_n5185_0[0]),.dinb(w_n3371_21[2]),.dout(n5526),.clk(gclk));
	jand g05279(.dina(n5526),.dinb(w_asqrt32_28[1]),.dout(n5527),.clk(gclk));
	jxor g05280(.dina(n5527),.dinb(w_n5191_0[0]),.dout(n5528),.clk(gclk));
	jand g05281(.dina(w_n5528_0[1]),.dinb(n5525),.dout(n5529),.clk(gclk));
	jor g05282(.dina(w_n5529_0[1]),.dinb(w_n5524_0[1]),.dout(n5530),.clk(gclk));
	jand g05283(.dina(n5530),.dinb(w_asqrt42_20[2]),.dout(n5531),.clk(gclk));
	jor g05284(.dina(w_n5524_0[0]),.dinb(w_asqrt42_20[1]),.dout(n5532),.clk(gclk));
	jor g05285(.dina(n5532),.dinb(w_n5529_0[0]),.dout(n5533),.clk(gclk));
	jnot g05286(.din(w_n5199_0[0]),.dout(n5534),.clk(gclk));
	jnot g05287(.din(w_n5201_0[0]),.dout(n5535),.clk(gclk));
	jand g05288(.dina(w_asqrt32_28[0]),.dinb(w_n5195_0[0]),.dout(n5536),.clk(gclk));
	jand g05289(.dina(w_n5536_0[1]),.dinb(n5535),.dout(n5537),.clk(gclk));
	jor g05290(.dina(n5537),.dinb(n5534),.dout(n5538),.clk(gclk));
	jnot g05291(.din(w_n5202_0[0]),.dout(n5539),.clk(gclk));
	jand g05292(.dina(w_n5536_0[0]),.dinb(n5539),.dout(n5540),.clk(gclk));
	jnot g05293(.din(n5540),.dout(n5541),.clk(gclk));
	jand g05294(.dina(n5541),.dinb(n5538),.dout(n5542),.clk(gclk));
	jand g05295(.dina(w_n5542_0[1]),.dinb(w_n5533_0[1]),.dout(n5543),.clk(gclk));
	jor g05296(.dina(n5543),.dinb(w_n5531_0[1]),.dout(n5544),.clk(gclk));
	jand g05297(.dina(w_n5544_0[1]),.dinb(w_asqrt43_18[1]),.dout(n5545),.clk(gclk));
	jxor g05298(.dina(w_n5203_0[0]),.dinb(w_n2870_21[2]),.dout(n5546),.clk(gclk));
	jand g05299(.dina(n5546),.dinb(w_asqrt32_27[2]),.dout(n5547),.clk(gclk));
	jxor g05300(.dina(n5547),.dinb(w_n5210_0[0]),.dout(n5548),.clk(gclk));
	jnot g05301(.din(n5548),.dout(n5549),.clk(gclk));
	jor g05302(.dina(w_n5544_0[0]),.dinb(w_asqrt43_18[0]),.dout(n5550),.clk(gclk));
	jand g05303(.dina(w_n5550_0[1]),.dinb(w_n5549_0[1]),.dout(n5551),.clk(gclk));
	jor g05304(.dina(w_n5551_0[2]),.dinb(w_n5545_0[2]),.dout(n5552),.clk(gclk));
	jand g05305(.dina(n5552),.dinb(w_asqrt44_20[2]),.dout(n5553),.clk(gclk));
	jnot g05306(.din(w_n5215_0[0]),.dout(n5554),.clk(gclk));
	jand g05307(.dina(n5554),.dinb(w_n5213_0[0]),.dout(n5555),.clk(gclk));
	jand g05308(.dina(n5555),.dinb(w_asqrt32_27[1]),.dout(n5556),.clk(gclk));
	jxor g05309(.dina(n5556),.dinb(w_n5223_0[0]),.dout(n5557),.clk(gclk));
	jnot g05310(.din(n5557),.dout(n5558),.clk(gclk));
	jor g05311(.dina(w_n5545_0[1]),.dinb(w_asqrt44_20[1]),.dout(n5559),.clk(gclk));
	jor g05312(.dina(n5559),.dinb(w_n5551_0[1]),.dout(n5560),.clk(gclk));
	jand g05313(.dina(w_n5560_0[1]),.dinb(w_n5558_0[1]),.dout(n5561),.clk(gclk));
	jor g05314(.dina(w_n5561_0[1]),.dinb(w_n5553_0[1]),.dout(n5562),.clk(gclk));
	jand g05315(.dina(w_n5562_0[2]),.dinb(w_asqrt45_18[2]),.dout(n5563),.clk(gclk));
	jor g05316(.dina(w_n5562_0[1]),.dinb(w_asqrt45_18[1]),.dout(n5564),.clk(gclk));
	jnot g05317(.din(w_n5229_0[0]),.dout(n5565),.clk(gclk));
	jnot g05318(.din(w_n5230_0[0]),.dout(n5566),.clk(gclk));
	jand g05319(.dina(w_asqrt32_27[0]),.dinb(w_n5226_0[0]),.dout(n5567),.clk(gclk));
	jand g05320(.dina(w_n5567_0[1]),.dinb(n5566),.dout(n5568),.clk(gclk));
	jor g05321(.dina(n5568),.dinb(n5565),.dout(n5569),.clk(gclk));
	jnot g05322(.din(w_n5231_0[0]),.dout(n5570),.clk(gclk));
	jand g05323(.dina(w_n5567_0[0]),.dinb(n5570),.dout(n5571),.clk(gclk));
	jnot g05324(.din(n5571),.dout(n5572),.clk(gclk));
	jand g05325(.dina(n5572),.dinb(n5569),.dout(n5573),.clk(gclk));
	jand g05326(.dina(w_n5573_0[1]),.dinb(n5564),.dout(n5574),.clk(gclk));
	jor g05327(.dina(w_n5574_0[1]),.dinb(w_n5563_0[1]),.dout(n5575),.clk(gclk));
	jand g05328(.dina(n5575),.dinb(w_asqrt46_20[2]),.dout(n5576),.clk(gclk));
	jor g05329(.dina(w_n5563_0[0]),.dinb(w_asqrt46_20[1]),.dout(n5577),.clk(gclk));
	jor g05330(.dina(n5577),.dinb(w_n5574_0[0]),.dout(n5578),.clk(gclk));
	jnot g05331(.din(w_n5237_0[0]),.dout(n5579),.clk(gclk));
	jnot g05332(.din(w_n5239_0[0]),.dout(n5580),.clk(gclk));
	jand g05333(.dina(w_asqrt32_26[2]),.dinb(w_n5233_0[0]),.dout(n5581),.clk(gclk));
	jand g05334(.dina(w_n5581_0[1]),.dinb(n5580),.dout(n5582),.clk(gclk));
	jor g05335(.dina(n5582),.dinb(n5579),.dout(n5583),.clk(gclk));
	jnot g05336(.din(w_n5240_0[0]),.dout(n5584),.clk(gclk));
	jand g05337(.dina(w_n5581_0[0]),.dinb(n5584),.dout(n5585),.clk(gclk));
	jnot g05338(.din(n5585),.dout(n5586),.clk(gclk));
	jand g05339(.dina(n5586),.dinb(n5583),.dout(n5587),.clk(gclk));
	jand g05340(.dina(w_n5587_0[1]),.dinb(w_n5578_0[1]),.dout(n5588),.clk(gclk));
	jor g05341(.dina(n5588),.dinb(w_n5576_0[1]),.dout(n5589),.clk(gclk));
	jand g05342(.dina(w_n5589_0[1]),.dinb(w_asqrt47_18[2]),.dout(n5590),.clk(gclk));
	jxor g05343(.dina(w_n5241_0[0]),.dinb(w_n2005_22[2]),.dout(n5591),.clk(gclk));
	jand g05344(.dina(n5591),.dinb(w_asqrt32_26[1]),.dout(n5592),.clk(gclk));
	jxor g05345(.dina(n5592),.dinb(w_n5251_0[0]),.dout(n5593),.clk(gclk));
	jnot g05346(.din(n5593),.dout(n5594),.clk(gclk));
	jor g05347(.dina(w_n5589_0[0]),.dinb(w_asqrt47_18[1]),.dout(n5595),.clk(gclk));
	jand g05348(.dina(w_n5595_0[1]),.dinb(w_n5594_0[1]),.dout(n5596),.clk(gclk));
	jor g05349(.dina(w_n5596_0[2]),.dinb(w_n5590_0[2]),.dout(n5597),.clk(gclk));
	jand g05350(.dina(n5597),.dinb(w_asqrt48_20[2]),.dout(n5598),.clk(gclk));
	jnot g05351(.din(w_n5256_0[0]),.dout(n5599),.clk(gclk));
	jand g05352(.dina(n5599),.dinb(w_n5254_0[0]),.dout(n5600),.clk(gclk));
	jand g05353(.dina(n5600),.dinb(w_asqrt32_26[0]),.dout(n5601),.clk(gclk));
	jxor g05354(.dina(n5601),.dinb(w_n5264_0[0]),.dout(n5602),.clk(gclk));
	jnot g05355(.din(n5602),.dout(n5603),.clk(gclk));
	jor g05356(.dina(w_n5590_0[1]),.dinb(w_asqrt48_20[1]),.dout(n5604),.clk(gclk));
	jor g05357(.dina(n5604),.dinb(w_n5596_0[1]),.dout(n5605),.clk(gclk));
	jand g05358(.dina(w_n5605_0[1]),.dinb(w_n5603_0[1]),.dout(n5606),.clk(gclk));
	jor g05359(.dina(w_n5606_0[1]),.dinb(w_n5598_0[1]),.dout(n5607),.clk(gclk));
	jand g05360(.dina(w_n5607_0[2]),.dinb(w_asqrt49_19[0]),.dout(n5608),.clk(gclk));
	jor g05361(.dina(w_n5607_0[1]),.dinb(w_asqrt49_18[2]),.dout(n5609),.clk(gclk));
	jnot g05362(.din(w_n5270_0[0]),.dout(n5610),.clk(gclk));
	jnot g05363(.din(w_n5271_0[0]),.dout(n5611),.clk(gclk));
	jand g05364(.dina(w_asqrt32_25[2]),.dinb(w_n5267_0[0]),.dout(n5612),.clk(gclk));
	jand g05365(.dina(w_n5612_0[1]),.dinb(n5611),.dout(n5613),.clk(gclk));
	jor g05366(.dina(n5613),.dinb(n5610),.dout(n5614),.clk(gclk));
	jnot g05367(.din(w_n5272_0[0]),.dout(n5615),.clk(gclk));
	jand g05368(.dina(w_n5612_0[0]),.dinb(n5615),.dout(n5616),.clk(gclk));
	jnot g05369(.din(n5616),.dout(n5617),.clk(gclk));
	jand g05370(.dina(n5617),.dinb(n5614),.dout(n5618),.clk(gclk));
	jand g05371(.dina(w_n5618_0[1]),.dinb(n5609),.dout(n5619),.clk(gclk));
	jor g05372(.dina(w_n5619_0[1]),.dinb(w_n5608_0[1]),.dout(n5620),.clk(gclk));
	jand g05373(.dina(n5620),.dinb(w_asqrt50_20[2]),.dout(n5621),.clk(gclk));
	jor g05374(.dina(w_n5608_0[0]),.dinb(w_asqrt50_20[1]),.dout(n5622),.clk(gclk));
	jor g05375(.dina(n5622),.dinb(w_n5619_0[0]),.dout(n5623),.clk(gclk));
	jnot g05376(.din(w_n5278_0[0]),.dout(n5624),.clk(gclk));
	jnot g05377(.din(w_n5280_0[0]),.dout(n5625),.clk(gclk));
	jand g05378(.dina(w_asqrt32_25[1]),.dinb(w_n5274_0[0]),.dout(n5626),.clk(gclk));
	jand g05379(.dina(w_n5626_0[1]),.dinb(n5625),.dout(n5627),.clk(gclk));
	jor g05380(.dina(n5627),.dinb(n5624),.dout(n5628),.clk(gclk));
	jnot g05381(.din(w_n5281_0[0]),.dout(n5629),.clk(gclk));
	jand g05382(.dina(w_n5626_0[0]),.dinb(n5629),.dout(n5630),.clk(gclk));
	jnot g05383(.din(n5630),.dout(n5631),.clk(gclk));
	jand g05384(.dina(n5631),.dinb(n5628),.dout(n5632),.clk(gclk));
	jand g05385(.dina(w_n5632_0[1]),.dinb(w_n5623_0[1]),.dout(n5633),.clk(gclk));
	jor g05386(.dina(n5633),.dinb(w_n5621_0[1]),.dout(n5634),.clk(gclk));
	jand g05387(.dina(w_n5634_0[1]),.dinb(w_asqrt51_19[0]),.dout(n5635),.clk(gclk));
	jxor g05388(.dina(w_n5282_0[0]),.dinb(w_n1312_23[1]),.dout(n5636),.clk(gclk));
	jand g05389(.dina(n5636),.dinb(w_asqrt32_25[0]),.dout(n5637),.clk(gclk));
	jxor g05390(.dina(n5637),.dinb(w_n5292_0[0]),.dout(n5638),.clk(gclk));
	jnot g05391(.din(n5638),.dout(n5639),.clk(gclk));
	jor g05392(.dina(w_n5634_0[0]),.dinb(w_asqrt51_18[2]),.dout(n5640),.clk(gclk));
	jand g05393(.dina(w_n5640_0[1]),.dinb(w_n5639_0[1]),.dout(n5641),.clk(gclk));
	jor g05394(.dina(w_n5641_0[2]),.dinb(w_n5635_0[2]),.dout(n5642),.clk(gclk));
	jand g05395(.dina(n5642),.dinb(w_asqrt52_20[2]),.dout(n5643),.clk(gclk));
	jnot g05396(.din(w_n5297_0[0]),.dout(n5644),.clk(gclk));
	jand g05397(.dina(n5644),.dinb(w_n5295_0[0]),.dout(n5645),.clk(gclk));
	jand g05398(.dina(n5645),.dinb(w_asqrt32_24[2]),.dout(n5646),.clk(gclk));
	jxor g05399(.dina(n5646),.dinb(w_n5305_0[0]),.dout(n5647),.clk(gclk));
	jnot g05400(.din(n5647),.dout(n5648),.clk(gclk));
	jor g05401(.dina(w_n5635_0[1]),.dinb(w_asqrt52_20[1]),.dout(n5649),.clk(gclk));
	jor g05402(.dina(n5649),.dinb(w_n5641_0[1]),.dout(n5650),.clk(gclk));
	jand g05403(.dina(w_n5650_0[1]),.dinb(w_n5648_0[1]),.dout(n5651),.clk(gclk));
	jor g05404(.dina(w_n5651_0[1]),.dinb(w_n5643_0[1]),.dout(n5652),.clk(gclk));
	jand g05405(.dina(w_n5652_0[2]),.dinb(w_asqrt53_19[1]),.dout(n5653),.clk(gclk));
	jor g05406(.dina(w_n5652_0[1]),.dinb(w_asqrt53_19[0]),.dout(n5654),.clk(gclk));
	jnot g05407(.din(w_n5311_0[0]),.dout(n5655),.clk(gclk));
	jnot g05408(.din(w_n5312_0[0]),.dout(n5656),.clk(gclk));
	jand g05409(.dina(w_asqrt32_24[1]),.dinb(w_n5308_0[0]),.dout(n5657),.clk(gclk));
	jand g05410(.dina(w_n5657_0[1]),.dinb(n5656),.dout(n5658),.clk(gclk));
	jor g05411(.dina(n5658),.dinb(n5655),.dout(n5659),.clk(gclk));
	jnot g05412(.din(w_n5313_0[0]),.dout(n5660),.clk(gclk));
	jand g05413(.dina(w_n5657_0[0]),.dinb(n5660),.dout(n5661),.clk(gclk));
	jnot g05414(.din(n5661),.dout(n5662),.clk(gclk));
	jand g05415(.dina(n5662),.dinb(n5659),.dout(n5663),.clk(gclk));
	jand g05416(.dina(w_n5663_0[1]),.dinb(n5654),.dout(n5664),.clk(gclk));
	jor g05417(.dina(w_n5664_0[1]),.dinb(w_n5653_0[1]),.dout(n5665),.clk(gclk));
	jand g05418(.dina(n5665),.dinb(w_asqrt54_20[2]),.dout(n5666),.clk(gclk));
	jor g05419(.dina(w_n5653_0[0]),.dinb(w_asqrt54_20[1]),.dout(n5667),.clk(gclk));
	jor g05420(.dina(n5667),.dinb(w_n5664_0[0]),.dout(n5668),.clk(gclk));
	jnot g05421(.din(w_n5319_0[0]),.dout(n5669),.clk(gclk));
	jnot g05422(.din(w_n5321_0[0]),.dout(n5670),.clk(gclk));
	jand g05423(.dina(w_asqrt32_24[0]),.dinb(w_n5315_0[0]),.dout(n5671),.clk(gclk));
	jand g05424(.dina(w_n5671_0[1]),.dinb(n5670),.dout(n5672),.clk(gclk));
	jor g05425(.dina(n5672),.dinb(n5669),.dout(n5673),.clk(gclk));
	jnot g05426(.din(w_n5322_0[0]),.dout(n5674),.clk(gclk));
	jand g05427(.dina(w_n5671_0[0]),.dinb(n5674),.dout(n5675),.clk(gclk));
	jnot g05428(.din(n5675),.dout(n5676),.clk(gclk));
	jand g05429(.dina(n5676),.dinb(n5673),.dout(n5677),.clk(gclk));
	jand g05430(.dina(w_n5677_0[1]),.dinb(w_n5668_0[1]),.dout(n5678),.clk(gclk));
	jor g05431(.dina(n5678),.dinb(w_n5666_0[1]),.dout(n5679),.clk(gclk));
	jand g05432(.dina(w_n5679_0[1]),.dinb(w_asqrt55_19[2]),.dout(n5680),.clk(gclk));
	jxor g05433(.dina(w_n5323_0[0]),.dinb(w_n791_24[1]),.dout(n5681),.clk(gclk));
	jand g05434(.dina(n5681),.dinb(w_asqrt32_23[2]),.dout(n5682),.clk(gclk));
	jxor g05435(.dina(n5682),.dinb(w_n5333_0[0]),.dout(n5683),.clk(gclk));
	jnot g05436(.din(n5683),.dout(n5684),.clk(gclk));
	jor g05437(.dina(w_n5679_0[0]),.dinb(w_asqrt55_19[1]),.dout(n5685),.clk(gclk));
	jand g05438(.dina(w_n5685_0[1]),.dinb(w_n5684_0[1]),.dout(n5686),.clk(gclk));
	jor g05439(.dina(w_n5686_0[2]),.dinb(w_n5680_0[2]),.dout(n5687),.clk(gclk));
	jand g05440(.dina(n5687),.dinb(w_asqrt56_20[2]),.dout(n5688),.clk(gclk));
	jnot g05441(.din(w_n5338_0[0]),.dout(n5689),.clk(gclk));
	jand g05442(.dina(n5689),.dinb(w_n5336_0[0]),.dout(n5690),.clk(gclk));
	jand g05443(.dina(n5690),.dinb(w_asqrt32_23[1]),.dout(n5691),.clk(gclk));
	jxor g05444(.dina(n5691),.dinb(w_n5346_0[0]),.dout(n5692),.clk(gclk));
	jnot g05445(.din(n5692),.dout(n5693),.clk(gclk));
	jor g05446(.dina(w_n5680_0[1]),.dinb(w_asqrt56_20[1]),.dout(n5694),.clk(gclk));
	jor g05447(.dina(n5694),.dinb(w_n5686_0[1]),.dout(n5695),.clk(gclk));
	jand g05448(.dina(w_n5695_0[1]),.dinb(w_n5693_0[1]),.dout(n5696),.clk(gclk));
	jor g05449(.dina(w_n5696_0[1]),.dinb(w_n5688_0[1]),.dout(n5697),.clk(gclk));
	jand g05450(.dina(w_n5697_0[2]),.dinb(w_asqrt57_20[0]),.dout(n5698),.clk(gclk));
	jor g05451(.dina(w_n5697_0[1]),.dinb(w_asqrt57_19[2]),.dout(n5699),.clk(gclk));
	jnot g05452(.din(w_n5352_0[0]),.dout(n5700),.clk(gclk));
	jnot g05453(.din(w_n5353_0[0]),.dout(n5701),.clk(gclk));
	jand g05454(.dina(w_asqrt32_23[0]),.dinb(w_n5349_0[0]),.dout(n5702),.clk(gclk));
	jand g05455(.dina(w_n5702_0[1]),.dinb(n5701),.dout(n5703),.clk(gclk));
	jor g05456(.dina(n5703),.dinb(n5700),.dout(n5704),.clk(gclk));
	jnot g05457(.din(w_n5354_0[0]),.dout(n5705),.clk(gclk));
	jand g05458(.dina(w_n5702_0[0]),.dinb(n5705),.dout(n5706),.clk(gclk));
	jnot g05459(.din(n5706),.dout(n5707),.clk(gclk));
	jand g05460(.dina(n5707),.dinb(n5704),.dout(n5708),.clk(gclk));
	jand g05461(.dina(w_n5708_0[1]),.dinb(n5699),.dout(n5709),.clk(gclk));
	jor g05462(.dina(w_n5709_0[1]),.dinb(w_n5698_0[1]),.dout(n5710),.clk(gclk));
	jand g05463(.dina(n5710),.dinb(w_asqrt58_20[2]),.dout(n5711),.clk(gclk));
	jor g05464(.dina(w_n5698_0[0]),.dinb(w_asqrt58_20[1]),.dout(n5712),.clk(gclk));
	jor g05465(.dina(n5712),.dinb(w_n5709_0[0]),.dout(n5713),.clk(gclk));
	jnot g05466(.din(w_n5360_0[0]),.dout(n5714),.clk(gclk));
	jnot g05467(.din(w_n5362_0[0]),.dout(n5715),.clk(gclk));
	jand g05468(.dina(w_asqrt32_22[2]),.dinb(w_n5356_0[0]),.dout(n5716),.clk(gclk));
	jand g05469(.dina(w_n5716_0[1]),.dinb(n5715),.dout(n5717),.clk(gclk));
	jor g05470(.dina(n5717),.dinb(n5714),.dout(n5718),.clk(gclk));
	jnot g05471(.din(w_n5363_0[0]),.dout(n5719),.clk(gclk));
	jand g05472(.dina(w_n5716_0[0]),.dinb(n5719),.dout(n5720),.clk(gclk));
	jnot g05473(.din(n5720),.dout(n5721),.clk(gclk));
	jand g05474(.dina(n5721),.dinb(n5718),.dout(n5722),.clk(gclk));
	jand g05475(.dina(w_n5722_0[1]),.dinb(w_n5713_0[1]),.dout(n5723),.clk(gclk));
	jor g05476(.dina(n5723),.dinb(w_n5711_0[1]),.dout(n5724),.clk(gclk));
	jand g05477(.dina(w_n5724_0[1]),.dinb(w_asqrt59_20[1]),.dout(n5725),.clk(gclk));
	jxor g05478(.dina(w_n5364_0[0]),.dinb(w_n425_25[0]),.dout(n5726),.clk(gclk));
	jand g05479(.dina(n5726),.dinb(w_asqrt32_22[1]),.dout(n5727),.clk(gclk));
	jxor g05480(.dina(n5727),.dinb(w_n5374_0[0]),.dout(n5728),.clk(gclk));
	jnot g05481(.din(n5728),.dout(n5729),.clk(gclk));
	jor g05482(.dina(w_n5724_0[0]),.dinb(w_asqrt59_20[0]),.dout(n5730),.clk(gclk));
	jand g05483(.dina(w_n5730_0[1]),.dinb(w_n5729_0[1]),.dout(n5731),.clk(gclk));
	jor g05484(.dina(w_n5731_0[2]),.dinb(w_n5725_0[2]),.dout(n5732),.clk(gclk));
	jand g05485(.dina(n5732),.dinb(w_asqrt60_20[1]),.dout(n5733),.clk(gclk));
	jnot g05486(.din(w_n5379_0[0]),.dout(n5734),.clk(gclk));
	jand g05487(.dina(n5734),.dinb(w_n5377_0[0]),.dout(n5735),.clk(gclk));
	jand g05488(.dina(n5735),.dinb(w_asqrt32_22[0]),.dout(n5736),.clk(gclk));
	jxor g05489(.dina(n5736),.dinb(w_n5387_0[0]),.dout(n5737),.clk(gclk));
	jnot g05490(.din(n5737),.dout(n5738),.clk(gclk));
	jor g05491(.dina(w_n5725_0[1]),.dinb(w_asqrt60_20[0]),.dout(n5739),.clk(gclk));
	jor g05492(.dina(n5739),.dinb(w_n5731_0[1]),.dout(n5740),.clk(gclk));
	jand g05493(.dina(w_n5740_0[1]),.dinb(w_n5738_0[1]),.dout(n5741),.clk(gclk));
	jor g05494(.dina(w_n5741_0[1]),.dinb(w_n5733_0[1]),.dout(n5742),.clk(gclk));
	jand g05495(.dina(w_n5742_0[2]),.dinb(w_asqrt61_20[2]),.dout(n5743),.clk(gclk));
	jor g05496(.dina(w_n5742_0[1]),.dinb(w_asqrt61_20[1]),.dout(n5744),.clk(gclk));
	jnot g05497(.din(w_n5393_0[0]),.dout(n5745),.clk(gclk));
	jnot g05498(.din(w_n5394_0[0]),.dout(n5746),.clk(gclk));
	jand g05499(.dina(w_asqrt32_21[2]),.dinb(w_n5390_0[0]),.dout(n5747),.clk(gclk));
	jand g05500(.dina(w_n5747_0[1]),.dinb(n5746),.dout(n5748),.clk(gclk));
	jor g05501(.dina(n5748),.dinb(n5745),.dout(n5749),.clk(gclk));
	jnot g05502(.din(w_n5395_0[0]),.dout(n5750),.clk(gclk));
	jand g05503(.dina(w_n5747_0[0]),.dinb(n5750),.dout(n5751),.clk(gclk));
	jnot g05504(.din(n5751),.dout(n5752),.clk(gclk));
	jand g05505(.dina(n5752),.dinb(n5749),.dout(n5753),.clk(gclk));
	jand g05506(.dina(w_n5753_0[1]),.dinb(n5744),.dout(n5754),.clk(gclk));
	jor g05507(.dina(w_n5754_0[1]),.dinb(w_n5743_0[1]),.dout(n5755),.clk(gclk));
	jand g05508(.dina(n5755),.dinb(w_asqrt62_20[2]),.dout(n5756),.clk(gclk));
	jor g05509(.dina(w_n5743_0[0]),.dinb(w_asqrt62_20[1]),.dout(n5757),.clk(gclk));
	jor g05510(.dina(n5757),.dinb(w_n5754_0[0]),.dout(n5758),.clk(gclk));
	jnot g05511(.din(w_n5401_0[0]),.dout(n5759),.clk(gclk));
	jnot g05512(.din(w_n5403_0[0]),.dout(n5760),.clk(gclk));
	jand g05513(.dina(w_asqrt32_21[1]),.dinb(w_n5397_0[0]),.dout(n5761),.clk(gclk));
	jand g05514(.dina(w_n5761_0[1]),.dinb(n5760),.dout(n5762),.clk(gclk));
	jor g05515(.dina(n5762),.dinb(n5759),.dout(n5763),.clk(gclk));
	jnot g05516(.din(w_n5404_0[0]),.dout(n5764),.clk(gclk));
	jand g05517(.dina(w_n5761_0[0]),.dinb(n5764),.dout(n5765),.clk(gclk));
	jnot g05518(.din(n5765),.dout(n5766),.clk(gclk));
	jand g05519(.dina(n5766),.dinb(n5763),.dout(n5767),.clk(gclk));
	jand g05520(.dina(w_n5767_0[1]),.dinb(w_n5758_0[1]),.dout(n5768),.clk(gclk));
	jor g05521(.dina(n5768),.dinb(w_n5756_0[1]),.dout(n5769),.clk(gclk));
	jxor g05522(.dina(w_n5405_0[0]),.dinb(w_n199_30[2]),.dout(n5770),.clk(gclk));
	jand g05523(.dina(n5770),.dinb(w_asqrt32_21[0]),.dout(n5771),.clk(gclk));
	jxor g05524(.dina(n5771),.dinb(w_n5415_0[0]),.dout(n5772),.clk(gclk));
	jnot g05525(.din(w_n5417_0[0]),.dout(n5773),.clk(gclk));
	jand g05526(.dina(w_asqrt32_20[2]),.dinb(w_n5424_0[1]),.dout(n5774),.clk(gclk));
	jand g05527(.dina(w_n5774_0[1]),.dinb(w_n5773_0[2]),.dout(n5775),.clk(gclk));
	jor g05528(.dina(n5775),.dinb(w_n5432_0[0]),.dout(n5776),.clk(gclk));
	jor g05529(.dina(n5776),.dinb(w_n5772_0[1]),.dout(n5777),.clk(gclk));
	jnot g05530(.din(n5777),.dout(n5778),.clk(gclk));
	jand g05531(.dina(n5778),.dinb(w_n5769_1[2]),.dout(n5779),.clk(gclk));
	jor g05532(.dina(n5779),.dinb(w_asqrt63_11[0]),.dout(n5780),.clk(gclk));
	jnot g05533(.din(w_n5772_0[0]),.dout(n5781),.clk(gclk));
	jor g05534(.dina(w_n5781_0[2]),.dinb(w_n5769_1[1]),.dout(n5782),.clk(gclk));
	jor g05535(.dina(w_n5774_0[0]),.dinb(w_n5773_0[1]),.dout(n5783),.clk(gclk));
	jand g05536(.dina(w_n5424_0[0]),.dinb(w_n5773_0[0]),.dout(n5784),.clk(gclk));
	jor g05537(.dina(n5784),.dinb(w_n194_29[2]),.dout(n5785),.clk(gclk));
	jnot g05538(.din(n5785),.dout(n5786),.clk(gclk));
	jand g05539(.dina(n5786),.dinb(n5783),.dout(n5787),.clk(gclk));
	jnot g05540(.din(w_asqrt32_20[1]),.dout(n5788),.clk(gclk));
	jnot g05541(.din(w_n5787_0[1]),.dout(n5791),.clk(gclk));
	jand g05542(.dina(n5791),.dinb(w_n5782_0[1]),.dout(n5792),.clk(gclk));
	jand g05543(.dina(n5792),.dinb(w_n5780_0[1]),.dout(n5793),.clk(gclk));
	jor g05544(.dina(w_n5793_29[2]),.dinb(w_a62_0[0]),.dout(n5794),.clk(gclk));
	jxor g05545(.dina(w_n5794_0[1]),.dinb(w_n200_0[0]),.dout(n5795),.clk(gclk));
	jor g05546(.dina(w_n5793_29[1]),.dinb(w_n5443_1[0]),.dout(n5796),.clk(gclk));
	jnot g05547(.din(w_a60_0[1]),.dout(n5797),.clk(gclk));
	jnot g05548(.din(a[61]),.dout(n5798),.clk(gclk));
	jand g05549(.dina(w_n5443_0[2]),.dinb(w_n5798_0[2]),.dout(n5799),.clk(gclk));
	jand g05550(.dina(n5799),.dinb(w_n5797_1[1]),.dout(n5800),.clk(gclk));
	jnot g05551(.din(n5800),.dout(n5801),.clk(gclk));
	jand g05552(.dina(n5801),.dinb(n5796),.dout(n5802),.clk(gclk));
	jor g05553(.dina(w_n5802_0[2]),.dinb(w_n5788_20[2]),.dout(n5803),.clk(gclk));
	jand g05554(.dina(w_n5802_0[1]),.dinb(w_n5788_20[1]),.dout(n5804),.clk(gclk));
	jor g05555(.dina(n5804),.dinb(w_n5795_0[1]),.dout(n5805),.clk(gclk));
	jand g05556(.dina(w_n5805_0[1]),.dinb(w_n5803_0[1]),.dout(n5806),.clk(gclk));
	jor g05557(.dina(n5806),.dinb(w_n5121_23[1]),.dout(n5807),.clk(gclk));
	jor g05558(.dina(w_n5794_0[0]),.dinb(w_a63_0[0]),.dout(n5808),.clk(gclk));
	jnot g05559(.din(w_n5780_0[0]),.dout(n5809),.clk(gclk));
	jnot g05560(.din(w_n5782_0[0]),.dout(n5810),.clk(gclk));
	jor g05561(.dina(w_n5787_0[0]),.dinb(w_n5788_20[0]),.dout(n5811),.clk(gclk));
	jor g05562(.dina(n5811),.dinb(w_n5810_0[1]),.dout(n5812),.clk(gclk));
	jor g05563(.dina(n5812),.dinb(n5809),.dout(n5813),.clk(gclk));
	jand g05564(.dina(n5813),.dinb(n5808),.dout(n5814),.clk(gclk));
	jxor g05565(.dina(n5814),.dinb(w_n5124_0[1]),.dout(n5815),.clk(gclk));
	jand g05566(.dina(w_n5803_0[0]),.dinb(w_n5121_23[0]),.dout(n5816),.clk(gclk));
	jand g05567(.dina(n5816),.dinb(w_n5805_0[0]),.dout(n5817),.clk(gclk));
	jor g05568(.dina(w_n5817_0[1]),.dinb(w_n5815_0[1]),.dout(n5818),.clk(gclk));
	jand g05569(.dina(w_n5818_0[1]),.dinb(w_n5807_0[1]),.dout(n5819),.clk(gclk));
	jor g05570(.dina(w_n5819_0[2]),.dinb(w_n5116_20[1]),.dout(n5820),.clk(gclk));
	jand g05571(.dina(w_n5819_0[1]),.dinb(w_n5116_20[0]),.dout(n5821),.clk(gclk));
	jxor g05572(.dina(w_n5446_0[0]),.dinb(w_n5121_22[2]),.dout(n5822),.clk(gclk));
	jor g05573(.dina(n5822),.dinb(w_n5793_29[0]),.dout(n5823),.clk(gclk));
	jxor g05574(.dina(n5823),.dinb(w_n5449_0[0]),.dout(n5824),.clk(gclk));
	jor g05575(.dina(w_n5824_0[1]),.dinb(n5821),.dout(n5825),.clk(gclk));
	jand g05576(.dina(w_n5825_0[1]),.dinb(w_n5820_0[1]),.dout(n5826),.clk(gclk));
	jor g05577(.dina(n5826),.dinb(w_n4499_24[0]),.dout(n5827),.clk(gclk));
	jnot g05578(.din(w_n5455_0[0]),.dout(n5828),.clk(gclk));
	jor g05579(.dina(n5828),.dinb(w_n5453_0[0]),.dout(n5829),.clk(gclk));
	jor g05580(.dina(n5829),.dinb(w_n5793_28[2]),.dout(n5830),.clk(gclk));
	jxor g05581(.dina(n5830),.dinb(w_n5464_0[0]),.dout(n5831),.clk(gclk));
	jand g05582(.dina(w_n5820_0[0]),.dinb(w_n4499_23[2]),.dout(n5832),.clk(gclk));
	jand g05583(.dina(n5832),.dinb(w_n5825_0[0]),.dout(n5833),.clk(gclk));
	jor g05584(.dina(w_n5833_0[1]),.dinb(w_n5831_0[1]),.dout(n5834),.clk(gclk));
	jand g05585(.dina(w_n5834_0[1]),.dinb(w_n5827_0[1]),.dout(n5835),.clk(gclk));
	jor g05586(.dina(w_n5835_0[2]),.dinb(w_n4494_21[0]),.dout(n5836),.clk(gclk));
	jand g05587(.dina(w_n5835_0[1]),.dinb(w_n4494_20[2]),.dout(n5837),.clk(gclk));
	jxor g05588(.dina(w_n5466_0[0]),.dinb(w_n4499_23[1]),.dout(n5838),.clk(gclk));
	jor g05589(.dina(n5838),.dinb(w_n5793_28[1]),.dout(n5839),.clk(gclk));
	jxor g05590(.dina(n5839),.dinb(w_n5471_0[0]),.dout(n5840),.clk(gclk));
	jnot g05591(.din(w_n5840_0[1]),.dout(n5841),.clk(gclk));
	jor g05592(.dina(n5841),.dinb(n5837),.dout(n5842),.clk(gclk));
	jand g05593(.dina(w_n5842_0[1]),.dinb(w_n5836_0[1]),.dout(n5843),.clk(gclk));
	jor g05594(.dina(n5843),.dinb(w_n3912_24[0]),.dout(n5844),.clk(gclk));
	jand g05595(.dina(w_n5836_0[0]),.dinb(w_n3912_23[2]),.dout(n5845),.clk(gclk));
	jand g05596(.dina(n5845),.dinb(w_n5842_0[0]),.dout(n5846),.clk(gclk));
	jnot g05597(.din(w_n5475_0[0]),.dout(n5847),.clk(gclk));
	jnot g05598(.din(w_n5793_28[0]),.dout(asqrt_fa_32),.clk(gclk));
	jand g05599(.dina(w_asqrt31_21[1]),.dinb(n5847),.dout(n5849),.clk(gclk));
	jand g05600(.dina(w_n5849_0[1]),.dinb(w_n5482_0[0]),.dout(n5850),.clk(gclk));
	jor g05601(.dina(n5850),.dinb(w_n5480_0[0]),.dout(n5851),.clk(gclk));
	jand g05602(.dina(w_n5849_0[0]),.dinb(w_n5483_0[0]),.dout(n5852),.clk(gclk));
	jnot g05603(.din(n5852),.dout(n5853),.clk(gclk));
	jand g05604(.dina(n5853),.dinb(n5851),.dout(n5854),.clk(gclk));
	jnot g05605(.din(n5854),.dout(n5855),.clk(gclk));
	jor g05606(.dina(w_n5855_0[1]),.dinb(w_n5846_0[1]),.dout(n5856),.clk(gclk));
	jand g05607(.dina(n5856),.dinb(w_n5844_0[1]),.dout(n5857),.clk(gclk));
	jor g05608(.dina(w_n5857_0[2]),.dinb(w_n3907_21[0]),.dout(n5858),.clk(gclk));
	jand g05609(.dina(w_n5857_0[1]),.dinb(w_n3907_20[2]),.dout(n5859),.clk(gclk));
	jnot g05610(.din(w_n5490_0[0]),.dout(n5860),.clk(gclk));
	jxor g05611(.dina(w_n5484_0[0]),.dinb(w_n3912_23[1]),.dout(n5861),.clk(gclk));
	jor g05612(.dina(n5861),.dinb(w_n5793_27[2]),.dout(n5862),.clk(gclk));
	jxor g05613(.dina(n5862),.dinb(n5860),.dout(n5863),.clk(gclk));
	jnot g05614(.din(w_n5863_0[1]),.dout(n5864),.clk(gclk));
	jor g05615(.dina(n5864),.dinb(n5859),.dout(n5865),.clk(gclk));
	jand g05616(.dina(w_n5865_0[1]),.dinb(w_n5858_0[1]),.dout(n5866),.clk(gclk));
	jor g05617(.dina(n5866),.dinb(w_n3376_24[2]),.dout(n5867),.clk(gclk));
	jnot g05618(.din(w_n5495_0[0]),.dout(n5868),.clk(gclk));
	jor g05619(.dina(n5868),.dinb(w_n5493_0[0]),.dout(n5869),.clk(gclk));
	jor g05620(.dina(n5869),.dinb(w_n5793_27[1]),.dout(n5870),.clk(gclk));
	jxor g05621(.dina(n5870),.dinb(w_n5504_0[0]),.dout(n5871),.clk(gclk));
	jand g05622(.dina(w_n5858_0[0]),.dinb(w_n3376_24[1]),.dout(n5872),.clk(gclk));
	jand g05623(.dina(n5872),.dinb(w_n5865_0[0]),.dout(n5873),.clk(gclk));
	jor g05624(.dina(w_n5873_0[1]),.dinb(w_n5871_0[1]),.dout(n5874),.clk(gclk));
	jand g05625(.dina(w_n5874_0[1]),.dinb(w_n5867_0[1]),.dout(n5875),.clk(gclk));
	jor g05626(.dina(w_n5875_0[2]),.dinb(w_n3371_21[1]),.dout(n5876),.clk(gclk));
	jand g05627(.dina(w_n5875_0[1]),.dinb(w_n3371_21[0]),.dout(n5877),.clk(gclk));
	jnot g05628(.din(w_n5511_0[0]),.dout(n5878),.clk(gclk));
	jxor g05629(.dina(w_n5506_0[0]),.dinb(w_n3376_24[0]),.dout(n5879),.clk(gclk));
	jor g05630(.dina(n5879),.dinb(w_n5793_27[0]),.dout(n5880),.clk(gclk));
	jxor g05631(.dina(n5880),.dinb(n5878),.dout(n5881),.clk(gclk));
	jnot g05632(.din(n5881),.dout(n5882),.clk(gclk));
	jor g05633(.dina(w_n5882_0[1]),.dinb(n5877),.dout(n5883),.clk(gclk));
	jand g05634(.dina(w_n5883_0[1]),.dinb(w_n5876_0[1]),.dout(n5884),.clk(gclk));
	jor g05635(.dina(n5884),.dinb(w_n2875_24[1]),.dout(n5885),.clk(gclk));
	jand g05636(.dina(w_n5876_0[0]),.dinb(w_n2875_24[0]),.dout(n5886),.clk(gclk));
	jand g05637(.dina(n5886),.dinb(w_n5883_0[0]),.dout(n5887),.clk(gclk));
	jnot g05638(.din(w_n5514_0[0]),.dout(n5888),.clk(gclk));
	jand g05639(.dina(w_asqrt31_21[0]),.dinb(n5888),.dout(n5889),.clk(gclk));
	jand g05640(.dina(w_n5889_0[1]),.dinb(w_n5521_0[0]),.dout(n5890),.clk(gclk));
	jor g05641(.dina(n5890),.dinb(w_n5519_0[0]),.dout(n5891),.clk(gclk));
	jand g05642(.dina(w_n5889_0[0]),.dinb(w_n5522_0[0]),.dout(n5892),.clk(gclk));
	jnot g05643(.din(n5892),.dout(n5893),.clk(gclk));
	jand g05644(.dina(n5893),.dinb(n5891),.dout(n5894),.clk(gclk));
	jnot g05645(.din(n5894),.dout(n5895),.clk(gclk));
	jor g05646(.dina(w_n5895_0[1]),.dinb(w_n5887_0[1]),.dout(n5896),.clk(gclk));
	jand g05647(.dina(n5896),.dinb(w_n5885_0[1]),.dout(n5897),.clk(gclk));
	jor g05648(.dina(w_n5897_0[1]),.dinb(w_n2870_21[1]),.dout(n5898),.clk(gclk));
	jxor g05649(.dina(w_n5523_0[0]),.dinb(w_n2875_23[2]),.dout(n5899),.clk(gclk));
	jor g05650(.dina(n5899),.dinb(w_n5793_26[2]),.dout(n5900),.clk(gclk));
	jxor g05651(.dina(n5900),.dinb(w_n5528_0[0]),.dout(n5901),.clk(gclk));
	jand g05652(.dina(w_n5897_0[0]),.dinb(w_n2870_21[0]),.dout(n5902),.clk(gclk));
	jor g05653(.dina(w_n5902_0[1]),.dinb(w_n5901_0[1]),.dout(n5903),.clk(gclk));
	jand g05654(.dina(w_n5903_0[2]),.dinb(w_n5898_0[2]),.dout(n5904),.clk(gclk));
	jor g05655(.dina(n5904),.dinb(w_n2425_24[2]),.dout(n5905),.clk(gclk));
	jnot g05656(.din(w_n5533_0[0]),.dout(n5906),.clk(gclk));
	jor g05657(.dina(n5906),.dinb(w_n5531_0[0]),.dout(n5907),.clk(gclk));
	jor g05658(.dina(n5907),.dinb(w_n5793_26[1]),.dout(n5908),.clk(gclk));
	jxor g05659(.dina(n5908),.dinb(w_n5542_0[0]),.dout(n5909),.clk(gclk));
	jand g05660(.dina(w_n5898_0[1]),.dinb(w_n2425_24[1]),.dout(n5910),.clk(gclk));
	jand g05661(.dina(n5910),.dinb(w_n5903_0[1]),.dout(n5911),.clk(gclk));
	jor g05662(.dina(w_n5911_0[1]),.dinb(w_n5909_0[1]),.dout(n5912),.clk(gclk));
	jand g05663(.dina(w_n5912_0[1]),.dinb(w_n5905_0[1]),.dout(n5913),.clk(gclk));
	jor g05664(.dina(w_n5913_0[2]),.dinb(w_n2420_22[1]),.dout(n5914),.clk(gclk));
	jand g05665(.dina(w_n5913_0[1]),.dinb(w_n2420_22[0]),.dout(n5915),.clk(gclk));
	jnot g05666(.din(w_n5545_0[0]),.dout(n5916),.clk(gclk));
	jand g05667(.dina(w_asqrt31_20[2]),.dinb(n5916),.dout(n5917),.clk(gclk));
	jand g05668(.dina(w_n5917_0[1]),.dinb(w_n5550_0[0]),.dout(n5918),.clk(gclk));
	jor g05669(.dina(n5918),.dinb(w_n5549_0[0]),.dout(n5919),.clk(gclk));
	jand g05670(.dina(w_n5917_0[0]),.dinb(w_n5551_0[0]),.dout(n5920),.clk(gclk));
	jnot g05671(.din(n5920),.dout(n5921),.clk(gclk));
	jand g05672(.dina(n5921),.dinb(n5919),.dout(n5922),.clk(gclk));
	jnot g05673(.din(n5922),.dout(n5923),.clk(gclk));
	jor g05674(.dina(w_n5923_0[1]),.dinb(n5915),.dout(n5924),.clk(gclk));
	jand g05675(.dina(w_n5924_0[1]),.dinb(w_n5914_0[1]),.dout(n5925),.clk(gclk));
	jor g05676(.dina(n5925),.dinb(w_n2010_24[2]),.dout(n5926),.clk(gclk));
	jand g05677(.dina(w_n5914_0[0]),.dinb(w_n2010_24[1]),.dout(n5927),.clk(gclk));
	jand g05678(.dina(n5927),.dinb(w_n5924_0[0]),.dout(n5928),.clk(gclk));
	jnot g05679(.din(w_n5553_0[0]),.dout(n5929),.clk(gclk));
	jand g05680(.dina(w_asqrt31_20[1]),.dinb(n5929),.dout(n5930),.clk(gclk));
	jand g05681(.dina(w_n5930_0[1]),.dinb(w_n5560_0[0]),.dout(n5931),.clk(gclk));
	jor g05682(.dina(n5931),.dinb(w_n5558_0[0]),.dout(n5932),.clk(gclk));
	jand g05683(.dina(w_n5930_0[0]),.dinb(w_n5561_0[0]),.dout(n5933),.clk(gclk));
	jnot g05684(.din(n5933),.dout(n5934),.clk(gclk));
	jand g05685(.dina(n5934),.dinb(n5932),.dout(n5935),.clk(gclk));
	jnot g05686(.din(n5935),.dout(n5936),.clk(gclk));
	jor g05687(.dina(w_n5936_0[1]),.dinb(w_n5928_0[1]),.dout(n5937),.clk(gclk));
	jand g05688(.dina(n5937),.dinb(w_n5926_0[1]),.dout(n5938),.clk(gclk));
	jor g05689(.dina(w_n5938_0[1]),.dinb(w_n2005_22[1]),.dout(n5939),.clk(gclk));
	jxor g05690(.dina(w_n5562_0[0]),.dinb(w_n2010_24[0]),.dout(n5940),.clk(gclk));
	jor g05691(.dina(n5940),.dinb(w_n5793_26[0]),.dout(n5941),.clk(gclk));
	jxor g05692(.dina(n5941),.dinb(w_n5573_0[0]),.dout(n5942),.clk(gclk));
	jand g05693(.dina(w_n5938_0[0]),.dinb(w_n2005_22[0]),.dout(n5943),.clk(gclk));
	jor g05694(.dina(w_n5943_0[1]),.dinb(w_n5942_0[1]),.dout(n5944),.clk(gclk));
	jand g05695(.dina(w_n5944_0[2]),.dinb(w_n5939_0[2]),.dout(n5945),.clk(gclk));
	jor g05696(.dina(n5945),.dinb(w_n1646_25[1]),.dout(n5946),.clk(gclk));
	jnot g05697(.din(w_n5578_0[0]),.dout(n5947),.clk(gclk));
	jor g05698(.dina(n5947),.dinb(w_n5576_0[0]),.dout(n5948),.clk(gclk));
	jor g05699(.dina(n5948),.dinb(w_n5793_25[2]),.dout(n5949),.clk(gclk));
	jxor g05700(.dina(n5949),.dinb(w_n5587_0[0]),.dout(n5950),.clk(gclk));
	jand g05701(.dina(w_n5939_0[1]),.dinb(w_n1646_25[0]),.dout(n5951),.clk(gclk));
	jand g05702(.dina(n5951),.dinb(w_n5944_0[1]),.dout(n5952),.clk(gclk));
	jor g05703(.dina(w_n5952_0[1]),.dinb(w_n5950_0[1]),.dout(n5953),.clk(gclk));
	jand g05704(.dina(w_n5953_0[1]),.dinb(w_n5946_0[1]),.dout(n5954),.clk(gclk));
	jor g05705(.dina(w_n5954_0[2]),.dinb(w_n1641_23[0]),.dout(n5955),.clk(gclk));
	jand g05706(.dina(w_n5954_0[1]),.dinb(w_n1641_22[2]),.dout(n5956),.clk(gclk));
	jnot g05707(.din(w_n5590_0[0]),.dout(n5957),.clk(gclk));
	jand g05708(.dina(w_asqrt31_20[0]),.dinb(n5957),.dout(n5958),.clk(gclk));
	jand g05709(.dina(w_n5958_0[1]),.dinb(w_n5595_0[0]),.dout(n5959),.clk(gclk));
	jor g05710(.dina(n5959),.dinb(w_n5594_0[0]),.dout(n5960),.clk(gclk));
	jand g05711(.dina(w_n5958_0[0]),.dinb(w_n5596_0[0]),.dout(n5961),.clk(gclk));
	jnot g05712(.din(n5961),.dout(n5962),.clk(gclk));
	jand g05713(.dina(n5962),.dinb(n5960),.dout(n5963),.clk(gclk));
	jnot g05714(.din(n5963),.dout(n5964),.clk(gclk));
	jor g05715(.dina(w_n5964_0[1]),.dinb(n5956),.dout(n5965),.clk(gclk));
	jand g05716(.dina(w_n5965_0[1]),.dinb(w_n5955_0[1]),.dout(n5966),.clk(gclk));
	jor g05717(.dina(n5966),.dinb(w_n1317_25[1]),.dout(n5967),.clk(gclk));
	jand g05718(.dina(w_n5955_0[0]),.dinb(w_n1317_25[0]),.dout(n5968),.clk(gclk));
	jand g05719(.dina(n5968),.dinb(w_n5965_0[0]),.dout(n5969),.clk(gclk));
	jnot g05720(.din(w_n5598_0[0]),.dout(n5970),.clk(gclk));
	jand g05721(.dina(w_asqrt31_19[2]),.dinb(n5970),.dout(n5971),.clk(gclk));
	jand g05722(.dina(w_n5971_0[1]),.dinb(w_n5605_0[0]),.dout(n5972),.clk(gclk));
	jor g05723(.dina(n5972),.dinb(w_n5603_0[0]),.dout(n5973),.clk(gclk));
	jand g05724(.dina(w_n5971_0[0]),.dinb(w_n5606_0[0]),.dout(n5974),.clk(gclk));
	jnot g05725(.din(n5974),.dout(n5975),.clk(gclk));
	jand g05726(.dina(n5975),.dinb(n5973),.dout(n5976),.clk(gclk));
	jnot g05727(.din(n5976),.dout(n5977),.clk(gclk));
	jor g05728(.dina(w_n5977_0[1]),.dinb(w_n5969_0[1]),.dout(n5978),.clk(gclk));
	jand g05729(.dina(n5978),.dinb(w_n5967_0[1]),.dout(n5979),.clk(gclk));
	jor g05730(.dina(w_n5979_0[1]),.dinb(w_n1312_23[0]),.dout(n5980),.clk(gclk));
	jxor g05731(.dina(w_n5607_0[0]),.dinb(w_n1317_24[2]),.dout(n5981),.clk(gclk));
	jor g05732(.dina(n5981),.dinb(w_n5793_25[1]),.dout(n5982),.clk(gclk));
	jxor g05733(.dina(n5982),.dinb(w_n5618_0[0]),.dout(n5983),.clk(gclk));
	jand g05734(.dina(w_n5979_0[0]),.dinb(w_n1312_22[2]),.dout(n5984),.clk(gclk));
	jor g05735(.dina(w_n5984_0[1]),.dinb(w_n5983_0[1]),.dout(n5985),.clk(gclk));
	jand g05736(.dina(w_n5985_0[2]),.dinb(w_n5980_0[2]),.dout(n5986),.clk(gclk));
	jor g05737(.dina(n5986),.dinb(w_n1039_25[2]),.dout(n5987),.clk(gclk));
	jnot g05738(.din(w_n5623_0[0]),.dout(n5988),.clk(gclk));
	jor g05739(.dina(n5988),.dinb(w_n5621_0[0]),.dout(n5989),.clk(gclk));
	jor g05740(.dina(n5989),.dinb(w_n5793_25[0]),.dout(n5990),.clk(gclk));
	jxor g05741(.dina(n5990),.dinb(w_n5632_0[0]),.dout(n5991),.clk(gclk));
	jand g05742(.dina(w_n5980_0[1]),.dinb(w_n1039_25[1]),.dout(n5992),.clk(gclk));
	jand g05743(.dina(n5992),.dinb(w_n5985_0[1]),.dout(n5993),.clk(gclk));
	jor g05744(.dina(w_n5993_0[1]),.dinb(w_n5991_0[1]),.dout(n5994),.clk(gclk));
	jand g05745(.dina(w_n5994_0[1]),.dinb(w_n5987_0[1]),.dout(n5995),.clk(gclk));
	jor g05746(.dina(w_n5995_0[2]),.dinb(w_n1034_24[0]),.dout(n5996),.clk(gclk));
	jand g05747(.dina(w_n5995_0[1]),.dinb(w_n1034_23[2]),.dout(n5997),.clk(gclk));
	jnot g05748(.din(w_n5635_0[0]),.dout(n5998),.clk(gclk));
	jand g05749(.dina(w_asqrt31_19[1]),.dinb(n5998),.dout(n5999),.clk(gclk));
	jand g05750(.dina(w_n5999_0[1]),.dinb(w_n5640_0[0]),.dout(n6000),.clk(gclk));
	jor g05751(.dina(n6000),.dinb(w_n5639_0[0]),.dout(n6001),.clk(gclk));
	jand g05752(.dina(w_n5999_0[0]),.dinb(w_n5641_0[0]),.dout(n6002),.clk(gclk));
	jnot g05753(.din(n6002),.dout(n6003),.clk(gclk));
	jand g05754(.dina(n6003),.dinb(n6001),.dout(n6004),.clk(gclk));
	jnot g05755(.din(n6004),.dout(n6005),.clk(gclk));
	jor g05756(.dina(w_n6005_0[1]),.dinb(n5997),.dout(n6006),.clk(gclk));
	jand g05757(.dina(w_n6006_0[1]),.dinb(w_n5996_0[1]),.dout(n6007),.clk(gclk));
	jor g05758(.dina(n6007),.dinb(w_n796_25[2]),.dout(n6008),.clk(gclk));
	jand g05759(.dina(w_n5996_0[0]),.dinb(w_n796_25[1]),.dout(n6009),.clk(gclk));
	jand g05760(.dina(n6009),.dinb(w_n6006_0[0]),.dout(n6010),.clk(gclk));
	jnot g05761(.din(w_n5643_0[0]),.dout(n6011),.clk(gclk));
	jand g05762(.dina(w_asqrt31_19[0]),.dinb(n6011),.dout(n6012),.clk(gclk));
	jand g05763(.dina(w_n6012_0[1]),.dinb(w_n5650_0[0]),.dout(n6013),.clk(gclk));
	jor g05764(.dina(n6013),.dinb(w_n5648_0[0]),.dout(n6014),.clk(gclk));
	jand g05765(.dina(w_n6012_0[0]),.dinb(w_n5651_0[0]),.dout(n6015),.clk(gclk));
	jnot g05766(.din(n6015),.dout(n6016),.clk(gclk));
	jand g05767(.dina(n6016),.dinb(n6014),.dout(n6017),.clk(gclk));
	jnot g05768(.din(n6017),.dout(n6018),.clk(gclk));
	jor g05769(.dina(w_n6018_0[1]),.dinb(w_n6010_0[1]),.dout(n6019),.clk(gclk));
	jand g05770(.dina(n6019),.dinb(w_n6008_0[1]),.dout(n6020),.clk(gclk));
	jor g05771(.dina(w_n6020_0[1]),.dinb(w_n791_24[0]),.dout(n6021),.clk(gclk));
	jxor g05772(.dina(w_n5652_0[0]),.dinb(w_n796_25[0]),.dout(n6022),.clk(gclk));
	jor g05773(.dina(n6022),.dinb(w_n5793_24[2]),.dout(n6023),.clk(gclk));
	jxor g05774(.dina(n6023),.dinb(w_n5663_0[0]),.dout(n6024),.clk(gclk));
	jand g05775(.dina(w_n6020_0[0]),.dinb(w_n791_23[2]),.dout(n6025),.clk(gclk));
	jor g05776(.dina(w_n6025_0[1]),.dinb(w_n6024_0[1]),.dout(n6026),.clk(gclk));
	jand g05777(.dina(w_n6026_0[2]),.dinb(w_n6021_0[2]),.dout(n6027),.clk(gclk));
	jor g05778(.dina(n6027),.dinb(w_n595_26[0]),.dout(n6028),.clk(gclk));
	jnot g05779(.din(w_n5668_0[0]),.dout(n6029),.clk(gclk));
	jor g05780(.dina(n6029),.dinb(w_n5666_0[0]),.dout(n6030),.clk(gclk));
	jor g05781(.dina(n6030),.dinb(w_n5793_24[1]),.dout(n6031),.clk(gclk));
	jxor g05782(.dina(n6031),.dinb(w_n5677_0[0]),.dout(n6032),.clk(gclk));
	jand g05783(.dina(w_n6021_0[1]),.dinb(w_n595_25[2]),.dout(n6033),.clk(gclk));
	jand g05784(.dina(n6033),.dinb(w_n6026_0[1]),.dout(n6034),.clk(gclk));
	jor g05785(.dina(w_n6034_0[1]),.dinb(w_n6032_0[1]),.dout(n6035),.clk(gclk));
	jand g05786(.dina(w_n6035_0[1]),.dinb(w_n6028_0[1]),.dout(n6036),.clk(gclk));
	jor g05787(.dina(w_n6036_0[2]),.dinb(w_n590_24[2]),.dout(n6037),.clk(gclk));
	jand g05788(.dina(w_n6036_0[1]),.dinb(w_n590_24[1]),.dout(n6038),.clk(gclk));
	jnot g05789(.din(w_n5680_0[0]),.dout(n6039),.clk(gclk));
	jand g05790(.dina(w_asqrt31_18[2]),.dinb(n6039),.dout(n6040),.clk(gclk));
	jand g05791(.dina(w_n6040_0[1]),.dinb(w_n5685_0[0]),.dout(n6041),.clk(gclk));
	jor g05792(.dina(n6041),.dinb(w_n5684_0[0]),.dout(n6042),.clk(gclk));
	jand g05793(.dina(w_n6040_0[0]),.dinb(w_n5686_0[0]),.dout(n6043),.clk(gclk));
	jnot g05794(.din(n6043),.dout(n6044),.clk(gclk));
	jand g05795(.dina(n6044),.dinb(n6042),.dout(n6045),.clk(gclk));
	jnot g05796(.din(n6045),.dout(n6046),.clk(gclk));
	jor g05797(.dina(w_n6046_0[1]),.dinb(n6038),.dout(n6047),.clk(gclk));
	jand g05798(.dina(w_n6047_0[1]),.dinb(w_n6037_0[1]),.dout(n6048),.clk(gclk));
	jor g05799(.dina(n6048),.dinb(w_n430_26[0]),.dout(n6049),.clk(gclk));
	jand g05800(.dina(w_n6037_0[0]),.dinb(w_n430_25[2]),.dout(n6050),.clk(gclk));
	jand g05801(.dina(n6050),.dinb(w_n6047_0[0]),.dout(n6051),.clk(gclk));
	jnot g05802(.din(w_n5688_0[0]),.dout(n6052),.clk(gclk));
	jand g05803(.dina(w_asqrt31_18[1]),.dinb(n6052),.dout(n6053),.clk(gclk));
	jand g05804(.dina(w_n6053_0[1]),.dinb(w_n5695_0[0]),.dout(n6054),.clk(gclk));
	jor g05805(.dina(n6054),.dinb(w_n5693_0[0]),.dout(n6055),.clk(gclk));
	jand g05806(.dina(w_n6053_0[0]),.dinb(w_n5696_0[0]),.dout(n6056),.clk(gclk));
	jnot g05807(.din(n6056),.dout(n6057),.clk(gclk));
	jand g05808(.dina(n6057),.dinb(n6055),.dout(n6058),.clk(gclk));
	jnot g05809(.din(n6058),.dout(n6059),.clk(gclk));
	jor g05810(.dina(w_n6059_0[1]),.dinb(w_n6051_0[1]),.dout(n6060),.clk(gclk));
	jand g05811(.dina(n6060),.dinb(w_n6049_0[1]),.dout(n6061),.clk(gclk));
	jor g05812(.dina(w_n6061_0[1]),.dinb(w_n425_24[2]),.dout(n6062),.clk(gclk));
	jxor g05813(.dina(w_n5697_0[0]),.dinb(w_n430_25[1]),.dout(n6063),.clk(gclk));
	jor g05814(.dina(n6063),.dinb(w_n5793_24[0]),.dout(n6064),.clk(gclk));
	jxor g05815(.dina(n6064),.dinb(w_n5708_0[0]),.dout(n6065),.clk(gclk));
	jand g05816(.dina(w_n6061_0[0]),.dinb(w_n425_24[1]),.dout(n6066),.clk(gclk));
	jor g05817(.dina(w_n6066_0[1]),.dinb(w_n6065_0[1]),.dout(n6067),.clk(gclk));
	jand g05818(.dina(w_n6067_0[2]),.dinb(w_n6062_0[2]),.dout(n6068),.clk(gclk));
	jor g05819(.dina(n6068),.dinb(w_n305_26[1]),.dout(n6069),.clk(gclk));
	jnot g05820(.din(w_n5713_0[0]),.dout(n6070),.clk(gclk));
	jor g05821(.dina(n6070),.dinb(w_n5711_0[0]),.dout(n6071),.clk(gclk));
	jor g05822(.dina(n6071),.dinb(w_n5793_23[2]),.dout(n6072),.clk(gclk));
	jxor g05823(.dina(n6072),.dinb(w_n5722_0[0]),.dout(n6073),.clk(gclk));
	jand g05824(.dina(w_n6062_0[1]),.dinb(w_n305_26[0]),.dout(n6074),.clk(gclk));
	jand g05825(.dina(n6074),.dinb(w_n6067_0[1]),.dout(n6075),.clk(gclk));
	jor g05826(.dina(w_n6075_0[1]),.dinb(w_n6073_0[1]),.dout(n6076),.clk(gclk));
	jand g05827(.dina(w_n6076_0[1]),.dinb(w_n6069_0[1]),.dout(n6077),.clk(gclk));
	jor g05828(.dina(w_n6077_0[2]),.dinb(w_n290_26[0]),.dout(n6078),.clk(gclk));
	jand g05829(.dina(w_n6077_0[1]),.dinb(w_n290_25[2]),.dout(n6079),.clk(gclk));
	jnot g05830(.din(w_n5725_0[0]),.dout(n6080),.clk(gclk));
	jand g05831(.dina(w_asqrt31_18[0]),.dinb(n6080),.dout(n6081),.clk(gclk));
	jand g05832(.dina(w_n6081_0[1]),.dinb(w_n5730_0[0]),.dout(n6082),.clk(gclk));
	jor g05833(.dina(n6082),.dinb(w_n5729_0[0]),.dout(n6083),.clk(gclk));
	jand g05834(.dina(w_n6081_0[0]),.dinb(w_n5731_0[0]),.dout(n6084),.clk(gclk));
	jnot g05835(.din(n6084),.dout(n6085),.clk(gclk));
	jand g05836(.dina(n6085),.dinb(n6083),.dout(n6086),.clk(gclk));
	jnot g05837(.din(n6086),.dout(n6087),.clk(gclk));
	jor g05838(.dina(w_n6087_0[1]),.dinb(n6079),.dout(n6088),.clk(gclk));
	jand g05839(.dina(w_n6088_0[1]),.dinb(w_n6078_0[1]),.dout(n6089),.clk(gclk));
	jor g05840(.dina(n6089),.dinb(w_n223_26[1]),.dout(n6090),.clk(gclk));
	jand g05841(.dina(w_n6078_0[0]),.dinb(w_n223_26[0]),.dout(n6091),.clk(gclk));
	jand g05842(.dina(n6091),.dinb(w_n6088_0[0]),.dout(n6092),.clk(gclk));
	jnot g05843(.din(w_n5733_0[0]),.dout(n6093),.clk(gclk));
	jand g05844(.dina(w_asqrt31_17[2]),.dinb(n6093),.dout(n6094),.clk(gclk));
	jand g05845(.dina(w_n6094_0[1]),.dinb(w_n5740_0[0]),.dout(n6095),.clk(gclk));
	jor g05846(.dina(n6095),.dinb(w_n5738_0[0]),.dout(n6096),.clk(gclk));
	jand g05847(.dina(w_n6094_0[0]),.dinb(w_n5741_0[0]),.dout(n6097),.clk(gclk));
	jnot g05848(.din(n6097),.dout(n6098),.clk(gclk));
	jand g05849(.dina(n6098),.dinb(n6096),.dout(n6099),.clk(gclk));
	jnot g05850(.din(n6099),.dout(n6100),.clk(gclk));
	jor g05851(.dina(w_n6100_0[1]),.dinb(w_n6092_0[1]),.dout(n6101),.clk(gclk));
	jand g05852(.dina(n6101),.dinb(w_n6090_0[1]),.dout(n6102),.clk(gclk));
	jor g05853(.dina(w_n6102_0[2]),.dinb(w_n199_30[1]),.dout(n6103),.clk(gclk));
	jand g05854(.dina(w_n6102_0[1]),.dinb(w_n199_30[0]),.dout(n6104),.clk(gclk));
	jxor g05855(.dina(w_n5742_0[0]),.dinb(w_n223_25[2]),.dout(n6105),.clk(gclk));
	jor g05856(.dina(n6105),.dinb(w_n5793_23[1]),.dout(n6106),.clk(gclk));
	jxor g05857(.dina(n6106),.dinb(w_n5753_0[0]),.dout(n6107),.clk(gclk));
	jor g05858(.dina(w_n6107_0[1]),.dinb(n6104),.dout(n6108),.clk(gclk));
	jand g05859(.dina(n6108),.dinb(n6103),.dout(n6109),.clk(gclk));
	jnot g05860(.din(w_n5758_0[0]),.dout(n6110),.clk(gclk));
	jor g05861(.dina(n6110),.dinb(w_n5756_0[0]),.dout(n6111),.clk(gclk));
	jor g05862(.dina(n6111),.dinb(w_n5793_23[0]),.dout(n6112),.clk(gclk));
	jxor g05863(.dina(n6112),.dinb(w_n5767_0[0]),.dout(n6113),.clk(gclk));
	jand g05864(.dina(w_asqrt31_17[1]),.dinb(w_n5781_0[1]),.dout(n6114),.clk(gclk));
	jand g05865(.dina(w_n6114_0[1]),.dinb(w_n5769_1[0]),.dout(n6115),.clk(gclk));
	jor g05866(.dina(n6115),.dinb(w_n5810_0[0]),.dout(n6116),.clk(gclk));
	jor g05867(.dina(n6116),.dinb(w_n6113_0[2]),.dout(n6117),.clk(gclk));
	jor g05868(.dina(n6117),.dinb(w_n6109_0[2]),.dout(n6118),.clk(gclk));
	jand g05869(.dina(n6118),.dinb(w_n194_29[1]),.dout(n6119),.clk(gclk));
	jand g05870(.dina(w_n6113_0[1]),.dinb(w_n6109_0[1]),.dout(n6120),.clk(gclk));
	jor g05871(.dina(w_n6114_0[0]),.dinb(w_n5769_0[2]),.dout(n6121),.clk(gclk));
	jand g05872(.dina(w_n5781_0[0]),.dinb(w_n5769_0[1]),.dout(n6122),.clk(gclk));
	jor g05873(.dina(n6122),.dinb(w_n194_29[0]),.dout(n6123),.clk(gclk));
	jnot g05874(.din(n6123),.dout(n6124),.clk(gclk));
	jand g05875(.dina(n6124),.dinb(n6121),.dout(n6125),.clk(gclk));
	jor g05876(.dina(w_n6125_0[1]),.dinb(w_n6120_0[2]),.dout(n6128),.clk(gclk));
	jor g05877(.dina(n6128),.dinb(w_n6119_0[1]),.dout(asqrt_fa_31),.clk(gclk));
	jxor g05878(.dina(w_n5802_0[0]),.dinb(w_n5788_19[2]),.dout(n6130),.clk(gclk));
	jand g05879(.dina(n6130),.dinb(w_asqrt30_31),.dout(n6131),.clk(gclk));
	jxor g05880(.dina(n6131),.dinb(w_n5795_0[0]),.dout(n6132),.clk(gclk));
	jand g05881(.dina(w_asqrt30_30[2]),.dinb(w_a60_0[0]),.dout(n6133),.clk(gclk));
	jnot g05882(.din(w_a58_0[1]),.dout(n6134),.clk(gclk));
	jnot g05883(.din(w_a59_0[1]),.dout(n6135),.clk(gclk));
	jand g05884(.dina(w_n5797_1[0]),.dinb(w_n6135_0[1]),.dout(n6136),.clk(gclk));
	jand g05885(.dina(n6136),.dinb(w_n6134_1[1]),.dout(n6137),.clk(gclk));
	jor g05886(.dina(n6137),.dinb(n6133),.dout(n6138),.clk(gclk));
	jand g05887(.dina(w_n6138_0[2]),.dinb(w_asqrt31_17[0]),.dout(n6139),.clk(gclk));
	jand g05888(.dina(w_asqrt30_30[1]),.dinb(w_n5797_0[2]),.dout(n6140),.clk(gclk));
	jxor g05889(.dina(w_n6140_0[1]),.dinb(w_n5798_0[1]),.dout(n6141),.clk(gclk));
	jor g05890(.dina(w_n6138_0[1]),.dinb(w_asqrt31_16[2]),.dout(n6142),.clk(gclk));
	jand g05891(.dina(n6142),.dinb(w_n6141_0[1]),.dout(n6143),.clk(gclk));
	jor g05892(.dina(w_n6143_0[1]),.dinb(w_n6139_0[1]),.dout(n6144),.clk(gclk));
	jand g05893(.dina(n6144),.dinb(w_asqrt32_20[0]),.dout(n6145),.clk(gclk));
	jand g05894(.dina(w_n6140_0[0]),.dinb(w_n5798_0[0]),.dout(n6146),.clk(gclk));
	jnot g05895(.din(w_n6119_0[0]),.dout(n6147),.clk(gclk));
	jnot g05896(.din(w_n6120_0[1]),.dout(n6148),.clk(gclk));
	jnot g05897(.din(w_n6125_0[0]),.dout(n6149),.clk(gclk));
	jand g05898(.dina(n6149),.dinb(w_asqrt31_16[1]),.dout(n6150),.clk(gclk));
	jand g05899(.dina(n6150),.dinb(n6148),.dout(n6151),.clk(gclk));
	jand g05900(.dina(n6151),.dinb(n6147),.dout(n6152),.clk(gclk));
	jor g05901(.dina(n6152),.dinb(n6146),.dout(n6153),.clk(gclk));
	jxor g05902(.dina(n6153),.dinb(w_n5443_0[1]),.dout(n6154),.clk(gclk));
	jor g05903(.dina(w_n6139_0[0]),.dinb(w_asqrt32_19[2]),.dout(n6155),.clk(gclk));
	jor g05904(.dina(n6155),.dinb(w_n6143_0[0]),.dout(n6156),.clk(gclk));
	jand g05905(.dina(w_n6156_0[1]),.dinb(w_n6154_0[1]),.dout(n6157),.clk(gclk));
	jor g05906(.dina(w_n6157_0[1]),.dinb(w_n6145_0[1]),.dout(n6158),.clk(gclk));
	jand g05907(.dina(w_n6158_0[2]),.dinb(w_asqrt33_17[0]),.dout(n6159),.clk(gclk));
	jnot g05908(.din(w_n6132_0[1]),.dout(n6160),.clk(gclk));
	jor g05909(.dina(w_n6158_0[1]),.dinb(w_asqrt33_16[2]),.dout(n6161),.clk(gclk));
	jand g05910(.dina(n6161),.dinb(n6160),.dout(n6162),.clk(gclk));
	jor g05911(.dina(w_n6162_0[1]),.dinb(w_n6159_0[1]),.dout(n6163),.clk(gclk));
	jand g05912(.dina(n6163),.dinb(w_asqrt34_20[0]),.dout(n6164),.clk(gclk));
	jor g05913(.dina(w_n6159_0[0]),.dinb(w_asqrt34_19[2]),.dout(n6165),.clk(gclk));
	jor g05914(.dina(n6165),.dinb(w_n6162_0[0]),.dout(n6166),.clk(gclk));
	jnot g05915(.din(w_n5815_0[0]),.dout(n6167),.clk(gclk));
	jnot g05916(.din(w_n5817_0[0]),.dout(n6168),.clk(gclk));
	jand g05917(.dina(w_asqrt30_30[0]),.dinb(w_n5807_0[0]),.dout(n6169),.clk(gclk));
	jand g05918(.dina(w_n6169_0[1]),.dinb(n6168),.dout(n6170),.clk(gclk));
	jor g05919(.dina(n6170),.dinb(n6167),.dout(n6171),.clk(gclk));
	jnot g05920(.din(w_n5818_0[0]),.dout(n6172),.clk(gclk));
	jand g05921(.dina(w_n6169_0[0]),.dinb(n6172),.dout(n6173),.clk(gclk));
	jnot g05922(.din(n6173),.dout(n6174),.clk(gclk));
	jand g05923(.dina(n6174),.dinb(n6171),.dout(n6175),.clk(gclk));
	jand g05924(.dina(w_n6175_0[1]),.dinb(w_n6166_0[1]),.dout(n6176),.clk(gclk));
	jor g05925(.dina(n6176),.dinb(w_n6164_0[1]),.dout(n6177),.clk(gclk));
	jand g05926(.dina(w_n6177_0[2]),.dinb(w_asqrt35_17[0]),.dout(n6178),.clk(gclk));
	jor g05927(.dina(w_n6177_0[1]),.dinb(w_asqrt35_16[2]),.dout(n6179),.clk(gclk));
	jnot g05928(.din(w_n5824_0[0]),.dout(n6180),.clk(gclk));
	jxor g05929(.dina(w_n5819_0[0]),.dinb(w_n5116_19[2]),.dout(n6181),.clk(gclk));
	jand g05930(.dina(n6181),.dinb(w_asqrt30_29[2]),.dout(n6182),.clk(gclk));
	jxor g05931(.dina(n6182),.dinb(n6180),.dout(n6183),.clk(gclk));
	jand g05932(.dina(w_n6183_0[1]),.dinb(n6179),.dout(n6184),.clk(gclk));
	jor g05933(.dina(w_n6184_0[1]),.dinb(w_n6178_0[1]),.dout(n6185),.clk(gclk));
	jand g05934(.dina(n6185),.dinb(w_asqrt36_20[0]),.dout(n6186),.clk(gclk));
	jor g05935(.dina(w_n6178_0[0]),.dinb(w_asqrt36_19[2]),.dout(n6187),.clk(gclk));
	jor g05936(.dina(n6187),.dinb(w_n6184_0[0]),.dout(n6188),.clk(gclk));
	jnot g05937(.din(w_n5831_0[0]),.dout(n6189),.clk(gclk));
	jnot g05938(.din(w_n5833_0[0]),.dout(n6190),.clk(gclk));
	jand g05939(.dina(w_asqrt30_29[1]),.dinb(w_n5827_0[0]),.dout(n6191),.clk(gclk));
	jand g05940(.dina(w_n6191_0[1]),.dinb(n6190),.dout(n6192),.clk(gclk));
	jor g05941(.dina(n6192),.dinb(n6189),.dout(n6193),.clk(gclk));
	jnot g05942(.din(w_n5834_0[0]),.dout(n6194),.clk(gclk));
	jand g05943(.dina(w_n6191_0[0]),.dinb(n6194),.dout(n6195),.clk(gclk));
	jnot g05944(.din(n6195),.dout(n6196),.clk(gclk));
	jand g05945(.dina(n6196),.dinb(n6193),.dout(n6197),.clk(gclk));
	jand g05946(.dina(w_n6197_0[1]),.dinb(w_n6188_0[1]),.dout(n6198),.clk(gclk));
	jor g05947(.dina(n6198),.dinb(w_n6186_0[1]),.dout(n6199),.clk(gclk));
	jand g05948(.dina(w_n6199_0[2]),.dinb(w_asqrt37_17[1]),.dout(n6200),.clk(gclk));
	jor g05949(.dina(w_n6199_0[1]),.dinb(w_asqrt37_17[0]),.dout(n6201),.clk(gclk));
	jxor g05950(.dina(w_n5835_0[0]),.dinb(w_n4494_20[1]),.dout(n6202),.clk(gclk));
	jand g05951(.dina(n6202),.dinb(w_asqrt30_29[0]),.dout(n6203),.clk(gclk));
	jxor g05952(.dina(n6203),.dinb(w_n5840_0[0]),.dout(n6204),.clk(gclk));
	jand g05953(.dina(w_n6204_0[1]),.dinb(n6201),.dout(n6205),.clk(gclk));
	jor g05954(.dina(w_n6205_0[1]),.dinb(w_n6200_0[1]),.dout(n6206),.clk(gclk));
	jand g05955(.dina(n6206),.dinb(w_asqrt38_20[0]),.dout(n6207),.clk(gclk));
	jnot g05956(.din(w_n5846_0[0]),.dout(n6208),.clk(gclk));
	jand g05957(.dina(n6208),.dinb(w_n5844_0[0]),.dout(n6209),.clk(gclk));
	jand g05958(.dina(n6209),.dinb(w_asqrt30_28[2]),.dout(n6210),.clk(gclk));
	jxor g05959(.dina(n6210),.dinb(w_n5855_0[0]),.dout(n6211),.clk(gclk));
	jnot g05960(.din(n6211),.dout(n6212),.clk(gclk));
	jor g05961(.dina(w_n6200_0[0]),.dinb(w_asqrt38_19[2]),.dout(n6213),.clk(gclk));
	jor g05962(.dina(n6213),.dinb(w_n6205_0[0]),.dout(n6214),.clk(gclk));
	jand g05963(.dina(w_n6214_0[1]),.dinb(w_n6212_0[1]),.dout(n6215),.clk(gclk));
	jor g05964(.dina(w_n6215_0[1]),.dinb(w_n6207_0[1]),.dout(n6216),.clk(gclk));
	jand g05965(.dina(w_n6216_0[2]),.dinb(w_asqrt39_17[1]),.dout(n6217),.clk(gclk));
	jor g05966(.dina(w_n6216_0[1]),.dinb(w_asqrt39_17[0]),.dout(n6218),.clk(gclk));
	jxor g05967(.dina(w_n5857_0[0]),.dinb(w_n3907_20[1]),.dout(n6219),.clk(gclk));
	jand g05968(.dina(n6219),.dinb(w_asqrt30_28[1]),.dout(n6220),.clk(gclk));
	jxor g05969(.dina(n6220),.dinb(w_n5863_0[0]),.dout(n6221),.clk(gclk));
	jand g05970(.dina(w_n6221_0[1]),.dinb(n6218),.dout(n6222),.clk(gclk));
	jor g05971(.dina(w_n6222_0[1]),.dinb(w_n6217_0[1]),.dout(n6223),.clk(gclk));
	jand g05972(.dina(n6223),.dinb(w_asqrt40_20[0]),.dout(n6224),.clk(gclk));
	jor g05973(.dina(w_n6217_0[0]),.dinb(w_asqrt40_19[2]),.dout(n6225),.clk(gclk));
	jor g05974(.dina(n6225),.dinb(w_n6222_0[0]),.dout(n6226),.clk(gclk));
	jnot g05975(.din(w_n5871_0[0]),.dout(n6227),.clk(gclk));
	jnot g05976(.din(w_n5873_0[0]),.dout(n6228),.clk(gclk));
	jand g05977(.dina(w_asqrt30_28[0]),.dinb(w_n5867_0[0]),.dout(n6229),.clk(gclk));
	jand g05978(.dina(w_n6229_0[1]),.dinb(n6228),.dout(n6230),.clk(gclk));
	jor g05979(.dina(n6230),.dinb(n6227),.dout(n6231),.clk(gclk));
	jnot g05980(.din(w_n5874_0[0]),.dout(n6232),.clk(gclk));
	jand g05981(.dina(w_n6229_0[0]),.dinb(n6232),.dout(n6233),.clk(gclk));
	jnot g05982(.din(n6233),.dout(n6234),.clk(gclk));
	jand g05983(.dina(n6234),.dinb(n6231),.dout(n6235),.clk(gclk));
	jand g05984(.dina(w_n6235_0[1]),.dinb(w_n6226_0[1]),.dout(n6236),.clk(gclk));
	jor g05985(.dina(n6236),.dinb(w_n6224_0[1]),.dout(n6237),.clk(gclk));
	jand g05986(.dina(w_n6237_0[1]),.dinb(w_asqrt41_17[2]),.dout(n6238),.clk(gclk));
	jxor g05987(.dina(w_n5875_0[0]),.dinb(w_n3371_20[2]),.dout(n6239),.clk(gclk));
	jand g05988(.dina(n6239),.dinb(w_asqrt30_27[2]),.dout(n6240),.clk(gclk));
	jxor g05989(.dina(n6240),.dinb(w_n5882_0[0]),.dout(n6241),.clk(gclk));
	jnot g05990(.din(n6241),.dout(n6242),.clk(gclk));
	jor g05991(.dina(w_n6237_0[0]),.dinb(w_asqrt41_17[1]),.dout(n6243),.clk(gclk));
	jand g05992(.dina(w_n6243_0[1]),.dinb(w_n6242_0[1]),.dout(n6244),.clk(gclk));
	jor g05993(.dina(w_n6244_0[2]),.dinb(w_n6238_0[2]),.dout(n6245),.clk(gclk));
	jand g05994(.dina(n6245),.dinb(w_asqrt42_20[0]),.dout(n6246),.clk(gclk));
	jnot g05995(.din(w_n5887_0[0]),.dout(n6247),.clk(gclk));
	jand g05996(.dina(n6247),.dinb(w_n5885_0[0]),.dout(n6248),.clk(gclk));
	jand g05997(.dina(n6248),.dinb(w_asqrt30_27[1]),.dout(n6249),.clk(gclk));
	jxor g05998(.dina(n6249),.dinb(w_n5895_0[0]),.dout(n6250),.clk(gclk));
	jnot g05999(.din(n6250),.dout(n6251),.clk(gclk));
	jor g06000(.dina(w_n6238_0[1]),.dinb(w_asqrt42_19[2]),.dout(n6252),.clk(gclk));
	jor g06001(.dina(n6252),.dinb(w_n6244_0[1]),.dout(n6253),.clk(gclk));
	jand g06002(.dina(w_n6253_0[1]),.dinb(w_n6251_0[1]),.dout(n6254),.clk(gclk));
	jor g06003(.dina(w_n6254_0[1]),.dinb(w_n6246_0[1]),.dout(n6255),.clk(gclk));
	jand g06004(.dina(w_n6255_0[2]),.dinb(w_asqrt43_17[2]),.dout(n6256),.clk(gclk));
	jor g06005(.dina(w_n6255_0[1]),.dinb(w_asqrt43_17[1]),.dout(n6257),.clk(gclk));
	jnot g06006(.din(w_n5901_0[0]),.dout(n6258),.clk(gclk));
	jnot g06007(.din(w_n5902_0[0]),.dout(n6259),.clk(gclk));
	jand g06008(.dina(w_asqrt30_27[0]),.dinb(w_n5898_0[0]),.dout(n6260),.clk(gclk));
	jand g06009(.dina(w_n6260_0[1]),.dinb(n6259),.dout(n6261),.clk(gclk));
	jor g06010(.dina(n6261),.dinb(n6258),.dout(n6262),.clk(gclk));
	jnot g06011(.din(w_n5903_0[0]),.dout(n6263),.clk(gclk));
	jand g06012(.dina(w_n6260_0[0]),.dinb(n6263),.dout(n6264),.clk(gclk));
	jnot g06013(.din(n6264),.dout(n6265),.clk(gclk));
	jand g06014(.dina(n6265),.dinb(n6262),.dout(n6266),.clk(gclk));
	jand g06015(.dina(w_n6266_0[1]),.dinb(n6257),.dout(n6267),.clk(gclk));
	jor g06016(.dina(w_n6267_0[1]),.dinb(w_n6256_0[1]),.dout(n6268),.clk(gclk));
	jand g06017(.dina(n6268),.dinb(w_asqrt44_20[0]),.dout(n6269),.clk(gclk));
	jor g06018(.dina(w_n6256_0[0]),.dinb(w_asqrt44_19[2]),.dout(n6270),.clk(gclk));
	jor g06019(.dina(n6270),.dinb(w_n6267_0[0]),.dout(n6271),.clk(gclk));
	jnot g06020(.din(w_n5909_0[0]),.dout(n6272),.clk(gclk));
	jnot g06021(.din(w_n5911_0[0]),.dout(n6273),.clk(gclk));
	jand g06022(.dina(w_asqrt30_26[2]),.dinb(w_n5905_0[0]),.dout(n6274),.clk(gclk));
	jand g06023(.dina(w_n6274_0[1]),.dinb(n6273),.dout(n6275),.clk(gclk));
	jor g06024(.dina(n6275),.dinb(n6272),.dout(n6276),.clk(gclk));
	jnot g06025(.din(w_n5912_0[0]),.dout(n6277),.clk(gclk));
	jand g06026(.dina(w_n6274_0[0]),.dinb(n6277),.dout(n6278),.clk(gclk));
	jnot g06027(.din(n6278),.dout(n6279),.clk(gclk));
	jand g06028(.dina(n6279),.dinb(n6276),.dout(n6280),.clk(gclk));
	jand g06029(.dina(w_n6280_0[1]),.dinb(w_n6271_0[1]),.dout(n6281),.clk(gclk));
	jor g06030(.dina(n6281),.dinb(w_n6269_0[1]),.dout(n6282),.clk(gclk));
	jand g06031(.dina(w_n6282_0[1]),.dinb(w_asqrt45_18[0]),.dout(n6283),.clk(gclk));
	jxor g06032(.dina(w_n5913_0[0]),.dinb(w_n2420_21[2]),.dout(n6284),.clk(gclk));
	jand g06033(.dina(n6284),.dinb(w_asqrt30_26[1]),.dout(n6285),.clk(gclk));
	jxor g06034(.dina(n6285),.dinb(w_n5923_0[0]),.dout(n6286),.clk(gclk));
	jnot g06035(.din(n6286),.dout(n6287),.clk(gclk));
	jor g06036(.dina(w_n6282_0[0]),.dinb(w_asqrt45_17[2]),.dout(n6288),.clk(gclk));
	jand g06037(.dina(w_n6288_0[1]),.dinb(w_n6287_0[1]),.dout(n6289),.clk(gclk));
	jor g06038(.dina(w_n6289_0[2]),.dinb(w_n6283_0[2]),.dout(n6290),.clk(gclk));
	jand g06039(.dina(n6290),.dinb(w_asqrt46_20[0]),.dout(n6291),.clk(gclk));
	jnot g06040(.din(w_n5928_0[0]),.dout(n6292),.clk(gclk));
	jand g06041(.dina(n6292),.dinb(w_n5926_0[0]),.dout(n6293),.clk(gclk));
	jand g06042(.dina(n6293),.dinb(w_asqrt30_26[0]),.dout(n6294),.clk(gclk));
	jxor g06043(.dina(n6294),.dinb(w_n5936_0[0]),.dout(n6295),.clk(gclk));
	jnot g06044(.din(n6295),.dout(n6296),.clk(gclk));
	jor g06045(.dina(w_n6283_0[1]),.dinb(w_asqrt46_19[2]),.dout(n6297),.clk(gclk));
	jor g06046(.dina(n6297),.dinb(w_n6289_0[1]),.dout(n6298),.clk(gclk));
	jand g06047(.dina(w_n6298_0[1]),.dinb(w_n6296_0[1]),.dout(n6299),.clk(gclk));
	jor g06048(.dina(w_n6299_0[1]),.dinb(w_n6291_0[1]),.dout(n6300),.clk(gclk));
	jand g06049(.dina(w_n6300_0[2]),.dinb(w_asqrt47_18[0]),.dout(n6301),.clk(gclk));
	jor g06050(.dina(w_n6300_0[1]),.dinb(w_asqrt47_17[2]),.dout(n6302),.clk(gclk));
	jnot g06051(.din(w_n5942_0[0]),.dout(n6303),.clk(gclk));
	jnot g06052(.din(w_n5943_0[0]),.dout(n6304),.clk(gclk));
	jand g06053(.dina(w_asqrt30_25[2]),.dinb(w_n5939_0[0]),.dout(n6305),.clk(gclk));
	jand g06054(.dina(w_n6305_0[1]),.dinb(n6304),.dout(n6306),.clk(gclk));
	jor g06055(.dina(n6306),.dinb(n6303),.dout(n6307),.clk(gclk));
	jnot g06056(.din(w_n5944_0[0]),.dout(n6308),.clk(gclk));
	jand g06057(.dina(w_n6305_0[0]),.dinb(n6308),.dout(n6309),.clk(gclk));
	jnot g06058(.din(n6309),.dout(n6310),.clk(gclk));
	jand g06059(.dina(n6310),.dinb(n6307),.dout(n6311),.clk(gclk));
	jand g06060(.dina(w_n6311_0[1]),.dinb(n6302),.dout(n6312),.clk(gclk));
	jor g06061(.dina(w_n6312_0[1]),.dinb(w_n6301_0[1]),.dout(n6313),.clk(gclk));
	jand g06062(.dina(n6313),.dinb(w_asqrt48_20[0]),.dout(n6314),.clk(gclk));
	jor g06063(.dina(w_n6301_0[0]),.dinb(w_asqrt48_19[2]),.dout(n6315),.clk(gclk));
	jor g06064(.dina(n6315),.dinb(w_n6312_0[0]),.dout(n6316),.clk(gclk));
	jnot g06065(.din(w_n5950_0[0]),.dout(n6317),.clk(gclk));
	jnot g06066(.din(w_n5952_0[0]),.dout(n6318),.clk(gclk));
	jand g06067(.dina(w_asqrt30_25[1]),.dinb(w_n5946_0[0]),.dout(n6319),.clk(gclk));
	jand g06068(.dina(w_n6319_0[1]),.dinb(n6318),.dout(n6320),.clk(gclk));
	jor g06069(.dina(n6320),.dinb(n6317),.dout(n6321),.clk(gclk));
	jnot g06070(.din(w_n5953_0[0]),.dout(n6322),.clk(gclk));
	jand g06071(.dina(w_n6319_0[0]),.dinb(n6322),.dout(n6323),.clk(gclk));
	jnot g06072(.din(n6323),.dout(n6324),.clk(gclk));
	jand g06073(.dina(n6324),.dinb(n6321),.dout(n6325),.clk(gclk));
	jand g06074(.dina(w_n6325_0[1]),.dinb(w_n6316_0[1]),.dout(n6326),.clk(gclk));
	jor g06075(.dina(n6326),.dinb(w_n6314_0[1]),.dout(n6327),.clk(gclk));
	jand g06076(.dina(w_n6327_0[1]),.dinb(w_asqrt49_18[1]),.dout(n6328),.clk(gclk));
	jxor g06077(.dina(w_n5954_0[0]),.dinb(w_n1641_22[1]),.dout(n6329),.clk(gclk));
	jand g06078(.dina(n6329),.dinb(w_asqrt30_25[0]),.dout(n6330),.clk(gclk));
	jxor g06079(.dina(n6330),.dinb(w_n5964_0[0]),.dout(n6331),.clk(gclk));
	jnot g06080(.din(n6331),.dout(n6332),.clk(gclk));
	jor g06081(.dina(w_n6327_0[0]),.dinb(w_asqrt49_18[0]),.dout(n6333),.clk(gclk));
	jand g06082(.dina(w_n6333_0[1]),.dinb(w_n6332_0[1]),.dout(n6334),.clk(gclk));
	jor g06083(.dina(w_n6334_0[2]),.dinb(w_n6328_0[2]),.dout(n6335),.clk(gclk));
	jand g06084(.dina(n6335),.dinb(w_asqrt50_20[0]),.dout(n6336),.clk(gclk));
	jnot g06085(.din(w_n5969_0[0]),.dout(n6337),.clk(gclk));
	jand g06086(.dina(n6337),.dinb(w_n5967_0[0]),.dout(n6338),.clk(gclk));
	jand g06087(.dina(n6338),.dinb(w_asqrt30_24[2]),.dout(n6339),.clk(gclk));
	jxor g06088(.dina(n6339),.dinb(w_n5977_0[0]),.dout(n6340),.clk(gclk));
	jnot g06089(.din(n6340),.dout(n6341),.clk(gclk));
	jor g06090(.dina(w_n6328_0[1]),.dinb(w_asqrt50_19[2]),.dout(n6342),.clk(gclk));
	jor g06091(.dina(n6342),.dinb(w_n6334_0[1]),.dout(n6343),.clk(gclk));
	jand g06092(.dina(w_n6343_0[1]),.dinb(w_n6341_0[1]),.dout(n6344),.clk(gclk));
	jor g06093(.dina(w_n6344_0[1]),.dinb(w_n6336_0[1]),.dout(n6345),.clk(gclk));
	jand g06094(.dina(w_n6345_0[2]),.dinb(w_asqrt51_18[1]),.dout(n6346),.clk(gclk));
	jor g06095(.dina(w_n6345_0[1]),.dinb(w_asqrt51_18[0]),.dout(n6347),.clk(gclk));
	jnot g06096(.din(w_n5983_0[0]),.dout(n6348),.clk(gclk));
	jnot g06097(.din(w_n5984_0[0]),.dout(n6349),.clk(gclk));
	jand g06098(.dina(w_asqrt30_24[1]),.dinb(w_n5980_0[0]),.dout(n6350),.clk(gclk));
	jand g06099(.dina(w_n6350_0[1]),.dinb(n6349),.dout(n6351),.clk(gclk));
	jor g06100(.dina(n6351),.dinb(n6348),.dout(n6352),.clk(gclk));
	jnot g06101(.din(w_n5985_0[0]),.dout(n6353),.clk(gclk));
	jand g06102(.dina(w_n6350_0[0]),.dinb(n6353),.dout(n6354),.clk(gclk));
	jnot g06103(.din(n6354),.dout(n6355),.clk(gclk));
	jand g06104(.dina(n6355),.dinb(n6352),.dout(n6356),.clk(gclk));
	jand g06105(.dina(w_n6356_0[1]),.dinb(n6347),.dout(n6357),.clk(gclk));
	jor g06106(.dina(w_n6357_0[1]),.dinb(w_n6346_0[1]),.dout(n6358),.clk(gclk));
	jand g06107(.dina(n6358),.dinb(w_asqrt52_20[0]),.dout(n6359),.clk(gclk));
	jor g06108(.dina(w_n6346_0[0]),.dinb(w_asqrt52_19[2]),.dout(n6360),.clk(gclk));
	jor g06109(.dina(n6360),.dinb(w_n6357_0[0]),.dout(n6361),.clk(gclk));
	jnot g06110(.din(w_n5991_0[0]),.dout(n6362),.clk(gclk));
	jnot g06111(.din(w_n5993_0[0]),.dout(n6363),.clk(gclk));
	jand g06112(.dina(w_asqrt30_24[0]),.dinb(w_n5987_0[0]),.dout(n6364),.clk(gclk));
	jand g06113(.dina(w_n6364_0[1]),.dinb(n6363),.dout(n6365),.clk(gclk));
	jor g06114(.dina(n6365),.dinb(n6362),.dout(n6366),.clk(gclk));
	jnot g06115(.din(w_n5994_0[0]),.dout(n6367),.clk(gclk));
	jand g06116(.dina(w_n6364_0[0]),.dinb(n6367),.dout(n6368),.clk(gclk));
	jnot g06117(.din(n6368),.dout(n6369),.clk(gclk));
	jand g06118(.dina(n6369),.dinb(n6366),.dout(n6370),.clk(gclk));
	jand g06119(.dina(w_n6370_0[1]),.dinb(w_n6361_0[1]),.dout(n6371),.clk(gclk));
	jor g06120(.dina(n6371),.dinb(w_n6359_0[1]),.dout(n6372),.clk(gclk));
	jand g06121(.dina(w_n6372_0[1]),.dinb(w_asqrt53_18[2]),.dout(n6373),.clk(gclk));
	jxor g06122(.dina(w_n5995_0[0]),.dinb(w_n1034_23[1]),.dout(n6374),.clk(gclk));
	jand g06123(.dina(n6374),.dinb(w_asqrt30_23[2]),.dout(n6375),.clk(gclk));
	jxor g06124(.dina(n6375),.dinb(w_n6005_0[0]),.dout(n6376),.clk(gclk));
	jnot g06125(.din(n6376),.dout(n6377),.clk(gclk));
	jor g06126(.dina(w_n6372_0[0]),.dinb(w_asqrt53_18[1]),.dout(n6378),.clk(gclk));
	jand g06127(.dina(w_n6378_0[1]),.dinb(w_n6377_0[1]),.dout(n6379),.clk(gclk));
	jor g06128(.dina(w_n6379_0[2]),.dinb(w_n6373_0[2]),.dout(n6380),.clk(gclk));
	jand g06129(.dina(n6380),.dinb(w_asqrt54_20[0]),.dout(n6381),.clk(gclk));
	jnot g06130(.din(w_n6010_0[0]),.dout(n6382),.clk(gclk));
	jand g06131(.dina(n6382),.dinb(w_n6008_0[0]),.dout(n6383),.clk(gclk));
	jand g06132(.dina(n6383),.dinb(w_asqrt30_23[1]),.dout(n6384),.clk(gclk));
	jxor g06133(.dina(n6384),.dinb(w_n6018_0[0]),.dout(n6385),.clk(gclk));
	jnot g06134(.din(n6385),.dout(n6386),.clk(gclk));
	jor g06135(.dina(w_n6373_0[1]),.dinb(w_asqrt54_19[2]),.dout(n6387),.clk(gclk));
	jor g06136(.dina(n6387),.dinb(w_n6379_0[1]),.dout(n6388),.clk(gclk));
	jand g06137(.dina(w_n6388_0[1]),.dinb(w_n6386_0[1]),.dout(n6389),.clk(gclk));
	jor g06138(.dina(w_n6389_0[1]),.dinb(w_n6381_0[1]),.dout(n6390),.clk(gclk));
	jand g06139(.dina(w_n6390_0[2]),.dinb(w_asqrt55_19[0]),.dout(n6391),.clk(gclk));
	jor g06140(.dina(w_n6390_0[1]),.dinb(w_asqrt55_18[2]),.dout(n6392),.clk(gclk));
	jnot g06141(.din(w_n6024_0[0]),.dout(n6393),.clk(gclk));
	jnot g06142(.din(w_n6025_0[0]),.dout(n6394),.clk(gclk));
	jand g06143(.dina(w_asqrt30_23[0]),.dinb(w_n6021_0[0]),.dout(n6395),.clk(gclk));
	jand g06144(.dina(w_n6395_0[1]),.dinb(n6394),.dout(n6396),.clk(gclk));
	jor g06145(.dina(n6396),.dinb(n6393),.dout(n6397),.clk(gclk));
	jnot g06146(.din(w_n6026_0[0]),.dout(n6398),.clk(gclk));
	jand g06147(.dina(w_n6395_0[0]),.dinb(n6398),.dout(n6399),.clk(gclk));
	jnot g06148(.din(n6399),.dout(n6400),.clk(gclk));
	jand g06149(.dina(n6400),.dinb(n6397),.dout(n6401),.clk(gclk));
	jand g06150(.dina(w_n6401_0[1]),.dinb(n6392),.dout(n6402),.clk(gclk));
	jor g06151(.dina(w_n6402_0[1]),.dinb(w_n6391_0[1]),.dout(n6403),.clk(gclk));
	jand g06152(.dina(n6403),.dinb(w_asqrt56_20[0]),.dout(n6404),.clk(gclk));
	jor g06153(.dina(w_n6391_0[0]),.dinb(w_asqrt56_19[2]),.dout(n6405),.clk(gclk));
	jor g06154(.dina(n6405),.dinb(w_n6402_0[0]),.dout(n6406),.clk(gclk));
	jnot g06155(.din(w_n6032_0[0]),.dout(n6407),.clk(gclk));
	jnot g06156(.din(w_n6034_0[0]),.dout(n6408),.clk(gclk));
	jand g06157(.dina(w_asqrt30_22[2]),.dinb(w_n6028_0[0]),.dout(n6409),.clk(gclk));
	jand g06158(.dina(w_n6409_0[1]),.dinb(n6408),.dout(n6410),.clk(gclk));
	jor g06159(.dina(n6410),.dinb(n6407),.dout(n6411),.clk(gclk));
	jnot g06160(.din(w_n6035_0[0]),.dout(n6412),.clk(gclk));
	jand g06161(.dina(w_n6409_0[0]),.dinb(n6412),.dout(n6413),.clk(gclk));
	jnot g06162(.din(n6413),.dout(n6414),.clk(gclk));
	jand g06163(.dina(n6414),.dinb(n6411),.dout(n6415),.clk(gclk));
	jand g06164(.dina(w_n6415_0[1]),.dinb(w_n6406_0[1]),.dout(n6416),.clk(gclk));
	jor g06165(.dina(n6416),.dinb(w_n6404_0[1]),.dout(n6417),.clk(gclk));
	jand g06166(.dina(w_n6417_0[1]),.dinb(w_asqrt57_19[1]),.dout(n6418),.clk(gclk));
	jxor g06167(.dina(w_n6036_0[0]),.dinb(w_n590_24[0]),.dout(n6419),.clk(gclk));
	jand g06168(.dina(n6419),.dinb(w_asqrt30_22[1]),.dout(n6420),.clk(gclk));
	jxor g06169(.dina(n6420),.dinb(w_n6046_0[0]),.dout(n6421),.clk(gclk));
	jnot g06170(.din(n6421),.dout(n6422),.clk(gclk));
	jor g06171(.dina(w_n6417_0[0]),.dinb(w_asqrt57_19[0]),.dout(n6423),.clk(gclk));
	jand g06172(.dina(w_n6423_0[1]),.dinb(w_n6422_0[1]),.dout(n6424),.clk(gclk));
	jor g06173(.dina(w_n6424_0[2]),.dinb(w_n6418_0[2]),.dout(n6425),.clk(gclk));
	jand g06174(.dina(n6425),.dinb(w_asqrt58_20[0]),.dout(n6426),.clk(gclk));
	jnot g06175(.din(w_n6051_0[0]),.dout(n6427),.clk(gclk));
	jand g06176(.dina(n6427),.dinb(w_n6049_0[0]),.dout(n6428),.clk(gclk));
	jand g06177(.dina(n6428),.dinb(w_asqrt30_22[0]),.dout(n6429),.clk(gclk));
	jxor g06178(.dina(n6429),.dinb(w_n6059_0[0]),.dout(n6430),.clk(gclk));
	jnot g06179(.din(n6430),.dout(n6431),.clk(gclk));
	jor g06180(.dina(w_n6418_0[1]),.dinb(w_asqrt58_19[2]),.dout(n6432),.clk(gclk));
	jor g06181(.dina(n6432),.dinb(w_n6424_0[1]),.dout(n6433),.clk(gclk));
	jand g06182(.dina(w_n6433_0[1]),.dinb(w_n6431_0[1]),.dout(n6434),.clk(gclk));
	jor g06183(.dina(w_n6434_0[1]),.dinb(w_n6426_0[1]),.dout(n6435),.clk(gclk));
	jand g06184(.dina(w_n6435_0[2]),.dinb(w_asqrt59_19[2]),.dout(n6436),.clk(gclk));
	jor g06185(.dina(w_n6435_0[1]),.dinb(w_asqrt59_19[1]),.dout(n6437),.clk(gclk));
	jnot g06186(.din(w_n6065_0[0]),.dout(n6438),.clk(gclk));
	jnot g06187(.din(w_n6066_0[0]),.dout(n6439),.clk(gclk));
	jand g06188(.dina(w_asqrt30_21[2]),.dinb(w_n6062_0[0]),.dout(n6440),.clk(gclk));
	jand g06189(.dina(w_n6440_0[1]),.dinb(n6439),.dout(n6441),.clk(gclk));
	jor g06190(.dina(n6441),.dinb(n6438),.dout(n6442),.clk(gclk));
	jnot g06191(.din(w_n6067_0[0]),.dout(n6443),.clk(gclk));
	jand g06192(.dina(w_n6440_0[0]),.dinb(n6443),.dout(n6444),.clk(gclk));
	jnot g06193(.din(n6444),.dout(n6445),.clk(gclk));
	jand g06194(.dina(n6445),.dinb(n6442),.dout(n6446),.clk(gclk));
	jand g06195(.dina(w_n6446_0[1]),.dinb(n6437),.dout(n6447),.clk(gclk));
	jor g06196(.dina(w_n6447_0[1]),.dinb(w_n6436_0[1]),.dout(n6448),.clk(gclk));
	jand g06197(.dina(n6448),.dinb(w_asqrt60_19[2]),.dout(n6449),.clk(gclk));
	jor g06198(.dina(w_n6436_0[0]),.dinb(w_asqrt60_19[1]),.dout(n6450),.clk(gclk));
	jor g06199(.dina(n6450),.dinb(w_n6447_0[0]),.dout(n6451),.clk(gclk));
	jnot g06200(.din(w_n6073_0[0]),.dout(n6452),.clk(gclk));
	jnot g06201(.din(w_n6075_0[0]),.dout(n6453),.clk(gclk));
	jand g06202(.dina(w_asqrt30_21[1]),.dinb(w_n6069_0[0]),.dout(n6454),.clk(gclk));
	jand g06203(.dina(w_n6454_0[1]),.dinb(n6453),.dout(n6455),.clk(gclk));
	jor g06204(.dina(n6455),.dinb(n6452),.dout(n6456),.clk(gclk));
	jnot g06205(.din(w_n6076_0[0]),.dout(n6457),.clk(gclk));
	jand g06206(.dina(w_n6454_0[0]),.dinb(n6457),.dout(n6458),.clk(gclk));
	jnot g06207(.din(n6458),.dout(n6459),.clk(gclk));
	jand g06208(.dina(n6459),.dinb(n6456),.dout(n6460),.clk(gclk));
	jand g06209(.dina(w_n6460_0[1]),.dinb(w_n6451_0[1]),.dout(n6461),.clk(gclk));
	jor g06210(.dina(n6461),.dinb(w_n6449_0[1]),.dout(n6462),.clk(gclk));
	jand g06211(.dina(w_n6462_0[1]),.dinb(w_asqrt61_20[0]),.dout(n6463),.clk(gclk));
	jxor g06212(.dina(w_n6077_0[0]),.dinb(w_n290_25[1]),.dout(n6464),.clk(gclk));
	jand g06213(.dina(n6464),.dinb(w_asqrt30_21[0]),.dout(n6465),.clk(gclk));
	jxor g06214(.dina(n6465),.dinb(w_n6087_0[0]),.dout(n6466),.clk(gclk));
	jnot g06215(.din(n6466),.dout(n6467),.clk(gclk));
	jor g06216(.dina(w_n6462_0[0]),.dinb(w_asqrt61_19[2]),.dout(n6468),.clk(gclk));
	jand g06217(.dina(w_n6468_0[1]),.dinb(w_n6467_0[1]),.dout(n6469),.clk(gclk));
	jor g06218(.dina(w_n6469_0[2]),.dinb(w_n6463_0[2]),.dout(n6470),.clk(gclk));
	jand g06219(.dina(n6470),.dinb(w_asqrt62_20[0]),.dout(n6471),.clk(gclk));
	jnot g06220(.din(w_n6092_0[0]),.dout(n6472),.clk(gclk));
	jand g06221(.dina(n6472),.dinb(w_n6090_0[0]),.dout(n6473),.clk(gclk));
	jand g06222(.dina(n6473),.dinb(w_asqrt30_20[2]),.dout(n6474),.clk(gclk));
	jxor g06223(.dina(n6474),.dinb(w_n6100_0[0]),.dout(n6475),.clk(gclk));
	jnot g06224(.din(n6475),.dout(n6476),.clk(gclk));
	jor g06225(.dina(w_n6463_0[1]),.dinb(w_asqrt62_19[2]),.dout(n6477),.clk(gclk));
	jor g06226(.dina(n6477),.dinb(w_n6469_0[1]),.dout(n6478),.clk(gclk));
	jand g06227(.dina(w_n6478_0[1]),.dinb(w_n6476_0[1]),.dout(n6479),.clk(gclk));
	jor g06228(.dina(w_n6479_0[1]),.dinb(w_n6471_0[1]),.dout(n6480),.clk(gclk));
	jxor g06229(.dina(w_n6102_0[0]),.dinb(w_n199_29[2]),.dout(n6481),.clk(gclk));
	jand g06230(.dina(n6481),.dinb(w_asqrt30_20[1]),.dout(n6482),.clk(gclk));
	jxor g06231(.dina(n6482),.dinb(w_n6107_0[0]),.dout(n6483),.clk(gclk));
	jnot g06232(.din(w_n6109_0[0]),.dout(n6484),.clk(gclk));
	jnot g06233(.din(w_n6113_0[0]),.dout(n6485),.clk(gclk));
	jand g06234(.dina(w_asqrt30_20[0]),.dinb(w_n6485_0[1]),.dout(n6486),.clk(gclk));
	jand g06235(.dina(w_n6486_0[1]),.dinb(w_n6484_0[2]),.dout(n6487),.clk(gclk));
	jor g06236(.dina(n6487),.dinb(w_n6120_0[0]),.dout(n6488),.clk(gclk));
	jor g06237(.dina(n6488),.dinb(w_n6483_0[1]),.dout(n6489),.clk(gclk));
	jnot g06238(.din(n6489),.dout(n6490),.clk(gclk));
	jand g06239(.dina(n6490),.dinb(w_n6480_1[2]),.dout(n6491),.clk(gclk));
	jor g06240(.dina(n6491),.dinb(w_asqrt63_10[2]),.dout(n6492),.clk(gclk));
	jnot g06241(.din(w_n6483_0[0]),.dout(n6493),.clk(gclk));
	jor g06242(.dina(w_n6493_0[2]),.dinb(w_n6480_1[1]),.dout(n6494),.clk(gclk));
	jor g06243(.dina(w_n6486_0[0]),.dinb(w_n6484_0[1]),.dout(n6495),.clk(gclk));
	jand g06244(.dina(w_n6485_0[0]),.dinb(w_n6484_0[0]),.dout(n6496),.clk(gclk));
	jor g06245(.dina(n6496),.dinb(w_n194_28[2]),.dout(n6497),.clk(gclk));
	jnot g06246(.din(n6497),.dout(n6498),.clk(gclk));
	jand g06247(.dina(n6498),.dinb(n6495),.dout(n6499),.clk(gclk));
	jnot g06248(.din(w_asqrt30_19[2]),.dout(n6500),.clk(gclk));
	jnot g06249(.din(w_n6499_0[1]),.dout(n6503),.clk(gclk));
	jand g06250(.dina(n6503),.dinb(w_n6494_0[1]),.dout(n6504),.clk(gclk));
	jand g06251(.dina(n6504),.dinb(w_n6492_0[1]),.dout(n6505),.clk(gclk));
	jxor g06252(.dina(w_n6158_0[0]),.dinb(w_n5121_22[1]),.dout(n6506),.clk(gclk));
	jor g06253(.dina(n6506),.dinb(w_n6505_28[1]),.dout(n6507),.clk(gclk));
	jxor g06254(.dina(n6507),.dinb(w_n6132_0[0]),.dout(n6508),.clk(gclk));
	jor g06255(.dina(w_n6505_28[0]),.dinb(w_n6134_1[0]),.dout(n6509),.clk(gclk));
	jnot g06256(.din(w_a56_0[1]),.dout(n6510),.clk(gclk));
	jnot g06257(.din(a[57]),.dout(n6511),.clk(gclk));
	jand g06258(.dina(w_n6134_0[2]),.dinb(w_n6511_0[2]),.dout(n6512),.clk(gclk));
	jand g06259(.dina(n6512),.dinb(w_n6510_1[1]),.dout(n6513),.clk(gclk));
	jnot g06260(.din(n6513),.dout(n6514),.clk(gclk));
	jand g06261(.dina(n6514),.dinb(n6509),.dout(n6515),.clk(gclk));
	jor g06262(.dina(w_n6515_0[2]),.dinb(w_n6500_19[1]),.dout(n6516),.clk(gclk));
	jor g06263(.dina(w_n6505_27[2]),.dinb(w_a58_0[0]),.dout(n6517),.clk(gclk));
	jxor g06264(.dina(w_n6517_0[1]),.dinb(w_n6135_0[0]),.dout(n6518),.clk(gclk));
	jand g06265(.dina(w_n6515_0[1]),.dinb(w_n6500_19[0]),.dout(n6519),.clk(gclk));
	jor g06266(.dina(n6519),.dinb(w_n6518_0[1]),.dout(n6520),.clk(gclk));
	jand g06267(.dina(w_n6520_0[1]),.dinb(w_n6516_0[1]),.dout(n6521),.clk(gclk));
	jor g06268(.dina(n6521),.dinb(w_n5793_22[2]),.dout(n6522),.clk(gclk));
	jand g06269(.dina(w_n6516_0[0]),.dinb(w_n5793_22[1]),.dout(n6523),.clk(gclk));
	jand g06270(.dina(n6523),.dinb(w_n6520_0[0]),.dout(n6524),.clk(gclk));
	jor g06271(.dina(w_n6517_0[0]),.dinb(w_a59_0[0]),.dout(n6525),.clk(gclk));
	jnot g06272(.din(w_n6492_0[0]),.dout(n6526),.clk(gclk));
	jnot g06273(.din(w_n6494_0[0]),.dout(n6527),.clk(gclk));
	jor g06274(.dina(w_n6499_0[0]),.dinb(w_n6500_18[2]),.dout(n6528),.clk(gclk));
	jor g06275(.dina(n6528),.dinb(w_n6527_0[1]),.dout(n6529),.clk(gclk));
	jor g06276(.dina(n6529),.dinb(n6526),.dout(n6530),.clk(gclk));
	jand g06277(.dina(n6530),.dinb(n6525),.dout(n6531),.clk(gclk));
	jxor g06278(.dina(n6531),.dinb(w_n5797_0[1]),.dout(n6532),.clk(gclk));
	jor g06279(.dina(w_n6532_0[1]),.dinb(w_n6524_0[1]),.dout(n6533),.clk(gclk));
	jand g06280(.dina(n6533),.dinb(w_n6522_0[1]),.dout(n6534),.clk(gclk));
	jor g06281(.dina(w_n6534_0[2]),.dinb(w_n5788_19[1]),.dout(n6535),.clk(gclk));
	jand g06282(.dina(w_n6534_0[1]),.dinb(w_n5788_19[0]),.dout(n6536),.clk(gclk));
	jxor g06283(.dina(w_n6138_0[0]),.dinb(w_n5793_22[0]),.dout(n6537),.clk(gclk));
	jor g06284(.dina(n6537),.dinb(w_n6505_27[1]),.dout(n6538),.clk(gclk));
	jxor g06285(.dina(n6538),.dinb(w_n6141_0[0]),.dout(n6539),.clk(gclk));
	jor g06286(.dina(w_n6539_0[1]),.dinb(n6536),.dout(n6540),.clk(gclk));
	jand g06287(.dina(w_n6540_0[1]),.dinb(w_n6535_0[1]),.dout(n6541),.clk(gclk));
	jor g06288(.dina(n6541),.dinb(w_n5121_22[0]),.dout(n6542),.clk(gclk));
	jand g06289(.dina(w_n6535_0[0]),.dinb(w_n5121_21[2]),.dout(n6543),.clk(gclk));
	jand g06290(.dina(n6543),.dinb(w_n6540_0[0]),.dout(n6544),.clk(gclk));
	jnot g06291(.din(w_n6145_0[0]),.dout(n6545),.clk(gclk));
	jnot g06292(.din(w_n6505_27[0]),.dout(asqrt_fa_30),.clk(gclk));
	jand g06293(.dina(w_asqrt29_21[1]),.dinb(n6545),.dout(n6547),.clk(gclk));
	jand g06294(.dina(w_n6547_0[1]),.dinb(w_n6156_0[0]),.dout(n6548),.clk(gclk));
	jor g06295(.dina(n6548),.dinb(w_n6154_0[0]),.dout(n6549),.clk(gclk));
	jand g06296(.dina(w_n6547_0[0]),.dinb(w_n6157_0[0]),.dout(n6550),.clk(gclk));
	jnot g06297(.din(n6550),.dout(n6551),.clk(gclk));
	jand g06298(.dina(n6551),.dinb(n6549),.dout(n6552),.clk(gclk));
	jnot g06299(.din(n6552),.dout(n6553),.clk(gclk));
	jor g06300(.dina(w_n6553_0[1]),.dinb(w_n6544_0[1]),.dout(n6554),.clk(gclk));
	jand g06301(.dina(n6554),.dinb(w_n6542_0[1]),.dout(n6555),.clk(gclk));
	jor g06302(.dina(w_n6555_0[2]),.dinb(w_n5116_19[1]),.dout(n6556),.clk(gclk));
	jnot g06303(.din(w_n6508_0[1]),.dout(n6557),.clk(gclk));
	jand g06304(.dina(w_n6555_0[1]),.dinb(w_n5116_19[0]),.dout(n6558),.clk(gclk));
	jor g06305(.dina(n6558),.dinb(n6557),.dout(n6559),.clk(gclk));
	jand g06306(.dina(w_n6559_0[1]),.dinb(w_n6556_0[1]),.dout(n6560),.clk(gclk));
	jor g06307(.dina(n6560),.dinb(w_n4499_23[0]),.dout(n6561),.clk(gclk));
	jnot g06308(.din(w_n6166_0[0]),.dout(n6562),.clk(gclk));
	jor g06309(.dina(n6562),.dinb(w_n6164_0[0]),.dout(n6563),.clk(gclk));
	jor g06310(.dina(n6563),.dinb(w_n6505_26[2]),.dout(n6564),.clk(gclk));
	jxor g06311(.dina(n6564),.dinb(w_n6175_0[0]),.dout(n6565),.clk(gclk));
	jand g06312(.dina(w_n6556_0[0]),.dinb(w_n4499_22[2]),.dout(n6566),.clk(gclk));
	jand g06313(.dina(n6566),.dinb(w_n6559_0[0]),.dout(n6567),.clk(gclk));
	jor g06314(.dina(w_n6567_0[1]),.dinb(w_n6565_0[1]),.dout(n6568),.clk(gclk));
	jand g06315(.dina(w_n6568_0[1]),.dinb(w_n6561_0[1]),.dout(n6569),.clk(gclk));
	jor g06316(.dina(w_n6569_0[2]),.dinb(w_n4494_20[0]),.dout(n6570),.clk(gclk));
	jand g06317(.dina(w_n6569_0[1]),.dinb(w_n4494_19[2]),.dout(n6571),.clk(gclk));
	jnot g06318(.din(w_n6183_0[0]),.dout(n6572),.clk(gclk));
	jxor g06319(.dina(w_n6177_0[0]),.dinb(w_n4499_22[1]),.dout(n6573),.clk(gclk));
	jor g06320(.dina(n6573),.dinb(w_n6505_26[1]),.dout(n6574),.clk(gclk));
	jxor g06321(.dina(n6574),.dinb(n6572),.dout(n6575),.clk(gclk));
	jnot g06322(.din(w_n6575_0[1]),.dout(n6576),.clk(gclk));
	jor g06323(.dina(n6576),.dinb(n6571),.dout(n6577),.clk(gclk));
	jand g06324(.dina(w_n6577_0[1]),.dinb(w_n6570_0[1]),.dout(n6578),.clk(gclk));
	jor g06325(.dina(n6578),.dinb(w_n3912_23[0]),.dout(n6579),.clk(gclk));
	jnot g06326(.din(w_n6188_0[0]),.dout(n6580),.clk(gclk));
	jor g06327(.dina(n6580),.dinb(w_n6186_0[0]),.dout(n6581),.clk(gclk));
	jor g06328(.dina(n6581),.dinb(w_n6505_26[0]),.dout(n6582),.clk(gclk));
	jxor g06329(.dina(n6582),.dinb(w_n6197_0[0]),.dout(n6583),.clk(gclk));
	jand g06330(.dina(w_n6570_0[0]),.dinb(w_n3912_22[2]),.dout(n6584),.clk(gclk));
	jand g06331(.dina(n6584),.dinb(w_n6577_0[0]),.dout(n6585),.clk(gclk));
	jor g06332(.dina(w_n6585_0[1]),.dinb(w_n6583_0[1]),.dout(n6586),.clk(gclk));
	jand g06333(.dina(w_n6586_0[1]),.dinb(w_n6579_0[1]),.dout(n6587),.clk(gclk));
	jor g06334(.dina(w_n6587_0[2]),.dinb(w_n3907_20[0]),.dout(n6588),.clk(gclk));
	jand g06335(.dina(w_n6587_0[1]),.dinb(w_n3907_19[2]),.dout(n6589),.clk(gclk));
	jnot g06336(.din(w_n6204_0[0]),.dout(n6590),.clk(gclk));
	jxor g06337(.dina(w_n6199_0[0]),.dinb(w_n3912_22[1]),.dout(n6591),.clk(gclk));
	jor g06338(.dina(n6591),.dinb(w_n6505_25[2]),.dout(n6592),.clk(gclk));
	jxor g06339(.dina(n6592),.dinb(n6590),.dout(n6593),.clk(gclk));
	jnot g06340(.din(n6593),.dout(n6594),.clk(gclk));
	jor g06341(.dina(w_n6594_0[1]),.dinb(n6589),.dout(n6595),.clk(gclk));
	jand g06342(.dina(w_n6595_0[1]),.dinb(w_n6588_0[1]),.dout(n6596),.clk(gclk));
	jor g06343(.dina(n6596),.dinb(w_n3376_23[2]),.dout(n6597),.clk(gclk));
	jand g06344(.dina(w_n6588_0[0]),.dinb(w_n3376_23[1]),.dout(n6598),.clk(gclk));
	jand g06345(.dina(n6598),.dinb(w_n6595_0[0]),.dout(n6599),.clk(gclk));
	jnot g06346(.din(w_n6207_0[0]),.dout(n6600),.clk(gclk));
	jand g06347(.dina(w_asqrt29_21[0]),.dinb(n6600),.dout(n6601),.clk(gclk));
	jand g06348(.dina(w_n6601_0[1]),.dinb(w_n6214_0[0]),.dout(n6602),.clk(gclk));
	jor g06349(.dina(n6602),.dinb(w_n6212_0[0]),.dout(n6603),.clk(gclk));
	jand g06350(.dina(w_n6601_0[0]),.dinb(w_n6215_0[0]),.dout(n6604),.clk(gclk));
	jnot g06351(.din(n6604),.dout(n6605),.clk(gclk));
	jand g06352(.dina(n6605),.dinb(n6603),.dout(n6606),.clk(gclk));
	jnot g06353(.din(n6606),.dout(n6607),.clk(gclk));
	jor g06354(.dina(w_n6607_0[1]),.dinb(w_n6599_0[1]),.dout(n6608),.clk(gclk));
	jand g06355(.dina(n6608),.dinb(w_n6597_0[1]),.dout(n6609),.clk(gclk));
	jor g06356(.dina(w_n6609_0[1]),.dinb(w_n3371_20[1]),.dout(n6610),.clk(gclk));
	jxor g06357(.dina(w_n6216_0[0]),.dinb(w_n3376_23[0]),.dout(n6611),.clk(gclk));
	jor g06358(.dina(n6611),.dinb(w_n6505_25[1]),.dout(n6612),.clk(gclk));
	jxor g06359(.dina(n6612),.dinb(w_n6221_0[0]),.dout(n6613),.clk(gclk));
	jand g06360(.dina(w_n6609_0[0]),.dinb(w_n3371_20[0]),.dout(n6614),.clk(gclk));
	jor g06361(.dina(w_n6614_0[1]),.dinb(w_n6613_0[1]),.dout(n6615),.clk(gclk));
	jand g06362(.dina(w_n6615_0[2]),.dinb(w_n6610_0[2]),.dout(n6616),.clk(gclk));
	jor g06363(.dina(n6616),.dinb(w_n2875_23[1]),.dout(n6617),.clk(gclk));
	jnot g06364(.din(w_n6226_0[0]),.dout(n6618),.clk(gclk));
	jor g06365(.dina(n6618),.dinb(w_n6224_0[0]),.dout(n6619),.clk(gclk));
	jor g06366(.dina(n6619),.dinb(w_n6505_25[0]),.dout(n6620),.clk(gclk));
	jxor g06367(.dina(n6620),.dinb(w_n6235_0[0]),.dout(n6621),.clk(gclk));
	jand g06368(.dina(w_n6610_0[1]),.dinb(w_n2875_23[0]),.dout(n6622),.clk(gclk));
	jand g06369(.dina(n6622),.dinb(w_n6615_0[1]),.dout(n6623),.clk(gclk));
	jor g06370(.dina(w_n6623_0[1]),.dinb(w_n6621_0[1]),.dout(n6624),.clk(gclk));
	jand g06371(.dina(w_n6624_0[1]),.dinb(w_n6617_0[1]),.dout(n6625),.clk(gclk));
	jor g06372(.dina(w_n6625_0[2]),.dinb(w_n2870_20[2]),.dout(n6626),.clk(gclk));
	jand g06373(.dina(w_n6625_0[1]),.dinb(w_n2870_20[1]),.dout(n6627),.clk(gclk));
	jnot g06374(.din(w_n6238_0[0]),.dout(n6628),.clk(gclk));
	jand g06375(.dina(w_asqrt29_20[2]),.dinb(n6628),.dout(n6629),.clk(gclk));
	jand g06376(.dina(w_n6629_0[1]),.dinb(w_n6243_0[0]),.dout(n6630),.clk(gclk));
	jor g06377(.dina(n6630),.dinb(w_n6242_0[0]),.dout(n6631),.clk(gclk));
	jand g06378(.dina(w_n6629_0[0]),.dinb(w_n6244_0[0]),.dout(n6632),.clk(gclk));
	jnot g06379(.din(n6632),.dout(n6633),.clk(gclk));
	jand g06380(.dina(n6633),.dinb(n6631),.dout(n6634),.clk(gclk));
	jnot g06381(.din(n6634),.dout(n6635),.clk(gclk));
	jor g06382(.dina(w_n6635_0[1]),.dinb(n6627),.dout(n6636),.clk(gclk));
	jand g06383(.dina(w_n6636_0[1]),.dinb(w_n6626_0[1]),.dout(n6637),.clk(gclk));
	jor g06384(.dina(n6637),.dinb(w_n2425_24[0]),.dout(n6638),.clk(gclk));
	jand g06385(.dina(w_n6626_0[0]),.dinb(w_n2425_23[2]),.dout(n6639),.clk(gclk));
	jand g06386(.dina(n6639),.dinb(w_n6636_0[0]),.dout(n6640),.clk(gclk));
	jnot g06387(.din(w_n6246_0[0]),.dout(n6641),.clk(gclk));
	jand g06388(.dina(w_asqrt29_20[1]),.dinb(n6641),.dout(n6642),.clk(gclk));
	jand g06389(.dina(w_n6642_0[1]),.dinb(w_n6253_0[0]),.dout(n6643),.clk(gclk));
	jor g06390(.dina(n6643),.dinb(w_n6251_0[0]),.dout(n6644),.clk(gclk));
	jand g06391(.dina(w_n6642_0[0]),.dinb(w_n6254_0[0]),.dout(n6645),.clk(gclk));
	jnot g06392(.din(n6645),.dout(n6646),.clk(gclk));
	jand g06393(.dina(n6646),.dinb(n6644),.dout(n6647),.clk(gclk));
	jnot g06394(.din(n6647),.dout(n6648),.clk(gclk));
	jor g06395(.dina(w_n6648_0[1]),.dinb(w_n6640_0[1]),.dout(n6649),.clk(gclk));
	jand g06396(.dina(n6649),.dinb(w_n6638_0[1]),.dout(n6650),.clk(gclk));
	jor g06397(.dina(w_n6650_0[1]),.dinb(w_n2420_21[1]),.dout(n6651),.clk(gclk));
	jxor g06398(.dina(w_n6255_0[0]),.dinb(w_n2425_23[1]),.dout(n6652),.clk(gclk));
	jor g06399(.dina(n6652),.dinb(w_n6505_24[2]),.dout(n6653),.clk(gclk));
	jxor g06400(.dina(n6653),.dinb(w_n6266_0[0]),.dout(n6654),.clk(gclk));
	jand g06401(.dina(w_n6650_0[0]),.dinb(w_n2420_21[0]),.dout(n6655),.clk(gclk));
	jor g06402(.dina(w_n6655_0[1]),.dinb(w_n6654_0[1]),.dout(n6656),.clk(gclk));
	jand g06403(.dina(w_n6656_0[2]),.dinb(w_n6651_0[2]),.dout(n6657),.clk(gclk));
	jor g06404(.dina(n6657),.dinb(w_n2010_23[2]),.dout(n6658),.clk(gclk));
	jnot g06405(.din(w_n6271_0[0]),.dout(n6659),.clk(gclk));
	jor g06406(.dina(n6659),.dinb(w_n6269_0[0]),.dout(n6660),.clk(gclk));
	jor g06407(.dina(n6660),.dinb(w_n6505_24[1]),.dout(n6661),.clk(gclk));
	jxor g06408(.dina(n6661),.dinb(w_n6280_0[0]),.dout(n6662),.clk(gclk));
	jand g06409(.dina(w_n6651_0[1]),.dinb(w_n2010_23[1]),.dout(n6663),.clk(gclk));
	jand g06410(.dina(n6663),.dinb(w_n6656_0[1]),.dout(n6664),.clk(gclk));
	jor g06411(.dina(w_n6664_0[1]),.dinb(w_n6662_0[1]),.dout(n6665),.clk(gclk));
	jand g06412(.dina(w_n6665_0[1]),.dinb(w_n6658_0[1]),.dout(n6666),.clk(gclk));
	jor g06413(.dina(w_n6666_0[2]),.dinb(w_n2005_21[2]),.dout(n6667),.clk(gclk));
	jand g06414(.dina(w_n6666_0[1]),.dinb(w_n2005_21[1]),.dout(n6668),.clk(gclk));
	jnot g06415(.din(w_n6283_0[0]),.dout(n6669),.clk(gclk));
	jand g06416(.dina(w_asqrt29_20[0]),.dinb(n6669),.dout(n6670),.clk(gclk));
	jand g06417(.dina(w_n6670_0[1]),.dinb(w_n6288_0[0]),.dout(n6671),.clk(gclk));
	jor g06418(.dina(n6671),.dinb(w_n6287_0[0]),.dout(n6672),.clk(gclk));
	jand g06419(.dina(w_n6670_0[0]),.dinb(w_n6289_0[0]),.dout(n6673),.clk(gclk));
	jnot g06420(.din(n6673),.dout(n6674),.clk(gclk));
	jand g06421(.dina(n6674),.dinb(n6672),.dout(n6675),.clk(gclk));
	jnot g06422(.din(n6675),.dout(n6676),.clk(gclk));
	jor g06423(.dina(w_n6676_0[1]),.dinb(n6668),.dout(n6677),.clk(gclk));
	jand g06424(.dina(w_n6677_0[1]),.dinb(w_n6667_0[1]),.dout(n6678),.clk(gclk));
	jor g06425(.dina(n6678),.dinb(w_n1646_24[2]),.dout(n6679),.clk(gclk));
	jand g06426(.dina(w_n6667_0[0]),.dinb(w_n1646_24[1]),.dout(n6680),.clk(gclk));
	jand g06427(.dina(n6680),.dinb(w_n6677_0[0]),.dout(n6681),.clk(gclk));
	jnot g06428(.din(w_n6291_0[0]),.dout(n6682),.clk(gclk));
	jand g06429(.dina(w_asqrt29_19[2]),.dinb(n6682),.dout(n6683),.clk(gclk));
	jand g06430(.dina(w_n6683_0[1]),.dinb(w_n6298_0[0]),.dout(n6684),.clk(gclk));
	jor g06431(.dina(n6684),.dinb(w_n6296_0[0]),.dout(n6685),.clk(gclk));
	jand g06432(.dina(w_n6683_0[0]),.dinb(w_n6299_0[0]),.dout(n6686),.clk(gclk));
	jnot g06433(.din(n6686),.dout(n6687),.clk(gclk));
	jand g06434(.dina(n6687),.dinb(n6685),.dout(n6688),.clk(gclk));
	jnot g06435(.din(n6688),.dout(n6689),.clk(gclk));
	jor g06436(.dina(w_n6689_0[1]),.dinb(w_n6681_0[1]),.dout(n6690),.clk(gclk));
	jand g06437(.dina(n6690),.dinb(w_n6679_0[1]),.dout(n6691),.clk(gclk));
	jor g06438(.dina(w_n6691_0[1]),.dinb(w_n1641_22[0]),.dout(n6692),.clk(gclk));
	jxor g06439(.dina(w_n6300_0[0]),.dinb(w_n1646_24[0]),.dout(n6693),.clk(gclk));
	jor g06440(.dina(n6693),.dinb(w_n6505_24[0]),.dout(n6694),.clk(gclk));
	jxor g06441(.dina(n6694),.dinb(w_n6311_0[0]),.dout(n6695),.clk(gclk));
	jand g06442(.dina(w_n6691_0[0]),.dinb(w_n1641_21[2]),.dout(n6696),.clk(gclk));
	jor g06443(.dina(w_n6696_0[1]),.dinb(w_n6695_0[1]),.dout(n6697),.clk(gclk));
	jand g06444(.dina(w_n6697_0[2]),.dinb(w_n6692_0[2]),.dout(n6698),.clk(gclk));
	jor g06445(.dina(n6698),.dinb(w_n1317_24[1]),.dout(n6699),.clk(gclk));
	jnot g06446(.din(w_n6316_0[0]),.dout(n6700),.clk(gclk));
	jor g06447(.dina(n6700),.dinb(w_n6314_0[0]),.dout(n6701),.clk(gclk));
	jor g06448(.dina(n6701),.dinb(w_n6505_23[2]),.dout(n6702),.clk(gclk));
	jxor g06449(.dina(n6702),.dinb(w_n6325_0[0]),.dout(n6703),.clk(gclk));
	jand g06450(.dina(w_n6692_0[1]),.dinb(w_n1317_24[0]),.dout(n6704),.clk(gclk));
	jand g06451(.dina(n6704),.dinb(w_n6697_0[1]),.dout(n6705),.clk(gclk));
	jor g06452(.dina(w_n6705_0[1]),.dinb(w_n6703_0[1]),.dout(n6706),.clk(gclk));
	jand g06453(.dina(w_n6706_0[1]),.dinb(w_n6699_0[1]),.dout(n6707),.clk(gclk));
	jor g06454(.dina(w_n6707_0[2]),.dinb(w_n1312_22[1]),.dout(n6708),.clk(gclk));
	jand g06455(.dina(w_n6707_0[1]),.dinb(w_n1312_22[0]),.dout(n6709),.clk(gclk));
	jnot g06456(.din(w_n6328_0[0]),.dout(n6710),.clk(gclk));
	jand g06457(.dina(w_asqrt29_19[1]),.dinb(n6710),.dout(n6711),.clk(gclk));
	jand g06458(.dina(w_n6711_0[1]),.dinb(w_n6333_0[0]),.dout(n6712),.clk(gclk));
	jor g06459(.dina(n6712),.dinb(w_n6332_0[0]),.dout(n6713),.clk(gclk));
	jand g06460(.dina(w_n6711_0[0]),.dinb(w_n6334_0[0]),.dout(n6714),.clk(gclk));
	jnot g06461(.din(n6714),.dout(n6715),.clk(gclk));
	jand g06462(.dina(n6715),.dinb(n6713),.dout(n6716),.clk(gclk));
	jnot g06463(.din(n6716),.dout(n6717),.clk(gclk));
	jor g06464(.dina(w_n6717_0[1]),.dinb(n6709),.dout(n6718),.clk(gclk));
	jand g06465(.dina(w_n6718_0[1]),.dinb(w_n6708_0[1]),.dout(n6719),.clk(gclk));
	jor g06466(.dina(n6719),.dinb(w_n1039_25[0]),.dout(n6720),.clk(gclk));
	jand g06467(.dina(w_n6708_0[0]),.dinb(w_n1039_24[2]),.dout(n6721),.clk(gclk));
	jand g06468(.dina(n6721),.dinb(w_n6718_0[0]),.dout(n6722),.clk(gclk));
	jnot g06469(.din(w_n6336_0[0]),.dout(n6723),.clk(gclk));
	jand g06470(.dina(w_asqrt29_19[0]),.dinb(n6723),.dout(n6724),.clk(gclk));
	jand g06471(.dina(w_n6724_0[1]),.dinb(w_n6343_0[0]),.dout(n6725),.clk(gclk));
	jor g06472(.dina(n6725),.dinb(w_n6341_0[0]),.dout(n6726),.clk(gclk));
	jand g06473(.dina(w_n6724_0[0]),.dinb(w_n6344_0[0]),.dout(n6727),.clk(gclk));
	jnot g06474(.din(n6727),.dout(n6728),.clk(gclk));
	jand g06475(.dina(n6728),.dinb(n6726),.dout(n6729),.clk(gclk));
	jnot g06476(.din(n6729),.dout(n6730),.clk(gclk));
	jor g06477(.dina(w_n6730_0[1]),.dinb(w_n6722_0[1]),.dout(n6731),.clk(gclk));
	jand g06478(.dina(n6731),.dinb(w_n6720_0[1]),.dout(n6732),.clk(gclk));
	jor g06479(.dina(w_n6732_0[1]),.dinb(w_n1034_23[0]),.dout(n6733),.clk(gclk));
	jxor g06480(.dina(w_n6345_0[0]),.dinb(w_n1039_24[1]),.dout(n6734),.clk(gclk));
	jor g06481(.dina(n6734),.dinb(w_n6505_23[1]),.dout(n6735),.clk(gclk));
	jxor g06482(.dina(n6735),.dinb(w_n6356_0[0]),.dout(n6736),.clk(gclk));
	jand g06483(.dina(w_n6732_0[0]),.dinb(w_n1034_22[2]),.dout(n6737),.clk(gclk));
	jor g06484(.dina(w_n6737_0[1]),.dinb(w_n6736_0[1]),.dout(n6738),.clk(gclk));
	jand g06485(.dina(w_n6738_0[2]),.dinb(w_n6733_0[2]),.dout(n6739),.clk(gclk));
	jor g06486(.dina(n6739),.dinb(w_n796_24[2]),.dout(n6740),.clk(gclk));
	jnot g06487(.din(w_n6361_0[0]),.dout(n6741),.clk(gclk));
	jor g06488(.dina(n6741),.dinb(w_n6359_0[0]),.dout(n6742),.clk(gclk));
	jor g06489(.dina(n6742),.dinb(w_n6505_23[0]),.dout(n6743),.clk(gclk));
	jxor g06490(.dina(n6743),.dinb(w_n6370_0[0]),.dout(n6744),.clk(gclk));
	jand g06491(.dina(w_n6733_0[1]),.dinb(w_n796_24[1]),.dout(n6745),.clk(gclk));
	jand g06492(.dina(n6745),.dinb(w_n6738_0[1]),.dout(n6746),.clk(gclk));
	jor g06493(.dina(w_n6746_0[1]),.dinb(w_n6744_0[1]),.dout(n6747),.clk(gclk));
	jand g06494(.dina(w_n6747_0[1]),.dinb(w_n6740_0[1]),.dout(n6748),.clk(gclk));
	jor g06495(.dina(w_n6748_0[2]),.dinb(w_n791_23[1]),.dout(n6749),.clk(gclk));
	jand g06496(.dina(w_n6748_0[1]),.dinb(w_n791_23[0]),.dout(n6750),.clk(gclk));
	jnot g06497(.din(w_n6373_0[0]),.dout(n6751),.clk(gclk));
	jand g06498(.dina(w_asqrt29_18[2]),.dinb(n6751),.dout(n6752),.clk(gclk));
	jand g06499(.dina(w_n6752_0[1]),.dinb(w_n6378_0[0]),.dout(n6753),.clk(gclk));
	jor g06500(.dina(n6753),.dinb(w_n6377_0[0]),.dout(n6754),.clk(gclk));
	jand g06501(.dina(w_n6752_0[0]),.dinb(w_n6379_0[0]),.dout(n6755),.clk(gclk));
	jnot g06502(.din(n6755),.dout(n6756),.clk(gclk));
	jand g06503(.dina(n6756),.dinb(n6754),.dout(n6757),.clk(gclk));
	jnot g06504(.din(n6757),.dout(n6758),.clk(gclk));
	jor g06505(.dina(w_n6758_0[1]),.dinb(n6750),.dout(n6759),.clk(gclk));
	jand g06506(.dina(w_n6759_0[1]),.dinb(w_n6749_0[1]),.dout(n6760),.clk(gclk));
	jor g06507(.dina(n6760),.dinb(w_n595_25[1]),.dout(n6761),.clk(gclk));
	jand g06508(.dina(w_n6749_0[0]),.dinb(w_n595_25[0]),.dout(n6762),.clk(gclk));
	jand g06509(.dina(n6762),.dinb(w_n6759_0[0]),.dout(n6763),.clk(gclk));
	jnot g06510(.din(w_n6381_0[0]),.dout(n6764),.clk(gclk));
	jand g06511(.dina(w_asqrt29_18[1]),.dinb(n6764),.dout(n6765),.clk(gclk));
	jand g06512(.dina(w_n6765_0[1]),.dinb(w_n6388_0[0]),.dout(n6766),.clk(gclk));
	jor g06513(.dina(n6766),.dinb(w_n6386_0[0]),.dout(n6767),.clk(gclk));
	jand g06514(.dina(w_n6765_0[0]),.dinb(w_n6389_0[0]),.dout(n6768),.clk(gclk));
	jnot g06515(.din(n6768),.dout(n6769),.clk(gclk));
	jand g06516(.dina(n6769),.dinb(n6767),.dout(n6770),.clk(gclk));
	jnot g06517(.din(n6770),.dout(n6771),.clk(gclk));
	jor g06518(.dina(w_n6771_0[1]),.dinb(w_n6763_0[1]),.dout(n6772),.clk(gclk));
	jand g06519(.dina(n6772),.dinb(w_n6761_0[1]),.dout(n6773),.clk(gclk));
	jor g06520(.dina(w_n6773_0[1]),.dinb(w_n590_23[2]),.dout(n6774),.clk(gclk));
	jxor g06521(.dina(w_n6390_0[0]),.dinb(w_n595_24[2]),.dout(n6775),.clk(gclk));
	jor g06522(.dina(n6775),.dinb(w_n6505_22[2]),.dout(n6776),.clk(gclk));
	jxor g06523(.dina(n6776),.dinb(w_n6401_0[0]),.dout(n6777),.clk(gclk));
	jand g06524(.dina(w_n6773_0[0]),.dinb(w_n590_23[1]),.dout(n6778),.clk(gclk));
	jor g06525(.dina(w_n6778_0[1]),.dinb(w_n6777_0[1]),.dout(n6779),.clk(gclk));
	jand g06526(.dina(w_n6779_0[2]),.dinb(w_n6774_0[2]),.dout(n6780),.clk(gclk));
	jor g06527(.dina(n6780),.dinb(w_n430_25[0]),.dout(n6781),.clk(gclk));
	jnot g06528(.din(w_n6406_0[0]),.dout(n6782),.clk(gclk));
	jor g06529(.dina(n6782),.dinb(w_n6404_0[0]),.dout(n6783),.clk(gclk));
	jor g06530(.dina(n6783),.dinb(w_n6505_22[1]),.dout(n6784),.clk(gclk));
	jxor g06531(.dina(n6784),.dinb(w_n6415_0[0]),.dout(n6785),.clk(gclk));
	jand g06532(.dina(w_n6774_0[1]),.dinb(w_n430_24[2]),.dout(n6786),.clk(gclk));
	jand g06533(.dina(n6786),.dinb(w_n6779_0[1]),.dout(n6787),.clk(gclk));
	jor g06534(.dina(w_n6787_0[1]),.dinb(w_n6785_0[1]),.dout(n6788),.clk(gclk));
	jand g06535(.dina(w_n6788_0[1]),.dinb(w_n6781_0[1]),.dout(n6789),.clk(gclk));
	jor g06536(.dina(w_n6789_0[2]),.dinb(w_n425_24[0]),.dout(n6790),.clk(gclk));
	jand g06537(.dina(w_n6789_0[1]),.dinb(w_n425_23[2]),.dout(n6791),.clk(gclk));
	jnot g06538(.din(w_n6418_0[0]),.dout(n6792),.clk(gclk));
	jand g06539(.dina(w_asqrt29_18[0]),.dinb(n6792),.dout(n6793),.clk(gclk));
	jand g06540(.dina(w_n6793_0[1]),.dinb(w_n6423_0[0]),.dout(n6794),.clk(gclk));
	jor g06541(.dina(n6794),.dinb(w_n6422_0[0]),.dout(n6795),.clk(gclk));
	jand g06542(.dina(w_n6793_0[0]),.dinb(w_n6424_0[0]),.dout(n6796),.clk(gclk));
	jnot g06543(.din(n6796),.dout(n6797),.clk(gclk));
	jand g06544(.dina(n6797),.dinb(n6795),.dout(n6798),.clk(gclk));
	jnot g06545(.din(n6798),.dout(n6799),.clk(gclk));
	jor g06546(.dina(w_n6799_0[1]),.dinb(n6791),.dout(n6800),.clk(gclk));
	jand g06547(.dina(w_n6800_0[1]),.dinb(w_n6790_0[1]),.dout(n6801),.clk(gclk));
	jor g06548(.dina(n6801),.dinb(w_n305_25[2]),.dout(n6802),.clk(gclk));
	jand g06549(.dina(w_n6790_0[0]),.dinb(w_n305_25[1]),.dout(n6803),.clk(gclk));
	jand g06550(.dina(n6803),.dinb(w_n6800_0[0]),.dout(n6804),.clk(gclk));
	jnot g06551(.din(w_n6426_0[0]),.dout(n6805),.clk(gclk));
	jand g06552(.dina(w_asqrt29_17[2]),.dinb(n6805),.dout(n6806),.clk(gclk));
	jand g06553(.dina(w_n6806_0[1]),.dinb(w_n6433_0[0]),.dout(n6807),.clk(gclk));
	jor g06554(.dina(n6807),.dinb(w_n6431_0[0]),.dout(n6808),.clk(gclk));
	jand g06555(.dina(w_n6806_0[0]),.dinb(w_n6434_0[0]),.dout(n6809),.clk(gclk));
	jnot g06556(.din(n6809),.dout(n6810),.clk(gclk));
	jand g06557(.dina(n6810),.dinb(n6808),.dout(n6811),.clk(gclk));
	jnot g06558(.din(n6811),.dout(n6812),.clk(gclk));
	jor g06559(.dina(w_n6812_0[1]),.dinb(w_n6804_0[1]),.dout(n6813),.clk(gclk));
	jand g06560(.dina(n6813),.dinb(w_n6802_0[1]),.dout(n6814),.clk(gclk));
	jor g06561(.dina(w_n6814_0[1]),.dinb(w_n290_25[0]),.dout(n6815),.clk(gclk));
	jxor g06562(.dina(w_n6435_0[0]),.dinb(w_n305_25[0]),.dout(n6816),.clk(gclk));
	jor g06563(.dina(n6816),.dinb(w_n6505_22[0]),.dout(n6817),.clk(gclk));
	jxor g06564(.dina(n6817),.dinb(w_n6446_0[0]),.dout(n6818),.clk(gclk));
	jand g06565(.dina(w_n6814_0[0]),.dinb(w_n290_24[2]),.dout(n6819),.clk(gclk));
	jor g06566(.dina(w_n6819_0[1]),.dinb(w_n6818_0[1]),.dout(n6820),.clk(gclk));
	jand g06567(.dina(w_n6820_0[2]),.dinb(w_n6815_0[2]),.dout(n6821),.clk(gclk));
	jor g06568(.dina(n6821),.dinb(w_n223_25[1]),.dout(n6822),.clk(gclk));
	jnot g06569(.din(w_n6451_0[0]),.dout(n6823),.clk(gclk));
	jor g06570(.dina(n6823),.dinb(w_n6449_0[0]),.dout(n6824),.clk(gclk));
	jor g06571(.dina(n6824),.dinb(w_n6505_21[2]),.dout(n6825),.clk(gclk));
	jxor g06572(.dina(n6825),.dinb(w_n6460_0[0]),.dout(n6826),.clk(gclk));
	jand g06573(.dina(w_n6815_0[1]),.dinb(w_n223_25[0]),.dout(n6827),.clk(gclk));
	jand g06574(.dina(n6827),.dinb(w_n6820_0[1]),.dout(n6828),.clk(gclk));
	jor g06575(.dina(w_n6828_0[1]),.dinb(w_n6826_0[1]),.dout(n6829),.clk(gclk));
	jand g06576(.dina(w_n6829_0[1]),.dinb(w_n6822_0[1]),.dout(n6830),.clk(gclk));
	jor g06577(.dina(w_n6830_0[2]),.dinb(w_n199_29[1]),.dout(n6831),.clk(gclk));
	jand g06578(.dina(w_n6830_0[1]),.dinb(w_n199_29[0]),.dout(n6832),.clk(gclk));
	jnot g06579(.din(w_n6463_0[0]),.dout(n6833),.clk(gclk));
	jand g06580(.dina(w_asqrt29_17[1]),.dinb(n6833),.dout(n6834),.clk(gclk));
	jand g06581(.dina(w_n6834_0[1]),.dinb(w_n6468_0[0]),.dout(n6835),.clk(gclk));
	jor g06582(.dina(n6835),.dinb(w_n6467_0[0]),.dout(n6836),.clk(gclk));
	jand g06583(.dina(w_n6834_0[0]),.dinb(w_n6469_0[0]),.dout(n6837),.clk(gclk));
	jnot g06584(.din(n6837),.dout(n6838),.clk(gclk));
	jand g06585(.dina(n6838),.dinb(n6836),.dout(n6839),.clk(gclk));
	jnot g06586(.din(n6839),.dout(n6840),.clk(gclk));
	jor g06587(.dina(w_n6840_0[1]),.dinb(n6832),.dout(n6841),.clk(gclk));
	jand g06588(.dina(n6841),.dinb(n6831),.dout(n6842),.clk(gclk));
	jnot g06589(.din(w_n6471_0[0]),.dout(n6843),.clk(gclk));
	jand g06590(.dina(w_asqrt29_17[0]),.dinb(n6843),.dout(n6844),.clk(gclk));
	jand g06591(.dina(w_n6844_0[1]),.dinb(w_n6478_0[0]),.dout(n6845),.clk(gclk));
	jor g06592(.dina(n6845),.dinb(w_n6476_0[0]),.dout(n6846),.clk(gclk));
	jand g06593(.dina(w_n6844_0[0]),.dinb(w_n6479_0[0]),.dout(n6847),.clk(gclk));
	jnot g06594(.din(n6847),.dout(n6848),.clk(gclk));
	jand g06595(.dina(n6848),.dinb(n6846),.dout(n6849),.clk(gclk));
	jnot g06596(.din(w_n6849_0[2]),.dout(n6850),.clk(gclk));
	jand g06597(.dina(w_asqrt29_16[2]),.dinb(w_n6493_0[1]),.dout(n6851),.clk(gclk));
	jand g06598(.dina(w_n6851_0[1]),.dinb(w_n6480_1[0]),.dout(n6852),.clk(gclk));
	jor g06599(.dina(n6852),.dinb(w_n6527_0[0]),.dout(n6853),.clk(gclk));
	jor g06600(.dina(n6853),.dinb(w_n6850_0[1]),.dout(n6854),.clk(gclk));
	jor g06601(.dina(n6854),.dinb(w_n6842_0[2]),.dout(n6855),.clk(gclk));
	jand g06602(.dina(n6855),.dinb(w_n194_28[1]),.dout(n6856),.clk(gclk));
	jand g06603(.dina(w_n6850_0[0]),.dinb(w_n6842_0[1]),.dout(n6857),.clk(gclk));
	jor g06604(.dina(w_n6851_0[0]),.dinb(w_n6480_0[2]),.dout(n6858),.clk(gclk));
	jand g06605(.dina(w_n6493_0[0]),.dinb(w_n6480_0[1]),.dout(n6859),.clk(gclk));
	jor g06606(.dina(n6859),.dinb(w_n194_28[0]),.dout(n6860),.clk(gclk));
	jnot g06607(.din(n6860),.dout(n6861),.clk(gclk));
	jand g06608(.dina(n6861),.dinb(n6858),.dout(n6862),.clk(gclk));
	jor g06609(.dina(w_n6862_0[1]),.dinb(w_n6857_0[2]),.dout(n6865),.clk(gclk));
	jor g06610(.dina(n6865),.dinb(w_n6856_0[1]),.dout(asqrt_fa_29),.clk(gclk));
	jxor g06611(.dina(w_n6555_0[0]),.dinb(w_n5116_18[2]),.dout(n6867),.clk(gclk));
	jand g06612(.dina(n6867),.dinb(w_asqrt28_31),.dout(n6868),.clk(gclk));
	jxor g06613(.dina(n6868),.dinb(w_n6508_0[0]),.dout(n6869),.clk(gclk));
	jnot g06614(.din(w_n6869_0[1]),.dout(n6870),.clk(gclk));
	jand g06615(.dina(w_asqrt28_30[2]),.dinb(w_a56_0[0]),.dout(n6871),.clk(gclk));
	jnot g06616(.din(w_a54_0[1]),.dout(n6872),.clk(gclk));
	jnot g06617(.din(w_a55_0[1]),.dout(n6873),.clk(gclk));
	jand g06618(.dina(w_n6510_1[0]),.dinb(w_n6873_0[1]),.dout(n6874),.clk(gclk));
	jand g06619(.dina(n6874),.dinb(w_n6872_1[1]),.dout(n6875),.clk(gclk));
	jor g06620(.dina(n6875),.dinb(n6871),.dout(n6876),.clk(gclk));
	jand g06621(.dina(w_n6876_0[2]),.dinb(w_asqrt29_16[1]),.dout(n6877),.clk(gclk));
	jand g06622(.dina(w_asqrt28_30[1]),.dinb(w_n6510_0[2]),.dout(n6878),.clk(gclk));
	jxor g06623(.dina(w_n6878_0[1]),.dinb(w_n6511_0[1]),.dout(n6879),.clk(gclk));
	jor g06624(.dina(w_n6876_0[1]),.dinb(w_asqrt29_16[0]),.dout(n6880),.clk(gclk));
	jand g06625(.dina(n6880),.dinb(w_n6879_0[1]),.dout(n6881),.clk(gclk));
	jor g06626(.dina(w_n6881_0[1]),.dinb(w_n6877_0[1]),.dout(n6882),.clk(gclk));
	jand g06627(.dina(n6882),.dinb(w_asqrt30_19[1]),.dout(n6883),.clk(gclk));
	jor g06628(.dina(w_n6877_0[0]),.dinb(w_asqrt30_19[0]),.dout(n6884),.clk(gclk));
	jor g06629(.dina(n6884),.dinb(w_n6881_0[0]),.dout(n6885),.clk(gclk));
	jand g06630(.dina(w_n6878_0[0]),.dinb(w_n6511_0[0]),.dout(n6886),.clk(gclk));
	jnot g06631(.din(w_n6856_0[0]),.dout(n6887),.clk(gclk));
	jnot g06632(.din(w_n6857_0[1]),.dout(n6888),.clk(gclk));
	jnot g06633(.din(w_n6862_0[0]),.dout(n6889),.clk(gclk));
	jand g06634(.dina(n6889),.dinb(w_asqrt29_15[2]),.dout(n6890),.clk(gclk));
	jand g06635(.dina(n6890),.dinb(n6888),.dout(n6891),.clk(gclk));
	jand g06636(.dina(n6891),.dinb(n6887),.dout(n6892),.clk(gclk));
	jor g06637(.dina(n6892),.dinb(n6886),.dout(n6893),.clk(gclk));
	jxor g06638(.dina(n6893),.dinb(w_n6134_0[1]),.dout(n6894),.clk(gclk));
	jand g06639(.dina(w_n6894_0[1]),.dinb(w_n6885_0[1]),.dout(n6895),.clk(gclk));
	jor g06640(.dina(n6895),.dinb(w_n6883_0[1]),.dout(n6896),.clk(gclk));
	jand g06641(.dina(w_n6896_0[2]),.dinb(w_asqrt31_16[0]),.dout(n6897),.clk(gclk));
	jor g06642(.dina(w_n6896_0[1]),.dinb(w_asqrt31_15[2]),.dout(n6898),.clk(gclk));
	jxor g06643(.dina(w_n6515_0[0]),.dinb(w_n6500_18[1]),.dout(n6899),.clk(gclk));
	jand g06644(.dina(n6899),.dinb(w_asqrt28_30[0]),.dout(n6900),.clk(gclk));
	jxor g06645(.dina(n6900),.dinb(w_n6518_0[0]),.dout(n6901),.clk(gclk));
	jnot g06646(.din(w_n6901_0[1]),.dout(n6902),.clk(gclk));
	jand g06647(.dina(n6902),.dinb(n6898),.dout(n6903),.clk(gclk));
	jor g06648(.dina(w_n6903_0[1]),.dinb(w_n6897_0[1]),.dout(n6904),.clk(gclk));
	jand g06649(.dina(n6904),.dinb(w_asqrt32_19[1]),.dout(n6905),.clk(gclk));
	jnot g06650(.din(w_n6524_0[0]),.dout(n6906),.clk(gclk));
	jand g06651(.dina(n6906),.dinb(w_n6522_0[0]),.dout(n6907),.clk(gclk));
	jand g06652(.dina(n6907),.dinb(w_asqrt28_29[2]),.dout(n6908),.clk(gclk));
	jxor g06653(.dina(n6908),.dinb(w_n6532_0[0]),.dout(n6909),.clk(gclk));
	jnot g06654(.din(n6909),.dout(n6910),.clk(gclk));
	jor g06655(.dina(w_n6897_0[0]),.dinb(w_asqrt32_19[0]),.dout(n6911),.clk(gclk));
	jor g06656(.dina(n6911),.dinb(w_n6903_0[0]),.dout(n6912),.clk(gclk));
	jand g06657(.dina(w_n6912_0[1]),.dinb(w_n6910_0[1]),.dout(n6913),.clk(gclk));
	jor g06658(.dina(w_n6913_0[1]),.dinb(w_n6905_0[1]),.dout(n6914),.clk(gclk));
	jand g06659(.dina(w_n6914_0[2]),.dinb(w_asqrt33_16[1]),.dout(n6915),.clk(gclk));
	jor g06660(.dina(w_n6914_0[1]),.dinb(w_asqrt33_16[0]),.dout(n6916),.clk(gclk));
	jnot g06661(.din(w_n6539_0[0]),.dout(n6917),.clk(gclk));
	jxor g06662(.dina(w_n6534_0[0]),.dinb(w_n5788_18[2]),.dout(n6918),.clk(gclk));
	jand g06663(.dina(n6918),.dinb(w_asqrt28_29[1]),.dout(n6919),.clk(gclk));
	jxor g06664(.dina(n6919),.dinb(n6917),.dout(n6920),.clk(gclk));
	jand g06665(.dina(w_n6920_0[1]),.dinb(n6916),.dout(n6921),.clk(gclk));
	jor g06666(.dina(w_n6921_0[1]),.dinb(w_n6915_0[1]),.dout(n6922),.clk(gclk));
	jand g06667(.dina(n6922),.dinb(w_asqrt34_19[1]),.dout(n6923),.clk(gclk));
	jnot g06668(.din(w_n6544_0[0]),.dout(n6924),.clk(gclk));
	jand g06669(.dina(n6924),.dinb(w_n6542_0[0]),.dout(n6925),.clk(gclk));
	jand g06670(.dina(n6925),.dinb(w_asqrt28_29[0]),.dout(n6926),.clk(gclk));
	jxor g06671(.dina(n6926),.dinb(w_n6553_0[0]),.dout(n6927),.clk(gclk));
	jnot g06672(.din(n6927),.dout(n6928),.clk(gclk));
	jor g06673(.dina(w_n6915_0[0]),.dinb(w_asqrt34_19[0]),.dout(n6929),.clk(gclk));
	jor g06674(.dina(n6929),.dinb(w_n6921_0[0]),.dout(n6930),.clk(gclk));
	jand g06675(.dina(w_n6930_0[1]),.dinb(w_n6928_0[1]),.dout(n6931),.clk(gclk));
	jor g06676(.dina(w_n6931_0[1]),.dinb(w_n6923_0[1]),.dout(n6932),.clk(gclk));
	jand g06677(.dina(w_n6932_0[2]),.dinb(w_asqrt35_16[1]),.dout(n6933),.clk(gclk));
	jor g06678(.dina(w_n6932_0[1]),.dinb(w_asqrt35_16[0]),.dout(n6934),.clk(gclk));
	jand g06679(.dina(n6934),.dinb(w_n6869_0[0]),.dout(n6935),.clk(gclk));
	jor g06680(.dina(w_n6935_0[1]),.dinb(w_n6933_0[1]),.dout(n6936),.clk(gclk));
	jand g06681(.dina(n6936),.dinb(w_asqrt36_19[1]),.dout(n6937),.clk(gclk));
	jor g06682(.dina(w_n6933_0[0]),.dinb(w_asqrt36_19[0]),.dout(n6938),.clk(gclk));
	jor g06683(.dina(n6938),.dinb(w_n6935_0[0]),.dout(n6939),.clk(gclk));
	jnot g06684(.din(w_n6565_0[0]),.dout(n6940),.clk(gclk));
	jnot g06685(.din(w_n6567_0[0]),.dout(n6941),.clk(gclk));
	jand g06686(.dina(w_asqrt28_28[2]),.dinb(w_n6561_0[0]),.dout(n6942),.clk(gclk));
	jand g06687(.dina(w_n6942_0[1]),.dinb(n6941),.dout(n6943),.clk(gclk));
	jor g06688(.dina(n6943),.dinb(n6940),.dout(n6944),.clk(gclk));
	jnot g06689(.din(w_n6568_0[0]),.dout(n6945),.clk(gclk));
	jand g06690(.dina(w_n6942_0[0]),.dinb(n6945),.dout(n6946),.clk(gclk));
	jnot g06691(.din(n6946),.dout(n6947),.clk(gclk));
	jand g06692(.dina(n6947),.dinb(n6944),.dout(n6948),.clk(gclk));
	jand g06693(.dina(w_n6948_0[1]),.dinb(w_n6939_0[1]),.dout(n6949),.clk(gclk));
	jor g06694(.dina(n6949),.dinb(w_n6937_0[1]),.dout(n6950),.clk(gclk));
	jand g06695(.dina(w_n6950_0[2]),.dinb(w_asqrt37_16[2]),.dout(n6951),.clk(gclk));
	jor g06696(.dina(w_n6950_0[1]),.dinb(w_asqrt37_16[1]),.dout(n6952),.clk(gclk));
	jxor g06697(.dina(w_n6569_0[0]),.dinb(w_n4494_19[1]),.dout(n6953),.clk(gclk));
	jand g06698(.dina(n6953),.dinb(w_asqrt28_28[1]),.dout(n6954),.clk(gclk));
	jxor g06699(.dina(n6954),.dinb(w_n6575_0[0]),.dout(n6955),.clk(gclk));
	jand g06700(.dina(w_n6955_0[1]),.dinb(n6952),.dout(n6956),.clk(gclk));
	jor g06701(.dina(w_n6956_0[1]),.dinb(w_n6951_0[1]),.dout(n6957),.clk(gclk));
	jand g06702(.dina(n6957),.dinb(w_asqrt38_19[1]),.dout(n6958),.clk(gclk));
	jor g06703(.dina(w_n6951_0[0]),.dinb(w_asqrt38_19[0]),.dout(n6959),.clk(gclk));
	jor g06704(.dina(n6959),.dinb(w_n6956_0[0]),.dout(n6960),.clk(gclk));
	jnot g06705(.din(w_n6583_0[0]),.dout(n6961),.clk(gclk));
	jnot g06706(.din(w_n6585_0[0]),.dout(n6962),.clk(gclk));
	jand g06707(.dina(w_asqrt28_28[0]),.dinb(w_n6579_0[0]),.dout(n6963),.clk(gclk));
	jand g06708(.dina(w_n6963_0[1]),.dinb(n6962),.dout(n6964),.clk(gclk));
	jor g06709(.dina(n6964),.dinb(n6961),.dout(n6965),.clk(gclk));
	jnot g06710(.din(w_n6586_0[0]),.dout(n6966),.clk(gclk));
	jand g06711(.dina(w_n6963_0[0]),.dinb(n6966),.dout(n6967),.clk(gclk));
	jnot g06712(.din(n6967),.dout(n6968),.clk(gclk));
	jand g06713(.dina(n6968),.dinb(n6965),.dout(n6969),.clk(gclk));
	jand g06714(.dina(w_n6969_0[1]),.dinb(w_n6960_0[1]),.dout(n6970),.clk(gclk));
	jor g06715(.dina(n6970),.dinb(w_n6958_0[1]),.dout(n6971),.clk(gclk));
	jand g06716(.dina(w_n6971_0[1]),.dinb(w_asqrt39_16[2]),.dout(n6972),.clk(gclk));
	jxor g06717(.dina(w_n6587_0[0]),.dinb(w_n3907_19[1]),.dout(n6973),.clk(gclk));
	jand g06718(.dina(n6973),.dinb(w_asqrt28_27[2]),.dout(n6974),.clk(gclk));
	jxor g06719(.dina(n6974),.dinb(w_n6594_0[0]),.dout(n6975),.clk(gclk));
	jnot g06720(.din(n6975),.dout(n6976),.clk(gclk));
	jor g06721(.dina(w_n6971_0[0]),.dinb(w_asqrt39_16[1]),.dout(n6977),.clk(gclk));
	jand g06722(.dina(w_n6977_0[1]),.dinb(w_n6976_0[1]),.dout(n6978),.clk(gclk));
	jor g06723(.dina(w_n6978_0[2]),.dinb(w_n6972_0[2]),.dout(n6979),.clk(gclk));
	jand g06724(.dina(n6979),.dinb(w_asqrt40_19[1]),.dout(n6980),.clk(gclk));
	jnot g06725(.din(w_n6599_0[0]),.dout(n6981),.clk(gclk));
	jand g06726(.dina(n6981),.dinb(w_n6597_0[0]),.dout(n6982),.clk(gclk));
	jand g06727(.dina(n6982),.dinb(w_asqrt28_27[1]),.dout(n6983),.clk(gclk));
	jxor g06728(.dina(n6983),.dinb(w_n6607_0[0]),.dout(n6984),.clk(gclk));
	jnot g06729(.din(n6984),.dout(n6985),.clk(gclk));
	jor g06730(.dina(w_n6972_0[1]),.dinb(w_asqrt40_19[0]),.dout(n6986),.clk(gclk));
	jor g06731(.dina(n6986),.dinb(w_n6978_0[1]),.dout(n6987),.clk(gclk));
	jand g06732(.dina(w_n6987_0[1]),.dinb(w_n6985_0[1]),.dout(n6988),.clk(gclk));
	jor g06733(.dina(w_n6988_0[1]),.dinb(w_n6980_0[1]),.dout(n6989),.clk(gclk));
	jand g06734(.dina(w_n6989_0[2]),.dinb(w_asqrt41_17[0]),.dout(n6990),.clk(gclk));
	jor g06735(.dina(w_n6989_0[1]),.dinb(w_asqrt41_16[2]),.dout(n6991),.clk(gclk));
	jnot g06736(.din(w_n6613_0[0]),.dout(n6992),.clk(gclk));
	jnot g06737(.din(w_n6614_0[0]),.dout(n6993),.clk(gclk));
	jand g06738(.dina(w_asqrt28_27[0]),.dinb(w_n6610_0[0]),.dout(n6994),.clk(gclk));
	jand g06739(.dina(w_n6994_0[1]),.dinb(n6993),.dout(n6995),.clk(gclk));
	jor g06740(.dina(n6995),.dinb(n6992),.dout(n6996),.clk(gclk));
	jnot g06741(.din(w_n6615_0[0]),.dout(n6997),.clk(gclk));
	jand g06742(.dina(w_n6994_0[0]),.dinb(n6997),.dout(n6998),.clk(gclk));
	jnot g06743(.din(n6998),.dout(n6999),.clk(gclk));
	jand g06744(.dina(n6999),.dinb(n6996),.dout(n7000),.clk(gclk));
	jand g06745(.dina(w_n7000_0[1]),.dinb(n6991),.dout(n7001),.clk(gclk));
	jor g06746(.dina(w_n7001_0[1]),.dinb(w_n6990_0[1]),.dout(n7002),.clk(gclk));
	jand g06747(.dina(n7002),.dinb(w_asqrt42_19[1]),.dout(n7003),.clk(gclk));
	jor g06748(.dina(w_n6990_0[0]),.dinb(w_asqrt42_19[0]),.dout(n7004),.clk(gclk));
	jor g06749(.dina(n7004),.dinb(w_n7001_0[0]),.dout(n7005),.clk(gclk));
	jnot g06750(.din(w_n6621_0[0]),.dout(n7006),.clk(gclk));
	jnot g06751(.din(w_n6623_0[0]),.dout(n7007),.clk(gclk));
	jand g06752(.dina(w_asqrt28_26[2]),.dinb(w_n6617_0[0]),.dout(n7008),.clk(gclk));
	jand g06753(.dina(w_n7008_0[1]),.dinb(n7007),.dout(n7009),.clk(gclk));
	jor g06754(.dina(n7009),.dinb(n7006),.dout(n7010),.clk(gclk));
	jnot g06755(.din(w_n6624_0[0]),.dout(n7011),.clk(gclk));
	jand g06756(.dina(w_n7008_0[0]),.dinb(n7011),.dout(n7012),.clk(gclk));
	jnot g06757(.din(n7012),.dout(n7013),.clk(gclk));
	jand g06758(.dina(n7013),.dinb(n7010),.dout(n7014),.clk(gclk));
	jand g06759(.dina(w_n7014_0[1]),.dinb(w_n7005_0[1]),.dout(n7015),.clk(gclk));
	jor g06760(.dina(n7015),.dinb(w_n7003_0[1]),.dout(n7016),.clk(gclk));
	jand g06761(.dina(w_n7016_0[1]),.dinb(w_asqrt43_17[0]),.dout(n7017),.clk(gclk));
	jxor g06762(.dina(w_n6625_0[0]),.dinb(w_n2870_20[0]),.dout(n7018),.clk(gclk));
	jand g06763(.dina(n7018),.dinb(w_asqrt28_26[1]),.dout(n7019),.clk(gclk));
	jxor g06764(.dina(n7019),.dinb(w_n6635_0[0]),.dout(n7020),.clk(gclk));
	jnot g06765(.din(n7020),.dout(n7021),.clk(gclk));
	jor g06766(.dina(w_n7016_0[0]),.dinb(w_asqrt43_16[2]),.dout(n7022),.clk(gclk));
	jand g06767(.dina(w_n7022_0[1]),.dinb(w_n7021_0[1]),.dout(n7023),.clk(gclk));
	jor g06768(.dina(w_n7023_0[2]),.dinb(w_n7017_0[2]),.dout(n7024),.clk(gclk));
	jand g06769(.dina(n7024),.dinb(w_asqrt44_19[1]),.dout(n7025),.clk(gclk));
	jnot g06770(.din(w_n6640_0[0]),.dout(n7026),.clk(gclk));
	jand g06771(.dina(n7026),.dinb(w_n6638_0[0]),.dout(n7027),.clk(gclk));
	jand g06772(.dina(n7027),.dinb(w_asqrt28_26[0]),.dout(n7028),.clk(gclk));
	jxor g06773(.dina(n7028),.dinb(w_n6648_0[0]),.dout(n7029),.clk(gclk));
	jnot g06774(.din(n7029),.dout(n7030),.clk(gclk));
	jor g06775(.dina(w_n7017_0[1]),.dinb(w_asqrt44_19[0]),.dout(n7031),.clk(gclk));
	jor g06776(.dina(n7031),.dinb(w_n7023_0[1]),.dout(n7032),.clk(gclk));
	jand g06777(.dina(w_n7032_0[1]),.dinb(w_n7030_0[1]),.dout(n7033),.clk(gclk));
	jor g06778(.dina(w_n7033_0[1]),.dinb(w_n7025_0[1]),.dout(n7034),.clk(gclk));
	jand g06779(.dina(w_n7034_0[2]),.dinb(w_asqrt45_17[1]),.dout(n7035),.clk(gclk));
	jor g06780(.dina(w_n7034_0[1]),.dinb(w_asqrt45_17[0]),.dout(n7036),.clk(gclk));
	jnot g06781(.din(w_n6654_0[0]),.dout(n7037),.clk(gclk));
	jnot g06782(.din(w_n6655_0[0]),.dout(n7038),.clk(gclk));
	jand g06783(.dina(w_asqrt28_25[2]),.dinb(w_n6651_0[0]),.dout(n7039),.clk(gclk));
	jand g06784(.dina(w_n7039_0[1]),.dinb(n7038),.dout(n7040),.clk(gclk));
	jor g06785(.dina(n7040),.dinb(n7037),.dout(n7041),.clk(gclk));
	jnot g06786(.din(w_n6656_0[0]),.dout(n7042),.clk(gclk));
	jand g06787(.dina(w_n7039_0[0]),.dinb(n7042),.dout(n7043),.clk(gclk));
	jnot g06788(.din(n7043),.dout(n7044),.clk(gclk));
	jand g06789(.dina(n7044),.dinb(n7041),.dout(n7045),.clk(gclk));
	jand g06790(.dina(w_n7045_0[1]),.dinb(n7036),.dout(n7046),.clk(gclk));
	jor g06791(.dina(w_n7046_0[1]),.dinb(w_n7035_0[1]),.dout(n7047),.clk(gclk));
	jand g06792(.dina(n7047),.dinb(w_asqrt46_19[1]),.dout(n7048),.clk(gclk));
	jor g06793(.dina(w_n7035_0[0]),.dinb(w_asqrt46_19[0]),.dout(n7049),.clk(gclk));
	jor g06794(.dina(n7049),.dinb(w_n7046_0[0]),.dout(n7050),.clk(gclk));
	jnot g06795(.din(w_n6662_0[0]),.dout(n7051),.clk(gclk));
	jnot g06796(.din(w_n6664_0[0]),.dout(n7052),.clk(gclk));
	jand g06797(.dina(w_asqrt28_25[1]),.dinb(w_n6658_0[0]),.dout(n7053),.clk(gclk));
	jand g06798(.dina(w_n7053_0[1]),.dinb(n7052),.dout(n7054),.clk(gclk));
	jor g06799(.dina(n7054),.dinb(n7051),.dout(n7055),.clk(gclk));
	jnot g06800(.din(w_n6665_0[0]),.dout(n7056),.clk(gclk));
	jand g06801(.dina(w_n7053_0[0]),.dinb(n7056),.dout(n7057),.clk(gclk));
	jnot g06802(.din(n7057),.dout(n7058),.clk(gclk));
	jand g06803(.dina(n7058),.dinb(n7055),.dout(n7059),.clk(gclk));
	jand g06804(.dina(w_n7059_0[1]),.dinb(w_n7050_0[1]),.dout(n7060),.clk(gclk));
	jor g06805(.dina(n7060),.dinb(w_n7048_0[1]),.dout(n7061),.clk(gclk));
	jand g06806(.dina(w_n7061_0[1]),.dinb(w_asqrt47_17[1]),.dout(n7062),.clk(gclk));
	jxor g06807(.dina(w_n6666_0[0]),.dinb(w_n2005_21[0]),.dout(n7063),.clk(gclk));
	jand g06808(.dina(n7063),.dinb(w_asqrt28_25[0]),.dout(n7064),.clk(gclk));
	jxor g06809(.dina(n7064),.dinb(w_n6676_0[0]),.dout(n7065),.clk(gclk));
	jnot g06810(.din(n7065),.dout(n7066),.clk(gclk));
	jor g06811(.dina(w_n7061_0[0]),.dinb(w_asqrt47_17[0]),.dout(n7067),.clk(gclk));
	jand g06812(.dina(w_n7067_0[1]),.dinb(w_n7066_0[1]),.dout(n7068),.clk(gclk));
	jor g06813(.dina(w_n7068_0[2]),.dinb(w_n7062_0[2]),.dout(n7069),.clk(gclk));
	jand g06814(.dina(n7069),.dinb(w_asqrt48_19[1]),.dout(n7070),.clk(gclk));
	jnot g06815(.din(w_n6681_0[0]),.dout(n7071),.clk(gclk));
	jand g06816(.dina(n7071),.dinb(w_n6679_0[0]),.dout(n7072),.clk(gclk));
	jand g06817(.dina(n7072),.dinb(w_asqrt28_24[2]),.dout(n7073),.clk(gclk));
	jxor g06818(.dina(n7073),.dinb(w_n6689_0[0]),.dout(n7074),.clk(gclk));
	jnot g06819(.din(n7074),.dout(n7075),.clk(gclk));
	jor g06820(.dina(w_n7062_0[1]),.dinb(w_asqrt48_19[0]),.dout(n7076),.clk(gclk));
	jor g06821(.dina(n7076),.dinb(w_n7068_0[1]),.dout(n7077),.clk(gclk));
	jand g06822(.dina(w_n7077_0[1]),.dinb(w_n7075_0[1]),.dout(n7078),.clk(gclk));
	jor g06823(.dina(w_n7078_0[1]),.dinb(w_n7070_0[1]),.dout(n7079),.clk(gclk));
	jand g06824(.dina(w_n7079_0[2]),.dinb(w_asqrt49_17[2]),.dout(n7080),.clk(gclk));
	jor g06825(.dina(w_n7079_0[1]),.dinb(w_asqrt49_17[1]),.dout(n7081),.clk(gclk));
	jnot g06826(.din(w_n6695_0[0]),.dout(n7082),.clk(gclk));
	jnot g06827(.din(w_n6696_0[0]),.dout(n7083),.clk(gclk));
	jand g06828(.dina(w_asqrt28_24[1]),.dinb(w_n6692_0[0]),.dout(n7084),.clk(gclk));
	jand g06829(.dina(w_n7084_0[1]),.dinb(n7083),.dout(n7085),.clk(gclk));
	jor g06830(.dina(n7085),.dinb(n7082),.dout(n7086),.clk(gclk));
	jnot g06831(.din(w_n6697_0[0]),.dout(n7087),.clk(gclk));
	jand g06832(.dina(w_n7084_0[0]),.dinb(n7087),.dout(n7088),.clk(gclk));
	jnot g06833(.din(n7088),.dout(n7089),.clk(gclk));
	jand g06834(.dina(n7089),.dinb(n7086),.dout(n7090),.clk(gclk));
	jand g06835(.dina(w_n7090_0[1]),.dinb(n7081),.dout(n7091),.clk(gclk));
	jor g06836(.dina(w_n7091_0[1]),.dinb(w_n7080_0[1]),.dout(n7092),.clk(gclk));
	jand g06837(.dina(n7092),.dinb(w_asqrt50_19[1]),.dout(n7093),.clk(gclk));
	jor g06838(.dina(w_n7080_0[0]),.dinb(w_asqrt50_19[0]),.dout(n7094),.clk(gclk));
	jor g06839(.dina(n7094),.dinb(w_n7091_0[0]),.dout(n7095),.clk(gclk));
	jnot g06840(.din(w_n6703_0[0]),.dout(n7096),.clk(gclk));
	jnot g06841(.din(w_n6705_0[0]),.dout(n7097),.clk(gclk));
	jand g06842(.dina(w_asqrt28_24[0]),.dinb(w_n6699_0[0]),.dout(n7098),.clk(gclk));
	jand g06843(.dina(w_n7098_0[1]),.dinb(n7097),.dout(n7099),.clk(gclk));
	jor g06844(.dina(n7099),.dinb(n7096),.dout(n7100),.clk(gclk));
	jnot g06845(.din(w_n6706_0[0]),.dout(n7101),.clk(gclk));
	jand g06846(.dina(w_n7098_0[0]),.dinb(n7101),.dout(n7102),.clk(gclk));
	jnot g06847(.din(n7102),.dout(n7103),.clk(gclk));
	jand g06848(.dina(n7103),.dinb(n7100),.dout(n7104),.clk(gclk));
	jand g06849(.dina(w_n7104_0[1]),.dinb(w_n7095_0[1]),.dout(n7105),.clk(gclk));
	jor g06850(.dina(n7105),.dinb(w_n7093_0[1]),.dout(n7106),.clk(gclk));
	jand g06851(.dina(w_n7106_0[1]),.dinb(w_asqrt51_17[2]),.dout(n7107),.clk(gclk));
	jxor g06852(.dina(w_n6707_0[0]),.dinb(w_n1312_21[2]),.dout(n7108),.clk(gclk));
	jand g06853(.dina(n7108),.dinb(w_asqrt28_23[2]),.dout(n7109),.clk(gclk));
	jxor g06854(.dina(n7109),.dinb(w_n6717_0[0]),.dout(n7110),.clk(gclk));
	jnot g06855(.din(n7110),.dout(n7111),.clk(gclk));
	jor g06856(.dina(w_n7106_0[0]),.dinb(w_asqrt51_17[1]),.dout(n7112),.clk(gclk));
	jand g06857(.dina(w_n7112_0[1]),.dinb(w_n7111_0[1]),.dout(n7113),.clk(gclk));
	jor g06858(.dina(w_n7113_0[2]),.dinb(w_n7107_0[2]),.dout(n7114),.clk(gclk));
	jand g06859(.dina(n7114),.dinb(w_asqrt52_19[1]),.dout(n7115),.clk(gclk));
	jnot g06860(.din(w_n6722_0[0]),.dout(n7116),.clk(gclk));
	jand g06861(.dina(n7116),.dinb(w_n6720_0[0]),.dout(n7117),.clk(gclk));
	jand g06862(.dina(n7117),.dinb(w_asqrt28_23[1]),.dout(n7118),.clk(gclk));
	jxor g06863(.dina(n7118),.dinb(w_n6730_0[0]),.dout(n7119),.clk(gclk));
	jnot g06864(.din(n7119),.dout(n7120),.clk(gclk));
	jor g06865(.dina(w_n7107_0[1]),.dinb(w_asqrt52_19[0]),.dout(n7121),.clk(gclk));
	jor g06866(.dina(n7121),.dinb(w_n7113_0[1]),.dout(n7122),.clk(gclk));
	jand g06867(.dina(w_n7122_0[1]),.dinb(w_n7120_0[1]),.dout(n7123),.clk(gclk));
	jor g06868(.dina(w_n7123_0[1]),.dinb(w_n7115_0[1]),.dout(n7124),.clk(gclk));
	jand g06869(.dina(w_n7124_0[2]),.dinb(w_asqrt53_18[0]),.dout(n7125),.clk(gclk));
	jor g06870(.dina(w_n7124_0[1]),.dinb(w_asqrt53_17[2]),.dout(n7126),.clk(gclk));
	jnot g06871(.din(w_n6736_0[0]),.dout(n7127),.clk(gclk));
	jnot g06872(.din(w_n6737_0[0]),.dout(n7128),.clk(gclk));
	jand g06873(.dina(w_asqrt28_23[0]),.dinb(w_n6733_0[0]),.dout(n7129),.clk(gclk));
	jand g06874(.dina(w_n7129_0[1]),.dinb(n7128),.dout(n7130),.clk(gclk));
	jor g06875(.dina(n7130),.dinb(n7127),.dout(n7131),.clk(gclk));
	jnot g06876(.din(w_n6738_0[0]),.dout(n7132),.clk(gclk));
	jand g06877(.dina(w_n7129_0[0]),.dinb(n7132),.dout(n7133),.clk(gclk));
	jnot g06878(.din(n7133),.dout(n7134),.clk(gclk));
	jand g06879(.dina(n7134),.dinb(n7131),.dout(n7135),.clk(gclk));
	jand g06880(.dina(w_n7135_0[1]),.dinb(n7126),.dout(n7136),.clk(gclk));
	jor g06881(.dina(w_n7136_0[1]),.dinb(w_n7125_0[1]),.dout(n7137),.clk(gclk));
	jand g06882(.dina(n7137),.dinb(w_asqrt54_19[1]),.dout(n7138),.clk(gclk));
	jor g06883(.dina(w_n7125_0[0]),.dinb(w_asqrt54_19[0]),.dout(n7139),.clk(gclk));
	jor g06884(.dina(n7139),.dinb(w_n7136_0[0]),.dout(n7140),.clk(gclk));
	jnot g06885(.din(w_n6744_0[0]),.dout(n7141),.clk(gclk));
	jnot g06886(.din(w_n6746_0[0]),.dout(n7142),.clk(gclk));
	jand g06887(.dina(w_asqrt28_22[2]),.dinb(w_n6740_0[0]),.dout(n7143),.clk(gclk));
	jand g06888(.dina(w_n7143_0[1]),.dinb(n7142),.dout(n7144),.clk(gclk));
	jor g06889(.dina(n7144),.dinb(n7141),.dout(n7145),.clk(gclk));
	jnot g06890(.din(w_n6747_0[0]),.dout(n7146),.clk(gclk));
	jand g06891(.dina(w_n7143_0[0]),.dinb(n7146),.dout(n7147),.clk(gclk));
	jnot g06892(.din(n7147),.dout(n7148),.clk(gclk));
	jand g06893(.dina(n7148),.dinb(n7145),.dout(n7149),.clk(gclk));
	jand g06894(.dina(w_n7149_0[1]),.dinb(w_n7140_0[1]),.dout(n7150),.clk(gclk));
	jor g06895(.dina(n7150),.dinb(w_n7138_0[1]),.dout(n7151),.clk(gclk));
	jand g06896(.dina(w_n7151_0[1]),.dinb(w_asqrt55_18[1]),.dout(n7152),.clk(gclk));
	jxor g06897(.dina(w_n6748_0[0]),.dinb(w_n791_22[2]),.dout(n7153),.clk(gclk));
	jand g06898(.dina(n7153),.dinb(w_asqrt28_22[1]),.dout(n7154),.clk(gclk));
	jxor g06899(.dina(n7154),.dinb(w_n6758_0[0]),.dout(n7155),.clk(gclk));
	jnot g06900(.din(n7155),.dout(n7156),.clk(gclk));
	jor g06901(.dina(w_n7151_0[0]),.dinb(w_asqrt55_18[0]),.dout(n7157),.clk(gclk));
	jand g06902(.dina(w_n7157_0[1]),.dinb(w_n7156_0[1]),.dout(n7158),.clk(gclk));
	jor g06903(.dina(w_n7158_0[2]),.dinb(w_n7152_0[2]),.dout(n7159),.clk(gclk));
	jand g06904(.dina(n7159),.dinb(w_asqrt56_19[1]),.dout(n7160),.clk(gclk));
	jnot g06905(.din(w_n6763_0[0]),.dout(n7161),.clk(gclk));
	jand g06906(.dina(n7161),.dinb(w_n6761_0[0]),.dout(n7162),.clk(gclk));
	jand g06907(.dina(n7162),.dinb(w_asqrt28_22[0]),.dout(n7163),.clk(gclk));
	jxor g06908(.dina(n7163),.dinb(w_n6771_0[0]),.dout(n7164),.clk(gclk));
	jnot g06909(.din(n7164),.dout(n7165),.clk(gclk));
	jor g06910(.dina(w_n7152_0[1]),.dinb(w_asqrt56_19[0]),.dout(n7166),.clk(gclk));
	jor g06911(.dina(n7166),.dinb(w_n7158_0[1]),.dout(n7167),.clk(gclk));
	jand g06912(.dina(w_n7167_0[1]),.dinb(w_n7165_0[1]),.dout(n7168),.clk(gclk));
	jor g06913(.dina(w_n7168_0[1]),.dinb(w_n7160_0[1]),.dout(n7169),.clk(gclk));
	jand g06914(.dina(w_n7169_0[2]),.dinb(w_asqrt57_18[2]),.dout(n7170),.clk(gclk));
	jor g06915(.dina(w_n7169_0[1]),.dinb(w_asqrt57_18[1]),.dout(n7171),.clk(gclk));
	jnot g06916(.din(w_n6777_0[0]),.dout(n7172),.clk(gclk));
	jnot g06917(.din(w_n6778_0[0]),.dout(n7173),.clk(gclk));
	jand g06918(.dina(w_asqrt28_21[2]),.dinb(w_n6774_0[0]),.dout(n7174),.clk(gclk));
	jand g06919(.dina(w_n7174_0[1]),.dinb(n7173),.dout(n7175),.clk(gclk));
	jor g06920(.dina(n7175),.dinb(n7172),.dout(n7176),.clk(gclk));
	jnot g06921(.din(w_n6779_0[0]),.dout(n7177),.clk(gclk));
	jand g06922(.dina(w_n7174_0[0]),.dinb(n7177),.dout(n7178),.clk(gclk));
	jnot g06923(.din(n7178),.dout(n7179),.clk(gclk));
	jand g06924(.dina(n7179),.dinb(n7176),.dout(n7180),.clk(gclk));
	jand g06925(.dina(w_n7180_0[1]),.dinb(n7171),.dout(n7181),.clk(gclk));
	jor g06926(.dina(w_n7181_0[1]),.dinb(w_n7170_0[1]),.dout(n7182),.clk(gclk));
	jand g06927(.dina(n7182),.dinb(w_asqrt58_19[1]),.dout(n7183),.clk(gclk));
	jor g06928(.dina(w_n7170_0[0]),.dinb(w_asqrt58_19[0]),.dout(n7184),.clk(gclk));
	jor g06929(.dina(n7184),.dinb(w_n7181_0[0]),.dout(n7185),.clk(gclk));
	jnot g06930(.din(w_n6785_0[0]),.dout(n7186),.clk(gclk));
	jnot g06931(.din(w_n6787_0[0]),.dout(n7187),.clk(gclk));
	jand g06932(.dina(w_asqrt28_21[1]),.dinb(w_n6781_0[0]),.dout(n7188),.clk(gclk));
	jand g06933(.dina(w_n7188_0[1]),.dinb(n7187),.dout(n7189),.clk(gclk));
	jor g06934(.dina(n7189),.dinb(n7186),.dout(n7190),.clk(gclk));
	jnot g06935(.din(w_n6788_0[0]),.dout(n7191),.clk(gclk));
	jand g06936(.dina(w_n7188_0[0]),.dinb(n7191),.dout(n7192),.clk(gclk));
	jnot g06937(.din(n7192),.dout(n7193),.clk(gclk));
	jand g06938(.dina(n7193),.dinb(n7190),.dout(n7194),.clk(gclk));
	jand g06939(.dina(w_n7194_0[1]),.dinb(w_n7185_0[1]),.dout(n7195),.clk(gclk));
	jor g06940(.dina(n7195),.dinb(w_n7183_0[1]),.dout(n7196),.clk(gclk));
	jand g06941(.dina(w_n7196_0[1]),.dinb(w_asqrt59_19[0]),.dout(n7197),.clk(gclk));
	jxor g06942(.dina(w_n6789_0[0]),.dinb(w_n425_23[1]),.dout(n7198),.clk(gclk));
	jand g06943(.dina(n7198),.dinb(w_asqrt28_21[0]),.dout(n7199),.clk(gclk));
	jxor g06944(.dina(n7199),.dinb(w_n6799_0[0]),.dout(n7200),.clk(gclk));
	jnot g06945(.din(n7200),.dout(n7201),.clk(gclk));
	jor g06946(.dina(w_n7196_0[0]),.dinb(w_asqrt59_18[2]),.dout(n7202),.clk(gclk));
	jand g06947(.dina(w_n7202_0[1]),.dinb(w_n7201_0[1]),.dout(n7203),.clk(gclk));
	jor g06948(.dina(w_n7203_0[2]),.dinb(w_n7197_0[2]),.dout(n7204),.clk(gclk));
	jand g06949(.dina(n7204),.dinb(w_asqrt60_19[0]),.dout(n7205),.clk(gclk));
	jnot g06950(.din(w_n6804_0[0]),.dout(n7206),.clk(gclk));
	jand g06951(.dina(n7206),.dinb(w_n6802_0[0]),.dout(n7207),.clk(gclk));
	jand g06952(.dina(n7207),.dinb(w_asqrt28_20[2]),.dout(n7208),.clk(gclk));
	jxor g06953(.dina(n7208),.dinb(w_n6812_0[0]),.dout(n7209),.clk(gclk));
	jnot g06954(.din(n7209),.dout(n7210),.clk(gclk));
	jor g06955(.dina(w_n7197_0[1]),.dinb(w_asqrt60_18[2]),.dout(n7211),.clk(gclk));
	jor g06956(.dina(n7211),.dinb(w_n7203_0[1]),.dout(n7212),.clk(gclk));
	jand g06957(.dina(w_n7212_0[1]),.dinb(w_n7210_0[1]),.dout(n7213),.clk(gclk));
	jor g06958(.dina(w_n7213_0[1]),.dinb(w_n7205_0[1]),.dout(n7214),.clk(gclk));
	jand g06959(.dina(w_n7214_0[2]),.dinb(w_asqrt61_19[1]),.dout(n7215),.clk(gclk));
	jor g06960(.dina(w_n7214_0[1]),.dinb(w_asqrt61_19[0]),.dout(n7216),.clk(gclk));
	jnot g06961(.din(w_n6818_0[0]),.dout(n7217),.clk(gclk));
	jnot g06962(.din(w_n6819_0[0]),.dout(n7218),.clk(gclk));
	jand g06963(.dina(w_asqrt28_20[1]),.dinb(w_n6815_0[0]),.dout(n7219),.clk(gclk));
	jand g06964(.dina(w_n7219_0[1]),.dinb(n7218),.dout(n7220),.clk(gclk));
	jor g06965(.dina(n7220),.dinb(n7217),.dout(n7221),.clk(gclk));
	jnot g06966(.din(w_n6820_0[0]),.dout(n7222),.clk(gclk));
	jand g06967(.dina(w_n7219_0[0]),.dinb(n7222),.dout(n7223),.clk(gclk));
	jnot g06968(.din(n7223),.dout(n7224),.clk(gclk));
	jand g06969(.dina(n7224),.dinb(n7221),.dout(n7225),.clk(gclk));
	jand g06970(.dina(w_n7225_0[1]),.dinb(n7216),.dout(n7226),.clk(gclk));
	jor g06971(.dina(w_n7226_0[1]),.dinb(w_n7215_0[1]),.dout(n7227),.clk(gclk));
	jand g06972(.dina(n7227),.dinb(w_asqrt62_19[1]),.dout(n7228),.clk(gclk));
	jor g06973(.dina(w_n7215_0[0]),.dinb(w_asqrt62_19[0]),.dout(n7229),.clk(gclk));
	jor g06974(.dina(n7229),.dinb(w_n7226_0[0]),.dout(n7230),.clk(gclk));
	jnot g06975(.din(w_n6826_0[0]),.dout(n7231),.clk(gclk));
	jnot g06976(.din(w_n6828_0[0]),.dout(n7232),.clk(gclk));
	jand g06977(.dina(w_asqrt28_20[0]),.dinb(w_n6822_0[0]),.dout(n7233),.clk(gclk));
	jand g06978(.dina(w_n7233_0[1]),.dinb(n7232),.dout(n7234),.clk(gclk));
	jor g06979(.dina(n7234),.dinb(n7231),.dout(n7235),.clk(gclk));
	jnot g06980(.din(w_n6829_0[0]),.dout(n7236),.clk(gclk));
	jand g06981(.dina(w_n7233_0[0]),.dinb(n7236),.dout(n7237),.clk(gclk));
	jnot g06982(.din(n7237),.dout(n7238),.clk(gclk));
	jand g06983(.dina(n7238),.dinb(n7235),.dout(n7239),.clk(gclk));
	jand g06984(.dina(w_n7239_0[1]),.dinb(w_n7230_0[1]),.dout(n7240),.clk(gclk));
	jor g06985(.dina(n7240),.dinb(w_n7228_0[1]),.dout(n7241),.clk(gclk));
	jxor g06986(.dina(w_n6830_0[0]),.dinb(w_n199_28[2]),.dout(n7242),.clk(gclk));
	jand g06987(.dina(n7242),.dinb(w_asqrt28_19[2]),.dout(n7243),.clk(gclk));
	jxor g06988(.dina(n7243),.dinb(w_n6840_0[0]),.dout(n7244),.clk(gclk));
	jnot g06989(.din(w_n6842_0[0]),.dout(n7245),.clk(gclk));
	jand g06990(.dina(w_asqrt28_19[1]),.dinb(w_n6849_0[1]),.dout(n7246),.clk(gclk));
	jand g06991(.dina(w_n7246_0[1]),.dinb(w_n7245_0[2]),.dout(n7247),.clk(gclk));
	jor g06992(.dina(n7247),.dinb(w_n6857_0[0]),.dout(n7248),.clk(gclk));
	jor g06993(.dina(n7248),.dinb(w_n7244_0[1]),.dout(n7249),.clk(gclk));
	jnot g06994(.din(n7249),.dout(n7250),.clk(gclk));
	jand g06995(.dina(n7250),.dinb(w_n7241_1[2]),.dout(n7251),.clk(gclk));
	jor g06996(.dina(n7251),.dinb(w_asqrt63_10[1]),.dout(n7252),.clk(gclk));
	jnot g06997(.din(w_n7244_0[0]),.dout(n7253),.clk(gclk));
	jor g06998(.dina(w_n7253_0[2]),.dinb(w_n7241_1[1]),.dout(n7254),.clk(gclk));
	jor g06999(.dina(w_n7246_0[0]),.dinb(w_n7245_0[1]),.dout(n7255),.clk(gclk));
	jand g07000(.dina(w_n6849_0[0]),.dinb(w_n7245_0[0]),.dout(n7256),.clk(gclk));
	jor g07001(.dina(n7256),.dinb(w_n194_27[2]),.dout(n7257),.clk(gclk));
	jnot g07002(.din(n7257),.dout(n7258),.clk(gclk));
	jand g07003(.dina(n7258),.dinb(n7255),.dout(n7259),.clk(gclk));
	jnot g07004(.din(w_asqrt28_19[0]),.dout(n7260),.clk(gclk));
	jnot g07005(.din(w_n7259_0[1]),.dout(n7263),.clk(gclk));
	jand g07006(.dina(n7263),.dinb(w_n7254_0[1]),.dout(n7264),.clk(gclk));
	jand g07007(.dina(n7264),.dinb(w_n7252_0[1]),.dout(n7265),.clk(gclk));
	jxor g07008(.dina(w_n6932_0[0]),.dinb(w_n4499_22[0]),.dout(n7266),.clk(gclk));
	jor g07009(.dina(n7266),.dinb(w_n7265_28[1]),.dout(n7267),.clk(gclk));
	jxor g07010(.dina(n7267),.dinb(n6870),.dout(n7268),.clk(gclk));
	jnot g07011(.din(n7268),.dout(n7269),.clk(gclk));
	jor g07012(.dina(w_n7265_28[0]),.dinb(w_n6872_1[0]),.dout(n7270),.clk(gclk));
	jnot g07013(.din(w_a52_0[1]),.dout(n7271),.clk(gclk));
	jnot g07014(.din(a[53]),.dout(n7272),.clk(gclk));
	jand g07015(.dina(w_n6872_0[2]),.dinb(w_n7272_0[2]),.dout(n7273),.clk(gclk));
	jand g07016(.dina(n7273),.dinb(w_n7271_1[1]),.dout(n7274),.clk(gclk));
	jnot g07017(.din(n7274),.dout(n7275),.clk(gclk));
	jand g07018(.dina(n7275),.dinb(n7270),.dout(n7276),.clk(gclk));
	jor g07019(.dina(w_n7276_0[2]),.dinb(w_n7260_18[1]),.dout(n7277),.clk(gclk));
	jor g07020(.dina(w_n7265_27[2]),.dinb(w_a54_0[0]),.dout(n7278),.clk(gclk));
	jxor g07021(.dina(w_n7278_0[1]),.dinb(w_n6873_0[0]),.dout(n7279),.clk(gclk));
	jand g07022(.dina(w_n7276_0[1]),.dinb(w_n7260_18[0]),.dout(n7280),.clk(gclk));
	jor g07023(.dina(n7280),.dinb(w_n7279_0[1]),.dout(n7281),.clk(gclk));
	jand g07024(.dina(w_n7281_0[1]),.dinb(w_n7277_0[1]),.dout(n7282),.clk(gclk));
	jor g07025(.dina(n7282),.dinb(w_n6505_21[1]),.dout(n7283),.clk(gclk));
	jand g07026(.dina(w_n7277_0[0]),.dinb(w_n6505_21[0]),.dout(n7284),.clk(gclk));
	jand g07027(.dina(n7284),.dinb(w_n7281_0[0]),.dout(n7285),.clk(gclk));
	jor g07028(.dina(w_n7278_0[0]),.dinb(w_a55_0[0]),.dout(n7286),.clk(gclk));
	jnot g07029(.din(w_n7252_0[0]),.dout(n7287),.clk(gclk));
	jnot g07030(.din(w_n7254_0[0]),.dout(n7288),.clk(gclk));
	jor g07031(.dina(w_n7259_0[0]),.dinb(w_n7260_17[2]),.dout(n7289),.clk(gclk));
	jor g07032(.dina(n7289),.dinb(w_n7288_0[1]),.dout(n7290),.clk(gclk));
	jor g07033(.dina(n7290),.dinb(n7287),.dout(n7291),.clk(gclk));
	jand g07034(.dina(n7291),.dinb(n7286),.dout(n7292),.clk(gclk));
	jxor g07035(.dina(n7292),.dinb(w_n6510_0[1]),.dout(n7293),.clk(gclk));
	jor g07036(.dina(w_n7293_0[1]),.dinb(w_n7285_0[1]),.dout(n7294),.clk(gclk));
	jand g07037(.dina(n7294),.dinb(w_n7283_0[1]),.dout(n7295),.clk(gclk));
	jor g07038(.dina(w_n7295_0[2]),.dinb(w_n6500_18[0]),.dout(n7296),.clk(gclk));
	jand g07039(.dina(w_n7295_0[1]),.dinb(w_n6500_17[2]),.dout(n7297),.clk(gclk));
	jxor g07040(.dina(w_n6876_0[0]),.dinb(w_n6505_20[2]),.dout(n7298),.clk(gclk));
	jor g07041(.dina(n7298),.dinb(w_n7265_27[1]),.dout(n7299),.clk(gclk));
	jxor g07042(.dina(n7299),.dinb(w_n6879_0[0]),.dout(n7300),.clk(gclk));
	jor g07043(.dina(w_n7300_0[1]),.dinb(n7297),.dout(n7301),.clk(gclk));
	jand g07044(.dina(w_n7301_0[1]),.dinb(w_n7296_0[1]),.dout(n7302),.clk(gclk));
	jor g07045(.dina(n7302),.dinb(w_n5793_21[2]),.dout(n7303),.clk(gclk));
	jnot g07046(.din(w_n6885_0[0]),.dout(n7304),.clk(gclk));
	jor g07047(.dina(n7304),.dinb(w_n6883_0[0]),.dout(n7305),.clk(gclk));
	jor g07048(.dina(n7305),.dinb(w_n7265_27[0]),.dout(n7306),.clk(gclk));
	jxor g07049(.dina(n7306),.dinb(w_n6894_0[0]),.dout(n7307),.clk(gclk));
	jand g07050(.dina(w_n7296_0[0]),.dinb(w_n5793_21[1]),.dout(n7308),.clk(gclk));
	jand g07051(.dina(n7308),.dinb(w_n7301_0[0]),.dout(n7309),.clk(gclk));
	jor g07052(.dina(w_n7309_0[1]),.dinb(w_n7307_0[1]),.dout(n7310),.clk(gclk));
	jand g07053(.dina(w_n7310_0[1]),.dinb(w_n7303_0[1]),.dout(n7311),.clk(gclk));
	jor g07054(.dina(w_n7311_0[2]),.dinb(w_n5788_18[1]),.dout(n7312),.clk(gclk));
	jand g07055(.dina(w_n7311_0[1]),.dinb(w_n5788_18[0]),.dout(n7313),.clk(gclk));
	jxor g07056(.dina(w_n6896_0[0]),.dinb(w_n5793_21[0]),.dout(n7314),.clk(gclk));
	jor g07057(.dina(n7314),.dinb(w_n7265_26[2]),.dout(n7315),.clk(gclk));
	jxor g07058(.dina(n7315),.dinb(w_n6901_0[0]),.dout(n7316),.clk(gclk));
	jnot g07059(.din(w_n7316_0[1]),.dout(n7317),.clk(gclk));
	jor g07060(.dina(n7317),.dinb(n7313),.dout(n7318),.clk(gclk));
	jand g07061(.dina(w_n7318_0[1]),.dinb(w_n7312_0[1]),.dout(n7319),.clk(gclk));
	jor g07062(.dina(n7319),.dinb(w_n5121_21[1]),.dout(n7320),.clk(gclk));
	jand g07063(.dina(w_n7312_0[0]),.dinb(w_n5121_21[0]),.dout(n7321),.clk(gclk));
	jand g07064(.dina(n7321),.dinb(w_n7318_0[0]),.dout(n7322),.clk(gclk));
	jnot g07065(.din(w_n6905_0[0]),.dout(n7323),.clk(gclk));
	jnot g07066(.din(w_n7265_26[1]),.dout(asqrt_fa_28),.clk(gclk));
	jand g07067(.dina(w_asqrt27_20[1]),.dinb(n7323),.dout(n7325),.clk(gclk));
	jand g07068(.dina(w_n7325_0[1]),.dinb(w_n6912_0[0]),.dout(n7326),.clk(gclk));
	jor g07069(.dina(n7326),.dinb(w_n6910_0[0]),.dout(n7327),.clk(gclk));
	jand g07070(.dina(w_n7325_0[0]),.dinb(w_n6913_0[0]),.dout(n7328),.clk(gclk));
	jnot g07071(.din(n7328),.dout(n7329),.clk(gclk));
	jand g07072(.dina(n7329),.dinb(n7327),.dout(n7330),.clk(gclk));
	jnot g07073(.din(n7330),.dout(n7331),.clk(gclk));
	jor g07074(.dina(w_n7331_0[1]),.dinb(w_n7322_0[1]),.dout(n7332),.clk(gclk));
	jand g07075(.dina(n7332),.dinb(w_n7320_0[1]),.dout(n7333),.clk(gclk));
	jor g07076(.dina(w_n7333_0[2]),.dinb(w_n5116_18[1]),.dout(n7334),.clk(gclk));
	jand g07077(.dina(w_n7333_0[1]),.dinb(w_n5116_18[0]),.dout(n7335),.clk(gclk));
	jnot g07078(.din(w_n6920_0[0]),.dout(n7336),.clk(gclk));
	jxor g07079(.dina(w_n6914_0[0]),.dinb(w_n5121_20[2]),.dout(n7337),.clk(gclk));
	jor g07080(.dina(n7337),.dinb(w_n7265_26[0]),.dout(n7338),.clk(gclk));
	jxor g07081(.dina(n7338),.dinb(n7336),.dout(n7339),.clk(gclk));
	jnot g07082(.din(w_n7339_0[1]),.dout(n7340),.clk(gclk));
	jor g07083(.dina(n7340),.dinb(n7335),.dout(n7341),.clk(gclk));
	jand g07084(.dina(w_n7341_0[1]),.dinb(w_n7334_0[1]),.dout(n7342),.clk(gclk));
	jor g07085(.dina(n7342),.dinb(w_n4499_21[2]),.dout(n7343),.clk(gclk));
	jand g07086(.dina(w_n7334_0[0]),.dinb(w_n4499_21[1]),.dout(n7344),.clk(gclk));
	jand g07087(.dina(n7344),.dinb(w_n7341_0[0]),.dout(n7345),.clk(gclk));
	jnot g07088(.din(w_n6923_0[0]),.dout(n7346),.clk(gclk));
	jand g07089(.dina(w_asqrt27_20[0]),.dinb(n7346),.dout(n7347),.clk(gclk));
	jand g07090(.dina(w_n7347_0[1]),.dinb(w_n6930_0[0]),.dout(n7348),.clk(gclk));
	jor g07091(.dina(n7348),.dinb(w_n6928_0[0]),.dout(n7349),.clk(gclk));
	jand g07092(.dina(w_n7347_0[0]),.dinb(w_n6931_0[0]),.dout(n7350),.clk(gclk));
	jnot g07093(.din(n7350),.dout(n7351),.clk(gclk));
	jand g07094(.dina(n7351),.dinb(n7349),.dout(n7352),.clk(gclk));
	jnot g07095(.din(n7352),.dout(n7353),.clk(gclk));
	jor g07096(.dina(w_n7353_0[1]),.dinb(w_n7345_0[1]),.dout(n7354),.clk(gclk));
	jand g07097(.dina(n7354),.dinb(w_n7343_0[1]),.dout(n7355),.clk(gclk));
	jor g07098(.dina(w_n7355_0[2]),.dinb(w_n4494_19[0]),.dout(n7356),.clk(gclk));
	jand g07099(.dina(w_n7355_0[1]),.dinb(w_n4494_18[2]),.dout(n7357),.clk(gclk));
	jor g07100(.dina(n7357),.dinb(w_n7269_0[1]),.dout(n7358),.clk(gclk));
	jand g07101(.dina(w_n7358_0[1]),.dinb(w_n7356_0[1]),.dout(n7359),.clk(gclk));
	jor g07102(.dina(n7359),.dinb(w_n3912_22[0]),.dout(n7360),.clk(gclk));
	jnot g07103(.din(w_n6939_0[0]),.dout(n7361),.clk(gclk));
	jor g07104(.dina(n7361),.dinb(w_n6937_0[0]),.dout(n7362),.clk(gclk));
	jor g07105(.dina(n7362),.dinb(w_n7265_25[2]),.dout(n7363),.clk(gclk));
	jxor g07106(.dina(n7363),.dinb(w_n6948_0[0]),.dout(n7364),.clk(gclk));
	jand g07107(.dina(w_n7356_0[0]),.dinb(w_n3912_21[2]),.dout(n7365),.clk(gclk));
	jand g07108(.dina(n7365),.dinb(w_n7358_0[0]),.dout(n7366),.clk(gclk));
	jor g07109(.dina(w_n7366_0[1]),.dinb(w_n7364_0[1]),.dout(n7367),.clk(gclk));
	jand g07110(.dina(w_n7367_0[1]),.dinb(w_n7360_0[1]),.dout(n7368),.clk(gclk));
	jor g07111(.dina(w_n7368_0[1]),.dinb(w_n3907_19[0]),.dout(n7369),.clk(gclk));
	jxor g07112(.dina(w_n6950_0[0]),.dinb(w_n3912_21[1]),.dout(n7370),.clk(gclk));
	jor g07113(.dina(n7370),.dinb(w_n7265_25[1]),.dout(n7371),.clk(gclk));
	jxor g07114(.dina(n7371),.dinb(w_n6955_0[0]),.dout(n7372),.clk(gclk));
	jand g07115(.dina(w_n7368_0[0]),.dinb(w_n3907_18[2]),.dout(n7373),.clk(gclk));
	jor g07116(.dina(w_n7373_0[1]),.dinb(w_n7372_0[1]),.dout(n7374),.clk(gclk));
	jand g07117(.dina(w_n7374_0[2]),.dinb(w_n7369_0[2]),.dout(n7375),.clk(gclk));
	jor g07118(.dina(n7375),.dinb(w_n3376_22[2]),.dout(n7376),.clk(gclk));
	jnot g07119(.din(w_n6960_0[0]),.dout(n7377),.clk(gclk));
	jor g07120(.dina(n7377),.dinb(w_n6958_0[0]),.dout(n7378),.clk(gclk));
	jor g07121(.dina(n7378),.dinb(w_n7265_25[0]),.dout(n7379),.clk(gclk));
	jxor g07122(.dina(n7379),.dinb(w_n6969_0[0]),.dout(n7380),.clk(gclk));
	jand g07123(.dina(w_n7369_0[1]),.dinb(w_n3376_22[1]),.dout(n7381),.clk(gclk));
	jand g07124(.dina(n7381),.dinb(w_n7374_0[1]),.dout(n7382),.clk(gclk));
	jor g07125(.dina(w_n7382_0[1]),.dinb(w_n7380_0[1]),.dout(n7383),.clk(gclk));
	jand g07126(.dina(w_n7383_0[1]),.dinb(w_n7376_0[1]),.dout(n7384),.clk(gclk));
	jor g07127(.dina(w_n7384_0[2]),.dinb(w_n3371_19[2]),.dout(n7385),.clk(gclk));
	jand g07128(.dina(w_n7384_0[1]),.dinb(w_n3371_19[1]),.dout(n7386),.clk(gclk));
	jnot g07129(.din(w_n6972_0[0]),.dout(n7387),.clk(gclk));
	jand g07130(.dina(w_asqrt27_19[2]),.dinb(n7387),.dout(n7388),.clk(gclk));
	jand g07131(.dina(w_n7388_0[1]),.dinb(w_n6977_0[0]),.dout(n7389),.clk(gclk));
	jor g07132(.dina(n7389),.dinb(w_n6976_0[0]),.dout(n7390),.clk(gclk));
	jand g07133(.dina(w_n7388_0[0]),.dinb(w_n6978_0[0]),.dout(n7391),.clk(gclk));
	jnot g07134(.din(n7391),.dout(n7392),.clk(gclk));
	jand g07135(.dina(n7392),.dinb(n7390),.dout(n7393),.clk(gclk));
	jnot g07136(.din(n7393),.dout(n7394),.clk(gclk));
	jor g07137(.dina(w_n7394_0[1]),.dinb(n7386),.dout(n7395),.clk(gclk));
	jand g07138(.dina(w_n7395_0[1]),.dinb(w_n7385_0[1]),.dout(n7396),.clk(gclk));
	jor g07139(.dina(n7396),.dinb(w_n2875_22[2]),.dout(n7397),.clk(gclk));
	jand g07140(.dina(w_n7385_0[0]),.dinb(w_n2875_22[1]),.dout(n7398),.clk(gclk));
	jand g07141(.dina(n7398),.dinb(w_n7395_0[0]),.dout(n7399),.clk(gclk));
	jnot g07142(.din(w_n6980_0[0]),.dout(n7400),.clk(gclk));
	jand g07143(.dina(w_asqrt27_19[1]),.dinb(n7400),.dout(n7401),.clk(gclk));
	jand g07144(.dina(w_n7401_0[1]),.dinb(w_n6987_0[0]),.dout(n7402),.clk(gclk));
	jor g07145(.dina(n7402),.dinb(w_n6985_0[0]),.dout(n7403),.clk(gclk));
	jand g07146(.dina(w_n7401_0[0]),.dinb(w_n6988_0[0]),.dout(n7404),.clk(gclk));
	jnot g07147(.din(n7404),.dout(n7405),.clk(gclk));
	jand g07148(.dina(n7405),.dinb(n7403),.dout(n7406),.clk(gclk));
	jnot g07149(.din(n7406),.dout(n7407),.clk(gclk));
	jor g07150(.dina(w_n7407_0[1]),.dinb(w_n7399_0[1]),.dout(n7408),.clk(gclk));
	jand g07151(.dina(n7408),.dinb(w_n7397_0[1]),.dout(n7409),.clk(gclk));
	jor g07152(.dina(w_n7409_0[1]),.dinb(w_n2870_19[2]),.dout(n7410),.clk(gclk));
	jxor g07153(.dina(w_n6989_0[0]),.dinb(w_n2875_22[0]),.dout(n7411),.clk(gclk));
	jor g07154(.dina(n7411),.dinb(w_n7265_24[2]),.dout(n7412),.clk(gclk));
	jxor g07155(.dina(n7412),.dinb(w_n7000_0[0]),.dout(n7413),.clk(gclk));
	jand g07156(.dina(w_n7409_0[0]),.dinb(w_n2870_19[1]),.dout(n7414),.clk(gclk));
	jor g07157(.dina(w_n7414_0[1]),.dinb(w_n7413_0[1]),.dout(n7415),.clk(gclk));
	jand g07158(.dina(w_n7415_0[2]),.dinb(w_n7410_0[2]),.dout(n7416),.clk(gclk));
	jor g07159(.dina(n7416),.dinb(w_n2425_23[0]),.dout(n7417),.clk(gclk));
	jnot g07160(.din(w_n7005_0[0]),.dout(n7418),.clk(gclk));
	jor g07161(.dina(n7418),.dinb(w_n7003_0[0]),.dout(n7419),.clk(gclk));
	jor g07162(.dina(n7419),.dinb(w_n7265_24[1]),.dout(n7420),.clk(gclk));
	jxor g07163(.dina(n7420),.dinb(w_n7014_0[0]),.dout(n7421),.clk(gclk));
	jand g07164(.dina(w_n7410_0[1]),.dinb(w_n2425_22[2]),.dout(n7422),.clk(gclk));
	jand g07165(.dina(n7422),.dinb(w_n7415_0[1]),.dout(n7423),.clk(gclk));
	jor g07166(.dina(w_n7423_0[1]),.dinb(w_n7421_0[1]),.dout(n7424),.clk(gclk));
	jand g07167(.dina(w_n7424_0[1]),.dinb(w_n7417_0[1]),.dout(n7425),.clk(gclk));
	jor g07168(.dina(w_n7425_0[2]),.dinb(w_n2420_20[2]),.dout(n7426),.clk(gclk));
	jand g07169(.dina(w_n7425_0[1]),.dinb(w_n2420_20[1]),.dout(n7427),.clk(gclk));
	jnot g07170(.din(w_n7017_0[0]),.dout(n7428),.clk(gclk));
	jand g07171(.dina(w_asqrt27_19[0]),.dinb(n7428),.dout(n7429),.clk(gclk));
	jand g07172(.dina(w_n7429_0[1]),.dinb(w_n7022_0[0]),.dout(n7430),.clk(gclk));
	jor g07173(.dina(n7430),.dinb(w_n7021_0[0]),.dout(n7431),.clk(gclk));
	jand g07174(.dina(w_n7429_0[0]),.dinb(w_n7023_0[0]),.dout(n7432),.clk(gclk));
	jnot g07175(.din(n7432),.dout(n7433),.clk(gclk));
	jand g07176(.dina(n7433),.dinb(n7431),.dout(n7434),.clk(gclk));
	jnot g07177(.din(n7434),.dout(n7435),.clk(gclk));
	jor g07178(.dina(w_n7435_0[1]),.dinb(n7427),.dout(n7436),.clk(gclk));
	jand g07179(.dina(w_n7436_0[1]),.dinb(w_n7426_0[1]),.dout(n7437),.clk(gclk));
	jor g07180(.dina(n7437),.dinb(w_n2010_23[0]),.dout(n7438),.clk(gclk));
	jand g07181(.dina(w_n7426_0[0]),.dinb(w_n2010_22[2]),.dout(n7439),.clk(gclk));
	jand g07182(.dina(n7439),.dinb(w_n7436_0[0]),.dout(n7440),.clk(gclk));
	jnot g07183(.din(w_n7025_0[0]),.dout(n7441),.clk(gclk));
	jand g07184(.dina(w_asqrt27_18[2]),.dinb(n7441),.dout(n7442),.clk(gclk));
	jand g07185(.dina(w_n7442_0[1]),.dinb(w_n7032_0[0]),.dout(n7443),.clk(gclk));
	jor g07186(.dina(n7443),.dinb(w_n7030_0[0]),.dout(n7444),.clk(gclk));
	jand g07187(.dina(w_n7442_0[0]),.dinb(w_n7033_0[0]),.dout(n7445),.clk(gclk));
	jnot g07188(.din(n7445),.dout(n7446),.clk(gclk));
	jand g07189(.dina(n7446),.dinb(n7444),.dout(n7447),.clk(gclk));
	jnot g07190(.din(n7447),.dout(n7448),.clk(gclk));
	jor g07191(.dina(w_n7448_0[1]),.dinb(w_n7440_0[1]),.dout(n7449),.clk(gclk));
	jand g07192(.dina(n7449),.dinb(w_n7438_0[1]),.dout(n7450),.clk(gclk));
	jor g07193(.dina(w_n7450_0[1]),.dinb(w_n2005_20[2]),.dout(n7451),.clk(gclk));
	jxor g07194(.dina(w_n7034_0[0]),.dinb(w_n2010_22[1]),.dout(n7452),.clk(gclk));
	jor g07195(.dina(n7452),.dinb(w_n7265_24[0]),.dout(n7453),.clk(gclk));
	jxor g07196(.dina(n7453),.dinb(w_n7045_0[0]),.dout(n7454),.clk(gclk));
	jand g07197(.dina(w_n7450_0[0]),.dinb(w_n2005_20[1]),.dout(n7455),.clk(gclk));
	jor g07198(.dina(w_n7455_0[1]),.dinb(w_n7454_0[1]),.dout(n7456),.clk(gclk));
	jand g07199(.dina(w_n7456_0[2]),.dinb(w_n7451_0[2]),.dout(n7457),.clk(gclk));
	jor g07200(.dina(n7457),.dinb(w_n1646_23[2]),.dout(n7458),.clk(gclk));
	jnot g07201(.din(w_n7050_0[0]),.dout(n7459),.clk(gclk));
	jor g07202(.dina(n7459),.dinb(w_n7048_0[0]),.dout(n7460),.clk(gclk));
	jor g07203(.dina(n7460),.dinb(w_n7265_23[2]),.dout(n7461),.clk(gclk));
	jxor g07204(.dina(n7461),.dinb(w_n7059_0[0]),.dout(n7462),.clk(gclk));
	jand g07205(.dina(w_n7451_0[1]),.dinb(w_n1646_23[1]),.dout(n7463),.clk(gclk));
	jand g07206(.dina(n7463),.dinb(w_n7456_0[1]),.dout(n7464),.clk(gclk));
	jor g07207(.dina(w_n7464_0[1]),.dinb(w_n7462_0[1]),.dout(n7465),.clk(gclk));
	jand g07208(.dina(w_n7465_0[1]),.dinb(w_n7458_0[1]),.dout(n7466),.clk(gclk));
	jor g07209(.dina(w_n7466_0[2]),.dinb(w_n1641_21[1]),.dout(n7467),.clk(gclk));
	jand g07210(.dina(w_n7466_0[1]),.dinb(w_n1641_21[0]),.dout(n7468),.clk(gclk));
	jnot g07211(.din(w_n7062_0[0]),.dout(n7469),.clk(gclk));
	jand g07212(.dina(w_asqrt27_18[1]),.dinb(n7469),.dout(n7470),.clk(gclk));
	jand g07213(.dina(w_n7470_0[1]),.dinb(w_n7067_0[0]),.dout(n7471),.clk(gclk));
	jor g07214(.dina(n7471),.dinb(w_n7066_0[0]),.dout(n7472),.clk(gclk));
	jand g07215(.dina(w_n7470_0[0]),.dinb(w_n7068_0[0]),.dout(n7473),.clk(gclk));
	jnot g07216(.din(n7473),.dout(n7474),.clk(gclk));
	jand g07217(.dina(n7474),.dinb(n7472),.dout(n7475),.clk(gclk));
	jnot g07218(.din(n7475),.dout(n7476),.clk(gclk));
	jor g07219(.dina(w_n7476_0[1]),.dinb(n7468),.dout(n7477),.clk(gclk));
	jand g07220(.dina(w_n7477_0[1]),.dinb(w_n7467_0[1]),.dout(n7478),.clk(gclk));
	jor g07221(.dina(n7478),.dinb(w_n1317_23[2]),.dout(n7479),.clk(gclk));
	jand g07222(.dina(w_n7467_0[0]),.dinb(w_n1317_23[1]),.dout(n7480),.clk(gclk));
	jand g07223(.dina(n7480),.dinb(w_n7477_0[0]),.dout(n7481),.clk(gclk));
	jnot g07224(.din(w_n7070_0[0]),.dout(n7482),.clk(gclk));
	jand g07225(.dina(w_asqrt27_18[0]),.dinb(n7482),.dout(n7483),.clk(gclk));
	jand g07226(.dina(w_n7483_0[1]),.dinb(w_n7077_0[0]),.dout(n7484),.clk(gclk));
	jor g07227(.dina(n7484),.dinb(w_n7075_0[0]),.dout(n7485),.clk(gclk));
	jand g07228(.dina(w_n7483_0[0]),.dinb(w_n7078_0[0]),.dout(n7486),.clk(gclk));
	jnot g07229(.din(n7486),.dout(n7487),.clk(gclk));
	jand g07230(.dina(n7487),.dinb(n7485),.dout(n7488),.clk(gclk));
	jnot g07231(.din(n7488),.dout(n7489),.clk(gclk));
	jor g07232(.dina(w_n7489_0[1]),.dinb(w_n7481_0[1]),.dout(n7490),.clk(gclk));
	jand g07233(.dina(n7490),.dinb(w_n7479_0[1]),.dout(n7491),.clk(gclk));
	jor g07234(.dina(w_n7491_0[1]),.dinb(w_n1312_21[1]),.dout(n7492),.clk(gclk));
	jxor g07235(.dina(w_n7079_0[0]),.dinb(w_n1317_23[0]),.dout(n7493),.clk(gclk));
	jor g07236(.dina(n7493),.dinb(w_n7265_23[1]),.dout(n7494),.clk(gclk));
	jxor g07237(.dina(n7494),.dinb(w_n7090_0[0]),.dout(n7495),.clk(gclk));
	jand g07238(.dina(w_n7491_0[0]),.dinb(w_n1312_21[0]),.dout(n7496),.clk(gclk));
	jor g07239(.dina(w_n7496_0[1]),.dinb(w_n7495_0[1]),.dout(n7497),.clk(gclk));
	jand g07240(.dina(w_n7497_0[2]),.dinb(w_n7492_0[2]),.dout(n7498),.clk(gclk));
	jor g07241(.dina(n7498),.dinb(w_n1039_24[0]),.dout(n7499),.clk(gclk));
	jnot g07242(.din(w_n7095_0[0]),.dout(n7500),.clk(gclk));
	jor g07243(.dina(n7500),.dinb(w_n7093_0[0]),.dout(n7501),.clk(gclk));
	jor g07244(.dina(n7501),.dinb(w_n7265_23[0]),.dout(n7502),.clk(gclk));
	jxor g07245(.dina(n7502),.dinb(w_n7104_0[0]),.dout(n7503),.clk(gclk));
	jand g07246(.dina(w_n7492_0[1]),.dinb(w_n1039_23[2]),.dout(n7504),.clk(gclk));
	jand g07247(.dina(n7504),.dinb(w_n7497_0[1]),.dout(n7505),.clk(gclk));
	jor g07248(.dina(w_n7505_0[1]),.dinb(w_n7503_0[1]),.dout(n7506),.clk(gclk));
	jand g07249(.dina(w_n7506_0[1]),.dinb(w_n7499_0[1]),.dout(n7507),.clk(gclk));
	jor g07250(.dina(w_n7507_0[2]),.dinb(w_n1034_22[1]),.dout(n7508),.clk(gclk));
	jand g07251(.dina(w_n7507_0[1]),.dinb(w_n1034_22[0]),.dout(n7509),.clk(gclk));
	jnot g07252(.din(w_n7107_0[0]),.dout(n7510),.clk(gclk));
	jand g07253(.dina(w_asqrt27_17[2]),.dinb(n7510),.dout(n7511),.clk(gclk));
	jand g07254(.dina(w_n7511_0[1]),.dinb(w_n7112_0[0]),.dout(n7512),.clk(gclk));
	jor g07255(.dina(n7512),.dinb(w_n7111_0[0]),.dout(n7513),.clk(gclk));
	jand g07256(.dina(w_n7511_0[0]),.dinb(w_n7113_0[0]),.dout(n7514),.clk(gclk));
	jnot g07257(.din(n7514),.dout(n7515),.clk(gclk));
	jand g07258(.dina(n7515),.dinb(n7513),.dout(n7516),.clk(gclk));
	jnot g07259(.din(n7516),.dout(n7517),.clk(gclk));
	jor g07260(.dina(w_n7517_0[1]),.dinb(n7509),.dout(n7518),.clk(gclk));
	jand g07261(.dina(w_n7518_0[1]),.dinb(w_n7508_0[1]),.dout(n7519),.clk(gclk));
	jor g07262(.dina(n7519),.dinb(w_n796_24[0]),.dout(n7520),.clk(gclk));
	jand g07263(.dina(w_n7508_0[0]),.dinb(w_n796_23[2]),.dout(n7521),.clk(gclk));
	jand g07264(.dina(n7521),.dinb(w_n7518_0[0]),.dout(n7522),.clk(gclk));
	jnot g07265(.din(w_n7115_0[0]),.dout(n7523),.clk(gclk));
	jand g07266(.dina(w_asqrt27_17[1]),.dinb(n7523),.dout(n7524),.clk(gclk));
	jand g07267(.dina(w_n7524_0[1]),.dinb(w_n7122_0[0]),.dout(n7525),.clk(gclk));
	jor g07268(.dina(n7525),.dinb(w_n7120_0[0]),.dout(n7526),.clk(gclk));
	jand g07269(.dina(w_n7524_0[0]),.dinb(w_n7123_0[0]),.dout(n7527),.clk(gclk));
	jnot g07270(.din(n7527),.dout(n7528),.clk(gclk));
	jand g07271(.dina(n7528),.dinb(n7526),.dout(n7529),.clk(gclk));
	jnot g07272(.din(n7529),.dout(n7530),.clk(gclk));
	jor g07273(.dina(w_n7530_0[1]),.dinb(w_n7522_0[1]),.dout(n7531),.clk(gclk));
	jand g07274(.dina(n7531),.dinb(w_n7520_0[1]),.dout(n7532),.clk(gclk));
	jor g07275(.dina(w_n7532_0[1]),.dinb(w_n791_22[1]),.dout(n7533),.clk(gclk));
	jxor g07276(.dina(w_n7124_0[0]),.dinb(w_n796_23[1]),.dout(n7534),.clk(gclk));
	jor g07277(.dina(n7534),.dinb(w_n7265_22[2]),.dout(n7535),.clk(gclk));
	jxor g07278(.dina(n7535),.dinb(w_n7135_0[0]),.dout(n7536),.clk(gclk));
	jand g07279(.dina(w_n7532_0[0]),.dinb(w_n791_22[0]),.dout(n7537),.clk(gclk));
	jor g07280(.dina(w_n7537_0[1]),.dinb(w_n7536_0[1]),.dout(n7538),.clk(gclk));
	jand g07281(.dina(w_n7538_0[2]),.dinb(w_n7533_0[2]),.dout(n7539),.clk(gclk));
	jor g07282(.dina(n7539),.dinb(w_n595_24[1]),.dout(n7540),.clk(gclk));
	jnot g07283(.din(w_n7140_0[0]),.dout(n7541),.clk(gclk));
	jor g07284(.dina(n7541),.dinb(w_n7138_0[0]),.dout(n7542),.clk(gclk));
	jor g07285(.dina(n7542),.dinb(w_n7265_22[1]),.dout(n7543),.clk(gclk));
	jxor g07286(.dina(n7543),.dinb(w_n7149_0[0]),.dout(n7544),.clk(gclk));
	jand g07287(.dina(w_n7533_0[1]),.dinb(w_n595_24[0]),.dout(n7545),.clk(gclk));
	jand g07288(.dina(n7545),.dinb(w_n7538_0[1]),.dout(n7546),.clk(gclk));
	jor g07289(.dina(w_n7546_0[1]),.dinb(w_n7544_0[1]),.dout(n7547),.clk(gclk));
	jand g07290(.dina(w_n7547_0[1]),.dinb(w_n7540_0[1]),.dout(n7548),.clk(gclk));
	jor g07291(.dina(w_n7548_0[2]),.dinb(w_n590_23[0]),.dout(n7549),.clk(gclk));
	jand g07292(.dina(w_n7548_0[1]),.dinb(w_n590_22[2]),.dout(n7550),.clk(gclk));
	jnot g07293(.din(w_n7152_0[0]),.dout(n7551),.clk(gclk));
	jand g07294(.dina(w_asqrt27_17[0]),.dinb(n7551),.dout(n7552),.clk(gclk));
	jand g07295(.dina(w_n7552_0[1]),.dinb(w_n7157_0[0]),.dout(n7553),.clk(gclk));
	jor g07296(.dina(n7553),.dinb(w_n7156_0[0]),.dout(n7554),.clk(gclk));
	jand g07297(.dina(w_n7552_0[0]),.dinb(w_n7158_0[0]),.dout(n7555),.clk(gclk));
	jnot g07298(.din(n7555),.dout(n7556),.clk(gclk));
	jand g07299(.dina(n7556),.dinb(n7554),.dout(n7557),.clk(gclk));
	jnot g07300(.din(n7557),.dout(n7558),.clk(gclk));
	jor g07301(.dina(w_n7558_0[1]),.dinb(n7550),.dout(n7559),.clk(gclk));
	jand g07302(.dina(w_n7559_0[1]),.dinb(w_n7549_0[1]),.dout(n7560),.clk(gclk));
	jor g07303(.dina(n7560),.dinb(w_n430_24[1]),.dout(n7561),.clk(gclk));
	jand g07304(.dina(w_n7549_0[0]),.dinb(w_n430_24[0]),.dout(n7562),.clk(gclk));
	jand g07305(.dina(n7562),.dinb(w_n7559_0[0]),.dout(n7563),.clk(gclk));
	jnot g07306(.din(w_n7160_0[0]),.dout(n7564),.clk(gclk));
	jand g07307(.dina(w_asqrt27_16[2]),.dinb(n7564),.dout(n7565),.clk(gclk));
	jand g07308(.dina(w_n7565_0[1]),.dinb(w_n7167_0[0]),.dout(n7566),.clk(gclk));
	jor g07309(.dina(n7566),.dinb(w_n7165_0[0]),.dout(n7567),.clk(gclk));
	jand g07310(.dina(w_n7565_0[0]),.dinb(w_n7168_0[0]),.dout(n7568),.clk(gclk));
	jnot g07311(.din(n7568),.dout(n7569),.clk(gclk));
	jand g07312(.dina(n7569),.dinb(n7567),.dout(n7570),.clk(gclk));
	jnot g07313(.din(n7570),.dout(n7571),.clk(gclk));
	jor g07314(.dina(w_n7571_0[1]),.dinb(w_n7563_0[1]),.dout(n7572),.clk(gclk));
	jand g07315(.dina(n7572),.dinb(w_n7561_0[1]),.dout(n7573),.clk(gclk));
	jor g07316(.dina(w_n7573_0[1]),.dinb(w_n425_23[0]),.dout(n7574),.clk(gclk));
	jxor g07317(.dina(w_n7169_0[0]),.dinb(w_n430_23[2]),.dout(n7575),.clk(gclk));
	jor g07318(.dina(n7575),.dinb(w_n7265_22[0]),.dout(n7576),.clk(gclk));
	jxor g07319(.dina(n7576),.dinb(w_n7180_0[0]),.dout(n7577),.clk(gclk));
	jand g07320(.dina(w_n7573_0[0]),.dinb(w_n425_22[2]),.dout(n7578),.clk(gclk));
	jor g07321(.dina(w_n7578_0[1]),.dinb(w_n7577_0[1]),.dout(n7579),.clk(gclk));
	jand g07322(.dina(w_n7579_0[2]),.dinb(w_n7574_0[2]),.dout(n7580),.clk(gclk));
	jor g07323(.dina(n7580),.dinb(w_n305_24[2]),.dout(n7581),.clk(gclk));
	jnot g07324(.din(w_n7185_0[0]),.dout(n7582),.clk(gclk));
	jor g07325(.dina(n7582),.dinb(w_n7183_0[0]),.dout(n7583),.clk(gclk));
	jor g07326(.dina(n7583),.dinb(w_n7265_21[2]),.dout(n7584),.clk(gclk));
	jxor g07327(.dina(n7584),.dinb(w_n7194_0[0]),.dout(n7585),.clk(gclk));
	jand g07328(.dina(w_n7574_0[1]),.dinb(w_n305_24[1]),.dout(n7586),.clk(gclk));
	jand g07329(.dina(n7586),.dinb(w_n7579_0[1]),.dout(n7587),.clk(gclk));
	jor g07330(.dina(w_n7587_0[1]),.dinb(w_n7585_0[1]),.dout(n7588),.clk(gclk));
	jand g07331(.dina(w_n7588_0[1]),.dinb(w_n7581_0[1]),.dout(n7589),.clk(gclk));
	jor g07332(.dina(w_n7589_0[2]),.dinb(w_n290_24[1]),.dout(n7590),.clk(gclk));
	jand g07333(.dina(w_n7589_0[1]),.dinb(w_n290_24[0]),.dout(n7591),.clk(gclk));
	jnot g07334(.din(w_n7197_0[0]),.dout(n7592),.clk(gclk));
	jand g07335(.dina(w_asqrt27_16[1]),.dinb(n7592),.dout(n7593),.clk(gclk));
	jand g07336(.dina(w_n7593_0[1]),.dinb(w_n7202_0[0]),.dout(n7594),.clk(gclk));
	jor g07337(.dina(n7594),.dinb(w_n7201_0[0]),.dout(n7595),.clk(gclk));
	jand g07338(.dina(w_n7593_0[0]),.dinb(w_n7203_0[0]),.dout(n7596),.clk(gclk));
	jnot g07339(.din(n7596),.dout(n7597),.clk(gclk));
	jand g07340(.dina(n7597),.dinb(n7595),.dout(n7598),.clk(gclk));
	jnot g07341(.din(n7598),.dout(n7599),.clk(gclk));
	jor g07342(.dina(w_n7599_0[1]),.dinb(n7591),.dout(n7600),.clk(gclk));
	jand g07343(.dina(w_n7600_0[1]),.dinb(w_n7590_0[1]),.dout(n7601),.clk(gclk));
	jor g07344(.dina(n7601),.dinb(w_n223_24[2]),.dout(n7602),.clk(gclk));
	jand g07345(.dina(w_n7590_0[0]),.dinb(w_n223_24[1]),.dout(n7603),.clk(gclk));
	jand g07346(.dina(n7603),.dinb(w_n7600_0[0]),.dout(n7604),.clk(gclk));
	jnot g07347(.din(w_n7205_0[0]),.dout(n7605),.clk(gclk));
	jand g07348(.dina(w_asqrt27_16[0]),.dinb(n7605),.dout(n7606),.clk(gclk));
	jand g07349(.dina(w_n7606_0[1]),.dinb(w_n7212_0[0]),.dout(n7607),.clk(gclk));
	jor g07350(.dina(n7607),.dinb(w_n7210_0[0]),.dout(n7608),.clk(gclk));
	jand g07351(.dina(w_n7606_0[0]),.dinb(w_n7213_0[0]),.dout(n7609),.clk(gclk));
	jnot g07352(.din(n7609),.dout(n7610),.clk(gclk));
	jand g07353(.dina(n7610),.dinb(n7608),.dout(n7611),.clk(gclk));
	jnot g07354(.din(n7611),.dout(n7612),.clk(gclk));
	jor g07355(.dina(w_n7612_0[1]),.dinb(w_n7604_0[1]),.dout(n7613),.clk(gclk));
	jand g07356(.dina(n7613),.dinb(w_n7602_0[1]),.dout(n7614),.clk(gclk));
	jor g07357(.dina(w_n7614_0[2]),.dinb(w_n199_28[1]),.dout(n7615),.clk(gclk));
	jand g07358(.dina(w_n7614_0[1]),.dinb(w_n199_28[0]),.dout(n7616),.clk(gclk));
	jxor g07359(.dina(w_n7214_0[0]),.dinb(w_n223_24[0]),.dout(n7617),.clk(gclk));
	jor g07360(.dina(n7617),.dinb(w_n7265_21[1]),.dout(n7618),.clk(gclk));
	jxor g07361(.dina(n7618),.dinb(w_n7225_0[0]),.dout(n7619),.clk(gclk));
	jor g07362(.dina(w_n7619_0[1]),.dinb(n7616),.dout(n7620),.clk(gclk));
	jand g07363(.dina(n7620),.dinb(n7615),.dout(n7621),.clk(gclk));
	jnot g07364(.din(w_n7230_0[0]),.dout(n7622),.clk(gclk));
	jor g07365(.dina(n7622),.dinb(w_n7228_0[0]),.dout(n7623),.clk(gclk));
	jor g07366(.dina(n7623),.dinb(w_n7265_21[0]),.dout(n7624),.clk(gclk));
	jxor g07367(.dina(n7624),.dinb(w_n7239_0[0]),.dout(n7625),.clk(gclk));
	jand g07368(.dina(w_asqrt27_15[2]),.dinb(w_n7253_0[1]),.dout(n7626),.clk(gclk));
	jand g07369(.dina(w_n7626_0[1]),.dinb(w_n7241_1[0]),.dout(n7627),.clk(gclk));
	jor g07370(.dina(n7627),.dinb(w_n7288_0[0]),.dout(n7628),.clk(gclk));
	jor g07371(.dina(n7628),.dinb(w_n7625_0[2]),.dout(n7629),.clk(gclk));
	jor g07372(.dina(n7629),.dinb(w_n7621_0[2]),.dout(n7630),.clk(gclk));
	jand g07373(.dina(n7630),.dinb(w_n194_27[1]),.dout(n7631),.clk(gclk));
	jand g07374(.dina(w_n7625_0[1]),.dinb(w_n7621_0[1]),.dout(n7632),.clk(gclk));
	jor g07375(.dina(w_n7626_0[0]),.dinb(w_n7241_0[2]),.dout(n7633),.clk(gclk));
	jand g07376(.dina(w_n7253_0[0]),.dinb(w_n7241_0[1]),.dout(n7634),.clk(gclk));
	jor g07377(.dina(n7634),.dinb(w_n194_27[0]),.dout(n7635),.clk(gclk));
	jnot g07378(.din(n7635),.dout(n7636),.clk(gclk));
	jand g07379(.dina(n7636),.dinb(n7633),.dout(n7637),.clk(gclk));
	jor g07380(.dina(w_n7637_0[1]),.dinb(w_n7632_0[2]),.dout(n7640),.clk(gclk));
	jor g07381(.dina(n7640),.dinb(w_n7631_0[1]),.dout(asqrt_fa_27),.clk(gclk));
	jxor g07382(.dina(w_n7355_0[0]),.dinb(w_n4494_18[1]),.dout(n7642),.clk(gclk));
	jand g07383(.dina(n7642),.dinb(w_asqrt26_31),.dout(n7643),.clk(gclk));
	jxor g07384(.dina(n7643),.dinb(w_n7269_0[0]),.dout(n7644),.clk(gclk));
	jnot g07385(.din(n7644),.dout(n7645),.clk(gclk));
	jand g07386(.dina(w_asqrt26_30[2]),.dinb(w_a52_0[0]),.dout(n7646),.clk(gclk));
	jnot g07387(.din(w_a50_0[1]),.dout(n7647),.clk(gclk));
	jnot g07388(.din(w_a51_0[1]),.dout(n7648),.clk(gclk));
	jand g07389(.dina(w_n7271_1[0]),.dinb(w_n7648_0[1]),.dout(n7649),.clk(gclk));
	jand g07390(.dina(n7649),.dinb(w_n7647_1[1]),.dout(n7650),.clk(gclk));
	jor g07391(.dina(n7650),.dinb(n7646),.dout(n7651),.clk(gclk));
	jand g07392(.dina(w_n7651_0[2]),.dinb(w_asqrt27_15[1]),.dout(n7652),.clk(gclk));
	jand g07393(.dina(w_asqrt26_30[1]),.dinb(w_n7271_0[2]),.dout(n7653),.clk(gclk));
	jxor g07394(.dina(w_n7653_0[1]),.dinb(w_n7272_0[1]),.dout(n7654),.clk(gclk));
	jor g07395(.dina(w_n7651_0[1]),.dinb(w_asqrt27_15[0]),.dout(n7655),.clk(gclk));
	jand g07396(.dina(n7655),.dinb(w_n7654_0[1]),.dout(n7656),.clk(gclk));
	jor g07397(.dina(w_n7656_0[1]),.dinb(w_n7652_0[1]),.dout(n7657),.clk(gclk));
	jand g07398(.dina(n7657),.dinb(w_asqrt28_18[2]),.dout(n7658),.clk(gclk));
	jor g07399(.dina(w_n7652_0[0]),.dinb(w_asqrt28_18[1]),.dout(n7659),.clk(gclk));
	jor g07400(.dina(n7659),.dinb(w_n7656_0[0]),.dout(n7660),.clk(gclk));
	jand g07401(.dina(w_n7653_0[0]),.dinb(w_n7272_0[0]),.dout(n7661),.clk(gclk));
	jnot g07402(.din(w_n7631_0[0]),.dout(n7662),.clk(gclk));
	jnot g07403(.din(w_n7632_0[1]),.dout(n7663),.clk(gclk));
	jnot g07404(.din(w_n7637_0[0]),.dout(n7664),.clk(gclk));
	jand g07405(.dina(n7664),.dinb(w_asqrt27_14[2]),.dout(n7665),.clk(gclk));
	jand g07406(.dina(n7665),.dinb(n7663),.dout(n7666),.clk(gclk));
	jand g07407(.dina(n7666),.dinb(n7662),.dout(n7667),.clk(gclk));
	jor g07408(.dina(n7667),.dinb(n7661),.dout(n7668),.clk(gclk));
	jxor g07409(.dina(n7668),.dinb(w_n6872_0[1]),.dout(n7669),.clk(gclk));
	jand g07410(.dina(w_n7669_0[1]),.dinb(w_n7660_0[1]),.dout(n7670),.clk(gclk));
	jor g07411(.dina(n7670),.dinb(w_n7658_0[1]),.dout(n7671),.clk(gclk));
	jand g07412(.dina(w_n7671_0[2]),.dinb(w_asqrt29_15[1]),.dout(n7672),.clk(gclk));
	jor g07413(.dina(w_n7671_0[1]),.dinb(w_asqrt29_15[0]),.dout(n7673),.clk(gclk));
	jxor g07414(.dina(w_n7276_0[0]),.dinb(w_n7260_17[1]),.dout(n7674),.clk(gclk));
	jand g07415(.dina(n7674),.dinb(w_asqrt26_30[0]),.dout(n7675),.clk(gclk));
	jxor g07416(.dina(n7675),.dinb(w_n7279_0[0]),.dout(n7676),.clk(gclk));
	jnot g07417(.din(w_n7676_0[1]),.dout(n7677),.clk(gclk));
	jand g07418(.dina(n7677),.dinb(n7673),.dout(n7678),.clk(gclk));
	jor g07419(.dina(w_n7678_0[1]),.dinb(w_n7672_0[1]),.dout(n7679),.clk(gclk));
	jand g07420(.dina(n7679),.dinb(w_asqrt30_18[2]),.dout(n7680),.clk(gclk));
	jnot g07421(.din(w_n7285_0[0]),.dout(n7681),.clk(gclk));
	jand g07422(.dina(n7681),.dinb(w_n7283_0[0]),.dout(n7682),.clk(gclk));
	jand g07423(.dina(n7682),.dinb(w_asqrt26_29[2]),.dout(n7683),.clk(gclk));
	jxor g07424(.dina(n7683),.dinb(w_n7293_0[0]),.dout(n7684),.clk(gclk));
	jnot g07425(.din(n7684),.dout(n7685),.clk(gclk));
	jor g07426(.dina(w_n7672_0[0]),.dinb(w_asqrt30_18[1]),.dout(n7686),.clk(gclk));
	jor g07427(.dina(n7686),.dinb(w_n7678_0[0]),.dout(n7687),.clk(gclk));
	jand g07428(.dina(w_n7687_0[1]),.dinb(w_n7685_0[1]),.dout(n7688),.clk(gclk));
	jor g07429(.dina(w_n7688_0[1]),.dinb(w_n7680_0[1]),.dout(n7689),.clk(gclk));
	jand g07430(.dina(w_n7689_0[2]),.dinb(w_asqrt31_15[1]),.dout(n7690),.clk(gclk));
	jor g07431(.dina(w_n7689_0[1]),.dinb(w_asqrt31_15[0]),.dout(n7691),.clk(gclk));
	jnot g07432(.din(w_n7300_0[0]),.dout(n7692),.clk(gclk));
	jxor g07433(.dina(w_n7295_0[0]),.dinb(w_n6500_17[1]),.dout(n7693),.clk(gclk));
	jand g07434(.dina(n7693),.dinb(w_asqrt26_29[1]),.dout(n7694),.clk(gclk));
	jxor g07435(.dina(n7694),.dinb(n7692),.dout(n7695),.clk(gclk));
	jand g07436(.dina(w_n7695_0[1]),.dinb(n7691),.dout(n7696),.clk(gclk));
	jor g07437(.dina(w_n7696_0[1]),.dinb(w_n7690_0[1]),.dout(n7697),.clk(gclk));
	jand g07438(.dina(n7697),.dinb(w_asqrt32_18[2]),.dout(n7698),.clk(gclk));
	jor g07439(.dina(w_n7690_0[0]),.dinb(w_asqrt32_18[1]),.dout(n7699),.clk(gclk));
	jor g07440(.dina(n7699),.dinb(w_n7696_0[0]),.dout(n7700),.clk(gclk));
	jnot g07441(.din(w_n7307_0[0]),.dout(n7701),.clk(gclk));
	jnot g07442(.din(w_n7309_0[0]),.dout(n7702),.clk(gclk));
	jand g07443(.dina(w_asqrt26_29[0]),.dinb(w_n7303_0[0]),.dout(n7703),.clk(gclk));
	jand g07444(.dina(w_n7703_0[1]),.dinb(n7702),.dout(n7704),.clk(gclk));
	jor g07445(.dina(n7704),.dinb(n7701),.dout(n7705),.clk(gclk));
	jnot g07446(.din(w_n7310_0[0]),.dout(n7706),.clk(gclk));
	jand g07447(.dina(w_n7703_0[0]),.dinb(n7706),.dout(n7707),.clk(gclk));
	jnot g07448(.din(n7707),.dout(n7708),.clk(gclk));
	jand g07449(.dina(n7708),.dinb(n7705),.dout(n7709),.clk(gclk));
	jand g07450(.dina(w_n7709_0[1]),.dinb(w_n7700_0[1]),.dout(n7710),.clk(gclk));
	jor g07451(.dina(n7710),.dinb(w_n7698_0[1]),.dout(n7711),.clk(gclk));
	jand g07452(.dina(w_n7711_0[2]),.dinb(w_asqrt33_15[2]),.dout(n7712),.clk(gclk));
	jor g07453(.dina(w_n7711_0[1]),.dinb(w_asqrt33_15[1]),.dout(n7713),.clk(gclk));
	jxor g07454(.dina(w_n7311_0[0]),.dinb(w_n5788_17[2]),.dout(n7714),.clk(gclk));
	jand g07455(.dina(n7714),.dinb(w_asqrt26_28[2]),.dout(n7715),.clk(gclk));
	jxor g07456(.dina(n7715),.dinb(w_n7316_0[0]),.dout(n7716),.clk(gclk));
	jand g07457(.dina(w_n7716_0[1]),.dinb(n7713),.dout(n7717),.clk(gclk));
	jor g07458(.dina(w_n7717_0[1]),.dinb(w_n7712_0[1]),.dout(n7718),.clk(gclk));
	jand g07459(.dina(n7718),.dinb(w_asqrt34_18[2]),.dout(n7719),.clk(gclk));
	jnot g07460(.din(w_n7322_0[0]),.dout(n7720),.clk(gclk));
	jand g07461(.dina(n7720),.dinb(w_n7320_0[0]),.dout(n7721),.clk(gclk));
	jand g07462(.dina(n7721),.dinb(w_asqrt26_28[1]),.dout(n7722),.clk(gclk));
	jxor g07463(.dina(n7722),.dinb(w_n7331_0[0]),.dout(n7723),.clk(gclk));
	jnot g07464(.din(n7723),.dout(n7724),.clk(gclk));
	jor g07465(.dina(w_n7712_0[0]),.dinb(w_asqrt34_18[1]),.dout(n7725),.clk(gclk));
	jor g07466(.dina(n7725),.dinb(w_n7717_0[0]),.dout(n7726),.clk(gclk));
	jand g07467(.dina(w_n7726_0[1]),.dinb(w_n7724_0[1]),.dout(n7727),.clk(gclk));
	jor g07468(.dina(w_n7727_0[1]),.dinb(w_n7719_0[1]),.dout(n7728),.clk(gclk));
	jand g07469(.dina(w_n7728_0[2]),.dinb(w_asqrt35_15[2]),.dout(n7729),.clk(gclk));
	jor g07470(.dina(w_n7728_0[1]),.dinb(w_asqrt35_15[1]),.dout(n7730),.clk(gclk));
	jxor g07471(.dina(w_n7333_0[0]),.dinb(w_n5116_17[2]),.dout(n7731),.clk(gclk));
	jand g07472(.dina(n7731),.dinb(w_asqrt26_28[0]),.dout(n7732),.clk(gclk));
	jxor g07473(.dina(n7732),.dinb(w_n7339_0[0]),.dout(n7733),.clk(gclk));
	jand g07474(.dina(w_n7733_0[1]),.dinb(n7730),.dout(n7734),.clk(gclk));
	jor g07475(.dina(w_n7734_0[1]),.dinb(w_n7729_0[1]),.dout(n7735),.clk(gclk));
	jand g07476(.dina(n7735),.dinb(w_asqrt36_18[2]),.dout(n7736),.clk(gclk));
	jnot g07477(.din(w_n7345_0[0]),.dout(n7737),.clk(gclk));
	jand g07478(.dina(n7737),.dinb(w_n7343_0[0]),.dout(n7738),.clk(gclk));
	jand g07479(.dina(n7738),.dinb(w_asqrt26_27[2]),.dout(n7739),.clk(gclk));
	jxor g07480(.dina(n7739),.dinb(w_n7353_0[0]),.dout(n7740),.clk(gclk));
	jnot g07481(.din(n7740),.dout(n7741),.clk(gclk));
	jor g07482(.dina(w_n7729_0[0]),.dinb(w_asqrt36_18[1]),.dout(n7742),.clk(gclk));
	jor g07483(.dina(n7742),.dinb(w_n7734_0[0]),.dout(n7743),.clk(gclk));
	jand g07484(.dina(w_n7743_0[1]),.dinb(w_n7741_0[1]),.dout(n7744),.clk(gclk));
	jor g07485(.dina(w_n7744_0[1]),.dinb(w_n7736_0[1]),.dout(n7745),.clk(gclk));
	jand g07486(.dina(w_n7745_0[2]),.dinb(w_asqrt37_16[0]),.dout(n7746),.clk(gclk));
	jor g07487(.dina(w_n7745_0[1]),.dinb(w_asqrt37_15[2]),.dout(n7747),.clk(gclk));
	jand g07488(.dina(n7747),.dinb(w_n7645_0[1]),.dout(n7748),.clk(gclk));
	jor g07489(.dina(w_n7748_0[1]),.dinb(w_n7746_0[1]),.dout(n7749),.clk(gclk));
	jand g07490(.dina(n7749),.dinb(w_asqrt38_18[2]),.dout(n7750),.clk(gclk));
	jor g07491(.dina(w_n7746_0[0]),.dinb(w_asqrt38_18[1]),.dout(n7751),.clk(gclk));
	jor g07492(.dina(n7751),.dinb(w_n7748_0[0]),.dout(n7752),.clk(gclk));
	jnot g07493(.din(w_n7364_0[0]),.dout(n7753),.clk(gclk));
	jnot g07494(.din(w_n7366_0[0]),.dout(n7754),.clk(gclk));
	jand g07495(.dina(w_asqrt26_27[1]),.dinb(w_n7360_0[0]),.dout(n7755),.clk(gclk));
	jand g07496(.dina(w_n7755_0[1]),.dinb(n7754),.dout(n7756),.clk(gclk));
	jor g07497(.dina(n7756),.dinb(n7753),.dout(n7757),.clk(gclk));
	jnot g07498(.din(w_n7367_0[0]),.dout(n7758),.clk(gclk));
	jand g07499(.dina(w_n7755_0[0]),.dinb(n7758),.dout(n7759),.clk(gclk));
	jnot g07500(.din(n7759),.dout(n7760),.clk(gclk));
	jand g07501(.dina(n7760),.dinb(n7757),.dout(n7761),.clk(gclk));
	jand g07502(.dina(w_n7761_0[1]),.dinb(w_n7752_0[1]),.dout(n7762),.clk(gclk));
	jor g07503(.dina(n7762),.dinb(w_n7750_0[1]),.dout(n7763),.clk(gclk));
	jand g07504(.dina(w_n7763_0[2]),.dinb(w_asqrt39_16[0]),.dout(n7764),.clk(gclk));
	jor g07505(.dina(w_n7763_0[1]),.dinb(w_asqrt39_15[2]),.dout(n7765),.clk(gclk));
	jnot g07506(.din(w_n7372_0[0]),.dout(n7766),.clk(gclk));
	jnot g07507(.din(w_n7373_0[0]),.dout(n7767),.clk(gclk));
	jand g07508(.dina(w_asqrt26_27[0]),.dinb(w_n7369_0[0]),.dout(n7768),.clk(gclk));
	jand g07509(.dina(w_n7768_0[1]),.dinb(n7767),.dout(n7769),.clk(gclk));
	jor g07510(.dina(n7769),.dinb(n7766),.dout(n7770),.clk(gclk));
	jnot g07511(.din(w_n7374_0[0]),.dout(n7771),.clk(gclk));
	jand g07512(.dina(w_n7768_0[0]),.dinb(n7771),.dout(n7772),.clk(gclk));
	jnot g07513(.din(n7772),.dout(n7773),.clk(gclk));
	jand g07514(.dina(n7773),.dinb(n7770),.dout(n7774),.clk(gclk));
	jand g07515(.dina(w_n7774_0[1]),.dinb(n7765),.dout(n7775),.clk(gclk));
	jor g07516(.dina(w_n7775_0[1]),.dinb(w_n7764_0[1]),.dout(n7776),.clk(gclk));
	jand g07517(.dina(n7776),.dinb(w_asqrt40_18[2]),.dout(n7777),.clk(gclk));
	jor g07518(.dina(w_n7764_0[0]),.dinb(w_asqrt40_18[1]),.dout(n7778),.clk(gclk));
	jor g07519(.dina(n7778),.dinb(w_n7775_0[0]),.dout(n7779),.clk(gclk));
	jnot g07520(.din(w_n7380_0[0]),.dout(n7780),.clk(gclk));
	jnot g07521(.din(w_n7382_0[0]),.dout(n7781),.clk(gclk));
	jand g07522(.dina(w_asqrt26_26[2]),.dinb(w_n7376_0[0]),.dout(n7782),.clk(gclk));
	jand g07523(.dina(w_n7782_0[1]),.dinb(n7781),.dout(n7783),.clk(gclk));
	jor g07524(.dina(n7783),.dinb(n7780),.dout(n7784),.clk(gclk));
	jnot g07525(.din(w_n7383_0[0]),.dout(n7785),.clk(gclk));
	jand g07526(.dina(w_n7782_0[0]),.dinb(n7785),.dout(n7786),.clk(gclk));
	jnot g07527(.din(n7786),.dout(n7787),.clk(gclk));
	jand g07528(.dina(n7787),.dinb(n7784),.dout(n7788),.clk(gclk));
	jand g07529(.dina(w_n7788_0[1]),.dinb(w_n7779_0[1]),.dout(n7789),.clk(gclk));
	jor g07530(.dina(n7789),.dinb(w_n7777_0[1]),.dout(n7790),.clk(gclk));
	jand g07531(.dina(w_n7790_0[1]),.dinb(w_asqrt41_16[1]),.dout(n7791),.clk(gclk));
	jxor g07532(.dina(w_n7384_0[0]),.dinb(w_n3371_19[0]),.dout(n7792),.clk(gclk));
	jand g07533(.dina(n7792),.dinb(w_asqrt26_26[1]),.dout(n7793),.clk(gclk));
	jxor g07534(.dina(n7793),.dinb(w_n7394_0[0]),.dout(n7794),.clk(gclk));
	jnot g07535(.din(n7794),.dout(n7795),.clk(gclk));
	jor g07536(.dina(w_n7790_0[0]),.dinb(w_asqrt41_16[0]),.dout(n7796),.clk(gclk));
	jand g07537(.dina(w_n7796_0[1]),.dinb(w_n7795_0[1]),.dout(n7797),.clk(gclk));
	jor g07538(.dina(w_n7797_0[2]),.dinb(w_n7791_0[2]),.dout(n7798),.clk(gclk));
	jand g07539(.dina(n7798),.dinb(w_asqrt42_18[2]),.dout(n7799),.clk(gclk));
	jnot g07540(.din(w_n7399_0[0]),.dout(n7800),.clk(gclk));
	jand g07541(.dina(n7800),.dinb(w_n7397_0[0]),.dout(n7801),.clk(gclk));
	jand g07542(.dina(n7801),.dinb(w_asqrt26_26[0]),.dout(n7802),.clk(gclk));
	jxor g07543(.dina(n7802),.dinb(w_n7407_0[0]),.dout(n7803),.clk(gclk));
	jnot g07544(.din(n7803),.dout(n7804),.clk(gclk));
	jor g07545(.dina(w_n7791_0[1]),.dinb(w_asqrt42_18[1]),.dout(n7805),.clk(gclk));
	jor g07546(.dina(n7805),.dinb(w_n7797_0[1]),.dout(n7806),.clk(gclk));
	jand g07547(.dina(w_n7806_0[1]),.dinb(w_n7804_0[1]),.dout(n7807),.clk(gclk));
	jor g07548(.dina(w_n7807_0[1]),.dinb(w_n7799_0[1]),.dout(n7808),.clk(gclk));
	jand g07549(.dina(w_n7808_0[2]),.dinb(w_asqrt43_16[1]),.dout(n7809),.clk(gclk));
	jor g07550(.dina(w_n7808_0[1]),.dinb(w_asqrt43_16[0]),.dout(n7810),.clk(gclk));
	jnot g07551(.din(w_n7413_0[0]),.dout(n7811),.clk(gclk));
	jnot g07552(.din(w_n7414_0[0]),.dout(n7812),.clk(gclk));
	jand g07553(.dina(w_asqrt26_25[2]),.dinb(w_n7410_0[0]),.dout(n7813),.clk(gclk));
	jand g07554(.dina(w_n7813_0[1]),.dinb(n7812),.dout(n7814),.clk(gclk));
	jor g07555(.dina(n7814),.dinb(n7811),.dout(n7815),.clk(gclk));
	jnot g07556(.din(w_n7415_0[0]),.dout(n7816),.clk(gclk));
	jand g07557(.dina(w_n7813_0[0]),.dinb(n7816),.dout(n7817),.clk(gclk));
	jnot g07558(.din(n7817),.dout(n7818),.clk(gclk));
	jand g07559(.dina(n7818),.dinb(n7815),.dout(n7819),.clk(gclk));
	jand g07560(.dina(w_n7819_0[1]),.dinb(n7810),.dout(n7820),.clk(gclk));
	jor g07561(.dina(w_n7820_0[1]),.dinb(w_n7809_0[1]),.dout(n7821),.clk(gclk));
	jand g07562(.dina(n7821),.dinb(w_asqrt44_18[2]),.dout(n7822),.clk(gclk));
	jor g07563(.dina(w_n7809_0[0]),.dinb(w_asqrt44_18[1]),.dout(n7823),.clk(gclk));
	jor g07564(.dina(n7823),.dinb(w_n7820_0[0]),.dout(n7824),.clk(gclk));
	jnot g07565(.din(w_n7421_0[0]),.dout(n7825),.clk(gclk));
	jnot g07566(.din(w_n7423_0[0]),.dout(n7826),.clk(gclk));
	jand g07567(.dina(w_asqrt26_25[1]),.dinb(w_n7417_0[0]),.dout(n7827),.clk(gclk));
	jand g07568(.dina(w_n7827_0[1]),.dinb(n7826),.dout(n7828),.clk(gclk));
	jor g07569(.dina(n7828),.dinb(n7825),.dout(n7829),.clk(gclk));
	jnot g07570(.din(w_n7424_0[0]),.dout(n7830),.clk(gclk));
	jand g07571(.dina(w_n7827_0[0]),.dinb(n7830),.dout(n7831),.clk(gclk));
	jnot g07572(.din(n7831),.dout(n7832),.clk(gclk));
	jand g07573(.dina(n7832),.dinb(n7829),.dout(n7833),.clk(gclk));
	jand g07574(.dina(w_n7833_0[1]),.dinb(w_n7824_0[1]),.dout(n7834),.clk(gclk));
	jor g07575(.dina(n7834),.dinb(w_n7822_0[1]),.dout(n7835),.clk(gclk));
	jand g07576(.dina(w_n7835_0[1]),.dinb(w_asqrt45_16[2]),.dout(n7836),.clk(gclk));
	jxor g07577(.dina(w_n7425_0[0]),.dinb(w_n2420_20[0]),.dout(n7837),.clk(gclk));
	jand g07578(.dina(n7837),.dinb(w_asqrt26_25[0]),.dout(n7838),.clk(gclk));
	jxor g07579(.dina(n7838),.dinb(w_n7435_0[0]),.dout(n7839),.clk(gclk));
	jnot g07580(.din(n7839),.dout(n7840),.clk(gclk));
	jor g07581(.dina(w_n7835_0[0]),.dinb(w_asqrt45_16[1]),.dout(n7841),.clk(gclk));
	jand g07582(.dina(w_n7841_0[1]),.dinb(w_n7840_0[1]),.dout(n7842),.clk(gclk));
	jor g07583(.dina(w_n7842_0[2]),.dinb(w_n7836_0[2]),.dout(n7843),.clk(gclk));
	jand g07584(.dina(n7843),.dinb(w_asqrt46_18[2]),.dout(n7844),.clk(gclk));
	jnot g07585(.din(w_n7440_0[0]),.dout(n7845),.clk(gclk));
	jand g07586(.dina(n7845),.dinb(w_n7438_0[0]),.dout(n7846),.clk(gclk));
	jand g07587(.dina(n7846),.dinb(w_asqrt26_24[2]),.dout(n7847),.clk(gclk));
	jxor g07588(.dina(n7847),.dinb(w_n7448_0[0]),.dout(n7848),.clk(gclk));
	jnot g07589(.din(n7848),.dout(n7849),.clk(gclk));
	jor g07590(.dina(w_n7836_0[1]),.dinb(w_asqrt46_18[1]),.dout(n7850),.clk(gclk));
	jor g07591(.dina(n7850),.dinb(w_n7842_0[1]),.dout(n7851),.clk(gclk));
	jand g07592(.dina(w_n7851_0[1]),.dinb(w_n7849_0[1]),.dout(n7852),.clk(gclk));
	jor g07593(.dina(w_n7852_0[1]),.dinb(w_n7844_0[1]),.dout(n7853),.clk(gclk));
	jand g07594(.dina(w_n7853_0[2]),.dinb(w_asqrt47_16[2]),.dout(n7854),.clk(gclk));
	jor g07595(.dina(w_n7853_0[1]),.dinb(w_asqrt47_16[1]),.dout(n7855),.clk(gclk));
	jnot g07596(.din(w_n7454_0[0]),.dout(n7856),.clk(gclk));
	jnot g07597(.din(w_n7455_0[0]),.dout(n7857),.clk(gclk));
	jand g07598(.dina(w_asqrt26_24[1]),.dinb(w_n7451_0[0]),.dout(n7858),.clk(gclk));
	jand g07599(.dina(w_n7858_0[1]),.dinb(n7857),.dout(n7859),.clk(gclk));
	jor g07600(.dina(n7859),.dinb(n7856),.dout(n7860),.clk(gclk));
	jnot g07601(.din(w_n7456_0[0]),.dout(n7861),.clk(gclk));
	jand g07602(.dina(w_n7858_0[0]),.dinb(n7861),.dout(n7862),.clk(gclk));
	jnot g07603(.din(n7862),.dout(n7863),.clk(gclk));
	jand g07604(.dina(n7863),.dinb(n7860),.dout(n7864),.clk(gclk));
	jand g07605(.dina(w_n7864_0[1]),.dinb(n7855),.dout(n7865),.clk(gclk));
	jor g07606(.dina(w_n7865_0[1]),.dinb(w_n7854_0[1]),.dout(n7866),.clk(gclk));
	jand g07607(.dina(n7866),.dinb(w_asqrt48_18[2]),.dout(n7867),.clk(gclk));
	jor g07608(.dina(w_n7854_0[0]),.dinb(w_asqrt48_18[1]),.dout(n7868),.clk(gclk));
	jor g07609(.dina(n7868),.dinb(w_n7865_0[0]),.dout(n7869),.clk(gclk));
	jnot g07610(.din(w_n7462_0[0]),.dout(n7870),.clk(gclk));
	jnot g07611(.din(w_n7464_0[0]),.dout(n7871),.clk(gclk));
	jand g07612(.dina(w_asqrt26_24[0]),.dinb(w_n7458_0[0]),.dout(n7872),.clk(gclk));
	jand g07613(.dina(w_n7872_0[1]),.dinb(n7871),.dout(n7873),.clk(gclk));
	jor g07614(.dina(n7873),.dinb(n7870),.dout(n7874),.clk(gclk));
	jnot g07615(.din(w_n7465_0[0]),.dout(n7875),.clk(gclk));
	jand g07616(.dina(w_n7872_0[0]),.dinb(n7875),.dout(n7876),.clk(gclk));
	jnot g07617(.din(n7876),.dout(n7877),.clk(gclk));
	jand g07618(.dina(n7877),.dinb(n7874),.dout(n7878),.clk(gclk));
	jand g07619(.dina(w_n7878_0[1]),.dinb(w_n7869_0[1]),.dout(n7879),.clk(gclk));
	jor g07620(.dina(n7879),.dinb(w_n7867_0[1]),.dout(n7880),.clk(gclk));
	jand g07621(.dina(w_n7880_0[1]),.dinb(w_asqrt49_17[0]),.dout(n7881),.clk(gclk));
	jxor g07622(.dina(w_n7466_0[0]),.dinb(w_n1641_20[2]),.dout(n7882),.clk(gclk));
	jand g07623(.dina(n7882),.dinb(w_asqrt26_23[2]),.dout(n7883),.clk(gclk));
	jxor g07624(.dina(n7883),.dinb(w_n7476_0[0]),.dout(n7884),.clk(gclk));
	jnot g07625(.din(n7884),.dout(n7885),.clk(gclk));
	jor g07626(.dina(w_n7880_0[0]),.dinb(w_asqrt49_16[2]),.dout(n7886),.clk(gclk));
	jand g07627(.dina(w_n7886_0[1]),.dinb(w_n7885_0[1]),.dout(n7887),.clk(gclk));
	jor g07628(.dina(w_n7887_0[2]),.dinb(w_n7881_0[2]),.dout(n7888),.clk(gclk));
	jand g07629(.dina(n7888),.dinb(w_asqrt50_18[2]),.dout(n7889),.clk(gclk));
	jnot g07630(.din(w_n7481_0[0]),.dout(n7890),.clk(gclk));
	jand g07631(.dina(n7890),.dinb(w_n7479_0[0]),.dout(n7891),.clk(gclk));
	jand g07632(.dina(n7891),.dinb(w_asqrt26_23[1]),.dout(n7892),.clk(gclk));
	jxor g07633(.dina(n7892),.dinb(w_n7489_0[0]),.dout(n7893),.clk(gclk));
	jnot g07634(.din(n7893),.dout(n7894),.clk(gclk));
	jor g07635(.dina(w_n7881_0[1]),.dinb(w_asqrt50_18[1]),.dout(n7895),.clk(gclk));
	jor g07636(.dina(n7895),.dinb(w_n7887_0[1]),.dout(n7896),.clk(gclk));
	jand g07637(.dina(w_n7896_0[1]),.dinb(w_n7894_0[1]),.dout(n7897),.clk(gclk));
	jor g07638(.dina(w_n7897_0[1]),.dinb(w_n7889_0[1]),.dout(n7898),.clk(gclk));
	jand g07639(.dina(w_n7898_0[2]),.dinb(w_asqrt51_17[0]),.dout(n7899),.clk(gclk));
	jor g07640(.dina(w_n7898_0[1]),.dinb(w_asqrt51_16[2]),.dout(n7900),.clk(gclk));
	jnot g07641(.din(w_n7495_0[0]),.dout(n7901),.clk(gclk));
	jnot g07642(.din(w_n7496_0[0]),.dout(n7902),.clk(gclk));
	jand g07643(.dina(w_asqrt26_23[0]),.dinb(w_n7492_0[0]),.dout(n7903),.clk(gclk));
	jand g07644(.dina(w_n7903_0[1]),.dinb(n7902),.dout(n7904),.clk(gclk));
	jor g07645(.dina(n7904),.dinb(n7901),.dout(n7905),.clk(gclk));
	jnot g07646(.din(w_n7497_0[0]),.dout(n7906),.clk(gclk));
	jand g07647(.dina(w_n7903_0[0]),.dinb(n7906),.dout(n7907),.clk(gclk));
	jnot g07648(.din(n7907),.dout(n7908),.clk(gclk));
	jand g07649(.dina(n7908),.dinb(n7905),.dout(n7909),.clk(gclk));
	jand g07650(.dina(w_n7909_0[1]),.dinb(n7900),.dout(n7910),.clk(gclk));
	jor g07651(.dina(w_n7910_0[1]),.dinb(w_n7899_0[1]),.dout(n7911),.clk(gclk));
	jand g07652(.dina(n7911),.dinb(w_asqrt52_18[2]),.dout(n7912),.clk(gclk));
	jor g07653(.dina(w_n7899_0[0]),.dinb(w_asqrt52_18[1]),.dout(n7913),.clk(gclk));
	jor g07654(.dina(n7913),.dinb(w_n7910_0[0]),.dout(n7914),.clk(gclk));
	jnot g07655(.din(w_n7503_0[0]),.dout(n7915),.clk(gclk));
	jnot g07656(.din(w_n7505_0[0]),.dout(n7916),.clk(gclk));
	jand g07657(.dina(w_asqrt26_22[2]),.dinb(w_n7499_0[0]),.dout(n7917),.clk(gclk));
	jand g07658(.dina(w_n7917_0[1]),.dinb(n7916),.dout(n7918),.clk(gclk));
	jor g07659(.dina(n7918),.dinb(n7915),.dout(n7919),.clk(gclk));
	jnot g07660(.din(w_n7506_0[0]),.dout(n7920),.clk(gclk));
	jand g07661(.dina(w_n7917_0[0]),.dinb(n7920),.dout(n7921),.clk(gclk));
	jnot g07662(.din(n7921),.dout(n7922),.clk(gclk));
	jand g07663(.dina(n7922),.dinb(n7919),.dout(n7923),.clk(gclk));
	jand g07664(.dina(w_n7923_0[1]),.dinb(w_n7914_0[1]),.dout(n7924),.clk(gclk));
	jor g07665(.dina(n7924),.dinb(w_n7912_0[1]),.dout(n7925),.clk(gclk));
	jand g07666(.dina(w_n7925_0[1]),.dinb(w_asqrt53_17[1]),.dout(n7926),.clk(gclk));
	jxor g07667(.dina(w_n7507_0[0]),.dinb(w_n1034_21[2]),.dout(n7927),.clk(gclk));
	jand g07668(.dina(n7927),.dinb(w_asqrt26_22[1]),.dout(n7928),.clk(gclk));
	jxor g07669(.dina(n7928),.dinb(w_n7517_0[0]),.dout(n7929),.clk(gclk));
	jnot g07670(.din(n7929),.dout(n7930),.clk(gclk));
	jor g07671(.dina(w_n7925_0[0]),.dinb(w_asqrt53_17[0]),.dout(n7931),.clk(gclk));
	jand g07672(.dina(w_n7931_0[1]),.dinb(w_n7930_0[1]),.dout(n7932),.clk(gclk));
	jor g07673(.dina(w_n7932_0[2]),.dinb(w_n7926_0[2]),.dout(n7933),.clk(gclk));
	jand g07674(.dina(n7933),.dinb(w_asqrt54_18[2]),.dout(n7934),.clk(gclk));
	jnot g07675(.din(w_n7522_0[0]),.dout(n7935),.clk(gclk));
	jand g07676(.dina(n7935),.dinb(w_n7520_0[0]),.dout(n7936),.clk(gclk));
	jand g07677(.dina(n7936),.dinb(w_asqrt26_22[0]),.dout(n7937),.clk(gclk));
	jxor g07678(.dina(n7937),.dinb(w_n7530_0[0]),.dout(n7938),.clk(gclk));
	jnot g07679(.din(n7938),.dout(n7939),.clk(gclk));
	jor g07680(.dina(w_n7926_0[1]),.dinb(w_asqrt54_18[1]),.dout(n7940),.clk(gclk));
	jor g07681(.dina(n7940),.dinb(w_n7932_0[1]),.dout(n7941),.clk(gclk));
	jand g07682(.dina(w_n7941_0[1]),.dinb(w_n7939_0[1]),.dout(n7942),.clk(gclk));
	jor g07683(.dina(w_n7942_0[1]),.dinb(w_n7934_0[1]),.dout(n7943),.clk(gclk));
	jand g07684(.dina(w_n7943_0[2]),.dinb(w_asqrt55_17[2]),.dout(n7944),.clk(gclk));
	jor g07685(.dina(w_n7943_0[1]),.dinb(w_asqrt55_17[1]),.dout(n7945),.clk(gclk));
	jnot g07686(.din(w_n7536_0[0]),.dout(n7946),.clk(gclk));
	jnot g07687(.din(w_n7537_0[0]),.dout(n7947),.clk(gclk));
	jand g07688(.dina(w_asqrt26_21[2]),.dinb(w_n7533_0[0]),.dout(n7948),.clk(gclk));
	jand g07689(.dina(w_n7948_0[1]),.dinb(n7947),.dout(n7949),.clk(gclk));
	jor g07690(.dina(n7949),.dinb(n7946),.dout(n7950),.clk(gclk));
	jnot g07691(.din(w_n7538_0[0]),.dout(n7951),.clk(gclk));
	jand g07692(.dina(w_n7948_0[0]),.dinb(n7951),.dout(n7952),.clk(gclk));
	jnot g07693(.din(n7952),.dout(n7953),.clk(gclk));
	jand g07694(.dina(n7953),.dinb(n7950),.dout(n7954),.clk(gclk));
	jand g07695(.dina(w_n7954_0[1]),.dinb(n7945),.dout(n7955),.clk(gclk));
	jor g07696(.dina(w_n7955_0[1]),.dinb(w_n7944_0[1]),.dout(n7956),.clk(gclk));
	jand g07697(.dina(n7956),.dinb(w_asqrt56_18[2]),.dout(n7957),.clk(gclk));
	jor g07698(.dina(w_n7944_0[0]),.dinb(w_asqrt56_18[1]),.dout(n7958),.clk(gclk));
	jor g07699(.dina(n7958),.dinb(w_n7955_0[0]),.dout(n7959),.clk(gclk));
	jnot g07700(.din(w_n7544_0[0]),.dout(n7960),.clk(gclk));
	jnot g07701(.din(w_n7546_0[0]),.dout(n7961),.clk(gclk));
	jand g07702(.dina(w_asqrt26_21[1]),.dinb(w_n7540_0[0]),.dout(n7962),.clk(gclk));
	jand g07703(.dina(w_n7962_0[1]),.dinb(n7961),.dout(n7963),.clk(gclk));
	jor g07704(.dina(n7963),.dinb(n7960),.dout(n7964),.clk(gclk));
	jnot g07705(.din(w_n7547_0[0]),.dout(n7965),.clk(gclk));
	jand g07706(.dina(w_n7962_0[0]),.dinb(n7965),.dout(n7966),.clk(gclk));
	jnot g07707(.din(n7966),.dout(n7967),.clk(gclk));
	jand g07708(.dina(n7967),.dinb(n7964),.dout(n7968),.clk(gclk));
	jand g07709(.dina(w_n7968_0[1]),.dinb(w_n7959_0[1]),.dout(n7969),.clk(gclk));
	jor g07710(.dina(n7969),.dinb(w_n7957_0[1]),.dout(n7970),.clk(gclk));
	jand g07711(.dina(w_n7970_0[1]),.dinb(w_asqrt57_18[0]),.dout(n7971),.clk(gclk));
	jxor g07712(.dina(w_n7548_0[0]),.dinb(w_n590_22[1]),.dout(n7972),.clk(gclk));
	jand g07713(.dina(n7972),.dinb(w_asqrt26_21[0]),.dout(n7973),.clk(gclk));
	jxor g07714(.dina(n7973),.dinb(w_n7558_0[0]),.dout(n7974),.clk(gclk));
	jnot g07715(.din(n7974),.dout(n7975),.clk(gclk));
	jor g07716(.dina(w_n7970_0[0]),.dinb(w_asqrt57_17[2]),.dout(n7976),.clk(gclk));
	jand g07717(.dina(w_n7976_0[1]),.dinb(w_n7975_0[1]),.dout(n7977),.clk(gclk));
	jor g07718(.dina(w_n7977_0[2]),.dinb(w_n7971_0[2]),.dout(n7978),.clk(gclk));
	jand g07719(.dina(n7978),.dinb(w_asqrt58_18[2]),.dout(n7979),.clk(gclk));
	jnot g07720(.din(w_n7563_0[0]),.dout(n7980),.clk(gclk));
	jand g07721(.dina(n7980),.dinb(w_n7561_0[0]),.dout(n7981),.clk(gclk));
	jand g07722(.dina(n7981),.dinb(w_asqrt26_20[2]),.dout(n7982),.clk(gclk));
	jxor g07723(.dina(n7982),.dinb(w_n7571_0[0]),.dout(n7983),.clk(gclk));
	jnot g07724(.din(n7983),.dout(n7984),.clk(gclk));
	jor g07725(.dina(w_n7971_0[1]),.dinb(w_asqrt58_18[1]),.dout(n7985),.clk(gclk));
	jor g07726(.dina(n7985),.dinb(w_n7977_0[1]),.dout(n7986),.clk(gclk));
	jand g07727(.dina(w_n7986_0[1]),.dinb(w_n7984_0[1]),.dout(n7987),.clk(gclk));
	jor g07728(.dina(w_n7987_0[1]),.dinb(w_n7979_0[1]),.dout(n7988),.clk(gclk));
	jand g07729(.dina(w_n7988_0[2]),.dinb(w_asqrt59_18[1]),.dout(n7989),.clk(gclk));
	jor g07730(.dina(w_n7988_0[1]),.dinb(w_asqrt59_18[0]),.dout(n7990),.clk(gclk));
	jnot g07731(.din(w_n7577_0[0]),.dout(n7991),.clk(gclk));
	jnot g07732(.din(w_n7578_0[0]),.dout(n7992),.clk(gclk));
	jand g07733(.dina(w_asqrt26_20[1]),.dinb(w_n7574_0[0]),.dout(n7993),.clk(gclk));
	jand g07734(.dina(w_n7993_0[1]),.dinb(n7992),.dout(n7994),.clk(gclk));
	jor g07735(.dina(n7994),.dinb(n7991),.dout(n7995),.clk(gclk));
	jnot g07736(.din(w_n7579_0[0]),.dout(n7996),.clk(gclk));
	jand g07737(.dina(w_n7993_0[0]),.dinb(n7996),.dout(n7997),.clk(gclk));
	jnot g07738(.din(n7997),.dout(n7998),.clk(gclk));
	jand g07739(.dina(n7998),.dinb(n7995),.dout(n7999),.clk(gclk));
	jand g07740(.dina(w_n7999_0[1]),.dinb(n7990),.dout(n8000),.clk(gclk));
	jor g07741(.dina(w_n8000_0[1]),.dinb(w_n7989_0[1]),.dout(n8001),.clk(gclk));
	jand g07742(.dina(n8001),.dinb(w_asqrt60_18[1]),.dout(n8002),.clk(gclk));
	jor g07743(.dina(w_n7989_0[0]),.dinb(w_asqrt60_18[0]),.dout(n8003),.clk(gclk));
	jor g07744(.dina(n8003),.dinb(w_n8000_0[0]),.dout(n8004),.clk(gclk));
	jnot g07745(.din(w_n7585_0[0]),.dout(n8005),.clk(gclk));
	jnot g07746(.din(w_n7587_0[0]),.dout(n8006),.clk(gclk));
	jand g07747(.dina(w_asqrt26_20[0]),.dinb(w_n7581_0[0]),.dout(n8007),.clk(gclk));
	jand g07748(.dina(w_n8007_0[1]),.dinb(n8006),.dout(n8008),.clk(gclk));
	jor g07749(.dina(n8008),.dinb(n8005),.dout(n8009),.clk(gclk));
	jnot g07750(.din(w_n7588_0[0]),.dout(n8010),.clk(gclk));
	jand g07751(.dina(w_n8007_0[0]),.dinb(n8010),.dout(n8011),.clk(gclk));
	jnot g07752(.din(n8011),.dout(n8012),.clk(gclk));
	jand g07753(.dina(n8012),.dinb(n8009),.dout(n8013),.clk(gclk));
	jand g07754(.dina(w_n8013_0[1]),.dinb(w_n8004_0[1]),.dout(n8014),.clk(gclk));
	jor g07755(.dina(n8014),.dinb(w_n8002_0[1]),.dout(n8015),.clk(gclk));
	jand g07756(.dina(w_n8015_0[1]),.dinb(w_asqrt61_18[2]),.dout(n8016),.clk(gclk));
	jxor g07757(.dina(w_n7589_0[0]),.dinb(w_n290_23[2]),.dout(n8017),.clk(gclk));
	jand g07758(.dina(n8017),.dinb(w_asqrt26_19[2]),.dout(n8018),.clk(gclk));
	jxor g07759(.dina(n8018),.dinb(w_n7599_0[0]),.dout(n8019),.clk(gclk));
	jnot g07760(.din(n8019),.dout(n8020),.clk(gclk));
	jor g07761(.dina(w_n8015_0[0]),.dinb(w_asqrt61_18[1]),.dout(n8021),.clk(gclk));
	jand g07762(.dina(w_n8021_0[1]),.dinb(w_n8020_0[1]),.dout(n8022),.clk(gclk));
	jor g07763(.dina(w_n8022_0[2]),.dinb(w_n8016_0[2]),.dout(n8023),.clk(gclk));
	jand g07764(.dina(n8023),.dinb(w_asqrt62_18[2]),.dout(n8024),.clk(gclk));
	jnot g07765(.din(w_n7604_0[0]),.dout(n8025),.clk(gclk));
	jand g07766(.dina(n8025),.dinb(w_n7602_0[0]),.dout(n8026),.clk(gclk));
	jand g07767(.dina(n8026),.dinb(w_asqrt26_19[1]),.dout(n8027),.clk(gclk));
	jxor g07768(.dina(n8027),.dinb(w_n7612_0[0]),.dout(n8028),.clk(gclk));
	jnot g07769(.din(n8028),.dout(n8029),.clk(gclk));
	jor g07770(.dina(w_n8016_0[1]),.dinb(w_asqrt62_18[1]),.dout(n8030),.clk(gclk));
	jor g07771(.dina(n8030),.dinb(w_n8022_0[1]),.dout(n8031),.clk(gclk));
	jand g07772(.dina(w_n8031_0[1]),.dinb(w_n8029_0[1]),.dout(n8032),.clk(gclk));
	jor g07773(.dina(w_n8032_0[1]),.dinb(w_n8024_0[1]),.dout(n8033),.clk(gclk));
	jxor g07774(.dina(w_n7614_0[0]),.dinb(w_n199_27[2]),.dout(n8034),.clk(gclk));
	jand g07775(.dina(n8034),.dinb(w_asqrt26_19[0]),.dout(n8035),.clk(gclk));
	jxor g07776(.dina(n8035),.dinb(w_n7619_0[0]),.dout(n8036),.clk(gclk));
	jnot g07777(.din(w_n7621_0[0]),.dout(n8037),.clk(gclk));
	jnot g07778(.din(w_n7625_0[0]),.dout(n8038),.clk(gclk));
	jand g07779(.dina(w_asqrt26_18[2]),.dinb(w_n8038_0[1]),.dout(n8039),.clk(gclk));
	jand g07780(.dina(w_n8039_0[1]),.dinb(w_n8037_0[2]),.dout(n8040),.clk(gclk));
	jor g07781(.dina(n8040),.dinb(w_n7632_0[0]),.dout(n8041),.clk(gclk));
	jor g07782(.dina(n8041),.dinb(w_n8036_0[1]),.dout(n8042),.clk(gclk));
	jnot g07783(.din(n8042),.dout(n8043),.clk(gclk));
	jand g07784(.dina(n8043),.dinb(w_n8033_1[2]),.dout(n8044),.clk(gclk));
	jor g07785(.dina(n8044),.dinb(w_asqrt63_10[0]),.dout(n8045),.clk(gclk));
	jnot g07786(.din(w_n8036_0[0]),.dout(n8046),.clk(gclk));
	jor g07787(.dina(w_n8046_0[2]),.dinb(w_n8033_1[1]),.dout(n8047),.clk(gclk));
	jor g07788(.dina(w_n8039_0[0]),.dinb(w_n8037_0[1]),.dout(n8048),.clk(gclk));
	jand g07789(.dina(w_n8038_0[0]),.dinb(w_n8037_0[0]),.dout(n8049),.clk(gclk));
	jor g07790(.dina(n8049),.dinb(w_n194_26[2]),.dout(n8050),.clk(gclk));
	jnot g07791(.din(n8050),.dout(n8051),.clk(gclk));
	jand g07792(.dina(n8051),.dinb(n8048),.dout(n8052),.clk(gclk));
	jnot g07793(.din(w_asqrt26_18[1]),.dout(n8053),.clk(gclk));
	jnot g07794(.din(w_n8052_0[1]),.dout(n8056),.clk(gclk));
	jand g07795(.dina(n8056),.dinb(w_n8047_0[1]),.dout(n8057),.clk(gclk));
	jand g07796(.dina(n8057),.dinb(w_n8045_0[1]),.dout(n8058),.clk(gclk));
	jxor g07797(.dina(w_n7745_0[0]),.dinb(w_n3912_21[0]),.dout(n8059),.clk(gclk));
	jor g07798(.dina(n8059),.dinb(w_n8058_27[1]),.dout(n8060),.clk(gclk));
	jxor g07799(.dina(n8060),.dinb(w_n7645_0[0]),.dout(n8061),.clk(gclk));
	jor g07800(.dina(w_n8058_27[0]),.dinb(w_n7647_1[0]),.dout(n8062),.clk(gclk));
	jnot g07801(.din(w_a48_0[1]),.dout(n8063),.clk(gclk));
	jnot g07802(.din(a[49]),.dout(n8064),.clk(gclk));
	jand g07803(.dina(w_n7647_0[2]),.dinb(w_n8064_0[2]),.dout(n8065),.clk(gclk));
	jand g07804(.dina(n8065),.dinb(w_n8063_1[1]),.dout(n8066),.clk(gclk));
	jnot g07805(.din(n8066),.dout(n8067),.clk(gclk));
	jand g07806(.dina(n8067),.dinb(n8062),.dout(n8068),.clk(gclk));
	jor g07807(.dina(w_n8068_0[2]),.dinb(w_n8053_16[2]),.dout(n8069),.clk(gclk));
	jor g07808(.dina(w_n8058_26[2]),.dinb(w_a50_0[0]),.dout(n8070),.clk(gclk));
	jxor g07809(.dina(w_n8070_0[1]),.dinb(w_n7648_0[0]),.dout(n8071),.clk(gclk));
	jand g07810(.dina(w_n8068_0[1]),.dinb(w_n8053_16[1]),.dout(n8072),.clk(gclk));
	jor g07811(.dina(n8072),.dinb(w_n8071_0[1]),.dout(n8073),.clk(gclk));
	jand g07812(.dina(w_n8073_0[1]),.dinb(w_n8069_0[1]),.dout(n8074),.clk(gclk));
	jor g07813(.dina(n8074),.dinb(w_n7265_20[2]),.dout(n8075),.clk(gclk));
	jand g07814(.dina(w_n8069_0[0]),.dinb(w_n7265_20[1]),.dout(n8076),.clk(gclk));
	jand g07815(.dina(n8076),.dinb(w_n8073_0[0]),.dout(n8077),.clk(gclk));
	jor g07816(.dina(w_n8070_0[0]),.dinb(w_a51_0[0]),.dout(n8078),.clk(gclk));
	jnot g07817(.din(w_n8045_0[0]),.dout(n8079),.clk(gclk));
	jnot g07818(.din(w_n8047_0[0]),.dout(n8080),.clk(gclk));
	jor g07819(.dina(w_n8052_0[0]),.dinb(w_n8053_16[0]),.dout(n8081),.clk(gclk));
	jor g07820(.dina(n8081),.dinb(w_n8080_0[1]),.dout(n8082),.clk(gclk));
	jor g07821(.dina(n8082),.dinb(n8079),.dout(n8083),.clk(gclk));
	jand g07822(.dina(n8083),.dinb(n8078),.dout(n8084),.clk(gclk));
	jxor g07823(.dina(n8084),.dinb(w_n7271_0[1]),.dout(n8085),.clk(gclk));
	jor g07824(.dina(w_n8085_0[1]),.dinb(w_n8077_0[1]),.dout(n8086),.clk(gclk));
	jand g07825(.dina(n8086),.dinb(w_n8075_0[1]),.dout(n8087),.clk(gclk));
	jor g07826(.dina(w_n8087_0[2]),.dinb(w_n7260_17[0]),.dout(n8088),.clk(gclk));
	jand g07827(.dina(w_n8087_0[1]),.dinb(w_n7260_16[2]),.dout(n8089),.clk(gclk));
	jxor g07828(.dina(w_n7651_0[0]),.dinb(w_n7265_20[0]),.dout(n8090),.clk(gclk));
	jor g07829(.dina(n8090),.dinb(w_n8058_26[1]),.dout(n8091),.clk(gclk));
	jxor g07830(.dina(n8091),.dinb(w_n7654_0[0]),.dout(n8092),.clk(gclk));
	jor g07831(.dina(w_n8092_0[1]),.dinb(n8089),.dout(n8093),.clk(gclk));
	jand g07832(.dina(w_n8093_0[1]),.dinb(w_n8088_0[1]),.dout(n8094),.clk(gclk));
	jor g07833(.dina(n8094),.dinb(w_n6505_20[1]),.dout(n8095),.clk(gclk));
	jnot g07834(.din(w_n7660_0[0]),.dout(n8096),.clk(gclk));
	jor g07835(.dina(n8096),.dinb(w_n7658_0[0]),.dout(n8097),.clk(gclk));
	jor g07836(.dina(n8097),.dinb(w_n8058_26[0]),.dout(n8098),.clk(gclk));
	jxor g07837(.dina(n8098),.dinb(w_n7669_0[0]),.dout(n8099),.clk(gclk));
	jand g07838(.dina(w_n8088_0[0]),.dinb(w_n6505_20[0]),.dout(n8100),.clk(gclk));
	jand g07839(.dina(n8100),.dinb(w_n8093_0[0]),.dout(n8101),.clk(gclk));
	jor g07840(.dina(w_n8101_0[1]),.dinb(w_n8099_0[1]),.dout(n8102),.clk(gclk));
	jand g07841(.dina(w_n8102_0[1]),.dinb(w_n8095_0[1]),.dout(n8103),.clk(gclk));
	jor g07842(.dina(w_n8103_0[2]),.dinb(w_n6500_17[0]),.dout(n8104),.clk(gclk));
	jand g07843(.dina(w_n8103_0[1]),.dinb(w_n6500_16[2]),.dout(n8105),.clk(gclk));
	jxor g07844(.dina(w_n7671_0[0]),.dinb(w_n6505_19[2]),.dout(n8106),.clk(gclk));
	jor g07845(.dina(n8106),.dinb(w_n8058_25[2]),.dout(n8107),.clk(gclk));
	jxor g07846(.dina(n8107),.dinb(w_n7676_0[0]),.dout(n8108),.clk(gclk));
	jnot g07847(.din(w_n8108_0[1]),.dout(n8109),.clk(gclk));
	jor g07848(.dina(n8109),.dinb(n8105),.dout(n8110),.clk(gclk));
	jand g07849(.dina(w_n8110_0[1]),.dinb(w_n8104_0[1]),.dout(n8111),.clk(gclk));
	jor g07850(.dina(n8111),.dinb(w_n5793_20[2]),.dout(n8112),.clk(gclk));
	jand g07851(.dina(w_n8104_0[0]),.dinb(w_n5793_20[1]),.dout(n8113),.clk(gclk));
	jand g07852(.dina(n8113),.dinb(w_n8110_0[0]),.dout(n8114),.clk(gclk));
	jnot g07853(.din(w_n7680_0[0]),.dout(n8115),.clk(gclk));
	jnot g07854(.din(w_n8058_25[1]),.dout(asqrt_fa_26),.clk(gclk));
	jand g07855(.dina(w_asqrt25_20),.dinb(n8115),.dout(n8117),.clk(gclk));
	jand g07856(.dina(w_n8117_0[1]),.dinb(w_n7687_0[0]),.dout(n8118),.clk(gclk));
	jor g07857(.dina(n8118),.dinb(w_n7685_0[0]),.dout(n8119),.clk(gclk));
	jand g07858(.dina(w_n8117_0[0]),.dinb(w_n7688_0[0]),.dout(n8120),.clk(gclk));
	jnot g07859(.din(n8120),.dout(n8121),.clk(gclk));
	jand g07860(.dina(n8121),.dinb(n8119),.dout(n8122),.clk(gclk));
	jnot g07861(.din(n8122),.dout(n8123),.clk(gclk));
	jor g07862(.dina(w_n8123_0[1]),.dinb(w_n8114_0[1]),.dout(n8124),.clk(gclk));
	jand g07863(.dina(n8124),.dinb(w_n8112_0[1]),.dout(n8125),.clk(gclk));
	jor g07864(.dina(w_n8125_0[2]),.dinb(w_n5788_17[1]),.dout(n8126),.clk(gclk));
	jand g07865(.dina(w_n8125_0[1]),.dinb(w_n5788_17[0]),.dout(n8127),.clk(gclk));
	jnot g07866(.din(w_n7695_0[0]),.dout(n8128),.clk(gclk));
	jxor g07867(.dina(w_n7689_0[0]),.dinb(w_n5793_20[0]),.dout(n8129),.clk(gclk));
	jor g07868(.dina(n8129),.dinb(w_n8058_25[0]),.dout(n8130),.clk(gclk));
	jxor g07869(.dina(n8130),.dinb(n8128),.dout(n8131),.clk(gclk));
	jnot g07870(.din(w_n8131_0[1]),.dout(n8132),.clk(gclk));
	jor g07871(.dina(n8132),.dinb(n8127),.dout(n8133),.clk(gclk));
	jand g07872(.dina(w_n8133_0[1]),.dinb(w_n8126_0[1]),.dout(n8134),.clk(gclk));
	jor g07873(.dina(n8134),.dinb(w_n5121_20[1]),.dout(n8135),.clk(gclk));
	jnot g07874(.din(w_n7700_0[0]),.dout(n8136),.clk(gclk));
	jor g07875(.dina(n8136),.dinb(w_n7698_0[0]),.dout(n8137),.clk(gclk));
	jor g07876(.dina(n8137),.dinb(w_n8058_24[2]),.dout(n8138),.clk(gclk));
	jxor g07877(.dina(n8138),.dinb(w_n7709_0[0]),.dout(n8139),.clk(gclk));
	jand g07878(.dina(w_n8126_0[0]),.dinb(w_n5121_20[0]),.dout(n8140),.clk(gclk));
	jand g07879(.dina(n8140),.dinb(w_n8133_0[0]),.dout(n8141),.clk(gclk));
	jor g07880(.dina(w_n8141_0[1]),.dinb(w_n8139_0[1]),.dout(n8142),.clk(gclk));
	jand g07881(.dina(w_n8142_0[1]),.dinb(w_n8135_0[1]),.dout(n8143),.clk(gclk));
	jor g07882(.dina(w_n8143_0[2]),.dinb(w_n5116_17[1]),.dout(n8144),.clk(gclk));
	jand g07883(.dina(w_n8143_0[1]),.dinb(w_n5116_17[0]),.dout(n8145),.clk(gclk));
	jnot g07884(.din(w_n7716_0[0]),.dout(n8146),.clk(gclk));
	jxor g07885(.dina(w_n7711_0[0]),.dinb(w_n5121_19[2]),.dout(n8147),.clk(gclk));
	jor g07886(.dina(n8147),.dinb(w_n8058_24[1]),.dout(n8148),.clk(gclk));
	jxor g07887(.dina(n8148),.dinb(n8146),.dout(n8149),.clk(gclk));
	jnot g07888(.din(n8149),.dout(n8150),.clk(gclk));
	jor g07889(.dina(w_n8150_0[1]),.dinb(n8145),.dout(n8151),.clk(gclk));
	jand g07890(.dina(w_n8151_0[1]),.dinb(w_n8144_0[1]),.dout(n8152),.clk(gclk));
	jor g07891(.dina(n8152),.dinb(w_n4499_21[0]),.dout(n8153),.clk(gclk));
	jand g07892(.dina(w_n8144_0[0]),.dinb(w_n4499_20[2]),.dout(n8154),.clk(gclk));
	jand g07893(.dina(n8154),.dinb(w_n8151_0[0]),.dout(n8155),.clk(gclk));
	jnot g07894(.din(w_n7719_0[0]),.dout(n8156),.clk(gclk));
	jand g07895(.dina(w_asqrt25_19[2]),.dinb(n8156),.dout(n8157),.clk(gclk));
	jand g07896(.dina(w_n8157_0[1]),.dinb(w_n7726_0[0]),.dout(n8158),.clk(gclk));
	jor g07897(.dina(n8158),.dinb(w_n7724_0[0]),.dout(n8159),.clk(gclk));
	jand g07898(.dina(w_n8157_0[0]),.dinb(w_n7727_0[0]),.dout(n8160),.clk(gclk));
	jnot g07899(.din(n8160),.dout(n8161),.clk(gclk));
	jand g07900(.dina(n8161),.dinb(n8159),.dout(n8162),.clk(gclk));
	jnot g07901(.din(n8162),.dout(n8163),.clk(gclk));
	jor g07902(.dina(w_n8163_0[1]),.dinb(w_n8155_0[1]),.dout(n8164),.clk(gclk));
	jand g07903(.dina(n8164),.dinb(w_n8153_0[1]),.dout(n8165),.clk(gclk));
	jor g07904(.dina(w_n8165_0[1]),.dinb(w_n4494_18[0]),.dout(n8166),.clk(gclk));
	jxor g07905(.dina(w_n7728_0[0]),.dinb(w_n4499_20[1]),.dout(n8167),.clk(gclk));
	jor g07906(.dina(n8167),.dinb(w_n8058_24[0]),.dout(n8168),.clk(gclk));
	jxor g07907(.dina(n8168),.dinb(w_n7733_0[0]),.dout(n8169),.clk(gclk));
	jand g07908(.dina(w_n8165_0[0]),.dinb(w_n4494_17[2]),.dout(n8170),.clk(gclk));
	jor g07909(.dina(w_n8170_0[1]),.dinb(w_n8169_0[1]),.dout(n8171),.clk(gclk));
	jand g07910(.dina(w_n8171_0[2]),.dinb(w_n8166_0[2]),.dout(n8172),.clk(gclk));
	jor g07911(.dina(n8172),.dinb(w_n3912_20[2]),.dout(n8173),.clk(gclk));
	jand g07912(.dina(w_n8166_0[1]),.dinb(w_n3912_20[1]),.dout(n8174),.clk(gclk));
	jand g07913(.dina(n8174),.dinb(w_n8171_0[1]),.dout(n8175),.clk(gclk));
	jnot g07914(.din(w_n7736_0[0]),.dout(n8176),.clk(gclk));
	jand g07915(.dina(w_asqrt25_19[1]),.dinb(n8176),.dout(n8177),.clk(gclk));
	jand g07916(.dina(w_n8177_0[1]),.dinb(w_n7743_0[0]),.dout(n8178),.clk(gclk));
	jor g07917(.dina(n8178),.dinb(w_n7741_0[0]),.dout(n8179),.clk(gclk));
	jand g07918(.dina(w_n8177_0[0]),.dinb(w_n7744_0[0]),.dout(n8180),.clk(gclk));
	jnot g07919(.din(n8180),.dout(n8181),.clk(gclk));
	jand g07920(.dina(n8181),.dinb(n8179),.dout(n8182),.clk(gclk));
	jnot g07921(.din(n8182),.dout(n8183),.clk(gclk));
	jor g07922(.dina(w_n8183_0[1]),.dinb(w_n8175_0[1]),.dout(n8184),.clk(gclk));
	jand g07923(.dina(n8184),.dinb(w_n8173_0[1]),.dout(n8185),.clk(gclk));
	jor g07924(.dina(w_n8185_0[2]),.dinb(w_n3907_18[1]),.dout(n8186),.clk(gclk));
	jand g07925(.dina(w_n8185_0[1]),.dinb(w_n3907_18[0]),.dout(n8187),.clk(gclk));
	jor g07926(.dina(n8187),.dinb(w_n8061_0[1]),.dout(n8188),.clk(gclk));
	jand g07927(.dina(w_n8188_0[1]),.dinb(w_n8186_0[1]),.dout(n8189),.clk(gclk));
	jor g07928(.dina(n8189),.dinb(w_n3376_22[0]),.dout(n8190),.clk(gclk));
	jnot g07929(.din(w_n7752_0[0]),.dout(n8191),.clk(gclk));
	jor g07930(.dina(n8191),.dinb(w_n7750_0[0]),.dout(n8192),.clk(gclk));
	jor g07931(.dina(n8192),.dinb(w_n8058_23[2]),.dout(n8193),.clk(gclk));
	jxor g07932(.dina(n8193),.dinb(w_n7761_0[0]),.dout(n8194),.clk(gclk));
	jand g07933(.dina(w_n8186_0[0]),.dinb(w_n3376_21[2]),.dout(n8195),.clk(gclk));
	jand g07934(.dina(n8195),.dinb(w_n8188_0[0]),.dout(n8196),.clk(gclk));
	jor g07935(.dina(w_n8196_0[1]),.dinb(w_n8194_0[1]),.dout(n8197),.clk(gclk));
	jand g07936(.dina(w_n8197_0[1]),.dinb(w_n8190_0[1]),.dout(n8198),.clk(gclk));
	jor g07937(.dina(w_n8198_0[1]),.dinb(w_n3371_18[2]),.dout(n8199),.clk(gclk));
	jxor g07938(.dina(w_n7763_0[0]),.dinb(w_n3376_21[1]),.dout(n8200),.clk(gclk));
	jor g07939(.dina(n8200),.dinb(w_n8058_23[1]),.dout(n8201),.clk(gclk));
	jxor g07940(.dina(n8201),.dinb(w_n7774_0[0]),.dout(n8202),.clk(gclk));
	jand g07941(.dina(w_n8198_0[0]),.dinb(w_n3371_18[1]),.dout(n8203),.clk(gclk));
	jor g07942(.dina(w_n8203_0[1]),.dinb(w_n8202_0[1]),.dout(n8204),.clk(gclk));
	jand g07943(.dina(w_n8204_0[2]),.dinb(w_n8199_0[2]),.dout(n8205),.clk(gclk));
	jor g07944(.dina(n8205),.dinb(w_n2875_21[2]),.dout(n8206),.clk(gclk));
	jnot g07945(.din(w_n7779_0[0]),.dout(n8207),.clk(gclk));
	jor g07946(.dina(n8207),.dinb(w_n7777_0[0]),.dout(n8208),.clk(gclk));
	jor g07947(.dina(n8208),.dinb(w_n8058_23[0]),.dout(n8209),.clk(gclk));
	jxor g07948(.dina(n8209),.dinb(w_n7788_0[0]),.dout(n8210),.clk(gclk));
	jand g07949(.dina(w_n8199_0[1]),.dinb(w_n2875_21[1]),.dout(n8211),.clk(gclk));
	jand g07950(.dina(n8211),.dinb(w_n8204_0[1]),.dout(n8212),.clk(gclk));
	jor g07951(.dina(w_n8212_0[1]),.dinb(w_n8210_0[1]),.dout(n8213),.clk(gclk));
	jand g07952(.dina(w_n8213_0[1]),.dinb(w_n8206_0[1]),.dout(n8214),.clk(gclk));
	jor g07953(.dina(w_n8214_0[2]),.dinb(w_n2870_19[0]),.dout(n8215),.clk(gclk));
	jand g07954(.dina(w_n8214_0[1]),.dinb(w_n2870_18[2]),.dout(n8216),.clk(gclk));
	jnot g07955(.din(w_n7791_0[0]),.dout(n8217),.clk(gclk));
	jand g07956(.dina(w_asqrt25_19[0]),.dinb(n8217),.dout(n8218),.clk(gclk));
	jand g07957(.dina(w_n8218_0[1]),.dinb(w_n7796_0[0]),.dout(n8219),.clk(gclk));
	jor g07958(.dina(n8219),.dinb(w_n7795_0[0]),.dout(n8220),.clk(gclk));
	jand g07959(.dina(w_n8218_0[0]),.dinb(w_n7797_0[0]),.dout(n8221),.clk(gclk));
	jnot g07960(.din(n8221),.dout(n8222),.clk(gclk));
	jand g07961(.dina(n8222),.dinb(n8220),.dout(n8223),.clk(gclk));
	jnot g07962(.din(n8223),.dout(n8224),.clk(gclk));
	jor g07963(.dina(w_n8224_0[1]),.dinb(n8216),.dout(n8225),.clk(gclk));
	jand g07964(.dina(w_n8225_0[1]),.dinb(w_n8215_0[1]),.dout(n8226),.clk(gclk));
	jor g07965(.dina(n8226),.dinb(w_n2425_22[1]),.dout(n8227),.clk(gclk));
	jand g07966(.dina(w_n8215_0[0]),.dinb(w_n2425_22[0]),.dout(n8228),.clk(gclk));
	jand g07967(.dina(n8228),.dinb(w_n8225_0[0]),.dout(n8229),.clk(gclk));
	jnot g07968(.din(w_n7799_0[0]),.dout(n8230),.clk(gclk));
	jand g07969(.dina(w_asqrt25_18[2]),.dinb(n8230),.dout(n8231),.clk(gclk));
	jand g07970(.dina(w_n8231_0[1]),.dinb(w_n7806_0[0]),.dout(n8232),.clk(gclk));
	jor g07971(.dina(n8232),.dinb(w_n7804_0[0]),.dout(n8233),.clk(gclk));
	jand g07972(.dina(w_n8231_0[0]),.dinb(w_n7807_0[0]),.dout(n8234),.clk(gclk));
	jnot g07973(.din(n8234),.dout(n8235),.clk(gclk));
	jand g07974(.dina(n8235),.dinb(n8233),.dout(n8236),.clk(gclk));
	jnot g07975(.din(n8236),.dout(n8237),.clk(gclk));
	jor g07976(.dina(w_n8237_0[1]),.dinb(w_n8229_0[1]),.dout(n8238),.clk(gclk));
	jand g07977(.dina(n8238),.dinb(w_n8227_0[1]),.dout(n8239),.clk(gclk));
	jor g07978(.dina(w_n8239_0[1]),.dinb(w_n2420_19[2]),.dout(n8240),.clk(gclk));
	jxor g07979(.dina(w_n7808_0[0]),.dinb(w_n2425_21[2]),.dout(n8241),.clk(gclk));
	jor g07980(.dina(n8241),.dinb(w_n8058_22[2]),.dout(n8242),.clk(gclk));
	jxor g07981(.dina(n8242),.dinb(w_n7819_0[0]),.dout(n8243),.clk(gclk));
	jand g07982(.dina(w_n8239_0[0]),.dinb(w_n2420_19[1]),.dout(n8244),.clk(gclk));
	jor g07983(.dina(w_n8244_0[1]),.dinb(w_n8243_0[1]),.dout(n8245),.clk(gclk));
	jand g07984(.dina(w_n8245_0[2]),.dinb(w_n8240_0[2]),.dout(n8246),.clk(gclk));
	jor g07985(.dina(n8246),.dinb(w_n2010_22[0]),.dout(n8247),.clk(gclk));
	jnot g07986(.din(w_n7824_0[0]),.dout(n8248),.clk(gclk));
	jor g07987(.dina(n8248),.dinb(w_n7822_0[0]),.dout(n8249),.clk(gclk));
	jor g07988(.dina(n8249),.dinb(w_n8058_22[1]),.dout(n8250),.clk(gclk));
	jxor g07989(.dina(n8250),.dinb(w_n7833_0[0]),.dout(n8251),.clk(gclk));
	jand g07990(.dina(w_n8240_0[1]),.dinb(w_n2010_21[2]),.dout(n8252),.clk(gclk));
	jand g07991(.dina(n8252),.dinb(w_n8245_0[1]),.dout(n8253),.clk(gclk));
	jor g07992(.dina(w_n8253_0[1]),.dinb(w_n8251_0[1]),.dout(n8254),.clk(gclk));
	jand g07993(.dina(w_n8254_0[1]),.dinb(w_n8247_0[1]),.dout(n8255),.clk(gclk));
	jor g07994(.dina(w_n8255_0[2]),.dinb(w_n2005_20[0]),.dout(n8256),.clk(gclk));
	jand g07995(.dina(w_n8255_0[1]),.dinb(w_n2005_19[2]),.dout(n8257),.clk(gclk));
	jnot g07996(.din(w_n7836_0[0]),.dout(n8258),.clk(gclk));
	jand g07997(.dina(w_asqrt25_18[1]),.dinb(n8258),.dout(n8259),.clk(gclk));
	jand g07998(.dina(w_n8259_0[1]),.dinb(w_n7841_0[0]),.dout(n8260),.clk(gclk));
	jor g07999(.dina(n8260),.dinb(w_n7840_0[0]),.dout(n8261),.clk(gclk));
	jand g08000(.dina(w_n8259_0[0]),.dinb(w_n7842_0[0]),.dout(n8262),.clk(gclk));
	jnot g08001(.din(n8262),.dout(n8263),.clk(gclk));
	jand g08002(.dina(n8263),.dinb(n8261),.dout(n8264),.clk(gclk));
	jnot g08003(.din(n8264),.dout(n8265),.clk(gclk));
	jor g08004(.dina(w_n8265_0[1]),.dinb(n8257),.dout(n8266),.clk(gclk));
	jand g08005(.dina(w_n8266_0[1]),.dinb(w_n8256_0[1]),.dout(n8267),.clk(gclk));
	jor g08006(.dina(n8267),.dinb(w_n1646_23[0]),.dout(n8268),.clk(gclk));
	jand g08007(.dina(w_n8256_0[0]),.dinb(w_n1646_22[2]),.dout(n8269),.clk(gclk));
	jand g08008(.dina(n8269),.dinb(w_n8266_0[0]),.dout(n8270),.clk(gclk));
	jnot g08009(.din(w_n7844_0[0]),.dout(n8271),.clk(gclk));
	jand g08010(.dina(w_asqrt25_18[0]),.dinb(n8271),.dout(n8272),.clk(gclk));
	jand g08011(.dina(w_n8272_0[1]),.dinb(w_n7851_0[0]),.dout(n8273),.clk(gclk));
	jor g08012(.dina(n8273),.dinb(w_n7849_0[0]),.dout(n8274),.clk(gclk));
	jand g08013(.dina(w_n8272_0[0]),.dinb(w_n7852_0[0]),.dout(n8275),.clk(gclk));
	jnot g08014(.din(n8275),.dout(n8276),.clk(gclk));
	jand g08015(.dina(n8276),.dinb(n8274),.dout(n8277),.clk(gclk));
	jnot g08016(.din(n8277),.dout(n8278),.clk(gclk));
	jor g08017(.dina(w_n8278_0[1]),.dinb(w_n8270_0[1]),.dout(n8279),.clk(gclk));
	jand g08018(.dina(n8279),.dinb(w_n8268_0[1]),.dout(n8280),.clk(gclk));
	jor g08019(.dina(w_n8280_0[1]),.dinb(w_n1641_20[1]),.dout(n8281),.clk(gclk));
	jxor g08020(.dina(w_n7853_0[0]),.dinb(w_n1646_22[1]),.dout(n8282),.clk(gclk));
	jor g08021(.dina(n8282),.dinb(w_n8058_22[0]),.dout(n8283),.clk(gclk));
	jxor g08022(.dina(n8283),.dinb(w_n7864_0[0]),.dout(n8284),.clk(gclk));
	jand g08023(.dina(w_n8280_0[0]),.dinb(w_n1641_20[0]),.dout(n8285),.clk(gclk));
	jor g08024(.dina(w_n8285_0[1]),.dinb(w_n8284_0[1]),.dout(n8286),.clk(gclk));
	jand g08025(.dina(w_n8286_0[2]),.dinb(w_n8281_0[2]),.dout(n8287),.clk(gclk));
	jor g08026(.dina(n8287),.dinb(w_n1317_22[2]),.dout(n8288),.clk(gclk));
	jnot g08027(.din(w_n7869_0[0]),.dout(n8289),.clk(gclk));
	jor g08028(.dina(n8289),.dinb(w_n7867_0[0]),.dout(n8290),.clk(gclk));
	jor g08029(.dina(n8290),.dinb(w_n8058_21[2]),.dout(n8291),.clk(gclk));
	jxor g08030(.dina(n8291),.dinb(w_n7878_0[0]),.dout(n8292),.clk(gclk));
	jand g08031(.dina(w_n8281_0[1]),.dinb(w_n1317_22[1]),.dout(n8293),.clk(gclk));
	jand g08032(.dina(n8293),.dinb(w_n8286_0[1]),.dout(n8294),.clk(gclk));
	jor g08033(.dina(w_n8294_0[1]),.dinb(w_n8292_0[1]),.dout(n8295),.clk(gclk));
	jand g08034(.dina(w_n8295_0[1]),.dinb(w_n8288_0[1]),.dout(n8296),.clk(gclk));
	jor g08035(.dina(w_n8296_0[2]),.dinb(w_n1312_20[2]),.dout(n8297),.clk(gclk));
	jand g08036(.dina(w_n8296_0[1]),.dinb(w_n1312_20[1]),.dout(n8298),.clk(gclk));
	jnot g08037(.din(w_n7881_0[0]),.dout(n8299),.clk(gclk));
	jand g08038(.dina(w_asqrt25_17[2]),.dinb(n8299),.dout(n8300),.clk(gclk));
	jand g08039(.dina(w_n8300_0[1]),.dinb(w_n7886_0[0]),.dout(n8301),.clk(gclk));
	jor g08040(.dina(n8301),.dinb(w_n7885_0[0]),.dout(n8302),.clk(gclk));
	jand g08041(.dina(w_n8300_0[0]),.dinb(w_n7887_0[0]),.dout(n8303),.clk(gclk));
	jnot g08042(.din(n8303),.dout(n8304),.clk(gclk));
	jand g08043(.dina(n8304),.dinb(n8302),.dout(n8305),.clk(gclk));
	jnot g08044(.din(n8305),.dout(n8306),.clk(gclk));
	jor g08045(.dina(w_n8306_0[1]),.dinb(n8298),.dout(n8307),.clk(gclk));
	jand g08046(.dina(w_n8307_0[1]),.dinb(w_n8297_0[1]),.dout(n8308),.clk(gclk));
	jor g08047(.dina(n8308),.dinb(w_n1039_23[1]),.dout(n8309),.clk(gclk));
	jand g08048(.dina(w_n8297_0[0]),.dinb(w_n1039_23[0]),.dout(n8310),.clk(gclk));
	jand g08049(.dina(n8310),.dinb(w_n8307_0[0]),.dout(n8311),.clk(gclk));
	jnot g08050(.din(w_n7889_0[0]),.dout(n8312),.clk(gclk));
	jand g08051(.dina(w_asqrt25_17[1]),.dinb(n8312),.dout(n8313),.clk(gclk));
	jand g08052(.dina(w_n8313_0[1]),.dinb(w_n7896_0[0]),.dout(n8314),.clk(gclk));
	jor g08053(.dina(n8314),.dinb(w_n7894_0[0]),.dout(n8315),.clk(gclk));
	jand g08054(.dina(w_n8313_0[0]),.dinb(w_n7897_0[0]),.dout(n8316),.clk(gclk));
	jnot g08055(.din(n8316),.dout(n8317),.clk(gclk));
	jand g08056(.dina(n8317),.dinb(n8315),.dout(n8318),.clk(gclk));
	jnot g08057(.din(n8318),.dout(n8319),.clk(gclk));
	jor g08058(.dina(w_n8319_0[1]),.dinb(w_n8311_0[1]),.dout(n8320),.clk(gclk));
	jand g08059(.dina(n8320),.dinb(w_n8309_0[1]),.dout(n8321),.clk(gclk));
	jor g08060(.dina(w_n8321_0[1]),.dinb(w_n1034_21[1]),.dout(n8322),.clk(gclk));
	jxor g08061(.dina(w_n7898_0[0]),.dinb(w_n1039_22[2]),.dout(n8323),.clk(gclk));
	jor g08062(.dina(n8323),.dinb(w_n8058_21[1]),.dout(n8324),.clk(gclk));
	jxor g08063(.dina(n8324),.dinb(w_n7909_0[0]),.dout(n8325),.clk(gclk));
	jand g08064(.dina(w_n8321_0[0]),.dinb(w_n1034_21[0]),.dout(n8326),.clk(gclk));
	jor g08065(.dina(w_n8326_0[1]),.dinb(w_n8325_0[1]),.dout(n8327),.clk(gclk));
	jand g08066(.dina(w_n8327_0[2]),.dinb(w_n8322_0[2]),.dout(n8328),.clk(gclk));
	jor g08067(.dina(n8328),.dinb(w_n796_23[0]),.dout(n8329),.clk(gclk));
	jnot g08068(.din(w_n7914_0[0]),.dout(n8330),.clk(gclk));
	jor g08069(.dina(n8330),.dinb(w_n7912_0[0]),.dout(n8331),.clk(gclk));
	jor g08070(.dina(n8331),.dinb(w_n8058_21[0]),.dout(n8332),.clk(gclk));
	jxor g08071(.dina(n8332),.dinb(w_n7923_0[0]),.dout(n8333),.clk(gclk));
	jand g08072(.dina(w_n8322_0[1]),.dinb(w_n796_22[2]),.dout(n8334),.clk(gclk));
	jand g08073(.dina(n8334),.dinb(w_n8327_0[1]),.dout(n8335),.clk(gclk));
	jor g08074(.dina(w_n8335_0[1]),.dinb(w_n8333_0[1]),.dout(n8336),.clk(gclk));
	jand g08075(.dina(w_n8336_0[1]),.dinb(w_n8329_0[1]),.dout(n8337),.clk(gclk));
	jor g08076(.dina(w_n8337_0[2]),.dinb(w_n791_21[2]),.dout(n8338),.clk(gclk));
	jand g08077(.dina(w_n8337_0[1]),.dinb(w_n791_21[1]),.dout(n8339),.clk(gclk));
	jnot g08078(.din(w_n7926_0[0]),.dout(n8340),.clk(gclk));
	jand g08079(.dina(w_asqrt25_17[0]),.dinb(n8340),.dout(n8341),.clk(gclk));
	jand g08080(.dina(w_n8341_0[1]),.dinb(w_n7931_0[0]),.dout(n8342),.clk(gclk));
	jor g08081(.dina(n8342),.dinb(w_n7930_0[0]),.dout(n8343),.clk(gclk));
	jand g08082(.dina(w_n8341_0[0]),.dinb(w_n7932_0[0]),.dout(n8344),.clk(gclk));
	jnot g08083(.din(n8344),.dout(n8345),.clk(gclk));
	jand g08084(.dina(n8345),.dinb(n8343),.dout(n8346),.clk(gclk));
	jnot g08085(.din(n8346),.dout(n8347),.clk(gclk));
	jor g08086(.dina(w_n8347_0[1]),.dinb(n8339),.dout(n8348),.clk(gclk));
	jand g08087(.dina(w_n8348_0[1]),.dinb(w_n8338_0[1]),.dout(n8349),.clk(gclk));
	jor g08088(.dina(n8349),.dinb(w_n595_23[2]),.dout(n8350),.clk(gclk));
	jand g08089(.dina(w_n8338_0[0]),.dinb(w_n595_23[1]),.dout(n8351),.clk(gclk));
	jand g08090(.dina(n8351),.dinb(w_n8348_0[0]),.dout(n8352),.clk(gclk));
	jnot g08091(.din(w_n7934_0[0]),.dout(n8353),.clk(gclk));
	jand g08092(.dina(w_asqrt25_16[2]),.dinb(n8353),.dout(n8354),.clk(gclk));
	jand g08093(.dina(w_n8354_0[1]),.dinb(w_n7941_0[0]),.dout(n8355),.clk(gclk));
	jor g08094(.dina(n8355),.dinb(w_n7939_0[0]),.dout(n8356),.clk(gclk));
	jand g08095(.dina(w_n8354_0[0]),.dinb(w_n7942_0[0]),.dout(n8357),.clk(gclk));
	jnot g08096(.din(n8357),.dout(n8358),.clk(gclk));
	jand g08097(.dina(n8358),.dinb(n8356),.dout(n8359),.clk(gclk));
	jnot g08098(.din(n8359),.dout(n8360),.clk(gclk));
	jor g08099(.dina(w_n8360_0[1]),.dinb(w_n8352_0[1]),.dout(n8361),.clk(gclk));
	jand g08100(.dina(n8361),.dinb(w_n8350_0[1]),.dout(n8362),.clk(gclk));
	jor g08101(.dina(w_n8362_0[1]),.dinb(w_n590_22[0]),.dout(n8363),.clk(gclk));
	jxor g08102(.dina(w_n7943_0[0]),.dinb(w_n595_23[0]),.dout(n8364),.clk(gclk));
	jor g08103(.dina(n8364),.dinb(w_n8058_20[2]),.dout(n8365),.clk(gclk));
	jxor g08104(.dina(n8365),.dinb(w_n7954_0[0]),.dout(n8366),.clk(gclk));
	jand g08105(.dina(w_n8362_0[0]),.dinb(w_n590_21[2]),.dout(n8367),.clk(gclk));
	jor g08106(.dina(w_n8367_0[1]),.dinb(w_n8366_0[1]),.dout(n8368),.clk(gclk));
	jand g08107(.dina(w_n8368_0[2]),.dinb(w_n8363_0[2]),.dout(n8369),.clk(gclk));
	jor g08108(.dina(n8369),.dinb(w_n430_23[1]),.dout(n8370),.clk(gclk));
	jnot g08109(.din(w_n7959_0[0]),.dout(n8371),.clk(gclk));
	jor g08110(.dina(n8371),.dinb(w_n7957_0[0]),.dout(n8372),.clk(gclk));
	jor g08111(.dina(n8372),.dinb(w_n8058_20[1]),.dout(n8373),.clk(gclk));
	jxor g08112(.dina(n8373),.dinb(w_n7968_0[0]),.dout(n8374),.clk(gclk));
	jand g08113(.dina(w_n8363_0[1]),.dinb(w_n430_23[0]),.dout(n8375),.clk(gclk));
	jand g08114(.dina(n8375),.dinb(w_n8368_0[1]),.dout(n8376),.clk(gclk));
	jor g08115(.dina(w_n8376_0[1]),.dinb(w_n8374_0[1]),.dout(n8377),.clk(gclk));
	jand g08116(.dina(w_n8377_0[1]),.dinb(w_n8370_0[1]),.dout(n8378),.clk(gclk));
	jor g08117(.dina(w_n8378_0[2]),.dinb(w_n425_22[1]),.dout(n8379),.clk(gclk));
	jand g08118(.dina(w_n8378_0[1]),.dinb(w_n425_22[0]),.dout(n8380),.clk(gclk));
	jnot g08119(.din(w_n7971_0[0]),.dout(n8381),.clk(gclk));
	jand g08120(.dina(w_asqrt25_16[1]),.dinb(n8381),.dout(n8382),.clk(gclk));
	jand g08121(.dina(w_n8382_0[1]),.dinb(w_n7976_0[0]),.dout(n8383),.clk(gclk));
	jor g08122(.dina(n8383),.dinb(w_n7975_0[0]),.dout(n8384),.clk(gclk));
	jand g08123(.dina(w_n8382_0[0]),.dinb(w_n7977_0[0]),.dout(n8385),.clk(gclk));
	jnot g08124(.din(n8385),.dout(n8386),.clk(gclk));
	jand g08125(.dina(n8386),.dinb(n8384),.dout(n8387),.clk(gclk));
	jnot g08126(.din(n8387),.dout(n8388),.clk(gclk));
	jor g08127(.dina(w_n8388_0[1]),.dinb(n8380),.dout(n8389),.clk(gclk));
	jand g08128(.dina(w_n8389_0[1]),.dinb(w_n8379_0[1]),.dout(n8390),.clk(gclk));
	jor g08129(.dina(n8390),.dinb(w_n305_24[0]),.dout(n8391),.clk(gclk));
	jand g08130(.dina(w_n8379_0[0]),.dinb(w_n305_23[2]),.dout(n8392),.clk(gclk));
	jand g08131(.dina(n8392),.dinb(w_n8389_0[0]),.dout(n8393),.clk(gclk));
	jnot g08132(.din(w_n7979_0[0]),.dout(n8394),.clk(gclk));
	jand g08133(.dina(w_asqrt25_16[0]),.dinb(n8394),.dout(n8395),.clk(gclk));
	jand g08134(.dina(w_n8395_0[1]),.dinb(w_n7986_0[0]),.dout(n8396),.clk(gclk));
	jor g08135(.dina(n8396),.dinb(w_n7984_0[0]),.dout(n8397),.clk(gclk));
	jand g08136(.dina(w_n8395_0[0]),.dinb(w_n7987_0[0]),.dout(n8398),.clk(gclk));
	jnot g08137(.din(n8398),.dout(n8399),.clk(gclk));
	jand g08138(.dina(n8399),.dinb(n8397),.dout(n8400),.clk(gclk));
	jnot g08139(.din(n8400),.dout(n8401),.clk(gclk));
	jor g08140(.dina(w_n8401_0[1]),.dinb(w_n8393_0[1]),.dout(n8402),.clk(gclk));
	jand g08141(.dina(n8402),.dinb(w_n8391_0[1]),.dout(n8403),.clk(gclk));
	jor g08142(.dina(w_n8403_0[1]),.dinb(w_n290_23[1]),.dout(n8404),.clk(gclk));
	jxor g08143(.dina(w_n7988_0[0]),.dinb(w_n305_23[1]),.dout(n8405),.clk(gclk));
	jor g08144(.dina(n8405),.dinb(w_n8058_20[0]),.dout(n8406),.clk(gclk));
	jxor g08145(.dina(n8406),.dinb(w_n7999_0[0]),.dout(n8407),.clk(gclk));
	jand g08146(.dina(w_n8403_0[0]),.dinb(w_n290_23[0]),.dout(n8408),.clk(gclk));
	jor g08147(.dina(w_n8408_0[1]),.dinb(w_n8407_0[1]),.dout(n8409),.clk(gclk));
	jand g08148(.dina(w_n8409_0[2]),.dinb(w_n8404_0[2]),.dout(n8410),.clk(gclk));
	jor g08149(.dina(n8410),.dinb(w_n223_23[2]),.dout(n8411),.clk(gclk));
	jnot g08150(.din(w_n8004_0[0]),.dout(n8412),.clk(gclk));
	jor g08151(.dina(n8412),.dinb(w_n8002_0[0]),.dout(n8413),.clk(gclk));
	jor g08152(.dina(n8413),.dinb(w_n8058_19[2]),.dout(n8414),.clk(gclk));
	jxor g08153(.dina(n8414),.dinb(w_n8013_0[0]),.dout(n8415),.clk(gclk));
	jand g08154(.dina(w_n8404_0[1]),.dinb(w_n223_23[1]),.dout(n8416),.clk(gclk));
	jand g08155(.dina(n8416),.dinb(w_n8409_0[1]),.dout(n8417),.clk(gclk));
	jor g08156(.dina(w_n8417_0[1]),.dinb(w_n8415_0[1]),.dout(n8418),.clk(gclk));
	jand g08157(.dina(w_n8418_0[1]),.dinb(w_n8411_0[1]),.dout(n8419),.clk(gclk));
	jor g08158(.dina(w_n8419_0[2]),.dinb(w_n199_27[1]),.dout(n8420),.clk(gclk));
	jand g08159(.dina(w_n8419_0[1]),.dinb(w_n199_27[0]),.dout(n8421),.clk(gclk));
	jnot g08160(.din(w_n8016_0[0]),.dout(n8422),.clk(gclk));
	jand g08161(.dina(w_asqrt25_15[2]),.dinb(n8422),.dout(n8423),.clk(gclk));
	jand g08162(.dina(w_n8423_0[1]),.dinb(w_n8021_0[0]),.dout(n8424),.clk(gclk));
	jor g08163(.dina(n8424),.dinb(w_n8020_0[0]),.dout(n8425),.clk(gclk));
	jand g08164(.dina(w_n8423_0[0]),.dinb(w_n8022_0[0]),.dout(n8426),.clk(gclk));
	jnot g08165(.din(n8426),.dout(n8427),.clk(gclk));
	jand g08166(.dina(n8427),.dinb(n8425),.dout(n8428),.clk(gclk));
	jnot g08167(.din(n8428),.dout(n8429),.clk(gclk));
	jor g08168(.dina(w_n8429_0[1]),.dinb(n8421),.dout(n8430),.clk(gclk));
	jand g08169(.dina(n8430),.dinb(n8420),.dout(n8431),.clk(gclk));
	jnot g08170(.din(w_n8024_0[0]),.dout(n8432),.clk(gclk));
	jand g08171(.dina(w_asqrt25_15[1]),.dinb(n8432),.dout(n8433),.clk(gclk));
	jand g08172(.dina(w_n8433_0[1]),.dinb(w_n8031_0[0]),.dout(n8434),.clk(gclk));
	jor g08173(.dina(n8434),.dinb(w_n8029_0[0]),.dout(n8435),.clk(gclk));
	jand g08174(.dina(w_n8433_0[0]),.dinb(w_n8032_0[0]),.dout(n8436),.clk(gclk));
	jnot g08175(.din(n8436),.dout(n8437),.clk(gclk));
	jand g08176(.dina(n8437),.dinb(n8435),.dout(n8438),.clk(gclk));
	jnot g08177(.din(w_n8438_0[2]),.dout(n8439),.clk(gclk));
	jand g08178(.dina(w_asqrt25_15[0]),.dinb(w_n8046_0[1]),.dout(n8440),.clk(gclk));
	jand g08179(.dina(w_n8440_0[1]),.dinb(w_n8033_1[0]),.dout(n8441),.clk(gclk));
	jor g08180(.dina(n8441),.dinb(w_n8080_0[0]),.dout(n8442),.clk(gclk));
	jor g08181(.dina(n8442),.dinb(w_n8439_0[1]),.dout(n8443),.clk(gclk));
	jor g08182(.dina(n8443),.dinb(w_n8431_0[2]),.dout(n8444),.clk(gclk));
	jand g08183(.dina(n8444),.dinb(w_n194_26[1]),.dout(n8445),.clk(gclk));
	jand g08184(.dina(w_n8439_0[0]),.dinb(w_n8431_0[1]),.dout(n8446),.clk(gclk));
	jor g08185(.dina(w_n8440_0[0]),.dinb(w_n8033_0[2]),.dout(n8447),.clk(gclk));
	jand g08186(.dina(w_n8046_0[0]),.dinb(w_n8033_0[1]),.dout(n8448),.clk(gclk));
	jor g08187(.dina(n8448),.dinb(w_n194_26[0]),.dout(n8449),.clk(gclk));
	jnot g08188(.din(n8449),.dout(n8450),.clk(gclk));
	jand g08189(.dina(n8450),.dinb(n8447),.dout(n8451),.clk(gclk));
	jor g08190(.dina(w_n8451_0[1]),.dinb(w_n8446_0[2]),.dout(n8454),.clk(gclk));
	jor g08191(.dina(n8454),.dinb(w_n8445_0[1]),.dout(asqrt_fa_25),.clk(gclk));
	jxor g08192(.dina(w_n8185_0[0]),.dinb(w_n3907_17[2]),.dout(n8456),.clk(gclk));
	jand g08193(.dina(n8456),.dinb(w_asqrt24_31),.dout(n8457),.clk(gclk));
	jxor g08194(.dina(n8457),.dinb(w_n8061_0[0]),.dout(n8458),.clk(gclk));
	jand g08195(.dina(w_asqrt24_30[2]),.dinb(w_a48_0[0]),.dout(n8459),.clk(gclk));
	jnot g08196(.din(w_a46_0[1]),.dout(n8460),.clk(gclk));
	jnot g08197(.din(w_a47_0[1]),.dout(n8461),.clk(gclk));
	jand g08198(.dina(w_n8063_1[0]),.dinb(w_n8461_0[1]),.dout(n8462),.clk(gclk));
	jand g08199(.dina(n8462),.dinb(w_n8460_1[1]),.dout(n8463),.clk(gclk));
	jor g08200(.dina(n8463),.dinb(n8459),.dout(n8464),.clk(gclk));
	jand g08201(.dina(w_n8464_0[2]),.dinb(w_asqrt25_14[2]),.dout(n8465),.clk(gclk));
	jand g08202(.dina(w_asqrt24_30[1]),.dinb(w_n8063_0[2]),.dout(n8466),.clk(gclk));
	jxor g08203(.dina(w_n8466_0[1]),.dinb(w_n8064_0[1]),.dout(n8467),.clk(gclk));
	jor g08204(.dina(w_n8464_0[1]),.dinb(w_asqrt25_14[1]),.dout(n8468),.clk(gclk));
	jand g08205(.dina(n8468),.dinb(w_n8467_0[1]),.dout(n8469),.clk(gclk));
	jor g08206(.dina(w_n8469_0[1]),.dinb(w_n8465_0[1]),.dout(n8470),.clk(gclk));
	jand g08207(.dina(n8470),.dinb(w_asqrt26_18[0]),.dout(n8471),.clk(gclk));
	jor g08208(.dina(w_n8465_0[0]),.dinb(w_asqrt26_17[2]),.dout(n8472),.clk(gclk));
	jor g08209(.dina(n8472),.dinb(w_n8469_0[0]),.dout(n8473),.clk(gclk));
	jand g08210(.dina(w_n8466_0[0]),.dinb(w_n8064_0[0]),.dout(n8474),.clk(gclk));
	jnot g08211(.din(w_n8445_0[0]),.dout(n8475),.clk(gclk));
	jnot g08212(.din(w_n8446_0[1]),.dout(n8476),.clk(gclk));
	jnot g08213(.din(w_n8451_0[0]),.dout(n8477),.clk(gclk));
	jand g08214(.dina(n8477),.dinb(w_asqrt25_14[0]),.dout(n8478),.clk(gclk));
	jand g08215(.dina(n8478),.dinb(n8476),.dout(n8479),.clk(gclk));
	jand g08216(.dina(n8479),.dinb(n8475),.dout(n8480),.clk(gclk));
	jor g08217(.dina(n8480),.dinb(n8474),.dout(n8481),.clk(gclk));
	jxor g08218(.dina(n8481),.dinb(w_n7647_0[1]),.dout(n8482),.clk(gclk));
	jand g08219(.dina(w_n8482_0[1]),.dinb(w_n8473_0[1]),.dout(n8483),.clk(gclk));
	jor g08220(.dina(n8483),.dinb(w_n8471_0[1]),.dout(n8484),.clk(gclk));
	jand g08221(.dina(w_n8484_0[2]),.dinb(w_asqrt27_14[1]),.dout(n8485),.clk(gclk));
	jor g08222(.dina(w_n8484_0[1]),.dinb(w_asqrt27_14[0]),.dout(n8486),.clk(gclk));
	jxor g08223(.dina(w_n8068_0[0]),.dinb(w_n8053_15[2]),.dout(n8487),.clk(gclk));
	jand g08224(.dina(n8487),.dinb(w_asqrt24_30[0]),.dout(n8488),.clk(gclk));
	jxor g08225(.dina(n8488),.dinb(w_n8071_0[0]),.dout(n8489),.clk(gclk));
	jnot g08226(.din(w_n8489_0[1]),.dout(n8490),.clk(gclk));
	jand g08227(.dina(n8490),.dinb(n8486),.dout(n8491),.clk(gclk));
	jor g08228(.dina(w_n8491_0[1]),.dinb(w_n8485_0[1]),.dout(n8492),.clk(gclk));
	jand g08229(.dina(n8492),.dinb(w_asqrt28_18[0]),.dout(n8493),.clk(gclk));
	jnot g08230(.din(w_n8077_0[0]),.dout(n8494),.clk(gclk));
	jand g08231(.dina(n8494),.dinb(w_n8075_0[0]),.dout(n8495),.clk(gclk));
	jand g08232(.dina(n8495),.dinb(w_asqrt24_29[2]),.dout(n8496),.clk(gclk));
	jxor g08233(.dina(n8496),.dinb(w_n8085_0[0]),.dout(n8497),.clk(gclk));
	jnot g08234(.din(n8497),.dout(n8498),.clk(gclk));
	jor g08235(.dina(w_n8485_0[0]),.dinb(w_asqrt28_17[2]),.dout(n8499),.clk(gclk));
	jor g08236(.dina(n8499),.dinb(w_n8491_0[0]),.dout(n8500),.clk(gclk));
	jand g08237(.dina(w_n8500_0[1]),.dinb(w_n8498_0[1]),.dout(n8501),.clk(gclk));
	jor g08238(.dina(w_n8501_0[1]),.dinb(w_n8493_0[1]),.dout(n8502),.clk(gclk));
	jand g08239(.dina(w_n8502_0[2]),.dinb(w_asqrt29_14[2]),.dout(n8503),.clk(gclk));
	jor g08240(.dina(w_n8502_0[1]),.dinb(w_asqrt29_14[1]),.dout(n8504),.clk(gclk));
	jnot g08241(.din(w_n8092_0[0]),.dout(n8505),.clk(gclk));
	jxor g08242(.dina(w_n8087_0[0]),.dinb(w_n7260_16[1]),.dout(n8506),.clk(gclk));
	jand g08243(.dina(n8506),.dinb(w_asqrt24_29[1]),.dout(n8507),.clk(gclk));
	jxor g08244(.dina(n8507),.dinb(n8505),.dout(n8508),.clk(gclk));
	jand g08245(.dina(w_n8508_0[1]),.dinb(n8504),.dout(n8509),.clk(gclk));
	jor g08246(.dina(w_n8509_0[1]),.dinb(w_n8503_0[1]),.dout(n8510),.clk(gclk));
	jand g08247(.dina(n8510),.dinb(w_asqrt30_18[0]),.dout(n8511),.clk(gclk));
	jor g08248(.dina(w_n8503_0[0]),.dinb(w_asqrt30_17[2]),.dout(n8512),.clk(gclk));
	jor g08249(.dina(n8512),.dinb(w_n8509_0[0]),.dout(n8513),.clk(gclk));
	jnot g08250(.din(w_n8099_0[0]),.dout(n8514),.clk(gclk));
	jnot g08251(.din(w_n8101_0[0]),.dout(n8515),.clk(gclk));
	jand g08252(.dina(w_asqrt24_29[0]),.dinb(w_n8095_0[0]),.dout(n8516),.clk(gclk));
	jand g08253(.dina(w_n8516_0[1]),.dinb(n8515),.dout(n8517),.clk(gclk));
	jor g08254(.dina(n8517),.dinb(n8514),.dout(n8518),.clk(gclk));
	jnot g08255(.din(w_n8102_0[0]),.dout(n8519),.clk(gclk));
	jand g08256(.dina(w_n8516_0[0]),.dinb(n8519),.dout(n8520),.clk(gclk));
	jnot g08257(.din(n8520),.dout(n8521),.clk(gclk));
	jand g08258(.dina(n8521),.dinb(n8518),.dout(n8522),.clk(gclk));
	jand g08259(.dina(w_n8522_0[1]),.dinb(w_n8513_0[1]),.dout(n8523),.clk(gclk));
	jor g08260(.dina(n8523),.dinb(w_n8511_0[1]),.dout(n8524),.clk(gclk));
	jand g08261(.dina(w_n8524_0[2]),.dinb(w_asqrt31_14[2]),.dout(n8525),.clk(gclk));
	jor g08262(.dina(w_n8524_0[1]),.dinb(w_asqrt31_14[1]),.dout(n8526),.clk(gclk));
	jxor g08263(.dina(w_n8103_0[0]),.dinb(w_n6500_16[1]),.dout(n8527),.clk(gclk));
	jand g08264(.dina(n8527),.dinb(w_asqrt24_28[2]),.dout(n8528),.clk(gclk));
	jxor g08265(.dina(n8528),.dinb(w_n8108_0[0]),.dout(n8529),.clk(gclk));
	jand g08266(.dina(w_n8529_0[1]),.dinb(n8526),.dout(n8530),.clk(gclk));
	jor g08267(.dina(w_n8530_0[1]),.dinb(w_n8525_0[1]),.dout(n8531),.clk(gclk));
	jand g08268(.dina(n8531),.dinb(w_asqrt32_18[0]),.dout(n8532),.clk(gclk));
	jnot g08269(.din(w_n8114_0[0]),.dout(n8533),.clk(gclk));
	jand g08270(.dina(n8533),.dinb(w_n8112_0[0]),.dout(n8534),.clk(gclk));
	jand g08271(.dina(n8534),.dinb(w_asqrt24_28[1]),.dout(n8535),.clk(gclk));
	jxor g08272(.dina(n8535),.dinb(w_n8123_0[0]),.dout(n8536),.clk(gclk));
	jnot g08273(.din(n8536),.dout(n8537),.clk(gclk));
	jor g08274(.dina(w_n8525_0[0]),.dinb(w_asqrt32_17[2]),.dout(n8538),.clk(gclk));
	jor g08275(.dina(n8538),.dinb(w_n8530_0[0]),.dout(n8539),.clk(gclk));
	jand g08276(.dina(w_n8539_0[1]),.dinb(w_n8537_0[1]),.dout(n8540),.clk(gclk));
	jor g08277(.dina(w_n8540_0[1]),.dinb(w_n8532_0[1]),.dout(n8541),.clk(gclk));
	jand g08278(.dina(w_n8541_0[2]),.dinb(w_asqrt33_15[0]),.dout(n8542),.clk(gclk));
	jor g08279(.dina(w_n8541_0[1]),.dinb(w_asqrt33_14[2]),.dout(n8543),.clk(gclk));
	jxor g08280(.dina(w_n8125_0[0]),.dinb(w_n5788_16[2]),.dout(n8544),.clk(gclk));
	jand g08281(.dina(n8544),.dinb(w_asqrt24_28[0]),.dout(n8545),.clk(gclk));
	jxor g08282(.dina(n8545),.dinb(w_n8131_0[0]),.dout(n8546),.clk(gclk));
	jand g08283(.dina(w_n8546_0[1]),.dinb(n8543),.dout(n8547),.clk(gclk));
	jor g08284(.dina(w_n8547_0[1]),.dinb(w_n8542_0[1]),.dout(n8548),.clk(gclk));
	jand g08285(.dina(n8548),.dinb(w_asqrt34_18[0]),.dout(n8549),.clk(gclk));
	jor g08286(.dina(w_n8542_0[0]),.dinb(w_asqrt34_17[2]),.dout(n8550),.clk(gclk));
	jor g08287(.dina(n8550),.dinb(w_n8547_0[0]),.dout(n8551),.clk(gclk));
	jnot g08288(.din(w_n8139_0[0]),.dout(n8552),.clk(gclk));
	jnot g08289(.din(w_n8141_0[0]),.dout(n8553),.clk(gclk));
	jand g08290(.dina(w_asqrt24_27[2]),.dinb(w_n8135_0[0]),.dout(n8554),.clk(gclk));
	jand g08291(.dina(w_n8554_0[1]),.dinb(n8553),.dout(n8555),.clk(gclk));
	jor g08292(.dina(n8555),.dinb(n8552),.dout(n8556),.clk(gclk));
	jnot g08293(.din(w_n8142_0[0]),.dout(n8557),.clk(gclk));
	jand g08294(.dina(w_n8554_0[0]),.dinb(n8557),.dout(n8558),.clk(gclk));
	jnot g08295(.din(n8558),.dout(n8559),.clk(gclk));
	jand g08296(.dina(n8559),.dinb(n8556),.dout(n8560),.clk(gclk));
	jand g08297(.dina(w_n8560_0[1]),.dinb(w_n8551_0[1]),.dout(n8561),.clk(gclk));
	jor g08298(.dina(n8561),.dinb(w_n8549_0[1]),.dout(n8562),.clk(gclk));
	jand g08299(.dina(w_n8562_0[1]),.dinb(w_asqrt35_15[0]),.dout(n8563),.clk(gclk));
	jxor g08300(.dina(w_n8143_0[0]),.dinb(w_n5116_16[2]),.dout(n8564),.clk(gclk));
	jand g08301(.dina(n8564),.dinb(w_asqrt24_27[1]),.dout(n8565),.clk(gclk));
	jxor g08302(.dina(n8565),.dinb(w_n8150_0[0]),.dout(n8566),.clk(gclk));
	jnot g08303(.din(n8566),.dout(n8567),.clk(gclk));
	jor g08304(.dina(w_n8562_0[0]),.dinb(w_asqrt35_14[2]),.dout(n8568),.clk(gclk));
	jand g08305(.dina(w_n8568_0[1]),.dinb(w_n8567_0[1]),.dout(n8569),.clk(gclk));
	jor g08306(.dina(w_n8569_0[2]),.dinb(w_n8563_0[2]),.dout(n8570),.clk(gclk));
	jand g08307(.dina(n8570),.dinb(w_asqrt36_18[0]),.dout(n8571),.clk(gclk));
	jnot g08308(.din(w_n8155_0[0]),.dout(n8572),.clk(gclk));
	jand g08309(.dina(n8572),.dinb(w_n8153_0[0]),.dout(n8573),.clk(gclk));
	jand g08310(.dina(n8573),.dinb(w_asqrt24_27[0]),.dout(n8574),.clk(gclk));
	jxor g08311(.dina(n8574),.dinb(w_n8163_0[0]),.dout(n8575),.clk(gclk));
	jnot g08312(.din(n8575),.dout(n8576),.clk(gclk));
	jor g08313(.dina(w_n8563_0[1]),.dinb(w_asqrt36_17[2]),.dout(n8577),.clk(gclk));
	jor g08314(.dina(n8577),.dinb(w_n8569_0[1]),.dout(n8578),.clk(gclk));
	jand g08315(.dina(w_n8578_0[1]),.dinb(w_n8576_0[1]),.dout(n8579),.clk(gclk));
	jor g08316(.dina(w_n8579_0[1]),.dinb(w_n8571_0[1]),.dout(n8580),.clk(gclk));
	jand g08317(.dina(w_n8580_0[2]),.dinb(w_asqrt37_15[1]),.dout(n8581),.clk(gclk));
	jor g08318(.dina(w_n8580_0[1]),.dinb(w_asqrt37_15[0]),.dout(n8582),.clk(gclk));
	jnot g08319(.din(w_n8169_0[0]),.dout(n8583),.clk(gclk));
	jnot g08320(.din(w_n8170_0[0]),.dout(n8584),.clk(gclk));
	jand g08321(.dina(w_asqrt24_26[2]),.dinb(w_n8166_0[0]),.dout(n8585),.clk(gclk));
	jand g08322(.dina(w_n8585_0[1]),.dinb(n8584),.dout(n8586),.clk(gclk));
	jor g08323(.dina(n8586),.dinb(n8583),.dout(n8587),.clk(gclk));
	jnot g08324(.din(w_n8171_0[0]),.dout(n8588),.clk(gclk));
	jand g08325(.dina(w_n8585_0[0]),.dinb(n8588),.dout(n8589),.clk(gclk));
	jnot g08326(.din(n8589),.dout(n8590),.clk(gclk));
	jand g08327(.dina(n8590),.dinb(n8587),.dout(n8591),.clk(gclk));
	jand g08328(.dina(w_n8591_0[1]),.dinb(n8582),.dout(n8592),.clk(gclk));
	jor g08329(.dina(w_n8592_0[1]),.dinb(w_n8581_0[1]),.dout(n8593),.clk(gclk));
	jand g08330(.dina(n8593),.dinb(w_asqrt38_18[0]),.dout(n8594),.clk(gclk));
	jnot g08331(.din(w_n8175_0[0]),.dout(n8595),.clk(gclk));
	jand g08332(.dina(n8595),.dinb(w_n8173_0[0]),.dout(n8596),.clk(gclk));
	jand g08333(.dina(n8596),.dinb(w_asqrt24_26[1]),.dout(n8597),.clk(gclk));
	jxor g08334(.dina(n8597),.dinb(w_n8183_0[0]),.dout(n8598),.clk(gclk));
	jnot g08335(.din(n8598),.dout(n8599),.clk(gclk));
	jor g08336(.dina(w_n8581_0[0]),.dinb(w_asqrt38_17[2]),.dout(n8600),.clk(gclk));
	jor g08337(.dina(n8600),.dinb(w_n8592_0[0]),.dout(n8601),.clk(gclk));
	jand g08338(.dina(w_n8601_0[1]),.dinb(w_n8599_0[1]),.dout(n8602),.clk(gclk));
	jor g08339(.dina(w_n8602_0[1]),.dinb(w_n8594_0[1]),.dout(n8603),.clk(gclk));
	jand g08340(.dina(w_n8603_0[2]),.dinb(w_asqrt39_15[1]),.dout(n8604),.clk(gclk));
	jnot g08341(.din(w_n8458_0[1]),.dout(n8605),.clk(gclk));
	jor g08342(.dina(w_n8603_0[1]),.dinb(w_asqrt39_15[0]),.dout(n8606),.clk(gclk));
	jand g08343(.dina(n8606),.dinb(n8605),.dout(n8607),.clk(gclk));
	jor g08344(.dina(w_n8607_0[1]),.dinb(w_n8604_0[1]),.dout(n8608),.clk(gclk));
	jand g08345(.dina(n8608),.dinb(w_asqrt40_18[0]),.dout(n8609),.clk(gclk));
	jor g08346(.dina(w_n8604_0[0]),.dinb(w_asqrt40_17[2]),.dout(n8610),.clk(gclk));
	jor g08347(.dina(n8610),.dinb(w_n8607_0[0]),.dout(n8611),.clk(gclk));
	jnot g08348(.din(w_n8194_0[0]),.dout(n8612),.clk(gclk));
	jnot g08349(.din(w_n8196_0[0]),.dout(n8613),.clk(gclk));
	jand g08350(.dina(w_asqrt24_26[0]),.dinb(w_n8190_0[0]),.dout(n8614),.clk(gclk));
	jand g08351(.dina(w_n8614_0[1]),.dinb(n8613),.dout(n8615),.clk(gclk));
	jor g08352(.dina(n8615),.dinb(n8612),.dout(n8616),.clk(gclk));
	jnot g08353(.din(w_n8197_0[0]),.dout(n8617),.clk(gclk));
	jand g08354(.dina(w_n8614_0[0]),.dinb(n8617),.dout(n8618),.clk(gclk));
	jnot g08355(.din(n8618),.dout(n8619),.clk(gclk));
	jand g08356(.dina(n8619),.dinb(n8616),.dout(n8620),.clk(gclk));
	jand g08357(.dina(w_n8620_0[1]),.dinb(w_n8611_0[1]),.dout(n8621),.clk(gclk));
	jor g08358(.dina(n8621),.dinb(w_n8609_0[1]),.dout(n8622),.clk(gclk));
	jand g08359(.dina(w_n8622_0[2]),.dinb(w_asqrt41_15[2]),.dout(n8623),.clk(gclk));
	jor g08360(.dina(w_n8622_0[1]),.dinb(w_asqrt41_15[1]),.dout(n8624),.clk(gclk));
	jnot g08361(.din(w_n8202_0[0]),.dout(n8625),.clk(gclk));
	jnot g08362(.din(w_n8203_0[0]),.dout(n8626),.clk(gclk));
	jand g08363(.dina(w_asqrt24_25[2]),.dinb(w_n8199_0[0]),.dout(n8627),.clk(gclk));
	jand g08364(.dina(w_n8627_0[1]),.dinb(n8626),.dout(n8628),.clk(gclk));
	jor g08365(.dina(n8628),.dinb(n8625),.dout(n8629),.clk(gclk));
	jnot g08366(.din(w_n8204_0[0]),.dout(n8630),.clk(gclk));
	jand g08367(.dina(w_n8627_0[0]),.dinb(n8630),.dout(n8631),.clk(gclk));
	jnot g08368(.din(n8631),.dout(n8632),.clk(gclk));
	jand g08369(.dina(n8632),.dinb(n8629),.dout(n8633),.clk(gclk));
	jand g08370(.dina(w_n8633_0[1]),.dinb(n8624),.dout(n8634),.clk(gclk));
	jor g08371(.dina(w_n8634_0[1]),.dinb(w_n8623_0[1]),.dout(n8635),.clk(gclk));
	jand g08372(.dina(n8635),.dinb(w_asqrt42_18[0]),.dout(n8636),.clk(gclk));
	jor g08373(.dina(w_n8623_0[0]),.dinb(w_asqrt42_17[2]),.dout(n8637),.clk(gclk));
	jor g08374(.dina(n8637),.dinb(w_n8634_0[0]),.dout(n8638),.clk(gclk));
	jnot g08375(.din(w_n8210_0[0]),.dout(n8639),.clk(gclk));
	jnot g08376(.din(w_n8212_0[0]),.dout(n8640),.clk(gclk));
	jand g08377(.dina(w_asqrt24_25[1]),.dinb(w_n8206_0[0]),.dout(n8641),.clk(gclk));
	jand g08378(.dina(w_n8641_0[1]),.dinb(n8640),.dout(n8642),.clk(gclk));
	jor g08379(.dina(n8642),.dinb(n8639),.dout(n8643),.clk(gclk));
	jnot g08380(.din(w_n8213_0[0]),.dout(n8644),.clk(gclk));
	jand g08381(.dina(w_n8641_0[0]),.dinb(n8644),.dout(n8645),.clk(gclk));
	jnot g08382(.din(n8645),.dout(n8646),.clk(gclk));
	jand g08383(.dina(n8646),.dinb(n8643),.dout(n8647),.clk(gclk));
	jand g08384(.dina(w_n8647_0[1]),.dinb(w_n8638_0[1]),.dout(n8648),.clk(gclk));
	jor g08385(.dina(n8648),.dinb(w_n8636_0[1]),.dout(n8649),.clk(gclk));
	jand g08386(.dina(w_n8649_0[1]),.dinb(w_asqrt43_15[2]),.dout(n8650),.clk(gclk));
	jxor g08387(.dina(w_n8214_0[0]),.dinb(w_n2870_18[1]),.dout(n8651),.clk(gclk));
	jand g08388(.dina(n8651),.dinb(w_asqrt24_25[0]),.dout(n8652),.clk(gclk));
	jxor g08389(.dina(n8652),.dinb(w_n8224_0[0]),.dout(n8653),.clk(gclk));
	jnot g08390(.din(n8653),.dout(n8654),.clk(gclk));
	jor g08391(.dina(w_n8649_0[0]),.dinb(w_asqrt43_15[1]),.dout(n8655),.clk(gclk));
	jand g08392(.dina(w_n8655_0[1]),.dinb(w_n8654_0[1]),.dout(n8656),.clk(gclk));
	jor g08393(.dina(w_n8656_0[2]),.dinb(w_n8650_0[2]),.dout(n8657),.clk(gclk));
	jand g08394(.dina(n8657),.dinb(w_asqrt44_18[0]),.dout(n8658),.clk(gclk));
	jnot g08395(.din(w_n8229_0[0]),.dout(n8659),.clk(gclk));
	jand g08396(.dina(n8659),.dinb(w_n8227_0[0]),.dout(n8660),.clk(gclk));
	jand g08397(.dina(n8660),.dinb(w_asqrt24_24[2]),.dout(n8661),.clk(gclk));
	jxor g08398(.dina(n8661),.dinb(w_n8237_0[0]),.dout(n8662),.clk(gclk));
	jnot g08399(.din(n8662),.dout(n8663),.clk(gclk));
	jor g08400(.dina(w_n8650_0[1]),.dinb(w_asqrt44_17[2]),.dout(n8664),.clk(gclk));
	jor g08401(.dina(n8664),.dinb(w_n8656_0[1]),.dout(n8665),.clk(gclk));
	jand g08402(.dina(w_n8665_0[1]),.dinb(w_n8663_0[1]),.dout(n8666),.clk(gclk));
	jor g08403(.dina(w_n8666_0[1]),.dinb(w_n8658_0[1]),.dout(n8667),.clk(gclk));
	jand g08404(.dina(w_n8667_0[2]),.dinb(w_asqrt45_16[0]),.dout(n8668),.clk(gclk));
	jor g08405(.dina(w_n8667_0[1]),.dinb(w_asqrt45_15[2]),.dout(n8669),.clk(gclk));
	jnot g08406(.din(w_n8243_0[0]),.dout(n8670),.clk(gclk));
	jnot g08407(.din(w_n8244_0[0]),.dout(n8671),.clk(gclk));
	jand g08408(.dina(w_asqrt24_24[1]),.dinb(w_n8240_0[0]),.dout(n8672),.clk(gclk));
	jand g08409(.dina(w_n8672_0[1]),.dinb(n8671),.dout(n8673),.clk(gclk));
	jor g08410(.dina(n8673),.dinb(n8670),.dout(n8674),.clk(gclk));
	jnot g08411(.din(w_n8245_0[0]),.dout(n8675),.clk(gclk));
	jand g08412(.dina(w_n8672_0[0]),.dinb(n8675),.dout(n8676),.clk(gclk));
	jnot g08413(.din(n8676),.dout(n8677),.clk(gclk));
	jand g08414(.dina(n8677),.dinb(n8674),.dout(n8678),.clk(gclk));
	jand g08415(.dina(w_n8678_0[1]),.dinb(n8669),.dout(n8679),.clk(gclk));
	jor g08416(.dina(w_n8679_0[1]),.dinb(w_n8668_0[1]),.dout(n8680),.clk(gclk));
	jand g08417(.dina(n8680),.dinb(w_asqrt46_18[0]),.dout(n8681),.clk(gclk));
	jor g08418(.dina(w_n8668_0[0]),.dinb(w_asqrt46_17[2]),.dout(n8682),.clk(gclk));
	jor g08419(.dina(n8682),.dinb(w_n8679_0[0]),.dout(n8683),.clk(gclk));
	jnot g08420(.din(w_n8251_0[0]),.dout(n8684),.clk(gclk));
	jnot g08421(.din(w_n8253_0[0]),.dout(n8685),.clk(gclk));
	jand g08422(.dina(w_asqrt24_24[0]),.dinb(w_n8247_0[0]),.dout(n8686),.clk(gclk));
	jand g08423(.dina(w_n8686_0[1]),.dinb(n8685),.dout(n8687),.clk(gclk));
	jor g08424(.dina(n8687),.dinb(n8684),.dout(n8688),.clk(gclk));
	jnot g08425(.din(w_n8254_0[0]),.dout(n8689),.clk(gclk));
	jand g08426(.dina(w_n8686_0[0]),.dinb(n8689),.dout(n8690),.clk(gclk));
	jnot g08427(.din(n8690),.dout(n8691),.clk(gclk));
	jand g08428(.dina(n8691),.dinb(n8688),.dout(n8692),.clk(gclk));
	jand g08429(.dina(w_n8692_0[1]),.dinb(w_n8683_0[1]),.dout(n8693),.clk(gclk));
	jor g08430(.dina(n8693),.dinb(w_n8681_0[1]),.dout(n8694),.clk(gclk));
	jand g08431(.dina(w_n8694_0[1]),.dinb(w_asqrt47_16[0]),.dout(n8695),.clk(gclk));
	jxor g08432(.dina(w_n8255_0[0]),.dinb(w_n2005_19[1]),.dout(n8696),.clk(gclk));
	jand g08433(.dina(n8696),.dinb(w_asqrt24_23[2]),.dout(n8697),.clk(gclk));
	jxor g08434(.dina(n8697),.dinb(w_n8265_0[0]),.dout(n8698),.clk(gclk));
	jnot g08435(.din(n8698),.dout(n8699),.clk(gclk));
	jor g08436(.dina(w_n8694_0[0]),.dinb(w_asqrt47_15[2]),.dout(n8700),.clk(gclk));
	jand g08437(.dina(w_n8700_0[1]),.dinb(w_n8699_0[1]),.dout(n8701),.clk(gclk));
	jor g08438(.dina(w_n8701_0[2]),.dinb(w_n8695_0[2]),.dout(n8702),.clk(gclk));
	jand g08439(.dina(n8702),.dinb(w_asqrt48_18[0]),.dout(n8703),.clk(gclk));
	jnot g08440(.din(w_n8270_0[0]),.dout(n8704),.clk(gclk));
	jand g08441(.dina(n8704),.dinb(w_n8268_0[0]),.dout(n8705),.clk(gclk));
	jand g08442(.dina(n8705),.dinb(w_asqrt24_23[1]),.dout(n8706),.clk(gclk));
	jxor g08443(.dina(n8706),.dinb(w_n8278_0[0]),.dout(n8707),.clk(gclk));
	jnot g08444(.din(n8707),.dout(n8708),.clk(gclk));
	jor g08445(.dina(w_n8695_0[1]),.dinb(w_asqrt48_17[2]),.dout(n8709),.clk(gclk));
	jor g08446(.dina(n8709),.dinb(w_n8701_0[1]),.dout(n8710),.clk(gclk));
	jand g08447(.dina(w_n8710_0[1]),.dinb(w_n8708_0[1]),.dout(n8711),.clk(gclk));
	jor g08448(.dina(w_n8711_0[1]),.dinb(w_n8703_0[1]),.dout(n8712),.clk(gclk));
	jand g08449(.dina(w_n8712_0[2]),.dinb(w_asqrt49_16[1]),.dout(n8713),.clk(gclk));
	jor g08450(.dina(w_n8712_0[1]),.dinb(w_asqrt49_16[0]),.dout(n8714),.clk(gclk));
	jnot g08451(.din(w_n8284_0[0]),.dout(n8715),.clk(gclk));
	jnot g08452(.din(w_n8285_0[0]),.dout(n8716),.clk(gclk));
	jand g08453(.dina(w_asqrt24_23[0]),.dinb(w_n8281_0[0]),.dout(n8717),.clk(gclk));
	jand g08454(.dina(w_n8717_0[1]),.dinb(n8716),.dout(n8718),.clk(gclk));
	jor g08455(.dina(n8718),.dinb(n8715),.dout(n8719),.clk(gclk));
	jnot g08456(.din(w_n8286_0[0]),.dout(n8720),.clk(gclk));
	jand g08457(.dina(w_n8717_0[0]),.dinb(n8720),.dout(n8721),.clk(gclk));
	jnot g08458(.din(n8721),.dout(n8722),.clk(gclk));
	jand g08459(.dina(n8722),.dinb(n8719),.dout(n8723),.clk(gclk));
	jand g08460(.dina(w_n8723_0[1]),.dinb(n8714),.dout(n8724),.clk(gclk));
	jor g08461(.dina(w_n8724_0[1]),.dinb(w_n8713_0[1]),.dout(n8725),.clk(gclk));
	jand g08462(.dina(n8725),.dinb(w_asqrt50_18[0]),.dout(n8726),.clk(gclk));
	jor g08463(.dina(w_n8713_0[0]),.dinb(w_asqrt50_17[2]),.dout(n8727),.clk(gclk));
	jor g08464(.dina(n8727),.dinb(w_n8724_0[0]),.dout(n8728),.clk(gclk));
	jnot g08465(.din(w_n8292_0[0]),.dout(n8729),.clk(gclk));
	jnot g08466(.din(w_n8294_0[0]),.dout(n8730),.clk(gclk));
	jand g08467(.dina(w_asqrt24_22[2]),.dinb(w_n8288_0[0]),.dout(n8731),.clk(gclk));
	jand g08468(.dina(w_n8731_0[1]),.dinb(n8730),.dout(n8732),.clk(gclk));
	jor g08469(.dina(n8732),.dinb(n8729),.dout(n8733),.clk(gclk));
	jnot g08470(.din(w_n8295_0[0]),.dout(n8734),.clk(gclk));
	jand g08471(.dina(w_n8731_0[0]),.dinb(n8734),.dout(n8735),.clk(gclk));
	jnot g08472(.din(n8735),.dout(n8736),.clk(gclk));
	jand g08473(.dina(n8736),.dinb(n8733),.dout(n8737),.clk(gclk));
	jand g08474(.dina(w_n8737_0[1]),.dinb(w_n8728_0[1]),.dout(n8738),.clk(gclk));
	jor g08475(.dina(n8738),.dinb(w_n8726_0[1]),.dout(n8739),.clk(gclk));
	jand g08476(.dina(w_n8739_0[1]),.dinb(w_asqrt51_16[1]),.dout(n8740),.clk(gclk));
	jxor g08477(.dina(w_n8296_0[0]),.dinb(w_n1312_20[0]),.dout(n8741),.clk(gclk));
	jand g08478(.dina(n8741),.dinb(w_asqrt24_22[1]),.dout(n8742),.clk(gclk));
	jxor g08479(.dina(n8742),.dinb(w_n8306_0[0]),.dout(n8743),.clk(gclk));
	jnot g08480(.din(n8743),.dout(n8744),.clk(gclk));
	jor g08481(.dina(w_n8739_0[0]),.dinb(w_asqrt51_16[0]),.dout(n8745),.clk(gclk));
	jand g08482(.dina(w_n8745_0[1]),.dinb(w_n8744_0[1]),.dout(n8746),.clk(gclk));
	jor g08483(.dina(w_n8746_0[2]),.dinb(w_n8740_0[2]),.dout(n8747),.clk(gclk));
	jand g08484(.dina(n8747),.dinb(w_asqrt52_18[0]),.dout(n8748),.clk(gclk));
	jnot g08485(.din(w_n8311_0[0]),.dout(n8749),.clk(gclk));
	jand g08486(.dina(n8749),.dinb(w_n8309_0[0]),.dout(n8750),.clk(gclk));
	jand g08487(.dina(n8750),.dinb(w_asqrt24_22[0]),.dout(n8751),.clk(gclk));
	jxor g08488(.dina(n8751),.dinb(w_n8319_0[0]),.dout(n8752),.clk(gclk));
	jnot g08489(.din(n8752),.dout(n8753),.clk(gclk));
	jor g08490(.dina(w_n8740_0[1]),.dinb(w_asqrt52_17[2]),.dout(n8754),.clk(gclk));
	jor g08491(.dina(n8754),.dinb(w_n8746_0[1]),.dout(n8755),.clk(gclk));
	jand g08492(.dina(w_n8755_0[1]),.dinb(w_n8753_0[1]),.dout(n8756),.clk(gclk));
	jor g08493(.dina(w_n8756_0[1]),.dinb(w_n8748_0[1]),.dout(n8757),.clk(gclk));
	jand g08494(.dina(w_n8757_0[2]),.dinb(w_asqrt53_16[2]),.dout(n8758),.clk(gclk));
	jor g08495(.dina(w_n8757_0[1]),.dinb(w_asqrt53_16[1]),.dout(n8759),.clk(gclk));
	jnot g08496(.din(w_n8325_0[0]),.dout(n8760),.clk(gclk));
	jnot g08497(.din(w_n8326_0[0]),.dout(n8761),.clk(gclk));
	jand g08498(.dina(w_asqrt24_21[2]),.dinb(w_n8322_0[0]),.dout(n8762),.clk(gclk));
	jand g08499(.dina(w_n8762_0[1]),.dinb(n8761),.dout(n8763),.clk(gclk));
	jor g08500(.dina(n8763),.dinb(n8760),.dout(n8764),.clk(gclk));
	jnot g08501(.din(w_n8327_0[0]),.dout(n8765),.clk(gclk));
	jand g08502(.dina(w_n8762_0[0]),.dinb(n8765),.dout(n8766),.clk(gclk));
	jnot g08503(.din(n8766),.dout(n8767),.clk(gclk));
	jand g08504(.dina(n8767),.dinb(n8764),.dout(n8768),.clk(gclk));
	jand g08505(.dina(w_n8768_0[1]),.dinb(n8759),.dout(n8769),.clk(gclk));
	jor g08506(.dina(w_n8769_0[1]),.dinb(w_n8758_0[1]),.dout(n8770),.clk(gclk));
	jand g08507(.dina(n8770),.dinb(w_asqrt54_18[0]),.dout(n8771),.clk(gclk));
	jor g08508(.dina(w_n8758_0[0]),.dinb(w_asqrt54_17[2]),.dout(n8772),.clk(gclk));
	jor g08509(.dina(n8772),.dinb(w_n8769_0[0]),.dout(n8773),.clk(gclk));
	jnot g08510(.din(w_n8333_0[0]),.dout(n8774),.clk(gclk));
	jnot g08511(.din(w_n8335_0[0]),.dout(n8775),.clk(gclk));
	jand g08512(.dina(w_asqrt24_21[1]),.dinb(w_n8329_0[0]),.dout(n8776),.clk(gclk));
	jand g08513(.dina(w_n8776_0[1]),.dinb(n8775),.dout(n8777),.clk(gclk));
	jor g08514(.dina(n8777),.dinb(n8774),.dout(n8778),.clk(gclk));
	jnot g08515(.din(w_n8336_0[0]),.dout(n8779),.clk(gclk));
	jand g08516(.dina(w_n8776_0[0]),.dinb(n8779),.dout(n8780),.clk(gclk));
	jnot g08517(.din(n8780),.dout(n8781),.clk(gclk));
	jand g08518(.dina(n8781),.dinb(n8778),.dout(n8782),.clk(gclk));
	jand g08519(.dina(w_n8782_0[1]),.dinb(w_n8773_0[1]),.dout(n8783),.clk(gclk));
	jor g08520(.dina(n8783),.dinb(w_n8771_0[1]),.dout(n8784),.clk(gclk));
	jand g08521(.dina(w_n8784_0[1]),.dinb(w_asqrt55_17[0]),.dout(n8785),.clk(gclk));
	jxor g08522(.dina(w_n8337_0[0]),.dinb(w_n791_21[0]),.dout(n8786),.clk(gclk));
	jand g08523(.dina(n8786),.dinb(w_asqrt24_21[0]),.dout(n8787),.clk(gclk));
	jxor g08524(.dina(n8787),.dinb(w_n8347_0[0]),.dout(n8788),.clk(gclk));
	jnot g08525(.din(n8788),.dout(n8789),.clk(gclk));
	jor g08526(.dina(w_n8784_0[0]),.dinb(w_asqrt55_16[2]),.dout(n8790),.clk(gclk));
	jand g08527(.dina(w_n8790_0[1]),.dinb(w_n8789_0[1]),.dout(n8791),.clk(gclk));
	jor g08528(.dina(w_n8791_0[2]),.dinb(w_n8785_0[2]),.dout(n8792),.clk(gclk));
	jand g08529(.dina(n8792),.dinb(w_asqrt56_18[0]),.dout(n8793),.clk(gclk));
	jnot g08530(.din(w_n8352_0[0]),.dout(n8794),.clk(gclk));
	jand g08531(.dina(n8794),.dinb(w_n8350_0[0]),.dout(n8795),.clk(gclk));
	jand g08532(.dina(n8795),.dinb(w_asqrt24_20[2]),.dout(n8796),.clk(gclk));
	jxor g08533(.dina(n8796),.dinb(w_n8360_0[0]),.dout(n8797),.clk(gclk));
	jnot g08534(.din(n8797),.dout(n8798),.clk(gclk));
	jor g08535(.dina(w_n8785_0[1]),.dinb(w_asqrt56_17[2]),.dout(n8799),.clk(gclk));
	jor g08536(.dina(n8799),.dinb(w_n8791_0[1]),.dout(n8800),.clk(gclk));
	jand g08537(.dina(w_n8800_0[1]),.dinb(w_n8798_0[1]),.dout(n8801),.clk(gclk));
	jor g08538(.dina(w_n8801_0[1]),.dinb(w_n8793_0[1]),.dout(n8802),.clk(gclk));
	jand g08539(.dina(w_n8802_0[2]),.dinb(w_asqrt57_17[1]),.dout(n8803),.clk(gclk));
	jor g08540(.dina(w_n8802_0[1]),.dinb(w_asqrt57_17[0]),.dout(n8804),.clk(gclk));
	jnot g08541(.din(w_n8366_0[0]),.dout(n8805),.clk(gclk));
	jnot g08542(.din(w_n8367_0[0]),.dout(n8806),.clk(gclk));
	jand g08543(.dina(w_asqrt24_20[1]),.dinb(w_n8363_0[0]),.dout(n8807),.clk(gclk));
	jand g08544(.dina(w_n8807_0[1]),.dinb(n8806),.dout(n8808),.clk(gclk));
	jor g08545(.dina(n8808),.dinb(n8805),.dout(n8809),.clk(gclk));
	jnot g08546(.din(w_n8368_0[0]),.dout(n8810),.clk(gclk));
	jand g08547(.dina(w_n8807_0[0]),.dinb(n8810),.dout(n8811),.clk(gclk));
	jnot g08548(.din(n8811),.dout(n8812),.clk(gclk));
	jand g08549(.dina(n8812),.dinb(n8809),.dout(n8813),.clk(gclk));
	jand g08550(.dina(w_n8813_0[1]),.dinb(n8804),.dout(n8814),.clk(gclk));
	jor g08551(.dina(w_n8814_0[1]),.dinb(w_n8803_0[1]),.dout(n8815),.clk(gclk));
	jand g08552(.dina(n8815),.dinb(w_asqrt58_18[0]),.dout(n8816),.clk(gclk));
	jor g08553(.dina(w_n8803_0[0]),.dinb(w_asqrt58_17[2]),.dout(n8817),.clk(gclk));
	jor g08554(.dina(n8817),.dinb(w_n8814_0[0]),.dout(n8818),.clk(gclk));
	jnot g08555(.din(w_n8374_0[0]),.dout(n8819),.clk(gclk));
	jnot g08556(.din(w_n8376_0[0]),.dout(n8820),.clk(gclk));
	jand g08557(.dina(w_asqrt24_20[0]),.dinb(w_n8370_0[0]),.dout(n8821),.clk(gclk));
	jand g08558(.dina(w_n8821_0[1]),.dinb(n8820),.dout(n8822),.clk(gclk));
	jor g08559(.dina(n8822),.dinb(n8819),.dout(n8823),.clk(gclk));
	jnot g08560(.din(w_n8377_0[0]),.dout(n8824),.clk(gclk));
	jand g08561(.dina(w_n8821_0[0]),.dinb(n8824),.dout(n8825),.clk(gclk));
	jnot g08562(.din(n8825),.dout(n8826),.clk(gclk));
	jand g08563(.dina(n8826),.dinb(n8823),.dout(n8827),.clk(gclk));
	jand g08564(.dina(w_n8827_0[1]),.dinb(w_n8818_0[1]),.dout(n8828),.clk(gclk));
	jor g08565(.dina(n8828),.dinb(w_n8816_0[1]),.dout(n8829),.clk(gclk));
	jand g08566(.dina(w_n8829_0[1]),.dinb(w_asqrt59_17[2]),.dout(n8830),.clk(gclk));
	jxor g08567(.dina(w_n8378_0[0]),.dinb(w_n425_21[2]),.dout(n8831),.clk(gclk));
	jand g08568(.dina(n8831),.dinb(w_asqrt24_19[2]),.dout(n8832),.clk(gclk));
	jxor g08569(.dina(n8832),.dinb(w_n8388_0[0]),.dout(n8833),.clk(gclk));
	jnot g08570(.din(n8833),.dout(n8834),.clk(gclk));
	jor g08571(.dina(w_n8829_0[0]),.dinb(w_asqrt59_17[1]),.dout(n8835),.clk(gclk));
	jand g08572(.dina(w_n8835_0[1]),.dinb(w_n8834_0[1]),.dout(n8836),.clk(gclk));
	jor g08573(.dina(w_n8836_0[2]),.dinb(w_n8830_0[2]),.dout(n8837),.clk(gclk));
	jand g08574(.dina(n8837),.dinb(w_asqrt60_17[2]),.dout(n8838),.clk(gclk));
	jnot g08575(.din(w_n8393_0[0]),.dout(n8839),.clk(gclk));
	jand g08576(.dina(n8839),.dinb(w_n8391_0[0]),.dout(n8840),.clk(gclk));
	jand g08577(.dina(n8840),.dinb(w_asqrt24_19[1]),.dout(n8841),.clk(gclk));
	jxor g08578(.dina(n8841),.dinb(w_n8401_0[0]),.dout(n8842),.clk(gclk));
	jnot g08579(.din(n8842),.dout(n8843),.clk(gclk));
	jor g08580(.dina(w_n8830_0[1]),.dinb(w_asqrt60_17[1]),.dout(n8844),.clk(gclk));
	jor g08581(.dina(n8844),.dinb(w_n8836_0[1]),.dout(n8845),.clk(gclk));
	jand g08582(.dina(w_n8845_0[1]),.dinb(w_n8843_0[1]),.dout(n8846),.clk(gclk));
	jor g08583(.dina(w_n8846_0[1]),.dinb(w_n8838_0[1]),.dout(n8847),.clk(gclk));
	jand g08584(.dina(w_n8847_0[2]),.dinb(w_asqrt61_18[0]),.dout(n8848),.clk(gclk));
	jor g08585(.dina(w_n8847_0[1]),.dinb(w_asqrt61_17[2]),.dout(n8849),.clk(gclk));
	jnot g08586(.din(w_n8407_0[0]),.dout(n8850),.clk(gclk));
	jnot g08587(.din(w_n8408_0[0]),.dout(n8851),.clk(gclk));
	jand g08588(.dina(w_asqrt24_19[0]),.dinb(w_n8404_0[0]),.dout(n8852),.clk(gclk));
	jand g08589(.dina(w_n8852_0[1]),.dinb(n8851),.dout(n8853),.clk(gclk));
	jor g08590(.dina(n8853),.dinb(n8850),.dout(n8854),.clk(gclk));
	jnot g08591(.din(w_n8409_0[0]),.dout(n8855),.clk(gclk));
	jand g08592(.dina(w_n8852_0[0]),.dinb(n8855),.dout(n8856),.clk(gclk));
	jnot g08593(.din(n8856),.dout(n8857),.clk(gclk));
	jand g08594(.dina(n8857),.dinb(n8854),.dout(n8858),.clk(gclk));
	jand g08595(.dina(w_n8858_0[1]),.dinb(n8849),.dout(n8859),.clk(gclk));
	jor g08596(.dina(w_n8859_0[1]),.dinb(w_n8848_0[1]),.dout(n8860),.clk(gclk));
	jand g08597(.dina(n8860),.dinb(w_asqrt62_18[0]),.dout(n8861),.clk(gclk));
	jor g08598(.dina(w_n8848_0[0]),.dinb(w_asqrt62_17[2]),.dout(n8862),.clk(gclk));
	jor g08599(.dina(n8862),.dinb(w_n8859_0[0]),.dout(n8863),.clk(gclk));
	jnot g08600(.din(w_n8415_0[0]),.dout(n8864),.clk(gclk));
	jnot g08601(.din(w_n8417_0[0]),.dout(n8865),.clk(gclk));
	jand g08602(.dina(w_asqrt24_18[2]),.dinb(w_n8411_0[0]),.dout(n8866),.clk(gclk));
	jand g08603(.dina(w_n8866_0[1]),.dinb(n8865),.dout(n8867),.clk(gclk));
	jor g08604(.dina(n8867),.dinb(n8864),.dout(n8868),.clk(gclk));
	jnot g08605(.din(w_n8418_0[0]),.dout(n8869),.clk(gclk));
	jand g08606(.dina(w_n8866_0[0]),.dinb(n8869),.dout(n8870),.clk(gclk));
	jnot g08607(.din(n8870),.dout(n8871),.clk(gclk));
	jand g08608(.dina(n8871),.dinb(n8868),.dout(n8872),.clk(gclk));
	jand g08609(.dina(w_n8872_0[1]),.dinb(w_n8863_0[1]),.dout(n8873),.clk(gclk));
	jor g08610(.dina(n8873),.dinb(w_n8861_0[1]),.dout(n8874),.clk(gclk));
	jxor g08611(.dina(w_n8419_0[0]),.dinb(w_n199_26[2]),.dout(n8875),.clk(gclk));
	jand g08612(.dina(n8875),.dinb(w_asqrt24_18[1]),.dout(n8876),.clk(gclk));
	jxor g08613(.dina(n8876),.dinb(w_n8429_0[0]),.dout(n8877),.clk(gclk));
	jnot g08614(.din(w_n8431_0[0]),.dout(n8878),.clk(gclk));
	jand g08615(.dina(w_asqrt24_18[0]),.dinb(w_n8438_0[1]),.dout(n8879),.clk(gclk));
	jand g08616(.dina(w_n8879_0[1]),.dinb(w_n8878_0[2]),.dout(n8880),.clk(gclk));
	jor g08617(.dina(n8880),.dinb(w_n8446_0[0]),.dout(n8881),.clk(gclk));
	jor g08618(.dina(n8881),.dinb(w_n8877_0[1]),.dout(n8882),.clk(gclk));
	jnot g08619(.din(n8882),.dout(n8883),.clk(gclk));
	jand g08620(.dina(n8883),.dinb(w_n8874_1[2]),.dout(n8884),.clk(gclk));
	jor g08621(.dina(n8884),.dinb(w_asqrt63_9[2]),.dout(n8885),.clk(gclk));
	jnot g08622(.din(w_n8877_0[0]),.dout(n8886),.clk(gclk));
	jor g08623(.dina(w_n8886_0[2]),.dinb(w_n8874_1[1]),.dout(n8887),.clk(gclk));
	jor g08624(.dina(w_n8879_0[0]),.dinb(w_n8878_0[1]),.dout(n8888),.clk(gclk));
	jand g08625(.dina(w_n8438_0[0]),.dinb(w_n8878_0[0]),.dout(n8889),.clk(gclk));
	jor g08626(.dina(n8889),.dinb(w_n194_25[2]),.dout(n8890),.clk(gclk));
	jnot g08627(.din(n8890),.dout(n8891),.clk(gclk));
	jand g08628(.dina(n8891),.dinb(n8888),.dout(n8892),.clk(gclk));
	jnot g08629(.din(w_asqrt24_17[2]),.dout(n8893),.clk(gclk));
	jnot g08630(.din(w_n8892_0[1]),.dout(n8896),.clk(gclk));
	jand g08631(.dina(n8896),.dinb(w_n8887_0[1]),.dout(n8897),.clk(gclk));
	jand g08632(.dina(n8897),.dinb(w_n8885_0[1]),.dout(n8898),.clk(gclk));
	jxor g08633(.dina(w_n8603_0[0]),.dinb(w_n3376_21[0]),.dout(n8899),.clk(gclk));
	jor g08634(.dina(n8899),.dinb(w_n8898_27[1]),.dout(n8900),.clk(gclk));
	jxor g08635(.dina(n8900),.dinb(w_n8458_0[0]),.dout(n8901),.clk(gclk));
	jor g08636(.dina(w_n8898_27[0]),.dinb(w_n8460_1[0]),.dout(n8902),.clk(gclk));
	jnot g08637(.din(w_a44_0[1]),.dout(n8903),.clk(gclk));
	jnot g08638(.din(a[45]),.dout(n8904),.clk(gclk));
	jand g08639(.dina(w_n8460_0[2]),.dinb(w_n8904_0[2]),.dout(n8905),.clk(gclk));
	jand g08640(.dina(n8905),.dinb(w_n8903_1[1]),.dout(n8906),.clk(gclk));
	jnot g08641(.din(n8906),.dout(n8907),.clk(gclk));
	jand g08642(.dina(n8907),.dinb(n8902),.dout(n8908),.clk(gclk));
	jor g08643(.dina(w_n8908_0[2]),.dinb(w_n8893_15[2]),.dout(n8909),.clk(gclk));
	jor g08644(.dina(w_n8898_26[2]),.dinb(w_a46_0[0]),.dout(n8910),.clk(gclk));
	jxor g08645(.dina(w_n8910_0[1]),.dinb(w_n8461_0[0]),.dout(n8911),.clk(gclk));
	jand g08646(.dina(w_n8908_0[1]),.dinb(w_n8893_15[1]),.dout(n8912),.clk(gclk));
	jor g08647(.dina(n8912),.dinb(w_n8911_0[1]),.dout(n8913),.clk(gclk));
	jand g08648(.dina(w_n8913_0[1]),.dinb(w_n8909_0[1]),.dout(n8914),.clk(gclk));
	jor g08649(.dina(n8914),.dinb(w_n8058_19[1]),.dout(n8915),.clk(gclk));
	jand g08650(.dina(w_n8909_0[0]),.dinb(w_n8058_19[0]),.dout(n8916),.clk(gclk));
	jand g08651(.dina(n8916),.dinb(w_n8913_0[0]),.dout(n8917),.clk(gclk));
	jor g08652(.dina(w_n8910_0[0]),.dinb(w_a47_0[0]),.dout(n8918),.clk(gclk));
	jnot g08653(.din(w_n8885_0[0]),.dout(n8919),.clk(gclk));
	jnot g08654(.din(w_n8887_0[0]),.dout(n8920),.clk(gclk));
	jor g08655(.dina(w_n8892_0[0]),.dinb(w_n8893_15[0]),.dout(n8921),.clk(gclk));
	jor g08656(.dina(n8921),.dinb(w_n8920_0[1]),.dout(n8922),.clk(gclk));
	jor g08657(.dina(n8922),.dinb(n8919),.dout(n8923),.clk(gclk));
	jand g08658(.dina(n8923),.dinb(n8918),.dout(n8924),.clk(gclk));
	jxor g08659(.dina(n8924),.dinb(w_n8063_0[1]),.dout(n8925),.clk(gclk));
	jor g08660(.dina(w_n8925_0[1]),.dinb(w_n8917_0[1]),.dout(n8926),.clk(gclk));
	jand g08661(.dina(n8926),.dinb(w_n8915_0[1]),.dout(n8927),.clk(gclk));
	jor g08662(.dina(w_n8927_0[2]),.dinb(w_n8053_15[1]),.dout(n8928),.clk(gclk));
	jand g08663(.dina(w_n8927_0[1]),.dinb(w_n8053_15[0]),.dout(n8929),.clk(gclk));
	jxor g08664(.dina(w_n8464_0[0]),.dinb(w_n8058_18[2]),.dout(n8930),.clk(gclk));
	jor g08665(.dina(n8930),.dinb(w_n8898_26[1]),.dout(n8931),.clk(gclk));
	jxor g08666(.dina(n8931),.dinb(w_n8467_0[0]),.dout(n8932),.clk(gclk));
	jor g08667(.dina(w_n8932_0[1]),.dinb(n8929),.dout(n8933),.clk(gclk));
	jand g08668(.dina(w_n8933_0[1]),.dinb(w_n8928_0[1]),.dout(n8934),.clk(gclk));
	jor g08669(.dina(n8934),.dinb(w_n7265_19[2]),.dout(n8935),.clk(gclk));
	jnot g08670(.din(w_n8473_0[0]),.dout(n8936),.clk(gclk));
	jor g08671(.dina(n8936),.dinb(w_n8471_0[0]),.dout(n8937),.clk(gclk));
	jor g08672(.dina(n8937),.dinb(w_n8898_26[0]),.dout(n8938),.clk(gclk));
	jxor g08673(.dina(n8938),.dinb(w_n8482_0[0]),.dout(n8939),.clk(gclk));
	jand g08674(.dina(w_n8928_0[0]),.dinb(w_n7265_19[1]),.dout(n8940),.clk(gclk));
	jand g08675(.dina(n8940),.dinb(w_n8933_0[0]),.dout(n8941),.clk(gclk));
	jor g08676(.dina(w_n8941_0[1]),.dinb(w_n8939_0[1]),.dout(n8942),.clk(gclk));
	jand g08677(.dina(w_n8942_0[1]),.dinb(w_n8935_0[1]),.dout(n8943),.clk(gclk));
	jor g08678(.dina(w_n8943_0[2]),.dinb(w_n7260_16[0]),.dout(n8944),.clk(gclk));
	jand g08679(.dina(w_n8943_0[1]),.dinb(w_n7260_15[2]),.dout(n8945),.clk(gclk));
	jxor g08680(.dina(w_n8484_0[0]),.dinb(w_n7265_19[0]),.dout(n8946),.clk(gclk));
	jor g08681(.dina(n8946),.dinb(w_n8898_25[2]),.dout(n8947),.clk(gclk));
	jxor g08682(.dina(n8947),.dinb(w_n8489_0[0]),.dout(n8948),.clk(gclk));
	jnot g08683(.din(w_n8948_0[1]),.dout(n8949),.clk(gclk));
	jor g08684(.dina(n8949),.dinb(n8945),.dout(n8950),.clk(gclk));
	jand g08685(.dina(w_n8950_0[1]),.dinb(w_n8944_0[1]),.dout(n8951),.clk(gclk));
	jor g08686(.dina(n8951),.dinb(w_n6505_19[1]),.dout(n8952),.clk(gclk));
	jand g08687(.dina(w_n8944_0[0]),.dinb(w_n6505_19[0]),.dout(n8953),.clk(gclk));
	jand g08688(.dina(n8953),.dinb(w_n8950_0[0]),.dout(n8954),.clk(gclk));
	jnot g08689(.din(w_n8493_0[0]),.dout(n8955),.clk(gclk));
	jnot g08690(.din(w_n8898_25[1]),.dout(asqrt_fa_24),.clk(gclk));
	jand g08691(.dina(w_asqrt23_19),.dinb(n8955),.dout(n8957),.clk(gclk));
	jand g08692(.dina(w_n8957_0[1]),.dinb(w_n8500_0[0]),.dout(n8958),.clk(gclk));
	jor g08693(.dina(n8958),.dinb(w_n8498_0[0]),.dout(n8959),.clk(gclk));
	jand g08694(.dina(w_n8957_0[0]),.dinb(w_n8501_0[0]),.dout(n8960),.clk(gclk));
	jnot g08695(.din(n8960),.dout(n8961),.clk(gclk));
	jand g08696(.dina(n8961),.dinb(n8959),.dout(n8962),.clk(gclk));
	jnot g08697(.din(n8962),.dout(n8963),.clk(gclk));
	jor g08698(.dina(w_n8963_0[1]),.dinb(w_n8954_0[1]),.dout(n8964),.clk(gclk));
	jand g08699(.dina(n8964),.dinb(w_n8952_0[1]),.dout(n8965),.clk(gclk));
	jor g08700(.dina(w_n8965_0[2]),.dinb(w_n6500_16[0]),.dout(n8966),.clk(gclk));
	jand g08701(.dina(w_n8965_0[1]),.dinb(w_n6500_15[2]),.dout(n8967),.clk(gclk));
	jnot g08702(.din(w_n8508_0[0]),.dout(n8968),.clk(gclk));
	jxor g08703(.dina(w_n8502_0[0]),.dinb(w_n6505_18[2]),.dout(n8969),.clk(gclk));
	jor g08704(.dina(n8969),.dinb(w_n8898_25[0]),.dout(n8970),.clk(gclk));
	jxor g08705(.dina(n8970),.dinb(n8968),.dout(n8971),.clk(gclk));
	jnot g08706(.din(w_n8971_0[1]),.dout(n8972),.clk(gclk));
	jor g08707(.dina(n8972),.dinb(n8967),.dout(n8973),.clk(gclk));
	jand g08708(.dina(w_n8973_0[1]),.dinb(w_n8966_0[1]),.dout(n8974),.clk(gclk));
	jor g08709(.dina(n8974),.dinb(w_n5793_19[2]),.dout(n8975),.clk(gclk));
	jnot g08710(.din(w_n8513_0[0]),.dout(n8976),.clk(gclk));
	jor g08711(.dina(n8976),.dinb(w_n8511_0[0]),.dout(n8977),.clk(gclk));
	jor g08712(.dina(n8977),.dinb(w_n8898_24[2]),.dout(n8978),.clk(gclk));
	jxor g08713(.dina(n8978),.dinb(w_n8522_0[0]),.dout(n8979),.clk(gclk));
	jand g08714(.dina(w_n8966_0[0]),.dinb(w_n5793_19[1]),.dout(n8980),.clk(gclk));
	jand g08715(.dina(n8980),.dinb(w_n8973_0[0]),.dout(n8981),.clk(gclk));
	jor g08716(.dina(w_n8981_0[1]),.dinb(w_n8979_0[1]),.dout(n8982),.clk(gclk));
	jand g08717(.dina(w_n8982_0[1]),.dinb(w_n8975_0[1]),.dout(n8983),.clk(gclk));
	jor g08718(.dina(w_n8983_0[2]),.dinb(w_n5788_16[1]),.dout(n8984),.clk(gclk));
	jand g08719(.dina(w_n8983_0[1]),.dinb(w_n5788_16[0]),.dout(n8985),.clk(gclk));
	jnot g08720(.din(w_n8529_0[0]),.dout(n8986),.clk(gclk));
	jxor g08721(.dina(w_n8524_0[0]),.dinb(w_n5793_19[0]),.dout(n8987),.clk(gclk));
	jor g08722(.dina(n8987),.dinb(w_n8898_24[1]),.dout(n8988),.clk(gclk));
	jxor g08723(.dina(n8988),.dinb(n8986),.dout(n8989),.clk(gclk));
	jnot g08724(.din(n8989),.dout(n8990),.clk(gclk));
	jor g08725(.dina(w_n8990_0[1]),.dinb(n8985),.dout(n8991),.clk(gclk));
	jand g08726(.dina(w_n8991_0[1]),.dinb(w_n8984_0[1]),.dout(n8992),.clk(gclk));
	jor g08727(.dina(n8992),.dinb(w_n5121_19[1]),.dout(n8993),.clk(gclk));
	jand g08728(.dina(w_n8984_0[0]),.dinb(w_n5121_19[0]),.dout(n8994),.clk(gclk));
	jand g08729(.dina(n8994),.dinb(w_n8991_0[0]),.dout(n8995),.clk(gclk));
	jnot g08730(.din(w_n8532_0[0]),.dout(n8996),.clk(gclk));
	jand g08731(.dina(w_asqrt23_18[2]),.dinb(n8996),.dout(n8997),.clk(gclk));
	jand g08732(.dina(w_n8997_0[1]),.dinb(w_n8539_0[0]),.dout(n8998),.clk(gclk));
	jor g08733(.dina(n8998),.dinb(w_n8537_0[0]),.dout(n8999),.clk(gclk));
	jand g08734(.dina(w_n8997_0[0]),.dinb(w_n8540_0[0]),.dout(n9000),.clk(gclk));
	jnot g08735(.din(n9000),.dout(n9001),.clk(gclk));
	jand g08736(.dina(n9001),.dinb(n8999),.dout(n9002),.clk(gclk));
	jnot g08737(.din(n9002),.dout(n9003),.clk(gclk));
	jor g08738(.dina(w_n9003_0[1]),.dinb(w_n8995_0[1]),.dout(n9004),.clk(gclk));
	jand g08739(.dina(n9004),.dinb(w_n8993_0[1]),.dout(n9005),.clk(gclk));
	jor g08740(.dina(w_n9005_0[1]),.dinb(w_n5116_16[1]),.dout(n9006),.clk(gclk));
	jxor g08741(.dina(w_n8541_0[0]),.dinb(w_n5121_18[2]),.dout(n9007),.clk(gclk));
	jor g08742(.dina(n9007),.dinb(w_n8898_24[0]),.dout(n9008),.clk(gclk));
	jxor g08743(.dina(n9008),.dinb(w_n8546_0[0]),.dout(n9009),.clk(gclk));
	jand g08744(.dina(w_n9005_0[0]),.dinb(w_n5116_16[0]),.dout(n9010),.clk(gclk));
	jor g08745(.dina(w_n9010_0[1]),.dinb(w_n9009_0[1]),.dout(n9011),.clk(gclk));
	jand g08746(.dina(w_n9011_0[2]),.dinb(w_n9006_0[2]),.dout(n9012),.clk(gclk));
	jor g08747(.dina(n9012),.dinb(w_n4499_20[0]),.dout(n9013),.clk(gclk));
	jnot g08748(.din(w_n8551_0[0]),.dout(n9014),.clk(gclk));
	jor g08749(.dina(n9014),.dinb(w_n8549_0[0]),.dout(n9015),.clk(gclk));
	jor g08750(.dina(n9015),.dinb(w_n8898_23[2]),.dout(n9016),.clk(gclk));
	jxor g08751(.dina(n9016),.dinb(w_n8560_0[0]),.dout(n9017),.clk(gclk));
	jand g08752(.dina(w_n9006_0[1]),.dinb(w_n4499_19[2]),.dout(n9018),.clk(gclk));
	jand g08753(.dina(n9018),.dinb(w_n9011_0[1]),.dout(n9019),.clk(gclk));
	jor g08754(.dina(w_n9019_0[1]),.dinb(w_n9017_0[1]),.dout(n9020),.clk(gclk));
	jand g08755(.dina(w_n9020_0[1]),.dinb(w_n9013_0[1]),.dout(n9021),.clk(gclk));
	jor g08756(.dina(w_n9021_0[2]),.dinb(w_n4494_17[1]),.dout(n9022),.clk(gclk));
	jand g08757(.dina(w_n9021_0[1]),.dinb(w_n4494_17[0]),.dout(n9023),.clk(gclk));
	jnot g08758(.din(w_n8563_0[0]),.dout(n9024),.clk(gclk));
	jand g08759(.dina(w_asqrt23_18[1]),.dinb(n9024),.dout(n9025),.clk(gclk));
	jand g08760(.dina(w_n9025_0[1]),.dinb(w_n8568_0[0]),.dout(n9026),.clk(gclk));
	jor g08761(.dina(n9026),.dinb(w_n8567_0[0]),.dout(n9027),.clk(gclk));
	jand g08762(.dina(w_n9025_0[0]),.dinb(w_n8569_0[0]),.dout(n9028),.clk(gclk));
	jnot g08763(.din(n9028),.dout(n9029),.clk(gclk));
	jand g08764(.dina(n9029),.dinb(n9027),.dout(n9030),.clk(gclk));
	jnot g08765(.din(n9030),.dout(n9031),.clk(gclk));
	jor g08766(.dina(w_n9031_0[1]),.dinb(n9023),.dout(n9032),.clk(gclk));
	jand g08767(.dina(w_n9032_0[1]),.dinb(w_n9022_0[1]),.dout(n9033),.clk(gclk));
	jor g08768(.dina(n9033),.dinb(w_n3912_20[0]),.dout(n9034),.clk(gclk));
	jand g08769(.dina(w_n9022_0[0]),.dinb(w_n3912_19[2]),.dout(n9035),.clk(gclk));
	jand g08770(.dina(n9035),.dinb(w_n9032_0[0]),.dout(n9036),.clk(gclk));
	jnot g08771(.din(w_n8571_0[0]),.dout(n9037),.clk(gclk));
	jand g08772(.dina(w_asqrt23_18[0]),.dinb(n9037),.dout(n9038),.clk(gclk));
	jand g08773(.dina(w_n9038_0[1]),.dinb(w_n8578_0[0]),.dout(n9039),.clk(gclk));
	jor g08774(.dina(n9039),.dinb(w_n8576_0[0]),.dout(n9040),.clk(gclk));
	jand g08775(.dina(w_n9038_0[0]),.dinb(w_n8579_0[0]),.dout(n9041),.clk(gclk));
	jnot g08776(.din(n9041),.dout(n9042),.clk(gclk));
	jand g08777(.dina(n9042),.dinb(n9040),.dout(n9043),.clk(gclk));
	jnot g08778(.din(n9043),.dout(n9044),.clk(gclk));
	jor g08779(.dina(w_n9044_0[1]),.dinb(w_n9036_0[1]),.dout(n9045),.clk(gclk));
	jand g08780(.dina(n9045),.dinb(w_n9034_0[1]),.dout(n9046),.clk(gclk));
	jor g08781(.dina(w_n9046_0[1]),.dinb(w_n3907_17[1]),.dout(n9047),.clk(gclk));
	jxor g08782(.dina(w_n8580_0[0]),.dinb(w_n3912_19[1]),.dout(n9048),.clk(gclk));
	jor g08783(.dina(n9048),.dinb(w_n8898_23[1]),.dout(n9049),.clk(gclk));
	jxor g08784(.dina(n9049),.dinb(w_n8591_0[0]),.dout(n9050),.clk(gclk));
	jand g08785(.dina(w_n9046_0[0]),.dinb(w_n3907_17[0]),.dout(n9051),.clk(gclk));
	jor g08786(.dina(w_n9051_0[1]),.dinb(w_n9050_0[1]),.dout(n9052),.clk(gclk));
	jand g08787(.dina(w_n9052_0[2]),.dinb(w_n9047_0[2]),.dout(n9053),.clk(gclk));
	jor g08788(.dina(n9053),.dinb(w_n3376_20[2]),.dout(n9054),.clk(gclk));
	jand g08789(.dina(w_n9047_0[1]),.dinb(w_n3376_20[1]),.dout(n9055),.clk(gclk));
	jand g08790(.dina(n9055),.dinb(w_n9052_0[1]),.dout(n9056),.clk(gclk));
	jnot g08791(.din(w_n8594_0[0]),.dout(n9057),.clk(gclk));
	jand g08792(.dina(w_asqrt23_17[2]),.dinb(n9057),.dout(n9058),.clk(gclk));
	jand g08793(.dina(w_n9058_0[1]),.dinb(w_n8601_0[0]),.dout(n9059),.clk(gclk));
	jor g08794(.dina(n9059),.dinb(w_n8599_0[0]),.dout(n9060),.clk(gclk));
	jand g08795(.dina(w_n9058_0[0]),.dinb(w_n8602_0[0]),.dout(n9061),.clk(gclk));
	jnot g08796(.din(n9061),.dout(n9062),.clk(gclk));
	jand g08797(.dina(n9062),.dinb(n9060),.dout(n9063),.clk(gclk));
	jnot g08798(.din(n9063),.dout(n9064),.clk(gclk));
	jor g08799(.dina(w_n9064_0[1]),.dinb(w_n9056_0[1]),.dout(n9065),.clk(gclk));
	jand g08800(.dina(n9065),.dinb(w_n9054_0[1]),.dout(n9066),.clk(gclk));
	jor g08801(.dina(w_n9066_0[2]),.dinb(w_n3371_18[0]),.dout(n9067),.clk(gclk));
	jnot g08802(.din(w_n8901_0[1]),.dout(n9068),.clk(gclk));
	jand g08803(.dina(w_n9066_0[1]),.dinb(w_n3371_17[2]),.dout(n9069),.clk(gclk));
	jor g08804(.dina(n9069),.dinb(n9068),.dout(n9070),.clk(gclk));
	jand g08805(.dina(w_n9070_0[1]),.dinb(w_n9067_0[1]),.dout(n9071),.clk(gclk));
	jor g08806(.dina(n9071),.dinb(w_n2875_21[0]),.dout(n9072),.clk(gclk));
	jnot g08807(.din(w_n8611_0[0]),.dout(n9073),.clk(gclk));
	jor g08808(.dina(n9073),.dinb(w_n8609_0[0]),.dout(n9074),.clk(gclk));
	jor g08809(.dina(n9074),.dinb(w_n8898_23[0]),.dout(n9075),.clk(gclk));
	jxor g08810(.dina(n9075),.dinb(w_n8620_0[0]),.dout(n9076),.clk(gclk));
	jand g08811(.dina(w_n9067_0[0]),.dinb(w_n2875_20[2]),.dout(n9077),.clk(gclk));
	jand g08812(.dina(n9077),.dinb(w_n9070_0[0]),.dout(n9078),.clk(gclk));
	jor g08813(.dina(w_n9078_0[1]),.dinb(w_n9076_0[1]),.dout(n9079),.clk(gclk));
	jand g08814(.dina(w_n9079_0[1]),.dinb(w_n9072_0[1]),.dout(n9080),.clk(gclk));
	jor g08815(.dina(w_n9080_0[1]),.dinb(w_n2870_18[0]),.dout(n9081),.clk(gclk));
	jxor g08816(.dina(w_n8622_0[0]),.dinb(w_n2875_20[1]),.dout(n9082),.clk(gclk));
	jor g08817(.dina(n9082),.dinb(w_n8898_22[2]),.dout(n9083),.clk(gclk));
	jxor g08818(.dina(n9083),.dinb(w_n8633_0[0]),.dout(n9084),.clk(gclk));
	jand g08819(.dina(w_n9080_0[0]),.dinb(w_n2870_17[2]),.dout(n9085),.clk(gclk));
	jor g08820(.dina(w_n9085_0[1]),.dinb(w_n9084_0[1]),.dout(n9086),.clk(gclk));
	jand g08821(.dina(w_n9086_0[2]),.dinb(w_n9081_0[2]),.dout(n9087),.clk(gclk));
	jor g08822(.dina(n9087),.dinb(w_n2425_21[1]),.dout(n9088),.clk(gclk));
	jnot g08823(.din(w_n8638_0[0]),.dout(n9089),.clk(gclk));
	jor g08824(.dina(n9089),.dinb(w_n8636_0[0]),.dout(n9090),.clk(gclk));
	jor g08825(.dina(n9090),.dinb(w_n8898_22[1]),.dout(n9091),.clk(gclk));
	jxor g08826(.dina(n9091),.dinb(w_n8647_0[0]),.dout(n9092),.clk(gclk));
	jand g08827(.dina(w_n9081_0[1]),.dinb(w_n2425_21[0]),.dout(n9093),.clk(gclk));
	jand g08828(.dina(n9093),.dinb(w_n9086_0[1]),.dout(n9094),.clk(gclk));
	jor g08829(.dina(w_n9094_0[1]),.dinb(w_n9092_0[1]),.dout(n9095),.clk(gclk));
	jand g08830(.dina(w_n9095_0[1]),.dinb(w_n9088_0[1]),.dout(n9096),.clk(gclk));
	jor g08831(.dina(w_n9096_0[2]),.dinb(w_n2420_19[0]),.dout(n9097),.clk(gclk));
	jand g08832(.dina(w_n9096_0[1]),.dinb(w_n2420_18[2]),.dout(n9098),.clk(gclk));
	jnot g08833(.din(w_n8650_0[0]),.dout(n9099),.clk(gclk));
	jand g08834(.dina(w_asqrt23_17[1]),.dinb(n9099),.dout(n9100),.clk(gclk));
	jand g08835(.dina(w_n9100_0[1]),.dinb(w_n8655_0[0]),.dout(n9101),.clk(gclk));
	jor g08836(.dina(n9101),.dinb(w_n8654_0[0]),.dout(n9102),.clk(gclk));
	jand g08837(.dina(w_n9100_0[0]),.dinb(w_n8656_0[0]),.dout(n9103),.clk(gclk));
	jnot g08838(.din(n9103),.dout(n9104),.clk(gclk));
	jand g08839(.dina(n9104),.dinb(n9102),.dout(n9105),.clk(gclk));
	jnot g08840(.din(n9105),.dout(n9106),.clk(gclk));
	jor g08841(.dina(w_n9106_0[1]),.dinb(n9098),.dout(n9107),.clk(gclk));
	jand g08842(.dina(w_n9107_0[1]),.dinb(w_n9097_0[1]),.dout(n9108),.clk(gclk));
	jor g08843(.dina(n9108),.dinb(w_n2010_21[1]),.dout(n9109),.clk(gclk));
	jand g08844(.dina(w_n9097_0[0]),.dinb(w_n2010_21[0]),.dout(n9110),.clk(gclk));
	jand g08845(.dina(n9110),.dinb(w_n9107_0[0]),.dout(n9111),.clk(gclk));
	jnot g08846(.din(w_n8658_0[0]),.dout(n9112),.clk(gclk));
	jand g08847(.dina(w_asqrt23_17[0]),.dinb(n9112),.dout(n9113),.clk(gclk));
	jand g08848(.dina(w_n9113_0[1]),.dinb(w_n8665_0[0]),.dout(n9114),.clk(gclk));
	jor g08849(.dina(n9114),.dinb(w_n8663_0[0]),.dout(n9115),.clk(gclk));
	jand g08850(.dina(w_n9113_0[0]),.dinb(w_n8666_0[0]),.dout(n9116),.clk(gclk));
	jnot g08851(.din(n9116),.dout(n9117),.clk(gclk));
	jand g08852(.dina(n9117),.dinb(n9115),.dout(n9118),.clk(gclk));
	jnot g08853(.din(n9118),.dout(n9119),.clk(gclk));
	jor g08854(.dina(w_n9119_0[1]),.dinb(w_n9111_0[1]),.dout(n9120),.clk(gclk));
	jand g08855(.dina(n9120),.dinb(w_n9109_0[1]),.dout(n9121),.clk(gclk));
	jor g08856(.dina(w_n9121_0[1]),.dinb(w_n2005_19[0]),.dout(n9122),.clk(gclk));
	jxor g08857(.dina(w_n8667_0[0]),.dinb(w_n2010_20[2]),.dout(n9123),.clk(gclk));
	jor g08858(.dina(n9123),.dinb(w_n8898_22[0]),.dout(n9124),.clk(gclk));
	jxor g08859(.dina(n9124),.dinb(w_n8678_0[0]),.dout(n9125),.clk(gclk));
	jand g08860(.dina(w_n9121_0[0]),.dinb(w_n2005_18[2]),.dout(n9126),.clk(gclk));
	jor g08861(.dina(w_n9126_0[1]),.dinb(w_n9125_0[1]),.dout(n9127),.clk(gclk));
	jand g08862(.dina(w_n9127_0[2]),.dinb(w_n9122_0[2]),.dout(n9128),.clk(gclk));
	jor g08863(.dina(n9128),.dinb(w_n1646_22[0]),.dout(n9129),.clk(gclk));
	jnot g08864(.din(w_n8683_0[0]),.dout(n9130),.clk(gclk));
	jor g08865(.dina(n9130),.dinb(w_n8681_0[0]),.dout(n9131),.clk(gclk));
	jor g08866(.dina(n9131),.dinb(w_n8898_21[2]),.dout(n9132),.clk(gclk));
	jxor g08867(.dina(n9132),.dinb(w_n8692_0[0]),.dout(n9133),.clk(gclk));
	jand g08868(.dina(w_n9122_0[1]),.dinb(w_n1646_21[2]),.dout(n9134),.clk(gclk));
	jand g08869(.dina(n9134),.dinb(w_n9127_0[1]),.dout(n9135),.clk(gclk));
	jor g08870(.dina(w_n9135_0[1]),.dinb(w_n9133_0[1]),.dout(n9136),.clk(gclk));
	jand g08871(.dina(w_n9136_0[1]),.dinb(w_n9129_0[1]),.dout(n9137),.clk(gclk));
	jor g08872(.dina(w_n9137_0[2]),.dinb(w_n1641_19[2]),.dout(n9138),.clk(gclk));
	jand g08873(.dina(w_n9137_0[1]),.dinb(w_n1641_19[1]),.dout(n9139),.clk(gclk));
	jnot g08874(.din(w_n8695_0[0]),.dout(n9140),.clk(gclk));
	jand g08875(.dina(w_asqrt23_16[2]),.dinb(n9140),.dout(n9141),.clk(gclk));
	jand g08876(.dina(w_n9141_0[1]),.dinb(w_n8700_0[0]),.dout(n9142),.clk(gclk));
	jor g08877(.dina(n9142),.dinb(w_n8699_0[0]),.dout(n9143),.clk(gclk));
	jand g08878(.dina(w_n9141_0[0]),.dinb(w_n8701_0[0]),.dout(n9144),.clk(gclk));
	jnot g08879(.din(n9144),.dout(n9145),.clk(gclk));
	jand g08880(.dina(n9145),.dinb(n9143),.dout(n9146),.clk(gclk));
	jnot g08881(.din(n9146),.dout(n9147),.clk(gclk));
	jor g08882(.dina(w_n9147_0[1]),.dinb(n9139),.dout(n9148),.clk(gclk));
	jand g08883(.dina(w_n9148_0[1]),.dinb(w_n9138_0[1]),.dout(n9149),.clk(gclk));
	jor g08884(.dina(n9149),.dinb(w_n1317_22[0]),.dout(n9150),.clk(gclk));
	jand g08885(.dina(w_n9138_0[0]),.dinb(w_n1317_21[2]),.dout(n9151),.clk(gclk));
	jand g08886(.dina(n9151),.dinb(w_n9148_0[0]),.dout(n9152),.clk(gclk));
	jnot g08887(.din(w_n8703_0[0]),.dout(n9153),.clk(gclk));
	jand g08888(.dina(w_asqrt23_16[1]),.dinb(n9153),.dout(n9154),.clk(gclk));
	jand g08889(.dina(w_n9154_0[1]),.dinb(w_n8710_0[0]),.dout(n9155),.clk(gclk));
	jor g08890(.dina(n9155),.dinb(w_n8708_0[0]),.dout(n9156),.clk(gclk));
	jand g08891(.dina(w_n9154_0[0]),.dinb(w_n8711_0[0]),.dout(n9157),.clk(gclk));
	jnot g08892(.din(n9157),.dout(n9158),.clk(gclk));
	jand g08893(.dina(n9158),.dinb(n9156),.dout(n9159),.clk(gclk));
	jnot g08894(.din(n9159),.dout(n9160),.clk(gclk));
	jor g08895(.dina(w_n9160_0[1]),.dinb(w_n9152_0[1]),.dout(n9161),.clk(gclk));
	jand g08896(.dina(n9161),.dinb(w_n9150_0[1]),.dout(n9162),.clk(gclk));
	jor g08897(.dina(w_n9162_0[1]),.dinb(w_n1312_19[2]),.dout(n9163),.clk(gclk));
	jxor g08898(.dina(w_n8712_0[0]),.dinb(w_n1317_21[1]),.dout(n9164),.clk(gclk));
	jor g08899(.dina(n9164),.dinb(w_n8898_21[1]),.dout(n9165),.clk(gclk));
	jxor g08900(.dina(n9165),.dinb(w_n8723_0[0]),.dout(n9166),.clk(gclk));
	jand g08901(.dina(w_n9162_0[0]),.dinb(w_n1312_19[1]),.dout(n9167),.clk(gclk));
	jor g08902(.dina(w_n9167_0[1]),.dinb(w_n9166_0[1]),.dout(n9168),.clk(gclk));
	jand g08903(.dina(w_n9168_0[2]),.dinb(w_n9163_0[2]),.dout(n9169),.clk(gclk));
	jor g08904(.dina(n9169),.dinb(w_n1039_22[1]),.dout(n9170),.clk(gclk));
	jnot g08905(.din(w_n8728_0[0]),.dout(n9171),.clk(gclk));
	jor g08906(.dina(n9171),.dinb(w_n8726_0[0]),.dout(n9172),.clk(gclk));
	jor g08907(.dina(n9172),.dinb(w_n8898_21[0]),.dout(n9173),.clk(gclk));
	jxor g08908(.dina(n9173),.dinb(w_n8737_0[0]),.dout(n9174),.clk(gclk));
	jand g08909(.dina(w_n9163_0[1]),.dinb(w_n1039_22[0]),.dout(n9175),.clk(gclk));
	jand g08910(.dina(n9175),.dinb(w_n9168_0[1]),.dout(n9176),.clk(gclk));
	jor g08911(.dina(w_n9176_0[1]),.dinb(w_n9174_0[1]),.dout(n9177),.clk(gclk));
	jand g08912(.dina(w_n9177_0[1]),.dinb(w_n9170_0[1]),.dout(n9178),.clk(gclk));
	jor g08913(.dina(w_n9178_0[2]),.dinb(w_n1034_20[2]),.dout(n9179),.clk(gclk));
	jand g08914(.dina(w_n9178_0[1]),.dinb(w_n1034_20[1]),.dout(n9180),.clk(gclk));
	jnot g08915(.din(w_n8740_0[0]),.dout(n9181),.clk(gclk));
	jand g08916(.dina(w_asqrt23_16[0]),.dinb(n9181),.dout(n9182),.clk(gclk));
	jand g08917(.dina(w_n9182_0[1]),.dinb(w_n8745_0[0]),.dout(n9183),.clk(gclk));
	jor g08918(.dina(n9183),.dinb(w_n8744_0[0]),.dout(n9184),.clk(gclk));
	jand g08919(.dina(w_n9182_0[0]),.dinb(w_n8746_0[0]),.dout(n9185),.clk(gclk));
	jnot g08920(.din(n9185),.dout(n9186),.clk(gclk));
	jand g08921(.dina(n9186),.dinb(n9184),.dout(n9187),.clk(gclk));
	jnot g08922(.din(n9187),.dout(n9188),.clk(gclk));
	jor g08923(.dina(w_n9188_0[1]),.dinb(n9180),.dout(n9189),.clk(gclk));
	jand g08924(.dina(w_n9189_0[1]),.dinb(w_n9179_0[1]),.dout(n9190),.clk(gclk));
	jor g08925(.dina(n9190),.dinb(w_n796_22[1]),.dout(n9191),.clk(gclk));
	jand g08926(.dina(w_n9179_0[0]),.dinb(w_n796_22[0]),.dout(n9192),.clk(gclk));
	jand g08927(.dina(n9192),.dinb(w_n9189_0[0]),.dout(n9193),.clk(gclk));
	jnot g08928(.din(w_n8748_0[0]),.dout(n9194),.clk(gclk));
	jand g08929(.dina(w_asqrt23_15[2]),.dinb(n9194),.dout(n9195),.clk(gclk));
	jand g08930(.dina(w_n9195_0[1]),.dinb(w_n8755_0[0]),.dout(n9196),.clk(gclk));
	jor g08931(.dina(n9196),.dinb(w_n8753_0[0]),.dout(n9197),.clk(gclk));
	jand g08932(.dina(w_n9195_0[0]),.dinb(w_n8756_0[0]),.dout(n9198),.clk(gclk));
	jnot g08933(.din(n9198),.dout(n9199),.clk(gclk));
	jand g08934(.dina(n9199),.dinb(n9197),.dout(n9200),.clk(gclk));
	jnot g08935(.din(n9200),.dout(n9201),.clk(gclk));
	jor g08936(.dina(w_n9201_0[1]),.dinb(w_n9193_0[1]),.dout(n9202),.clk(gclk));
	jand g08937(.dina(n9202),.dinb(w_n9191_0[1]),.dout(n9203),.clk(gclk));
	jor g08938(.dina(w_n9203_0[1]),.dinb(w_n791_20[2]),.dout(n9204),.clk(gclk));
	jxor g08939(.dina(w_n8757_0[0]),.dinb(w_n796_21[2]),.dout(n9205),.clk(gclk));
	jor g08940(.dina(n9205),.dinb(w_n8898_20[2]),.dout(n9206),.clk(gclk));
	jxor g08941(.dina(n9206),.dinb(w_n8768_0[0]),.dout(n9207),.clk(gclk));
	jand g08942(.dina(w_n9203_0[0]),.dinb(w_n791_20[1]),.dout(n9208),.clk(gclk));
	jor g08943(.dina(w_n9208_0[1]),.dinb(w_n9207_0[1]),.dout(n9209),.clk(gclk));
	jand g08944(.dina(w_n9209_0[2]),.dinb(w_n9204_0[2]),.dout(n9210),.clk(gclk));
	jor g08945(.dina(n9210),.dinb(w_n595_22[2]),.dout(n9211),.clk(gclk));
	jnot g08946(.din(w_n8773_0[0]),.dout(n9212),.clk(gclk));
	jor g08947(.dina(n9212),.dinb(w_n8771_0[0]),.dout(n9213),.clk(gclk));
	jor g08948(.dina(n9213),.dinb(w_n8898_20[1]),.dout(n9214),.clk(gclk));
	jxor g08949(.dina(n9214),.dinb(w_n8782_0[0]),.dout(n9215),.clk(gclk));
	jand g08950(.dina(w_n9204_0[1]),.dinb(w_n595_22[1]),.dout(n9216),.clk(gclk));
	jand g08951(.dina(n9216),.dinb(w_n9209_0[1]),.dout(n9217),.clk(gclk));
	jor g08952(.dina(w_n9217_0[1]),.dinb(w_n9215_0[1]),.dout(n9218),.clk(gclk));
	jand g08953(.dina(w_n9218_0[1]),.dinb(w_n9211_0[1]),.dout(n9219),.clk(gclk));
	jor g08954(.dina(w_n9219_0[2]),.dinb(w_n590_21[1]),.dout(n9220),.clk(gclk));
	jand g08955(.dina(w_n9219_0[1]),.dinb(w_n590_21[0]),.dout(n9221),.clk(gclk));
	jnot g08956(.din(w_n8785_0[0]),.dout(n9222),.clk(gclk));
	jand g08957(.dina(w_asqrt23_15[1]),.dinb(n9222),.dout(n9223),.clk(gclk));
	jand g08958(.dina(w_n9223_0[1]),.dinb(w_n8790_0[0]),.dout(n9224),.clk(gclk));
	jor g08959(.dina(n9224),.dinb(w_n8789_0[0]),.dout(n9225),.clk(gclk));
	jand g08960(.dina(w_n9223_0[0]),.dinb(w_n8791_0[0]),.dout(n9226),.clk(gclk));
	jnot g08961(.din(n9226),.dout(n9227),.clk(gclk));
	jand g08962(.dina(n9227),.dinb(n9225),.dout(n9228),.clk(gclk));
	jnot g08963(.din(n9228),.dout(n9229),.clk(gclk));
	jor g08964(.dina(w_n9229_0[1]),.dinb(n9221),.dout(n9230),.clk(gclk));
	jand g08965(.dina(w_n9230_0[1]),.dinb(w_n9220_0[1]),.dout(n9231),.clk(gclk));
	jor g08966(.dina(n9231),.dinb(w_n430_22[2]),.dout(n9232),.clk(gclk));
	jand g08967(.dina(w_n9220_0[0]),.dinb(w_n430_22[1]),.dout(n9233),.clk(gclk));
	jand g08968(.dina(n9233),.dinb(w_n9230_0[0]),.dout(n9234),.clk(gclk));
	jnot g08969(.din(w_n8793_0[0]),.dout(n9235),.clk(gclk));
	jand g08970(.dina(w_asqrt23_15[0]),.dinb(n9235),.dout(n9236),.clk(gclk));
	jand g08971(.dina(w_n9236_0[1]),.dinb(w_n8800_0[0]),.dout(n9237),.clk(gclk));
	jor g08972(.dina(n9237),.dinb(w_n8798_0[0]),.dout(n9238),.clk(gclk));
	jand g08973(.dina(w_n9236_0[0]),.dinb(w_n8801_0[0]),.dout(n9239),.clk(gclk));
	jnot g08974(.din(n9239),.dout(n9240),.clk(gclk));
	jand g08975(.dina(n9240),.dinb(n9238),.dout(n9241),.clk(gclk));
	jnot g08976(.din(n9241),.dout(n9242),.clk(gclk));
	jor g08977(.dina(w_n9242_0[1]),.dinb(w_n9234_0[1]),.dout(n9243),.clk(gclk));
	jand g08978(.dina(n9243),.dinb(w_n9232_0[1]),.dout(n9244),.clk(gclk));
	jor g08979(.dina(w_n9244_0[1]),.dinb(w_n425_21[1]),.dout(n9245),.clk(gclk));
	jxor g08980(.dina(w_n8802_0[0]),.dinb(w_n430_22[0]),.dout(n9246),.clk(gclk));
	jor g08981(.dina(n9246),.dinb(w_n8898_20[0]),.dout(n9247),.clk(gclk));
	jxor g08982(.dina(n9247),.dinb(w_n8813_0[0]),.dout(n9248),.clk(gclk));
	jand g08983(.dina(w_n9244_0[0]),.dinb(w_n425_21[0]),.dout(n9249),.clk(gclk));
	jor g08984(.dina(w_n9249_0[1]),.dinb(w_n9248_0[1]),.dout(n9250),.clk(gclk));
	jand g08985(.dina(w_n9250_0[2]),.dinb(w_n9245_0[2]),.dout(n9251),.clk(gclk));
	jor g08986(.dina(n9251),.dinb(w_n305_23[0]),.dout(n9252),.clk(gclk));
	jnot g08987(.din(w_n8818_0[0]),.dout(n9253),.clk(gclk));
	jor g08988(.dina(n9253),.dinb(w_n8816_0[0]),.dout(n9254),.clk(gclk));
	jor g08989(.dina(n9254),.dinb(w_n8898_19[2]),.dout(n9255),.clk(gclk));
	jxor g08990(.dina(n9255),.dinb(w_n8827_0[0]),.dout(n9256),.clk(gclk));
	jand g08991(.dina(w_n9245_0[1]),.dinb(w_n305_22[2]),.dout(n9257),.clk(gclk));
	jand g08992(.dina(n9257),.dinb(w_n9250_0[1]),.dout(n9258),.clk(gclk));
	jor g08993(.dina(w_n9258_0[1]),.dinb(w_n9256_0[1]),.dout(n9259),.clk(gclk));
	jand g08994(.dina(w_n9259_0[1]),.dinb(w_n9252_0[1]),.dout(n9260),.clk(gclk));
	jor g08995(.dina(w_n9260_0[2]),.dinb(w_n290_22[2]),.dout(n9261),.clk(gclk));
	jand g08996(.dina(w_n9260_0[1]),.dinb(w_n290_22[1]),.dout(n9262),.clk(gclk));
	jnot g08997(.din(w_n8830_0[0]),.dout(n9263),.clk(gclk));
	jand g08998(.dina(w_asqrt23_14[2]),.dinb(n9263),.dout(n9264),.clk(gclk));
	jand g08999(.dina(w_n9264_0[1]),.dinb(w_n8835_0[0]),.dout(n9265),.clk(gclk));
	jor g09000(.dina(n9265),.dinb(w_n8834_0[0]),.dout(n9266),.clk(gclk));
	jand g09001(.dina(w_n9264_0[0]),.dinb(w_n8836_0[0]),.dout(n9267),.clk(gclk));
	jnot g09002(.din(n9267),.dout(n9268),.clk(gclk));
	jand g09003(.dina(n9268),.dinb(n9266),.dout(n9269),.clk(gclk));
	jnot g09004(.din(n9269),.dout(n9270),.clk(gclk));
	jor g09005(.dina(w_n9270_0[1]),.dinb(n9262),.dout(n9271),.clk(gclk));
	jand g09006(.dina(w_n9271_0[1]),.dinb(w_n9261_0[1]),.dout(n9272),.clk(gclk));
	jor g09007(.dina(n9272),.dinb(w_n223_23[0]),.dout(n9273),.clk(gclk));
	jand g09008(.dina(w_n9261_0[0]),.dinb(w_n223_22[2]),.dout(n9274),.clk(gclk));
	jand g09009(.dina(n9274),.dinb(w_n9271_0[0]),.dout(n9275),.clk(gclk));
	jnot g09010(.din(w_n8838_0[0]),.dout(n9276),.clk(gclk));
	jand g09011(.dina(w_asqrt23_14[1]),.dinb(n9276),.dout(n9277),.clk(gclk));
	jand g09012(.dina(w_n9277_0[1]),.dinb(w_n8845_0[0]),.dout(n9278),.clk(gclk));
	jor g09013(.dina(n9278),.dinb(w_n8843_0[0]),.dout(n9279),.clk(gclk));
	jand g09014(.dina(w_n9277_0[0]),.dinb(w_n8846_0[0]),.dout(n9280),.clk(gclk));
	jnot g09015(.din(n9280),.dout(n9281),.clk(gclk));
	jand g09016(.dina(n9281),.dinb(n9279),.dout(n9282),.clk(gclk));
	jnot g09017(.din(n9282),.dout(n9283),.clk(gclk));
	jor g09018(.dina(w_n9283_0[1]),.dinb(w_n9275_0[1]),.dout(n9284),.clk(gclk));
	jand g09019(.dina(n9284),.dinb(w_n9273_0[1]),.dout(n9285),.clk(gclk));
	jor g09020(.dina(w_n9285_0[2]),.dinb(w_n199_26[1]),.dout(n9286),.clk(gclk));
	jand g09021(.dina(w_n9285_0[1]),.dinb(w_n199_26[0]),.dout(n9287),.clk(gclk));
	jxor g09022(.dina(w_n8847_0[0]),.dinb(w_n223_22[1]),.dout(n9288),.clk(gclk));
	jor g09023(.dina(n9288),.dinb(w_n8898_19[1]),.dout(n9289),.clk(gclk));
	jxor g09024(.dina(n9289),.dinb(w_n8858_0[0]),.dout(n9290),.clk(gclk));
	jor g09025(.dina(w_n9290_0[1]),.dinb(n9287),.dout(n9291),.clk(gclk));
	jand g09026(.dina(n9291),.dinb(n9286),.dout(n9292),.clk(gclk));
	jnot g09027(.din(w_n8863_0[0]),.dout(n9293),.clk(gclk));
	jor g09028(.dina(n9293),.dinb(w_n8861_0[0]),.dout(n9294),.clk(gclk));
	jor g09029(.dina(n9294),.dinb(w_n8898_19[0]),.dout(n9295),.clk(gclk));
	jxor g09030(.dina(n9295),.dinb(w_n8872_0[0]),.dout(n9296),.clk(gclk));
	jand g09031(.dina(w_asqrt23_14[0]),.dinb(w_n8886_0[1]),.dout(n9297),.clk(gclk));
	jand g09032(.dina(w_n9297_0[1]),.dinb(w_n8874_1[0]),.dout(n9298),.clk(gclk));
	jor g09033(.dina(n9298),.dinb(w_n8920_0[0]),.dout(n9299),.clk(gclk));
	jor g09034(.dina(n9299),.dinb(w_n9296_0[2]),.dout(n9300),.clk(gclk));
	jor g09035(.dina(n9300),.dinb(w_n9292_0[2]),.dout(n9301),.clk(gclk));
	jand g09036(.dina(n9301),.dinb(w_n194_25[1]),.dout(n9302),.clk(gclk));
	jand g09037(.dina(w_n9296_0[1]),.dinb(w_n9292_0[1]),.dout(n9303),.clk(gclk));
	jor g09038(.dina(w_n9297_0[0]),.dinb(w_n8874_0[2]),.dout(n9304),.clk(gclk));
	jand g09039(.dina(w_n8886_0[0]),.dinb(w_n8874_0[1]),.dout(n9305),.clk(gclk));
	jor g09040(.dina(n9305),.dinb(w_n194_25[0]),.dout(n9306),.clk(gclk));
	jnot g09041(.din(n9306),.dout(n9307),.clk(gclk));
	jand g09042(.dina(n9307),.dinb(n9304),.dout(n9308),.clk(gclk));
	jor g09043(.dina(w_n9308_0[1]),.dinb(w_n9303_0[2]),.dout(n9311),.clk(gclk));
	jor g09044(.dina(n9311),.dinb(w_n9302_0[1]),.dout(asqrt_fa_23),.clk(gclk));
	jxor g09045(.dina(w_n9066_0[0]),.dinb(w_n3371_17[1]),.dout(n9313),.clk(gclk));
	jand g09046(.dina(n9313),.dinb(w_asqrt22_31),.dout(n9314),.clk(gclk));
	jxor g09047(.dina(n9314),.dinb(w_n8901_0[0]),.dout(n9315),.clk(gclk));
	jnot g09048(.din(w_n9315_0[1]),.dout(n9316),.clk(gclk));
	jand g09049(.dina(w_asqrt22_30[2]),.dinb(w_a44_0[0]),.dout(n9317),.clk(gclk));
	jnot g09050(.din(w_a42_0[1]),.dout(n9318),.clk(gclk));
	jnot g09051(.din(w_a43_0[1]),.dout(n9319),.clk(gclk));
	jand g09052(.dina(w_n8903_1[0]),.dinb(w_n9319_0[1]),.dout(n9320),.clk(gclk));
	jand g09053(.dina(n9320),.dinb(w_n9318_1[1]),.dout(n9321),.clk(gclk));
	jor g09054(.dina(n9321),.dinb(n9317),.dout(n9322),.clk(gclk));
	jand g09055(.dina(w_n9322_0[2]),.dinb(w_asqrt23_13[2]),.dout(n9323),.clk(gclk));
	jand g09056(.dina(w_asqrt22_30[1]),.dinb(w_n8903_0[2]),.dout(n9324),.clk(gclk));
	jxor g09057(.dina(w_n9324_0[1]),.dinb(w_n8904_0[1]),.dout(n9325),.clk(gclk));
	jor g09058(.dina(w_n9322_0[1]),.dinb(w_asqrt23_13[1]),.dout(n9326),.clk(gclk));
	jand g09059(.dina(n9326),.dinb(w_n9325_0[1]),.dout(n9327),.clk(gclk));
	jor g09060(.dina(w_n9327_0[1]),.dinb(w_n9323_0[1]),.dout(n9328),.clk(gclk));
	jand g09061(.dina(n9328),.dinb(w_asqrt24_17[1]),.dout(n9329),.clk(gclk));
	jor g09062(.dina(w_n9323_0[0]),.dinb(w_asqrt24_17[0]),.dout(n9330),.clk(gclk));
	jor g09063(.dina(n9330),.dinb(w_n9327_0[0]),.dout(n9331),.clk(gclk));
	jand g09064(.dina(w_n9324_0[0]),.dinb(w_n8904_0[0]),.dout(n9332),.clk(gclk));
	jnot g09065(.din(w_n9302_0[0]),.dout(n9333),.clk(gclk));
	jnot g09066(.din(w_n9303_0[1]),.dout(n9334),.clk(gclk));
	jnot g09067(.din(w_n9308_0[0]),.dout(n9335),.clk(gclk));
	jand g09068(.dina(n9335),.dinb(w_asqrt23_13[0]),.dout(n9336),.clk(gclk));
	jand g09069(.dina(n9336),.dinb(n9334),.dout(n9337),.clk(gclk));
	jand g09070(.dina(n9337),.dinb(n9333),.dout(n9338),.clk(gclk));
	jor g09071(.dina(n9338),.dinb(n9332),.dout(n9339),.clk(gclk));
	jxor g09072(.dina(n9339),.dinb(w_n8460_0[1]),.dout(n9340),.clk(gclk));
	jand g09073(.dina(w_n9340_0[1]),.dinb(w_n9331_0[1]),.dout(n9341),.clk(gclk));
	jor g09074(.dina(n9341),.dinb(w_n9329_0[1]),.dout(n9342),.clk(gclk));
	jand g09075(.dina(w_n9342_0[2]),.dinb(w_asqrt25_13[2]),.dout(n9343),.clk(gclk));
	jor g09076(.dina(w_n9342_0[1]),.dinb(w_asqrt25_13[1]),.dout(n9344),.clk(gclk));
	jxor g09077(.dina(w_n8908_0[0]),.dinb(w_n8893_14[2]),.dout(n9345),.clk(gclk));
	jand g09078(.dina(n9345),.dinb(w_asqrt22_30[0]),.dout(n9346),.clk(gclk));
	jxor g09079(.dina(n9346),.dinb(w_n8911_0[0]),.dout(n9347),.clk(gclk));
	jnot g09080(.din(w_n9347_0[1]),.dout(n9348),.clk(gclk));
	jand g09081(.dina(n9348),.dinb(n9344),.dout(n9349),.clk(gclk));
	jor g09082(.dina(w_n9349_0[1]),.dinb(w_n9343_0[1]),.dout(n9350),.clk(gclk));
	jand g09083(.dina(n9350),.dinb(w_asqrt26_17[1]),.dout(n9351),.clk(gclk));
	jnot g09084(.din(w_n8917_0[0]),.dout(n9352),.clk(gclk));
	jand g09085(.dina(n9352),.dinb(w_n8915_0[0]),.dout(n9353),.clk(gclk));
	jand g09086(.dina(n9353),.dinb(w_asqrt22_29[2]),.dout(n9354),.clk(gclk));
	jxor g09087(.dina(n9354),.dinb(w_n8925_0[0]),.dout(n9355),.clk(gclk));
	jnot g09088(.din(n9355),.dout(n9356),.clk(gclk));
	jor g09089(.dina(w_n9343_0[0]),.dinb(w_asqrt26_17[0]),.dout(n9357),.clk(gclk));
	jor g09090(.dina(n9357),.dinb(w_n9349_0[0]),.dout(n9358),.clk(gclk));
	jand g09091(.dina(w_n9358_0[1]),.dinb(w_n9356_0[1]),.dout(n9359),.clk(gclk));
	jor g09092(.dina(w_n9359_0[1]),.dinb(w_n9351_0[1]),.dout(n9360),.clk(gclk));
	jand g09093(.dina(w_n9360_0[2]),.dinb(w_asqrt27_13[2]),.dout(n9361),.clk(gclk));
	jor g09094(.dina(w_n9360_0[1]),.dinb(w_asqrt27_13[1]),.dout(n9362),.clk(gclk));
	jnot g09095(.din(w_n8932_0[0]),.dout(n9363),.clk(gclk));
	jxor g09096(.dina(w_n8927_0[0]),.dinb(w_n8053_14[2]),.dout(n9364),.clk(gclk));
	jand g09097(.dina(n9364),.dinb(w_asqrt22_29[1]),.dout(n9365),.clk(gclk));
	jxor g09098(.dina(n9365),.dinb(n9363),.dout(n9366),.clk(gclk));
	jand g09099(.dina(w_n9366_0[1]),.dinb(n9362),.dout(n9367),.clk(gclk));
	jor g09100(.dina(w_n9367_0[1]),.dinb(w_n9361_0[1]),.dout(n9368),.clk(gclk));
	jand g09101(.dina(n9368),.dinb(w_asqrt28_17[1]),.dout(n9369),.clk(gclk));
	jor g09102(.dina(w_n9361_0[0]),.dinb(w_asqrt28_17[0]),.dout(n9370),.clk(gclk));
	jor g09103(.dina(n9370),.dinb(w_n9367_0[0]),.dout(n9371),.clk(gclk));
	jnot g09104(.din(w_n8939_0[0]),.dout(n9372),.clk(gclk));
	jnot g09105(.din(w_n8941_0[0]),.dout(n9373),.clk(gclk));
	jand g09106(.dina(w_asqrt22_29[0]),.dinb(w_n8935_0[0]),.dout(n9374),.clk(gclk));
	jand g09107(.dina(w_n9374_0[1]),.dinb(n9373),.dout(n9375),.clk(gclk));
	jor g09108(.dina(n9375),.dinb(n9372),.dout(n9376),.clk(gclk));
	jnot g09109(.din(w_n8942_0[0]),.dout(n9377),.clk(gclk));
	jand g09110(.dina(w_n9374_0[0]),.dinb(n9377),.dout(n9378),.clk(gclk));
	jnot g09111(.din(n9378),.dout(n9379),.clk(gclk));
	jand g09112(.dina(n9379),.dinb(n9376),.dout(n9380),.clk(gclk));
	jand g09113(.dina(w_n9380_0[1]),.dinb(w_n9371_0[1]),.dout(n9381),.clk(gclk));
	jor g09114(.dina(n9381),.dinb(w_n9369_0[1]),.dout(n9382),.clk(gclk));
	jand g09115(.dina(w_n9382_0[2]),.dinb(w_asqrt29_14[0]),.dout(n9383),.clk(gclk));
	jor g09116(.dina(w_n9382_0[1]),.dinb(w_asqrt29_13[2]),.dout(n9384),.clk(gclk));
	jxor g09117(.dina(w_n8943_0[0]),.dinb(w_n7260_15[1]),.dout(n9385),.clk(gclk));
	jand g09118(.dina(n9385),.dinb(w_asqrt22_28[2]),.dout(n9386),.clk(gclk));
	jxor g09119(.dina(n9386),.dinb(w_n8948_0[0]),.dout(n9387),.clk(gclk));
	jand g09120(.dina(w_n9387_0[1]),.dinb(n9384),.dout(n9388),.clk(gclk));
	jor g09121(.dina(w_n9388_0[1]),.dinb(w_n9383_0[1]),.dout(n9389),.clk(gclk));
	jand g09122(.dina(n9389),.dinb(w_asqrt30_17[1]),.dout(n9390),.clk(gclk));
	jnot g09123(.din(w_n8954_0[0]),.dout(n9391),.clk(gclk));
	jand g09124(.dina(n9391),.dinb(w_n8952_0[0]),.dout(n9392),.clk(gclk));
	jand g09125(.dina(n9392),.dinb(w_asqrt22_28[1]),.dout(n9393),.clk(gclk));
	jxor g09126(.dina(n9393),.dinb(w_n8963_0[0]),.dout(n9394),.clk(gclk));
	jnot g09127(.din(n9394),.dout(n9395),.clk(gclk));
	jor g09128(.dina(w_n9383_0[0]),.dinb(w_asqrt30_17[0]),.dout(n9396),.clk(gclk));
	jor g09129(.dina(n9396),.dinb(w_n9388_0[0]),.dout(n9397),.clk(gclk));
	jand g09130(.dina(w_n9397_0[1]),.dinb(w_n9395_0[1]),.dout(n9398),.clk(gclk));
	jor g09131(.dina(w_n9398_0[1]),.dinb(w_n9390_0[1]),.dout(n9399),.clk(gclk));
	jand g09132(.dina(w_n9399_0[2]),.dinb(w_asqrt31_14[0]),.dout(n9400),.clk(gclk));
	jor g09133(.dina(w_n9399_0[1]),.dinb(w_asqrt31_13[2]),.dout(n9401),.clk(gclk));
	jxor g09134(.dina(w_n8965_0[0]),.dinb(w_n6500_15[1]),.dout(n9402),.clk(gclk));
	jand g09135(.dina(n9402),.dinb(w_asqrt22_28[0]),.dout(n9403),.clk(gclk));
	jxor g09136(.dina(n9403),.dinb(w_n8971_0[0]),.dout(n9404),.clk(gclk));
	jand g09137(.dina(w_n9404_0[1]),.dinb(n9401),.dout(n9405),.clk(gclk));
	jor g09138(.dina(w_n9405_0[1]),.dinb(w_n9400_0[1]),.dout(n9406),.clk(gclk));
	jand g09139(.dina(n9406),.dinb(w_asqrt32_17[1]),.dout(n9407),.clk(gclk));
	jor g09140(.dina(w_n9400_0[0]),.dinb(w_asqrt32_17[0]),.dout(n9408),.clk(gclk));
	jor g09141(.dina(n9408),.dinb(w_n9405_0[0]),.dout(n9409),.clk(gclk));
	jnot g09142(.din(w_n8979_0[0]),.dout(n9410),.clk(gclk));
	jnot g09143(.din(w_n8981_0[0]),.dout(n9411),.clk(gclk));
	jand g09144(.dina(w_asqrt22_27[2]),.dinb(w_n8975_0[0]),.dout(n9412),.clk(gclk));
	jand g09145(.dina(w_n9412_0[1]),.dinb(n9411),.dout(n9413),.clk(gclk));
	jor g09146(.dina(n9413),.dinb(n9410),.dout(n9414),.clk(gclk));
	jnot g09147(.din(w_n8982_0[0]),.dout(n9415),.clk(gclk));
	jand g09148(.dina(w_n9412_0[0]),.dinb(n9415),.dout(n9416),.clk(gclk));
	jnot g09149(.din(n9416),.dout(n9417),.clk(gclk));
	jand g09150(.dina(n9417),.dinb(n9414),.dout(n9418),.clk(gclk));
	jand g09151(.dina(w_n9418_0[1]),.dinb(w_n9409_0[1]),.dout(n9419),.clk(gclk));
	jor g09152(.dina(n9419),.dinb(w_n9407_0[1]),.dout(n9420),.clk(gclk));
	jand g09153(.dina(w_n9420_0[1]),.dinb(w_asqrt33_14[1]),.dout(n9421),.clk(gclk));
	jxor g09154(.dina(w_n8983_0[0]),.dinb(w_n5788_15[2]),.dout(n9422),.clk(gclk));
	jand g09155(.dina(n9422),.dinb(w_asqrt22_27[1]),.dout(n9423),.clk(gclk));
	jxor g09156(.dina(n9423),.dinb(w_n8990_0[0]),.dout(n9424),.clk(gclk));
	jnot g09157(.din(n9424),.dout(n9425),.clk(gclk));
	jor g09158(.dina(w_n9420_0[0]),.dinb(w_asqrt33_14[0]),.dout(n9426),.clk(gclk));
	jand g09159(.dina(w_n9426_0[1]),.dinb(w_n9425_0[1]),.dout(n9427),.clk(gclk));
	jor g09160(.dina(w_n9427_0[2]),.dinb(w_n9421_0[2]),.dout(n9428),.clk(gclk));
	jand g09161(.dina(n9428),.dinb(w_asqrt34_17[1]),.dout(n9429),.clk(gclk));
	jnot g09162(.din(w_n8995_0[0]),.dout(n9430),.clk(gclk));
	jand g09163(.dina(n9430),.dinb(w_n8993_0[0]),.dout(n9431),.clk(gclk));
	jand g09164(.dina(n9431),.dinb(w_asqrt22_27[0]),.dout(n9432),.clk(gclk));
	jxor g09165(.dina(n9432),.dinb(w_n9003_0[0]),.dout(n9433),.clk(gclk));
	jnot g09166(.din(n9433),.dout(n9434),.clk(gclk));
	jor g09167(.dina(w_n9421_0[1]),.dinb(w_asqrt34_17[0]),.dout(n9435),.clk(gclk));
	jor g09168(.dina(n9435),.dinb(w_n9427_0[1]),.dout(n9436),.clk(gclk));
	jand g09169(.dina(w_n9436_0[1]),.dinb(w_n9434_0[1]),.dout(n9437),.clk(gclk));
	jor g09170(.dina(w_n9437_0[1]),.dinb(w_n9429_0[1]),.dout(n9438),.clk(gclk));
	jand g09171(.dina(w_n9438_0[2]),.dinb(w_asqrt35_14[1]),.dout(n9439),.clk(gclk));
	jor g09172(.dina(w_n9438_0[1]),.dinb(w_asqrt35_14[0]),.dout(n9440),.clk(gclk));
	jnot g09173(.din(w_n9009_0[0]),.dout(n9441),.clk(gclk));
	jnot g09174(.din(w_n9010_0[0]),.dout(n9442),.clk(gclk));
	jand g09175(.dina(w_asqrt22_26[2]),.dinb(w_n9006_0[0]),.dout(n9443),.clk(gclk));
	jand g09176(.dina(w_n9443_0[1]),.dinb(n9442),.dout(n9444),.clk(gclk));
	jor g09177(.dina(n9444),.dinb(n9441),.dout(n9445),.clk(gclk));
	jnot g09178(.din(w_n9011_0[0]),.dout(n9446),.clk(gclk));
	jand g09179(.dina(w_n9443_0[0]),.dinb(n9446),.dout(n9447),.clk(gclk));
	jnot g09180(.din(n9447),.dout(n9448),.clk(gclk));
	jand g09181(.dina(n9448),.dinb(n9445),.dout(n9449),.clk(gclk));
	jand g09182(.dina(w_n9449_0[1]),.dinb(n9440),.dout(n9450),.clk(gclk));
	jor g09183(.dina(w_n9450_0[1]),.dinb(w_n9439_0[1]),.dout(n9451),.clk(gclk));
	jand g09184(.dina(n9451),.dinb(w_asqrt36_17[1]),.dout(n9452),.clk(gclk));
	jor g09185(.dina(w_n9439_0[0]),.dinb(w_asqrt36_17[0]),.dout(n9453),.clk(gclk));
	jor g09186(.dina(n9453),.dinb(w_n9450_0[0]),.dout(n9454),.clk(gclk));
	jnot g09187(.din(w_n9017_0[0]),.dout(n9455),.clk(gclk));
	jnot g09188(.din(w_n9019_0[0]),.dout(n9456),.clk(gclk));
	jand g09189(.dina(w_asqrt22_26[1]),.dinb(w_n9013_0[0]),.dout(n9457),.clk(gclk));
	jand g09190(.dina(w_n9457_0[1]),.dinb(n9456),.dout(n9458),.clk(gclk));
	jor g09191(.dina(n9458),.dinb(n9455),.dout(n9459),.clk(gclk));
	jnot g09192(.din(w_n9020_0[0]),.dout(n9460),.clk(gclk));
	jand g09193(.dina(w_n9457_0[0]),.dinb(n9460),.dout(n9461),.clk(gclk));
	jnot g09194(.din(n9461),.dout(n9462),.clk(gclk));
	jand g09195(.dina(n9462),.dinb(n9459),.dout(n9463),.clk(gclk));
	jand g09196(.dina(w_n9463_0[1]),.dinb(w_n9454_0[1]),.dout(n9464),.clk(gclk));
	jor g09197(.dina(n9464),.dinb(w_n9452_0[1]),.dout(n9465),.clk(gclk));
	jand g09198(.dina(w_n9465_0[1]),.dinb(w_asqrt37_14[2]),.dout(n9466),.clk(gclk));
	jxor g09199(.dina(w_n9021_0[0]),.dinb(w_n4494_16[2]),.dout(n9467),.clk(gclk));
	jand g09200(.dina(n9467),.dinb(w_asqrt22_26[0]),.dout(n9468),.clk(gclk));
	jxor g09201(.dina(n9468),.dinb(w_n9031_0[0]),.dout(n9469),.clk(gclk));
	jnot g09202(.din(n9469),.dout(n9470),.clk(gclk));
	jor g09203(.dina(w_n9465_0[0]),.dinb(w_asqrt37_14[1]),.dout(n9471),.clk(gclk));
	jand g09204(.dina(w_n9471_0[1]),.dinb(w_n9470_0[1]),.dout(n9472),.clk(gclk));
	jor g09205(.dina(w_n9472_0[2]),.dinb(w_n9466_0[2]),.dout(n9473),.clk(gclk));
	jand g09206(.dina(n9473),.dinb(w_asqrt38_17[1]),.dout(n9474),.clk(gclk));
	jnot g09207(.din(w_n9036_0[0]),.dout(n9475),.clk(gclk));
	jand g09208(.dina(n9475),.dinb(w_n9034_0[0]),.dout(n9476),.clk(gclk));
	jand g09209(.dina(n9476),.dinb(w_asqrt22_25[2]),.dout(n9477),.clk(gclk));
	jxor g09210(.dina(n9477),.dinb(w_n9044_0[0]),.dout(n9478),.clk(gclk));
	jnot g09211(.din(n9478),.dout(n9479),.clk(gclk));
	jor g09212(.dina(w_n9466_0[1]),.dinb(w_asqrt38_17[0]),.dout(n9480),.clk(gclk));
	jor g09213(.dina(n9480),.dinb(w_n9472_0[1]),.dout(n9481),.clk(gclk));
	jand g09214(.dina(w_n9481_0[1]),.dinb(w_n9479_0[1]),.dout(n9482),.clk(gclk));
	jor g09215(.dina(w_n9482_0[1]),.dinb(w_n9474_0[1]),.dout(n9483),.clk(gclk));
	jand g09216(.dina(w_n9483_0[2]),.dinb(w_asqrt39_14[2]),.dout(n9484),.clk(gclk));
	jor g09217(.dina(w_n9483_0[1]),.dinb(w_asqrt39_14[1]),.dout(n9485),.clk(gclk));
	jnot g09218(.din(w_n9050_0[0]),.dout(n9486),.clk(gclk));
	jnot g09219(.din(w_n9051_0[0]),.dout(n9487),.clk(gclk));
	jand g09220(.dina(w_asqrt22_25[1]),.dinb(w_n9047_0[0]),.dout(n9488),.clk(gclk));
	jand g09221(.dina(w_n9488_0[1]),.dinb(n9487),.dout(n9489),.clk(gclk));
	jor g09222(.dina(n9489),.dinb(n9486),.dout(n9490),.clk(gclk));
	jnot g09223(.din(w_n9052_0[0]),.dout(n9491),.clk(gclk));
	jand g09224(.dina(w_n9488_0[0]),.dinb(n9491),.dout(n9492),.clk(gclk));
	jnot g09225(.din(n9492),.dout(n9493),.clk(gclk));
	jand g09226(.dina(n9493),.dinb(n9490),.dout(n9494),.clk(gclk));
	jand g09227(.dina(w_n9494_0[1]),.dinb(n9485),.dout(n9495),.clk(gclk));
	jor g09228(.dina(w_n9495_0[1]),.dinb(w_n9484_0[1]),.dout(n9496),.clk(gclk));
	jand g09229(.dina(n9496),.dinb(w_asqrt40_17[1]),.dout(n9497),.clk(gclk));
	jnot g09230(.din(w_n9056_0[0]),.dout(n9498),.clk(gclk));
	jand g09231(.dina(n9498),.dinb(w_n9054_0[0]),.dout(n9499),.clk(gclk));
	jand g09232(.dina(n9499),.dinb(w_asqrt22_25[0]),.dout(n9500),.clk(gclk));
	jxor g09233(.dina(n9500),.dinb(w_n9064_0[0]),.dout(n9501),.clk(gclk));
	jnot g09234(.din(n9501),.dout(n9502),.clk(gclk));
	jor g09235(.dina(w_n9484_0[0]),.dinb(w_asqrt40_17[0]),.dout(n9503),.clk(gclk));
	jor g09236(.dina(n9503),.dinb(w_n9495_0[0]),.dout(n9504),.clk(gclk));
	jand g09237(.dina(w_n9504_0[1]),.dinb(w_n9502_0[1]),.dout(n9505),.clk(gclk));
	jor g09238(.dina(w_n9505_0[1]),.dinb(w_n9497_0[1]),.dout(n9506),.clk(gclk));
	jand g09239(.dina(w_n9506_0[2]),.dinb(w_asqrt41_15[0]),.dout(n9507),.clk(gclk));
	jor g09240(.dina(w_n9506_0[1]),.dinb(w_asqrt41_14[2]),.dout(n9508),.clk(gclk));
	jand g09241(.dina(n9508),.dinb(w_n9315_0[0]),.dout(n9509),.clk(gclk));
	jor g09242(.dina(w_n9509_0[1]),.dinb(w_n9507_0[1]),.dout(n9510),.clk(gclk));
	jand g09243(.dina(n9510),.dinb(w_asqrt42_17[1]),.dout(n9511),.clk(gclk));
	jor g09244(.dina(w_n9507_0[0]),.dinb(w_asqrt42_17[0]),.dout(n9512),.clk(gclk));
	jor g09245(.dina(n9512),.dinb(w_n9509_0[0]),.dout(n9513),.clk(gclk));
	jnot g09246(.din(w_n9076_0[0]),.dout(n9514),.clk(gclk));
	jnot g09247(.din(w_n9078_0[0]),.dout(n9515),.clk(gclk));
	jand g09248(.dina(w_asqrt22_24[2]),.dinb(w_n9072_0[0]),.dout(n9516),.clk(gclk));
	jand g09249(.dina(w_n9516_0[1]),.dinb(n9515),.dout(n9517),.clk(gclk));
	jor g09250(.dina(n9517),.dinb(n9514),.dout(n9518),.clk(gclk));
	jnot g09251(.din(w_n9079_0[0]),.dout(n9519),.clk(gclk));
	jand g09252(.dina(w_n9516_0[0]),.dinb(n9519),.dout(n9520),.clk(gclk));
	jnot g09253(.din(n9520),.dout(n9521),.clk(gclk));
	jand g09254(.dina(n9521),.dinb(n9518),.dout(n9522),.clk(gclk));
	jand g09255(.dina(w_n9522_0[1]),.dinb(w_n9513_0[1]),.dout(n9523),.clk(gclk));
	jor g09256(.dina(n9523),.dinb(w_n9511_0[1]),.dout(n9524),.clk(gclk));
	jand g09257(.dina(w_n9524_0[2]),.dinb(w_asqrt43_15[0]),.dout(n9525),.clk(gclk));
	jor g09258(.dina(w_n9524_0[1]),.dinb(w_asqrt43_14[2]),.dout(n9526),.clk(gclk));
	jnot g09259(.din(w_n9084_0[0]),.dout(n9527),.clk(gclk));
	jnot g09260(.din(w_n9085_0[0]),.dout(n9528),.clk(gclk));
	jand g09261(.dina(w_asqrt22_24[1]),.dinb(w_n9081_0[0]),.dout(n9529),.clk(gclk));
	jand g09262(.dina(w_n9529_0[1]),.dinb(n9528),.dout(n9530),.clk(gclk));
	jor g09263(.dina(n9530),.dinb(n9527),.dout(n9531),.clk(gclk));
	jnot g09264(.din(w_n9086_0[0]),.dout(n9532),.clk(gclk));
	jand g09265(.dina(w_n9529_0[0]),.dinb(n9532),.dout(n9533),.clk(gclk));
	jnot g09266(.din(n9533),.dout(n9534),.clk(gclk));
	jand g09267(.dina(n9534),.dinb(n9531),.dout(n9535),.clk(gclk));
	jand g09268(.dina(w_n9535_0[1]),.dinb(n9526),.dout(n9536),.clk(gclk));
	jor g09269(.dina(w_n9536_0[1]),.dinb(w_n9525_0[1]),.dout(n9537),.clk(gclk));
	jand g09270(.dina(n9537),.dinb(w_asqrt44_17[1]),.dout(n9538),.clk(gclk));
	jor g09271(.dina(w_n9525_0[0]),.dinb(w_asqrt44_17[0]),.dout(n9539),.clk(gclk));
	jor g09272(.dina(n9539),.dinb(w_n9536_0[0]),.dout(n9540),.clk(gclk));
	jnot g09273(.din(w_n9092_0[0]),.dout(n9541),.clk(gclk));
	jnot g09274(.din(w_n9094_0[0]),.dout(n9542),.clk(gclk));
	jand g09275(.dina(w_asqrt22_24[0]),.dinb(w_n9088_0[0]),.dout(n9543),.clk(gclk));
	jand g09276(.dina(w_n9543_0[1]),.dinb(n9542),.dout(n9544),.clk(gclk));
	jor g09277(.dina(n9544),.dinb(n9541),.dout(n9545),.clk(gclk));
	jnot g09278(.din(w_n9095_0[0]),.dout(n9546),.clk(gclk));
	jand g09279(.dina(w_n9543_0[0]),.dinb(n9546),.dout(n9547),.clk(gclk));
	jnot g09280(.din(n9547),.dout(n9548),.clk(gclk));
	jand g09281(.dina(n9548),.dinb(n9545),.dout(n9549),.clk(gclk));
	jand g09282(.dina(w_n9549_0[1]),.dinb(w_n9540_0[1]),.dout(n9550),.clk(gclk));
	jor g09283(.dina(n9550),.dinb(w_n9538_0[1]),.dout(n9551),.clk(gclk));
	jand g09284(.dina(w_n9551_0[1]),.dinb(w_asqrt45_15[1]),.dout(n9552),.clk(gclk));
	jxor g09285(.dina(w_n9096_0[0]),.dinb(w_n2420_18[1]),.dout(n9553),.clk(gclk));
	jand g09286(.dina(n9553),.dinb(w_asqrt22_23[2]),.dout(n9554),.clk(gclk));
	jxor g09287(.dina(n9554),.dinb(w_n9106_0[0]),.dout(n9555),.clk(gclk));
	jnot g09288(.din(n9555),.dout(n9556),.clk(gclk));
	jor g09289(.dina(w_n9551_0[0]),.dinb(w_asqrt45_15[0]),.dout(n9557),.clk(gclk));
	jand g09290(.dina(w_n9557_0[1]),.dinb(w_n9556_0[1]),.dout(n9558),.clk(gclk));
	jor g09291(.dina(w_n9558_0[2]),.dinb(w_n9552_0[2]),.dout(n9559),.clk(gclk));
	jand g09292(.dina(n9559),.dinb(w_asqrt46_17[1]),.dout(n9560),.clk(gclk));
	jnot g09293(.din(w_n9111_0[0]),.dout(n9561),.clk(gclk));
	jand g09294(.dina(n9561),.dinb(w_n9109_0[0]),.dout(n9562),.clk(gclk));
	jand g09295(.dina(n9562),.dinb(w_asqrt22_23[1]),.dout(n9563),.clk(gclk));
	jxor g09296(.dina(n9563),.dinb(w_n9119_0[0]),.dout(n9564),.clk(gclk));
	jnot g09297(.din(n9564),.dout(n9565),.clk(gclk));
	jor g09298(.dina(w_n9552_0[1]),.dinb(w_asqrt46_17[0]),.dout(n9566),.clk(gclk));
	jor g09299(.dina(n9566),.dinb(w_n9558_0[1]),.dout(n9567),.clk(gclk));
	jand g09300(.dina(w_n9567_0[1]),.dinb(w_n9565_0[1]),.dout(n9568),.clk(gclk));
	jor g09301(.dina(w_n9568_0[1]),.dinb(w_n9560_0[1]),.dout(n9569),.clk(gclk));
	jand g09302(.dina(w_n9569_0[2]),.dinb(w_asqrt47_15[1]),.dout(n9570),.clk(gclk));
	jor g09303(.dina(w_n9569_0[1]),.dinb(w_asqrt47_15[0]),.dout(n9571),.clk(gclk));
	jnot g09304(.din(w_n9125_0[0]),.dout(n9572),.clk(gclk));
	jnot g09305(.din(w_n9126_0[0]),.dout(n9573),.clk(gclk));
	jand g09306(.dina(w_asqrt22_23[0]),.dinb(w_n9122_0[0]),.dout(n9574),.clk(gclk));
	jand g09307(.dina(w_n9574_0[1]),.dinb(n9573),.dout(n9575),.clk(gclk));
	jor g09308(.dina(n9575),.dinb(n9572),.dout(n9576),.clk(gclk));
	jnot g09309(.din(w_n9127_0[0]),.dout(n9577),.clk(gclk));
	jand g09310(.dina(w_n9574_0[0]),.dinb(n9577),.dout(n9578),.clk(gclk));
	jnot g09311(.din(n9578),.dout(n9579),.clk(gclk));
	jand g09312(.dina(n9579),.dinb(n9576),.dout(n9580),.clk(gclk));
	jand g09313(.dina(w_n9580_0[1]),.dinb(n9571),.dout(n9581),.clk(gclk));
	jor g09314(.dina(w_n9581_0[1]),.dinb(w_n9570_0[1]),.dout(n9582),.clk(gclk));
	jand g09315(.dina(n9582),.dinb(w_asqrt48_17[1]),.dout(n9583),.clk(gclk));
	jor g09316(.dina(w_n9570_0[0]),.dinb(w_asqrt48_17[0]),.dout(n9584),.clk(gclk));
	jor g09317(.dina(n9584),.dinb(w_n9581_0[0]),.dout(n9585),.clk(gclk));
	jnot g09318(.din(w_n9133_0[0]),.dout(n9586),.clk(gclk));
	jnot g09319(.din(w_n9135_0[0]),.dout(n9587),.clk(gclk));
	jand g09320(.dina(w_asqrt22_22[2]),.dinb(w_n9129_0[0]),.dout(n9588),.clk(gclk));
	jand g09321(.dina(w_n9588_0[1]),.dinb(n9587),.dout(n9589),.clk(gclk));
	jor g09322(.dina(n9589),.dinb(n9586),.dout(n9590),.clk(gclk));
	jnot g09323(.din(w_n9136_0[0]),.dout(n9591),.clk(gclk));
	jand g09324(.dina(w_n9588_0[0]),.dinb(n9591),.dout(n9592),.clk(gclk));
	jnot g09325(.din(n9592),.dout(n9593),.clk(gclk));
	jand g09326(.dina(n9593),.dinb(n9590),.dout(n9594),.clk(gclk));
	jand g09327(.dina(w_n9594_0[1]),.dinb(w_n9585_0[1]),.dout(n9595),.clk(gclk));
	jor g09328(.dina(n9595),.dinb(w_n9583_0[1]),.dout(n9596),.clk(gclk));
	jand g09329(.dina(w_n9596_0[1]),.dinb(w_asqrt49_15[2]),.dout(n9597),.clk(gclk));
	jxor g09330(.dina(w_n9137_0[0]),.dinb(w_n1641_19[0]),.dout(n9598),.clk(gclk));
	jand g09331(.dina(n9598),.dinb(w_asqrt22_22[1]),.dout(n9599),.clk(gclk));
	jxor g09332(.dina(n9599),.dinb(w_n9147_0[0]),.dout(n9600),.clk(gclk));
	jnot g09333(.din(n9600),.dout(n9601),.clk(gclk));
	jor g09334(.dina(w_n9596_0[0]),.dinb(w_asqrt49_15[1]),.dout(n9602),.clk(gclk));
	jand g09335(.dina(w_n9602_0[1]),.dinb(w_n9601_0[1]),.dout(n9603),.clk(gclk));
	jor g09336(.dina(w_n9603_0[2]),.dinb(w_n9597_0[2]),.dout(n9604),.clk(gclk));
	jand g09337(.dina(n9604),.dinb(w_asqrt50_17[1]),.dout(n9605),.clk(gclk));
	jnot g09338(.din(w_n9152_0[0]),.dout(n9606),.clk(gclk));
	jand g09339(.dina(n9606),.dinb(w_n9150_0[0]),.dout(n9607),.clk(gclk));
	jand g09340(.dina(n9607),.dinb(w_asqrt22_22[0]),.dout(n9608),.clk(gclk));
	jxor g09341(.dina(n9608),.dinb(w_n9160_0[0]),.dout(n9609),.clk(gclk));
	jnot g09342(.din(n9609),.dout(n9610),.clk(gclk));
	jor g09343(.dina(w_n9597_0[1]),.dinb(w_asqrt50_17[0]),.dout(n9611),.clk(gclk));
	jor g09344(.dina(n9611),.dinb(w_n9603_0[1]),.dout(n9612),.clk(gclk));
	jand g09345(.dina(w_n9612_0[1]),.dinb(w_n9610_0[1]),.dout(n9613),.clk(gclk));
	jor g09346(.dina(w_n9613_0[1]),.dinb(w_n9605_0[1]),.dout(n9614),.clk(gclk));
	jand g09347(.dina(w_n9614_0[2]),.dinb(w_asqrt51_15[2]),.dout(n9615),.clk(gclk));
	jor g09348(.dina(w_n9614_0[1]),.dinb(w_asqrt51_15[1]),.dout(n9616),.clk(gclk));
	jnot g09349(.din(w_n9166_0[0]),.dout(n9617),.clk(gclk));
	jnot g09350(.din(w_n9167_0[0]),.dout(n9618),.clk(gclk));
	jand g09351(.dina(w_asqrt22_21[2]),.dinb(w_n9163_0[0]),.dout(n9619),.clk(gclk));
	jand g09352(.dina(w_n9619_0[1]),.dinb(n9618),.dout(n9620),.clk(gclk));
	jor g09353(.dina(n9620),.dinb(n9617),.dout(n9621),.clk(gclk));
	jnot g09354(.din(w_n9168_0[0]),.dout(n9622),.clk(gclk));
	jand g09355(.dina(w_n9619_0[0]),.dinb(n9622),.dout(n9623),.clk(gclk));
	jnot g09356(.din(n9623),.dout(n9624),.clk(gclk));
	jand g09357(.dina(n9624),.dinb(n9621),.dout(n9625),.clk(gclk));
	jand g09358(.dina(w_n9625_0[1]),.dinb(n9616),.dout(n9626),.clk(gclk));
	jor g09359(.dina(w_n9626_0[1]),.dinb(w_n9615_0[1]),.dout(n9627),.clk(gclk));
	jand g09360(.dina(n9627),.dinb(w_asqrt52_17[1]),.dout(n9628),.clk(gclk));
	jor g09361(.dina(w_n9615_0[0]),.dinb(w_asqrt52_17[0]),.dout(n9629),.clk(gclk));
	jor g09362(.dina(n9629),.dinb(w_n9626_0[0]),.dout(n9630),.clk(gclk));
	jnot g09363(.din(w_n9174_0[0]),.dout(n9631),.clk(gclk));
	jnot g09364(.din(w_n9176_0[0]),.dout(n9632),.clk(gclk));
	jand g09365(.dina(w_asqrt22_21[1]),.dinb(w_n9170_0[0]),.dout(n9633),.clk(gclk));
	jand g09366(.dina(w_n9633_0[1]),.dinb(n9632),.dout(n9634),.clk(gclk));
	jor g09367(.dina(n9634),.dinb(n9631),.dout(n9635),.clk(gclk));
	jnot g09368(.din(w_n9177_0[0]),.dout(n9636),.clk(gclk));
	jand g09369(.dina(w_n9633_0[0]),.dinb(n9636),.dout(n9637),.clk(gclk));
	jnot g09370(.din(n9637),.dout(n9638),.clk(gclk));
	jand g09371(.dina(n9638),.dinb(n9635),.dout(n9639),.clk(gclk));
	jand g09372(.dina(w_n9639_0[1]),.dinb(w_n9630_0[1]),.dout(n9640),.clk(gclk));
	jor g09373(.dina(n9640),.dinb(w_n9628_0[1]),.dout(n9641),.clk(gclk));
	jand g09374(.dina(w_n9641_0[1]),.dinb(w_asqrt53_16[0]),.dout(n9642),.clk(gclk));
	jxor g09375(.dina(w_n9178_0[0]),.dinb(w_n1034_20[0]),.dout(n9643),.clk(gclk));
	jand g09376(.dina(n9643),.dinb(w_asqrt22_21[0]),.dout(n9644),.clk(gclk));
	jxor g09377(.dina(n9644),.dinb(w_n9188_0[0]),.dout(n9645),.clk(gclk));
	jnot g09378(.din(n9645),.dout(n9646),.clk(gclk));
	jor g09379(.dina(w_n9641_0[0]),.dinb(w_asqrt53_15[2]),.dout(n9647),.clk(gclk));
	jand g09380(.dina(w_n9647_0[1]),.dinb(w_n9646_0[1]),.dout(n9648),.clk(gclk));
	jor g09381(.dina(w_n9648_0[2]),.dinb(w_n9642_0[2]),.dout(n9649),.clk(gclk));
	jand g09382(.dina(n9649),.dinb(w_asqrt54_17[1]),.dout(n9650),.clk(gclk));
	jnot g09383(.din(w_n9193_0[0]),.dout(n9651),.clk(gclk));
	jand g09384(.dina(n9651),.dinb(w_n9191_0[0]),.dout(n9652),.clk(gclk));
	jand g09385(.dina(n9652),.dinb(w_asqrt22_20[2]),.dout(n9653),.clk(gclk));
	jxor g09386(.dina(n9653),.dinb(w_n9201_0[0]),.dout(n9654),.clk(gclk));
	jnot g09387(.din(n9654),.dout(n9655),.clk(gclk));
	jor g09388(.dina(w_n9642_0[1]),.dinb(w_asqrt54_17[0]),.dout(n9656),.clk(gclk));
	jor g09389(.dina(n9656),.dinb(w_n9648_0[1]),.dout(n9657),.clk(gclk));
	jand g09390(.dina(w_n9657_0[1]),.dinb(w_n9655_0[1]),.dout(n9658),.clk(gclk));
	jor g09391(.dina(w_n9658_0[1]),.dinb(w_n9650_0[1]),.dout(n9659),.clk(gclk));
	jand g09392(.dina(w_n9659_0[2]),.dinb(w_asqrt55_16[1]),.dout(n9660),.clk(gclk));
	jor g09393(.dina(w_n9659_0[1]),.dinb(w_asqrt55_16[0]),.dout(n9661),.clk(gclk));
	jnot g09394(.din(w_n9207_0[0]),.dout(n9662),.clk(gclk));
	jnot g09395(.din(w_n9208_0[0]),.dout(n9663),.clk(gclk));
	jand g09396(.dina(w_asqrt22_20[1]),.dinb(w_n9204_0[0]),.dout(n9664),.clk(gclk));
	jand g09397(.dina(w_n9664_0[1]),.dinb(n9663),.dout(n9665),.clk(gclk));
	jor g09398(.dina(n9665),.dinb(n9662),.dout(n9666),.clk(gclk));
	jnot g09399(.din(w_n9209_0[0]),.dout(n9667),.clk(gclk));
	jand g09400(.dina(w_n9664_0[0]),.dinb(n9667),.dout(n9668),.clk(gclk));
	jnot g09401(.din(n9668),.dout(n9669),.clk(gclk));
	jand g09402(.dina(n9669),.dinb(n9666),.dout(n9670),.clk(gclk));
	jand g09403(.dina(w_n9670_0[1]),.dinb(n9661),.dout(n9671),.clk(gclk));
	jor g09404(.dina(w_n9671_0[1]),.dinb(w_n9660_0[1]),.dout(n9672),.clk(gclk));
	jand g09405(.dina(n9672),.dinb(w_asqrt56_17[1]),.dout(n9673),.clk(gclk));
	jor g09406(.dina(w_n9660_0[0]),.dinb(w_asqrt56_17[0]),.dout(n9674),.clk(gclk));
	jor g09407(.dina(n9674),.dinb(w_n9671_0[0]),.dout(n9675),.clk(gclk));
	jnot g09408(.din(w_n9215_0[0]),.dout(n9676),.clk(gclk));
	jnot g09409(.din(w_n9217_0[0]),.dout(n9677),.clk(gclk));
	jand g09410(.dina(w_asqrt22_20[0]),.dinb(w_n9211_0[0]),.dout(n9678),.clk(gclk));
	jand g09411(.dina(w_n9678_0[1]),.dinb(n9677),.dout(n9679),.clk(gclk));
	jor g09412(.dina(n9679),.dinb(n9676),.dout(n9680),.clk(gclk));
	jnot g09413(.din(w_n9218_0[0]),.dout(n9681),.clk(gclk));
	jand g09414(.dina(w_n9678_0[0]),.dinb(n9681),.dout(n9682),.clk(gclk));
	jnot g09415(.din(n9682),.dout(n9683),.clk(gclk));
	jand g09416(.dina(n9683),.dinb(n9680),.dout(n9684),.clk(gclk));
	jand g09417(.dina(w_n9684_0[1]),.dinb(w_n9675_0[1]),.dout(n9685),.clk(gclk));
	jor g09418(.dina(n9685),.dinb(w_n9673_0[1]),.dout(n9686),.clk(gclk));
	jand g09419(.dina(w_n9686_0[1]),.dinb(w_asqrt57_16[2]),.dout(n9687),.clk(gclk));
	jxor g09420(.dina(w_n9219_0[0]),.dinb(w_n590_20[2]),.dout(n9688),.clk(gclk));
	jand g09421(.dina(n9688),.dinb(w_asqrt22_19[2]),.dout(n9689),.clk(gclk));
	jxor g09422(.dina(n9689),.dinb(w_n9229_0[0]),.dout(n9690),.clk(gclk));
	jnot g09423(.din(n9690),.dout(n9691),.clk(gclk));
	jor g09424(.dina(w_n9686_0[0]),.dinb(w_asqrt57_16[1]),.dout(n9692),.clk(gclk));
	jand g09425(.dina(w_n9692_0[1]),.dinb(w_n9691_0[1]),.dout(n9693),.clk(gclk));
	jor g09426(.dina(w_n9693_0[2]),.dinb(w_n9687_0[2]),.dout(n9694),.clk(gclk));
	jand g09427(.dina(n9694),.dinb(w_asqrt58_17[1]),.dout(n9695),.clk(gclk));
	jnot g09428(.din(w_n9234_0[0]),.dout(n9696),.clk(gclk));
	jand g09429(.dina(n9696),.dinb(w_n9232_0[0]),.dout(n9697),.clk(gclk));
	jand g09430(.dina(n9697),.dinb(w_asqrt22_19[1]),.dout(n9698),.clk(gclk));
	jxor g09431(.dina(n9698),.dinb(w_n9242_0[0]),.dout(n9699),.clk(gclk));
	jnot g09432(.din(n9699),.dout(n9700),.clk(gclk));
	jor g09433(.dina(w_n9687_0[1]),.dinb(w_asqrt58_17[0]),.dout(n9701),.clk(gclk));
	jor g09434(.dina(n9701),.dinb(w_n9693_0[1]),.dout(n9702),.clk(gclk));
	jand g09435(.dina(w_n9702_0[1]),.dinb(w_n9700_0[1]),.dout(n9703),.clk(gclk));
	jor g09436(.dina(w_n9703_0[1]),.dinb(w_n9695_0[1]),.dout(n9704),.clk(gclk));
	jand g09437(.dina(w_n9704_0[2]),.dinb(w_asqrt59_17[0]),.dout(n9705),.clk(gclk));
	jor g09438(.dina(w_n9704_0[1]),.dinb(w_asqrt59_16[2]),.dout(n9706),.clk(gclk));
	jnot g09439(.din(w_n9248_0[0]),.dout(n9707),.clk(gclk));
	jnot g09440(.din(w_n9249_0[0]),.dout(n9708),.clk(gclk));
	jand g09441(.dina(w_asqrt22_19[0]),.dinb(w_n9245_0[0]),.dout(n9709),.clk(gclk));
	jand g09442(.dina(w_n9709_0[1]),.dinb(n9708),.dout(n9710),.clk(gclk));
	jor g09443(.dina(n9710),.dinb(n9707),.dout(n9711),.clk(gclk));
	jnot g09444(.din(w_n9250_0[0]),.dout(n9712),.clk(gclk));
	jand g09445(.dina(w_n9709_0[0]),.dinb(n9712),.dout(n9713),.clk(gclk));
	jnot g09446(.din(n9713),.dout(n9714),.clk(gclk));
	jand g09447(.dina(n9714),.dinb(n9711),.dout(n9715),.clk(gclk));
	jand g09448(.dina(w_n9715_0[1]),.dinb(n9706),.dout(n9716),.clk(gclk));
	jor g09449(.dina(w_n9716_0[1]),.dinb(w_n9705_0[1]),.dout(n9717),.clk(gclk));
	jand g09450(.dina(n9717),.dinb(w_asqrt60_17[0]),.dout(n9718),.clk(gclk));
	jor g09451(.dina(w_n9705_0[0]),.dinb(w_asqrt60_16[2]),.dout(n9719),.clk(gclk));
	jor g09452(.dina(n9719),.dinb(w_n9716_0[0]),.dout(n9720),.clk(gclk));
	jnot g09453(.din(w_n9256_0[0]),.dout(n9721),.clk(gclk));
	jnot g09454(.din(w_n9258_0[0]),.dout(n9722),.clk(gclk));
	jand g09455(.dina(w_asqrt22_18[2]),.dinb(w_n9252_0[0]),.dout(n9723),.clk(gclk));
	jand g09456(.dina(w_n9723_0[1]),.dinb(n9722),.dout(n9724),.clk(gclk));
	jor g09457(.dina(n9724),.dinb(n9721),.dout(n9725),.clk(gclk));
	jnot g09458(.din(w_n9259_0[0]),.dout(n9726),.clk(gclk));
	jand g09459(.dina(w_n9723_0[0]),.dinb(n9726),.dout(n9727),.clk(gclk));
	jnot g09460(.din(n9727),.dout(n9728),.clk(gclk));
	jand g09461(.dina(n9728),.dinb(n9725),.dout(n9729),.clk(gclk));
	jand g09462(.dina(w_n9729_0[1]),.dinb(w_n9720_0[1]),.dout(n9730),.clk(gclk));
	jor g09463(.dina(n9730),.dinb(w_n9718_0[1]),.dout(n9731),.clk(gclk));
	jand g09464(.dina(w_n9731_0[1]),.dinb(w_asqrt61_17[1]),.dout(n9732),.clk(gclk));
	jxor g09465(.dina(w_n9260_0[0]),.dinb(w_n290_22[0]),.dout(n9733),.clk(gclk));
	jand g09466(.dina(n9733),.dinb(w_asqrt22_18[1]),.dout(n9734),.clk(gclk));
	jxor g09467(.dina(n9734),.dinb(w_n9270_0[0]),.dout(n9735),.clk(gclk));
	jnot g09468(.din(n9735),.dout(n9736),.clk(gclk));
	jor g09469(.dina(w_n9731_0[0]),.dinb(w_asqrt61_17[0]),.dout(n9737),.clk(gclk));
	jand g09470(.dina(w_n9737_0[1]),.dinb(w_n9736_0[1]),.dout(n9738),.clk(gclk));
	jor g09471(.dina(w_n9738_0[2]),.dinb(w_n9732_0[2]),.dout(n9739),.clk(gclk));
	jand g09472(.dina(n9739),.dinb(w_asqrt62_17[1]),.dout(n9740),.clk(gclk));
	jnot g09473(.din(w_n9275_0[0]),.dout(n9741),.clk(gclk));
	jand g09474(.dina(n9741),.dinb(w_n9273_0[0]),.dout(n9742),.clk(gclk));
	jand g09475(.dina(n9742),.dinb(w_asqrt22_18[0]),.dout(n9743),.clk(gclk));
	jxor g09476(.dina(n9743),.dinb(w_n9283_0[0]),.dout(n9744),.clk(gclk));
	jnot g09477(.din(n9744),.dout(n9745),.clk(gclk));
	jor g09478(.dina(w_n9732_0[1]),.dinb(w_asqrt62_17[0]),.dout(n9746),.clk(gclk));
	jor g09479(.dina(n9746),.dinb(w_n9738_0[1]),.dout(n9747),.clk(gclk));
	jand g09480(.dina(w_n9747_0[1]),.dinb(w_n9745_0[1]),.dout(n9748),.clk(gclk));
	jor g09481(.dina(w_n9748_0[1]),.dinb(w_n9740_0[1]),.dout(n9749),.clk(gclk));
	jxor g09482(.dina(w_n9285_0[0]),.dinb(w_n199_25[2]),.dout(n9750),.clk(gclk));
	jand g09483(.dina(n9750),.dinb(w_asqrt22_17[2]),.dout(n9751),.clk(gclk));
	jxor g09484(.dina(n9751),.dinb(w_n9290_0[0]),.dout(n9752),.clk(gclk));
	jnot g09485(.din(w_n9292_0[0]),.dout(n9753),.clk(gclk));
	jnot g09486(.din(w_n9296_0[0]),.dout(n9754),.clk(gclk));
	jand g09487(.dina(w_asqrt22_17[1]),.dinb(w_n9754_0[1]),.dout(n9755),.clk(gclk));
	jand g09488(.dina(w_n9755_0[1]),.dinb(w_n9753_0[2]),.dout(n9756),.clk(gclk));
	jor g09489(.dina(n9756),.dinb(w_n9303_0[0]),.dout(n9757),.clk(gclk));
	jor g09490(.dina(n9757),.dinb(w_n9752_0[1]),.dout(n9758),.clk(gclk));
	jnot g09491(.din(n9758),.dout(n9759),.clk(gclk));
	jand g09492(.dina(n9759),.dinb(w_n9749_1[2]),.dout(n9760),.clk(gclk));
	jor g09493(.dina(n9760),.dinb(w_asqrt63_9[1]),.dout(n9761),.clk(gclk));
	jnot g09494(.din(w_n9752_0[0]),.dout(n9762),.clk(gclk));
	jor g09495(.dina(w_n9762_0[2]),.dinb(w_n9749_1[1]),.dout(n9763),.clk(gclk));
	jor g09496(.dina(w_n9755_0[0]),.dinb(w_n9753_0[1]),.dout(n9764),.clk(gclk));
	jand g09497(.dina(w_n9754_0[0]),.dinb(w_n9753_0[0]),.dout(n9765),.clk(gclk));
	jor g09498(.dina(n9765),.dinb(w_n194_24[2]),.dout(n9766),.clk(gclk));
	jnot g09499(.din(n9766),.dout(n9767),.clk(gclk));
	jand g09500(.dina(n9767),.dinb(n9764),.dout(n9768),.clk(gclk));
	jnot g09501(.din(w_asqrt22_17[0]),.dout(n9769),.clk(gclk));
	jnot g09502(.din(w_n9768_0[1]),.dout(n9772),.clk(gclk));
	jand g09503(.dina(n9772),.dinb(w_n9763_0[1]),.dout(n9773),.clk(gclk));
	jand g09504(.dina(n9773),.dinb(w_n9761_0[1]),.dout(n9774),.clk(gclk));
	jxor g09505(.dina(w_n9506_0[0]),.dinb(w_n2875_20[0]),.dout(n9775),.clk(gclk));
	jor g09506(.dina(n9775),.dinb(w_n9774_25[2]),.dout(n9776),.clk(gclk));
	jxor g09507(.dina(n9776),.dinb(n9316),.dout(n9777),.clk(gclk));
	jnot g09508(.din(n9777),.dout(n9778),.clk(gclk));
	jor g09509(.dina(w_n9774_25[1]),.dinb(w_n9318_1[0]),.dout(n9779),.clk(gclk));
	jnot g09510(.din(w_a40_0[1]),.dout(n9780),.clk(gclk));
	jnot g09511(.din(a[41]),.dout(n9781),.clk(gclk));
	jand g09512(.dina(w_n9318_0[2]),.dinb(w_n9781_0[2]),.dout(n9782),.clk(gclk));
	jand g09513(.dina(n9782),.dinb(w_n9780_1[1]),.dout(n9783),.clk(gclk));
	jnot g09514(.din(n9783),.dout(n9784),.clk(gclk));
	jand g09515(.dina(n9784),.dinb(n9779),.dout(n9785),.clk(gclk));
	jor g09516(.dina(w_n9785_0[2]),.dinb(w_n9769_14[1]),.dout(n9786),.clk(gclk));
	jor g09517(.dina(w_n9774_25[0]),.dinb(w_a42_0[0]),.dout(n9787),.clk(gclk));
	jxor g09518(.dina(w_n9787_0[1]),.dinb(w_n9319_0[0]),.dout(n9788),.clk(gclk));
	jand g09519(.dina(w_n9785_0[1]),.dinb(w_n9769_14[0]),.dout(n9789),.clk(gclk));
	jor g09520(.dina(n9789),.dinb(w_n9788_0[1]),.dout(n9790),.clk(gclk));
	jand g09521(.dina(w_n9790_0[1]),.dinb(w_n9786_0[1]),.dout(n9791),.clk(gclk));
	jor g09522(.dina(n9791),.dinb(w_n8898_18[2]),.dout(n9792),.clk(gclk));
	jand g09523(.dina(w_n9786_0[0]),.dinb(w_n8898_18[1]),.dout(n9793),.clk(gclk));
	jand g09524(.dina(n9793),.dinb(w_n9790_0[0]),.dout(n9794),.clk(gclk));
	jor g09525(.dina(w_n9787_0[0]),.dinb(w_a43_0[0]),.dout(n9795),.clk(gclk));
	jnot g09526(.din(w_n9761_0[0]),.dout(n9796),.clk(gclk));
	jnot g09527(.din(w_n9763_0[0]),.dout(n9797),.clk(gclk));
	jor g09528(.dina(w_n9768_0[0]),.dinb(w_n9769_13[2]),.dout(n9798),.clk(gclk));
	jor g09529(.dina(n9798),.dinb(w_n9797_0[1]),.dout(n9799),.clk(gclk));
	jor g09530(.dina(n9799),.dinb(n9796),.dout(n9800),.clk(gclk));
	jand g09531(.dina(n9800),.dinb(n9795),.dout(n9801),.clk(gclk));
	jxor g09532(.dina(n9801),.dinb(w_n8903_0[1]),.dout(n9802),.clk(gclk));
	jor g09533(.dina(w_n9802_0[1]),.dinb(w_n9794_0[1]),.dout(n9803),.clk(gclk));
	jand g09534(.dina(n9803),.dinb(w_n9792_0[1]),.dout(n9804),.clk(gclk));
	jor g09535(.dina(w_n9804_0[2]),.dinb(w_n8893_14[1]),.dout(n9805),.clk(gclk));
	jand g09536(.dina(w_n9804_0[1]),.dinb(w_n8893_14[0]),.dout(n9806),.clk(gclk));
	jxor g09537(.dina(w_n9322_0[0]),.dinb(w_n8898_18[0]),.dout(n9807),.clk(gclk));
	jor g09538(.dina(n9807),.dinb(w_n9774_24[2]),.dout(n9808),.clk(gclk));
	jxor g09539(.dina(n9808),.dinb(w_n9325_0[0]),.dout(n9809),.clk(gclk));
	jor g09540(.dina(w_n9809_0[1]),.dinb(n9806),.dout(n9810),.clk(gclk));
	jand g09541(.dina(w_n9810_0[1]),.dinb(w_n9805_0[1]),.dout(n9811),.clk(gclk));
	jor g09542(.dina(n9811),.dinb(w_n8058_18[1]),.dout(n9812),.clk(gclk));
	jnot g09543(.din(w_n9331_0[0]),.dout(n9813),.clk(gclk));
	jor g09544(.dina(n9813),.dinb(w_n9329_0[0]),.dout(n9814),.clk(gclk));
	jor g09545(.dina(n9814),.dinb(w_n9774_24[1]),.dout(n9815),.clk(gclk));
	jxor g09546(.dina(n9815),.dinb(w_n9340_0[0]),.dout(n9816),.clk(gclk));
	jand g09547(.dina(w_n9805_0[0]),.dinb(w_n8058_18[0]),.dout(n9817),.clk(gclk));
	jand g09548(.dina(n9817),.dinb(w_n9810_0[0]),.dout(n9818),.clk(gclk));
	jor g09549(.dina(w_n9818_0[1]),.dinb(w_n9816_0[1]),.dout(n9819),.clk(gclk));
	jand g09550(.dina(w_n9819_0[1]),.dinb(w_n9812_0[1]),.dout(n9820),.clk(gclk));
	jor g09551(.dina(w_n9820_0[2]),.dinb(w_n8053_14[1]),.dout(n9821),.clk(gclk));
	jand g09552(.dina(w_n9820_0[1]),.dinb(w_n8053_14[0]),.dout(n9822),.clk(gclk));
	jxor g09553(.dina(w_n9342_0[0]),.dinb(w_n8058_17[2]),.dout(n9823),.clk(gclk));
	jor g09554(.dina(n9823),.dinb(w_n9774_24[0]),.dout(n9824),.clk(gclk));
	jxor g09555(.dina(n9824),.dinb(w_n9347_0[0]),.dout(n9825),.clk(gclk));
	jnot g09556(.din(w_n9825_0[1]),.dout(n9826),.clk(gclk));
	jor g09557(.dina(n9826),.dinb(n9822),.dout(n9827),.clk(gclk));
	jand g09558(.dina(w_n9827_0[1]),.dinb(w_n9821_0[1]),.dout(n9828),.clk(gclk));
	jor g09559(.dina(n9828),.dinb(w_n7265_18[2]),.dout(n9829),.clk(gclk));
	jand g09560(.dina(w_n9821_0[0]),.dinb(w_n7265_18[1]),.dout(n9830),.clk(gclk));
	jand g09561(.dina(n9830),.dinb(w_n9827_0[0]),.dout(n9831),.clk(gclk));
	jnot g09562(.din(w_n9351_0[0]),.dout(n9832),.clk(gclk));
	jnot g09563(.din(w_n9774_23[2]),.dout(asqrt_fa_22),.clk(gclk));
	jand g09564(.dina(w_asqrt21_19),.dinb(n9832),.dout(n9834),.clk(gclk));
	jand g09565(.dina(w_n9834_0[1]),.dinb(w_n9358_0[0]),.dout(n9835),.clk(gclk));
	jor g09566(.dina(n9835),.dinb(w_n9356_0[0]),.dout(n9836),.clk(gclk));
	jand g09567(.dina(w_n9834_0[0]),.dinb(w_n9359_0[0]),.dout(n9837),.clk(gclk));
	jnot g09568(.din(n9837),.dout(n9838),.clk(gclk));
	jand g09569(.dina(n9838),.dinb(n9836),.dout(n9839),.clk(gclk));
	jnot g09570(.din(n9839),.dout(n9840),.clk(gclk));
	jor g09571(.dina(w_n9840_0[1]),.dinb(w_n9831_0[1]),.dout(n9841),.clk(gclk));
	jand g09572(.dina(n9841),.dinb(w_n9829_0[1]),.dout(n9842),.clk(gclk));
	jor g09573(.dina(w_n9842_0[2]),.dinb(w_n7260_15[0]),.dout(n9843),.clk(gclk));
	jand g09574(.dina(w_n9842_0[1]),.dinb(w_n7260_14[2]),.dout(n9844),.clk(gclk));
	jnot g09575(.din(w_n9366_0[0]),.dout(n9845),.clk(gclk));
	jxor g09576(.dina(w_n9360_0[0]),.dinb(w_n7265_18[0]),.dout(n9846),.clk(gclk));
	jor g09577(.dina(n9846),.dinb(w_n9774_23[1]),.dout(n9847),.clk(gclk));
	jxor g09578(.dina(n9847),.dinb(n9845),.dout(n9848),.clk(gclk));
	jnot g09579(.din(w_n9848_0[1]),.dout(n9849),.clk(gclk));
	jor g09580(.dina(n9849),.dinb(n9844),.dout(n9850),.clk(gclk));
	jand g09581(.dina(w_n9850_0[1]),.dinb(w_n9843_0[1]),.dout(n9851),.clk(gclk));
	jor g09582(.dina(n9851),.dinb(w_n6505_18[1]),.dout(n9852),.clk(gclk));
	jnot g09583(.din(w_n9371_0[0]),.dout(n9853),.clk(gclk));
	jor g09584(.dina(n9853),.dinb(w_n9369_0[0]),.dout(n9854),.clk(gclk));
	jor g09585(.dina(n9854),.dinb(w_n9774_23[0]),.dout(n9855),.clk(gclk));
	jxor g09586(.dina(n9855),.dinb(w_n9380_0[0]),.dout(n9856),.clk(gclk));
	jand g09587(.dina(w_n9843_0[0]),.dinb(w_n6505_18[0]),.dout(n9857),.clk(gclk));
	jand g09588(.dina(n9857),.dinb(w_n9850_0[0]),.dout(n9858),.clk(gclk));
	jor g09589(.dina(w_n9858_0[1]),.dinb(w_n9856_0[1]),.dout(n9859),.clk(gclk));
	jand g09590(.dina(w_n9859_0[1]),.dinb(w_n9852_0[1]),.dout(n9860),.clk(gclk));
	jor g09591(.dina(w_n9860_0[2]),.dinb(w_n6500_15[0]),.dout(n9861),.clk(gclk));
	jand g09592(.dina(w_n9860_0[1]),.dinb(w_n6500_14[2]),.dout(n9862),.clk(gclk));
	jnot g09593(.din(w_n9387_0[0]),.dout(n9863),.clk(gclk));
	jxor g09594(.dina(w_n9382_0[0]),.dinb(w_n6505_17[2]),.dout(n9864),.clk(gclk));
	jor g09595(.dina(n9864),.dinb(w_n9774_22[2]),.dout(n9865),.clk(gclk));
	jxor g09596(.dina(n9865),.dinb(n9863),.dout(n9866),.clk(gclk));
	jnot g09597(.din(n9866),.dout(n9867),.clk(gclk));
	jor g09598(.dina(w_n9867_0[1]),.dinb(n9862),.dout(n9868),.clk(gclk));
	jand g09599(.dina(w_n9868_0[1]),.dinb(w_n9861_0[1]),.dout(n9869),.clk(gclk));
	jor g09600(.dina(n9869),.dinb(w_n5793_18[2]),.dout(n9870),.clk(gclk));
	jand g09601(.dina(w_n9861_0[0]),.dinb(w_n5793_18[1]),.dout(n9871),.clk(gclk));
	jand g09602(.dina(n9871),.dinb(w_n9868_0[0]),.dout(n9872),.clk(gclk));
	jnot g09603(.din(w_n9390_0[0]),.dout(n9873),.clk(gclk));
	jand g09604(.dina(w_asqrt21_18[2]),.dinb(n9873),.dout(n9874),.clk(gclk));
	jand g09605(.dina(w_n9874_0[1]),.dinb(w_n9397_0[0]),.dout(n9875),.clk(gclk));
	jor g09606(.dina(n9875),.dinb(w_n9395_0[0]),.dout(n9876),.clk(gclk));
	jand g09607(.dina(w_n9874_0[0]),.dinb(w_n9398_0[0]),.dout(n9877),.clk(gclk));
	jnot g09608(.din(n9877),.dout(n9878),.clk(gclk));
	jand g09609(.dina(n9878),.dinb(n9876),.dout(n9879),.clk(gclk));
	jnot g09610(.din(n9879),.dout(n9880),.clk(gclk));
	jor g09611(.dina(w_n9880_0[1]),.dinb(w_n9872_0[1]),.dout(n9881),.clk(gclk));
	jand g09612(.dina(n9881),.dinb(w_n9870_0[1]),.dout(n9882),.clk(gclk));
	jor g09613(.dina(w_n9882_0[1]),.dinb(w_n5788_15[1]),.dout(n9883),.clk(gclk));
	jxor g09614(.dina(w_n9399_0[0]),.dinb(w_n5793_18[0]),.dout(n9884),.clk(gclk));
	jor g09615(.dina(n9884),.dinb(w_n9774_22[1]),.dout(n9885),.clk(gclk));
	jxor g09616(.dina(n9885),.dinb(w_n9404_0[0]),.dout(n9886),.clk(gclk));
	jand g09617(.dina(w_n9882_0[0]),.dinb(w_n5788_15[0]),.dout(n9887),.clk(gclk));
	jor g09618(.dina(w_n9887_0[1]),.dinb(w_n9886_0[1]),.dout(n9888),.clk(gclk));
	jand g09619(.dina(w_n9888_0[2]),.dinb(w_n9883_0[2]),.dout(n9889),.clk(gclk));
	jor g09620(.dina(n9889),.dinb(w_n5121_18[1]),.dout(n9890),.clk(gclk));
	jnot g09621(.din(w_n9409_0[0]),.dout(n9891),.clk(gclk));
	jor g09622(.dina(n9891),.dinb(w_n9407_0[0]),.dout(n9892),.clk(gclk));
	jor g09623(.dina(n9892),.dinb(w_n9774_22[0]),.dout(n9893),.clk(gclk));
	jxor g09624(.dina(n9893),.dinb(w_n9418_0[0]),.dout(n9894),.clk(gclk));
	jand g09625(.dina(w_n9883_0[1]),.dinb(w_n5121_18[0]),.dout(n9895),.clk(gclk));
	jand g09626(.dina(n9895),.dinb(w_n9888_0[1]),.dout(n9896),.clk(gclk));
	jor g09627(.dina(w_n9896_0[1]),.dinb(w_n9894_0[1]),.dout(n9897),.clk(gclk));
	jand g09628(.dina(w_n9897_0[1]),.dinb(w_n9890_0[1]),.dout(n9898),.clk(gclk));
	jor g09629(.dina(w_n9898_0[2]),.dinb(w_n5116_15[2]),.dout(n9899),.clk(gclk));
	jand g09630(.dina(w_n9898_0[1]),.dinb(w_n5116_15[1]),.dout(n9900),.clk(gclk));
	jnot g09631(.din(w_n9421_0[0]),.dout(n9901),.clk(gclk));
	jand g09632(.dina(w_asqrt21_18[1]),.dinb(n9901),.dout(n9902),.clk(gclk));
	jand g09633(.dina(w_n9902_0[1]),.dinb(w_n9426_0[0]),.dout(n9903),.clk(gclk));
	jor g09634(.dina(n9903),.dinb(w_n9425_0[0]),.dout(n9904),.clk(gclk));
	jand g09635(.dina(w_n9902_0[0]),.dinb(w_n9427_0[0]),.dout(n9905),.clk(gclk));
	jnot g09636(.din(n9905),.dout(n9906),.clk(gclk));
	jand g09637(.dina(n9906),.dinb(n9904),.dout(n9907),.clk(gclk));
	jnot g09638(.din(n9907),.dout(n9908),.clk(gclk));
	jor g09639(.dina(w_n9908_0[1]),.dinb(n9900),.dout(n9909),.clk(gclk));
	jand g09640(.dina(w_n9909_0[1]),.dinb(w_n9899_0[1]),.dout(n9910),.clk(gclk));
	jor g09641(.dina(n9910),.dinb(w_n4499_19[1]),.dout(n9911),.clk(gclk));
	jand g09642(.dina(w_n9899_0[0]),.dinb(w_n4499_19[0]),.dout(n9912),.clk(gclk));
	jand g09643(.dina(n9912),.dinb(w_n9909_0[0]),.dout(n9913),.clk(gclk));
	jnot g09644(.din(w_n9429_0[0]),.dout(n9914),.clk(gclk));
	jand g09645(.dina(w_asqrt21_18[0]),.dinb(n9914),.dout(n9915),.clk(gclk));
	jand g09646(.dina(w_n9915_0[1]),.dinb(w_n9436_0[0]),.dout(n9916),.clk(gclk));
	jor g09647(.dina(n9916),.dinb(w_n9434_0[0]),.dout(n9917),.clk(gclk));
	jand g09648(.dina(w_n9915_0[0]),.dinb(w_n9437_0[0]),.dout(n9918),.clk(gclk));
	jnot g09649(.din(n9918),.dout(n9919),.clk(gclk));
	jand g09650(.dina(n9919),.dinb(n9917),.dout(n9920),.clk(gclk));
	jnot g09651(.din(n9920),.dout(n9921),.clk(gclk));
	jor g09652(.dina(w_n9921_0[1]),.dinb(w_n9913_0[1]),.dout(n9922),.clk(gclk));
	jand g09653(.dina(n9922),.dinb(w_n9911_0[1]),.dout(n9923),.clk(gclk));
	jor g09654(.dina(w_n9923_0[1]),.dinb(w_n4494_16[1]),.dout(n9924),.clk(gclk));
	jxor g09655(.dina(w_n9438_0[0]),.dinb(w_n4499_18[2]),.dout(n9925),.clk(gclk));
	jor g09656(.dina(n9925),.dinb(w_n9774_21[2]),.dout(n9926),.clk(gclk));
	jxor g09657(.dina(n9926),.dinb(w_n9449_0[0]),.dout(n9927),.clk(gclk));
	jand g09658(.dina(w_n9923_0[0]),.dinb(w_n4494_16[0]),.dout(n9928),.clk(gclk));
	jor g09659(.dina(w_n9928_0[1]),.dinb(w_n9927_0[1]),.dout(n9929),.clk(gclk));
	jand g09660(.dina(w_n9929_0[2]),.dinb(w_n9924_0[2]),.dout(n9930),.clk(gclk));
	jor g09661(.dina(n9930),.dinb(w_n3912_19[0]),.dout(n9931),.clk(gclk));
	jnot g09662(.din(w_n9454_0[0]),.dout(n9932),.clk(gclk));
	jor g09663(.dina(n9932),.dinb(w_n9452_0[0]),.dout(n9933),.clk(gclk));
	jor g09664(.dina(n9933),.dinb(w_n9774_21[1]),.dout(n9934),.clk(gclk));
	jxor g09665(.dina(n9934),.dinb(w_n9463_0[0]),.dout(n9935),.clk(gclk));
	jand g09666(.dina(w_n9924_0[1]),.dinb(w_n3912_18[2]),.dout(n9936),.clk(gclk));
	jand g09667(.dina(n9936),.dinb(w_n9929_0[1]),.dout(n9937),.clk(gclk));
	jor g09668(.dina(w_n9937_0[1]),.dinb(w_n9935_0[1]),.dout(n9938),.clk(gclk));
	jand g09669(.dina(w_n9938_0[1]),.dinb(w_n9931_0[1]),.dout(n9939),.clk(gclk));
	jor g09670(.dina(w_n9939_0[2]),.dinb(w_n3907_16[2]),.dout(n9940),.clk(gclk));
	jand g09671(.dina(w_n9939_0[1]),.dinb(w_n3907_16[1]),.dout(n9941),.clk(gclk));
	jnot g09672(.din(w_n9466_0[0]),.dout(n9942),.clk(gclk));
	jand g09673(.dina(w_asqrt21_17[2]),.dinb(n9942),.dout(n9943),.clk(gclk));
	jand g09674(.dina(w_n9943_0[1]),.dinb(w_n9471_0[0]),.dout(n9944),.clk(gclk));
	jor g09675(.dina(n9944),.dinb(w_n9470_0[0]),.dout(n9945),.clk(gclk));
	jand g09676(.dina(w_n9943_0[0]),.dinb(w_n9472_0[0]),.dout(n9946),.clk(gclk));
	jnot g09677(.din(n9946),.dout(n9947),.clk(gclk));
	jand g09678(.dina(n9947),.dinb(n9945),.dout(n9948),.clk(gclk));
	jnot g09679(.din(n9948),.dout(n9949),.clk(gclk));
	jor g09680(.dina(w_n9949_0[1]),.dinb(n9941),.dout(n9950),.clk(gclk));
	jand g09681(.dina(w_n9950_0[1]),.dinb(w_n9940_0[1]),.dout(n9951),.clk(gclk));
	jor g09682(.dina(n9951),.dinb(w_n3376_20[0]),.dout(n9952),.clk(gclk));
	jand g09683(.dina(w_n9940_0[0]),.dinb(w_n3376_19[2]),.dout(n9953),.clk(gclk));
	jand g09684(.dina(n9953),.dinb(w_n9950_0[0]),.dout(n9954),.clk(gclk));
	jnot g09685(.din(w_n9474_0[0]),.dout(n9955),.clk(gclk));
	jand g09686(.dina(w_asqrt21_17[1]),.dinb(n9955),.dout(n9956),.clk(gclk));
	jand g09687(.dina(w_n9956_0[1]),.dinb(w_n9481_0[0]),.dout(n9957),.clk(gclk));
	jor g09688(.dina(n9957),.dinb(w_n9479_0[0]),.dout(n9958),.clk(gclk));
	jand g09689(.dina(w_n9956_0[0]),.dinb(w_n9482_0[0]),.dout(n9959),.clk(gclk));
	jnot g09690(.din(n9959),.dout(n9960),.clk(gclk));
	jand g09691(.dina(n9960),.dinb(n9958),.dout(n9961),.clk(gclk));
	jnot g09692(.din(n9961),.dout(n9962),.clk(gclk));
	jor g09693(.dina(w_n9962_0[1]),.dinb(w_n9954_0[1]),.dout(n9963),.clk(gclk));
	jand g09694(.dina(n9963),.dinb(w_n9952_0[1]),.dout(n9964),.clk(gclk));
	jor g09695(.dina(w_n9964_0[1]),.dinb(w_n3371_17[0]),.dout(n9965),.clk(gclk));
	jxor g09696(.dina(w_n9483_0[0]),.dinb(w_n3376_19[1]),.dout(n9966),.clk(gclk));
	jor g09697(.dina(n9966),.dinb(w_n9774_21[0]),.dout(n9967),.clk(gclk));
	jxor g09698(.dina(n9967),.dinb(w_n9494_0[0]),.dout(n9968),.clk(gclk));
	jand g09699(.dina(w_n9964_0[0]),.dinb(w_n3371_16[2]),.dout(n9969),.clk(gclk));
	jor g09700(.dina(w_n9969_0[1]),.dinb(w_n9968_0[1]),.dout(n9970),.clk(gclk));
	jand g09701(.dina(w_n9970_0[2]),.dinb(w_n9965_0[2]),.dout(n9971),.clk(gclk));
	jor g09702(.dina(n9971),.dinb(w_n2875_19[2]),.dout(n9972),.clk(gclk));
	jand g09703(.dina(w_n9965_0[1]),.dinb(w_n2875_19[1]),.dout(n9973),.clk(gclk));
	jand g09704(.dina(n9973),.dinb(w_n9970_0[1]),.dout(n9974),.clk(gclk));
	jnot g09705(.din(w_n9497_0[0]),.dout(n9975),.clk(gclk));
	jand g09706(.dina(w_asqrt21_17[0]),.dinb(n9975),.dout(n9976),.clk(gclk));
	jand g09707(.dina(w_n9976_0[1]),.dinb(w_n9504_0[0]),.dout(n9977),.clk(gclk));
	jor g09708(.dina(n9977),.dinb(w_n9502_0[0]),.dout(n9978),.clk(gclk));
	jand g09709(.dina(w_n9976_0[0]),.dinb(w_n9505_0[0]),.dout(n9979),.clk(gclk));
	jnot g09710(.din(n9979),.dout(n9980),.clk(gclk));
	jand g09711(.dina(n9980),.dinb(n9978),.dout(n9981),.clk(gclk));
	jnot g09712(.din(n9981),.dout(n9982),.clk(gclk));
	jor g09713(.dina(w_n9982_0[1]),.dinb(w_n9974_0[1]),.dout(n9983),.clk(gclk));
	jand g09714(.dina(n9983),.dinb(w_n9972_0[1]),.dout(n9984),.clk(gclk));
	jor g09715(.dina(w_n9984_0[2]),.dinb(w_n2870_17[1]),.dout(n9985),.clk(gclk));
	jand g09716(.dina(w_n9984_0[1]),.dinb(w_n2870_17[0]),.dout(n9986),.clk(gclk));
	jor g09717(.dina(n9986),.dinb(w_n9778_0[1]),.dout(n9987),.clk(gclk));
	jand g09718(.dina(w_n9987_0[1]),.dinb(w_n9985_0[1]),.dout(n9988),.clk(gclk));
	jor g09719(.dina(n9988),.dinb(w_n2425_20[2]),.dout(n9989),.clk(gclk));
	jnot g09720(.din(w_n9513_0[0]),.dout(n9990),.clk(gclk));
	jor g09721(.dina(n9990),.dinb(w_n9511_0[0]),.dout(n9991),.clk(gclk));
	jor g09722(.dina(n9991),.dinb(w_n9774_20[2]),.dout(n9992),.clk(gclk));
	jxor g09723(.dina(n9992),.dinb(w_n9522_0[0]),.dout(n9993),.clk(gclk));
	jand g09724(.dina(w_n9985_0[0]),.dinb(w_n2425_20[1]),.dout(n9994),.clk(gclk));
	jand g09725(.dina(n9994),.dinb(w_n9987_0[0]),.dout(n9995),.clk(gclk));
	jor g09726(.dina(w_n9995_0[1]),.dinb(w_n9993_0[1]),.dout(n9996),.clk(gclk));
	jand g09727(.dina(w_n9996_0[1]),.dinb(w_n9989_0[1]),.dout(n9997),.clk(gclk));
	jor g09728(.dina(w_n9997_0[1]),.dinb(w_n2420_18[0]),.dout(n9998),.clk(gclk));
	jxor g09729(.dina(w_n9524_0[0]),.dinb(w_n2425_20[0]),.dout(n9999),.clk(gclk));
	jor g09730(.dina(n9999),.dinb(w_n9774_20[1]),.dout(n10000),.clk(gclk));
	jxor g09731(.dina(n10000),.dinb(w_n9535_0[0]),.dout(n10001),.clk(gclk));
	jand g09732(.dina(w_n9997_0[0]),.dinb(w_n2420_17[2]),.dout(n10002),.clk(gclk));
	jor g09733(.dina(w_n10002_0[1]),.dinb(w_n10001_0[1]),.dout(n10003),.clk(gclk));
	jand g09734(.dina(w_n10003_0[2]),.dinb(w_n9998_0[2]),.dout(n10004),.clk(gclk));
	jor g09735(.dina(n10004),.dinb(w_n2010_20[1]),.dout(n10005),.clk(gclk));
	jnot g09736(.din(w_n9540_0[0]),.dout(n10006),.clk(gclk));
	jor g09737(.dina(n10006),.dinb(w_n9538_0[0]),.dout(n10007),.clk(gclk));
	jor g09738(.dina(n10007),.dinb(w_n9774_20[0]),.dout(n10008),.clk(gclk));
	jxor g09739(.dina(n10008),.dinb(w_n9549_0[0]),.dout(n10009),.clk(gclk));
	jand g09740(.dina(w_n9998_0[1]),.dinb(w_n2010_20[0]),.dout(n10010),.clk(gclk));
	jand g09741(.dina(n10010),.dinb(w_n10003_0[1]),.dout(n10011),.clk(gclk));
	jor g09742(.dina(w_n10011_0[1]),.dinb(w_n10009_0[1]),.dout(n10012),.clk(gclk));
	jand g09743(.dina(w_n10012_0[1]),.dinb(w_n10005_0[1]),.dout(n10013),.clk(gclk));
	jor g09744(.dina(w_n10013_0[2]),.dinb(w_n2005_18[1]),.dout(n10014),.clk(gclk));
	jand g09745(.dina(w_n10013_0[1]),.dinb(w_n2005_18[0]),.dout(n10015),.clk(gclk));
	jnot g09746(.din(w_n9552_0[0]),.dout(n10016),.clk(gclk));
	jand g09747(.dina(w_asqrt21_16[2]),.dinb(n10016),.dout(n10017),.clk(gclk));
	jand g09748(.dina(w_n10017_0[1]),.dinb(w_n9557_0[0]),.dout(n10018),.clk(gclk));
	jor g09749(.dina(n10018),.dinb(w_n9556_0[0]),.dout(n10019),.clk(gclk));
	jand g09750(.dina(w_n10017_0[0]),.dinb(w_n9558_0[0]),.dout(n10020),.clk(gclk));
	jnot g09751(.din(n10020),.dout(n10021),.clk(gclk));
	jand g09752(.dina(n10021),.dinb(n10019),.dout(n10022),.clk(gclk));
	jnot g09753(.din(n10022),.dout(n10023),.clk(gclk));
	jor g09754(.dina(w_n10023_0[1]),.dinb(n10015),.dout(n10024),.clk(gclk));
	jand g09755(.dina(w_n10024_0[1]),.dinb(w_n10014_0[1]),.dout(n10025),.clk(gclk));
	jor g09756(.dina(n10025),.dinb(w_n1646_21[1]),.dout(n10026),.clk(gclk));
	jand g09757(.dina(w_n10014_0[0]),.dinb(w_n1646_21[0]),.dout(n10027),.clk(gclk));
	jand g09758(.dina(n10027),.dinb(w_n10024_0[0]),.dout(n10028),.clk(gclk));
	jnot g09759(.din(w_n9560_0[0]),.dout(n10029),.clk(gclk));
	jand g09760(.dina(w_asqrt21_16[1]),.dinb(n10029),.dout(n10030),.clk(gclk));
	jand g09761(.dina(w_n10030_0[1]),.dinb(w_n9567_0[0]),.dout(n10031),.clk(gclk));
	jor g09762(.dina(n10031),.dinb(w_n9565_0[0]),.dout(n10032),.clk(gclk));
	jand g09763(.dina(w_n10030_0[0]),.dinb(w_n9568_0[0]),.dout(n10033),.clk(gclk));
	jnot g09764(.din(n10033),.dout(n10034),.clk(gclk));
	jand g09765(.dina(n10034),.dinb(n10032),.dout(n10035),.clk(gclk));
	jnot g09766(.din(n10035),.dout(n10036),.clk(gclk));
	jor g09767(.dina(w_n10036_0[1]),.dinb(w_n10028_0[1]),.dout(n10037),.clk(gclk));
	jand g09768(.dina(n10037),.dinb(w_n10026_0[1]),.dout(n10038),.clk(gclk));
	jor g09769(.dina(w_n10038_0[1]),.dinb(w_n1641_18[2]),.dout(n10039),.clk(gclk));
	jxor g09770(.dina(w_n9569_0[0]),.dinb(w_n1646_20[2]),.dout(n10040),.clk(gclk));
	jor g09771(.dina(n10040),.dinb(w_n9774_19[2]),.dout(n10041),.clk(gclk));
	jxor g09772(.dina(n10041),.dinb(w_n9580_0[0]),.dout(n10042),.clk(gclk));
	jand g09773(.dina(w_n10038_0[0]),.dinb(w_n1641_18[1]),.dout(n10043),.clk(gclk));
	jor g09774(.dina(w_n10043_0[1]),.dinb(w_n10042_0[1]),.dout(n10044),.clk(gclk));
	jand g09775(.dina(w_n10044_0[2]),.dinb(w_n10039_0[2]),.dout(n10045),.clk(gclk));
	jor g09776(.dina(n10045),.dinb(w_n1317_21[0]),.dout(n10046),.clk(gclk));
	jnot g09777(.din(w_n9585_0[0]),.dout(n10047),.clk(gclk));
	jor g09778(.dina(n10047),.dinb(w_n9583_0[0]),.dout(n10048),.clk(gclk));
	jor g09779(.dina(n10048),.dinb(w_n9774_19[1]),.dout(n10049),.clk(gclk));
	jxor g09780(.dina(n10049),.dinb(w_n9594_0[0]),.dout(n10050),.clk(gclk));
	jand g09781(.dina(w_n10039_0[1]),.dinb(w_n1317_20[2]),.dout(n10051),.clk(gclk));
	jand g09782(.dina(n10051),.dinb(w_n10044_0[1]),.dout(n10052),.clk(gclk));
	jor g09783(.dina(w_n10052_0[1]),.dinb(w_n10050_0[1]),.dout(n10053),.clk(gclk));
	jand g09784(.dina(w_n10053_0[1]),.dinb(w_n10046_0[1]),.dout(n10054),.clk(gclk));
	jor g09785(.dina(w_n10054_0[2]),.dinb(w_n1312_19[0]),.dout(n10055),.clk(gclk));
	jand g09786(.dina(w_n10054_0[1]),.dinb(w_n1312_18[2]),.dout(n10056),.clk(gclk));
	jnot g09787(.din(w_n9597_0[0]),.dout(n10057),.clk(gclk));
	jand g09788(.dina(w_asqrt21_16[0]),.dinb(n10057),.dout(n10058),.clk(gclk));
	jand g09789(.dina(w_n10058_0[1]),.dinb(w_n9602_0[0]),.dout(n10059),.clk(gclk));
	jor g09790(.dina(n10059),.dinb(w_n9601_0[0]),.dout(n10060),.clk(gclk));
	jand g09791(.dina(w_n10058_0[0]),.dinb(w_n9603_0[0]),.dout(n10061),.clk(gclk));
	jnot g09792(.din(n10061),.dout(n10062),.clk(gclk));
	jand g09793(.dina(n10062),.dinb(n10060),.dout(n10063),.clk(gclk));
	jnot g09794(.din(n10063),.dout(n10064),.clk(gclk));
	jor g09795(.dina(w_n10064_0[1]),.dinb(n10056),.dout(n10065),.clk(gclk));
	jand g09796(.dina(w_n10065_0[1]),.dinb(w_n10055_0[1]),.dout(n10066),.clk(gclk));
	jor g09797(.dina(n10066),.dinb(w_n1039_21[2]),.dout(n10067),.clk(gclk));
	jand g09798(.dina(w_n10055_0[0]),.dinb(w_n1039_21[1]),.dout(n10068),.clk(gclk));
	jand g09799(.dina(n10068),.dinb(w_n10065_0[0]),.dout(n10069),.clk(gclk));
	jnot g09800(.din(w_n9605_0[0]),.dout(n10070),.clk(gclk));
	jand g09801(.dina(w_asqrt21_15[2]),.dinb(n10070),.dout(n10071),.clk(gclk));
	jand g09802(.dina(w_n10071_0[1]),.dinb(w_n9612_0[0]),.dout(n10072),.clk(gclk));
	jor g09803(.dina(n10072),.dinb(w_n9610_0[0]),.dout(n10073),.clk(gclk));
	jand g09804(.dina(w_n10071_0[0]),.dinb(w_n9613_0[0]),.dout(n10074),.clk(gclk));
	jnot g09805(.din(n10074),.dout(n10075),.clk(gclk));
	jand g09806(.dina(n10075),.dinb(n10073),.dout(n10076),.clk(gclk));
	jnot g09807(.din(n10076),.dout(n10077),.clk(gclk));
	jor g09808(.dina(w_n10077_0[1]),.dinb(w_n10069_0[1]),.dout(n10078),.clk(gclk));
	jand g09809(.dina(n10078),.dinb(w_n10067_0[1]),.dout(n10079),.clk(gclk));
	jor g09810(.dina(w_n10079_0[1]),.dinb(w_n1034_19[2]),.dout(n10080),.clk(gclk));
	jxor g09811(.dina(w_n9614_0[0]),.dinb(w_n1039_21[0]),.dout(n10081),.clk(gclk));
	jor g09812(.dina(n10081),.dinb(w_n9774_19[0]),.dout(n10082),.clk(gclk));
	jxor g09813(.dina(n10082),.dinb(w_n9625_0[0]),.dout(n10083),.clk(gclk));
	jand g09814(.dina(w_n10079_0[0]),.dinb(w_n1034_19[1]),.dout(n10084),.clk(gclk));
	jor g09815(.dina(w_n10084_0[1]),.dinb(w_n10083_0[1]),.dout(n10085),.clk(gclk));
	jand g09816(.dina(w_n10085_0[2]),.dinb(w_n10080_0[2]),.dout(n10086),.clk(gclk));
	jor g09817(.dina(n10086),.dinb(w_n796_21[1]),.dout(n10087),.clk(gclk));
	jnot g09818(.din(w_n9630_0[0]),.dout(n10088),.clk(gclk));
	jor g09819(.dina(n10088),.dinb(w_n9628_0[0]),.dout(n10089),.clk(gclk));
	jor g09820(.dina(n10089),.dinb(w_n9774_18[2]),.dout(n10090),.clk(gclk));
	jxor g09821(.dina(n10090),.dinb(w_n9639_0[0]),.dout(n10091),.clk(gclk));
	jand g09822(.dina(w_n10080_0[1]),.dinb(w_n796_21[0]),.dout(n10092),.clk(gclk));
	jand g09823(.dina(n10092),.dinb(w_n10085_0[1]),.dout(n10093),.clk(gclk));
	jor g09824(.dina(w_n10093_0[1]),.dinb(w_n10091_0[1]),.dout(n10094),.clk(gclk));
	jand g09825(.dina(w_n10094_0[1]),.dinb(w_n10087_0[1]),.dout(n10095),.clk(gclk));
	jor g09826(.dina(w_n10095_0[2]),.dinb(w_n791_20[0]),.dout(n10096),.clk(gclk));
	jand g09827(.dina(w_n10095_0[1]),.dinb(w_n791_19[2]),.dout(n10097),.clk(gclk));
	jnot g09828(.din(w_n9642_0[0]),.dout(n10098),.clk(gclk));
	jand g09829(.dina(w_asqrt21_15[1]),.dinb(n10098),.dout(n10099),.clk(gclk));
	jand g09830(.dina(w_n10099_0[1]),.dinb(w_n9647_0[0]),.dout(n10100),.clk(gclk));
	jor g09831(.dina(n10100),.dinb(w_n9646_0[0]),.dout(n10101),.clk(gclk));
	jand g09832(.dina(w_n10099_0[0]),.dinb(w_n9648_0[0]),.dout(n10102),.clk(gclk));
	jnot g09833(.din(n10102),.dout(n10103),.clk(gclk));
	jand g09834(.dina(n10103),.dinb(n10101),.dout(n10104),.clk(gclk));
	jnot g09835(.din(n10104),.dout(n10105),.clk(gclk));
	jor g09836(.dina(w_n10105_0[1]),.dinb(n10097),.dout(n10106),.clk(gclk));
	jand g09837(.dina(w_n10106_0[1]),.dinb(w_n10096_0[1]),.dout(n10107),.clk(gclk));
	jor g09838(.dina(n10107),.dinb(w_n595_22[0]),.dout(n10108),.clk(gclk));
	jand g09839(.dina(w_n10096_0[0]),.dinb(w_n595_21[2]),.dout(n10109),.clk(gclk));
	jand g09840(.dina(n10109),.dinb(w_n10106_0[0]),.dout(n10110),.clk(gclk));
	jnot g09841(.din(w_n9650_0[0]),.dout(n10111),.clk(gclk));
	jand g09842(.dina(w_asqrt21_15[0]),.dinb(n10111),.dout(n10112),.clk(gclk));
	jand g09843(.dina(w_n10112_0[1]),.dinb(w_n9657_0[0]),.dout(n10113),.clk(gclk));
	jor g09844(.dina(n10113),.dinb(w_n9655_0[0]),.dout(n10114),.clk(gclk));
	jand g09845(.dina(w_n10112_0[0]),.dinb(w_n9658_0[0]),.dout(n10115),.clk(gclk));
	jnot g09846(.din(n10115),.dout(n10116),.clk(gclk));
	jand g09847(.dina(n10116),.dinb(n10114),.dout(n10117),.clk(gclk));
	jnot g09848(.din(n10117),.dout(n10118),.clk(gclk));
	jor g09849(.dina(w_n10118_0[1]),.dinb(w_n10110_0[1]),.dout(n10119),.clk(gclk));
	jand g09850(.dina(n10119),.dinb(w_n10108_0[1]),.dout(n10120),.clk(gclk));
	jor g09851(.dina(w_n10120_0[1]),.dinb(w_n590_20[1]),.dout(n10121),.clk(gclk));
	jxor g09852(.dina(w_n9659_0[0]),.dinb(w_n595_21[1]),.dout(n10122),.clk(gclk));
	jor g09853(.dina(n10122),.dinb(w_n9774_18[1]),.dout(n10123),.clk(gclk));
	jxor g09854(.dina(n10123),.dinb(w_n9670_0[0]),.dout(n10124),.clk(gclk));
	jand g09855(.dina(w_n10120_0[0]),.dinb(w_n590_20[0]),.dout(n10125),.clk(gclk));
	jor g09856(.dina(w_n10125_0[1]),.dinb(w_n10124_0[1]),.dout(n10126),.clk(gclk));
	jand g09857(.dina(w_n10126_0[2]),.dinb(w_n10121_0[2]),.dout(n10127),.clk(gclk));
	jor g09858(.dina(n10127),.dinb(w_n430_21[2]),.dout(n10128),.clk(gclk));
	jnot g09859(.din(w_n9675_0[0]),.dout(n10129),.clk(gclk));
	jor g09860(.dina(n10129),.dinb(w_n9673_0[0]),.dout(n10130),.clk(gclk));
	jor g09861(.dina(n10130),.dinb(w_n9774_18[0]),.dout(n10131),.clk(gclk));
	jxor g09862(.dina(n10131),.dinb(w_n9684_0[0]),.dout(n10132),.clk(gclk));
	jand g09863(.dina(w_n10121_0[1]),.dinb(w_n430_21[1]),.dout(n10133),.clk(gclk));
	jand g09864(.dina(n10133),.dinb(w_n10126_0[1]),.dout(n10134),.clk(gclk));
	jor g09865(.dina(w_n10134_0[1]),.dinb(w_n10132_0[1]),.dout(n10135),.clk(gclk));
	jand g09866(.dina(w_n10135_0[1]),.dinb(w_n10128_0[1]),.dout(n10136),.clk(gclk));
	jor g09867(.dina(w_n10136_0[2]),.dinb(w_n425_20[2]),.dout(n10137),.clk(gclk));
	jand g09868(.dina(w_n10136_0[1]),.dinb(w_n425_20[1]),.dout(n10138),.clk(gclk));
	jnot g09869(.din(w_n9687_0[0]),.dout(n10139),.clk(gclk));
	jand g09870(.dina(w_asqrt21_14[2]),.dinb(n10139),.dout(n10140),.clk(gclk));
	jand g09871(.dina(w_n10140_0[1]),.dinb(w_n9692_0[0]),.dout(n10141),.clk(gclk));
	jor g09872(.dina(n10141),.dinb(w_n9691_0[0]),.dout(n10142),.clk(gclk));
	jand g09873(.dina(w_n10140_0[0]),.dinb(w_n9693_0[0]),.dout(n10143),.clk(gclk));
	jnot g09874(.din(n10143),.dout(n10144),.clk(gclk));
	jand g09875(.dina(n10144),.dinb(n10142),.dout(n10145),.clk(gclk));
	jnot g09876(.din(n10145),.dout(n10146),.clk(gclk));
	jor g09877(.dina(w_n10146_0[1]),.dinb(n10138),.dout(n10147),.clk(gclk));
	jand g09878(.dina(w_n10147_0[1]),.dinb(w_n10137_0[1]),.dout(n10148),.clk(gclk));
	jor g09879(.dina(n10148),.dinb(w_n305_22[1]),.dout(n10149),.clk(gclk));
	jand g09880(.dina(w_n10137_0[0]),.dinb(w_n305_22[0]),.dout(n10150),.clk(gclk));
	jand g09881(.dina(n10150),.dinb(w_n10147_0[0]),.dout(n10151),.clk(gclk));
	jnot g09882(.din(w_n9695_0[0]),.dout(n10152),.clk(gclk));
	jand g09883(.dina(w_asqrt21_14[1]),.dinb(n10152),.dout(n10153),.clk(gclk));
	jand g09884(.dina(w_n10153_0[1]),.dinb(w_n9702_0[0]),.dout(n10154),.clk(gclk));
	jor g09885(.dina(n10154),.dinb(w_n9700_0[0]),.dout(n10155),.clk(gclk));
	jand g09886(.dina(w_n10153_0[0]),.dinb(w_n9703_0[0]),.dout(n10156),.clk(gclk));
	jnot g09887(.din(n10156),.dout(n10157),.clk(gclk));
	jand g09888(.dina(n10157),.dinb(n10155),.dout(n10158),.clk(gclk));
	jnot g09889(.din(n10158),.dout(n10159),.clk(gclk));
	jor g09890(.dina(w_n10159_0[1]),.dinb(w_n10151_0[1]),.dout(n10160),.clk(gclk));
	jand g09891(.dina(n10160),.dinb(w_n10149_0[1]),.dout(n10161),.clk(gclk));
	jor g09892(.dina(w_n10161_0[1]),.dinb(w_n290_21[2]),.dout(n10162),.clk(gclk));
	jxor g09893(.dina(w_n9704_0[0]),.dinb(w_n305_21[2]),.dout(n10163),.clk(gclk));
	jor g09894(.dina(n10163),.dinb(w_n9774_17[2]),.dout(n10164),.clk(gclk));
	jxor g09895(.dina(n10164),.dinb(w_n9715_0[0]),.dout(n10165),.clk(gclk));
	jand g09896(.dina(w_n10161_0[0]),.dinb(w_n290_21[1]),.dout(n10166),.clk(gclk));
	jor g09897(.dina(w_n10166_0[1]),.dinb(w_n10165_0[1]),.dout(n10167),.clk(gclk));
	jand g09898(.dina(w_n10167_0[2]),.dinb(w_n10162_0[2]),.dout(n10168),.clk(gclk));
	jor g09899(.dina(n10168),.dinb(w_n223_22[0]),.dout(n10169),.clk(gclk));
	jnot g09900(.din(w_n9720_0[0]),.dout(n10170),.clk(gclk));
	jor g09901(.dina(n10170),.dinb(w_n9718_0[0]),.dout(n10171),.clk(gclk));
	jor g09902(.dina(n10171),.dinb(w_n9774_17[1]),.dout(n10172),.clk(gclk));
	jxor g09903(.dina(n10172),.dinb(w_n9729_0[0]),.dout(n10173),.clk(gclk));
	jand g09904(.dina(w_n10162_0[1]),.dinb(w_n223_21[2]),.dout(n10174),.clk(gclk));
	jand g09905(.dina(n10174),.dinb(w_n10167_0[1]),.dout(n10175),.clk(gclk));
	jor g09906(.dina(w_n10175_0[1]),.dinb(w_n10173_0[1]),.dout(n10176),.clk(gclk));
	jand g09907(.dina(w_n10176_0[1]),.dinb(w_n10169_0[1]),.dout(n10177),.clk(gclk));
	jor g09908(.dina(w_n10177_0[2]),.dinb(w_n199_25[1]),.dout(n10178),.clk(gclk));
	jand g09909(.dina(w_n10177_0[1]),.dinb(w_n199_25[0]),.dout(n10179),.clk(gclk));
	jnot g09910(.din(w_n9732_0[0]),.dout(n10180),.clk(gclk));
	jand g09911(.dina(w_asqrt21_14[0]),.dinb(n10180),.dout(n10181),.clk(gclk));
	jand g09912(.dina(w_n10181_0[1]),.dinb(w_n9737_0[0]),.dout(n10182),.clk(gclk));
	jor g09913(.dina(n10182),.dinb(w_n9736_0[0]),.dout(n10183),.clk(gclk));
	jand g09914(.dina(w_n10181_0[0]),.dinb(w_n9738_0[0]),.dout(n10184),.clk(gclk));
	jnot g09915(.din(n10184),.dout(n10185),.clk(gclk));
	jand g09916(.dina(n10185),.dinb(n10183),.dout(n10186),.clk(gclk));
	jnot g09917(.din(n10186),.dout(n10187),.clk(gclk));
	jor g09918(.dina(w_n10187_0[1]),.dinb(n10179),.dout(n10188),.clk(gclk));
	jand g09919(.dina(n10188),.dinb(n10178),.dout(n10189),.clk(gclk));
	jnot g09920(.din(w_n9740_0[0]),.dout(n10190),.clk(gclk));
	jand g09921(.dina(w_asqrt21_13[2]),.dinb(n10190),.dout(n10191),.clk(gclk));
	jand g09922(.dina(w_n10191_0[1]),.dinb(w_n9747_0[0]),.dout(n10192),.clk(gclk));
	jor g09923(.dina(n10192),.dinb(w_n9745_0[0]),.dout(n10193),.clk(gclk));
	jand g09924(.dina(w_n10191_0[0]),.dinb(w_n9748_0[0]),.dout(n10194),.clk(gclk));
	jnot g09925(.din(n10194),.dout(n10195),.clk(gclk));
	jand g09926(.dina(n10195),.dinb(n10193),.dout(n10196),.clk(gclk));
	jnot g09927(.din(w_n10196_0[2]),.dout(n10197),.clk(gclk));
	jand g09928(.dina(w_asqrt21_13[1]),.dinb(w_n9762_0[1]),.dout(n10198),.clk(gclk));
	jand g09929(.dina(w_n10198_0[1]),.dinb(w_n9749_1[0]),.dout(n10199),.clk(gclk));
	jor g09930(.dina(n10199),.dinb(w_n9797_0[0]),.dout(n10200),.clk(gclk));
	jor g09931(.dina(n10200),.dinb(w_n10197_0[1]),.dout(n10201),.clk(gclk));
	jor g09932(.dina(n10201),.dinb(w_n10189_0[2]),.dout(n10202),.clk(gclk));
	jand g09933(.dina(n10202),.dinb(w_n194_24[1]),.dout(n10203),.clk(gclk));
	jand g09934(.dina(w_n10197_0[0]),.dinb(w_n10189_0[1]),.dout(n10204),.clk(gclk));
	jor g09935(.dina(w_n10198_0[0]),.dinb(w_n9749_0[2]),.dout(n10205),.clk(gclk));
	jand g09936(.dina(w_n9762_0[0]),.dinb(w_n9749_0[1]),.dout(n10206),.clk(gclk));
	jor g09937(.dina(n10206),.dinb(w_n194_24[0]),.dout(n10207),.clk(gclk));
	jnot g09938(.din(n10207),.dout(n10208),.clk(gclk));
	jand g09939(.dina(n10208),.dinb(n10205),.dout(n10209),.clk(gclk));
	jor g09940(.dina(w_n10209_0[1]),.dinb(w_n10204_0[2]),.dout(n10212),.clk(gclk));
	jor g09941(.dina(n10212),.dinb(w_n10203_0[1]),.dout(asqrt_fa_21),.clk(gclk));
	jxor g09942(.dina(w_n9984_0[0]),.dinb(w_n2870_16[2]),.dout(n10214),.clk(gclk));
	jand g09943(.dina(n10214),.dinb(w_asqrt20_31),.dout(n10215),.clk(gclk));
	jxor g09944(.dina(n10215),.dinb(w_n9778_0[0]),.dout(n10216),.clk(gclk));
	jnot g09945(.din(n10216),.dout(n10217),.clk(gclk));
	jand g09946(.dina(w_asqrt20_30[2]),.dinb(w_a40_0[0]),.dout(n10218),.clk(gclk));
	jnot g09947(.din(w_a38_0[1]),.dout(n10219),.clk(gclk));
	jnot g09948(.din(w_a39_0[1]),.dout(n10220),.clk(gclk));
	jand g09949(.dina(w_n9780_1[0]),.dinb(w_n10220_0[1]),.dout(n10221),.clk(gclk));
	jand g09950(.dina(n10221),.dinb(w_n10219_1[1]),.dout(n10222),.clk(gclk));
	jor g09951(.dina(n10222),.dinb(n10218),.dout(n10223),.clk(gclk));
	jand g09952(.dina(w_n10223_0[2]),.dinb(w_asqrt21_13[0]),.dout(n10224),.clk(gclk));
	jand g09953(.dina(w_asqrt20_30[1]),.dinb(w_n9780_0[2]),.dout(n10225),.clk(gclk));
	jxor g09954(.dina(w_n10225_0[1]),.dinb(w_n9781_0[1]),.dout(n10226),.clk(gclk));
	jor g09955(.dina(w_n10223_0[1]),.dinb(w_asqrt21_12[2]),.dout(n10227),.clk(gclk));
	jand g09956(.dina(n10227),.dinb(w_n10226_0[1]),.dout(n10228),.clk(gclk));
	jor g09957(.dina(w_n10228_0[1]),.dinb(w_n10224_0[1]),.dout(n10229),.clk(gclk));
	jand g09958(.dina(n10229),.dinb(w_asqrt22_16[2]),.dout(n10230),.clk(gclk));
	jor g09959(.dina(w_n10224_0[0]),.dinb(w_asqrt22_16[1]),.dout(n10231),.clk(gclk));
	jor g09960(.dina(n10231),.dinb(w_n10228_0[0]),.dout(n10232),.clk(gclk));
	jand g09961(.dina(w_n10225_0[0]),.dinb(w_n9781_0[0]),.dout(n10233),.clk(gclk));
	jnot g09962(.din(w_n10203_0[0]),.dout(n10234),.clk(gclk));
	jnot g09963(.din(w_n10204_0[1]),.dout(n10235),.clk(gclk));
	jnot g09964(.din(w_n10209_0[0]),.dout(n10236),.clk(gclk));
	jand g09965(.dina(n10236),.dinb(w_asqrt21_12[1]),.dout(n10237),.clk(gclk));
	jand g09966(.dina(n10237),.dinb(n10235),.dout(n10238),.clk(gclk));
	jand g09967(.dina(n10238),.dinb(n10234),.dout(n10239),.clk(gclk));
	jor g09968(.dina(n10239),.dinb(n10233),.dout(n10240),.clk(gclk));
	jxor g09969(.dina(n10240),.dinb(w_n9318_0[1]),.dout(n10241),.clk(gclk));
	jand g09970(.dina(w_n10241_0[1]),.dinb(w_n10232_0[1]),.dout(n10242),.clk(gclk));
	jor g09971(.dina(n10242),.dinb(w_n10230_0[1]),.dout(n10243),.clk(gclk));
	jand g09972(.dina(w_n10243_0[2]),.dinb(w_asqrt23_12[2]),.dout(n10244),.clk(gclk));
	jor g09973(.dina(w_n10243_0[1]),.dinb(w_asqrt23_12[1]),.dout(n10245),.clk(gclk));
	jxor g09974(.dina(w_n9785_0[0]),.dinb(w_n9769_13[1]),.dout(n10246),.clk(gclk));
	jand g09975(.dina(n10246),.dinb(w_asqrt20_30[0]),.dout(n10247),.clk(gclk));
	jxor g09976(.dina(n10247),.dinb(w_n9788_0[0]),.dout(n10248),.clk(gclk));
	jnot g09977(.din(w_n10248_0[1]),.dout(n10249),.clk(gclk));
	jand g09978(.dina(n10249),.dinb(n10245),.dout(n10250),.clk(gclk));
	jor g09979(.dina(w_n10250_0[1]),.dinb(w_n10244_0[1]),.dout(n10251),.clk(gclk));
	jand g09980(.dina(n10251),.dinb(w_asqrt24_16[2]),.dout(n10252),.clk(gclk));
	jnot g09981(.din(w_n9794_0[0]),.dout(n10253),.clk(gclk));
	jand g09982(.dina(n10253),.dinb(w_n9792_0[0]),.dout(n10254),.clk(gclk));
	jand g09983(.dina(n10254),.dinb(w_asqrt20_29[2]),.dout(n10255),.clk(gclk));
	jxor g09984(.dina(n10255),.dinb(w_n9802_0[0]),.dout(n10256),.clk(gclk));
	jnot g09985(.din(n10256),.dout(n10257),.clk(gclk));
	jor g09986(.dina(w_n10244_0[0]),.dinb(w_asqrt24_16[1]),.dout(n10258),.clk(gclk));
	jor g09987(.dina(n10258),.dinb(w_n10250_0[0]),.dout(n10259),.clk(gclk));
	jand g09988(.dina(w_n10259_0[1]),.dinb(w_n10257_0[1]),.dout(n10260),.clk(gclk));
	jor g09989(.dina(w_n10260_0[1]),.dinb(w_n10252_0[1]),.dout(n10261),.clk(gclk));
	jand g09990(.dina(w_n10261_0[2]),.dinb(w_asqrt25_13[0]),.dout(n10262),.clk(gclk));
	jor g09991(.dina(w_n10261_0[1]),.dinb(w_asqrt25_12[2]),.dout(n10263),.clk(gclk));
	jnot g09992(.din(w_n9809_0[0]),.dout(n10264),.clk(gclk));
	jxor g09993(.dina(w_n9804_0[0]),.dinb(w_n8893_13[2]),.dout(n10265),.clk(gclk));
	jand g09994(.dina(n10265),.dinb(w_asqrt20_29[1]),.dout(n10266),.clk(gclk));
	jxor g09995(.dina(n10266),.dinb(n10264),.dout(n10267),.clk(gclk));
	jand g09996(.dina(w_n10267_0[1]),.dinb(n10263),.dout(n10268),.clk(gclk));
	jor g09997(.dina(w_n10268_0[1]),.dinb(w_n10262_0[1]),.dout(n10269),.clk(gclk));
	jand g09998(.dina(n10269),.dinb(w_asqrt26_16[2]),.dout(n10270),.clk(gclk));
	jor g09999(.dina(w_n10262_0[0]),.dinb(w_asqrt26_16[1]),.dout(n10271),.clk(gclk));
	jor g10000(.dina(n10271),.dinb(w_n10268_0[0]),.dout(n10272),.clk(gclk));
	jnot g10001(.din(w_n9816_0[0]),.dout(n10273),.clk(gclk));
	jnot g10002(.din(w_n9818_0[0]),.dout(n10274),.clk(gclk));
	jand g10003(.dina(w_asqrt20_29[0]),.dinb(w_n9812_0[0]),.dout(n10275),.clk(gclk));
	jand g10004(.dina(w_n10275_0[1]),.dinb(n10274),.dout(n10276),.clk(gclk));
	jor g10005(.dina(n10276),.dinb(n10273),.dout(n10277),.clk(gclk));
	jnot g10006(.din(w_n9819_0[0]),.dout(n10278),.clk(gclk));
	jand g10007(.dina(w_n10275_0[0]),.dinb(n10278),.dout(n10279),.clk(gclk));
	jnot g10008(.din(n10279),.dout(n10280),.clk(gclk));
	jand g10009(.dina(n10280),.dinb(n10277),.dout(n10281),.clk(gclk));
	jand g10010(.dina(w_n10281_0[1]),.dinb(w_n10272_0[1]),.dout(n10282),.clk(gclk));
	jor g10011(.dina(n10282),.dinb(w_n10270_0[1]),.dout(n10283),.clk(gclk));
	jand g10012(.dina(w_n10283_0[2]),.dinb(w_asqrt27_13[0]),.dout(n10284),.clk(gclk));
	jor g10013(.dina(w_n10283_0[1]),.dinb(w_asqrt27_12[2]),.dout(n10285),.clk(gclk));
	jxor g10014(.dina(w_n9820_0[0]),.dinb(w_n8053_13[2]),.dout(n10286),.clk(gclk));
	jand g10015(.dina(n10286),.dinb(w_asqrt20_28[2]),.dout(n10287),.clk(gclk));
	jxor g10016(.dina(n10287),.dinb(w_n9825_0[0]),.dout(n10288),.clk(gclk));
	jand g10017(.dina(w_n10288_0[1]),.dinb(n10285),.dout(n10289),.clk(gclk));
	jor g10018(.dina(w_n10289_0[1]),.dinb(w_n10284_0[1]),.dout(n10290),.clk(gclk));
	jand g10019(.dina(n10290),.dinb(w_asqrt28_16[2]),.dout(n10291),.clk(gclk));
	jnot g10020(.din(w_n9831_0[0]),.dout(n10292),.clk(gclk));
	jand g10021(.dina(n10292),.dinb(w_n9829_0[0]),.dout(n10293),.clk(gclk));
	jand g10022(.dina(n10293),.dinb(w_asqrt20_28[1]),.dout(n10294),.clk(gclk));
	jxor g10023(.dina(n10294),.dinb(w_n9840_0[0]),.dout(n10295),.clk(gclk));
	jnot g10024(.din(n10295),.dout(n10296),.clk(gclk));
	jor g10025(.dina(w_n10284_0[0]),.dinb(w_asqrt28_16[1]),.dout(n10297),.clk(gclk));
	jor g10026(.dina(n10297),.dinb(w_n10289_0[0]),.dout(n10298),.clk(gclk));
	jand g10027(.dina(w_n10298_0[1]),.dinb(w_n10296_0[1]),.dout(n10299),.clk(gclk));
	jor g10028(.dina(w_n10299_0[1]),.dinb(w_n10291_0[1]),.dout(n10300),.clk(gclk));
	jand g10029(.dina(w_n10300_0[2]),.dinb(w_asqrt29_13[1]),.dout(n10301),.clk(gclk));
	jor g10030(.dina(w_n10300_0[1]),.dinb(w_asqrt29_13[0]),.dout(n10302),.clk(gclk));
	jxor g10031(.dina(w_n9842_0[0]),.dinb(w_n7260_14[1]),.dout(n10303),.clk(gclk));
	jand g10032(.dina(n10303),.dinb(w_asqrt20_28[0]),.dout(n10304),.clk(gclk));
	jxor g10033(.dina(n10304),.dinb(w_n9848_0[0]),.dout(n10305),.clk(gclk));
	jand g10034(.dina(w_n10305_0[1]),.dinb(n10302),.dout(n10306),.clk(gclk));
	jor g10035(.dina(w_n10306_0[1]),.dinb(w_n10301_0[1]),.dout(n10307),.clk(gclk));
	jand g10036(.dina(n10307),.dinb(w_asqrt30_16[2]),.dout(n10308),.clk(gclk));
	jor g10037(.dina(w_n10301_0[0]),.dinb(w_asqrt30_16[1]),.dout(n10309),.clk(gclk));
	jor g10038(.dina(n10309),.dinb(w_n10306_0[0]),.dout(n10310),.clk(gclk));
	jnot g10039(.din(w_n9856_0[0]),.dout(n10311),.clk(gclk));
	jnot g10040(.din(w_n9858_0[0]),.dout(n10312),.clk(gclk));
	jand g10041(.dina(w_asqrt20_27[2]),.dinb(w_n9852_0[0]),.dout(n10313),.clk(gclk));
	jand g10042(.dina(w_n10313_0[1]),.dinb(n10312),.dout(n10314),.clk(gclk));
	jor g10043(.dina(n10314),.dinb(n10311),.dout(n10315),.clk(gclk));
	jnot g10044(.din(w_n9859_0[0]),.dout(n10316),.clk(gclk));
	jand g10045(.dina(w_n10313_0[0]),.dinb(n10316),.dout(n10317),.clk(gclk));
	jnot g10046(.din(n10317),.dout(n10318),.clk(gclk));
	jand g10047(.dina(n10318),.dinb(n10315),.dout(n10319),.clk(gclk));
	jand g10048(.dina(w_n10319_0[1]),.dinb(w_n10310_0[1]),.dout(n10320),.clk(gclk));
	jor g10049(.dina(n10320),.dinb(w_n10308_0[1]),.dout(n10321),.clk(gclk));
	jand g10050(.dina(w_n10321_0[1]),.dinb(w_asqrt31_13[1]),.dout(n10322),.clk(gclk));
	jxor g10051(.dina(w_n9860_0[0]),.dinb(w_n6500_14[1]),.dout(n10323),.clk(gclk));
	jand g10052(.dina(n10323),.dinb(w_asqrt20_27[1]),.dout(n10324),.clk(gclk));
	jxor g10053(.dina(n10324),.dinb(w_n9867_0[0]),.dout(n10325),.clk(gclk));
	jnot g10054(.din(n10325),.dout(n10326),.clk(gclk));
	jor g10055(.dina(w_n10321_0[0]),.dinb(w_asqrt31_13[0]),.dout(n10327),.clk(gclk));
	jand g10056(.dina(w_n10327_0[1]),.dinb(w_n10326_0[1]),.dout(n10328),.clk(gclk));
	jor g10057(.dina(w_n10328_0[2]),.dinb(w_n10322_0[2]),.dout(n10329),.clk(gclk));
	jand g10058(.dina(n10329),.dinb(w_asqrt32_16[2]),.dout(n10330),.clk(gclk));
	jnot g10059(.din(w_n9872_0[0]),.dout(n10331),.clk(gclk));
	jand g10060(.dina(n10331),.dinb(w_n9870_0[0]),.dout(n10332),.clk(gclk));
	jand g10061(.dina(n10332),.dinb(w_asqrt20_27[0]),.dout(n10333),.clk(gclk));
	jxor g10062(.dina(n10333),.dinb(w_n9880_0[0]),.dout(n10334),.clk(gclk));
	jnot g10063(.din(n10334),.dout(n10335),.clk(gclk));
	jor g10064(.dina(w_n10322_0[1]),.dinb(w_asqrt32_16[1]),.dout(n10336),.clk(gclk));
	jor g10065(.dina(n10336),.dinb(w_n10328_0[1]),.dout(n10337),.clk(gclk));
	jand g10066(.dina(w_n10337_0[1]),.dinb(w_n10335_0[1]),.dout(n10338),.clk(gclk));
	jor g10067(.dina(w_n10338_0[1]),.dinb(w_n10330_0[1]),.dout(n10339),.clk(gclk));
	jand g10068(.dina(w_n10339_0[2]),.dinb(w_asqrt33_13[2]),.dout(n10340),.clk(gclk));
	jor g10069(.dina(w_n10339_0[1]),.dinb(w_asqrt33_13[1]),.dout(n10341),.clk(gclk));
	jnot g10070(.din(w_n9886_0[0]),.dout(n10342),.clk(gclk));
	jnot g10071(.din(w_n9887_0[0]),.dout(n10343),.clk(gclk));
	jand g10072(.dina(w_asqrt20_26[2]),.dinb(w_n9883_0[0]),.dout(n10344),.clk(gclk));
	jand g10073(.dina(w_n10344_0[1]),.dinb(n10343),.dout(n10345),.clk(gclk));
	jor g10074(.dina(n10345),.dinb(n10342),.dout(n10346),.clk(gclk));
	jnot g10075(.din(w_n9888_0[0]),.dout(n10347),.clk(gclk));
	jand g10076(.dina(w_n10344_0[0]),.dinb(n10347),.dout(n10348),.clk(gclk));
	jnot g10077(.din(n10348),.dout(n10349),.clk(gclk));
	jand g10078(.dina(n10349),.dinb(n10346),.dout(n10350),.clk(gclk));
	jand g10079(.dina(w_n10350_0[1]),.dinb(n10341),.dout(n10351),.clk(gclk));
	jor g10080(.dina(w_n10351_0[1]),.dinb(w_n10340_0[1]),.dout(n10352),.clk(gclk));
	jand g10081(.dina(n10352),.dinb(w_asqrt34_16[2]),.dout(n10353),.clk(gclk));
	jor g10082(.dina(w_n10340_0[0]),.dinb(w_asqrt34_16[1]),.dout(n10354),.clk(gclk));
	jor g10083(.dina(n10354),.dinb(w_n10351_0[0]),.dout(n10355),.clk(gclk));
	jnot g10084(.din(w_n9894_0[0]),.dout(n10356),.clk(gclk));
	jnot g10085(.din(w_n9896_0[0]),.dout(n10357),.clk(gclk));
	jand g10086(.dina(w_asqrt20_26[1]),.dinb(w_n9890_0[0]),.dout(n10358),.clk(gclk));
	jand g10087(.dina(w_n10358_0[1]),.dinb(n10357),.dout(n10359),.clk(gclk));
	jor g10088(.dina(n10359),.dinb(n10356),.dout(n10360),.clk(gclk));
	jnot g10089(.din(w_n9897_0[0]),.dout(n10361),.clk(gclk));
	jand g10090(.dina(w_n10358_0[0]),.dinb(n10361),.dout(n10362),.clk(gclk));
	jnot g10091(.din(n10362),.dout(n10363),.clk(gclk));
	jand g10092(.dina(n10363),.dinb(n10360),.dout(n10364),.clk(gclk));
	jand g10093(.dina(w_n10364_0[1]),.dinb(w_n10355_0[1]),.dout(n10365),.clk(gclk));
	jor g10094(.dina(n10365),.dinb(w_n10353_0[1]),.dout(n10366),.clk(gclk));
	jand g10095(.dina(w_n10366_0[1]),.dinb(w_asqrt35_13[2]),.dout(n10367),.clk(gclk));
	jxor g10096(.dina(w_n9898_0[0]),.dinb(w_n5116_15[0]),.dout(n10368),.clk(gclk));
	jand g10097(.dina(n10368),.dinb(w_asqrt20_26[0]),.dout(n10369),.clk(gclk));
	jxor g10098(.dina(n10369),.dinb(w_n9908_0[0]),.dout(n10370),.clk(gclk));
	jnot g10099(.din(n10370),.dout(n10371),.clk(gclk));
	jor g10100(.dina(w_n10366_0[0]),.dinb(w_asqrt35_13[1]),.dout(n10372),.clk(gclk));
	jand g10101(.dina(w_n10372_0[1]),.dinb(w_n10371_0[1]),.dout(n10373),.clk(gclk));
	jor g10102(.dina(w_n10373_0[2]),.dinb(w_n10367_0[2]),.dout(n10374),.clk(gclk));
	jand g10103(.dina(n10374),.dinb(w_asqrt36_16[2]),.dout(n10375),.clk(gclk));
	jnot g10104(.din(w_n9913_0[0]),.dout(n10376),.clk(gclk));
	jand g10105(.dina(n10376),.dinb(w_n9911_0[0]),.dout(n10377),.clk(gclk));
	jand g10106(.dina(n10377),.dinb(w_asqrt20_25[2]),.dout(n10378),.clk(gclk));
	jxor g10107(.dina(n10378),.dinb(w_n9921_0[0]),.dout(n10379),.clk(gclk));
	jnot g10108(.din(n10379),.dout(n10380),.clk(gclk));
	jor g10109(.dina(w_n10367_0[1]),.dinb(w_asqrt36_16[1]),.dout(n10381),.clk(gclk));
	jor g10110(.dina(n10381),.dinb(w_n10373_0[1]),.dout(n10382),.clk(gclk));
	jand g10111(.dina(w_n10382_0[1]),.dinb(w_n10380_0[1]),.dout(n10383),.clk(gclk));
	jor g10112(.dina(w_n10383_0[1]),.dinb(w_n10375_0[1]),.dout(n10384),.clk(gclk));
	jand g10113(.dina(w_n10384_0[2]),.dinb(w_asqrt37_14[0]),.dout(n10385),.clk(gclk));
	jor g10114(.dina(w_n10384_0[1]),.dinb(w_asqrt37_13[2]),.dout(n10386),.clk(gclk));
	jnot g10115(.din(w_n9927_0[0]),.dout(n10387),.clk(gclk));
	jnot g10116(.din(w_n9928_0[0]),.dout(n10388),.clk(gclk));
	jand g10117(.dina(w_asqrt20_25[1]),.dinb(w_n9924_0[0]),.dout(n10389),.clk(gclk));
	jand g10118(.dina(w_n10389_0[1]),.dinb(n10388),.dout(n10390),.clk(gclk));
	jor g10119(.dina(n10390),.dinb(n10387),.dout(n10391),.clk(gclk));
	jnot g10120(.din(w_n9929_0[0]),.dout(n10392),.clk(gclk));
	jand g10121(.dina(w_n10389_0[0]),.dinb(n10392),.dout(n10393),.clk(gclk));
	jnot g10122(.din(n10393),.dout(n10394),.clk(gclk));
	jand g10123(.dina(n10394),.dinb(n10391),.dout(n10395),.clk(gclk));
	jand g10124(.dina(w_n10395_0[1]),.dinb(n10386),.dout(n10396),.clk(gclk));
	jor g10125(.dina(w_n10396_0[1]),.dinb(w_n10385_0[1]),.dout(n10397),.clk(gclk));
	jand g10126(.dina(n10397),.dinb(w_asqrt38_16[2]),.dout(n10398),.clk(gclk));
	jor g10127(.dina(w_n10385_0[0]),.dinb(w_asqrt38_16[1]),.dout(n10399),.clk(gclk));
	jor g10128(.dina(n10399),.dinb(w_n10396_0[0]),.dout(n10400),.clk(gclk));
	jnot g10129(.din(w_n9935_0[0]),.dout(n10401),.clk(gclk));
	jnot g10130(.din(w_n9937_0[0]),.dout(n10402),.clk(gclk));
	jand g10131(.dina(w_asqrt20_25[0]),.dinb(w_n9931_0[0]),.dout(n10403),.clk(gclk));
	jand g10132(.dina(w_n10403_0[1]),.dinb(n10402),.dout(n10404),.clk(gclk));
	jor g10133(.dina(n10404),.dinb(n10401),.dout(n10405),.clk(gclk));
	jnot g10134(.din(w_n9938_0[0]),.dout(n10406),.clk(gclk));
	jand g10135(.dina(w_n10403_0[0]),.dinb(n10406),.dout(n10407),.clk(gclk));
	jnot g10136(.din(n10407),.dout(n10408),.clk(gclk));
	jand g10137(.dina(n10408),.dinb(n10405),.dout(n10409),.clk(gclk));
	jand g10138(.dina(w_n10409_0[1]),.dinb(w_n10400_0[1]),.dout(n10410),.clk(gclk));
	jor g10139(.dina(n10410),.dinb(w_n10398_0[1]),.dout(n10411),.clk(gclk));
	jand g10140(.dina(w_n10411_0[1]),.dinb(w_asqrt39_14[0]),.dout(n10412),.clk(gclk));
	jxor g10141(.dina(w_n9939_0[0]),.dinb(w_n3907_16[0]),.dout(n10413),.clk(gclk));
	jand g10142(.dina(n10413),.dinb(w_asqrt20_24[2]),.dout(n10414),.clk(gclk));
	jxor g10143(.dina(n10414),.dinb(w_n9949_0[0]),.dout(n10415),.clk(gclk));
	jnot g10144(.din(n10415),.dout(n10416),.clk(gclk));
	jor g10145(.dina(w_n10411_0[0]),.dinb(w_asqrt39_13[2]),.dout(n10417),.clk(gclk));
	jand g10146(.dina(w_n10417_0[1]),.dinb(w_n10416_0[1]),.dout(n10418),.clk(gclk));
	jor g10147(.dina(w_n10418_0[2]),.dinb(w_n10412_0[2]),.dout(n10419),.clk(gclk));
	jand g10148(.dina(n10419),.dinb(w_asqrt40_16[2]),.dout(n10420),.clk(gclk));
	jnot g10149(.din(w_n9954_0[0]),.dout(n10421),.clk(gclk));
	jand g10150(.dina(n10421),.dinb(w_n9952_0[0]),.dout(n10422),.clk(gclk));
	jand g10151(.dina(n10422),.dinb(w_asqrt20_24[1]),.dout(n10423),.clk(gclk));
	jxor g10152(.dina(n10423),.dinb(w_n9962_0[0]),.dout(n10424),.clk(gclk));
	jnot g10153(.din(n10424),.dout(n10425),.clk(gclk));
	jor g10154(.dina(w_n10412_0[1]),.dinb(w_asqrt40_16[1]),.dout(n10426),.clk(gclk));
	jor g10155(.dina(n10426),.dinb(w_n10418_0[1]),.dout(n10427),.clk(gclk));
	jand g10156(.dina(w_n10427_0[1]),.dinb(w_n10425_0[1]),.dout(n10428),.clk(gclk));
	jor g10157(.dina(w_n10428_0[1]),.dinb(w_n10420_0[1]),.dout(n10429),.clk(gclk));
	jand g10158(.dina(w_n10429_0[2]),.dinb(w_asqrt41_14[1]),.dout(n10430),.clk(gclk));
	jor g10159(.dina(w_n10429_0[1]),.dinb(w_asqrt41_14[0]),.dout(n10431),.clk(gclk));
	jnot g10160(.din(w_n9968_0[0]),.dout(n10432),.clk(gclk));
	jnot g10161(.din(w_n9969_0[0]),.dout(n10433),.clk(gclk));
	jand g10162(.dina(w_asqrt20_24[0]),.dinb(w_n9965_0[0]),.dout(n10434),.clk(gclk));
	jand g10163(.dina(w_n10434_0[1]),.dinb(n10433),.dout(n10435),.clk(gclk));
	jor g10164(.dina(n10435),.dinb(n10432),.dout(n10436),.clk(gclk));
	jnot g10165(.din(w_n9970_0[0]),.dout(n10437),.clk(gclk));
	jand g10166(.dina(w_n10434_0[0]),.dinb(n10437),.dout(n10438),.clk(gclk));
	jnot g10167(.din(n10438),.dout(n10439),.clk(gclk));
	jand g10168(.dina(n10439),.dinb(n10436),.dout(n10440),.clk(gclk));
	jand g10169(.dina(w_n10440_0[1]),.dinb(n10431),.dout(n10441),.clk(gclk));
	jor g10170(.dina(w_n10441_0[1]),.dinb(w_n10430_0[1]),.dout(n10442),.clk(gclk));
	jand g10171(.dina(n10442),.dinb(w_asqrt42_16[2]),.dout(n10443),.clk(gclk));
	jnot g10172(.din(w_n9974_0[0]),.dout(n10444),.clk(gclk));
	jand g10173(.dina(n10444),.dinb(w_n9972_0[0]),.dout(n10445),.clk(gclk));
	jand g10174(.dina(n10445),.dinb(w_asqrt20_23[2]),.dout(n10446),.clk(gclk));
	jxor g10175(.dina(n10446),.dinb(w_n9982_0[0]),.dout(n10447),.clk(gclk));
	jnot g10176(.din(n10447),.dout(n10448),.clk(gclk));
	jor g10177(.dina(w_n10430_0[0]),.dinb(w_asqrt42_16[1]),.dout(n10449),.clk(gclk));
	jor g10178(.dina(n10449),.dinb(w_n10441_0[0]),.dout(n10450),.clk(gclk));
	jand g10179(.dina(w_n10450_0[1]),.dinb(w_n10448_0[1]),.dout(n10451),.clk(gclk));
	jor g10180(.dina(w_n10451_0[1]),.dinb(w_n10443_0[1]),.dout(n10452),.clk(gclk));
	jand g10181(.dina(w_n10452_0[2]),.dinb(w_asqrt43_14[1]),.dout(n10453),.clk(gclk));
	jor g10182(.dina(w_n10452_0[1]),.dinb(w_asqrt43_14[0]),.dout(n10454),.clk(gclk));
	jand g10183(.dina(n10454),.dinb(w_n10217_0[1]),.dout(n10455),.clk(gclk));
	jor g10184(.dina(w_n10455_0[1]),.dinb(w_n10453_0[1]),.dout(n10456),.clk(gclk));
	jand g10185(.dina(n10456),.dinb(w_asqrt44_16[2]),.dout(n10457),.clk(gclk));
	jor g10186(.dina(w_n10453_0[0]),.dinb(w_asqrt44_16[1]),.dout(n10458),.clk(gclk));
	jor g10187(.dina(n10458),.dinb(w_n10455_0[0]),.dout(n10459),.clk(gclk));
	jnot g10188(.din(w_n9993_0[0]),.dout(n10460),.clk(gclk));
	jnot g10189(.din(w_n9995_0[0]),.dout(n10461),.clk(gclk));
	jand g10190(.dina(w_asqrt20_23[1]),.dinb(w_n9989_0[0]),.dout(n10462),.clk(gclk));
	jand g10191(.dina(w_n10462_0[1]),.dinb(n10461),.dout(n10463),.clk(gclk));
	jor g10192(.dina(n10463),.dinb(n10460),.dout(n10464),.clk(gclk));
	jnot g10193(.din(w_n9996_0[0]),.dout(n10465),.clk(gclk));
	jand g10194(.dina(w_n10462_0[0]),.dinb(n10465),.dout(n10466),.clk(gclk));
	jnot g10195(.din(n10466),.dout(n10467),.clk(gclk));
	jand g10196(.dina(n10467),.dinb(n10464),.dout(n10468),.clk(gclk));
	jand g10197(.dina(w_n10468_0[1]),.dinb(w_n10459_0[1]),.dout(n10469),.clk(gclk));
	jor g10198(.dina(n10469),.dinb(w_n10457_0[1]),.dout(n10470),.clk(gclk));
	jand g10199(.dina(w_n10470_0[2]),.dinb(w_asqrt45_14[2]),.dout(n10471),.clk(gclk));
	jor g10200(.dina(w_n10470_0[1]),.dinb(w_asqrt45_14[1]),.dout(n10472),.clk(gclk));
	jnot g10201(.din(w_n10001_0[0]),.dout(n10473),.clk(gclk));
	jnot g10202(.din(w_n10002_0[0]),.dout(n10474),.clk(gclk));
	jand g10203(.dina(w_asqrt20_23[0]),.dinb(w_n9998_0[0]),.dout(n10475),.clk(gclk));
	jand g10204(.dina(w_n10475_0[1]),.dinb(n10474),.dout(n10476),.clk(gclk));
	jor g10205(.dina(n10476),.dinb(n10473),.dout(n10477),.clk(gclk));
	jnot g10206(.din(w_n10003_0[0]),.dout(n10478),.clk(gclk));
	jand g10207(.dina(w_n10475_0[0]),.dinb(n10478),.dout(n10479),.clk(gclk));
	jnot g10208(.din(n10479),.dout(n10480),.clk(gclk));
	jand g10209(.dina(n10480),.dinb(n10477),.dout(n10481),.clk(gclk));
	jand g10210(.dina(w_n10481_0[1]),.dinb(n10472),.dout(n10482),.clk(gclk));
	jor g10211(.dina(w_n10482_0[1]),.dinb(w_n10471_0[1]),.dout(n10483),.clk(gclk));
	jand g10212(.dina(n10483),.dinb(w_asqrt46_16[2]),.dout(n10484),.clk(gclk));
	jor g10213(.dina(w_n10471_0[0]),.dinb(w_asqrt46_16[1]),.dout(n10485),.clk(gclk));
	jor g10214(.dina(n10485),.dinb(w_n10482_0[0]),.dout(n10486),.clk(gclk));
	jnot g10215(.din(w_n10009_0[0]),.dout(n10487),.clk(gclk));
	jnot g10216(.din(w_n10011_0[0]),.dout(n10488),.clk(gclk));
	jand g10217(.dina(w_asqrt20_22[2]),.dinb(w_n10005_0[0]),.dout(n10489),.clk(gclk));
	jand g10218(.dina(w_n10489_0[1]),.dinb(n10488),.dout(n10490),.clk(gclk));
	jor g10219(.dina(n10490),.dinb(n10487),.dout(n10491),.clk(gclk));
	jnot g10220(.din(w_n10012_0[0]),.dout(n10492),.clk(gclk));
	jand g10221(.dina(w_n10489_0[0]),.dinb(n10492),.dout(n10493),.clk(gclk));
	jnot g10222(.din(n10493),.dout(n10494),.clk(gclk));
	jand g10223(.dina(n10494),.dinb(n10491),.dout(n10495),.clk(gclk));
	jand g10224(.dina(w_n10495_0[1]),.dinb(w_n10486_0[1]),.dout(n10496),.clk(gclk));
	jor g10225(.dina(n10496),.dinb(w_n10484_0[1]),.dout(n10497),.clk(gclk));
	jand g10226(.dina(w_n10497_0[1]),.dinb(w_asqrt47_14[2]),.dout(n10498),.clk(gclk));
	jxor g10227(.dina(w_n10013_0[0]),.dinb(w_n2005_17[2]),.dout(n10499),.clk(gclk));
	jand g10228(.dina(n10499),.dinb(w_asqrt20_22[1]),.dout(n10500),.clk(gclk));
	jxor g10229(.dina(n10500),.dinb(w_n10023_0[0]),.dout(n10501),.clk(gclk));
	jnot g10230(.din(n10501),.dout(n10502),.clk(gclk));
	jor g10231(.dina(w_n10497_0[0]),.dinb(w_asqrt47_14[1]),.dout(n10503),.clk(gclk));
	jand g10232(.dina(w_n10503_0[1]),.dinb(w_n10502_0[1]),.dout(n10504),.clk(gclk));
	jor g10233(.dina(w_n10504_0[2]),.dinb(w_n10498_0[2]),.dout(n10505),.clk(gclk));
	jand g10234(.dina(n10505),.dinb(w_asqrt48_16[2]),.dout(n10506),.clk(gclk));
	jnot g10235(.din(w_n10028_0[0]),.dout(n10507),.clk(gclk));
	jand g10236(.dina(n10507),.dinb(w_n10026_0[0]),.dout(n10508),.clk(gclk));
	jand g10237(.dina(n10508),.dinb(w_asqrt20_22[0]),.dout(n10509),.clk(gclk));
	jxor g10238(.dina(n10509),.dinb(w_n10036_0[0]),.dout(n10510),.clk(gclk));
	jnot g10239(.din(n10510),.dout(n10511),.clk(gclk));
	jor g10240(.dina(w_n10498_0[1]),.dinb(w_asqrt48_16[1]),.dout(n10512),.clk(gclk));
	jor g10241(.dina(n10512),.dinb(w_n10504_0[1]),.dout(n10513),.clk(gclk));
	jand g10242(.dina(w_n10513_0[1]),.dinb(w_n10511_0[1]),.dout(n10514),.clk(gclk));
	jor g10243(.dina(w_n10514_0[1]),.dinb(w_n10506_0[1]),.dout(n10515),.clk(gclk));
	jand g10244(.dina(w_n10515_0[2]),.dinb(w_asqrt49_15[0]),.dout(n10516),.clk(gclk));
	jor g10245(.dina(w_n10515_0[1]),.dinb(w_asqrt49_14[2]),.dout(n10517),.clk(gclk));
	jnot g10246(.din(w_n10042_0[0]),.dout(n10518),.clk(gclk));
	jnot g10247(.din(w_n10043_0[0]),.dout(n10519),.clk(gclk));
	jand g10248(.dina(w_asqrt20_21[2]),.dinb(w_n10039_0[0]),.dout(n10520),.clk(gclk));
	jand g10249(.dina(w_n10520_0[1]),.dinb(n10519),.dout(n10521),.clk(gclk));
	jor g10250(.dina(n10521),.dinb(n10518),.dout(n10522),.clk(gclk));
	jnot g10251(.din(w_n10044_0[0]),.dout(n10523),.clk(gclk));
	jand g10252(.dina(w_n10520_0[0]),.dinb(n10523),.dout(n10524),.clk(gclk));
	jnot g10253(.din(n10524),.dout(n10525),.clk(gclk));
	jand g10254(.dina(n10525),.dinb(n10522),.dout(n10526),.clk(gclk));
	jand g10255(.dina(w_n10526_0[1]),.dinb(n10517),.dout(n10527),.clk(gclk));
	jor g10256(.dina(w_n10527_0[1]),.dinb(w_n10516_0[1]),.dout(n10528),.clk(gclk));
	jand g10257(.dina(n10528),.dinb(w_asqrt50_16[2]),.dout(n10529),.clk(gclk));
	jor g10258(.dina(w_n10516_0[0]),.dinb(w_asqrt50_16[1]),.dout(n10530),.clk(gclk));
	jor g10259(.dina(n10530),.dinb(w_n10527_0[0]),.dout(n10531),.clk(gclk));
	jnot g10260(.din(w_n10050_0[0]),.dout(n10532),.clk(gclk));
	jnot g10261(.din(w_n10052_0[0]),.dout(n10533),.clk(gclk));
	jand g10262(.dina(w_asqrt20_21[1]),.dinb(w_n10046_0[0]),.dout(n10534),.clk(gclk));
	jand g10263(.dina(w_n10534_0[1]),.dinb(n10533),.dout(n10535),.clk(gclk));
	jor g10264(.dina(n10535),.dinb(n10532),.dout(n10536),.clk(gclk));
	jnot g10265(.din(w_n10053_0[0]),.dout(n10537),.clk(gclk));
	jand g10266(.dina(w_n10534_0[0]),.dinb(n10537),.dout(n10538),.clk(gclk));
	jnot g10267(.din(n10538),.dout(n10539),.clk(gclk));
	jand g10268(.dina(n10539),.dinb(n10536),.dout(n10540),.clk(gclk));
	jand g10269(.dina(w_n10540_0[1]),.dinb(w_n10531_0[1]),.dout(n10541),.clk(gclk));
	jor g10270(.dina(n10541),.dinb(w_n10529_0[1]),.dout(n10542),.clk(gclk));
	jand g10271(.dina(w_n10542_0[1]),.dinb(w_asqrt51_15[0]),.dout(n10543),.clk(gclk));
	jxor g10272(.dina(w_n10054_0[0]),.dinb(w_n1312_18[1]),.dout(n10544),.clk(gclk));
	jand g10273(.dina(n10544),.dinb(w_asqrt20_21[0]),.dout(n10545),.clk(gclk));
	jxor g10274(.dina(n10545),.dinb(w_n10064_0[0]),.dout(n10546),.clk(gclk));
	jnot g10275(.din(n10546),.dout(n10547),.clk(gclk));
	jor g10276(.dina(w_n10542_0[0]),.dinb(w_asqrt51_14[2]),.dout(n10548),.clk(gclk));
	jand g10277(.dina(w_n10548_0[1]),.dinb(w_n10547_0[1]),.dout(n10549),.clk(gclk));
	jor g10278(.dina(w_n10549_0[2]),.dinb(w_n10543_0[2]),.dout(n10550),.clk(gclk));
	jand g10279(.dina(n10550),.dinb(w_asqrt52_16[2]),.dout(n10551),.clk(gclk));
	jnot g10280(.din(w_n10069_0[0]),.dout(n10552),.clk(gclk));
	jand g10281(.dina(n10552),.dinb(w_n10067_0[0]),.dout(n10553),.clk(gclk));
	jand g10282(.dina(n10553),.dinb(w_asqrt20_20[2]),.dout(n10554),.clk(gclk));
	jxor g10283(.dina(n10554),.dinb(w_n10077_0[0]),.dout(n10555),.clk(gclk));
	jnot g10284(.din(n10555),.dout(n10556),.clk(gclk));
	jor g10285(.dina(w_n10543_0[1]),.dinb(w_asqrt52_16[1]),.dout(n10557),.clk(gclk));
	jor g10286(.dina(n10557),.dinb(w_n10549_0[1]),.dout(n10558),.clk(gclk));
	jand g10287(.dina(w_n10558_0[1]),.dinb(w_n10556_0[1]),.dout(n10559),.clk(gclk));
	jor g10288(.dina(w_n10559_0[1]),.dinb(w_n10551_0[1]),.dout(n10560),.clk(gclk));
	jand g10289(.dina(w_n10560_0[2]),.dinb(w_asqrt53_15[1]),.dout(n10561),.clk(gclk));
	jor g10290(.dina(w_n10560_0[1]),.dinb(w_asqrt53_15[0]),.dout(n10562),.clk(gclk));
	jnot g10291(.din(w_n10083_0[0]),.dout(n10563),.clk(gclk));
	jnot g10292(.din(w_n10084_0[0]),.dout(n10564),.clk(gclk));
	jand g10293(.dina(w_asqrt20_20[1]),.dinb(w_n10080_0[0]),.dout(n10565),.clk(gclk));
	jand g10294(.dina(w_n10565_0[1]),.dinb(n10564),.dout(n10566),.clk(gclk));
	jor g10295(.dina(n10566),.dinb(n10563),.dout(n10567),.clk(gclk));
	jnot g10296(.din(w_n10085_0[0]),.dout(n10568),.clk(gclk));
	jand g10297(.dina(w_n10565_0[0]),.dinb(n10568),.dout(n10569),.clk(gclk));
	jnot g10298(.din(n10569),.dout(n10570),.clk(gclk));
	jand g10299(.dina(n10570),.dinb(n10567),.dout(n10571),.clk(gclk));
	jand g10300(.dina(w_n10571_0[1]),.dinb(n10562),.dout(n10572),.clk(gclk));
	jor g10301(.dina(w_n10572_0[1]),.dinb(w_n10561_0[1]),.dout(n10573),.clk(gclk));
	jand g10302(.dina(n10573),.dinb(w_asqrt54_16[2]),.dout(n10574),.clk(gclk));
	jor g10303(.dina(w_n10561_0[0]),.dinb(w_asqrt54_16[1]),.dout(n10575),.clk(gclk));
	jor g10304(.dina(n10575),.dinb(w_n10572_0[0]),.dout(n10576),.clk(gclk));
	jnot g10305(.din(w_n10091_0[0]),.dout(n10577),.clk(gclk));
	jnot g10306(.din(w_n10093_0[0]),.dout(n10578),.clk(gclk));
	jand g10307(.dina(w_asqrt20_20[0]),.dinb(w_n10087_0[0]),.dout(n10579),.clk(gclk));
	jand g10308(.dina(w_n10579_0[1]),.dinb(n10578),.dout(n10580),.clk(gclk));
	jor g10309(.dina(n10580),.dinb(n10577),.dout(n10581),.clk(gclk));
	jnot g10310(.din(w_n10094_0[0]),.dout(n10582),.clk(gclk));
	jand g10311(.dina(w_n10579_0[0]),.dinb(n10582),.dout(n10583),.clk(gclk));
	jnot g10312(.din(n10583),.dout(n10584),.clk(gclk));
	jand g10313(.dina(n10584),.dinb(n10581),.dout(n10585),.clk(gclk));
	jand g10314(.dina(w_n10585_0[1]),.dinb(w_n10576_0[1]),.dout(n10586),.clk(gclk));
	jor g10315(.dina(n10586),.dinb(w_n10574_0[1]),.dout(n10587),.clk(gclk));
	jand g10316(.dina(w_n10587_0[1]),.dinb(w_asqrt55_15[2]),.dout(n10588),.clk(gclk));
	jxor g10317(.dina(w_n10095_0[0]),.dinb(w_n791_19[1]),.dout(n10589),.clk(gclk));
	jand g10318(.dina(n10589),.dinb(w_asqrt20_19[2]),.dout(n10590),.clk(gclk));
	jxor g10319(.dina(n10590),.dinb(w_n10105_0[0]),.dout(n10591),.clk(gclk));
	jnot g10320(.din(n10591),.dout(n10592),.clk(gclk));
	jor g10321(.dina(w_n10587_0[0]),.dinb(w_asqrt55_15[1]),.dout(n10593),.clk(gclk));
	jand g10322(.dina(w_n10593_0[1]),.dinb(w_n10592_0[1]),.dout(n10594),.clk(gclk));
	jor g10323(.dina(w_n10594_0[2]),.dinb(w_n10588_0[2]),.dout(n10595),.clk(gclk));
	jand g10324(.dina(n10595),.dinb(w_asqrt56_16[2]),.dout(n10596),.clk(gclk));
	jnot g10325(.din(w_n10110_0[0]),.dout(n10597),.clk(gclk));
	jand g10326(.dina(n10597),.dinb(w_n10108_0[0]),.dout(n10598),.clk(gclk));
	jand g10327(.dina(n10598),.dinb(w_asqrt20_19[1]),.dout(n10599),.clk(gclk));
	jxor g10328(.dina(n10599),.dinb(w_n10118_0[0]),.dout(n10600),.clk(gclk));
	jnot g10329(.din(n10600),.dout(n10601),.clk(gclk));
	jor g10330(.dina(w_n10588_0[1]),.dinb(w_asqrt56_16[1]),.dout(n10602),.clk(gclk));
	jor g10331(.dina(n10602),.dinb(w_n10594_0[1]),.dout(n10603),.clk(gclk));
	jand g10332(.dina(w_n10603_0[1]),.dinb(w_n10601_0[1]),.dout(n10604),.clk(gclk));
	jor g10333(.dina(w_n10604_0[1]),.dinb(w_n10596_0[1]),.dout(n10605),.clk(gclk));
	jand g10334(.dina(w_n10605_0[2]),.dinb(w_asqrt57_16[0]),.dout(n10606),.clk(gclk));
	jor g10335(.dina(w_n10605_0[1]),.dinb(w_asqrt57_15[2]),.dout(n10607),.clk(gclk));
	jnot g10336(.din(w_n10124_0[0]),.dout(n10608),.clk(gclk));
	jnot g10337(.din(w_n10125_0[0]),.dout(n10609),.clk(gclk));
	jand g10338(.dina(w_asqrt20_19[0]),.dinb(w_n10121_0[0]),.dout(n10610),.clk(gclk));
	jand g10339(.dina(w_n10610_0[1]),.dinb(n10609),.dout(n10611),.clk(gclk));
	jor g10340(.dina(n10611),.dinb(n10608),.dout(n10612),.clk(gclk));
	jnot g10341(.din(w_n10126_0[0]),.dout(n10613),.clk(gclk));
	jand g10342(.dina(w_n10610_0[0]),.dinb(n10613),.dout(n10614),.clk(gclk));
	jnot g10343(.din(n10614),.dout(n10615),.clk(gclk));
	jand g10344(.dina(n10615),.dinb(n10612),.dout(n10616),.clk(gclk));
	jand g10345(.dina(w_n10616_0[1]),.dinb(n10607),.dout(n10617),.clk(gclk));
	jor g10346(.dina(w_n10617_0[1]),.dinb(w_n10606_0[1]),.dout(n10618),.clk(gclk));
	jand g10347(.dina(n10618),.dinb(w_asqrt58_16[2]),.dout(n10619),.clk(gclk));
	jor g10348(.dina(w_n10606_0[0]),.dinb(w_asqrt58_16[1]),.dout(n10620),.clk(gclk));
	jor g10349(.dina(n10620),.dinb(w_n10617_0[0]),.dout(n10621),.clk(gclk));
	jnot g10350(.din(w_n10132_0[0]),.dout(n10622),.clk(gclk));
	jnot g10351(.din(w_n10134_0[0]),.dout(n10623),.clk(gclk));
	jand g10352(.dina(w_asqrt20_18[2]),.dinb(w_n10128_0[0]),.dout(n10624),.clk(gclk));
	jand g10353(.dina(w_n10624_0[1]),.dinb(n10623),.dout(n10625),.clk(gclk));
	jor g10354(.dina(n10625),.dinb(n10622),.dout(n10626),.clk(gclk));
	jnot g10355(.din(w_n10135_0[0]),.dout(n10627),.clk(gclk));
	jand g10356(.dina(w_n10624_0[0]),.dinb(n10627),.dout(n10628),.clk(gclk));
	jnot g10357(.din(n10628),.dout(n10629),.clk(gclk));
	jand g10358(.dina(n10629),.dinb(n10626),.dout(n10630),.clk(gclk));
	jand g10359(.dina(w_n10630_0[1]),.dinb(w_n10621_0[1]),.dout(n10631),.clk(gclk));
	jor g10360(.dina(n10631),.dinb(w_n10619_0[1]),.dout(n10632),.clk(gclk));
	jand g10361(.dina(w_n10632_0[1]),.dinb(w_asqrt59_16[1]),.dout(n10633),.clk(gclk));
	jxor g10362(.dina(w_n10136_0[0]),.dinb(w_n425_20[0]),.dout(n10634),.clk(gclk));
	jand g10363(.dina(n10634),.dinb(w_asqrt20_18[1]),.dout(n10635),.clk(gclk));
	jxor g10364(.dina(n10635),.dinb(w_n10146_0[0]),.dout(n10636),.clk(gclk));
	jnot g10365(.din(n10636),.dout(n10637),.clk(gclk));
	jor g10366(.dina(w_n10632_0[0]),.dinb(w_asqrt59_16[0]),.dout(n10638),.clk(gclk));
	jand g10367(.dina(w_n10638_0[1]),.dinb(w_n10637_0[1]),.dout(n10639),.clk(gclk));
	jor g10368(.dina(w_n10639_0[2]),.dinb(w_n10633_0[2]),.dout(n10640),.clk(gclk));
	jand g10369(.dina(n10640),.dinb(w_asqrt60_16[1]),.dout(n10641),.clk(gclk));
	jnot g10370(.din(w_n10151_0[0]),.dout(n10642),.clk(gclk));
	jand g10371(.dina(n10642),.dinb(w_n10149_0[0]),.dout(n10643),.clk(gclk));
	jand g10372(.dina(n10643),.dinb(w_asqrt20_18[0]),.dout(n10644),.clk(gclk));
	jxor g10373(.dina(n10644),.dinb(w_n10159_0[0]),.dout(n10645),.clk(gclk));
	jnot g10374(.din(n10645),.dout(n10646),.clk(gclk));
	jor g10375(.dina(w_n10633_0[1]),.dinb(w_asqrt60_16[0]),.dout(n10647),.clk(gclk));
	jor g10376(.dina(n10647),.dinb(w_n10639_0[1]),.dout(n10648),.clk(gclk));
	jand g10377(.dina(w_n10648_0[1]),.dinb(w_n10646_0[1]),.dout(n10649),.clk(gclk));
	jor g10378(.dina(w_n10649_0[1]),.dinb(w_n10641_0[1]),.dout(n10650),.clk(gclk));
	jand g10379(.dina(w_n10650_0[2]),.dinb(w_asqrt61_16[2]),.dout(n10651),.clk(gclk));
	jor g10380(.dina(w_n10650_0[1]),.dinb(w_asqrt61_16[1]),.dout(n10652),.clk(gclk));
	jnot g10381(.din(w_n10165_0[0]),.dout(n10653),.clk(gclk));
	jnot g10382(.din(w_n10166_0[0]),.dout(n10654),.clk(gclk));
	jand g10383(.dina(w_asqrt20_17[2]),.dinb(w_n10162_0[0]),.dout(n10655),.clk(gclk));
	jand g10384(.dina(w_n10655_0[1]),.dinb(n10654),.dout(n10656),.clk(gclk));
	jor g10385(.dina(n10656),.dinb(n10653),.dout(n10657),.clk(gclk));
	jnot g10386(.din(w_n10167_0[0]),.dout(n10658),.clk(gclk));
	jand g10387(.dina(w_n10655_0[0]),.dinb(n10658),.dout(n10659),.clk(gclk));
	jnot g10388(.din(n10659),.dout(n10660),.clk(gclk));
	jand g10389(.dina(n10660),.dinb(n10657),.dout(n10661),.clk(gclk));
	jand g10390(.dina(w_n10661_0[1]),.dinb(n10652),.dout(n10662),.clk(gclk));
	jor g10391(.dina(w_n10662_0[1]),.dinb(w_n10651_0[1]),.dout(n10663),.clk(gclk));
	jand g10392(.dina(n10663),.dinb(w_asqrt62_16[2]),.dout(n10664),.clk(gclk));
	jor g10393(.dina(w_n10651_0[0]),.dinb(w_asqrt62_16[1]),.dout(n10665),.clk(gclk));
	jor g10394(.dina(n10665),.dinb(w_n10662_0[0]),.dout(n10666),.clk(gclk));
	jnot g10395(.din(w_n10173_0[0]),.dout(n10667),.clk(gclk));
	jnot g10396(.din(w_n10175_0[0]),.dout(n10668),.clk(gclk));
	jand g10397(.dina(w_asqrt20_17[1]),.dinb(w_n10169_0[0]),.dout(n10669),.clk(gclk));
	jand g10398(.dina(w_n10669_0[1]),.dinb(n10668),.dout(n10670),.clk(gclk));
	jor g10399(.dina(n10670),.dinb(n10667),.dout(n10671),.clk(gclk));
	jnot g10400(.din(w_n10176_0[0]),.dout(n10672),.clk(gclk));
	jand g10401(.dina(w_n10669_0[0]),.dinb(n10672),.dout(n10673),.clk(gclk));
	jnot g10402(.din(n10673),.dout(n10674),.clk(gclk));
	jand g10403(.dina(n10674),.dinb(n10671),.dout(n10675),.clk(gclk));
	jand g10404(.dina(w_n10675_0[1]),.dinb(w_n10666_0[1]),.dout(n10676),.clk(gclk));
	jor g10405(.dina(n10676),.dinb(w_n10664_0[1]),.dout(n10677),.clk(gclk));
	jxor g10406(.dina(w_n10177_0[0]),.dinb(w_n199_24[2]),.dout(n10678),.clk(gclk));
	jand g10407(.dina(n10678),.dinb(w_asqrt20_17[0]),.dout(n10679),.clk(gclk));
	jxor g10408(.dina(n10679),.dinb(w_n10187_0[0]),.dout(n10680),.clk(gclk));
	jnot g10409(.din(w_n10189_0[0]),.dout(n10681),.clk(gclk));
	jand g10410(.dina(w_asqrt20_16[2]),.dinb(w_n10196_0[1]),.dout(n10682),.clk(gclk));
	jand g10411(.dina(w_n10682_0[1]),.dinb(w_n10681_0[2]),.dout(n10683),.clk(gclk));
	jor g10412(.dina(n10683),.dinb(w_n10204_0[0]),.dout(n10684),.clk(gclk));
	jor g10413(.dina(n10684),.dinb(w_n10680_0[1]),.dout(n10685),.clk(gclk));
	jnot g10414(.din(n10685),.dout(n10686),.clk(gclk));
	jand g10415(.dina(n10686),.dinb(w_n10677_1[2]),.dout(n10687),.clk(gclk));
	jor g10416(.dina(n10687),.dinb(w_asqrt63_9[0]),.dout(n10688),.clk(gclk));
	jnot g10417(.din(w_n10680_0[0]),.dout(n10689),.clk(gclk));
	jor g10418(.dina(w_n10689_0[2]),.dinb(w_n10677_1[1]),.dout(n10690),.clk(gclk));
	jor g10419(.dina(w_n10682_0[0]),.dinb(w_n10681_0[1]),.dout(n10691),.clk(gclk));
	jand g10420(.dina(w_n10196_0[0]),.dinb(w_n10681_0[0]),.dout(n10692),.clk(gclk));
	jor g10421(.dina(n10692),.dinb(w_n194_23[2]),.dout(n10693),.clk(gclk));
	jnot g10422(.din(n10693),.dout(n10694),.clk(gclk));
	jand g10423(.dina(n10694),.dinb(n10691),.dout(n10695),.clk(gclk));
	jnot g10424(.din(w_asqrt20_16[1]),.dout(n10696),.clk(gclk));
	jnot g10425(.din(w_n10695_0[1]),.dout(n10699),.clk(gclk));
	jand g10426(.dina(n10699),.dinb(w_n10690_0[1]),.dout(n10700),.clk(gclk));
	jand g10427(.dina(n10700),.dinb(w_n10688_0[1]),.dout(n10701),.clk(gclk));
	jxor g10428(.dina(w_n10452_0[0]),.dinb(w_n2425_19[2]),.dout(n10702),.clk(gclk));
	jor g10429(.dina(n10702),.dinb(w_n10701_25[2]),.dout(n10703),.clk(gclk));
	jxor g10430(.dina(n10703),.dinb(w_n10217_0[0]),.dout(n10704),.clk(gclk));
	jor g10431(.dina(w_n10701_25[1]),.dinb(w_n10219_1[0]),.dout(n10705),.clk(gclk));
	jnot g10432(.din(w_a36_0[1]),.dout(n10706),.clk(gclk));
	jnot g10433(.din(a[37]),.dout(n10707),.clk(gclk));
	jand g10434(.dina(w_n10219_0[2]),.dinb(w_n10707_0[2]),.dout(n10708),.clk(gclk));
	jand g10435(.dina(n10708),.dinb(w_n10706_1[1]),.dout(n10709),.clk(gclk));
	jnot g10436(.din(n10709),.dout(n10710),.clk(gclk));
	jand g10437(.dina(n10710),.dinb(n10705),.dout(n10711),.clk(gclk));
	jor g10438(.dina(w_n10711_0[2]),.dinb(w_n10696_13[1]),.dout(n10712),.clk(gclk));
	jor g10439(.dina(w_n10701_25[0]),.dinb(w_a38_0[0]),.dout(n10713),.clk(gclk));
	jxor g10440(.dina(w_n10713_0[1]),.dinb(w_n10220_0[0]),.dout(n10714),.clk(gclk));
	jand g10441(.dina(w_n10711_0[1]),.dinb(w_n10696_13[0]),.dout(n10715),.clk(gclk));
	jor g10442(.dina(n10715),.dinb(w_n10714_0[1]),.dout(n10716),.clk(gclk));
	jand g10443(.dina(w_n10716_0[1]),.dinb(w_n10712_0[1]),.dout(n10717),.clk(gclk));
	jor g10444(.dina(n10717),.dinb(w_n9774_17[0]),.dout(n10718),.clk(gclk));
	jand g10445(.dina(w_n10712_0[0]),.dinb(w_n9774_16[2]),.dout(n10719),.clk(gclk));
	jand g10446(.dina(n10719),.dinb(w_n10716_0[0]),.dout(n10720),.clk(gclk));
	jor g10447(.dina(w_n10713_0[0]),.dinb(w_a39_0[0]),.dout(n10721),.clk(gclk));
	jnot g10448(.din(w_n10688_0[0]),.dout(n10722),.clk(gclk));
	jnot g10449(.din(w_n10690_0[0]),.dout(n10723),.clk(gclk));
	jor g10450(.dina(w_n10695_0[0]),.dinb(w_n10696_12[2]),.dout(n10724),.clk(gclk));
	jor g10451(.dina(n10724),.dinb(w_n10723_0[1]),.dout(n10725),.clk(gclk));
	jor g10452(.dina(n10725),.dinb(n10722),.dout(n10726),.clk(gclk));
	jand g10453(.dina(n10726),.dinb(n10721),.dout(n10727),.clk(gclk));
	jxor g10454(.dina(n10727),.dinb(w_n9780_0[1]),.dout(n10728),.clk(gclk));
	jor g10455(.dina(w_n10728_0[1]),.dinb(w_n10720_0[1]),.dout(n10729),.clk(gclk));
	jand g10456(.dina(n10729),.dinb(w_n10718_0[1]),.dout(n10730),.clk(gclk));
	jor g10457(.dina(w_n10730_0[2]),.dinb(w_n9769_13[0]),.dout(n10731),.clk(gclk));
	jand g10458(.dina(w_n10730_0[1]),.dinb(w_n9769_12[2]),.dout(n10732),.clk(gclk));
	jxor g10459(.dina(w_n10223_0[0]),.dinb(w_n9774_16[1]),.dout(n10733),.clk(gclk));
	jor g10460(.dina(n10733),.dinb(w_n10701_24[2]),.dout(n10734),.clk(gclk));
	jxor g10461(.dina(n10734),.dinb(w_n10226_0[0]),.dout(n10735),.clk(gclk));
	jor g10462(.dina(w_n10735_0[1]),.dinb(n10732),.dout(n10736),.clk(gclk));
	jand g10463(.dina(w_n10736_0[1]),.dinb(w_n10731_0[1]),.dout(n10737),.clk(gclk));
	jor g10464(.dina(n10737),.dinb(w_n8898_17[2]),.dout(n10738),.clk(gclk));
	jnot g10465(.din(w_n10232_0[0]),.dout(n10739),.clk(gclk));
	jor g10466(.dina(n10739),.dinb(w_n10230_0[0]),.dout(n10740),.clk(gclk));
	jor g10467(.dina(n10740),.dinb(w_n10701_24[1]),.dout(n10741),.clk(gclk));
	jxor g10468(.dina(n10741),.dinb(w_n10241_0[0]),.dout(n10742),.clk(gclk));
	jand g10469(.dina(w_n10731_0[0]),.dinb(w_n8898_17[1]),.dout(n10743),.clk(gclk));
	jand g10470(.dina(n10743),.dinb(w_n10736_0[0]),.dout(n10744),.clk(gclk));
	jor g10471(.dina(w_n10744_0[1]),.dinb(w_n10742_0[1]),.dout(n10745),.clk(gclk));
	jand g10472(.dina(w_n10745_0[1]),.dinb(w_n10738_0[1]),.dout(n10746),.clk(gclk));
	jor g10473(.dina(w_n10746_0[2]),.dinb(w_n8893_13[1]),.dout(n10747),.clk(gclk));
	jand g10474(.dina(w_n10746_0[1]),.dinb(w_n8893_13[0]),.dout(n10748),.clk(gclk));
	jxor g10475(.dina(w_n10243_0[0]),.dinb(w_n8898_17[0]),.dout(n10749),.clk(gclk));
	jor g10476(.dina(n10749),.dinb(w_n10701_24[0]),.dout(n10750),.clk(gclk));
	jxor g10477(.dina(n10750),.dinb(w_n10248_0[0]),.dout(n10751),.clk(gclk));
	jnot g10478(.din(w_n10751_0[1]),.dout(n10752),.clk(gclk));
	jor g10479(.dina(n10752),.dinb(n10748),.dout(n10753),.clk(gclk));
	jand g10480(.dina(w_n10753_0[1]),.dinb(w_n10747_0[1]),.dout(n10754),.clk(gclk));
	jor g10481(.dina(n10754),.dinb(w_n8058_17[1]),.dout(n10755),.clk(gclk));
	jand g10482(.dina(w_n10747_0[0]),.dinb(w_n8058_17[0]),.dout(n10756),.clk(gclk));
	jand g10483(.dina(n10756),.dinb(w_n10753_0[0]),.dout(n10757),.clk(gclk));
	jnot g10484(.din(w_n10252_0[0]),.dout(n10758),.clk(gclk));
	jnot g10485(.din(w_n10701_23[2]),.dout(asqrt_fa_20),.clk(gclk));
	jand g10486(.dina(w_asqrt19_18),.dinb(n10758),.dout(n10760),.clk(gclk));
	jand g10487(.dina(w_n10760_0[1]),.dinb(w_n10259_0[0]),.dout(n10761),.clk(gclk));
	jor g10488(.dina(n10761),.dinb(w_n10257_0[0]),.dout(n10762),.clk(gclk));
	jand g10489(.dina(w_n10760_0[0]),.dinb(w_n10260_0[0]),.dout(n10763),.clk(gclk));
	jnot g10490(.din(n10763),.dout(n10764),.clk(gclk));
	jand g10491(.dina(n10764),.dinb(n10762),.dout(n10765),.clk(gclk));
	jnot g10492(.din(n10765),.dout(n10766),.clk(gclk));
	jor g10493(.dina(w_n10766_0[1]),.dinb(w_n10757_0[1]),.dout(n10767),.clk(gclk));
	jand g10494(.dina(n10767),.dinb(w_n10755_0[1]),.dout(n10768),.clk(gclk));
	jor g10495(.dina(w_n10768_0[2]),.dinb(w_n8053_13[1]),.dout(n10769),.clk(gclk));
	jand g10496(.dina(w_n10768_0[1]),.dinb(w_n8053_13[0]),.dout(n10770),.clk(gclk));
	jnot g10497(.din(w_n10267_0[0]),.dout(n10771),.clk(gclk));
	jxor g10498(.dina(w_n10261_0[0]),.dinb(w_n8058_16[2]),.dout(n10772),.clk(gclk));
	jor g10499(.dina(n10772),.dinb(w_n10701_23[1]),.dout(n10773),.clk(gclk));
	jxor g10500(.dina(n10773),.dinb(n10771),.dout(n10774),.clk(gclk));
	jnot g10501(.din(w_n10774_0[1]),.dout(n10775),.clk(gclk));
	jor g10502(.dina(n10775),.dinb(n10770),.dout(n10776),.clk(gclk));
	jand g10503(.dina(w_n10776_0[1]),.dinb(w_n10769_0[1]),.dout(n10777),.clk(gclk));
	jor g10504(.dina(n10777),.dinb(w_n7265_17[2]),.dout(n10778),.clk(gclk));
	jnot g10505(.din(w_n10272_0[0]),.dout(n10779),.clk(gclk));
	jor g10506(.dina(n10779),.dinb(w_n10270_0[0]),.dout(n10780),.clk(gclk));
	jor g10507(.dina(n10780),.dinb(w_n10701_23[0]),.dout(n10781),.clk(gclk));
	jxor g10508(.dina(n10781),.dinb(w_n10281_0[0]),.dout(n10782),.clk(gclk));
	jand g10509(.dina(w_n10769_0[0]),.dinb(w_n7265_17[1]),.dout(n10783),.clk(gclk));
	jand g10510(.dina(n10783),.dinb(w_n10776_0[0]),.dout(n10784),.clk(gclk));
	jor g10511(.dina(w_n10784_0[1]),.dinb(w_n10782_0[1]),.dout(n10785),.clk(gclk));
	jand g10512(.dina(w_n10785_0[1]),.dinb(w_n10778_0[1]),.dout(n10786),.clk(gclk));
	jor g10513(.dina(w_n10786_0[2]),.dinb(w_n7260_14[0]),.dout(n10787),.clk(gclk));
	jand g10514(.dina(w_n10786_0[1]),.dinb(w_n7260_13[2]),.dout(n10788),.clk(gclk));
	jnot g10515(.din(w_n10288_0[0]),.dout(n10789),.clk(gclk));
	jxor g10516(.dina(w_n10283_0[0]),.dinb(w_n7265_17[0]),.dout(n10790),.clk(gclk));
	jor g10517(.dina(n10790),.dinb(w_n10701_22[2]),.dout(n10791),.clk(gclk));
	jxor g10518(.dina(n10791),.dinb(n10789),.dout(n10792),.clk(gclk));
	jnot g10519(.din(n10792),.dout(n10793),.clk(gclk));
	jor g10520(.dina(w_n10793_0[1]),.dinb(n10788),.dout(n10794),.clk(gclk));
	jand g10521(.dina(w_n10794_0[1]),.dinb(w_n10787_0[1]),.dout(n10795),.clk(gclk));
	jor g10522(.dina(n10795),.dinb(w_n6505_17[1]),.dout(n10796),.clk(gclk));
	jand g10523(.dina(w_n10787_0[0]),.dinb(w_n6505_17[0]),.dout(n10797),.clk(gclk));
	jand g10524(.dina(n10797),.dinb(w_n10794_0[0]),.dout(n10798),.clk(gclk));
	jnot g10525(.din(w_n10291_0[0]),.dout(n10799),.clk(gclk));
	jand g10526(.dina(w_asqrt19_17[2]),.dinb(n10799),.dout(n10800),.clk(gclk));
	jand g10527(.dina(w_n10800_0[1]),.dinb(w_n10298_0[0]),.dout(n10801),.clk(gclk));
	jor g10528(.dina(n10801),.dinb(w_n10296_0[0]),.dout(n10802),.clk(gclk));
	jand g10529(.dina(w_n10800_0[0]),.dinb(w_n10299_0[0]),.dout(n10803),.clk(gclk));
	jnot g10530(.din(n10803),.dout(n10804),.clk(gclk));
	jand g10531(.dina(n10804),.dinb(n10802),.dout(n10805),.clk(gclk));
	jnot g10532(.din(n10805),.dout(n10806),.clk(gclk));
	jor g10533(.dina(w_n10806_0[1]),.dinb(w_n10798_0[1]),.dout(n10807),.clk(gclk));
	jand g10534(.dina(n10807),.dinb(w_n10796_0[1]),.dout(n10808),.clk(gclk));
	jor g10535(.dina(w_n10808_0[1]),.dinb(w_n6500_14[0]),.dout(n10809),.clk(gclk));
	jxor g10536(.dina(w_n10300_0[0]),.dinb(w_n6505_16[2]),.dout(n10810),.clk(gclk));
	jor g10537(.dina(n10810),.dinb(w_n10701_22[1]),.dout(n10811),.clk(gclk));
	jxor g10538(.dina(n10811),.dinb(w_n10305_0[0]),.dout(n10812),.clk(gclk));
	jand g10539(.dina(w_n10808_0[0]),.dinb(w_n6500_13[2]),.dout(n10813),.clk(gclk));
	jor g10540(.dina(w_n10813_0[1]),.dinb(w_n10812_0[1]),.dout(n10814),.clk(gclk));
	jand g10541(.dina(w_n10814_0[2]),.dinb(w_n10809_0[2]),.dout(n10815),.clk(gclk));
	jor g10542(.dina(n10815),.dinb(w_n5793_17[2]),.dout(n10816),.clk(gclk));
	jnot g10543(.din(w_n10310_0[0]),.dout(n10817),.clk(gclk));
	jor g10544(.dina(n10817),.dinb(w_n10308_0[0]),.dout(n10818),.clk(gclk));
	jor g10545(.dina(n10818),.dinb(w_n10701_22[0]),.dout(n10819),.clk(gclk));
	jxor g10546(.dina(n10819),.dinb(w_n10319_0[0]),.dout(n10820),.clk(gclk));
	jand g10547(.dina(w_n10809_0[1]),.dinb(w_n5793_17[1]),.dout(n10821),.clk(gclk));
	jand g10548(.dina(n10821),.dinb(w_n10814_0[1]),.dout(n10822),.clk(gclk));
	jor g10549(.dina(w_n10822_0[1]),.dinb(w_n10820_0[1]),.dout(n10823),.clk(gclk));
	jand g10550(.dina(w_n10823_0[1]),.dinb(w_n10816_0[1]),.dout(n10824),.clk(gclk));
	jor g10551(.dina(w_n10824_0[2]),.dinb(w_n5788_14[2]),.dout(n10825),.clk(gclk));
	jand g10552(.dina(w_n10824_0[1]),.dinb(w_n5788_14[1]),.dout(n10826),.clk(gclk));
	jnot g10553(.din(w_n10322_0[0]),.dout(n10827),.clk(gclk));
	jand g10554(.dina(w_asqrt19_17[1]),.dinb(n10827),.dout(n10828),.clk(gclk));
	jand g10555(.dina(w_n10828_0[1]),.dinb(w_n10327_0[0]),.dout(n10829),.clk(gclk));
	jor g10556(.dina(n10829),.dinb(w_n10326_0[0]),.dout(n10830),.clk(gclk));
	jand g10557(.dina(w_n10828_0[0]),.dinb(w_n10328_0[0]),.dout(n10831),.clk(gclk));
	jnot g10558(.din(n10831),.dout(n10832),.clk(gclk));
	jand g10559(.dina(n10832),.dinb(n10830),.dout(n10833),.clk(gclk));
	jnot g10560(.din(n10833),.dout(n10834),.clk(gclk));
	jor g10561(.dina(w_n10834_0[1]),.dinb(n10826),.dout(n10835),.clk(gclk));
	jand g10562(.dina(w_n10835_0[1]),.dinb(w_n10825_0[1]),.dout(n10836),.clk(gclk));
	jor g10563(.dina(n10836),.dinb(w_n5121_17[2]),.dout(n10837),.clk(gclk));
	jand g10564(.dina(w_n10825_0[0]),.dinb(w_n5121_17[1]),.dout(n10838),.clk(gclk));
	jand g10565(.dina(n10838),.dinb(w_n10835_0[0]),.dout(n10839),.clk(gclk));
	jnot g10566(.din(w_n10330_0[0]),.dout(n10840),.clk(gclk));
	jand g10567(.dina(w_asqrt19_17[0]),.dinb(n10840),.dout(n10841),.clk(gclk));
	jand g10568(.dina(w_n10841_0[1]),.dinb(w_n10337_0[0]),.dout(n10842),.clk(gclk));
	jor g10569(.dina(n10842),.dinb(w_n10335_0[0]),.dout(n10843),.clk(gclk));
	jand g10570(.dina(w_n10841_0[0]),.dinb(w_n10338_0[0]),.dout(n10844),.clk(gclk));
	jnot g10571(.din(n10844),.dout(n10845),.clk(gclk));
	jand g10572(.dina(n10845),.dinb(n10843),.dout(n10846),.clk(gclk));
	jnot g10573(.din(n10846),.dout(n10847),.clk(gclk));
	jor g10574(.dina(w_n10847_0[1]),.dinb(w_n10839_0[1]),.dout(n10848),.clk(gclk));
	jand g10575(.dina(n10848),.dinb(w_n10837_0[1]),.dout(n10849),.clk(gclk));
	jor g10576(.dina(w_n10849_0[1]),.dinb(w_n5116_14[2]),.dout(n10850),.clk(gclk));
	jxor g10577(.dina(w_n10339_0[0]),.dinb(w_n5121_17[0]),.dout(n10851),.clk(gclk));
	jor g10578(.dina(n10851),.dinb(w_n10701_21[2]),.dout(n10852),.clk(gclk));
	jxor g10579(.dina(n10852),.dinb(w_n10350_0[0]),.dout(n10853),.clk(gclk));
	jand g10580(.dina(w_n10849_0[0]),.dinb(w_n5116_14[1]),.dout(n10854),.clk(gclk));
	jor g10581(.dina(w_n10854_0[1]),.dinb(w_n10853_0[1]),.dout(n10855),.clk(gclk));
	jand g10582(.dina(w_n10855_0[2]),.dinb(w_n10850_0[2]),.dout(n10856),.clk(gclk));
	jor g10583(.dina(n10856),.dinb(w_n4499_18[1]),.dout(n10857),.clk(gclk));
	jnot g10584(.din(w_n10355_0[0]),.dout(n10858),.clk(gclk));
	jor g10585(.dina(n10858),.dinb(w_n10353_0[0]),.dout(n10859),.clk(gclk));
	jor g10586(.dina(n10859),.dinb(w_n10701_21[1]),.dout(n10860),.clk(gclk));
	jxor g10587(.dina(n10860),.dinb(w_n10364_0[0]),.dout(n10861),.clk(gclk));
	jand g10588(.dina(w_n10850_0[1]),.dinb(w_n4499_18[0]),.dout(n10862),.clk(gclk));
	jand g10589(.dina(n10862),.dinb(w_n10855_0[1]),.dout(n10863),.clk(gclk));
	jor g10590(.dina(w_n10863_0[1]),.dinb(w_n10861_0[1]),.dout(n10864),.clk(gclk));
	jand g10591(.dina(w_n10864_0[1]),.dinb(w_n10857_0[1]),.dout(n10865),.clk(gclk));
	jor g10592(.dina(w_n10865_0[2]),.dinb(w_n4494_15[2]),.dout(n10866),.clk(gclk));
	jand g10593(.dina(w_n10865_0[1]),.dinb(w_n4494_15[1]),.dout(n10867),.clk(gclk));
	jnot g10594(.din(w_n10367_0[0]),.dout(n10868),.clk(gclk));
	jand g10595(.dina(w_asqrt19_16[2]),.dinb(n10868),.dout(n10869),.clk(gclk));
	jand g10596(.dina(w_n10869_0[1]),.dinb(w_n10372_0[0]),.dout(n10870),.clk(gclk));
	jor g10597(.dina(n10870),.dinb(w_n10371_0[0]),.dout(n10871),.clk(gclk));
	jand g10598(.dina(w_n10869_0[0]),.dinb(w_n10373_0[0]),.dout(n10872),.clk(gclk));
	jnot g10599(.din(n10872),.dout(n10873),.clk(gclk));
	jand g10600(.dina(n10873),.dinb(n10871),.dout(n10874),.clk(gclk));
	jnot g10601(.din(n10874),.dout(n10875),.clk(gclk));
	jor g10602(.dina(w_n10875_0[1]),.dinb(n10867),.dout(n10876),.clk(gclk));
	jand g10603(.dina(w_n10876_0[1]),.dinb(w_n10866_0[1]),.dout(n10877),.clk(gclk));
	jor g10604(.dina(n10877),.dinb(w_n3912_18[1]),.dout(n10878),.clk(gclk));
	jand g10605(.dina(w_n10866_0[0]),.dinb(w_n3912_18[0]),.dout(n10879),.clk(gclk));
	jand g10606(.dina(n10879),.dinb(w_n10876_0[0]),.dout(n10880),.clk(gclk));
	jnot g10607(.din(w_n10375_0[0]),.dout(n10881),.clk(gclk));
	jand g10608(.dina(w_asqrt19_16[1]),.dinb(n10881),.dout(n10882),.clk(gclk));
	jand g10609(.dina(w_n10882_0[1]),.dinb(w_n10382_0[0]),.dout(n10883),.clk(gclk));
	jor g10610(.dina(n10883),.dinb(w_n10380_0[0]),.dout(n10884),.clk(gclk));
	jand g10611(.dina(w_n10882_0[0]),.dinb(w_n10383_0[0]),.dout(n10885),.clk(gclk));
	jnot g10612(.din(n10885),.dout(n10886),.clk(gclk));
	jand g10613(.dina(n10886),.dinb(n10884),.dout(n10887),.clk(gclk));
	jnot g10614(.din(n10887),.dout(n10888),.clk(gclk));
	jor g10615(.dina(w_n10888_0[1]),.dinb(w_n10880_0[1]),.dout(n10889),.clk(gclk));
	jand g10616(.dina(n10889),.dinb(w_n10878_0[1]),.dout(n10890),.clk(gclk));
	jor g10617(.dina(w_n10890_0[1]),.dinb(w_n3907_15[2]),.dout(n10891),.clk(gclk));
	jxor g10618(.dina(w_n10384_0[0]),.dinb(w_n3912_17[2]),.dout(n10892),.clk(gclk));
	jor g10619(.dina(n10892),.dinb(w_n10701_21[0]),.dout(n10893),.clk(gclk));
	jxor g10620(.dina(n10893),.dinb(w_n10395_0[0]),.dout(n10894),.clk(gclk));
	jand g10621(.dina(w_n10890_0[0]),.dinb(w_n3907_15[1]),.dout(n10895),.clk(gclk));
	jor g10622(.dina(w_n10895_0[1]),.dinb(w_n10894_0[1]),.dout(n10896),.clk(gclk));
	jand g10623(.dina(w_n10896_0[2]),.dinb(w_n10891_0[2]),.dout(n10897),.clk(gclk));
	jor g10624(.dina(n10897),.dinb(w_n3376_19[0]),.dout(n10898),.clk(gclk));
	jnot g10625(.din(w_n10400_0[0]),.dout(n10899),.clk(gclk));
	jor g10626(.dina(n10899),.dinb(w_n10398_0[0]),.dout(n10900),.clk(gclk));
	jor g10627(.dina(n10900),.dinb(w_n10701_20[2]),.dout(n10901),.clk(gclk));
	jxor g10628(.dina(n10901),.dinb(w_n10409_0[0]),.dout(n10902),.clk(gclk));
	jand g10629(.dina(w_n10891_0[1]),.dinb(w_n3376_18[2]),.dout(n10903),.clk(gclk));
	jand g10630(.dina(n10903),.dinb(w_n10896_0[1]),.dout(n10904),.clk(gclk));
	jor g10631(.dina(w_n10904_0[1]),.dinb(w_n10902_0[1]),.dout(n10905),.clk(gclk));
	jand g10632(.dina(w_n10905_0[1]),.dinb(w_n10898_0[1]),.dout(n10906),.clk(gclk));
	jor g10633(.dina(w_n10906_0[2]),.dinb(w_n3371_16[1]),.dout(n10907),.clk(gclk));
	jand g10634(.dina(w_n10906_0[1]),.dinb(w_n3371_16[0]),.dout(n10908),.clk(gclk));
	jnot g10635(.din(w_n10412_0[0]),.dout(n10909),.clk(gclk));
	jand g10636(.dina(w_asqrt19_16[0]),.dinb(n10909),.dout(n10910),.clk(gclk));
	jand g10637(.dina(w_n10910_0[1]),.dinb(w_n10417_0[0]),.dout(n10911),.clk(gclk));
	jor g10638(.dina(n10911),.dinb(w_n10416_0[0]),.dout(n10912),.clk(gclk));
	jand g10639(.dina(w_n10910_0[0]),.dinb(w_n10418_0[0]),.dout(n10913),.clk(gclk));
	jnot g10640(.din(n10913),.dout(n10914),.clk(gclk));
	jand g10641(.dina(n10914),.dinb(n10912),.dout(n10915),.clk(gclk));
	jnot g10642(.din(n10915),.dout(n10916),.clk(gclk));
	jor g10643(.dina(w_n10916_0[1]),.dinb(n10908),.dout(n10917),.clk(gclk));
	jand g10644(.dina(w_n10917_0[1]),.dinb(w_n10907_0[1]),.dout(n10918),.clk(gclk));
	jor g10645(.dina(n10918),.dinb(w_n2875_19[0]),.dout(n10919),.clk(gclk));
	jand g10646(.dina(w_n10907_0[0]),.dinb(w_n2875_18[2]),.dout(n10920),.clk(gclk));
	jand g10647(.dina(n10920),.dinb(w_n10917_0[0]),.dout(n10921),.clk(gclk));
	jnot g10648(.din(w_n10420_0[0]),.dout(n10922),.clk(gclk));
	jand g10649(.dina(w_asqrt19_15[2]),.dinb(n10922),.dout(n10923),.clk(gclk));
	jand g10650(.dina(w_n10923_0[1]),.dinb(w_n10427_0[0]),.dout(n10924),.clk(gclk));
	jor g10651(.dina(n10924),.dinb(w_n10425_0[0]),.dout(n10925),.clk(gclk));
	jand g10652(.dina(w_n10923_0[0]),.dinb(w_n10428_0[0]),.dout(n10926),.clk(gclk));
	jnot g10653(.din(n10926),.dout(n10927),.clk(gclk));
	jand g10654(.dina(n10927),.dinb(n10925),.dout(n10928),.clk(gclk));
	jnot g10655(.din(n10928),.dout(n10929),.clk(gclk));
	jor g10656(.dina(w_n10929_0[1]),.dinb(w_n10921_0[1]),.dout(n10930),.clk(gclk));
	jand g10657(.dina(n10930),.dinb(w_n10919_0[1]),.dout(n10931),.clk(gclk));
	jor g10658(.dina(w_n10931_0[1]),.dinb(w_n2870_16[1]),.dout(n10932),.clk(gclk));
	jxor g10659(.dina(w_n10429_0[0]),.dinb(w_n2875_18[1]),.dout(n10933),.clk(gclk));
	jor g10660(.dina(n10933),.dinb(w_n10701_20[1]),.dout(n10934),.clk(gclk));
	jxor g10661(.dina(n10934),.dinb(w_n10440_0[0]),.dout(n10935),.clk(gclk));
	jand g10662(.dina(w_n10931_0[0]),.dinb(w_n2870_16[0]),.dout(n10936),.clk(gclk));
	jor g10663(.dina(w_n10936_0[1]),.dinb(w_n10935_0[1]),.dout(n10937),.clk(gclk));
	jand g10664(.dina(w_n10937_0[2]),.dinb(w_n10932_0[2]),.dout(n10938),.clk(gclk));
	jor g10665(.dina(n10938),.dinb(w_n2425_19[1]),.dout(n10939),.clk(gclk));
	jand g10666(.dina(w_n10932_0[1]),.dinb(w_n2425_19[0]),.dout(n10940),.clk(gclk));
	jand g10667(.dina(n10940),.dinb(w_n10937_0[1]),.dout(n10941),.clk(gclk));
	jnot g10668(.din(w_n10443_0[0]),.dout(n10942),.clk(gclk));
	jand g10669(.dina(w_asqrt19_15[1]),.dinb(n10942),.dout(n10943),.clk(gclk));
	jand g10670(.dina(w_n10943_0[1]),.dinb(w_n10450_0[0]),.dout(n10944),.clk(gclk));
	jor g10671(.dina(n10944),.dinb(w_n10448_0[0]),.dout(n10945),.clk(gclk));
	jand g10672(.dina(w_n10943_0[0]),.dinb(w_n10451_0[0]),.dout(n10946),.clk(gclk));
	jnot g10673(.din(n10946),.dout(n10947),.clk(gclk));
	jand g10674(.dina(n10947),.dinb(n10945),.dout(n10948),.clk(gclk));
	jnot g10675(.din(n10948),.dout(n10949),.clk(gclk));
	jor g10676(.dina(w_n10949_0[1]),.dinb(w_n10941_0[1]),.dout(n10950),.clk(gclk));
	jand g10677(.dina(n10950),.dinb(w_n10939_0[1]),.dout(n10951),.clk(gclk));
	jor g10678(.dina(w_n10951_0[2]),.dinb(w_n2420_17[1]),.dout(n10952),.clk(gclk));
	jand g10679(.dina(w_n10951_0[1]),.dinb(w_n2420_17[0]),.dout(n10953),.clk(gclk));
	jor g10680(.dina(n10953),.dinb(w_n10704_0[1]),.dout(n10954),.clk(gclk));
	jand g10681(.dina(w_n10954_0[1]),.dinb(w_n10952_0[1]),.dout(n10955),.clk(gclk));
	jor g10682(.dina(n10955),.dinb(w_n2010_19[2]),.dout(n10956),.clk(gclk));
	jnot g10683(.din(w_n10459_0[0]),.dout(n10957),.clk(gclk));
	jor g10684(.dina(n10957),.dinb(w_n10457_0[0]),.dout(n10958),.clk(gclk));
	jor g10685(.dina(n10958),.dinb(w_n10701_20[0]),.dout(n10959),.clk(gclk));
	jxor g10686(.dina(n10959),.dinb(w_n10468_0[0]),.dout(n10960),.clk(gclk));
	jand g10687(.dina(w_n10952_0[0]),.dinb(w_n2010_19[1]),.dout(n10961),.clk(gclk));
	jand g10688(.dina(n10961),.dinb(w_n10954_0[0]),.dout(n10962),.clk(gclk));
	jor g10689(.dina(w_n10962_0[1]),.dinb(w_n10960_0[1]),.dout(n10963),.clk(gclk));
	jand g10690(.dina(w_n10963_0[1]),.dinb(w_n10956_0[1]),.dout(n10964),.clk(gclk));
	jor g10691(.dina(w_n10964_0[1]),.dinb(w_n2005_17[1]),.dout(n10965),.clk(gclk));
	jxor g10692(.dina(w_n10470_0[0]),.dinb(w_n2010_19[0]),.dout(n10966),.clk(gclk));
	jor g10693(.dina(n10966),.dinb(w_n10701_19[2]),.dout(n10967),.clk(gclk));
	jxor g10694(.dina(n10967),.dinb(w_n10481_0[0]),.dout(n10968),.clk(gclk));
	jand g10695(.dina(w_n10964_0[0]),.dinb(w_n2005_17[0]),.dout(n10969),.clk(gclk));
	jor g10696(.dina(w_n10969_0[1]),.dinb(w_n10968_0[1]),.dout(n10970),.clk(gclk));
	jand g10697(.dina(w_n10970_0[2]),.dinb(w_n10965_0[2]),.dout(n10971),.clk(gclk));
	jor g10698(.dina(n10971),.dinb(w_n1646_20[1]),.dout(n10972),.clk(gclk));
	jnot g10699(.din(w_n10486_0[0]),.dout(n10973),.clk(gclk));
	jor g10700(.dina(n10973),.dinb(w_n10484_0[0]),.dout(n10974),.clk(gclk));
	jor g10701(.dina(n10974),.dinb(w_n10701_19[1]),.dout(n10975),.clk(gclk));
	jxor g10702(.dina(n10975),.dinb(w_n10495_0[0]),.dout(n10976),.clk(gclk));
	jand g10703(.dina(w_n10965_0[1]),.dinb(w_n1646_20[0]),.dout(n10977),.clk(gclk));
	jand g10704(.dina(n10977),.dinb(w_n10970_0[1]),.dout(n10978),.clk(gclk));
	jor g10705(.dina(w_n10978_0[1]),.dinb(w_n10976_0[1]),.dout(n10979),.clk(gclk));
	jand g10706(.dina(w_n10979_0[1]),.dinb(w_n10972_0[1]),.dout(n10980),.clk(gclk));
	jor g10707(.dina(w_n10980_0[2]),.dinb(w_n1641_18[0]),.dout(n10981),.clk(gclk));
	jand g10708(.dina(w_n10980_0[1]),.dinb(w_n1641_17[2]),.dout(n10982),.clk(gclk));
	jnot g10709(.din(w_n10498_0[0]),.dout(n10983),.clk(gclk));
	jand g10710(.dina(w_asqrt19_15[0]),.dinb(n10983),.dout(n10984),.clk(gclk));
	jand g10711(.dina(w_n10984_0[1]),.dinb(w_n10503_0[0]),.dout(n10985),.clk(gclk));
	jor g10712(.dina(n10985),.dinb(w_n10502_0[0]),.dout(n10986),.clk(gclk));
	jand g10713(.dina(w_n10984_0[0]),.dinb(w_n10504_0[0]),.dout(n10987),.clk(gclk));
	jnot g10714(.din(n10987),.dout(n10988),.clk(gclk));
	jand g10715(.dina(n10988),.dinb(n10986),.dout(n10989),.clk(gclk));
	jnot g10716(.din(n10989),.dout(n10990),.clk(gclk));
	jor g10717(.dina(w_n10990_0[1]),.dinb(n10982),.dout(n10991),.clk(gclk));
	jand g10718(.dina(w_n10991_0[1]),.dinb(w_n10981_0[1]),.dout(n10992),.clk(gclk));
	jor g10719(.dina(n10992),.dinb(w_n1317_20[1]),.dout(n10993),.clk(gclk));
	jand g10720(.dina(w_n10981_0[0]),.dinb(w_n1317_20[0]),.dout(n10994),.clk(gclk));
	jand g10721(.dina(n10994),.dinb(w_n10991_0[0]),.dout(n10995),.clk(gclk));
	jnot g10722(.din(w_n10506_0[0]),.dout(n10996),.clk(gclk));
	jand g10723(.dina(w_asqrt19_14[2]),.dinb(n10996),.dout(n10997),.clk(gclk));
	jand g10724(.dina(w_n10997_0[1]),.dinb(w_n10513_0[0]),.dout(n10998),.clk(gclk));
	jor g10725(.dina(n10998),.dinb(w_n10511_0[0]),.dout(n10999),.clk(gclk));
	jand g10726(.dina(w_n10997_0[0]),.dinb(w_n10514_0[0]),.dout(n11000),.clk(gclk));
	jnot g10727(.din(n11000),.dout(n11001),.clk(gclk));
	jand g10728(.dina(n11001),.dinb(n10999),.dout(n11002),.clk(gclk));
	jnot g10729(.din(n11002),.dout(n11003),.clk(gclk));
	jor g10730(.dina(w_n11003_0[1]),.dinb(w_n10995_0[1]),.dout(n11004),.clk(gclk));
	jand g10731(.dina(n11004),.dinb(w_n10993_0[1]),.dout(n11005),.clk(gclk));
	jor g10732(.dina(w_n11005_0[1]),.dinb(w_n1312_18[0]),.dout(n11006),.clk(gclk));
	jxor g10733(.dina(w_n10515_0[0]),.dinb(w_n1317_19[2]),.dout(n11007),.clk(gclk));
	jor g10734(.dina(n11007),.dinb(w_n10701_19[0]),.dout(n11008),.clk(gclk));
	jxor g10735(.dina(n11008),.dinb(w_n10526_0[0]),.dout(n11009),.clk(gclk));
	jand g10736(.dina(w_n11005_0[0]),.dinb(w_n1312_17[2]),.dout(n11010),.clk(gclk));
	jor g10737(.dina(w_n11010_0[1]),.dinb(w_n11009_0[1]),.dout(n11011),.clk(gclk));
	jand g10738(.dina(w_n11011_0[2]),.dinb(w_n11006_0[2]),.dout(n11012),.clk(gclk));
	jor g10739(.dina(n11012),.dinb(w_n1039_20[2]),.dout(n11013),.clk(gclk));
	jnot g10740(.din(w_n10531_0[0]),.dout(n11014),.clk(gclk));
	jor g10741(.dina(n11014),.dinb(w_n10529_0[0]),.dout(n11015),.clk(gclk));
	jor g10742(.dina(n11015),.dinb(w_n10701_18[2]),.dout(n11016),.clk(gclk));
	jxor g10743(.dina(n11016),.dinb(w_n10540_0[0]),.dout(n11017),.clk(gclk));
	jand g10744(.dina(w_n11006_0[1]),.dinb(w_n1039_20[1]),.dout(n11018),.clk(gclk));
	jand g10745(.dina(n11018),.dinb(w_n11011_0[1]),.dout(n11019),.clk(gclk));
	jor g10746(.dina(w_n11019_0[1]),.dinb(w_n11017_0[1]),.dout(n11020),.clk(gclk));
	jand g10747(.dina(w_n11020_0[1]),.dinb(w_n11013_0[1]),.dout(n11021),.clk(gclk));
	jor g10748(.dina(w_n11021_0[2]),.dinb(w_n1034_19[0]),.dout(n11022),.clk(gclk));
	jand g10749(.dina(w_n11021_0[1]),.dinb(w_n1034_18[2]),.dout(n11023),.clk(gclk));
	jnot g10750(.din(w_n10543_0[0]),.dout(n11024),.clk(gclk));
	jand g10751(.dina(w_asqrt19_14[1]),.dinb(n11024),.dout(n11025),.clk(gclk));
	jand g10752(.dina(w_n11025_0[1]),.dinb(w_n10548_0[0]),.dout(n11026),.clk(gclk));
	jor g10753(.dina(n11026),.dinb(w_n10547_0[0]),.dout(n11027),.clk(gclk));
	jand g10754(.dina(w_n11025_0[0]),.dinb(w_n10549_0[0]),.dout(n11028),.clk(gclk));
	jnot g10755(.din(n11028),.dout(n11029),.clk(gclk));
	jand g10756(.dina(n11029),.dinb(n11027),.dout(n11030),.clk(gclk));
	jnot g10757(.din(n11030),.dout(n11031),.clk(gclk));
	jor g10758(.dina(w_n11031_0[1]),.dinb(n11023),.dout(n11032),.clk(gclk));
	jand g10759(.dina(w_n11032_0[1]),.dinb(w_n11022_0[1]),.dout(n11033),.clk(gclk));
	jor g10760(.dina(n11033),.dinb(w_n796_20[2]),.dout(n11034),.clk(gclk));
	jand g10761(.dina(w_n11022_0[0]),.dinb(w_n796_20[1]),.dout(n11035),.clk(gclk));
	jand g10762(.dina(n11035),.dinb(w_n11032_0[0]),.dout(n11036),.clk(gclk));
	jnot g10763(.din(w_n10551_0[0]),.dout(n11037),.clk(gclk));
	jand g10764(.dina(w_asqrt19_14[0]),.dinb(n11037),.dout(n11038),.clk(gclk));
	jand g10765(.dina(w_n11038_0[1]),.dinb(w_n10558_0[0]),.dout(n11039),.clk(gclk));
	jor g10766(.dina(n11039),.dinb(w_n10556_0[0]),.dout(n11040),.clk(gclk));
	jand g10767(.dina(w_n11038_0[0]),.dinb(w_n10559_0[0]),.dout(n11041),.clk(gclk));
	jnot g10768(.din(n11041),.dout(n11042),.clk(gclk));
	jand g10769(.dina(n11042),.dinb(n11040),.dout(n11043),.clk(gclk));
	jnot g10770(.din(n11043),.dout(n11044),.clk(gclk));
	jor g10771(.dina(w_n11044_0[1]),.dinb(w_n11036_0[1]),.dout(n11045),.clk(gclk));
	jand g10772(.dina(n11045),.dinb(w_n11034_0[1]),.dout(n11046),.clk(gclk));
	jor g10773(.dina(w_n11046_0[1]),.dinb(w_n791_19[0]),.dout(n11047),.clk(gclk));
	jxor g10774(.dina(w_n10560_0[0]),.dinb(w_n796_20[0]),.dout(n11048),.clk(gclk));
	jor g10775(.dina(n11048),.dinb(w_n10701_18[1]),.dout(n11049),.clk(gclk));
	jxor g10776(.dina(n11049),.dinb(w_n10571_0[0]),.dout(n11050),.clk(gclk));
	jand g10777(.dina(w_n11046_0[0]),.dinb(w_n791_18[2]),.dout(n11051),.clk(gclk));
	jor g10778(.dina(w_n11051_0[1]),.dinb(w_n11050_0[1]),.dout(n11052),.clk(gclk));
	jand g10779(.dina(w_n11052_0[2]),.dinb(w_n11047_0[2]),.dout(n11053),.clk(gclk));
	jor g10780(.dina(n11053),.dinb(w_n595_21[0]),.dout(n11054),.clk(gclk));
	jnot g10781(.din(w_n10576_0[0]),.dout(n11055),.clk(gclk));
	jor g10782(.dina(n11055),.dinb(w_n10574_0[0]),.dout(n11056),.clk(gclk));
	jor g10783(.dina(n11056),.dinb(w_n10701_18[0]),.dout(n11057),.clk(gclk));
	jxor g10784(.dina(n11057),.dinb(w_n10585_0[0]),.dout(n11058),.clk(gclk));
	jand g10785(.dina(w_n11047_0[1]),.dinb(w_n595_20[2]),.dout(n11059),.clk(gclk));
	jand g10786(.dina(n11059),.dinb(w_n11052_0[1]),.dout(n11060),.clk(gclk));
	jor g10787(.dina(w_n11060_0[1]),.dinb(w_n11058_0[1]),.dout(n11061),.clk(gclk));
	jand g10788(.dina(w_n11061_0[1]),.dinb(w_n11054_0[1]),.dout(n11062),.clk(gclk));
	jor g10789(.dina(w_n11062_0[2]),.dinb(w_n590_19[2]),.dout(n11063),.clk(gclk));
	jand g10790(.dina(w_n11062_0[1]),.dinb(w_n590_19[1]),.dout(n11064),.clk(gclk));
	jnot g10791(.din(w_n10588_0[0]),.dout(n11065),.clk(gclk));
	jand g10792(.dina(w_asqrt19_13[2]),.dinb(n11065),.dout(n11066),.clk(gclk));
	jand g10793(.dina(w_n11066_0[1]),.dinb(w_n10593_0[0]),.dout(n11067),.clk(gclk));
	jor g10794(.dina(n11067),.dinb(w_n10592_0[0]),.dout(n11068),.clk(gclk));
	jand g10795(.dina(w_n11066_0[0]),.dinb(w_n10594_0[0]),.dout(n11069),.clk(gclk));
	jnot g10796(.din(n11069),.dout(n11070),.clk(gclk));
	jand g10797(.dina(n11070),.dinb(n11068),.dout(n11071),.clk(gclk));
	jnot g10798(.din(n11071),.dout(n11072),.clk(gclk));
	jor g10799(.dina(w_n11072_0[1]),.dinb(n11064),.dout(n11073),.clk(gclk));
	jand g10800(.dina(w_n11073_0[1]),.dinb(w_n11063_0[1]),.dout(n11074),.clk(gclk));
	jor g10801(.dina(n11074),.dinb(w_n430_21[0]),.dout(n11075),.clk(gclk));
	jand g10802(.dina(w_n11063_0[0]),.dinb(w_n430_20[2]),.dout(n11076),.clk(gclk));
	jand g10803(.dina(n11076),.dinb(w_n11073_0[0]),.dout(n11077),.clk(gclk));
	jnot g10804(.din(w_n10596_0[0]),.dout(n11078),.clk(gclk));
	jand g10805(.dina(w_asqrt19_13[1]),.dinb(n11078),.dout(n11079),.clk(gclk));
	jand g10806(.dina(w_n11079_0[1]),.dinb(w_n10603_0[0]),.dout(n11080),.clk(gclk));
	jor g10807(.dina(n11080),.dinb(w_n10601_0[0]),.dout(n11081),.clk(gclk));
	jand g10808(.dina(w_n11079_0[0]),.dinb(w_n10604_0[0]),.dout(n11082),.clk(gclk));
	jnot g10809(.din(n11082),.dout(n11083),.clk(gclk));
	jand g10810(.dina(n11083),.dinb(n11081),.dout(n11084),.clk(gclk));
	jnot g10811(.din(n11084),.dout(n11085),.clk(gclk));
	jor g10812(.dina(w_n11085_0[1]),.dinb(w_n11077_0[1]),.dout(n11086),.clk(gclk));
	jand g10813(.dina(n11086),.dinb(w_n11075_0[1]),.dout(n11087),.clk(gclk));
	jor g10814(.dina(w_n11087_0[1]),.dinb(w_n425_19[2]),.dout(n11088),.clk(gclk));
	jxor g10815(.dina(w_n10605_0[0]),.dinb(w_n430_20[1]),.dout(n11089),.clk(gclk));
	jor g10816(.dina(n11089),.dinb(w_n10701_17[2]),.dout(n11090),.clk(gclk));
	jxor g10817(.dina(n11090),.dinb(w_n10616_0[0]),.dout(n11091),.clk(gclk));
	jand g10818(.dina(w_n11087_0[0]),.dinb(w_n425_19[1]),.dout(n11092),.clk(gclk));
	jor g10819(.dina(w_n11092_0[1]),.dinb(w_n11091_0[1]),.dout(n11093),.clk(gclk));
	jand g10820(.dina(w_n11093_0[2]),.dinb(w_n11088_0[2]),.dout(n11094),.clk(gclk));
	jor g10821(.dina(n11094),.dinb(w_n305_21[1]),.dout(n11095),.clk(gclk));
	jnot g10822(.din(w_n10621_0[0]),.dout(n11096),.clk(gclk));
	jor g10823(.dina(n11096),.dinb(w_n10619_0[0]),.dout(n11097),.clk(gclk));
	jor g10824(.dina(n11097),.dinb(w_n10701_17[1]),.dout(n11098),.clk(gclk));
	jxor g10825(.dina(n11098),.dinb(w_n10630_0[0]),.dout(n11099),.clk(gclk));
	jand g10826(.dina(w_n11088_0[1]),.dinb(w_n305_21[0]),.dout(n11100),.clk(gclk));
	jand g10827(.dina(n11100),.dinb(w_n11093_0[1]),.dout(n11101),.clk(gclk));
	jor g10828(.dina(w_n11101_0[1]),.dinb(w_n11099_0[1]),.dout(n11102),.clk(gclk));
	jand g10829(.dina(w_n11102_0[1]),.dinb(w_n11095_0[1]),.dout(n11103),.clk(gclk));
	jor g10830(.dina(w_n11103_0[2]),.dinb(w_n290_21[0]),.dout(n11104),.clk(gclk));
	jand g10831(.dina(w_n11103_0[1]),.dinb(w_n290_20[2]),.dout(n11105),.clk(gclk));
	jnot g10832(.din(w_n10633_0[0]),.dout(n11106),.clk(gclk));
	jand g10833(.dina(w_asqrt19_13[0]),.dinb(n11106),.dout(n11107),.clk(gclk));
	jand g10834(.dina(w_n11107_0[1]),.dinb(w_n10638_0[0]),.dout(n11108),.clk(gclk));
	jor g10835(.dina(n11108),.dinb(w_n10637_0[0]),.dout(n11109),.clk(gclk));
	jand g10836(.dina(w_n11107_0[0]),.dinb(w_n10639_0[0]),.dout(n11110),.clk(gclk));
	jnot g10837(.din(n11110),.dout(n11111),.clk(gclk));
	jand g10838(.dina(n11111),.dinb(n11109),.dout(n11112),.clk(gclk));
	jnot g10839(.din(n11112),.dout(n11113),.clk(gclk));
	jor g10840(.dina(w_n11113_0[1]),.dinb(n11105),.dout(n11114),.clk(gclk));
	jand g10841(.dina(w_n11114_0[1]),.dinb(w_n11104_0[1]),.dout(n11115),.clk(gclk));
	jor g10842(.dina(n11115),.dinb(w_n223_21[1]),.dout(n11116),.clk(gclk));
	jand g10843(.dina(w_n11104_0[0]),.dinb(w_n223_21[0]),.dout(n11117),.clk(gclk));
	jand g10844(.dina(n11117),.dinb(w_n11114_0[0]),.dout(n11118),.clk(gclk));
	jnot g10845(.din(w_n10641_0[0]),.dout(n11119),.clk(gclk));
	jand g10846(.dina(w_asqrt19_12[2]),.dinb(n11119),.dout(n11120),.clk(gclk));
	jand g10847(.dina(w_n11120_0[1]),.dinb(w_n10648_0[0]),.dout(n11121),.clk(gclk));
	jor g10848(.dina(n11121),.dinb(w_n10646_0[0]),.dout(n11122),.clk(gclk));
	jand g10849(.dina(w_n11120_0[0]),.dinb(w_n10649_0[0]),.dout(n11123),.clk(gclk));
	jnot g10850(.din(n11123),.dout(n11124),.clk(gclk));
	jand g10851(.dina(n11124),.dinb(n11122),.dout(n11125),.clk(gclk));
	jnot g10852(.din(n11125),.dout(n11126),.clk(gclk));
	jor g10853(.dina(w_n11126_0[1]),.dinb(w_n11118_0[1]),.dout(n11127),.clk(gclk));
	jand g10854(.dina(n11127),.dinb(w_n11116_0[1]),.dout(n11128),.clk(gclk));
	jor g10855(.dina(w_n11128_0[2]),.dinb(w_n199_24[1]),.dout(n11129),.clk(gclk));
	jand g10856(.dina(w_n11128_0[1]),.dinb(w_n199_24[0]),.dout(n11130),.clk(gclk));
	jxor g10857(.dina(w_n10650_0[0]),.dinb(w_n223_20[2]),.dout(n11131),.clk(gclk));
	jor g10858(.dina(n11131),.dinb(w_n10701_17[0]),.dout(n11132),.clk(gclk));
	jxor g10859(.dina(n11132),.dinb(w_n10661_0[0]),.dout(n11133),.clk(gclk));
	jor g10860(.dina(w_n11133_0[1]),.dinb(n11130),.dout(n11134),.clk(gclk));
	jand g10861(.dina(n11134),.dinb(n11129),.dout(n11135),.clk(gclk));
	jnot g10862(.din(w_n10666_0[0]),.dout(n11136),.clk(gclk));
	jor g10863(.dina(n11136),.dinb(w_n10664_0[0]),.dout(n11137),.clk(gclk));
	jor g10864(.dina(n11137),.dinb(w_n10701_16[2]),.dout(n11138),.clk(gclk));
	jxor g10865(.dina(n11138),.dinb(w_n10675_0[0]),.dout(n11139),.clk(gclk));
	jand g10866(.dina(w_asqrt19_12[1]),.dinb(w_n10689_0[1]),.dout(n11140),.clk(gclk));
	jand g10867(.dina(w_n11140_0[1]),.dinb(w_n10677_1[0]),.dout(n11141),.clk(gclk));
	jor g10868(.dina(n11141),.dinb(w_n10723_0[0]),.dout(n11142),.clk(gclk));
	jor g10869(.dina(n11142),.dinb(w_n11139_0[2]),.dout(n11143),.clk(gclk));
	jor g10870(.dina(n11143),.dinb(w_n11135_0[2]),.dout(n11144),.clk(gclk));
	jand g10871(.dina(n11144),.dinb(w_n194_23[1]),.dout(n11145),.clk(gclk));
	jand g10872(.dina(w_n11139_0[1]),.dinb(w_n11135_0[1]),.dout(n11146),.clk(gclk));
	jor g10873(.dina(w_n11140_0[0]),.dinb(w_n10677_0[2]),.dout(n11147),.clk(gclk));
	jand g10874(.dina(w_n10689_0[0]),.dinb(w_n10677_0[1]),.dout(n11148),.clk(gclk));
	jor g10875(.dina(n11148),.dinb(w_n194_23[0]),.dout(n11149),.clk(gclk));
	jnot g10876(.din(n11149),.dout(n11150),.clk(gclk));
	jand g10877(.dina(n11150),.dinb(n11147),.dout(n11151),.clk(gclk));
	jor g10878(.dina(w_n11151_0[1]),.dinb(w_n11146_0[2]),.dout(n11154),.clk(gclk));
	jor g10879(.dina(n11154),.dinb(w_n11145_0[1]),.dout(asqrt_fa_19),.clk(gclk));
	jxor g10880(.dina(w_n10951_0[0]),.dinb(w_n2420_16[2]),.dout(n11156),.clk(gclk));
	jand g10881(.dina(n11156),.dinb(w_asqrt18_31),.dout(n11157),.clk(gclk));
	jxor g10882(.dina(n11157),.dinb(w_n10704_0[0]),.dout(n11158),.clk(gclk));
	jand g10883(.dina(w_asqrt18_30[2]),.dinb(w_a36_0[0]),.dout(n11159),.clk(gclk));
	jnot g10884(.din(w_a34_0[1]),.dout(n11160),.clk(gclk));
	jnot g10885(.din(w_a35_0[1]),.dout(n11161),.clk(gclk));
	jand g10886(.dina(w_n10706_1[0]),.dinb(w_n11161_0[1]),.dout(n11162),.clk(gclk));
	jand g10887(.dina(n11162),.dinb(w_n11160_1[1]),.dout(n11163),.clk(gclk));
	jor g10888(.dina(n11163),.dinb(n11159),.dout(n11164),.clk(gclk));
	jand g10889(.dina(w_n11164_0[2]),.dinb(w_asqrt19_12[0]),.dout(n11165),.clk(gclk));
	jand g10890(.dina(w_asqrt18_30[1]),.dinb(w_n10706_0[2]),.dout(n11166),.clk(gclk));
	jxor g10891(.dina(w_n11166_0[1]),.dinb(w_n10707_0[1]),.dout(n11167),.clk(gclk));
	jor g10892(.dina(w_n11164_0[1]),.dinb(w_asqrt19_11[2]),.dout(n11168),.clk(gclk));
	jand g10893(.dina(n11168),.dinb(w_n11167_0[1]),.dout(n11169),.clk(gclk));
	jor g10894(.dina(w_n11169_0[1]),.dinb(w_n11165_0[1]),.dout(n11170),.clk(gclk));
	jand g10895(.dina(n11170),.dinb(w_asqrt20_16[0]),.dout(n11171),.clk(gclk));
	jor g10896(.dina(w_n11165_0[0]),.dinb(w_asqrt20_15[2]),.dout(n11172),.clk(gclk));
	jor g10897(.dina(n11172),.dinb(w_n11169_0[0]),.dout(n11173),.clk(gclk));
	jand g10898(.dina(w_n11166_0[0]),.dinb(w_n10707_0[0]),.dout(n11174),.clk(gclk));
	jnot g10899(.din(w_n11145_0[0]),.dout(n11175),.clk(gclk));
	jnot g10900(.din(w_n11146_0[1]),.dout(n11176),.clk(gclk));
	jnot g10901(.din(w_n11151_0[0]),.dout(n11177),.clk(gclk));
	jand g10902(.dina(n11177),.dinb(w_asqrt19_11[1]),.dout(n11178),.clk(gclk));
	jand g10903(.dina(n11178),.dinb(n11176),.dout(n11179),.clk(gclk));
	jand g10904(.dina(n11179),.dinb(n11175),.dout(n11180),.clk(gclk));
	jor g10905(.dina(n11180),.dinb(n11174),.dout(n11181),.clk(gclk));
	jxor g10906(.dina(n11181),.dinb(w_n10219_0[1]),.dout(n11182),.clk(gclk));
	jand g10907(.dina(w_n11182_0[1]),.dinb(w_n11173_0[1]),.dout(n11183),.clk(gclk));
	jor g10908(.dina(n11183),.dinb(w_n11171_0[1]),.dout(n11184),.clk(gclk));
	jand g10909(.dina(w_n11184_0[2]),.dinb(w_asqrt21_12[0]),.dout(n11185),.clk(gclk));
	jor g10910(.dina(w_n11184_0[1]),.dinb(w_asqrt21_11[2]),.dout(n11186),.clk(gclk));
	jxor g10911(.dina(w_n10711_0[0]),.dinb(w_n10696_12[1]),.dout(n11187),.clk(gclk));
	jand g10912(.dina(n11187),.dinb(w_asqrt18_30[0]),.dout(n11188),.clk(gclk));
	jxor g10913(.dina(n11188),.dinb(w_n10714_0[0]),.dout(n11189),.clk(gclk));
	jnot g10914(.din(w_n11189_0[1]),.dout(n11190),.clk(gclk));
	jand g10915(.dina(n11190),.dinb(n11186),.dout(n11191),.clk(gclk));
	jor g10916(.dina(w_n11191_0[1]),.dinb(w_n11185_0[1]),.dout(n11192),.clk(gclk));
	jand g10917(.dina(n11192),.dinb(w_asqrt22_16[0]),.dout(n11193),.clk(gclk));
	jnot g10918(.din(w_n10720_0[0]),.dout(n11194),.clk(gclk));
	jand g10919(.dina(n11194),.dinb(w_n10718_0[0]),.dout(n11195),.clk(gclk));
	jand g10920(.dina(n11195),.dinb(w_asqrt18_29[2]),.dout(n11196),.clk(gclk));
	jxor g10921(.dina(n11196),.dinb(w_n10728_0[0]),.dout(n11197),.clk(gclk));
	jnot g10922(.din(n11197),.dout(n11198),.clk(gclk));
	jor g10923(.dina(w_n11185_0[0]),.dinb(w_asqrt22_15[2]),.dout(n11199),.clk(gclk));
	jor g10924(.dina(n11199),.dinb(w_n11191_0[0]),.dout(n11200),.clk(gclk));
	jand g10925(.dina(w_n11200_0[1]),.dinb(w_n11198_0[1]),.dout(n11201),.clk(gclk));
	jor g10926(.dina(w_n11201_0[1]),.dinb(w_n11193_0[1]),.dout(n11202),.clk(gclk));
	jand g10927(.dina(w_n11202_0[2]),.dinb(w_asqrt23_12[0]),.dout(n11203),.clk(gclk));
	jor g10928(.dina(w_n11202_0[1]),.dinb(w_asqrt23_11[2]),.dout(n11204),.clk(gclk));
	jnot g10929(.din(w_n10735_0[0]),.dout(n11205),.clk(gclk));
	jxor g10930(.dina(w_n10730_0[0]),.dinb(w_n9769_12[1]),.dout(n11206),.clk(gclk));
	jand g10931(.dina(n11206),.dinb(w_asqrt18_29[1]),.dout(n11207),.clk(gclk));
	jxor g10932(.dina(n11207),.dinb(n11205),.dout(n11208),.clk(gclk));
	jand g10933(.dina(w_n11208_0[1]),.dinb(n11204),.dout(n11209),.clk(gclk));
	jor g10934(.dina(w_n11209_0[1]),.dinb(w_n11203_0[1]),.dout(n11210),.clk(gclk));
	jand g10935(.dina(n11210),.dinb(w_asqrt24_16[0]),.dout(n11211),.clk(gclk));
	jor g10936(.dina(w_n11203_0[0]),.dinb(w_asqrt24_15[2]),.dout(n11212),.clk(gclk));
	jor g10937(.dina(n11212),.dinb(w_n11209_0[0]),.dout(n11213),.clk(gclk));
	jnot g10938(.din(w_n10742_0[0]),.dout(n11214),.clk(gclk));
	jnot g10939(.din(w_n10744_0[0]),.dout(n11215),.clk(gclk));
	jand g10940(.dina(w_asqrt18_29[0]),.dinb(w_n10738_0[0]),.dout(n11216),.clk(gclk));
	jand g10941(.dina(w_n11216_0[1]),.dinb(n11215),.dout(n11217),.clk(gclk));
	jor g10942(.dina(n11217),.dinb(n11214),.dout(n11218),.clk(gclk));
	jnot g10943(.din(w_n10745_0[0]),.dout(n11219),.clk(gclk));
	jand g10944(.dina(w_n11216_0[0]),.dinb(n11219),.dout(n11220),.clk(gclk));
	jnot g10945(.din(n11220),.dout(n11221),.clk(gclk));
	jand g10946(.dina(n11221),.dinb(n11218),.dout(n11222),.clk(gclk));
	jand g10947(.dina(w_n11222_0[1]),.dinb(w_n11213_0[1]),.dout(n11223),.clk(gclk));
	jor g10948(.dina(n11223),.dinb(w_n11211_0[1]),.dout(n11224),.clk(gclk));
	jand g10949(.dina(w_n11224_0[2]),.dinb(w_asqrt25_12[1]),.dout(n11225),.clk(gclk));
	jor g10950(.dina(w_n11224_0[1]),.dinb(w_asqrt25_12[0]),.dout(n11226),.clk(gclk));
	jxor g10951(.dina(w_n10746_0[0]),.dinb(w_n8893_12[2]),.dout(n11227),.clk(gclk));
	jand g10952(.dina(n11227),.dinb(w_asqrt18_28[2]),.dout(n11228),.clk(gclk));
	jxor g10953(.dina(n11228),.dinb(w_n10751_0[0]),.dout(n11229),.clk(gclk));
	jand g10954(.dina(w_n11229_0[1]),.dinb(n11226),.dout(n11230),.clk(gclk));
	jor g10955(.dina(w_n11230_0[1]),.dinb(w_n11225_0[1]),.dout(n11231),.clk(gclk));
	jand g10956(.dina(n11231),.dinb(w_asqrt26_16[0]),.dout(n11232),.clk(gclk));
	jnot g10957(.din(w_n10757_0[0]),.dout(n11233),.clk(gclk));
	jand g10958(.dina(n11233),.dinb(w_n10755_0[0]),.dout(n11234),.clk(gclk));
	jand g10959(.dina(n11234),.dinb(w_asqrt18_28[1]),.dout(n11235),.clk(gclk));
	jxor g10960(.dina(n11235),.dinb(w_n10766_0[0]),.dout(n11236),.clk(gclk));
	jnot g10961(.din(n11236),.dout(n11237),.clk(gclk));
	jor g10962(.dina(w_n11225_0[0]),.dinb(w_asqrt26_15[2]),.dout(n11238),.clk(gclk));
	jor g10963(.dina(n11238),.dinb(w_n11230_0[0]),.dout(n11239),.clk(gclk));
	jand g10964(.dina(w_n11239_0[1]),.dinb(w_n11237_0[1]),.dout(n11240),.clk(gclk));
	jor g10965(.dina(w_n11240_0[1]),.dinb(w_n11232_0[1]),.dout(n11241),.clk(gclk));
	jand g10966(.dina(w_n11241_0[2]),.dinb(w_asqrt27_12[1]),.dout(n11242),.clk(gclk));
	jor g10967(.dina(w_n11241_0[1]),.dinb(w_asqrt27_12[0]),.dout(n11243),.clk(gclk));
	jxor g10968(.dina(w_n10768_0[0]),.dinb(w_n8053_12[2]),.dout(n11244),.clk(gclk));
	jand g10969(.dina(n11244),.dinb(w_asqrt18_28[0]),.dout(n11245),.clk(gclk));
	jxor g10970(.dina(n11245),.dinb(w_n10774_0[0]),.dout(n11246),.clk(gclk));
	jand g10971(.dina(w_n11246_0[1]),.dinb(n11243),.dout(n11247),.clk(gclk));
	jor g10972(.dina(w_n11247_0[1]),.dinb(w_n11242_0[1]),.dout(n11248),.clk(gclk));
	jand g10973(.dina(n11248),.dinb(w_asqrt28_16[0]),.dout(n11249),.clk(gclk));
	jor g10974(.dina(w_n11242_0[0]),.dinb(w_asqrt28_15[2]),.dout(n11250),.clk(gclk));
	jor g10975(.dina(n11250),.dinb(w_n11247_0[0]),.dout(n11251),.clk(gclk));
	jnot g10976(.din(w_n10782_0[0]),.dout(n11252),.clk(gclk));
	jnot g10977(.din(w_n10784_0[0]),.dout(n11253),.clk(gclk));
	jand g10978(.dina(w_asqrt18_27[2]),.dinb(w_n10778_0[0]),.dout(n11254),.clk(gclk));
	jand g10979(.dina(w_n11254_0[1]),.dinb(n11253),.dout(n11255),.clk(gclk));
	jor g10980(.dina(n11255),.dinb(n11252),.dout(n11256),.clk(gclk));
	jnot g10981(.din(w_n10785_0[0]),.dout(n11257),.clk(gclk));
	jand g10982(.dina(w_n11254_0[0]),.dinb(n11257),.dout(n11258),.clk(gclk));
	jnot g10983(.din(n11258),.dout(n11259),.clk(gclk));
	jand g10984(.dina(n11259),.dinb(n11256),.dout(n11260),.clk(gclk));
	jand g10985(.dina(w_n11260_0[1]),.dinb(w_n11251_0[1]),.dout(n11261),.clk(gclk));
	jor g10986(.dina(n11261),.dinb(w_n11249_0[1]),.dout(n11262),.clk(gclk));
	jand g10987(.dina(w_n11262_0[1]),.dinb(w_asqrt29_12[2]),.dout(n11263),.clk(gclk));
	jxor g10988(.dina(w_n10786_0[0]),.dinb(w_n7260_13[1]),.dout(n11264),.clk(gclk));
	jand g10989(.dina(n11264),.dinb(w_asqrt18_27[1]),.dout(n11265),.clk(gclk));
	jxor g10990(.dina(n11265),.dinb(w_n10793_0[0]),.dout(n11266),.clk(gclk));
	jnot g10991(.din(n11266),.dout(n11267),.clk(gclk));
	jor g10992(.dina(w_n11262_0[0]),.dinb(w_asqrt29_12[1]),.dout(n11268),.clk(gclk));
	jand g10993(.dina(w_n11268_0[1]),.dinb(w_n11267_0[1]),.dout(n11269),.clk(gclk));
	jor g10994(.dina(w_n11269_0[2]),.dinb(w_n11263_0[2]),.dout(n11270),.clk(gclk));
	jand g10995(.dina(n11270),.dinb(w_asqrt30_16[0]),.dout(n11271),.clk(gclk));
	jnot g10996(.din(w_n10798_0[0]),.dout(n11272),.clk(gclk));
	jand g10997(.dina(n11272),.dinb(w_n10796_0[0]),.dout(n11273),.clk(gclk));
	jand g10998(.dina(n11273),.dinb(w_asqrt18_27[0]),.dout(n11274),.clk(gclk));
	jxor g10999(.dina(n11274),.dinb(w_n10806_0[0]),.dout(n11275),.clk(gclk));
	jnot g11000(.din(n11275),.dout(n11276),.clk(gclk));
	jor g11001(.dina(w_n11263_0[1]),.dinb(w_asqrt30_15[2]),.dout(n11277),.clk(gclk));
	jor g11002(.dina(n11277),.dinb(w_n11269_0[1]),.dout(n11278),.clk(gclk));
	jand g11003(.dina(w_n11278_0[1]),.dinb(w_n11276_0[1]),.dout(n11279),.clk(gclk));
	jor g11004(.dina(w_n11279_0[1]),.dinb(w_n11271_0[1]),.dout(n11280),.clk(gclk));
	jand g11005(.dina(w_n11280_0[2]),.dinb(w_asqrt31_12[2]),.dout(n11281),.clk(gclk));
	jor g11006(.dina(w_n11280_0[1]),.dinb(w_asqrt31_12[1]),.dout(n11282),.clk(gclk));
	jnot g11007(.din(w_n10812_0[0]),.dout(n11283),.clk(gclk));
	jnot g11008(.din(w_n10813_0[0]),.dout(n11284),.clk(gclk));
	jand g11009(.dina(w_asqrt18_26[2]),.dinb(w_n10809_0[0]),.dout(n11285),.clk(gclk));
	jand g11010(.dina(w_n11285_0[1]),.dinb(n11284),.dout(n11286),.clk(gclk));
	jor g11011(.dina(n11286),.dinb(n11283),.dout(n11287),.clk(gclk));
	jnot g11012(.din(w_n10814_0[0]),.dout(n11288),.clk(gclk));
	jand g11013(.dina(w_n11285_0[0]),.dinb(n11288),.dout(n11289),.clk(gclk));
	jnot g11014(.din(n11289),.dout(n11290),.clk(gclk));
	jand g11015(.dina(n11290),.dinb(n11287),.dout(n11291),.clk(gclk));
	jand g11016(.dina(w_n11291_0[1]),.dinb(n11282),.dout(n11292),.clk(gclk));
	jor g11017(.dina(w_n11292_0[1]),.dinb(w_n11281_0[1]),.dout(n11293),.clk(gclk));
	jand g11018(.dina(n11293),.dinb(w_asqrt32_16[0]),.dout(n11294),.clk(gclk));
	jor g11019(.dina(w_n11281_0[0]),.dinb(w_asqrt32_15[2]),.dout(n11295),.clk(gclk));
	jor g11020(.dina(n11295),.dinb(w_n11292_0[0]),.dout(n11296),.clk(gclk));
	jnot g11021(.din(w_n10820_0[0]),.dout(n11297),.clk(gclk));
	jnot g11022(.din(w_n10822_0[0]),.dout(n11298),.clk(gclk));
	jand g11023(.dina(w_asqrt18_26[1]),.dinb(w_n10816_0[0]),.dout(n11299),.clk(gclk));
	jand g11024(.dina(w_n11299_0[1]),.dinb(n11298),.dout(n11300),.clk(gclk));
	jor g11025(.dina(n11300),.dinb(n11297),.dout(n11301),.clk(gclk));
	jnot g11026(.din(w_n10823_0[0]),.dout(n11302),.clk(gclk));
	jand g11027(.dina(w_n11299_0[0]),.dinb(n11302),.dout(n11303),.clk(gclk));
	jnot g11028(.din(n11303),.dout(n11304),.clk(gclk));
	jand g11029(.dina(n11304),.dinb(n11301),.dout(n11305),.clk(gclk));
	jand g11030(.dina(w_n11305_0[1]),.dinb(w_n11296_0[1]),.dout(n11306),.clk(gclk));
	jor g11031(.dina(n11306),.dinb(w_n11294_0[1]),.dout(n11307),.clk(gclk));
	jand g11032(.dina(w_n11307_0[1]),.dinb(w_asqrt33_13[0]),.dout(n11308),.clk(gclk));
	jxor g11033(.dina(w_n10824_0[0]),.dinb(w_n5788_14[0]),.dout(n11309),.clk(gclk));
	jand g11034(.dina(n11309),.dinb(w_asqrt18_26[0]),.dout(n11310),.clk(gclk));
	jxor g11035(.dina(n11310),.dinb(w_n10834_0[0]),.dout(n11311),.clk(gclk));
	jnot g11036(.din(n11311),.dout(n11312),.clk(gclk));
	jor g11037(.dina(w_n11307_0[0]),.dinb(w_asqrt33_12[2]),.dout(n11313),.clk(gclk));
	jand g11038(.dina(w_n11313_0[1]),.dinb(w_n11312_0[1]),.dout(n11314),.clk(gclk));
	jor g11039(.dina(w_n11314_0[2]),.dinb(w_n11308_0[2]),.dout(n11315),.clk(gclk));
	jand g11040(.dina(n11315),.dinb(w_asqrt34_16[0]),.dout(n11316),.clk(gclk));
	jnot g11041(.din(w_n10839_0[0]),.dout(n11317),.clk(gclk));
	jand g11042(.dina(n11317),.dinb(w_n10837_0[0]),.dout(n11318),.clk(gclk));
	jand g11043(.dina(n11318),.dinb(w_asqrt18_25[2]),.dout(n11319),.clk(gclk));
	jxor g11044(.dina(n11319),.dinb(w_n10847_0[0]),.dout(n11320),.clk(gclk));
	jnot g11045(.din(n11320),.dout(n11321),.clk(gclk));
	jor g11046(.dina(w_n11308_0[1]),.dinb(w_asqrt34_15[2]),.dout(n11322),.clk(gclk));
	jor g11047(.dina(n11322),.dinb(w_n11314_0[1]),.dout(n11323),.clk(gclk));
	jand g11048(.dina(w_n11323_0[1]),.dinb(w_n11321_0[1]),.dout(n11324),.clk(gclk));
	jor g11049(.dina(w_n11324_0[1]),.dinb(w_n11316_0[1]),.dout(n11325),.clk(gclk));
	jand g11050(.dina(w_n11325_0[2]),.dinb(w_asqrt35_13[0]),.dout(n11326),.clk(gclk));
	jor g11051(.dina(w_n11325_0[1]),.dinb(w_asqrt35_12[2]),.dout(n11327),.clk(gclk));
	jnot g11052(.din(w_n10853_0[0]),.dout(n11328),.clk(gclk));
	jnot g11053(.din(w_n10854_0[0]),.dout(n11329),.clk(gclk));
	jand g11054(.dina(w_asqrt18_25[1]),.dinb(w_n10850_0[0]),.dout(n11330),.clk(gclk));
	jand g11055(.dina(w_n11330_0[1]),.dinb(n11329),.dout(n11331),.clk(gclk));
	jor g11056(.dina(n11331),.dinb(n11328),.dout(n11332),.clk(gclk));
	jnot g11057(.din(w_n10855_0[0]),.dout(n11333),.clk(gclk));
	jand g11058(.dina(w_n11330_0[0]),.dinb(n11333),.dout(n11334),.clk(gclk));
	jnot g11059(.din(n11334),.dout(n11335),.clk(gclk));
	jand g11060(.dina(n11335),.dinb(n11332),.dout(n11336),.clk(gclk));
	jand g11061(.dina(w_n11336_0[1]),.dinb(n11327),.dout(n11337),.clk(gclk));
	jor g11062(.dina(w_n11337_0[1]),.dinb(w_n11326_0[1]),.dout(n11338),.clk(gclk));
	jand g11063(.dina(n11338),.dinb(w_asqrt36_16[0]),.dout(n11339),.clk(gclk));
	jor g11064(.dina(w_n11326_0[0]),.dinb(w_asqrt36_15[2]),.dout(n11340),.clk(gclk));
	jor g11065(.dina(n11340),.dinb(w_n11337_0[0]),.dout(n11341),.clk(gclk));
	jnot g11066(.din(w_n10861_0[0]),.dout(n11342),.clk(gclk));
	jnot g11067(.din(w_n10863_0[0]),.dout(n11343),.clk(gclk));
	jand g11068(.dina(w_asqrt18_25[0]),.dinb(w_n10857_0[0]),.dout(n11344),.clk(gclk));
	jand g11069(.dina(w_n11344_0[1]),.dinb(n11343),.dout(n11345),.clk(gclk));
	jor g11070(.dina(n11345),.dinb(n11342),.dout(n11346),.clk(gclk));
	jnot g11071(.din(w_n10864_0[0]),.dout(n11347),.clk(gclk));
	jand g11072(.dina(w_n11344_0[0]),.dinb(n11347),.dout(n11348),.clk(gclk));
	jnot g11073(.din(n11348),.dout(n11349),.clk(gclk));
	jand g11074(.dina(n11349),.dinb(n11346),.dout(n11350),.clk(gclk));
	jand g11075(.dina(w_n11350_0[1]),.dinb(w_n11341_0[1]),.dout(n11351),.clk(gclk));
	jor g11076(.dina(n11351),.dinb(w_n11339_0[1]),.dout(n11352),.clk(gclk));
	jand g11077(.dina(w_n11352_0[1]),.dinb(w_asqrt37_13[1]),.dout(n11353),.clk(gclk));
	jxor g11078(.dina(w_n10865_0[0]),.dinb(w_n4494_15[0]),.dout(n11354),.clk(gclk));
	jand g11079(.dina(n11354),.dinb(w_asqrt18_24[2]),.dout(n11355),.clk(gclk));
	jxor g11080(.dina(n11355),.dinb(w_n10875_0[0]),.dout(n11356),.clk(gclk));
	jnot g11081(.din(n11356),.dout(n11357),.clk(gclk));
	jor g11082(.dina(w_n11352_0[0]),.dinb(w_asqrt37_13[0]),.dout(n11358),.clk(gclk));
	jand g11083(.dina(w_n11358_0[1]),.dinb(w_n11357_0[1]),.dout(n11359),.clk(gclk));
	jor g11084(.dina(w_n11359_0[2]),.dinb(w_n11353_0[2]),.dout(n11360),.clk(gclk));
	jand g11085(.dina(n11360),.dinb(w_asqrt38_16[0]),.dout(n11361),.clk(gclk));
	jnot g11086(.din(w_n10880_0[0]),.dout(n11362),.clk(gclk));
	jand g11087(.dina(n11362),.dinb(w_n10878_0[0]),.dout(n11363),.clk(gclk));
	jand g11088(.dina(n11363),.dinb(w_asqrt18_24[1]),.dout(n11364),.clk(gclk));
	jxor g11089(.dina(n11364),.dinb(w_n10888_0[0]),.dout(n11365),.clk(gclk));
	jnot g11090(.din(n11365),.dout(n11366),.clk(gclk));
	jor g11091(.dina(w_n11353_0[1]),.dinb(w_asqrt38_15[2]),.dout(n11367),.clk(gclk));
	jor g11092(.dina(n11367),.dinb(w_n11359_0[1]),.dout(n11368),.clk(gclk));
	jand g11093(.dina(w_n11368_0[1]),.dinb(w_n11366_0[1]),.dout(n11369),.clk(gclk));
	jor g11094(.dina(w_n11369_0[1]),.dinb(w_n11361_0[1]),.dout(n11370),.clk(gclk));
	jand g11095(.dina(w_n11370_0[2]),.dinb(w_asqrt39_13[1]),.dout(n11371),.clk(gclk));
	jor g11096(.dina(w_n11370_0[1]),.dinb(w_asqrt39_13[0]),.dout(n11372),.clk(gclk));
	jnot g11097(.din(w_n10894_0[0]),.dout(n11373),.clk(gclk));
	jnot g11098(.din(w_n10895_0[0]),.dout(n11374),.clk(gclk));
	jand g11099(.dina(w_asqrt18_24[0]),.dinb(w_n10891_0[0]),.dout(n11375),.clk(gclk));
	jand g11100(.dina(w_n11375_0[1]),.dinb(n11374),.dout(n11376),.clk(gclk));
	jor g11101(.dina(n11376),.dinb(n11373),.dout(n11377),.clk(gclk));
	jnot g11102(.din(w_n10896_0[0]),.dout(n11378),.clk(gclk));
	jand g11103(.dina(w_n11375_0[0]),.dinb(n11378),.dout(n11379),.clk(gclk));
	jnot g11104(.din(n11379),.dout(n11380),.clk(gclk));
	jand g11105(.dina(n11380),.dinb(n11377),.dout(n11381),.clk(gclk));
	jand g11106(.dina(w_n11381_0[1]),.dinb(n11372),.dout(n11382),.clk(gclk));
	jor g11107(.dina(w_n11382_0[1]),.dinb(w_n11371_0[1]),.dout(n11383),.clk(gclk));
	jand g11108(.dina(n11383),.dinb(w_asqrt40_16[0]),.dout(n11384),.clk(gclk));
	jor g11109(.dina(w_n11371_0[0]),.dinb(w_asqrt40_15[2]),.dout(n11385),.clk(gclk));
	jor g11110(.dina(n11385),.dinb(w_n11382_0[0]),.dout(n11386),.clk(gclk));
	jnot g11111(.din(w_n10902_0[0]),.dout(n11387),.clk(gclk));
	jnot g11112(.din(w_n10904_0[0]),.dout(n11388),.clk(gclk));
	jand g11113(.dina(w_asqrt18_23[2]),.dinb(w_n10898_0[0]),.dout(n11389),.clk(gclk));
	jand g11114(.dina(w_n11389_0[1]),.dinb(n11388),.dout(n11390),.clk(gclk));
	jor g11115(.dina(n11390),.dinb(n11387),.dout(n11391),.clk(gclk));
	jnot g11116(.din(w_n10905_0[0]),.dout(n11392),.clk(gclk));
	jand g11117(.dina(w_n11389_0[0]),.dinb(n11392),.dout(n11393),.clk(gclk));
	jnot g11118(.din(n11393),.dout(n11394),.clk(gclk));
	jand g11119(.dina(n11394),.dinb(n11391),.dout(n11395),.clk(gclk));
	jand g11120(.dina(w_n11395_0[1]),.dinb(w_n11386_0[1]),.dout(n11396),.clk(gclk));
	jor g11121(.dina(n11396),.dinb(w_n11384_0[1]),.dout(n11397),.clk(gclk));
	jand g11122(.dina(w_n11397_0[1]),.dinb(w_asqrt41_13[2]),.dout(n11398),.clk(gclk));
	jxor g11123(.dina(w_n10906_0[0]),.dinb(w_n3371_15[2]),.dout(n11399),.clk(gclk));
	jand g11124(.dina(n11399),.dinb(w_asqrt18_23[1]),.dout(n11400),.clk(gclk));
	jxor g11125(.dina(n11400),.dinb(w_n10916_0[0]),.dout(n11401),.clk(gclk));
	jnot g11126(.din(n11401),.dout(n11402),.clk(gclk));
	jor g11127(.dina(w_n11397_0[0]),.dinb(w_asqrt41_13[1]),.dout(n11403),.clk(gclk));
	jand g11128(.dina(w_n11403_0[1]),.dinb(w_n11402_0[1]),.dout(n11404),.clk(gclk));
	jor g11129(.dina(w_n11404_0[2]),.dinb(w_n11398_0[2]),.dout(n11405),.clk(gclk));
	jand g11130(.dina(n11405),.dinb(w_asqrt42_16[0]),.dout(n11406),.clk(gclk));
	jnot g11131(.din(w_n10921_0[0]),.dout(n11407),.clk(gclk));
	jand g11132(.dina(n11407),.dinb(w_n10919_0[0]),.dout(n11408),.clk(gclk));
	jand g11133(.dina(n11408),.dinb(w_asqrt18_23[0]),.dout(n11409),.clk(gclk));
	jxor g11134(.dina(n11409),.dinb(w_n10929_0[0]),.dout(n11410),.clk(gclk));
	jnot g11135(.din(n11410),.dout(n11411),.clk(gclk));
	jor g11136(.dina(w_n11398_0[1]),.dinb(w_asqrt42_15[2]),.dout(n11412),.clk(gclk));
	jor g11137(.dina(n11412),.dinb(w_n11404_0[1]),.dout(n11413),.clk(gclk));
	jand g11138(.dina(w_n11413_0[1]),.dinb(w_n11411_0[1]),.dout(n11414),.clk(gclk));
	jor g11139(.dina(w_n11414_0[1]),.dinb(w_n11406_0[1]),.dout(n11415),.clk(gclk));
	jand g11140(.dina(w_n11415_0[2]),.dinb(w_asqrt43_13[2]),.dout(n11416),.clk(gclk));
	jor g11141(.dina(w_n11415_0[1]),.dinb(w_asqrt43_13[1]),.dout(n11417),.clk(gclk));
	jnot g11142(.din(w_n10935_0[0]),.dout(n11418),.clk(gclk));
	jnot g11143(.din(w_n10936_0[0]),.dout(n11419),.clk(gclk));
	jand g11144(.dina(w_asqrt18_22[2]),.dinb(w_n10932_0[0]),.dout(n11420),.clk(gclk));
	jand g11145(.dina(w_n11420_0[1]),.dinb(n11419),.dout(n11421),.clk(gclk));
	jor g11146(.dina(n11421),.dinb(n11418),.dout(n11422),.clk(gclk));
	jnot g11147(.din(w_n10937_0[0]),.dout(n11423),.clk(gclk));
	jand g11148(.dina(w_n11420_0[0]),.dinb(n11423),.dout(n11424),.clk(gclk));
	jnot g11149(.din(n11424),.dout(n11425),.clk(gclk));
	jand g11150(.dina(n11425),.dinb(n11422),.dout(n11426),.clk(gclk));
	jand g11151(.dina(w_n11426_0[1]),.dinb(n11417),.dout(n11427),.clk(gclk));
	jor g11152(.dina(w_n11427_0[1]),.dinb(w_n11416_0[1]),.dout(n11428),.clk(gclk));
	jand g11153(.dina(n11428),.dinb(w_asqrt44_16[0]),.dout(n11429),.clk(gclk));
	jnot g11154(.din(w_n10941_0[0]),.dout(n11430),.clk(gclk));
	jand g11155(.dina(n11430),.dinb(w_n10939_0[0]),.dout(n11431),.clk(gclk));
	jand g11156(.dina(n11431),.dinb(w_asqrt18_22[1]),.dout(n11432),.clk(gclk));
	jxor g11157(.dina(n11432),.dinb(w_n10949_0[0]),.dout(n11433),.clk(gclk));
	jnot g11158(.din(n11433),.dout(n11434),.clk(gclk));
	jor g11159(.dina(w_n11416_0[0]),.dinb(w_asqrt44_15[2]),.dout(n11435),.clk(gclk));
	jor g11160(.dina(n11435),.dinb(w_n11427_0[0]),.dout(n11436),.clk(gclk));
	jand g11161(.dina(w_n11436_0[1]),.dinb(w_n11434_0[1]),.dout(n11437),.clk(gclk));
	jor g11162(.dina(w_n11437_0[1]),.dinb(w_n11429_0[1]),.dout(n11438),.clk(gclk));
	jand g11163(.dina(w_n11438_0[2]),.dinb(w_asqrt45_14[0]),.dout(n11439),.clk(gclk));
	jnot g11164(.din(w_n11158_0[1]),.dout(n11440),.clk(gclk));
	jor g11165(.dina(w_n11438_0[1]),.dinb(w_asqrt45_13[2]),.dout(n11441),.clk(gclk));
	jand g11166(.dina(n11441),.dinb(n11440),.dout(n11442),.clk(gclk));
	jor g11167(.dina(w_n11442_0[1]),.dinb(w_n11439_0[1]),.dout(n11443),.clk(gclk));
	jand g11168(.dina(n11443),.dinb(w_asqrt46_16[0]),.dout(n11444),.clk(gclk));
	jor g11169(.dina(w_n11439_0[0]),.dinb(w_asqrt46_15[2]),.dout(n11445),.clk(gclk));
	jor g11170(.dina(n11445),.dinb(w_n11442_0[0]),.dout(n11446),.clk(gclk));
	jnot g11171(.din(w_n10960_0[0]),.dout(n11447),.clk(gclk));
	jnot g11172(.din(w_n10962_0[0]),.dout(n11448),.clk(gclk));
	jand g11173(.dina(w_asqrt18_22[0]),.dinb(w_n10956_0[0]),.dout(n11449),.clk(gclk));
	jand g11174(.dina(w_n11449_0[1]),.dinb(n11448),.dout(n11450),.clk(gclk));
	jor g11175(.dina(n11450),.dinb(n11447),.dout(n11451),.clk(gclk));
	jnot g11176(.din(w_n10963_0[0]),.dout(n11452),.clk(gclk));
	jand g11177(.dina(w_n11449_0[0]),.dinb(n11452),.dout(n11453),.clk(gclk));
	jnot g11178(.din(n11453),.dout(n11454),.clk(gclk));
	jand g11179(.dina(n11454),.dinb(n11451),.dout(n11455),.clk(gclk));
	jand g11180(.dina(w_n11455_0[1]),.dinb(w_n11446_0[1]),.dout(n11456),.clk(gclk));
	jor g11181(.dina(n11456),.dinb(w_n11444_0[1]),.dout(n11457),.clk(gclk));
	jand g11182(.dina(w_n11457_0[2]),.dinb(w_asqrt47_14[0]),.dout(n11458),.clk(gclk));
	jor g11183(.dina(w_n11457_0[1]),.dinb(w_asqrt47_13[2]),.dout(n11459),.clk(gclk));
	jnot g11184(.din(w_n10968_0[0]),.dout(n11460),.clk(gclk));
	jnot g11185(.din(w_n10969_0[0]),.dout(n11461),.clk(gclk));
	jand g11186(.dina(w_asqrt18_21[2]),.dinb(w_n10965_0[0]),.dout(n11462),.clk(gclk));
	jand g11187(.dina(w_n11462_0[1]),.dinb(n11461),.dout(n11463),.clk(gclk));
	jor g11188(.dina(n11463),.dinb(n11460),.dout(n11464),.clk(gclk));
	jnot g11189(.din(w_n10970_0[0]),.dout(n11465),.clk(gclk));
	jand g11190(.dina(w_n11462_0[0]),.dinb(n11465),.dout(n11466),.clk(gclk));
	jnot g11191(.din(n11466),.dout(n11467),.clk(gclk));
	jand g11192(.dina(n11467),.dinb(n11464),.dout(n11468),.clk(gclk));
	jand g11193(.dina(w_n11468_0[1]),.dinb(n11459),.dout(n11469),.clk(gclk));
	jor g11194(.dina(w_n11469_0[1]),.dinb(w_n11458_0[1]),.dout(n11470),.clk(gclk));
	jand g11195(.dina(n11470),.dinb(w_asqrt48_16[0]),.dout(n11471),.clk(gclk));
	jor g11196(.dina(w_n11458_0[0]),.dinb(w_asqrt48_15[2]),.dout(n11472),.clk(gclk));
	jor g11197(.dina(n11472),.dinb(w_n11469_0[0]),.dout(n11473),.clk(gclk));
	jnot g11198(.din(w_n10976_0[0]),.dout(n11474),.clk(gclk));
	jnot g11199(.din(w_n10978_0[0]),.dout(n11475),.clk(gclk));
	jand g11200(.dina(w_asqrt18_21[1]),.dinb(w_n10972_0[0]),.dout(n11476),.clk(gclk));
	jand g11201(.dina(w_n11476_0[1]),.dinb(n11475),.dout(n11477),.clk(gclk));
	jor g11202(.dina(n11477),.dinb(n11474),.dout(n11478),.clk(gclk));
	jnot g11203(.din(w_n10979_0[0]),.dout(n11479),.clk(gclk));
	jand g11204(.dina(w_n11476_0[0]),.dinb(n11479),.dout(n11480),.clk(gclk));
	jnot g11205(.din(n11480),.dout(n11481),.clk(gclk));
	jand g11206(.dina(n11481),.dinb(n11478),.dout(n11482),.clk(gclk));
	jand g11207(.dina(w_n11482_0[1]),.dinb(w_n11473_0[1]),.dout(n11483),.clk(gclk));
	jor g11208(.dina(n11483),.dinb(w_n11471_0[1]),.dout(n11484),.clk(gclk));
	jand g11209(.dina(w_n11484_0[1]),.dinb(w_asqrt49_14[1]),.dout(n11485),.clk(gclk));
	jxor g11210(.dina(w_n10980_0[0]),.dinb(w_n1641_17[1]),.dout(n11486),.clk(gclk));
	jand g11211(.dina(n11486),.dinb(w_asqrt18_21[0]),.dout(n11487),.clk(gclk));
	jxor g11212(.dina(n11487),.dinb(w_n10990_0[0]),.dout(n11488),.clk(gclk));
	jnot g11213(.din(n11488),.dout(n11489),.clk(gclk));
	jor g11214(.dina(w_n11484_0[0]),.dinb(w_asqrt49_14[0]),.dout(n11490),.clk(gclk));
	jand g11215(.dina(w_n11490_0[1]),.dinb(w_n11489_0[1]),.dout(n11491),.clk(gclk));
	jor g11216(.dina(w_n11491_0[2]),.dinb(w_n11485_0[2]),.dout(n11492),.clk(gclk));
	jand g11217(.dina(n11492),.dinb(w_asqrt50_16[0]),.dout(n11493),.clk(gclk));
	jnot g11218(.din(w_n10995_0[0]),.dout(n11494),.clk(gclk));
	jand g11219(.dina(n11494),.dinb(w_n10993_0[0]),.dout(n11495),.clk(gclk));
	jand g11220(.dina(n11495),.dinb(w_asqrt18_20[2]),.dout(n11496),.clk(gclk));
	jxor g11221(.dina(n11496),.dinb(w_n11003_0[0]),.dout(n11497),.clk(gclk));
	jnot g11222(.din(n11497),.dout(n11498),.clk(gclk));
	jor g11223(.dina(w_n11485_0[1]),.dinb(w_asqrt50_15[2]),.dout(n11499),.clk(gclk));
	jor g11224(.dina(n11499),.dinb(w_n11491_0[1]),.dout(n11500),.clk(gclk));
	jand g11225(.dina(w_n11500_0[1]),.dinb(w_n11498_0[1]),.dout(n11501),.clk(gclk));
	jor g11226(.dina(w_n11501_0[1]),.dinb(w_n11493_0[1]),.dout(n11502),.clk(gclk));
	jand g11227(.dina(w_n11502_0[2]),.dinb(w_asqrt51_14[1]),.dout(n11503),.clk(gclk));
	jor g11228(.dina(w_n11502_0[1]),.dinb(w_asqrt51_14[0]),.dout(n11504),.clk(gclk));
	jnot g11229(.din(w_n11009_0[0]),.dout(n11505),.clk(gclk));
	jnot g11230(.din(w_n11010_0[0]),.dout(n11506),.clk(gclk));
	jand g11231(.dina(w_asqrt18_20[1]),.dinb(w_n11006_0[0]),.dout(n11507),.clk(gclk));
	jand g11232(.dina(w_n11507_0[1]),.dinb(n11506),.dout(n11508),.clk(gclk));
	jor g11233(.dina(n11508),.dinb(n11505),.dout(n11509),.clk(gclk));
	jnot g11234(.din(w_n11011_0[0]),.dout(n11510),.clk(gclk));
	jand g11235(.dina(w_n11507_0[0]),.dinb(n11510),.dout(n11511),.clk(gclk));
	jnot g11236(.din(n11511),.dout(n11512),.clk(gclk));
	jand g11237(.dina(n11512),.dinb(n11509),.dout(n11513),.clk(gclk));
	jand g11238(.dina(w_n11513_0[1]),.dinb(n11504),.dout(n11514),.clk(gclk));
	jor g11239(.dina(w_n11514_0[1]),.dinb(w_n11503_0[1]),.dout(n11515),.clk(gclk));
	jand g11240(.dina(n11515),.dinb(w_asqrt52_16[0]),.dout(n11516),.clk(gclk));
	jor g11241(.dina(w_n11503_0[0]),.dinb(w_asqrt52_15[2]),.dout(n11517),.clk(gclk));
	jor g11242(.dina(n11517),.dinb(w_n11514_0[0]),.dout(n11518),.clk(gclk));
	jnot g11243(.din(w_n11017_0[0]),.dout(n11519),.clk(gclk));
	jnot g11244(.din(w_n11019_0[0]),.dout(n11520),.clk(gclk));
	jand g11245(.dina(w_asqrt18_20[0]),.dinb(w_n11013_0[0]),.dout(n11521),.clk(gclk));
	jand g11246(.dina(w_n11521_0[1]),.dinb(n11520),.dout(n11522),.clk(gclk));
	jor g11247(.dina(n11522),.dinb(n11519),.dout(n11523),.clk(gclk));
	jnot g11248(.din(w_n11020_0[0]),.dout(n11524),.clk(gclk));
	jand g11249(.dina(w_n11521_0[0]),.dinb(n11524),.dout(n11525),.clk(gclk));
	jnot g11250(.din(n11525),.dout(n11526),.clk(gclk));
	jand g11251(.dina(n11526),.dinb(n11523),.dout(n11527),.clk(gclk));
	jand g11252(.dina(w_n11527_0[1]),.dinb(w_n11518_0[1]),.dout(n11528),.clk(gclk));
	jor g11253(.dina(n11528),.dinb(w_n11516_0[1]),.dout(n11529),.clk(gclk));
	jand g11254(.dina(w_n11529_0[1]),.dinb(w_asqrt53_14[2]),.dout(n11530),.clk(gclk));
	jxor g11255(.dina(w_n11021_0[0]),.dinb(w_n1034_18[1]),.dout(n11531),.clk(gclk));
	jand g11256(.dina(n11531),.dinb(w_asqrt18_19[2]),.dout(n11532),.clk(gclk));
	jxor g11257(.dina(n11532),.dinb(w_n11031_0[0]),.dout(n11533),.clk(gclk));
	jnot g11258(.din(n11533),.dout(n11534),.clk(gclk));
	jor g11259(.dina(w_n11529_0[0]),.dinb(w_asqrt53_14[1]),.dout(n11535),.clk(gclk));
	jand g11260(.dina(w_n11535_0[1]),.dinb(w_n11534_0[1]),.dout(n11536),.clk(gclk));
	jor g11261(.dina(w_n11536_0[2]),.dinb(w_n11530_0[2]),.dout(n11537),.clk(gclk));
	jand g11262(.dina(n11537),.dinb(w_asqrt54_16[0]),.dout(n11538),.clk(gclk));
	jnot g11263(.din(w_n11036_0[0]),.dout(n11539),.clk(gclk));
	jand g11264(.dina(n11539),.dinb(w_n11034_0[0]),.dout(n11540),.clk(gclk));
	jand g11265(.dina(n11540),.dinb(w_asqrt18_19[1]),.dout(n11541),.clk(gclk));
	jxor g11266(.dina(n11541),.dinb(w_n11044_0[0]),.dout(n11542),.clk(gclk));
	jnot g11267(.din(n11542),.dout(n11543),.clk(gclk));
	jor g11268(.dina(w_n11530_0[1]),.dinb(w_asqrt54_15[2]),.dout(n11544),.clk(gclk));
	jor g11269(.dina(n11544),.dinb(w_n11536_0[1]),.dout(n11545),.clk(gclk));
	jand g11270(.dina(w_n11545_0[1]),.dinb(w_n11543_0[1]),.dout(n11546),.clk(gclk));
	jor g11271(.dina(w_n11546_0[1]),.dinb(w_n11538_0[1]),.dout(n11547),.clk(gclk));
	jand g11272(.dina(w_n11547_0[2]),.dinb(w_asqrt55_15[0]),.dout(n11548),.clk(gclk));
	jor g11273(.dina(w_n11547_0[1]),.dinb(w_asqrt55_14[2]),.dout(n11549),.clk(gclk));
	jnot g11274(.din(w_n11050_0[0]),.dout(n11550),.clk(gclk));
	jnot g11275(.din(w_n11051_0[0]),.dout(n11551),.clk(gclk));
	jand g11276(.dina(w_asqrt18_19[0]),.dinb(w_n11047_0[0]),.dout(n11552),.clk(gclk));
	jand g11277(.dina(w_n11552_0[1]),.dinb(n11551),.dout(n11553),.clk(gclk));
	jor g11278(.dina(n11553),.dinb(n11550),.dout(n11554),.clk(gclk));
	jnot g11279(.din(w_n11052_0[0]),.dout(n11555),.clk(gclk));
	jand g11280(.dina(w_n11552_0[0]),.dinb(n11555),.dout(n11556),.clk(gclk));
	jnot g11281(.din(n11556),.dout(n11557),.clk(gclk));
	jand g11282(.dina(n11557),.dinb(n11554),.dout(n11558),.clk(gclk));
	jand g11283(.dina(w_n11558_0[1]),.dinb(n11549),.dout(n11559),.clk(gclk));
	jor g11284(.dina(w_n11559_0[1]),.dinb(w_n11548_0[1]),.dout(n11560),.clk(gclk));
	jand g11285(.dina(n11560),.dinb(w_asqrt56_16[0]),.dout(n11561),.clk(gclk));
	jor g11286(.dina(w_n11548_0[0]),.dinb(w_asqrt56_15[2]),.dout(n11562),.clk(gclk));
	jor g11287(.dina(n11562),.dinb(w_n11559_0[0]),.dout(n11563),.clk(gclk));
	jnot g11288(.din(w_n11058_0[0]),.dout(n11564),.clk(gclk));
	jnot g11289(.din(w_n11060_0[0]),.dout(n11565),.clk(gclk));
	jand g11290(.dina(w_asqrt18_18[2]),.dinb(w_n11054_0[0]),.dout(n11566),.clk(gclk));
	jand g11291(.dina(w_n11566_0[1]),.dinb(n11565),.dout(n11567),.clk(gclk));
	jor g11292(.dina(n11567),.dinb(n11564),.dout(n11568),.clk(gclk));
	jnot g11293(.din(w_n11061_0[0]),.dout(n11569),.clk(gclk));
	jand g11294(.dina(w_n11566_0[0]),.dinb(n11569),.dout(n11570),.clk(gclk));
	jnot g11295(.din(n11570),.dout(n11571),.clk(gclk));
	jand g11296(.dina(n11571),.dinb(n11568),.dout(n11572),.clk(gclk));
	jand g11297(.dina(w_n11572_0[1]),.dinb(w_n11563_0[1]),.dout(n11573),.clk(gclk));
	jor g11298(.dina(n11573),.dinb(w_n11561_0[1]),.dout(n11574),.clk(gclk));
	jand g11299(.dina(w_n11574_0[1]),.dinb(w_asqrt57_15[1]),.dout(n11575),.clk(gclk));
	jxor g11300(.dina(w_n11062_0[0]),.dinb(w_n590_19[0]),.dout(n11576),.clk(gclk));
	jand g11301(.dina(n11576),.dinb(w_asqrt18_18[1]),.dout(n11577),.clk(gclk));
	jxor g11302(.dina(n11577),.dinb(w_n11072_0[0]),.dout(n11578),.clk(gclk));
	jnot g11303(.din(n11578),.dout(n11579),.clk(gclk));
	jor g11304(.dina(w_n11574_0[0]),.dinb(w_asqrt57_15[0]),.dout(n11580),.clk(gclk));
	jand g11305(.dina(w_n11580_0[1]),.dinb(w_n11579_0[1]),.dout(n11581),.clk(gclk));
	jor g11306(.dina(w_n11581_0[2]),.dinb(w_n11575_0[2]),.dout(n11582),.clk(gclk));
	jand g11307(.dina(n11582),.dinb(w_asqrt58_16[0]),.dout(n11583),.clk(gclk));
	jnot g11308(.din(w_n11077_0[0]),.dout(n11584),.clk(gclk));
	jand g11309(.dina(n11584),.dinb(w_n11075_0[0]),.dout(n11585),.clk(gclk));
	jand g11310(.dina(n11585),.dinb(w_asqrt18_18[0]),.dout(n11586),.clk(gclk));
	jxor g11311(.dina(n11586),.dinb(w_n11085_0[0]),.dout(n11587),.clk(gclk));
	jnot g11312(.din(n11587),.dout(n11588),.clk(gclk));
	jor g11313(.dina(w_n11575_0[1]),.dinb(w_asqrt58_15[2]),.dout(n11589),.clk(gclk));
	jor g11314(.dina(n11589),.dinb(w_n11581_0[1]),.dout(n11590),.clk(gclk));
	jand g11315(.dina(w_n11590_0[1]),.dinb(w_n11588_0[1]),.dout(n11591),.clk(gclk));
	jor g11316(.dina(w_n11591_0[1]),.dinb(w_n11583_0[1]),.dout(n11592),.clk(gclk));
	jand g11317(.dina(w_n11592_0[2]),.dinb(w_asqrt59_15[2]),.dout(n11593),.clk(gclk));
	jor g11318(.dina(w_n11592_0[1]),.dinb(w_asqrt59_15[1]),.dout(n11594),.clk(gclk));
	jnot g11319(.din(w_n11091_0[0]),.dout(n11595),.clk(gclk));
	jnot g11320(.din(w_n11092_0[0]),.dout(n11596),.clk(gclk));
	jand g11321(.dina(w_asqrt18_17[2]),.dinb(w_n11088_0[0]),.dout(n11597),.clk(gclk));
	jand g11322(.dina(w_n11597_0[1]),.dinb(n11596),.dout(n11598),.clk(gclk));
	jor g11323(.dina(n11598),.dinb(n11595),.dout(n11599),.clk(gclk));
	jnot g11324(.din(w_n11093_0[0]),.dout(n11600),.clk(gclk));
	jand g11325(.dina(w_n11597_0[0]),.dinb(n11600),.dout(n11601),.clk(gclk));
	jnot g11326(.din(n11601),.dout(n11602),.clk(gclk));
	jand g11327(.dina(n11602),.dinb(n11599),.dout(n11603),.clk(gclk));
	jand g11328(.dina(w_n11603_0[1]),.dinb(n11594),.dout(n11604),.clk(gclk));
	jor g11329(.dina(w_n11604_0[1]),.dinb(w_n11593_0[1]),.dout(n11605),.clk(gclk));
	jand g11330(.dina(n11605),.dinb(w_asqrt60_15[2]),.dout(n11606),.clk(gclk));
	jor g11331(.dina(w_n11593_0[0]),.dinb(w_asqrt60_15[1]),.dout(n11607),.clk(gclk));
	jor g11332(.dina(n11607),.dinb(w_n11604_0[0]),.dout(n11608),.clk(gclk));
	jnot g11333(.din(w_n11099_0[0]),.dout(n11609),.clk(gclk));
	jnot g11334(.din(w_n11101_0[0]),.dout(n11610),.clk(gclk));
	jand g11335(.dina(w_asqrt18_17[1]),.dinb(w_n11095_0[0]),.dout(n11611),.clk(gclk));
	jand g11336(.dina(w_n11611_0[1]),.dinb(n11610),.dout(n11612),.clk(gclk));
	jor g11337(.dina(n11612),.dinb(n11609),.dout(n11613),.clk(gclk));
	jnot g11338(.din(w_n11102_0[0]),.dout(n11614),.clk(gclk));
	jand g11339(.dina(w_n11611_0[0]),.dinb(n11614),.dout(n11615),.clk(gclk));
	jnot g11340(.din(n11615),.dout(n11616),.clk(gclk));
	jand g11341(.dina(n11616),.dinb(n11613),.dout(n11617),.clk(gclk));
	jand g11342(.dina(w_n11617_0[1]),.dinb(w_n11608_0[1]),.dout(n11618),.clk(gclk));
	jor g11343(.dina(n11618),.dinb(w_n11606_0[1]),.dout(n11619),.clk(gclk));
	jand g11344(.dina(w_n11619_0[1]),.dinb(w_asqrt61_16[0]),.dout(n11620),.clk(gclk));
	jxor g11345(.dina(w_n11103_0[0]),.dinb(w_n290_20[1]),.dout(n11621),.clk(gclk));
	jand g11346(.dina(n11621),.dinb(w_asqrt18_17[0]),.dout(n11622),.clk(gclk));
	jxor g11347(.dina(n11622),.dinb(w_n11113_0[0]),.dout(n11623),.clk(gclk));
	jnot g11348(.din(n11623),.dout(n11624),.clk(gclk));
	jor g11349(.dina(w_n11619_0[0]),.dinb(w_asqrt61_15[2]),.dout(n11625),.clk(gclk));
	jand g11350(.dina(w_n11625_0[1]),.dinb(w_n11624_0[1]),.dout(n11626),.clk(gclk));
	jor g11351(.dina(w_n11626_0[2]),.dinb(w_n11620_0[2]),.dout(n11627),.clk(gclk));
	jand g11352(.dina(n11627),.dinb(w_asqrt62_16[0]),.dout(n11628),.clk(gclk));
	jnot g11353(.din(w_n11118_0[0]),.dout(n11629),.clk(gclk));
	jand g11354(.dina(n11629),.dinb(w_n11116_0[0]),.dout(n11630),.clk(gclk));
	jand g11355(.dina(n11630),.dinb(w_asqrt18_16[2]),.dout(n11631),.clk(gclk));
	jxor g11356(.dina(n11631),.dinb(w_n11126_0[0]),.dout(n11632),.clk(gclk));
	jnot g11357(.din(n11632),.dout(n11633),.clk(gclk));
	jor g11358(.dina(w_n11620_0[1]),.dinb(w_asqrt62_15[2]),.dout(n11634),.clk(gclk));
	jor g11359(.dina(n11634),.dinb(w_n11626_0[1]),.dout(n11635),.clk(gclk));
	jand g11360(.dina(w_n11635_0[1]),.dinb(w_n11633_0[1]),.dout(n11636),.clk(gclk));
	jor g11361(.dina(w_n11636_0[1]),.dinb(w_n11628_0[1]),.dout(n11637),.clk(gclk));
	jxor g11362(.dina(w_n11128_0[0]),.dinb(w_n199_23[2]),.dout(n11638),.clk(gclk));
	jand g11363(.dina(n11638),.dinb(w_asqrt18_16[1]),.dout(n11639),.clk(gclk));
	jxor g11364(.dina(n11639),.dinb(w_n11133_0[0]),.dout(n11640),.clk(gclk));
	jnot g11365(.din(w_n11135_0[0]),.dout(n11641),.clk(gclk));
	jnot g11366(.din(w_n11139_0[0]),.dout(n11642),.clk(gclk));
	jand g11367(.dina(w_asqrt18_16[0]),.dinb(w_n11642_0[1]),.dout(n11643),.clk(gclk));
	jand g11368(.dina(w_n11643_0[1]),.dinb(w_n11641_0[2]),.dout(n11644),.clk(gclk));
	jor g11369(.dina(n11644),.dinb(w_n11146_0[0]),.dout(n11645),.clk(gclk));
	jor g11370(.dina(n11645),.dinb(w_n11640_0[1]),.dout(n11646),.clk(gclk));
	jnot g11371(.din(n11646),.dout(n11647),.clk(gclk));
	jand g11372(.dina(n11647),.dinb(w_n11637_1[2]),.dout(n11648),.clk(gclk));
	jor g11373(.dina(n11648),.dinb(w_asqrt63_8[2]),.dout(n11649),.clk(gclk));
	jnot g11374(.din(w_n11640_0[0]),.dout(n11650),.clk(gclk));
	jor g11375(.dina(w_n11650_0[2]),.dinb(w_n11637_1[1]),.dout(n11651),.clk(gclk));
	jor g11376(.dina(w_n11643_0[0]),.dinb(w_n11641_0[1]),.dout(n11652),.clk(gclk));
	jand g11377(.dina(w_n11642_0[0]),.dinb(w_n11641_0[0]),.dout(n11653),.clk(gclk));
	jor g11378(.dina(n11653),.dinb(w_n194_22[2]),.dout(n11654),.clk(gclk));
	jnot g11379(.din(n11654),.dout(n11655),.clk(gclk));
	jand g11380(.dina(n11655),.dinb(n11652),.dout(n11656),.clk(gclk));
	jnot g11381(.din(w_asqrt18_15[2]),.dout(n11657),.clk(gclk));
	jnot g11382(.din(w_n11656_0[1]),.dout(n11660),.clk(gclk));
	jand g11383(.dina(n11660),.dinb(w_n11651_0[1]),.dout(n11661),.clk(gclk));
	jand g11384(.dina(n11661),.dinb(w_n11649_0[1]),.dout(n11662),.clk(gclk));
	jxor g11385(.dina(w_n11438_0[0]),.dinb(w_n2010_18[2]),.dout(n11663),.clk(gclk));
	jor g11386(.dina(n11663),.dinb(w_n11662_24[1]),.dout(n11664),.clk(gclk));
	jxor g11387(.dina(n11664),.dinb(w_n11158_0[0]),.dout(n11665),.clk(gclk));
	jor g11388(.dina(w_n11662_24[0]),.dinb(w_n11160_1[0]),.dout(n11666),.clk(gclk));
	jnot g11389(.din(w_a32_0[1]),.dout(n11667),.clk(gclk));
	jnot g11390(.din(a[33]),.dout(n11668),.clk(gclk));
	jand g11391(.dina(w_n11160_0[2]),.dinb(w_n11668_0[2]),.dout(n11669),.clk(gclk));
	jand g11392(.dina(n11669),.dinb(w_n11667_1[1]),.dout(n11670),.clk(gclk));
	jnot g11393(.din(n11670),.dout(n11671),.clk(gclk));
	jand g11394(.dina(n11671),.dinb(n11666),.dout(n11672),.clk(gclk));
	jor g11395(.dina(w_n11672_0[2]),.dinb(w_n11657_11[2]),.dout(n11673),.clk(gclk));
	jor g11396(.dina(w_n11662_23[2]),.dinb(w_a34_0[0]),.dout(n11674),.clk(gclk));
	jxor g11397(.dina(w_n11674_0[1]),.dinb(w_n11161_0[0]),.dout(n11675),.clk(gclk));
	jand g11398(.dina(w_n11672_0[1]),.dinb(w_n11657_11[1]),.dout(n11676),.clk(gclk));
	jor g11399(.dina(n11676),.dinb(w_n11675_0[1]),.dout(n11677),.clk(gclk));
	jand g11400(.dina(w_n11677_0[1]),.dinb(w_n11673_0[1]),.dout(n11678),.clk(gclk));
	jor g11401(.dina(n11678),.dinb(w_n10701_16[1]),.dout(n11679),.clk(gclk));
	jand g11402(.dina(w_n11673_0[0]),.dinb(w_n10701_16[0]),.dout(n11680),.clk(gclk));
	jand g11403(.dina(n11680),.dinb(w_n11677_0[0]),.dout(n11681),.clk(gclk));
	jor g11404(.dina(w_n11674_0[0]),.dinb(w_a35_0[0]),.dout(n11682),.clk(gclk));
	jnot g11405(.din(w_n11649_0[0]),.dout(n11683),.clk(gclk));
	jnot g11406(.din(w_n11651_0[0]),.dout(n11684),.clk(gclk));
	jor g11407(.dina(w_n11656_0[0]),.dinb(w_n11657_11[0]),.dout(n11685),.clk(gclk));
	jor g11408(.dina(n11685),.dinb(w_n11684_0[1]),.dout(n11686),.clk(gclk));
	jor g11409(.dina(n11686),.dinb(n11683),.dout(n11687),.clk(gclk));
	jand g11410(.dina(n11687),.dinb(n11682),.dout(n11688),.clk(gclk));
	jxor g11411(.dina(n11688),.dinb(w_n10706_0[1]),.dout(n11689),.clk(gclk));
	jor g11412(.dina(w_n11689_0[1]),.dinb(w_n11681_0[1]),.dout(n11690),.clk(gclk));
	jand g11413(.dina(n11690),.dinb(w_n11679_0[1]),.dout(n11691),.clk(gclk));
	jor g11414(.dina(w_n11691_0[2]),.dinb(w_n10696_12[0]),.dout(n11692),.clk(gclk));
	jand g11415(.dina(w_n11691_0[1]),.dinb(w_n10696_11[2]),.dout(n11693),.clk(gclk));
	jxor g11416(.dina(w_n11164_0[0]),.dinb(w_n10701_15[2]),.dout(n11694),.clk(gclk));
	jor g11417(.dina(n11694),.dinb(w_n11662_23[1]),.dout(n11695),.clk(gclk));
	jxor g11418(.dina(n11695),.dinb(w_n11167_0[0]),.dout(n11696),.clk(gclk));
	jor g11419(.dina(w_n11696_0[1]),.dinb(n11693),.dout(n11697),.clk(gclk));
	jand g11420(.dina(w_n11697_0[1]),.dinb(w_n11692_0[1]),.dout(n11698),.clk(gclk));
	jor g11421(.dina(n11698),.dinb(w_n9774_16[0]),.dout(n11699),.clk(gclk));
	jnot g11422(.din(w_n11173_0[0]),.dout(n11700),.clk(gclk));
	jor g11423(.dina(n11700),.dinb(w_n11171_0[0]),.dout(n11701),.clk(gclk));
	jor g11424(.dina(n11701),.dinb(w_n11662_23[0]),.dout(n11702),.clk(gclk));
	jxor g11425(.dina(n11702),.dinb(w_n11182_0[0]),.dout(n11703),.clk(gclk));
	jand g11426(.dina(w_n11692_0[0]),.dinb(w_n9774_15[2]),.dout(n11704),.clk(gclk));
	jand g11427(.dina(n11704),.dinb(w_n11697_0[0]),.dout(n11705),.clk(gclk));
	jor g11428(.dina(w_n11705_0[1]),.dinb(w_n11703_0[1]),.dout(n11706),.clk(gclk));
	jand g11429(.dina(w_n11706_0[1]),.dinb(w_n11699_0[1]),.dout(n11707),.clk(gclk));
	jor g11430(.dina(w_n11707_0[2]),.dinb(w_n9769_12[0]),.dout(n11708),.clk(gclk));
	jand g11431(.dina(w_n11707_0[1]),.dinb(w_n9769_11[2]),.dout(n11709),.clk(gclk));
	jxor g11432(.dina(w_n11184_0[0]),.dinb(w_n9774_15[1]),.dout(n11710),.clk(gclk));
	jor g11433(.dina(n11710),.dinb(w_n11662_22[2]),.dout(n11711),.clk(gclk));
	jxor g11434(.dina(n11711),.dinb(w_n11189_0[0]),.dout(n11712),.clk(gclk));
	jnot g11435(.din(w_n11712_0[1]),.dout(n11713),.clk(gclk));
	jor g11436(.dina(n11713),.dinb(n11709),.dout(n11714),.clk(gclk));
	jand g11437(.dina(w_n11714_0[1]),.dinb(w_n11708_0[1]),.dout(n11715),.clk(gclk));
	jor g11438(.dina(n11715),.dinb(w_n8898_16[2]),.dout(n11716),.clk(gclk));
	jand g11439(.dina(w_n11708_0[0]),.dinb(w_n8898_16[1]),.dout(n11717),.clk(gclk));
	jand g11440(.dina(n11717),.dinb(w_n11714_0[0]),.dout(n11718),.clk(gclk));
	jnot g11441(.din(w_n11193_0[0]),.dout(n11719),.clk(gclk));
	jnot g11442(.din(w_n11662_22[1]),.dout(asqrt_fa_18),.clk(gclk));
	jand g11443(.dina(w_asqrt17_18),.dinb(n11719),.dout(n11721),.clk(gclk));
	jand g11444(.dina(w_n11721_0[1]),.dinb(w_n11200_0[0]),.dout(n11722),.clk(gclk));
	jor g11445(.dina(n11722),.dinb(w_n11198_0[0]),.dout(n11723),.clk(gclk));
	jand g11446(.dina(w_n11721_0[0]),.dinb(w_n11201_0[0]),.dout(n11724),.clk(gclk));
	jnot g11447(.din(n11724),.dout(n11725),.clk(gclk));
	jand g11448(.dina(n11725),.dinb(n11723),.dout(n11726),.clk(gclk));
	jnot g11449(.din(n11726),.dout(n11727),.clk(gclk));
	jor g11450(.dina(w_n11727_0[1]),.dinb(w_n11718_0[1]),.dout(n11728),.clk(gclk));
	jand g11451(.dina(n11728),.dinb(w_n11716_0[1]),.dout(n11729),.clk(gclk));
	jor g11452(.dina(w_n11729_0[2]),.dinb(w_n8893_12[1]),.dout(n11730),.clk(gclk));
	jand g11453(.dina(w_n11729_0[1]),.dinb(w_n8893_12[0]),.dout(n11731),.clk(gclk));
	jnot g11454(.din(w_n11208_0[0]),.dout(n11732),.clk(gclk));
	jxor g11455(.dina(w_n11202_0[0]),.dinb(w_n8898_16[0]),.dout(n11733),.clk(gclk));
	jor g11456(.dina(n11733),.dinb(w_n11662_22[0]),.dout(n11734),.clk(gclk));
	jxor g11457(.dina(n11734),.dinb(n11732),.dout(n11735),.clk(gclk));
	jnot g11458(.din(w_n11735_0[1]),.dout(n11736),.clk(gclk));
	jor g11459(.dina(n11736),.dinb(n11731),.dout(n11737),.clk(gclk));
	jand g11460(.dina(w_n11737_0[1]),.dinb(w_n11730_0[1]),.dout(n11738),.clk(gclk));
	jor g11461(.dina(n11738),.dinb(w_n8058_16[1]),.dout(n11739),.clk(gclk));
	jnot g11462(.din(w_n11213_0[0]),.dout(n11740),.clk(gclk));
	jor g11463(.dina(n11740),.dinb(w_n11211_0[0]),.dout(n11741),.clk(gclk));
	jor g11464(.dina(n11741),.dinb(w_n11662_21[2]),.dout(n11742),.clk(gclk));
	jxor g11465(.dina(n11742),.dinb(w_n11222_0[0]),.dout(n11743),.clk(gclk));
	jand g11466(.dina(w_n11730_0[0]),.dinb(w_n8058_16[0]),.dout(n11744),.clk(gclk));
	jand g11467(.dina(n11744),.dinb(w_n11737_0[0]),.dout(n11745),.clk(gclk));
	jor g11468(.dina(w_n11745_0[1]),.dinb(w_n11743_0[1]),.dout(n11746),.clk(gclk));
	jand g11469(.dina(w_n11746_0[1]),.dinb(w_n11739_0[1]),.dout(n11747),.clk(gclk));
	jor g11470(.dina(w_n11747_0[2]),.dinb(w_n8053_12[1]),.dout(n11748),.clk(gclk));
	jand g11471(.dina(w_n11747_0[1]),.dinb(w_n8053_12[0]),.dout(n11749),.clk(gclk));
	jnot g11472(.din(w_n11229_0[0]),.dout(n11750),.clk(gclk));
	jxor g11473(.dina(w_n11224_0[0]),.dinb(w_n8058_15[2]),.dout(n11751),.clk(gclk));
	jor g11474(.dina(n11751),.dinb(w_n11662_21[1]),.dout(n11752),.clk(gclk));
	jxor g11475(.dina(n11752),.dinb(n11750),.dout(n11753),.clk(gclk));
	jnot g11476(.din(n11753),.dout(n11754),.clk(gclk));
	jor g11477(.dina(w_n11754_0[1]),.dinb(n11749),.dout(n11755),.clk(gclk));
	jand g11478(.dina(w_n11755_0[1]),.dinb(w_n11748_0[1]),.dout(n11756),.clk(gclk));
	jor g11479(.dina(n11756),.dinb(w_n7265_16[2]),.dout(n11757),.clk(gclk));
	jand g11480(.dina(w_n11748_0[0]),.dinb(w_n7265_16[1]),.dout(n11758),.clk(gclk));
	jand g11481(.dina(n11758),.dinb(w_n11755_0[0]),.dout(n11759),.clk(gclk));
	jnot g11482(.din(w_n11232_0[0]),.dout(n11760),.clk(gclk));
	jand g11483(.dina(w_asqrt17_17[2]),.dinb(n11760),.dout(n11761),.clk(gclk));
	jand g11484(.dina(w_n11761_0[1]),.dinb(w_n11239_0[0]),.dout(n11762),.clk(gclk));
	jor g11485(.dina(n11762),.dinb(w_n11237_0[0]),.dout(n11763),.clk(gclk));
	jand g11486(.dina(w_n11761_0[0]),.dinb(w_n11240_0[0]),.dout(n11764),.clk(gclk));
	jnot g11487(.din(n11764),.dout(n11765),.clk(gclk));
	jand g11488(.dina(n11765),.dinb(n11763),.dout(n11766),.clk(gclk));
	jnot g11489(.din(n11766),.dout(n11767),.clk(gclk));
	jor g11490(.dina(w_n11767_0[1]),.dinb(w_n11759_0[1]),.dout(n11768),.clk(gclk));
	jand g11491(.dina(n11768),.dinb(w_n11757_0[1]),.dout(n11769),.clk(gclk));
	jor g11492(.dina(w_n11769_0[1]),.dinb(w_n7260_13[0]),.dout(n11770),.clk(gclk));
	jxor g11493(.dina(w_n11241_0[0]),.dinb(w_n7265_16[0]),.dout(n11771),.clk(gclk));
	jor g11494(.dina(n11771),.dinb(w_n11662_21[0]),.dout(n11772),.clk(gclk));
	jxor g11495(.dina(n11772),.dinb(w_n11246_0[0]),.dout(n11773),.clk(gclk));
	jand g11496(.dina(w_n11769_0[0]),.dinb(w_n7260_12[2]),.dout(n11774),.clk(gclk));
	jor g11497(.dina(w_n11774_0[1]),.dinb(w_n11773_0[1]),.dout(n11775),.clk(gclk));
	jand g11498(.dina(w_n11775_0[2]),.dinb(w_n11770_0[2]),.dout(n11776),.clk(gclk));
	jor g11499(.dina(n11776),.dinb(w_n6505_16[1]),.dout(n11777),.clk(gclk));
	jnot g11500(.din(w_n11251_0[0]),.dout(n11778),.clk(gclk));
	jor g11501(.dina(n11778),.dinb(w_n11249_0[0]),.dout(n11779),.clk(gclk));
	jor g11502(.dina(n11779),.dinb(w_n11662_20[2]),.dout(n11780),.clk(gclk));
	jxor g11503(.dina(n11780),.dinb(w_n11260_0[0]),.dout(n11781),.clk(gclk));
	jand g11504(.dina(w_n11770_0[1]),.dinb(w_n6505_16[0]),.dout(n11782),.clk(gclk));
	jand g11505(.dina(n11782),.dinb(w_n11775_0[1]),.dout(n11783),.clk(gclk));
	jor g11506(.dina(w_n11783_0[1]),.dinb(w_n11781_0[1]),.dout(n11784),.clk(gclk));
	jand g11507(.dina(w_n11784_0[1]),.dinb(w_n11777_0[1]),.dout(n11785),.clk(gclk));
	jor g11508(.dina(w_n11785_0[2]),.dinb(w_n6500_13[1]),.dout(n11786),.clk(gclk));
	jand g11509(.dina(w_n11785_0[1]),.dinb(w_n6500_13[0]),.dout(n11787),.clk(gclk));
	jnot g11510(.din(w_n11263_0[0]),.dout(n11788),.clk(gclk));
	jand g11511(.dina(w_asqrt17_17[1]),.dinb(n11788),.dout(n11789),.clk(gclk));
	jand g11512(.dina(w_n11789_0[1]),.dinb(w_n11268_0[0]),.dout(n11790),.clk(gclk));
	jor g11513(.dina(n11790),.dinb(w_n11267_0[0]),.dout(n11791),.clk(gclk));
	jand g11514(.dina(w_n11789_0[0]),.dinb(w_n11269_0[0]),.dout(n11792),.clk(gclk));
	jnot g11515(.din(n11792),.dout(n11793),.clk(gclk));
	jand g11516(.dina(n11793),.dinb(n11791),.dout(n11794),.clk(gclk));
	jnot g11517(.din(n11794),.dout(n11795),.clk(gclk));
	jor g11518(.dina(w_n11795_0[1]),.dinb(n11787),.dout(n11796),.clk(gclk));
	jand g11519(.dina(w_n11796_0[1]),.dinb(w_n11786_0[1]),.dout(n11797),.clk(gclk));
	jor g11520(.dina(n11797),.dinb(w_n5793_17[0]),.dout(n11798),.clk(gclk));
	jand g11521(.dina(w_n11786_0[0]),.dinb(w_n5793_16[2]),.dout(n11799),.clk(gclk));
	jand g11522(.dina(n11799),.dinb(w_n11796_0[0]),.dout(n11800),.clk(gclk));
	jnot g11523(.din(w_n11271_0[0]),.dout(n11801),.clk(gclk));
	jand g11524(.dina(w_asqrt17_17[0]),.dinb(n11801),.dout(n11802),.clk(gclk));
	jand g11525(.dina(w_n11802_0[1]),.dinb(w_n11278_0[0]),.dout(n11803),.clk(gclk));
	jor g11526(.dina(n11803),.dinb(w_n11276_0[0]),.dout(n11804),.clk(gclk));
	jand g11527(.dina(w_n11802_0[0]),.dinb(w_n11279_0[0]),.dout(n11805),.clk(gclk));
	jnot g11528(.din(n11805),.dout(n11806),.clk(gclk));
	jand g11529(.dina(n11806),.dinb(n11804),.dout(n11807),.clk(gclk));
	jnot g11530(.din(n11807),.dout(n11808),.clk(gclk));
	jor g11531(.dina(w_n11808_0[1]),.dinb(w_n11800_0[1]),.dout(n11809),.clk(gclk));
	jand g11532(.dina(n11809),.dinb(w_n11798_0[1]),.dout(n11810),.clk(gclk));
	jor g11533(.dina(w_n11810_0[1]),.dinb(w_n5788_13[2]),.dout(n11811),.clk(gclk));
	jxor g11534(.dina(w_n11280_0[0]),.dinb(w_n5793_16[1]),.dout(n11812),.clk(gclk));
	jor g11535(.dina(n11812),.dinb(w_n11662_20[1]),.dout(n11813),.clk(gclk));
	jxor g11536(.dina(n11813),.dinb(w_n11291_0[0]),.dout(n11814),.clk(gclk));
	jand g11537(.dina(w_n11810_0[0]),.dinb(w_n5788_13[1]),.dout(n11815),.clk(gclk));
	jor g11538(.dina(w_n11815_0[1]),.dinb(w_n11814_0[1]),.dout(n11816),.clk(gclk));
	jand g11539(.dina(w_n11816_0[2]),.dinb(w_n11811_0[2]),.dout(n11817),.clk(gclk));
	jor g11540(.dina(n11817),.dinb(w_n5121_16[2]),.dout(n11818),.clk(gclk));
	jnot g11541(.din(w_n11296_0[0]),.dout(n11819),.clk(gclk));
	jor g11542(.dina(n11819),.dinb(w_n11294_0[0]),.dout(n11820),.clk(gclk));
	jor g11543(.dina(n11820),.dinb(w_n11662_20[0]),.dout(n11821),.clk(gclk));
	jxor g11544(.dina(n11821),.dinb(w_n11305_0[0]),.dout(n11822),.clk(gclk));
	jand g11545(.dina(w_n11811_0[1]),.dinb(w_n5121_16[1]),.dout(n11823),.clk(gclk));
	jand g11546(.dina(n11823),.dinb(w_n11816_0[1]),.dout(n11824),.clk(gclk));
	jor g11547(.dina(w_n11824_0[1]),.dinb(w_n11822_0[1]),.dout(n11825),.clk(gclk));
	jand g11548(.dina(w_n11825_0[1]),.dinb(w_n11818_0[1]),.dout(n11826),.clk(gclk));
	jor g11549(.dina(w_n11826_0[2]),.dinb(w_n5116_14[0]),.dout(n11827),.clk(gclk));
	jand g11550(.dina(w_n11826_0[1]),.dinb(w_n5116_13[2]),.dout(n11828),.clk(gclk));
	jnot g11551(.din(w_n11308_0[0]),.dout(n11829),.clk(gclk));
	jand g11552(.dina(w_asqrt17_16[2]),.dinb(n11829),.dout(n11830),.clk(gclk));
	jand g11553(.dina(w_n11830_0[1]),.dinb(w_n11313_0[0]),.dout(n11831),.clk(gclk));
	jor g11554(.dina(n11831),.dinb(w_n11312_0[0]),.dout(n11832),.clk(gclk));
	jand g11555(.dina(w_n11830_0[0]),.dinb(w_n11314_0[0]),.dout(n11833),.clk(gclk));
	jnot g11556(.din(n11833),.dout(n11834),.clk(gclk));
	jand g11557(.dina(n11834),.dinb(n11832),.dout(n11835),.clk(gclk));
	jnot g11558(.din(n11835),.dout(n11836),.clk(gclk));
	jor g11559(.dina(w_n11836_0[1]),.dinb(n11828),.dout(n11837),.clk(gclk));
	jand g11560(.dina(w_n11837_0[1]),.dinb(w_n11827_0[1]),.dout(n11838),.clk(gclk));
	jor g11561(.dina(n11838),.dinb(w_n4499_17[2]),.dout(n11839),.clk(gclk));
	jand g11562(.dina(w_n11827_0[0]),.dinb(w_n4499_17[1]),.dout(n11840),.clk(gclk));
	jand g11563(.dina(n11840),.dinb(w_n11837_0[0]),.dout(n11841),.clk(gclk));
	jnot g11564(.din(w_n11316_0[0]),.dout(n11842),.clk(gclk));
	jand g11565(.dina(w_asqrt17_16[1]),.dinb(n11842),.dout(n11843),.clk(gclk));
	jand g11566(.dina(w_n11843_0[1]),.dinb(w_n11323_0[0]),.dout(n11844),.clk(gclk));
	jor g11567(.dina(n11844),.dinb(w_n11321_0[0]),.dout(n11845),.clk(gclk));
	jand g11568(.dina(w_n11843_0[0]),.dinb(w_n11324_0[0]),.dout(n11846),.clk(gclk));
	jnot g11569(.din(n11846),.dout(n11847),.clk(gclk));
	jand g11570(.dina(n11847),.dinb(n11845),.dout(n11848),.clk(gclk));
	jnot g11571(.din(n11848),.dout(n11849),.clk(gclk));
	jor g11572(.dina(w_n11849_0[1]),.dinb(w_n11841_0[1]),.dout(n11850),.clk(gclk));
	jand g11573(.dina(n11850),.dinb(w_n11839_0[1]),.dout(n11851),.clk(gclk));
	jor g11574(.dina(w_n11851_0[1]),.dinb(w_n4494_14[2]),.dout(n11852),.clk(gclk));
	jxor g11575(.dina(w_n11325_0[0]),.dinb(w_n4499_17[0]),.dout(n11853),.clk(gclk));
	jor g11576(.dina(n11853),.dinb(w_n11662_19[2]),.dout(n11854),.clk(gclk));
	jxor g11577(.dina(n11854),.dinb(w_n11336_0[0]),.dout(n11855),.clk(gclk));
	jand g11578(.dina(w_n11851_0[0]),.dinb(w_n4494_14[1]),.dout(n11856),.clk(gclk));
	jor g11579(.dina(w_n11856_0[1]),.dinb(w_n11855_0[1]),.dout(n11857),.clk(gclk));
	jand g11580(.dina(w_n11857_0[2]),.dinb(w_n11852_0[2]),.dout(n11858),.clk(gclk));
	jor g11581(.dina(n11858),.dinb(w_n3912_17[1]),.dout(n11859),.clk(gclk));
	jnot g11582(.din(w_n11341_0[0]),.dout(n11860),.clk(gclk));
	jor g11583(.dina(n11860),.dinb(w_n11339_0[0]),.dout(n11861),.clk(gclk));
	jor g11584(.dina(n11861),.dinb(w_n11662_19[1]),.dout(n11862),.clk(gclk));
	jxor g11585(.dina(n11862),.dinb(w_n11350_0[0]),.dout(n11863),.clk(gclk));
	jand g11586(.dina(w_n11852_0[1]),.dinb(w_n3912_17[0]),.dout(n11864),.clk(gclk));
	jand g11587(.dina(n11864),.dinb(w_n11857_0[1]),.dout(n11865),.clk(gclk));
	jor g11588(.dina(w_n11865_0[1]),.dinb(w_n11863_0[1]),.dout(n11866),.clk(gclk));
	jand g11589(.dina(w_n11866_0[1]),.dinb(w_n11859_0[1]),.dout(n11867),.clk(gclk));
	jor g11590(.dina(w_n11867_0[2]),.dinb(w_n3907_15[0]),.dout(n11868),.clk(gclk));
	jand g11591(.dina(w_n11867_0[1]),.dinb(w_n3907_14[2]),.dout(n11869),.clk(gclk));
	jnot g11592(.din(w_n11353_0[0]),.dout(n11870),.clk(gclk));
	jand g11593(.dina(w_asqrt17_16[0]),.dinb(n11870),.dout(n11871),.clk(gclk));
	jand g11594(.dina(w_n11871_0[1]),.dinb(w_n11358_0[0]),.dout(n11872),.clk(gclk));
	jor g11595(.dina(n11872),.dinb(w_n11357_0[0]),.dout(n11873),.clk(gclk));
	jand g11596(.dina(w_n11871_0[0]),.dinb(w_n11359_0[0]),.dout(n11874),.clk(gclk));
	jnot g11597(.din(n11874),.dout(n11875),.clk(gclk));
	jand g11598(.dina(n11875),.dinb(n11873),.dout(n11876),.clk(gclk));
	jnot g11599(.din(n11876),.dout(n11877),.clk(gclk));
	jor g11600(.dina(w_n11877_0[1]),.dinb(n11869),.dout(n11878),.clk(gclk));
	jand g11601(.dina(w_n11878_0[1]),.dinb(w_n11868_0[1]),.dout(n11879),.clk(gclk));
	jor g11602(.dina(n11879),.dinb(w_n3376_18[1]),.dout(n11880),.clk(gclk));
	jand g11603(.dina(w_n11868_0[0]),.dinb(w_n3376_18[0]),.dout(n11881),.clk(gclk));
	jand g11604(.dina(n11881),.dinb(w_n11878_0[0]),.dout(n11882),.clk(gclk));
	jnot g11605(.din(w_n11361_0[0]),.dout(n11883),.clk(gclk));
	jand g11606(.dina(w_asqrt17_15[2]),.dinb(n11883),.dout(n11884),.clk(gclk));
	jand g11607(.dina(w_n11884_0[1]),.dinb(w_n11368_0[0]),.dout(n11885),.clk(gclk));
	jor g11608(.dina(n11885),.dinb(w_n11366_0[0]),.dout(n11886),.clk(gclk));
	jand g11609(.dina(w_n11884_0[0]),.dinb(w_n11369_0[0]),.dout(n11887),.clk(gclk));
	jnot g11610(.din(n11887),.dout(n11888),.clk(gclk));
	jand g11611(.dina(n11888),.dinb(n11886),.dout(n11889),.clk(gclk));
	jnot g11612(.din(n11889),.dout(n11890),.clk(gclk));
	jor g11613(.dina(w_n11890_0[1]),.dinb(w_n11882_0[1]),.dout(n11891),.clk(gclk));
	jand g11614(.dina(n11891),.dinb(w_n11880_0[1]),.dout(n11892),.clk(gclk));
	jor g11615(.dina(w_n11892_0[1]),.dinb(w_n3371_15[1]),.dout(n11893),.clk(gclk));
	jxor g11616(.dina(w_n11370_0[0]),.dinb(w_n3376_17[2]),.dout(n11894),.clk(gclk));
	jor g11617(.dina(n11894),.dinb(w_n11662_19[0]),.dout(n11895),.clk(gclk));
	jxor g11618(.dina(n11895),.dinb(w_n11381_0[0]),.dout(n11896),.clk(gclk));
	jand g11619(.dina(w_n11892_0[0]),.dinb(w_n3371_15[0]),.dout(n11897),.clk(gclk));
	jor g11620(.dina(w_n11897_0[1]),.dinb(w_n11896_0[1]),.dout(n11898),.clk(gclk));
	jand g11621(.dina(w_n11898_0[2]),.dinb(w_n11893_0[2]),.dout(n11899),.clk(gclk));
	jor g11622(.dina(n11899),.dinb(w_n2875_18[0]),.dout(n11900),.clk(gclk));
	jnot g11623(.din(w_n11386_0[0]),.dout(n11901),.clk(gclk));
	jor g11624(.dina(n11901),.dinb(w_n11384_0[0]),.dout(n11902),.clk(gclk));
	jor g11625(.dina(n11902),.dinb(w_n11662_18[2]),.dout(n11903),.clk(gclk));
	jxor g11626(.dina(n11903),.dinb(w_n11395_0[0]),.dout(n11904),.clk(gclk));
	jand g11627(.dina(w_n11893_0[1]),.dinb(w_n2875_17[2]),.dout(n11905),.clk(gclk));
	jand g11628(.dina(n11905),.dinb(w_n11898_0[1]),.dout(n11906),.clk(gclk));
	jor g11629(.dina(w_n11906_0[1]),.dinb(w_n11904_0[1]),.dout(n11907),.clk(gclk));
	jand g11630(.dina(w_n11907_0[1]),.dinb(w_n11900_0[1]),.dout(n11908),.clk(gclk));
	jor g11631(.dina(w_n11908_0[2]),.dinb(w_n2870_15[2]),.dout(n11909),.clk(gclk));
	jand g11632(.dina(w_n11908_0[1]),.dinb(w_n2870_15[1]),.dout(n11910),.clk(gclk));
	jnot g11633(.din(w_n11398_0[0]),.dout(n11911),.clk(gclk));
	jand g11634(.dina(w_asqrt17_15[1]),.dinb(n11911),.dout(n11912),.clk(gclk));
	jand g11635(.dina(w_n11912_0[1]),.dinb(w_n11403_0[0]),.dout(n11913),.clk(gclk));
	jor g11636(.dina(n11913),.dinb(w_n11402_0[0]),.dout(n11914),.clk(gclk));
	jand g11637(.dina(w_n11912_0[0]),.dinb(w_n11404_0[0]),.dout(n11915),.clk(gclk));
	jnot g11638(.din(n11915),.dout(n11916),.clk(gclk));
	jand g11639(.dina(n11916),.dinb(n11914),.dout(n11917),.clk(gclk));
	jnot g11640(.din(n11917),.dout(n11918),.clk(gclk));
	jor g11641(.dina(w_n11918_0[1]),.dinb(n11910),.dout(n11919),.clk(gclk));
	jand g11642(.dina(w_n11919_0[1]),.dinb(w_n11909_0[1]),.dout(n11920),.clk(gclk));
	jor g11643(.dina(n11920),.dinb(w_n2425_18[2]),.dout(n11921),.clk(gclk));
	jand g11644(.dina(w_n11909_0[0]),.dinb(w_n2425_18[1]),.dout(n11922),.clk(gclk));
	jand g11645(.dina(n11922),.dinb(w_n11919_0[0]),.dout(n11923),.clk(gclk));
	jnot g11646(.din(w_n11406_0[0]),.dout(n11924),.clk(gclk));
	jand g11647(.dina(w_asqrt17_15[0]),.dinb(n11924),.dout(n11925),.clk(gclk));
	jand g11648(.dina(w_n11925_0[1]),.dinb(w_n11413_0[0]),.dout(n11926),.clk(gclk));
	jor g11649(.dina(n11926),.dinb(w_n11411_0[0]),.dout(n11927),.clk(gclk));
	jand g11650(.dina(w_n11925_0[0]),.dinb(w_n11414_0[0]),.dout(n11928),.clk(gclk));
	jnot g11651(.din(n11928),.dout(n11929),.clk(gclk));
	jand g11652(.dina(n11929),.dinb(n11927),.dout(n11930),.clk(gclk));
	jnot g11653(.din(n11930),.dout(n11931),.clk(gclk));
	jor g11654(.dina(w_n11931_0[1]),.dinb(w_n11923_0[1]),.dout(n11932),.clk(gclk));
	jand g11655(.dina(n11932),.dinb(w_n11921_0[1]),.dout(n11933),.clk(gclk));
	jor g11656(.dina(w_n11933_0[1]),.dinb(w_n2420_16[1]),.dout(n11934),.clk(gclk));
	jxor g11657(.dina(w_n11415_0[0]),.dinb(w_n2425_18[0]),.dout(n11935),.clk(gclk));
	jor g11658(.dina(n11935),.dinb(w_n11662_18[1]),.dout(n11936),.clk(gclk));
	jxor g11659(.dina(n11936),.dinb(w_n11426_0[0]),.dout(n11937),.clk(gclk));
	jand g11660(.dina(w_n11933_0[0]),.dinb(w_n2420_16[0]),.dout(n11938),.clk(gclk));
	jor g11661(.dina(w_n11938_0[1]),.dinb(w_n11937_0[1]),.dout(n11939),.clk(gclk));
	jand g11662(.dina(w_n11939_0[2]),.dinb(w_n11934_0[2]),.dout(n11940),.clk(gclk));
	jor g11663(.dina(n11940),.dinb(w_n2010_18[1]),.dout(n11941),.clk(gclk));
	jand g11664(.dina(w_n11934_0[1]),.dinb(w_n2010_18[0]),.dout(n11942),.clk(gclk));
	jand g11665(.dina(n11942),.dinb(w_n11939_0[1]),.dout(n11943),.clk(gclk));
	jnot g11666(.din(w_n11429_0[0]),.dout(n11944),.clk(gclk));
	jand g11667(.dina(w_asqrt17_14[2]),.dinb(n11944),.dout(n11945),.clk(gclk));
	jand g11668(.dina(w_n11945_0[1]),.dinb(w_n11436_0[0]),.dout(n11946),.clk(gclk));
	jor g11669(.dina(n11946),.dinb(w_n11434_0[0]),.dout(n11947),.clk(gclk));
	jand g11670(.dina(w_n11945_0[0]),.dinb(w_n11437_0[0]),.dout(n11948),.clk(gclk));
	jnot g11671(.din(n11948),.dout(n11949),.clk(gclk));
	jand g11672(.dina(n11949),.dinb(n11947),.dout(n11950),.clk(gclk));
	jnot g11673(.din(n11950),.dout(n11951),.clk(gclk));
	jor g11674(.dina(w_n11951_0[1]),.dinb(w_n11943_0[1]),.dout(n11952),.clk(gclk));
	jand g11675(.dina(n11952),.dinb(w_n11941_0[1]),.dout(n11953),.clk(gclk));
	jor g11676(.dina(w_n11953_0[2]),.dinb(w_n2005_16[2]),.dout(n11954),.clk(gclk));
	jnot g11677(.din(w_n11665_0[1]),.dout(n11955),.clk(gclk));
	jand g11678(.dina(w_n11953_0[1]),.dinb(w_n2005_16[1]),.dout(n11956),.clk(gclk));
	jor g11679(.dina(n11956),.dinb(n11955),.dout(n11957),.clk(gclk));
	jand g11680(.dina(w_n11957_0[1]),.dinb(w_n11954_0[1]),.dout(n11958),.clk(gclk));
	jor g11681(.dina(n11958),.dinb(w_n1646_19[2]),.dout(n11959),.clk(gclk));
	jnot g11682(.din(w_n11446_0[0]),.dout(n11960),.clk(gclk));
	jor g11683(.dina(n11960),.dinb(w_n11444_0[0]),.dout(n11961),.clk(gclk));
	jor g11684(.dina(n11961),.dinb(w_n11662_18[0]),.dout(n11962),.clk(gclk));
	jxor g11685(.dina(n11962),.dinb(w_n11455_0[0]),.dout(n11963),.clk(gclk));
	jand g11686(.dina(w_n11954_0[0]),.dinb(w_n1646_19[1]),.dout(n11964),.clk(gclk));
	jand g11687(.dina(n11964),.dinb(w_n11957_0[0]),.dout(n11965),.clk(gclk));
	jor g11688(.dina(w_n11965_0[1]),.dinb(w_n11963_0[1]),.dout(n11966),.clk(gclk));
	jand g11689(.dina(w_n11966_0[1]),.dinb(w_n11959_0[1]),.dout(n11967),.clk(gclk));
	jor g11690(.dina(w_n11967_0[1]),.dinb(w_n1641_17[0]),.dout(n11968),.clk(gclk));
	jxor g11691(.dina(w_n11457_0[0]),.dinb(w_n1646_19[0]),.dout(n11969),.clk(gclk));
	jor g11692(.dina(n11969),.dinb(w_n11662_17[2]),.dout(n11970),.clk(gclk));
	jxor g11693(.dina(n11970),.dinb(w_n11468_0[0]),.dout(n11971),.clk(gclk));
	jand g11694(.dina(w_n11967_0[0]),.dinb(w_n1641_16[2]),.dout(n11972),.clk(gclk));
	jor g11695(.dina(w_n11972_0[1]),.dinb(w_n11971_0[1]),.dout(n11973),.clk(gclk));
	jand g11696(.dina(w_n11973_0[2]),.dinb(w_n11968_0[2]),.dout(n11974),.clk(gclk));
	jor g11697(.dina(n11974),.dinb(w_n1317_19[1]),.dout(n11975),.clk(gclk));
	jnot g11698(.din(w_n11473_0[0]),.dout(n11976),.clk(gclk));
	jor g11699(.dina(n11976),.dinb(w_n11471_0[0]),.dout(n11977),.clk(gclk));
	jor g11700(.dina(n11977),.dinb(w_n11662_17[1]),.dout(n11978),.clk(gclk));
	jxor g11701(.dina(n11978),.dinb(w_n11482_0[0]),.dout(n11979),.clk(gclk));
	jand g11702(.dina(w_n11968_0[1]),.dinb(w_n1317_19[0]),.dout(n11980),.clk(gclk));
	jand g11703(.dina(n11980),.dinb(w_n11973_0[1]),.dout(n11981),.clk(gclk));
	jor g11704(.dina(w_n11981_0[1]),.dinb(w_n11979_0[1]),.dout(n11982),.clk(gclk));
	jand g11705(.dina(w_n11982_0[1]),.dinb(w_n11975_0[1]),.dout(n11983),.clk(gclk));
	jor g11706(.dina(w_n11983_0[2]),.dinb(w_n1312_17[1]),.dout(n11984),.clk(gclk));
	jand g11707(.dina(w_n11983_0[1]),.dinb(w_n1312_17[0]),.dout(n11985),.clk(gclk));
	jnot g11708(.din(w_n11485_0[0]),.dout(n11986),.clk(gclk));
	jand g11709(.dina(w_asqrt17_14[1]),.dinb(n11986),.dout(n11987),.clk(gclk));
	jand g11710(.dina(w_n11987_0[1]),.dinb(w_n11490_0[0]),.dout(n11988),.clk(gclk));
	jor g11711(.dina(n11988),.dinb(w_n11489_0[0]),.dout(n11989),.clk(gclk));
	jand g11712(.dina(w_n11987_0[0]),.dinb(w_n11491_0[0]),.dout(n11990),.clk(gclk));
	jnot g11713(.din(n11990),.dout(n11991),.clk(gclk));
	jand g11714(.dina(n11991),.dinb(n11989),.dout(n11992),.clk(gclk));
	jnot g11715(.din(n11992),.dout(n11993),.clk(gclk));
	jor g11716(.dina(w_n11993_0[1]),.dinb(n11985),.dout(n11994),.clk(gclk));
	jand g11717(.dina(w_n11994_0[1]),.dinb(w_n11984_0[1]),.dout(n11995),.clk(gclk));
	jor g11718(.dina(n11995),.dinb(w_n1039_20[0]),.dout(n11996),.clk(gclk));
	jand g11719(.dina(w_n11984_0[0]),.dinb(w_n1039_19[2]),.dout(n11997),.clk(gclk));
	jand g11720(.dina(n11997),.dinb(w_n11994_0[0]),.dout(n11998),.clk(gclk));
	jnot g11721(.din(w_n11493_0[0]),.dout(n11999),.clk(gclk));
	jand g11722(.dina(w_asqrt17_14[0]),.dinb(n11999),.dout(n12000),.clk(gclk));
	jand g11723(.dina(w_n12000_0[1]),.dinb(w_n11500_0[0]),.dout(n12001),.clk(gclk));
	jor g11724(.dina(n12001),.dinb(w_n11498_0[0]),.dout(n12002),.clk(gclk));
	jand g11725(.dina(w_n12000_0[0]),.dinb(w_n11501_0[0]),.dout(n12003),.clk(gclk));
	jnot g11726(.din(n12003),.dout(n12004),.clk(gclk));
	jand g11727(.dina(n12004),.dinb(n12002),.dout(n12005),.clk(gclk));
	jnot g11728(.din(n12005),.dout(n12006),.clk(gclk));
	jor g11729(.dina(w_n12006_0[1]),.dinb(w_n11998_0[1]),.dout(n12007),.clk(gclk));
	jand g11730(.dina(n12007),.dinb(w_n11996_0[1]),.dout(n12008),.clk(gclk));
	jor g11731(.dina(w_n12008_0[1]),.dinb(w_n1034_18[0]),.dout(n12009),.clk(gclk));
	jxor g11732(.dina(w_n11502_0[0]),.dinb(w_n1039_19[1]),.dout(n12010),.clk(gclk));
	jor g11733(.dina(n12010),.dinb(w_n11662_17[0]),.dout(n12011),.clk(gclk));
	jxor g11734(.dina(n12011),.dinb(w_n11513_0[0]),.dout(n12012),.clk(gclk));
	jand g11735(.dina(w_n12008_0[0]),.dinb(w_n1034_17[2]),.dout(n12013),.clk(gclk));
	jor g11736(.dina(w_n12013_0[1]),.dinb(w_n12012_0[1]),.dout(n12014),.clk(gclk));
	jand g11737(.dina(w_n12014_0[2]),.dinb(w_n12009_0[2]),.dout(n12015),.clk(gclk));
	jor g11738(.dina(n12015),.dinb(w_n796_19[2]),.dout(n12016),.clk(gclk));
	jnot g11739(.din(w_n11518_0[0]),.dout(n12017),.clk(gclk));
	jor g11740(.dina(n12017),.dinb(w_n11516_0[0]),.dout(n12018),.clk(gclk));
	jor g11741(.dina(n12018),.dinb(w_n11662_16[2]),.dout(n12019),.clk(gclk));
	jxor g11742(.dina(n12019),.dinb(w_n11527_0[0]),.dout(n12020),.clk(gclk));
	jand g11743(.dina(w_n12009_0[1]),.dinb(w_n796_19[1]),.dout(n12021),.clk(gclk));
	jand g11744(.dina(n12021),.dinb(w_n12014_0[1]),.dout(n12022),.clk(gclk));
	jor g11745(.dina(w_n12022_0[1]),.dinb(w_n12020_0[1]),.dout(n12023),.clk(gclk));
	jand g11746(.dina(w_n12023_0[1]),.dinb(w_n12016_0[1]),.dout(n12024),.clk(gclk));
	jor g11747(.dina(w_n12024_0[2]),.dinb(w_n791_18[1]),.dout(n12025),.clk(gclk));
	jand g11748(.dina(w_n12024_0[1]),.dinb(w_n791_18[0]),.dout(n12026),.clk(gclk));
	jnot g11749(.din(w_n11530_0[0]),.dout(n12027),.clk(gclk));
	jand g11750(.dina(w_asqrt17_13[2]),.dinb(n12027),.dout(n12028),.clk(gclk));
	jand g11751(.dina(w_n12028_0[1]),.dinb(w_n11535_0[0]),.dout(n12029),.clk(gclk));
	jor g11752(.dina(n12029),.dinb(w_n11534_0[0]),.dout(n12030),.clk(gclk));
	jand g11753(.dina(w_n12028_0[0]),.dinb(w_n11536_0[0]),.dout(n12031),.clk(gclk));
	jnot g11754(.din(n12031),.dout(n12032),.clk(gclk));
	jand g11755(.dina(n12032),.dinb(n12030),.dout(n12033),.clk(gclk));
	jnot g11756(.din(n12033),.dout(n12034),.clk(gclk));
	jor g11757(.dina(w_n12034_0[1]),.dinb(n12026),.dout(n12035),.clk(gclk));
	jand g11758(.dina(w_n12035_0[1]),.dinb(w_n12025_0[1]),.dout(n12036),.clk(gclk));
	jor g11759(.dina(n12036),.dinb(w_n595_20[1]),.dout(n12037),.clk(gclk));
	jand g11760(.dina(w_n12025_0[0]),.dinb(w_n595_20[0]),.dout(n12038),.clk(gclk));
	jand g11761(.dina(n12038),.dinb(w_n12035_0[0]),.dout(n12039),.clk(gclk));
	jnot g11762(.din(w_n11538_0[0]),.dout(n12040),.clk(gclk));
	jand g11763(.dina(w_asqrt17_13[1]),.dinb(n12040),.dout(n12041),.clk(gclk));
	jand g11764(.dina(w_n12041_0[1]),.dinb(w_n11545_0[0]),.dout(n12042),.clk(gclk));
	jor g11765(.dina(n12042),.dinb(w_n11543_0[0]),.dout(n12043),.clk(gclk));
	jand g11766(.dina(w_n12041_0[0]),.dinb(w_n11546_0[0]),.dout(n12044),.clk(gclk));
	jnot g11767(.din(n12044),.dout(n12045),.clk(gclk));
	jand g11768(.dina(n12045),.dinb(n12043),.dout(n12046),.clk(gclk));
	jnot g11769(.din(n12046),.dout(n12047),.clk(gclk));
	jor g11770(.dina(w_n12047_0[1]),.dinb(w_n12039_0[1]),.dout(n12048),.clk(gclk));
	jand g11771(.dina(n12048),.dinb(w_n12037_0[1]),.dout(n12049),.clk(gclk));
	jor g11772(.dina(w_n12049_0[1]),.dinb(w_n590_18[2]),.dout(n12050),.clk(gclk));
	jxor g11773(.dina(w_n11547_0[0]),.dinb(w_n595_19[2]),.dout(n12051),.clk(gclk));
	jor g11774(.dina(n12051),.dinb(w_n11662_16[1]),.dout(n12052),.clk(gclk));
	jxor g11775(.dina(n12052),.dinb(w_n11558_0[0]),.dout(n12053),.clk(gclk));
	jand g11776(.dina(w_n12049_0[0]),.dinb(w_n590_18[1]),.dout(n12054),.clk(gclk));
	jor g11777(.dina(w_n12054_0[1]),.dinb(w_n12053_0[1]),.dout(n12055),.clk(gclk));
	jand g11778(.dina(w_n12055_0[2]),.dinb(w_n12050_0[2]),.dout(n12056),.clk(gclk));
	jor g11779(.dina(n12056),.dinb(w_n430_20[0]),.dout(n12057),.clk(gclk));
	jnot g11780(.din(w_n11563_0[0]),.dout(n12058),.clk(gclk));
	jor g11781(.dina(n12058),.dinb(w_n11561_0[0]),.dout(n12059),.clk(gclk));
	jor g11782(.dina(n12059),.dinb(w_n11662_16[0]),.dout(n12060),.clk(gclk));
	jxor g11783(.dina(n12060),.dinb(w_n11572_0[0]),.dout(n12061),.clk(gclk));
	jand g11784(.dina(w_n12050_0[1]),.dinb(w_n430_19[2]),.dout(n12062),.clk(gclk));
	jand g11785(.dina(n12062),.dinb(w_n12055_0[1]),.dout(n12063),.clk(gclk));
	jor g11786(.dina(w_n12063_0[1]),.dinb(w_n12061_0[1]),.dout(n12064),.clk(gclk));
	jand g11787(.dina(w_n12064_0[1]),.dinb(w_n12057_0[1]),.dout(n12065),.clk(gclk));
	jor g11788(.dina(w_n12065_0[2]),.dinb(w_n425_19[0]),.dout(n12066),.clk(gclk));
	jand g11789(.dina(w_n12065_0[1]),.dinb(w_n425_18[2]),.dout(n12067),.clk(gclk));
	jnot g11790(.din(w_n11575_0[0]),.dout(n12068),.clk(gclk));
	jand g11791(.dina(w_asqrt17_13[0]),.dinb(n12068),.dout(n12069),.clk(gclk));
	jand g11792(.dina(w_n12069_0[1]),.dinb(w_n11580_0[0]),.dout(n12070),.clk(gclk));
	jor g11793(.dina(n12070),.dinb(w_n11579_0[0]),.dout(n12071),.clk(gclk));
	jand g11794(.dina(w_n12069_0[0]),.dinb(w_n11581_0[0]),.dout(n12072),.clk(gclk));
	jnot g11795(.din(n12072),.dout(n12073),.clk(gclk));
	jand g11796(.dina(n12073),.dinb(n12071),.dout(n12074),.clk(gclk));
	jnot g11797(.din(n12074),.dout(n12075),.clk(gclk));
	jor g11798(.dina(w_n12075_0[1]),.dinb(n12067),.dout(n12076),.clk(gclk));
	jand g11799(.dina(w_n12076_0[1]),.dinb(w_n12066_0[1]),.dout(n12077),.clk(gclk));
	jor g11800(.dina(n12077),.dinb(w_n305_20[2]),.dout(n12078),.clk(gclk));
	jand g11801(.dina(w_n12066_0[0]),.dinb(w_n305_20[1]),.dout(n12079),.clk(gclk));
	jand g11802(.dina(n12079),.dinb(w_n12076_0[0]),.dout(n12080),.clk(gclk));
	jnot g11803(.din(w_n11583_0[0]),.dout(n12081),.clk(gclk));
	jand g11804(.dina(w_asqrt17_12[2]),.dinb(n12081),.dout(n12082),.clk(gclk));
	jand g11805(.dina(w_n12082_0[1]),.dinb(w_n11590_0[0]),.dout(n12083),.clk(gclk));
	jor g11806(.dina(n12083),.dinb(w_n11588_0[0]),.dout(n12084),.clk(gclk));
	jand g11807(.dina(w_n12082_0[0]),.dinb(w_n11591_0[0]),.dout(n12085),.clk(gclk));
	jnot g11808(.din(n12085),.dout(n12086),.clk(gclk));
	jand g11809(.dina(n12086),.dinb(n12084),.dout(n12087),.clk(gclk));
	jnot g11810(.din(n12087),.dout(n12088),.clk(gclk));
	jor g11811(.dina(w_n12088_0[1]),.dinb(w_n12080_0[1]),.dout(n12089),.clk(gclk));
	jand g11812(.dina(n12089),.dinb(w_n12078_0[1]),.dout(n12090),.clk(gclk));
	jor g11813(.dina(w_n12090_0[1]),.dinb(w_n290_20[0]),.dout(n12091),.clk(gclk));
	jxor g11814(.dina(w_n11592_0[0]),.dinb(w_n305_20[0]),.dout(n12092),.clk(gclk));
	jor g11815(.dina(n12092),.dinb(w_n11662_15[2]),.dout(n12093),.clk(gclk));
	jxor g11816(.dina(n12093),.dinb(w_n11603_0[0]),.dout(n12094),.clk(gclk));
	jand g11817(.dina(w_n12090_0[0]),.dinb(w_n290_19[2]),.dout(n12095),.clk(gclk));
	jor g11818(.dina(w_n12095_0[1]),.dinb(w_n12094_0[1]),.dout(n12096),.clk(gclk));
	jand g11819(.dina(w_n12096_0[2]),.dinb(w_n12091_0[2]),.dout(n12097),.clk(gclk));
	jor g11820(.dina(n12097),.dinb(w_n223_20[1]),.dout(n12098),.clk(gclk));
	jnot g11821(.din(w_n11608_0[0]),.dout(n12099),.clk(gclk));
	jor g11822(.dina(n12099),.dinb(w_n11606_0[0]),.dout(n12100),.clk(gclk));
	jor g11823(.dina(n12100),.dinb(w_n11662_15[1]),.dout(n12101),.clk(gclk));
	jxor g11824(.dina(n12101),.dinb(w_n11617_0[0]),.dout(n12102),.clk(gclk));
	jand g11825(.dina(w_n12091_0[1]),.dinb(w_n223_20[0]),.dout(n12103),.clk(gclk));
	jand g11826(.dina(n12103),.dinb(w_n12096_0[1]),.dout(n12104),.clk(gclk));
	jor g11827(.dina(w_n12104_0[1]),.dinb(w_n12102_0[1]),.dout(n12105),.clk(gclk));
	jand g11828(.dina(w_n12105_0[1]),.dinb(w_n12098_0[1]),.dout(n12106),.clk(gclk));
	jor g11829(.dina(w_n12106_0[2]),.dinb(w_n199_23[1]),.dout(n12107),.clk(gclk));
	jand g11830(.dina(w_n12106_0[1]),.dinb(w_n199_23[0]),.dout(n12108),.clk(gclk));
	jnot g11831(.din(w_n11620_0[0]),.dout(n12109),.clk(gclk));
	jand g11832(.dina(w_asqrt17_12[1]),.dinb(n12109),.dout(n12110),.clk(gclk));
	jand g11833(.dina(w_n12110_0[1]),.dinb(w_n11625_0[0]),.dout(n12111),.clk(gclk));
	jor g11834(.dina(n12111),.dinb(w_n11624_0[0]),.dout(n12112),.clk(gclk));
	jand g11835(.dina(w_n12110_0[0]),.dinb(w_n11626_0[0]),.dout(n12113),.clk(gclk));
	jnot g11836(.din(n12113),.dout(n12114),.clk(gclk));
	jand g11837(.dina(n12114),.dinb(n12112),.dout(n12115),.clk(gclk));
	jnot g11838(.din(n12115),.dout(n12116),.clk(gclk));
	jor g11839(.dina(w_n12116_0[1]),.dinb(n12108),.dout(n12117),.clk(gclk));
	jand g11840(.dina(n12117),.dinb(n12107),.dout(n12118),.clk(gclk));
	jnot g11841(.din(w_n11628_0[0]),.dout(n12119),.clk(gclk));
	jand g11842(.dina(w_asqrt17_12[0]),.dinb(n12119),.dout(n12120),.clk(gclk));
	jand g11843(.dina(w_n12120_0[1]),.dinb(w_n11635_0[0]),.dout(n12121),.clk(gclk));
	jor g11844(.dina(n12121),.dinb(w_n11633_0[0]),.dout(n12122),.clk(gclk));
	jand g11845(.dina(w_n12120_0[0]),.dinb(w_n11636_0[0]),.dout(n12123),.clk(gclk));
	jnot g11846(.din(n12123),.dout(n12124),.clk(gclk));
	jand g11847(.dina(n12124),.dinb(n12122),.dout(n12125),.clk(gclk));
	jnot g11848(.din(w_n12125_0[2]),.dout(n12126),.clk(gclk));
	jand g11849(.dina(w_asqrt17_11[2]),.dinb(w_n11650_0[1]),.dout(n12127),.clk(gclk));
	jand g11850(.dina(w_n12127_0[1]),.dinb(w_n11637_1[0]),.dout(n12128),.clk(gclk));
	jor g11851(.dina(n12128),.dinb(w_n11684_0[0]),.dout(n12129),.clk(gclk));
	jor g11852(.dina(n12129),.dinb(w_n12126_0[1]),.dout(n12130),.clk(gclk));
	jor g11853(.dina(n12130),.dinb(w_n12118_0[2]),.dout(n12131),.clk(gclk));
	jand g11854(.dina(n12131),.dinb(w_n194_22[1]),.dout(n12132),.clk(gclk));
	jand g11855(.dina(w_n12126_0[0]),.dinb(w_n12118_0[1]),.dout(n12133),.clk(gclk));
	jor g11856(.dina(w_n12127_0[0]),.dinb(w_n11637_0[2]),.dout(n12134),.clk(gclk));
	jand g11857(.dina(w_n11650_0[0]),.dinb(w_n11637_0[1]),.dout(n12135),.clk(gclk));
	jor g11858(.dina(n12135),.dinb(w_n194_22[0]),.dout(n12136),.clk(gclk));
	jnot g11859(.din(n12136),.dout(n12137),.clk(gclk));
	jand g11860(.dina(n12137),.dinb(n12134),.dout(n12138),.clk(gclk));
	jor g11861(.dina(w_n12138_0[1]),.dinb(w_n12133_0[2]),.dout(n12141),.clk(gclk));
	jor g11862(.dina(n12141),.dinb(w_n12132_0[1]),.dout(asqrt_fa_17),.clk(gclk));
	jxor g11863(.dina(w_n11953_0[0]),.dinb(w_n2005_16[0]),.dout(n12143),.clk(gclk));
	jand g11864(.dina(n12143),.dinb(w_asqrt16_31),.dout(n12144),.clk(gclk));
	jxor g11865(.dina(n12144),.dinb(w_n11665_0[0]),.dout(n12145),.clk(gclk));
	jnot g11866(.din(w_n12145_0[1]),.dout(n12146),.clk(gclk));
	jand g11867(.dina(w_asqrt16_30[2]),.dinb(w_a32_0[0]),.dout(n12147),.clk(gclk));
	jnot g11868(.din(w_a30_0[1]),.dout(n12148),.clk(gclk));
	jnot g11869(.din(w_a31_0[1]),.dout(n12149),.clk(gclk));
	jand g11870(.dina(w_n11667_1[0]),.dinb(w_n12149_0[1]),.dout(n12150),.clk(gclk));
	jand g11871(.dina(n12150),.dinb(w_n12148_1[1]),.dout(n12151),.clk(gclk));
	jor g11872(.dina(n12151),.dinb(n12147),.dout(n12152),.clk(gclk));
	jand g11873(.dina(w_n12152_0[2]),.dinb(w_asqrt17_11[1]),.dout(n12153),.clk(gclk));
	jand g11874(.dina(w_asqrt16_30[1]),.dinb(w_n11667_0[2]),.dout(n12154),.clk(gclk));
	jxor g11875(.dina(w_n12154_0[1]),.dinb(w_n11668_0[1]),.dout(n12155),.clk(gclk));
	jor g11876(.dina(w_n12152_0[1]),.dinb(w_asqrt17_11[0]),.dout(n12156),.clk(gclk));
	jand g11877(.dina(n12156),.dinb(w_n12155_0[1]),.dout(n12157),.clk(gclk));
	jor g11878(.dina(w_n12157_0[1]),.dinb(w_n12153_0[1]),.dout(n12158),.clk(gclk));
	jand g11879(.dina(n12158),.dinb(w_asqrt18_15[1]),.dout(n12159),.clk(gclk));
	jor g11880(.dina(w_n12153_0[0]),.dinb(w_asqrt18_15[0]),.dout(n12160),.clk(gclk));
	jor g11881(.dina(n12160),.dinb(w_n12157_0[0]),.dout(n12161),.clk(gclk));
	jand g11882(.dina(w_n12154_0[0]),.dinb(w_n11668_0[0]),.dout(n12162),.clk(gclk));
	jnot g11883(.din(w_n12132_0[0]),.dout(n12163),.clk(gclk));
	jnot g11884(.din(w_n12133_0[1]),.dout(n12164),.clk(gclk));
	jnot g11885(.din(w_n12138_0[0]),.dout(n12165),.clk(gclk));
	jand g11886(.dina(n12165),.dinb(w_asqrt17_10[2]),.dout(n12166),.clk(gclk));
	jand g11887(.dina(n12166),.dinb(n12164),.dout(n12167),.clk(gclk));
	jand g11888(.dina(n12167),.dinb(n12163),.dout(n12168),.clk(gclk));
	jor g11889(.dina(n12168),.dinb(n12162),.dout(n12169),.clk(gclk));
	jxor g11890(.dina(n12169),.dinb(w_n11160_0[1]),.dout(n12170),.clk(gclk));
	jand g11891(.dina(w_n12170_0[1]),.dinb(w_n12161_0[1]),.dout(n12171),.clk(gclk));
	jor g11892(.dina(n12171),.dinb(w_n12159_0[1]),.dout(n12172),.clk(gclk));
	jand g11893(.dina(w_n12172_0[2]),.dinb(w_asqrt19_11[0]),.dout(n12173),.clk(gclk));
	jor g11894(.dina(w_n12172_0[1]),.dinb(w_asqrt19_10[2]),.dout(n12174),.clk(gclk));
	jxor g11895(.dina(w_n11672_0[0]),.dinb(w_n11657_10[2]),.dout(n12175),.clk(gclk));
	jand g11896(.dina(n12175),.dinb(w_asqrt16_30[0]),.dout(n12176),.clk(gclk));
	jxor g11897(.dina(n12176),.dinb(w_n11675_0[0]),.dout(n12177),.clk(gclk));
	jnot g11898(.din(w_n12177_0[1]),.dout(n12178),.clk(gclk));
	jand g11899(.dina(n12178),.dinb(n12174),.dout(n12179),.clk(gclk));
	jor g11900(.dina(w_n12179_0[1]),.dinb(w_n12173_0[1]),.dout(n12180),.clk(gclk));
	jand g11901(.dina(n12180),.dinb(w_asqrt20_15[1]),.dout(n12181),.clk(gclk));
	jnot g11902(.din(w_n11681_0[0]),.dout(n12182),.clk(gclk));
	jand g11903(.dina(n12182),.dinb(w_n11679_0[0]),.dout(n12183),.clk(gclk));
	jand g11904(.dina(n12183),.dinb(w_asqrt16_29[2]),.dout(n12184),.clk(gclk));
	jxor g11905(.dina(n12184),.dinb(w_n11689_0[0]),.dout(n12185),.clk(gclk));
	jnot g11906(.din(n12185),.dout(n12186),.clk(gclk));
	jor g11907(.dina(w_n12173_0[0]),.dinb(w_asqrt20_15[0]),.dout(n12187),.clk(gclk));
	jor g11908(.dina(n12187),.dinb(w_n12179_0[0]),.dout(n12188),.clk(gclk));
	jand g11909(.dina(w_n12188_0[1]),.dinb(w_n12186_0[1]),.dout(n12189),.clk(gclk));
	jor g11910(.dina(w_n12189_0[1]),.dinb(w_n12181_0[1]),.dout(n12190),.clk(gclk));
	jand g11911(.dina(w_n12190_0[2]),.dinb(w_asqrt21_11[1]),.dout(n12191),.clk(gclk));
	jor g11912(.dina(w_n12190_0[1]),.dinb(w_asqrt21_11[0]),.dout(n12192),.clk(gclk));
	jnot g11913(.din(w_n11696_0[0]),.dout(n12193),.clk(gclk));
	jxor g11914(.dina(w_n11691_0[0]),.dinb(w_n10696_11[1]),.dout(n12194),.clk(gclk));
	jand g11915(.dina(n12194),.dinb(w_asqrt16_29[1]),.dout(n12195),.clk(gclk));
	jxor g11916(.dina(n12195),.dinb(n12193),.dout(n12196),.clk(gclk));
	jand g11917(.dina(w_n12196_0[1]),.dinb(n12192),.dout(n12197),.clk(gclk));
	jor g11918(.dina(w_n12197_0[1]),.dinb(w_n12191_0[1]),.dout(n12198),.clk(gclk));
	jand g11919(.dina(n12198),.dinb(w_asqrt22_15[1]),.dout(n12199),.clk(gclk));
	jor g11920(.dina(w_n12191_0[0]),.dinb(w_asqrt22_15[0]),.dout(n12200),.clk(gclk));
	jor g11921(.dina(n12200),.dinb(w_n12197_0[0]),.dout(n12201),.clk(gclk));
	jnot g11922(.din(w_n11703_0[0]),.dout(n12202),.clk(gclk));
	jnot g11923(.din(w_n11705_0[0]),.dout(n12203),.clk(gclk));
	jand g11924(.dina(w_asqrt16_29[0]),.dinb(w_n11699_0[0]),.dout(n12204),.clk(gclk));
	jand g11925(.dina(w_n12204_0[1]),.dinb(n12203),.dout(n12205),.clk(gclk));
	jor g11926(.dina(n12205),.dinb(n12202),.dout(n12206),.clk(gclk));
	jnot g11927(.din(w_n11706_0[0]),.dout(n12207),.clk(gclk));
	jand g11928(.dina(w_n12204_0[0]),.dinb(n12207),.dout(n12208),.clk(gclk));
	jnot g11929(.din(n12208),.dout(n12209),.clk(gclk));
	jand g11930(.dina(n12209),.dinb(n12206),.dout(n12210),.clk(gclk));
	jand g11931(.dina(w_n12210_0[1]),.dinb(w_n12201_0[1]),.dout(n12211),.clk(gclk));
	jor g11932(.dina(n12211),.dinb(w_n12199_0[1]),.dout(n12212),.clk(gclk));
	jand g11933(.dina(w_n12212_0[2]),.dinb(w_asqrt23_11[1]),.dout(n12213),.clk(gclk));
	jor g11934(.dina(w_n12212_0[1]),.dinb(w_asqrt23_11[0]),.dout(n12214),.clk(gclk));
	jxor g11935(.dina(w_n11707_0[0]),.dinb(w_n9769_11[1]),.dout(n12215),.clk(gclk));
	jand g11936(.dina(n12215),.dinb(w_asqrt16_28[2]),.dout(n12216),.clk(gclk));
	jxor g11937(.dina(n12216),.dinb(w_n11712_0[0]),.dout(n12217),.clk(gclk));
	jand g11938(.dina(w_n12217_0[1]),.dinb(n12214),.dout(n12218),.clk(gclk));
	jor g11939(.dina(w_n12218_0[1]),.dinb(w_n12213_0[1]),.dout(n12219),.clk(gclk));
	jand g11940(.dina(n12219),.dinb(w_asqrt24_15[1]),.dout(n12220),.clk(gclk));
	jnot g11941(.din(w_n11718_0[0]),.dout(n12221),.clk(gclk));
	jand g11942(.dina(n12221),.dinb(w_n11716_0[0]),.dout(n12222),.clk(gclk));
	jand g11943(.dina(n12222),.dinb(w_asqrt16_28[1]),.dout(n12223),.clk(gclk));
	jxor g11944(.dina(n12223),.dinb(w_n11727_0[0]),.dout(n12224),.clk(gclk));
	jnot g11945(.din(n12224),.dout(n12225),.clk(gclk));
	jor g11946(.dina(w_n12213_0[0]),.dinb(w_asqrt24_15[0]),.dout(n12226),.clk(gclk));
	jor g11947(.dina(n12226),.dinb(w_n12218_0[0]),.dout(n12227),.clk(gclk));
	jand g11948(.dina(w_n12227_0[1]),.dinb(w_n12225_0[1]),.dout(n12228),.clk(gclk));
	jor g11949(.dina(w_n12228_0[1]),.dinb(w_n12220_0[1]),.dout(n12229),.clk(gclk));
	jand g11950(.dina(w_n12229_0[2]),.dinb(w_asqrt25_11[2]),.dout(n12230),.clk(gclk));
	jor g11951(.dina(w_n12229_0[1]),.dinb(w_asqrt25_11[1]),.dout(n12231),.clk(gclk));
	jxor g11952(.dina(w_n11729_0[0]),.dinb(w_n8893_11[2]),.dout(n12232),.clk(gclk));
	jand g11953(.dina(n12232),.dinb(w_asqrt16_28[0]),.dout(n12233),.clk(gclk));
	jxor g11954(.dina(n12233),.dinb(w_n11735_0[0]),.dout(n12234),.clk(gclk));
	jand g11955(.dina(w_n12234_0[1]),.dinb(n12231),.dout(n12235),.clk(gclk));
	jor g11956(.dina(w_n12235_0[1]),.dinb(w_n12230_0[1]),.dout(n12236),.clk(gclk));
	jand g11957(.dina(n12236),.dinb(w_asqrt26_15[1]),.dout(n12237),.clk(gclk));
	jor g11958(.dina(w_n12230_0[0]),.dinb(w_asqrt26_15[0]),.dout(n12238),.clk(gclk));
	jor g11959(.dina(n12238),.dinb(w_n12235_0[0]),.dout(n12239),.clk(gclk));
	jnot g11960(.din(w_n11743_0[0]),.dout(n12240),.clk(gclk));
	jnot g11961(.din(w_n11745_0[0]),.dout(n12241),.clk(gclk));
	jand g11962(.dina(w_asqrt16_27[2]),.dinb(w_n11739_0[0]),.dout(n12242),.clk(gclk));
	jand g11963(.dina(w_n12242_0[1]),.dinb(n12241),.dout(n12243),.clk(gclk));
	jor g11964(.dina(n12243),.dinb(n12240),.dout(n12244),.clk(gclk));
	jnot g11965(.din(w_n11746_0[0]),.dout(n12245),.clk(gclk));
	jand g11966(.dina(w_n12242_0[0]),.dinb(n12245),.dout(n12246),.clk(gclk));
	jnot g11967(.din(n12246),.dout(n12247),.clk(gclk));
	jand g11968(.dina(n12247),.dinb(n12244),.dout(n12248),.clk(gclk));
	jand g11969(.dina(w_n12248_0[1]),.dinb(w_n12239_0[1]),.dout(n12249),.clk(gclk));
	jor g11970(.dina(n12249),.dinb(w_n12237_0[1]),.dout(n12250),.clk(gclk));
	jand g11971(.dina(w_n12250_0[1]),.dinb(w_asqrt27_11[2]),.dout(n12251),.clk(gclk));
	jxor g11972(.dina(w_n11747_0[0]),.dinb(w_n8053_11[2]),.dout(n12252),.clk(gclk));
	jand g11973(.dina(n12252),.dinb(w_asqrt16_27[1]),.dout(n12253),.clk(gclk));
	jxor g11974(.dina(n12253),.dinb(w_n11754_0[0]),.dout(n12254),.clk(gclk));
	jnot g11975(.din(n12254),.dout(n12255),.clk(gclk));
	jor g11976(.dina(w_n12250_0[0]),.dinb(w_asqrt27_11[1]),.dout(n12256),.clk(gclk));
	jand g11977(.dina(w_n12256_0[1]),.dinb(w_n12255_0[1]),.dout(n12257),.clk(gclk));
	jor g11978(.dina(w_n12257_0[2]),.dinb(w_n12251_0[2]),.dout(n12258),.clk(gclk));
	jand g11979(.dina(n12258),.dinb(w_asqrt28_15[1]),.dout(n12259),.clk(gclk));
	jnot g11980(.din(w_n11759_0[0]),.dout(n12260),.clk(gclk));
	jand g11981(.dina(n12260),.dinb(w_n11757_0[0]),.dout(n12261),.clk(gclk));
	jand g11982(.dina(n12261),.dinb(w_asqrt16_27[0]),.dout(n12262),.clk(gclk));
	jxor g11983(.dina(n12262),.dinb(w_n11767_0[0]),.dout(n12263),.clk(gclk));
	jnot g11984(.din(n12263),.dout(n12264),.clk(gclk));
	jor g11985(.dina(w_n12251_0[1]),.dinb(w_asqrt28_15[0]),.dout(n12265),.clk(gclk));
	jor g11986(.dina(n12265),.dinb(w_n12257_0[1]),.dout(n12266),.clk(gclk));
	jand g11987(.dina(w_n12266_0[1]),.dinb(w_n12264_0[1]),.dout(n12267),.clk(gclk));
	jor g11988(.dina(w_n12267_0[1]),.dinb(w_n12259_0[1]),.dout(n12268),.clk(gclk));
	jand g11989(.dina(w_n12268_0[2]),.dinb(w_asqrt29_12[0]),.dout(n12269),.clk(gclk));
	jor g11990(.dina(w_n12268_0[1]),.dinb(w_asqrt29_11[2]),.dout(n12270),.clk(gclk));
	jnot g11991(.din(w_n11773_0[0]),.dout(n12271),.clk(gclk));
	jnot g11992(.din(w_n11774_0[0]),.dout(n12272),.clk(gclk));
	jand g11993(.dina(w_asqrt16_26[2]),.dinb(w_n11770_0[0]),.dout(n12273),.clk(gclk));
	jand g11994(.dina(w_n12273_0[1]),.dinb(n12272),.dout(n12274),.clk(gclk));
	jor g11995(.dina(n12274),.dinb(n12271),.dout(n12275),.clk(gclk));
	jnot g11996(.din(w_n11775_0[0]),.dout(n12276),.clk(gclk));
	jand g11997(.dina(w_n12273_0[0]),.dinb(n12276),.dout(n12277),.clk(gclk));
	jnot g11998(.din(n12277),.dout(n12278),.clk(gclk));
	jand g11999(.dina(n12278),.dinb(n12275),.dout(n12279),.clk(gclk));
	jand g12000(.dina(w_n12279_0[1]),.dinb(n12270),.dout(n12280),.clk(gclk));
	jor g12001(.dina(w_n12280_0[1]),.dinb(w_n12269_0[1]),.dout(n12281),.clk(gclk));
	jand g12002(.dina(n12281),.dinb(w_asqrt30_15[1]),.dout(n12282),.clk(gclk));
	jor g12003(.dina(w_n12269_0[0]),.dinb(w_asqrt30_15[0]),.dout(n12283),.clk(gclk));
	jor g12004(.dina(n12283),.dinb(w_n12280_0[0]),.dout(n12284),.clk(gclk));
	jnot g12005(.din(w_n11781_0[0]),.dout(n12285),.clk(gclk));
	jnot g12006(.din(w_n11783_0[0]),.dout(n12286),.clk(gclk));
	jand g12007(.dina(w_asqrt16_26[1]),.dinb(w_n11777_0[0]),.dout(n12287),.clk(gclk));
	jand g12008(.dina(w_n12287_0[1]),.dinb(n12286),.dout(n12288),.clk(gclk));
	jor g12009(.dina(n12288),.dinb(n12285),.dout(n12289),.clk(gclk));
	jnot g12010(.din(w_n11784_0[0]),.dout(n12290),.clk(gclk));
	jand g12011(.dina(w_n12287_0[0]),.dinb(n12290),.dout(n12291),.clk(gclk));
	jnot g12012(.din(n12291),.dout(n12292),.clk(gclk));
	jand g12013(.dina(n12292),.dinb(n12289),.dout(n12293),.clk(gclk));
	jand g12014(.dina(w_n12293_0[1]),.dinb(w_n12284_0[1]),.dout(n12294),.clk(gclk));
	jor g12015(.dina(n12294),.dinb(w_n12282_0[1]),.dout(n12295),.clk(gclk));
	jand g12016(.dina(w_n12295_0[1]),.dinb(w_asqrt31_12[0]),.dout(n12296),.clk(gclk));
	jxor g12017(.dina(w_n11785_0[0]),.dinb(w_n6500_12[2]),.dout(n12297),.clk(gclk));
	jand g12018(.dina(n12297),.dinb(w_asqrt16_26[0]),.dout(n12298),.clk(gclk));
	jxor g12019(.dina(n12298),.dinb(w_n11795_0[0]),.dout(n12299),.clk(gclk));
	jnot g12020(.din(n12299),.dout(n12300),.clk(gclk));
	jor g12021(.dina(w_n12295_0[0]),.dinb(w_asqrt31_11[2]),.dout(n12301),.clk(gclk));
	jand g12022(.dina(w_n12301_0[1]),.dinb(w_n12300_0[1]),.dout(n12302),.clk(gclk));
	jor g12023(.dina(w_n12302_0[2]),.dinb(w_n12296_0[2]),.dout(n12303),.clk(gclk));
	jand g12024(.dina(n12303),.dinb(w_asqrt32_15[1]),.dout(n12304),.clk(gclk));
	jnot g12025(.din(w_n11800_0[0]),.dout(n12305),.clk(gclk));
	jand g12026(.dina(n12305),.dinb(w_n11798_0[0]),.dout(n12306),.clk(gclk));
	jand g12027(.dina(n12306),.dinb(w_asqrt16_25[2]),.dout(n12307),.clk(gclk));
	jxor g12028(.dina(n12307),.dinb(w_n11808_0[0]),.dout(n12308),.clk(gclk));
	jnot g12029(.din(n12308),.dout(n12309),.clk(gclk));
	jor g12030(.dina(w_n12296_0[1]),.dinb(w_asqrt32_15[0]),.dout(n12310),.clk(gclk));
	jor g12031(.dina(n12310),.dinb(w_n12302_0[1]),.dout(n12311),.clk(gclk));
	jand g12032(.dina(w_n12311_0[1]),.dinb(w_n12309_0[1]),.dout(n12312),.clk(gclk));
	jor g12033(.dina(w_n12312_0[1]),.dinb(w_n12304_0[1]),.dout(n12313),.clk(gclk));
	jand g12034(.dina(w_n12313_0[2]),.dinb(w_asqrt33_12[1]),.dout(n12314),.clk(gclk));
	jor g12035(.dina(w_n12313_0[1]),.dinb(w_asqrt33_12[0]),.dout(n12315),.clk(gclk));
	jnot g12036(.din(w_n11814_0[0]),.dout(n12316),.clk(gclk));
	jnot g12037(.din(w_n11815_0[0]),.dout(n12317),.clk(gclk));
	jand g12038(.dina(w_asqrt16_25[1]),.dinb(w_n11811_0[0]),.dout(n12318),.clk(gclk));
	jand g12039(.dina(w_n12318_0[1]),.dinb(n12317),.dout(n12319),.clk(gclk));
	jor g12040(.dina(n12319),.dinb(n12316),.dout(n12320),.clk(gclk));
	jnot g12041(.din(w_n11816_0[0]),.dout(n12321),.clk(gclk));
	jand g12042(.dina(w_n12318_0[0]),.dinb(n12321),.dout(n12322),.clk(gclk));
	jnot g12043(.din(n12322),.dout(n12323),.clk(gclk));
	jand g12044(.dina(n12323),.dinb(n12320),.dout(n12324),.clk(gclk));
	jand g12045(.dina(w_n12324_0[1]),.dinb(n12315),.dout(n12325),.clk(gclk));
	jor g12046(.dina(w_n12325_0[1]),.dinb(w_n12314_0[1]),.dout(n12326),.clk(gclk));
	jand g12047(.dina(n12326),.dinb(w_asqrt34_15[1]),.dout(n12327),.clk(gclk));
	jor g12048(.dina(w_n12314_0[0]),.dinb(w_asqrt34_15[0]),.dout(n12328),.clk(gclk));
	jor g12049(.dina(n12328),.dinb(w_n12325_0[0]),.dout(n12329),.clk(gclk));
	jnot g12050(.din(w_n11822_0[0]),.dout(n12330),.clk(gclk));
	jnot g12051(.din(w_n11824_0[0]),.dout(n12331),.clk(gclk));
	jand g12052(.dina(w_asqrt16_25[0]),.dinb(w_n11818_0[0]),.dout(n12332),.clk(gclk));
	jand g12053(.dina(w_n12332_0[1]),.dinb(n12331),.dout(n12333),.clk(gclk));
	jor g12054(.dina(n12333),.dinb(n12330),.dout(n12334),.clk(gclk));
	jnot g12055(.din(w_n11825_0[0]),.dout(n12335),.clk(gclk));
	jand g12056(.dina(w_n12332_0[0]),.dinb(n12335),.dout(n12336),.clk(gclk));
	jnot g12057(.din(n12336),.dout(n12337),.clk(gclk));
	jand g12058(.dina(n12337),.dinb(n12334),.dout(n12338),.clk(gclk));
	jand g12059(.dina(w_n12338_0[1]),.dinb(w_n12329_0[1]),.dout(n12339),.clk(gclk));
	jor g12060(.dina(n12339),.dinb(w_n12327_0[1]),.dout(n12340),.clk(gclk));
	jand g12061(.dina(w_n12340_0[1]),.dinb(w_asqrt35_12[1]),.dout(n12341),.clk(gclk));
	jxor g12062(.dina(w_n11826_0[0]),.dinb(w_n5116_13[1]),.dout(n12342),.clk(gclk));
	jand g12063(.dina(n12342),.dinb(w_asqrt16_24[2]),.dout(n12343),.clk(gclk));
	jxor g12064(.dina(n12343),.dinb(w_n11836_0[0]),.dout(n12344),.clk(gclk));
	jnot g12065(.din(n12344),.dout(n12345),.clk(gclk));
	jor g12066(.dina(w_n12340_0[0]),.dinb(w_asqrt35_12[0]),.dout(n12346),.clk(gclk));
	jand g12067(.dina(w_n12346_0[1]),.dinb(w_n12345_0[1]),.dout(n12347),.clk(gclk));
	jor g12068(.dina(w_n12347_0[2]),.dinb(w_n12341_0[2]),.dout(n12348),.clk(gclk));
	jand g12069(.dina(n12348),.dinb(w_asqrt36_15[1]),.dout(n12349),.clk(gclk));
	jnot g12070(.din(w_n11841_0[0]),.dout(n12350),.clk(gclk));
	jand g12071(.dina(n12350),.dinb(w_n11839_0[0]),.dout(n12351),.clk(gclk));
	jand g12072(.dina(n12351),.dinb(w_asqrt16_24[1]),.dout(n12352),.clk(gclk));
	jxor g12073(.dina(n12352),.dinb(w_n11849_0[0]),.dout(n12353),.clk(gclk));
	jnot g12074(.din(n12353),.dout(n12354),.clk(gclk));
	jor g12075(.dina(w_n12341_0[1]),.dinb(w_asqrt36_15[0]),.dout(n12355),.clk(gclk));
	jor g12076(.dina(n12355),.dinb(w_n12347_0[1]),.dout(n12356),.clk(gclk));
	jand g12077(.dina(w_n12356_0[1]),.dinb(w_n12354_0[1]),.dout(n12357),.clk(gclk));
	jor g12078(.dina(w_n12357_0[1]),.dinb(w_n12349_0[1]),.dout(n12358),.clk(gclk));
	jand g12079(.dina(w_n12358_0[2]),.dinb(w_asqrt37_12[2]),.dout(n12359),.clk(gclk));
	jor g12080(.dina(w_n12358_0[1]),.dinb(w_asqrt37_12[1]),.dout(n12360),.clk(gclk));
	jnot g12081(.din(w_n11855_0[0]),.dout(n12361),.clk(gclk));
	jnot g12082(.din(w_n11856_0[0]),.dout(n12362),.clk(gclk));
	jand g12083(.dina(w_asqrt16_24[0]),.dinb(w_n11852_0[0]),.dout(n12363),.clk(gclk));
	jand g12084(.dina(w_n12363_0[1]),.dinb(n12362),.dout(n12364),.clk(gclk));
	jor g12085(.dina(n12364),.dinb(n12361),.dout(n12365),.clk(gclk));
	jnot g12086(.din(w_n11857_0[0]),.dout(n12366),.clk(gclk));
	jand g12087(.dina(w_n12363_0[0]),.dinb(n12366),.dout(n12367),.clk(gclk));
	jnot g12088(.din(n12367),.dout(n12368),.clk(gclk));
	jand g12089(.dina(n12368),.dinb(n12365),.dout(n12369),.clk(gclk));
	jand g12090(.dina(w_n12369_0[1]),.dinb(n12360),.dout(n12370),.clk(gclk));
	jor g12091(.dina(w_n12370_0[1]),.dinb(w_n12359_0[1]),.dout(n12371),.clk(gclk));
	jand g12092(.dina(n12371),.dinb(w_asqrt38_15[1]),.dout(n12372),.clk(gclk));
	jor g12093(.dina(w_n12359_0[0]),.dinb(w_asqrt38_15[0]),.dout(n12373),.clk(gclk));
	jor g12094(.dina(n12373),.dinb(w_n12370_0[0]),.dout(n12374),.clk(gclk));
	jnot g12095(.din(w_n11863_0[0]),.dout(n12375),.clk(gclk));
	jnot g12096(.din(w_n11865_0[0]),.dout(n12376),.clk(gclk));
	jand g12097(.dina(w_asqrt16_23[2]),.dinb(w_n11859_0[0]),.dout(n12377),.clk(gclk));
	jand g12098(.dina(w_n12377_0[1]),.dinb(n12376),.dout(n12378),.clk(gclk));
	jor g12099(.dina(n12378),.dinb(n12375),.dout(n12379),.clk(gclk));
	jnot g12100(.din(w_n11866_0[0]),.dout(n12380),.clk(gclk));
	jand g12101(.dina(w_n12377_0[0]),.dinb(n12380),.dout(n12381),.clk(gclk));
	jnot g12102(.din(n12381),.dout(n12382),.clk(gclk));
	jand g12103(.dina(n12382),.dinb(n12379),.dout(n12383),.clk(gclk));
	jand g12104(.dina(w_n12383_0[1]),.dinb(w_n12374_0[1]),.dout(n12384),.clk(gclk));
	jor g12105(.dina(n12384),.dinb(w_n12372_0[1]),.dout(n12385),.clk(gclk));
	jand g12106(.dina(w_n12385_0[1]),.dinb(w_asqrt39_12[2]),.dout(n12386),.clk(gclk));
	jxor g12107(.dina(w_n11867_0[0]),.dinb(w_n3907_14[1]),.dout(n12387),.clk(gclk));
	jand g12108(.dina(n12387),.dinb(w_asqrt16_23[1]),.dout(n12388),.clk(gclk));
	jxor g12109(.dina(n12388),.dinb(w_n11877_0[0]),.dout(n12389),.clk(gclk));
	jnot g12110(.din(n12389),.dout(n12390),.clk(gclk));
	jor g12111(.dina(w_n12385_0[0]),.dinb(w_asqrt39_12[1]),.dout(n12391),.clk(gclk));
	jand g12112(.dina(w_n12391_0[1]),.dinb(w_n12390_0[1]),.dout(n12392),.clk(gclk));
	jor g12113(.dina(w_n12392_0[2]),.dinb(w_n12386_0[2]),.dout(n12393),.clk(gclk));
	jand g12114(.dina(n12393),.dinb(w_asqrt40_15[1]),.dout(n12394),.clk(gclk));
	jnot g12115(.din(w_n11882_0[0]),.dout(n12395),.clk(gclk));
	jand g12116(.dina(n12395),.dinb(w_n11880_0[0]),.dout(n12396),.clk(gclk));
	jand g12117(.dina(n12396),.dinb(w_asqrt16_23[0]),.dout(n12397),.clk(gclk));
	jxor g12118(.dina(n12397),.dinb(w_n11890_0[0]),.dout(n12398),.clk(gclk));
	jnot g12119(.din(n12398),.dout(n12399),.clk(gclk));
	jor g12120(.dina(w_n12386_0[1]),.dinb(w_asqrt40_15[0]),.dout(n12400),.clk(gclk));
	jor g12121(.dina(n12400),.dinb(w_n12392_0[1]),.dout(n12401),.clk(gclk));
	jand g12122(.dina(w_n12401_0[1]),.dinb(w_n12399_0[1]),.dout(n12402),.clk(gclk));
	jor g12123(.dina(w_n12402_0[1]),.dinb(w_n12394_0[1]),.dout(n12403),.clk(gclk));
	jand g12124(.dina(w_n12403_0[2]),.dinb(w_asqrt41_13[0]),.dout(n12404),.clk(gclk));
	jor g12125(.dina(w_n12403_0[1]),.dinb(w_asqrt41_12[2]),.dout(n12405),.clk(gclk));
	jnot g12126(.din(w_n11896_0[0]),.dout(n12406),.clk(gclk));
	jnot g12127(.din(w_n11897_0[0]),.dout(n12407),.clk(gclk));
	jand g12128(.dina(w_asqrt16_22[2]),.dinb(w_n11893_0[0]),.dout(n12408),.clk(gclk));
	jand g12129(.dina(w_n12408_0[1]),.dinb(n12407),.dout(n12409),.clk(gclk));
	jor g12130(.dina(n12409),.dinb(n12406),.dout(n12410),.clk(gclk));
	jnot g12131(.din(w_n11898_0[0]),.dout(n12411),.clk(gclk));
	jand g12132(.dina(w_n12408_0[0]),.dinb(n12411),.dout(n12412),.clk(gclk));
	jnot g12133(.din(n12412),.dout(n12413),.clk(gclk));
	jand g12134(.dina(n12413),.dinb(n12410),.dout(n12414),.clk(gclk));
	jand g12135(.dina(w_n12414_0[1]),.dinb(n12405),.dout(n12415),.clk(gclk));
	jor g12136(.dina(w_n12415_0[1]),.dinb(w_n12404_0[1]),.dout(n12416),.clk(gclk));
	jand g12137(.dina(n12416),.dinb(w_asqrt42_15[1]),.dout(n12417),.clk(gclk));
	jor g12138(.dina(w_n12404_0[0]),.dinb(w_asqrt42_15[0]),.dout(n12418),.clk(gclk));
	jor g12139(.dina(n12418),.dinb(w_n12415_0[0]),.dout(n12419),.clk(gclk));
	jnot g12140(.din(w_n11904_0[0]),.dout(n12420),.clk(gclk));
	jnot g12141(.din(w_n11906_0[0]),.dout(n12421),.clk(gclk));
	jand g12142(.dina(w_asqrt16_22[1]),.dinb(w_n11900_0[0]),.dout(n12422),.clk(gclk));
	jand g12143(.dina(w_n12422_0[1]),.dinb(n12421),.dout(n12423),.clk(gclk));
	jor g12144(.dina(n12423),.dinb(n12420),.dout(n12424),.clk(gclk));
	jnot g12145(.din(w_n11907_0[0]),.dout(n12425),.clk(gclk));
	jand g12146(.dina(w_n12422_0[0]),.dinb(n12425),.dout(n12426),.clk(gclk));
	jnot g12147(.din(n12426),.dout(n12427),.clk(gclk));
	jand g12148(.dina(n12427),.dinb(n12424),.dout(n12428),.clk(gclk));
	jand g12149(.dina(w_n12428_0[1]),.dinb(w_n12419_0[1]),.dout(n12429),.clk(gclk));
	jor g12150(.dina(n12429),.dinb(w_n12417_0[1]),.dout(n12430),.clk(gclk));
	jand g12151(.dina(w_n12430_0[1]),.dinb(w_asqrt43_13[0]),.dout(n12431),.clk(gclk));
	jxor g12152(.dina(w_n11908_0[0]),.dinb(w_n2870_15[0]),.dout(n12432),.clk(gclk));
	jand g12153(.dina(n12432),.dinb(w_asqrt16_22[0]),.dout(n12433),.clk(gclk));
	jxor g12154(.dina(n12433),.dinb(w_n11918_0[0]),.dout(n12434),.clk(gclk));
	jnot g12155(.din(n12434),.dout(n12435),.clk(gclk));
	jor g12156(.dina(w_n12430_0[0]),.dinb(w_asqrt43_12[2]),.dout(n12436),.clk(gclk));
	jand g12157(.dina(w_n12436_0[1]),.dinb(w_n12435_0[1]),.dout(n12437),.clk(gclk));
	jor g12158(.dina(w_n12437_0[2]),.dinb(w_n12431_0[2]),.dout(n12438),.clk(gclk));
	jand g12159(.dina(n12438),.dinb(w_asqrt44_15[1]),.dout(n12439),.clk(gclk));
	jnot g12160(.din(w_n11923_0[0]),.dout(n12440),.clk(gclk));
	jand g12161(.dina(n12440),.dinb(w_n11921_0[0]),.dout(n12441),.clk(gclk));
	jand g12162(.dina(n12441),.dinb(w_asqrt16_21[2]),.dout(n12442),.clk(gclk));
	jxor g12163(.dina(n12442),.dinb(w_n11931_0[0]),.dout(n12443),.clk(gclk));
	jnot g12164(.din(n12443),.dout(n12444),.clk(gclk));
	jor g12165(.dina(w_n12431_0[1]),.dinb(w_asqrt44_15[0]),.dout(n12445),.clk(gclk));
	jor g12166(.dina(n12445),.dinb(w_n12437_0[1]),.dout(n12446),.clk(gclk));
	jand g12167(.dina(w_n12446_0[1]),.dinb(w_n12444_0[1]),.dout(n12447),.clk(gclk));
	jor g12168(.dina(w_n12447_0[1]),.dinb(w_n12439_0[1]),.dout(n12448),.clk(gclk));
	jand g12169(.dina(w_n12448_0[2]),.dinb(w_asqrt45_13[1]),.dout(n12449),.clk(gclk));
	jor g12170(.dina(w_n12448_0[1]),.dinb(w_asqrt45_13[0]),.dout(n12450),.clk(gclk));
	jnot g12171(.din(w_n11937_0[0]),.dout(n12451),.clk(gclk));
	jnot g12172(.din(w_n11938_0[0]),.dout(n12452),.clk(gclk));
	jand g12173(.dina(w_asqrt16_21[1]),.dinb(w_n11934_0[0]),.dout(n12453),.clk(gclk));
	jand g12174(.dina(w_n12453_0[1]),.dinb(n12452),.dout(n12454),.clk(gclk));
	jor g12175(.dina(n12454),.dinb(n12451),.dout(n12455),.clk(gclk));
	jnot g12176(.din(w_n11939_0[0]),.dout(n12456),.clk(gclk));
	jand g12177(.dina(w_n12453_0[0]),.dinb(n12456),.dout(n12457),.clk(gclk));
	jnot g12178(.din(n12457),.dout(n12458),.clk(gclk));
	jand g12179(.dina(n12458),.dinb(n12455),.dout(n12459),.clk(gclk));
	jand g12180(.dina(w_n12459_0[1]),.dinb(n12450),.dout(n12460),.clk(gclk));
	jor g12181(.dina(w_n12460_0[1]),.dinb(w_n12449_0[1]),.dout(n12461),.clk(gclk));
	jand g12182(.dina(n12461),.dinb(w_asqrt46_15[1]),.dout(n12462),.clk(gclk));
	jnot g12183(.din(w_n11943_0[0]),.dout(n12463),.clk(gclk));
	jand g12184(.dina(n12463),.dinb(w_n11941_0[0]),.dout(n12464),.clk(gclk));
	jand g12185(.dina(n12464),.dinb(w_asqrt16_21[0]),.dout(n12465),.clk(gclk));
	jxor g12186(.dina(n12465),.dinb(w_n11951_0[0]),.dout(n12466),.clk(gclk));
	jnot g12187(.din(n12466),.dout(n12467),.clk(gclk));
	jor g12188(.dina(w_n12449_0[0]),.dinb(w_asqrt46_15[0]),.dout(n12468),.clk(gclk));
	jor g12189(.dina(n12468),.dinb(w_n12460_0[0]),.dout(n12469),.clk(gclk));
	jand g12190(.dina(w_n12469_0[1]),.dinb(w_n12467_0[1]),.dout(n12470),.clk(gclk));
	jor g12191(.dina(w_n12470_0[1]),.dinb(w_n12462_0[1]),.dout(n12471),.clk(gclk));
	jand g12192(.dina(w_n12471_0[2]),.dinb(w_asqrt47_13[1]),.dout(n12472),.clk(gclk));
	jor g12193(.dina(w_n12471_0[1]),.dinb(w_asqrt47_13[0]),.dout(n12473),.clk(gclk));
	jand g12194(.dina(n12473),.dinb(w_n12145_0[0]),.dout(n12474),.clk(gclk));
	jor g12195(.dina(w_n12474_0[1]),.dinb(w_n12472_0[1]),.dout(n12475),.clk(gclk));
	jand g12196(.dina(n12475),.dinb(w_asqrt48_15[1]),.dout(n12476),.clk(gclk));
	jor g12197(.dina(w_n12472_0[0]),.dinb(w_asqrt48_15[0]),.dout(n12477),.clk(gclk));
	jor g12198(.dina(n12477),.dinb(w_n12474_0[0]),.dout(n12478),.clk(gclk));
	jnot g12199(.din(w_n11963_0[0]),.dout(n12479),.clk(gclk));
	jnot g12200(.din(w_n11965_0[0]),.dout(n12480),.clk(gclk));
	jand g12201(.dina(w_asqrt16_20[2]),.dinb(w_n11959_0[0]),.dout(n12481),.clk(gclk));
	jand g12202(.dina(w_n12481_0[1]),.dinb(n12480),.dout(n12482),.clk(gclk));
	jor g12203(.dina(n12482),.dinb(n12479),.dout(n12483),.clk(gclk));
	jnot g12204(.din(w_n11966_0[0]),.dout(n12484),.clk(gclk));
	jand g12205(.dina(w_n12481_0[0]),.dinb(n12484),.dout(n12485),.clk(gclk));
	jnot g12206(.din(n12485),.dout(n12486),.clk(gclk));
	jand g12207(.dina(n12486),.dinb(n12483),.dout(n12487),.clk(gclk));
	jand g12208(.dina(w_n12487_0[1]),.dinb(w_n12478_0[1]),.dout(n12488),.clk(gclk));
	jor g12209(.dina(n12488),.dinb(w_n12476_0[1]),.dout(n12489),.clk(gclk));
	jand g12210(.dina(w_n12489_0[2]),.dinb(w_asqrt49_13[2]),.dout(n12490),.clk(gclk));
	jor g12211(.dina(w_n12489_0[1]),.dinb(w_asqrt49_13[1]),.dout(n12491),.clk(gclk));
	jnot g12212(.din(w_n11971_0[0]),.dout(n12492),.clk(gclk));
	jnot g12213(.din(w_n11972_0[0]),.dout(n12493),.clk(gclk));
	jand g12214(.dina(w_asqrt16_20[1]),.dinb(w_n11968_0[0]),.dout(n12494),.clk(gclk));
	jand g12215(.dina(w_n12494_0[1]),.dinb(n12493),.dout(n12495),.clk(gclk));
	jor g12216(.dina(n12495),.dinb(n12492),.dout(n12496),.clk(gclk));
	jnot g12217(.din(w_n11973_0[0]),.dout(n12497),.clk(gclk));
	jand g12218(.dina(w_n12494_0[0]),.dinb(n12497),.dout(n12498),.clk(gclk));
	jnot g12219(.din(n12498),.dout(n12499),.clk(gclk));
	jand g12220(.dina(n12499),.dinb(n12496),.dout(n12500),.clk(gclk));
	jand g12221(.dina(w_n12500_0[1]),.dinb(n12491),.dout(n12501),.clk(gclk));
	jor g12222(.dina(w_n12501_0[1]),.dinb(w_n12490_0[1]),.dout(n12502),.clk(gclk));
	jand g12223(.dina(n12502),.dinb(w_asqrt50_15[1]),.dout(n12503),.clk(gclk));
	jor g12224(.dina(w_n12490_0[0]),.dinb(w_asqrt50_15[0]),.dout(n12504),.clk(gclk));
	jor g12225(.dina(n12504),.dinb(w_n12501_0[0]),.dout(n12505),.clk(gclk));
	jnot g12226(.din(w_n11979_0[0]),.dout(n12506),.clk(gclk));
	jnot g12227(.din(w_n11981_0[0]),.dout(n12507),.clk(gclk));
	jand g12228(.dina(w_asqrt16_20[0]),.dinb(w_n11975_0[0]),.dout(n12508),.clk(gclk));
	jand g12229(.dina(w_n12508_0[1]),.dinb(n12507),.dout(n12509),.clk(gclk));
	jor g12230(.dina(n12509),.dinb(n12506),.dout(n12510),.clk(gclk));
	jnot g12231(.din(w_n11982_0[0]),.dout(n12511),.clk(gclk));
	jand g12232(.dina(w_n12508_0[0]),.dinb(n12511),.dout(n12512),.clk(gclk));
	jnot g12233(.din(n12512),.dout(n12513),.clk(gclk));
	jand g12234(.dina(n12513),.dinb(n12510),.dout(n12514),.clk(gclk));
	jand g12235(.dina(w_n12514_0[1]),.dinb(w_n12505_0[1]),.dout(n12515),.clk(gclk));
	jor g12236(.dina(n12515),.dinb(w_n12503_0[1]),.dout(n12516),.clk(gclk));
	jand g12237(.dina(w_n12516_0[1]),.dinb(w_asqrt51_13[2]),.dout(n12517),.clk(gclk));
	jxor g12238(.dina(w_n11983_0[0]),.dinb(w_n1312_16[2]),.dout(n12518),.clk(gclk));
	jand g12239(.dina(n12518),.dinb(w_asqrt16_19[2]),.dout(n12519),.clk(gclk));
	jxor g12240(.dina(n12519),.dinb(w_n11993_0[0]),.dout(n12520),.clk(gclk));
	jnot g12241(.din(n12520),.dout(n12521),.clk(gclk));
	jor g12242(.dina(w_n12516_0[0]),.dinb(w_asqrt51_13[1]),.dout(n12522),.clk(gclk));
	jand g12243(.dina(w_n12522_0[1]),.dinb(w_n12521_0[1]),.dout(n12523),.clk(gclk));
	jor g12244(.dina(w_n12523_0[2]),.dinb(w_n12517_0[2]),.dout(n12524),.clk(gclk));
	jand g12245(.dina(n12524),.dinb(w_asqrt52_15[1]),.dout(n12525),.clk(gclk));
	jnot g12246(.din(w_n11998_0[0]),.dout(n12526),.clk(gclk));
	jand g12247(.dina(n12526),.dinb(w_n11996_0[0]),.dout(n12527),.clk(gclk));
	jand g12248(.dina(n12527),.dinb(w_asqrt16_19[1]),.dout(n12528),.clk(gclk));
	jxor g12249(.dina(n12528),.dinb(w_n12006_0[0]),.dout(n12529),.clk(gclk));
	jnot g12250(.din(n12529),.dout(n12530),.clk(gclk));
	jor g12251(.dina(w_n12517_0[1]),.dinb(w_asqrt52_15[0]),.dout(n12531),.clk(gclk));
	jor g12252(.dina(n12531),.dinb(w_n12523_0[1]),.dout(n12532),.clk(gclk));
	jand g12253(.dina(w_n12532_0[1]),.dinb(w_n12530_0[1]),.dout(n12533),.clk(gclk));
	jor g12254(.dina(w_n12533_0[1]),.dinb(w_n12525_0[1]),.dout(n12534),.clk(gclk));
	jand g12255(.dina(w_n12534_0[2]),.dinb(w_asqrt53_14[0]),.dout(n12535),.clk(gclk));
	jor g12256(.dina(w_n12534_0[1]),.dinb(w_asqrt53_13[2]),.dout(n12536),.clk(gclk));
	jnot g12257(.din(w_n12012_0[0]),.dout(n12537),.clk(gclk));
	jnot g12258(.din(w_n12013_0[0]),.dout(n12538),.clk(gclk));
	jand g12259(.dina(w_asqrt16_19[0]),.dinb(w_n12009_0[0]),.dout(n12539),.clk(gclk));
	jand g12260(.dina(w_n12539_0[1]),.dinb(n12538),.dout(n12540),.clk(gclk));
	jor g12261(.dina(n12540),.dinb(n12537),.dout(n12541),.clk(gclk));
	jnot g12262(.din(w_n12014_0[0]),.dout(n12542),.clk(gclk));
	jand g12263(.dina(w_n12539_0[0]),.dinb(n12542),.dout(n12543),.clk(gclk));
	jnot g12264(.din(n12543),.dout(n12544),.clk(gclk));
	jand g12265(.dina(n12544),.dinb(n12541),.dout(n12545),.clk(gclk));
	jand g12266(.dina(w_n12545_0[1]),.dinb(n12536),.dout(n12546),.clk(gclk));
	jor g12267(.dina(w_n12546_0[1]),.dinb(w_n12535_0[1]),.dout(n12547),.clk(gclk));
	jand g12268(.dina(n12547),.dinb(w_asqrt54_15[1]),.dout(n12548),.clk(gclk));
	jor g12269(.dina(w_n12535_0[0]),.dinb(w_asqrt54_15[0]),.dout(n12549),.clk(gclk));
	jor g12270(.dina(n12549),.dinb(w_n12546_0[0]),.dout(n12550),.clk(gclk));
	jnot g12271(.din(w_n12020_0[0]),.dout(n12551),.clk(gclk));
	jnot g12272(.din(w_n12022_0[0]),.dout(n12552),.clk(gclk));
	jand g12273(.dina(w_asqrt16_18[2]),.dinb(w_n12016_0[0]),.dout(n12553),.clk(gclk));
	jand g12274(.dina(w_n12553_0[1]),.dinb(n12552),.dout(n12554),.clk(gclk));
	jor g12275(.dina(n12554),.dinb(n12551),.dout(n12555),.clk(gclk));
	jnot g12276(.din(w_n12023_0[0]),.dout(n12556),.clk(gclk));
	jand g12277(.dina(w_n12553_0[0]),.dinb(n12556),.dout(n12557),.clk(gclk));
	jnot g12278(.din(n12557),.dout(n12558),.clk(gclk));
	jand g12279(.dina(n12558),.dinb(n12555),.dout(n12559),.clk(gclk));
	jand g12280(.dina(w_n12559_0[1]),.dinb(w_n12550_0[1]),.dout(n12560),.clk(gclk));
	jor g12281(.dina(n12560),.dinb(w_n12548_0[1]),.dout(n12561),.clk(gclk));
	jand g12282(.dina(w_n12561_0[1]),.dinb(w_asqrt55_14[1]),.dout(n12562),.clk(gclk));
	jxor g12283(.dina(w_n12024_0[0]),.dinb(w_n791_17[2]),.dout(n12563),.clk(gclk));
	jand g12284(.dina(n12563),.dinb(w_asqrt16_18[1]),.dout(n12564),.clk(gclk));
	jxor g12285(.dina(n12564),.dinb(w_n12034_0[0]),.dout(n12565),.clk(gclk));
	jnot g12286(.din(n12565),.dout(n12566),.clk(gclk));
	jor g12287(.dina(w_n12561_0[0]),.dinb(w_asqrt55_14[0]),.dout(n12567),.clk(gclk));
	jand g12288(.dina(w_n12567_0[1]),.dinb(w_n12566_0[1]),.dout(n12568),.clk(gclk));
	jor g12289(.dina(w_n12568_0[2]),.dinb(w_n12562_0[2]),.dout(n12569),.clk(gclk));
	jand g12290(.dina(n12569),.dinb(w_asqrt56_15[1]),.dout(n12570),.clk(gclk));
	jnot g12291(.din(w_n12039_0[0]),.dout(n12571),.clk(gclk));
	jand g12292(.dina(n12571),.dinb(w_n12037_0[0]),.dout(n12572),.clk(gclk));
	jand g12293(.dina(n12572),.dinb(w_asqrt16_18[0]),.dout(n12573),.clk(gclk));
	jxor g12294(.dina(n12573),.dinb(w_n12047_0[0]),.dout(n12574),.clk(gclk));
	jnot g12295(.din(n12574),.dout(n12575),.clk(gclk));
	jor g12296(.dina(w_n12562_0[1]),.dinb(w_asqrt56_15[0]),.dout(n12576),.clk(gclk));
	jor g12297(.dina(n12576),.dinb(w_n12568_0[1]),.dout(n12577),.clk(gclk));
	jand g12298(.dina(w_n12577_0[1]),.dinb(w_n12575_0[1]),.dout(n12578),.clk(gclk));
	jor g12299(.dina(w_n12578_0[1]),.dinb(w_n12570_0[1]),.dout(n12579),.clk(gclk));
	jand g12300(.dina(w_n12579_0[2]),.dinb(w_asqrt57_14[2]),.dout(n12580),.clk(gclk));
	jor g12301(.dina(w_n12579_0[1]),.dinb(w_asqrt57_14[1]),.dout(n12581),.clk(gclk));
	jnot g12302(.din(w_n12053_0[0]),.dout(n12582),.clk(gclk));
	jnot g12303(.din(w_n12054_0[0]),.dout(n12583),.clk(gclk));
	jand g12304(.dina(w_asqrt16_17[2]),.dinb(w_n12050_0[0]),.dout(n12584),.clk(gclk));
	jand g12305(.dina(w_n12584_0[1]),.dinb(n12583),.dout(n12585),.clk(gclk));
	jor g12306(.dina(n12585),.dinb(n12582),.dout(n12586),.clk(gclk));
	jnot g12307(.din(w_n12055_0[0]),.dout(n12587),.clk(gclk));
	jand g12308(.dina(w_n12584_0[0]),.dinb(n12587),.dout(n12588),.clk(gclk));
	jnot g12309(.din(n12588),.dout(n12589),.clk(gclk));
	jand g12310(.dina(n12589),.dinb(n12586),.dout(n12590),.clk(gclk));
	jand g12311(.dina(w_n12590_0[1]),.dinb(n12581),.dout(n12591),.clk(gclk));
	jor g12312(.dina(w_n12591_0[1]),.dinb(w_n12580_0[1]),.dout(n12592),.clk(gclk));
	jand g12313(.dina(n12592),.dinb(w_asqrt58_15[1]),.dout(n12593),.clk(gclk));
	jor g12314(.dina(w_n12580_0[0]),.dinb(w_asqrt58_15[0]),.dout(n12594),.clk(gclk));
	jor g12315(.dina(n12594),.dinb(w_n12591_0[0]),.dout(n12595),.clk(gclk));
	jnot g12316(.din(w_n12061_0[0]),.dout(n12596),.clk(gclk));
	jnot g12317(.din(w_n12063_0[0]),.dout(n12597),.clk(gclk));
	jand g12318(.dina(w_asqrt16_17[1]),.dinb(w_n12057_0[0]),.dout(n12598),.clk(gclk));
	jand g12319(.dina(w_n12598_0[1]),.dinb(n12597),.dout(n12599),.clk(gclk));
	jor g12320(.dina(n12599),.dinb(n12596),.dout(n12600),.clk(gclk));
	jnot g12321(.din(w_n12064_0[0]),.dout(n12601),.clk(gclk));
	jand g12322(.dina(w_n12598_0[0]),.dinb(n12601),.dout(n12602),.clk(gclk));
	jnot g12323(.din(n12602),.dout(n12603),.clk(gclk));
	jand g12324(.dina(n12603),.dinb(n12600),.dout(n12604),.clk(gclk));
	jand g12325(.dina(w_n12604_0[1]),.dinb(w_n12595_0[1]),.dout(n12605),.clk(gclk));
	jor g12326(.dina(n12605),.dinb(w_n12593_0[1]),.dout(n12606),.clk(gclk));
	jand g12327(.dina(w_n12606_0[1]),.dinb(w_asqrt59_15[0]),.dout(n12607),.clk(gclk));
	jxor g12328(.dina(w_n12065_0[0]),.dinb(w_n425_18[1]),.dout(n12608),.clk(gclk));
	jand g12329(.dina(n12608),.dinb(w_asqrt16_17[0]),.dout(n12609),.clk(gclk));
	jxor g12330(.dina(n12609),.dinb(w_n12075_0[0]),.dout(n12610),.clk(gclk));
	jnot g12331(.din(n12610),.dout(n12611),.clk(gclk));
	jor g12332(.dina(w_n12606_0[0]),.dinb(w_asqrt59_14[2]),.dout(n12612),.clk(gclk));
	jand g12333(.dina(w_n12612_0[1]),.dinb(w_n12611_0[1]),.dout(n12613),.clk(gclk));
	jor g12334(.dina(w_n12613_0[2]),.dinb(w_n12607_0[2]),.dout(n12614),.clk(gclk));
	jand g12335(.dina(n12614),.dinb(w_asqrt60_15[0]),.dout(n12615),.clk(gclk));
	jnot g12336(.din(w_n12080_0[0]),.dout(n12616),.clk(gclk));
	jand g12337(.dina(n12616),.dinb(w_n12078_0[0]),.dout(n12617),.clk(gclk));
	jand g12338(.dina(n12617),.dinb(w_asqrt16_16[2]),.dout(n12618),.clk(gclk));
	jxor g12339(.dina(n12618),.dinb(w_n12088_0[0]),.dout(n12619),.clk(gclk));
	jnot g12340(.din(n12619),.dout(n12620),.clk(gclk));
	jor g12341(.dina(w_n12607_0[1]),.dinb(w_asqrt60_14[2]),.dout(n12621),.clk(gclk));
	jor g12342(.dina(n12621),.dinb(w_n12613_0[1]),.dout(n12622),.clk(gclk));
	jand g12343(.dina(w_n12622_0[1]),.dinb(w_n12620_0[1]),.dout(n12623),.clk(gclk));
	jor g12344(.dina(w_n12623_0[1]),.dinb(w_n12615_0[1]),.dout(n12624),.clk(gclk));
	jand g12345(.dina(w_n12624_0[2]),.dinb(w_asqrt61_15[1]),.dout(n12625),.clk(gclk));
	jor g12346(.dina(w_n12624_0[1]),.dinb(w_asqrt61_15[0]),.dout(n12626),.clk(gclk));
	jnot g12347(.din(w_n12094_0[0]),.dout(n12627),.clk(gclk));
	jnot g12348(.din(w_n12095_0[0]),.dout(n12628),.clk(gclk));
	jand g12349(.dina(w_asqrt16_16[1]),.dinb(w_n12091_0[0]),.dout(n12629),.clk(gclk));
	jand g12350(.dina(w_n12629_0[1]),.dinb(n12628),.dout(n12630),.clk(gclk));
	jor g12351(.dina(n12630),.dinb(n12627),.dout(n12631),.clk(gclk));
	jnot g12352(.din(w_n12096_0[0]),.dout(n12632),.clk(gclk));
	jand g12353(.dina(w_n12629_0[0]),.dinb(n12632),.dout(n12633),.clk(gclk));
	jnot g12354(.din(n12633),.dout(n12634),.clk(gclk));
	jand g12355(.dina(n12634),.dinb(n12631),.dout(n12635),.clk(gclk));
	jand g12356(.dina(w_n12635_0[1]),.dinb(n12626),.dout(n12636),.clk(gclk));
	jor g12357(.dina(w_n12636_0[1]),.dinb(w_n12625_0[1]),.dout(n12637),.clk(gclk));
	jand g12358(.dina(n12637),.dinb(w_asqrt62_15[1]),.dout(n12638),.clk(gclk));
	jor g12359(.dina(w_n12625_0[0]),.dinb(w_asqrt62_15[0]),.dout(n12639),.clk(gclk));
	jor g12360(.dina(n12639),.dinb(w_n12636_0[0]),.dout(n12640),.clk(gclk));
	jnot g12361(.din(w_n12102_0[0]),.dout(n12641),.clk(gclk));
	jnot g12362(.din(w_n12104_0[0]),.dout(n12642),.clk(gclk));
	jand g12363(.dina(w_asqrt16_16[0]),.dinb(w_n12098_0[0]),.dout(n12643),.clk(gclk));
	jand g12364(.dina(w_n12643_0[1]),.dinb(n12642),.dout(n12644),.clk(gclk));
	jor g12365(.dina(n12644),.dinb(n12641),.dout(n12645),.clk(gclk));
	jnot g12366(.din(w_n12105_0[0]),.dout(n12646),.clk(gclk));
	jand g12367(.dina(w_n12643_0[0]),.dinb(n12646),.dout(n12647),.clk(gclk));
	jnot g12368(.din(n12647),.dout(n12648),.clk(gclk));
	jand g12369(.dina(n12648),.dinb(n12645),.dout(n12649),.clk(gclk));
	jand g12370(.dina(w_n12649_0[1]),.dinb(w_n12640_0[1]),.dout(n12650),.clk(gclk));
	jor g12371(.dina(n12650),.dinb(w_n12638_0[1]),.dout(n12651),.clk(gclk));
	jxor g12372(.dina(w_n12106_0[0]),.dinb(w_n199_22[2]),.dout(n12652),.clk(gclk));
	jand g12373(.dina(n12652),.dinb(w_asqrt16_15[2]),.dout(n12653),.clk(gclk));
	jxor g12374(.dina(n12653),.dinb(w_n12116_0[0]),.dout(n12654),.clk(gclk));
	jnot g12375(.din(w_n12118_0[0]),.dout(n12655),.clk(gclk));
	jand g12376(.dina(w_asqrt16_15[1]),.dinb(w_n12125_0[1]),.dout(n12656),.clk(gclk));
	jand g12377(.dina(w_n12656_0[1]),.dinb(w_n12655_0[2]),.dout(n12657),.clk(gclk));
	jor g12378(.dina(n12657),.dinb(w_n12133_0[0]),.dout(n12658),.clk(gclk));
	jor g12379(.dina(n12658),.dinb(w_n12654_0[1]),.dout(n12659),.clk(gclk));
	jnot g12380(.din(n12659),.dout(n12660),.clk(gclk));
	jand g12381(.dina(n12660),.dinb(w_n12651_1[2]),.dout(n12661),.clk(gclk));
	jor g12382(.dina(n12661),.dinb(w_asqrt63_8[1]),.dout(n12662),.clk(gclk));
	jnot g12383(.din(w_n12654_0[0]),.dout(n12663),.clk(gclk));
	jor g12384(.dina(w_n12663_0[2]),.dinb(w_n12651_1[1]),.dout(n12664),.clk(gclk));
	jor g12385(.dina(w_n12656_0[0]),.dinb(w_n12655_0[1]),.dout(n12665),.clk(gclk));
	jand g12386(.dina(w_n12125_0[0]),.dinb(w_n12655_0[0]),.dout(n12666),.clk(gclk));
	jor g12387(.dina(n12666),.dinb(w_n194_21[2]),.dout(n12667),.clk(gclk));
	jnot g12388(.din(n12667),.dout(n12668),.clk(gclk));
	jand g12389(.dina(n12668),.dinb(n12665),.dout(n12669),.clk(gclk));
	jnot g12390(.din(w_asqrt16_15[0]),.dout(n12670),.clk(gclk));
	jnot g12391(.din(w_n12669_0[1]),.dout(n12673),.clk(gclk));
	jand g12392(.dina(n12673),.dinb(w_n12664_0[1]),.dout(n12674),.clk(gclk));
	jand g12393(.dina(n12674),.dinb(w_n12662_0[1]),.dout(n12675),.clk(gclk));
	jxor g12394(.dina(w_n12471_0[0]),.dinb(w_n1646_18[2]),.dout(n12676),.clk(gclk));
	jor g12395(.dina(n12676),.dinb(w_n12675_24[1]),.dout(n12677),.clk(gclk));
	jxor g12396(.dina(n12677),.dinb(n12146),.dout(n12678),.clk(gclk));
	jnot g12397(.din(n12678),.dout(n12679),.clk(gclk));
	jor g12398(.dina(w_n12675_24[0]),.dinb(w_n12148_1[0]),.dout(n12680),.clk(gclk));
	jnot g12399(.din(w_a28_0[1]),.dout(n12681),.clk(gclk));
	jnot g12400(.din(a[29]),.dout(n12682),.clk(gclk));
	jand g12401(.dina(w_n12148_0[2]),.dinb(w_n12682_0[2]),.dout(n12683),.clk(gclk));
	jand g12402(.dina(n12683),.dinb(w_n12681_1[1]),.dout(n12684),.clk(gclk));
	jnot g12403(.din(n12684),.dout(n12685),.clk(gclk));
	jand g12404(.dina(n12685),.dinb(n12680),.dout(n12686),.clk(gclk));
	jor g12405(.dina(w_n12686_0[2]),.dinb(w_n12670_10[2]),.dout(n12687),.clk(gclk));
	jor g12406(.dina(w_n12675_23[2]),.dinb(w_a30_0[0]),.dout(n12688),.clk(gclk));
	jxor g12407(.dina(w_n12688_0[1]),.dinb(w_n12149_0[0]),.dout(n12689),.clk(gclk));
	jand g12408(.dina(w_n12686_0[1]),.dinb(w_n12670_10[1]),.dout(n12690),.clk(gclk));
	jor g12409(.dina(n12690),.dinb(w_n12689_0[1]),.dout(n12691),.clk(gclk));
	jand g12410(.dina(w_n12691_0[1]),.dinb(w_n12687_0[1]),.dout(n12692),.clk(gclk));
	jor g12411(.dina(n12692),.dinb(w_n11662_15[0]),.dout(n12693),.clk(gclk));
	jand g12412(.dina(w_n12687_0[0]),.dinb(w_n11662_14[2]),.dout(n12694),.clk(gclk));
	jand g12413(.dina(n12694),.dinb(w_n12691_0[0]),.dout(n12695),.clk(gclk));
	jor g12414(.dina(w_n12688_0[0]),.dinb(w_a31_0[0]),.dout(n12696),.clk(gclk));
	jnot g12415(.din(w_n12662_0[0]),.dout(n12697),.clk(gclk));
	jnot g12416(.din(w_n12664_0[0]),.dout(n12698),.clk(gclk));
	jor g12417(.dina(w_n12669_0[0]),.dinb(w_n12670_10[0]),.dout(n12699),.clk(gclk));
	jor g12418(.dina(n12699),.dinb(w_n12698_0[1]),.dout(n12700),.clk(gclk));
	jor g12419(.dina(n12700),.dinb(n12697),.dout(n12701),.clk(gclk));
	jand g12420(.dina(n12701),.dinb(n12696),.dout(n12702),.clk(gclk));
	jxor g12421(.dina(n12702),.dinb(w_n11667_0[1]),.dout(n12703),.clk(gclk));
	jor g12422(.dina(w_n12703_0[1]),.dinb(w_n12695_0[1]),.dout(n12704),.clk(gclk));
	jand g12423(.dina(n12704),.dinb(w_n12693_0[1]),.dout(n12705),.clk(gclk));
	jor g12424(.dina(w_n12705_0[2]),.dinb(w_n11657_10[1]),.dout(n12706),.clk(gclk));
	jand g12425(.dina(w_n12705_0[1]),.dinb(w_n11657_10[0]),.dout(n12707),.clk(gclk));
	jxor g12426(.dina(w_n12152_0[0]),.dinb(w_n11662_14[1]),.dout(n12708),.clk(gclk));
	jor g12427(.dina(n12708),.dinb(w_n12675_23[1]),.dout(n12709),.clk(gclk));
	jxor g12428(.dina(n12709),.dinb(w_n12155_0[0]),.dout(n12710),.clk(gclk));
	jor g12429(.dina(w_n12710_0[1]),.dinb(n12707),.dout(n12711),.clk(gclk));
	jand g12430(.dina(w_n12711_0[1]),.dinb(w_n12706_0[1]),.dout(n12712),.clk(gclk));
	jor g12431(.dina(n12712),.dinb(w_n10701_15[1]),.dout(n12713),.clk(gclk));
	jnot g12432(.din(w_n12161_0[0]),.dout(n12714),.clk(gclk));
	jor g12433(.dina(n12714),.dinb(w_n12159_0[0]),.dout(n12715),.clk(gclk));
	jor g12434(.dina(n12715),.dinb(w_n12675_23[0]),.dout(n12716),.clk(gclk));
	jxor g12435(.dina(n12716),.dinb(w_n12170_0[0]),.dout(n12717),.clk(gclk));
	jand g12436(.dina(w_n12706_0[0]),.dinb(w_n10701_15[0]),.dout(n12718),.clk(gclk));
	jand g12437(.dina(n12718),.dinb(w_n12711_0[0]),.dout(n12719),.clk(gclk));
	jor g12438(.dina(w_n12719_0[1]),.dinb(w_n12717_0[1]),.dout(n12720),.clk(gclk));
	jand g12439(.dina(w_n12720_0[1]),.dinb(w_n12713_0[1]),.dout(n12721),.clk(gclk));
	jor g12440(.dina(w_n12721_0[2]),.dinb(w_n10696_11[0]),.dout(n12722),.clk(gclk));
	jand g12441(.dina(w_n12721_0[1]),.dinb(w_n10696_10[2]),.dout(n12723),.clk(gclk));
	jxor g12442(.dina(w_n12172_0[0]),.dinb(w_n10701_14[2]),.dout(n12724),.clk(gclk));
	jor g12443(.dina(n12724),.dinb(w_n12675_22[2]),.dout(n12725),.clk(gclk));
	jxor g12444(.dina(n12725),.dinb(w_n12177_0[0]),.dout(n12726),.clk(gclk));
	jnot g12445(.din(w_n12726_0[1]),.dout(n12727),.clk(gclk));
	jor g12446(.dina(n12727),.dinb(n12723),.dout(n12728),.clk(gclk));
	jand g12447(.dina(w_n12728_0[1]),.dinb(w_n12722_0[1]),.dout(n12729),.clk(gclk));
	jor g12448(.dina(n12729),.dinb(w_n9774_15[0]),.dout(n12730),.clk(gclk));
	jand g12449(.dina(w_n12722_0[0]),.dinb(w_n9774_14[2]),.dout(n12731),.clk(gclk));
	jand g12450(.dina(n12731),.dinb(w_n12728_0[0]),.dout(n12732),.clk(gclk));
	jnot g12451(.din(w_n12181_0[0]),.dout(n12733),.clk(gclk));
	jnot g12452(.din(w_n12675_22[1]),.dout(asqrt_fa_16),.clk(gclk));
	jand g12453(.dina(w_asqrt15_17),.dinb(n12733),.dout(n12735),.clk(gclk));
	jand g12454(.dina(w_n12735_0[1]),.dinb(w_n12188_0[0]),.dout(n12736),.clk(gclk));
	jor g12455(.dina(n12736),.dinb(w_n12186_0[0]),.dout(n12737),.clk(gclk));
	jand g12456(.dina(w_n12735_0[0]),.dinb(w_n12189_0[0]),.dout(n12738),.clk(gclk));
	jnot g12457(.din(n12738),.dout(n12739),.clk(gclk));
	jand g12458(.dina(n12739),.dinb(n12737),.dout(n12740),.clk(gclk));
	jnot g12459(.din(n12740),.dout(n12741),.clk(gclk));
	jor g12460(.dina(w_n12741_0[1]),.dinb(w_n12732_0[1]),.dout(n12742),.clk(gclk));
	jand g12461(.dina(n12742),.dinb(w_n12730_0[1]),.dout(n12743),.clk(gclk));
	jor g12462(.dina(w_n12743_0[2]),.dinb(w_n9769_11[0]),.dout(n12744),.clk(gclk));
	jand g12463(.dina(w_n12743_0[1]),.dinb(w_n9769_10[2]),.dout(n12745),.clk(gclk));
	jnot g12464(.din(w_n12196_0[0]),.dout(n12746),.clk(gclk));
	jxor g12465(.dina(w_n12190_0[0]),.dinb(w_n9774_14[1]),.dout(n12747),.clk(gclk));
	jor g12466(.dina(n12747),.dinb(w_n12675_22[0]),.dout(n12748),.clk(gclk));
	jxor g12467(.dina(n12748),.dinb(n12746),.dout(n12749),.clk(gclk));
	jnot g12468(.din(w_n12749_0[1]),.dout(n12750),.clk(gclk));
	jor g12469(.dina(n12750),.dinb(n12745),.dout(n12751),.clk(gclk));
	jand g12470(.dina(w_n12751_0[1]),.dinb(w_n12744_0[1]),.dout(n12752),.clk(gclk));
	jor g12471(.dina(n12752),.dinb(w_n8898_15[2]),.dout(n12753),.clk(gclk));
	jnot g12472(.din(w_n12201_0[0]),.dout(n12754),.clk(gclk));
	jor g12473(.dina(n12754),.dinb(w_n12199_0[0]),.dout(n12755),.clk(gclk));
	jor g12474(.dina(n12755),.dinb(w_n12675_21[2]),.dout(n12756),.clk(gclk));
	jxor g12475(.dina(n12756),.dinb(w_n12210_0[0]),.dout(n12757),.clk(gclk));
	jand g12476(.dina(w_n12744_0[0]),.dinb(w_n8898_15[1]),.dout(n12758),.clk(gclk));
	jand g12477(.dina(n12758),.dinb(w_n12751_0[0]),.dout(n12759),.clk(gclk));
	jor g12478(.dina(w_n12759_0[1]),.dinb(w_n12757_0[1]),.dout(n12760),.clk(gclk));
	jand g12479(.dina(w_n12760_0[1]),.dinb(w_n12753_0[1]),.dout(n12761),.clk(gclk));
	jor g12480(.dina(w_n12761_0[2]),.dinb(w_n8893_11[1]),.dout(n12762),.clk(gclk));
	jand g12481(.dina(w_n12761_0[1]),.dinb(w_n8893_11[0]),.dout(n12763),.clk(gclk));
	jnot g12482(.din(w_n12217_0[0]),.dout(n12764),.clk(gclk));
	jxor g12483(.dina(w_n12212_0[0]),.dinb(w_n8898_15[0]),.dout(n12765),.clk(gclk));
	jor g12484(.dina(n12765),.dinb(w_n12675_21[1]),.dout(n12766),.clk(gclk));
	jxor g12485(.dina(n12766),.dinb(n12764),.dout(n12767),.clk(gclk));
	jnot g12486(.din(n12767),.dout(n12768),.clk(gclk));
	jor g12487(.dina(w_n12768_0[1]),.dinb(n12763),.dout(n12769),.clk(gclk));
	jand g12488(.dina(w_n12769_0[1]),.dinb(w_n12762_0[1]),.dout(n12770),.clk(gclk));
	jor g12489(.dina(n12770),.dinb(w_n8058_15[1]),.dout(n12771),.clk(gclk));
	jand g12490(.dina(w_n12762_0[0]),.dinb(w_n8058_15[0]),.dout(n12772),.clk(gclk));
	jand g12491(.dina(n12772),.dinb(w_n12769_0[0]),.dout(n12773),.clk(gclk));
	jnot g12492(.din(w_n12220_0[0]),.dout(n12774),.clk(gclk));
	jand g12493(.dina(w_asqrt15_16[2]),.dinb(n12774),.dout(n12775),.clk(gclk));
	jand g12494(.dina(w_n12775_0[1]),.dinb(w_n12227_0[0]),.dout(n12776),.clk(gclk));
	jor g12495(.dina(n12776),.dinb(w_n12225_0[0]),.dout(n12777),.clk(gclk));
	jand g12496(.dina(w_n12775_0[0]),.dinb(w_n12228_0[0]),.dout(n12778),.clk(gclk));
	jnot g12497(.din(n12778),.dout(n12779),.clk(gclk));
	jand g12498(.dina(n12779),.dinb(n12777),.dout(n12780),.clk(gclk));
	jnot g12499(.din(n12780),.dout(n12781),.clk(gclk));
	jor g12500(.dina(w_n12781_0[1]),.dinb(w_n12773_0[1]),.dout(n12782),.clk(gclk));
	jand g12501(.dina(n12782),.dinb(w_n12771_0[1]),.dout(n12783),.clk(gclk));
	jor g12502(.dina(w_n12783_0[1]),.dinb(w_n8053_11[1]),.dout(n12784),.clk(gclk));
	jxor g12503(.dina(w_n12229_0[0]),.dinb(w_n8058_14[2]),.dout(n12785),.clk(gclk));
	jor g12504(.dina(n12785),.dinb(w_n12675_21[0]),.dout(n12786),.clk(gclk));
	jxor g12505(.dina(n12786),.dinb(w_n12234_0[0]),.dout(n12787),.clk(gclk));
	jand g12506(.dina(w_n12783_0[0]),.dinb(w_n8053_11[0]),.dout(n12788),.clk(gclk));
	jor g12507(.dina(w_n12788_0[1]),.dinb(w_n12787_0[1]),.dout(n12789),.clk(gclk));
	jand g12508(.dina(w_n12789_0[2]),.dinb(w_n12784_0[2]),.dout(n12790),.clk(gclk));
	jor g12509(.dina(n12790),.dinb(w_n7265_15[2]),.dout(n12791),.clk(gclk));
	jnot g12510(.din(w_n12239_0[0]),.dout(n12792),.clk(gclk));
	jor g12511(.dina(n12792),.dinb(w_n12237_0[0]),.dout(n12793),.clk(gclk));
	jor g12512(.dina(n12793),.dinb(w_n12675_20[2]),.dout(n12794),.clk(gclk));
	jxor g12513(.dina(n12794),.dinb(w_n12248_0[0]),.dout(n12795),.clk(gclk));
	jand g12514(.dina(w_n12784_0[1]),.dinb(w_n7265_15[1]),.dout(n12796),.clk(gclk));
	jand g12515(.dina(n12796),.dinb(w_n12789_0[1]),.dout(n12797),.clk(gclk));
	jor g12516(.dina(w_n12797_0[1]),.dinb(w_n12795_0[1]),.dout(n12798),.clk(gclk));
	jand g12517(.dina(w_n12798_0[1]),.dinb(w_n12791_0[1]),.dout(n12799),.clk(gclk));
	jor g12518(.dina(w_n12799_0[2]),.dinb(w_n7260_12[1]),.dout(n12800),.clk(gclk));
	jand g12519(.dina(w_n12799_0[1]),.dinb(w_n7260_12[0]),.dout(n12801),.clk(gclk));
	jnot g12520(.din(w_n12251_0[0]),.dout(n12802),.clk(gclk));
	jand g12521(.dina(w_asqrt15_16[1]),.dinb(n12802),.dout(n12803),.clk(gclk));
	jand g12522(.dina(w_n12803_0[1]),.dinb(w_n12256_0[0]),.dout(n12804),.clk(gclk));
	jor g12523(.dina(n12804),.dinb(w_n12255_0[0]),.dout(n12805),.clk(gclk));
	jand g12524(.dina(w_n12803_0[0]),.dinb(w_n12257_0[0]),.dout(n12806),.clk(gclk));
	jnot g12525(.din(n12806),.dout(n12807),.clk(gclk));
	jand g12526(.dina(n12807),.dinb(n12805),.dout(n12808),.clk(gclk));
	jnot g12527(.din(n12808),.dout(n12809),.clk(gclk));
	jor g12528(.dina(w_n12809_0[1]),.dinb(n12801),.dout(n12810),.clk(gclk));
	jand g12529(.dina(w_n12810_0[1]),.dinb(w_n12800_0[1]),.dout(n12811),.clk(gclk));
	jor g12530(.dina(n12811),.dinb(w_n6505_15[2]),.dout(n12812),.clk(gclk));
	jand g12531(.dina(w_n12800_0[0]),.dinb(w_n6505_15[1]),.dout(n12813),.clk(gclk));
	jand g12532(.dina(n12813),.dinb(w_n12810_0[0]),.dout(n12814),.clk(gclk));
	jnot g12533(.din(w_n12259_0[0]),.dout(n12815),.clk(gclk));
	jand g12534(.dina(w_asqrt15_16[0]),.dinb(n12815),.dout(n12816),.clk(gclk));
	jand g12535(.dina(w_n12816_0[1]),.dinb(w_n12266_0[0]),.dout(n12817),.clk(gclk));
	jor g12536(.dina(n12817),.dinb(w_n12264_0[0]),.dout(n12818),.clk(gclk));
	jand g12537(.dina(w_n12816_0[0]),.dinb(w_n12267_0[0]),.dout(n12819),.clk(gclk));
	jnot g12538(.din(n12819),.dout(n12820),.clk(gclk));
	jand g12539(.dina(n12820),.dinb(n12818),.dout(n12821),.clk(gclk));
	jnot g12540(.din(n12821),.dout(n12822),.clk(gclk));
	jor g12541(.dina(w_n12822_0[1]),.dinb(w_n12814_0[1]),.dout(n12823),.clk(gclk));
	jand g12542(.dina(n12823),.dinb(w_n12812_0[1]),.dout(n12824),.clk(gclk));
	jor g12543(.dina(w_n12824_0[1]),.dinb(w_n6500_12[1]),.dout(n12825),.clk(gclk));
	jxor g12544(.dina(w_n12268_0[0]),.dinb(w_n6505_15[0]),.dout(n12826),.clk(gclk));
	jor g12545(.dina(n12826),.dinb(w_n12675_20[1]),.dout(n12827),.clk(gclk));
	jxor g12546(.dina(n12827),.dinb(w_n12279_0[0]),.dout(n12828),.clk(gclk));
	jand g12547(.dina(w_n12824_0[0]),.dinb(w_n6500_12[0]),.dout(n12829),.clk(gclk));
	jor g12548(.dina(w_n12829_0[1]),.dinb(w_n12828_0[1]),.dout(n12830),.clk(gclk));
	jand g12549(.dina(w_n12830_0[2]),.dinb(w_n12825_0[2]),.dout(n12831),.clk(gclk));
	jor g12550(.dina(n12831),.dinb(w_n5793_16[0]),.dout(n12832),.clk(gclk));
	jnot g12551(.din(w_n12284_0[0]),.dout(n12833),.clk(gclk));
	jor g12552(.dina(n12833),.dinb(w_n12282_0[0]),.dout(n12834),.clk(gclk));
	jor g12553(.dina(n12834),.dinb(w_n12675_20[0]),.dout(n12835),.clk(gclk));
	jxor g12554(.dina(n12835),.dinb(w_n12293_0[0]),.dout(n12836),.clk(gclk));
	jand g12555(.dina(w_n12825_0[1]),.dinb(w_n5793_15[2]),.dout(n12837),.clk(gclk));
	jand g12556(.dina(n12837),.dinb(w_n12830_0[1]),.dout(n12838),.clk(gclk));
	jor g12557(.dina(w_n12838_0[1]),.dinb(w_n12836_0[1]),.dout(n12839),.clk(gclk));
	jand g12558(.dina(w_n12839_0[1]),.dinb(w_n12832_0[1]),.dout(n12840),.clk(gclk));
	jor g12559(.dina(w_n12840_0[2]),.dinb(w_n5788_13[0]),.dout(n12841),.clk(gclk));
	jand g12560(.dina(w_n12840_0[1]),.dinb(w_n5788_12[2]),.dout(n12842),.clk(gclk));
	jnot g12561(.din(w_n12296_0[0]),.dout(n12843),.clk(gclk));
	jand g12562(.dina(w_asqrt15_15[2]),.dinb(n12843),.dout(n12844),.clk(gclk));
	jand g12563(.dina(w_n12844_0[1]),.dinb(w_n12301_0[0]),.dout(n12845),.clk(gclk));
	jor g12564(.dina(n12845),.dinb(w_n12300_0[0]),.dout(n12846),.clk(gclk));
	jand g12565(.dina(w_n12844_0[0]),.dinb(w_n12302_0[0]),.dout(n12847),.clk(gclk));
	jnot g12566(.din(n12847),.dout(n12848),.clk(gclk));
	jand g12567(.dina(n12848),.dinb(n12846),.dout(n12849),.clk(gclk));
	jnot g12568(.din(n12849),.dout(n12850),.clk(gclk));
	jor g12569(.dina(w_n12850_0[1]),.dinb(n12842),.dout(n12851),.clk(gclk));
	jand g12570(.dina(w_n12851_0[1]),.dinb(w_n12841_0[1]),.dout(n12852),.clk(gclk));
	jor g12571(.dina(n12852),.dinb(w_n5121_16[0]),.dout(n12853),.clk(gclk));
	jand g12572(.dina(w_n12841_0[0]),.dinb(w_n5121_15[2]),.dout(n12854),.clk(gclk));
	jand g12573(.dina(n12854),.dinb(w_n12851_0[0]),.dout(n12855),.clk(gclk));
	jnot g12574(.din(w_n12304_0[0]),.dout(n12856),.clk(gclk));
	jand g12575(.dina(w_asqrt15_15[1]),.dinb(n12856),.dout(n12857),.clk(gclk));
	jand g12576(.dina(w_n12857_0[1]),.dinb(w_n12311_0[0]),.dout(n12858),.clk(gclk));
	jor g12577(.dina(n12858),.dinb(w_n12309_0[0]),.dout(n12859),.clk(gclk));
	jand g12578(.dina(w_n12857_0[0]),.dinb(w_n12312_0[0]),.dout(n12860),.clk(gclk));
	jnot g12579(.din(n12860),.dout(n12861),.clk(gclk));
	jand g12580(.dina(n12861),.dinb(n12859),.dout(n12862),.clk(gclk));
	jnot g12581(.din(n12862),.dout(n12863),.clk(gclk));
	jor g12582(.dina(w_n12863_0[1]),.dinb(w_n12855_0[1]),.dout(n12864),.clk(gclk));
	jand g12583(.dina(n12864),.dinb(w_n12853_0[1]),.dout(n12865),.clk(gclk));
	jor g12584(.dina(w_n12865_0[1]),.dinb(w_n5116_13[0]),.dout(n12866),.clk(gclk));
	jxor g12585(.dina(w_n12313_0[0]),.dinb(w_n5121_15[1]),.dout(n12867),.clk(gclk));
	jor g12586(.dina(n12867),.dinb(w_n12675_19[2]),.dout(n12868),.clk(gclk));
	jxor g12587(.dina(n12868),.dinb(w_n12324_0[0]),.dout(n12869),.clk(gclk));
	jand g12588(.dina(w_n12865_0[0]),.dinb(w_n5116_12[2]),.dout(n12870),.clk(gclk));
	jor g12589(.dina(w_n12870_0[1]),.dinb(w_n12869_0[1]),.dout(n12871),.clk(gclk));
	jand g12590(.dina(w_n12871_0[2]),.dinb(w_n12866_0[2]),.dout(n12872),.clk(gclk));
	jor g12591(.dina(n12872),.dinb(w_n4499_16[2]),.dout(n12873),.clk(gclk));
	jnot g12592(.din(w_n12329_0[0]),.dout(n12874),.clk(gclk));
	jor g12593(.dina(n12874),.dinb(w_n12327_0[0]),.dout(n12875),.clk(gclk));
	jor g12594(.dina(n12875),.dinb(w_n12675_19[1]),.dout(n12876),.clk(gclk));
	jxor g12595(.dina(n12876),.dinb(w_n12338_0[0]),.dout(n12877),.clk(gclk));
	jand g12596(.dina(w_n12866_0[1]),.dinb(w_n4499_16[1]),.dout(n12878),.clk(gclk));
	jand g12597(.dina(n12878),.dinb(w_n12871_0[1]),.dout(n12879),.clk(gclk));
	jor g12598(.dina(w_n12879_0[1]),.dinb(w_n12877_0[1]),.dout(n12880),.clk(gclk));
	jand g12599(.dina(w_n12880_0[1]),.dinb(w_n12873_0[1]),.dout(n12881),.clk(gclk));
	jor g12600(.dina(w_n12881_0[2]),.dinb(w_n4494_14[0]),.dout(n12882),.clk(gclk));
	jand g12601(.dina(w_n12881_0[1]),.dinb(w_n4494_13[2]),.dout(n12883),.clk(gclk));
	jnot g12602(.din(w_n12341_0[0]),.dout(n12884),.clk(gclk));
	jand g12603(.dina(w_asqrt15_15[0]),.dinb(n12884),.dout(n12885),.clk(gclk));
	jand g12604(.dina(w_n12885_0[1]),.dinb(w_n12346_0[0]),.dout(n12886),.clk(gclk));
	jor g12605(.dina(n12886),.dinb(w_n12345_0[0]),.dout(n12887),.clk(gclk));
	jand g12606(.dina(w_n12885_0[0]),.dinb(w_n12347_0[0]),.dout(n12888),.clk(gclk));
	jnot g12607(.din(n12888),.dout(n12889),.clk(gclk));
	jand g12608(.dina(n12889),.dinb(n12887),.dout(n12890),.clk(gclk));
	jnot g12609(.din(n12890),.dout(n12891),.clk(gclk));
	jor g12610(.dina(w_n12891_0[1]),.dinb(n12883),.dout(n12892),.clk(gclk));
	jand g12611(.dina(w_n12892_0[1]),.dinb(w_n12882_0[1]),.dout(n12893),.clk(gclk));
	jor g12612(.dina(n12893),.dinb(w_n3912_16[2]),.dout(n12894),.clk(gclk));
	jand g12613(.dina(w_n12882_0[0]),.dinb(w_n3912_16[1]),.dout(n12895),.clk(gclk));
	jand g12614(.dina(n12895),.dinb(w_n12892_0[0]),.dout(n12896),.clk(gclk));
	jnot g12615(.din(w_n12349_0[0]),.dout(n12897),.clk(gclk));
	jand g12616(.dina(w_asqrt15_14[2]),.dinb(n12897),.dout(n12898),.clk(gclk));
	jand g12617(.dina(w_n12898_0[1]),.dinb(w_n12356_0[0]),.dout(n12899),.clk(gclk));
	jor g12618(.dina(n12899),.dinb(w_n12354_0[0]),.dout(n12900),.clk(gclk));
	jand g12619(.dina(w_n12898_0[0]),.dinb(w_n12357_0[0]),.dout(n12901),.clk(gclk));
	jnot g12620(.din(n12901),.dout(n12902),.clk(gclk));
	jand g12621(.dina(n12902),.dinb(n12900),.dout(n12903),.clk(gclk));
	jnot g12622(.din(n12903),.dout(n12904),.clk(gclk));
	jor g12623(.dina(w_n12904_0[1]),.dinb(w_n12896_0[1]),.dout(n12905),.clk(gclk));
	jand g12624(.dina(n12905),.dinb(w_n12894_0[1]),.dout(n12906),.clk(gclk));
	jor g12625(.dina(w_n12906_0[1]),.dinb(w_n3907_14[0]),.dout(n12907),.clk(gclk));
	jxor g12626(.dina(w_n12358_0[0]),.dinb(w_n3912_16[0]),.dout(n12908),.clk(gclk));
	jor g12627(.dina(n12908),.dinb(w_n12675_19[0]),.dout(n12909),.clk(gclk));
	jxor g12628(.dina(n12909),.dinb(w_n12369_0[0]),.dout(n12910),.clk(gclk));
	jand g12629(.dina(w_n12906_0[0]),.dinb(w_n3907_13[2]),.dout(n12911),.clk(gclk));
	jor g12630(.dina(w_n12911_0[1]),.dinb(w_n12910_0[1]),.dout(n12912),.clk(gclk));
	jand g12631(.dina(w_n12912_0[2]),.dinb(w_n12907_0[2]),.dout(n12913),.clk(gclk));
	jor g12632(.dina(n12913),.dinb(w_n3376_17[1]),.dout(n12914),.clk(gclk));
	jnot g12633(.din(w_n12374_0[0]),.dout(n12915),.clk(gclk));
	jor g12634(.dina(n12915),.dinb(w_n12372_0[0]),.dout(n12916),.clk(gclk));
	jor g12635(.dina(n12916),.dinb(w_n12675_18[2]),.dout(n12917),.clk(gclk));
	jxor g12636(.dina(n12917),.dinb(w_n12383_0[0]),.dout(n12918),.clk(gclk));
	jand g12637(.dina(w_n12907_0[1]),.dinb(w_n3376_17[0]),.dout(n12919),.clk(gclk));
	jand g12638(.dina(n12919),.dinb(w_n12912_0[1]),.dout(n12920),.clk(gclk));
	jor g12639(.dina(w_n12920_0[1]),.dinb(w_n12918_0[1]),.dout(n12921),.clk(gclk));
	jand g12640(.dina(w_n12921_0[1]),.dinb(w_n12914_0[1]),.dout(n12922),.clk(gclk));
	jor g12641(.dina(w_n12922_0[2]),.dinb(w_n3371_14[2]),.dout(n12923),.clk(gclk));
	jand g12642(.dina(w_n12922_0[1]),.dinb(w_n3371_14[1]),.dout(n12924),.clk(gclk));
	jnot g12643(.din(w_n12386_0[0]),.dout(n12925),.clk(gclk));
	jand g12644(.dina(w_asqrt15_14[1]),.dinb(n12925),.dout(n12926),.clk(gclk));
	jand g12645(.dina(w_n12926_0[1]),.dinb(w_n12391_0[0]),.dout(n12927),.clk(gclk));
	jor g12646(.dina(n12927),.dinb(w_n12390_0[0]),.dout(n12928),.clk(gclk));
	jand g12647(.dina(w_n12926_0[0]),.dinb(w_n12392_0[0]),.dout(n12929),.clk(gclk));
	jnot g12648(.din(n12929),.dout(n12930),.clk(gclk));
	jand g12649(.dina(n12930),.dinb(n12928),.dout(n12931),.clk(gclk));
	jnot g12650(.din(n12931),.dout(n12932),.clk(gclk));
	jor g12651(.dina(w_n12932_0[1]),.dinb(n12924),.dout(n12933),.clk(gclk));
	jand g12652(.dina(w_n12933_0[1]),.dinb(w_n12923_0[1]),.dout(n12934),.clk(gclk));
	jor g12653(.dina(n12934),.dinb(w_n2875_17[1]),.dout(n12935),.clk(gclk));
	jand g12654(.dina(w_n12923_0[0]),.dinb(w_n2875_17[0]),.dout(n12936),.clk(gclk));
	jand g12655(.dina(n12936),.dinb(w_n12933_0[0]),.dout(n12937),.clk(gclk));
	jnot g12656(.din(w_n12394_0[0]),.dout(n12938),.clk(gclk));
	jand g12657(.dina(w_asqrt15_14[0]),.dinb(n12938),.dout(n12939),.clk(gclk));
	jand g12658(.dina(w_n12939_0[1]),.dinb(w_n12401_0[0]),.dout(n12940),.clk(gclk));
	jor g12659(.dina(n12940),.dinb(w_n12399_0[0]),.dout(n12941),.clk(gclk));
	jand g12660(.dina(w_n12939_0[0]),.dinb(w_n12402_0[0]),.dout(n12942),.clk(gclk));
	jnot g12661(.din(n12942),.dout(n12943),.clk(gclk));
	jand g12662(.dina(n12943),.dinb(n12941),.dout(n12944),.clk(gclk));
	jnot g12663(.din(n12944),.dout(n12945),.clk(gclk));
	jor g12664(.dina(w_n12945_0[1]),.dinb(w_n12937_0[1]),.dout(n12946),.clk(gclk));
	jand g12665(.dina(n12946),.dinb(w_n12935_0[1]),.dout(n12947),.clk(gclk));
	jor g12666(.dina(w_n12947_0[1]),.dinb(w_n2870_14[2]),.dout(n12948),.clk(gclk));
	jxor g12667(.dina(w_n12403_0[0]),.dinb(w_n2875_16[2]),.dout(n12949),.clk(gclk));
	jor g12668(.dina(n12949),.dinb(w_n12675_18[1]),.dout(n12950),.clk(gclk));
	jxor g12669(.dina(n12950),.dinb(w_n12414_0[0]),.dout(n12951),.clk(gclk));
	jand g12670(.dina(w_n12947_0[0]),.dinb(w_n2870_14[1]),.dout(n12952),.clk(gclk));
	jor g12671(.dina(w_n12952_0[1]),.dinb(w_n12951_0[1]),.dout(n12953),.clk(gclk));
	jand g12672(.dina(w_n12953_0[2]),.dinb(w_n12948_0[2]),.dout(n12954),.clk(gclk));
	jor g12673(.dina(n12954),.dinb(w_n2425_17[2]),.dout(n12955),.clk(gclk));
	jnot g12674(.din(w_n12419_0[0]),.dout(n12956),.clk(gclk));
	jor g12675(.dina(n12956),.dinb(w_n12417_0[0]),.dout(n12957),.clk(gclk));
	jor g12676(.dina(n12957),.dinb(w_n12675_18[0]),.dout(n12958),.clk(gclk));
	jxor g12677(.dina(n12958),.dinb(w_n12428_0[0]),.dout(n12959),.clk(gclk));
	jand g12678(.dina(w_n12948_0[1]),.dinb(w_n2425_17[1]),.dout(n12960),.clk(gclk));
	jand g12679(.dina(n12960),.dinb(w_n12953_0[1]),.dout(n12961),.clk(gclk));
	jor g12680(.dina(w_n12961_0[1]),.dinb(w_n12959_0[1]),.dout(n12962),.clk(gclk));
	jand g12681(.dina(w_n12962_0[1]),.dinb(w_n12955_0[1]),.dout(n12963),.clk(gclk));
	jor g12682(.dina(w_n12963_0[2]),.dinb(w_n2420_15[2]),.dout(n12964),.clk(gclk));
	jand g12683(.dina(w_n12963_0[1]),.dinb(w_n2420_15[1]),.dout(n12965),.clk(gclk));
	jnot g12684(.din(w_n12431_0[0]),.dout(n12966),.clk(gclk));
	jand g12685(.dina(w_asqrt15_13[2]),.dinb(n12966),.dout(n12967),.clk(gclk));
	jand g12686(.dina(w_n12967_0[1]),.dinb(w_n12436_0[0]),.dout(n12968),.clk(gclk));
	jor g12687(.dina(n12968),.dinb(w_n12435_0[0]),.dout(n12969),.clk(gclk));
	jand g12688(.dina(w_n12967_0[0]),.dinb(w_n12437_0[0]),.dout(n12970),.clk(gclk));
	jnot g12689(.din(n12970),.dout(n12971),.clk(gclk));
	jand g12690(.dina(n12971),.dinb(n12969),.dout(n12972),.clk(gclk));
	jnot g12691(.din(n12972),.dout(n12973),.clk(gclk));
	jor g12692(.dina(w_n12973_0[1]),.dinb(n12965),.dout(n12974),.clk(gclk));
	jand g12693(.dina(w_n12974_0[1]),.dinb(w_n12964_0[1]),.dout(n12975),.clk(gclk));
	jor g12694(.dina(n12975),.dinb(w_n2010_17[2]),.dout(n12976),.clk(gclk));
	jand g12695(.dina(w_n12964_0[0]),.dinb(w_n2010_17[1]),.dout(n12977),.clk(gclk));
	jand g12696(.dina(n12977),.dinb(w_n12974_0[0]),.dout(n12978),.clk(gclk));
	jnot g12697(.din(w_n12439_0[0]),.dout(n12979),.clk(gclk));
	jand g12698(.dina(w_asqrt15_13[1]),.dinb(n12979),.dout(n12980),.clk(gclk));
	jand g12699(.dina(w_n12980_0[1]),.dinb(w_n12446_0[0]),.dout(n12981),.clk(gclk));
	jor g12700(.dina(n12981),.dinb(w_n12444_0[0]),.dout(n12982),.clk(gclk));
	jand g12701(.dina(w_n12980_0[0]),.dinb(w_n12447_0[0]),.dout(n12983),.clk(gclk));
	jnot g12702(.din(n12983),.dout(n12984),.clk(gclk));
	jand g12703(.dina(n12984),.dinb(n12982),.dout(n12985),.clk(gclk));
	jnot g12704(.din(n12985),.dout(n12986),.clk(gclk));
	jor g12705(.dina(w_n12986_0[1]),.dinb(w_n12978_0[1]),.dout(n12987),.clk(gclk));
	jand g12706(.dina(n12987),.dinb(w_n12976_0[1]),.dout(n12988),.clk(gclk));
	jor g12707(.dina(w_n12988_0[1]),.dinb(w_n2005_15[2]),.dout(n12989),.clk(gclk));
	jxor g12708(.dina(w_n12448_0[0]),.dinb(w_n2010_17[0]),.dout(n12990),.clk(gclk));
	jor g12709(.dina(n12990),.dinb(w_n12675_17[2]),.dout(n12991),.clk(gclk));
	jxor g12710(.dina(n12991),.dinb(w_n12459_0[0]),.dout(n12992),.clk(gclk));
	jand g12711(.dina(w_n12988_0[0]),.dinb(w_n2005_15[1]),.dout(n12993),.clk(gclk));
	jor g12712(.dina(w_n12993_0[1]),.dinb(w_n12992_0[1]),.dout(n12994),.clk(gclk));
	jand g12713(.dina(w_n12994_0[2]),.dinb(w_n12989_0[2]),.dout(n12995),.clk(gclk));
	jor g12714(.dina(n12995),.dinb(w_n1646_18[1]),.dout(n12996),.clk(gclk));
	jand g12715(.dina(w_n12989_0[1]),.dinb(w_n1646_18[0]),.dout(n12997),.clk(gclk));
	jand g12716(.dina(n12997),.dinb(w_n12994_0[1]),.dout(n12998),.clk(gclk));
	jnot g12717(.din(w_n12462_0[0]),.dout(n12999),.clk(gclk));
	jand g12718(.dina(w_asqrt15_13[0]),.dinb(n12999),.dout(n13000),.clk(gclk));
	jand g12719(.dina(w_n13000_0[1]),.dinb(w_n12469_0[0]),.dout(n13001),.clk(gclk));
	jor g12720(.dina(n13001),.dinb(w_n12467_0[0]),.dout(n13002),.clk(gclk));
	jand g12721(.dina(w_n13000_0[0]),.dinb(w_n12470_0[0]),.dout(n13003),.clk(gclk));
	jnot g12722(.din(n13003),.dout(n13004),.clk(gclk));
	jand g12723(.dina(n13004),.dinb(n13002),.dout(n13005),.clk(gclk));
	jnot g12724(.din(n13005),.dout(n13006),.clk(gclk));
	jor g12725(.dina(w_n13006_0[1]),.dinb(w_n12998_0[1]),.dout(n13007),.clk(gclk));
	jand g12726(.dina(n13007),.dinb(w_n12996_0[1]),.dout(n13008),.clk(gclk));
	jor g12727(.dina(w_n13008_0[2]),.dinb(w_n1641_16[1]),.dout(n13009),.clk(gclk));
	jand g12728(.dina(w_n13008_0[1]),.dinb(w_n1641_16[0]),.dout(n13010),.clk(gclk));
	jor g12729(.dina(n13010),.dinb(w_n12679_0[1]),.dout(n13011),.clk(gclk));
	jand g12730(.dina(w_n13011_0[1]),.dinb(w_n13009_0[1]),.dout(n13012),.clk(gclk));
	jor g12731(.dina(n13012),.dinb(w_n1317_18[2]),.dout(n13013),.clk(gclk));
	jnot g12732(.din(w_n12478_0[0]),.dout(n13014),.clk(gclk));
	jor g12733(.dina(n13014),.dinb(w_n12476_0[0]),.dout(n13015),.clk(gclk));
	jor g12734(.dina(n13015),.dinb(w_n12675_17[1]),.dout(n13016),.clk(gclk));
	jxor g12735(.dina(n13016),.dinb(w_n12487_0[0]),.dout(n13017),.clk(gclk));
	jand g12736(.dina(w_n13009_0[0]),.dinb(w_n1317_18[1]),.dout(n13018),.clk(gclk));
	jand g12737(.dina(n13018),.dinb(w_n13011_0[0]),.dout(n13019),.clk(gclk));
	jor g12738(.dina(w_n13019_0[1]),.dinb(w_n13017_0[1]),.dout(n13020),.clk(gclk));
	jand g12739(.dina(w_n13020_0[1]),.dinb(w_n13013_0[1]),.dout(n13021),.clk(gclk));
	jor g12740(.dina(w_n13021_0[1]),.dinb(w_n1312_16[1]),.dout(n13022),.clk(gclk));
	jxor g12741(.dina(w_n12489_0[0]),.dinb(w_n1317_18[0]),.dout(n13023),.clk(gclk));
	jor g12742(.dina(n13023),.dinb(w_n12675_17[0]),.dout(n13024),.clk(gclk));
	jxor g12743(.dina(n13024),.dinb(w_n12500_0[0]),.dout(n13025),.clk(gclk));
	jand g12744(.dina(w_n13021_0[0]),.dinb(w_n1312_16[0]),.dout(n13026),.clk(gclk));
	jor g12745(.dina(w_n13026_0[1]),.dinb(w_n13025_0[1]),.dout(n13027),.clk(gclk));
	jand g12746(.dina(w_n13027_0[2]),.dinb(w_n13022_0[2]),.dout(n13028),.clk(gclk));
	jor g12747(.dina(n13028),.dinb(w_n1039_19[0]),.dout(n13029),.clk(gclk));
	jnot g12748(.din(w_n12505_0[0]),.dout(n13030),.clk(gclk));
	jor g12749(.dina(n13030),.dinb(w_n12503_0[0]),.dout(n13031),.clk(gclk));
	jor g12750(.dina(n13031),.dinb(w_n12675_16[2]),.dout(n13032),.clk(gclk));
	jxor g12751(.dina(n13032),.dinb(w_n12514_0[0]),.dout(n13033),.clk(gclk));
	jand g12752(.dina(w_n13022_0[1]),.dinb(w_n1039_18[2]),.dout(n13034),.clk(gclk));
	jand g12753(.dina(n13034),.dinb(w_n13027_0[1]),.dout(n13035),.clk(gclk));
	jor g12754(.dina(w_n13035_0[1]),.dinb(w_n13033_0[1]),.dout(n13036),.clk(gclk));
	jand g12755(.dina(w_n13036_0[1]),.dinb(w_n13029_0[1]),.dout(n13037),.clk(gclk));
	jor g12756(.dina(w_n13037_0[2]),.dinb(w_n1034_17[1]),.dout(n13038),.clk(gclk));
	jand g12757(.dina(w_n13037_0[1]),.dinb(w_n1034_17[0]),.dout(n13039),.clk(gclk));
	jnot g12758(.din(w_n12517_0[0]),.dout(n13040),.clk(gclk));
	jand g12759(.dina(w_asqrt15_12[2]),.dinb(n13040),.dout(n13041),.clk(gclk));
	jand g12760(.dina(w_n13041_0[1]),.dinb(w_n12522_0[0]),.dout(n13042),.clk(gclk));
	jor g12761(.dina(n13042),.dinb(w_n12521_0[0]),.dout(n13043),.clk(gclk));
	jand g12762(.dina(w_n13041_0[0]),.dinb(w_n12523_0[0]),.dout(n13044),.clk(gclk));
	jnot g12763(.din(n13044),.dout(n13045),.clk(gclk));
	jand g12764(.dina(n13045),.dinb(n13043),.dout(n13046),.clk(gclk));
	jnot g12765(.din(n13046),.dout(n13047),.clk(gclk));
	jor g12766(.dina(w_n13047_0[1]),.dinb(n13039),.dout(n13048),.clk(gclk));
	jand g12767(.dina(w_n13048_0[1]),.dinb(w_n13038_0[1]),.dout(n13049),.clk(gclk));
	jor g12768(.dina(n13049),.dinb(w_n796_19[0]),.dout(n13050),.clk(gclk));
	jand g12769(.dina(w_n13038_0[0]),.dinb(w_n796_18[2]),.dout(n13051),.clk(gclk));
	jand g12770(.dina(n13051),.dinb(w_n13048_0[0]),.dout(n13052),.clk(gclk));
	jnot g12771(.din(w_n12525_0[0]),.dout(n13053),.clk(gclk));
	jand g12772(.dina(w_asqrt15_12[1]),.dinb(n13053),.dout(n13054),.clk(gclk));
	jand g12773(.dina(w_n13054_0[1]),.dinb(w_n12532_0[0]),.dout(n13055),.clk(gclk));
	jor g12774(.dina(n13055),.dinb(w_n12530_0[0]),.dout(n13056),.clk(gclk));
	jand g12775(.dina(w_n13054_0[0]),.dinb(w_n12533_0[0]),.dout(n13057),.clk(gclk));
	jnot g12776(.din(n13057),.dout(n13058),.clk(gclk));
	jand g12777(.dina(n13058),.dinb(n13056),.dout(n13059),.clk(gclk));
	jnot g12778(.din(n13059),.dout(n13060),.clk(gclk));
	jor g12779(.dina(w_n13060_0[1]),.dinb(w_n13052_0[1]),.dout(n13061),.clk(gclk));
	jand g12780(.dina(n13061),.dinb(w_n13050_0[1]),.dout(n13062),.clk(gclk));
	jor g12781(.dina(w_n13062_0[1]),.dinb(w_n791_17[1]),.dout(n13063),.clk(gclk));
	jxor g12782(.dina(w_n12534_0[0]),.dinb(w_n796_18[1]),.dout(n13064),.clk(gclk));
	jor g12783(.dina(n13064),.dinb(w_n12675_16[1]),.dout(n13065),.clk(gclk));
	jxor g12784(.dina(n13065),.dinb(w_n12545_0[0]),.dout(n13066),.clk(gclk));
	jand g12785(.dina(w_n13062_0[0]),.dinb(w_n791_17[0]),.dout(n13067),.clk(gclk));
	jor g12786(.dina(w_n13067_0[1]),.dinb(w_n13066_0[1]),.dout(n13068),.clk(gclk));
	jand g12787(.dina(w_n13068_0[2]),.dinb(w_n13063_0[2]),.dout(n13069),.clk(gclk));
	jor g12788(.dina(n13069),.dinb(w_n595_19[1]),.dout(n13070),.clk(gclk));
	jnot g12789(.din(w_n12550_0[0]),.dout(n13071),.clk(gclk));
	jor g12790(.dina(n13071),.dinb(w_n12548_0[0]),.dout(n13072),.clk(gclk));
	jor g12791(.dina(n13072),.dinb(w_n12675_16[0]),.dout(n13073),.clk(gclk));
	jxor g12792(.dina(n13073),.dinb(w_n12559_0[0]),.dout(n13074),.clk(gclk));
	jand g12793(.dina(w_n13063_0[1]),.dinb(w_n595_19[0]),.dout(n13075),.clk(gclk));
	jand g12794(.dina(n13075),.dinb(w_n13068_0[1]),.dout(n13076),.clk(gclk));
	jor g12795(.dina(w_n13076_0[1]),.dinb(w_n13074_0[1]),.dout(n13077),.clk(gclk));
	jand g12796(.dina(w_n13077_0[1]),.dinb(w_n13070_0[1]),.dout(n13078),.clk(gclk));
	jor g12797(.dina(w_n13078_0[2]),.dinb(w_n590_18[0]),.dout(n13079),.clk(gclk));
	jand g12798(.dina(w_n13078_0[1]),.dinb(w_n590_17[2]),.dout(n13080),.clk(gclk));
	jnot g12799(.din(w_n12562_0[0]),.dout(n13081),.clk(gclk));
	jand g12800(.dina(w_asqrt15_12[0]),.dinb(n13081),.dout(n13082),.clk(gclk));
	jand g12801(.dina(w_n13082_0[1]),.dinb(w_n12567_0[0]),.dout(n13083),.clk(gclk));
	jor g12802(.dina(n13083),.dinb(w_n12566_0[0]),.dout(n13084),.clk(gclk));
	jand g12803(.dina(w_n13082_0[0]),.dinb(w_n12568_0[0]),.dout(n13085),.clk(gclk));
	jnot g12804(.din(n13085),.dout(n13086),.clk(gclk));
	jand g12805(.dina(n13086),.dinb(n13084),.dout(n13087),.clk(gclk));
	jnot g12806(.din(n13087),.dout(n13088),.clk(gclk));
	jor g12807(.dina(w_n13088_0[1]),.dinb(n13080),.dout(n13089),.clk(gclk));
	jand g12808(.dina(w_n13089_0[1]),.dinb(w_n13079_0[1]),.dout(n13090),.clk(gclk));
	jor g12809(.dina(n13090),.dinb(w_n430_19[1]),.dout(n13091),.clk(gclk));
	jand g12810(.dina(w_n13079_0[0]),.dinb(w_n430_19[0]),.dout(n13092),.clk(gclk));
	jand g12811(.dina(n13092),.dinb(w_n13089_0[0]),.dout(n13093),.clk(gclk));
	jnot g12812(.din(w_n12570_0[0]),.dout(n13094),.clk(gclk));
	jand g12813(.dina(w_asqrt15_11[2]),.dinb(n13094),.dout(n13095),.clk(gclk));
	jand g12814(.dina(w_n13095_0[1]),.dinb(w_n12577_0[0]),.dout(n13096),.clk(gclk));
	jor g12815(.dina(n13096),.dinb(w_n12575_0[0]),.dout(n13097),.clk(gclk));
	jand g12816(.dina(w_n13095_0[0]),.dinb(w_n12578_0[0]),.dout(n13098),.clk(gclk));
	jnot g12817(.din(n13098),.dout(n13099),.clk(gclk));
	jand g12818(.dina(n13099),.dinb(n13097),.dout(n13100),.clk(gclk));
	jnot g12819(.din(n13100),.dout(n13101),.clk(gclk));
	jor g12820(.dina(w_n13101_0[1]),.dinb(w_n13093_0[1]),.dout(n13102),.clk(gclk));
	jand g12821(.dina(n13102),.dinb(w_n13091_0[1]),.dout(n13103),.clk(gclk));
	jor g12822(.dina(w_n13103_0[1]),.dinb(w_n425_18[0]),.dout(n13104),.clk(gclk));
	jxor g12823(.dina(w_n12579_0[0]),.dinb(w_n430_18[2]),.dout(n13105),.clk(gclk));
	jor g12824(.dina(n13105),.dinb(w_n12675_15[2]),.dout(n13106),.clk(gclk));
	jxor g12825(.dina(n13106),.dinb(w_n12590_0[0]),.dout(n13107),.clk(gclk));
	jand g12826(.dina(w_n13103_0[0]),.dinb(w_n425_17[2]),.dout(n13108),.clk(gclk));
	jor g12827(.dina(w_n13108_0[1]),.dinb(w_n13107_0[1]),.dout(n13109),.clk(gclk));
	jand g12828(.dina(w_n13109_0[2]),.dinb(w_n13104_0[2]),.dout(n13110),.clk(gclk));
	jor g12829(.dina(n13110),.dinb(w_n305_19[2]),.dout(n13111),.clk(gclk));
	jnot g12830(.din(w_n12595_0[0]),.dout(n13112),.clk(gclk));
	jor g12831(.dina(n13112),.dinb(w_n12593_0[0]),.dout(n13113),.clk(gclk));
	jor g12832(.dina(n13113),.dinb(w_n12675_15[1]),.dout(n13114),.clk(gclk));
	jxor g12833(.dina(n13114),.dinb(w_n12604_0[0]),.dout(n13115),.clk(gclk));
	jand g12834(.dina(w_n13104_0[1]),.dinb(w_n305_19[1]),.dout(n13116),.clk(gclk));
	jand g12835(.dina(n13116),.dinb(w_n13109_0[1]),.dout(n13117),.clk(gclk));
	jor g12836(.dina(w_n13117_0[1]),.dinb(w_n13115_0[1]),.dout(n13118),.clk(gclk));
	jand g12837(.dina(w_n13118_0[1]),.dinb(w_n13111_0[1]),.dout(n13119),.clk(gclk));
	jor g12838(.dina(w_n13119_0[2]),.dinb(w_n290_19[1]),.dout(n13120),.clk(gclk));
	jand g12839(.dina(w_n13119_0[1]),.dinb(w_n290_19[0]),.dout(n13121),.clk(gclk));
	jnot g12840(.din(w_n12607_0[0]),.dout(n13122),.clk(gclk));
	jand g12841(.dina(w_asqrt15_11[1]),.dinb(n13122),.dout(n13123),.clk(gclk));
	jand g12842(.dina(w_n13123_0[1]),.dinb(w_n12612_0[0]),.dout(n13124),.clk(gclk));
	jor g12843(.dina(n13124),.dinb(w_n12611_0[0]),.dout(n13125),.clk(gclk));
	jand g12844(.dina(w_n13123_0[0]),.dinb(w_n12613_0[0]),.dout(n13126),.clk(gclk));
	jnot g12845(.din(n13126),.dout(n13127),.clk(gclk));
	jand g12846(.dina(n13127),.dinb(n13125),.dout(n13128),.clk(gclk));
	jnot g12847(.din(n13128),.dout(n13129),.clk(gclk));
	jor g12848(.dina(w_n13129_0[1]),.dinb(n13121),.dout(n13130),.clk(gclk));
	jand g12849(.dina(w_n13130_0[1]),.dinb(w_n13120_0[1]),.dout(n13131),.clk(gclk));
	jor g12850(.dina(n13131),.dinb(w_n223_19[2]),.dout(n13132),.clk(gclk));
	jand g12851(.dina(w_n13120_0[0]),.dinb(w_n223_19[1]),.dout(n13133),.clk(gclk));
	jand g12852(.dina(n13133),.dinb(w_n13130_0[0]),.dout(n13134),.clk(gclk));
	jnot g12853(.din(w_n12615_0[0]),.dout(n13135),.clk(gclk));
	jand g12854(.dina(w_asqrt15_11[0]),.dinb(n13135),.dout(n13136),.clk(gclk));
	jand g12855(.dina(w_n13136_0[1]),.dinb(w_n12622_0[0]),.dout(n13137),.clk(gclk));
	jor g12856(.dina(n13137),.dinb(w_n12620_0[0]),.dout(n13138),.clk(gclk));
	jand g12857(.dina(w_n13136_0[0]),.dinb(w_n12623_0[0]),.dout(n13139),.clk(gclk));
	jnot g12858(.din(n13139),.dout(n13140),.clk(gclk));
	jand g12859(.dina(n13140),.dinb(n13138),.dout(n13141),.clk(gclk));
	jnot g12860(.din(n13141),.dout(n13142),.clk(gclk));
	jor g12861(.dina(w_n13142_0[1]),.dinb(w_n13134_0[1]),.dout(n13143),.clk(gclk));
	jand g12862(.dina(n13143),.dinb(w_n13132_0[1]),.dout(n13144),.clk(gclk));
	jor g12863(.dina(w_n13144_0[2]),.dinb(w_n199_22[1]),.dout(n13145),.clk(gclk));
	jand g12864(.dina(w_n13144_0[1]),.dinb(w_n199_22[0]),.dout(n13146),.clk(gclk));
	jxor g12865(.dina(w_n12624_0[0]),.dinb(w_n223_19[0]),.dout(n13147),.clk(gclk));
	jor g12866(.dina(n13147),.dinb(w_n12675_15[0]),.dout(n13148),.clk(gclk));
	jxor g12867(.dina(n13148),.dinb(w_n12635_0[0]),.dout(n13149),.clk(gclk));
	jor g12868(.dina(w_n13149_0[1]),.dinb(n13146),.dout(n13150),.clk(gclk));
	jand g12869(.dina(n13150),.dinb(n13145),.dout(n13151),.clk(gclk));
	jnot g12870(.din(w_n12640_0[0]),.dout(n13152),.clk(gclk));
	jor g12871(.dina(n13152),.dinb(w_n12638_0[0]),.dout(n13153),.clk(gclk));
	jor g12872(.dina(n13153),.dinb(w_n12675_14[2]),.dout(n13154),.clk(gclk));
	jxor g12873(.dina(n13154),.dinb(w_n12649_0[0]),.dout(n13155),.clk(gclk));
	jand g12874(.dina(w_asqrt15_10[2]),.dinb(w_n12663_0[1]),.dout(n13156),.clk(gclk));
	jand g12875(.dina(w_n13156_0[1]),.dinb(w_n12651_1[0]),.dout(n13157),.clk(gclk));
	jor g12876(.dina(n13157),.dinb(w_n12698_0[0]),.dout(n13158),.clk(gclk));
	jor g12877(.dina(n13158),.dinb(w_n13155_0[2]),.dout(n13159),.clk(gclk));
	jor g12878(.dina(n13159),.dinb(w_n13151_0[2]),.dout(n13160),.clk(gclk));
	jand g12879(.dina(n13160),.dinb(w_n194_21[1]),.dout(n13161),.clk(gclk));
	jand g12880(.dina(w_n13155_0[1]),.dinb(w_n13151_0[1]),.dout(n13162),.clk(gclk));
	jor g12881(.dina(w_n13156_0[0]),.dinb(w_n12651_0[2]),.dout(n13163),.clk(gclk));
	jand g12882(.dina(w_n12663_0[0]),.dinb(w_n12651_0[1]),.dout(n13164),.clk(gclk));
	jor g12883(.dina(n13164),.dinb(w_n194_21[0]),.dout(n13165),.clk(gclk));
	jnot g12884(.din(n13165),.dout(n13166),.clk(gclk));
	jand g12885(.dina(n13166),.dinb(n13163),.dout(n13167),.clk(gclk));
	jor g12886(.dina(w_n13167_0[1]),.dinb(w_n13162_0[2]),.dout(n13170),.clk(gclk));
	jor g12887(.dina(n13170),.dinb(w_n13161_0[1]),.dout(asqrt_fa_15),.clk(gclk));
	jxor g12888(.dina(w_n13008_0[0]),.dinb(w_n1641_15[2]),.dout(n13172),.clk(gclk));
	jand g12889(.dina(n13172),.dinb(w_asqrt14_31),.dout(n13173),.clk(gclk));
	jxor g12890(.dina(n13173),.dinb(w_n12679_0[0]),.dout(n13174),.clk(gclk));
	jnot g12891(.din(n13174),.dout(n13175),.clk(gclk));
	jand g12892(.dina(w_asqrt14_30[2]),.dinb(w_a28_0[0]),.dout(n13176),.clk(gclk));
	jnot g12893(.din(w_a26_0[1]),.dout(n13177),.clk(gclk));
	jnot g12894(.din(w_a27_0[1]),.dout(n13178),.clk(gclk));
	jand g12895(.dina(w_n12681_1[0]),.dinb(w_n13178_0[1]),.dout(n13179),.clk(gclk));
	jand g12896(.dina(n13179),.dinb(w_n13177_1[1]),.dout(n13180),.clk(gclk));
	jor g12897(.dina(n13180),.dinb(n13176),.dout(n13181),.clk(gclk));
	jand g12898(.dina(w_n13181_0[2]),.dinb(w_asqrt15_10[1]),.dout(n13182),.clk(gclk));
	jand g12899(.dina(w_asqrt14_30[1]),.dinb(w_n12681_0[2]),.dout(n13183),.clk(gclk));
	jxor g12900(.dina(w_n13183_0[1]),.dinb(w_n12682_0[1]),.dout(n13184),.clk(gclk));
	jor g12901(.dina(w_n13181_0[1]),.dinb(w_asqrt15_10[0]),.dout(n13185),.clk(gclk));
	jand g12902(.dina(n13185),.dinb(w_n13184_0[1]),.dout(n13186),.clk(gclk));
	jor g12903(.dina(w_n13186_0[1]),.dinb(w_n13182_0[1]),.dout(n13187),.clk(gclk));
	jand g12904(.dina(n13187),.dinb(w_asqrt16_14[2]),.dout(n13188),.clk(gclk));
	jor g12905(.dina(w_n13182_0[0]),.dinb(w_asqrt16_14[1]),.dout(n13189),.clk(gclk));
	jor g12906(.dina(n13189),.dinb(w_n13186_0[0]),.dout(n13190),.clk(gclk));
	jand g12907(.dina(w_n13183_0[0]),.dinb(w_n12682_0[0]),.dout(n13191),.clk(gclk));
	jnot g12908(.din(w_n13161_0[0]),.dout(n13192),.clk(gclk));
	jnot g12909(.din(w_n13162_0[1]),.dout(n13193),.clk(gclk));
	jnot g12910(.din(w_n13167_0[0]),.dout(n13194),.clk(gclk));
	jand g12911(.dina(n13194),.dinb(w_asqrt15_9[2]),.dout(n13195),.clk(gclk));
	jand g12912(.dina(n13195),.dinb(n13193),.dout(n13196),.clk(gclk));
	jand g12913(.dina(n13196),.dinb(n13192),.dout(n13197),.clk(gclk));
	jor g12914(.dina(n13197),.dinb(n13191),.dout(n13198),.clk(gclk));
	jxor g12915(.dina(n13198),.dinb(w_n12148_0[1]),.dout(n13199),.clk(gclk));
	jand g12916(.dina(w_n13199_0[1]),.dinb(w_n13190_0[1]),.dout(n13200),.clk(gclk));
	jor g12917(.dina(n13200),.dinb(w_n13188_0[1]),.dout(n13201),.clk(gclk));
	jand g12918(.dina(w_n13201_0[2]),.dinb(w_asqrt17_10[1]),.dout(n13202),.clk(gclk));
	jor g12919(.dina(w_n13201_0[1]),.dinb(w_asqrt17_10[0]),.dout(n13203),.clk(gclk));
	jxor g12920(.dina(w_n12686_0[0]),.dinb(w_n12670_9[2]),.dout(n13204),.clk(gclk));
	jand g12921(.dina(n13204),.dinb(w_asqrt14_30[0]),.dout(n13205),.clk(gclk));
	jxor g12922(.dina(n13205),.dinb(w_n12689_0[0]),.dout(n13206),.clk(gclk));
	jnot g12923(.din(w_n13206_0[1]),.dout(n13207),.clk(gclk));
	jand g12924(.dina(n13207),.dinb(n13203),.dout(n13208),.clk(gclk));
	jor g12925(.dina(w_n13208_0[1]),.dinb(w_n13202_0[1]),.dout(n13209),.clk(gclk));
	jand g12926(.dina(n13209),.dinb(w_asqrt18_14[2]),.dout(n13210),.clk(gclk));
	jnot g12927(.din(w_n12695_0[0]),.dout(n13211),.clk(gclk));
	jand g12928(.dina(n13211),.dinb(w_n12693_0[0]),.dout(n13212),.clk(gclk));
	jand g12929(.dina(n13212),.dinb(w_asqrt14_29[2]),.dout(n13213),.clk(gclk));
	jxor g12930(.dina(n13213),.dinb(w_n12703_0[0]),.dout(n13214),.clk(gclk));
	jnot g12931(.din(n13214),.dout(n13215),.clk(gclk));
	jor g12932(.dina(w_n13202_0[0]),.dinb(w_asqrt18_14[1]),.dout(n13216),.clk(gclk));
	jor g12933(.dina(n13216),.dinb(w_n13208_0[0]),.dout(n13217),.clk(gclk));
	jand g12934(.dina(w_n13217_0[1]),.dinb(w_n13215_0[1]),.dout(n13218),.clk(gclk));
	jor g12935(.dina(w_n13218_0[1]),.dinb(w_n13210_0[1]),.dout(n13219),.clk(gclk));
	jand g12936(.dina(w_n13219_0[2]),.dinb(w_asqrt19_10[1]),.dout(n13220),.clk(gclk));
	jor g12937(.dina(w_n13219_0[1]),.dinb(w_asqrt19_10[0]),.dout(n13221),.clk(gclk));
	jnot g12938(.din(w_n12710_0[0]),.dout(n13222),.clk(gclk));
	jxor g12939(.dina(w_n12705_0[0]),.dinb(w_n11657_9[2]),.dout(n13223),.clk(gclk));
	jand g12940(.dina(n13223),.dinb(w_asqrt14_29[1]),.dout(n13224),.clk(gclk));
	jxor g12941(.dina(n13224),.dinb(n13222),.dout(n13225),.clk(gclk));
	jand g12942(.dina(w_n13225_0[1]),.dinb(n13221),.dout(n13226),.clk(gclk));
	jor g12943(.dina(w_n13226_0[1]),.dinb(w_n13220_0[1]),.dout(n13227),.clk(gclk));
	jand g12944(.dina(n13227),.dinb(w_asqrt20_14[2]),.dout(n13228),.clk(gclk));
	jor g12945(.dina(w_n13220_0[0]),.dinb(w_asqrt20_14[1]),.dout(n13229),.clk(gclk));
	jor g12946(.dina(n13229),.dinb(w_n13226_0[0]),.dout(n13230),.clk(gclk));
	jnot g12947(.din(w_n12717_0[0]),.dout(n13231),.clk(gclk));
	jnot g12948(.din(w_n12719_0[0]),.dout(n13232),.clk(gclk));
	jand g12949(.dina(w_asqrt14_29[0]),.dinb(w_n12713_0[0]),.dout(n13233),.clk(gclk));
	jand g12950(.dina(w_n13233_0[1]),.dinb(n13232),.dout(n13234),.clk(gclk));
	jor g12951(.dina(n13234),.dinb(n13231),.dout(n13235),.clk(gclk));
	jnot g12952(.din(w_n12720_0[0]),.dout(n13236),.clk(gclk));
	jand g12953(.dina(w_n13233_0[0]),.dinb(n13236),.dout(n13237),.clk(gclk));
	jnot g12954(.din(n13237),.dout(n13238),.clk(gclk));
	jand g12955(.dina(n13238),.dinb(n13235),.dout(n13239),.clk(gclk));
	jand g12956(.dina(w_n13239_0[1]),.dinb(w_n13230_0[1]),.dout(n13240),.clk(gclk));
	jor g12957(.dina(n13240),.dinb(w_n13228_0[1]),.dout(n13241),.clk(gclk));
	jand g12958(.dina(w_n13241_0[2]),.dinb(w_asqrt21_10[2]),.dout(n13242),.clk(gclk));
	jor g12959(.dina(w_n13241_0[1]),.dinb(w_asqrt21_10[1]),.dout(n13243),.clk(gclk));
	jxor g12960(.dina(w_n12721_0[0]),.dinb(w_n10696_10[1]),.dout(n13244),.clk(gclk));
	jand g12961(.dina(n13244),.dinb(w_asqrt14_28[2]),.dout(n13245),.clk(gclk));
	jxor g12962(.dina(n13245),.dinb(w_n12726_0[0]),.dout(n13246),.clk(gclk));
	jand g12963(.dina(w_n13246_0[1]),.dinb(n13243),.dout(n13247),.clk(gclk));
	jor g12964(.dina(w_n13247_0[1]),.dinb(w_n13242_0[1]),.dout(n13248),.clk(gclk));
	jand g12965(.dina(n13248),.dinb(w_asqrt22_14[2]),.dout(n13249),.clk(gclk));
	jnot g12966(.din(w_n12732_0[0]),.dout(n13250),.clk(gclk));
	jand g12967(.dina(n13250),.dinb(w_n12730_0[0]),.dout(n13251),.clk(gclk));
	jand g12968(.dina(n13251),.dinb(w_asqrt14_28[1]),.dout(n13252),.clk(gclk));
	jxor g12969(.dina(n13252),.dinb(w_n12741_0[0]),.dout(n13253),.clk(gclk));
	jnot g12970(.din(n13253),.dout(n13254),.clk(gclk));
	jor g12971(.dina(w_n13242_0[0]),.dinb(w_asqrt22_14[1]),.dout(n13255),.clk(gclk));
	jor g12972(.dina(n13255),.dinb(w_n13247_0[0]),.dout(n13256),.clk(gclk));
	jand g12973(.dina(w_n13256_0[1]),.dinb(w_n13254_0[1]),.dout(n13257),.clk(gclk));
	jor g12974(.dina(w_n13257_0[1]),.dinb(w_n13249_0[1]),.dout(n13258),.clk(gclk));
	jand g12975(.dina(w_n13258_0[2]),.dinb(w_asqrt23_10[2]),.dout(n13259),.clk(gclk));
	jor g12976(.dina(w_n13258_0[1]),.dinb(w_asqrt23_10[1]),.dout(n13260),.clk(gclk));
	jxor g12977(.dina(w_n12743_0[0]),.dinb(w_n9769_10[1]),.dout(n13261),.clk(gclk));
	jand g12978(.dina(n13261),.dinb(w_asqrt14_28[0]),.dout(n13262),.clk(gclk));
	jxor g12979(.dina(n13262),.dinb(w_n12749_0[0]),.dout(n13263),.clk(gclk));
	jand g12980(.dina(w_n13263_0[1]),.dinb(n13260),.dout(n13264),.clk(gclk));
	jor g12981(.dina(w_n13264_0[1]),.dinb(w_n13259_0[1]),.dout(n13265),.clk(gclk));
	jand g12982(.dina(n13265),.dinb(w_asqrt24_14[2]),.dout(n13266),.clk(gclk));
	jor g12983(.dina(w_n13259_0[0]),.dinb(w_asqrt24_14[1]),.dout(n13267),.clk(gclk));
	jor g12984(.dina(n13267),.dinb(w_n13264_0[0]),.dout(n13268),.clk(gclk));
	jnot g12985(.din(w_n12757_0[0]),.dout(n13269),.clk(gclk));
	jnot g12986(.din(w_n12759_0[0]),.dout(n13270),.clk(gclk));
	jand g12987(.dina(w_asqrt14_27[2]),.dinb(w_n12753_0[0]),.dout(n13271),.clk(gclk));
	jand g12988(.dina(w_n13271_0[1]),.dinb(n13270),.dout(n13272),.clk(gclk));
	jor g12989(.dina(n13272),.dinb(n13269),.dout(n13273),.clk(gclk));
	jnot g12990(.din(w_n12760_0[0]),.dout(n13274),.clk(gclk));
	jand g12991(.dina(w_n13271_0[0]),.dinb(n13274),.dout(n13275),.clk(gclk));
	jnot g12992(.din(n13275),.dout(n13276),.clk(gclk));
	jand g12993(.dina(n13276),.dinb(n13273),.dout(n13277),.clk(gclk));
	jand g12994(.dina(w_n13277_0[1]),.dinb(w_n13268_0[1]),.dout(n13278),.clk(gclk));
	jor g12995(.dina(n13278),.dinb(w_n13266_0[1]),.dout(n13279),.clk(gclk));
	jand g12996(.dina(w_n13279_0[1]),.dinb(w_asqrt25_11[0]),.dout(n13280),.clk(gclk));
	jxor g12997(.dina(w_n12761_0[0]),.dinb(w_n8893_10[2]),.dout(n13281),.clk(gclk));
	jand g12998(.dina(n13281),.dinb(w_asqrt14_27[1]),.dout(n13282),.clk(gclk));
	jxor g12999(.dina(n13282),.dinb(w_n12768_0[0]),.dout(n13283),.clk(gclk));
	jnot g13000(.din(n13283),.dout(n13284),.clk(gclk));
	jor g13001(.dina(w_n13279_0[0]),.dinb(w_asqrt25_10[2]),.dout(n13285),.clk(gclk));
	jand g13002(.dina(w_n13285_0[1]),.dinb(w_n13284_0[1]),.dout(n13286),.clk(gclk));
	jor g13003(.dina(w_n13286_0[2]),.dinb(w_n13280_0[2]),.dout(n13287),.clk(gclk));
	jand g13004(.dina(n13287),.dinb(w_asqrt26_14[2]),.dout(n13288),.clk(gclk));
	jnot g13005(.din(w_n12773_0[0]),.dout(n13289),.clk(gclk));
	jand g13006(.dina(n13289),.dinb(w_n12771_0[0]),.dout(n13290),.clk(gclk));
	jand g13007(.dina(n13290),.dinb(w_asqrt14_27[0]),.dout(n13291),.clk(gclk));
	jxor g13008(.dina(n13291),.dinb(w_n12781_0[0]),.dout(n13292),.clk(gclk));
	jnot g13009(.din(n13292),.dout(n13293),.clk(gclk));
	jor g13010(.dina(w_n13280_0[1]),.dinb(w_asqrt26_14[1]),.dout(n13294),.clk(gclk));
	jor g13011(.dina(n13294),.dinb(w_n13286_0[1]),.dout(n13295),.clk(gclk));
	jand g13012(.dina(w_n13295_0[1]),.dinb(w_n13293_0[1]),.dout(n13296),.clk(gclk));
	jor g13013(.dina(w_n13296_0[1]),.dinb(w_n13288_0[1]),.dout(n13297),.clk(gclk));
	jand g13014(.dina(w_n13297_0[2]),.dinb(w_asqrt27_11[0]),.dout(n13298),.clk(gclk));
	jor g13015(.dina(w_n13297_0[1]),.dinb(w_asqrt27_10[2]),.dout(n13299),.clk(gclk));
	jnot g13016(.din(w_n12787_0[0]),.dout(n13300),.clk(gclk));
	jnot g13017(.din(w_n12788_0[0]),.dout(n13301),.clk(gclk));
	jand g13018(.dina(w_asqrt14_26[2]),.dinb(w_n12784_0[0]),.dout(n13302),.clk(gclk));
	jand g13019(.dina(w_n13302_0[1]),.dinb(n13301),.dout(n13303),.clk(gclk));
	jor g13020(.dina(n13303),.dinb(n13300),.dout(n13304),.clk(gclk));
	jnot g13021(.din(w_n12789_0[0]),.dout(n13305),.clk(gclk));
	jand g13022(.dina(w_n13302_0[0]),.dinb(n13305),.dout(n13306),.clk(gclk));
	jnot g13023(.din(n13306),.dout(n13307),.clk(gclk));
	jand g13024(.dina(n13307),.dinb(n13304),.dout(n13308),.clk(gclk));
	jand g13025(.dina(w_n13308_0[1]),.dinb(n13299),.dout(n13309),.clk(gclk));
	jor g13026(.dina(w_n13309_0[1]),.dinb(w_n13298_0[1]),.dout(n13310),.clk(gclk));
	jand g13027(.dina(n13310),.dinb(w_asqrt28_14[2]),.dout(n13311),.clk(gclk));
	jor g13028(.dina(w_n13298_0[0]),.dinb(w_asqrt28_14[1]),.dout(n13312),.clk(gclk));
	jor g13029(.dina(n13312),.dinb(w_n13309_0[0]),.dout(n13313),.clk(gclk));
	jnot g13030(.din(w_n12795_0[0]),.dout(n13314),.clk(gclk));
	jnot g13031(.din(w_n12797_0[0]),.dout(n13315),.clk(gclk));
	jand g13032(.dina(w_asqrt14_26[1]),.dinb(w_n12791_0[0]),.dout(n13316),.clk(gclk));
	jand g13033(.dina(w_n13316_0[1]),.dinb(n13315),.dout(n13317),.clk(gclk));
	jor g13034(.dina(n13317),.dinb(n13314),.dout(n13318),.clk(gclk));
	jnot g13035(.din(w_n12798_0[0]),.dout(n13319),.clk(gclk));
	jand g13036(.dina(w_n13316_0[0]),.dinb(n13319),.dout(n13320),.clk(gclk));
	jnot g13037(.din(n13320),.dout(n13321),.clk(gclk));
	jand g13038(.dina(n13321),.dinb(n13318),.dout(n13322),.clk(gclk));
	jand g13039(.dina(w_n13322_0[1]),.dinb(w_n13313_0[1]),.dout(n13323),.clk(gclk));
	jor g13040(.dina(n13323),.dinb(w_n13311_0[1]),.dout(n13324),.clk(gclk));
	jand g13041(.dina(w_n13324_0[1]),.dinb(w_asqrt29_11[1]),.dout(n13325),.clk(gclk));
	jxor g13042(.dina(w_n12799_0[0]),.dinb(w_n7260_11[2]),.dout(n13326),.clk(gclk));
	jand g13043(.dina(n13326),.dinb(w_asqrt14_26[0]),.dout(n13327),.clk(gclk));
	jxor g13044(.dina(n13327),.dinb(w_n12809_0[0]),.dout(n13328),.clk(gclk));
	jnot g13045(.din(n13328),.dout(n13329),.clk(gclk));
	jor g13046(.dina(w_n13324_0[0]),.dinb(w_asqrt29_11[0]),.dout(n13330),.clk(gclk));
	jand g13047(.dina(w_n13330_0[1]),.dinb(w_n13329_0[1]),.dout(n13331),.clk(gclk));
	jor g13048(.dina(w_n13331_0[2]),.dinb(w_n13325_0[2]),.dout(n13332),.clk(gclk));
	jand g13049(.dina(n13332),.dinb(w_asqrt30_14[2]),.dout(n13333),.clk(gclk));
	jnot g13050(.din(w_n12814_0[0]),.dout(n13334),.clk(gclk));
	jand g13051(.dina(n13334),.dinb(w_n12812_0[0]),.dout(n13335),.clk(gclk));
	jand g13052(.dina(n13335),.dinb(w_asqrt14_25[2]),.dout(n13336),.clk(gclk));
	jxor g13053(.dina(n13336),.dinb(w_n12822_0[0]),.dout(n13337),.clk(gclk));
	jnot g13054(.din(n13337),.dout(n13338),.clk(gclk));
	jor g13055(.dina(w_n13325_0[1]),.dinb(w_asqrt30_14[1]),.dout(n13339),.clk(gclk));
	jor g13056(.dina(n13339),.dinb(w_n13331_0[1]),.dout(n13340),.clk(gclk));
	jand g13057(.dina(w_n13340_0[1]),.dinb(w_n13338_0[1]),.dout(n13341),.clk(gclk));
	jor g13058(.dina(w_n13341_0[1]),.dinb(w_n13333_0[1]),.dout(n13342),.clk(gclk));
	jand g13059(.dina(w_n13342_0[2]),.dinb(w_asqrt31_11[1]),.dout(n13343),.clk(gclk));
	jor g13060(.dina(w_n13342_0[1]),.dinb(w_asqrt31_11[0]),.dout(n13344),.clk(gclk));
	jnot g13061(.din(w_n12828_0[0]),.dout(n13345),.clk(gclk));
	jnot g13062(.din(w_n12829_0[0]),.dout(n13346),.clk(gclk));
	jand g13063(.dina(w_asqrt14_25[1]),.dinb(w_n12825_0[0]),.dout(n13347),.clk(gclk));
	jand g13064(.dina(w_n13347_0[1]),.dinb(n13346),.dout(n13348),.clk(gclk));
	jor g13065(.dina(n13348),.dinb(n13345),.dout(n13349),.clk(gclk));
	jnot g13066(.din(w_n12830_0[0]),.dout(n13350),.clk(gclk));
	jand g13067(.dina(w_n13347_0[0]),.dinb(n13350),.dout(n13351),.clk(gclk));
	jnot g13068(.din(n13351),.dout(n13352),.clk(gclk));
	jand g13069(.dina(n13352),.dinb(n13349),.dout(n13353),.clk(gclk));
	jand g13070(.dina(w_n13353_0[1]),.dinb(n13344),.dout(n13354),.clk(gclk));
	jor g13071(.dina(w_n13354_0[1]),.dinb(w_n13343_0[1]),.dout(n13355),.clk(gclk));
	jand g13072(.dina(n13355),.dinb(w_asqrt32_14[2]),.dout(n13356),.clk(gclk));
	jor g13073(.dina(w_n13343_0[0]),.dinb(w_asqrt32_14[1]),.dout(n13357),.clk(gclk));
	jor g13074(.dina(n13357),.dinb(w_n13354_0[0]),.dout(n13358),.clk(gclk));
	jnot g13075(.din(w_n12836_0[0]),.dout(n13359),.clk(gclk));
	jnot g13076(.din(w_n12838_0[0]),.dout(n13360),.clk(gclk));
	jand g13077(.dina(w_asqrt14_25[0]),.dinb(w_n12832_0[0]),.dout(n13361),.clk(gclk));
	jand g13078(.dina(w_n13361_0[1]),.dinb(n13360),.dout(n13362),.clk(gclk));
	jor g13079(.dina(n13362),.dinb(n13359),.dout(n13363),.clk(gclk));
	jnot g13080(.din(w_n12839_0[0]),.dout(n13364),.clk(gclk));
	jand g13081(.dina(w_n13361_0[0]),.dinb(n13364),.dout(n13365),.clk(gclk));
	jnot g13082(.din(n13365),.dout(n13366),.clk(gclk));
	jand g13083(.dina(n13366),.dinb(n13363),.dout(n13367),.clk(gclk));
	jand g13084(.dina(w_n13367_0[1]),.dinb(w_n13358_0[1]),.dout(n13368),.clk(gclk));
	jor g13085(.dina(n13368),.dinb(w_n13356_0[1]),.dout(n13369),.clk(gclk));
	jand g13086(.dina(w_n13369_0[1]),.dinb(w_asqrt33_11[2]),.dout(n13370),.clk(gclk));
	jxor g13087(.dina(w_n12840_0[0]),.dinb(w_n5788_12[1]),.dout(n13371),.clk(gclk));
	jand g13088(.dina(n13371),.dinb(w_asqrt14_24[2]),.dout(n13372),.clk(gclk));
	jxor g13089(.dina(n13372),.dinb(w_n12850_0[0]),.dout(n13373),.clk(gclk));
	jnot g13090(.din(n13373),.dout(n13374),.clk(gclk));
	jor g13091(.dina(w_n13369_0[0]),.dinb(w_asqrt33_11[1]),.dout(n13375),.clk(gclk));
	jand g13092(.dina(w_n13375_0[1]),.dinb(w_n13374_0[1]),.dout(n13376),.clk(gclk));
	jor g13093(.dina(w_n13376_0[2]),.dinb(w_n13370_0[2]),.dout(n13377),.clk(gclk));
	jand g13094(.dina(n13377),.dinb(w_asqrt34_14[2]),.dout(n13378),.clk(gclk));
	jnot g13095(.din(w_n12855_0[0]),.dout(n13379),.clk(gclk));
	jand g13096(.dina(n13379),.dinb(w_n12853_0[0]),.dout(n13380),.clk(gclk));
	jand g13097(.dina(n13380),.dinb(w_asqrt14_24[1]),.dout(n13381),.clk(gclk));
	jxor g13098(.dina(n13381),.dinb(w_n12863_0[0]),.dout(n13382),.clk(gclk));
	jnot g13099(.din(n13382),.dout(n13383),.clk(gclk));
	jor g13100(.dina(w_n13370_0[1]),.dinb(w_asqrt34_14[1]),.dout(n13384),.clk(gclk));
	jor g13101(.dina(n13384),.dinb(w_n13376_0[1]),.dout(n13385),.clk(gclk));
	jand g13102(.dina(w_n13385_0[1]),.dinb(w_n13383_0[1]),.dout(n13386),.clk(gclk));
	jor g13103(.dina(w_n13386_0[1]),.dinb(w_n13378_0[1]),.dout(n13387),.clk(gclk));
	jand g13104(.dina(w_n13387_0[2]),.dinb(w_asqrt35_11[2]),.dout(n13388),.clk(gclk));
	jor g13105(.dina(w_n13387_0[1]),.dinb(w_asqrt35_11[1]),.dout(n13389),.clk(gclk));
	jnot g13106(.din(w_n12869_0[0]),.dout(n13390),.clk(gclk));
	jnot g13107(.din(w_n12870_0[0]),.dout(n13391),.clk(gclk));
	jand g13108(.dina(w_asqrt14_24[0]),.dinb(w_n12866_0[0]),.dout(n13392),.clk(gclk));
	jand g13109(.dina(w_n13392_0[1]),.dinb(n13391),.dout(n13393),.clk(gclk));
	jor g13110(.dina(n13393),.dinb(n13390),.dout(n13394),.clk(gclk));
	jnot g13111(.din(w_n12871_0[0]),.dout(n13395),.clk(gclk));
	jand g13112(.dina(w_n13392_0[0]),.dinb(n13395),.dout(n13396),.clk(gclk));
	jnot g13113(.din(n13396),.dout(n13397),.clk(gclk));
	jand g13114(.dina(n13397),.dinb(n13394),.dout(n13398),.clk(gclk));
	jand g13115(.dina(w_n13398_0[1]),.dinb(n13389),.dout(n13399),.clk(gclk));
	jor g13116(.dina(w_n13399_0[1]),.dinb(w_n13388_0[1]),.dout(n13400),.clk(gclk));
	jand g13117(.dina(n13400),.dinb(w_asqrt36_14[2]),.dout(n13401),.clk(gclk));
	jor g13118(.dina(w_n13388_0[0]),.dinb(w_asqrt36_14[1]),.dout(n13402),.clk(gclk));
	jor g13119(.dina(n13402),.dinb(w_n13399_0[0]),.dout(n13403),.clk(gclk));
	jnot g13120(.din(w_n12877_0[0]),.dout(n13404),.clk(gclk));
	jnot g13121(.din(w_n12879_0[0]),.dout(n13405),.clk(gclk));
	jand g13122(.dina(w_asqrt14_23[2]),.dinb(w_n12873_0[0]),.dout(n13406),.clk(gclk));
	jand g13123(.dina(w_n13406_0[1]),.dinb(n13405),.dout(n13407),.clk(gclk));
	jor g13124(.dina(n13407),.dinb(n13404),.dout(n13408),.clk(gclk));
	jnot g13125(.din(w_n12880_0[0]),.dout(n13409),.clk(gclk));
	jand g13126(.dina(w_n13406_0[0]),.dinb(n13409),.dout(n13410),.clk(gclk));
	jnot g13127(.din(n13410),.dout(n13411),.clk(gclk));
	jand g13128(.dina(n13411),.dinb(n13408),.dout(n13412),.clk(gclk));
	jand g13129(.dina(w_n13412_0[1]),.dinb(w_n13403_0[1]),.dout(n13413),.clk(gclk));
	jor g13130(.dina(n13413),.dinb(w_n13401_0[1]),.dout(n13414),.clk(gclk));
	jand g13131(.dina(w_n13414_0[1]),.dinb(w_asqrt37_12[0]),.dout(n13415),.clk(gclk));
	jxor g13132(.dina(w_n12881_0[0]),.dinb(w_n4494_13[1]),.dout(n13416),.clk(gclk));
	jand g13133(.dina(n13416),.dinb(w_asqrt14_23[1]),.dout(n13417),.clk(gclk));
	jxor g13134(.dina(n13417),.dinb(w_n12891_0[0]),.dout(n13418),.clk(gclk));
	jnot g13135(.din(n13418),.dout(n13419),.clk(gclk));
	jor g13136(.dina(w_n13414_0[0]),.dinb(w_asqrt37_11[2]),.dout(n13420),.clk(gclk));
	jand g13137(.dina(w_n13420_0[1]),.dinb(w_n13419_0[1]),.dout(n13421),.clk(gclk));
	jor g13138(.dina(w_n13421_0[2]),.dinb(w_n13415_0[2]),.dout(n13422),.clk(gclk));
	jand g13139(.dina(n13422),.dinb(w_asqrt38_14[2]),.dout(n13423),.clk(gclk));
	jnot g13140(.din(w_n12896_0[0]),.dout(n13424),.clk(gclk));
	jand g13141(.dina(n13424),.dinb(w_n12894_0[0]),.dout(n13425),.clk(gclk));
	jand g13142(.dina(n13425),.dinb(w_asqrt14_23[0]),.dout(n13426),.clk(gclk));
	jxor g13143(.dina(n13426),.dinb(w_n12904_0[0]),.dout(n13427),.clk(gclk));
	jnot g13144(.din(n13427),.dout(n13428),.clk(gclk));
	jor g13145(.dina(w_n13415_0[1]),.dinb(w_asqrt38_14[1]),.dout(n13429),.clk(gclk));
	jor g13146(.dina(n13429),.dinb(w_n13421_0[1]),.dout(n13430),.clk(gclk));
	jand g13147(.dina(w_n13430_0[1]),.dinb(w_n13428_0[1]),.dout(n13431),.clk(gclk));
	jor g13148(.dina(w_n13431_0[1]),.dinb(w_n13423_0[1]),.dout(n13432),.clk(gclk));
	jand g13149(.dina(w_n13432_0[2]),.dinb(w_asqrt39_12[0]),.dout(n13433),.clk(gclk));
	jor g13150(.dina(w_n13432_0[1]),.dinb(w_asqrt39_11[2]),.dout(n13434),.clk(gclk));
	jnot g13151(.din(w_n12910_0[0]),.dout(n13435),.clk(gclk));
	jnot g13152(.din(w_n12911_0[0]),.dout(n13436),.clk(gclk));
	jand g13153(.dina(w_asqrt14_22[2]),.dinb(w_n12907_0[0]),.dout(n13437),.clk(gclk));
	jand g13154(.dina(w_n13437_0[1]),.dinb(n13436),.dout(n13438),.clk(gclk));
	jor g13155(.dina(n13438),.dinb(n13435),.dout(n13439),.clk(gclk));
	jnot g13156(.din(w_n12912_0[0]),.dout(n13440),.clk(gclk));
	jand g13157(.dina(w_n13437_0[0]),.dinb(n13440),.dout(n13441),.clk(gclk));
	jnot g13158(.din(n13441),.dout(n13442),.clk(gclk));
	jand g13159(.dina(n13442),.dinb(n13439),.dout(n13443),.clk(gclk));
	jand g13160(.dina(w_n13443_0[1]),.dinb(n13434),.dout(n13444),.clk(gclk));
	jor g13161(.dina(w_n13444_0[1]),.dinb(w_n13433_0[1]),.dout(n13445),.clk(gclk));
	jand g13162(.dina(n13445),.dinb(w_asqrt40_14[2]),.dout(n13446),.clk(gclk));
	jor g13163(.dina(w_n13433_0[0]),.dinb(w_asqrt40_14[1]),.dout(n13447),.clk(gclk));
	jor g13164(.dina(n13447),.dinb(w_n13444_0[0]),.dout(n13448),.clk(gclk));
	jnot g13165(.din(w_n12918_0[0]),.dout(n13449),.clk(gclk));
	jnot g13166(.din(w_n12920_0[0]),.dout(n13450),.clk(gclk));
	jand g13167(.dina(w_asqrt14_22[1]),.dinb(w_n12914_0[0]),.dout(n13451),.clk(gclk));
	jand g13168(.dina(w_n13451_0[1]),.dinb(n13450),.dout(n13452),.clk(gclk));
	jor g13169(.dina(n13452),.dinb(n13449),.dout(n13453),.clk(gclk));
	jnot g13170(.din(w_n12921_0[0]),.dout(n13454),.clk(gclk));
	jand g13171(.dina(w_n13451_0[0]),.dinb(n13454),.dout(n13455),.clk(gclk));
	jnot g13172(.din(n13455),.dout(n13456),.clk(gclk));
	jand g13173(.dina(n13456),.dinb(n13453),.dout(n13457),.clk(gclk));
	jand g13174(.dina(w_n13457_0[1]),.dinb(w_n13448_0[1]),.dout(n13458),.clk(gclk));
	jor g13175(.dina(n13458),.dinb(w_n13446_0[1]),.dout(n13459),.clk(gclk));
	jand g13176(.dina(w_n13459_0[1]),.dinb(w_asqrt41_12[1]),.dout(n13460),.clk(gclk));
	jxor g13177(.dina(w_n12922_0[0]),.dinb(w_n3371_14[0]),.dout(n13461),.clk(gclk));
	jand g13178(.dina(n13461),.dinb(w_asqrt14_22[0]),.dout(n13462),.clk(gclk));
	jxor g13179(.dina(n13462),.dinb(w_n12932_0[0]),.dout(n13463),.clk(gclk));
	jnot g13180(.din(n13463),.dout(n13464),.clk(gclk));
	jor g13181(.dina(w_n13459_0[0]),.dinb(w_asqrt41_12[0]),.dout(n13465),.clk(gclk));
	jand g13182(.dina(w_n13465_0[1]),.dinb(w_n13464_0[1]),.dout(n13466),.clk(gclk));
	jor g13183(.dina(w_n13466_0[2]),.dinb(w_n13460_0[2]),.dout(n13467),.clk(gclk));
	jand g13184(.dina(n13467),.dinb(w_asqrt42_14[2]),.dout(n13468),.clk(gclk));
	jnot g13185(.din(w_n12937_0[0]),.dout(n13469),.clk(gclk));
	jand g13186(.dina(n13469),.dinb(w_n12935_0[0]),.dout(n13470),.clk(gclk));
	jand g13187(.dina(n13470),.dinb(w_asqrt14_21[2]),.dout(n13471),.clk(gclk));
	jxor g13188(.dina(n13471),.dinb(w_n12945_0[0]),.dout(n13472),.clk(gclk));
	jnot g13189(.din(n13472),.dout(n13473),.clk(gclk));
	jor g13190(.dina(w_n13460_0[1]),.dinb(w_asqrt42_14[1]),.dout(n13474),.clk(gclk));
	jor g13191(.dina(n13474),.dinb(w_n13466_0[1]),.dout(n13475),.clk(gclk));
	jand g13192(.dina(w_n13475_0[1]),.dinb(w_n13473_0[1]),.dout(n13476),.clk(gclk));
	jor g13193(.dina(w_n13476_0[1]),.dinb(w_n13468_0[1]),.dout(n13477),.clk(gclk));
	jand g13194(.dina(w_n13477_0[2]),.dinb(w_asqrt43_12[1]),.dout(n13478),.clk(gclk));
	jor g13195(.dina(w_n13477_0[1]),.dinb(w_asqrt43_12[0]),.dout(n13479),.clk(gclk));
	jnot g13196(.din(w_n12951_0[0]),.dout(n13480),.clk(gclk));
	jnot g13197(.din(w_n12952_0[0]),.dout(n13481),.clk(gclk));
	jand g13198(.dina(w_asqrt14_21[1]),.dinb(w_n12948_0[0]),.dout(n13482),.clk(gclk));
	jand g13199(.dina(w_n13482_0[1]),.dinb(n13481),.dout(n13483),.clk(gclk));
	jor g13200(.dina(n13483),.dinb(n13480),.dout(n13484),.clk(gclk));
	jnot g13201(.din(w_n12953_0[0]),.dout(n13485),.clk(gclk));
	jand g13202(.dina(w_n13482_0[0]),.dinb(n13485),.dout(n13486),.clk(gclk));
	jnot g13203(.din(n13486),.dout(n13487),.clk(gclk));
	jand g13204(.dina(n13487),.dinb(n13484),.dout(n13488),.clk(gclk));
	jand g13205(.dina(w_n13488_0[1]),.dinb(n13479),.dout(n13489),.clk(gclk));
	jor g13206(.dina(w_n13489_0[1]),.dinb(w_n13478_0[1]),.dout(n13490),.clk(gclk));
	jand g13207(.dina(n13490),.dinb(w_asqrt44_14[2]),.dout(n13491),.clk(gclk));
	jor g13208(.dina(w_n13478_0[0]),.dinb(w_asqrt44_14[1]),.dout(n13492),.clk(gclk));
	jor g13209(.dina(n13492),.dinb(w_n13489_0[0]),.dout(n13493),.clk(gclk));
	jnot g13210(.din(w_n12959_0[0]),.dout(n13494),.clk(gclk));
	jnot g13211(.din(w_n12961_0[0]),.dout(n13495),.clk(gclk));
	jand g13212(.dina(w_asqrt14_21[0]),.dinb(w_n12955_0[0]),.dout(n13496),.clk(gclk));
	jand g13213(.dina(w_n13496_0[1]),.dinb(n13495),.dout(n13497),.clk(gclk));
	jor g13214(.dina(n13497),.dinb(n13494),.dout(n13498),.clk(gclk));
	jnot g13215(.din(w_n12962_0[0]),.dout(n13499),.clk(gclk));
	jand g13216(.dina(w_n13496_0[0]),.dinb(n13499),.dout(n13500),.clk(gclk));
	jnot g13217(.din(n13500),.dout(n13501),.clk(gclk));
	jand g13218(.dina(n13501),.dinb(n13498),.dout(n13502),.clk(gclk));
	jand g13219(.dina(w_n13502_0[1]),.dinb(w_n13493_0[1]),.dout(n13503),.clk(gclk));
	jor g13220(.dina(n13503),.dinb(w_n13491_0[1]),.dout(n13504),.clk(gclk));
	jand g13221(.dina(w_n13504_0[1]),.dinb(w_asqrt45_12[2]),.dout(n13505),.clk(gclk));
	jxor g13222(.dina(w_n12963_0[0]),.dinb(w_n2420_15[0]),.dout(n13506),.clk(gclk));
	jand g13223(.dina(n13506),.dinb(w_asqrt14_20[2]),.dout(n13507),.clk(gclk));
	jxor g13224(.dina(n13507),.dinb(w_n12973_0[0]),.dout(n13508),.clk(gclk));
	jnot g13225(.din(n13508),.dout(n13509),.clk(gclk));
	jor g13226(.dina(w_n13504_0[0]),.dinb(w_asqrt45_12[1]),.dout(n13510),.clk(gclk));
	jand g13227(.dina(w_n13510_0[1]),.dinb(w_n13509_0[1]),.dout(n13511),.clk(gclk));
	jor g13228(.dina(w_n13511_0[2]),.dinb(w_n13505_0[2]),.dout(n13512),.clk(gclk));
	jand g13229(.dina(n13512),.dinb(w_asqrt46_14[2]),.dout(n13513),.clk(gclk));
	jnot g13230(.din(w_n12978_0[0]),.dout(n13514),.clk(gclk));
	jand g13231(.dina(n13514),.dinb(w_n12976_0[0]),.dout(n13515),.clk(gclk));
	jand g13232(.dina(n13515),.dinb(w_asqrt14_20[1]),.dout(n13516),.clk(gclk));
	jxor g13233(.dina(n13516),.dinb(w_n12986_0[0]),.dout(n13517),.clk(gclk));
	jnot g13234(.din(n13517),.dout(n13518),.clk(gclk));
	jor g13235(.dina(w_n13505_0[1]),.dinb(w_asqrt46_14[1]),.dout(n13519),.clk(gclk));
	jor g13236(.dina(n13519),.dinb(w_n13511_0[1]),.dout(n13520),.clk(gclk));
	jand g13237(.dina(w_n13520_0[1]),.dinb(w_n13518_0[1]),.dout(n13521),.clk(gclk));
	jor g13238(.dina(w_n13521_0[1]),.dinb(w_n13513_0[1]),.dout(n13522),.clk(gclk));
	jand g13239(.dina(w_n13522_0[2]),.dinb(w_asqrt47_12[2]),.dout(n13523),.clk(gclk));
	jor g13240(.dina(w_n13522_0[1]),.dinb(w_asqrt47_12[1]),.dout(n13524),.clk(gclk));
	jnot g13241(.din(w_n12992_0[0]),.dout(n13525),.clk(gclk));
	jnot g13242(.din(w_n12993_0[0]),.dout(n13526),.clk(gclk));
	jand g13243(.dina(w_asqrt14_20[0]),.dinb(w_n12989_0[0]),.dout(n13527),.clk(gclk));
	jand g13244(.dina(w_n13527_0[1]),.dinb(n13526),.dout(n13528),.clk(gclk));
	jor g13245(.dina(n13528),.dinb(n13525),.dout(n13529),.clk(gclk));
	jnot g13246(.din(w_n12994_0[0]),.dout(n13530),.clk(gclk));
	jand g13247(.dina(w_n13527_0[0]),.dinb(n13530),.dout(n13531),.clk(gclk));
	jnot g13248(.din(n13531),.dout(n13532),.clk(gclk));
	jand g13249(.dina(n13532),.dinb(n13529),.dout(n13533),.clk(gclk));
	jand g13250(.dina(w_n13533_0[1]),.dinb(n13524),.dout(n13534),.clk(gclk));
	jor g13251(.dina(w_n13534_0[1]),.dinb(w_n13523_0[1]),.dout(n13535),.clk(gclk));
	jand g13252(.dina(n13535),.dinb(w_asqrt48_14[2]),.dout(n13536),.clk(gclk));
	jnot g13253(.din(w_n12998_0[0]),.dout(n13537),.clk(gclk));
	jand g13254(.dina(n13537),.dinb(w_n12996_0[0]),.dout(n13538),.clk(gclk));
	jand g13255(.dina(n13538),.dinb(w_asqrt14_19[2]),.dout(n13539),.clk(gclk));
	jxor g13256(.dina(n13539),.dinb(w_n13006_0[0]),.dout(n13540),.clk(gclk));
	jnot g13257(.din(n13540),.dout(n13541),.clk(gclk));
	jor g13258(.dina(w_n13523_0[0]),.dinb(w_asqrt48_14[1]),.dout(n13542),.clk(gclk));
	jor g13259(.dina(n13542),.dinb(w_n13534_0[0]),.dout(n13543),.clk(gclk));
	jand g13260(.dina(w_n13543_0[1]),.dinb(w_n13541_0[1]),.dout(n13544),.clk(gclk));
	jor g13261(.dina(w_n13544_0[1]),.dinb(w_n13536_0[1]),.dout(n13545),.clk(gclk));
	jand g13262(.dina(w_n13545_0[2]),.dinb(w_asqrt49_13[0]),.dout(n13546),.clk(gclk));
	jor g13263(.dina(w_n13545_0[1]),.dinb(w_asqrt49_12[2]),.dout(n13547),.clk(gclk));
	jand g13264(.dina(n13547),.dinb(w_n13175_0[1]),.dout(n13548),.clk(gclk));
	jor g13265(.dina(w_n13548_0[1]),.dinb(w_n13546_0[1]),.dout(n13549),.clk(gclk));
	jand g13266(.dina(n13549),.dinb(w_asqrt50_14[2]),.dout(n13550),.clk(gclk));
	jor g13267(.dina(w_n13546_0[0]),.dinb(w_asqrt50_14[1]),.dout(n13551),.clk(gclk));
	jor g13268(.dina(n13551),.dinb(w_n13548_0[0]),.dout(n13552),.clk(gclk));
	jnot g13269(.din(w_n13017_0[0]),.dout(n13553),.clk(gclk));
	jnot g13270(.din(w_n13019_0[0]),.dout(n13554),.clk(gclk));
	jand g13271(.dina(w_asqrt14_19[1]),.dinb(w_n13013_0[0]),.dout(n13555),.clk(gclk));
	jand g13272(.dina(w_n13555_0[1]),.dinb(n13554),.dout(n13556),.clk(gclk));
	jor g13273(.dina(n13556),.dinb(n13553),.dout(n13557),.clk(gclk));
	jnot g13274(.din(w_n13020_0[0]),.dout(n13558),.clk(gclk));
	jand g13275(.dina(w_n13555_0[0]),.dinb(n13558),.dout(n13559),.clk(gclk));
	jnot g13276(.din(n13559),.dout(n13560),.clk(gclk));
	jand g13277(.dina(n13560),.dinb(n13557),.dout(n13561),.clk(gclk));
	jand g13278(.dina(w_n13561_0[1]),.dinb(w_n13552_0[1]),.dout(n13562),.clk(gclk));
	jor g13279(.dina(n13562),.dinb(w_n13550_0[1]),.dout(n13563),.clk(gclk));
	jand g13280(.dina(w_n13563_0[2]),.dinb(w_asqrt51_13[0]),.dout(n13564),.clk(gclk));
	jor g13281(.dina(w_n13563_0[1]),.dinb(w_asqrt51_12[2]),.dout(n13565),.clk(gclk));
	jnot g13282(.din(w_n13025_0[0]),.dout(n13566),.clk(gclk));
	jnot g13283(.din(w_n13026_0[0]),.dout(n13567),.clk(gclk));
	jand g13284(.dina(w_asqrt14_19[0]),.dinb(w_n13022_0[0]),.dout(n13568),.clk(gclk));
	jand g13285(.dina(w_n13568_0[1]),.dinb(n13567),.dout(n13569),.clk(gclk));
	jor g13286(.dina(n13569),.dinb(n13566),.dout(n13570),.clk(gclk));
	jnot g13287(.din(w_n13027_0[0]),.dout(n13571),.clk(gclk));
	jand g13288(.dina(w_n13568_0[0]),.dinb(n13571),.dout(n13572),.clk(gclk));
	jnot g13289(.din(n13572),.dout(n13573),.clk(gclk));
	jand g13290(.dina(n13573),.dinb(n13570),.dout(n13574),.clk(gclk));
	jand g13291(.dina(w_n13574_0[1]),.dinb(n13565),.dout(n13575),.clk(gclk));
	jor g13292(.dina(w_n13575_0[1]),.dinb(w_n13564_0[1]),.dout(n13576),.clk(gclk));
	jand g13293(.dina(n13576),.dinb(w_asqrt52_14[2]),.dout(n13577),.clk(gclk));
	jor g13294(.dina(w_n13564_0[0]),.dinb(w_asqrt52_14[1]),.dout(n13578),.clk(gclk));
	jor g13295(.dina(n13578),.dinb(w_n13575_0[0]),.dout(n13579),.clk(gclk));
	jnot g13296(.din(w_n13033_0[0]),.dout(n13580),.clk(gclk));
	jnot g13297(.din(w_n13035_0[0]),.dout(n13581),.clk(gclk));
	jand g13298(.dina(w_asqrt14_18[2]),.dinb(w_n13029_0[0]),.dout(n13582),.clk(gclk));
	jand g13299(.dina(w_n13582_0[1]),.dinb(n13581),.dout(n13583),.clk(gclk));
	jor g13300(.dina(n13583),.dinb(n13580),.dout(n13584),.clk(gclk));
	jnot g13301(.din(w_n13036_0[0]),.dout(n13585),.clk(gclk));
	jand g13302(.dina(w_n13582_0[0]),.dinb(n13585),.dout(n13586),.clk(gclk));
	jnot g13303(.din(n13586),.dout(n13587),.clk(gclk));
	jand g13304(.dina(n13587),.dinb(n13584),.dout(n13588),.clk(gclk));
	jand g13305(.dina(w_n13588_0[1]),.dinb(w_n13579_0[1]),.dout(n13589),.clk(gclk));
	jor g13306(.dina(n13589),.dinb(w_n13577_0[1]),.dout(n13590),.clk(gclk));
	jand g13307(.dina(w_n13590_0[1]),.dinb(w_asqrt53_13[1]),.dout(n13591),.clk(gclk));
	jxor g13308(.dina(w_n13037_0[0]),.dinb(w_n1034_16[2]),.dout(n13592),.clk(gclk));
	jand g13309(.dina(n13592),.dinb(w_asqrt14_18[1]),.dout(n13593),.clk(gclk));
	jxor g13310(.dina(n13593),.dinb(w_n13047_0[0]),.dout(n13594),.clk(gclk));
	jnot g13311(.din(n13594),.dout(n13595),.clk(gclk));
	jor g13312(.dina(w_n13590_0[0]),.dinb(w_asqrt53_13[0]),.dout(n13596),.clk(gclk));
	jand g13313(.dina(w_n13596_0[1]),.dinb(w_n13595_0[1]),.dout(n13597),.clk(gclk));
	jor g13314(.dina(w_n13597_0[2]),.dinb(w_n13591_0[2]),.dout(n13598),.clk(gclk));
	jand g13315(.dina(n13598),.dinb(w_asqrt54_14[2]),.dout(n13599),.clk(gclk));
	jnot g13316(.din(w_n13052_0[0]),.dout(n13600),.clk(gclk));
	jand g13317(.dina(n13600),.dinb(w_n13050_0[0]),.dout(n13601),.clk(gclk));
	jand g13318(.dina(n13601),.dinb(w_asqrt14_18[0]),.dout(n13602),.clk(gclk));
	jxor g13319(.dina(n13602),.dinb(w_n13060_0[0]),.dout(n13603),.clk(gclk));
	jnot g13320(.din(n13603),.dout(n13604),.clk(gclk));
	jor g13321(.dina(w_n13591_0[1]),.dinb(w_asqrt54_14[1]),.dout(n13605),.clk(gclk));
	jor g13322(.dina(n13605),.dinb(w_n13597_0[1]),.dout(n13606),.clk(gclk));
	jand g13323(.dina(w_n13606_0[1]),.dinb(w_n13604_0[1]),.dout(n13607),.clk(gclk));
	jor g13324(.dina(w_n13607_0[1]),.dinb(w_n13599_0[1]),.dout(n13608),.clk(gclk));
	jand g13325(.dina(w_n13608_0[2]),.dinb(w_asqrt55_13[2]),.dout(n13609),.clk(gclk));
	jor g13326(.dina(w_n13608_0[1]),.dinb(w_asqrt55_13[1]),.dout(n13610),.clk(gclk));
	jnot g13327(.din(w_n13066_0[0]),.dout(n13611),.clk(gclk));
	jnot g13328(.din(w_n13067_0[0]),.dout(n13612),.clk(gclk));
	jand g13329(.dina(w_asqrt14_17[2]),.dinb(w_n13063_0[0]),.dout(n13613),.clk(gclk));
	jand g13330(.dina(w_n13613_0[1]),.dinb(n13612),.dout(n13614),.clk(gclk));
	jor g13331(.dina(n13614),.dinb(n13611),.dout(n13615),.clk(gclk));
	jnot g13332(.din(w_n13068_0[0]),.dout(n13616),.clk(gclk));
	jand g13333(.dina(w_n13613_0[0]),.dinb(n13616),.dout(n13617),.clk(gclk));
	jnot g13334(.din(n13617),.dout(n13618),.clk(gclk));
	jand g13335(.dina(n13618),.dinb(n13615),.dout(n13619),.clk(gclk));
	jand g13336(.dina(w_n13619_0[1]),.dinb(n13610),.dout(n13620),.clk(gclk));
	jor g13337(.dina(w_n13620_0[1]),.dinb(w_n13609_0[1]),.dout(n13621),.clk(gclk));
	jand g13338(.dina(n13621),.dinb(w_asqrt56_14[2]),.dout(n13622),.clk(gclk));
	jor g13339(.dina(w_n13609_0[0]),.dinb(w_asqrt56_14[1]),.dout(n13623),.clk(gclk));
	jor g13340(.dina(n13623),.dinb(w_n13620_0[0]),.dout(n13624),.clk(gclk));
	jnot g13341(.din(w_n13074_0[0]),.dout(n13625),.clk(gclk));
	jnot g13342(.din(w_n13076_0[0]),.dout(n13626),.clk(gclk));
	jand g13343(.dina(w_asqrt14_17[1]),.dinb(w_n13070_0[0]),.dout(n13627),.clk(gclk));
	jand g13344(.dina(w_n13627_0[1]),.dinb(n13626),.dout(n13628),.clk(gclk));
	jor g13345(.dina(n13628),.dinb(n13625),.dout(n13629),.clk(gclk));
	jnot g13346(.din(w_n13077_0[0]),.dout(n13630),.clk(gclk));
	jand g13347(.dina(w_n13627_0[0]),.dinb(n13630),.dout(n13631),.clk(gclk));
	jnot g13348(.din(n13631),.dout(n13632),.clk(gclk));
	jand g13349(.dina(n13632),.dinb(n13629),.dout(n13633),.clk(gclk));
	jand g13350(.dina(w_n13633_0[1]),.dinb(w_n13624_0[1]),.dout(n13634),.clk(gclk));
	jor g13351(.dina(n13634),.dinb(w_n13622_0[1]),.dout(n13635),.clk(gclk));
	jand g13352(.dina(w_n13635_0[1]),.dinb(w_asqrt57_14[0]),.dout(n13636),.clk(gclk));
	jxor g13353(.dina(w_n13078_0[0]),.dinb(w_n590_17[1]),.dout(n13637),.clk(gclk));
	jand g13354(.dina(n13637),.dinb(w_asqrt14_17[0]),.dout(n13638),.clk(gclk));
	jxor g13355(.dina(n13638),.dinb(w_n13088_0[0]),.dout(n13639),.clk(gclk));
	jnot g13356(.din(n13639),.dout(n13640),.clk(gclk));
	jor g13357(.dina(w_n13635_0[0]),.dinb(w_asqrt57_13[2]),.dout(n13641),.clk(gclk));
	jand g13358(.dina(w_n13641_0[1]),.dinb(w_n13640_0[1]),.dout(n13642),.clk(gclk));
	jor g13359(.dina(w_n13642_0[2]),.dinb(w_n13636_0[2]),.dout(n13643),.clk(gclk));
	jand g13360(.dina(n13643),.dinb(w_asqrt58_14[2]),.dout(n13644),.clk(gclk));
	jnot g13361(.din(w_n13093_0[0]),.dout(n13645),.clk(gclk));
	jand g13362(.dina(n13645),.dinb(w_n13091_0[0]),.dout(n13646),.clk(gclk));
	jand g13363(.dina(n13646),.dinb(w_asqrt14_16[2]),.dout(n13647),.clk(gclk));
	jxor g13364(.dina(n13647),.dinb(w_n13101_0[0]),.dout(n13648),.clk(gclk));
	jnot g13365(.din(n13648),.dout(n13649),.clk(gclk));
	jor g13366(.dina(w_n13636_0[1]),.dinb(w_asqrt58_14[1]),.dout(n13650),.clk(gclk));
	jor g13367(.dina(n13650),.dinb(w_n13642_0[1]),.dout(n13651),.clk(gclk));
	jand g13368(.dina(w_n13651_0[1]),.dinb(w_n13649_0[1]),.dout(n13652),.clk(gclk));
	jor g13369(.dina(w_n13652_0[1]),.dinb(w_n13644_0[1]),.dout(n13653),.clk(gclk));
	jand g13370(.dina(w_n13653_0[2]),.dinb(w_asqrt59_14[1]),.dout(n13654),.clk(gclk));
	jor g13371(.dina(w_n13653_0[1]),.dinb(w_asqrt59_14[0]),.dout(n13655),.clk(gclk));
	jnot g13372(.din(w_n13107_0[0]),.dout(n13656),.clk(gclk));
	jnot g13373(.din(w_n13108_0[0]),.dout(n13657),.clk(gclk));
	jand g13374(.dina(w_asqrt14_16[1]),.dinb(w_n13104_0[0]),.dout(n13658),.clk(gclk));
	jand g13375(.dina(w_n13658_0[1]),.dinb(n13657),.dout(n13659),.clk(gclk));
	jor g13376(.dina(n13659),.dinb(n13656),.dout(n13660),.clk(gclk));
	jnot g13377(.din(w_n13109_0[0]),.dout(n13661),.clk(gclk));
	jand g13378(.dina(w_n13658_0[0]),.dinb(n13661),.dout(n13662),.clk(gclk));
	jnot g13379(.din(n13662),.dout(n13663),.clk(gclk));
	jand g13380(.dina(n13663),.dinb(n13660),.dout(n13664),.clk(gclk));
	jand g13381(.dina(w_n13664_0[1]),.dinb(n13655),.dout(n13665),.clk(gclk));
	jor g13382(.dina(w_n13665_0[1]),.dinb(w_n13654_0[1]),.dout(n13666),.clk(gclk));
	jand g13383(.dina(n13666),.dinb(w_asqrt60_14[1]),.dout(n13667),.clk(gclk));
	jor g13384(.dina(w_n13654_0[0]),.dinb(w_asqrt60_14[0]),.dout(n13668),.clk(gclk));
	jor g13385(.dina(n13668),.dinb(w_n13665_0[0]),.dout(n13669),.clk(gclk));
	jnot g13386(.din(w_n13115_0[0]),.dout(n13670),.clk(gclk));
	jnot g13387(.din(w_n13117_0[0]),.dout(n13671),.clk(gclk));
	jand g13388(.dina(w_asqrt14_16[0]),.dinb(w_n13111_0[0]),.dout(n13672),.clk(gclk));
	jand g13389(.dina(w_n13672_0[1]),.dinb(n13671),.dout(n13673),.clk(gclk));
	jor g13390(.dina(n13673),.dinb(n13670),.dout(n13674),.clk(gclk));
	jnot g13391(.din(w_n13118_0[0]),.dout(n13675),.clk(gclk));
	jand g13392(.dina(w_n13672_0[0]),.dinb(n13675),.dout(n13676),.clk(gclk));
	jnot g13393(.din(n13676),.dout(n13677),.clk(gclk));
	jand g13394(.dina(n13677),.dinb(n13674),.dout(n13678),.clk(gclk));
	jand g13395(.dina(w_n13678_0[1]),.dinb(w_n13669_0[1]),.dout(n13679),.clk(gclk));
	jor g13396(.dina(n13679),.dinb(w_n13667_0[1]),.dout(n13680),.clk(gclk));
	jand g13397(.dina(w_n13680_0[1]),.dinb(w_asqrt61_14[2]),.dout(n13681),.clk(gclk));
	jxor g13398(.dina(w_n13119_0[0]),.dinb(w_n290_18[2]),.dout(n13682),.clk(gclk));
	jand g13399(.dina(n13682),.dinb(w_asqrt14_15[2]),.dout(n13683),.clk(gclk));
	jxor g13400(.dina(n13683),.dinb(w_n13129_0[0]),.dout(n13684),.clk(gclk));
	jnot g13401(.din(n13684),.dout(n13685),.clk(gclk));
	jor g13402(.dina(w_n13680_0[0]),.dinb(w_asqrt61_14[1]),.dout(n13686),.clk(gclk));
	jand g13403(.dina(w_n13686_0[1]),.dinb(w_n13685_0[1]),.dout(n13687),.clk(gclk));
	jor g13404(.dina(w_n13687_0[2]),.dinb(w_n13681_0[2]),.dout(n13688),.clk(gclk));
	jand g13405(.dina(n13688),.dinb(w_asqrt62_14[2]),.dout(n13689),.clk(gclk));
	jnot g13406(.din(w_n13134_0[0]),.dout(n13690),.clk(gclk));
	jand g13407(.dina(n13690),.dinb(w_n13132_0[0]),.dout(n13691),.clk(gclk));
	jand g13408(.dina(n13691),.dinb(w_asqrt14_15[1]),.dout(n13692),.clk(gclk));
	jxor g13409(.dina(n13692),.dinb(w_n13142_0[0]),.dout(n13693),.clk(gclk));
	jnot g13410(.din(n13693),.dout(n13694),.clk(gclk));
	jor g13411(.dina(w_n13681_0[1]),.dinb(w_asqrt62_14[1]),.dout(n13695),.clk(gclk));
	jor g13412(.dina(n13695),.dinb(w_n13687_0[1]),.dout(n13696),.clk(gclk));
	jand g13413(.dina(w_n13696_0[1]),.dinb(w_n13694_0[1]),.dout(n13697),.clk(gclk));
	jor g13414(.dina(w_n13697_0[1]),.dinb(w_n13689_0[1]),.dout(n13698),.clk(gclk));
	jxor g13415(.dina(w_n13144_0[0]),.dinb(w_n199_21[2]),.dout(n13699),.clk(gclk));
	jand g13416(.dina(n13699),.dinb(w_asqrt14_15[0]),.dout(n13700),.clk(gclk));
	jxor g13417(.dina(n13700),.dinb(w_n13149_0[0]),.dout(n13701),.clk(gclk));
	jnot g13418(.din(w_n13151_0[0]),.dout(n13702),.clk(gclk));
	jnot g13419(.din(w_n13155_0[0]),.dout(n13703),.clk(gclk));
	jand g13420(.dina(w_asqrt14_14[2]),.dinb(w_n13703_0[1]),.dout(n13704),.clk(gclk));
	jand g13421(.dina(w_n13704_0[1]),.dinb(w_n13702_0[2]),.dout(n13705),.clk(gclk));
	jor g13422(.dina(n13705),.dinb(w_n13162_0[0]),.dout(n13706),.clk(gclk));
	jor g13423(.dina(n13706),.dinb(w_n13701_0[1]),.dout(n13707),.clk(gclk));
	jnot g13424(.din(n13707),.dout(n13708),.clk(gclk));
	jand g13425(.dina(n13708),.dinb(w_n13698_1[2]),.dout(n13709),.clk(gclk));
	jor g13426(.dina(n13709),.dinb(w_asqrt63_8[0]),.dout(n13710),.clk(gclk));
	jnot g13427(.din(w_n13701_0[0]),.dout(n13711),.clk(gclk));
	jor g13428(.dina(w_n13711_0[2]),.dinb(w_n13698_1[1]),.dout(n13712),.clk(gclk));
	jor g13429(.dina(w_n13704_0[0]),.dinb(w_n13702_0[1]),.dout(n13713),.clk(gclk));
	jand g13430(.dina(w_n13703_0[0]),.dinb(w_n13702_0[0]),.dout(n13714),.clk(gclk));
	jor g13431(.dina(n13714),.dinb(w_n194_20[2]),.dout(n13715),.clk(gclk));
	jnot g13432(.din(n13715),.dout(n13716),.clk(gclk));
	jand g13433(.dina(n13716),.dinb(n13713),.dout(n13717),.clk(gclk));
	jnot g13434(.din(w_asqrt14_14[1]),.dout(n13718),.clk(gclk));
	jnot g13435(.din(w_n13717_0[1]),.dout(n13721),.clk(gclk));
	jand g13436(.dina(n13721),.dinb(w_n13712_0[1]),.dout(n13722),.clk(gclk));
	jand g13437(.dina(n13722),.dinb(w_n13710_0[1]),.dout(n13723),.clk(gclk));
	jxor g13438(.dina(w_n13545_0[0]),.dinb(w_n1317_17[2]),.dout(n13724),.clk(gclk));
	jor g13439(.dina(n13724),.dinb(w_n13723_22[2]),.dout(n13725),.clk(gclk));
	jxor g13440(.dina(n13725),.dinb(w_n13175_0[0]),.dout(n13726),.clk(gclk));
	jor g13441(.dina(w_n13723_22[1]),.dinb(w_n13177_1[0]),.dout(n13727),.clk(gclk));
	jnot g13442(.din(w_a24_0[1]),.dout(n13728),.clk(gclk));
	jnot g13443(.din(a[25]),.dout(n13729),.clk(gclk));
	jand g13444(.dina(w_n13177_0[2]),.dinb(w_n13729_0[2]),.dout(n13730),.clk(gclk));
	jand g13445(.dina(n13730),.dinb(w_n13728_1[1]),.dout(n13731),.clk(gclk));
	jnot g13446(.din(n13731),.dout(n13732),.clk(gclk));
	jand g13447(.dina(n13732),.dinb(n13727),.dout(n13733),.clk(gclk));
	jor g13448(.dina(w_n13733_0[2]),.dinb(w_n13718_9[1]),.dout(n13734),.clk(gclk));
	jor g13449(.dina(w_n13723_22[0]),.dinb(w_a26_0[0]),.dout(n13735),.clk(gclk));
	jxor g13450(.dina(w_n13735_0[1]),.dinb(w_n13178_0[0]),.dout(n13736),.clk(gclk));
	jand g13451(.dina(w_n13733_0[1]),.dinb(w_n13718_9[0]),.dout(n13737),.clk(gclk));
	jor g13452(.dina(n13737),.dinb(w_n13736_0[1]),.dout(n13738),.clk(gclk));
	jand g13453(.dina(w_n13738_0[1]),.dinb(w_n13734_0[1]),.dout(n13739),.clk(gclk));
	jor g13454(.dina(n13739),.dinb(w_n12675_14[1]),.dout(n13740),.clk(gclk));
	jand g13455(.dina(w_n13734_0[0]),.dinb(w_n12675_14[0]),.dout(n13741),.clk(gclk));
	jand g13456(.dina(n13741),.dinb(w_n13738_0[0]),.dout(n13742),.clk(gclk));
	jor g13457(.dina(w_n13735_0[0]),.dinb(w_a27_0[0]),.dout(n13743),.clk(gclk));
	jnot g13458(.din(w_n13710_0[0]),.dout(n13744),.clk(gclk));
	jnot g13459(.din(w_n13712_0[0]),.dout(n13745),.clk(gclk));
	jor g13460(.dina(w_n13717_0[0]),.dinb(w_n13718_8[2]),.dout(n13746),.clk(gclk));
	jor g13461(.dina(n13746),.dinb(w_n13745_0[1]),.dout(n13747),.clk(gclk));
	jor g13462(.dina(n13747),.dinb(n13744),.dout(n13748),.clk(gclk));
	jand g13463(.dina(n13748),.dinb(n13743),.dout(n13749),.clk(gclk));
	jxor g13464(.dina(n13749),.dinb(w_n12681_0[1]),.dout(n13750),.clk(gclk));
	jor g13465(.dina(w_n13750_0[1]),.dinb(w_n13742_0[1]),.dout(n13751),.clk(gclk));
	jand g13466(.dina(n13751),.dinb(w_n13740_0[1]),.dout(n13752),.clk(gclk));
	jor g13467(.dina(w_n13752_0[2]),.dinb(w_n12670_9[1]),.dout(n13753),.clk(gclk));
	jand g13468(.dina(w_n13752_0[1]),.dinb(w_n12670_9[0]),.dout(n13754),.clk(gclk));
	jxor g13469(.dina(w_n13181_0[0]),.dinb(w_n12675_13[2]),.dout(n13755),.clk(gclk));
	jor g13470(.dina(n13755),.dinb(w_n13723_21[2]),.dout(n13756),.clk(gclk));
	jxor g13471(.dina(n13756),.dinb(w_n13184_0[0]),.dout(n13757),.clk(gclk));
	jor g13472(.dina(w_n13757_0[1]),.dinb(n13754),.dout(n13758),.clk(gclk));
	jand g13473(.dina(w_n13758_0[1]),.dinb(w_n13753_0[1]),.dout(n13759),.clk(gclk));
	jor g13474(.dina(n13759),.dinb(w_n11662_14[0]),.dout(n13760),.clk(gclk));
	jnot g13475(.din(w_n13190_0[0]),.dout(n13761),.clk(gclk));
	jor g13476(.dina(n13761),.dinb(w_n13188_0[0]),.dout(n13762),.clk(gclk));
	jor g13477(.dina(n13762),.dinb(w_n13723_21[1]),.dout(n13763),.clk(gclk));
	jxor g13478(.dina(n13763),.dinb(w_n13199_0[0]),.dout(n13764),.clk(gclk));
	jand g13479(.dina(w_n13753_0[0]),.dinb(w_n11662_13[2]),.dout(n13765),.clk(gclk));
	jand g13480(.dina(n13765),.dinb(w_n13758_0[0]),.dout(n13766),.clk(gclk));
	jor g13481(.dina(w_n13766_0[1]),.dinb(w_n13764_0[1]),.dout(n13767),.clk(gclk));
	jand g13482(.dina(w_n13767_0[1]),.dinb(w_n13760_0[1]),.dout(n13768),.clk(gclk));
	jor g13483(.dina(w_n13768_0[2]),.dinb(w_n11657_9[1]),.dout(n13769),.clk(gclk));
	jand g13484(.dina(w_n13768_0[1]),.dinb(w_n11657_9[0]),.dout(n13770),.clk(gclk));
	jxor g13485(.dina(w_n13201_0[0]),.dinb(w_n11662_13[1]),.dout(n13771),.clk(gclk));
	jor g13486(.dina(n13771),.dinb(w_n13723_21[0]),.dout(n13772),.clk(gclk));
	jxor g13487(.dina(n13772),.dinb(w_n13206_0[0]),.dout(n13773),.clk(gclk));
	jnot g13488(.din(w_n13773_0[1]),.dout(n13774),.clk(gclk));
	jor g13489(.dina(n13774),.dinb(n13770),.dout(n13775),.clk(gclk));
	jand g13490(.dina(w_n13775_0[1]),.dinb(w_n13769_0[1]),.dout(n13776),.clk(gclk));
	jor g13491(.dina(n13776),.dinb(w_n10701_14[1]),.dout(n13777),.clk(gclk));
	jand g13492(.dina(w_n13769_0[0]),.dinb(w_n10701_14[0]),.dout(n13778),.clk(gclk));
	jand g13493(.dina(n13778),.dinb(w_n13775_0[0]),.dout(n13779),.clk(gclk));
	jnot g13494(.din(w_n13210_0[0]),.dout(n13780),.clk(gclk));
	jnot g13495(.din(w_n13723_20[2]),.dout(asqrt_fa_14),.clk(gclk));
	jand g13496(.dina(w_asqrt13_17),.dinb(n13780),.dout(n13782),.clk(gclk));
	jand g13497(.dina(w_n13782_0[1]),.dinb(w_n13217_0[0]),.dout(n13783),.clk(gclk));
	jor g13498(.dina(n13783),.dinb(w_n13215_0[0]),.dout(n13784),.clk(gclk));
	jand g13499(.dina(w_n13782_0[0]),.dinb(w_n13218_0[0]),.dout(n13785),.clk(gclk));
	jnot g13500(.din(n13785),.dout(n13786),.clk(gclk));
	jand g13501(.dina(n13786),.dinb(n13784),.dout(n13787),.clk(gclk));
	jnot g13502(.din(n13787),.dout(n13788),.clk(gclk));
	jor g13503(.dina(w_n13788_0[1]),.dinb(w_n13779_0[1]),.dout(n13789),.clk(gclk));
	jand g13504(.dina(n13789),.dinb(w_n13777_0[1]),.dout(n13790),.clk(gclk));
	jor g13505(.dina(w_n13790_0[2]),.dinb(w_n10696_10[0]),.dout(n13791),.clk(gclk));
	jand g13506(.dina(w_n13790_0[1]),.dinb(w_n10696_9[2]),.dout(n13792),.clk(gclk));
	jnot g13507(.din(w_n13225_0[0]),.dout(n13793),.clk(gclk));
	jxor g13508(.dina(w_n13219_0[0]),.dinb(w_n10701_13[2]),.dout(n13794),.clk(gclk));
	jor g13509(.dina(n13794),.dinb(w_n13723_20[1]),.dout(n13795),.clk(gclk));
	jxor g13510(.dina(n13795),.dinb(n13793),.dout(n13796),.clk(gclk));
	jnot g13511(.din(w_n13796_0[1]),.dout(n13797),.clk(gclk));
	jor g13512(.dina(n13797),.dinb(n13792),.dout(n13798),.clk(gclk));
	jand g13513(.dina(w_n13798_0[1]),.dinb(w_n13791_0[1]),.dout(n13799),.clk(gclk));
	jor g13514(.dina(n13799),.dinb(w_n9774_14[0]),.dout(n13800),.clk(gclk));
	jnot g13515(.din(w_n13230_0[0]),.dout(n13801),.clk(gclk));
	jor g13516(.dina(n13801),.dinb(w_n13228_0[0]),.dout(n13802),.clk(gclk));
	jor g13517(.dina(n13802),.dinb(w_n13723_20[0]),.dout(n13803),.clk(gclk));
	jxor g13518(.dina(n13803),.dinb(w_n13239_0[0]),.dout(n13804),.clk(gclk));
	jand g13519(.dina(w_n13791_0[0]),.dinb(w_n9774_13[2]),.dout(n13805),.clk(gclk));
	jand g13520(.dina(n13805),.dinb(w_n13798_0[0]),.dout(n13806),.clk(gclk));
	jor g13521(.dina(w_n13806_0[1]),.dinb(w_n13804_0[1]),.dout(n13807),.clk(gclk));
	jand g13522(.dina(w_n13807_0[1]),.dinb(w_n13800_0[1]),.dout(n13808),.clk(gclk));
	jor g13523(.dina(w_n13808_0[2]),.dinb(w_n9769_10[0]),.dout(n13809),.clk(gclk));
	jand g13524(.dina(w_n13808_0[1]),.dinb(w_n9769_9[2]),.dout(n13810),.clk(gclk));
	jnot g13525(.din(w_n13246_0[0]),.dout(n13811),.clk(gclk));
	jxor g13526(.dina(w_n13241_0[0]),.dinb(w_n9774_13[1]),.dout(n13812),.clk(gclk));
	jor g13527(.dina(n13812),.dinb(w_n13723_19[2]),.dout(n13813),.clk(gclk));
	jxor g13528(.dina(n13813),.dinb(n13811),.dout(n13814),.clk(gclk));
	jnot g13529(.din(n13814),.dout(n13815),.clk(gclk));
	jor g13530(.dina(w_n13815_0[1]),.dinb(n13810),.dout(n13816),.clk(gclk));
	jand g13531(.dina(w_n13816_0[1]),.dinb(w_n13809_0[1]),.dout(n13817),.clk(gclk));
	jor g13532(.dina(n13817),.dinb(w_n8898_14[2]),.dout(n13818),.clk(gclk));
	jand g13533(.dina(w_n13809_0[0]),.dinb(w_n8898_14[1]),.dout(n13819),.clk(gclk));
	jand g13534(.dina(n13819),.dinb(w_n13816_0[0]),.dout(n13820),.clk(gclk));
	jnot g13535(.din(w_n13249_0[0]),.dout(n13821),.clk(gclk));
	jand g13536(.dina(w_asqrt13_16[2]),.dinb(n13821),.dout(n13822),.clk(gclk));
	jand g13537(.dina(w_n13822_0[1]),.dinb(w_n13256_0[0]),.dout(n13823),.clk(gclk));
	jor g13538(.dina(n13823),.dinb(w_n13254_0[0]),.dout(n13824),.clk(gclk));
	jand g13539(.dina(w_n13822_0[0]),.dinb(w_n13257_0[0]),.dout(n13825),.clk(gclk));
	jnot g13540(.din(n13825),.dout(n13826),.clk(gclk));
	jand g13541(.dina(n13826),.dinb(n13824),.dout(n13827),.clk(gclk));
	jnot g13542(.din(n13827),.dout(n13828),.clk(gclk));
	jor g13543(.dina(w_n13828_0[1]),.dinb(w_n13820_0[1]),.dout(n13829),.clk(gclk));
	jand g13544(.dina(n13829),.dinb(w_n13818_0[1]),.dout(n13830),.clk(gclk));
	jor g13545(.dina(w_n13830_0[1]),.dinb(w_n8893_10[1]),.dout(n13831),.clk(gclk));
	jxor g13546(.dina(w_n13258_0[0]),.dinb(w_n8898_14[0]),.dout(n13832),.clk(gclk));
	jor g13547(.dina(n13832),.dinb(w_n13723_19[1]),.dout(n13833),.clk(gclk));
	jxor g13548(.dina(n13833),.dinb(w_n13263_0[0]),.dout(n13834),.clk(gclk));
	jand g13549(.dina(w_n13830_0[0]),.dinb(w_n8893_10[0]),.dout(n13835),.clk(gclk));
	jor g13550(.dina(w_n13835_0[1]),.dinb(w_n13834_0[1]),.dout(n13836),.clk(gclk));
	jand g13551(.dina(w_n13836_0[2]),.dinb(w_n13831_0[2]),.dout(n13837),.clk(gclk));
	jor g13552(.dina(n13837),.dinb(w_n8058_14[1]),.dout(n13838),.clk(gclk));
	jnot g13553(.din(w_n13268_0[0]),.dout(n13839),.clk(gclk));
	jor g13554(.dina(n13839),.dinb(w_n13266_0[0]),.dout(n13840),.clk(gclk));
	jor g13555(.dina(n13840),.dinb(w_n13723_19[0]),.dout(n13841),.clk(gclk));
	jxor g13556(.dina(n13841),.dinb(w_n13277_0[0]),.dout(n13842),.clk(gclk));
	jand g13557(.dina(w_n13831_0[1]),.dinb(w_n8058_14[0]),.dout(n13843),.clk(gclk));
	jand g13558(.dina(n13843),.dinb(w_n13836_0[1]),.dout(n13844),.clk(gclk));
	jor g13559(.dina(w_n13844_0[1]),.dinb(w_n13842_0[1]),.dout(n13845),.clk(gclk));
	jand g13560(.dina(w_n13845_0[1]),.dinb(w_n13838_0[1]),.dout(n13846),.clk(gclk));
	jor g13561(.dina(w_n13846_0[2]),.dinb(w_n8053_10[2]),.dout(n13847),.clk(gclk));
	jand g13562(.dina(w_n13846_0[1]),.dinb(w_n8053_10[1]),.dout(n13848),.clk(gclk));
	jnot g13563(.din(w_n13280_0[0]),.dout(n13849),.clk(gclk));
	jand g13564(.dina(w_asqrt13_16[1]),.dinb(n13849),.dout(n13850),.clk(gclk));
	jand g13565(.dina(w_n13850_0[1]),.dinb(w_n13285_0[0]),.dout(n13851),.clk(gclk));
	jor g13566(.dina(n13851),.dinb(w_n13284_0[0]),.dout(n13852),.clk(gclk));
	jand g13567(.dina(w_n13850_0[0]),.dinb(w_n13286_0[0]),.dout(n13853),.clk(gclk));
	jnot g13568(.din(n13853),.dout(n13854),.clk(gclk));
	jand g13569(.dina(n13854),.dinb(n13852),.dout(n13855),.clk(gclk));
	jnot g13570(.din(n13855),.dout(n13856),.clk(gclk));
	jor g13571(.dina(w_n13856_0[1]),.dinb(n13848),.dout(n13857),.clk(gclk));
	jand g13572(.dina(w_n13857_0[1]),.dinb(w_n13847_0[1]),.dout(n13858),.clk(gclk));
	jor g13573(.dina(n13858),.dinb(w_n7265_15[0]),.dout(n13859),.clk(gclk));
	jand g13574(.dina(w_n13847_0[0]),.dinb(w_n7265_14[2]),.dout(n13860),.clk(gclk));
	jand g13575(.dina(n13860),.dinb(w_n13857_0[0]),.dout(n13861),.clk(gclk));
	jnot g13576(.din(w_n13288_0[0]),.dout(n13862),.clk(gclk));
	jand g13577(.dina(w_asqrt13_16[0]),.dinb(n13862),.dout(n13863),.clk(gclk));
	jand g13578(.dina(w_n13863_0[1]),.dinb(w_n13295_0[0]),.dout(n13864),.clk(gclk));
	jor g13579(.dina(n13864),.dinb(w_n13293_0[0]),.dout(n13865),.clk(gclk));
	jand g13580(.dina(w_n13863_0[0]),.dinb(w_n13296_0[0]),.dout(n13866),.clk(gclk));
	jnot g13581(.din(n13866),.dout(n13867),.clk(gclk));
	jand g13582(.dina(n13867),.dinb(n13865),.dout(n13868),.clk(gclk));
	jnot g13583(.din(n13868),.dout(n13869),.clk(gclk));
	jor g13584(.dina(w_n13869_0[1]),.dinb(w_n13861_0[1]),.dout(n13870),.clk(gclk));
	jand g13585(.dina(n13870),.dinb(w_n13859_0[1]),.dout(n13871),.clk(gclk));
	jor g13586(.dina(w_n13871_0[1]),.dinb(w_n7260_11[1]),.dout(n13872),.clk(gclk));
	jxor g13587(.dina(w_n13297_0[0]),.dinb(w_n7265_14[1]),.dout(n13873),.clk(gclk));
	jor g13588(.dina(n13873),.dinb(w_n13723_18[2]),.dout(n13874),.clk(gclk));
	jxor g13589(.dina(n13874),.dinb(w_n13308_0[0]),.dout(n13875),.clk(gclk));
	jand g13590(.dina(w_n13871_0[0]),.dinb(w_n7260_11[0]),.dout(n13876),.clk(gclk));
	jor g13591(.dina(w_n13876_0[1]),.dinb(w_n13875_0[1]),.dout(n13877),.clk(gclk));
	jand g13592(.dina(w_n13877_0[2]),.dinb(w_n13872_0[2]),.dout(n13878),.clk(gclk));
	jor g13593(.dina(n13878),.dinb(w_n6505_14[2]),.dout(n13879),.clk(gclk));
	jnot g13594(.din(w_n13313_0[0]),.dout(n13880),.clk(gclk));
	jor g13595(.dina(n13880),.dinb(w_n13311_0[0]),.dout(n13881),.clk(gclk));
	jor g13596(.dina(n13881),.dinb(w_n13723_18[1]),.dout(n13882),.clk(gclk));
	jxor g13597(.dina(n13882),.dinb(w_n13322_0[0]),.dout(n13883),.clk(gclk));
	jand g13598(.dina(w_n13872_0[1]),.dinb(w_n6505_14[1]),.dout(n13884),.clk(gclk));
	jand g13599(.dina(n13884),.dinb(w_n13877_0[1]),.dout(n13885),.clk(gclk));
	jor g13600(.dina(w_n13885_0[1]),.dinb(w_n13883_0[1]),.dout(n13886),.clk(gclk));
	jand g13601(.dina(w_n13886_0[1]),.dinb(w_n13879_0[1]),.dout(n13887),.clk(gclk));
	jor g13602(.dina(w_n13887_0[2]),.dinb(w_n6500_11[2]),.dout(n13888),.clk(gclk));
	jand g13603(.dina(w_n13887_0[1]),.dinb(w_n6500_11[1]),.dout(n13889),.clk(gclk));
	jnot g13604(.din(w_n13325_0[0]),.dout(n13890),.clk(gclk));
	jand g13605(.dina(w_asqrt13_15[2]),.dinb(n13890),.dout(n13891),.clk(gclk));
	jand g13606(.dina(w_n13891_0[1]),.dinb(w_n13330_0[0]),.dout(n13892),.clk(gclk));
	jor g13607(.dina(n13892),.dinb(w_n13329_0[0]),.dout(n13893),.clk(gclk));
	jand g13608(.dina(w_n13891_0[0]),.dinb(w_n13331_0[0]),.dout(n13894),.clk(gclk));
	jnot g13609(.din(n13894),.dout(n13895),.clk(gclk));
	jand g13610(.dina(n13895),.dinb(n13893),.dout(n13896),.clk(gclk));
	jnot g13611(.din(n13896),.dout(n13897),.clk(gclk));
	jor g13612(.dina(w_n13897_0[1]),.dinb(n13889),.dout(n13898),.clk(gclk));
	jand g13613(.dina(w_n13898_0[1]),.dinb(w_n13888_0[1]),.dout(n13899),.clk(gclk));
	jor g13614(.dina(n13899),.dinb(w_n5793_15[1]),.dout(n13900),.clk(gclk));
	jand g13615(.dina(w_n13888_0[0]),.dinb(w_n5793_15[0]),.dout(n13901),.clk(gclk));
	jand g13616(.dina(n13901),.dinb(w_n13898_0[0]),.dout(n13902),.clk(gclk));
	jnot g13617(.din(w_n13333_0[0]),.dout(n13903),.clk(gclk));
	jand g13618(.dina(w_asqrt13_15[1]),.dinb(n13903),.dout(n13904),.clk(gclk));
	jand g13619(.dina(w_n13904_0[1]),.dinb(w_n13340_0[0]),.dout(n13905),.clk(gclk));
	jor g13620(.dina(n13905),.dinb(w_n13338_0[0]),.dout(n13906),.clk(gclk));
	jand g13621(.dina(w_n13904_0[0]),.dinb(w_n13341_0[0]),.dout(n13907),.clk(gclk));
	jnot g13622(.din(n13907),.dout(n13908),.clk(gclk));
	jand g13623(.dina(n13908),.dinb(n13906),.dout(n13909),.clk(gclk));
	jnot g13624(.din(n13909),.dout(n13910),.clk(gclk));
	jor g13625(.dina(w_n13910_0[1]),.dinb(w_n13902_0[1]),.dout(n13911),.clk(gclk));
	jand g13626(.dina(n13911),.dinb(w_n13900_0[1]),.dout(n13912),.clk(gclk));
	jor g13627(.dina(w_n13912_0[1]),.dinb(w_n5788_12[0]),.dout(n13913),.clk(gclk));
	jxor g13628(.dina(w_n13342_0[0]),.dinb(w_n5793_14[2]),.dout(n13914),.clk(gclk));
	jor g13629(.dina(n13914),.dinb(w_n13723_18[0]),.dout(n13915),.clk(gclk));
	jxor g13630(.dina(n13915),.dinb(w_n13353_0[0]),.dout(n13916),.clk(gclk));
	jand g13631(.dina(w_n13912_0[0]),.dinb(w_n5788_11[2]),.dout(n13917),.clk(gclk));
	jor g13632(.dina(w_n13917_0[1]),.dinb(w_n13916_0[1]),.dout(n13918),.clk(gclk));
	jand g13633(.dina(w_n13918_0[2]),.dinb(w_n13913_0[2]),.dout(n13919),.clk(gclk));
	jor g13634(.dina(n13919),.dinb(w_n5121_15[0]),.dout(n13920),.clk(gclk));
	jnot g13635(.din(w_n13358_0[0]),.dout(n13921),.clk(gclk));
	jor g13636(.dina(n13921),.dinb(w_n13356_0[0]),.dout(n13922),.clk(gclk));
	jor g13637(.dina(n13922),.dinb(w_n13723_17[2]),.dout(n13923),.clk(gclk));
	jxor g13638(.dina(n13923),.dinb(w_n13367_0[0]),.dout(n13924),.clk(gclk));
	jand g13639(.dina(w_n13913_0[1]),.dinb(w_n5121_14[2]),.dout(n13925),.clk(gclk));
	jand g13640(.dina(n13925),.dinb(w_n13918_0[1]),.dout(n13926),.clk(gclk));
	jor g13641(.dina(w_n13926_0[1]),.dinb(w_n13924_0[1]),.dout(n13927),.clk(gclk));
	jand g13642(.dina(w_n13927_0[1]),.dinb(w_n13920_0[1]),.dout(n13928),.clk(gclk));
	jor g13643(.dina(w_n13928_0[2]),.dinb(w_n5116_12[1]),.dout(n13929),.clk(gclk));
	jand g13644(.dina(w_n13928_0[1]),.dinb(w_n5116_12[0]),.dout(n13930),.clk(gclk));
	jnot g13645(.din(w_n13370_0[0]),.dout(n13931),.clk(gclk));
	jand g13646(.dina(w_asqrt13_15[0]),.dinb(n13931),.dout(n13932),.clk(gclk));
	jand g13647(.dina(w_n13932_0[1]),.dinb(w_n13375_0[0]),.dout(n13933),.clk(gclk));
	jor g13648(.dina(n13933),.dinb(w_n13374_0[0]),.dout(n13934),.clk(gclk));
	jand g13649(.dina(w_n13932_0[0]),.dinb(w_n13376_0[0]),.dout(n13935),.clk(gclk));
	jnot g13650(.din(n13935),.dout(n13936),.clk(gclk));
	jand g13651(.dina(n13936),.dinb(n13934),.dout(n13937),.clk(gclk));
	jnot g13652(.din(n13937),.dout(n13938),.clk(gclk));
	jor g13653(.dina(w_n13938_0[1]),.dinb(n13930),.dout(n13939),.clk(gclk));
	jand g13654(.dina(w_n13939_0[1]),.dinb(w_n13929_0[1]),.dout(n13940),.clk(gclk));
	jor g13655(.dina(n13940),.dinb(w_n4499_16[0]),.dout(n13941),.clk(gclk));
	jand g13656(.dina(w_n13929_0[0]),.dinb(w_n4499_15[2]),.dout(n13942),.clk(gclk));
	jand g13657(.dina(n13942),.dinb(w_n13939_0[0]),.dout(n13943),.clk(gclk));
	jnot g13658(.din(w_n13378_0[0]),.dout(n13944),.clk(gclk));
	jand g13659(.dina(w_asqrt13_14[2]),.dinb(n13944),.dout(n13945),.clk(gclk));
	jand g13660(.dina(w_n13945_0[1]),.dinb(w_n13385_0[0]),.dout(n13946),.clk(gclk));
	jor g13661(.dina(n13946),.dinb(w_n13383_0[0]),.dout(n13947),.clk(gclk));
	jand g13662(.dina(w_n13945_0[0]),.dinb(w_n13386_0[0]),.dout(n13948),.clk(gclk));
	jnot g13663(.din(n13948),.dout(n13949),.clk(gclk));
	jand g13664(.dina(n13949),.dinb(n13947),.dout(n13950),.clk(gclk));
	jnot g13665(.din(n13950),.dout(n13951),.clk(gclk));
	jor g13666(.dina(w_n13951_0[1]),.dinb(w_n13943_0[1]),.dout(n13952),.clk(gclk));
	jand g13667(.dina(n13952),.dinb(w_n13941_0[1]),.dout(n13953),.clk(gclk));
	jor g13668(.dina(w_n13953_0[1]),.dinb(w_n4494_13[0]),.dout(n13954),.clk(gclk));
	jxor g13669(.dina(w_n13387_0[0]),.dinb(w_n4499_15[1]),.dout(n13955),.clk(gclk));
	jor g13670(.dina(n13955),.dinb(w_n13723_17[1]),.dout(n13956),.clk(gclk));
	jxor g13671(.dina(n13956),.dinb(w_n13398_0[0]),.dout(n13957),.clk(gclk));
	jand g13672(.dina(w_n13953_0[0]),.dinb(w_n4494_12[2]),.dout(n13958),.clk(gclk));
	jor g13673(.dina(w_n13958_0[1]),.dinb(w_n13957_0[1]),.dout(n13959),.clk(gclk));
	jand g13674(.dina(w_n13959_0[2]),.dinb(w_n13954_0[2]),.dout(n13960),.clk(gclk));
	jor g13675(.dina(n13960),.dinb(w_n3912_15[2]),.dout(n13961),.clk(gclk));
	jnot g13676(.din(w_n13403_0[0]),.dout(n13962),.clk(gclk));
	jor g13677(.dina(n13962),.dinb(w_n13401_0[0]),.dout(n13963),.clk(gclk));
	jor g13678(.dina(n13963),.dinb(w_n13723_17[0]),.dout(n13964),.clk(gclk));
	jxor g13679(.dina(n13964),.dinb(w_n13412_0[0]),.dout(n13965),.clk(gclk));
	jand g13680(.dina(w_n13954_0[1]),.dinb(w_n3912_15[1]),.dout(n13966),.clk(gclk));
	jand g13681(.dina(n13966),.dinb(w_n13959_0[1]),.dout(n13967),.clk(gclk));
	jor g13682(.dina(w_n13967_0[1]),.dinb(w_n13965_0[1]),.dout(n13968),.clk(gclk));
	jand g13683(.dina(w_n13968_0[1]),.dinb(w_n13961_0[1]),.dout(n13969),.clk(gclk));
	jor g13684(.dina(w_n13969_0[2]),.dinb(w_n3907_13[1]),.dout(n13970),.clk(gclk));
	jand g13685(.dina(w_n13969_0[1]),.dinb(w_n3907_13[0]),.dout(n13971),.clk(gclk));
	jnot g13686(.din(w_n13415_0[0]),.dout(n13972),.clk(gclk));
	jand g13687(.dina(w_asqrt13_14[1]),.dinb(n13972),.dout(n13973),.clk(gclk));
	jand g13688(.dina(w_n13973_0[1]),.dinb(w_n13420_0[0]),.dout(n13974),.clk(gclk));
	jor g13689(.dina(n13974),.dinb(w_n13419_0[0]),.dout(n13975),.clk(gclk));
	jand g13690(.dina(w_n13973_0[0]),.dinb(w_n13421_0[0]),.dout(n13976),.clk(gclk));
	jnot g13691(.din(n13976),.dout(n13977),.clk(gclk));
	jand g13692(.dina(n13977),.dinb(n13975),.dout(n13978),.clk(gclk));
	jnot g13693(.din(n13978),.dout(n13979),.clk(gclk));
	jor g13694(.dina(w_n13979_0[1]),.dinb(n13971),.dout(n13980),.clk(gclk));
	jand g13695(.dina(w_n13980_0[1]),.dinb(w_n13970_0[1]),.dout(n13981),.clk(gclk));
	jor g13696(.dina(n13981),.dinb(w_n3376_16[2]),.dout(n13982),.clk(gclk));
	jand g13697(.dina(w_n13970_0[0]),.dinb(w_n3376_16[1]),.dout(n13983),.clk(gclk));
	jand g13698(.dina(n13983),.dinb(w_n13980_0[0]),.dout(n13984),.clk(gclk));
	jnot g13699(.din(w_n13423_0[0]),.dout(n13985),.clk(gclk));
	jand g13700(.dina(w_asqrt13_14[0]),.dinb(n13985),.dout(n13986),.clk(gclk));
	jand g13701(.dina(w_n13986_0[1]),.dinb(w_n13430_0[0]),.dout(n13987),.clk(gclk));
	jor g13702(.dina(n13987),.dinb(w_n13428_0[0]),.dout(n13988),.clk(gclk));
	jand g13703(.dina(w_n13986_0[0]),.dinb(w_n13431_0[0]),.dout(n13989),.clk(gclk));
	jnot g13704(.din(n13989),.dout(n13990),.clk(gclk));
	jand g13705(.dina(n13990),.dinb(n13988),.dout(n13991),.clk(gclk));
	jnot g13706(.din(n13991),.dout(n13992),.clk(gclk));
	jor g13707(.dina(w_n13992_0[1]),.dinb(w_n13984_0[1]),.dout(n13993),.clk(gclk));
	jand g13708(.dina(n13993),.dinb(w_n13982_0[1]),.dout(n13994),.clk(gclk));
	jor g13709(.dina(w_n13994_0[1]),.dinb(w_n3371_13[2]),.dout(n13995),.clk(gclk));
	jxor g13710(.dina(w_n13432_0[0]),.dinb(w_n3376_16[0]),.dout(n13996),.clk(gclk));
	jor g13711(.dina(n13996),.dinb(w_n13723_16[2]),.dout(n13997),.clk(gclk));
	jxor g13712(.dina(n13997),.dinb(w_n13443_0[0]),.dout(n13998),.clk(gclk));
	jand g13713(.dina(w_n13994_0[0]),.dinb(w_n3371_13[1]),.dout(n13999),.clk(gclk));
	jor g13714(.dina(w_n13999_0[1]),.dinb(w_n13998_0[1]),.dout(n14000),.clk(gclk));
	jand g13715(.dina(w_n14000_0[2]),.dinb(w_n13995_0[2]),.dout(n14001),.clk(gclk));
	jor g13716(.dina(n14001),.dinb(w_n2875_16[1]),.dout(n14002),.clk(gclk));
	jnot g13717(.din(w_n13448_0[0]),.dout(n14003),.clk(gclk));
	jor g13718(.dina(n14003),.dinb(w_n13446_0[0]),.dout(n14004),.clk(gclk));
	jor g13719(.dina(n14004),.dinb(w_n13723_16[1]),.dout(n14005),.clk(gclk));
	jxor g13720(.dina(n14005),.dinb(w_n13457_0[0]),.dout(n14006),.clk(gclk));
	jand g13721(.dina(w_n13995_0[1]),.dinb(w_n2875_16[0]),.dout(n14007),.clk(gclk));
	jand g13722(.dina(n14007),.dinb(w_n14000_0[1]),.dout(n14008),.clk(gclk));
	jor g13723(.dina(w_n14008_0[1]),.dinb(w_n14006_0[1]),.dout(n14009),.clk(gclk));
	jand g13724(.dina(w_n14009_0[1]),.dinb(w_n14002_0[1]),.dout(n14010),.clk(gclk));
	jor g13725(.dina(w_n14010_0[2]),.dinb(w_n2870_14[0]),.dout(n14011),.clk(gclk));
	jand g13726(.dina(w_n14010_0[1]),.dinb(w_n2870_13[2]),.dout(n14012),.clk(gclk));
	jnot g13727(.din(w_n13460_0[0]),.dout(n14013),.clk(gclk));
	jand g13728(.dina(w_asqrt13_13[2]),.dinb(n14013),.dout(n14014),.clk(gclk));
	jand g13729(.dina(w_n14014_0[1]),.dinb(w_n13465_0[0]),.dout(n14015),.clk(gclk));
	jor g13730(.dina(n14015),.dinb(w_n13464_0[0]),.dout(n14016),.clk(gclk));
	jand g13731(.dina(w_n14014_0[0]),.dinb(w_n13466_0[0]),.dout(n14017),.clk(gclk));
	jnot g13732(.din(n14017),.dout(n14018),.clk(gclk));
	jand g13733(.dina(n14018),.dinb(n14016),.dout(n14019),.clk(gclk));
	jnot g13734(.din(n14019),.dout(n14020),.clk(gclk));
	jor g13735(.dina(w_n14020_0[1]),.dinb(n14012),.dout(n14021),.clk(gclk));
	jand g13736(.dina(w_n14021_0[1]),.dinb(w_n14011_0[1]),.dout(n14022),.clk(gclk));
	jor g13737(.dina(n14022),.dinb(w_n2425_17[0]),.dout(n14023),.clk(gclk));
	jand g13738(.dina(w_n14011_0[0]),.dinb(w_n2425_16[2]),.dout(n14024),.clk(gclk));
	jand g13739(.dina(n14024),.dinb(w_n14021_0[0]),.dout(n14025),.clk(gclk));
	jnot g13740(.din(w_n13468_0[0]),.dout(n14026),.clk(gclk));
	jand g13741(.dina(w_asqrt13_13[1]),.dinb(n14026),.dout(n14027),.clk(gclk));
	jand g13742(.dina(w_n14027_0[1]),.dinb(w_n13475_0[0]),.dout(n14028),.clk(gclk));
	jor g13743(.dina(n14028),.dinb(w_n13473_0[0]),.dout(n14029),.clk(gclk));
	jand g13744(.dina(w_n14027_0[0]),.dinb(w_n13476_0[0]),.dout(n14030),.clk(gclk));
	jnot g13745(.din(n14030),.dout(n14031),.clk(gclk));
	jand g13746(.dina(n14031),.dinb(n14029),.dout(n14032),.clk(gclk));
	jnot g13747(.din(n14032),.dout(n14033),.clk(gclk));
	jor g13748(.dina(w_n14033_0[1]),.dinb(w_n14025_0[1]),.dout(n14034),.clk(gclk));
	jand g13749(.dina(n14034),.dinb(w_n14023_0[1]),.dout(n14035),.clk(gclk));
	jor g13750(.dina(w_n14035_0[1]),.dinb(w_n2420_14[2]),.dout(n14036),.clk(gclk));
	jxor g13751(.dina(w_n13477_0[0]),.dinb(w_n2425_16[1]),.dout(n14037),.clk(gclk));
	jor g13752(.dina(n14037),.dinb(w_n13723_16[0]),.dout(n14038),.clk(gclk));
	jxor g13753(.dina(n14038),.dinb(w_n13488_0[0]),.dout(n14039),.clk(gclk));
	jand g13754(.dina(w_n14035_0[0]),.dinb(w_n2420_14[1]),.dout(n14040),.clk(gclk));
	jor g13755(.dina(w_n14040_0[1]),.dinb(w_n14039_0[1]),.dout(n14041),.clk(gclk));
	jand g13756(.dina(w_n14041_0[2]),.dinb(w_n14036_0[2]),.dout(n14042),.clk(gclk));
	jor g13757(.dina(n14042),.dinb(w_n2010_16[2]),.dout(n14043),.clk(gclk));
	jnot g13758(.din(w_n13493_0[0]),.dout(n14044),.clk(gclk));
	jor g13759(.dina(n14044),.dinb(w_n13491_0[0]),.dout(n14045),.clk(gclk));
	jor g13760(.dina(n14045),.dinb(w_n13723_15[2]),.dout(n14046),.clk(gclk));
	jxor g13761(.dina(n14046),.dinb(w_n13502_0[0]),.dout(n14047),.clk(gclk));
	jand g13762(.dina(w_n14036_0[1]),.dinb(w_n2010_16[1]),.dout(n14048),.clk(gclk));
	jand g13763(.dina(n14048),.dinb(w_n14041_0[1]),.dout(n14049),.clk(gclk));
	jor g13764(.dina(w_n14049_0[1]),.dinb(w_n14047_0[1]),.dout(n14050),.clk(gclk));
	jand g13765(.dina(w_n14050_0[1]),.dinb(w_n14043_0[1]),.dout(n14051),.clk(gclk));
	jor g13766(.dina(w_n14051_0[2]),.dinb(w_n2005_15[0]),.dout(n14052),.clk(gclk));
	jand g13767(.dina(w_n14051_0[1]),.dinb(w_n2005_14[2]),.dout(n14053),.clk(gclk));
	jnot g13768(.din(w_n13505_0[0]),.dout(n14054),.clk(gclk));
	jand g13769(.dina(w_asqrt13_13[0]),.dinb(n14054),.dout(n14055),.clk(gclk));
	jand g13770(.dina(w_n14055_0[1]),.dinb(w_n13510_0[0]),.dout(n14056),.clk(gclk));
	jor g13771(.dina(n14056),.dinb(w_n13509_0[0]),.dout(n14057),.clk(gclk));
	jand g13772(.dina(w_n14055_0[0]),.dinb(w_n13511_0[0]),.dout(n14058),.clk(gclk));
	jnot g13773(.din(n14058),.dout(n14059),.clk(gclk));
	jand g13774(.dina(n14059),.dinb(n14057),.dout(n14060),.clk(gclk));
	jnot g13775(.din(n14060),.dout(n14061),.clk(gclk));
	jor g13776(.dina(w_n14061_0[1]),.dinb(n14053),.dout(n14062),.clk(gclk));
	jand g13777(.dina(w_n14062_0[1]),.dinb(w_n14052_0[1]),.dout(n14063),.clk(gclk));
	jor g13778(.dina(n14063),.dinb(w_n1646_17[2]),.dout(n14064),.clk(gclk));
	jand g13779(.dina(w_n14052_0[0]),.dinb(w_n1646_17[1]),.dout(n14065),.clk(gclk));
	jand g13780(.dina(n14065),.dinb(w_n14062_0[0]),.dout(n14066),.clk(gclk));
	jnot g13781(.din(w_n13513_0[0]),.dout(n14067),.clk(gclk));
	jand g13782(.dina(w_asqrt13_12[2]),.dinb(n14067),.dout(n14068),.clk(gclk));
	jand g13783(.dina(w_n14068_0[1]),.dinb(w_n13520_0[0]),.dout(n14069),.clk(gclk));
	jor g13784(.dina(n14069),.dinb(w_n13518_0[0]),.dout(n14070),.clk(gclk));
	jand g13785(.dina(w_n14068_0[0]),.dinb(w_n13521_0[0]),.dout(n14071),.clk(gclk));
	jnot g13786(.din(n14071),.dout(n14072),.clk(gclk));
	jand g13787(.dina(n14072),.dinb(n14070),.dout(n14073),.clk(gclk));
	jnot g13788(.din(n14073),.dout(n14074),.clk(gclk));
	jor g13789(.dina(w_n14074_0[1]),.dinb(w_n14066_0[1]),.dout(n14075),.clk(gclk));
	jand g13790(.dina(n14075),.dinb(w_n14064_0[1]),.dout(n14076),.clk(gclk));
	jor g13791(.dina(w_n14076_0[1]),.dinb(w_n1641_15[1]),.dout(n14077),.clk(gclk));
	jxor g13792(.dina(w_n13522_0[0]),.dinb(w_n1646_17[0]),.dout(n14078),.clk(gclk));
	jor g13793(.dina(n14078),.dinb(w_n13723_15[1]),.dout(n14079),.clk(gclk));
	jxor g13794(.dina(n14079),.dinb(w_n13533_0[0]),.dout(n14080),.clk(gclk));
	jand g13795(.dina(w_n14076_0[0]),.dinb(w_n1641_15[0]),.dout(n14081),.clk(gclk));
	jor g13796(.dina(w_n14081_0[1]),.dinb(w_n14080_0[1]),.dout(n14082),.clk(gclk));
	jand g13797(.dina(w_n14082_0[2]),.dinb(w_n14077_0[2]),.dout(n14083),.clk(gclk));
	jor g13798(.dina(n14083),.dinb(w_n1317_17[1]),.dout(n14084),.clk(gclk));
	jand g13799(.dina(w_n14077_0[1]),.dinb(w_n1317_17[0]),.dout(n14085),.clk(gclk));
	jand g13800(.dina(n14085),.dinb(w_n14082_0[1]),.dout(n14086),.clk(gclk));
	jnot g13801(.din(w_n13536_0[0]),.dout(n14087),.clk(gclk));
	jand g13802(.dina(w_asqrt13_12[1]),.dinb(n14087),.dout(n14088),.clk(gclk));
	jand g13803(.dina(w_n14088_0[1]),.dinb(w_n13543_0[0]),.dout(n14089),.clk(gclk));
	jor g13804(.dina(n14089),.dinb(w_n13541_0[0]),.dout(n14090),.clk(gclk));
	jand g13805(.dina(w_n14088_0[0]),.dinb(w_n13544_0[0]),.dout(n14091),.clk(gclk));
	jnot g13806(.din(n14091),.dout(n14092),.clk(gclk));
	jand g13807(.dina(n14092),.dinb(n14090),.dout(n14093),.clk(gclk));
	jnot g13808(.din(n14093),.dout(n14094),.clk(gclk));
	jor g13809(.dina(w_n14094_0[1]),.dinb(w_n14086_0[1]),.dout(n14095),.clk(gclk));
	jand g13810(.dina(n14095),.dinb(w_n14084_0[1]),.dout(n14096),.clk(gclk));
	jor g13811(.dina(w_n14096_0[2]),.dinb(w_n1312_15[2]),.dout(n14097),.clk(gclk));
	jand g13812(.dina(w_n14096_0[1]),.dinb(w_n1312_15[1]),.dout(n14098),.clk(gclk));
	jor g13813(.dina(n14098),.dinb(w_n13726_0[1]),.dout(n14099),.clk(gclk));
	jand g13814(.dina(w_n14099_0[1]),.dinb(w_n14097_0[1]),.dout(n14100),.clk(gclk));
	jor g13815(.dina(n14100),.dinb(w_n1039_18[1]),.dout(n14101),.clk(gclk));
	jnot g13816(.din(w_n13552_0[0]),.dout(n14102),.clk(gclk));
	jor g13817(.dina(n14102),.dinb(w_n13550_0[0]),.dout(n14103),.clk(gclk));
	jor g13818(.dina(n14103),.dinb(w_n13723_15[0]),.dout(n14104),.clk(gclk));
	jxor g13819(.dina(n14104),.dinb(w_n13561_0[0]),.dout(n14105),.clk(gclk));
	jand g13820(.dina(w_n14097_0[0]),.dinb(w_n1039_18[0]),.dout(n14106),.clk(gclk));
	jand g13821(.dina(n14106),.dinb(w_n14099_0[0]),.dout(n14107),.clk(gclk));
	jor g13822(.dina(w_n14107_0[1]),.dinb(w_n14105_0[1]),.dout(n14108),.clk(gclk));
	jand g13823(.dina(w_n14108_0[1]),.dinb(w_n14101_0[1]),.dout(n14109),.clk(gclk));
	jor g13824(.dina(w_n14109_0[1]),.dinb(w_n1034_16[1]),.dout(n14110),.clk(gclk));
	jxor g13825(.dina(w_n13563_0[0]),.dinb(w_n1039_17[2]),.dout(n14111),.clk(gclk));
	jor g13826(.dina(n14111),.dinb(w_n13723_14[2]),.dout(n14112),.clk(gclk));
	jxor g13827(.dina(n14112),.dinb(w_n13574_0[0]),.dout(n14113),.clk(gclk));
	jand g13828(.dina(w_n14109_0[0]),.dinb(w_n1034_16[0]),.dout(n14114),.clk(gclk));
	jor g13829(.dina(w_n14114_0[1]),.dinb(w_n14113_0[1]),.dout(n14115),.clk(gclk));
	jand g13830(.dina(w_n14115_0[2]),.dinb(w_n14110_0[2]),.dout(n14116),.clk(gclk));
	jor g13831(.dina(n14116),.dinb(w_n796_18[0]),.dout(n14117),.clk(gclk));
	jnot g13832(.din(w_n13579_0[0]),.dout(n14118),.clk(gclk));
	jor g13833(.dina(n14118),.dinb(w_n13577_0[0]),.dout(n14119),.clk(gclk));
	jor g13834(.dina(n14119),.dinb(w_n13723_14[1]),.dout(n14120),.clk(gclk));
	jxor g13835(.dina(n14120),.dinb(w_n13588_0[0]),.dout(n14121),.clk(gclk));
	jand g13836(.dina(w_n14110_0[1]),.dinb(w_n796_17[2]),.dout(n14122),.clk(gclk));
	jand g13837(.dina(n14122),.dinb(w_n14115_0[1]),.dout(n14123),.clk(gclk));
	jor g13838(.dina(w_n14123_0[1]),.dinb(w_n14121_0[1]),.dout(n14124),.clk(gclk));
	jand g13839(.dina(w_n14124_0[1]),.dinb(w_n14117_0[1]),.dout(n14125),.clk(gclk));
	jor g13840(.dina(w_n14125_0[2]),.dinb(w_n791_16[2]),.dout(n14126),.clk(gclk));
	jand g13841(.dina(w_n14125_0[1]),.dinb(w_n791_16[1]),.dout(n14127),.clk(gclk));
	jnot g13842(.din(w_n13591_0[0]),.dout(n14128),.clk(gclk));
	jand g13843(.dina(w_asqrt13_12[0]),.dinb(n14128),.dout(n14129),.clk(gclk));
	jand g13844(.dina(w_n14129_0[1]),.dinb(w_n13596_0[0]),.dout(n14130),.clk(gclk));
	jor g13845(.dina(n14130),.dinb(w_n13595_0[0]),.dout(n14131),.clk(gclk));
	jand g13846(.dina(w_n14129_0[0]),.dinb(w_n13597_0[0]),.dout(n14132),.clk(gclk));
	jnot g13847(.din(n14132),.dout(n14133),.clk(gclk));
	jand g13848(.dina(n14133),.dinb(n14131),.dout(n14134),.clk(gclk));
	jnot g13849(.din(n14134),.dout(n14135),.clk(gclk));
	jor g13850(.dina(w_n14135_0[1]),.dinb(n14127),.dout(n14136),.clk(gclk));
	jand g13851(.dina(w_n14136_0[1]),.dinb(w_n14126_0[1]),.dout(n14137),.clk(gclk));
	jor g13852(.dina(n14137),.dinb(w_n595_18[2]),.dout(n14138),.clk(gclk));
	jand g13853(.dina(w_n14126_0[0]),.dinb(w_n595_18[1]),.dout(n14139),.clk(gclk));
	jand g13854(.dina(n14139),.dinb(w_n14136_0[0]),.dout(n14140),.clk(gclk));
	jnot g13855(.din(w_n13599_0[0]),.dout(n14141),.clk(gclk));
	jand g13856(.dina(w_asqrt13_11[2]),.dinb(n14141),.dout(n14142),.clk(gclk));
	jand g13857(.dina(w_n14142_0[1]),.dinb(w_n13606_0[0]),.dout(n14143),.clk(gclk));
	jor g13858(.dina(n14143),.dinb(w_n13604_0[0]),.dout(n14144),.clk(gclk));
	jand g13859(.dina(w_n14142_0[0]),.dinb(w_n13607_0[0]),.dout(n14145),.clk(gclk));
	jnot g13860(.din(n14145),.dout(n14146),.clk(gclk));
	jand g13861(.dina(n14146),.dinb(n14144),.dout(n14147),.clk(gclk));
	jnot g13862(.din(n14147),.dout(n14148),.clk(gclk));
	jor g13863(.dina(w_n14148_0[1]),.dinb(w_n14140_0[1]),.dout(n14149),.clk(gclk));
	jand g13864(.dina(n14149),.dinb(w_n14138_0[1]),.dout(n14150),.clk(gclk));
	jor g13865(.dina(w_n14150_0[1]),.dinb(w_n590_17[0]),.dout(n14151),.clk(gclk));
	jxor g13866(.dina(w_n13608_0[0]),.dinb(w_n595_18[0]),.dout(n14152),.clk(gclk));
	jor g13867(.dina(n14152),.dinb(w_n13723_14[0]),.dout(n14153),.clk(gclk));
	jxor g13868(.dina(n14153),.dinb(w_n13619_0[0]),.dout(n14154),.clk(gclk));
	jand g13869(.dina(w_n14150_0[0]),.dinb(w_n590_16[2]),.dout(n14155),.clk(gclk));
	jor g13870(.dina(w_n14155_0[1]),.dinb(w_n14154_0[1]),.dout(n14156),.clk(gclk));
	jand g13871(.dina(w_n14156_0[2]),.dinb(w_n14151_0[2]),.dout(n14157),.clk(gclk));
	jor g13872(.dina(n14157),.dinb(w_n430_18[1]),.dout(n14158),.clk(gclk));
	jnot g13873(.din(w_n13624_0[0]),.dout(n14159),.clk(gclk));
	jor g13874(.dina(n14159),.dinb(w_n13622_0[0]),.dout(n14160),.clk(gclk));
	jor g13875(.dina(n14160),.dinb(w_n13723_13[2]),.dout(n14161),.clk(gclk));
	jxor g13876(.dina(n14161),.dinb(w_n13633_0[0]),.dout(n14162),.clk(gclk));
	jand g13877(.dina(w_n14151_0[1]),.dinb(w_n430_18[0]),.dout(n14163),.clk(gclk));
	jand g13878(.dina(n14163),.dinb(w_n14156_0[1]),.dout(n14164),.clk(gclk));
	jor g13879(.dina(w_n14164_0[1]),.dinb(w_n14162_0[1]),.dout(n14165),.clk(gclk));
	jand g13880(.dina(w_n14165_0[1]),.dinb(w_n14158_0[1]),.dout(n14166),.clk(gclk));
	jor g13881(.dina(w_n14166_0[2]),.dinb(w_n425_17[1]),.dout(n14167),.clk(gclk));
	jand g13882(.dina(w_n14166_0[1]),.dinb(w_n425_17[0]),.dout(n14168),.clk(gclk));
	jnot g13883(.din(w_n13636_0[0]),.dout(n14169),.clk(gclk));
	jand g13884(.dina(w_asqrt13_11[1]),.dinb(n14169),.dout(n14170),.clk(gclk));
	jand g13885(.dina(w_n14170_0[1]),.dinb(w_n13641_0[0]),.dout(n14171),.clk(gclk));
	jor g13886(.dina(n14171),.dinb(w_n13640_0[0]),.dout(n14172),.clk(gclk));
	jand g13887(.dina(w_n14170_0[0]),.dinb(w_n13642_0[0]),.dout(n14173),.clk(gclk));
	jnot g13888(.din(n14173),.dout(n14174),.clk(gclk));
	jand g13889(.dina(n14174),.dinb(n14172),.dout(n14175),.clk(gclk));
	jnot g13890(.din(n14175),.dout(n14176),.clk(gclk));
	jor g13891(.dina(w_n14176_0[1]),.dinb(n14168),.dout(n14177),.clk(gclk));
	jand g13892(.dina(w_n14177_0[1]),.dinb(w_n14167_0[1]),.dout(n14178),.clk(gclk));
	jor g13893(.dina(n14178),.dinb(w_n305_19[0]),.dout(n14179),.clk(gclk));
	jand g13894(.dina(w_n14167_0[0]),.dinb(w_n305_18[2]),.dout(n14180),.clk(gclk));
	jand g13895(.dina(n14180),.dinb(w_n14177_0[0]),.dout(n14181),.clk(gclk));
	jnot g13896(.din(w_n13644_0[0]),.dout(n14182),.clk(gclk));
	jand g13897(.dina(w_asqrt13_11[0]),.dinb(n14182),.dout(n14183),.clk(gclk));
	jand g13898(.dina(w_n14183_0[1]),.dinb(w_n13651_0[0]),.dout(n14184),.clk(gclk));
	jor g13899(.dina(n14184),.dinb(w_n13649_0[0]),.dout(n14185),.clk(gclk));
	jand g13900(.dina(w_n14183_0[0]),.dinb(w_n13652_0[0]),.dout(n14186),.clk(gclk));
	jnot g13901(.din(n14186),.dout(n14187),.clk(gclk));
	jand g13902(.dina(n14187),.dinb(n14185),.dout(n14188),.clk(gclk));
	jnot g13903(.din(n14188),.dout(n14189),.clk(gclk));
	jor g13904(.dina(w_n14189_0[1]),.dinb(w_n14181_0[1]),.dout(n14190),.clk(gclk));
	jand g13905(.dina(n14190),.dinb(w_n14179_0[1]),.dout(n14191),.clk(gclk));
	jor g13906(.dina(w_n14191_0[1]),.dinb(w_n290_18[1]),.dout(n14192),.clk(gclk));
	jxor g13907(.dina(w_n13653_0[0]),.dinb(w_n305_18[1]),.dout(n14193),.clk(gclk));
	jor g13908(.dina(n14193),.dinb(w_n13723_13[1]),.dout(n14194),.clk(gclk));
	jxor g13909(.dina(n14194),.dinb(w_n13664_0[0]),.dout(n14195),.clk(gclk));
	jand g13910(.dina(w_n14191_0[0]),.dinb(w_n290_18[0]),.dout(n14196),.clk(gclk));
	jor g13911(.dina(w_n14196_0[1]),.dinb(w_n14195_0[1]),.dout(n14197),.clk(gclk));
	jand g13912(.dina(w_n14197_0[2]),.dinb(w_n14192_0[2]),.dout(n14198),.clk(gclk));
	jor g13913(.dina(n14198),.dinb(w_n223_18[2]),.dout(n14199),.clk(gclk));
	jnot g13914(.din(w_n13669_0[0]),.dout(n14200),.clk(gclk));
	jor g13915(.dina(n14200),.dinb(w_n13667_0[0]),.dout(n14201),.clk(gclk));
	jor g13916(.dina(n14201),.dinb(w_n13723_13[0]),.dout(n14202),.clk(gclk));
	jxor g13917(.dina(n14202),.dinb(w_n13678_0[0]),.dout(n14203),.clk(gclk));
	jand g13918(.dina(w_n14192_0[1]),.dinb(w_n223_18[1]),.dout(n14204),.clk(gclk));
	jand g13919(.dina(n14204),.dinb(w_n14197_0[1]),.dout(n14205),.clk(gclk));
	jor g13920(.dina(w_n14205_0[1]),.dinb(w_n14203_0[1]),.dout(n14206),.clk(gclk));
	jand g13921(.dina(w_n14206_0[1]),.dinb(w_n14199_0[1]),.dout(n14207),.clk(gclk));
	jor g13922(.dina(w_n14207_0[2]),.dinb(w_n199_21[1]),.dout(n14208),.clk(gclk));
	jand g13923(.dina(w_n14207_0[1]),.dinb(w_n199_21[0]),.dout(n14209),.clk(gclk));
	jnot g13924(.din(w_n13681_0[0]),.dout(n14210),.clk(gclk));
	jand g13925(.dina(w_asqrt13_10[2]),.dinb(n14210),.dout(n14211),.clk(gclk));
	jand g13926(.dina(w_n14211_0[1]),.dinb(w_n13686_0[0]),.dout(n14212),.clk(gclk));
	jor g13927(.dina(n14212),.dinb(w_n13685_0[0]),.dout(n14213),.clk(gclk));
	jand g13928(.dina(w_n14211_0[0]),.dinb(w_n13687_0[0]),.dout(n14214),.clk(gclk));
	jnot g13929(.din(n14214),.dout(n14215),.clk(gclk));
	jand g13930(.dina(n14215),.dinb(n14213),.dout(n14216),.clk(gclk));
	jnot g13931(.din(n14216),.dout(n14217),.clk(gclk));
	jor g13932(.dina(w_n14217_0[1]),.dinb(n14209),.dout(n14218),.clk(gclk));
	jand g13933(.dina(n14218),.dinb(n14208),.dout(n14219),.clk(gclk));
	jnot g13934(.din(w_n13689_0[0]),.dout(n14220),.clk(gclk));
	jand g13935(.dina(w_asqrt13_10[1]),.dinb(n14220),.dout(n14221),.clk(gclk));
	jand g13936(.dina(w_n14221_0[1]),.dinb(w_n13696_0[0]),.dout(n14222),.clk(gclk));
	jor g13937(.dina(n14222),.dinb(w_n13694_0[0]),.dout(n14223),.clk(gclk));
	jand g13938(.dina(w_n14221_0[0]),.dinb(w_n13697_0[0]),.dout(n14224),.clk(gclk));
	jnot g13939(.din(n14224),.dout(n14225),.clk(gclk));
	jand g13940(.dina(n14225),.dinb(n14223),.dout(n14226),.clk(gclk));
	jnot g13941(.din(w_n14226_0[2]),.dout(n14227),.clk(gclk));
	jand g13942(.dina(w_asqrt13_10[0]),.dinb(w_n13711_0[1]),.dout(n14228),.clk(gclk));
	jand g13943(.dina(w_n14228_0[1]),.dinb(w_n13698_1[0]),.dout(n14229),.clk(gclk));
	jor g13944(.dina(n14229),.dinb(w_n13745_0[0]),.dout(n14230),.clk(gclk));
	jor g13945(.dina(n14230),.dinb(w_n14227_0[1]),.dout(n14231),.clk(gclk));
	jor g13946(.dina(n14231),.dinb(w_n14219_0[2]),.dout(n14232),.clk(gclk));
	jand g13947(.dina(n14232),.dinb(w_n194_20[1]),.dout(n14233),.clk(gclk));
	jand g13948(.dina(w_n14227_0[0]),.dinb(w_n14219_0[1]),.dout(n14234),.clk(gclk));
	jor g13949(.dina(w_n14228_0[0]),.dinb(w_n13698_0[2]),.dout(n14235),.clk(gclk));
	jand g13950(.dina(w_n13711_0[0]),.dinb(w_n13698_0[1]),.dout(n14236),.clk(gclk));
	jor g13951(.dina(n14236),.dinb(w_n194_20[0]),.dout(n14237),.clk(gclk));
	jnot g13952(.din(n14237),.dout(n14238),.clk(gclk));
	jand g13953(.dina(n14238),.dinb(n14235),.dout(n14239),.clk(gclk));
	jor g13954(.dina(w_n14239_0[1]),.dinb(w_n14234_0[2]),.dout(n14242),.clk(gclk));
	jor g13955(.dina(n14242),.dinb(w_n14233_0[1]),.dout(asqrt_fa_13),.clk(gclk));
	jxor g13956(.dina(w_n14096_0[0]),.dinb(w_n1312_15[0]),.dout(n14244),.clk(gclk));
	jand g13957(.dina(n14244),.dinb(w_asqrt12_31),.dout(n14245),.clk(gclk));
	jxor g13958(.dina(n14245),.dinb(w_n13726_0[0]),.dout(n14246),.clk(gclk));
	jand g13959(.dina(w_asqrt12_30[2]),.dinb(w_a24_0[0]),.dout(n14247),.clk(gclk));
	jnot g13960(.din(w_a22_0[1]),.dout(n14248),.clk(gclk));
	jnot g13961(.din(w_a23_0[1]),.dout(n14249),.clk(gclk));
	jand g13962(.dina(w_n13728_1[0]),.dinb(w_n14249_0[1]),.dout(n14250),.clk(gclk));
	jand g13963(.dina(n14250),.dinb(w_n14248_1[1]),.dout(n14251),.clk(gclk));
	jor g13964(.dina(n14251),.dinb(n14247),.dout(n14252),.clk(gclk));
	jand g13965(.dina(w_n14252_0[2]),.dinb(w_asqrt13_9[2]),.dout(n14253),.clk(gclk));
	jand g13966(.dina(w_asqrt12_30[1]),.dinb(w_n13728_0[2]),.dout(n14254),.clk(gclk));
	jxor g13967(.dina(w_n14254_0[1]),.dinb(w_n13729_0[1]),.dout(n14255),.clk(gclk));
	jor g13968(.dina(w_n14252_0[1]),.dinb(w_asqrt13_9[1]),.dout(n14256),.clk(gclk));
	jand g13969(.dina(n14256),.dinb(w_n14255_0[1]),.dout(n14257),.clk(gclk));
	jor g13970(.dina(w_n14257_0[1]),.dinb(w_n14253_0[1]),.dout(n14258),.clk(gclk));
	jand g13971(.dina(n14258),.dinb(w_asqrt14_14[0]),.dout(n14259),.clk(gclk));
	jor g13972(.dina(w_n14253_0[0]),.dinb(w_asqrt14_13[2]),.dout(n14260),.clk(gclk));
	jor g13973(.dina(n14260),.dinb(w_n14257_0[0]),.dout(n14261),.clk(gclk));
	jand g13974(.dina(w_n14254_0[0]),.dinb(w_n13729_0[0]),.dout(n14262),.clk(gclk));
	jnot g13975(.din(w_n14233_0[0]),.dout(n14263),.clk(gclk));
	jnot g13976(.din(w_n14234_0[1]),.dout(n14264),.clk(gclk));
	jnot g13977(.din(w_n14239_0[0]),.dout(n14265),.clk(gclk));
	jand g13978(.dina(n14265),.dinb(w_asqrt13_9[0]),.dout(n14266),.clk(gclk));
	jand g13979(.dina(n14266),.dinb(n14264),.dout(n14267),.clk(gclk));
	jand g13980(.dina(n14267),.dinb(n14263),.dout(n14268),.clk(gclk));
	jor g13981(.dina(n14268),.dinb(n14262),.dout(n14269),.clk(gclk));
	jxor g13982(.dina(n14269),.dinb(w_n13177_0[1]),.dout(n14270),.clk(gclk));
	jand g13983(.dina(w_n14270_0[1]),.dinb(w_n14261_0[1]),.dout(n14271),.clk(gclk));
	jor g13984(.dina(n14271),.dinb(w_n14259_0[1]),.dout(n14272),.clk(gclk));
	jand g13985(.dina(w_n14272_0[2]),.dinb(w_asqrt15_9[1]),.dout(n14273),.clk(gclk));
	jor g13986(.dina(w_n14272_0[1]),.dinb(w_asqrt15_9[0]),.dout(n14274),.clk(gclk));
	jxor g13987(.dina(w_n13733_0[0]),.dinb(w_n13718_8[1]),.dout(n14275),.clk(gclk));
	jand g13988(.dina(n14275),.dinb(w_asqrt12_30[0]),.dout(n14276),.clk(gclk));
	jxor g13989(.dina(n14276),.dinb(w_n13736_0[0]),.dout(n14277),.clk(gclk));
	jnot g13990(.din(w_n14277_0[1]),.dout(n14278),.clk(gclk));
	jand g13991(.dina(n14278),.dinb(n14274),.dout(n14279),.clk(gclk));
	jor g13992(.dina(w_n14279_0[1]),.dinb(w_n14273_0[1]),.dout(n14280),.clk(gclk));
	jand g13993(.dina(n14280),.dinb(w_asqrt16_14[0]),.dout(n14281),.clk(gclk));
	jnot g13994(.din(w_n13742_0[0]),.dout(n14282),.clk(gclk));
	jand g13995(.dina(n14282),.dinb(w_n13740_0[0]),.dout(n14283),.clk(gclk));
	jand g13996(.dina(n14283),.dinb(w_asqrt12_29[2]),.dout(n14284),.clk(gclk));
	jxor g13997(.dina(n14284),.dinb(w_n13750_0[0]),.dout(n14285),.clk(gclk));
	jnot g13998(.din(n14285),.dout(n14286),.clk(gclk));
	jor g13999(.dina(w_n14273_0[0]),.dinb(w_asqrt16_13[2]),.dout(n14287),.clk(gclk));
	jor g14000(.dina(n14287),.dinb(w_n14279_0[0]),.dout(n14288),.clk(gclk));
	jand g14001(.dina(w_n14288_0[1]),.dinb(w_n14286_0[1]),.dout(n14289),.clk(gclk));
	jor g14002(.dina(w_n14289_0[1]),.dinb(w_n14281_0[1]),.dout(n14290),.clk(gclk));
	jand g14003(.dina(w_n14290_0[2]),.dinb(w_asqrt17_9[2]),.dout(n14291),.clk(gclk));
	jor g14004(.dina(w_n14290_0[1]),.dinb(w_asqrt17_9[1]),.dout(n14292),.clk(gclk));
	jnot g14005(.din(w_n13757_0[0]),.dout(n14293),.clk(gclk));
	jxor g14006(.dina(w_n13752_0[0]),.dinb(w_n12670_8[2]),.dout(n14294),.clk(gclk));
	jand g14007(.dina(n14294),.dinb(w_asqrt12_29[1]),.dout(n14295),.clk(gclk));
	jxor g14008(.dina(n14295),.dinb(n14293),.dout(n14296),.clk(gclk));
	jand g14009(.dina(w_n14296_0[1]),.dinb(n14292),.dout(n14297),.clk(gclk));
	jor g14010(.dina(w_n14297_0[1]),.dinb(w_n14291_0[1]),.dout(n14298),.clk(gclk));
	jand g14011(.dina(n14298),.dinb(w_asqrt18_14[0]),.dout(n14299),.clk(gclk));
	jor g14012(.dina(w_n14291_0[0]),.dinb(w_asqrt18_13[2]),.dout(n14300),.clk(gclk));
	jor g14013(.dina(n14300),.dinb(w_n14297_0[0]),.dout(n14301),.clk(gclk));
	jnot g14014(.din(w_n13764_0[0]),.dout(n14302),.clk(gclk));
	jnot g14015(.din(w_n13766_0[0]),.dout(n14303),.clk(gclk));
	jand g14016(.dina(w_asqrt12_29[0]),.dinb(w_n13760_0[0]),.dout(n14304),.clk(gclk));
	jand g14017(.dina(w_n14304_0[1]),.dinb(n14303),.dout(n14305),.clk(gclk));
	jor g14018(.dina(n14305),.dinb(n14302),.dout(n14306),.clk(gclk));
	jnot g14019(.din(w_n13767_0[0]),.dout(n14307),.clk(gclk));
	jand g14020(.dina(w_n14304_0[0]),.dinb(n14307),.dout(n14308),.clk(gclk));
	jnot g14021(.din(n14308),.dout(n14309),.clk(gclk));
	jand g14022(.dina(n14309),.dinb(n14306),.dout(n14310),.clk(gclk));
	jand g14023(.dina(w_n14310_0[1]),.dinb(w_n14301_0[1]),.dout(n14311),.clk(gclk));
	jor g14024(.dina(n14311),.dinb(w_n14299_0[1]),.dout(n14312),.clk(gclk));
	jand g14025(.dina(w_n14312_0[2]),.dinb(w_asqrt19_9[2]),.dout(n14313),.clk(gclk));
	jor g14026(.dina(w_n14312_0[1]),.dinb(w_asqrt19_9[1]),.dout(n14314),.clk(gclk));
	jxor g14027(.dina(w_n13768_0[0]),.dinb(w_n11657_8[2]),.dout(n14315),.clk(gclk));
	jand g14028(.dina(n14315),.dinb(w_asqrt12_28[2]),.dout(n14316),.clk(gclk));
	jxor g14029(.dina(n14316),.dinb(w_n13773_0[0]),.dout(n14317),.clk(gclk));
	jand g14030(.dina(w_n14317_0[1]),.dinb(n14314),.dout(n14318),.clk(gclk));
	jor g14031(.dina(w_n14318_0[1]),.dinb(w_n14313_0[1]),.dout(n14319),.clk(gclk));
	jand g14032(.dina(n14319),.dinb(w_asqrt20_14[0]),.dout(n14320),.clk(gclk));
	jnot g14033(.din(w_n13779_0[0]),.dout(n14321),.clk(gclk));
	jand g14034(.dina(n14321),.dinb(w_n13777_0[0]),.dout(n14322),.clk(gclk));
	jand g14035(.dina(n14322),.dinb(w_asqrt12_28[1]),.dout(n14323),.clk(gclk));
	jxor g14036(.dina(n14323),.dinb(w_n13788_0[0]),.dout(n14324),.clk(gclk));
	jnot g14037(.din(n14324),.dout(n14325),.clk(gclk));
	jor g14038(.dina(w_n14313_0[0]),.dinb(w_asqrt20_13[2]),.dout(n14326),.clk(gclk));
	jor g14039(.dina(n14326),.dinb(w_n14318_0[0]),.dout(n14327),.clk(gclk));
	jand g14040(.dina(w_n14327_0[1]),.dinb(w_n14325_0[1]),.dout(n14328),.clk(gclk));
	jor g14041(.dina(w_n14328_0[1]),.dinb(w_n14320_0[1]),.dout(n14329),.clk(gclk));
	jand g14042(.dina(w_n14329_0[2]),.dinb(w_asqrt21_10[0]),.dout(n14330),.clk(gclk));
	jor g14043(.dina(w_n14329_0[1]),.dinb(w_asqrt21_9[2]),.dout(n14331),.clk(gclk));
	jxor g14044(.dina(w_n13790_0[0]),.dinb(w_n10696_9[1]),.dout(n14332),.clk(gclk));
	jand g14045(.dina(n14332),.dinb(w_asqrt12_28[0]),.dout(n14333),.clk(gclk));
	jxor g14046(.dina(n14333),.dinb(w_n13796_0[0]),.dout(n14334),.clk(gclk));
	jand g14047(.dina(w_n14334_0[1]),.dinb(n14331),.dout(n14335),.clk(gclk));
	jor g14048(.dina(w_n14335_0[1]),.dinb(w_n14330_0[1]),.dout(n14336),.clk(gclk));
	jand g14049(.dina(n14336),.dinb(w_asqrt22_14[0]),.dout(n14337),.clk(gclk));
	jor g14050(.dina(w_n14330_0[0]),.dinb(w_asqrt22_13[2]),.dout(n14338),.clk(gclk));
	jor g14051(.dina(n14338),.dinb(w_n14335_0[0]),.dout(n14339),.clk(gclk));
	jnot g14052(.din(w_n13804_0[0]),.dout(n14340),.clk(gclk));
	jnot g14053(.din(w_n13806_0[0]),.dout(n14341),.clk(gclk));
	jand g14054(.dina(w_asqrt12_27[2]),.dinb(w_n13800_0[0]),.dout(n14342),.clk(gclk));
	jand g14055(.dina(w_n14342_0[1]),.dinb(n14341),.dout(n14343),.clk(gclk));
	jor g14056(.dina(n14343),.dinb(n14340),.dout(n14344),.clk(gclk));
	jnot g14057(.din(w_n13807_0[0]),.dout(n14345),.clk(gclk));
	jand g14058(.dina(w_n14342_0[0]),.dinb(n14345),.dout(n14346),.clk(gclk));
	jnot g14059(.din(n14346),.dout(n14347),.clk(gclk));
	jand g14060(.dina(n14347),.dinb(n14344),.dout(n14348),.clk(gclk));
	jand g14061(.dina(w_n14348_0[1]),.dinb(w_n14339_0[1]),.dout(n14349),.clk(gclk));
	jor g14062(.dina(n14349),.dinb(w_n14337_0[1]),.dout(n14350),.clk(gclk));
	jand g14063(.dina(w_n14350_0[1]),.dinb(w_asqrt23_10[0]),.dout(n14351),.clk(gclk));
	jxor g14064(.dina(w_n13808_0[0]),.dinb(w_n9769_9[1]),.dout(n14352),.clk(gclk));
	jand g14065(.dina(n14352),.dinb(w_asqrt12_27[1]),.dout(n14353),.clk(gclk));
	jxor g14066(.dina(n14353),.dinb(w_n13815_0[0]),.dout(n14354),.clk(gclk));
	jnot g14067(.din(n14354),.dout(n14355),.clk(gclk));
	jor g14068(.dina(w_n14350_0[0]),.dinb(w_asqrt23_9[2]),.dout(n14356),.clk(gclk));
	jand g14069(.dina(w_n14356_0[1]),.dinb(w_n14355_0[1]),.dout(n14357),.clk(gclk));
	jor g14070(.dina(w_n14357_0[2]),.dinb(w_n14351_0[2]),.dout(n14358),.clk(gclk));
	jand g14071(.dina(n14358),.dinb(w_asqrt24_14[0]),.dout(n14359),.clk(gclk));
	jnot g14072(.din(w_n13820_0[0]),.dout(n14360),.clk(gclk));
	jand g14073(.dina(n14360),.dinb(w_n13818_0[0]),.dout(n14361),.clk(gclk));
	jand g14074(.dina(n14361),.dinb(w_asqrt12_27[0]),.dout(n14362),.clk(gclk));
	jxor g14075(.dina(n14362),.dinb(w_n13828_0[0]),.dout(n14363),.clk(gclk));
	jnot g14076(.din(n14363),.dout(n14364),.clk(gclk));
	jor g14077(.dina(w_n14351_0[1]),.dinb(w_asqrt24_13[2]),.dout(n14365),.clk(gclk));
	jor g14078(.dina(n14365),.dinb(w_n14357_0[1]),.dout(n14366),.clk(gclk));
	jand g14079(.dina(w_n14366_0[1]),.dinb(w_n14364_0[1]),.dout(n14367),.clk(gclk));
	jor g14080(.dina(w_n14367_0[1]),.dinb(w_n14359_0[1]),.dout(n14368),.clk(gclk));
	jand g14081(.dina(w_n14368_0[2]),.dinb(w_asqrt25_10[1]),.dout(n14369),.clk(gclk));
	jor g14082(.dina(w_n14368_0[1]),.dinb(w_asqrt25_10[0]),.dout(n14370),.clk(gclk));
	jnot g14083(.din(w_n13834_0[0]),.dout(n14371),.clk(gclk));
	jnot g14084(.din(w_n13835_0[0]),.dout(n14372),.clk(gclk));
	jand g14085(.dina(w_asqrt12_26[2]),.dinb(w_n13831_0[0]),.dout(n14373),.clk(gclk));
	jand g14086(.dina(w_n14373_0[1]),.dinb(n14372),.dout(n14374),.clk(gclk));
	jor g14087(.dina(n14374),.dinb(n14371),.dout(n14375),.clk(gclk));
	jnot g14088(.din(w_n13836_0[0]),.dout(n14376),.clk(gclk));
	jand g14089(.dina(w_n14373_0[0]),.dinb(n14376),.dout(n14377),.clk(gclk));
	jnot g14090(.din(n14377),.dout(n14378),.clk(gclk));
	jand g14091(.dina(n14378),.dinb(n14375),.dout(n14379),.clk(gclk));
	jand g14092(.dina(w_n14379_0[1]),.dinb(n14370),.dout(n14380),.clk(gclk));
	jor g14093(.dina(w_n14380_0[1]),.dinb(w_n14369_0[1]),.dout(n14381),.clk(gclk));
	jand g14094(.dina(n14381),.dinb(w_asqrt26_14[0]),.dout(n14382),.clk(gclk));
	jor g14095(.dina(w_n14369_0[0]),.dinb(w_asqrt26_13[2]),.dout(n14383),.clk(gclk));
	jor g14096(.dina(n14383),.dinb(w_n14380_0[0]),.dout(n14384),.clk(gclk));
	jnot g14097(.din(w_n13842_0[0]),.dout(n14385),.clk(gclk));
	jnot g14098(.din(w_n13844_0[0]),.dout(n14386),.clk(gclk));
	jand g14099(.dina(w_asqrt12_26[1]),.dinb(w_n13838_0[0]),.dout(n14387),.clk(gclk));
	jand g14100(.dina(w_n14387_0[1]),.dinb(n14386),.dout(n14388),.clk(gclk));
	jor g14101(.dina(n14388),.dinb(n14385),.dout(n14389),.clk(gclk));
	jnot g14102(.din(w_n13845_0[0]),.dout(n14390),.clk(gclk));
	jand g14103(.dina(w_n14387_0[0]),.dinb(n14390),.dout(n14391),.clk(gclk));
	jnot g14104(.din(n14391),.dout(n14392),.clk(gclk));
	jand g14105(.dina(n14392),.dinb(n14389),.dout(n14393),.clk(gclk));
	jand g14106(.dina(w_n14393_0[1]),.dinb(w_n14384_0[1]),.dout(n14394),.clk(gclk));
	jor g14107(.dina(n14394),.dinb(w_n14382_0[1]),.dout(n14395),.clk(gclk));
	jand g14108(.dina(w_n14395_0[1]),.dinb(w_asqrt27_10[1]),.dout(n14396),.clk(gclk));
	jxor g14109(.dina(w_n13846_0[0]),.dinb(w_n8053_10[0]),.dout(n14397),.clk(gclk));
	jand g14110(.dina(n14397),.dinb(w_asqrt12_26[0]),.dout(n14398),.clk(gclk));
	jxor g14111(.dina(n14398),.dinb(w_n13856_0[0]),.dout(n14399),.clk(gclk));
	jnot g14112(.din(n14399),.dout(n14400),.clk(gclk));
	jor g14113(.dina(w_n14395_0[0]),.dinb(w_asqrt27_10[0]),.dout(n14401),.clk(gclk));
	jand g14114(.dina(w_n14401_0[1]),.dinb(w_n14400_0[1]),.dout(n14402),.clk(gclk));
	jor g14115(.dina(w_n14402_0[2]),.dinb(w_n14396_0[2]),.dout(n14403),.clk(gclk));
	jand g14116(.dina(n14403),.dinb(w_asqrt28_14[0]),.dout(n14404),.clk(gclk));
	jnot g14117(.din(w_n13861_0[0]),.dout(n14405),.clk(gclk));
	jand g14118(.dina(n14405),.dinb(w_n13859_0[0]),.dout(n14406),.clk(gclk));
	jand g14119(.dina(n14406),.dinb(w_asqrt12_25[2]),.dout(n14407),.clk(gclk));
	jxor g14120(.dina(n14407),.dinb(w_n13869_0[0]),.dout(n14408),.clk(gclk));
	jnot g14121(.din(n14408),.dout(n14409),.clk(gclk));
	jor g14122(.dina(w_n14396_0[1]),.dinb(w_asqrt28_13[2]),.dout(n14410),.clk(gclk));
	jor g14123(.dina(n14410),.dinb(w_n14402_0[1]),.dout(n14411),.clk(gclk));
	jand g14124(.dina(w_n14411_0[1]),.dinb(w_n14409_0[1]),.dout(n14412),.clk(gclk));
	jor g14125(.dina(w_n14412_0[1]),.dinb(w_n14404_0[1]),.dout(n14413),.clk(gclk));
	jand g14126(.dina(w_n14413_0[2]),.dinb(w_asqrt29_10[2]),.dout(n14414),.clk(gclk));
	jor g14127(.dina(w_n14413_0[1]),.dinb(w_asqrt29_10[1]),.dout(n14415),.clk(gclk));
	jnot g14128(.din(w_n13875_0[0]),.dout(n14416),.clk(gclk));
	jnot g14129(.din(w_n13876_0[0]),.dout(n14417),.clk(gclk));
	jand g14130(.dina(w_asqrt12_25[1]),.dinb(w_n13872_0[0]),.dout(n14418),.clk(gclk));
	jand g14131(.dina(w_n14418_0[1]),.dinb(n14417),.dout(n14419),.clk(gclk));
	jor g14132(.dina(n14419),.dinb(n14416),.dout(n14420),.clk(gclk));
	jnot g14133(.din(w_n13877_0[0]),.dout(n14421),.clk(gclk));
	jand g14134(.dina(w_n14418_0[0]),.dinb(n14421),.dout(n14422),.clk(gclk));
	jnot g14135(.din(n14422),.dout(n14423),.clk(gclk));
	jand g14136(.dina(n14423),.dinb(n14420),.dout(n14424),.clk(gclk));
	jand g14137(.dina(w_n14424_0[1]),.dinb(n14415),.dout(n14425),.clk(gclk));
	jor g14138(.dina(w_n14425_0[1]),.dinb(w_n14414_0[1]),.dout(n14426),.clk(gclk));
	jand g14139(.dina(n14426),.dinb(w_asqrt30_14[0]),.dout(n14427),.clk(gclk));
	jor g14140(.dina(w_n14414_0[0]),.dinb(w_asqrt30_13[2]),.dout(n14428),.clk(gclk));
	jor g14141(.dina(n14428),.dinb(w_n14425_0[0]),.dout(n14429),.clk(gclk));
	jnot g14142(.din(w_n13883_0[0]),.dout(n14430),.clk(gclk));
	jnot g14143(.din(w_n13885_0[0]),.dout(n14431),.clk(gclk));
	jand g14144(.dina(w_asqrt12_25[0]),.dinb(w_n13879_0[0]),.dout(n14432),.clk(gclk));
	jand g14145(.dina(w_n14432_0[1]),.dinb(n14431),.dout(n14433),.clk(gclk));
	jor g14146(.dina(n14433),.dinb(n14430),.dout(n14434),.clk(gclk));
	jnot g14147(.din(w_n13886_0[0]),.dout(n14435),.clk(gclk));
	jand g14148(.dina(w_n14432_0[0]),.dinb(n14435),.dout(n14436),.clk(gclk));
	jnot g14149(.din(n14436),.dout(n14437),.clk(gclk));
	jand g14150(.dina(n14437),.dinb(n14434),.dout(n14438),.clk(gclk));
	jand g14151(.dina(w_n14438_0[1]),.dinb(w_n14429_0[1]),.dout(n14439),.clk(gclk));
	jor g14152(.dina(n14439),.dinb(w_n14427_0[1]),.dout(n14440),.clk(gclk));
	jand g14153(.dina(w_n14440_0[1]),.dinb(w_asqrt31_10[2]),.dout(n14441),.clk(gclk));
	jxor g14154(.dina(w_n13887_0[0]),.dinb(w_n6500_11[0]),.dout(n14442),.clk(gclk));
	jand g14155(.dina(n14442),.dinb(w_asqrt12_24[2]),.dout(n14443),.clk(gclk));
	jxor g14156(.dina(n14443),.dinb(w_n13897_0[0]),.dout(n14444),.clk(gclk));
	jnot g14157(.din(n14444),.dout(n14445),.clk(gclk));
	jor g14158(.dina(w_n14440_0[0]),.dinb(w_asqrt31_10[1]),.dout(n14446),.clk(gclk));
	jand g14159(.dina(w_n14446_0[1]),.dinb(w_n14445_0[1]),.dout(n14447),.clk(gclk));
	jor g14160(.dina(w_n14447_0[2]),.dinb(w_n14441_0[2]),.dout(n14448),.clk(gclk));
	jand g14161(.dina(n14448),.dinb(w_asqrt32_14[0]),.dout(n14449),.clk(gclk));
	jnot g14162(.din(w_n13902_0[0]),.dout(n14450),.clk(gclk));
	jand g14163(.dina(n14450),.dinb(w_n13900_0[0]),.dout(n14451),.clk(gclk));
	jand g14164(.dina(n14451),.dinb(w_asqrt12_24[1]),.dout(n14452),.clk(gclk));
	jxor g14165(.dina(n14452),.dinb(w_n13910_0[0]),.dout(n14453),.clk(gclk));
	jnot g14166(.din(n14453),.dout(n14454),.clk(gclk));
	jor g14167(.dina(w_n14441_0[1]),.dinb(w_asqrt32_13[2]),.dout(n14455),.clk(gclk));
	jor g14168(.dina(n14455),.dinb(w_n14447_0[1]),.dout(n14456),.clk(gclk));
	jand g14169(.dina(w_n14456_0[1]),.dinb(w_n14454_0[1]),.dout(n14457),.clk(gclk));
	jor g14170(.dina(w_n14457_0[1]),.dinb(w_n14449_0[1]),.dout(n14458),.clk(gclk));
	jand g14171(.dina(w_n14458_0[2]),.dinb(w_asqrt33_11[0]),.dout(n14459),.clk(gclk));
	jor g14172(.dina(w_n14458_0[1]),.dinb(w_asqrt33_10[2]),.dout(n14460),.clk(gclk));
	jnot g14173(.din(w_n13916_0[0]),.dout(n14461),.clk(gclk));
	jnot g14174(.din(w_n13917_0[0]),.dout(n14462),.clk(gclk));
	jand g14175(.dina(w_asqrt12_24[0]),.dinb(w_n13913_0[0]),.dout(n14463),.clk(gclk));
	jand g14176(.dina(w_n14463_0[1]),.dinb(n14462),.dout(n14464),.clk(gclk));
	jor g14177(.dina(n14464),.dinb(n14461),.dout(n14465),.clk(gclk));
	jnot g14178(.din(w_n13918_0[0]),.dout(n14466),.clk(gclk));
	jand g14179(.dina(w_n14463_0[0]),.dinb(n14466),.dout(n14467),.clk(gclk));
	jnot g14180(.din(n14467),.dout(n14468),.clk(gclk));
	jand g14181(.dina(n14468),.dinb(n14465),.dout(n14469),.clk(gclk));
	jand g14182(.dina(w_n14469_0[1]),.dinb(n14460),.dout(n14470),.clk(gclk));
	jor g14183(.dina(w_n14470_0[1]),.dinb(w_n14459_0[1]),.dout(n14471),.clk(gclk));
	jand g14184(.dina(n14471),.dinb(w_asqrt34_14[0]),.dout(n14472),.clk(gclk));
	jor g14185(.dina(w_n14459_0[0]),.dinb(w_asqrt34_13[2]),.dout(n14473),.clk(gclk));
	jor g14186(.dina(n14473),.dinb(w_n14470_0[0]),.dout(n14474),.clk(gclk));
	jnot g14187(.din(w_n13924_0[0]),.dout(n14475),.clk(gclk));
	jnot g14188(.din(w_n13926_0[0]),.dout(n14476),.clk(gclk));
	jand g14189(.dina(w_asqrt12_23[2]),.dinb(w_n13920_0[0]),.dout(n14477),.clk(gclk));
	jand g14190(.dina(w_n14477_0[1]),.dinb(n14476),.dout(n14478),.clk(gclk));
	jor g14191(.dina(n14478),.dinb(n14475),.dout(n14479),.clk(gclk));
	jnot g14192(.din(w_n13927_0[0]),.dout(n14480),.clk(gclk));
	jand g14193(.dina(w_n14477_0[0]),.dinb(n14480),.dout(n14481),.clk(gclk));
	jnot g14194(.din(n14481),.dout(n14482),.clk(gclk));
	jand g14195(.dina(n14482),.dinb(n14479),.dout(n14483),.clk(gclk));
	jand g14196(.dina(w_n14483_0[1]),.dinb(w_n14474_0[1]),.dout(n14484),.clk(gclk));
	jor g14197(.dina(n14484),.dinb(w_n14472_0[1]),.dout(n14485),.clk(gclk));
	jand g14198(.dina(w_n14485_0[1]),.dinb(w_asqrt35_11[0]),.dout(n14486),.clk(gclk));
	jxor g14199(.dina(w_n13928_0[0]),.dinb(w_n5116_11[2]),.dout(n14487),.clk(gclk));
	jand g14200(.dina(n14487),.dinb(w_asqrt12_23[1]),.dout(n14488),.clk(gclk));
	jxor g14201(.dina(n14488),.dinb(w_n13938_0[0]),.dout(n14489),.clk(gclk));
	jnot g14202(.din(n14489),.dout(n14490),.clk(gclk));
	jor g14203(.dina(w_n14485_0[0]),.dinb(w_asqrt35_10[2]),.dout(n14491),.clk(gclk));
	jand g14204(.dina(w_n14491_0[1]),.dinb(w_n14490_0[1]),.dout(n14492),.clk(gclk));
	jor g14205(.dina(w_n14492_0[2]),.dinb(w_n14486_0[2]),.dout(n14493),.clk(gclk));
	jand g14206(.dina(n14493),.dinb(w_asqrt36_14[0]),.dout(n14494),.clk(gclk));
	jnot g14207(.din(w_n13943_0[0]),.dout(n14495),.clk(gclk));
	jand g14208(.dina(n14495),.dinb(w_n13941_0[0]),.dout(n14496),.clk(gclk));
	jand g14209(.dina(n14496),.dinb(w_asqrt12_23[0]),.dout(n14497),.clk(gclk));
	jxor g14210(.dina(n14497),.dinb(w_n13951_0[0]),.dout(n14498),.clk(gclk));
	jnot g14211(.din(n14498),.dout(n14499),.clk(gclk));
	jor g14212(.dina(w_n14486_0[1]),.dinb(w_asqrt36_13[2]),.dout(n14500),.clk(gclk));
	jor g14213(.dina(n14500),.dinb(w_n14492_0[1]),.dout(n14501),.clk(gclk));
	jand g14214(.dina(w_n14501_0[1]),.dinb(w_n14499_0[1]),.dout(n14502),.clk(gclk));
	jor g14215(.dina(w_n14502_0[1]),.dinb(w_n14494_0[1]),.dout(n14503),.clk(gclk));
	jand g14216(.dina(w_n14503_0[2]),.dinb(w_asqrt37_11[1]),.dout(n14504),.clk(gclk));
	jor g14217(.dina(w_n14503_0[1]),.dinb(w_asqrt37_11[0]),.dout(n14505),.clk(gclk));
	jnot g14218(.din(w_n13957_0[0]),.dout(n14506),.clk(gclk));
	jnot g14219(.din(w_n13958_0[0]),.dout(n14507),.clk(gclk));
	jand g14220(.dina(w_asqrt12_22[2]),.dinb(w_n13954_0[0]),.dout(n14508),.clk(gclk));
	jand g14221(.dina(w_n14508_0[1]),.dinb(n14507),.dout(n14509),.clk(gclk));
	jor g14222(.dina(n14509),.dinb(n14506),.dout(n14510),.clk(gclk));
	jnot g14223(.din(w_n13959_0[0]),.dout(n14511),.clk(gclk));
	jand g14224(.dina(w_n14508_0[0]),.dinb(n14511),.dout(n14512),.clk(gclk));
	jnot g14225(.din(n14512),.dout(n14513),.clk(gclk));
	jand g14226(.dina(n14513),.dinb(n14510),.dout(n14514),.clk(gclk));
	jand g14227(.dina(w_n14514_0[1]),.dinb(n14505),.dout(n14515),.clk(gclk));
	jor g14228(.dina(w_n14515_0[1]),.dinb(w_n14504_0[1]),.dout(n14516),.clk(gclk));
	jand g14229(.dina(n14516),.dinb(w_asqrt38_14[0]),.dout(n14517),.clk(gclk));
	jor g14230(.dina(w_n14504_0[0]),.dinb(w_asqrt38_13[2]),.dout(n14518),.clk(gclk));
	jor g14231(.dina(n14518),.dinb(w_n14515_0[0]),.dout(n14519),.clk(gclk));
	jnot g14232(.din(w_n13965_0[0]),.dout(n14520),.clk(gclk));
	jnot g14233(.din(w_n13967_0[0]),.dout(n14521),.clk(gclk));
	jand g14234(.dina(w_asqrt12_22[1]),.dinb(w_n13961_0[0]),.dout(n14522),.clk(gclk));
	jand g14235(.dina(w_n14522_0[1]),.dinb(n14521),.dout(n14523),.clk(gclk));
	jor g14236(.dina(n14523),.dinb(n14520),.dout(n14524),.clk(gclk));
	jnot g14237(.din(w_n13968_0[0]),.dout(n14525),.clk(gclk));
	jand g14238(.dina(w_n14522_0[0]),.dinb(n14525),.dout(n14526),.clk(gclk));
	jnot g14239(.din(n14526),.dout(n14527),.clk(gclk));
	jand g14240(.dina(n14527),.dinb(n14524),.dout(n14528),.clk(gclk));
	jand g14241(.dina(w_n14528_0[1]),.dinb(w_n14519_0[1]),.dout(n14529),.clk(gclk));
	jor g14242(.dina(n14529),.dinb(w_n14517_0[1]),.dout(n14530),.clk(gclk));
	jand g14243(.dina(w_n14530_0[1]),.dinb(w_asqrt39_11[1]),.dout(n14531),.clk(gclk));
	jxor g14244(.dina(w_n13969_0[0]),.dinb(w_n3907_12[2]),.dout(n14532),.clk(gclk));
	jand g14245(.dina(n14532),.dinb(w_asqrt12_22[0]),.dout(n14533),.clk(gclk));
	jxor g14246(.dina(n14533),.dinb(w_n13979_0[0]),.dout(n14534),.clk(gclk));
	jnot g14247(.din(n14534),.dout(n14535),.clk(gclk));
	jor g14248(.dina(w_n14530_0[0]),.dinb(w_asqrt39_11[0]),.dout(n14536),.clk(gclk));
	jand g14249(.dina(w_n14536_0[1]),.dinb(w_n14535_0[1]),.dout(n14537),.clk(gclk));
	jor g14250(.dina(w_n14537_0[2]),.dinb(w_n14531_0[2]),.dout(n14538),.clk(gclk));
	jand g14251(.dina(n14538),.dinb(w_asqrt40_14[0]),.dout(n14539),.clk(gclk));
	jnot g14252(.din(w_n13984_0[0]),.dout(n14540),.clk(gclk));
	jand g14253(.dina(n14540),.dinb(w_n13982_0[0]),.dout(n14541),.clk(gclk));
	jand g14254(.dina(n14541),.dinb(w_asqrt12_21[2]),.dout(n14542),.clk(gclk));
	jxor g14255(.dina(n14542),.dinb(w_n13992_0[0]),.dout(n14543),.clk(gclk));
	jnot g14256(.din(n14543),.dout(n14544),.clk(gclk));
	jor g14257(.dina(w_n14531_0[1]),.dinb(w_asqrt40_13[2]),.dout(n14545),.clk(gclk));
	jor g14258(.dina(n14545),.dinb(w_n14537_0[1]),.dout(n14546),.clk(gclk));
	jand g14259(.dina(w_n14546_0[1]),.dinb(w_n14544_0[1]),.dout(n14547),.clk(gclk));
	jor g14260(.dina(w_n14547_0[1]),.dinb(w_n14539_0[1]),.dout(n14548),.clk(gclk));
	jand g14261(.dina(w_n14548_0[2]),.dinb(w_asqrt41_11[2]),.dout(n14549),.clk(gclk));
	jor g14262(.dina(w_n14548_0[1]),.dinb(w_asqrt41_11[1]),.dout(n14550),.clk(gclk));
	jnot g14263(.din(w_n13998_0[0]),.dout(n14551),.clk(gclk));
	jnot g14264(.din(w_n13999_0[0]),.dout(n14552),.clk(gclk));
	jand g14265(.dina(w_asqrt12_21[1]),.dinb(w_n13995_0[0]),.dout(n14553),.clk(gclk));
	jand g14266(.dina(w_n14553_0[1]),.dinb(n14552),.dout(n14554),.clk(gclk));
	jor g14267(.dina(n14554),.dinb(n14551),.dout(n14555),.clk(gclk));
	jnot g14268(.din(w_n14000_0[0]),.dout(n14556),.clk(gclk));
	jand g14269(.dina(w_n14553_0[0]),.dinb(n14556),.dout(n14557),.clk(gclk));
	jnot g14270(.din(n14557),.dout(n14558),.clk(gclk));
	jand g14271(.dina(n14558),.dinb(n14555),.dout(n14559),.clk(gclk));
	jand g14272(.dina(w_n14559_0[1]),.dinb(n14550),.dout(n14560),.clk(gclk));
	jor g14273(.dina(w_n14560_0[1]),.dinb(w_n14549_0[1]),.dout(n14561),.clk(gclk));
	jand g14274(.dina(n14561),.dinb(w_asqrt42_14[0]),.dout(n14562),.clk(gclk));
	jor g14275(.dina(w_n14549_0[0]),.dinb(w_asqrt42_13[2]),.dout(n14563),.clk(gclk));
	jor g14276(.dina(n14563),.dinb(w_n14560_0[0]),.dout(n14564),.clk(gclk));
	jnot g14277(.din(w_n14006_0[0]),.dout(n14565),.clk(gclk));
	jnot g14278(.din(w_n14008_0[0]),.dout(n14566),.clk(gclk));
	jand g14279(.dina(w_asqrt12_21[0]),.dinb(w_n14002_0[0]),.dout(n14567),.clk(gclk));
	jand g14280(.dina(w_n14567_0[1]),.dinb(n14566),.dout(n14568),.clk(gclk));
	jor g14281(.dina(n14568),.dinb(n14565),.dout(n14569),.clk(gclk));
	jnot g14282(.din(w_n14009_0[0]),.dout(n14570),.clk(gclk));
	jand g14283(.dina(w_n14567_0[0]),.dinb(n14570),.dout(n14571),.clk(gclk));
	jnot g14284(.din(n14571),.dout(n14572),.clk(gclk));
	jand g14285(.dina(n14572),.dinb(n14569),.dout(n14573),.clk(gclk));
	jand g14286(.dina(w_n14573_0[1]),.dinb(w_n14564_0[1]),.dout(n14574),.clk(gclk));
	jor g14287(.dina(n14574),.dinb(w_n14562_0[1]),.dout(n14575),.clk(gclk));
	jand g14288(.dina(w_n14575_0[1]),.dinb(w_asqrt43_11[2]),.dout(n14576),.clk(gclk));
	jxor g14289(.dina(w_n14010_0[0]),.dinb(w_n2870_13[1]),.dout(n14577),.clk(gclk));
	jand g14290(.dina(n14577),.dinb(w_asqrt12_20[2]),.dout(n14578),.clk(gclk));
	jxor g14291(.dina(n14578),.dinb(w_n14020_0[0]),.dout(n14579),.clk(gclk));
	jnot g14292(.din(n14579),.dout(n14580),.clk(gclk));
	jor g14293(.dina(w_n14575_0[0]),.dinb(w_asqrt43_11[1]),.dout(n14581),.clk(gclk));
	jand g14294(.dina(w_n14581_0[1]),.dinb(w_n14580_0[1]),.dout(n14582),.clk(gclk));
	jor g14295(.dina(w_n14582_0[2]),.dinb(w_n14576_0[2]),.dout(n14583),.clk(gclk));
	jand g14296(.dina(n14583),.dinb(w_asqrt44_14[0]),.dout(n14584),.clk(gclk));
	jnot g14297(.din(w_n14025_0[0]),.dout(n14585),.clk(gclk));
	jand g14298(.dina(n14585),.dinb(w_n14023_0[0]),.dout(n14586),.clk(gclk));
	jand g14299(.dina(n14586),.dinb(w_asqrt12_20[1]),.dout(n14587),.clk(gclk));
	jxor g14300(.dina(n14587),.dinb(w_n14033_0[0]),.dout(n14588),.clk(gclk));
	jnot g14301(.din(n14588),.dout(n14589),.clk(gclk));
	jor g14302(.dina(w_n14576_0[1]),.dinb(w_asqrt44_13[2]),.dout(n14590),.clk(gclk));
	jor g14303(.dina(n14590),.dinb(w_n14582_0[1]),.dout(n14591),.clk(gclk));
	jand g14304(.dina(w_n14591_0[1]),.dinb(w_n14589_0[1]),.dout(n14592),.clk(gclk));
	jor g14305(.dina(w_n14592_0[1]),.dinb(w_n14584_0[1]),.dout(n14593),.clk(gclk));
	jand g14306(.dina(w_n14593_0[2]),.dinb(w_asqrt45_12[0]),.dout(n14594),.clk(gclk));
	jor g14307(.dina(w_n14593_0[1]),.dinb(w_asqrt45_11[2]),.dout(n14595),.clk(gclk));
	jnot g14308(.din(w_n14039_0[0]),.dout(n14596),.clk(gclk));
	jnot g14309(.din(w_n14040_0[0]),.dout(n14597),.clk(gclk));
	jand g14310(.dina(w_asqrt12_20[0]),.dinb(w_n14036_0[0]),.dout(n14598),.clk(gclk));
	jand g14311(.dina(w_n14598_0[1]),.dinb(n14597),.dout(n14599),.clk(gclk));
	jor g14312(.dina(n14599),.dinb(n14596),.dout(n14600),.clk(gclk));
	jnot g14313(.din(w_n14041_0[0]),.dout(n14601),.clk(gclk));
	jand g14314(.dina(w_n14598_0[0]),.dinb(n14601),.dout(n14602),.clk(gclk));
	jnot g14315(.din(n14602),.dout(n14603),.clk(gclk));
	jand g14316(.dina(n14603),.dinb(n14600),.dout(n14604),.clk(gclk));
	jand g14317(.dina(w_n14604_0[1]),.dinb(n14595),.dout(n14605),.clk(gclk));
	jor g14318(.dina(w_n14605_0[1]),.dinb(w_n14594_0[1]),.dout(n14606),.clk(gclk));
	jand g14319(.dina(n14606),.dinb(w_asqrt46_14[0]),.dout(n14607),.clk(gclk));
	jor g14320(.dina(w_n14594_0[0]),.dinb(w_asqrt46_13[2]),.dout(n14608),.clk(gclk));
	jor g14321(.dina(n14608),.dinb(w_n14605_0[0]),.dout(n14609),.clk(gclk));
	jnot g14322(.din(w_n14047_0[0]),.dout(n14610),.clk(gclk));
	jnot g14323(.din(w_n14049_0[0]),.dout(n14611),.clk(gclk));
	jand g14324(.dina(w_asqrt12_19[2]),.dinb(w_n14043_0[0]),.dout(n14612),.clk(gclk));
	jand g14325(.dina(w_n14612_0[1]),.dinb(n14611),.dout(n14613),.clk(gclk));
	jor g14326(.dina(n14613),.dinb(n14610),.dout(n14614),.clk(gclk));
	jnot g14327(.din(w_n14050_0[0]),.dout(n14615),.clk(gclk));
	jand g14328(.dina(w_n14612_0[0]),.dinb(n14615),.dout(n14616),.clk(gclk));
	jnot g14329(.din(n14616),.dout(n14617),.clk(gclk));
	jand g14330(.dina(n14617),.dinb(n14614),.dout(n14618),.clk(gclk));
	jand g14331(.dina(w_n14618_0[1]),.dinb(w_n14609_0[1]),.dout(n14619),.clk(gclk));
	jor g14332(.dina(n14619),.dinb(w_n14607_0[1]),.dout(n14620),.clk(gclk));
	jand g14333(.dina(w_n14620_0[1]),.dinb(w_asqrt47_12[0]),.dout(n14621),.clk(gclk));
	jxor g14334(.dina(w_n14051_0[0]),.dinb(w_n2005_14[1]),.dout(n14622),.clk(gclk));
	jand g14335(.dina(n14622),.dinb(w_asqrt12_19[1]),.dout(n14623),.clk(gclk));
	jxor g14336(.dina(n14623),.dinb(w_n14061_0[0]),.dout(n14624),.clk(gclk));
	jnot g14337(.din(n14624),.dout(n14625),.clk(gclk));
	jor g14338(.dina(w_n14620_0[0]),.dinb(w_asqrt47_11[2]),.dout(n14626),.clk(gclk));
	jand g14339(.dina(w_n14626_0[1]),.dinb(w_n14625_0[1]),.dout(n14627),.clk(gclk));
	jor g14340(.dina(w_n14627_0[2]),.dinb(w_n14621_0[2]),.dout(n14628),.clk(gclk));
	jand g14341(.dina(n14628),.dinb(w_asqrt48_14[0]),.dout(n14629),.clk(gclk));
	jnot g14342(.din(w_n14066_0[0]),.dout(n14630),.clk(gclk));
	jand g14343(.dina(n14630),.dinb(w_n14064_0[0]),.dout(n14631),.clk(gclk));
	jand g14344(.dina(n14631),.dinb(w_asqrt12_19[0]),.dout(n14632),.clk(gclk));
	jxor g14345(.dina(n14632),.dinb(w_n14074_0[0]),.dout(n14633),.clk(gclk));
	jnot g14346(.din(n14633),.dout(n14634),.clk(gclk));
	jor g14347(.dina(w_n14621_0[1]),.dinb(w_asqrt48_13[2]),.dout(n14635),.clk(gclk));
	jor g14348(.dina(n14635),.dinb(w_n14627_0[1]),.dout(n14636),.clk(gclk));
	jand g14349(.dina(w_n14636_0[1]),.dinb(w_n14634_0[1]),.dout(n14637),.clk(gclk));
	jor g14350(.dina(w_n14637_0[1]),.dinb(w_n14629_0[1]),.dout(n14638),.clk(gclk));
	jand g14351(.dina(w_n14638_0[2]),.dinb(w_asqrt49_12[1]),.dout(n14639),.clk(gclk));
	jor g14352(.dina(w_n14638_0[1]),.dinb(w_asqrt49_12[0]),.dout(n14640),.clk(gclk));
	jnot g14353(.din(w_n14080_0[0]),.dout(n14641),.clk(gclk));
	jnot g14354(.din(w_n14081_0[0]),.dout(n14642),.clk(gclk));
	jand g14355(.dina(w_asqrt12_18[2]),.dinb(w_n14077_0[0]),.dout(n14643),.clk(gclk));
	jand g14356(.dina(w_n14643_0[1]),.dinb(n14642),.dout(n14644),.clk(gclk));
	jor g14357(.dina(n14644),.dinb(n14641),.dout(n14645),.clk(gclk));
	jnot g14358(.din(w_n14082_0[0]),.dout(n14646),.clk(gclk));
	jand g14359(.dina(w_n14643_0[0]),.dinb(n14646),.dout(n14647),.clk(gclk));
	jnot g14360(.din(n14647),.dout(n14648),.clk(gclk));
	jand g14361(.dina(n14648),.dinb(n14645),.dout(n14649),.clk(gclk));
	jand g14362(.dina(w_n14649_0[1]),.dinb(n14640),.dout(n14650),.clk(gclk));
	jor g14363(.dina(w_n14650_0[1]),.dinb(w_n14639_0[1]),.dout(n14651),.clk(gclk));
	jand g14364(.dina(n14651),.dinb(w_asqrt50_14[0]),.dout(n14652),.clk(gclk));
	jnot g14365(.din(w_n14086_0[0]),.dout(n14653),.clk(gclk));
	jand g14366(.dina(n14653),.dinb(w_n14084_0[0]),.dout(n14654),.clk(gclk));
	jand g14367(.dina(n14654),.dinb(w_asqrt12_18[1]),.dout(n14655),.clk(gclk));
	jxor g14368(.dina(n14655),.dinb(w_n14094_0[0]),.dout(n14656),.clk(gclk));
	jnot g14369(.din(n14656),.dout(n14657),.clk(gclk));
	jor g14370(.dina(w_n14639_0[0]),.dinb(w_asqrt50_13[2]),.dout(n14658),.clk(gclk));
	jor g14371(.dina(n14658),.dinb(w_n14650_0[0]),.dout(n14659),.clk(gclk));
	jand g14372(.dina(w_n14659_0[1]),.dinb(w_n14657_0[1]),.dout(n14660),.clk(gclk));
	jor g14373(.dina(w_n14660_0[1]),.dinb(w_n14652_0[1]),.dout(n14661),.clk(gclk));
	jand g14374(.dina(w_n14661_0[2]),.dinb(w_asqrt51_12[1]),.dout(n14662),.clk(gclk));
	jnot g14375(.din(w_n14246_0[1]),.dout(n14663),.clk(gclk));
	jor g14376(.dina(w_n14661_0[1]),.dinb(w_asqrt51_12[0]),.dout(n14664),.clk(gclk));
	jand g14377(.dina(n14664),.dinb(n14663),.dout(n14665),.clk(gclk));
	jor g14378(.dina(w_n14665_0[1]),.dinb(w_n14662_0[1]),.dout(n14666),.clk(gclk));
	jand g14379(.dina(n14666),.dinb(w_asqrt52_14[0]),.dout(n14667),.clk(gclk));
	jor g14380(.dina(w_n14662_0[0]),.dinb(w_asqrt52_13[2]),.dout(n14668),.clk(gclk));
	jor g14381(.dina(n14668),.dinb(w_n14665_0[0]),.dout(n14669),.clk(gclk));
	jnot g14382(.din(w_n14105_0[0]),.dout(n14670),.clk(gclk));
	jnot g14383(.din(w_n14107_0[0]),.dout(n14671),.clk(gclk));
	jand g14384(.dina(w_asqrt12_18[0]),.dinb(w_n14101_0[0]),.dout(n14672),.clk(gclk));
	jand g14385(.dina(w_n14672_0[1]),.dinb(n14671),.dout(n14673),.clk(gclk));
	jor g14386(.dina(n14673),.dinb(n14670),.dout(n14674),.clk(gclk));
	jnot g14387(.din(w_n14108_0[0]),.dout(n14675),.clk(gclk));
	jand g14388(.dina(w_n14672_0[0]),.dinb(n14675),.dout(n14676),.clk(gclk));
	jnot g14389(.din(n14676),.dout(n14677),.clk(gclk));
	jand g14390(.dina(n14677),.dinb(n14674),.dout(n14678),.clk(gclk));
	jand g14391(.dina(w_n14678_0[1]),.dinb(w_n14669_0[1]),.dout(n14679),.clk(gclk));
	jor g14392(.dina(n14679),.dinb(w_n14667_0[1]),.dout(n14680),.clk(gclk));
	jand g14393(.dina(w_n14680_0[2]),.dinb(w_asqrt53_12[2]),.dout(n14681),.clk(gclk));
	jor g14394(.dina(w_n14680_0[1]),.dinb(w_asqrt53_12[1]),.dout(n14682),.clk(gclk));
	jnot g14395(.din(w_n14113_0[0]),.dout(n14683),.clk(gclk));
	jnot g14396(.din(w_n14114_0[0]),.dout(n14684),.clk(gclk));
	jand g14397(.dina(w_asqrt12_17[2]),.dinb(w_n14110_0[0]),.dout(n14685),.clk(gclk));
	jand g14398(.dina(w_n14685_0[1]),.dinb(n14684),.dout(n14686),.clk(gclk));
	jor g14399(.dina(n14686),.dinb(n14683),.dout(n14687),.clk(gclk));
	jnot g14400(.din(w_n14115_0[0]),.dout(n14688),.clk(gclk));
	jand g14401(.dina(w_n14685_0[0]),.dinb(n14688),.dout(n14689),.clk(gclk));
	jnot g14402(.din(n14689),.dout(n14690),.clk(gclk));
	jand g14403(.dina(n14690),.dinb(n14687),.dout(n14691),.clk(gclk));
	jand g14404(.dina(w_n14691_0[1]),.dinb(n14682),.dout(n14692),.clk(gclk));
	jor g14405(.dina(w_n14692_0[1]),.dinb(w_n14681_0[1]),.dout(n14693),.clk(gclk));
	jand g14406(.dina(n14693),.dinb(w_asqrt54_14[0]),.dout(n14694),.clk(gclk));
	jor g14407(.dina(w_n14681_0[0]),.dinb(w_asqrt54_13[2]),.dout(n14695),.clk(gclk));
	jor g14408(.dina(n14695),.dinb(w_n14692_0[0]),.dout(n14696),.clk(gclk));
	jnot g14409(.din(w_n14121_0[0]),.dout(n14697),.clk(gclk));
	jnot g14410(.din(w_n14123_0[0]),.dout(n14698),.clk(gclk));
	jand g14411(.dina(w_asqrt12_17[1]),.dinb(w_n14117_0[0]),.dout(n14699),.clk(gclk));
	jand g14412(.dina(w_n14699_0[1]),.dinb(n14698),.dout(n14700),.clk(gclk));
	jor g14413(.dina(n14700),.dinb(n14697),.dout(n14701),.clk(gclk));
	jnot g14414(.din(w_n14124_0[0]),.dout(n14702),.clk(gclk));
	jand g14415(.dina(w_n14699_0[0]),.dinb(n14702),.dout(n14703),.clk(gclk));
	jnot g14416(.din(n14703),.dout(n14704),.clk(gclk));
	jand g14417(.dina(n14704),.dinb(n14701),.dout(n14705),.clk(gclk));
	jand g14418(.dina(w_n14705_0[1]),.dinb(w_n14696_0[1]),.dout(n14706),.clk(gclk));
	jor g14419(.dina(n14706),.dinb(w_n14694_0[1]),.dout(n14707),.clk(gclk));
	jand g14420(.dina(w_n14707_0[1]),.dinb(w_asqrt55_13[0]),.dout(n14708),.clk(gclk));
	jxor g14421(.dina(w_n14125_0[0]),.dinb(w_n791_16[0]),.dout(n14709),.clk(gclk));
	jand g14422(.dina(n14709),.dinb(w_asqrt12_17[0]),.dout(n14710),.clk(gclk));
	jxor g14423(.dina(n14710),.dinb(w_n14135_0[0]),.dout(n14711),.clk(gclk));
	jnot g14424(.din(n14711),.dout(n14712),.clk(gclk));
	jor g14425(.dina(w_n14707_0[0]),.dinb(w_asqrt55_12[2]),.dout(n14713),.clk(gclk));
	jand g14426(.dina(w_n14713_0[1]),.dinb(w_n14712_0[1]),.dout(n14714),.clk(gclk));
	jor g14427(.dina(w_n14714_0[2]),.dinb(w_n14708_0[2]),.dout(n14715),.clk(gclk));
	jand g14428(.dina(n14715),.dinb(w_asqrt56_14[0]),.dout(n14716),.clk(gclk));
	jnot g14429(.din(w_n14140_0[0]),.dout(n14717),.clk(gclk));
	jand g14430(.dina(n14717),.dinb(w_n14138_0[0]),.dout(n14718),.clk(gclk));
	jand g14431(.dina(n14718),.dinb(w_asqrt12_16[2]),.dout(n14719),.clk(gclk));
	jxor g14432(.dina(n14719),.dinb(w_n14148_0[0]),.dout(n14720),.clk(gclk));
	jnot g14433(.din(n14720),.dout(n14721),.clk(gclk));
	jor g14434(.dina(w_n14708_0[1]),.dinb(w_asqrt56_13[2]),.dout(n14722),.clk(gclk));
	jor g14435(.dina(n14722),.dinb(w_n14714_0[1]),.dout(n14723),.clk(gclk));
	jand g14436(.dina(w_n14723_0[1]),.dinb(w_n14721_0[1]),.dout(n14724),.clk(gclk));
	jor g14437(.dina(w_n14724_0[1]),.dinb(w_n14716_0[1]),.dout(n14725),.clk(gclk));
	jand g14438(.dina(w_n14725_0[2]),.dinb(w_asqrt57_13[1]),.dout(n14726),.clk(gclk));
	jor g14439(.dina(w_n14725_0[1]),.dinb(w_asqrt57_13[0]),.dout(n14727),.clk(gclk));
	jnot g14440(.din(w_n14154_0[0]),.dout(n14728),.clk(gclk));
	jnot g14441(.din(w_n14155_0[0]),.dout(n14729),.clk(gclk));
	jand g14442(.dina(w_asqrt12_16[1]),.dinb(w_n14151_0[0]),.dout(n14730),.clk(gclk));
	jand g14443(.dina(w_n14730_0[1]),.dinb(n14729),.dout(n14731),.clk(gclk));
	jor g14444(.dina(n14731),.dinb(n14728),.dout(n14732),.clk(gclk));
	jnot g14445(.din(w_n14156_0[0]),.dout(n14733),.clk(gclk));
	jand g14446(.dina(w_n14730_0[0]),.dinb(n14733),.dout(n14734),.clk(gclk));
	jnot g14447(.din(n14734),.dout(n14735),.clk(gclk));
	jand g14448(.dina(n14735),.dinb(n14732),.dout(n14736),.clk(gclk));
	jand g14449(.dina(w_n14736_0[1]),.dinb(n14727),.dout(n14737),.clk(gclk));
	jor g14450(.dina(w_n14737_0[1]),.dinb(w_n14726_0[1]),.dout(n14738),.clk(gclk));
	jand g14451(.dina(n14738),.dinb(w_asqrt58_14[0]),.dout(n14739),.clk(gclk));
	jor g14452(.dina(w_n14726_0[0]),.dinb(w_asqrt58_13[2]),.dout(n14740),.clk(gclk));
	jor g14453(.dina(n14740),.dinb(w_n14737_0[0]),.dout(n14741),.clk(gclk));
	jnot g14454(.din(w_n14162_0[0]),.dout(n14742),.clk(gclk));
	jnot g14455(.din(w_n14164_0[0]),.dout(n14743),.clk(gclk));
	jand g14456(.dina(w_asqrt12_16[0]),.dinb(w_n14158_0[0]),.dout(n14744),.clk(gclk));
	jand g14457(.dina(w_n14744_0[1]),.dinb(n14743),.dout(n14745),.clk(gclk));
	jor g14458(.dina(n14745),.dinb(n14742),.dout(n14746),.clk(gclk));
	jnot g14459(.din(w_n14165_0[0]),.dout(n14747),.clk(gclk));
	jand g14460(.dina(w_n14744_0[0]),.dinb(n14747),.dout(n14748),.clk(gclk));
	jnot g14461(.din(n14748),.dout(n14749),.clk(gclk));
	jand g14462(.dina(n14749),.dinb(n14746),.dout(n14750),.clk(gclk));
	jand g14463(.dina(w_n14750_0[1]),.dinb(w_n14741_0[1]),.dout(n14751),.clk(gclk));
	jor g14464(.dina(n14751),.dinb(w_n14739_0[1]),.dout(n14752),.clk(gclk));
	jand g14465(.dina(w_n14752_0[1]),.dinb(w_asqrt59_13[2]),.dout(n14753),.clk(gclk));
	jxor g14466(.dina(w_n14166_0[0]),.dinb(w_n425_16[2]),.dout(n14754),.clk(gclk));
	jand g14467(.dina(n14754),.dinb(w_asqrt12_15[2]),.dout(n14755),.clk(gclk));
	jxor g14468(.dina(n14755),.dinb(w_n14176_0[0]),.dout(n14756),.clk(gclk));
	jnot g14469(.din(n14756),.dout(n14757),.clk(gclk));
	jor g14470(.dina(w_n14752_0[0]),.dinb(w_asqrt59_13[1]),.dout(n14758),.clk(gclk));
	jand g14471(.dina(w_n14758_0[1]),.dinb(w_n14757_0[1]),.dout(n14759),.clk(gclk));
	jor g14472(.dina(w_n14759_0[2]),.dinb(w_n14753_0[2]),.dout(n14760),.clk(gclk));
	jand g14473(.dina(n14760),.dinb(w_asqrt60_13[2]),.dout(n14761),.clk(gclk));
	jnot g14474(.din(w_n14181_0[0]),.dout(n14762),.clk(gclk));
	jand g14475(.dina(n14762),.dinb(w_n14179_0[0]),.dout(n14763),.clk(gclk));
	jand g14476(.dina(n14763),.dinb(w_asqrt12_15[1]),.dout(n14764),.clk(gclk));
	jxor g14477(.dina(n14764),.dinb(w_n14189_0[0]),.dout(n14765),.clk(gclk));
	jnot g14478(.din(n14765),.dout(n14766),.clk(gclk));
	jor g14479(.dina(w_n14753_0[1]),.dinb(w_asqrt60_13[1]),.dout(n14767),.clk(gclk));
	jor g14480(.dina(n14767),.dinb(w_n14759_0[1]),.dout(n14768),.clk(gclk));
	jand g14481(.dina(w_n14768_0[1]),.dinb(w_n14766_0[1]),.dout(n14769),.clk(gclk));
	jor g14482(.dina(w_n14769_0[1]),.dinb(w_n14761_0[1]),.dout(n14770),.clk(gclk));
	jand g14483(.dina(w_n14770_0[2]),.dinb(w_asqrt61_14[0]),.dout(n14771),.clk(gclk));
	jor g14484(.dina(w_n14770_0[1]),.dinb(w_asqrt61_13[2]),.dout(n14772),.clk(gclk));
	jnot g14485(.din(w_n14195_0[0]),.dout(n14773),.clk(gclk));
	jnot g14486(.din(w_n14196_0[0]),.dout(n14774),.clk(gclk));
	jand g14487(.dina(w_asqrt12_15[0]),.dinb(w_n14192_0[0]),.dout(n14775),.clk(gclk));
	jand g14488(.dina(w_n14775_0[1]),.dinb(n14774),.dout(n14776),.clk(gclk));
	jor g14489(.dina(n14776),.dinb(n14773),.dout(n14777),.clk(gclk));
	jnot g14490(.din(w_n14197_0[0]),.dout(n14778),.clk(gclk));
	jand g14491(.dina(w_n14775_0[0]),.dinb(n14778),.dout(n14779),.clk(gclk));
	jnot g14492(.din(n14779),.dout(n14780),.clk(gclk));
	jand g14493(.dina(n14780),.dinb(n14777),.dout(n14781),.clk(gclk));
	jand g14494(.dina(w_n14781_0[1]),.dinb(n14772),.dout(n14782),.clk(gclk));
	jor g14495(.dina(w_n14782_0[1]),.dinb(w_n14771_0[1]),.dout(n14783),.clk(gclk));
	jand g14496(.dina(n14783),.dinb(w_asqrt62_14[0]),.dout(n14784),.clk(gclk));
	jor g14497(.dina(w_n14771_0[0]),.dinb(w_asqrt62_13[2]),.dout(n14785),.clk(gclk));
	jor g14498(.dina(n14785),.dinb(w_n14782_0[0]),.dout(n14786),.clk(gclk));
	jnot g14499(.din(w_n14203_0[0]),.dout(n14787),.clk(gclk));
	jnot g14500(.din(w_n14205_0[0]),.dout(n14788),.clk(gclk));
	jand g14501(.dina(w_asqrt12_14[2]),.dinb(w_n14199_0[0]),.dout(n14789),.clk(gclk));
	jand g14502(.dina(w_n14789_0[1]),.dinb(n14788),.dout(n14790),.clk(gclk));
	jor g14503(.dina(n14790),.dinb(n14787),.dout(n14791),.clk(gclk));
	jnot g14504(.din(w_n14206_0[0]),.dout(n14792),.clk(gclk));
	jand g14505(.dina(w_n14789_0[0]),.dinb(n14792),.dout(n14793),.clk(gclk));
	jnot g14506(.din(n14793),.dout(n14794),.clk(gclk));
	jand g14507(.dina(n14794),.dinb(n14791),.dout(n14795),.clk(gclk));
	jand g14508(.dina(w_n14795_0[1]),.dinb(w_n14786_0[1]),.dout(n14796),.clk(gclk));
	jor g14509(.dina(n14796),.dinb(w_n14784_0[1]),.dout(n14797),.clk(gclk));
	jxor g14510(.dina(w_n14207_0[0]),.dinb(w_n199_20[2]),.dout(n14798),.clk(gclk));
	jand g14511(.dina(n14798),.dinb(w_asqrt12_14[1]),.dout(n14799),.clk(gclk));
	jxor g14512(.dina(n14799),.dinb(w_n14217_0[0]),.dout(n14800),.clk(gclk));
	jnot g14513(.din(w_n14219_0[0]),.dout(n14801),.clk(gclk));
	jand g14514(.dina(w_asqrt12_14[0]),.dinb(w_n14226_0[1]),.dout(n14802),.clk(gclk));
	jand g14515(.dina(w_n14802_0[1]),.dinb(w_n14801_0[2]),.dout(n14803),.clk(gclk));
	jor g14516(.dina(n14803),.dinb(w_n14234_0[0]),.dout(n14804),.clk(gclk));
	jor g14517(.dina(n14804),.dinb(w_n14800_0[1]),.dout(n14805),.clk(gclk));
	jnot g14518(.din(n14805),.dout(n14806),.clk(gclk));
	jand g14519(.dina(n14806),.dinb(w_n14797_1[2]),.dout(n14807),.clk(gclk));
	jor g14520(.dina(n14807),.dinb(w_asqrt63_7[2]),.dout(n14808),.clk(gclk));
	jnot g14521(.din(w_n14800_0[0]),.dout(n14809),.clk(gclk));
	jor g14522(.dina(w_n14809_0[2]),.dinb(w_n14797_1[1]),.dout(n14810),.clk(gclk));
	jor g14523(.dina(w_n14802_0[0]),.dinb(w_n14801_0[1]),.dout(n14811),.clk(gclk));
	jand g14524(.dina(w_n14226_0[0]),.dinb(w_n14801_0[0]),.dout(n14812),.clk(gclk));
	jor g14525(.dina(n14812),.dinb(w_n194_19[2]),.dout(n14813),.clk(gclk));
	jnot g14526(.din(n14813),.dout(n14814),.clk(gclk));
	jand g14527(.dina(n14814),.dinb(n14811),.dout(n14815),.clk(gclk));
	jnot g14528(.din(w_asqrt12_13[2]),.dout(n14816),.clk(gclk));
	jnot g14529(.din(w_n14815_0[1]),.dout(n14819),.clk(gclk));
	jand g14530(.dina(n14819),.dinb(w_n14810_0[1]),.dout(n14820),.clk(gclk));
	jand g14531(.dina(n14820),.dinb(w_n14808_0[1]),.dout(n14821),.clk(gclk));
	jxor g14532(.dina(w_n14661_0[0]),.dinb(w_n1039_17[1]),.dout(n14822),.clk(gclk));
	jor g14533(.dina(n14822),.dinb(w_n14821_22[2]),.dout(n14823),.clk(gclk));
	jxor g14534(.dina(n14823),.dinb(w_n14246_0[0]),.dout(n14824),.clk(gclk));
	jor g14535(.dina(w_n14821_22[1]),.dinb(w_n14248_1[0]),.dout(n14825),.clk(gclk));
	jnot g14536(.din(w_a20_0[1]),.dout(n14826),.clk(gclk));
	jnot g14537(.din(a[21]),.dout(n14827),.clk(gclk));
	jand g14538(.dina(w_n14248_0[2]),.dinb(w_n14827_0[2]),.dout(n14828),.clk(gclk));
	jand g14539(.dina(n14828),.dinb(w_n14826_1[1]),.dout(n14829),.clk(gclk));
	jnot g14540(.din(n14829),.dout(n14830),.clk(gclk));
	jand g14541(.dina(n14830),.dinb(n14825),.dout(n14831),.clk(gclk));
	jor g14542(.dina(w_n14831_0[2]),.dinb(w_n14816_8[1]),.dout(n14832),.clk(gclk));
	jor g14543(.dina(w_n14821_22[0]),.dinb(w_a22_0[0]),.dout(n14833),.clk(gclk));
	jxor g14544(.dina(w_n14833_0[1]),.dinb(w_n14249_0[0]),.dout(n14834),.clk(gclk));
	jand g14545(.dina(w_n14831_0[1]),.dinb(w_n14816_8[0]),.dout(n14835),.clk(gclk));
	jor g14546(.dina(n14835),.dinb(w_n14834_0[1]),.dout(n14836),.clk(gclk));
	jand g14547(.dina(w_n14836_0[1]),.dinb(w_n14832_0[1]),.dout(n14837),.clk(gclk));
	jor g14548(.dina(n14837),.dinb(w_n13723_12[2]),.dout(n14838),.clk(gclk));
	jand g14549(.dina(w_n14832_0[0]),.dinb(w_n13723_12[1]),.dout(n14839),.clk(gclk));
	jand g14550(.dina(n14839),.dinb(w_n14836_0[0]),.dout(n14840),.clk(gclk));
	jor g14551(.dina(w_n14833_0[0]),.dinb(w_a23_0[0]),.dout(n14841),.clk(gclk));
	jnot g14552(.din(w_n14808_0[0]),.dout(n14842),.clk(gclk));
	jnot g14553(.din(w_n14810_0[0]),.dout(n14843),.clk(gclk));
	jor g14554(.dina(w_n14815_0[0]),.dinb(w_n14816_7[2]),.dout(n14844),.clk(gclk));
	jor g14555(.dina(n14844),.dinb(w_n14843_0[1]),.dout(n14845),.clk(gclk));
	jor g14556(.dina(n14845),.dinb(n14842),.dout(n14846),.clk(gclk));
	jand g14557(.dina(n14846),.dinb(n14841),.dout(n14847),.clk(gclk));
	jxor g14558(.dina(n14847),.dinb(w_n13728_0[1]),.dout(n14848),.clk(gclk));
	jor g14559(.dina(w_n14848_0[1]),.dinb(w_n14840_0[1]),.dout(n14849),.clk(gclk));
	jand g14560(.dina(n14849),.dinb(w_n14838_0[1]),.dout(n14850),.clk(gclk));
	jor g14561(.dina(w_n14850_0[2]),.dinb(w_n13718_8[0]),.dout(n14851),.clk(gclk));
	jand g14562(.dina(w_n14850_0[1]),.dinb(w_n13718_7[2]),.dout(n14852),.clk(gclk));
	jxor g14563(.dina(w_n14252_0[0]),.dinb(w_n13723_12[0]),.dout(n14853),.clk(gclk));
	jor g14564(.dina(n14853),.dinb(w_n14821_21[2]),.dout(n14854),.clk(gclk));
	jxor g14565(.dina(n14854),.dinb(w_n14255_0[0]),.dout(n14855),.clk(gclk));
	jor g14566(.dina(w_n14855_0[1]),.dinb(n14852),.dout(n14856),.clk(gclk));
	jand g14567(.dina(w_n14856_0[1]),.dinb(w_n14851_0[1]),.dout(n14857),.clk(gclk));
	jor g14568(.dina(n14857),.dinb(w_n12675_13[1]),.dout(n14858),.clk(gclk));
	jnot g14569(.din(w_n14261_0[0]),.dout(n14859),.clk(gclk));
	jor g14570(.dina(n14859),.dinb(w_n14259_0[0]),.dout(n14860),.clk(gclk));
	jor g14571(.dina(n14860),.dinb(w_n14821_21[1]),.dout(n14861),.clk(gclk));
	jxor g14572(.dina(n14861),.dinb(w_n14270_0[0]),.dout(n14862),.clk(gclk));
	jand g14573(.dina(w_n14851_0[0]),.dinb(w_n12675_13[0]),.dout(n14863),.clk(gclk));
	jand g14574(.dina(n14863),.dinb(w_n14856_0[0]),.dout(n14864),.clk(gclk));
	jor g14575(.dina(w_n14864_0[1]),.dinb(w_n14862_0[1]),.dout(n14865),.clk(gclk));
	jand g14576(.dina(w_n14865_0[1]),.dinb(w_n14858_0[1]),.dout(n14866),.clk(gclk));
	jor g14577(.dina(w_n14866_0[2]),.dinb(w_n12670_8[1]),.dout(n14867),.clk(gclk));
	jand g14578(.dina(w_n14866_0[1]),.dinb(w_n12670_8[0]),.dout(n14868),.clk(gclk));
	jxor g14579(.dina(w_n14272_0[0]),.dinb(w_n12675_12[2]),.dout(n14869),.clk(gclk));
	jor g14580(.dina(n14869),.dinb(w_n14821_21[0]),.dout(n14870),.clk(gclk));
	jxor g14581(.dina(n14870),.dinb(w_n14277_0[0]),.dout(n14871),.clk(gclk));
	jnot g14582(.din(w_n14871_0[1]),.dout(n14872),.clk(gclk));
	jor g14583(.dina(n14872),.dinb(n14868),.dout(n14873),.clk(gclk));
	jand g14584(.dina(w_n14873_0[1]),.dinb(w_n14867_0[1]),.dout(n14874),.clk(gclk));
	jor g14585(.dina(n14874),.dinb(w_n11662_13[0]),.dout(n14875),.clk(gclk));
	jand g14586(.dina(w_n14867_0[0]),.dinb(w_n11662_12[2]),.dout(n14876),.clk(gclk));
	jand g14587(.dina(n14876),.dinb(w_n14873_0[0]),.dout(n14877),.clk(gclk));
	jnot g14588(.din(w_n14281_0[0]),.dout(n14878),.clk(gclk));
	jnot g14589(.din(w_n14821_20[2]),.dout(asqrt_fa_12),.clk(gclk));
	jand g14590(.dina(w_asqrt11_16),.dinb(n14878),.dout(n14880),.clk(gclk));
	jand g14591(.dina(w_n14880_0[1]),.dinb(w_n14288_0[0]),.dout(n14881),.clk(gclk));
	jor g14592(.dina(n14881),.dinb(w_n14286_0[0]),.dout(n14882),.clk(gclk));
	jand g14593(.dina(w_n14880_0[0]),.dinb(w_n14289_0[0]),.dout(n14883),.clk(gclk));
	jnot g14594(.din(n14883),.dout(n14884),.clk(gclk));
	jand g14595(.dina(n14884),.dinb(n14882),.dout(n14885),.clk(gclk));
	jnot g14596(.din(n14885),.dout(n14886),.clk(gclk));
	jor g14597(.dina(w_n14886_0[1]),.dinb(w_n14877_0[1]),.dout(n14887),.clk(gclk));
	jand g14598(.dina(n14887),.dinb(w_n14875_0[1]),.dout(n14888),.clk(gclk));
	jor g14599(.dina(w_n14888_0[2]),.dinb(w_n11657_8[1]),.dout(n14889),.clk(gclk));
	jand g14600(.dina(w_n14888_0[1]),.dinb(w_n11657_8[0]),.dout(n14890),.clk(gclk));
	jnot g14601(.din(w_n14296_0[0]),.dout(n14891),.clk(gclk));
	jxor g14602(.dina(w_n14290_0[0]),.dinb(w_n11662_12[1]),.dout(n14892),.clk(gclk));
	jor g14603(.dina(n14892),.dinb(w_n14821_20[1]),.dout(n14893),.clk(gclk));
	jxor g14604(.dina(n14893),.dinb(n14891),.dout(n14894),.clk(gclk));
	jnot g14605(.din(w_n14894_0[1]),.dout(n14895),.clk(gclk));
	jor g14606(.dina(n14895),.dinb(n14890),.dout(n14896),.clk(gclk));
	jand g14607(.dina(w_n14896_0[1]),.dinb(w_n14889_0[1]),.dout(n14897),.clk(gclk));
	jor g14608(.dina(n14897),.dinb(w_n10701_13[1]),.dout(n14898),.clk(gclk));
	jnot g14609(.din(w_n14301_0[0]),.dout(n14899),.clk(gclk));
	jor g14610(.dina(n14899),.dinb(w_n14299_0[0]),.dout(n14900),.clk(gclk));
	jor g14611(.dina(n14900),.dinb(w_n14821_20[0]),.dout(n14901),.clk(gclk));
	jxor g14612(.dina(n14901),.dinb(w_n14310_0[0]),.dout(n14902),.clk(gclk));
	jand g14613(.dina(w_n14889_0[0]),.dinb(w_n10701_13[0]),.dout(n14903),.clk(gclk));
	jand g14614(.dina(n14903),.dinb(w_n14896_0[0]),.dout(n14904),.clk(gclk));
	jor g14615(.dina(w_n14904_0[1]),.dinb(w_n14902_0[1]),.dout(n14905),.clk(gclk));
	jand g14616(.dina(w_n14905_0[1]),.dinb(w_n14898_0[1]),.dout(n14906),.clk(gclk));
	jor g14617(.dina(w_n14906_0[2]),.dinb(w_n10696_9[0]),.dout(n14907),.clk(gclk));
	jand g14618(.dina(w_n14906_0[1]),.dinb(w_n10696_8[2]),.dout(n14908),.clk(gclk));
	jnot g14619(.din(w_n14317_0[0]),.dout(n14909),.clk(gclk));
	jxor g14620(.dina(w_n14312_0[0]),.dinb(w_n10701_12[2]),.dout(n14910),.clk(gclk));
	jor g14621(.dina(n14910),.dinb(w_n14821_19[2]),.dout(n14911),.clk(gclk));
	jxor g14622(.dina(n14911),.dinb(n14909),.dout(n14912),.clk(gclk));
	jnot g14623(.din(n14912),.dout(n14913),.clk(gclk));
	jor g14624(.dina(w_n14913_0[1]),.dinb(n14908),.dout(n14914),.clk(gclk));
	jand g14625(.dina(w_n14914_0[1]),.dinb(w_n14907_0[1]),.dout(n14915),.clk(gclk));
	jor g14626(.dina(n14915),.dinb(w_n9774_13[0]),.dout(n14916),.clk(gclk));
	jand g14627(.dina(w_n14907_0[0]),.dinb(w_n9774_12[2]),.dout(n14917),.clk(gclk));
	jand g14628(.dina(n14917),.dinb(w_n14914_0[0]),.dout(n14918),.clk(gclk));
	jnot g14629(.din(w_n14320_0[0]),.dout(n14919),.clk(gclk));
	jand g14630(.dina(w_asqrt11_15[2]),.dinb(n14919),.dout(n14920),.clk(gclk));
	jand g14631(.dina(w_n14920_0[1]),.dinb(w_n14327_0[0]),.dout(n14921),.clk(gclk));
	jor g14632(.dina(n14921),.dinb(w_n14325_0[0]),.dout(n14922),.clk(gclk));
	jand g14633(.dina(w_n14920_0[0]),.dinb(w_n14328_0[0]),.dout(n14923),.clk(gclk));
	jnot g14634(.din(n14923),.dout(n14924),.clk(gclk));
	jand g14635(.dina(n14924),.dinb(n14922),.dout(n14925),.clk(gclk));
	jnot g14636(.din(n14925),.dout(n14926),.clk(gclk));
	jor g14637(.dina(w_n14926_0[1]),.dinb(w_n14918_0[1]),.dout(n14927),.clk(gclk));
	jand g14638(.dina(n14927),.dinb(w_n14916_0[1]),.dout(n14928),.clk(gclk));
	jor g14639(.dina(w_n14928_0[1]),.dinb(w_n9769_9[0]),.dout(n14929),.clk(gclk));
	jxor g14640(.dina(w_n14329_0[0]),.dinb(w_n9774_12[1]),.dout(n14930),.clk(gclk));
	jor g14641(.dina(n14930),.dinb(w_n14821_19[1]),.dout(n14931),.clk(gclk));
	jxor g14642(.dina(n14931),.dinb(w_n14334_0[0]),.dout(n14932),.clk(gclk));
	jand g14643(.dina(w_n14928_0[0]),.dinb(w_n9769_8[2]),.dout(n14933),.clk(gclk));
	jor g14644(.dina(w_n14933_0[1]),.dinb(w_n14932_0[1]),.dout(n14934),.clk(gclk));
	jand g14645(.dina(w_n14934_0[2]),.dinb(w_n14929_0[2]),.dout(n14935),.clk(gclk));
	jor g14646(.dina(n14935),.dinb(w_n8898_13[2]),.dout(n14936),.clk(gclk));
	jnot g14647(.din(w_n14339_0[0]),.dout(n14937),.clk(gclk));
	jor g14648(.dina(n14937),.dinb(w_n14337_0[0]),.dout(n14938),.clk(gclk));
	jor g14649(.dina(n14938),.dinb(w_n14821_19[0]),.dout(n14939),.clk(gclk));
	jxor g14650(.dina(n14939),.dinb(w_n14348_0[0]),.dout(n14940),.clk(gclk));
	jand g14651(.dina(w_n14929_0[1]),.dinb(w_n8898_13[1]),.dout(n14941),.clk(gclk));
	jand g14652(.dina(n14941),.dinb(w_n14934_0[1]),.dout(n14942),.clk(gclk));
	jor g14653(.dina(w_n14942_0[1]),.dinb(w_n14940_0[1]),.dout(n14943),.clk(gclk));
	jand g14654(.dina(w_n14943_0[1]),.dinb(w_n14936_0[1]),.dout(n14944),.clk(gclk));
	jor g14655(.dina(w_n14944_0[2]),.dinb(w_n8893_9[2]),.dout(n14945),.clk(gclk));
	jand g14656(.dina(w_n14944_0[1]),.dinb(w_n8893_9[1]),.dout(n14946),.clk(gclk));
	jnot g14657(.din(w_n14351_0[0]),.dout(n14947),.clk(gclk));
	jand g14658(.dina(w_asqrt11_15[1]),.dinb(n14947),.dout(n14948),.clk(gclk));
	jand g14659(.dina(w_n14948_0[1]),.dinb(w_n14356_0[0]),.dout(n14949),.clk(gclk));
	jor g14660(.dina(n14949),.dinb(w_n14355_0[0]),.dout(n14950),.clk(gclk));
	jand g14661(.dina(w_n14948_0[0]),.dinb(w_n14357_0[0]),.dout(n14951),.clk(gclk));
	jnot g14662(.din(n14951),.dout(n14952),.clk(gclk));
	jand g14663(.dina(n14952),.dinb(n14950),.dout(n14953),.clk(gclk));
	jnot g14664(.din(n14953),.dout(n14954),.clk(gclk));
	jor g14665(.dina(w_n14954_0[1]),.dinb(n14946),.dout(n14955),.clk(gclk));
	jand g14666(.dina(w_n14955_0[1]),.dinb(w_n14945_0[1]),.dout(n14956),.clk(gclk));
	jor g14667(.dina(n14956),.dinb(w_n8058_13[2]),.dout(n14957),.clk(gclk));
	jand g14668(.dina(w_n14945_0[0]),.dinb(w_n8058_13[1]),.dout(n14958),.clk(gclk));
	jand g14669(.dina(n14958),.dinb(w_n14955_0[0]),.dout(n14959),.clk(gclk));
	jnot g14670(.din(w_n14359_0[0]),.dout(n14960),.clk(gclk));
	jand g14671(.dina(w_asqrt11_15[0]),.dinb(n14960),.dout(n14961),.clk(gclk));
	jand g14672(.dina(w_n14961_0[1]),.dinb(w_n14366_0[0]),.dout(n14962),.clk(gclk));
	jor g14673(.dina(n14962),.dinb(w_n14364_0[0]),.dout(n14963),.clk(gclk));
	jand g14674(.dina(w_n14961_0[0]),.dinb(w_n14367_0[0]),.dout(n14964),.clk(gclk));
	jnot g14675(.din(n14964),.dout(n14965),.clk(gclk));
	jand g14676(.dina(n14965),.dinb(n14963),.dout(n14966),.clk(gclk));
	jnot g14677(.din(n14966),.dout(n14967),.clk(gclk));
	jor g14678(.dina(w_n14967_0[1]),.dinb(w_n14959_0[1]),.dout(n14968),.clk(gclk));
	jand g14679(.dina(n14968),.dinb(w_n14957_0[1]),.dout(n14969),.clk(gclk));
	jor g14680(.dina(w_n14969_0[1]),.dinb(w_n8053_9[2]),.dout(n14970),.clk(gclk));
	jxor g14681(.dina(w_n14368_0[0]),.dinb(w_n8058_13[0]),.dout(n14971),.clk(gclk));
	jor g14682(.dina(n14971),.dinb(w_n14821_18[2]),.dout(n14972),.clk(gclk));
	jxor g14683(.dina(n14972),.dinb(w_n14379_0[0]),.dout(n14973),.clk(gclk));
	jand g14684(.dina(w_n14969_0[0]),.dinb(w_n8053_9[1]),.dout(n14974),.clk(gclk));
	jor g14685(.dina(w_n14974_0[1]),.dinb(w_n14973_0[1]),.dout(n14975),.clk(gclk));
	jand g14686(.dina(w_n14975_0[2]),.dinb(w_n14970_0[2]),.dout(n14976),.clk(gclk));
	jor g14687(.dina(n14976),.dinb(w_n7265_14[0]),.dout(n14977),.clk(gclk));
	jnot g14688(.din(w_n14384_0[0]),.dout(n14978),.clk(gclk));
	jor g14689(.dina(n14978),.dinb(w_n14382_0[0]),.dout(n14979),.clk(gclk));
	jor g14690(.dina(n14979),.dinb(w_n14821_18[1]),.dout(n14980),.clk(gclk));
	jxor g14691(.dina(n14980),.dinb(w_n14393_0[0]),.dout(n14981),.clk(gclk));
	jand g14692(.dina(w_n14970_0[1]),.dinb(w_n7265_13[2]),.dout(n14982),.clk(gclk));
	jand g14693(.dina(n14982),.dinb(w_n14975_0[1]),.dout(n14983),.clk(gclk));
	jor g14694(.dina(w_n14983_0[1]),.dinb(w_n14981_0[1]),.dout(n14984),.clk(gclk));
	jand g14695(.dina(w_n14984_0[1]),.dinb(w_n14977_0[1]),.dout(n14985),.clk(gclk));
	jor g14696(.dina(w_n14985_0[2]),.dinb(w_n7260_10[2]),.dout(n14986),.clk(gclk));
	jand g14697(.dina(w_n14985_0[1]),.dinb(w_n7260_10[1]),.dout(n14987),.clk(gclk));
	jnot g14698(.din(w_n14396_0[0]),.dout(n14988),.clk(gclk));
	jand g14699(.dina(w_asqrt11_14[2]),.dinb(n14988),.dout(n14989),.clk(gclk));
	jand g14700(.dina(w_n14989_0[1]),.dinb(w_n14401_0[0]),.dout(n14990),.clk(gclk));
	jor g14701(.dina(n14990),.dinb(w_n14400_0[0]),.dout(n14991),.clk(gclk));
	jand g14702(.dina(w_n14989_0[0]),.dinb(w_n14402_0[0]),.dout(n14992),.clk(gclk));
	jnot g14703(.din(n14992),.dout(n14993),.clk(gclk));
	jand g14704(.dina(n14993),.dinb(n14991),.dout(n14994),.clk(gclk));
	jnot g14705(.din(n14994),.dout(n14995),.clk(gclk));
	jor g14706(.dina(w_n14995_0[1]),.dinb(n14987),.dout(n14996),.clk(gclk));
	jand g14707(.dina(w_n14996_0[1]),.dinb(w_n14986_0[1]),.dout(n14997),.clk(gclk));
	jor g14708(.dina(n14997),.dinb(w_n6505_14[0]),.dout(n14998),.clk(gclk));
	jand g14709(.dina(w_n14986_0[0]),.dinb(w_n6505_13[2]),.dout(n14999),.clk(gclk));
	jand g14710(.dina(n14999),.dinb(w_n14996_0[0]),.dout(n15000),.clk(gclk));
	jnot g14711(.din(w_n14404_0[0]),.dout(n15001),.clk(gclk));
	jand g14712(.dina(w_asqrt11_14[1]),.dinb(n15001),.dout(n15002),.clk(gclk));
	jand g14713(.dina(w_n15002_0[1]),.dinb(w_n14411_0[0]),.dout(n15003),.clk(gclk));
	jor g14714(.dina(n15003),.dinb(w_n14409_0[0]),.dout(n15004),.clk(gclk));
	jand g14715(.dina(w_n15002_0[0]),.dinb(w_n14412_0[0]),.dout(n15005),.clk(gclk));
	jnot g14716(.din(n15005),.dout(n15006),.clk(gclk));
	jand g14717(.dina(n15006),.dinb(n15004),.dout(n15007),.clk(gclk));
	jnot g14718(.din(n15007),.dout(n15008),.clk(gclk));
	jor g14719(.dina(w_n15008_0[1]),.dinb(w_n15000_0[1]),.dout(n15009),.clk(gclk));
	jand g14720(.dina(n15009),.dinb(w_n14998_0[1]),.dout(n15010),.clk(gclk));
	jor g14721(.dina(w_n15010_0[1]),.dinb(w_n6500_10[2]),.dout(n15011),.clk(gclk));
	jxor g14722(.dina(w_n14413_0[0]),.dinb(w_n6505_13[1]),.dout(n15012),.clk(gclk));
	jor g14723(.dina(n15012),.dinb(w_n14821_18[0]),.dout(n15013),.clk(gclk));
	jxor g14724(.dina(n15013),.dinb(w_n14424_0[0]),.dout(n15014),.clk(gclk));
	jand g14725(.dina(w_n15010_0[0]),.dinb(w_n6500_10[1]),.dout(n15015),.clk(gclk));
	jor g14726(.dina(w_n15015_0[1]),.dinb(w_n15014_0[1]),.dout(n15016),.clk(gclk));
	jand g14727(.dina(w_n15016_0[2]),.dinb(w_n15011_0[2]),.dout(n15017),.clk(gclk));
	jor g14728(.dina(n15017),.dinb(w_n5793_14[1]),.dout(n15018),.clk(gclk));
	jnot g14729(.din(w_n14429_0[0]),.dout(n15019),.clk(gclk));
	jor g14730(.dina(n15019),.dinb(w_n14427_0[0]),.dout(n15020),.clk(gclk));
	jor g14731(.dina(n15020),.dinb(w_n14821_17[2]),.dout(n15021),.clk(gclk));
	jxor g14732(.dina(n15021),.dinb(w_n14438_0[0]),.dout(n15022),.clk(gclk));
	jand g14733(.dina(w_n15011_0[1]),.dinb(w_n5793_14[0]),.dout(n15023),.clk(gclk));
	jand g14734(.dina(n15023),.dinb(w_n15016_0[1]),.dout(n15024),.clk(gclk));
	jor g14735(.dina(w_n15024_0[1]),.dinb(w_n15022_0[1]),.dout(n15025),.clk(gclk));
	jand g14736(.dina(w_n15025_0[1]),.dinb(w_n15018_0[1]),.dout(n15026),.clk(gclk));
	jor g14737(.dina(w_n15026_0[2]),.dinb(w_n5788_11[1]),.dout(n15027),.clk(gclk));
	jand g14738(.dina(w_n15026_0[1]),.dinb(w_n5788_11[0]),.dout(n15028),.clk(gclk));
	jnot g14739(.din(w_n14441_0[0]),.dout(n15029),.clk(gclk));
	jand g14740(.dina(w_asqrt11_14[0]),.dinb(n15029),.dout(n15030),.clk(gclk));
	jand g14741(.dina(w_n15030_0[1]),.dinb(w_n14446_0[0]),.dout(n15031),.clk(gclk));
	jor g14742(.dina(n15031),.dinb(w_n14445_0[0]),.dout(n15032),.clk(gclk));
	jand g14743(.dina(w_n15030_0[0]),.dinb(w_n14447_0[0]),.dout(n15033),.clk(gclk));
	jnot g14744(.din(n15033),.dout(n15034),.clk(gclk));
	jand g14745(.dina(n15034),.dinb(n15032),.dout(n15035),.clk(gclk));
	jnot g14746(.din(n15035),.dout(n15036),.clk(gclk));
	jor g14747(.dina(w_n15036_0[1]),.dinb(n15028),.dout(n15037),.clk(gclk));
	jand g14748(.dina(w_n15037_0[1]),.dinb(w_n15027_0[1]),.dout(n15038),.clk(gclk));
	jor g14749(.dina(n15038),.dinb(w_n5121_14[1]),.dout(n15039),.clk(gclk));
	jand g14750(.dina(w_n15027_0[0]),.dinb(w_n5121_14[0]),.dout(n15040),.clk(gclk));
	jand g14751(.dina(n15040),.dinb(w_n15037_0[0]),.dout(n15041),.clk(gclk));
	jnot g14752(.din(w_n14449_0[0]),.dout(n15042),.clk(gclk));
	jand g14753(.dina(w_asqrt11_13[2]),.dinb(n15042),.dout(n15043),.clk(gclk));
	jand g14754(.dina(w_n15043_0[1]),.dinb(w_n14456_0[0]),.dout(n15044),.clk(gclk));
	jor g14755(.dina(n15044),.dinb(w_n14454_0[0]),.dout(n15045),.clk(gclk));
	jand g14756(.dina(w_n15043_0[0]),.dinb(w_n14457_0[0]),.dout(n15046),.clk(gclk));
	jnot g14757(.din(n15046),.dout(n15047),.clk(gclk));
	jand g14758(.dina(n15047),.dinb(n15045),.dout(n15048),.clk(gclk));
	jnot g14759(.din(n15048),.dout(n15049),.clk(gclk));
	jor g14760(.dina(w_n15049_0[1]),.dinb(w_n15041_0[1]),.dout(n15050),.clk(gclk));
	jand g14761(.dina(n15050),.dinb(w_n15039_0[1]),.dout(n15051),.clk(gclk));
	jor g14762(.dina(w_n15051_0[1]),.dinb(w_n5116_11[1]),.dout(n15052),.clk(gclk));
	jxor g14763(.dina(w_n14458_0[0]),.dinb(w_n5121_13[2]),.dout(n15053),.clk(gclk));
	jor g14764(.dina(n15053),.dinb(w_n14821_17[1]),.dout(n15054),.clk(gclk));
	jxor g14765(.dina(n15054),.dinb(w_n14469_0[0]),.dout(n15055),.clk(gclk));
	jand g14766(.dina(w_n15051_0[0]),.dinb(w_n5116_11[0]),.dout(n15056),.clk(gclk));
	jor g14767(.dina(w_n15056_0[1]),.dinb(w_n15055_0[1]),.dout(n15057),.clk(gclk));
	jand g14768(.dina(w_n15057_0[2]),.dinb(w_n15052_0[2]),.dout(n15058),.clk(gclk));
	jor g14769(.dina(n15058),.dinb(w_n4499_15[0]),.dout(n15059),.clk(gclk));
	jnot g14770(.din(w_n14474_0[0]),.dout(n15060),.clk(gclk));
	jor g14771(.dina(n15060),.dinb(w_n14472_0[0]),.dout(n15061),.clk(gclk));
	jor g14772(.dina(n15061),.dinb(w_n14821_17[0]),.dout(n15062),.clk(gclk));
	jxor g14773(.dina(n15062),.dinb(w_n14483_0[0]),.dout(n15063),.clk(gclk));
	jand g14774(.dina(w_n15052_0[1]),.dinb(w_n4499_14[2]),.dout(n15064),.clk(gclk));
	jand g14775(.dina(n15064),.dinb(w_n15057_0[1]),.dout(n15065),.clk(gclk));
	jor g14776(.dina(w_n15065_0[1]),.dinb(w_n15063_0[1]),.dout(n15066),.clk(gclk));
	jand g14777(.dina(w_n15066_0[1]),.dinb(w_n15059_0[1]),.dout(n15067),.clk(gclk));
	jor g14778(.dina(w_n15067_0[2]),.dinb(w_n4494_12[1]),.dout(n15068),.clk(gclk));
	jand g14779(.dina(w_n15067_0[1]),.dinb(w_n4494_12[0]),.dout(n15069),.clk(gclk));
	jnot g14780(.din(w_n14486_0[0]),.dout(n15070),.clk(gclk));
	jand g14781(.dina(w_asqrt11_13[1]),.dinb(n15070),.dout(n15071),.clk(gclk));
	jand g14782(.dina(w_n15071_0[1]),.dinb(w_n14491_0[0]),.dout(n15072),.clk(gclk));
	jor g14783(.dina(n15072),.dinb(w_n14490_0[0]),.dout(n15073),.clk(gclk));
	jand g14784(.dina(w_n15071_0[0]),.dinb(w_n14492_0[0]),.dout(n15074),.clk(gclk));
	jnot g14785(.din(n15074),.dout(n15075),.clk(gclk));
	jand g14786(.dina(n15075),.dinb(n15073),.dout(n15076),.clk(gclk));
	jnot g14787(.din(n15076),.dout(n15077),.clk(gclk));
	jor g14788(.dina(w_n15077_0[1]),.dinb(n15069),.dout(n15078),.clk(gclk));
	jand g14789(.dina(w_n15078_0[1]),.dinb(w_n15068_0[1]),.dout(n15079),.clk(gclk));
	jor g14790(.dina(n15079),.dinb(w_n3912_15[0]),.dout(n15080),.clk(gclk));
	jand g14791(.dina(w_n15068_0[0]),.dinb(w_n3912_14[2]),.dout(n15081),.clk(gclk));
	jand g14792(.dina(n15081),.dinb(w_n15078_0[0]),.dout(n15082),.clk(gclk));
	jnot g14793(.din(w_n14494_0[0]),.dout(n15083),.clk(gclk));
	jand g14794(.dina(w_asqrt11_13[0]),.dinb(n15083),.dout(n15084),.clk(gclk));
	jand g14795(.dina(w_n15084_0[1]),.dinb(w_n14501_0[0]),.dout(n15085),.clk(gclk));
	jor g14796(.dina(n15085),.dinb(w_n14499_0[0]),.dout(n15086),.clk(gclk));
	jand g14797(.dina(w_n15084_0[0]),.dinb(w_n14502_0[0]),.dout(n15087),.clk(gclk));
	jnot g14798(.din(n15087),.dout(n15088),.clk(gclk));
	jand g14799(.dina(n15088),.dinb(n15086),.dout(n15089),.clk(gclk));
	jnot g14800(.din(n15089),.dout(n15090),.clk(gclk));
	jor g14801(.dina(w_n15090_0[1]),.dinb(w_n15082_0[1]),.dout(n15091),.clk(gclk));
	jand g14802(.dina(n15091),.dinb(w_n15080_0[1]),.dout(n15092),.clk(gclk));
	jor g14803(.dina(w_n15092_0[1]),.dinb(w_n3907_12[1]),.dout(n15093),.clk(gclk));
	jxor g14804(.dina(w_n14503_0[0]),.dinb(w_n3912_14[1]),.dout(n15094),.clk(gclk));
	jor g14805(.dina(n15094),.dinb(w_n14821_16[2]),.dout(n15095),.clk(gclk));
	jxor g14806(.dina(n15095),.dinb(w_n14514_0[0]),.dout(n15096),.clk(gclk));
	jand g14807(.dina(w_n15092_0[0]),.dinb(w_n3907_12[0]),.dout(n15097),.clk(gclk));
	jor g14808(.dina(w_n15097_0[1]),.dinb(w_n15096_0[1]),.dout(n15098),.clk(gclk));
	jand g14809(.dina(w_n15098_0[2]),.dinb(w_n15093_0[2]),.dout(n15099),.clk(gclk));
	jor g14810(.dina(n15099),.dinb(w_n3376_15[2]),.dout(n15100),.clk(gclk));
	jnot g14811(.din(w_n14519_0[0]),.dout(n15101),.clk(gclk));
	jor g14812(.dina(n15101),.dinb(w_n14517_0[0]),.dout(n15102),.clk(gclk));
	jor g14813(.dina(n15102),.dinb(w_n14821_16[1]),.dout(n15103),.clk(gclk));
	jxor g14814(.dina(n15103),.dinb(w_n14528_0[0]),.dout(n15104),.clk(gclk));
	jand g14815(.dina(w_n15093_0[1]),.dinb(w_n3376_15[1]),.dout(n15105),.clk(gclk));
	jand g14816(.dina(n15105),.dinb(w_n15098_0[1]),.dout(n15106),.clk(gclk));
	jor g14817(.dina(w_n15106_0[1]),.dinb(w_n15104_0[1]),.dout(n15107),.clk(gclk));
	jand g14818(.dina(w_n15107_0[1]),.dinb(w_n15100_0[1]),.dout(n15108),.clk(gclk));
	jor g14819(.dina(w_n15108_0[2]),.dinb(w_n3371_13[0]),.dout(n15109),.clk(gclk));
	jand g14820(.dina(w_n15108_0[1]),.dinb(w_n3371_12[2]),.dout(n15110),.clk(gclk));
	jnot g14821(.din(w_n14531_0[0]),.dout(n15111),.clk(gclk));
	jand g14822(.dina(w_asqrt11_12[2]),.dinb(n15111),.dout(n15112),.clk(gclk));
	jand g14823(.dina(w_n15112_0[1]),.dinb(w_n14536_0[0]),.dout(n15113),.clk(gclk));
	jor g14824(.dina(n15113),.dinb(w_n14535_0[0]),.dout(n15114),.clk(gclk));
	jand g14825(.dina(w_n15112_0[0]),.dinb(w_n14537_0[0]),.dout(n15115),.clk(gclk));
	jnot g14826(.din(n15115),.dout(n15116),.clk(gclk));
	jand g14827(.dina(n15116),.dinb(n15114),.dout(n15117),.clk(gclk));
	jnot g14828(.din(n15117),.dout(n15118),.clk(gclk));
	jor g14829(.dina(w_n15118_0[1]),.dinb(n15110),.dout(n15119),.clk(gclk));
	jand g14830(.dina(w_n15119_0[1]),.dinb(w_n15109_0[1]),.dout(n15120),.clk(gclk));
	jor g14831(.dina(n15120),.dinb(w_n2875_15[2]),.dout(n15121),.clk(gclk));
	jand g14832(.dina(w_n15109_0[0]),.dinb(w_n2875_15[1]),.dout(n15122),.clk(gclk));
	jand g14833(.dina(n15122),.dinb(w_n15119_0[0]),.dout(n15123),.clk(gclk));
	jnot g14834(.din(w_n14539_0[0]),.dout(n15124),.clk(gclk));
	jand g14835(.dina(w_asqrt11_12[1]),.dinb(n15124),.dout(n15125),.clk(gclk));
	jand g14836(.dina(w_n15125_0[1]),.dinb(w_n14546_0[0]),.dout(n15126),.clk(gclk));
	jor g14837(.dina(n15126),.dinb(w_n14544_0[0]),.dout(n15127),.clk(gclk));
	jand g14838(.dina(w_n15125_0[0]),.dinb(w_n14547_0[0]),.dout(n15128),.clk(gclk));
	jnot g14839(.din(n15128),.dout(n15129),.clk(gclk));
	jand g14840(.dina(n15129),.dinb(n15127),.dout(n15130),.clk(gclk));
	jnot g14841(.din(n15130),.dout(n15131),.clk(gclk));
	jor g14842(.dina(w_n15131_0[1]),.dinb(w_n15123_0[1]),.dout(n15132),.clk(gclk));
	jand g14843(.dina(n15132),.dinb(w_n15121_0[1]),.dout(n15133),.clk(gclk));
	jor g14844(.dina(w_n15133_0[1]),.dinb(w_n2870_13[0]),.dout(n15134),.clk(gclk));
	jxor g14845(.dina(w_n14548_0[0]),.dinb(w_n2875_15[0]),.dout(n15135),.clk(gclk));
	jor g14846(.dina(n15135),.dinb(w_n14821_16[0]),.dout(n15136),.clk(gclk));
	jxor g14847(.dina(n15136),.dinb(w_n14559_0[0]),.dout(n15137),.clk(gclk));
	jand g14848(.dina(w_n15133_0[0]),.dinb(w_n2870_12[2]),.dout(n15138),.clk(gclk));
	jor g14849(.dina(w_n15138_0[1]),.dinb(w_n15137_0[1]),.dout(n15139),.clk(gclk));
	jand g14850(.dina(w_n15139_0[2]),.dinb(w_n15134_0[2]),.dout(n15140),.clk(gclk));
	jor g14851(.dina(n15140),.dinb(w_n2425_16[0]),.dout(n15141),.clk(gclk));
	jnot g14852(.din(w_n14564_0[0]),.dout(n15142),.clk(gclk));
	jor g14853(.dina(n15142),.dinb(w_n14562_0[0]),.dout(n15143),.clk(gclk));
	jor g14854(.dina(n15143),.dinb(w_n14821_15[2]),.dout(n15144),.clk(gclk));
	jxor g14855(.dina(n15144),.dinb(w_n14573_0[0]),.dout(n15145),.clk(gclk));
	jand g14856(.dina(w_n15134_0[1]),.dinb(w_n2425_15[2]),.dout(n15146),.clk(gclk));
	jand g14857(.dina(n15146),.dinb(w_n15139_0[1]),.dout(n15147),.clk(gclk));
	jor g14858(.dina(w_n15147_0[1]),.dinb(w_n15145_0[1]),.dout(n15148),.clk(gclk));
	jand g14859(.dina(w_n15148_0[1]),.dinb(w_n15141_0[1]),.dout(n15149),.clk(gclk));
	jor g14860(.dina(w_n15149_0[2]),.dinb(w_n2420_14[0]),.dout(n15150),.clk(gclk));
	jand g14861(.dina(w_n15149_0[1]),.dinb(w_n2420_13[2]),.dout(n15151),.clk(gclk));
	jnot g14862(.din(w_n14576_0[0]),.dout(n15152),.clk(gclk));
	jand g14863(.dina(w_asqrt11_12[0]),.dinb(n15152),.dout(n15153),.clk(gclk));
	jand g14864(.dina(w_n15153_0[1]),.dinb(w_n14581_0[0]),.dout(n15154),.clk(gclk));
	jor g14865(.dina(n15154),.dinb(w_n14580_0[0]),.dout(n15155),.clk(gclk));
	jand g14866(.dina(w_n15153_0[0]),.dinb(w_n14582_0[0]),.dout(n15156),.clk(gclk));
	jnot g14867(.din(n15156),.dout(n15157),.clk(gclk));
	jand g14868(.dina(n15157),.dinb(n15155),.dout(n15158),.clk(gclk));
	jnot g14869(.din(n15158),.dout(n15159),.clk(gclk));
	jor g14870(.dina(w_n15159_0[1]),.dinb(n15151),.dout(n15160),.clk(gclk));
	jand g14871(.dina(w_n15160_0[1]),.dinb(w_n15150_0[1]),.dout(n15161),.clk(gclk));
	jor g14872(.dina(n15161),.dinb(w_n2010_16[0]),.dout(n15162),.clk(gclk));
	jand g14873(.dina(w_n15150_0[0]),.dinb(w_n2010_15[2]),.dout(n15163),.clk(gclk));
	jand g14874(.dina(n15163),.dinb(w_n15160_0[0]),.dout(n15164),.clk(gclk));
	jnot g14875(.din(w_n14584_0[0]),.dout(n15165),.clk(gclk));
	jand g14876(.dina(w_asqrt11_11[2]),.dinb(n15165),.dout(n15166),.clk(gclk));
	jand g14877(.dina(w_n15166_0[1]),.dinb(w_n14591_0[0]),.dout(n15167),.clk(gclk));
	jor g14878(.dina(n15167),.dinb(w_n14589_0[0]),.dout(n15168),.clk(gclk));
	jand g14879(.dina(w_n15166_0[0]),.dinb(w_n14592_0[0]),.dout(n15169),.clk(gclk));
	jnot g14880(.din(n15169),.dout(n15170),.clk(gclk));
	jand g14881(.dina(n15170),.dinb(n15168),.dout(n15171),.clk(gclk));
	jnot g14882(.din(n15171),.dout(n15172),.clk(gclk));
	jor g14883(.dina(w_n15172_0[1]),.dinb(w_n15164_0[1]),.dout(n15173),.clk(gclk));
	jand g14884(.dina(n15173),.dinb(w_n15162_0[1]),.dout(n15174),.clk(gclk));
	jor g14885(.dina(w_n15174_0[1]),.dinb(w_n2005_14[0]),.dout(n15175),.clk(gclk));
	jxor g14886(.dina(w_n14593_0[0]),.dinb(w_n2010_15[1]),.dout(n15176),.clk(gclk));
	jor g14887(.dina(n15176),.dinb(w_n14821_15[1]),.dout(n15177),.clk(gclk));
	jxor g14888(.dina(n15177),.dinb(w_n14604_0[0]),.dout(n15178),.clk(gclk));
	jand g14889(.dina(w_n15174_0[0]),.dinb(w_n2005_13[2]),.dout(n15179),.clk(gclk));
	jor g14890(.dina(w_n15179_0[1]),.dinb(w_n15178_0[1]),.dout(n15180),.clk(gclk));
	jand g14891(.dina(w_n15180_0[2]),.dinb(w_n15175_0[2]),.dout(n15181),.clk(gclk));
	jor g14892(.dina(n15181),.dinb(w_n1646_16[2]),.dout(n15182),.clk(gclk));
	jnot g14893(.din(w_n14609_0[0]),.dout(n15183),.clk(gclk));
	jor g14894(.dina(n15183),.dinb(w_n14607_0[0]),.dout(n15184),.clk(gclk));
	jor g14895(.dina(n15184),.dinb(w_n14821_15[0]),.dout(n15185),.clk(gclk));
	jxor g14896(.dina(n15185),.dinb(w_n14618_0[0]),.dout(n15186),.clk(gclk));
	jand g14897(.dina(w_n15175_0[1]),.dinb(w_n1646_16[1]),.dout(n15187),.clk(gclk));
	jand g14898(.dina(n15187),.dinb(w_n15180_0[1]),.dout(n15188),.clk(gclk));
	jor g14899(.dina(w_n15188_0[1]),.dinb(w_n15186_0[1]),.dout(n15189),.clk(gclk));
	jand g14900(.dina(w_n15189_0[1]),.dinb(w_n15182_0[1]),.dout(n15190),.clk(gclk));
	jor g14901(.dina(w_n15190_0[2]),.dinb(w_n1641_14[2]),.dout(n15191),.clk(gclk));
	jand g14902(.dina(w_n15190_0[1]),.dinb(w_n1641_14[1]),.dout(n15192),.clk(gclk));
	jnot g14903(.din(w_n14621_0[0]),.dout(n15193),.clk(gclk));
	jand g14904(.dina(w_asqrt11_11[1]),.dinb(n15193),.dout(n15194),.clk(gclk));
	jand g14905(.dina(w_n15194_0[1]),.dinb(w_n14626_0[0]),.dout(n15195),.clk(gclk));
	jor g14906(.dina(n15195),.dinb(w_n14625_0[0]),.dout(n15196),.clk(gclk));
	jand g14907(.dina(w_n15194_0[0]),.dinb(w_n14627_0[0]),.dout(n15197),.clk(gclk));
	jnot g14908(.din(n15197),.dout(n15198),.clk(gclk));
	jand g14909(.dina(n15198),.dinb(n15196),.dout(n15199),.clk(gclk));
	jnot g14910(.din(n15199),.dout(n15200),.clk(gclk));
	jor g14911(.dina(w_n15200_0[1]),.dinb(n15192),.dout(n15201),.clk(gclk));
	jand g14912(.dina(w_n15201_0[1]),.dinb(w_n15191_0[1]),.dout(n15202),.clk(gclk));
	jor g14913(.dina(n15202),.dinb(w_n1317_16[2]),.dout(n15203),.clk(gclk));
	jand g14914(.dina(w_n15191_0[0]),.dinb(w_n1317_16[1]),.dout(n15204),.clk(gclk));
	jand g14915(.dina(n15204),.dinb(w_n15201_0[0]),.dout(n15205),.clk(gclk));
	jnot g14916(.din(w_n14629_0[0]),.dout(n15206),.clk(gclk));
	jand g14917(.dina(w_asqrt11_11[0]),.dinb(n15206),.dout(n15207),.clk(gclk));
	jand g14918(.dina(w_n15207_0[1]),.dinb(w_n14636_0[0]),.dout(n15208),.clk(gclk));
	jor g14919(.dina(n15208),.dinb(w_n14634_0[0]),.dout(n15209),.clk(gclk));
	jand g14920(.dina(w_n15207_0[0]),.dinb(w_n14637_0[0]),.dout(n15210),.clk(gclk));
	jnot g14921(.din(n15210),.dout(n15211),.clk(gclk));
	jand g14922(.dina(n15211),.dinb(n15209),.dout(n15212),.clk(gclk));
	jnot g14923(.din(n15212),.dout(n15213),.clk(gclk));
	jor g14924(.dina(w_n15213_0[1]),.dinb(w_n15205_0[1]),.dout(n15214),.clk(gclk));
	jand g14925(.dina(n15214),.dinb(w_n15203_0[1]),.dout(n15215),.clk(gclk));
	jor g14926(.dina(w_n15215_0[1]),.dinb(w_n1312_14[2]),.dout(n15216),.clk(gclk));
	jxor g14927(.dina(w_n14638_0[0]),.dinb(w_n1317_16[0]),.dout(n15217),.clk(gclk));
	jor g14928(.dina(n15217),.dinb(w_n14821_14[2]),.dout(n15218),.clk(gclk));
	jxor g14929(.dina(n15218),.dinb(w_n14649_0[0]),.dout(n15219),.clk(gclk));
	jand g14930(.dina(w_n15215_0[0]),.dinb(w_n1312_14[1]),.dout(n15220),.clk(gclk));
	jor g14931(.dina(w_n15220_0[1]),.dinb(w_n15219_0[1]),.dout(n15221),.clk(gclk));
	jand g14932(.dina(w_n15221_0[2]),.dinb(w_n15216_0[2]),.dout(n15222),.clk(gclk));
	jor g14933(.dina(n15222),.dinb(w_n1039_17[0]),.dout(n15223),.clk(gclk));
	jand g14934(.dina(w_n15216_0[1]),.dinb(w_n1039_16[2]),.dout(n15224),.clk(gclk));
	jand g14935(.dina(n15224),.dinb(w_n15221_0[1]),.dout(n15225),.clk(gclk));
	jnot g14936(.din(w_n14652_0[0]),.dout(n15226),.clk(gclk));
	jand g14937(.dina(w_asqrt11_10[2]),.dinb(n15226),.dout(n15227),.clk(gclk));
	jand g14938(.dina(w_n15227_0[1]),.dinb(w_n14659_0[0]),.dout(n15228),.clk(gclk));
	jor g14939(.dina(n15228),.dinb(w_n14657_0[0]),.dout(n15229),.clk(gclk));
	jand g14940(.dina(w_n15227_0[0]),.dinb(w_n14660_0[0]),.dout(n15230),.clk(gclk));
	jnot g14941(.din(n15230),.dout(n15231),.clk(gclk));
	jand g14942(.dina(n15231),.dinb(n15229),.dout(n15232),.clk(gclk));
	jnot g14943(.din(n15232),.dout(n15233),.clk(gclk));
	jor g14944(.dina(w_n15233_0[1]),.dinb(w_n15225_0[1]),.dout(n15234),.clk(gclk));
	jand g14945(.dina(n15234),.dinb(w_n15223_0[1]),.dout(n15235),.clk(gclk));
	jor g14946(.dina(w_n15235_0[2]),.dinb(w_n1034_15[2]),.dout(n15236),.clk(gclk));
	jnot g14947(.din(w_n14824_0[1]),.dout(n15237),.clk(gclk));
	jand g14948(.dina(w_n15235_0[1]),.dinb(w_n1034_15[1]),.dout(n15238),.clk(gclk));
	jor g14949(.dina(n15238),.dinb(n15237),.dout(n15239),.clk(gclk));
	jand g14950(.dina(w_n15239_0[1]),.dinb(w_n15236_0[1]),.dout(n15240),.clk(gclk));
	jor g14951(.dina(n15240),.dinb(w_n796_17[1]),.dout(n15241),.clk(gclk));
	jnot g14952(.din(w_n14669_0[0]),.dout(n15242),.clk(gclk));
	jor g14953(.dina(n15242),.dinb(w_n14667_0[0]),.dout(n15243),.clk(gclk));
	jor g14954(.dina(n15243),.dinb(w_n14821_14[1]),.dout(n15244),.clk(gclk));
	jxor g14955(.dina(n15244),.dinb(w_n14678_0[0]),.dout(n15245),.clk(gclk));
	jand g14956(.dina(w_n15236_0[0]),.dinb(w_n796_17[0]),.dout(n15246),.clk(gclk));
	jand g14957(.dina(n15246),.dinb(w_n15239_0[0]),.dout(n15247),.clk(gclk));
	jor g14958(.dina(w_n15247_0[1]),.dinb(w_n15245_0[1]),.dout(n15248),.clk(gclk));
	jand g14959(.dina(w_n15248_0[1]),.dinb(w_n15241_0[1]),.dout(n15249),.clk(gclk));
	jor g14960(.dina(w_n15249_0[1]),.dinb(w_n791_15[2]),.dout(n15250),.clk(gclk));
	jxor g14961(.dina(w_n14680_0[0]),.dinb(w_n796_16[2]),.dout(n15251),.clk(gclk));
	jor g14962(.dina(n15251),.dinb(w_n14821_14[0]),.dout(n15252),.clk(gclk));
	jxor g14963(.dina(n15252),.dinb(w_n14691_0[0]),.dout(n15253),.clk(gclk));
	jand g14964(.dina(w_n15249_0[0]),.dinb(w_n791_15[1]),.dout(n15254),.clk(gclk));
	jor g14965(.dina(w_n15254_0[1]),.dinb(w_n15253_0[1]),.dout(n15255),.clk(gclk));
	jand g14966(.dina(w_n15255_0[2]),.dinb(w_n15250_0[2]),.dout(n15256),.clk(gclk));
	jor g14967(.dina(n15256),.dinb(w_n595_17[2]),.dout(n15257),.clk(gclk));
	jnot g14968(.din(w_n14696_0[0]),.dout(n15258),.clk(gclk));
	jor g14969(.dina(n15258),.dinb(w_n14694_0[0]),.dout(n15259),.clk(gclk));
	jor g14970(.dina(n15259),.dinb(w_n14821_13[2]),.dout(n15260),.clk(gclk));
	jxor g14971(.dina(n15260),.dinb(w_n14705_0[0]),.dout(n15261),.clk(gclk));
	jand g14972(.dina(w_n15250_0[1]),.dinb(w_n595_17[1]),.dout(n15262),.clk(gclk));
	jand g14973(.dina(n15262),.dinb(w_n15255_0[1]),.dout(n15263),.clk(gclk));
	jor g14974(.dina(w_n15263_0[1]),.dinb(w_n15261_0[1]),.dout(n15264),.clk(gclk));
	jand g14975(.dina(w_n15264_0[1]),.dinb(w_n15257_0[1]),.dout(n15265),.clk(gclk));
	jor g14976(.dina(w_n15265_0[2]),.dinb(w_n590_16[1]),.dout(n15266),.clk(gclk));
	jand g14977(.dina(w_n15265_0[1]),.dinb(w_n590_16[0]),.dout(n15267),.clk(gclk));
	jnot g14978(.din(w_n14708_0[0]),.dout(n15268),.clk(gclk));
	jand g14979(.dina(w_asqrt11_10[1]),.dinb(n15268),.dout(n15269),.clk(gclk));
	jand g14980(.dina(w_n15269_0[1]),.dinb(w_n14713_0[0]),.dout(n15270),.clk(gclk));
	jor g14981(.dina(n15270),.dinb(w_n14712_0[0]),.dout(n15271),.clk(gclk));
	jand g14982(.dina(w_n15269_0[0]),.dinb(w_n14714_0[0]),.dout(n15272),.clk(gclk));
	jnot g14983(.din(n15272),.dout(n15273),.clk(gclk));
	jand g14984(.dina(n15273),.dinb(n15271),.dout(n15274),.clk(gclk));
	jnot g14985(.din(n15274),.dout(n15275),.clk(gclk));
	jor g14986(.dina(w_n15275_0[1]),.dinb(n15267),.dout(n15276),.clk(gclk));
	jand g14987(.dina(w_n15276_0[1]),.dinb(w_n15266_0[1]),.dout(n15277),.clk(gclk));
	jor g14988(.dina(n15277),.dinb(w_n430_17[2]),.dout(n15278),.clk(gclk));
	jand g14989(.dina(w_n15266_0[0]),.dinb(w_n430_17[1]),.dout(n15279),.clk(gclk));
	jand g14990(.dina(n15279),.dinb(w_n15276_0[0]),.dout(n15280),.clk(gclk));
	jnot g14991(.din(w_n14716_0[0]),.dout(n15281),.clk(gclk));
	jand g14992(.dina(w_asqrt11_10[0]),.dinb(n15281),.dout(n15282),.clk(gclk));
	jand g14993(.dina(w_n15282_0[1]),.dinb(w_n14723_0[0]),.dout(n15283),.clk(gclk));
	jor g14994(.dina(n15283),.dinb(w_n14721_0[0]),.dout(n15284),.clk(gclk));
	jand g14995(.dina(w_n15282_0[0]),.dinb(w_n14724_0[0]),.dout(n15285),.clk(gclk));
	jnot g14996(.din(n15285),.dout(n15286),.clk(gclk));
	jand g14997(.dina(n15286),.dinb(n15284),.dout(n15287),.clk(gclk));
	jnot g14998(.din(n15287),.dout(n15288),.clk(gclk));
	jor g14999(.dina(w_n15288_0[1]),.dinb(w_n15280_0[1]),.dout(n15289),.clk(gclk));
	jand g15000(.dina(n15289),.dinb(w_n15278_0[1]),.dout(n15290),.clk(gclk));
	jor g15001(.dina(w_n15290_0[1]),.dinb(w_n425_16[1]),.dout(n15291),.clk(gclk));
	jxor g15002(.dina(w_n14725_0[0]),.dinb(w_n430_17[0]),.dout(n15292),.clk(gclk));
	jor g15003(.dina(n15292),.dinb(w_n14821_13[1]),.dout(n15293),.clk(gclk));
	jxor g15004(.dina(n15293),.dinb(w_n14736_0[0]),.dout(n15294),.clk(gclk));
	jand g15005(.dina(w_n15290_0[0]),.dinb(w_n425_16[0]),.dout(n15295),.clk(gclk));
	jor g15006(.dina(w_n15295_0[1]),.dinb(w_n15294_0[1]),.dout(n15296),.clk(gclk));
	jand g15007(.dina(w_n15296_0[2]),.dinb(w_n15291_0[2]),.dout(n15297),.clk(gclk));
	jor g15008(.dina(n15297),.dinb(w_n305_18[0]),.dout(n15298),.clk(gclk));
	jnot g15009(.din(w_n14741_0[0]),.dout(n15299),.clk(gclk));
	jor g15010(.dina(n15299),.dinb(w_n14739_0[0]),.dout(n15300),.clk(gclk));
	jor g15011(.dina(n15300),.dinb(w_n14821_13[0]),.dout(n15301),.clk(gclk));
	jxor g15012(.dina(n15301),.dinb(w_n14750_0[0]),.dout(n15302),.clk(gclk));
	jand g15013(.dina(w_n15291_0[1]),.dinb(w_n305_17[2]),.dout(n15303),.clk(gclk));
	jand g15014(.dina(n15303),.dinb(w_n15296_0[1]),.dout(n15304),.clk(gclk));
	jor g15015(.dina(w_n15304_0[1]),.dinb(w_n15302_0[1]),.dout(n15305),.clk(gclk));
	jand g15016(.dina(w_n15305_0[1]),.dinb(w_n15298_0[1]),.dout(n15306),.clk(gclk));
	jor g15017(.dina(w_n15306_0[2]),.dinb(w_n290_17[2]),.dout(n15307),.clk(gclk));
	jand g15018(.dina(w_n15306_0[1]),.dinb(w_n290_17[1]),.dout(n15308),.clk(gclk));
	jnot g15019(.din(w_n14753_0[0]),.dout(n15309),.clk(gclk));
	jand g15020(.dina(w_asqrt11_9[2]),.dinb(n15309),.dout(n15310),.clk(gclk));
	jand g15021(.dina(w_n15310_0[1]),.dinb(w_n14758_0[0]),.dout(n15311),.clk(gclk));
	jor g15022(.dina(n15311),.dinb(w_n14757_0[0]),.dout(n15312),.clk(gclk));
	jand g15023(.dina(w_n15310_0[0]),.dinb(w_n14759_0[0]),.dout(n15313),.clk(gclk));
	jnot g15024(.din(n15313),.dout(n15314),.clk(gclk));
	jand g15025(.dina(n15314),.dinb(n15312),.dout(n15315),.clk(gclk));
	jnot g15026(.din(n15315),.dout(n15316),.clk(gclk));
	jor g15027(.dina(w_n15316_0[1]),.dinb(n15308),.dout(n15317),.clk(gclk));
	jand g15028(.dina(w_n15317_0[1]),.dinb(w_n15307_0[1]),.dout(n15318),.clk(gclk));
	jor g15029(.dina(n15318),.dinb(w_n223_18[0]),.dout(n15319),.clk(gclk));
	jand g15030(.dina(w_n15307_0[0]),.dinb(w_n223_17[2]),.dout(n15320),.clk(gclk));
	jand g15031(.dina(n15320),.dinb(w_n15317_0[0]),.dout(n15321),.clk(gclk));
	jnot g15032(.din(w_n14761_0[0]),.dout(n15322),.clk(gclk));
	jand g15033(.dina(w_asqrt11_9[1]),.dinb(n15322),.dout(n15323),.clk(gclk));
	jand g15034(.dina(w_n15323_0[1]),.dinb(w_n14768_0[0]),.dout(n15324),.clk(gclk));
	jor g15035(.dina(n15324),.dinb(w_n14766_0[0]),.dout(n15325),.clk(gclk));
	jand g15036(.dina(w_n15323_0[0]),.dinb(w_n14769_0[0]),.dout(n15326),.clk(gclk));
	jnot g15037(.din(n15326),.dout(n15327),.clk(gclk));
	jand g15038(.dina(n15327),.dinb(n15325),.dout(n15328),.clk(gclk));
	jnot g15039(.din(n15328),.dout(n15329),.clk(gclk));
	jor g15040(.dina(w_n15329_0[1]),.dinb(w_n15321_0[1]),.dout(n15330),.clk(gclk));
	jand g15041(.dina(n15330),.dinb(w_n15319_0[1]),.dout(n15331),.clk(gclk));
	jor g15042(.dina(w_n15331_0[2]),.dinb(w_n199_20[1]),.dout(n15332),.clk(gclk));
	jand g15043(.dina(w_n15331_0[1]),.dinb(w_n199_20[0]),.dout(n15333),.clk(gclk));
	jxor g15044(.dina(w_n14770_0[0]),.dinb(w_n223_17[1]),.dout(n15334),.clk(gclk));
	jor g15045(.dina(n15334),.dinb(w_n14821_12[2]),.dout(n15335),.clk(gclk));
	jxor g15046(.dina(n15335),.dinb(w_n14781_0[0]),.dout(n15336),.clk(gclk));
	jor g15047(.dina(w_n15336_0[1]),.dinb(n15333),.dout(n15337),.clk(gclk));
	jand g15048(.dina(n15337),.dinb(n15332),.dout(n15338),.clk(gclk));
	jnot g15049(.din(w_n14786_0[0]),.dout(n15339),.clk(gclk));
	jor g15050(.dina(n15339),.dinb(w_n14784_0[0]),.dout(n15340),.clk(gclk));
	jor g15051(.dina(n15340),.dinb(w_n14821_12[1]),.dout(n15341),.clk(gclk));
	jxor g15052(.dina(n15341),.dinb(w_n14795_0[0]),.dout(n15342),.clk(gclk));
	jand g15053(.dina(w_asqrt11_9[0]),.dinb(w_n14809_0[1]),.dout(n15343),.clk(gclk));
	jand g15054(.dina(w_n15343_0[1]),.dinb(w_n14797_1[0]),.dout(n15344),.clk(gclk));
	jor g15055(.dina(n15344),.dinb(w_n14843_0[0]),.dout(n15345),.clk(gclk));
	jor g15056(.dina(n15345),.dinb(w_n15342_0[2]),.dout(n15346),.clk(gclk));
	jor g15057(.dina(n15346),.dinb(w_n15338_0[2]),.dout(n15347),.clk(gclk));
	jand g15058(.dina(n15347),.dinb(w_n194_19[1]),.dout(n15348),.clk(gclk));
	jand g15059(.dina(w_n15342_0[1]),.dinb(w_n15338_0[1]),.dout(n15349),.clk(gclk));
	jor g15060(.dina(w_n15343_0[0]),.dinb(w_n14797_0[2]),.dout(n15350),.clk(gclk));
	jand g15061(.dina(w_n14809_0[0]),.dinb(w_n14797_0[1]),.dout(n15351),.clk(gclk));
	jor g15062(.dina(n15351),.dinb(w_n194_19[0]),.dout(n15352),.clk(gclk));
	jnot g15063(.din(n15352),.dout(n15353),.clk(gclk));
	jand g15064(.dina(n15353),.dinb(n15350),.dout(n15354),.clk(gclk));
	jor g15065(.dina(w_n15354_0[1]),.dinb(w_n15349_0[2]),.dout(n15357),.clk(gclk));
	jor g15066(.dina(n15357),.dinb(w_n15348_0[1]),.dout(asqrt_fa_11),.clk(gclk));
	jxor g15067(.dina(w_n15235_0[0]),.dinb(w_n1034_15[0]),.dout(n15359),.clk(gclk));
	jand g15068(.dina(n15359),.dinb(w_asqrt10_31),.dout(n15360),.clk(gclk));
	jxor g15069(.dina(n15360),.dinb(w_n14824_0[0]),.dout(n15361),.clk(gclk));
	jnot g15070(.din(w_n15361_0[1]),.dout(n15362),.clk(gclk));
	jand g15071(.dina(w_asqrt10_30[2]),.dinb(w_a20_0[0]),.dout(n15363),.clk(gclk));
	jnot g15072(.din(w_a18_0[1]),.dout(n15364),.clk(gclk));
	jnot g15073(.din(w_a19_0[1]),.dout(n15365),.clk(gclk));
	jand g15074(.dina(w_n14826_1[0]),.dinb(w_n15365_0[1]),.dout(n15366),.clk(gclk));
	jand g15075(.dina(n15366),.dinb(w_n15364_1[1]),.dout(n15367),.clk(gclk));
	jor g15076(.dina(n15367),.dinb(n15363),.dout(n15368),.clk(gclk));
	jand g15077(.dina(w_n15368_0[2]),.dinb(w_asqrt11_8[2]),.dout(n15369),.clk(gclk));
	jand g15078(.dina(w_asqrt10_30[1]),.dinb(w_n14826_0[2]),.dout(n15370),.clk(gclk));
	jxor g15079(.dina(w_n15370_0[1]),.dinb(w_n14827_0[1]),.dout(n15371),.clk(gclk));
	jor g15080(.dina(w_n15368_0[1]),.dinb(w_asqrt11_8[1]),.dout(n15372),.clk(gclk));
	jand g15081(.dina(n15372),.dinb(w_n15371_0[1]),.dout(n15373),.clk(gclk));
	jor g15082(.dina(w_n15373_0[1]),.dinb(w_n15369_0[1]),.dout(n15374),.clk(gclk));
	jand g15083(.dina(n15374),.dinb(w_asqrt12_13[1]),.dout(n15375),.clk(gclk));
	jor g15084(.dina(w_n15369_0[0]),.dinb(w_asqrt12_13[0]),.dout(n15376),.clk(gclk));
	jor g15085(.dina(n15376),.dinb(w_n15373_0[0]),.dout(n15377),.clk(gclk));
	jand g15086(.dina(w_n15370_0[0]),.dinb(w_n14827_0[0]),.dout(n15378),.clk(gclk));
	jnot g15087(.din(w_n15348_0[0]),.dout(n15379),.clk(gclk));
	jnot g15088(.din(w_n15349_0[1]),.dout(n15380),.clk(gclk));
	jnot g15089(.din(w_n15354_0[0]),.dout(n15381),.clk(gclk));
	jand g15090(.dina(n15381),.dinb(w_asqrt11_8[0]),.dout(n15382),.clk(gclk));
	jand g15091(.dina(n15382),.dinb(n15380),.dout(n15383),.clk(gclk));
	jand g15092(.dina(n15383),.dinb(n15379),.dout(n15384),.clk(gclk));
	jor g15093(.dina(n15384),.dinb(n15378),.dout(n15385),.clk(gclk));
	jxor g15094(.dina(n15385),.dinb(w_n14248_0[1]),.dout(n15386),.clk(gclk));
	jand g15095(.dina(w_n15386_0[1]),.dinb(w_n15377_0[1]),.dout(n15387),.clk(gclk));
	jor g15096(.dina(n15387),.dinb(w_n15375_0[1]),.dout(n15388),.clk(gclk));
	jand g15097(.dina(w_n15388_0[2]),.dinb(w_asqrt13_8[2]),.dout(n15389),.clk(gclk));
	jor g15098(.dina(w_n15388_0[1]),.dinb(w_asqrt13_8[1]),.dout(n15390),.clk(gclk));
	jxor g15099(.dina(w_n14831_0[0]),.dinb(w_n14816_7[1]),.dout(n15391),.clk(gclk));
	jand g15100(.dina(n15391),.dinb(w_asqrt10_30[0]),.dout(n15392),.clk(gclk));
	jxor g15101(.dina(n15392),.dinb(w_n14834_0[0]),.dout(n15393),.clk(gclk));
	jnot g15102(.din(w_n15393_0[1]),.dout(n15394),.clk(gclk));
	jand g15103(.dina(n15394),.dinb(n15390),.dout(n15395),.clk(gclk));
	jor g15104(.dina(w_n15395_0[1]),.dinb(w_n15389_0[1]),.dout(n15396),.clk(gclk));
	jand g15105(.dina(n15396),.dinb(w_asqrt14_13[1]),.dout(n15397),.clk(gclk));
	jnot g15106(.din(w_n14840_0[0]),.dout(n15398),.clk(gclk));
	jand g15107(.dina(n15398),.dinb(w_n14838_0[0]),.dout(n15399),.clk(gclk));
	jand g15108(.dina(n15399),.dinb(w_asqrt10_29[2]),.dout(n15400),.clk(gclk));
	jxor g15109(.dina(n15400),.dinb(w_n14848_0[0]),.dout(n15401),.clk(gclk));
	jnot g15110(.din(n15401),.dout(n15402),.clk(gclk));
	jor g15111(.dina(w_n15389_0[0]),.dinb(w_asqrt14_13[0]),.dout(n15403),.clk(gclk));
	jor g15112(.dina(n15403),.dinb(w_n15395_0[0]),.dout(n15404),.clk(gclk));
	jand g15113(.dina(w_n15404_0[1]),.dinb(w_n15402_0[1]),.dout(n15405),.clk(gclk));
	jor g15114(.dina(w_n15405_0[1]),.dinb(w_n15397_0[1]),.dout(n15406),.clk(gclk));
	jand g15115(.dina(w_n15406_0[2]),.dinb(w_asqrt15_8[2]),.dout(n15407),.clk(gclk));
	jor g15116(.dina(w_n15406_0[1]),.dinb(w_asqrt15_8[1]),.dout(n15408),.clk(gclk));
	jnot g15117(.din(w_n14855_0[0]),.dout(n15409),.clk(gclk));
	jxor g15118(.dina(w_n14850_0[0]),.dinb(w_n13718_7[1]),.dout(n15410),.clk(gclk));
	jand g15119(.dina(n15410),.dinb(w_asqrt10_29[1]),.dout(n15411),.clk(gclk));
	jxor g15120(.dina(n15411),.dinb(n15409),.dout(n15412),.clk(gclk));
	jand g15121(.dina(w_n15412_0[1]),.dinb(n15408),.dout(n15413),.clk(gclk));
	jor g15122(.dina(w_n15413_0[1]),.dinb(w_n15407_0[1]),.dout(n15414),.clk(gclk));
	jand g15123(.dina(n15414),.dinb(w_asqrt16_13[1]),.dout(n15415),.clk(gclk));
	jor g15124(.dina(w_n15407_0[0]),.dinb(w_asqrt16_13[0]),.dout(n15416),.clk(gclk));
	jor g15125(.dina(n15416),.dinb(w_n15413_0[0]),.dout(n15417),.clk(gclk));
	jnot g15126(.din(w_n14862_0[0]),.dout(n15418),.clk(gclk));
	jnot g15127(.din(w_n14864_0[0]),.dout(n15419),.clk(gclk));
	jand g15128(.dina(w_asqrt10_29[0]),.dinb(w_n14858_0[0]),.dout(n15420),.clk(gclk));
	jand g15129(.dina(w_n15420_0[1]),.dinb(n15419),.dout(n15421),.clk(gclk));
	jor g15130(.dina(n15421),.dinb(n15418),.dout(n15422),.clk(gclk));
	jnot g15131(.din(w_n14865_0[0]),.dout(n15423),.clk(gclk));
	jand g15132(.dina(w_n15420_0[0]),.dinb(n15423),.dout(n15424),.clk(gclk));
	jnot g15133(.din(n15424),.dout(n15425),.clk(gclk));
	jand g15134(.dina(n15425),.dinb(n15422),.dout(n15426),.clk(gclk));
	jand g15135(.dina(w_n15426_0[1]),.dinb(w_n15417_0[1]),.dout(n15427),.clk(gclk));
	jor g15136(.dina(n15427),.dinb(w_n15415_0[1]),.dout(n15428),.clk(gclk));
	jand g15137(.dina(w_n15428_0[2]),.dinb(w_asqrt17_9[0]),.dout(n15429),.clk(gclk));
	jor g15138(.dina(w_n15428_0[1]),.dinb(w_asqrt17_8[2]),.dout(n15430),.clk(gclk));
	jxor g15139(.dina(w_n14866_0[0]),.dinb(w_n12670_7[2]),.dout(n15431),.clk(gclk));
	jand g15140(.dina(n15431),.dinb(w_asqrt10_28[2]),.dout(n15432),.clk(gclk));
	jxor g15141(.dina(n15432),.dinb(w_n14871_0[0]),.dout(n15433),.clk(gclk));
	jand g15142(.dina(w_n15433_0[1]),.dinb(n15430),.dout(n15434),.clk(gclk));
	jor g15143(.dina(w_n15434_0[1]),.dinb(w_n15429_0[1]),.dout(n15435),.clk(gclk));
	jand g15144(.dina(n15435),.dinb(w_asqrt18_13[1]),.dout(n15436),.clk(gclk));
	jnot g15145(.din(w_n14877_0[0]),.dout(n15437),.clk(gclk));
	jand g15146(.dina(n15437),.dinb(w_n14875_0[0]),.dout(n15438),.clk(gclk));
	jand g15147(.dina(n15438),.dinb(w_asqrt10_28[1]),.dout(n15439),.clk(gclk));
	jxor g15148(.dina(n15439),.dinb(w_n14886_0[0]),.dout(n15440),.clk(gclk));
	jnot g15149(.din(n15440),.dout(n15441),.clk(gclk));
	jor g15150(.dina(w_n15429_0[0]),.dinb(w_asqrt18_13[0]),.dout(n15442),.clk(gclk));
	jor g15151(.dina(n15442),.dinb(w_n15434_0[0]),.dout(n15443),.clk(gclk));
	jand g15152(.dina(w_n15443_0[1]),.dinb(w_n15441_0[1]),.dout(n15444),.clk(gclk));
	jor g15153(.dina(w_n15444_0[1]),.dinb(w_n15436_0[1]),.dout(n15445),.clk(gclk));
	jand g15154(.dina(w_n15445_0[2]),.dinb(w_asqrt19_9[0]),.dout(n15446),.clk(gclk));
	jor g15155(.dina(w_n15445_0[1]),.dinb(w_asqrt19_8[2]),.dout(n15447),.clk(gclk));
	jxor g15156(.dina(w_n14888_0[0]),.dinb(w_n11657_7[2]),.dout(n15448),.clk(gclk));
	jand g15157(.dina(n15448),.dinb(w_asqrt10_28[0]),.dout(n15449),.clk(gclk));
	jxor g15158(.dina(n15449),.dinb(w_n14894_0[0]),.dout(n15450),.clk(gclk));
	jand g15159(.dina(w_n15450_0[1]),.dinb(n15447),.dout(n15451),.clk(gclk));
	jor g15160(.dina(w_n15451_0[1]),.dinb(w_n15446_0[1]),.dout(n15452),.clk(gclk));
	jand g15161(.dina(n15452),.dinb(w_asqrt20_13[1]),.dout(n15453),.clk(gclk));
	jor g15162(.dina(w_n15446_0[0]),.dinb(w_asqrt20_13[0]),.dout(n15454),.clk(gclk));
	jor g15163(.dina(n15454),.dinb(w_n15451_0[0]),.dout(n15455),.clk(gclk));
	jnot g15164(.din(w_n14902_0[0]),.dout(n15456),.clk(gclk));
	jnot g15165(.din(w_n14904_0[0]),.dout(n15457),.clk(gclk));
	jand g15166(.dina(w_asqrt10_27[2]),.dinb(w_n14898_0[0]),.dout(n15458),.clk(gclk));
	jand g15167(.dina(w_n15458_0[1]),.dinb(n15457),.dout(n15459),.clk(gclk));
	jor g15168(.dina(n15459),.dinb(n15456),.dout(n15460),.clk(gclk));
	jnot g15169(.din(w_n14905_0[0]),.dout(n15461),.clk(gclk));
	jand g15170(.dina(w_n15458_0[0]),.dinb(n15461),.dout(n15462),.clk(gclk));
	jnot g15171(.din(n15462),.dout(n15463),.clk(gclk));
	jand g15172(.dina(n15463),.dinb(n15460),.dout(n15464),.clk(gclk));
	jand g15173(.dina(w_n15464_0[1]),.dinb(w_n15455_0[1]),.dout(n15465),.clk(gclk));
	jor g15174(.dina(n15465),.dinb(w_n15453_0[1]),.dout(n15466),.clk(gclk));
	jand g15175(.dina(w_n15466_0[1]),.dinb(w_asqrt21_9[1]),.dout(n15467),.clk(gclk));
	jxor g15176(.dina(w_n14906_0[0]),.dinb(w_n10696_8[1]),.dout(n15468),.clk(gclk));
	jand g15177(.dina(n15468),.dinb(w_asqrt10_27[1]),.dout(n15469),.clk(gclk));
	jxor g15178(.dina(n15469),.dinb(w_n14913_0[0]),.dout(n15470),.clk(gclk));
	jnot g15179(.din(n15470),.dout(n15471),.clk(gclk));
	jor g15180(.dina(w_n15466_0[0]),.dinb(w_asqrt21_9[0]),.dout(n15472),.clk(gclk));
	jand g15181(.dina(w_n15472_0[1]),.dinb(w_n15471_0[1]),.dout(n15473),.clk(gclk));
	jor g15182(.dina(w_n15473_0[2]),.dinb(w_n15467_0[2]),.dout(n15474),.clk(gclk));
	jand g15183(.dina(n15474),.dinb(w_asqrt22_13[1]),.dout(n15475),.clk(gclk));
	jnot g15184(.din(w_n14918_0[0]),.dout(n15476),.clk(gclk));
	jand g15185(.dina(n15476),.dinb(w_n14916_0[0]),.dout(n15477),.clk(gclk));
	jand g15186(.dina(n15477),.dinb(w_asqrt10_27[0]),.dout(n15478),.clk(gclk));
	jxor g15187(.dina(n15478),.dinb(w_n14926_0[0]),.dout(n15479),.clk(gclk));
	jnot g15188(.din(n15479),.dout(n15480),.clk(gclk));
	jor g15189(.dina(w_n15467_0[1]),.dinb(w_asqrt22_13[0]),.dout(n15481),.clk(gclk));
	jor g15190(.dina(n15481),.dinb(w_n15473_0[1]),.dout(n15482),.clk(gclk));
	jand g15191(.dina(w_n15482_0[1]),.dinb(w_n15480_0[1]),.dout(n15483),.clk(gclk));
	jor g15192(.dina(w_n15483_0[1]),.dinb(w_n15475_0[1]),.dout(n15484),.clk(gclk));
	jand g15193(.dina(w_n15484_0[2]),.dinb(w_asqrt23_9[1]),.dout(n15485),.clk(gclk));
	jor g15194(.dina(w_n15484_0[1]),.dinb(w_asqrt23_9[0]),.dout(n15486),.clk(gclk));
	jnot g15195(.din(w_n14932_0[0]),.dout(n15487),.clk(gclk));
	jnot g15196(.din(w_n14933_0[0]),.dout(n15488),.clk(gclk));
	jand g15197(.dina(w_asqrt10_26[2]),.dinb(w_n14929_0[0]),.dout(n15489),.clk(gclk));
	jand g15198(.dina(w_n15489_0[1]),.dinb(n15488),.dout(n15490),.clk(gclk));
	jor g15199(.dina(n15490),.dinb(n15487),.dout(n15491),.clk(gclk));
	jnot g15200(.din(w_n14934_0[0]),.dout(n15492),.clk(gclk));
	jand g15201(.dina(w_n15489_0[0]),.dinb(n15492),.dout(n15493),.clk(gclk));
	jnot g15202(.din(n15493),.dout(n15494),.clk(gclk));
	jand g15203(.dina(n15494),.dinb(n15491),.dout(n15495),.clk(gclk));
	jand g15204(.dina(w_n15495_0[1]),.dinb(n15486),.dout(n15496),.clk(gclk));
	jor g15205(.dina(w_n15496_0[1]),.dinb(w_n15485_0[1]),.dout(n15497),.clk(gclk));
	jand g15206(.dina(n15497),.dinb(w_asqrt24_13[1]),.dout(n15498),.clk(gclk));
	jor g15207(.dina(w_n15485_0[0]),.dinb(w_asqrt24_13[0]),.dout(n15499),.clk(gclk));
	jor g15208(.dina(n15499),.dinb(w_n15496_0[0]),.dout(n15500),.clk(gclk));
	jnot g15209(.din(w_n14940_0[0]),.dout(n15501),.clk(gclk));
	jnot g15210(.din(w_n14942_0[0]),.dout(n15502),.clk(gclk));
	jand g15211(.dina(w_asqrt10_26[1]),.dinb(w_n14936_0[0]),.dout(n15503),.clk(gclk));
	jand g15212(.dina(w_n15503_0[1]),.dinb(n15502),.dout(n15504),.clk(gclk));
	jor g15213(.dina(n15504),.dinb(n15501),.dout(n15505),.clk(gclk));
	jnot g15214(.din(w_n14943_0[0]),.dout(n15506),.clk(gclk));
	jand g15215(.dina(w_n15503_0[0]),.dinb(n15506),.dout(n15507),.clk(gclk));
	jnot g15216(.din(n15507),.dout(n15508),.clk(gclk));
	jand g15217(.dina(n15508),.dinb(n15505),.dout(n15509),.clk(gclk));
	jand g15218(.dina(w_n15509_0[1]),.dinb(w_n15500_0[1]),.dout(n15510),.clk(gclk));
	jor g15219(.dina(n15510),.dinb(w_n15498_0[1]),.dout(n15511),.clk(gclk));
	jand g15220(.dina(w_n15511_0[1]),.dinb(w_asqrt25_9[2]),.dout(n15512),.clk(gclk));
	jxor g15221(.dina(w_n14944_0[0]),.dinb(w_n8893_9[0]),.dout(n15513),.clk(gclk));
	jand g15222(.dina(n15513),.dinb(w_asqrt10_26[0]),.dout(n15514),.clk(gclk));
	jxor g15223(.dina(n15514),.dinb(w_n14954_0[0]),.dout(n15515),.clk(gclk));
	jnot g15224(.din(n15515),.dout(n15516),.clk(gclk));
	jor g15225(.dina(w_n15511_0[0]),.dinb(w_asqrt25_9[1]),.dout(n15517),.clk(gclk));
	jand g15226(.dina(w_n15517_0[1]),.dinb(w_n15516_0[1]),.dout(n15518),.clk(gclk));
	jor g15227(.dina(w_n15518_0[2]),.dinb(w_n15512_0[2]),.dout(n15519),.clk(gclk));
	jand g15228(.dina(n15519),.dinb(w_asqrt26_13[1]),.dout(n15520),.clk(gclk));
	jnot g15229(.din(w_n14959_0[0]),.dout(n15521),.clk(gclk));
	jand g15230(.dina(n15521),.dinb(w_n14957_0[0]),.dout(n15522),.clk(gclk));
	jand g15231(.dina(n15522),.dinb(w_asqrt10_25[2]),.dout(n15523),.clk(gclk));
	jxor g15232(.dina(n15523),.dinb(w_n14967_0[0]),.dout(n15524),.clk(gclk));
	jnot g15233(.din(n15524),.dout(n15525),.clk(gclk));
	jor g15234(.dina(w_n15512_0[1]),.dinb(w_asqrt26_13[0]),.dout(n15526),.clk(gclk));
	jor g15235(.dina(n15526),.dinb(w_n15518_0[1]),.dout(n15527),.clk(gclk));
	jand g15236(.dina(w_n15527_0[1]),.dinb(w_n15525_0[1]),.dout(n15528),.clk(gclk));
	jor g15237(.dina(w_n15528_0[1]),.dinb(w_n15520_0[1]),.dout(n15529),.clk(gclk));
	jand g15238(.dina(w_n15529_0[2]),.dinb(w_asqrt27_9[2]),.dout(n15530),.clk(gclk));
	jor g15239(.dina(w_n15529_0[1]),.dinb(w_asqrt27_9[1]),.dout(n15531),.clk(gclk));
	jnot g15240(.din(w_n14973_0[0]),.dout(n15532),.clk(gclk));
	jnot g15241(.din(w_n14974_0[0]),.dout(n15533),.clk(gclk));
	jand g15242(.dina(w_asqrt10_25[1]),.dinb(w_n14970_0[0]),.dout(n15534),.clk(gclk));
	jand g15243(.dina(w_n15534_0[1]),.dinb(n15533),.dout(n15535),.clk(gclk));
	jor g15244(.dina(n15535),.dinb(n15532),.dout(n15536),.clk(gclk));
	jnot g15245(.din(w_n14975_0[0]),.dout(n15537),.clk(gclk));
	jand g15246(.dina(w_n15534_0[0]),.dinb(n15537),.dout(n15538),.clk(gclk));
	jnot g15247(.din(n15538),.dout(n15539),.clk(gclk));
	jand g15248(.dina(n15539),.dinb(n15536),.dout(n15540),.clk(gclk));
	jand g15249(.dina(w_n15540_0[1]),.dinb(n15531),.dout(n15541),.clk(gclk));
	jor g15250(.dina(w_n15541_0[1]),.dinb(w_n15530_0[1]),.dout(n15542),.clk(gclk));
	jand g15251(.dina(n15542),.dinb(w_asqrt28_13[1]),.dout(n15543),.clk(gclk));
	jor g15252(.dina(w_n15530_0[0]),.dinb(w_asqrt28_13[0]),.dout(n15544),.clk(gclk));
	jor g15253(.dina(n15544),.dinb(w_n15541_0[0]),.dout(n15545),.clk(gclk));
	jnot g15254(.din(w_n14981_0[0]),.dout(n15546),.clk(gclk));
	jnot g15255(.din(w_n14983_0[0]),.dout(n15547),.clk(gclk));
	jand g15256(.dina(w_asqrt10_25[0]),.dinb(w_n14977_0[0]),.dout(n15548),.clk(gclk));
	jand g15257(.dina(w_n15548_0[1]),.dinb(n15547),.dout(n15549),.clk(gclk));
	jor g15258(.dina(n15549),.dinb(n15546),.dout(n15550),.clk(gclk));
	jnot g15259(.din(w_n14984_0[0]),.dout(n15551),.clk(gclk));
	jand g15260(.dina(w_n15548_0[0]),.dinb(n15551),.dout(n15552),.clk(gclk));
	jnot g15261(.din(n15552),.dout(n15553),.clk(gclk));
	jand g15262(.dina(n15553),.dinb(n15550),.dout(n15554),.clk(gclk));
	jand g15263(.dina(w_n15554_0[1]),.dinb(w_n15545_0[1]),.dout(n15555),.clk(gclk));
	jor g15264(.dina(n15555),.dinb(w_n15543_0[1]),.dout(n15556),.clk(gclk));
	jand g15265(.dina(w_n15556_0[1]),.dinb(w_asqrt29_10[0]),.dout(n15557),.clk(gclk));
	jxor g15266(.dina(w_n14985_0[0]),.dinb(w_n7260_10[0]),.dout(n15558),.clk(gclk));
	jand g15267(.dina(n15558),.dinb(w_asqrt10_24[2]),.dout(n15559),.clk(gclk));
	jxor g15268(.dina(n15559),.dinb(w_n14995_0[0]),.dout(n15560),.clk(gclk));
	jnot g15269(.din(n15560),.dout(n15561),.clk(gclk));
	jor g15270(.dina(w_n15556_0[0]),.dinb(w_asqrt29_9[2]),.dout(n15562),.clk(gclk));
	jand g15271(.dina(w_n15562_0[1]),.dinb(w_n15561_0[1]),.dout(n15563),.clk(gclk));
	jor g15272(.dina(w_n15563_0[2]),.dinb(w_n15557_0[2]),.dout(n15564),.clk(gclk));
	jand g15273(.dina(n15564),.dinb(w_asqrt30_13[1]),.dout(n15565),.clk(gclk));
	jnot g15274(.din(w_n15000_0[0]),.dout(n15566),.clk(gclk));
	jand g15275(.dina(n15566),.dinb(w_n14998_0[0]),.dout(n15567),.clk(gclk));
	jand g15276(.dina(n15567),.dinb(w_asqrt10_24[1]),.dout(n15568),.clk(gclk));
	jxor g15277(.dina(n15568),.dinb(w_n15008_0[0]),.dout(n15569),.clk(gclk));
	jnot g15278(.din(n15569),.dout(n15570),.clk(gclk));
	jor g15279(.dina(w_n15557_0[1]),.dinb(w_asqrt30_13[0]),.dout(n15571),.clk(gclk));
	jor g15280(.dina(n15571),.dinb(w_n15563_0[1]),.dout(n15572),.clk(gclk));
	jand g15281(.dina(w_n15572_0[1]),.dinb(w_n15570_0[1]),.dout(n15573),.clk(gclk));
	jor g15282(.dina(w_n15573_0[1]),.dinb(w_n15565_0[1]),.dout(n15574),.clk(gclk));
	jand g15283(.dina(w_n15574_0[2]),.dinb(w_asqrt31_10[0]),.dout(n15575),.clk(gclk));
	jor g15284(.dina(w_n15574_0[1]),.dinb(w_asqrt31_9[2]),.dout(n15576),.clk(gclk));
	jnot g15285(.din(w_n15014_0[0]),.dout(n15577),.clk(gclk));
	jnot g15286(.din(w_n15015_0[0]),.dout(n15578),.clk(gclk));
	jand g15287(.dina(w_asqrt10_24[0]),.dinb(w_n15011_0[0]),.dout(n15579),.clk(gclk));
	jand g15288(.dina(w_n15579_0[1]),.dinb(n15578),.dout(n15580),.clk(gclk));
	jor g15289(.dina(n15580),.dinb(n15577),.dout(n15581),.clk(gclk));
	jnot g15290(.din(w_n15016_0[0]),.dout(n15582),.clk(gclk));
	jand g15291(.dina(w_n15579_0[0]),.dinb(n15582),.dout(n15583),.clk(gclk));
	jnot g15292(.din(n15583),.dout(n15584),.clk(gclk));
	jand g15293(.dina(n15584),.dinb(n15581),.dout(n15585),.clk(gclk));
	jand g15294(.dina(w_n15585_0[1]),.dinb(n15576),.dout(n15586),.clk(gclk));
	jor g15295(.dina(w_n15586_0[1]),.dinb(w_n15575_0[1]),.dout(n15587),.clk(gclk));
	jand g15296(.dina(n15587),.dinb(w_asqrt32_13[1]),.dout(n15588),.clk(gclk));
	jor g15297(.dina(w_n15575_0[0]),.dinb(w_asqrt32_13[0]),.dout(n15589),.clk(gclk));
	jor g15298(.dina(n15589),.dinb(w_n15586_0[0]),.dout(n15590),.clk(gclk));
	jnot g15299(.din(w_n15022_0[0]),.dout(n15591),.clk(gclk));
	jnot g15300(.din(w_n15024_0[0]),.dout(n15592),.clk(gclk));
	jand g15301(.dina(w_asqrt10_23[2]),.dinb(w_n15018_0[0]),.dout(n15593),.clk(gclk));
	jand g15302(.dina(w_n15593_0[1]),.dinb(n15592),.dout(n15594),.clk(gclk));
	jor g15303(.dina(n15594),.dinb(n15591),.dout(n15595),.clk(gclk));
	jnot g15304(.din(w_n15025_0[0]),.dout(n15596),.clk(gclk));
	jand g15305(.dina(w_n15593_0[0]),.dinb(n15596),.dout(n15597),.clk(gclk));
	jnot g15306(.din(n15597),.dout(n15598),.clk(gclk));
	jand g15307(.dina(n15598),.dinb(n15595),.dout(n15599),.clk(gclk));
	jand g15308(.dina(w_n15599_0[1]),.dinb(w_n15590_0[1]),.dout(n15600),.clk(gclk));
	jor g15309(.dina(n15600),.dinb(w_n15588_0[1]),.dout(n15601),.clk(gclk));
	jand g15310(.dina(w_n15601_0[1]),.dinb(w_asqrt33_10[1]),.dout(n15602),.clk(gclk));
	jxor g15311(.dina(w_n15026_0[0]),.dinb(w_n5788_10[2]),.dout(n15603),.clk(gclk));
	jand g15312(.dina(n15603),.dinb(w_asqrt10_23[1]),.dout(n15604),.clk(gclk));
	jxor g15313(.dina(n15604),.dinb(w_n15036_0[0]),.dout(n15605),.clk(gclk));
	jnot g15314(.din(n15605),.dout(n15606),.clk(gclk));
	jor g15315(.dina(w_n15601_0[0]),.dinb(w_asqrt33_10[0]),.dout(n15607),.clk(gclk));
	jand g15316(.dina(w_n15607_0[1]),.dinb(w_n15606_0[1]),.dout(n15608),.clk(gclk));
	jor g15317(.dina(w_n15608_0[2]),.dinb(w_n15602_0[2]),.dout(n15609),.clk(gclk));
	jand g15318(.dina(n15609),.dinb(w_asqrt34_13[1]),.dout(n15610),.clk(gclk));
	jnot g15319(.din(w_n15041_0[0]),.dout(n15611),.clk(gclk));
	jand g15320(.dina(n15611),.dinb(w_n15039_0[0]),.dout(n15612),.clk(gclk));
	jand g15321(.dina(n15612),.dinb(w_asqrt10_23[0]),.dout(n15613),.clk(gclk));
	jxor g15322(.dina(n15613),.dinb(w_n15049_0[0]),.dout(n15614),.clk(gclk));
	jnot g15323(.din(n15614),.dout(n15615),.clk(gclk));
	jor g15324(.dina(w_n15602_0[1]),.dinb(w_asqrt34_13[0]),.dout(n15616),.clk(gclk));
	jor g15325(.dina(n15616),.dinb(w_n15608_0[1]),.dout(n15617),.clk(gclk));
	jand g15326(.dina(w_n15617_0[1]),.dinb(w_n15615_0[1]),.dout(n15618),.clk(gclk));
	jor g15327(.dina(w_n15618_0[1]),.dinb(w_n15610_0[1]),.dout(n15619),.clk(gclk));
	jand g15328(.dina(w_n15619_0[2]),.dinb(w_asqrt35_10[1]),.dout(n15620),.clk(gclk));
	jor g15329(.dina(w_n15619_0[1]),.dinb(w_asqrt35_10[0]),.dout(n15621),.clk(gclk));
	jnot g15330(.din(w_n15055_0[0]),.dout(n15622),.clk(gclk));
	jnot g15331(.din(w_n15056_0[0]),.dout(n15623),.clk(gclk));
	jand g15332(.dina(w_asqrt10_22[2]),.dinb(w_n15052_0[0]),.dout(n15624),.clk(gclk));
	jand g15333(.dina(w_n15624_0[1]),.dinb(n15623),.dout(n15625),.clk(gclk));
	jor g15334(.dina(n15625),.dinb(n15622),.dout(n15626),.clk(gclk));
	jnot g15335(.din(w_n15057_0[0]),.dout(n15627),.clk(gclk));
	jand g15336(.dina(w_n15624_0[0]),.dinb(n15627),.dout(n15628),.clk(gclk));
	jnot g15337(.din(n15628),.dout(n15629),.clk(gclk));
	jand g15338(.dina(n15629),.dinb(n15626),.dout(n15630),.clk(gclk));
	jand g15339(.dina(w_n15630_0[1]),.dinb(n15621),.dout(n15631),.clk(gclk));
	jor g15340(.dina(w_n15631_0[1]),.dinb(w_n15620_0[1]),.dout(n15632),.clk(gclk));
	jand g15341(.dina(n15632),.dinb(w_asqrt36_13[1]),.dout(n15633),.clk(gclk));
	jor g15342(.dina(w_n15620_0[0]),.dinb(w_asqrt36_13[0]),.dout(n15634),.clk(gclk));
	jor g15343(.dina(n15634),.dinb(w_n15631_0[0]),.dout(n15635),.clk(gclk));
	jnot g15344(.din(w_n15063_0[0]),.dout(n15636),.clk(gclk));
	jnot g15345(.din(w_n15065_0[0]),.dout(n15637),.clk(gclk));
	jand g15346(.dina(w_asqrt10_22[1]),.dinb(w_n15059_0[0]),.dout(n15638),.clk(gclk));
	jand g15347(.dina(w_n15638_0[1]),.dinb(n15637),.dout(n15639),.clk(gclk));
	jor g15348(.dina(n15639),.dinb(n15636),.dout(n15640),.clk(gclk));
	jnot g15349(.din(w_n15066_0[0]),.dout(n15641),.clk(gclk));
	jand g15350(.dina(w_n15638_0[0]),.dinb(n15641),.dout(n15642),.clk(gclk));
	jnot g15351(.din(n15642),.dout(n15643),.clk(gclk));
	jand g15352(.dina(n15643),.dinb(n15640),.dout(n15644),.clk(gclk));
	jand g15353(.dina(w_n15644_0[1]),.dinb(w_n15635_0[1]),.dout(n15645),.clk(gclk));
	jor g15354(.dina(n15645),.dinb(w_n15633_0[1]),.dout(n15646),.clk(gclk));
	jand g15355(.dina(w_n15646_0[1]),.dinb(w_asqrt37_10[2]),.dout(n15647),.clk(gclk));
	jxor g15356(.dina(w_n15067_0[0]),.dinb(w_n4494_11[2]),.dout(n15648),.clk(gclk));
	jand g15357(.dina(n15648),.dinb(w_asqrt10_22[0]),.dout(n15649),.clk(gclk));
	jxor g15358(.dina(n15649),.dinb(w_n15077_0[0]),.dout(n15650),.clk(gclk));
	jnot g15359(.din(n15650),.dout(n15651),.clk(gclk));
	jor g15360(.dina(w_n15646_0[0]),.dinb(w_asqrt37_10[1]),.dout(n15652),.clk(gclk));
	jand g15361(.dina(w_n15652_0[1]),.dinb(w_n15651_0[1]),.dout(n15653),.clk(gclk));
	jor g15362(.dina(w_n15653_0[2]),.dinb(w_n15647_0[2]),.dout(n15654),.clk(gclk));
	jand g15363(.dina(n15654),.dinb(w_asqrt38_13[1]),.dout(n15655),.clk(gclk));
	jnot g15364(.din(w_n15082_0[0]),.dout(n15656),.clk(gclk));
	jand g15365(.dina(n15656),.dinb(w_n15080_0[0]),.dout(n15657),.clk(gclk));
	jand g15366(.dina(n15657),.dinb(w_asqrt10_21[2]),.dout(n15658),.clk(gclk));
	jxor g15367(.dina(n15658),.dinb(w_n15090_0[0]),.dout(n15659),.clk(gclk));
	jnot g15368(.din(n15659),.dout(n15660),.clk(gclk));
	jor g15369(.dina(w_n15647_0[1]),.dinb(w_asqrt38_13[0]),.dout(n15661),.clk(gclk));
	jor g15370(.dina(n15661),.dinb(w_n15653_0[1]),.dout(n15662),.clk(gclk));
	jand g15371(.dina(w_n15662_0[1]),.dinb(w_n15660_0[1]),.dout(n15663),.clk(gclk));
	jor g15372(.dina(w_n15663_0[1]),.dinb(w_n15655_0[1]),.dout(n15664),.clk(gclk));
	jand g15373(.dina(w_n15664_0[2]),.dinb(w_asqrt39_10[2]),.dout(n15665),.clk(gclk));
	jor g15374(.dina(w_n15664_0[1]),.dinb(w_asqrt39_10[1]),.dout(n15666),.clk(gclk));
	jnot g15375(.din(w_n15096_0[0]),.dout(n15667),.clk(gclk));
	jnot g15376(.din(w_n15097_0[0]),.dout(n15668),.clk(gclk));
	jand g15377(.dina(w_asqrt10_21[1]),.dinb(w_n15093_0[0]),.dout(n15669),.clk(gclk));
	jand g15378(.dina(w_n15669_0[1]),.dinb(n15668),.dout(n15670),.clk(gclk));
	jor g15379(.dina(n15670),.dinb(n15667),.dout(n15671),.clk(gclk));
	jnot g15380(.din(w_n15098_0[0]),.dout(n15672),.clk(gclk));
	jand g15381(.dina(w_n15669_0[0]),.dinb(n15672),.dout(n15673),.clk(gclk));
	jnot g15382(.din(n15673),.dout(n15674),.clk(gclk));
	jand g15383(.dina(n15674),.dinb(n15671),.dout(n15675),.clk(gclk));
	jand g15384(.dina(w_n15675_0[1]),.dinb(n15666),.dout(n15676),.clk(gclk));
	jor g15385(.dina(w_n15676_0[1]),.dinb(w_n15665_0[1]),.dout(n15677),.clk(gclk));
	jand g15386(.dina(n15677),.dinb(w_asqrt40_13[1]),.dout(n15678),.clk(gclk));
	jor g15387(.dina(w_n15665_0[0]),.dinb(w_asqrt40_13[0]),.dout(n15679),.clk(gclk));
	jor g15388(.dina(n15679),.dinb(w_n15676_0[0]),.dout(n15680),.clk(gclk));
	jnot g15389(.din(w_n15104_0[0]),.dout(n15681),.clk(gclk));
	jnot g15390(.din(w_n15106_0[0]),.dout(n15682),.clk(gclk));
	jand g15391(.dina(w_asqrt10_21[0]),.dinb(w_n15100_0[0]),.dout(n15683),.clk(gclk));
	jand g15392(.dina(w_n15683_0[1]),.dinb(n15682),.dout(n15684),.clk(gclk));
	jor g15393(.dina(n15684),.dinb(n15681),.dout(n15685),.clk(gclk));
	jnot g15394(.din(w_n15107_0[0]),.dout(n15686),.clk(gclk));
	jand g15395(.dina(w_n15683_0[0]),.dinb(n15686),.dout(n15687),.clk(gclk));
	jnot g15396(.din(n15687),.dout(n15688),.clk(gclk));
	jand g15397(.dina(n15688),.dinb(n15685),.dout(n15689),.clk(gclk));
	jand g15398(.dina(w_n15689_0[1]),.dinb(w_n15680_0[1]),.dout(n15690),.clk(gclk));
	jor g15399(.dina(n15690),.dinb(w_n15678_0[1]),.dout(n15691),.clk(gclk));
	jand g15400(.dina(w_n15691_0[1]),.dinb(w_asqrt41_11[0]),.dout(n15692),.clk(gclk));
	jxor g15401(.dina(w_n15108_0[0]),.dinb(w_n3371_12[1]),.dout(n15693),.clk(gclk));
	jand g15402(.dina(n15693),.dinb(w_asqrt10_20[2]),.dout(n15694),.clk(gclk));
	jxor g15403(.dina(n15694),.dinb(w_n15118_0[0]),.dout(n15695),.clk(gclk));
	jnot g15404(.din(n15695),.dout(n15696),.clk(gclk));
	jor g15405(.dina(w_n15691_0[0]),.dinb(w_asqrt41_10[2]),.dout(n15697),.clk(gclk));
	jand g15406(.dina(w_n15697_0[1]),.dinb(w_n15696_0[1]),.dout(n15698),.clk(gclk));
	jor g15407(.dina(w_n15698_0[2]),.dinb(w_n15692_0[2]),.dout(n15699),.clk(gclk));
	jand g15408(.dina(n15699),.dinb(w_asqrt42_13[1]),.dout(n15700),.clk(gclk));
	jnot g15409(.din(w_n15123_0[0]),.dout(n15701),.clk(gclk));
	jand g15410(.dina(n15701),.dinb(w_n15121_0[0]),.dout(n15702),.clk(gclk));
	jand g15411(.dina(n15702),.dinb(w_asqrt10_20[1]),.dout(n15703),.clk(gclk));
	jxor g15412(.dina(n15703),.dinb(w_n15131_0[0]),.dout(n15704),.clk(gclk));
	jnot g15413(.din(n15704),.dout(n15705),.clk(gclk));
	jor g15414(.dina(w_n15692_0[1]),.dinb(w_asqrt42_13[0]),.dout(n15706),.clk(gclk));
	jor g15415(.dina(n15706),.dinb(w_n15698_0[1]),.dout(n15707),.clk(gclk));
	jand g15416(.dina(w_n15707_0[1]),.dinb(w_n15705_0[1]),.dout(n15708),.clk(gclk));
	jor g15417(.dina(w_n15708_0[1]),.dinb(w_n15700_0[1]),.dout(n15709),.clk(gclk));
	jand g15418(.dina(w_n15709_0[2]),.dinb(w_asqrt43_11[0]),.dout(n15710),.clk(gclk));
	jor g15419(.dina(w_n15709_0[1]),.dinb(w_asqrt43_10[2]),.dout(n15711),.clk(gclk));
	jnot g15420(.din(w_n15137_0[0]),.dout(n15712),.clk(gclk));
	jnot g15421(.din(w_n15138_0[0]),.dout(n15713),.clk(gclk));
	jand g15422(.dina(w_asqrt10_20[0]),.dinb(w_n15134_0[0]),.dout(n15714),.clk(gclk));
	jand g15423(.dina(w_n15714_0[1]),.dinb(n15713),.dout(n15715),.clk(gclk));
	jor g15424(.dina(n15715),.dinb(n15712),.dout(n15716),.clk(gclk));
	jnot g15425(.din(w_n15139_0[0]),.dout(n15717),.clk(gclk));
	jand g15426(.dina(w_n15714_0[0]),.dinb(n15717),.dout(n15718),.clk(gclk));
	jnot g15427(.din(n15718),.dout(n15719),.clk(gclk));
	jand g15428(.dina(n15719),.dinb(n15716),.dout(n15720),.clk(gclk));
	jand g15429(.dina(w_n15720_0[1]),.dinb(n15711),.dout(n15721),.clk(gclk));
	jor g15430(.dina(w_n15721_0[1]),.dinb(w_n15710_0[1]),.dout(n15722),.clk(gclk));
	jand g15431(.dina(n15722),.dinb(w_asqrt44_13[1]),.dout(n15723),.clk(gclk));
	jor g15432(.dina(w_n15710_0[0]),.dinb(w_asqrt44_13[0]),.dout(n15724),.clk(gclk));
	jor g15433(.dina(n15724),.dinb(w_n15721_0[0]),.dout(n15725),.clk(gclk));
	jnot g15434(.din(w_n15145_0[0]),.dout(n15726),.clk(gclk));
	jnot g15435(.din(w_n15147_0[0]),.dout(n15727),.clk(gclk));
	jand g15436(.dina(w_asqrt10_19[2]),.dinb(w_n15141_0[0]),.dout(n15728),.clk(gclk));
	jand g15437(.dina(w_n15728_0[1]),.dinb(n15727),.dout(n15729),.clk(gclk));
	jor g15438(.dina(n15729),.dinb(n15726),.dout(n15730),.clk(gclk));
	jnot g15439(.din(w_n15148_0[0]),.dout(n15731),.clk(gclk));
	jand g15440(.dina(w_n15728_0[0]),.dinb(n15731),.dout(n15732),.clk(gclk));
	jnot g15441(.din(n15732),.dout(n15733),.clk(gclk));
	jand g15442(.dina(n15733),.dinb(n15730),.dout(n15734),.clk(gclk));
	jand g15443(.dina(w_n15734_0[1]),.dinb(w_n15725_0[1]),.dout(n15735),.clk(gclk));
	jor g15444(.dina(n15735),.dinb(w_n15723_0[1]),.dout(n15736),.clk(gclk));
	jand g15445(.dina(w_n15736_0[1]),.dinb(w_asqrt45_11[1]),.dout(n15737),.clk(gclk));
	jxor g15446(.dina(w_n15149_0[0]),.dinb(w_n2420_13[1]),.dout(n15738),.clk(gclk));
	jand g15447(.dina(n15738),.dinb(w_asqrt10_19[1]),.dout(n15739),.clk(gclk));
	jxor g15448(.dina(n15739),.dinb(w_n15159_0[0]),.dout(n15740),.clk(gclk));
	jnot g15449(.din(n15740),.dout(n15741),.clk(gclk));
	jor g15450(.dina(w_n15736_0[0]),.dinb(w_asqrt45_11[0]),.dout(n15742),.clk(gclk));
	jand g15451(.dina(w_n15742_0[1]),.dinb(w_n15741_0[1]),.dout(n15743),.clk(gclk));
	jor g15452(.dina(w_n15743_0[2]),.dinb(w_n15737_0[2]),.dout(n15744),.clk(gclk));
	jand g15453(.dina(n15744),.dinb(w_asqrt46_13[1]),.dout(n15745),.clk(gclk));
	jnot g15454(.din(w_n15164_0[0]),.dout(n15746),.clk(gclk));
	jand g15455(.dina(n15746),.dinb(w_n15162_0[0]),.dout(n15747),.clk(gclk));
	jand g15456(.dina(n15747),.dinb(w_asqrt10_19[0]),.dout(n15748),.clk(gclk));
	jxor g15457(.dina(n15748),.dinb(w_n15172_0[0]),.dout(n15749),.clk(gclk));
	jnot g15458(.din(n15749),.dout(n15750),.clk(gclk));
	jor g15459(.dina(w_n15737_0[1]),.dinb(w_asqrt46_13[0]),.dout(n15751),.clk(gclk));
	jor g15460(.dina(n15751),.dinb(w_n15743_0[1]),.dout(n15752),.clk(gclk));
	jand g15461(.dina(w_n15752_0[1]),.dinb(w_n15750_0[1]),.dout(n15753),.clk(gclk));
	jor g15462(.dina(w_n15753_0[1]),.dinb(w_n15745_0[1]),.dout(n15754),.clk(gclk));
	jand g15463(.dina(w_n15754_0[2]),.dinb(w_asqrt47_11[1]),.dout(n15755),.clk(gclk));
	jor g15464(.dina(w_n15754_0[1]),.dinb(w_asqrt47_11[0]),.dout(n15756),.clk(gclk));
	jnot g15465(.din(w_n15178_0[0]),.dout(n15757),.clk(gclk));
	jnot g15466(.din(w_n15179_0[0]),.dout(n15758),.clk(gclk));
	jand g15467(.dina(w_asqrt10_18[2]),.dinb(w_n15175_0[0]),.dout(n15759),.clk(gclk));
	jand g15468(.dina(w_n15759_0[1]),.dinb(n15758),.dout(n15760),.clk(gclk));
	jor g15469(.dina(n15760),.dinb(n15757),.dout(n15761),.clk(gclk));
	jnot g15470(.din(w_n15180_0[0]),.dout(n15762),.clk(gclk));
	jand g15471(.dina(w_n15759_0[0]),.dinb(n15762),.dout(n15763),.clk(gclk));
	jnot g15472(.din(n15763),.dout(n15764),.clk(gclk));
	jand g15473(.dina(n15764),.dinb(n15761),.dout(n15765),.clk(gclk));
	jand g15474(.dina(w_n15765_0[1]),.dinb(n15756),.dout(n15766),.clk(gclk));
	jor g15475(.dina(w_n15766_0[1]),.dinb(w_n15755_0[1]),.dout(n15767),.clk(gclk));
	jand g15476(.dina(n15767),.dinb(w_asqrt48_13[1]),.dout(n15768),.clk(gclk));
	jor g15477(.dina(w_n15755_0[0]),.dinb(w_asqrt48_13[0]),.dout(n15769),.clk(gclk));
	jor g15478(.dina(n15769),.dinb(w_n15766_0[0]),.dout(n15770),.clk(gclk));
	jnot g15479(.din(w_n15186_0[0]),.dout(n15771),.clk(gclk));
	jnot g15480(.din(w_n15188_0[0]),.dout(n15772),.clk(gclk));
	jand g15481(.dina(w_asqrt10_18[1]),.dinb(w_n15182_0[0]),.dout(n15773),.clk(gclk));
	jand g15482(.dina(w_n15773_0[1]),.dinb(n15772),.dout(n15774),.clk(gclk));
	jor g15483(.dina(n15774),.dinb(n15771),.dout(n15775),.clk(gclk));
	jnot g15484(.din(w_n15189_0[0]),.dout(n15776),.clk(gclk));
	jand g15485(.dina(w_n15773_0[0]),.dinb(n15776),.dout(n15777),.clk(gclk));
	jnot g15486(.din(n15777),.dout(n15778),.clk(gclk));
	jand g15487(.dina(n15778),.dinb(n15775),.dout(n15779),.clk(gclk));
	jand g15488(.dina(w_n15779_0[1]),.dinb(w_n15770_0[1]),.dout(n15780),.clk(gclk));
	jor g15489(.dina(n15780),.dinb(w_n15768_0[1]),.dout(n15781),.clk(gclk));
	jand g15490(.dina(w_n15781_0[1]),.dinb(w_asqrt49_11[2]),.dout(n15782),.clk(gclk));
	jxor g15491(.dina(w_n15190_0[0]),.dinb(w_n1641_14[0]),.dout(n15783),.clk(gclk));
	jand g15492(.dina(n15783),.dinb(w_asqrt10_18[0]),.dout(n15784),.clk(gclk));
	jxor g15493(.dina(n15784),.dinb(w_n15200_0[0]),.dout(n15785),.clk(gclk));
	jnot g15494(.din(n15785),.dout(n15786),.clk(gclk));
	jor g15495(.dina(w_n15781_0[0]),.dinb(w_asqrt49_11[1]),.dout(n15787),.clk(gclk));
	jand g15496(.dina(w_n15787_0[1]),.dinb(w_n15786_0[1]),.dout(n15788),.clk(gclk));
	jor g15497(.dina(w_n15788_0[2]),.dinb(w_n15782_0[2]),.dout(n15789),.clk(gclk));
	jand g15498(.dina(n15789),.dinb(w_asqrt50_13[1]),.dout(n15790),.clk(gclk));
	jnot g15499(.din(w_n15205_0[0]),.dout(n15791),.clk(gclk));
	jand g15500(.dina(n15791),.dinb(w_n15203_0[0]),.dout(n15792),.clk(gclk));
	jand g15501(.dina(n15792),.dinb(w_asqrt10_17[2]),.dout(n15793),.clk(gclk));
	jxor g15502(.dina(n15793),.dinb(w_n15213_0[0]),.dout(n15794),.clk(gclk));
	jnot g15503(.din(n15794),.dout(n15795),.clk(gclk));
	jor g15504(.dina(w_n15782_0[1]),.dinb(w_asqrt50_13[0]),.dout(n15796),.clk(gclk));
	jor g15505(.dina(n15796),.dinb(w_n15788_0[1]),.dout(n15797),.clk(gclk));
	jand g15506(.dina(w_n15797_0[1]),.dinb(w_n15795_0[1]),.dout(n15798),.clk(gclk));
	jor g15507(.dina(w_n15798_0[1]),.dinb(w_n15790_0[1]),.dout(n15799),.clk(gclk));
	jand g15508(.dina(w_n15799_0[2]),.dinb(w_asqrt51_11[2]),.dout(n15800),.clk(gclk));
	jor g15509(.dina(w_n15799_0[1]),.dinb(w_asqrt51_11[1]),.dout(n15801),.clk(gclk));
	jnot g15510(.din(w_n15219_0[0]),.dout(n15802),.clk(gclk));
	jnot g15511(.din(w_n15220_0[0]),.dout(n15803),.clk(gclk));
	jand g15512(.dina(w_asqrt10_17[1]),.dinb(w_n15216_0[0]),.dout(n15804),.clk(gclk));
	jand g15513(.dina(w_n15804_0[1]),.dinb(n15803),.dout(n15805),.clk(gclk));
	jor g15514(.dina(n15805),.dinb(n15802),.dout(n15806),.clk(gclk));
	jnot g15515(.din(w_n15221_0[0]),.dout(n15807),.clk(gclk));
	jand g15516(.dina(w_n15804_0[0]),.dinb(n15807),.dout(n15808),.clk(gclk));
	jnot g15517(.din(n15808),.dout(n15809),.clk(gclk));
	jand g15518(.dina(n15809),.dinb(n15806),.dout(n15810),.clk(gclk));
	jand g15519(.dina(w_n15810_0[1]),.dinb(n15801),.dout(n15811),.clk(gclk));
	jor g15520(.dina(w_n15811_0[1]),.dinb(w_n15800_0[1]),.dout(n15812),.clk(gclk));
	jand g15521(.dina(n15812),.dinb(w_asqrt52_13[1]),.dout(n15813),.clk(gclk));
	jnot g15522(.din(w_n15225_0[0]),.dout(n15814),.clk(gclk));
	jand g15523(.dina(n15814),.dinb(w_n15223_0[0]),.dout(n15815),.clk(gclk));
	jand g15524(.dina(n15815),.dinb(w_asqrt10_17[0]),.dout(n15816),.clk(gclk));
	jxor g15525(.dina(n15816),.dinb(w_n15233_0[0]),.dout(n15817),.clk(gclk));
	jnot g15526(.din(n15817),.dout(n15818),.clk(gclk));
	jor g15527(.dina(w_n15800_0[0]),.dinb(w_asqrt52_13[0]),.dout(n15819),.clk(gclk));
	jor g15528(.dina(n15819),.dinb(w_n15811_0[0]),.dout(n15820),.clk(gclk));
	jand g15529(.dina(w_n15820_0[1]),.dinb(w_n15818_0[1]),.dout(n15821),.clk(gclk));
	jor g15530(.dina(w_n15821_0[1]),.dinb(w_n15813_0[1]),.dout(n15822),.clk(gclk));
	jand g15531(.dina(w_n15822_0[2]),.dinb(w_asqrt53_12[0]),.dout(n15823),.clk(gclk));
	jor g15532(.dina(w_n15822_0[1]),.dinb(w_asqrt53_11[2]),.dout(n15824),.clk(gclk));
	jand g15533(.dina(n15824),.dinb(w_n15361_0[0]),.dout(n15825),.clk(gclk));
	jor g15534(.dina(w_n15825_0[1]),.dinb(w_n15823_0[1]),.dout(n15826),.clk(gclk));
	jand g15535(.dina(n15826),.dinb(w_asqrt54_13[1]),.dout(n15827),.clk(gclk));
	jor g15536(.dina(w_n15823_0[0]),.dinb(w_asqrt54_13[0]),.dout(n15828),.clk(gclk));
	jor g15537(.dina(n15828),.dinb(w_n15825_0[0]),.dout(n15829),.clk(gclk));
	jnot g15538(.din(w_n15245_0[0]),.dout(n15830),.clk(gclk));
	jnot g15539(.din(w_n15247_0[0]),.dout(n15831),.clk(gclk));
	jand g15540(.dina(w_asqrt10_16[2]),.dinb(w_n15241_0[0]),.dout(n15832),.clk(gclk));
	jand g15541(.dina(w_n15832_0[1]),.dinb(n15831),.dout(n15833),.clk(gclk));
	jor g15542(.dina(n15833),.dinb(n15830),.dout(n15834),.clk(gclk));
	jnot g15543(.din(w_n15248_0[0]),.dout(n15835),.clk(gclk));
	jand g15544(.dina(w_n15832_0[0]),.dinb(n15835),.dout(n15836),.clk(gclk));
	jnot g15545(.din(n15836),.dout(n15837),.clk(gclk));
	jand g15546(.dina(n15837),.dinb(n15834),.dout(n15838),.clk(gclk));
	jand g15547(.dina(w_n15838_0[1]),.dinb(w_n15829_0[1]),.dout(n15839),.clk(gclk));
	jor g15548(.dina(n15839),.dinb(w_n15827_0[1]),.dout(n15840),.clk(gclk));
	jand g15549(.dina(w_n15840_0[2]),.dinb(w_asqrt55_12[1]),.dout(n15841),.clk(gclk));
	jor g15550(.dina(w_n15840_0[1]),.dinb(w_asqrt55_12[0]),.dout(n15842),.clk(gclk));
	jnot g15551(.din(w_n15253_0[0]),.dout(n15843),.clk(gclk));
	jnot g15552(.din(w_n15254_0[0]),.dout(n15844),.clk(gclk));
	jand g15553(.dina(w_asqrt10_16[1]),.dinb(w_n15250_0[0]),.dout(n15845),.clk(gclk));
	jand g15554(.dina(w_n15845_0[1]),.dinb(n15844),.dout(n15846),.clk(gclk));
	jor g15555(.dina(n15846),.dinb(n15843),.dout(n15847),.clk(gclk));
	jnot g15556(.din(w_n15255_0[0]),.dout(n15848),.clk(gclk));
	jand g15557(.dina(w_n15845_0[0]),.dinb(n15848),.dout(n15849),.clk(gclk));
	jnot g15558(.din(n15849),.dout(n15850),.clk(gclk));
	jand g15559(.dina(n15850),.dinb(n15847),.dout(n15851),.clk(gclk));
	jand g15560(.dina(w_n15851_0[1]),.dinb(n15842),.dout(n15852),.clk(gclk));
	jor g15561(.dina(w_n15852_0[1]),.dinb(w_n15841_0[1]),.dout(n15853),.clk(gclk));
	jand g15562(.dina(n15853),.dinb(w_asqrt56_13[1]),.dout(n15854),.clk(gclk));
	jor g15563(.dina(w_n15841_0[0]),.dinb(w_asqrt56_13[0]),.dout(n15855),.clk(gclk));
	jor g15564(.dina(n15855),.dinb(w_n15852_0[0]),.dout(n15856),.clk(gclk));
	jnot g15565(.din(w_n15261_0[0]),.dout(n15857),.clk(gclk));
	jnot g15566(.din(w_n15263_0[0]),.dout(n15858),.clk(gclk));
	jand g15567(.dina(w_asqrt10_16[0]),.dinb(w_n15257_0[0]),.dout(n15859),.clk(gclk));
	jand g15568(.dina(w_n15859_0[1]),.dinb(n15858),.dout(n15860),.clk(gclk));
	jor g15569(.dina(n15860),.dinb(n15857),.dout(n15861),.clk(gclk));
	jnot g15570(.din(w_n15264_0[0]),.dout(n15862),.clk(gclk));
	jand g15571(.dina(w_n15859_0[0]),.dinb(n15862),.dout(n15863),.clk(gclk));
	jnot g15572(.din(n15863),.dout(n15864),.clk(gclk));
	jand g15573(.dina(n15864),.dinb(n15861),.dout(n15865),.clk(gclk));
	jand g15574(.dina(w_n15865_0[1]),.dinb(w_n15856_0[1]),.dout(n15866),.clk(gclk));
	jor g15575(.dina(n15866),.dinb(w_n15854_0[1]),.dout(n15867),.clk(gclk));
	jand g15576(.dina(w_n15867_0[1]),.dinb(w_asqrt57_12[2]),.dout(n15868),.clk(gclk));
	jxor g15577(.dina(w_n15265_0[0]),.dinb(w_n590_15[2]),.dout(n15869),.clk(gclk));
	jand g15578(.dina(n15869),.dinb(w_asqrt10_15[2]),.dout(n15870),.clk(gclk));
	jxor g15579(.dina(n15870),.dinb(w_n15275_0[0]),.dout(n15871),.clk(gclk));
	jnot g15580(.din(n15871),.dout(n15872),.clk(gclk));
	jor g15581(.dina(w_n15867_0[0]),.dinb(w_asqrt57_12[1]),.dout(n15873),.clk(gclk));
	jand g15582(.dina(w_n15873_0[1]),.dinb(w_n15872_0[1]),.dout(n15874),.clk(gclk));
	jor g15583(.dina(w_n15874_0[2]),.dinb(w_n15868_0[2]),.dout(n15875),.clk(gclk));
	jand g15584(.dina(n15875),.dinb(w_asqrt58_13[1]),.dout(n15876),.clk(gclk));
	jnot g15585(.din(w_n15280_0[0]),.dout(n15877),.clk(gclk));
	jand g15586(.dina(n15877),.dinb(w_n15278_0[0]),.dout(n15878),.clk(gclk));
	jand g15587(.dina(n15878),.dinb(w_asqrt10_15[1]),.dout(n15879),.clk(gclk));
	jxor g15588(.dina(n15879),.dinb(w_n15288_0[0]),.dout(n15880),.clk(gclk));
	jnot g15589(.din(n15880),.dout(n15881),.clk(gclk));
	jor g15590(.dina(w_n15868_0[1]),.dinb(w_asqrt58_13[0]),.dout(n15882),.clk(gclk));
	jor g15591(.dina(n15882),.dinb(w_n15874_0[1]),.dout(n15883),.clk(gclk));
	jand g15592(.dina(w_n15883_0[1]),.dinb(w_n15881_0[1]),.dout(n15884),.clk(gclk));
	jor g15593(.dina(w_n15884_0[1]),.dinb(w_n15876_0[1]),.dout(n15885),.clk(gclk));
	jand g15594(.dina(w_n15885_0[2]),.dinb(w_asqrt59_13[0]),.dout(n15886),.clk(gclk));
	jor g15595(.dina(w_n15885_0[1]),.dinb(w_asqrt59_12[2]),.dout(n15887),.clk(gclk));
	jnot g15596(.din(w_n15294_0[0]),.dout(n15888),.clk(gclk));
	jnot g15597(.din(w_n15295_0[0]),.dout(n15889),.clk(gclk));
	jand g15598(.dina(w_asqrt10_15[0]),.dinb(w_n15291_0[0]),.dout(n15890),.clk(gclk));
	jand g15599(.dina(w_n15890_0[1]),.dinb(n15889),.dout(n15891),.clk(gclk));
	jor g15600(.dina(n15891),.dinb(n15888),.dout(n15892),.clk(gclk));
	jnot g15601(.din(w_n15296_0[0]),.dout(n15893),.clk(gclk));
	jand g15602(.dina(w_n15890_0[0]),.dinb(n15893),.dout(n15894),.clk(gclk));
	jnot g15603(.din(n15894),.dout(n15895),.clk(gclk));
	jand g15604(.dina(n15895),.dinb(n15892),.dout(n15896),.clk(gclk));
	jand g15605(.dina(w_n15896_0[1]),.dinb(n15887),.dout(n15897),.clk(gclk));
	jor g15606(.dina(w_n15897_0[1]),.dinb(w_n15886_0[1]),.dout(n15898),.clk(gclk));
	jand g15607(.dina(n15898),.dinb(w_asqrt60_13[0]),.dout(n15899),.clk(gclk));
	jor g15608(.dina(w_n15886_0[0]),.dinb(w_asqrt60_12[2]),.dout(n15900),.clk(gclk));
	jor g15609(.dina(n15900),.dinb(w_n15897_0[0]),.dout(n15901),.clk(gclk));
	jnot g15610(.din(w_n15302_0[0]),.dout(n15902),.clk(gclk));
	jnot g15611(.din(w_n15304_0[0]),.dout(n15903),.clk(gclk));
	jand g15612(.dina(w_asqrt10_14[2]),.dinb(w_n15298_0[0]),.dout(n15904),.clk(gclk));
	jand g15613(.dina(w_n15904_0[1]),.dinb(n15903),.dout(n15905),.clk(gclk));
	jor g15614(.dina(n15905),.dinb(n15902),.dout(n15906),.clk(gclk));
	jnot g15615(.din(w_n15305_0[0]),.dout(n15907),.clk(gclk));
	jand g15616(.dina(w_n15904_0[0]),.dinb(n15907),.dout(n15908),.clk(gclk));
	jnot g15617(.din(n15908),.dout(n15909),.clk(gclk));
	jand g15618(.dina(n15909),.dinb(n15906),.dout(n15910),.clk(gclk));
	jand g15619(.dina(w_n15910_0[1]),.dinb(w_n15901_0[1]),.dout(n15911),.clk(gclk));
	jor g15620(.dina(n15911),.dinb(w_n15899_0[1]),.dout(n15912),.clk(gclk));
	jand g15621(.dina(w_n15912_0[1]),.dinb(w_asqrt61_13[1]),.dout(n15913),.clk(gclk));
	jxor g15622(.dina(w_n15306_0[0]),.dinb(w_n290_17[0]),.dout(n15914),.clk(gclk));
	jand g15623(.dina(n15914),.dinb(w_asqrt10_14[1]),.dout(n15915),.clk(gclk));
	jxor g15624(.dina(n15915),.dinb(w_n15316_0[0]),.dout(n15916),.clk(gclk));
	jnot g15625(.din(n15916),.dout(n15917),.clk(gclk));
	jor g15626(.dina(w_n15912_0[0]),.dinb(w_asqrt61_13[0]),.dout(n15918),.clk(gclk));
	jand g15627(.dina(w_n15918_0[1]),.dinb(w_n15917_0[1]),.dout(n15919),.clk(gclk));
	jor g15628(.dina(w_n15919_0[2]),.dinb(w_n15913_0[2]),.dout(n15920),.clk(gclk));
	jand g15629(.dina(n15920),.dinb(w_asqrt62_13[1]),.dout(n15921),.clk(gclk));
	jnot g15630(.din(w_n15321_0[0]),.dout(n15922),.clk(gclk));
	jand g15631(.dina(n15922),.dinb(w_n15319_0[0]),.dout(n15923),.clk(gclk));
	jand g15632(.dina(n15923),.dinb(w_asqrt10_14[0]),.dout(n15924),.clk(gclk));
	jxor g15633(.dina(n15924),.dinb(w_n15329_0[0]),.dout(n15925),.clk(gclk));
	jnot g15634(.din(n15925),.dout(n15926),.clk(gclk));
	jor g15635(.dina(w_n15913_0[1]),.dinb(w_asqrt62_13[0]),.dout(n15927),.clk(gclk));
	jor g15636(.dina(n15927),.dinb(w_n15919_0[1]),.dout(n15928),.clk(gclk));
	jand g15637(.dina(w_n15928_0[1]),.dinb(w_n15926_0[1]),.dout(n15929),.clk(gclk));
	jor g15638(.dina(w_n15929_0[1]),.dinb(w_n15921_0[1]),.dout(n15930),.clk(gclk));
	jxor g15639(.dina(w_n15331_0[0]),.dinb(w_n199_19[2]),.dout(n15931),.clk(gclk));
	jand g15640(.dina(n15931),.dinb(w_asqrt10_13[2]),.dout(n15932),.clk(gclk));
	jxor g15641(.dina(n15932),.dinb(w_n15336_0[0]),.dout(n15933),.clk(gclk));
	jnot g15642(.din(w_n15338_0[0]),.dout(n15934),.clk(gclk));
	jnot g15643(.din(w_n15342_0[0]),.dout(n15935),.clk(gclk));
	jand g15644(.dina(w_asqrt10_13[1]),.dinb(w_n15935_0[1]),.dout(n15936),.clk(gclk));
	jand g15645(.dina(w_n15936_0[1]),.dinb(w_n15934_0[2]),.dout(n15937),.clk(gclk));
	jor g15646(.dina(n15937),.dinb(w_n15349_0[0]),.dout(n15938),.clk(gclk));
	jor g15647(.dina(n15938),.dinb(w_n15933_0[1]),.dout(n15939),.clk(gclk));
	jnot g15648(.din(n15939),.dout(n15940),.clk(gclk));
	jand g15649(.dina(n15940),.dinb(w_n15930_1[2]),.dout(n15941),.clk(gclk));
	jor g15650(.dina(n15941),.dinb(w_asqrt63_7[1]),.dout(n15942),.clk(gclk));
	jnot g15651(.din(w_n15933_0[0]),.dout(n15943),.clk(gclk));
	jor g15652(.dina(w_n15943_0[2]),.dinb(w_n15930_1[1]),.dout(n15944),.clk(gclk));
	jor g15653(.dina(w_n15936_0[0]),.dinb(w_n15934_0[1]),.dout(n15945),.clk(gclk));
	jand g15654(.dina(w_n15935_0[0]),.dinb(w_n15934_0[0]),.dout(n15946),.clk(gclk));
	jor g15655(.dina(n15946),.dinb(w_n194_18[2]),.dout(n15947),.clk(gclk));
	jnot g15656(.din(n15947),.dout(n15948),.clk(gclk));
	jand g15657(.dina(n15948),.dinb(n15945),.dout(n15949),.clk(gclk));
	jnot g15658(.din(w_asqrt10_13[0]),.dout(n15950),.clk(gclk));
	jnot g15659(.din(w_n15949_0[1]),.dout(n15953),.clk(gclk));
	jand g15660(.dina(n15953),.dinb(w_n15944_0[1]),.dout(n15954),.clk(gclk));
	jand g15661(.dina(n15954),.dinb(w_n15942_0[1]),.dout(n15955),.clk(gclk));
	jxor g15662(.dina(w_n15822_0[0]),.dinb(w_n796_16[1]),.dout(n15956),.clk(gclk));
	jor g15663(.dina(n15956),.dinb(w_n15955_21[1]),.dout(n15957),.clk(gclk));
	jxor g15664(.dina(n15957),.dinb(n15362),.dout(n15958),.clk(gclk));
	jnot g15665(.din(n15958),.dout(n15959),.clk(gclk));
	jor g15666(.dina(w_n15955_21[0]),.dinb(w_n15364_1[0]),.dout(n15960),.clk(gclk));
	jnot g15667(.din(w_a16_0[1]),.dout(n15961),.clk(gclk));
	jnot g15668(.din(a[17]),.dout(n15962),.clk(gclk));
	jand g15669(.dina(w_n15364_0[2]),.dinb(w_n15962_0[2]),.dout(n15963),.clk(gclk));
	jand g15670(.dina(n15963),.dinb(w_n15961_1[1]),.dout(n15964),.clk(gclk));
	jnot g15671(.din(n15964),.dout(n15965),.clk(gclk));
	jand g15672(.dina(n15965),.dinb(n15960),.dout(n15966),.clk(gclk));
	jor g15673(.dina(w_n15966_0[2]),.dinb(w_n15950_6[2]),.dout(n15967),.clk(gclk));
	jor g15674(.dina(w_n15955_20[2]),.dinb(w_a18_0[0]),.dout(n15968),.clk(gclk));
	jxor g15675(.dina(w_n15968_0[1]),.dinb(w_n15365_0[0]),.dout(n15969),.clk(gclk));
	jand g15676(.dina(w_n15966_0[1]),.dinb(w_n15950_6[1]),.dout(n15970),.clk(gclk));
	jor g15677(.dina(n15970),.dinb(w_n15969_0[1]),.dout(n15971),.clk(gclk));
	jand g15678(.dina(w_n15971_0[1]),.dinb(w_n15967_0[1]),.dout(n15972),.clk(gclk));
	jor g15679(.dina(n15972),.dinb(w_n14821_12[0]),.dout(n15973),.clk(gclk));
	jand g15680(.dina(w_n15967_0[0]),.dinb(w_n14821_11[2]),.dout(n15974),.clk(gclk));
	jand g15681(.dina(n15974),.dinb(w_n15971_0[0]),.dout(n15975),.clk(gclk));
	jor g15682(.dina(w_n15968_0[0]),.dinb(w_a19_0[0]),.dout(n15976),.clk(gclk));
	jnot g15683(.din(w_n15942_0[0]),.dout(n15977),.clk(gclk));
	jnot g15684(.din(w_n15944_0[0]),.dout(n15978),.clk(gclk));
	jor g15685(.dina(w_n15949_0[0]),.dinb(w_n15950_6[0]),.dout(n15979),.clk(gclk));
	jor g15686(.dina(n15979),.dinb(w_n15978_0[1]),.dout(n15980),.clk(gclk));
	jor g15687(.dina(n15980),.dinb(n15977),.dout(n15981),.clk(gclk));
	jand g15688(.dina(n15981),.dinb(n15976),.dout(n15982),.clk(gclk));
	jxor g15689(.dina(n15982),.dinb(w_n14826_0[1]),.dout(n15983),.clk(gclk));
	jor g15690(.dina(w_n15983_0[1]),.dinb(w_n15975_0[1]),.dout(n15984),.clk(gclk));
	jand g15691(.dina(n15984),.dinb(w_n15973_0[1]),.dout(n15985),.clk(gclk));
	jor g15692(.dina(w_n15985_0[2]),.dinb(w_n14816_7[0]),.dout(n15986),.clk(gclk));
	jand g15693(.dina(w_n15985_0[1]),.dinb(w_n14816_6[2]),.dout(n15987),.clk(gclk));
	jxor g15694(.dina(w_n15368_0[0]),.dinb(w_n14821_11[1]),.dout(n15988),.clk(gclk));
	jor g15695(.dina(n15988),.dinb(w_n15955_20[1]),.dout(n15989),.clk(gclk));
	jxor g15696(.dina(n15989),.dinb(w_n15371_0[0]),.dout(n15990),.clk(gclk));
	jor g15697(.dina(w_n15990_0[1]),.dinb(n15987),.dout(n15991),.clk(gclk));
	jand g15698(.dina(w_n15991_0[1]),.dinb(w_n15986_0[1]),.dout(n15992),.clk(gclk));
	jor g15699(.dina(n15992),.dinb(w_n13723_11[2]),.dout(n15993),.clk(gclk));
	jnot g15700(.din(w_n15377_0[0]),.dout(n15994),.clk(gclk));
	jor g15701(.dina(n15994),.dinb(w_n15375_0[0]),.dout(n15995),.clk(gclk));
	jor g15702(.dina(n15995),.dinb(w_n15955_20[0]),.dout(n15996),.clk(gclk));
	jxor g15703(.dina(n15996),.dinb(w_n15386_0[0]),.dout(n15997),.clk(gclk));
	jand g15704(.dina(w_n15986_0[0]),.dinb(w_n13723_11[1]),.dout(n15998),.clk(gclk));
	jand g15705(.dina(n15998),.dinb(w_n15991_0[0]),.dout(n15999),.clk(gclk));
	jor g15706(.dina(w_n15999_0[1]),.dinb(w_n15997_0[1]),.dout(n16000),.clk(gclk));
	jand g15707(.dina(w_n16000_0[1]),.dinb(w_n15993_0[1]),.dout(n16001),.clk(gclk));
	jor g15708(.dina(w_n16001_0[2]),.dinb(w_n13718_7[0]),.dout(n16002),.clk(gclk));
	jand g15709(.dina(w_n16001_0[1]),.dinb(w_n13718_6[2]),.dout(n16003),.clk(gclk));
	jxor g15710(.dina(w_n15388_0[0]),.dinb(w_n13723_11[0]),.dout(n16004),.clk(gclk));
	jor g15711(.dina(n16004),.dinb(w_n15955_19[2]),.dout(n16005),.clk(gclk));
	jxor g15712(.dina(n16005),.dinb(w_n15393_0[0]),.dout(n16006),.clk(gclk));
	jnot g15713(.din(w_n16006_0[1]),.dout(n16007),.clk(gclk));
	jor g15714(.dina(n16007),.dinb(n16003),.dout(n16008),.clk(gclk));
	jand g15715(.dina(w_n16008_0[1]),.dinb(w_n16002_0[1]),.dout(n16009),.clk(gclk));
	jor g15716(.dina(n16009),.dinb(w_n12675_12[1]),.dout(n16010),.clk(gclk));
	jand g15717(.dina(w_n16002_0[0]),.dinb(w_n12675_12[0]),.dout(n16011),.clk(gclk));
	jand g15718(.dina(n16011),.dinb(w_n16008_0[0]),.dout(n16012),.clk(gclk));
	jnot g15719(.din(w_n15397_0[0]),.dout(n16013),.clk(gclk));
	jnot g15720(.din(w_n15955_19[1]),.dout(asqrt_fa_10),.clk(gclk));
	jand g15721(.dina(w_asqrt9_16),.dinb(n16013),.dout(n16015),.clk(gclk));
	jand g15722(.dina(w_n16015_0[1]),.dinb(w_n15404_0[0]),.dout(n16016),.clk(gclk));
	jor g15723(.dina(n16016),.dinb(w_n15402_0[0]),.dout(n16017),.clk(gclk));
	jand g15724(.dina(w_n16015_0[0]),.dinb(w_n15405_0[0]),.dout(n16018),.clk(gclk));
	jnot g15725(.din(n16018),.dout(n16019),.clk(gclk));
	jand g15726(.dina(n16019),.dinb(n16017),.dout(n16020),.clk(gclk));
	jnot g15727(.din(n16020),.dout(n16021),.clk(gclk));
	jor g15728(.dina(w_n16021_0[1]),.dinb(w_n16012_0[1]),.dout(n16022),.clk(gclk));
	jand g15729(.dina(n16022),.dinb(w_n16010_0[1]),.dout(n16023),.clk(gclk));
	jor g15730(.dina(w_n16023_0[2]),.dinb(w_n12670_7[1]),.dout(n16024),.clk(gclk));
	jand g15731(.dina(w_n16023_0[1]),.dinb(w_n12670_7[0]),.dout(n16025),.clk(gclk));
	jnot g15732(.din(w_n15412_0[0]),.dout(n16026),.clk(gclk));
	jxor g15733(.dina(w_n15406_0[0]),.dinb(w_n12675_11[2]),.dout(n16027),.clk(gclk));
	jor g15734(.dina(n16027),.dinb(w_n15955_19[0]),.dout(n16028),.clk(gclk));
	jxor g15735(.dina(n16028),.dinb(n16026),.dout(n16029),.clk(gclk));
	jnot g15736(.din(w_n16029_0[1]),.dout(n16030),.clk(gclk));
	jor g15737(.dina(n16030),.dinb(n16025),.dout(n16031),.clk(gclk));
	jand g15738(.dina(w_n16031_0[1]),.dinb(w_n16024_0[1]),.dout(n16032),.clk(gclk));
	jor g15739(.dina(n16032),.dinb(w_n11662_12[0]),.dout(n16033),.clk(gclk));
	jnot g15740(.din(w_n15417_0[0]),.dout(n16034),.clk(gclk));
	jor g15741(.dina(n16034),.dinb(w_n15415_0[0]),.dout(n16035),.clk(gclk));
	jor g15742(.dina(n16035),.dinb(w_n15955_18[2]),.dout(n16036),.clk(gclk));
	jxor g15743(.dina(n16036),.dinb(w_n15426_0[0]),.dout(n16037),.clk(gclk));
	jand g15744(.dina(w_n16024_0[0]),.dinb(w_n11662_11[2]),.dout(n16038),.clk(gclk));
	jand g15745(.dina(n16038),.dinb(w_n16031_0[0]),.dout(n16039),.clk(gclk));
	jor g15746(.dina(w_n16039_0[1]),.dinb(w_n16037_0[1]),.dout(n16040),.clk(gclk));
	jand g15747(.dina(w_n16040_0[1]),.dinb(w_n16033_0[1]),.dout(n16041),.clk(gclk));
	jor g15748(.dina(w_n16041_0[2]),.dinb(w_n11657_7[1]),.dout(n16042),.clk(gclk));
	jand g15749(.dina(w_n16041_0[1]),.dinb(w_n11657_7[0]),.dout(n16043),.clk(gclk));
	jnot g15750(.din(w_n15433_0[0]),.dout(n16044),.clk(gclk));
	jxor g15751(.dina(w_n15428_0[0]),.dinb(w_n11662_11[1]),.dout(n16045),.clk(gclk));
	jor g15752(.dina(n16045),.dinb(w_n15955_18[1]),.dout(n16046),.clk(gclk));
	jxor g15753(.dina(n16046),.dinb(n16044),.dout(n16047),.clk(gclk));
	jnot g15754(.din(n16047),.dout(n16048),.clk(gclk));
	jor g15755(.dina(w_n16048_0[1]),.dinb(n16043),.dout(n16049),.clk(gclk));
	jand g15756(.dina(w_n16049_0[1]),.dinb(w_n16042_0[1]),.dout(n16050),.clk(gclk));
	jor g15757(.dina(n16050),.dinb(w_n10701_12[1]),.dout(n16051),.clk(gclk));
	jand g15758(.dina(w_n16042_0[0]),.dinb(w_n10701_12[0]),.dout(n16052),.clk(gclk));
	jand g15759(.dina(n16052),.dinb(w_n16049_0[0]),.dout(n16053),.clk(gclk));
	jnot g15760(.din(w_n15436_0[0]),.dout(n16054),.clk(gclk));
	jand g15761(.dina(w_asqrt9_15[2]),.dinb(n16054),.dout(n16055),.clk(gclk));
	jand g15762(.dina(w_n16055_0[1]),.dinb(w_n15443_0[0]),.dout(n16056),.clk(gclk));
	jor g15763(.dina(n16056),.dinb(w_n15441_0[0]),.dout(n16057),.clk(gclk));
	jand g15764(.dina(w_n16055_0[0]),.dinb(w_n15444_0[0]),.dout(n16058),.clk(gclk));
	jnot g15765(.din(n16058),.dout(n16059),.clk(gclk));
	jand g15766(.dina(n16059),.dinb(n16057),.dout(n16060),.clk(gclk));
	jnot g15767(.din(n16060),.dout(n16061),.clk(gclk));
	jor g15768(.dina(w_n16061_0[1]),.dinb(w_n16053_0[1]),.dout(n16062),.clk(gclk));
	jand g15769(.dina(n16062),.dinb(w_n16051_0[1]),.dout(n16063),.clk(gclk));
	jor g15770(.dina(w_n16063_0[1]),.dinb(w_n10696_8[0]),.dout(n16064),.clk(gclk));
	jxor g15771(.dina(w_n15445_0[0]),.dinb(w_n10701_11[2]),.dout(n16065),.clk(gclk));
	jor g15772(.dina(n16065),.dinb(w_n15955_18[0]),.dout(n16066),.clk(gclk));
	jxor g15773(.dina(n16066),.dinb(w_n15450_0[0]),.dout(n16067),.clk(gclk));
	jand g15774(.dina(w_n16063_0[0]),.dinb(w_n10696_7[2]),.dout(n16068),.clk(gclk));
	jor g15775(.dina(w_n16068_0[1]),.dinb(w_n16067_0[1]),.dout(n16069),.clk(gclk));
	jand g15776(.dina(w_n16069_0[2]),.dinb(w_n16064_0[2]),.dout(n16070),.clk(gclk));
	jor g15777(.dina(n16070),.dinb(w_n9774_12[0]),.dout(n16071),.clk(gclk));
	jnot g15778(.din(w_n15455_0[0]),.dout(n16072),.clk(gclk));
	jor g15779(.dina(n16072),.dinb(w_n15453_0[0]),.dout(n16073),.clk(gclk));
	jor g15780(.dina(n16073),.dinb(w_n15955_17[2]),.dout(n16074),.clk(gclk));
	jxor g15781(.dina(n16074),.dinb(w_n15464_0[0]),.dout(n16075),.clk(gclk));
	jand g15782(.dina(w_n16064_0[1]),.dinb(w_n9774_11[2]),.dout(n16076),.clk(gclk));
	jand g15783(.dina(n16076),.dinb(w_n16069_0[1]),.dout(n16077),.clk(gclk));
	jor g15784(.dina(w_n16077_0[1]),.dinb(w_n16075_0[1]),.dout(n16078),.clk(gclk));
	jand g15785(.dina(w_n16078_0[1]),.dinb(w_n16071_0[1]),.dout(n16079),.clk(gclk));
	jor g15786(.dina(w_n16079_0[2]),.dinb(w_n9769_8[1]),.dout(n16080),.clk(gclk));
	jand g15787(.dina(w_n16079_0[1]),.dinb(w_n9769_8[0]),.dout(n16081),.clk(gclk));
	jnot g15788(.din(w_n15467_0[0]),.dout(n16082),.clk(gclk));
	jand g15789(.dina(w_asqrt9_15[1]),.dinb(n16082),.dout(n16083),.clk(gclk));
	jand g15790(.dina(w_n16083_0[1]),.dinb(w_n15472_0[0]),.dout(n16084),.clk(gclk));
	jor g15791(.dina(n16084),.dinb(w_n15471_0[0]),.dout(n16085),.clk(gclk));
	jand g15792(.dina(w_n16083_0[0]),.dinb(w_n15473_0[0]),.dout(n16086),.clk(gclk));
	jnot g15793(.din(n16086),.dout(n16087),.clk(gclk));
	jand g15794(.dina(n16087),.dinb(n16085),.dout(n16088),.clk(gclk));
	jnot g15795(.din(n16088),.dout(n16089),.clk(gclk));
	jor g15796(.dina(w_n16089_0[1]),.dinb(n16081),.dout(n16090),.clk(gclk));
	jand g15797(.dina(w_n16090_0[1]),.dinb(w_n16080_0[1]),.dout(n16091),.clk(gclk));
	jor g15798(.dina(n16091),.dinb(w_n8898_13[0]),.dout(n16092),.clk(gclk));
	jand g15799(.dina(w_n16080_0[0]),.dinb(w_n8898_12[2]),.dout(n16093),.clk(gclk));
	jand g15800(.dina(n16093),.dinb(w_n16090_0[0]),.dout(n16094),.clk(gclk));
	jnot g15801(.din(w_n15475_0[0]),.dout(n16095),.clk(gclk));
	jand g15802(.dina(w_asqrt9_15[0]),.dinb(n16095),.dout(n16096),.clk(gclk));
	jand g15803(.dina(w_n16096_0[1]),.dinb(w_n15482_0[0]),.dout(n16097),.clk(gclk));
	jor g15804(.dina(n16097),.dinb(w_n15480_0[0]),.dout(n16098),.clk(gclk));
	jand g15805(.dina(w_n16096_0[0]),.dinb(w_n15483_0[0]),.dout(n16099),.clk(gclk));
	jnot g15806(.din(n16099),.dout(n16100),.clk(gclk));
	jand g15807(.dina(n16100),.dinb(n16098),.dout(n16101),.clk(gclk));
	jnot g15808(.din(n16101),.dout(n16102),.clk(gclk));
	jor g15809(.dina(w_n16102_0[1]),.dinb(w_n16094_0[1]),.dout(n16103),.clk(gclk));
	jand g15810(.dina(n16103),.dinb(w_n16092_0[1]),.dout(n16104),.clk(gclk));
	jor g15811(.dina(w_n16104_0[1]),.dinb(w_n8893_8[2]),.dout(n16105),.clk(gclk));
	jxor g15812(.dina(w_n15484_0[0]),.dinb(w_n8898_12[1]),.dout(n16106),.clk(gclk));
	jor g15813(.dina(n16106),.dinb(w_n15955_17[1]),.dout(n16107),.clk(gclk));
	jxor g15814(.dina(n16107),.dinb(w_n15495_0[0]),.dout(n16108),.clk(gclk));
	jand g15815(.dina(w_n16104_0[0]),.dinb(w_n8893_8[1]),.dout(n16109),.clk(gclk));
	jor g15816(.dina(w_n16109_0[1]),.dinb(w_n16108_0[1]),.dout(n16110),.clk(gclk));
	jand g15817(.dina(w_n16110_0[2]),.dinb(w_n16105_0[2]),.dout(n16111),.clk(gclk));
	jor g15818(.dina(n16111),.dinb(w_n8058_12[2]),.dout(n16112),.clk(gclk));
	jnot g15819(.din(w_n15500_0[0]),.dout(n16113),.clk(gclk));
	jor g15820(.dina(n16113),.dinb(w_n15498_0[0]),.dout(n16114),.clk(gclk));
	jor g15821(.dina(n16114),.dinb(w_n15955_17[0]),.dout(n16115),.clk(gclk));
	jxor g15822(.dina(n16115),.dinb(w_n15509_0[0]),.dout(n16116),.clk(gclk));
	jand g15823(.dina(w_n16105_0[1]),.dinb(w_n8058_12[1]),.dout(n16117),.clk(gclk));
	jand g15824(.dina(n16117),.dinb(w_n16110_0[1]),.dout(n16118),.clk(gclk));
	jor g15825(.dina(w_n16118_0[1]),.dinb(w_n16116_0[1]),.dout(n16119),.clk(gclk));
	jand g15826(.dina(w_n16119_0[1]),.dinb(w_n16112_0[1]),.dout(n16120),.clk(gclk));
	jor g15827(.dina(w_n16120_0[2]),.dinb(w_n8053_9[0]),.dout(n16121),.clk(gclk));
	jand g15828(.dina(w_n16120_0[1]),.dinb(w_n8053_8[2]),.dout(n16122),.clk(gclk));
	jnot g15829(.din(w_n15512_0[0]),.dout(n16123),.clk(gclk));
	jand g15830(.dina(w_asqrt9_14[2]),.dinb(n16123),.dout(n16124),.clk(gclk));
	jand g15831(.dina(w_n16124_0[1]),.dinb(w_n15517_0[0]),.dout(n16125),.clk(gclk));
	jor g15832(.dina(n16125),.dinb(w_n15516_0[0]),.dout(n16126),.clk(gclk));
	jand g15833(.dina(w_n16124_0[0]),.dinb(w_n15518_0[0]),.dout(n16127),.clk(gclk));
	jnot g15834(.din(n16127),.dout(n16128),.clk(gclk));
	jand g15835(.dina(n16128),.dinb(n16126),.dout(n16129),.clk(gclk));
	jnot g15836(.din(n16129),.dout(n16130),.clk(gclk));
	jor g15837(.dina(w_n16130_0[1]),.dinb(n16122),.dout(n16131),.clk(gclk));
	jand g15838(.dina(w_n16131_0[1]),.dinb(w_n16121_0[1]),.dout(n16132),.clk(gclk));
	jor g15839(.dina(n16132),.dinb(w_n7265_13[1]),.dout(n16133),.clk(gclk));
	jand g15840(.dina(w_n16121_0[0]),.dinb(w_n7265_13[0]),.dout(n16134),.clk(gclk));
	jand g15841(.dina(n16134),.dinb(w_n16131_0[0]),.dout(n16135),.clk(gclk));
	jnot g15842(.din(w_n15520_0[0]),.dout(n16136),.clk(gclk));
	jand g15843(.dina(w_asqrt9_14[1]),.dinb(n16136),.dout(n16137),.clk(gclk));
	jand g15844(.dina(w_n16137_0[1]),.dinb(w_n15527_0[0]),.dout(n16138),.clk(gclk));
	jor g15845(.dina(n16138),.dinb(w_n15525_0[0]),.dout(n16139),.clk(gclk));
	jand g15846(.dina(w_n16137_0[0]),.dinb(w_n15528_0[0]),.dout(n16140),.clk(gclk));
	jnot g15847(.din(n16140),.dout(n16141),.clk(gclk));
	jand g15848(.dina(n16141),.dinb(n16139),.dout(n16142),.clk(gclk));
	jnot g15849(.din(n16142),.dout(n16143),.clk(gclk));
	jor g15850(.dina(w_n16143_0[1]),.dinb(w_n16135_0[1]),.dout(n16144),.clk(gclk));
	jand g15851(.dina(n16144),.dinb(w_n16133_0[1]),.dout(n16145),.clk(gclk));
	jor g15852(.dina(w_n16145_0[1]),.dinb(w_n7260_9[2]),.dout(n16146),.clk(gclk));
	jxor g15853(.dina(w_n15529_0[0]),.dinb(w_n7265_12[2]),.dout(n16147),.clk(gclk));
	jor g15854(.dina(n16147),.dinb(w_n15955_16[2]),.dout(n16148),.clk(gclk));
	jxor g15855(.dina(n16148),.dinb(w_n15540_0[0]),.dout(n16149),.clk(gclk));
	jand g15856(.dina(w_n16145_0[0]),.dinb(w_n7260_9[1]),.dout(n16150),.clk(gclk));
	jor g15857(.dina(w_n16150_0[1]),.dinb(w_n16149_0[1]),.dout(n16151),.clk(gclk));
	jand g15858(.dina(w_n16151_0[2]),.dinb(w_n16146_0[2]),.dout(n16152),.clk(gclk));
	jor g15859(.dina(n16152),.dinb(w_n6505_13[0]),.dout(n16153),.clk(gclk));
	jnot g15860(.din(w_n15545_0[0]),.dout(n16154),.clk(gclk));
	jor g15861(.dina(n16154),.dinb(w_n15543_0[0]),.dout(n16155),.clk(gclk));
	jor g15862(.dina(n16155),.dinb(w_n15955_16[1]),.dout(n16156),.clk(gclk));
	jxor g15863(.dina(n16156),.dinb(w_n15554_0[0]),.dout(n16157),.clk(gclk));
	jand g15864(.dina(w_n16146_0[1]),.dinb(w_n6505_12[2]),.dout(n16158),.clk(gclk));
	jand g15865(.dina(n16158),.dinb(w_n16151_0[1]),.dout(n16159),.clk(gclk));
	jor g15866(.dina(w_n16159_0[1]),.dinb(w_n16157_0[1]),.dout(n16160),.clk(gclk));
	jand g15867(.dina(w_n16160_0[1]),.dinb(w_n16153_0[1]),.dout(n16161),.clk(gclk));
	jor g15868(.dina(w_n16161_0[2]),.dinb(w_n6500_10[0]),.dout(n16162),.clk(gclk));
	jand g15869(.dina(w_n16161_0[1]),.dinb(w_n6500_9[2]),.dout(n16163),.clk(gclk));
	jnot g15870(.din(w_n15557_0[0]),.dout(n16164),.clk(gclk));
	jand g15871(.dina(w_asqrt9_14[0]),.dinb(n16164),.dout(n16165),.clk(gclk));
	jand g15872(.dina(w_n16165_0[1]),.dinb(w_n15562_0[0]),.dout(n16166),.clk(gclk));
	jor g15873(.dina(n16166),.dinb(w_n15561_0[0]),.dout(n16167),.clk(gclk));
	jand g15874(.dina(w_n16165_0[0]),.dinb(w_n15563_0[0]),.dout(n16168),.clk(gclk));
	jnot g15875(.din(n16168),.dout(n16169),.clk(gclk));
	jand g15876(.dina(n16169),.dinb(n16167),.dout(n16170),.clk(gclk));
	jnot g15877(.din(n16170),.dout(n16171),.clk(gclk));
	jor g15878(.dina(w_n16171_0[1]),.dinb(n16163),.dout(n16172),.clk(gclk));
	jand g15879(.dina(w_n16172_0[1]),.dinb(w_n16162_0[1]),.dout(n16173),.clk(gclk));
	jor g15880(.dina(n16173),.dinb(w_n5793_13[2]),.dout(n16174),.clk(gclk));
	jand g15881(.dina(w_n16162_0[0]),.dinb(w_n5793_13[1]),.dout(n16175),.clk(gclk));
	jand g15882(.dina(n16175),.dinb(w_n16172_0[0]),.dout(n16176),.clk(gclk));
	jnot g15883(.din(w_n15565_0[0]),.dout(n16177),.clk(gclk));
	jand g15884(.dina(w_asqrt9_13[2]),.dinb(n16177),.dout(n16178),.clk(gclk));
	jand g15885(.dina(w_n16178_0[1]),.dinb(w_n15572_0[0]),.dout(n16179),.clk(gclk));
	jor g15886(.dina(n16179),.dinb(w_n15570_0[0]),.dout(n16180),.clk(gclk));
	jand g15887(.dina(w_n16178_0[0]),.dinb(w_n15573_0[0]),.dout(n16181),.clk(gclk));
	jnot g15888(.din(n16181),.dout(n16182),.clk(gclk));
	jand g15889(.dina(n16182),.dinb(n16180),.dout(n16183),.clk(gclk));
	jnot g15890(.din(n16183),.dout(n16184),.clk(gclk));
	jor g15891(.dina(w_n16184_0[1]),.dinb(w_n16176_0[1]),.dout(n16185),.clk(gclk));
	jand g15892(.dina(n16185),.dinb(w_n16174_0[1]),.dout(n16186),.clk(gclk));
	jor g15893(.dina(w_n16186_0[1]),.dinb(w_n5788_10[1]),.dout(n16187),.clk(gclk));
	jxor g15894(.dina(w_n15574_0[0]),.dinb(w_n5793_13[0]),.dout(n16188),.clk(gclk));
	jor g15895(.dina(n16188),.dinb(w_n15955_16[0]),.dout(n16189),.clk(gclk));
	jxor g15896(.dina(n16189),.dinb(w_n15585_0[0]),.dout(n16190),.clk(gclk));
	jand g15897(.dina(w_n16186_0[0]),.dinb(w_n5788_10[0]),.dout(n16191),.clk(gclk));
	jor g15898(.dina(w_n16191_0[1]),.dinb(w_n16190_0[1]),.dout(n16192),.clk(gclk));
	jand g15899(.dina(w_n16192_0[2]),.dinb(w_n16187_0[2]),.dout(n16193),.clk(gclk));
	jor g15900(.dina(n16193),.dinb(w_n5121_13[1]),.dout(n16194),.clk(gclk));
	jnot g15901(.din(w_n15590_0[0]),.dout(n16195),.clk(gclk));
	jor g15902(.dina(n16195),.dinb(w_n15588_0[0]),.dout(n16196),.clk(gclk));
	jor g15903(.dina(n16196),.dinb(w_n15955_15[2]),.dout(n16197),.clk(gclk));
	jxor g15904(.dina(n16197),.dinb(w_n15599_0[0]),.dout(n16198),.clk(gclk));
	jand g15905(.dina(w_n16187_0[1]),.dinb(w_n5121_13[0]),.dout(n16199),.clk(gclk));
	jand g15906(.dina(n16199),.dinb(w_n16192_0[1]),.dout(n16200),.clk(gclk));
	jor g15907(.dina(w_n16200_0[1]),.dinb(w_n16198_0[1]),.dout(n16201),.clk(gclk));
	jand g15908(.dina(w_n16201_0[1]),.dinb(w_n16194_0[1]),.dout(n16202),.clk(gclk));
	jor g15909(.dina(w_n16202_0[2]),.dinb(w_n5116_10[2]),.dout(n16203),.clk(gclk));
	jand g15910(.dina(w_n16202_0[1]),.dinb(w_n5116_10[1]),.dout(n16204),.clk(gclk));
	jnot g15911(.din(w_n15602_0[0]),.dout(n16205),.clk(gclk));
	jand g15912(.dina(w_asqrt9_13[1]),.dinb(n16205),.dout(n16206),.clk(gclk));
	jand g15913(.dina(w_n16206_0[1]),.dinb(w_n15607_0[0]),.dout(n16207),.clk(gclk));
	jor g15914(.dina(n16207),.dinb(w_n15606_0[0]),.dout(n16208),.clk(gclk));
	jand g15915(.dina(w_n16206_0[0]),.dinb(w_n15608_0[0]),.dout(n16209),.clk(gclk));
	jnot g15916(.din(n16209),.dout(n16210),.clk(gclk));
	jand g15917(.dina(n16210),.dinb(n16208),.dout(n16211),.clk(gclk));
	jnot g15918(.din(n16211),.dout(n16212),.clk(gclk));
	jor g15919(.dina(w_n16212_0[1]),.dinb(n16204),.dout(n16213),.clk(gclk));
	jand g15920(.dina(w_n16213_0[1]),.dinb(w_n16203_0[1]),.dout(n16214),.clk(gclk));
	jor g15921(.dina(n16214),.dinb(w_n4499_14[1]),.dout(n16215),.clk(gclk));
	jand g15922(.dina(w_n16203_0[0]),.dinb(w_n4499_14[0]),.dout(n16216),.clk(gclk));
	jand g15923(.dina(n16216),.dinb(w_n16213_0[0]),.dout(n16217),.clk(gclk));
	jnot g15924(.din(w_n15610_0[0]),.dout(n16218),.clk(gclk));
	jand g15925(.dina(w_asqrt9_13[0]),.dinb(n16218),.dout(n16219),.clk(gclk));
	jand g15926(.dina(w_n16219_0[1]),.dinb(w_n15617_0[0]),.dout(n16220),.clk(gclk));
	jor g15927(.dina(n16220),.dinb(w_n15615_0[0]),.dout(n16221),.clk(gclk));
	jand g15928(.dina(w_n16219_0[0]),.dinb(w_n15618_0[0]),.dout(n16222),.clk(gclk));
	jnot g15929(.din(n16222),.dout(n16223),.clk(gclk));
	jand g15930(.dina(n16223),.dinb(n16221),.dout(n16224),.clk(gclk));
	jnot g15931(.din(n16224),.dout(n16225),.clk(gclk));
	jor g15932(.dina(w_n16225_0[1]),.dinb(w_n16217_0[1]),.dout(n16226),.clk(gclk));
	jand g15933(.dina(n16226),.dinb(w_n16215_0[1]),.dout(n16227),.clk(gclk));
	jor g15934(.dina(w_n16227_0[1]),.dinb(w_n4494_11[1]),.dout(n16228),.clk(gclk));
	jxor g15935(.dina(w_n15619_0[0]),.dinb(w_n4499_13[2]),.dout(n16229),.clk(gclk));
	jor g15936(.dina(n16229),.dinb(w_n15955_15[1]),.dout(n16230),.clk(gclk));
	jxor g15937(.dina(n16230),.dinb(w_n15630_0[0]),.dout(n16231),.clk(gclk));
	jand g15938(.dina(w_n16227_0[0]),.dinb(w_n4494_11[0]),.dout(n16232),.clk(gclk));
	jor g15939(.dina(w_n16232_0[1]),.dinb(w_n16231_0[1]),.dout(n16233),.clk(gclk));
	jand g15940(.dina(w_n16233_0[2]),.dinb(w_n16228_0[2]),.dout(n16234),.clk(gclk));
	jor g15941(.dina(n16234),.dinb(w_n3912_14[0]),.dout(n16235),.clk(gclk));
	jnot g15942(.din(w_n15635_0[0]),.dout(n16236),.clk(gclk));
	jor g15943(.dina(n16236),.dinb(w_n15633_0[0]),.dout(n16237),.clk(gclk));
	jor g15944(.dina(n16237),.dinb(w_n15955_15[0]),.dout(n16238),.clk(gclk));
	jxor g15945(.dina(n16238),.dinb(w_n15644_0[0]),.dout(n16239),.clk(gclk));
	jand g15946(.dina(w_n16228_0[1]),.dinb(w_n3912_13[2]),.dout(n16240),.clk(gclk));
	jand g15947(.dina(n16240),.dinb(w_n16233_0[1]),.dout(n16241),.clk(gclk));
	jor g15948(.dina(w_n16241_0[1]),.dinb(w_n16239_0[1]),.dout(n16242),.clk(gclk));
	jand g15949(.dina(w_n16242_0[1]),.dinb(w_n16235_0[1]),.dout(n16243),.clk(gclk));
	jor g15950(.dina(w_n16243_0[2]),.dinb(w_n3907_11[2]),.dout(n16244),.clk(gclk));
	jand g15951(.dina(w_n16243_0[1]),.dinb(w_n3907_11[1]),.dout(n16245),.clk(gclk));
	jnot g15952(.din(w_n15647_0[0]),.dout(n16246),.clk(gclk));
	jand g15953(.dina(w_asqrt9_12[2]),.dinb(n16246),.dout(n16247),.clk(gclk));
	jand g15954(.dina(w_n16247_0[1]),.dinb(w_n15652_0[0]),.dout(n16248),.clk(gclk));
	jor g15955(.dina(n16248),.dinb(w_n15651_0[0]),.dout(n16249),.clk(gclk));
	jand g15956(.dina(w_n16247_0[0]),.dinb(w_n15653_0[0]),.dout(n16250),.clk(gclk));
	jnot g15957(.din(n16250),.dout(n16251),.clk(gclk));
	jand g15958(.dina(n16251),.dinb(n16249),.dout(n16252),.clk(gclk));
	jnot g15959(.din(n16252),.dout(n16253),.clk(gclk));
	jor g15960(.dina(w_n16253_0[1]),.dinb(n16245),.dout(n16254),.clk(gclk));
	jand g15961(.dina(w_n16254_0[1]),.dinb(w_n16244_0[1]),.dout(n16255),.clk(gclk));
	jor g15962(.dina(n16255),.dinb(w_n3376_15[0]),.dout(n16256),.clk(gclk));
	jand g15963(.dina(w_n16244_0[0]),.dinb(w_n3376_14[2]),.dout(n16257),.clk(gclk));
	jand g15964(.dina(n16257),.dinb(w_n16254_0[0]),.dout(n16258),.clk(gclk));
	jnot g15965(.din(w_n15655_0[0]),.dout(n16259),.clk(gclk));
	jand g15966(.dina(w_asqrt9_12[1]),.dinb(n16259),.dout(n16260),.clk(gclk));
	jand g15967(.dina(w_n16260_0[1]),.dinb(w_n15662_0[0]),.dout(n16261),.clk(gclk));
	jor g15968(.dina(n16261),.dinb(w_n15660_0[0]),.dout(n16262),.clk(gclk));
	jand g15969(.dina(w_n16260_0[0]),.dinb(w_n15663_0[0]),.dout(n16263),.clk(gclk));
	jnot g15970(.din(n16263),.dout(n16264),.clk(gclk));
	jand g15971(.dina(n16264),.dinb(n16262),.dout(n16265),.clk(gclk));
	jnot g15972(.din(n16265),.dout(n16266),.clk(gclk));
	jor g15973(.dina(w_n16266_0[1]),.dinb(w_n16258_0[1]),.dout(n16267),.clk(gclk));
	jand g15974(.dina(n16267),.dinb(w_n16256_0[1]),.dout(n16268),.clk(gclk));
	jor g15975(.dina(w_n16268_0[1]),.dinb(w_n3371_12[0]),.dout(n16269),.clk(gclk));
	jxor g15976(.dina(w_n15664_0[0]),.dinb(w_n3376_14[1]),.dout(n16270),.clk(gclk));
	jor g15977(.dina(n16270),.dinb(w_n15955_14[2]),.dout(n16271),.clk(gclk));
	jxor g15978(.dina(n16271),.dinb(w_n15675_0[0]),.dout(n16272),.clk(gclk));
	jand g15979(.dina(w_n16268_0[0]),.dinb(w_n3371_11[2]),.dout(n16273),.clk(gclk));
	jor g15980(.dina(w_n16273_0[1]),.dinb(w_n16272_0[1]),.dout(n16274),.clk(gclk));
	jand g15981(.dina(w_n16274_0[2]),.dinb(w_n16269_0[2]),.dout(n16275),.clk(gclk));
	jor g15982(.dina(n16275),.dinb(w_n2875_14[2]),.dout(n16276),.clk(gclk));
	jnot g15983(.din(w_n15680_0[0]),.dout(n16277),.clk(gclk));
	jor g15984(.dina(n16277),.dinb(w_n15678_0[0]),.dout(n16278),.clk(gclk));
	jor g15985(.dina(n16278),.dinb(w_n15955_14[1]),.dout(n16279),.clk(gclk));
	jxor g15986(.dina(n16279),.dinb(w_n15689_0[0]),.dout(n16280),.clk(gclk));
	jand g15987(.dina(w_n16269_0[1]),.dinb(w_n2875_14[1]),.dout(n16281),.clk(gclk));
	jand g15988(.dina(n16281),.dinb(w_n16274_0[1]),.dout(n16282),.clk(gclk));
	jor g15989(.dina(w_n16282_0[1]),.dinb(w_n16280_0[1]),.dout(n16283),.clk(gclk));
	jand g15990(.dina(w_n16283_0[1]),.dinb(w_n16276_0[1]),.dout(n16284),.clk(gclk));
	jor g15991(.dina(w_n16284_0[2]),.dinb(w_n2870_12[1]),.dout(n16285),.clk(gclk));
	jand g15992(.dina(w_n16284_0[1]),.dinb(w_n2870_12[0]),.dout(n16286),.clk(gclk));
	jnot g15993(.din(w_n15692_0[0]),.dout(n16287),.clk(gclk));
	jand g15994(.dina(w_asqrt9_12[0]),.dinb(n16287),.dout(n16288),.clk(gclk));
	jand g15995(.dina(w_n16288_0[1]),.dinb(w_n15697_0[0]),.dout(n16289),.clk(gclk));
	jor g15996(.dina(n16289),.dinb(w_n15696_0[0]),.dout(n16290),.clk(gclk));
	jand g15997(.dina(w_n16288_0[0]),.dinb(w_n15698_0[0]),.dout(n16291),.clk(gclk));
	jnot g15998(.din(n16291),.dout(n16292),.clk(gclk));
	jand g15999(.dina(n16292),.dinb(n16290),.dout(n16293),.clk(gclk));
	jnot g16000(.din(n16293),.dout(n16294),.clk(gclk));
	jor g16001(.dina(w_n16294_0[1]),.dinb(n16286),.dout(n16295),.clk(gclk));
	jand g16002(.dina(w_n16295_0[1]),.dinb(w_n16285_0[1]),.dout(n16296),.clk(gclk));
	jor g16003(.dina(n16296),.dinb(w_n2425_15[1]),.dout(n16297),.clk(gclk));
	jand g16004(.dina(w_n16285_0[0]),.dinb(w_n2425_15[0]),.dout(n16298),.clk(gclk));
	jand g16005(.dina(n16298),.dinb(w_n16295_0[0]),.dout(n16299),.clk(gclk));
	jnot g16006(.din(w_n15700_0[0]),.dout(n16300),.clk(gclk));
	jand g16007(.dina(w_asqrt9_11[2]),.dinb(n16300),.dout(n16301),.clk(gclk));
	jand g16008(.dina(w_n16301_0[1]),.dinb(w_n15707_0[0]),.dout(n16302),.clk(gclk));
	jor g16009(.dina(n16302),.dinb(w_n15705_0[0]),.dout(n16303),.clk(gclk));
	jand g16010(.dina(w_n16301_0[0]),.dinb(w_n15708_0[0]),.dout(n16304),.clk(gclk));
	jnot g16011(.din(n16304),.dout(n16305),.clk(gclk));
	jand g16012(.dina(n16305),.dinb(n16303),.dout(n16306),.clk(gclk));
	jnot g16013(.din(n16306),.dout(n16307),.clk(gclk));
	jor g16014(.dina(w_n16307_0[1]),.dinb(w_n16299_0[1]),.dout(n16308),.clk(gclk));
	jand g16015(.dina(n16308),.dinb(w_n16297_0[1]),.dout(n16309),.clk(gclk));
	jor g16016(.dina(w_n16309_0[1]),.dinb(w_n2420_13[0]),.dout(n16310),.clk(gclk));
	jxor g16017(.dina(w_n15709_0[0]),.dinb(w_n2425_14[2]),.dout(n16311),.clk(gclk));
	jor g16018(.dina(n16311),.dinb(w_n15955_14[0]),.dout(n16312),.clk(gclk));
	jxor g16019(.dina(n16312),.dinb(w_n15720_0[0]),.dout(n16313),.clk(gclk));
	jand g16020(.dina(w_n16309_0[0]),.dinb(w_n2420_12[2]),.dout(n16314),.clk(gclk));
	jor g16021(.dina(w_n16314_0[1]),.dinb(w_n16313_0[1]),.dout(n16315),.clk(gclk));
	jand g16022(.dina(w_n16315_0[2]),.dinb(w_n16310_0[2]),.dout(n16316),.clk(gclk));
	jor g16023(.dina(n16316),.dinb(w_n2010_15[0]),.dout(n16317),.clk(gclk));
	jnot g16024(.din(w_n15725_0[0]),.dout(n16318),.clk(gclk));
	jor g16025(.dina(n16318),.dinb(w_n15723_0[0]),.dout(n16319),.clk(gclk));
	jor g16026(.dina(n16319),.dinb(w_n15955_13[2]),.dout(n16320),.clk(gclk));
	jxor g16027(.dina(n16320),.dinb(w_n15734_0[0]),.dout(n16321),.clk(gclk));
	jand g16028(.dina(w_n16310_0[1]),.dinb(w_n2010_14[2]),.dout(n16322),.clk(gclk));
	jand g16029(.dina(n16322),.dinb(w_n16315_0[1]),.dout(n16323),.clk(gclk));
	jor g16030(.dina(w_n16323_0[1]),.dinb(w_n16321_0[1]),.dout(n16324),.clk(gclk));
	jand g16031(.dina(w_n16324_0[1]),.dinb(w_n16317_0[1]),.dout(n16325),.clk(gclk));
	jor g16032(.dina(w_n16325_0[2]),.dinb(w_n2005_13[1]),.dout(n16326),.clk(gclk));
	jand g16033(.dina(w_n16325_0[1]),.dinb(w_n2005_13[0]),.dout(n16327),.clk(gclk));
	jnot g16034(.din(w_n15737_0[0]),.dout(n16328),.clk(gclk));
	jand g16035(.dina(w_asqrt9_11[1]),.dinb(n16328),.dout(n16329),.clk(gclk));
	jand g16036(.dina(w_n16329_0[1]),.dinb(w_n15742_0[0]),.dout(n16330),.clk(gclk));
	jor g16037(.dina(n16330),.dinb(w_n15741_0[0]),.dout(n16331),.clk(gclk));
	jand g16038(.dina(w_n16329_0[0]),.dinb(w_n15743_0[0]),.dout(n16332),.clk(gclk));
	jnot g16039(.din(n16332),.dout(n16333),.clk(gclk));
	jand g16040(.dina(n16333),.dinb(n16331),.dout(n16334),.clk(gclk));
	jnot g16041(.din(n16334),.dout(n16335),.clk(gclk));
	jor g16042(.dina(w_n16335_0[1]),.dinb(n16327),.dout(n16336),.clk(gclk));
	jand g16043(.dina(w_n16336_0[1]),.dinb(w_n16326_0[1]),.dout(n16337),.clk(gclk));
	jor g16044(.dina(n16337),.dinb(w_n1646_16[0]),.dout(n16338),.clk(gclk));
	jand g16045(.dina(w_n16326_0[0]),.dinb(w_n1646_15[2]),.dout(n16339),.clk(gclk));
	jand g16046(.dina(n16339),.dinb(w_n16336_0[0]),.dout(n16340),.clk(gclk));
	jnot g16047(.din(w_n15745_0[0]),.dout(n16341),.clk(gclk));
	jand g16048(.dina(w_asqrt9_11[0]),.dinb(n16341),.dout(n16342),.clk(gclk));
	jand g16049(.dina(w_n16342_0[1]),.dinb(w_n15752_0[0]),.dout(n16343),.clk(gclk));
	jor g16050(.dina(n16343),.dinb(w_n15750_0[0]),.dout(n16344),.clk(gclk));
	jand g16051(.dina(w_n16342_0[0]),.dinb(w_n15753_0[0]),.dout(n16345),.clk(gclk));
	jnot g16052(.din(n16345),.dout(n16346),.clk(gclk));
	jand g16053(.dina(n16346),.dinb(n16344),.dout(n16347),.clk(gclk));
	jnot g16054(.din(n16347),.dout(n16348),.clk(gclk));
	jor g16055(.dina(w_n16348_0[1]),.dinb(w_n16340_0[1]),.dout(n16349),.clk(gclk));
	jand g16056(.dina(n16349),.dinb(w_n16338_0[1]),.dout(n16350),.clk(gclk));
	jor g16057(.dina(w_n16350_0[1]),.dinb(w_n1641_13[2]),.dout(n16351),.clk(gclk));
	jxor g16058(.dina(w_n15754_0[0]),.dinb(w_n1646_15[1]),.dout(n16352),.clk(gclk));
	jor g16059(.dina(n16352),.dinb(w_n15955_13[1]),.dout(n16353),.clk(gclk));
	jxor g16060(.dina(n16353),.dinb(w_n15765_0[0]),.dout(n16354),.clk(gclk));
	jand g16061(.dina(w_n16350_0[0]),.dinb(w_n1641_13[1]),.dout(n16355),.clk(gclk));
	jor g16062(.dina(w_n16355_0[1]),.dinb(w_n16354_0[1]),.dout(n16356),.clk(gclk));
	jand g16063(.dina(w_n16356_0[2]),.dinb(w_n16351_0[2]),.dout(n16357),.clk(gclk));
	jor g16064(.dina(n16357),.dinb(w_n1317_15[2]),.dout(n16358),.clk(gclk));
	jnot g16065(.din(w_n15770_0[0]),.dout(n16359),.clk(gclk));
	jor g16066(.dina(n16359),.dinb(w_n15768_0[0]),.dout(n16360),.clk(gclk));
	jor g16067(.dina(n16360),.dinb(w_n15955_13[0]),.dout(n16361),.clk(gclk));
	jxor g16068(.dina(n16361),.dinb(w_n15779_0[0]),.dout(n16362),.clk(gclk));
	jand g16069(.dina(w_n16351_0[1]),.dinb(w_n1317_15[1]),.dout(n16363),.clk(gclk));
	jand g16070(.dina(n16363),.dinb(w_n16356_0[1]),.dout(n16364),.clk(gclk));
	jor g16071(.dina(w_n16364_0[1]),.dinb(w_n16362_0[1]),.dout(n16365),.clk(gclk));
	jand g16072(.dina(w_n16365_0[1]),.dinb(w_n16358_0[1]),.dout(n16366),.clk(gclk));
	jor g16073(.dina(w_n16366_0[2]),.dinb(w_n1312_14[0]),.dout(n16367),.clk(gclk));
	jand g16074(.dina(w_n16366_0[1]),.dinb(w_n1312_13[2]),.dout(n16368),.clk(gclk));
	jnot g16075(.din(w_n15782_0[0]),.dout(n16369),.clk(gclk));
	jand g16076(.dina(w_asqrt9_10[2]),.dinb(n16369),.dout(n16370),.clk(gclk));
	jand g16077(.dina(w_n16370_0[1]),.dinb(w_n15787_0[0]),.dout(n16371),.clk(gclk));
	jor g16078(.dina(n16371),.dinb(w_n15786_0[0]),.dout(n16372),.clk(gclk));
	jand g16079(.dina(w_n16370_0[0]),.dinb(w_n15788_0[0]),.dout(n16373),.clk(gclk));
	jnot g16080(.din(n16373),.dout(n16374),.clk(gclk));
	jand g16081(.dina(n16374),.dinb(n16372),.dout(n16375),.clk(gclk));
	jnot g16082(.din(n16375),.dout(n16376),.clk(gclk));
	jor g16083(.dina(w_n16376_0[1]),.dinb(n16368),.dout(n16377),.clk(gclk));
	jand g16084(.dina(w_n16377_0[1]),.dinb(w_n16367_0[1]),.dout(n16378),.clk(gclk));
	jor g16085(.dina(n16378),.dinb(w_n1039_16[1]),.dout(n16379),.clk(gclk));
	jand g16086(.dina(w_n16367_0[0]),.dinb(w_n1039_16[0]),.dout(n16380),.clk(gclk));
	jand g16087(.dina(n16380),.dinb(w_n16377_0[0]),.dout(n16381),.clk(gclk));
	jnot g16088(.din(w_n15790_0[0]),.dout(n16382),.clk(gclk));
	jand g16089(.dina(w_asqrt9_10[1]),.dinb(n16382),.dout(n16383),.clk(gclk));
	jand g16090(.dina(w_n16383_0[1]),.dinb(w_n15797_0[0]),.dout(n16384),.clk(gclk));
	jor g16091(.dina(n16384),.dinb(w_n15795_0[0]),.dout(n16385),.clk(gclk));
	jand g16092(.dina(w_n16383_0[0]),.dinb(w_n15798_0[0]),.dout(n16386),.clk(gclk));
	jnot g16093(.din(n16386),.dout(n16387),.clk(gclk));
	jand g16094(.dina(n16387),.dinb(n16385),.dout(n16388),.clk(gclk));
	jnot g16095(.din(n16388),.dout(n16389),.clk(gclk));
	jor g16096(.dina(w_n16389_0[1]),.dinb(w_n16381_0[1]),.dout(n16390),.clk(gclk));
	jand g16097(.dina(n16390),.dinb(w_n16379_0[1]),.dout(n16391),.clk(gclk));
	jor g16098(.dina(w_n16391_0[1]),.dinb(w_n1034_14[2]),.dout(n16392),.clk(gclk));
	jxor g16099(.dina(w_n15799_0[0]),.dinb(w_n1039_15[2]),.dout(n16393),.clk(gclk));
	jor g16100(.dina(n16393),.dinb(w_n15955_12[2]),.dout(n16394),.clk(gclk));
	jxor g16101(.dina(n16394),.dinb(w_n15810_0[0]),.dout(n16395),.clk(gclk));
	jand g16102(.dina(w_n16391_0[0]),.dinb(w_n1034_14[1]),.dout(n16396),.clk(gclk));
	jor g16103(.dina(w_n16396_0[1]),.dinb(w_n16395_0[1]),.dout(n16397),.clk(gclk));
	jand g16104(.dina(w_n16397_0[2]),.dinb(w_n16392_0[2]),.dout(n16398),.clk(gclk));
	jor g16105(.dina(n16398),.dinb(w_n796_16[0]),.dout(n16399),.clk(gclk));
	jand g16106(.dina(w_n16392_0[1]),.dinb(w_n796_15[2]),.dout(n16400),.clk(gclk));
	jand g16107(.dina(n16400),.dinb(w_n16397_0[1]),.dout(n16401),.clk(gclk));
	jnot g16108(.din(w_n15813_0[0]),.dout(n16402),.clk(gclk));
	jand g16109(.dina(w_asqrt9_10[0]),.dinb(n16402),.dout(n16403),.clk(gclk));
	jand g16110(.dina(w_n16403_0[1]),.dinb(w_n15820_0[0]),.dout(n16404),.clk(gclk));
	jor g16111(.dina(n16404),.dinb(w_n15818_0[0]),.dout(n16405),.clk(gclk));
	jand g16112(.dina(w_n16403_0[0]),.dinb(w_n15821_0[0]),.dout(n16406),.clk(gclk));
	jnot g16113(.din(n16406),.dout(n16407),.clk(gclk));
	jand g16114(.dina(n16407),.dinb(n16405),.dout(n16408),.clk(gclk));
	jnot g16115(.din(n16408),.dout(n16409),.clk(gclk));
	jor g16116(.dina(w_n16409_0[1]),.dinb(w_n16401_0[1]),.dout(n16410),.clk(gclk));
	jand g16117(.dina(n16410),.dinb(w_n16399_0[1]),.dout(n16411),.clk(gclk));
	jor g16118(.dina(w_n16411_0[2]),.dinb(w_n791_15[0]),.dout(n16412),.clk(gclk));
	jand g16119(.dina(w_n16411_0[1]),.dinb(w_n791_14[2]),.dout(n16413),.clk(gclk));
	jor g16120(.dina(n16413),.dinb(w_n15959_0[1]),.dout(n16414),.clk(gclk));
	jand g16121(.dina(w_n16414_0[1]),.dinb(w_n16412_0[1]),.dout(n16415),.clk(gclk));
	jor g16122(.dina(n16415),.dinb(w_n595_17[0]),.dout(n16416),.clk(gclk));
	jnot g16123(.din(w_n15829_0[0]),.dout(n16417),.clk(gclk));
	jor g16124(.dina(n16417),.dinb(w_n15827_0[0]),.dout(n16418),.clk(gclk));
	jor g16125(.dina(n16418),.dinb(w_n15955_12[1]),.dout(n16419),.clk(gclk));
	jxor g16126(.dina(n16419),.dinb(w_n15838_0[0]),.dout(n16420),.clk(gclk));
	jand g16127(.dina(w_n16412_0[0]),.dinb(w_n595_16[2]),.dout(n16421),.clk(gclk));
	jand g16128(.dina(n16421),.dinb(w_n16414_0[0]),.dout(n16422),.clk(gclk));
	jor g16129(.dina(w_n16422_0[1]),.dinb(w_n16420_0[1]),.dout(n16423),.clk(gclk));
	jand g16130(.dina(w_n16423_0[1]),.dinb(w_n16416_0[1]),.dout(n16424),.clk(gclk));
	jor g16131(.dina(w_n16424_0[1]),.dinb(w_n590_15[1]),.dout(n16425),.clk(gclk));
	jxor g16132(.dina(w_n15840_0[0]),.dinb(w_n595_16[1]),.dout(n16426),.clk(gclk));
	jor g16133(.dina(n16426),.dinb(w_n15955_12[0]),.dout(n16427),.clk(gclk));
	jxor g16134(.dina(n16427),.dinb(w_n15851_0[0]),.dout(n16428),.clk(gclk));
	jand g16135(.dina(w_n16424_0[0]),.dinb(w_n590_15[0]),.dout(n16429),.clk(gclk));
	jor g16136(.dina(w_n16429_0[1]),.dinb(w_n16428_0[1]),.dout(n16430),.clk(gclk));
	jand g16137(.dina(w_n16430_0[2]),.dinb(w_n16425_0[2]),.dout(n16431),.clk(gclk));
	jor g16138(.dina(n16431),.dinb(w_n430_16[2]),.dout(n16432),.clk(gclk));
	jnot g16139(.din(w_n15856_0[0]),.dout(n16433),.clk(gclk));
	jor g16140(.dina(n16433),.dinb(w_n15854_0[0]),.dout(n16434),.clk(gclk));
	jor g16141(.dina(n16434),.dinb(w_n15955_11[2]),.dout(n16435),.clk(gclk));
	jxor g16142(.dina(n16435),.dinb(w_n15865_0[0]),.dout(n16436),.clk(gclk));
	jand g16143(.dina(w_n16425_0[1]),.dinb(w_n430_16[1]),.dout(n16437),.clk(gclk));
	jand g16144(.dina(n16437),.dinb(w_n16430_0[1]),.dout(n16438),.clk(gclk));
	jor g16145(.dina(w_n16438_0[1]),.dinb(w_n16436_0[1]),.dout(n16439),.clk(gclk));
	jand g16146(.dina(w_n16439_0[1]),.dinb(w_n16432_0[1]),.dout(n16440),.clk(gclk));
	jor g16147(.dina(w_n16440_0[2]),.dinb(w_n425_15[2]),.dout(n16441),.clk(gclk));
	jand g16148(.dina(w_n16440_0[1]),.dinb(w_n425_15[1]),.dout(n16442),.clk(gclk));
	jnot g16149(.din(w_n15868_0[0]),.dout(n16443),.clk(gclk));
	jand g16150(.dina(w_asqrt9_9[2]),.dinb(n16443),.dout(n16444),.clk(gclk));
	jand g16151(.dina(w_n16444_0[1]),.dinb(w_n15873_0[0]),.dout(n16445),.clk(gclk));
	jor g16152(.dina(n16445),.dinb(w_n15872_0[0]),.dout(n16446),.clk(gclk));
	jand g16153(.dina(w_n16444_0[0]),.dinb(w_n15874_0[0]),.dout(n16447),.clk(gclk));
	jnot g16154(.din(n16447),.dout(n16448),.clk(gclk));
	jand g16155(.dina(n16448),.dinb(n16446),.dout(n16449),.clk(gclk));
	jnot g16156(.din(n16449),.dout(n16450),.clk(gclk));
	jor g16157(.dina(w_n16450_0[1]),.dinb(n16442),.dout(n16451),.clk(gclk));
	jand g16158(.dina(w_n16451_0[1]),.dinb(w_n16441_0[1]),.dout(n16452),.clk(gclk));
	jor g16159(.dina(n16452),.dinb(w_n305_17[1]),.dout(n16453),.clk(gclk));
	jand g16160(.dina(w_n16441_0[0]),.dinb(w_n305_17[0]),.dout(n16454),.clk(gclk));
	jand g16161(.dina(n16454),.dinb(w_n16451_0[0]),.dout(n16455),.clk(gclk));
	jnot g16162(.din(w_n15876_0[0]),.dout(n16456),.clk(gclk));
	jand g16163(.dina(w_asqrt9_9[1]),.dinb(n16456),.dout(n16457),.clk(gclk));
	jand g16164(.dina(w_n16457_0[1]),.dinb(w_n15883_0[0]),.dout(n16458),.clk(gclk));
	jor g16165(.dina(n16458),.dinb(w_n15881_0[0]),.dout(n16459),.clk(gclk));
	jand g16166(.dina(w_n16457_0[0]),.dinb(w_n15884_0[0]),.dout(n16460),.clk(gclk));
	jnot g16167(.din(n16460),.dout(n16461),.clk(gclk));
	jand g16168(.dina(n16461),.dinb(n16459),.dout(n16462),.clk(gclk));
	jnot g16169(.din(n16462),.dout(n16463),.clk(gclk));
	jor g16170(.dina(w_n16463_0[1]),.dinb(w_n16455_0[1]),.dout(n16464),.clk(gclk));
	jand g16171(.dina(n16464),.dinb(w_n16453_0[1]),.dout(n16465),.clk(gclk));
	jor g16172(.dina(w_n16465_0[1]),.dinb(w_n290_16[2]),.dout(n16466),.clk(gclk));
	jxor g16173(.dina(w_n15885_0[0]),.dinb(w_n305_16[2]),.dout(n16467),.clk(gclk));
	jor g16174(.dina(n16467),.dinb(w_n15955_11[1]),.dout(n16468),.clk(gclk));
	jxor g16175(.dina(n16468),.dinb(w_n15896_0[0]),.dout(n16469),.clk(gclk));
	jand g16176(.dina(w_n16465_0[0]),.dinb(w_n290_16[1]),.dout(n16470),.clk(gclk));
	jor g16177(.dina(w_n16470_0[1]),.dinb(w_n16469_0[1]),.dout(n16471),.clk(gclk));
	jand g16178(.dina(w_n16471_0[2]),.dinb(w_n16466_0[2]),.dout(n16472),.clk(gclk));
	jor g16179(.dina(n16472),.dinb(w_n223_17[0]),.dout(n16473),.clk(gclk));
	jnot g16180(.din(w_n15901_0[0]),.dout(n16474),.clk(gclk));
	jor g16181(.dina(n16474),.dinb(w_n15899_0[0]),.dout(n16475),.clk(gclk));
	jor g16182(.dina(n16475),.dinb(w_n15955_11[0]),.dout(n16476),.clk(gclk));
	jxor g16183(.dina(n16476),.dinb(w_n15910_0[0]),.dout(n16477),.clk(gclk));
	jand g16184(.dina(w_n16466_0[1]),.dinb(w_n223_16[2]),.dout(n16478),.clk(gclk));
	jand g16185(.dina(n16478),.dinb(w_n16471_0[1]),.dout(n16479),.clk(gclk));
	jor g16186(.dina(w_n16479_0[1]),.dinb(w_n16477_0[1]),.dout(n16480),.clk(gclk));
	jand g16187(.dina(w_n16480_0[1]),.dinb(w_n16473_0[1]),.dout(n16481),.clk(gclk));
	jor g16188(.dina(w_n16481_0[2]),.dinb(w_n199_19[1]),.dout(n16482),.clk(gclk));
	jand g16189(.dina(w_n16481_0[1]),.dinb(w_n199_19[0]),.dout(n16483),.clk(gclk));
	jnot g16190(.din(w_n15913_0[0]),.dout(n16484),.clk(gclk));
	jand g16191(.dina(w_asqrt9_9[0]),.dinb(n16484),.dout(n16485),.clk(gclk));
	jand g16192(.dina(w_n16485_0[1]),.dinb(w_n15918_0[0]),.dout(n16486),.clk(gclk));
	jor g16193(.dina(n16486),.dinb(w_n15917_0[0]),.dout(n16487),.clk(gclk));
	jand g16194(.dina(w_n16485_0[0]),.dinb(w_n15919_0[0]),.dout(n16488),.clk(gclk));
	jnot g16195(.din(n16488),.dout(n16489),.clk(gclk));
	jand g16196(.dina(n16489),.dinb(n16487),.dout(n16490),.clk(gclk));
	jnot g16197(.din(n16490),.dout(n16491),.clk(gclk));
	jor g16198(.dina(w_n16491_0[1]),.dinb(n16483),.dout(n16492),.clk(gclk));
	jand g16199(.dina(n16492),.dinb(n16482),.dout(n16493),.clk(gclk));
	jnot g16200(.din(w_n15921_0[0]),.dout(n16494),.clk(gclk));
	jand g16201(.dina(w_asqrt9_8[2]),.dinb(n16494),.dout(n16495),.clk(gclk));
	jand g16202(.dina(w_n16495_0[1]),.dinb(w_n15928_0[0]),.dout(n16496),.clk(gclk));
	jor g16203(.dina(n16496),.dinb(w_n15926_0[0]),.dout(n16497),.clk(gclk));
	jand g16204(.dina(w_n16495_0[0]),.dinb(w_n15929_0[0]),.dout(n16498),.clk(gclk));
	jnot g16205(.din(n16498),.dout(n16499),.clk(gclk));
	jand g16206(.dina(n16499),.dinb(n16497),.dout(n16500),.clk(gclk));
	jnot g16207(.din(w_n16500_0[2]),.dout(n16501),.clk(gclk));
	jand g16208(.dina(w_asqrt9_8[1]),.dinb(w_n15943_0[1]),.dout(n16502),.clk(gclk));
	jand g16209(.dina(w_n16502_0[1]),.dinb(w_n15930_1[0]),.dout(n16503),.clk(gclk));
	jor g16210(.dina(n16503),.dinb(w_n15978_0[0]),.dout(n16504),.clk(gclk));
	jor g16211(.dina(n16504),.dinb(w_n16501_0[1]),.dout(n16505),.clk(gclk));
	jor g16212(.dina(n16505),.dinb(w_n16493_0[2]),.dout(n16506),.clk(gclk));
	jand g16213(.dina(n16506),.dinb(w_n194_18[1]),.dout(n16507),.clk(gclk));
	jand g16214(.dina(w_n16501_0[0]),.dinb(w_n16493_0[1]),.dout(n16508),.clk(gclk));
	jor g16215(.dina(w_n16502_0[0]),.dinb(w_n15930_0[2]),.dout(n16509),.clk(gclk));
	jand g16216(.dina(w_n15943_0[0]),.dinb(w_n15930_0[1]),.dout(n16510),.clk(gclk));
	jor g16217(.dina(n16510),.dinb(w_n194_18[0]),.dout(n16511),.clk(gclk));
	jnot g16218(.din(n16511),.dout(n16512),.clk(gclk));
	jand g16219(.dina(n16512),.dinb(n16509),.dout(n16513),.clk(gclk));
	jor g16220(.dina(w_n16513_0[1]),.dinb(w_n16508_0[2]),.dout(n16516),.clk(gclk));
	jor g16221(.dina(n16516),.dinb(w_n16507_0[1]),.dout(asqrt_fa_9),.clk(gclk));
	jxor g16222(.dina(w_n16411_0[0]),.dinb(w_n791_14[1]),.dout(n16518),.clk(gclk));
	jand g16223(.dina(n16518),.dinb(w_asqrt8_31),.dout(n16519),.clk(gclk));
	jxor g16224(.dina(n16519),.dinb(w_n15959_0[0]),.dout(n16520),.clk(gclk));
	jnot g16225(.din(n16520),.dout(n16521),.clk(gclk));
	jand g16226(.dina(w_asqrt8_30[2]),.dinb(w_a16_0[0]),.dout(n16522),.clk(gclk));
	jnot g16227(.din(w_a14_0[1]),.dout(n16523),.clk(gclk));
	jnot g16228(.din(w_a15_0[1]),.dout(n16524),.clk(gclk));
	jand g16229(.dina(w_n15961_1[0]),.dinb(w_n16524_0[1]),.dout(n16525),.clk(gclk));
	jand g16230(.dina(n16525),.dinb(w_n16523_1[1]),.dout(n16526),.clk(gclk));
	jor g16231(.dina(n16526),.dinb(n16522),.dout(n16527),.clk(gclk));
	jand g16232(.dina(w_n16527_0[2]),.dinb(w_asqrt9_8[0]),.dout(n16528),.clk(gclk));
	jand g16233(.dina(w_asqrt8_30[1]),.dinb(w_n15961_0[2]),.dout(n16529),.clk(gclk));
	jxor g16234(.dina(w_n16529_0[1]),.dinb(w_n15962_0[1]),.dout(n16530),.clk(gclk));
	jor g16235(.dina(w_n16527_0[1]),.dinb(w_asqrt9_7[2]),.dout(n16531),.clk(gclk));
	jand g16236(.dina(n16531),.dinb(w_n16530_0[1]),.dout(n16532),.clk(gclk));
	jor g16237(.dina(w_n16532_0[1]),.dinb(w_n16528_0[1]),.dout(n16533),.clk(gclk));
	jand g16238(.dina(n16533),.dinb(w_asqrt10_12[2]),.dout(n16534),.clk(gclk));
	jor g16239(.dina(w_n16528_0[0]),.dinb(w_asqrt10_12[1]),.dout(n16535),.clk(gclk));
	jor g16240(.dina(n16535),.dinb(w_n16532_0[0]),.dout(n16536),.clk(gclk));
	jand g16241(.dina(w_n16529_0[0]),.dinb(w_n15962_0[0]),.dout(n16537),.clk(gclk));
	jnot g16242(.din(w_n16507_0[0]),.dout(n16538),.clk(gclk));
	jnot g16243(.din(w_n16508_0[1]),.dout(n16539),.clk(gclk));
	jnot g16244(.din(w_n16513_0[0]),.dout(n16540),.clk(gclk));
	jand g16245(.dina(n16540),.dinb(w_asqrt9_7[1]),.dout(n16541),.clk(gclk));
	jand g16246(.dina(n16541),.dinb(n16539),.dout(n16542),.clk(gclk));
	jand g16247(.dina(n16542),.dinb(n16538),.dout(n16543),.clk(gclk));
	jor g16248(.dina(n16543),.dinb(n16537),.dout(n16544),.clk(gclk));
	jxor g16249(.dina(n16544),.dinb(w_n15364_0[1]),.dout(n16545),.clk(gclk));
	jand g16250(.dina(w_n16545_0[1]),.dinb(w_n16536_0[1]),.dout(n16546),.clk(gclk));
	jor g16251(.dina(n16546),.dinb(w_n16534_0[1]),.dout(n16547),.clk(gclk));
	jand g16252(.dina(w_n16547_0[2]),.dinb(w_asqrt11_7[2]),.dout(n16548),.clk(gclk));
	jor g16253(.dina(w_n16547_0[1]),.dinb(w_asqrt11_7[1]),.dout(n16549),.clk(gclk));
	jxor g16254(.dina(w_n15966_0[0]),.dinb(w_n15950_5[2]),.dout(n16550),.clk(gclk));
	jand g16255(.dina(n16550),.dinb(w_asqrt8_30[0]),.dout(n16551),.clk(gclk));
	jxor g16256(.dina(n16551),.dinb(w_n15969_0[0]),.dout(n16552),.clk(gclk));
	jnot g16257(.din(w_n16552_0[1]),.dout(n16553),.clk(gclk));
	jand g16258(.dina(n16553),.dinb(n16549),.dout(n16554),.clk(gclk));
	jor g16259(.dina(w_n16554_0[1]),.dinb(w_n16548_0[1]),.dout(n16555),.clk(gclk));
	jand g16260(.dina(n16555),.dinb(w_asqrt12_12[2]),.dout(n16556),.clk(gclk));
	jnot g16261(.din(w_n15975_0[0]),.dout(n16557),.clk(gclk));
	jand g16262(.dina(n16557),.dinb(w_n15973_0[0]),.dout(n16558),.clk(gclk));
	jand g16263(.dina(n16558),.dinb(w_asqrt8_29[2]),.dout(n16559),.clk(gclk));
	jxor g16264(.dina(n16559),.dinb(w_n15983_0[0]),.dout(n16560),.clk(gclk));
	jnot g16265(.din(n16560),.dout(n16561),.clk(gclk));
	jor g16266(.dina(w_n16548_0[0]),.dinb(w_asqrt12_12[1]),.dout(n16562),.clk(gclk));
	jor g16267(.dina(n16562),.dinb(w_n16554_0[0]),.dout(n16563),.clk(gclk));
	jand g16268(.dina(w_n16563_0[1]),.dinb(w_n16561_0[1]),.dout(n16564),.clk(gclk));
	jor g16269(.dina(w_n16564_0[1]),.dinb(w_n16556_0[1]),.dout(n16565),.clk(gclk));
	jand g16270(.dina(w_n16565_0[2]),.dinb(w_asqrt13_8[0]),.dout(n16566),.clk(gclk));
	jor g16271(.dina(w_n16565_0[1]),.dinb(w_asqrt13_7[2]),.dout(n16567),.clk(gclk));
	jnot g16272(.din(w_n15990_0[0]),.dout(n16568),.clk(gclk));
	jxor g16273(.dina(w_n15985_0[0]),.dinb(w_n14816_6[1]),.dout(n16569),.clk(gclk));
	jand g16274(.dina(n16569),.dinb(w_asqrt8_29[1]),.dout(n16570),.clk(gclk));
	jxor g16275(.dina(n16570),.dinb(n16568),.dout(n16571),.clk(gclk));
	jand g16276(.dina(w_n16571_0[1]),.dinb(n16567),.dout(n16572),.clk(gclk));
	jor g16277(.dina(w_n16572_0[1]),.dinb(w_n16566_0[1]),.dout(n16573),.clk(gclk));
	jand g16278(.dina(n16573),.dinb(w_asqrt14_12[2]),.dout(n16574),.clk(gclk));
	jor g16279(.dina(w_n16566_0[0]),.dinb(w_asqrt14_12[1]),.dout(n16575),.clk(gclk));
	jor g16280(.dina(n16575),.dinb(w_n16572_0[0]),.dout(n16576),.clk(gclk));
	jnot g16281(.din(w_n15997_0[0]),.dout(n16577),.clk(gclk));
	jnot g16282(.din(w_n15999_0[0]),.dout(n16578),.clk(gclk));
	jand g16283(.dina(w_asqrt8_29[0]),.dinb(w_n15993_0[0]),.dout(n16579),.clk(gclk));
	jand g16284(.dina(w_n16579_0[1]),.dinb(n16578),.dout(n16580),.clk(gclk));
	jor g16285(.dina(n16580),.dinb(n16577),.dout(n16581),.clk(gclk));
	jnot g16286(.din(w_n16000_0[0]),.dout(n16582),.clk(gclk));
	jand g16287(.dina(w_n16579_0[0]),.dinb(n16582),.dout(n16583),.clk(gclk));
	jnot g16288(.din(n16583),.dout(n16584),.clk(gclk));
	jand g16289(.dina(n16584),.dinb(n16581),.dout(n16585),.clk(gclk));
	jand g16290(.dina(w_n16585_0[1]),.dinb(w_n16576_0[1]),.dout(n16586),.clk(gclk));
	jor g16291(.dina(n16586),.dinb(w_n16574_0[1]),.dout(n16587),.clk(gclk));
	jand g16292(.dina(w_n16587_0[2]),.dinb(w_asqrt15_8[0]),.dout(n16588),.clk(gclk));
	jor g16293(.dina(w_n16587_0[1]),.dinb(w_asqrt15_7[2]),.dout(n16589),.clk(gclk));
	jxor g16294(.dina(w_n16001_0[0]),.dinb(w_n13718_6[1]),.dout(n16590),.clk(gclk));
	jand g16295(.dina(n16590),.dinb(w_asqrt8_28[2]),.dout(n16591),.clk(gclk));
	jxor g16296(.dina(n16591),.dinb(w_n16006_0[0]),.dout(n16592),.clk(gclk));
	jand g16297(.dina(w_n16592_0[1]),.dinb(n16589),.dout(n16593),.clk(gclk));
	jor g16298(.dina(w_n16593_0[1]),.dinb(w_n16588_0[1]),.dout(n16594),.clk(gclk));
	jand g16299(.dina(n16594),.dinb(w_asqrt16_12[2]),.dout(n16595),.clk(gclk));
	jnot g16300(.din(w_n16012_0[0]),.dout(n16596),.clk(gclk));
	jand g16301(.dina(n16596),.dinb(w_n16010_0[0]),.dout(n16597),.clk(gclk));
	jand g16302(.dina(n16597),.dinb(w_asqrt8_28[1]),.dout(n16598),.clk(gclk));
	jxor g16303(.dina(n16598),.dinb(w_n16021_0[0]),.dout(n16599),.clk(gclk));
	jnot g16304(.din(n16599),.dout(n16600),.clk(gclk));
	jor g16305(.dina(w_n16588_0[0]),.dinb(w_asqrt16_12[1]),.dout(n16601),.clk(gclk));
	jor g16306(.dina(n16601),.dinb(w_n16593_0[0]),.dout(n16602),.clk(gclk));
	jand g16307(.dina(w_n16602_0[1]),.dinb(w_n16600_0[1]),.dout(n16603),.clk(gclk));
	jor g16308(.dina(w_n16603_0[1]),.dinb(w_n16595_0[1]),.dout(n16604),.clk(gclk));
	jand g16309(.dina(w_n16604_0[2]),.dinb(w_asqrt17_8[1]),.dout(n16605),.clk(gclk));
	jor g16310(.dina(w_n16604_0[1]),.dinb(w_asqrt17_8[0]),.dout(n16606),.clk(gclk));
	jxor g16311(.dina(w_n16023_0[0]),.dinb(w_n12670_6[2]),.dout(n16607),.clk(gclk));
	jand g16312(.dina(n16607),.dinb(w_asqrt8_28[0]),.dout(n16608),.clk(gclk));
	jxor g16313(.dina(n16608),.dinb(w_n16029_0[0]),.dout(n16609),.clk(gclk));
	jand g16314(.dina(w_n16609_0[1]),.dinb(n16606),.dout(n16610),.clk(gclk));
	jor g16315(.dina(w_n16610_0[1]),.dinb(w_n16605_0[1]),.dout(n16611),.clk(gclk));
	jand g16316(.dina(n16611),.dinb(w_asqrt18_12[2]),.dout(n16612),.clk(gclk));
	jor g16317(.dina(w_n16605_0[0]),.dinb(w_asqrt18_12[1]),.dout(n16613),.clk(gclk));
	jor g16318(.dina(n16613),.dinb(w_n16610_0[0]),.dout(n16614),.clk(gclk));
	jnot g16319(.din(w_n16037_0[0]),.dout(n16615),.clk(gclk));
	jnot g16320(.din(w_n16039_0[0]),.dout(n16616),.clk(gclk));
	jand g16321(.dina(w_asqrt8_27[2]),.dinb(w_n16033_0[0]),.dout(n16617),.clk(gclk));
	jand g16322(.dina(w_n16617_0[1]),.dinb(n16616),.dout(n16618),.clk(gclk));
	jor g16323(.dina(n16618),.dinb(n16615),.dout(n16619),.clk(gclk));
	jnot g16324(.din(w_n16040_0[0]),.dout(n16620),.clk(gclk));
	jand g16325(.dina(w_n16617_0[0]),.dinb(n16620),.dout(n16621),.clk(gclk));
	jnot g16326(.din(n16621),.dout(n16622),.clk(gclk));
	jand g16327(.dina(n16622),.dinb(n16619),.dout(n16623),.clk(gclk));
	jand g16328(.dina(w_n16623_0[1]),.dinb(w_n16614_0[1]),.dout(n16624),.clk(gclk));
	jor g16329(.dina(n16624),.dinb(w_n16612_0[1]),.dout(n16625),.clk(gclk));
	jand g16330(.dina(w_n16625_0[1]),.dinb(w_asqrt19_8[1]),.dout(n16626),.clk(gclk));
	jxor g16331(.dina(w_n16041_0[0]),.dinb(w_n11657_6[2]),.dout(n16627),.clk(gclk));
	jand g16332(.dina(n16627),.dinb(w_asqrt8_27[1]),.dout(n16628),.clk(gclk));
	jxor g16333(.dina(n16628),.dinb(w_n16048_0[0]),.dout(n16629),.clk(gclk));
	jnot g16334(.din(n16629),.dout(n16630),.clk(gclk));
	jor g16335(.dina(w_n16625_0[0]),.dinb(w_asqrt19_8[0]),.dout(n16631),.clk(gclk));
	jand g16336(.dina(w_n16631_0[1]),.dinb(w_n16630_0[1]),.dout(n16632),.clk(gclk));
	jor g16337(.dina(w_n16632_0[2]),.dinb(w_n16626_0[2]),.dout(n16633),.clk(gclk));
	jand g16338(.dina(n16633),.dinb(w_asqrt20_12[2]),.dout(n16634),.clk(gclk));
	jnot g16339(.din(w_n16053_0[0]),.dout(n16635),.clk(gclk));
	jand g16340(.dina(n16635),.dinb(w_n16051_0[0]),.dout(n16636),.clk(gclk));
	jand g16341(.dina(n16636),.dinb(w_asqrt8_27[0]),.dout(n16637),.clk(gclk));
	jxor g16342(.dina(n16637),.dinb(w_n16061_0[0]),.dout(n16638),.clk(gclk));
	jnot g16343(.din(n16638),.dout(n16639),.clk(gclk));
	jor g16344(.dina(w_n16626_0[1]),.dinb(w_asqrt20_12[1]),.dout(n16640),.clk(gclk));
	jor g16345(.dina(n16640),.dinb(w_n16632_0[1]),.dout(n16641),.clk(gclk));
	jand g16346(.dina(w_n16641_0[1]),.dinb(w_n16639_0[1]),.dout(n16642),.clk(gclk));
	jor g16347(.dina(w_n16642_0[1]),.dinb(w_n16634_0[1]),.dout(n16643),.clk(gclk));
	jand g16348(.dina(w_n16643_0[2]),.dinb(w_asqrt21_8[2]),.dout(n16644),.clk(gclk));
	jor g16349(.dina(w_n16643_0[1]),.dinb(w_asqrt21_8[1]),.dout(n16645),.clk(gclk));
	jnot g16350(.din(w_n16067_0[0]),.dout(n16646),.clk(gclk));
	jnot g16351(.din(w_n16068_0[0]),.dout(n16647),.clk(gclk));
	jand g16352(.dina(w_asqrt8_26[2]),.dinb(w_n16064_0[0]),.dout(n16648),.clk(gclk));
	jand g16353(.dina(w_n16648_0[1]),.dinb(n16647),.dout(n16649),.clk(gclk));
	jor g16354(.dina(n16649),.dinb(n16646),.dout(n16650),.clk(gclk));
	jnot g16355(.din(w_n16069_0[0]),.dout(n16651),.clk(gclk));
	jand g16356(.dina(w_n16648_0[0]),.dinb(n16651),.dout(n16652),.clk(gclk));
	jnot g16357(.din(n16652),.dout(n16653),.clk(gclk));
	jand g16358(.dina(n16653),.dinb(n16650),.dout(n16654),.clk(gclk));
	jand g16359(.dina(w_n16654_0[1]),.dinb(n16645),.dout(n16655),.clk(gclk));
	jor g16360(.dina(w_n16655_0[1]),.dinb(w_n16644_0[1]),.dout(n16656),.clk(gclk));
	jand g16361(.dina(n16656),.dinb(w_asqrt22_12[2]),.dout(n16657),.clk(gclk));
	jor g16362(.dina(w_n16644_0[0]),.dinb(w_asqrt22_12[1]),.dout(n16658),.clk(gclk));
	jor g16363(.dina(n16658),.dinb(w_n16655_0[0]),.dout(n16659),.clk(gclk));
	jnot g16364(.din(w_n16075_0[0]),.dout(n16660),.clk(gclk));
	jnot g16365(.din(w_n16077_0[0]),.dout(n16661),.clk(gclk));
	jand g16366(.dina(w_asqrt8_26[1]),.dinb(w_n16071_0[0]),.dout(n16662),.clk(gclk));
	jand g16367(.dina(w_n16662_0[1]),.dinb(n16661),.dout(n16663),.clk(gclk));
	jor g16368(.dina(n16663),.dinb(n16660),.dout(n16664),.clk(gclk));
	jnot g16369(.din(w_n16078_0[0]),.dout(n16665),.clk(gclk));
	jand g16370(.dina(w_n16662_0[0]),.dinb(n16665),.dout(n16666),.clk(gclk));
	jnot g16371(.din(n16666),.dout(n16667),.clk(gclk));
	jand g16372(.dina(n16667),.dinb(n16664),.dout(n16668),.clk(gclk));
	jand g16373(.dina(w_n16668_0[1]),.dinb(w_n16659_0[1]),.dout(n16669),.clk(gclk));
	jor g16374(.dina(n16669),.dinb(w_n16657_0[1]),.dout(n16670),.clk(gclk));
	jand g16375(.dina(w_n16670_0[1]),.dinb(w_asqrt23_8[2]),.dout(n16671),.clk(gclk));
	jxor g16376(.dina(w_n16079_0[0]),.dinb(w_n9769_7[2]),.dout(n16672),.clk(gclk));
	jand g16377(.dina(n16672),.dinb(w_asqrt8_26[0]),.dout(n16673),.clk(gclk));
	jxor g16378(.dina(n16673),.dinb(w_n16089_0[0]),.dout(n16674),.clk(gclk));
	jnot g16379(.din(n16674),.dout(n16675),.clk(gclk));
	jor g16380(.dina(w_n16670_0[0]),.dinb(w_asqrt23_8[1]),.dout(n16676),.clk(gclk));
	jand g16381(.dina(w_n16676_0[1]),.dinb(w_n16675_0[1]),.dout(n16677),.clk(gclk));
	jor g16382(.dina(w_n16677_0[2]),.dinb(w_n16671_0[2]),.dout(n16678),.clk(gclk));
	jand g16383(.dina(n16678),.dinb(w_asqrt24_12[2]),.dout(n16679),.clk(gclk));
	jnot g16384(.din(w_n16094_0[0]),.dout(n16680),.clk(gclk));
	jand g16385(.dina(n16680),.dinb(w_n16092_0[0]),.dout(n16681),.clk(gclk));
	jand g16386(.dina(n16681),.dinb(w_asqrt8_25[2]),.dout(n16682),.clk(gclk));
	jxor g16387(.dina(n16682),.dinb(w_n16102_0[0]),.dout(n16683),.clk(gclk));
	jnot g16388(.din(n16683),.dout(n16684),.clk(gclk));
	jor g16389(.dina(w_n16671_0[1]),.dinb(w_asqrt24_12[1]),.dout(n16685),.clk(gclk));
	jor g16390(.dina(n16685),.dinb(w_n16677_0[1]),.dout(n16686),.clk(gclk));
	jand g16391(.dina(w_n16686_0[1]),.dinb(w_n16684_0[1]),.dout(n16687),.clk(gclk));
	jor g16392(.dina(w_n16687_0[1]),.dinb(w_n16679_0[1]),.dout(n16688),.clk(gclk));
	jand g16393(.dina(w_n16688_0[2]),.dinb(w_asqrt25_9[0]),.dout(n16689),.clk(gclk));
	jor g16394(.dina(w_n16688_0[1]),.dinb(w_asqrt25_8[2]),.dout(n16690),.clk(gclk));
	jnot g16395(.din(w_n16108_0[0]),.dout(n16691),.clk(gclk));
	jnot g16396(.din(w_n16109_0[0]),.dout(n16692),.clk(gclk));
	jand g16397(.dina(w_asqrt8_25[1]),.dinb(w_n16105_0[0]),.dout(n16693),.clk(gclk));
	jand g16398(.dina(w_n16693_0[1]),.dinb(n16692),.dout(n16694),.clk(gclk));
	jor g16399(.dina(n16694),.dinb(n16691),.dout(n16695),.clk(gclk));
	jnot g16400(.din(w_n16110_0[0]),.dout(n16696),.clk(gclk));
	jand g16401(.dina(w_n16693_0[0]),.dinb(n16696),.dout(n16697),.clk(gclk));
	jnot g16402(.din(n16697),.dout(n16698),.clk(gclk));
	jand g16403(.dina(n16698),.dinb(n16695),.dout(n16699),.clk(gclk));
	jand g16404(.dina(w_n16699_0[1]),.dinb(n16690),.dout(n16700),.clk(gclk));
	jor g16405(.dina(w_n16700_0[1]),.dinb(w_n16689_0[1]),.dout(n16701),.clk(gclk));
	jand g16406(.dina(n16701),.dinb(w_asqrt26_12[2]),.dout(n16702),.clk(gclk));
	jor g16407(.dina(w_n16689_0[0]),.dinb(w_asqrt26_12[1]),.dout(n16703),.clk(gclk));
	jor g16408(.dina(n16703),.dinb(w_n16700_0[0]),.dout(n16704),.clk(gclk));
	jnot g16409(.din(w_n16116_0[0]),.dout(n16705),.clk(gclk));
	jnot g16410(.din(w_n16118_0[0]),.dout(n16706),.clk(gclk));
	jand g16411(.dina(w_asqrt8_25[0]),.dinb(w_n16112_0[0]),.dout(n16707),.clk(gclk));
	jand g16412(.dina(w_n16707_0[1]),.dinb(n16706),.dout(n16708),.clk(gclk));
	jor g16413(.dina(n16708),.dinb(n16705),.dout(n16709),.clk(gclk));
	jnot g16414(.din(w_n16119_0[0]),.dout(n16710),.clk(gclk));
	jand g16415(.dina(w_n16707_0[0]),.dinb(n16710),.dout(n16711),.clk(gclk));
	jnot g16416(.din(n16711),.dout(n16712),.clk(gclk));
	jand g16417(.dina(n16712),.dinb(n16709),.dout(n16713),.clk(gclk));
	jand g16418(.dina(w_n16713_0[1]),.dinb(w_n16704_0[1]),.dout(n16714),.clk(gclk));
	jor g16419(.dina(n16714),.dinb(w_n16702_0[1]),.dout(n16715),.clk(gclk));
	jand g16420(.dina(w_n16715_0[1]),.dinb(w_asqrt27_9[0]),.dout(n16716),.clk(gclk));
	jxor g16421(.dina(w_n16120_0[0]),.dinb(w_n8053_8[1]),.dout(n16717),.clk(gclk));
	jand g16422(.dina(n16717),.dinb(w_asqrt8_24[2]),.dout(n16718),.clk(gclk));
	jxor g16423(.dina(n16718),.dinb(w_n16130_0[0]),.dout(n16719),.clk(gclk));
	jnot g16424(.din(n16719),.dout(n16720),.clk(gclk));
	jor g16425(.dina(w_n16715_0[0]),.dinb(w_asqrt27_8[2]),.dout(n16721),.clk(gclk));
	jand g16426(.dina(w_n16721_0[1]),.dinb(w_n16720_0[1]),.dout(n16722),.clk(gclk));
	jor g16427(.dina(w_n16722_0[2]),.dinb(w_n16716_0[2]),.dout(n16723),.clk(gclk));
	jand g16428(.dina(n16723),.dinb(w_asqrt28_12[2]),.dout(n16724),.clk(gclk));
	jnot g16429(.din(w_n16135_0[0]),.dout(n16725),.clk(gclk));
	jand g16430(.dina(n16725),.dinb(w_n16133_0[0]),.dout(n16726),.clk(gclk));
	jand g16431(.dina(n16726),.dinb(w_asqrt8_24[1]),.dout(n16727),.clk(gclk));
	jxor g16432(.dina(n16727),.dinb(w_n16143_0[0]),.dout(n16728),.clk(gclk));
	jnot g16433(.din(n16728),.dout(n16729),.clk(gclk));
	jor g16434(.dina(w_n16716_0[1]),.dinb(w_asqrt28_12[1]),.dout(n16730),.clk(gclk));
	jor g16435(.dina(n16730),.dinb(w_n16722_0[1]),.dout(n16731),.clk(gclk));
	jand g16436(.dina(w_n16731_0[1]),.dinb(w_n16729_0[1]),.dout(n16732),.clk(gclk));
	jor g16437(.dina(w_n16732_0[1]),.dinb(w_n16724_0[1]),.dout(n16733),.clk(gclk));
	jand g16438(.dina(w_n16733_0[2]),.dinb(w_asqrt29_9[1]),.dout(n16734),.clk(gclk));
	jor g16439(.dina(w_n16733_0[1]),.dinb(w_asqrt29_9[0]),.dout(n16735),.clk(gclk));
	jnot g16440(.din(w_n16149_0[0]),.dout(n16736),.clk(gclk));
	jnot g16441(.din(w_n16150_0[0]),.dout(n16737),.clk(gclk));
	jand g16442(.dina(w_asqrt8_24[0]),.dinb(w_n16146_0[0]),.dout(n16738),.clk(gclk));
	jand g16443(.dina(w_n16738_0[1]),.dinb(n16737),.dout(n16739),.clk(gclk));
	jor g16444(.dina(n16739),.dinb(n16736),.dout(n16740),.clk(gclk));
	jnot g16445(.din(w_n16151_0[0]),.dout(n16741),.clk(gclk));
	jand g16446(.dina(w_n16738_0[0]),.dinb(n16741),.dout(n16742),.clk(gclk));
	jnot g16447(.din(n16742),.dout(n16743),.clk(gclk));
	jand g16448(.dina(n16743),.dinb(n16740),.dout(n16744),.clk(gclk));
	jand g16449(.dina(w_n16744_0[1]),.dinb(n16735),.dout(n16745),.clk(gclk));
	jor g16450(.dina(w_n16745_0[1]),.dinb(w_n16734_0[1]),.dout(n16746),.clk(gclk));
	jand g16451(.dina(n16746),.dinb(w_asqrt30_12[2]),.dout(n16747),.clk(gclk));
	jor g16452(.dina(w_n16734_0[0]),.dinb(w_asqrt30_12[1]),.dout(n16748),.clk(gclk));
	jor g16453(.dina(n16748),.dinb(w_n16745_0[0]),.dout(n16749),.clk(gclk));
	jnot g16454(.din(w_n16157_0[0]),.dout(n16750),.clk(gclk));
	jnot g16455(.din(w_n16159_0[0]),.dout(n16751),.clk(gclk));
	jand g16456(.dina(w_asqrt8_23[2]),.dinb(w_n16153_0[0]),.dout(n16752),.clk(gclk));
	jand g16457(.dina(w_n16752_0[1]),.dinb(n16751),.dout(n16753),.clk(gclk));
	jor g16458(.dina(n16753),.dinb(n16750),.dout(n16754),.clk(gclk));
	jnot g16459(.din(w_n16160_0[0]),.dout(n16755),.clk(gclk));
	jand g16460(.dina(w_n16752_0[0]),.dinb(n16755),.dout(n16756),.clk(gclk));
	jnot g16461(.din(n16756),.dout(n16757),.clk(gclk));
	jand g16462(.dina(n16757),.dinb(n16754),.dout(n16758),.clk(gclk));
	jand g16463(.dina(w_n16758_0[1]),.dinb(w_n16749_0[1]),.dout(n16759),.clk(gclk));
	jor g16464(.dina(n16759),.dinb(w_n16747_0[1]),.dout(n16760),.clk(gclk));
	jand g16465(.dina(w_n16760_0[1]),.dinb(w_asqrt31_9[1]),.dout(n16761),.clk(gclk));
	jxor g16466(.dina(w_n16161_0[0]),.dinb(w_n6500_9[1]),.dout(n16762),.clk(gclk));
	jand g16467(.dina(n16762),.dinb(w_asqrt8_23[1]),.dout(n16763),.clk(gclk));
	jxor g16468(.dina(n16763),.dinb(w_n16171_0[0]),.dout(n16764),.clk(gclk));
	jnot g16469(.din(n16764),.dout(n16765),.clk(gclk));
	jor g16470(.dina(w_n16760_0[0]),.dinb(w_asqrt31_9[0]),.dout(n16766),.clk(gclk));
	jand g16471(.dina(w_n16766_0[1]),.dinb(w_n16765_0[1]),.dout(n16767),.clk(gclk));
	jor g16472(.dina(w_n16767_0[2]),.dinb(w_n16761_0[2]),.dout(n16768),.clk(gclk));
	jand g16473(.dina(n16768),.dinb(w_asqrt32_12[2]),.dout(n16769),.clk(gclk));
	jnot g16474(.din(w_n16176_0[0]),.dout(n16770),.clk(gclk));
	jand g16475(.dina(n16770),.dinb(w_n16174_0[0]),.dout(n16771),.clk(gclk));
	jand g16476(.dina(n16771),.dinb(w_asqrt8_23[0]),.dout(n16772),.clk(gclk));
	jxor g16477(.dina(n16772),.dinb(w_n16184_0[0]),.dout(n16773),.clk(gclk));
	jnot g16478(.din(n16773),.dout(n16774),.clk(gclk));
	jor g16479(.dina(w_n16761_0[1]),.dinb(w_asqrt32_12[1]),.dout(n16775),.clk(gclk));
	jor g16480(.dina(n16775),.dinb(w_n16767_0[1]),.dout(n16776),.clk(gclk));
	jand g16481(.dina(w_n16776_0[1]),.dinb(w_n16774_0[1]),.dout(n16777),.clk(gclk));
	jor g16482(.dina(w_n16777_0[1]),.dinb(w_n16769_0[1]),.dout(n16778),.clk(gclk));
	jand g16483(.dina(w_n16778_0[2]),.dinb(w_asqrt33_9[2]),.dout(n16779),.clk(gclk));
	jor g16484(.dina(w_n16778_0[1]),.dinb(w_asqrt33_9[1]),.dout(n16780),.clk(gclk));
	jnot g16485(.din(w_n16190_0[0]),.dout(n16781),.clk(gclk));
	jnot g16486(.din(w_n16191_0[0]),.dout(n16782),.clk(gclk));
	jand g16487(.dina(w_asqrt8_22[2]),.dinb(w_n16187_0[0]),.dout(n16783),.clk(gclk));
	jand g16488(.dina(w_n16783_0[1]),.dinb(n16782),.dout(n16784),.clk(gclk));
	jor g16489(.dina(n16784),.dinb(n16781),.dout(n16785),.clk(gclk));
	jnot g16490(.din(w_n16192_0[0]),.dout(n16786),.clk(gclk));
	jand g16491(.dina(w_n16783_0[0]),.dinb(n16786),.dout(n16787),.clk(gclk));
	jnot g16492(.din(n16787),.dout(n16788),.clk(gclk));
	jand g16493(.dina(n16788),.dinb(n16785),.dout(n16789),.clk(gclk));
	jand g16494(.dina(w_n16789_0[1]),.dinb(n16780),.dout(n16790),.clk(gclk));
	jor g16495(.dina(w_n16790_0[1]),.dinb(w_n16779_0[1]),.dout(n16791),.clk(gclk));
	jand g16496(.dina(n16791),.dinb(w_asqrt34_12[2]),.dout(n16792),.clk(gclk));
	jor g16497(.dina(w_n16779_0[0]),.dinb(w_asqrt34_12[1]),.dout(n16793),.clk(gclk));
	jor g16498(.dina(n16793),.dinb(w_n16790_0[0]),.dout(n16794),.clk(gclk));
	jnot g16499(.din(w_n16198_0[0]),.dout(n16795),.clk(gclk));
	jnot g16500(.din(w_n16200_0[0]),.dout(n16796),.clk(gclk));
	jand g16501(.dina(w_asqrt8_22[1]),.dinb(w_n16194_0[0]),.dout(n16797),.clk(gclk));
	jand g16502(.dina(w_n16797_0[1]),.dinb(n16796),.dout(n16798),.clk(gclk));
	jor g16503(.dina(n16798),.dinb(n16795),.dout(n16799),.clk(gclk));
	jnot g16504(.din(w_n16201_0[0]),.dout(n16800),.clk(gclk));
	jand g16505(.dina(w_n16797_0[0]),.dinb(n16800),.dout(n16801),.clk(gclk));
	jnot g16506(.din(n16801),.dout(n16802),.clk(gclk));
	jand g16507(.dina(n16802),.dinb(n16799),.dout(n16803),.clk(gclk));
	jand g16508(.dina(w_n16803_0[1]),.dinb(w_n16794_0[1]),.dout(n16804),.clk(gclk));
	jor g16509(.dina(n16804),.dinb(w_n16792_0[1]),.dout(n16805),.clk(gclk));
	jand g16510(.dina(w_n16805_0[1]),.dinb(w_asqrt35_9[2]),.dout(n16806),.clk(gclk));
	jxor g16511(.dina(w_n16202_0[0]),.dinb(w_n5116_10[0]),.dout(n16807),.clk(gclk));
	jand g16512(.dina(n16807),.dinb(w_asqrt8_22[0]),.dout(n16808),.clk(gclk));
	jxor g16513(.dina(n16808),.dinb(w_n16212_0[0]),.dout(n16809),.clk(gclk));
	jnot g16514(.din(n16809),.dout(n16810),.clk(gclk));
	jor g16515(.dina(w_n16805_0[0]),.dinb(w_asqrt35_9[1]),.dout(n16811),.clk(gclk));
	jand g16516(.dina(w_n16811_0[1]),.dinb(w_n16810_0[1]),.dout(n16812),.clk(gclk));
	jor g16517(.dina(w_n16812_0[2]),.dinb(w_n16806_0[2]),.dout(n16813),.clk(gclk));
	jand g16518(.dina(n16813),.dinb(w_asqrt36_12[2]),.dout(n16814),.clk(gclk));
	jnot g16519(.din(w_n16217_0[0]),.dout(n16815),.clk(gclk));
	jand g16520(.dina(n16815),.dinb(w_n16215_0[0]),.dout(n16816),.clk(gclk));
	jand g16521(.dina(n16816),.dinb(w_asqrt8_21[2]),.dout(n16817),.clk(gclk));
	jxor g16522(.dina(n16817),.dinb(w_n16225_0[0]),.dout(n16818),.clk(gclk));
	jnot g16523(.din(n16818),.dout(n16819),.clk(gclk));
	jor g16524(.dina(w_n16806_0[1]),.dinb(w_asqrt36_12[1]),.dout(n16820),.clk(gclk));
	jor g16525(.dina(n16820),.dinb(w_n16812_0[1]),.dout(n16821),.clk(gclk));
	jand g16526(.dina(w_n16821_0[1]),.dinb(w_n16819_0[1]),.dout(n16822),.clk(gclk));
	jor g16527(.dina(w_n16822_0[1]),.dinb(w_n16814_0[1]),.dout(n16823),.clk(gclk));
	jand g16528(.dina(w_n16823_0[2]),.dinb(w_asqrt37_10[0]),.dout(n16824),.clk(gclk));
	jor g16529(.dina(w_n16823_0[1]),.dinb(w_asqrt37_9[2]),.dout(n16825),.clk(gclk));
	jnot g16530(.din(w_n16231_0[0]),.dout(n16826),.clk(gclk));
	jnot g16531(.din(w_n16232_0[0]),.dout(n16827),.clk(gclk));
	jand g16532(.dina(w_asqrt8_21[1]),.dinb(w_n16228_0[0]),.dout(n16828),.clk(gclk));
	jand g16533(.dina(w_n16828_0[1]),.dinb(n16827),.dout(n16829),.clk(gclk));
	jor g16534(.dina(n16829),.dinb(n16826),.dout(n16830),.clk(gclk));
	jnot g16535(.din(w_n16233_0[0]),.dout(n16831),.clk(gclk));
	jand g16536(.dina(w_n16828_0[0]),.dinb(n16831),.dout(n16832),.clk(gclk));
	jnot g16537(.din(n16832),.dout(n16833),.clk(gclk));
	jand g16538(.dina(n16833),.dinb(n16830),.dout(n16834),.clk(gclk));
	jand g16539(.dina(w_n16834_0[1]),.dinb(n16825),.dout(n16835),.clk(gclk));
	jor g16540(.dina(w_n16835_0[1]),.dinb(w_n16824_0[1]),.dout(n16836),.clk(gclk));
	jand g16541(.dina(n16836),.dinb(w_asqrt38_12[2]),.dout(n16837),.clk(gclk));
	jor g16542(.dina(w_n16824_0[0]),.dinb(w_asqrt38_12[1]),.dout(n16838),.clk(gclk));
	jor g16543(.dina(n16838),.dinb(w_n16835_0[0]),.dout(n16839),.clk(gclk));
	jnot g16544(.din(w_n16239_0[0]),.dout(n16840),.clk(gclk));
	jnot g16545(.din(w_n16241_0[0]),.dout(n16841),.clk(gclk));
	jand g16546(.dina(w_asqrt8_21[0]),.dinb(w_n16235_0[0]),.dout(n16842),.clk(gclk));
	jand g16547(.dina(w_n16842_0[1]),.dinb(n16841),.dout(n16843),.clk(gclk));
	jor g16548(.dina(n16843),.dinb(n16840),.dout(n16844),.clk(gclk));
	jnot g16549(.din(w_n16242_0[0]),.dout(n16845),.clk(gclk));
	jand g16550(.dina(w_n16842_0[0]),.dinb(n16845),.dout(n16846),.clk(gclk));
	jnot g16551(.din(n16846),.dout(n16847),.clk(gclk));
	jand g16552(.dina(n16847),.dinb(n16844),.dout(n16848),.clk(gclk));
	jand g16553(.dina(w_n16848_0[1]),.dinb(w_n16839_0[1]),.dout(n16849),.clk(gclk));
	jor g16554(.dina(n16849),.dinb(w_n16837_0[1]),.dout(n16850),.clk(gclk));
	jand g16555(.dina(w_n16850_0[1]),.dinb(w_asqrt39_10[0]),.dout(n16851),.clk(gclk));
	jxor g16556(.dina(w_n16243_0[0]),.dinb(w_n3907_11[0]),.dout(n16852),.clk(gclk));
	jand g16557(.dina(n16852),.dinb(w_asqrt8_20[2]),.dout(n16853),.clk(gclk));
	jxor g16558(.dina(n16853),.dinb(w_n16253_0[0]),.dout(n16854),.clk(gclk));
	jnot g16559(.din(n16854),.dout(n16855),.clk(gclk));
	jor g16560(.dina(w_n16850_0[0]),.dinb(w_asqrt39_9[2]),.dout(n16856),.clk(gclk));
	jand g16561(.dina(w_n16856_0[1]),.dinb(w_n16855_0[1]),.dout(n16857),.clk(gclk));
	jor g16562(.dina(w_n16857_0[2]),.dinb(w_n16851_0[2]),.dout(n16858),.clk(gclk));
	jand g16563(.dina(n16858),.dinb(w_asqrt40_12[2]),.dout(n16859),.clk(gclk));
	jnot g16564(.din(w_n16258_0[0]),.dout(n16860),.clk(gclk));
	jand g16565(.dina(n16860),.dinb(w_n16256_0[0]),.dout(n16861),.clk(gclk));
	jand g16566(.dina(n16861),.dinb(w_asqrt8_20[1]),.dout(n16862),.clk(gclk));
	jxor g16567(.dina(n16862),.dinb(w_n16266_0[0]),.dout(n16863),.clk(gclk));
	jnot g16568(.din(n16863),.dout(n16864),.clk(gclk));
	jor g16569(.dina(w_n16851_0[1]),.dinb(w_asqrt40_12[1]),.dout(n16865),.clk(gclk));
	jor g16570(.dina(n16865),.dinb(w_n16857_0[1]),.dout(n16866),.clk(gclk));
	jand g16571(.dina(w_n16866_0[1]),.dinb(w_n16864_0[1]),.dout(n16867),.clk(gclk));
	jor g16572(.dina(w_n16867_0[1]),.dinb(w_n16859_0[1]),.dout(n16868),.clk(gclk));
	jand g16573(.dina(w_n16868_0[2]),.dinb(w_asqrt41_10[1]),.dout(n16869),.clk(gclk));
	jor g16574(.dina(w_n16868_0[1]),.dinb(w_asqrt41_10[0]),.dout(n16870),.clk(gclk));
	jnot g16575(.din(w_n16272_0[0]),.dout(n16871),.clk(gclk));
	jnot g16576(.din(w_n16273_0[0]),.dout(n16872),.clk(gclk));
	jand g16577(.dina(w_asqrt8_20[0]),.dinb(w_n16269_0[0]),.dout(n16873),.clk(gclk));
	jand g16578(.dina(w_n16873_0[1]),.dinb(n16872),.dout(n16874),.clk(gclk));
	jor g16579(.dina(n16874),.dinb(n16871),.dout(n16875),.clk(gclk));
	jnot g16580(.din(w_n16274_0[0]),.dout(n16876),.clk(gclk));
	jand g16581(.dina(w_n16873_0[0]),.dinb(n16876),.dout(n16877),.clk(gclk));
	jnot g16582(.din(n16877),.dout(n16878),.clk(gclk));
	jand g16583(.dina(n16878),.dinb(n16875),.dout(n16879),.clk(gclk));
	jand g16584(.dina(w_n16879_0[1]),.dinb(n16870),.dout(n16880),.clk(gclk));
	jor g16585(.dina(w_n16880_0[1]),.dinb(w_n16869_0[1]),.dout(n16881),.clk(gclk));
	jand g16586(.dina(n16881),.dinb(w_asqrt42_12[2]),.dout(n16882),.clk(gclk));
	jor g16587(.dina(w_n16869_0[0]),.dinb(w_asqrt42_12[1]),.dout(n16883),.clk(gclk));
	jor g16588(.dina(n16883),.dinb(w_n16880_0[0]),.dout(n16884),.clk(gclk));
	jnot g16589(.din(w_n16280_0[0]),.dout(n16885),.clk(gclk));
	jnot g16590(.din(w_n16282_0[0]),.dout(n16886),.clk(gclk));
	jand g16591(.dina(w_asqrt8_19[2]),.dinb(w_n16276_0[0]),.dout(n16887),.clk(gclk));
	jand g16592(.dina(w_n16887_0[1]),.dinb(n16886),.dout(n16888),.clk(gclk));
	jor g16593(.dina(n16888),.dinb(n16885),.dout(n16889),.clk(gclk));
	jnot g16594(.din(w_n16283_0[0]),.dout(n16890),.clk(gclk));
	jand g16595(.dina(w_n16887_0[0]),.dinb(n16890),.dout(n16891),.clk(gclk));
	jnot g16596(.din(n16891),.dout(n16892),.clk(gclk));
	jand g16597(.dina(n16892),.dinb(n16889),.dout(n16893),.clk(gclk));
	jand g16598(.dina(w_n16893_0[1]),.dinb(w_n16884_0[1]),.dout(n16894),.clk(gclk));
	jor g16599(.dina(n16894),.dinb(w_n16882_0[1]),.dout(n16895),.clk(gclk));
	jand g16600(.dina(w_n16895_0[1]),.dinb(w_asqrt43_10[1]),.dout(n16896),.clk(gclk));
	jxor g16601(.dina(w_n16284_0[0]),.dinb(w_n2870_11[2]),.dout(n16897),.clk(gclk));
	jand g16602(.dina(n16897),.dinb(w_asqrt8_19[1]),.dout(n16898),.clk(gclk));
	jxor g16603(.dina(n16898),.dinb(w_n16294_0[0]),.dout(n16899),.clk(gclk));
	jnot g16604(.din(n16899),.dout(n16900),.clk(gclk));
	jor g16605(.dina(w_n16895_0[0]),.dinb(w_asqrt43_10[0]),.dout(n16901),.clk(gclk));
	jand g16606(.dina(w_n16901_0[1]),.dinb(w_n16900_0[1]),.dout(n16902),.clk(gclk));
	jor g16607(.dina(w_n16902_0[2]),.dinb(w_n16896_0[2]),.dout(n16903),.clk(gclk));
	jand g16608(.dina(n16903),.dinb(w_asqrt44_12[2]),.dout(n16904),.clk(gclk));
	jnot g16609(.din(w_n16299_0[0]),.dout(n16905),.clk(gclk));
	jand g16610(.dina(n16905),.dinb(w_n16297_0[0]),.dout(n16906),.clk(gclk));
	jand g16611(.dina(n16906),.dinb(w_asqrt8_19[0]),.dout(n16907),.clk(gclk));
	jxor g16612(.dina(n16907),.dinb(w_n16307_0[0]),.dout(n16908),.clk(gclk));
	jnot g16613(.din(n16908),.dout(n16909),.clk(gclk));
	jor g16614(.dina(w_n16896_0[1]),.dinb(w_asqrt44_12[1]),.dout(n16910),.clk(gclk));
	jor g16615(.dina(n16910),.dinb(w_n16902_0[1]),.dout(n16911),.clk(gclk));
	jand g16616(.dina(w_n16911_0[1]),.dinb(w_n16909_0[1]),.dout(n16912),.clk(gclk));
	jor g16617(.dina(w_n16912_0[1]),.dinb(w_n16904_0[1]),.dout(n16913),.clk(gclk));
	jand g16618(.dina(w_n16913_0[2]),.dinb(w_asqrt45_10[2]),.dout(n16914),.clk(gclk));
	jor g16619(.dina(w_n16913_0[1]),.dinb(w_asqrt45_10[1]),.dout(n16915),.clk(gclk));
	jnot g16620(.din(w_n16313_0[0]),.dout(n16916),.clk(gclk));
	jnot g16621(.din(w_n16314_0[0]),.dout(n16917),.clk(gclk));
	jand g16622(.dina(w_asqrt8_18[2]),.dinb(w_n16310_0[0]),.dout(n16918),.clk(gclk));
	jand g16623(.dina(w_n16918_0[1]),.dinb(n16917),.dout(n16919),.clk(gclk));
	jor g16624(.dina(n16919),.dinb(n16916),.dout(n16920),.clk(gclk));
	jnot g16625(.din(w_n16315_0[0]),.dout(n16921),.clk(gclk));
	jand g16626(.dina(w_n16918_0[0]),.dinb(n16921),.dout(n16922),.clk(gclk));
	jnot g16627(.din(n16922),.dout(n16923),.clk(gclk));
	jand g16628(.dina(n16923),.dinb(n16920),.dout(n16924),.clk(gclk));
	jand g16629(.dina(w_n16924_0[1]),.dinb(n16915),.dout(n16925),.clk(gclk));
	jor g16630(.dina(w_n16925_0[1]),.dinb(w_n16914_0[1]),.dout(n16926),.clk(gclk));
	jand g16631(.dina(n16926),.dinb(w_asqrt46_12[2]),.dout(n16927),.clk(gclk));
	jor g16632(.dina(w_n16914_0[0]),.dinb(w_asqrt46_12[1]),.dout(n16928),.clk(gclk));
	jor g16633(.dina(n16928),.dinb(w_n16925_0[0]),.dout(n16929),.clk(gclk));
	jnot g16634(.din(w_n16321_0[0]),.dout(n16930),.clk(gclk));
	jnot g16635(.din(w_n16323_0[0]),.dout(n16931),.clk(gclk));
	jand g16636(.dina(w_asqrt8_18[1]),.dinb(w_n16317_0[0]),.dout(n16932),.clk(gclk));
	jand g16637(.dina(w_n16932_0[1]),.dinb(n16931),.dout(n16933),.clk(gclk));
	jor g16638(.dina(n16933),.dinb(n16930),.dout(n16934),.clk(gclk));
	jnot g16639(.din(w_n16324_0[0]),.dout(n16935),.clk(gclk));
	jand g16640(.dina(w_n16932_0[0]),.dinb(n16935),.dout(n16936),.clk(gclk));
	jnot g16641(.din(n16936),.dout(n16937),.clk(gclk));
	jand g16642(.dina(n16937),.dinb(n16934),.dout(n16938),.clk(gclk));
	jand g16643(.dina(w_n16938_0[1]),.dinb(w_n16929_0[1]),.dout(n16939),.clk(gclk));
	jor g16644(.dina(n16939),.dinb(w_n16927_0[1]),.dout(n16940),.clk(gclk));
	jand g16645(.dina(w_n16940_0[1]),.dinb(w_asqrt47_10[2]),.dout(n16941),.clk(gclk));
	jxor g16646(.dina(w_n16325_0[0]),.dinb(w_n2005_12[2]),.dout(n16942),.clk(gclk));
	jand g16647(.dina(n16942),.dinb(w_asqrt8_18[0]),.dout(n16943),.clk(gclk));
	jxor g16648(.dina(n16943),.dinb(w_n16335_0[0]),.dout(n16944),.clk(gclk));
	jnot g16649(.din(n16944),.dout(n16945),.clk(gclk));
	jor g16650(.dina(w_n16940_0[0]),.dinb(w_asqrt47_10[1]),.dout(n16946),.clk(gclk));
	jand g16651(.dina(w_n16946_0[1]),.dinb(w_n16945_0[1]),.dout(n16947),.clk(gclk));
	jor g16652(.dina(w_n16947_0[2]),.dinb(w_n16941_0[2]),.dout(n16948),.clk(gclk));
	jand g16653(.dina(n16948),.dinb(w_asqrt48_12[2]),.dout(n16949),.clk(gclk));
	jnot g16654(.din(w_n16340_0[0]),.dout(n16950),.clk(gclk));
	jand g16655(.dina(n16950),.dinb(w_n16338_0[0]),.dout(n16951),.clk(gclk));
	jand g16656(.dina(n16951),.dinb(w_asqrt8_17[2]),.dout(n16952),.clk(gclk));
	jxor g16657(.dina(n16952),.dinb(w_n16348_0[0]),.dout(n16953),.clk(gclk));
	jnot g16658(.din(n16953),.dout(n16954),.clk(gclk));
	jor g16659(.dina(w_n16941_0[1]),.dinb(w_asqrt48_12[1]),.dout(n16955),.clk(gclk));
	jor g16660(.dina(n16955),.dinb(w_n16947_0[1]),.dout(n16956),.clk(gclk));
	jand g16661(.dina(w_n16956_0[1]),.dinb(w_n16954_0[1]),.dout(n16957),.clk(gclk));
	jor g16662(.dina(w_n16957_0[1]),.dinb(w_n16949_0[1]),.dout(n16958),.clk(gclk));
	jand g16663(.dina(w_n16958_0[2]),.dinb(w_asqrt49_11[0]),.dout(n16959),.clk(gclk));
	jor g16664(.dina(w_n16958_0[1]),.dinb(w_asqrt49_10[2]),.dout(n16960),.clk(gclk));
	jnot g16665(.din(w_n16354_0[0]),.dout(n16961),.clk(gclk));
	jnot g16666(.din(w_n16355_0[0]),.dout(n16962),.clk(gclk));
	jand g16667(.dina(w_asqrt8_17[1]),.dinb(w_n16351_0[0]),.dout(n16963),.clk(gclk));
	jand g16668(.dina(w_n16963_0[1]),.dinb(n16962),.dout(n16964),.clk(gclk));
	jor g16669(.dina(n16964),.dinb(n16961),.dout(n16965),.clk(gclk));
	jnot g16670(.din(w_n16356_0[0]),.dout(n16966),.clk(gclk));
	jand g16671(.dina(w_n16963_0[0]),.dinb(n16966),.dout(n16967),.clk(gclk));
	jnot g16672(.din(n16967),.dout(n16968),.clk(gclk));
	jand g16673(.dina(n16968),.dinb(n16965),.dout(n16969),.clk(gclk));
	jand g16674(.dina(w_n16969_0[1]),.dinb(n16960),.dout(n16970),.clk(gclk));
	jor g16675(.dina(w_n16970_0[1]),.dinb(w_n16959_0[1]),.dout(n16971),.clk(gclk));
	jand g16676(.dina(n16971),.dinb(w_asqrt50_12[2]),.dout(n16972),.clk(gclk));
	jor g16677(.dina(w_n16959_0[0]),.dinb(w_asqrt50_12[1]),.dout(n16973),.clk(gclk));
	jor g16678(.dina(n16973),.dinb(w_n16970_0[0]),.dout(n16974),.clk(gclk));
	jnot g16679(.din(w_n16362_0[0]),.dout(n16975),.clk(gclk));
	jnot g16680(.din(w_n16364_0[0]),.dout(n16976),.clk(gclk));
	jand g16681(.dina(w_asqrt8_17[0]),.dinb(w_n16358_0[0]),.dout(n16977),.clk(gclk));
	jand g16682(.dina(w_n16977_0[1]),.dinb(n16976),.dout(n16978),.clk(gclk));
	jor g16683(.dina(n16978),.dinb(n16975),.dout(n16979),.clk(gclk));
	jnot g16684(.din(w_n16365_0[0]),.dout(n16980),.clk(gclk));
	jand g16685(.dina(w_n16977_0[0]),.dinb(n16980),.dout(n16981),.clk(gclk));
	jnot g16686(.din(n16981),.dout(n16982),.clk(gclk));
	jand g16687(.dina(n16982),.dinb(n16979),.dout(n16983),.clk(gclk));
	jand g16688(.dina(w_n16983_0[1]),.dinb(w_n16974_0[1]),.dout(n16984),.clk(gclk));
	jor g16689(.dina(n16984),.dinb(w_n16972_0[1]),.dout(n16985),.clk(gclk));
	jand g16690(.dina(w_n16985_0[1]),.dinb(w_asqrt51_11[0]),.dout(n16986),.clk(gclk));
	jxor g16691(.dina(w_n16366_0[0]),.dinb(w_n1312_13[1]),.dout(n16987),.clk(gclk));
	jand g16692(.dina(n16987),.dinb(w_asqrt8_16[2]),.dout(n16988),.clk(gclk));
	jxor g16693(.dina(n16988),.dinb(w_n16376_0[0]),.dout(n16989),.clk(gclk));
	jnot g16694(.din(n16989),.dout(n16990),.clk(gclk));
	jor g16695(.dina(w_n16985_0[0]),.dinb(w_asqrt51_10[2]),.dout(n16991),.clk(gclk));
	jand g16696(.dina(w_n16991_0[1]),.dinb(w_n16990_0[1]),.dout(n16992),.clk(gclk));
	jor g16697(.dina(w_n16992_0[2]),.dinb(w_n16986_0[2]),.dout(n16993),.clk(gclk));
	jand g16698(.dina(n16993),.dinb(w_asqrt52_12[2]),.dout(n16994),.clk(gclk));
	jnot g16699(.din(w_n16381_0[0]),.dout(n16995),.clk(gclk));
	jand g16700(.dina(n16995),.dinb(w_n16379_0[0]),.dout(n16996),.clk(gclk));
	jand g16701(.dina(n16996),.dinb(w_asqrt8_16[1]),.dout(n16997),.clk(gclk));
	jxor g16702(.dina(n16997),.dinb(w_n16389_0[0]),.dout(n16998),.clk(gclk));
	jnot g16703(.din(n16998),.dout(n16999),.clk(gclk));
	jor g16704(.dina(w_n16986_0[1]),.dinb(w_asqrt52_12[1]),.dout(n17000),.clk(gclk));
	jor g16705(.dina(n17000),.dinb(w_n16992_0[1]),.dout(n17001),.clk(gclk));
	jand g16706(.dina(w_n17001_0[1]),.dinb(w_n16999_0[1]),.dout(n17002),.clk(gclk));
	jor g16707(.dina(w_n17002_0[1]),.dinb(w_n16994_0[1]),.dout(n17003),.clk(gclk));
	jand g16708(.dina(w_n17003_0[2]),.dinb(w_asqrt53_11[1]),.dout(n17004),.clk(gclk));
	jor g16709(.dina(w_n17003_0[1]),.dinb(w_asqrt53_11[0]),.dout(n17005),.clk(gclk));
	jnot g16710(.din(w_n16395_0[0]),.dout(n17006),.clk(gclk));
	jnot g16711(.din(w_n16396_0[0]),.dout(n17007),.clk(gclk));
	jand g16712(.dina(w_asqrt8_16[0]),.dinb(w_n16392_0[0]),.dout(n17008),.clk(gclk));
	jand g16713(.dina(w_n17008_0[1]),.dinb(n17007),.dout(n17009),.clk(gclk));
	jor g16714(.dina(n17009),.dinb(n17006),.dout(n17010),.clk(gclk));
	jnot g16715(.din(w_n16397_0[0]),.dout(n17011),.clk(gclk));
	jand g16716(.dina(w_n17008_0[0]),.dinb(n17011),.dout(n17012),.clk(gclk));
	jnot g16717(.din(n17012),.dout(n17013),.clk(gclk));
	jand g16718(.dina(n17013),.dinb(n17010),.dout(n17014),.clk(gclk));
	jand g16719(.dina(w_n17014_0[1]),.dinb(n17005),.dout(n17015),.clk(gclk));
	jor g16720(.dina(w_n17015_0[1]),.dinb(w_n17004_0[1]),.dout(n17016),.clk(gclk));
	jand g16721(.dina(n17016),.dinb(w_asqrt54_12[2]),.dout(n17017),.clk(gclk));
	jnot g16722(.din(w_n16401_0[0]),.dout(n17018),.clk(gclk));
	jand g16723(.dina(n17018),.dinb(w_n16399_0[0]),.dout(n17019),.clk(gclk));
	jand g16724(.dina(n17019),.dinb(w_asqrt8_15[2]),.dout(n17020),.clk(gclk));
	jxor g16725(.dina(n17020),.dinb(w_n16409_0[0]),.dout(n17021),.clk(gclk));
	jnot g16726(.din(n17021),.dout(n17022),.clk(gclk));
	jor g16727(.dina(w_n17004_0[0]),.dinb(w_asqrt54_12[1]),.dout(n17023),.clk(gclk));
	jor g16728(.dina(n17023),.dinb(w_n17015_0[0]),.dout(n17024),.clk(gclk));
	jand g16729(.dina(w_n17024_0[1]),.dinb(w_n17022_0[1]),.dout(n17025),.clk(gclk));
	jor g16730(.dina(w_n17025_0[1]),.dinb(w_n17017_0[1]),.dout(n17026),.clk(gclk));
	jand g16731(.dina(w_n17026_0[2]),.dinb(w_asqrt55_11[2]),.dout(n17027),.clk(gclk));
	jor g16732(.dina(w_n17026_0[1]),.dinb(w_asqrt55_11[1]),.dout(n17028),.clk(gclk));
	jand g16733(.dina(n17028),.dinb(w_n16521_0[1]),.dout(n17029),.clk(gclk));
	jor g16734(.dina(w_n17029_0[1]),.dinb(w_n17027_0[1]),.dout(n17030),.clk(gclk));
	jand g16735(.dina(n17030),.dinb(w_asqrt56_12[2]),.dout(n17031),.clk(gclk));
	jor g16736(.dina(w_n17027_0[0]),.dinb(w_asqrt56_12[1]),.dout(n17032),.clk(gclk));
	jor g16737(.dina(n17032),.dinb(w_n17029_0[0]),.dout(n17033),.clk(gclk));
	jnot g16738(.din(w_n16420_0[0]),.dout(n17034),.clk(gclk));
	jnot g16739(.din(w_n16422_0[0]),.dout(n17035),.clk(gclk));
	jand g16740(.dina(w_asqrt8_15[1]),.dinb(w_n16416_0[0]),.dout(n17036),.clk(gclk));
	jand g16741(.dina(w_n17036_0[1]),.dinb(n17035),.dout(n17037),.clk(gclk));
	jor g16742(.dina(n17037),.dinb(n17034),.dout(n17038),.clk(gclk));
	jnot g16743(.din(w_n16423_0[0]),.dout(n17039),.clk(gclk));
	jand g16744(.dina(w_n17036_0[0]),.dinb(n17039),.dout(n17040),.clk(gclk));
	jnot g16745(.din(n17040),.dout(n17041),.clk(gclk));
	jand g16746(.dina(n17041),.dinb(n17038),.dout(n17042),.clk(gclk));
	jand g16747(.dina(w_n17042_0[1]),.dinb(w_n17033_0[1]),.dout(n17043),.clk(gclk));
	jor g16748(.dina(n17043),.dinb(w_n17031_0[1]),.dout(n17044),.clk(gclk));
	jand g16749(.dina(w_n17044_0[2]),.dinb(w_asqrt57_12[0]),.dout(n17045),.clk(gclk));
	jor g16750(.dina(w_n17044_0[1]),.dinb(w_asqrt57_11[2]),.dout(n17046),.clk(gclk));
	jnot g16751(.din(w_n16428_0[0]),.dout(n17047),.clk(gclk));
	jnot g16752(.din(w_n16429_0[0]),.dout(n17048),.clk(gclk));
	jand g16753(.dina(w_asqrt8_15[0]),.dinb(w_n16425_0[0]),.dout(n17049),.clk(gclk));
	jand g16754(.dina(w_n17049_0[1]),.dinb(n17048),.dout(n17050),.clk(gclk));
	jor g16755(.dina(n17050),.dinb(n17047),.dout(n17051),.clk(gclk));
	jnot g16756(.din(w_n16430_0[0]),.dout(n17052),.clk(gclk));
	jand g16757(.dina(w_n17049_0[0]),.dinb(n17052),.dout(n17053),.clk(gclk));
	jnot g16758(.din(n17053),.dout(n17054),.clk(gclk));
	jand g16759(.dina(n17054),.dinb(n17051),.dout(n17055),.clk(gclk));
	jand g16760(.dina(w_n17055_0[1]),.dinb(n17046),.dout(n17056),.clk(gclk));
	jor g16761(.dina(w_n17056_0[1]),.dinb(w_n17045_0[1]),.dout(n17057),.clk(gclk));
	jand g16762(.dina(n17057),.dinb(w_asqrt58_12[2]),.dout(n17058),.clk(gclk));
	jor g16763(.dina(w_n17045_0[0]),.dinb(w_asqrt58_12[1]),.dout(n17059),.clk(gclk));
	jor g16764(.dina(n17059),.dinb(w_n17056_0[0]),.dout(n17060),.clk(gclk));
	jnot g16765(.din(w_n16436_0[0]),.dout(n17061),.clk(gclk));
	jnot g16766(.din(w_n16438_0[0]),.dout(n17062),.clk(gclk));
	jand g16767(.dina(w_asqrt8_14[2]),.dinb(w_n16432_0[0]),.dout(n17063),.clk(gclk));
	jand g16768(.dina(w_n17063_0[1]),.dinb(n17062),.dout(n17064),.clk(gclk));
	jor g16769(.dina(n17064),.dinb(n17061),.dout(n17065),.clk(gclk));
	jnot g16770(.din(w_n16439_0[0]),.dout(n17066),.clk(gclk));
	jand g16771(.dina(w_n17063_0[0]),.dinb(n17066),.dout(n17067),.clk(gclk));
	jnot g16772(.din(n17067),.dout(n17068),.clk(gclk));
	jand g16773(.dina(n17068),.dinb(n17065),.dout(n17069),.clk(gclk));
	jand g16774(.dina(w_n17069_0[1]),.dinb(w_n17060_0[1]),.dout(n17070),.clk(gclk));
	jor g16775(.dina(n17070),.dinb(w_n17058_0[1]),.dout(n17071),.clk(gclk));
	jand g16776(.dina(w_n17071_0[1]),.dinb(w_asqrt59_12[1]),.dout(n17072),.clk(gclk));
	jxor g16777(.dina(w_n16440_0[0]),.dinb(w_n425_15[0]),.dout(n17073),.clk(gclk));
	jand g16778(.dina(n17073),.dinb(w_asqrt8_14[1]),.dout(n17074),.clk(gclk));
	jxor g16779(.dina(n17074),.dinb(w_n16450_0[0]),.dout(n17075),.clk(gclk));
	jnot g16780(.din(n17075),.dout(n17076),.clk(gclk));
	jor g16781(.dina(w_n17071_0[0]),.dinb(w_asqrt59_12[0]),.dout(n17077),.clk(gclk));
	jand g16782(.dina(w_n17077_0[1]),.dinb(w_n17076_0[1]),.dout(n17078),.clk(gclk));
	jor g16783(.dina(w_n17078_0[2]),.dinb(w_n17072_0[2]),.dout(n17079),.clk(gclk));
	jand g16784(.dina(n17079),.dinb(w_asqrt60_12[1]),.dout(n17080),.clk(gclk));
	jnot g16785(.din(w_n16455_0[0]),.dout(n17081),.clk(gclk));
	jand g16786(.dina(n17081),.dinb(w_n16453_0[0]),.dout(n17082),.clk(gclk));
	jand g16787(.dina(n17082),.dinb(w_asqrt8_14[0]),.dout(n17083),.clk(gclk));
	jxor g16788(.dina(n17083),.dinb(w_n16463_0[0]),.dout(n17084),.clk(gclk));
	jnot g16789(.din(n17084),.dout(n17085),.clk(gclk));
	jor g16790(.dina(w_n17072_0[1]),.dinb(w_asqrt60_12[0]),.dout(n17086),.clk(gclk));
	jor g16791(.dina(n17086),.dinb(w_n17078_0[1]),.dout(n17087),.clk(gclk));
	jand g16792(.dina(w_n17087_0[1]),.dinb(w_n17085_0[1]),.dout(n17088),.clk(gclk));
	jor g16793(.dina(w_n17088_0[1]),.dinb(w_n17080_0[1]),.dout(n17089),.clk(gclk));
	jand g16794(.dina(w_n17089_0[2]),.dinb(w_asqrt61_12[2]),.dout(n17090),.clk(gclk));
	jor g16795(.dina(w_n17089_0[1]),.dinb(w_asqrt61_12[1]),.dout(n17091),.clk(gclk));
	jnot g16796(.din(w_n16469_0[0]),.dout(n17092),.clk(gclk));
	jnot g16797(.din(w_n16470_0[0]),.dout(n17093),.clk(gclk));
	jand g16798(.dina(w_asqrt8_13[2]),.dinb(w_n16466_0[0]),.dout(n17094),.clk(gclk));
	jand g16799(.dina(w_n17094_0[1]),.dinb(n17093),.dout(n17095),.clk(gclk));
	jor g16800(.dina(n17095),.dinb(n17092),.dout(n17096),.clk(gclk));
	jnot g16801(.din(w_n16471_0[0]),.dout(n17097),.clk(gclk));
	jand g16802(.dina(w_n17094_0[0]),.dinb(n17097),.dout(n17098),.clk(gclk));
	jnot g16803(.din(n17098),.dout(n17099),.clk(gclk));
	jand g16804(.dina(n17099),.dinb(n17096),.dout(n17100),.clk(gclk));
	jand g16805(.dina(w_n17100_0[1]),.dinb(n17091),.dout(n17101),.clk(gclk));
	jor g16806(.dina(w_n17101_0[1]),.dinb(w_n17090_0[1]),.dout(n17102),.clk(gclk));
	jand g16807(.dina(n17102),.dinb(w_asqrt62_12[2]),.dout(n17103),.clk(gclk));
	jor g16808(.dina(w_n17090_0[0]),.dinb(w_asqrt62_12[1]),.dout(n17104),.clk(gclk));
	jor g16809(.dina(n17104),.dinb(w_n17101_0[0]),.dout(n17105),.clk(gclk));
	jnot g16810(.din(w_n16477_0[0]),.dout(n17106),.clk(gclk));
	jnot g16811(.din(w_n16479_0[0]),.dout(n17107),.clk(gclk));
	jand g16812(.dina(w_asqrt8_13[1]),.dinb(w_n16473_0[0]),.dout(n17108),.clk(gclk));
	jand g16813(.dina(w_n17108_0[1]),.dinb(n17107),.dout(n17109),.clk(gclk));
	jor g16814(.dina(n17109),.dinb(n17106),.dout(n17110),.clk(gclk));
	jnot g16815(.din(w_n16480_0[0]),.dout(n17111),.clk(gclk));
	jand g16816(.dina(w_n17108_0[0]),.dinb(n17111),.dout(n17112),.clk(gclk));
	jnot g16817(.din(n17112),.dout(n17113),.clk(gclk));
	jand g16818(.dina(n17113),.dinb(n17110),.dout(n17114),.clk(gclk));
	jand g16819(.dina(w_n17114_0[1]),.dinb(w_n17105_0[1]),.dout(n17115),.clk(gclk));
	jor g16820(.dina(n17115),.dinb(w_n17103_0[1]),.dout(n17116),.clk(gclk));
	jxor g16821(.dina(w_n16481_0[0]),.dinb(w_n199_18[2]),.dout(n17117),.clk(gclk));
	jand g16822(.dina(n17117),.dinb(w_asqrt8_13[0]),.dout(n17118),.clk(gclk));
	jxor g16823(.dina(n17118),.dinb(w_n16491_0[0]),.dout(n17119),.clk(gclk));
	jnot g16824(.din(w_n16493_0[0]),.dout(n17120),.clk(gclk));
	jand g16825(.dina(w_asqrt8_12[2]),.dinb(w_n16500_0[1]),.dout(n17121),.clk(gclk));
	jand g16826(.dina(w_n17121_0[1]),.dinb(w_n17120_0[2]),.dout(n17122),.clk(gclk));
	jor g16827(.dina(n17122),.dinb(w_n16508_0[0]),.dout(n17123),.clk(gclk));
	jor g16828(.dina(n17123),.dinb(w_n17119_0[1]),.dout(n17124),.clk(gclk));
	jnot g16829(.din(n17124),.dout(n17125),.clk(gclk));
	jand g16830(.dina(n17125),.dinb(w_n17116_1[2]),.dout(n17126),.clk(gclk));
	jor g16831(.dina(n17126),.dinb(w_asqrt63_7[0]),.dout(n17127),.clk(gclk));
	jnot g16832(.din(w_n17119_0[0]),.dout(n17128),.clk(gclk));
	jor g16833(.dina(w_n17128_0[2]),.dinb(w_n17116_1[1]),.dout(n17129),.clk(gclk));
	jor g16834(.dina(w_n17121_0[0]),.dinb(w_n17120_0[1]),.dout(n17130),.clk(gclk));
	jand g16835(.dina(w_n16500_0[0]),.dinb(w_n17120_0[0]),.dout(n17131),.clk(gclk));
	jor g16836(.dina(n17131),.dinb(w_n194_17[2]),.dout(n17132),.clk(gclk));
	jnot g16837(.din(n17132),.dout(n17133),.clk(gclk));
	jand g16838(.dina(n17133),.dinb(n17130),.dout(n17134),.clk(gclk));
	jnot g16839(.din(w_asqrt8_12[1]),.dout(n17135),.clk(gclk));
	jnot g16840(.din(w_n17134_0[1]),.dout(n17138),.clk(gclk));
	jand g16841(.dina(n17138),.dinb(w_n17129_0[1]),.dout(n17139),.clk(gclk));
	jand g16842(.dina(n17139),.dinb(w_n17127_0[1]),.dout(n17140),.clk(gclk));
	jxor g16843(.dina(w_n17026_0[0]),.dinb(w_n595_16[0]),.dout(n17141),.clk(gclk));
	jor g16844(.dina(n17141),.dinb(w_n17140_20[2]),.dout(n17142),.clk(gclk));
	jxor g16845(.dina(n17142),.dinb(w_n16521_0[0]),.dout(n17143),.clk(gclk));
	jor g16846(.dina(w_n17140_20[1]),.dinb(w_n16523_1[0]),.dout(n17144),.clk(gclk));
	jnot g16847(.din(w_a12_0[1]),.dout(n17145),.clk(gclk));
	jnot g16848(.din(a[13]),.dout(n17146),.clk(gclk));
	jand g16849(.dina(w_n16523_0[2]),.dinb(w_n17146_0[2]),.dout(n17147),.clk(gclk));
	jand g16850(.dina(n17147),.dinb(w_n17145_1[1]),.dout(n17148),.clk(gclk));
	jnot g16851(.din(n17148),.dout(n17149),.clk(gclk));
	jand g16852(.dina(n17149),.dinb(n17144),.dout(n17150),.clk(gclk));
	jor g16853(.dina(w_n17150_0[2]),.dinb(w_n17135_5[1]),.dout(n17151),.clk(gclk));
	jor g16854(.dina(w_n17140_20[0]),.dinb(w_a14_0[0]),.dout(n17152),.clk(gclk));
	jxor g16855(.dina(w_n17152_0[1]),.dinb(w_n16524_0[0]),.dout(n17153),.clk(gclk));
	jand g16856(.dina(w_n17150_0[1]),.dinb(w_n17135_5[0]),.dout(n17154),.clk(gclk));
	jor g16857(.dina(n17154),.dinb(w_n17153_0[1]),.dout(n17155),.clk(gclk));
	jand g16858(.dina(w_n17155_0[1]),.dinb(w_n17151_0[1]),.dout(n17156),.clk(gclk));
	jor g16859(.dina(n17156),.dinb(w_n15955_10[2]),.dout(n17157),.clk(gclk));
	jand g16860(.dina(w_n17151_0[0]),.dinb(w_n15955_10[1]),.dout(n17158),.clk(gclk));
	jand g16861(.dina(n17158),.dinb(w_n17155_0[0]),.dout(n17159),.clk(gclk));
	jor g16862(.dina(w_n17152_0[0]),.dinb(w_a15_0[0]),.dout(n17160),.clk(gclk));
	jnot g16863(.din(w_n17127_0[0]),.dout(n17161),.clk(gclk));
	jnot g16864(.din(w_n17129_0[0]),.dout(n17162),.clk(gclk));
	jor g16865(.dina(w_n17134_0[0]),.dinb(w_n17135_4[2]),.dout(n17163),.clk(gclk));
	jor g16866(.dina(n17163),.dinb(w_n17162_0[1]),.dout(n17164),.clk(gclk));
	jor g16867(.dina(n17164),.dinb(n17161),.dout(n17165),.clk(gclk));
	jand g16868(.dina(n17165),.dinb(n17160),.dout(n17166),.clk(gclk));
	jxor g16869(.dina(n17166),.dinb(w_n15961_0[1]),.dout(n17167),.clk(gclk));
	jor g16870(.dina(w_n17167_0[1]),.dinb(w_n17159_0[1]),.dout(n17168),.clk(gclk));
	jand g16871(.dina(n17168),.dinb(w_n17157_0[1]),.dout(n17169),.clk(gclk));
	jor g16872(.dina(w_n17169_0[2]),.dinb(w_n15950_5[1]),.dout(n17170),.clk(gclk));
	jand g16873(.dina(w_n17169_0[1]),.dinb(w_n15950_5[0]),.dout(n17171),.clk(gclk));
	jxor g16874(.dina(w_n16527_0[0]),.dinb(w_n15955_10[0]),.dout(n17172),.clk(gclk));
	jor g16875(.dina(n17172),.dinb(w_n17140_19[2]),.dout(n17173),.clk(gclk));
	jxor g16876(.dina(n17173),.dinb(w_n16530_0[0]),.dout(n17174),.clk(gclk));
	jor g16877(.dina(w_n17174_0[1]),.dinb(n17171),.dout(n17175),.clk(gclk));
	jand g16878(.dina(w_n17175_0[1]),.dinb(w_n17170_0[1]),.dout(n17176),.clk(gclk));
	jor g16879(.dina(n17176),.dinb(w_n14821_11[0]),.dout(n17177),.clk(gclk));
	jnot g16880(.din(w_n16536_0[0]),.dout(n17178),.clk(gclk));
	jor g16881(.dina(n17178),.dinb(w_n16534_0[0]),.dout(n17179),.clk(gclk));
	jor g16882(.dina(n17179),.dinb(w_n17140_19[1]),.dout(n17180),.clk(gclk));
	jxor g16883(.dina(n17180),.dinb(w_n16545_0[0]),.dout(n17181),.clk(gclk));
	jand g16884(.dina(w_n17170_0[0]),.dinb(w_n14821_10[2]),.dout(n17182),.clk(gclk));
	jand g16885(.dina(n17182),.dinb(w_n17175_0[0]),.dout(n17183),.clk(gclk));
	jor g16886(.dina(w_n17183_0[1]),.dinb(w_n17181_0[1]),.dout(n17184),.clk(gclk));
	jand g16887(.dina(w_n17184_0[1]),.dinb(w_n17177_0[1]),.dout(n17185),.clk(gclk));
	jor g16888(.dina(w_n17185_0[2]),.dinb(w_n14816_6[0]),.dout(n17186),.clk(gclk));
	jand g16889(.dina(w_n17185_0[1]),.dinb(w_n14816_5[2]),.dout(n17187),.clk(gclk));
	jxor g16890(.dina(w_n16547_0[0]),.dinb(w_n14821_10[1]),.dout(n17188),.clk(gclk));
	jor g16891(.dina(n17188),.dinb(w_n17140_19[0]),.dout(n17189),.clk(gclk));
	jxor g16892(.dina(n17189),.dinb(w_n16552_0[0]),.dout(n17190),.clk(gclk));
	jnot g16893(.din(w_n17190_0[1]),.dout(n17191),.clk(gclk));
	jor g16894(.dina(n17191),.dinb(n17187),.dout(n17192),.clk(gclk));
	jand g16895(.dina(w_n17192_0[1]),.dinb(w_n17186_0[1]),.dout(n17193),.clk(gclk));
	jor g16896(.dina(n17193),.dinb(w_n13723_10[2]),.dout(n17194),.clk(gclk));
	jand g16897(.dina(w_n17186_0[0]),.dinb(w_n13723_10[1]),.dout(n17195),.clk(gclk));
	jand g16898(.dina(n17195),.dinb(w_n17192_0[0]),.dout(n17196),.clk(gclk));
	jnot g16899(.din(w_n16556_0[0]),.dout(n17197),.clk(gclk));
	jnot g16900(.din(w_n17140_18[2]),.dout(asqrt_fa_8),.clk(gclk));
	jand g16901(.dina(w_asqrt7_15),.dinb(n17197),.dout(n17199),.clk(gclk));
	jand g16902(.dina(w_n17199_0[1]),.dinb(w_n16563_0[0]),.dout(n17200),.clk(gclk));
	jor g16903(.dina(n17200),.dinb(w_n16561_0[0]),.dout(n17201),.clk(gclk));
	jand g16904(.dina(w_n17199_0[0]),.dinb(w_n16564_0[0]),.dout(n17202),.clk(gclk));
	jnot g16905(.din(n17202),.dout(n17203),.clk(gclk));
	jand g16906(.dina(n17203),.dinb(n17201),.dout(n17204),.clk(gclk));
	jnot g16907(.din(n17204),.dout(n17205),.clk(gclk));
	jor g16908(.dina(w_n17205_0[1]),.dinb(w_n17196_0[1]),.dout(n17206),.clk(gclk));
	jand g16909(.dina(n17206),.dinb(w_n17194_0[1]),.dout(n17207),.clk(gclk));
	jor g16910(.dina(w_n17207_0[2]),.dinb(w_n13718_6[0]),.dout(n17208),.clk(gclk));
	jand g16911(.dina(w_n17207_0[1]),.dinb(w_n13718_5[2]),.dout(n17209),.clk(gclk));
	jnot g16912(.din(w_n16571_0[0]),.dout(n17210),.clk(gclk));
	jxor g16913(.dina(w_n16565_0[0]),.dinb(w_n13723_10[0]),.dout(n17211),.clk(gclk));
	jor g16914(.dina(n17211),.dinb(w_n17140_18[1]),.dout(n17212),.clk(gclk));
	jxor g16915(.dina(n17212),.dinb(n17210),.dout(n17213),.clk(gclk));
	jnot g16916(.din(w_n17213_0[1]),.dout(n17214),.clk(gclk));
	jor g16917(.dina(n17214),.dinb(n17209),.dout(n17215),.clk(gclk));
	jand g16918(.dina(w_n17215_0[1]),.dinb(w_n17208_0[1]),.dout(n17216),.clk(gclk));
	jor g16919(.dina(n17216),.dinb(w_n12675_11[1]),.dout(n17217),.clk(gclk));
	jnot g16920(.din(w_n16576_0[0]),.dout(n17218),.clk(gclk));
	jor g16921(.dina(n17218),.dinb(w_n16574_0[0]),.dout(n17219),.clk(gclk));
	jor g16922(.dina(n17219),.dinb(w_n17140_18[0]),.dout(n17220),.clk(gclk));
	jxor g16923(.dina(n17220),.dinb(w_n16585_0[0]),.dout(n17221),.clk(gclk));
	jand g16924(.dina(w_n17208_0[0]),.dinb(w_n12675_11[0]),.dout(n17222),.clk(gclk));
	jand g16925(.dina(n17222),.dinb(w_n17215_0[0]),.dout(n17223),.clk(gclk));
	jor g16926(.dina(w_n17223_0[1]),.dinb(w_n17221_0[1]),.dout(n17224),.clk(gclk));
	jand g16927(.dina(w_n17224_0[1]),.dinb(w_n17217_0[1]),.dout(n17225),.clk(gclk));
	jor g16928(.dina(w_n17225_0[2]),.dinb(w_n12670_6[1]),.dout(n17226),.clk(gclk));
	jand g16929(.dina(w_n17225_0[1]),.dinb(w_n12670_6[0]),.dout(n17227),.clk(gclk));
	jnot g16930(.din(w_n16592_0[0]),.dout(n17228),.clk(gclk));
	jxor g16931(.dina(w_n16587_0[0]),.dinb(w_n12675_10[2]),.dout(n17229),.clk(gclk));
	jor g16932(.dina(n17229),.dinb(w_n17140_17[2]),.dout(n17230),.clk(gclk));
	jxor g16933(.dina(n17230),.dinb(n17228),.dout(n17231),.clk(gclk));
	jnot g16934(.din(n17231),.dout(n17232),.clk(gclk));
	jor g16935(.dina(w_n17232_0[1]),.dinb(n17227),.dout(n17233),.clk(gclk));
	jand g16936(.dina(w_n17233_0[1]),.dinb(w_n17226_0[1]),.dout(n17234),.clk(gclk));
	jor g16937(.dina(n17234),.dinb(w_n11662_11[0]),.dout(n17235),.clk(gclk));
	jand g16938(.dina(w_n17226_0[0]),.dinb(w_n11662_10[2]),.dout(n17236),.clk(gclk));
	jand g16939(.dina(n17236),.dinb(w_n17233_0[0]),.dout(n17237),.clk(gclk));
	jnot g16940(.din(w_n16595_0[0]),.dout(n17238),.clk(gclk));
	jand g16941(.dina(w_asqrt7_14[2]),.dinb(n17238),.dout(n17239),.clk(gclk));
	jand g16942(.dina(w_n17239_0[1]),.dinb(w_n16602_0[0]),.dout(n17240),.clk(gclk));
	jor g16943(.dina(n17240),.dinb(w_n16600_0[0]),.dout(n17241),.clk(gclk));
	jand g16944(.dina(w_n17239_0[0]),.dinb(w_n16603_0[0]),.dout(n17242),.clk(gclk));
	jnot g16945(.din(n17242),.dout(n17243),.clk(gclk));
	jand g16946(.dina(n17243),.dinb(n17241),.dout(n17244),.clk(gclk));
	jnot g16947(.din(n17244),.dout(n17245),.clk(gclk));
	jor g16948(.dina(w_n17245_0[1]),.dinb(w_n17237_0[1]),.dout(n17246),.clk(gclk));
	jand g16949(.dina(n17246),.dinb(w_n17235_0[1]),.dout(n17247),.clk(gclk));
	jor g16950(.dina(w_n17247_0[1]),.dinb(w_n11657_6[1]),.dout(n17248),.clk(gclk));
	jxor g16951(.dina(w_n16604_0[0]),.dinb(w_n11662_10[1]),.dout(n17249),.clk(gclk));
	jor g16952(.dina(n17249),.dinb(w_n17140_17[1]),.dout(n17250),.clk(gclk));
	jxor g16953(.dina(n17250),.dinb(w_n16609_0[0]),.dout(n17251),.clk(gclk));
	jand g16954(.dina(w_n17247_0[0]),.dinb(w_n11657_6[0]),.dout(n17252),.clk(gclk));
	jor g16955(.dina(w_n17252_0[1]),.dinb(w_n17251_0[1]),.dout(n17253),.clk(gclk));
	jand g16956(.dina(w_n17253_0[2]),.dinb(w_n17248_0[2]),.dout(n17254),.clk(gclk));
	jor g16957(.dina(n17254),.dinb(w_n10701_11[1]),.dout(n17255),.clk(gclk));
	jnot g16958(.din(w_n16614_0[0]),.dout(n17256),.clk(gclk));
	jor g16959(.dina(n17256),.dinb(w_n16612_0[0]),.dout(n17257),.clk(gclk));
	jor g16960(.dina(n17257),.dinb(w_n17140_17[0]),.dout(n17258),.clk(gclk));
	jxor g16961(.dina(n17258),.dinb(w_n16623_0[0]),.dout(n17259),.clk(gclk));
	jand g16962(.dina(w_n17248_0[1]),.dinb(w_n10701_11[0]),.dout(n17260),.clk(gclk));
	jand g16963(.dina(n17260),.dinb(w_n17253_0[1]),.dout(n17261),.clk(gclk));
	jor g16964(.dina(w_n17261_0[1]),.dinb(w_n17259_0[1]),.dout(n17262),.clk(gclk));
	jand g16965(.dina(w_n17262_0[1]),.dinb(w_n17255_0[1]),.dout(n17263),.clk(gclk));
	jor g16966(.dina(w_n17263_0[2]),.dinb(w_n10696_7[1]),.dout(n17264),.clk(gclk));
	jand g16967(.dina(w_n17263_0[1]),.dinb(w_n10696_7[0]),.dout(n17265),.clk(gclk));
	jnot g16968(.din(w_n16626_0[0]),.dout(n17266),.clk(gclk));
	jand g16969(.dina(w_asqrt7_14[1]),.dinb(n17266),.dout(n17267),.clk(gclk));
	jand g16970(.dina(w_n17267_0[1]),.dinb(w_n16631_0[0]),.dout(n17268),.clk(gclk));
	jor g16971(.dina(n17268),.dinb(w_n16630_0[0]),.dout(n17269),.clk(gclk));
	jand g16972(.dina(w_n17267_0[0]),.dinb(w_n16632_0[0]),.dout(n17270),.clk(gclk));
	jnot g16973(.din(n17270),.dout(n17271),.clk(gclk));
	jand g16974(.dina(n17271),.dinb(n17269),.dout(n17272),.clk(gclk));
	jnot g16975(.din(n17272),.dout(n17273),.clk(gclk));
	jor g16976(.dina(w_n17273_0[1]),.dinb(n17265),.dout(n17274),.clk(gclk));
	jand g16977(.dina(w_n17274_0[1]),.dinb(w_n17264_0[1]),.dout(n17275),.clk(gclk));
	jor g16978(.dina(n17275),.dinb(w_n9774_11[1]),.dout(n17276),.clk(gclk));
	jand g16979(.dina(w_n17264_0[0]),.dinb(w_n9774_11[0]),.dout(n17277),.clk(gclk));
	jand g16980(.dina(n17277),.dinb(w_n17274_0[0]),.dout(n17278),.clk(gclk));
	jnot g16981(.din(w_n16634_0[0]),.dout(n17279),.clk(gclk));
	jand g16982(.dina(w_asqrt7_14[0]),.dinb(n17279),.dout(n17280),.clk(gclk));
	jand g16983(.dina(w_n17280_0[1]),.dinb(w_n16641_0[0]),.dout(n17281),.clk(gclk));
	jor g16984(.dina(n17281),.dinb(w_n16639_0[0]),.dout(n17282),.clk(gclk));
	jand g16985(.dina(w_n17280_0[0]),.dinb(w_n16642_0[0]),.dout(n17283),.clk(gclk));
	jnot g16986(.din(n17283),.dout(n17284),.clk(gclk));
	jand g16987(.dina(n17284),.dinb(n17282),.dout(n17285),.clk(gclk));
	jnot g16988(.din(n17285),.dout(n17286),.clk(gclk));
	jor g16989(.dina(w_n17286_0[1]),.dinb(w_n17278_0[1]),.dout(n17287),.clk(gclk));
	jand g16990(.dina(n17287),.dinb(w_n17276_0[1]),.dout(n17288),.clk(gclk));
	jor g16991(.dina(w_n17288_0[1]),.dinb(w_n9769_7[1]),.dout(n17289),.clk(gclk));
	jxor g16992(.dina(w_n16643_0[0]),.dinb(w_n9774_10[2]),.dout(n17290),.clk(gclk));
	jor g16993(.dina(n17290),.dinb(w_n17140_16[2]),.dout(n17291),.clk(gclk));
	jxor g16994(.dina(n17291),.dinb(w_n16654_0[0]),.dout(n17292),.clk(gclk));
	jand g16995(.dina(w_n17288_0[0]),.dinb(w_n9769_7[0]),.dout(n17293),.clk(gclk));
	jor g16996(.dina(w_n17293_0[1]),.dinb(w_n17292_0[1]),.dout(n17294),.clk(gclk));
	jand g16997(.dina(w_n17294_0[2]),.dinb(w_n17289_0[2]),.dout(n17295),.clk(gclk));
	jor g16998(.dina(n17295),.dinb(w_n8898_12[0]),.dout(n17296),.clk(gclk));
	jnot g16999(.din(w_n16659_0[0]),.dout(n17297),.clk(gclk));
	jor g17000(.dina(n17297),.dinb(w_n16657_0[0]),.dout(n17298),.clk(gclk));
	jor g17001(.dina(n17298),.dinb(w_n17140_16[1]),.dout(n17299),.clk(gclk));
	jxor g17002(.dina(n17299),.dinb(w_n16668_0[0]),.dout(n17300),.clk(gclk));
	jand g17003(.dina(w_n17289_0[1]),.dinb(w_n8898_11[2]),.dout(n17301),.clk(gclk));
	jand g17004(.dina(n17301),.dinb(w_n17294_0[1]),.dout(n17302),.clk(gclk));
	jor g17005(.dina(w_n17302_0[1]),.dinb(w_n17300_0[1]),.dout(n17303),.clk(gclk));
	jand g17006(.dina(w_n17303_0[1]),.dinb(w_n17296_0[1]),.dout(n17304),.clk(gclk));
	jor g17007(.dina(w_n17304_0[2]),.dinb(w_n8893_8[0]),.dout(n17305),.clk(gclk));
	jand g17008(.dina(w_n17304_0[1]),.dinb(w_n8893_7[2]),.dout(n17306),.clk(gclk));
	jnot g17009(.din(w_n16671_0[0]),.dout(n17307),.clk(gclk));
	jand g17010(.dina(w_asqrt7_13[2]),.dinb(n17307),.dout(n17308),.clk(gclk));
	jand g17011(.dina(w_n17308_0[1]),.dinb(w_n16676_0[0]),.dout(n17309),.clk(gclk));
	jor g17012(.dina(n17309),.dinb(w_n16675_0[0]),.dout(n17310),.clk(gclk));
	jand g17013(.dina(w_n17308_0[0]),.dinb(w_n16677_0[0]),.dout(n17311),.clk(gclk));
	jnot g17014(.din(n17311),.dout(n17312),.clk(gclk));
	jand g17015(.dina(n17312),.dinb(n17310),.dout(n17313),.clk(gclk));
	jnot g17016(.din(n17313),.dout(n17314),.clk(gclk));
	jor g17017(.dina(w_n17314_0[1]),.dinb(n17306),.dout(n17315),.clk(gclk));
	jand g17018(.dina(w_n17315_0[1]),.dinb(w_n17305_0[1]),.dout(n17316),.clk(gclk));
	jor g17019(.dina(n17316),.dinb(w_n8058_12[0]),.dout(n17317),.clk(gclk));
	jand g17020(.dina(w_n17305_0[0]),.dinb(w_n8058_11[2]),.dout(n17318),.clk(gclk));
	jand g17021(.dina(n17318),.dinb(w_n17315_0[0]),.dout(n17319),.clk(gclk));
	jnot g17022(.din(w_n16679_0[0]),.dout(n17320),.clk(gclk));
	jand g17023(.dina(w_asqrt7_13[1]),.dinb(n17320),.dout(n17321),.clk(gclk));
	jand g17024(.dina(w_n17321_0[1]),.dinb(w_n16686_0[0]),.dout(n17322),.clk(gclk));
	jor g17025(.dina(n17322),.dinb(w_n16684_0[0]),.dout(n17323),.clk(gclk));
	jand g17026(.dina(w_n17321_0[0]),.dinb(w_n16687_0[0]),.dout(n17324),.clk(gclk));
	jnot g17027(.din(n17324),.dout(n17325),.clk(gclk));
	jand g17028(.dina(n17325),.dinb(n17323),.dout(n17326),.clk(gclk));
	jnot g17029(.din(n17326),.dout(n17327),.clk(gclk));
	jor g17030(.dina(w_n17327_0[1]),.dinb(w_n17319_0[1]),.dout(n17328),.clk(gclk));
	jand g17031(.dina(n17328),.dinb(w_n17317_0[1]),.dout(n17329),.clk(gclk));
	jor g17032(.dina(w_n17329_0[1]),.dinb(w_n8053_8[0]),.dout(n17330),.clk(gclk));
	jxor g17033(.dina(w_n16688_0[0]),.dinb(w_n8058_11[1]),.dout(n17331),.clk(gclk));
	jor g17034(.dina(n17331),.dinb(w_n17140_16[0]),.dout(n17332),.clk(gclk));
	jxor g17035(.dina(n17332),.dinb(w_n16699_0[0]),.dout(n17333),.clk(gclk));
	jand g17036(.dina(w_n17329_0[0]),.dinb(w_n8053_7[2]),.dout(n17334),.clk(gclk));
	jor g17037(.dina(w_n17334_0[1]),.dinb(w_n17333_0[1]),.dout(n17335),.clk(gclk));
	jand g17038(.dina(w_n17335_0[2]),.dinb(w_n17330_0[2]),.dout(n17336),.clk(gclk));
	jor g17039(.dina(n17336),.dinb(w_n7265_12[1]),.dout(n17337),.clk(gclk));
	jnot g17040(.din(w_n16704_0[0]),.dout(n17338),.clk(gclk));
	jor g17041(.dina(n17338),.dinb(w_n16702_0[0]),.dout(n17339),.clk(gclk));
	jor g17042(.dina(n17339),.dinb(w_n17140_15[2]),.dout(n17340),.clk(gclk));
	jxor g17043(.dina(n17340),.dinb(w_n16713_0[0]),.dout(n17341),.clk(gclk));
	jand g17044(.dina(w_n17330_0[1]),.dinb(w_n7265_12[0]),.dout(n17342),.clk(gclk));
	jand g17045(.dina(n17342),.dinb(w_n17335_0[1]),.dout(n17343),.clk(gclk));
	jor g17046(.dina(w_n17343_0[1]),.dinb(w_n17341_0[1]),.dout(n17344),.clk(gclk));
	jand g17047(.dina(w_n17344_0[1]),.dinb(w_n17337_0[1]),.dout(n17345),.clk(gclk));
	jor g17048(.dina(w_n17345_0[2]),.dinb(w_n7260_9[0]),.dout(n17346),.clk(gclk));
	jand g17049(.dina(w_n17345_0[1]),.dinb(w_n7260_8[2]),.dout(n17347),.clk(gclk));
	jnot g17050(.din(w_n16716_0[0]),.dout(n17348),.clk(gclk));
	jand g17051(.dina(w_asqrt7_13[0]),.dinb(n17348),.dout(n17349),.clk(gclk));
	jand g17052(.dina(w_n17349_0[1]),.dinb(w_n16721_0[0]),.dout(n17350),.clk(gclk));
	jor g17053(.dina(n17350),.dinb(w_n16720_0[0]),.dout(n17351),.clk(gclk));
	jand g17054(.dina(w_n17349_0[0]),.dinb(w_n16722_0[0]),.dout(n17352),.clk(gclk));
	jnot g17055(.din(n17352),.dout(n17353),.clk(gclk));
	jand g17056(.dina(n17353),.dinb(n17351),.dout(n17354),.clk(gclk));
	jnot g17057(.din(n17354),.dout(n17355),.clk(gclk));
	jor g17058(.dina(w_n17355_0[1]),.dinb(n17347),.dout(n17356),.clk(gclk));
	jand g17059(.dina(w_n17356_0[1]),.dinb(w_n17346_0[1]),.dout(n17357),.clk(gclk));
	jor g17060(.dina(n17357),.dinb(w_n6505_12[1]),.dout(n17358),.clk(gclk));
	jand g17061(.dina(w_n17346_0[0]),.dinb(w_n6505_12[0]),.dout(n17359),.clk(gclk));
	jand g17062(.dina(n17359),.dinb(w_n17356_0[0]),.dout(n17360),.clk(gclk));
	jnot g17063(.din(w_n16724_0[0]),.dout(n17361),.clk(gclk));
	jand g17064(.dina(w_asqrt7_12[2]),.dinb(n17361),.dout(n17362),.clk(gclk));
	jand g17065(.dina(w_n17362_0[1]),.dinb(w_n16731_0[0]),.dout(n17363),.clk(gclk));
	jor g17066(.dina(n17363),.dinb(w_n16729_0[0]),.dout(n17364),.clk(gclk));
	jand g17067(.dina(w_n17362_0[0]),.dinb(w_n16732_0[0]),.dout(n17365),.clk(gclk));
	jnot g17068(.din(n17365),.dout(n17366),.clk(gclk));
	jand g17069(.dina(n17366),.dinb(n17364),.dout(n17367),.clk(gclk));
	jnot g17070(.din(n17367),.dout(n17368),.clk(gclk));
	jor g17071(.dina(w_n17368_0[1]),.dinb(w_n17360_0[1]),.dout(n17369),.clk(gclk));
	jand g17072(.dina(n17369),.dinb(w_n17358_0[1]),.dout(n17370),.clk(gclk));
	jor g17073(.dina(w_n17370_0[1]),.dinb(w_n6500_9[0]),.dout(n17371),.clk(gclk));
	jxor g17074(.dina(w_n16733_0[0]),.dinb(w_n6505_11[2]),.dout(n17372),.clk(gclk));
	jor g17075(.dina(n17372),.dinb(w_n17140_15[1]),.dout(n17373),.clk(gclk));
	jxor g17076(.dina(n17373),.dinb(w_n16744_0[0]),.dout(n17374),.clk(gclk));
	jand g17077(.dina(w_n17370_0[0]),.dinb(w_n6500_8[2]),.dout(n17375),.clk(gclk));
	jor g17078(.dina(w_n17375_0[1]),.dinb(w_n17374_0[1]),.dout(n17376),.clk(gclk));
	jand g17079(.dina(w_n17376_0[2]),.dinb(w_n17371_0[2]),.dout(n17377),.clk(gclk));
	jor g17080(.dina(n17377),.dinb(w_n5793_12[2]),.dout(n17378),.clk(gclk));
	jnot g17081(.din(w_n16749_0[0]),.dout(n17379),.clk(gclk));
	jor g17082(.dina(n17379),.dinb(w_n16747_0[0]),.dout(n17380),.clk(gclk));
	jor g17083(.dina(n17380),.dinb(w_n17140_15[0]),.dout(n17381),.clk(gclk));
	jxor g17084(.dina(n17381),.dinb(w_n16758_0[0]),.dout(n17382),.clk(gclk));
	jand g17085(.dina(w_n17371_0[1]),.dinb(w_n5793_12[1]),.dout(n17383),.clk(gclk));
	jand g17086(.dina(n17383),.dinb(w_n17376_0[1]),.dout(n17384),.clk(gclk));
	jor g17087(.dina(w_n17384_0[1]),.dinb(w_n17382_0[1]),.dout(n17385),.clk(gclk));
	jand g17088(.dina(w_n17385_0[1]),.dinb(w_n17378_0[1]),.dout(n17386),.clk(gclk));
	jor g17089(.dina(w_n17386_0[2]),.dinb(w_n5788_9[2]),.dout(n17387),.clk(gclk));
	jand g17090(.dina(w_n17386_0[1]),.dinb(w_n5788_9[1]),.dout(n17388),.clk(gclk));
	jnot g17091(.din(w_n16761_0[0]),.dout(n17389),.clk(gclk));
	jand g17092(.dina(w_asqrt7_12[1]),.dinb(n17389),.dout(n17390),.clk(gclk));
	jand g17093(.dina(w_n17390_0[1]),.dinb(w_n16766_0[0]),.dout(n17391),.clk(gclk));
	jor g17094(.dina(n17391),.dinb(w_n16765_0[0]),.dout(n17392),.clk(gclk));
	jand g17095(.dina(w_n17390_0[0]),.dinb(w_n16767_0[0]),.dout(n17393),.clk(gclk));
	jnot g17096(.din(n17393),.dout(n17394),.clk(gclk));
	jand g17097(.dina(n17394),.dinb(n17392),.dout(n17395),.clk(gclk));
	jnot g17098(.din(n17395),.dout(n17396),.clk(gclk));
	jor g17099(.dina(w_n17396_0[1]),.dinb(n17388),.dout(n17397),.clk(gclk));
	jand g17100(.dina(w_n17397_0[1]),.dinb(w_n17387_0[1]),.dout(n17398),.clk(gclk));
	jor g17101(.dina(n17398),.dinb(w_n5121_12[2]),.dout(n17399),.clk(gclk));
	jand g17102(.dina(w_n17387_0[0]),.dinb(w_n5121_12[1]),.dout(n17400),.clk(gclk));
	jand g17103(.dina(n17400),.dinb(w_n17397_0[0]),.dout(n17401),.clk(gclk));
	jnot g17104(.din(w_n16769_0[0]),.dout(n17402),.clk(gclk));
	jand g17105(.dina(w_asqrt7_12[0]),.dinb(n17402),.dout(n17403),.clk(gclk));
	jand g17106(.dina(w_n17403_0[1]),.dinb(w_n16776_0[0]),.dout(n17404),.clk(gclk));
	jor g17107(.dina(n17404),.dinb(w_n16774_0[0]),.dout(n17405),.clk(gclk));
	jand g17108(.dina(w_n17403_0[0]),.dinb(w_n16777_0[0]),.dout(n17406),.clk(gclk));
	jnot g17109(.din(n17406),.dout(n17407),.clk(gclk));
	jand g17110(.dina(n17407),.dinb(n17405),.dout(n17408),.clk(gclk));
	jnot g17111(.din(n17408),.dout(n17409),.clk(gclk));
	jor g17112(.dina(w_n17409_0[1]),.dinb(w_n17401_0[1]),.dout(n17410),.clk(gclk));
	jand g17113(.dina(n17410),.dinb(w_n17399_0[1]),.dout(n17411),.clk(gclk));
	jor g17114(.dina(w_n17411_0[1]),.dinb(w_n5116_9[2]),.dout(n17412),.clk(gclk));
	jxor g17115(.dina(w_n16778_0[0]),.dinb(w_n5121_12[0]),.dout(n17413),.clk(gclk));
	jor g17116(.dina(n17413),.dinb(w_n17140_14[2]),.dout(n17414),.clk(gclk));
	jxor g17117(.dina(n17414),.dinb(w_n16789_0[0]),.dout(n17415),.clk(gclk));
	jand g17118(.dina(w_n17411_0[0]),.dinb(w_n5116_9[1]),.dout(n17416),.clk(gclk));
	jor g17119(.dina(w_n17416_0[1]),.dinb(w_n17415_0[1]),.dout(n17417),.clk(gclk));
	jand g17120(.dina(w_n17417_0[2]),.dinb(w_n17412_0[2]),.dout(n17418),.clk(gclk));
	jor g17121(.dina(n17418),.dinb(w_n4499_13[1]),.dout(n17419),.clk(gclk));
	jnot g17122(.din(w_n16794_0[0]),.dout(n17420),.clk(gclk));
	jor g17123(.dina(n17420),.dinb(w_n16792_0[0]),.dout(n17421),.clk(gclk));
	jor g17124(.dina(n17421),.dinb(w_n17140_14[1]),.dout(n17422),.clk(gclk));
	jxor g17125(.dina(n17422),.dinb(w_n16803_0[0]),.dout(n17423),.clk(gclk));
	jand g17126(.dina(w_n17412_0[1]),.dinb(w_n4499_13[0]),.dout(n17424),.clk(gclk));
	jand g17127(.dina(n17424),.dinb(w_n17417_0[1]),.dout(n17425),.clk(gclk));
	jor g17128(.dina(w_n17425_0[1]),.dinb(w_n17423_0[1]),.dout(n17426),.clk(gclk));
	jand g17129(.dina(w_n17426_0[1]),.dinb(w_n17419_0[1]),.dout(n17427),.clk(gclk));
	jor g17130(.dina(w_n17427_0[2]),.dinb(w_n4494_10[2]),.dout(n17428),.clk(gclk));
	jand g17131(.dina(w_n17427_0[1]),.dinb(w_n4494_10[1]),.dout(n17429),.clk(gclk));
	jnot g17132(.din(w_n16806_0[0]),.dout(n17430),.clk(gclk));
	jand g17133(.dina(w_asqrt7_11[2]),.dinb(n17430),.dout(n17431),.clk(gclk));
	jand g17134(.dina(w_n17431_0[1]),.dinb(w_n16811_0[0]),.dout(n17432),.clk(gclk));
	jor g17135(.dina(n17432),.dinb(w_n16810_0[0]),.dout(n17433),.clk(gclk));
	jand g17136(.dina(w_n17431_0[0]),.dinb(w_n16812_0[0]),.dout(n17434),.clk(gclk));
	jnot g17137(.din(n17434),.dout(n17435),.clk(gclk));
	jand g17138(.dina(n17435),.dinb(n17433),.dout(n17436),.clk(gclk));
	jnot g17139(.din(n17436),.dout(n17437),.clk(gclk));
	jor g17140(.dina(w_n17437_0[1]),.dinb(n17429),.dout(n17438),.clk(gclk));
	jand g17141(.dina(w_n17438_0[1]),.dinb(w_n17428_0[1]),.dout(n17439),.clk(gclk));
	jor g17142(.dina(n17439),.dinb(w_n3912_13[1]),.dout(n17440),.clk(gclk));
	jand g17143(.dina(w_n17428_0[0]),.dinb(w_n3912_13[0]),.dout(n17441),.clk(gclk));
	jand g17144(.dina(n17441),.dinb(w_n17438_0[0]),.dout(n17442),.clk(gclk));
	jnot g17145(.din(w_n16814_0[0]),.dout(n17443),.clk(gclk));
	jand g17146(.dina(w_asqrt7_11[1]),.dinb(n17443),.dout(n17444),.clk(gclk));
	jand g17147(.dina(w_n17444_0[1]),.dinb(w_n16821_0[0]),.dout(n17445),.clk(gclk));
	jor g17148(.dina(n17445),.dinb(w_n16819_0[0]),.dout(n17446),.clk(gclk));
	jand g17149(.dina(w_n17444_0[0]),.dinb(w_n16822_0[0]),.dout(n17447),.clk(gclk));
	jnot g17150(.din(n17447),.dout(n17448),.clk(gclk));
	jand g17151(.dina(n17448),.dinb(n17446),.dout(n17449),.clk(gclk));
	jnot g17152(.din(n17449),.dout(n17450),.clk(gclk));
	jor g17153(.dina(w_n17450_0[1]),.dinb(w_n17442_0[1]),.dout(n17451),.clk(gclk));
	jand g17154(.dina(n17451),.dinb(w_n17440_0[1]),.dout(n17452),.clk(gclk));
	jor g17155(.dina(w_n17452_0[1]),.dinb(w_n3907_10[2]),.dout(n17453),.clk(gclk));
	jxor g17156(.dina(w_n16823_0[0]),.dinb(w_n3912_12[2]),.dout(n17454),.clk(gclk));
	jor g17157(.dina(n17454),.dinb(w_n17140_14[0]),.dout(n17455),.clk(gclk));
	jxor g17158(.dina(n17455),.dinb(w_n16834_0[0]),.dout(n17456),.clk(gclk));
	jand g17159(.dina(w_n17452_0[0]),.dinb(w_n3907_10[1]),.dout(n17457),.clk(gclk));
	jor g17160(.dina(w_n17457_0[1]),.dinb(w_n17456_0[1]),.dout(n17458),.clk(gclk));
	jand g17161(.dina(w_n17458_0[2]),.dinb(w_n17453_0[2]),.dout(n17459),.clk(gclk));
	jor g17162(.dina(n17459),.dinb(w_n3376_14[0]),.dout(n17460),.clk(gclk));
	jnot g17163(.din(w_n16839_0[0]),.dout(n17461),.clk(gclk));
	jor g17164(.dina(n17461),.dinb(w_n16837_0[0]),.dout(n17462),.clk(gclk));
	jor g17165(.dina(n17462),.dinb(w_n17140_13[2]),.dout(n17463),.clk(gclk));
	jxor g17166(.dina(n17463),.dinb(w_n16848_0[0]),.dout(n17464),.clk(gclk));
	jand g17167(.dina(w_n17453_0[1]),.dinb(w_n3376_13[2]),.dout(n17465),.clk(gclk));
	jand g17168(.dina(n17465),.dinb(w_n17458_0[1]),.dout(n17466),.clk(gclk));
	jor g17169(.dina(w_n17466_0[1]),.dinb(w_n17464_0[1]),.dout(n17467),.clk(gclk));
	jand g17170(.dina(w_n17467_0[1]),.dinb(w_n17460_0[1]),.dout(n17468),.clk(gclk));
	jor g17171(.dina(w_n17468_0[2]),.dinb(w_n3371_11[1]),.dout(n17469),.clk(gclk));
	jand g17172(.dina(w_n17468_0[1]),.dinb(w_n3371_11[0]),.dout(n17470),.clk(gclk));
	jnot g17173(.din(w_n16851_0[0]),.dout(n17471),.clk(gclk));
	jand g17174(.dina(w_asqrt7_11[0]),.dinb(n17471),.dout(n17472),.clk(gclk));
	jand g17175(.dina(w_n17472_0[1]),.dinb(w_n16856_0[0]),.dout(n17473),.clk(gclk));
	jor g17176(.dina(n17473),.dinb(w_n16855_0[0]),.dout(n17474),.clk(gclk));
	jand g17177(.dina(w_n17472_0[0]),.dinb(w_n16857_0[0]),.dout(n17475),.clk(gclk));
	jnot g17178(.din(n17475),.dout(n17476),.clk(gclk));
	jand g17179(.dina(n17476),.dinb(n17474),.dout(n17477),.clk(gclk));
	jnot g17180(.din(n17477),.dout(n17478),.clk(gclk));
	jor g17181(.dina(w_n17478_0[1]),.dinb(n17470),.dout(n17479),.clk(gclk));
	jand g17182(.dina(w_n17479_0[1]),.dinb(w_n17469_0[1]),.dout(n17480),.clk(gclk));
	jor g17183(.dina(n17480),.dinb(w_n2875_14[0]),.dout(n17481),.clk(gclk));
	jand g17184(.dina(w_n17469_0[0]),.dinb(w_n2875_13[2]),.dout(n17482),.clk(gclk));
	jand g17185(.dina(n17482),.dinb(w_n17479_0[0]),.dout(n17483),.clk(gclk));
	jnot g17186(.din(w_n16859_0[0]),.dout(n17484),.clk(gclk));
	jand g17187(.dina(w_asqrt7_10[2]),.dinb(n17484),.dout(n17485),.clk(gclk));
	jand g17188(.dina(w_n17485_0[1]),.dinb(w_n16866_0[0]),.dout(n17486),.clk(gclk));
	jor g17189(.dina(n17486),.dinb(w_n16864_0[0]),.dout(n17487),.clk(gclk));
	jand g17190(.dina(w_n17485_0[0]),.dinb(w_n16867_0[0]),.dout(n17488),.clk(gclk));
	jnot g17191(.din(n17488),.dout(n17489),.clk(gclk));
	jand g17192(.dina(n17489),.dinb(n17487),.dout(n17490),.clk(gclk));
	jnot g17193(.din(n17490),.dout(n17491),.clk(gclk));
	jor g17194(.dina(w_n17491_0[1]),.dinb(w_n17483_0[1]),.dout(n17492),.clk(gclk));
	jand g17195(.dina(n17492),.dinb(w_n17481_0[1]),.dout(n17493),.clk(gclk));
	jor g17196(.dina(w_n17493_0[1]),.dinb(w_n2870_11[1]),.dout(n17494),.clk(gclk));
	jxor g17197(.dina(w_n16868_0[0]),.dinb(w_n2875_13[1]),.dout(n17495),.clk(gclk));
	jor g17198(.dina(n17495),.dinb(w_n17140_13[1]),.dout(n17496),.clk(gclk));
	jxor g17199(.dina(n17496),.dinb(w_n16879_0[0]),.dout(n17497),.clk(gclk));
	jand g17200(.dina(w_n17493_0[0]),.dinb(w_n2870_11[0]),.dout(n17498),.clk(gclk));
	jor g17201(.dina(w_n17498_0[1]),.dinb(w_n17497_0[1]),.dout(n17499),.clk(gclk));
	jand g17202(.dina(w_n17499_0[2]),.dinb(w_n17494_0[2]),.dout(n17500),.clk(gclk));
	jor g17203(.dina(n17500),.dinb(w_n2425_14[1]),.dout(n17501),.clk(gclk));
	jnot g17204(.din(w_n16884_0[0]),.dout(n17502),.clk(gclk));
	jor g17205(.dina(n17502),.dinb(w_n16882_0[0]),.dout(n17503),.clk(gclk));
	jor g17206(.dina(n17503),.dinb(w_n17140_13[0]),.dout(n17504),.clk(gclk));
	jxor g17207(.dina(n17504),.dinb(w_n16893_0[0]),.dout(n17505),.clk(gclk));
	jand g17208(.dina(w_n17494_0[1]),.dinb(w_n2425_14[0]),.dout(n17506),.clk(gclk));
	jand g17209(.dina(n17506),.dinb(w_n17499_0[1]),.dout(n17507),.clk(gclk));
	jor g17210(.dina(w_n17507_0[1]),.dinb(w_n17505_0[1]),.dout(n17508),.clk(gclk));
	jand g17211(.dina(w_n17508_0[1]),.dinb(w_n17501_0[1]),.dout(n17509),.clk(gclk));
	jor g17212(.dina(w_n17509_0[2]),.dinb(w_n2420_12[1]),.dout(n17510),.clk(gclk));
	jand g17213(.dina(w_n17509_0[1]),.dinb(w_n2420_12[0]),.dout(n17511),.clk(gclk));
	jnot g17214(.din(w_n16896_0[0]),.dout(n17512),.clk(gclk));
	jand g17215(.dina(w_asqrt7_10[1]),.dinb(n17512),.dout(n17513),.clk(gclk));
	jand g17216(.dina(w_n17513_0[1]),.dinb(w_n16901_0[0]),.dout(n17514),.clk(gclk));
	jor g17217(.dina(n17514),.dinb(w_n16900_0[0]),.dout(n17515),.clk(gclk));
	jand g17218(.dina(w_n17513_0[0]),.dinb(w_n16902_0[0]),.dout(n17516),.clk(gclk));
	jnot g17219(.din(n17516),.dout(n17517),.clk(gclk));
	jand g17220(.dina(n17517),.dinb(n17515),.dout(n17518),.clk(gclk));
	jnot g17221(.din(n17518),.dout(n17519),.clk(gclk));
	jor g17222(.dina(w_n17519_0[1]),.dinb(n17511),.dout(n17520),.clk(gclk));
	jand g17223(.dina(w_n17520_0[1]),.dinb(w_n17510_0[1]),.dout(n17521),.clk(gclk));
	jor g17224(.dina(n17521),.dinb(w_n2010_14[1]),.dout(n17522),.clk(gclk));
	jand g17225(.dina(w_n17510_0[0]),.dinb(w_n2010_14[0]),.dout(n17523),.clk(gclk));
	jand g17226(.dina(n17523),.dinb(w_n17520_0[0]),.dout(n17524),.clk(gclk));
	jnot g17227(.din(w_n16904_0[0]),.dout(n17525),.clk(gclk));
	jand g17228(.dina(w_asqrt7_10[0]),.dinb(n17525),.dout(n17526),.clk(gclk));
	jand g17229(.dina(w_n17526_0[1]),.dinb(w_n16911_0[0]),.dout(n17527),.clk(gclk));
	jor g17230(.dina(n17527),.dinb(w_n16909_0[0]),.dout(n17528),.clk(gclk));
	jand g17231(.dina(w_n17526_0[0]),.dinb(w_n16912_0[0]),.dout(n17529),.clk(gclk));
	jnot g17232(.din(n17529),.dout(n17530),.clk(gclk));
	jand g17233(.dina(n17530),.dinb(n17528),.dout(n17531),.clk(gclk));
	jnot g17234(.din(n17531),.dout(n17532),.clk(gclk));
	jor g17235(.dina(w_n17532_0[1]),.dinb(w_n17524_0[1]),.dout(n17533),.clk(gclk));
	jand g17236(.dina(n17533),.dinb(w_n17522_0[1]),.dout(n17534),.clk(gclk));
	jor g17237(.dina(w_n17534_0[1]),.dinb(w_n2005_12[1]),.dout(n17535),.clk(gclk));
	jxor g17238(.dina(w_n16913_0[0]),.dinb(w_n2010_13[2]),.dout(n17536),.clk(gclk));
	jor g17239(.dina(n17536),.dinb(w_n17140_12[2]),.dout(n17537),.clk(gclk));
	jxor g17240(.dina(n17537),.dinb(w_n16924_0[0]),.dout(n17538),.clk(gclk));
	jand g17241(.dina(w_n17534_0[0]),.dinb(w_n2005_12[0]),.dout(n17539),.clk(gclk));
	jor g17242(.dina(w_n17539_0[1]),.dinb(w_n17538_0[1]),.dout(n17540),.clk(gclk));
	jand g17243(.dina(w_n17540_0[2]),.dinb(w_n17535_0[2]),.dout(n17541),.clk(gclk));
	jor g17244(.dina(n17541),.dinb(w_n1646_15[0]),.dout(n17542),.clk(gclk));
	jnot g17245(.din(w_n16929_0[0]),.dout(n17543),.clk(gclk));
	jor g17246(.dina(n17543),.dinb(w_n16927_0[0]),.dout(n17544),.clk(gclk));
	jor g17247(.dina(n17544),.dinb(w_n17140_12[1]),.dout(n17545),.clk(gclk));
	jxor g17248(.dina(n17545),.dinb(w_n16938_0[0]),.dout(n17546),.clk(gclk));
	jand g17249(.dina(w_n17535_0[1]),.dinb(w_n1646_14[2]),.dout(n17547),.clk(gclk));
	jand g17250(.dina(n17547),.dinb(w_n17540_0[1]),.dout(n17548),.clk(gclk));
	jor g17251(.dina(w_n17548_0[1]),.dinb(w_n17546_0[1]),.dout(n17549),.clk(gclk));
	jand g17252(.dina(w_n17549_0[1]),.dinb(w_n17542_0[1]),.dout(n17550),.clk(gclk));
	jor g17253(.dina(w_n17550_0[2]),.dinb(w_n1641_13[0]),.dout(n17551),.clk(gclk));
	jand g17254(.dina(w_n17550_0[1]),.dinb(w_n1641_12[2]),.dout(n17552),.clk(gclk));
	jnot g17255(.din(w_n16941_0[0]),.dout(n17553),.clk(gclk));
	jand g17256(.dina(w_asqrt7_9[2]),.dinb(n17553),.dout(n17554),.clk(gclk));
	jand g17257(.dina(w_n17554_0[1]),.dinb(w_n16946_0[0]),.dout(n17555),.clk(gclk));
	jor g17258(.dina(n17555),.dinb(w_n16945_0[0]),.dout(n17556),.clk(gclk));
	jand g17259(.dina(w_n17554_0[0]),.dinb(w_n16947_0[0]),.dout(n17557),.clk(gclk));
	jnot g17260(.din(n17557),.dout(n17558),.clk(gclk));
	jand g17261(.dina(n17558),.dinb(n17556),.dout(n17559),.clk(gclk));
	jnot g17262(.din(n17559),.dout(n17560),.clk(gclk));
	jor g17263(.dina(w_n17560_0[1]),.dinb(n17552),.dout(n17561),.clk(gclk));
	jand g17264(.dina(w_n17561_0[1]),.dinb(w_n17551_0[1]),.dout(n17562),.clk(gclk));
	jor g17265(.dina(n17562),.dinb(w_n1317_15[0]),.dout(n17563),.clk(gclk));
	jand g17266(.dina(w_n17551_0[0]),.dinb(w_n1317_14[2]),.dout(n17564),.clk(gclk));
	jand g17267(.dina(n17564),.dinb(w_n17561_0[0]),.dout(n17565),.clk(gclk));
	jnot g17268(.din(w_n16949_0[0]),.dout(n17566),.clk(gclk));
	jand g17269(.dina(w_asqrt7_9[1]),.dinb(n17566),.dout(n17567),.clk(gclk));
	jand g17270(.dina(w_n17567_0[1]),.dinb(w_n16956_0[0]),.dout(n17568),.clk(gclk));
	jor g17271(.dina(n17568),.dinb(w_n16954_0[0]),.dout(n17569),.clk(gclk));
	jand g17272(.dina(w_n17567_0[0]),.dinb(w_n16957_0[0]),.dout(n17570),.clk(gclk));
	jnot g17273(.din(n17570),.dout(n17571),.clk(gclk));
	jand g17274(.dina(n17571),.dinb(n17569),.dout(n17572),.clk(gclk));
	jnot g17275(.din(n17572),.dout(n17573),.clk(gclk));
	jor g17276(.dina(w_n17573_0[1]),.dinb(w_n17565_0[1]),.dout(n17574),.clk(gclk));
	jand g17277(.dina(n17574),.dinb(w_n17563_0[1]),.dout(n17575),.clk(gclk));
	jor g17278(.dina(w_n17575_0[1]),.dinb(w_n1312_13[0]),.dout(n17576),.clk(gclk));
	jxor g17279(.dina(w_n16958_0[0]),.dinb(w_n1317_14[1]),.dout(n17577),.clk(gclk));
	jor g17280(.dina(n17577),.dinb(w_n17140_12[0]),.dout(n17578),.clk(gclk));
	jxor g17281(.dina(n17578),.dinb(w_n16969_0[0]),.dout(n17579),.clk(gclk));
	jand g17282(.dina(w_n17575_0[0]),.dinb(w_n1312_12[2]),.dout(n17580),.clk(gclk));
	jor g17283(.dina(w_n17580_0[1]),.dinb(w_n17579_0[1]),.dout(n17581),.clk(gclk));
	jand g17284(.dina(w_n17581_0[2]),.dinb(w_n17576_0[2]),.dout(n17582),.clk(gclk));
	jor g17285(.dina(n17582),.dinb(w_n1039_15[1]),.dout(n17583),.clk(gclk));
	jnot g17286(.din(w_n16974_0[0]),.dout(n17584),.clk(gclk));
	jor g17287(.dina(n17584),.dinb(w_n16972_0[0]),.dout(n17585),.clk(gclk));
	jor g17288(.dina(n17585),.dinb(w_n17140_11[2]),.dout(n17586),.clk(gclk));
	jxor g17289(.dina(n17586),.dinb(w_n16983_0[0]),.dout(n17587),.clk(gclk));
	jand g17290(.dina(w_n17576_0[1]),.dinb(w_n1039_15[0]),.dout(n17588),.clk(gclk));
	jand g17291(.dina(n17588),.dinb(w_n17581_0[1]),.dout(n17589),.clk(gclk));
	jor g17292(.dina(w_n17589_0[1]),.dinb(w_n17587_0[1]),.dout(n17590),.clk(gclk));
	jand g17293(.dina(w_n17590_0[1]),.dinb(w_n17583_0[1]),.dout(n17591),.clk(gclk));
	jor g17294(.dina(w_n17591_0[2]),.dinb(w_n1034_14[0]),.dout(n17592),.clk(gclk));
	jand g17295(.dina(w_n17591_0[1]),.dinb(w_n1034_13[2]),.dout(n17593),.clk(gclk));
	jnot g17296(.din(w_n16986_0[0]),.dout(n17594),.clk(gclk));
	jand g17297(.dina(w_asqrt7_9[0]),.dinb(n17594),.dout(n17595),.clk(gclk));
	jand g17298(.dina(w_n17595_0[1]),.dinb(w_n16991_0[0]),.dout(n17596),.clk(gclk));
	jor g17299(.dina(n17596),.dinb(w_n16990_0[0]),.dout(n17597),.clk(gclk));
	jand g17300(.dina(w_n17595_0[0]),.dinb(w_n16992_0[0]),.dout(n17598),.clk(gclk));
	jnot g17301(.din(n17598),.dout(n17599),.clk(gclk));
	jand g17302(.dina(n17599),.dinb(n17597),.dout(n17600),.clk(gclk));
	jnot g17303(.din(n17600),.dout(n17601),.clk(gclk));
	jor g17304(.dina(w_n17601_0[1]),.dinb(n17593),.dout(n17602),.clk(gclk));
	jand g17305(.dina(w_n17602_0[1]),.dinb(w_n17592_0[1]),.dout(n17603),.clk(gclk));
	jor g17306(.dina(n17603),.dinb(w_n796_15[1]),.dout(n17604),.clk(gclk));
	jand g17307(.dina(w_n17592_0[0]),.dinb(w_n796_15[0]),.dout(n17605),.clk(gclk));
	jand g17308(.dina(n17605),.dinb(w_n17602_0[0]),.dout(n17606),.clk(gclk));
	jnot g17309(.din(w_n16994_0[0]),.dout(n17607),.clk(gclk));
	jand g17310(.dina(w_asqrt7_8[2]),.dinb(n17607),.dout(n17608),.clk(gclk));
	jand g17311(.dina(w_n17608_0[1]),.dinb(w_n17001_0[0]),.dout(n17609),.clk(gclk));
	jor g17312(.dina(n17609),.dinb(w_n16999_0[0]),.dout(n17610),.clk(gclk));
	jand g17313(.dina(w_n17608_0[0]),.dinb(w_n17002_0[0]),.dout(n17611),.clk(gclk));
	jnot g17314(.din(n17611),.dout(n17612),.clk(gclk));
	jand g17315(.dina(n17612),.dinb(n17610),.dout(n17613),.clk(gclk));
	jnot g17316(.din(n17613),.dout(n17614),.clk(gclk));
	jor g17317(.dina(w_n17614_0[1]),.dinb(w_n17606_0[1]),.dout(n17615),.clk(gclk));
	jand g17318(.dina(n17615),.dinb(w_n17604_0[1]),.dout(n17616),.clk(gclk));
	jor g17319(.dina(w_n17616_0[1]),.dinb(w_n791_14[0]),.dout(n17617),.clk(gclk));
	jxor g17320(.dina(w_n17003_0[0]),.dinb(w_n796_14[2]),.dout(n17618),.clk(gclk));
	jor g17321(.dina(n17618),.dinb(w_n17140_11[1]),.dout(n17619),.clk(gclk));
	jxor g17322(.dina(n17619),.dinb(w_n17014_0[0]),.dout(n17620),.clk(gclk));
	jand g17323(.dina(w_n17616_0[0]),.dinb(w_n791_13[2]),.dout(n17621),.clk(gclk));
	jor g17324(.dina(w_n17621_0[1]),.dinb(w_n17620_0[1]),.dout(n17622),.clk(gclk));
	jand g17325(.dina(w_n17622_0[2]),.dinb(w_n17617_0[2]),.dout(n17623),.clk(gclk));
	jor g17326(.dina(n17623),.dinb(w_n595_15[2]),.dout(n17624),.clk(gclk));
	jand g17327(.dina(w_n17617_0[1]),.dinb(w_n595_15[1]),.dout(n17625),.clk(gclk));
	jand g17328(.dina(n17625),.dinb(w_n17622_0[1]),.dout(n17626),.clk(gclk));
	jnot g17329(.din(w_n17017_0[0]),.dout(n17627),.clk(gclk));
	jand g17330(.dina(w_asqrt7_8[1]),.dinb(n17627),.dout(n17628),.clk(gclk));
	jand g17331(.dina(w_n17628_0[1]),.dinb(w_n17024_0[0]),.dout(n17629),.clk(gclk));
	jor g17332(.dina(n17629),.dinb(w_n17022_0[0]),.dout(n17630),.clk(gclk));
	jand g17333(.dina(w_n17628_0[0]),.dinb(w_n17025_0[0]),.dout(n17631),.clk(gclk));
	jnot g17334(.din(n17631),.dout(n17632),.clk(gclk));
	jand g17335(.dina(n17632),.dinb(n17630),.dout(n17633),.clk(gclk));
	jnot g17336(.din(n17633),.dout(n17634),.clk(gclk));
	jor g17337(.dina(w_n17634_0[1]),.dinb(w_n17626_0[1]),.dout(n17635),.clk(gclk));
	jand g17338(.dina(n17635),.dinb(w_n17624_0[1]),.dout(n17636),.clk(gclk));
	jor g17339(.dina(w_n17636_0[2]),.dinb(w_n590_14[2]),.dout(n17637),.clk(gclk));
	jand g17340(.dina(w_n17636_0[1]),.dinb(w_n590_14[1]),.dout(n17638),.clk(gclk));
	jor g17341(.dina(n17638),.dinb(w_n17143_0[1]),.dout(n17639),.clk(gclk));
	jand g17342(.dina(w_n17639_0[1]),.dinb(w_n17637_0[1]),.dout(n17640),.clk(gclk));
	jor g17343(.dina(n17640),.dinb(w_n430_16[0]),.dout(n17641),.clk(gclk));
	jnot g17344(.din(w_n17033_0[0]),.dout(n17642),.clk(gclk));
	jor g17345(.dina(n17642),.dinb(w_n17031_0[0]),.dout(n17643),.clk(gclk));
	jor g17346(.dina(n17643),.dinb(w_n17140_11[0]),.dout(n17644),.clk(gclk));
	jxor g17347(.dina(n17644),.dinb(w_n17042_0[0]),.dout(n17645),.clk(gclk));
	jand g17348(.dina(w_n17637_0[0]),.dinb(w_n430_15[2]),.dout(n17646),.clk(gclk));
	jand g17349(.dina(n17646),.dinb(w_n17639_0[0]),.dout(n17647),.clk(gclk));
	jor g17350(.dina(w_n17647_0[1]),.dinb(w_n17645_0[1]),.dout(n17648),.clk(gclk));
	jand g17351(.dina(w_n17648_0[1]),.dinb(w_n17641_0[1]),.dout(n17649),.clk(gclk));
	jor g17352(.dina(w_n17649_0[1]),.dinb(w_n425_14[2]),.dout(n17650),.clk(gclk));
	jxor g17353(.dina(w_n17044_0[0]),.dinb(w_n430_15[1]),.dout(n17651),.clk(gclk));
	jor g17354(.dina(n17651),.dinb(w_n17140_10[2]),.dout(n17652),.clk(gclk));
	jxor g17355(.dina(n17652),.dinb(w_n17055_0[0]),.dout(n17653),.clk(gclk));
	jand g17356(.dina(w_n17649_0[0]),.dinb(w_n425_14[1]),.dout(n17654),.clk(gclk));
	jor g17357(.dina(w_n17654_0[1]),.dinb(w_n17653_0[1]),.dout(n17655),.clk(gclk));
	jand g17358(.dina(w_n17655_0[2]),.dinb(w_n17650_0[2]),.dout(n17656),.clk(gclk));
	jor g17359(.dina(n17656),.dinb(w_n305_16[1]),.dout(n17657),.clk(gclk));
	jnot g17360(.din(w_n17060_0[0]),.dout(n17658),.clk(gclk));
	jor g17361(.dina(n17658),.dinb(w_n17058_0[0]),.dout(n17659),.clk(gclk));
	jor g17362(.dina(n17659),.dinb(w_n17140_10[1]),.dout(n17660),.clk(gclk));
	jxor g17363(.dina(n17660),.dinb(w_n17069_0[0]),.dout(n17661),.clk(gclk));
	jand g17364(.dina(w_n17650_0[1]),.dinb(w_n305_16[0]),.dout(n17662),.clk(gclk));
	jand g17365(.dina(n17662),.dinb(w_n17655_0[1]),.dout(n17663),.clk(gclk));
	jor g17366(.dina(w_n17663_0[1]),.dinb(w_n17661_0[1]),.dout(n17664),.clk(gclk));
	jand g17367(.dina(w_n17664_0[1]),.dinb(w_n17657_0[1]),.dout(n17665),.clk(gclk));
	jor g17368(.dina(w_n17665_0[2]),.dinb(w_n290_16[0]),.dout(n17666),.clk(gclk));
	jand g17369(.dina(w_n17665_0[1]),.dinb(w_n290_15[2]),.dout(n17667),.clk(gclk));
	jnot g17370(.din(w_n17072_0[0]),.dout(n17668),.clk(gclk));
	jand g17371(.dina(w_asqrt7_8[0]),.dinb(n17668),.dout(n17669),.clk(gclk));
	jand g17372(.dina(w_n17669_0[1]),.dinb(w_n17077_0[0]),.dout(n17670),.clk(gclk));
	jor g17373(.dina(n17670),.dinb(w_n17076_0[0]),.dout(n17671),.clk(gclk));
	jand g17374(.dina(w_n17669_0[0]),.dinb(w_n17078_0[0]),.dout(n17672),.clk(gclk));
	jnot g17375(.din(n17672),.dout(n17673),.clk(gclk));
	jand g17376(.dina(n17673),.dinb(n17671),.dout(n17674),.clk(gclk));
	jnot g17377(.din(n17674),.dout(n17675),.clk(gclk));
	jor g17378(.dina(w_n17675_0[1]),.dinb(n17667),.dout(n17676),.clk(gclk));
	jand g17379(.dina(w_n17676_0[1]),.dinb(w_n17666_0[1]),.dout(n17677),.clk(gclk));
	jor g17380(.dina(n17677),.dinb(w_n223_16[1]),.dout(n17678),.clk(gclk));
	jand g17381(.dina(w_n17666_0[0]),.dinb(w_n223_16[0]),.dout(n17679),.clk(gclk));
	jand g17382(.dina(n17679),.dinb(w_n17676_0[0]),.dout(n17680),.clk(gclk));
	jnot g17383(.din(w_n17080_0[0]),.dout(n17681),.clk(gclk));
	jand g17384(.dina(w_asqrt7_7[2]),.dinb(n17681),.dout(n17682),.clk(gclk));
	jand g17385(.dina(w_n17682_0[1]),.dinb(w_n17087_0[0]),.dout(n17683),.clk(gclk));
	jor g17386(.dina(n17683),.dinb(w_n17085_0[0]),.dout(n17684),.clk(gclk));
	jand g17387(.dina(w_n17682_0[0]),.dinb(w_n17088_0[0]),.dout(n17685),.clk(gclk));
	jnot g17388(.din(n17685),.dout(n17686),.clk(gclk));
	jand g17389(.dina(n17686),.dinb(n17684),.dout(n17687),.clk(gclk));
	jnot g17390(.din(n17687),.dout(n17688),.clk(gclk));
	jor g17391(.dina(w_n17688_0[1]),.dinb(w_n17680_0[1]),.dout(n17689),.clk(gclk));
	jand g17392(.dina(n17689),.dinb(w_n17678_0[1]),.dout(n17690),.clk(gclk));
	jor g17393(.dina(w_n17690_0[2]),.dinb(w_n199_18[1]),.dout(n17691),.clk(gclk));
	jand g17394(.dina(w_n17690_0[1]),.dinb(w_n199_18[0]),.dout(n17692),.clk(gclk));
	jxor g17395(.dina(w_n17089_0[0]),.dinb(w_n223_15[2]),.dout(n17693),.clk(gclk));
	jor g17396(.dina(n17693),.dinb(w_n17140_10[0]),.dout(n17694),.clk(gclk));
	jxor g17397(.dina(n17694),.dinb(w_n17100_0[0]),.dout(n17695),.clk(gclk));
	jor g17398(.dina(w_n17695_0[1]),.dinb(n17692),.dout(n17696),.clk(gclk));
	jand g17399(.dina(n17696),.dinb(n17691),.dout(n17697),.clk(gclk));
	jnot g17400(.din(w_n17105_0[0]),.dout(n17698),.clk(gclk));
	jor g17401(.dina(n17698),.dinb(w_n17103_0[0]),.dout(n17699),.clk(gclk));
	jor g17402(.dina(n17699),.dinb(w_n17140_9[2]),.dout(n17700),.clk(gclk));
	jxor g17403(.dina(n17700),.dinb(w_n17114_0[0]),.dout(n17701),.clk(gclk));
	jand g17404(.dina(w_asqrt7_7[1]),.dinb(w_n17128_0[1]),.dout(n17702),.clk(gclk));
	jand g17405(.dina(w_n17702_0[1]),.dinb(w_n17116_1[0]),.dout(n17703),.clk(gclk));
	jor g17406(.dina(n17703),.dinb(w_n17162_0[0]),.dout(n17704),.clk(gclk));
	jor g17407(.dina(n17704),.dinb(w_n17701_0[2]),.dout(n17705),.clk(gclk));
	jor g17408(.dina(n17705),.dinb(w_n17697_0[2]),.dout(n17706),.clk(gclk));
	jand g17409(.dina(n17706),.dinb(w_n194_17[1]),.dout(n17707),.clk(gclk));
	jand g17410(.dina(w_n17701_0[1]),.dinb(w_n17697_0[1]),.dout(n17708),.clk(gclk));
	jor g17411(.dina(w_n17702_0[0]),.dinb(w_n17116_0[2]),.dout(n17709),.clk(gclk));
	jand g17412(.dina(w_n17128_0[0]),.dinb(w_n17116_0[1]),.dout(n17710),.clk(gclk));
	jor g17413(.dina(n17710),.dinb(w_n194_17[0]),.dout(n17711),.clk(gclk));
	jnot g17414(.din(n17711),.dout(n17712),.clk(gclk));
	jand g17415(.dina(n17712),.dinb(n17709),.dout(n17713),.clk(gclk));
	jor g17416(.dina(w_n17713_0[1]),.dinb(w_n17708_0[2]),.dout(n17716),.clk(gclk));
	jor g17417(.dina(n17716),.dinb(w_n17707_0[1]),.dout(asqrt_fa_7),.clk(gclk));
	jxor g17418(.dina(w_n17636_0[0]),.dinb(w_n590_14[0]),.dout(n17718),.clk(gclk));
	jand g17419(.dina(n17718),.dinb(w_asqrt6_31),.dout(n17719),.clk(gclk));
	jxor g17420(.dina(n17719),.dinb(w_n17143_0[0]),.dout(n17720),.clk(gclk));
	jand g17421(.dina(w_asqrt6_30[2]),.dinb(w_a12_0[0]),.dout(n17721),.clk(gclk));
	jnot g17422(.din(w_a10_0[1]),.dout(n17722),.clk(gclk));
	jnot g17423(.din(w_a11_0[1]),.dout(n17723),.clk(gclk));
	jand g17424(.dina(w_n17145_1[0]),.dinb(w_n17723_0[1]),.dout(n17724),.clk(gclk));
	jand g17425(.dina(n17724),.dinb(w_n17722_1[1]),.dout(n17725),.clk(gclk));
	jor g17426(.dina(n17725),.dinb(n17721),.dout(n17726),.clk(gclk));
	jand g17427(.dina(w_n17726_0[2]),.dinb(w_asqrt7_7[0]),.dout(n17727),.clk(gclk));
	jand g17428(.dina(w_asqrt6_30[1]),.dinb(w_n17145_0[2]),.dout(n17728),.clk(gclk));
	jxor g17429(.dina(w_n17728_0[1]),.dinb(w_n17146_0[1]),.dout(n17729),.clk(gclk));
	jor g17430(.dina(w_n17726_0[1]),.dinb(w_asqrt7_6[2]),.dout(n17730),.clk(gclk));
	jand g17431(.dina(n17730),.dinb(w_n17729_0[1]),.dout(n17731),.clk(gclk));
	jor g17432(.dina(w_n17731_0[1]),.dinb(w_n17727_0[1]),.dout(n17732),.clk(gclk));
	jand g17433(.dina(n17732),.dinb(w_asqrt8_12[0]),.dout(n17733),.clk(gclk));
	jor g17434(.dina(w_n17727_0[0]),.dinb(w_asqrt8_11[2]),.dout(n17734),.clk(gclk));
	jor g17435(.dina(n17734),.dinb(w_n17731_0[0]),.dout(n17735),.clk(gclk));
	jand g17436(.dina(w_n17728_0[0]),.dinb(w_n17146_0[0]),.dout(n17736),.clk(gclk));
	jnot g17437(.din(w_n17707_0[0]),.dout(n17737),.clk(gclk));
	jnot g17438(.din(w_n17708_0[1]),.dout(n17738),.clk(gclk));
	jnot g17439(.din(w_n17713_0[0]),.dout(n17739),.clk(gclk));
	jand g17440(.dina(n17739),.dinb(w_asqrt7_6[1]),.dout(n17740),.clk(gclk));
	jand g17441(.dina(n17740),.dinb(n17738),.dout(n17741),.clk(gclk));
	jand g17442(.dina(n17741),.dinb(n17737),.dout(n17742),.clk(gclk));
	jor g17443(.dina(n17742),.dinb(n17736),.dout(n17743),.clk(gclk));
	jxor g17444(.dina(n17743),.dinb(w_n16523_0[1]),.dout(n17744),.clk(gclk));
	jand g17445(.dina(w_n17744_0[1]),.dinb(w_n17735_0[1]),.dout(n17745),.clk(gclk));
	jor g17446(.dina(n17745),.dinb(w_n17733_0[1]),.dout(n17746),.clk(gclk));
	jand g17447(.dina(w_n17746_0[2]),.dinb(w_asqrt9_7[0]),.dout(n17747),.clk(gclk));
	jor g17448(.dina(w_n17746_0[1]),.dinb(w_asqrt9_6[2]),.dout(n17748),.clk(gclk));
	jxor g17449(.dina(w_n17150_0[0]),.dinb(w_n17135_4[1]),.dout(n17749),.clk(gclk));
	jand g17450(.dina(n17749),.dinb(w_asqrt6_30[0]),.dout(n17750),.clk(gclk));
	jxor g17451(.dina(n17750),.dinb(w_n17153_0[0]),.dout(n17751),.clk(gclk));
	jnot g17452(.din(w_n17751_0[1]),.dout(n17752),.clk(gclk));
	jand g17453(.dina(n17752),.dinb(n17748),.dout(n17753),.clk(gclk));
	jor g17454(.dina(w_n17753_0[1]),.dinb(w_n17747_0[1]),.dout(n17754),.clk(gclk));
	jand g17455(.dina(n17754),.dinb(w_asqrt10_12[0]),.dout(n17755),.clk(gclk));
	jnot g17456(.din(w_n17159_0[0]),.dout(n17756),.clk(gclk));
	jand g17457(.dina(n17756),.dinb(w_n17157_0[0]),.dout(n17757),.clk(gclk));
	jand g17458(.dina(n17757),.dinb(w_asqrt6_29[2]),.dout(n17758),.clk(gclk));
	jxor g17459(.dina(n17758),.dinb(w_n17167_0[0]),.dout(n17759),.clk(gclk));
	jnot g17460(.din(n17759),.dout(n17760),.clk(gclk));
	jor g17461(.dina(w_n17747_0[0]),.dinb(w_asqrt10_11[2]),.dout(n17761),.clk(gclk));
	jor g17462(.dina(n17761),.dinb(w_n17753_0[0]),.dout(n17762),.clk(gclk));
	jand g17463(.dina(w_n17762_0[1]),.dinb(w_n17760_0[1]),.dout(n17763),.clk(gclk));
	jor g17464(.dina(w_n17763_0[1]),.dinb(w_n17755_0[1]),.dout(n17764),.clk(gclk));
	jand g17465(.dina(w_n17764_0[2]),.dinb(w_asqrt11_7[0]),.dout(n17765),.clk(gclk));
	jor g17466(.dina(w_n17764_0[1]),.dinb(w_asqrt11_6[2]),.dout(n17766),.clk(gclk));
	jnot g17467(.din(w_n17174_0[0]),.dout(n17767),.clk(gclk));
	jxor g17468(.dina(w_n17169_0[0]),.dinb(w_n15950_4[2]),.dout(n17768),.clk(gclk));
	jand g17469(.dina(n17768),.dinb(w_asqrt6_29[1]),.dout(n17769),.clk(gclk));
	jxor g17470(.dina(n17769),.dinb(n17767),.dout(n17770),.clk(gclk));
	jand g17471(.dina(w_n17770_0[1]),.dinb(n17766),.dout(n17771),.clk(gclk));
	jor g17472(.dina(w_n17771_0[1]),.dinb(w_n17765_0[1]),.dout(n17772),.clk(gclk));
	jand g17473(.dina(n17772),.dinb(w_asqrt12_12[0]),.dout(n17773),.clk(gclk));
	jor g17474(.dina(w_n17765_0[0]),.dinb(w_asqrt12_11[2]),.dout(n17774),.clk(gclk));
	jor g17475(.dina(n17774),.dinb(w_n17771_0[0]),.dout(n17775),.clk(gclk));
	jnot g17476(.din(w_n17181_0[0]),.dout(n17776),.clk(gclk));
	jnot g17477(.din(w_n17183_0[0]),.dout(n17777),.clk(gclk));
	jand g17478(.dina(w_asqrt6_29[0]),.dinb(w_n17177_0[0]),.dout(n17778),.clk(gclk));
	jand g17479(.dina(w_n17778_0[1]),.dinb(n17777),.dout(n17779),.clk(gclk));
	jor g17480(.dina(n17779),.dinb(n17776),.dout(n17780),.clk(gclk));
	jnot g17481(.din(w_n17184_0[0]),.dout(n17781),.clk(gclk));
	jand g17482(.dina(w_n17778_0[0]),.dinb(n17781),.dout(n17782),.clk(gclk));
	jnot g17483(.din(n17782),.dout(n17783),.clk(gclk));
	jand g17484(.dina(n17783),.dinb(n17780),.dout(n17784),.clk(gclk));
	jand g17485(.dina(w_n17784_0[1]),.dinb(w_n17775_0[1]),.dout(n17785),.clk(gclk));
	jor g17486(.dina(n17785),.dinb(w_n17773_0[1]),.dout(n17786),.clk(gclk));
	jand g17487(.dina(w_n17786_0[2]),.dinb(w_asqrt13_7[1]),.dout(n17787),.clk(gclk));
	jor g17488(.dina(w_n17786_0[1]),.dinb(w_asqrt13_7[0]),.dout(n17788),.clk(gclk));
	jxor g17489(.dina(w_n17185_0[0]),.dinb(w_n14816_5[1]),.dout(n17789),.clk(gclk));
	jand g17490(.dina(n17789),.dinb(w_asqrt6_28[2]),.dout(n17790),.clk(gclk));
	jxor g17491(.dina(n17790),.dinb(w_n17190_0[0]),.dout(n17791),.clk(gclk));
	jand g17492(.dina(w_n17791_0[1]),.dinb(n17788),.dout(n17792),.clk(gclk));
	jor g17493(.dina(w_n17792_0[1]),.dinb(w_n17787_0[1]),.dout(n17793),.clk(gclk));
	jand g17494(.dina(n17793),.dinb(w_asqrt14_12[0]),.dout(n17794),.clk(gclk));
	jnot g17495(.din(w_n17196_0[0]),.dout(n17795),.clk(gclk));
	jand g17496(.dina(n17795),.dinb(w_n17194_0[0]),.dout(n17796),.clk(gclk));
	jand g17497(.dina(n17796),.dinb(w_asqrt6_28[1]),.dout(n17797),.clk(gclk));
	jxor g17498(.dina(n17797),.dinb(w_n17205_0[0]),.dout(n17798),.clk(gclk));
	jnot g17499(.din(n17798),.dout(n17799),.clk(gclk));
	jor g17500(.dina(w_n17787_0[0]),.dinb(w_asqrt14_11[2]),.dout(n17800),.clk(gclk));
	jor g17501(.dina(n17800),.dinb(w_n17792_0[0]),.dout(n17801),.clk(gclk));
	jand g17502(.dina(w_n17801_0[1]),.dinb(w_n17799_0[1]),.dout(n17802),.clk(gclk));
	jor g17503(.dina(w_n17802_0[1]),.dinb(w_n17794_0[1]),.dout(n17803),.clk(gclk));
	jand g17504(.dina(w_n17803_0[2]),.dinb(w_asqrt15_7[1]),.dout(n17804),.clk(gclk));
	jor g17505(.dina(w_n17803_0[1]),.dinb(w_asqrt15_7[0]),.dout(n17805),.clk(gclk));
	jxor g17506(.dina(w_n17207_0[0]),.dinb(w_n13718_5[1]),.dout(n17806),.clk(gclk));
	jand g17507(.dina(n17806),.dinb(w_asqrt6_28[0]),.dout(n17807),.clk(gclk));
	jxor g17508(.dina(n17807),.dinb(w_n17213_0[0]),.dout(n17808),.clk(gclk));
	jand g17509(.dina(w_n17808_0[1]),.dinb(n17805),.dout(n17809),.clk(gclk));
	jor g17510(.dina(w_n17809_0[1]),.dinb(w_n17804_0[1]),.dout(n17810),.clk(gclk));
	jand g17511(.dina(n17810),.dinb(w_asqrt16_12[0]),.dout(n17811),.clk(gclk));
	jor g17512(.dina(w_n17804_0[0]),.dinb(w_asqrt16_11[2]),.dout(n17812),.clk(gclk));
	jor g17513(.dina(n17812),.dinb(w_n17809_0[0]),.dout(n17813),.clk(gclk));
	jnot g17514(.din(w_n17221_0[0]),.dout(n17814),.clk(gclk));
	jnot g17515(.din(w_n17223_0[0]),.dout(n17815),.clk(gclk));
	jand g17516(.dina(w_asqrt6_27[2]),.dinb(w_n17217_0[0]),.dout(n17816),.clk(gclk));
	jand g17517(.dina(w_n17816_0[1]),.dinb(n17815),.dout(n17817),.clk(gclk));
	jor g17518(.dina(n17817),.dinb(n17814),.dout(n17818),.clk(gclk));
	jnot g17519(.din(w_n17224_0[0]),.dout(n17819),.clk(gclk));
	jand g17520(.dina(w_n17816_0[0]),.dinb(n17819),.dout(n17820),.clk(gclk));
	jnot g17521(.din(n17820),.dout(n17821),.clk(gclk));
	jand g17522(.dina(n17821),.dinb(n17818),.dout(n17822),.clk(gclk));
	jand g17523(.dina(w_n17822_0[1]),.dinb(w_n17813_0[1]),.dout(n17823),.clk(gclk));
	jor g17524(.dina(n17823),.dinb(w_n17811_0[1]),.dout(n17824),.clk(gclk));
	jand g17525(.dina(w_n17824_0[1]),.dinb(w_asqrt17_7[2]),.dout(n17825),.clk(gclk));
	jxor g17526(.dina(w_n17225_0[0]),.dinb(w_n12670_5[2]),.dout(n17826),.clk(gclk));
	jand g17527(.dina(n17826),.dinb(w_asqrt6_27[1]),.dout(n17827),.clk(gclk));
	jxor g17528(.dina(n17827),.dinb(w_n17232_0[0]),.dout(n17828),.clk(gclk));
	jnot g17529(.din(n17828),.dout(n17829),.clk(gclk));
	jor g17530(.dina(w_n17824_0[0]),.dinb(w_asqrt17_7[1]),.dout(n17830),.clk(gclk));
	jand g17531(.dina(w_n17830_0[1]),.dinb(w_n17829_0[1]),.dout(n17831),.clk(gclk));
	jor g17532(.dina(w_n17831_0[2]),.dinb(w_n17825_0[2]),.dout(n17832),.clk(gclk));
	jand g17533(.dina(n17832),.dinb(w_asqrt18_12[0]),.dout(n17833),.clk(gclk));
	jnot g17534(.din(w_n17237_0[0]),.dout(n17834),.clk(gclk));
	jand g17535(.dina(n17834),.dinb(w_n17235_0[0]),.dout(n17835),.clk(gclk));
	jand g17536(.dina(n17835),.dinb(w_asqrt6_27[0]),.dout(n17836),.clk(gclk));
	jxor g17537(.dina(n17836),.dinb(w_n17245_0[0]),.dout(n17837),.clk(gclk));
	jnot g17538(.din(n17837),.dout(n17838),.clk(gclk));
	jor g17539(.dina(w_n17825_0[1]),.dinb(w_asqrt18_11[2]),.dout(n17839),.clk(gclk));
	jor g17540(.dina(n17839),.dinb(w_n17831_0[1]),.dout(n17840),.clk(gclk));
	jand g17541(.dina(w_n17840_0[1]),.dinb(w_n17838_0[1]),.dout(n17841),.clk(gclk));
	jor g17542(.dina(w_n17841_0[1]),.dinb(w_n17833_0[1]),.dout(n17842),.clk(gclk));
	jand g17543(.dina(w_n17842_0[2]),.dinb(w_asqrt19_7[2]),.dout(n17843),.clk(gclk));
	jor g17544(.dina(w_n17842_0[1]),.dinb(w_asqrt19_7[1]),.dout(n17844),.clk(gclk));
	jnot g17545(.din(w_n17251_0[0]),.dout(n17845),.clk(gclk));
	jnot g17546(.din(w_n17252_0[0]),.dout(n17846),.clk(gclk));
	jand g17547(.dina(w_asqrt6_26[2]),.dinb(w_n17248_0[0]),.dout(n17847),.clk(gclk));
	jand g17548(.dina(w_n17847_0[1]),.dinb(n17846),.dout(n17848),.clk(gclk));
	jor g17549(.dina(n17848),.dinb(n17845),.dout(n17849),.clk(gclk));
	jnot g17550(.din(w_n17253_0[0]),.dout(n17850),.clk(gclk));
	jand g17551(.dina(w_n17847_0[0]),.dinb(n17850),.dout(n17851),.clk(gclk));
	jnot g17552(.din(n17851),.dout(n17852),.clk(gclk));
	jand g17553(.dina(n17852),.dinb(n17849),.dout(n17853),.clk(gclk));
	jand g17554(.dina(w_n17853_0[1]),.dinb(n17844),.dout(n17854),.clk(gclk));
	jor g17555(.dina(w_n17854_0[1]),.dinb(w_n17843_0[1]),.dout(n17855),.clk(gclk));
	jand g17556(.dina(n17855),.dinb(w_asqrt20_12[0]),.dout(n17856),.clk(gclk));
	jor g17557(.dina(w_n17843_0[0]),.dinb(w_asqrt20_11[2]),.dout(n17857),.clk(gclk));
	jor g17558(.dina(n17857),.dinb(w_n17854_0[0]),.dout(n17858),.clk(gclk));
	jnot g17559(.din(w_n17259_0[0]),.dout(n17859),.clk(gclk));
	jnot g17560(.din(w_n17261_0[0]),.dout(n17860),.clk(gclk));
	jand g17561(.dina(w_asqrt6_26[1]),.dinb(w_n17255_0[0]),.dout(n17861),.clk(gclk));
	jand g17562(.dina(w_n17861_0[1]),.dinb(n17860),.dout(n17862),.clk(gclk));
	jor g17563(.dina(n17862),.dinb(n17859),.dout(n17863),.clk(gclk));
	jnot g17564(.din(w_n17262_0[0]),.dout(n17864),.clk(gclk));
	jand g17565(.dina(w_n17861_0[0]),.dinb(n17864),.dout(n17865),.clk(gclk));
	jnot g17566(.din(n17865),.dout(n17866),.clk(gclk));
	jand g17567(.dina(n17866),.dinb(n17863),.dout(n17867),.clk(gclk));
	jand g17568(.dina(w_n17867_0[1]),.dinb(w_n17858_0[1]),.dout(n17868),.clk(gclk));
	jor g17569(.dina(n17868),.dinb(w_n17856_0[1]),.dout(n17869),.clk(gclk));
	jand g17570(.dina(w_n17869_0[1]),.dinb(w_asqrt21_8[0]),.dout(n17870),.clk(gclk));
	jxor g17571(.dina(w_n17263_0[0]),.dinb(w_n10696_6[2]),.dout(n17871),.clk(gclk));
	jand g17572(.dina(n17871),.dinb(w_asqrt6_26[0]),.dout(n17872),.clk(gclk));
	jxor g17573(.dina(n17872),.dinb(w_n17273_0[0]),.dout(n17873),.clk(gclk));
	jnot g17574(.din(n17873),.dout(n17874),.clk(gclk));
	jor g17575(.dina(w_n17869_0[0]),.dinb(w_asqrt21_7[2]),.dout(n17875),.clk(gclk));
	jand g17576(.dina(w_n17875_0[1]),.dinb(w_n17874_0[1]),.dout(n17876),.clk(gclk));
	jor g17577(.dina(w_n17876_0[2]),.dinb(w_n17870_0[2]),.dout(n17877),.clk(gclk));
	jand g17578(.dina(n17877),.dinb(w_asqrt22_12[0]),.dout(n17878),.clk(gclk));
	jnot g17579(.din(w_n17278_0[0]),.dout(n17879),.clk(gclk));
	jand g17580(.dina(n17879),.dinb(w_n17276_0[0]),.dout(n17880),.clk(gclk));
	jand g17581(.dina(n17880),.dinb(w_asqrt6_25[2]),.dout(n17881),.clk(gclk));
	jxor g17582(.dina(n17881),.dinb(w_n17286_0[0]),.dout(n17882),.clk(gclk));
	jnot g17583(.din(n17882),.dout(n17883),.clk(gclk));
	jor g17584(.dina(w_n17870_0[1]),.dinb(w_asqrt22_11[2]),.dout(n17884),.clk(gclk));
	jor g17585(.dina(n17884),.dinb(w_n17876_0[1]),.dout(n17885),.clk(gclk));
	jand g17586(.dina(w_n17885_0[1]),.dinb(w_n17883_0[1]),.dout(n17886),.clk(gclk));
	jor g17587(.dina(w_n17886_0[1]),.dinb(w_n17878_0[1]),.dout(n17887),.clk(gclk));
	jand g17588(.dina(w_n17887_0[2]),.dinb(w_asqrt23_8[0]),.dout(n17888),.clk(gclk));
	jor g17589(.dina(w_n17887_0[1]),.dinb(w_asqrt23_7[2]),.dout(n17889),.clk(gclk));
	jnot g17590(.din(w_n17292_0[0]),.dout(n17890),.clk(gclk));
	jnot g17591(.din(w_n17293_0[0]),.dout(n17891),.clk(gclk));
	jand g17592(.dina(w_asqrt6_25[1]),.dinb(w_n17289_0[0]),.dout(n17892),.clk(gclk));
	jand g17593(.dina(w_n17892_0[1]),.dinb(n17891),.dout(n17893),.clk(gclk));
	jor g17594(.dina(n17893),.dinb(n17890),.dout(n17894),.clk(gclk));
	jnot g17595(.din(w_n17294_0[0]),.dout(n17895),.clk(gclk));
	jand g17596(.dina(w_n17892_0[0]),.dinb(n17895),.dout(n17896),.clk(gclk));
	jnot g17597(.din(n17896),.dout(n17897),.clk(gclk));
	jand g17598(.dina(n17897),.dinb(n17894),.dout(n17898),.clk(gclk));
	jand g17599(.dina(w_n17898_0[1]),.dinb(n17889),.dout(n17899),.clk(gclk));
	jor g17600(.dina(w_n17899_0[1]),.dinb(w_n17888_0[1]),.dout(n17900),.clk(gclk));
	jand g17601(.dina(n17900),.dinb(w_asqrt24_12[0]),.dout(n17901),.clk(gclk));
	jor g17602(.dina(w_n17888_0[0]),.dinb(w_asqrt24_11[2]),.dout(n17902),.clk(gclk));
	jor g17603(.dina(n17902),.dinb(w_n17899_0[0]),.dout(n17903),.clk(gclk));
	jnot g17604(.din(w_n17300_0[0]),.dout(n17904),.clk(gclk));
	jnot g17605(.din(w_n17302_0[0]),.dout(n17905),.clk(gclk));
	jand g17606(.dina(w_asqrt6_25[0]),.dinb(w_n17296_0[0]),.dout(n17906),.clk(gclk));
	jand g17607(.dina(w_n17906_0[1]),.dinb(n17905),.dout(n17907),.clk(gclk));
	jor g17608(.dina(n17907),.dinb(n17904),.dout(n17908),.clk(gclk));
	jnot g17609(.din(w_n17303_0[0]),.dout(n17909),.clk(gclk));
	jand g17610(.dina(w_n17906_0[0]),.dinb(n17909),.dout(n17910),.clk(gclk));
	jnot g17611(.din(n17910),.dout(n17911),.clk(gclk));
	jand g17612(.dina(n17911),.dinb(n17908),.dout(n17912),.clk(gclk));
	jand g17613(.dina(w_n17912_0[1]),.dinb(w_n17903_0[1]),.dout(n17913),.clk(gclk));
	jor g17614(.dina(n17913),.dinb(w_n17901_0[1]),.dout(n17914),.clk(gclk));
	jand g17615(.dina(w_n17914_0[1]),.dinb(w_asqrt25_8[1]),.dout(n17915),.clk(gclk));
	jxor g17616(.dina(w_n17304_0[0]),.dinb(w_n8893_7[1]),.dout(n17916),.clk(gclk));
	jand g17617(.dina(n17916),.dinb(w_asqrt6_24[2]),.dout(n17917),.clk(gclk));
	jxor g17618(.dina(n17917),.dinb(w_n17314_0[0]),.dout(n17918),.clk(gclk));
	jnot g17619(.din(n17918),.dout(n17919),.clk(gclk));
	jor g17620(.dina(w_n17914_0[0]),.dinb(w_asqrt25_8[0]),.dout(n17920),.clk(gclk));
	jand g17621(.dina(w_n17920_0[1]),.dinb(w_n17919_0[1]),.dout(n17921),.clk(gclk));
	jor g17622(.dina(w_n17921_0[2]),.dinb(w_n17915_0[2]),.dout(n17922),.clk(gclk));
	jand g17623(.dina(n17922),.dinb(w_asqrt26_12[0]),.dout(n17923),.clk(gclk));
	jnot g17624(.din(w_n17319_0[0]),.dout(n17924),.clk(gclk));
	jand g17625(.dina(n17924),.dinb(w_n17317_0[0]),.dout(n17925),.clk(gclk));
	jand g17626(.dina(n17925),.dinb(w_asqrt6_24[1]),.dout(n17926),.clk(gclk));
	jxor g17627(.dina(n17926),.dinb(w_n17327_0[0]),.dout(n17927),.clk(gclk));
	jnot g17628(.din(n17927),.dout(n17928),.clk(gclk));
	jor g17629(.dina(w_n17915_0[1]),.dinb(w_asqrt26_11[2]),.dout(n17929),.clk(gclk));
	jor g17630(.dina(n17929),.dinb(w_n17921_0[1]),.dout(n17930),.clk(gclk));
	jand g17631(.dina(w_n17930_0[1]),.dinb(w_n17928_0[1]),.dout(n17931),.clk(gclk));
	jor g17632(.dina(w_n17931_0[1]),.dinb(w_n17923_0[1]),.dout(n17932),.clk(gclk));
	jand g17633(.dina(w_n17932_0[2]),.dinb(w_asqrt27_8[1]),.dout(n17933),.clk(gclk));
	jor g17634(.dina(w_n17932_0[1]),.dinb(w_asqrt27_8[0]),.dout(n17934),.clk(gclk));
	jnot g17635(.din(w_n17333_0[0]),.dout(n17935),.clk(gclk));
	jnot g17636(.din(w_n17334_0[0]),.dout(n17936),.clk(gclk));
	jand g17637(.dina(w_asqrt6_24[0]),.dinb(w_n17330_0[0]),.dout(n17937),.clk(gclk));
	jand g17638(.dina(w_n17937_0[1]),.dinb(n17936),.dout(n17938),.clk(gclk));
	jor g17639(.dina(n17938),.dinb(n17935),.dout(n17939),.clk(gclk));
	jnot g17640(.din(w_n17335_0[0]),.dout(n17940),.clk(gclk));
	jand g17641(.dina(w_n17937_0[0]),.dinb(n17940),.dout(n17941),.clk(gclk));
	jnot g17642(.din(n17941),.dout(n17942),.clk(gclk));
	jand g17643(.dina(n17942),.dinb(n17939),.dout(n17943),.clk(gclk));
	jand g17644(.dina(w_n17943_0[1]),.dinb(n17934),.dout(n17944),.clk(gclk));
	jor g17645(.dina(w_n17944_0[1]),.dinb(w_n17933_0[1]),.dout(n17945),.clk(gclk));
	jand g17646(.dina(n17945),.dinb(w_asqrt28_12[0]),.dout(n17946),.clk(gclk));
	jor g17647(.dina(w_n17933_0[0]),.dinb(w_asqrt28_11[2]),.dout(n17947),.clk(gclk));
	jor g17648(.dina(n17947),.dinb(w_n17944_0[0]),.dout(n17948),.clk(gclk));
	jnot g17649(.din(w_n17341_0[0]),.dout(n17949),.clk(gclk));
	jnot g17650(.din(w_n17343_0[0]),.dout(n17950),.clk(gclk));
	jand g17651(.dina(w_asqrt6_23[2]),.dinb(w_n17337_0[0]),.dout(n17951),.clk(gclk));
	jand g17652(.dina(w_n17951_0[1]),.dinb(n17950),.dout(n17952),.clk(gclk));
	jor g17653(.dina(n17952),.dinb(n17949),.dout(n17953),.clk(gclk));
	jnot g17654(.din(w_n17344_0[0]),.dout(n17954),.clk(gclk));
	jand g17655(.dina(w_n17951_0[0]),.dinb(n17954),.dout(n17955),.clk(gclk));
	jnot g17656(.din(n17955),.dout(n17956),.clk(gclk));
	jand g17657(.dina(n17956),.dinb(n17953),.dout(n17957),.clk(gclk));
	jand g17658(.dina(w_n17957_0[1]),.dinb(w_n17948_0[1]),.dout(n17958),.clk(gclk));
	jor g17659(.dina(n17958),.dinb(w_n17946_0[1]),.dout(n17959),.clk(gclk));
	jand g17660(.dina(w_n17959_0[1]),.dinb(w_asqrt29_8[2]),.dout(n17960),.clk(gclk));
	jxor g17661(.dina(w_n17345_0[0]),.dinb(w_n7260_8[1]),.dout(n17961),.clk(gclk));
	jand g17662(.dina(n17961),.dinb(w_asqrt6_23[1]),.dout(n17962),.clk(gclk));
	jxor g17663(.dina(n17962),.dinb(w_n17355_0[0]),.dout(n17963),.clk(gclk));
	jnot g17664(.din(n17963),.dout(n17964),.clk(gclk));
	jor g17665(.dina(w_n17959_0[0]),.dinb(w_asqrt29_8[1]),.dout(n17965),.clk(gclk));
	jand g17666(.dina(w_n17965_0[1]),.dinb(w_n17964_0[1]),.dout(n17966),.clk(gclk));
	jor g17667(.dina(w_n17966_0[2]),.dinb(w_n17960_0[2]),.dout(n17967),.clk(gclk));
	jand g17668(.dina(n17967),.dinb(w_asqrt30_12[0]),.dout(n17968),.clk(gclk));
	jnot g17669(.din(w_n17360_0[0]),.dout(n17969),.clk(gclk));
	jand g17670(.dina(n17969),.dinb(w_n17358_0[0]),.dout(n17970),.clk(gclk));
	jand g17671(.dina(n17970),.dinb(w_asqrt6_23[0]),.dout(n17971),.clk(gclk));
	jxor g17672(.dina(n17971),.dinb(w_n17368_0[0]),.dout(n17972),.clk(gclk));
	jnot g17673(.din(n17972),.dout(n17973),.clk(gclk));
	jor g17674(.dina(w_n17960_0[1]),.dinb(w_asqrt30_11[2]),.dout(n17974),.clk(gclk));
	jor g17675(.dina(n17974),.dinb(w_n17966_0[1]),.dout(n17975),.clk(gclk));
	jand g17676(.dina(w_n17975_0[1]),.dinb(w_n17973_0[1]),.dout(n17976),.clk(gclk));
	jor g17677(.dina(w_n17976_0[1]),.dinb(w_n17968_0[1]),.dout(n17977),.clk(gclk));
	jand g17678(.dina(w_n17977_0[2]),.dinb(w_asqrt31_8[2]),.dout(n17978),.clk(gclk));
	jor g17679(.dina(w_n17977_0[1]),.dinb(w_asqrt31_8[1]),.dout(n17979),.clk(gclk));
	jnot g17680(.din(w_n17374_0[0]),.dout(n17980),.clk(gclk));
	jnot g17681(.din(w_n17375_0[0]),.dout(n17981),.clk(gclk));
	jand g17682(.dina(w_asqrt6_22[2]),.dinb(w_n17371_0[0]),.dout(n17982),.clk(gclk));
	jand g17683(.dina(w_n17982_0[1]),.dinb(n17981),.dout(n17983),.clk(gclk));
	jor g17684(.dina(n17983),.dinb(n17980),.dout(n17984),.clk(gclk));
	jnot g17685(.din(w_n17376_0[0]),.dout(n17985),.clk(gclk));
	jand g17686(.dina(w_n17982_0[0]),.dinb(n17985),.dout(n17986),.clk(gclk));
	jnot g17687(.din(n17986),.dout(n17987),.clk(gclk));
	jand g17688(.dina(n17987),.dinb(n17984),.dout(n17988),.clk(gclk));
	jand g17689(.dina(w_n17988_0[1]),.dinb(n17979),.dout(n17989),.clk(gclk));
	jor g17690(.dina(w_n17989_0[1]),.dinb(w_n17978_0[1]),.dout(n17990),.clk(gclk));
	jand g17691(.dina(n17990),.dinb(w_asqrt32_12[0]),.dout(n17991),.clk(gclk));
	jor g17692(.dina(w_n17978_0[0]),.dinb(w_asqrt32_11[2]),.dout(n17992),.clk(gclk));
	jor g17693(.dina(n17992),.dinb(w_n17989_0[0]),.dout(n17993),.clk(gclk));
	jnot g17694(.din(w_n17382_0[0]),.dout(n17994),.clk(gclk));
	jnot g17695(.din(w_n17384_0[0]),.dout(n17995),.clk(gclk));
	jand g17696(.dina(w_asqrt6_22[1]),.dinb(w_n17378_0[0]),.dout(n17996),.clk(gclk));
	jand g17697(.dina(w_n17996_0[1]),.dinb(n17995),.dout(n17997),.clk(gclk));
	jor g17698(.dina(n17997),.dinb(n17994),.dout(n17998),.clk(gclk));
	jnot g17699(.din(w_n17385_0[0]),.dout(n17999),.clk(gclk));
	jand g17700(.dina(w_n17996_0[0]),.dinb(n17999),.dout(n18000),.clk(gclk));
	jnot g17701(.din(n18000),.dout(n18001),.clk(gclk));
	jand g17702(.dina(n18001),.dinb(n17998),.dout(n18002),.clk(gclk));
	jand g17703(.dina(w_n18002_0[1]),.dinb(w_n17993_0[1]),.dout(n18003),.clk(gclk));
	jor g17704(.dina(n18003),.dinb(w_n17991_0[1]),.dout(n18004),.clk(gclk));
	jand g17705(.dina(w_n18004_0[1]),.dinb(w_asqrt33_9[0]),.dout(n18005),.clk(gclk));
	jxor g17706(.dina(w_n17386_0[0]),.dinb(w_n5788_9[0]),.dout(n18006),.clk(gclk));
	jand g17707(.dina(n18006),.dinb(w_asqrt6_22[0]),.dout(n18007),.clk(gclk));
	jxor g17708(.dina(n18007),.dinb(w_n17396_0[0]),.dout(n18008),.clk(gclk));
	jnot g17709(.din(n18008),.dout(n18009),.clk(gclk));
	jor g17710(.dina(w_n18004_0[0]),.dinb(w_asqrt33_8[2]),.dout(n18010),.clk(gclk));
	jand g17711(.dina(w_n18010_0[1]),.dinb(w_n18009_0[1]),.dout(n18011),.clk(gclk));
	jor g17712(.dina(w_n18011_0[2]),.dinb(w_n18005_0[2]),.dout(n18012),.clk(gclk));
	jand g17713(.dina(n18012),.dinb(w_asqrt34_12[0]),.dout(n18013),.clk(gclk));
	jnot g17714(.din(w_n17401_0[0]),.dout(n18014),.clk(gclk));
	jand g17715(.dina(n18014),.dinb(w_n17399_0[0]),.dout(n18015),.clk(gclk));
	jand g17716(.dina(n18015),.dinb(w_asqrt6_21[2]),.dout(n18016),.clk(gclk));
	jxor g17717(.dina(n18016),.dinb(w_n17409_0[0]),.dout(n18017),.clk(gclk));
	jnot g17718(.din(n18017),.dout(n18018),.clk(gclk));
	jor g17719(.dina(w_n18005_0[1]),.dinb(w_asqrt34_11[2]),.dout(n18019),.clk(gclk));
	jor g17720(.dina(n18019),.dinb(w_n18011_0[1]),.dout(n18020),.clk(gclk));
	jand g17721(.dina(w_n18020_0[1]),.dinb(w_n18018_0[1]),.dout(n18021),.clk(gclk));
	jor g17722(.dina(w_n18021_0[1]),.dinb(w_n18013_0[1]),.dout(n18022),.clk(gclk));
	jand g17723(.dina(w_n18022_0[2]),.dinb(w_asqrt35_9[0]),.dout(n18023),.clk(gclk));
	jor g17724(.dina(w_n18022_0[1]),.dinb(w_asqrt35_8[2]),.dout(n18024),.clk(gclk));
	jnot g17725(.din(w_n17415_0[0]),.dout(n18025),.clk(gclk));
	jnot g17726(.din(w_n17416_0[0]),.dout(n18026),.clk(gclk));
	jand g17727(.dina(w_asqrt6_21[1]),.dinb(w_n17412_0[0]),.dout(n18027),.clk(gclk));
	jand g17728(.dina(w_n18027_0[1]),.dinb(n18026),.dout(n18028),.clk(gclk));
	jor g17729(.dina(n18028),.dinb(n18025),.dout(n18029),.clk(gclk));
	jnot g17730(.din(w_n17417_0[0]),.dout(n18030),.clk(gclk));
	jand g17731(.dina(w_n18027_0[0]),.dinb(n18030),.dout(n18031),.clk(gclk));
	jnot g17732(.din(n18031),.dout(n18032),.clk(gclk));
	jand g17733(.dina(n18032),.dinb(n18029),.dout(n18033),.clk(gclk));
	jand g17734(.dina(w_n18033_0[1]),.dinb(n18024),.dout(n18034),.clk(gclk));
	jor g17735(.dina(w_n18034_0[1]),.dinb(w_n18023_0[1]),.dout(n18035),.clk(gclk));
	jand g17736(.dina(n18035),.dinb(w_asqrt36_12[0]),.dout(n18036),.clk(gclk));
	jor g17737(.dina(w_n18023_0[0]),.dinb(w_asqrt36_11[2]),.dout(n18037),.clk(gclk));
	jor g17738(.dina(n18037),.dinb(w_n18034_0[0]),.dout(n18038),.clk(gclk));
	jnot g17739(.din(w_n17423_0[0]),.dout(n18039),.clk(gclk));
	jnot g17740(.din(w_n17425_0[0]),.dout(n18040),.clk(gclk));
	jand g17741(.dina(w_asqrt6_21[0]),.dinb(w_n17419_0[0]),.dout(n18041),.clk(gclk));
	jand g17742(.dina(w_n18041_0[1]),.dinb(n18040),.dout(n18042),.clk(gclk));
	jor g17743(.dina(n18042),.dinb(n18039),.dout(n18043),.clk(gclk));
	jnot g17744(.din(w_n17426_0[0]),.dout(n18044),.clk(gclk));
	jand g17745(.dina(w_n18041_0[0]),.dinb(n18044),.dout(n18045),.clk(gclk));
	jnot g17746(.din(n18045),.dout(n18046),.clk(gclk));
	jand g17747(.dina(n18046),.dinb(n18043),.dout(n18047),.clk(gclk));
	jand g17748(.dina(w_n18047_0[1]),.dinb(w_n18038_0[1]),.dout(n18048),.clk(gclk));
	jor g17749(.dina(n18048),.dinb(w_n18036_0[1]),.dout(n18049),.clk(gclk));
	jand g17750(.dina(w_n18049_0[1]),.dinb(w_asqrt37_9[1]),.dout(n18050),.clk(gclk));
	jxor g17751(.dina(w_n17427_0[0]),.dinb(w_n4494_10[0]),.dout(n18051),.clk(gclk));
	jand g17752(.dina(n18051),.dinb(w_asqrt6_20[2]),.dout(n18052),.clk(gclk));
	jxor g17753(.dina(n18052),.dinb(w_n17437_0[0]),.dout(n18053),.clk(gclk));
	jnot g17754(.din(n18053),.dout(n18054),.clk(gclk));
	jor g17755(.dina(w_n18049_0[0]),.dinb(w_asqrt37_9[0]),.dout(n18055),.clk(gclk));
	jand g17756(.dina(w_n18055_0[1]),.dinb(w_n18054_0[1]),.dout(n18056),.clk(gclk));
	jor g17757(.dina(w_n18056_0[2]),.dinb(w_n18050_0[2]),.dout(n18057),.clk(gclk));
	jand g17758(.dina(n18057),.dinb(w_asqrt38_12[0]),.dout(n18058),.clk(gclk));
	jnot g17759(.din(w_n17442_0[0]),.dout(n18059),.clk(gclk));
	jand g17760(.dina(n18059),.dinb(w_n17440_0[0]),.dout(n18060),.clk(gclk));
	jand g17761(.dina(n18060),.dinb(w_asqrt6_20[1]),.dout(n18061),.clk(gclk));
	jxor g17762(.dina(n18061),.dinb(w_n17450_0[0]),.dout(n18062),.clk(gclk));
	jnot g17763(.din(n18062),.dout(n18063),.clk(gclk));
	jor g17764(.dina(w_n18050_0[1]),.dinb(w_asqrt38_11[2]),.dout(n18064),.clk(gclk));
	jor g17765(.dina(n18064),.dinb(w_n18056_0[1]),.dout(n18065),.clk(gclk));
	jand g17766(.dina(w_n18065_0[1]),.dinb(w_n18063_0[1]),.dout(n18066),.clk(gclk));
	jor g17767(.dina(w_n18066_0[1]),.dinb(w_n18058_0[1]),.dout(n18067),.clk(gclk));
	jand g17768(.dina(w_n18067_0[2]),.dinb(w_asqrt39_9[1]),.dout(n18068),.clk(gclk));
	jor g17769(.dina(w_n18067_0[1]),.dinb(w_asqrt39_9[0]),.dout(n18069),.clk(gclk));
	jnot g17770(.din(w_n17456_0[0]),.dout(n18070),.clk(gclk));
	jnot g17771(.din(w_n17457_0[0]),.dout(n18071),.clk(gclk));
	jand g17772(.dina(w_asqrt6_20[0]),.dinb(w_n17453_0[0]),.dout(n18072),.clk(gclk));
	jand g17773(.dina(w_n18072_0[1]),.dinb(n18071),.dout(n18073),.clk(gclk));
	jor g17774(.dina(n18073),.dinb(n18070),.dout(n18074),.clk(gclk));
	jnot g17775(.din(w_n17458_0[0]),.dout(n18075),.clk(gclk));
	jand g17776(.dina(w_n18072_0[0]),.dinb(n18075),.dout(n18076),.clk(gclk));
	jnot g17777(.din(n18076),.dout(n18077),.clk(gclk));
	jand g17778(.dina(n18077),.dinb(n18074),.dout(n18078),.clk(gclk));
	jand g17779(.dina(w_n18078_0[1]),.dinb(n18069),.dout(n18079),.clk(gclk));
	jor g17780(.dina(w_n18079_0[1]),.dinb(w_n18068_0[1]),.dout(n18080),.clk(gclk));
	jand g17781(.dina(n18080),.dinb(w_asqrt40_12[0]),.dout(n18081),.clk(gclk));
	jor g17782(.dina(w_n18068_0[0]),.dinb(w_asqrt40_11[2]),.dout(n18082),.clk(gclk));
	jor g17783(.dina(n18082),.dinb(w_n18079_0[0]),.dout(n18083),.clk(gclk));
	jnot g17784(.din(w_n17464_0[0]),.dout(n18084),.clk(gclk));
	jnot g17785(.din(w_n17466_0[0]),.dout(n18085),.clk(gclk));
	jand g17786(.dina(w_asqrt6_19[2]),.dinb(w_n17460_0[0]),.dout(n18086),.clk(gclk));
	jand g17787(.dina(w_n18086_0[1]),.dinb(n18085),.dout(n18087),.clk(gclk));
	jor g17788(.dina(n18087),.dinb(n18084),.dout(n18088),.clk(gclk));
	jnot g17789(.din(w_n17467_0[0]),.dout(n18089),.clk(gclk));
	jand g17790(.dina(w_n18086_0[0]),.dinb(n18089),.dout(n18090),.clk(gclk));
	jnot g17791(.din(n18090),.dout(n18091),.clk(gclk));
	jand g17792(.dina(n18091),.dinb(n18088),.dout(n18092),.clk(gclk));
	jand g17793(.dina(w_n18092_0[1]),.dinb(w_n18083_0[1]),.dout(n18093),.clk(gclk));
	jor g17794(.dina(n18093),.dinb(w_n18081_0[1]),.dout(n18094),.clk(gclk));
	jand g17795(.dina(w_n18094_0[1]),.dinb(w_asqrt41_9[2]),.dout(n18095),.clk(gclk));
	jxor g17796(.dina(w_n17468_0[0]),.dinb(w_n3371_10[2]),.dout(n18096),.clk(gclk));
	jand g17797(.dina(n18096),.dinb(w_asqrt6_19[1]),.dout(n18097),.clk(gclk));
	jxor g17798(.dina(n18097),.dinb(w_n17478_0[0]),.dout(n18098),.clk(gclk));
	jnot g17799(.din(n18098),.dout(n18099),.clk(gclk));
	jor g17800(.dina(w_n18094_0[0]),.dinb(w_asqrt41_9[1]),.dout(n18100),.clk(gclk));
	jand g17801(.dina(w_n18100_0[1]),.dinb(w_n18099_0[1]),.dout(n18101),.clk(gclk));
	jor g17802(.dina(w_n18101_0[2]),.dinb(w_n18095_0[2]),.dout(n18102),.clk(gclk));
	jand g17803(.dina(n18102),.dinb(w_asqrt42_12[0]),.dout(n18103),.clk(gclk));
	jnot g17804(.din(w_n17483_0[0]),.dout(n18104),.clk(gclk));
	jand g17805(.dina(n18104),.dinb(w_n17481_0[0]),.dout(n18105),.clk(gclk));
	jand g17806(.dina(n18105),.dinb(w_asqrt6_19[0]),.dout(n18106),.clk(gclk));
	jxor g17807(.dina(n18106),.dinb(w_n17491_0[0]),.dout(n18107),.clk(gclk));
	jnot g17808(.din(n18107),.dout(n18108),.clk(gclk));
	jor g17809(.dina(w_n18095_0[1]),.dinb(w_asqrt42_11[2]),.dout(n18109),.clk(gclk));
	jor g17810(.dina(n18109),.dinb(w_n18101_0[1]),.dout(n18110),.clk(gclk));
	jand g17811(.dina(w_n18110_0[1]),.dinb(w_n18108_0[1]),.dout(n18111),.clk(gclk));
	jor g17812(.dina(w_n18111_0[1]),.dinb(w_n18103_0[1]),.dout(n18112),.clk(gclk));
	jand g17813(.dina(w_n18112_0[2]),.dinb(w_asqrt43_9[2]),.dout(n18113),.clk(gclk));
	jor g17814(.dina(w_n18112_0[1]),.dinb(w_asqrt43_9[1]),.dout(n18114),.clk(gclk));
	jnot g17815(.din(w_n17497_0[0]),.dout(n18115),.clk(gclk));
	jnot g17816(.din(w_n17498_0[0]),.dout(n18116),.clk(gclk));
	jand g17817(.dina(w_asqrt6_18[2]),.dinb(w_n17494_0[0]),.dout(n18117),.clk(gclk));
	jand g17818(.dina(w_n18117_0[1]),.dinb(n18116),.dout(n18118),.clk(gclk));
	jor g17819(.dina(n18118),.dinb(n18115),.dout(n18119),.clk(gclk));
	jnot g17820(.din(w_n17499_0[0]),.dout(n18120),.clk(gclk));
	jand g17821(.dina(w_n18117_0[0]),.dinb(n18120),.dout(n18121),.clk(gclk));
	jnot g17822(.din(n18121),.dout(n18122),.clk(gclk));
	jand g17823(.dina(n18122),.dinb(n18119),.dout(n18123),.clk(gclk));
	jand g17824(.dina(w_n18123_0[1]),.dinb(n18114),.dout(n18124),.clk(gclk));
	jor g17825(.dina(w_n18124_0[1]),.dinb(w_n18113_0[1]),.dout(n18125),.clk(gclk));
	jand g17826(.dina(n18125),.dinb(w_asqrt44_12[0]),.dout(n18126),.clk(gclk));
	jor g17827(.dina(w_n18113_0[0]),.dinb(w_asqrt44_11[2]),.dout(n18127),.clk(gclk));
	jor g17828(.dina(n18127),.dinb(w_n18124_0[0]),.dout(n18128),.clk(gclk));
	jnot g17829(.din(w_n17505_0[0]),.dout(n18129),.clk(gclk));
	jnot g17830(.din(w_n17507_0[0]),.dout(n18130),.clk(gclk));
	jand g17831(.dina(w_asqrt6_18[1]),.dinb(w_n17501_0[0]),.dout(n18131),.clk(gclk));
	jand g17832(.dina(w_n18131_0[1]),.dinb(n18130),.dout(n18132),.clk(gclk));
	jor g17833(.dina(n18132),.dinb(n18129),.dout(n18133),.clk(gclk));
	jnot g17834(.din(w_n17508_0[0]),.dout(n18134),.clk(gclk));
	jand g17835(.dina(w_n18131_0[0]),.dinb(n18134),.dout(n18135),.clk(gclk));
	jnot g17836(.din(n18135),.dout(n18136),.clk(gclk));
	jand g17837(.dina(n18136),.dinb(n18133),.dout(n18137),.clk(gclk));
	jand g17838(.dina(w_n18137_0[1]),.dinb(w_n18128_0[1]),.dout(n18138),.clk(gclk));
	jor g17839(.dina(n18138),.dinb(w_n18126_0[1]),.dout(n18139),.clk(gclk));
	jand g17840(.dina(w_n18139_0[1]),.dinb(w_asqrt45_10[0]),.dout(n18140),.clk(gclk));
	jxor g17841(.dina(w_n17509_0[0]),.dinb(w_n2420_11[2]),.dout(n18141),.clk(gclk));
	jand g17842(.dina(n18141),.dinb(w_asqrt6_18[0]),.dout(n18142),.clk(gclk));
	jxor g17843(.dina(n18142),.dinb(w_n17519_0[0]),.dout(n18143),.clk(gclk));
	jnot g17844(.din(n18143),.dout(n18144),.clk(gclk));
	jor g17845(.dina(w_n18139_0[0]),.dinb(w_asqrt45_9[2]),.dout(n18145),.clk(gclk));
	jand g17846(.dina(w_n18145_0[1]),.dinb(w_n18144_0[1]),.dout(n18146),.clk(gclk));
	jor g17847(.dina(w_n18146_0[2]),.dinb(w_n18140_0[2]),.dout(n18147),.clk(gclk));
	jand g17848(.dina(n18147),.dinb(w_asqrt46_12[0]),.dout(n18148),.clk(gclk));
	jnot g17849(.din(w_n17524_0[0]),.dout(n18149),.clk(gclk));
	jand g17850(.dina(n18149),.dinb(w_n17522_0[0]),.dout(n18150),.clk(gclk));
	jand g17851(.dina(n18150),.dinb(w_asqrt6_17[2]),.dout(n18151),.clk(gclk));
	jxor g17852(.dina(n18151),.dinb(w_n17532_0[0]),.dout(n18152),.clk(gclk));
	jnot g17853(.din(n18152),.dout(n18153),.clk(gclk));
	jor g17854(.dina(w_n18140_0[1]),.dinb(w_asqrt46_11[2]),.dout(n18154),.clk(gclk));
	jor g17855(.dina(n18154),.dinb(w_n18146_0[1]),.dout(n18155),.clk(gclk));
	jand g17856(.dina(w_n18155_0[1]),.dinb(w_n18153_0[1]),.dout(n18156),.clk(gclk));
	jor g17857(.dina(w_n18156_0[1]),.dinb(w_n18148_0[1]),.dout(n18157),.clk(gclk));
	jand g17858(.dina(w_n18157_0[2]),.dinb(w_asqrt47_10[0]),.dout(n18158),.clk(gclk));
	jor g17859(.dina(w_n18157_0[1]),.dinb(w_asqrt47_9[2]),.dout(n18159),.clk(gclk));
	jnot g17860(.din(w_n17538_0[0]),.dout(n18160),.clk(gclk));
	jnot g17861(.din(w_n17539_0[0]),.dout(n18161),.clk(gclk));
	jand g17862(.dina(w_asqrt6_17[1]),.dinb(w_n17535_0[0]),.dout(n18162),.clk(gclk));
	jand g17863(.dina(w_n18162_0[1]),.dinb(n18161),.dout(n18163),.clk(gclk));
	jor g17864(.dina(n18163),.dinb(n18160),.dout(n18164),.clk(gclk));
	jnot g17865(.din(w_n17540_0[0]),.dout(n18165),.clk(gclk));
	jand g17866(.dina(w_n18162_0[0]),.dinb(n18165),.dout(n18166),.clk(gclk));
	jnot g17867(.din(n18166),.dout(n18167),.clk(gclk));
	jand g17868(.dina(n18167),.dinb(n18164),.dout(n18168),.clk(gclk));
	jand g17869(.dina(w_n18168_0[1]),.dinb(n18159),.dout(n18169),.clk(gclk));
	jor g17870(.dina(w_n18169_0[1]),.dinb(w_n18158_0[1]),.dout(n18170),.clk(gclk));
	jand g17871(.dina(n18170),.dinb(w_asqrt48_12[0]),.dout(n18171),.clk(gclk));
	jor g17872(.dina(w_n18158_0[0]),.dinb(w_asqrt48_11[2]),.dout(n18172),.clk(gclk));
	jor g17873(.dina(n18172),.dinb(w_n18169_0[0]),.dout(n18173),.clk(gclk));
	jnot g17874(.din(w_n17546_0[0]),.dout(n18174),.clk(gclk));
	jnot g17875(.din(w_n17548_0[0]),.dout(n18175),.clk(gclk));
	jand g17876(.dina(w_asqrt6_17[0]),.dinb(w_n17542_0[0]),.dout(n18176),.clk(gclk));
	jand g17877(.dina(w_n18176_0[1]),.dinb(n18175),.dout(n18177),.clk(gclk));
	jor g17878(.dina(n18177),.dinb(n18174),.dout(n18178),.clk(gclk));
	jnot g17879(.din(w_n17549_0[0]),.dout(n18179),.clk(gclk));
	jand g17880(.dina(w_n18176_0[0]),.dinb(n18179),.dout(n18180),.clk(gclk));
	jnot g17881(.din(n18180),.dout(n18181),.clk(gclk));
	jand g17882(.dina(n18181),.dinb(n18178),.dout(n18182),.clk(gclk));
	jand g17883(.dina(w_n18182_0[1]),.dinb(w_n18173_0[1]),.dout(n18183),.clk(gclk));
	jor g17884(.dina(n18183),.dinb(w_n18171_0[1]),.dout(n18184),.clk(gclk));
	jand g17885(.dina(w_n18184_0[1]),.dinb(w_asqrt49_10[1]),.dout(n18185),.clk(gclk));
	jxor g17886(.dina(w_n17550_0[0]),.dinb(w_n1641_12[1]),.dout(n18186),.clk(gclk));
	jand g17887(.dina(n18186),.dinb(w_asqrt6_16[2]),.dout(n18187),.clk(gclk));
	jxor g17888(.dina(n18187),.dinb(w_n17560_0[0]),.dout(n18188),.clk(gclk));
	jnot g17889(.din(n18188),.dout(n18189),.clk(gclk));
	jor g17890(.dina(w_n18184_0[0]),.dinb(w_asqrt49_10[0]),.dout(n18190),.clk(gclk));
	jand g17891(.dina(w_n18190_0[1]),.dinb(w_n18189_0[1]),.dout(n18191),.clk(gclk));
	jor g17892(.dina(w_n18191_0[2]),.dinb(w_n18185_0[2]),.dout(n18192),.clk(gclk));
	jand g17893(.dina(n18192),.dinb(w_asqrt50_12[0]),.dout(n18193),.clk(gclk));
	jnot g17894(.din(w_n17565_0[0]),.dout(n18194),.clk(gclk));
	jand g17895(.dina(n18194),.dinb(w_n17563_0[0]),.dout(n18195),.clk(gclk));
	jand g17896(.dina(n18195),.dinb(w_asqrt6_16[1]),.dout(n18196),.clk(gclk));
	jxor g17897(.dina(n18196),.dinb(w_n17573_0[0]),.dout(n18197),.clk(gclk));
	jnot g17898(.din(n18197),.dout(n18198),.clk(gclk));
	jor g17899(.dina(w_n18185_0[1]),.dinb(w_asqrt50_11[2]),.dout(n18199),.clk(gclk));
	jor g17900(.dina(n18199),.dinb(w_n18191_0[1]),.dout(n18200),.clk(gclk));
	jand g17901(.dina(w_n18200_0[1]),.dinb(w_n18198_0[1]),.dout(n18201),.clk(gclk));
	jor g17902(.dina(w_n18201_0[1]),.dinb(w_n18193_0[1]),.dout(n18202),.clk(gclk));
	jand g17903(.dina(w_n18202_0[2]),.dinb(w_asqrt51_10[1]),.dout(n18203),.clk(gclk));
	jor g17904(.dina(w_n18202_0[1]),.dinb(w_asqrt51_10[0]),.dout(n18204),.clk(gclk));
	jnot g17905(.din(w_n17579_0[0]),.dout(n18205),.clk(gclk));
	jnot g17906(.din(w_n17580_0[0]),.dout(n18206),.clk(gclk));
	jand g17907(.dina(w_asqrt6_16[0]),.dinb(w_n17576_0[0]),.dout(n18207),.clk(gclk));
	jand g17908(.dina(w_n18207_0[1]),.dinb(n18206),.dout(n18208),.clk(gclk));
	jor g17909(.dina(n18208),.dinb(n18205),.dout(n18209),.clk(gclk));
	jnot g17910(.din(w_n17581_0[0]),.dout(n18210),.clk(gclk));
	jand g17911(.dina(w_n18207_0[0]),.dinb(n18210),.dout(n18211),.clk(gclk));
	jnot g17912(.din(n18211),.dout(n18212),.clk(gclk));
	jand g17913(.dina(n18212),.dinb(n18209),.dout(n18213),.clk(gclk));
	jand g17914(.dina(w_n18213_0[1]),.dinb(n18204),.dout(n18214),.clk(gclk));
	jor g17915(.dina(w_n18214_0[1]),.dinb(w_n18203_0[1]),.dout(n18215),.clk(gclk));
	jand g17916(.dina(n18215),.dinb(w_asqrt52_12[0]),.dout(n18216),.clk(gclk));
	jor g17917(.dina(w_n18203_0[0]),.dinb(w_asqrt52_11[2]),.dout(n18217),.clk(gclk));
	jor g17918(.dina(n18217),.dinb(w_n18214_0[0]),.dout(n18218),.clk(gclk));
	jnot g17919(.din(w_n17587_0[0]),.dout(n18219),.clk(gclk));
	jnot g17920(.din(w_n17589_0[0]),.dout(n18220),.clk(gclk));
	jand g17921(.dina(w_asqrt6_15[2]),.dinb(w_n17583_0[0]),.dout(n18221),.clk(gclk));
	jand g17922(.dina(w_n18221_0[1]),.dinb(n18220),.dout(n18222),.clk(gclk));
	jor g17923(.dina(n18222),.dinb(n18219),.dout(n18223),.clk(gclk));
	jnot g17924(.din(w_n17590_0[0]),.dout(n18224),.clk(gclk));
	jand g17925(.dina(w_n18221_0[0]),.dinb(n18224),.dout(n18225),.clk(gclk));
	jnot g17926(.din(n18225),.dout(n18226),.clk(gclk));
	jand g17927(.dina(n18226),.dinb(n18223),.dout(n18227),.clk(gclk));
	jand g17928(.dina(w_n18227_0[1]),.dinb(w_n18218_0[1]),.dout(n18228),.clk(gclk));
	jor g17929(.dina(n18228),.dinb(w_n18216_0[1]),.dout(n18229),.clk(gclk));
	jand g17930(.dina(w_n18229_0[1]),.dinb(w_asqrt53_10[2]),.dout(n18230),.clk(gclk));
	jxor g17931(.dina(w_n17591_0[0]),.dinb(w_n1034_13[1]),.dout(n18231),.clk(gclk));
	jand g17932(.dina(n18231),.dinb(w_asqrt6_15[1]),.dout(n18232),.clk(gclk));
	jxor g17933(.dina(n18232),.dinb(w_n17601_0[0]),.dout(n18233),.clk(gclk));
	jnot g17934(.din(n18233),.dout(n18234),.clk(gclk));
	jor g17935(.dina(w_n18229_0[0]),.dinb(w_asqrt53_10[1]),.dout(n18235),.clk(gclk));
	jand g17936(.dina(w_n18235_0[1]),.dinb(w_n18234_0[1]),.dout(n18236),.clk(gclk));
	jor g17937(.dina(w_n18236_0[2]),.dinb(w_n18230_0[2]),.dout(n18237),.clk(gclk));
	jand g17938(.dina(n18237),.dinb(w_asqrt54_12[0]),.dout(n18238),.clk(gclk));
	jnot g17939(.din(w_n17606_0[0]),.dout(n18239),.clk(gclk));
	jand g17940(.dina(n18239),.dinb(w_n17604_0[0]),.dout(n18240),.clk(gclk));
	jand g17941(.dina(n18240),.dinb(w_asqrt6_15[0]),.dout(n18241),.clk(gclk));
	jxor g17942(.dina(n18241),.dinb(w_n17614_0[0]),.dout(n18242),.clk(gclk));
	jnot g17943(.din(n18242),.dout(n18243),.clk(gclk));
	jor g17944(.dina(w_n18230_0[1]),.dinb(w_asqrt54_11[2]),.dout(n18244),.clk(gclk));
	jor g17945(.dina(n18244),.dinb(w_n18236_0[1]),.dout(n18245),.clk(gclk));
	jand g17946(.dina(w_n18245_0[1]),.dinb(w_n18243_0[1]),.dout(n18246),.clk(gclk));
	jor g17947(.dina(w_n18246_0[1]),.dinb(w_n18238_0[1]),.dout(n18247),.clk(gclk));
	jand g17948(.dina(w_n18247_0[2]),.dinb(w_asqrt55_11[0]),.dout(n18248),.clk(gclk));
	jor g17949(.dina(w_n18247_0[1]),.dinb(w_asqrt55_10[2]),.dout(n18249),.clk(gclk));
	jnot g17950(.din(w_n17620_0[0]),.dout(n18250),.clk(gclk));
	jnot g17951(.din(w_n17621_0[0]),.dout(n18251),.clk(gclk));
	jand g17952(.dina(w_asqrt6_14[2]),.dinb(w_n17617_0[0]),.dout(n18252),.clk(gclk));
	jand g17953(.dina(w_n18252_0[1]),.dinb(n18251),.dout(n18253),.clk(gclk));
	jor g17954(.dina(n18253),.dinb(n18250),.dout(n18254),.clk(gclk));
	jnot g17955(.din(w_n17622_0[0]),.dout(n18255),.clk(gclk));
	jand g17956(.dina(w_n18252_0[0]),.dinb(n18255),.dout(n18256),.clk(gclk));
	jnot g17957(.din(n18256),.dout(n18257),.clk(gclk));
	jand g17958(.dina(n18257),.dinb(n18254),.dout(n18258),.clk(gclk));
	jand g17959(.dina(w_n18258_0[1]),.dinb(n18249),.dout(n18259),.clk(gclk));
	jor g17960(.dina(w_n18259_0[1]),.dinb(w_n18248_0[1]),.dout(n18260),.clk(gclk));
	jand g17961(.dina(n18260),.dinb(w_asqrt56_12[0]),.dout(n18261),.clk(gclk));
	jnot g17962(.din(w_n17626_0[0]),.dout(n18262),.clk(gclk));
	jand g17963(.dina(n18262),.dinb(w_n17624_0[0]),.dout(n18263),.clk(gclk));
	jand g17964(.dina(n18263),.dinb(w_asqrt6_14[1]),.dout(n18264),.clk(gclk));
	jxor g17965(.dina(n18264),.dinb(w_n17634_0[0]),.dout(n18265),.clk(gclk));
	jnot g17966(.din(n18265),.dout(n18266),.clk(gclk));
	jor g17967(.dina(w_n18248_0[0]),.dinb(w_asqrt56_11[2]),.dout(n18267),.clk(gclk));
	jor g17968(.dina(n18267),.dinb(w_n18259_0[0]),.dout(n18268),.clk(gclk));
	jand g17969(.dina(w_n18268_0[1]),.dinb(w_n18266_0[1]),.dout(n18269),.clk(gclk));
	jor g17970(.dina(w_n18269_0[1]),.dinb(w_n18261_0[1]),.dout(n18270),.clk(gclk));
	jand g17971(.dina(w_n18270_0[2]),.dinb(w_asqrt57_11[1]),.dout(n18271),.clk(gclk));
	jnot g17972(.din(w_n17720_0[1]),.dout(n18272),.clk(gclk));
	jor g17973(.dina(w_n18270_0[1]),.dinb(w_asqrt57_11[0]),.dout(n18273),.clk(gclk));
	jand g17974(.dina(n18273),.dinb(n18272),.dout(n18274),.clk(gclk));
	jor g17975(.dina(w_n18274_0[1]),.dinb(w_n18271_0[1]),.dout(n18275),.clk(gclk));
	jand g17976(.dina(n18275),.dinb(w_asqrt58_12[0]),.dout(n18276),.clk(gclk));
	jor g17977(.dina(w_n18271_0[0]),.dinb(w_asqrt58_11[2]),.dout(n18277),.clk(gclk));
	jor g17978(.dina(n18277),.dinb(w_n18274_0[0]),.dout(n18278),.clk(gclk));
	jnot g17979(.din(w_n17645_0[0]),.dout(n18279),.clk(gclk));
	jnot g17980(.din(w_n17647_0[0]),.dout(n18280),.clk(gclk));
	jand g17981(.dina(w_asqrt6_14[0]),.dinb(w_n17641_0[0]),.dout(n18281),.clk(gclk));
	jand g17982(.dina(w_n18281_0[1]),.dinb(n18280),.dout(n18282),.clk(gclk));
	jor g17983(.dina(n18282),.dinb(n18279),.dout(n18283),.clk(gclk));
	jnot g17984(.din(w_n17648_0[0]),.dout(n18284),.clk(gclk));
	jand g17985(.dina(w_n18281_0[0]),.dinb(n18284),.dout(n18285),.clk(gclk));
	jnot g17986(.din(n18285),.dout(n18286),.clk(gclk));
	jand g17987(.dina(n18286),.dinb(n18283),.dout(n18287),.clk(gclk));
	jand g17988(.dina(w_n18287_0[1]),.dinb(w_n18278_0[1]),.dout(n18288),.clk(gclk));
	jor g17989(.dina(n18288),.dinb(w_n18276_0[1]),.dout(n18289),.clk(gclk));
	jand g17990(.dina(w_n18289_0[2]),.dinb(w_asqrt59_11[2]),.dout(n18290),.clk(gclk));
	jor g17991(.dina(w_n18289_0[1]),.dinb(w_asqrt59_11[1]),.dout(n18291),.clk(gclk));
	jnot g17992(.din(w_n17653_0[0]),.dout(n18292),.clk(gclk));
	jnot g17993(.din(w_n17654_0[0]),.dout(n18293),.clk(gclk));
	jand g17994(.dina(w_asqrt6_13[2]),.dinb(w_n17650_0[0]),.dout(n18294),.clk(gclk));
	jand g17995(.dina(w_n18294_0[1]),.dinb(n18293),.dout(n18295),.clk(gclk));
	jor g17996(.dina(n18295),.dinb(n18292),.dout(n18296),.clk(gclk));
	jnot g17997(.din(w_n17655_0[0]),.dout(n18297),.clk(gclk));
	jand g17998(.dina(w_n18294_0[0]),.dinb(n18297),.dout(n18298),.clk(gclk));
	jnot g17999(.din(n18298),.dout(n18299),.clk(gclk));
	jand g18000(.dina(n18299),.dinb(n18296),.dout(n18300),.clk(gclk));
	jand g18001(.dina(w_n18300_0[1]),.dinb(n18291),.dout(n18301),.clk(gclk));
	jor g18002(.dina(w_n18301_0[1]),.dinb(w_n18290_0[1]),.dout(n18302),.clk(gclk));
	jand g18003(.dina(n18302),.dinb(w_asqrt60_11[2]),.dout(n18303),.clk(gclk));
	jor g18004(.dina(w_n18290_0[0]),.dinb(w_asqrt60_11[1]),.dout(n18304),.clk(gclk));
	jor g18005(.dina(n18304),.dinb(w_n18301_0[0]),.dout(n18305),.clk(gclk));
	jnot g18006(.din(w_n17661_0[0]),.dout(n18306),.clk(gclk));
	jnot g18007(.din(w_n17663_0[0]),.dout(n18307),.clk(gclk));
	jand g18008(.dina(w_asqrt6_13[1]),.dinb(w_n17657_0[0]),.dout(n18308),.clk(gclk));
	jand g18009(.dina(w_n18308_0[1]),.dinb(n18307),.dout(n18309),.clk(gclk));
	jor g18010(.dina(n18309),.dinb(n18306),.dout(n18310),.clk(gclk));
	jnot g18011(.din(w_n17664_0[0]),.dout(n18311),.clk(gclk));
	jand g18012(.dina(w_n18308_0[0]),.dinb(n18311),.dout(n18312),.clk(gclk));
	jnot g18013(.din(n18312),.dout(n18313),.clk(gclk));
	jand g18014(.dina(n18313),.dinb(n18310),.dout(n18314),.clk(gclk));
	jand g18015(.dina(w_n18314_0[1]),.dinb(w_n18305_0[1]),.dout(n18315),.clk(gclk));
	jor g18016(.dina(n18315),.dinb(w_n18303_0[1]),.dout(n18316),.clk(gclk));
	jand g18017(.dina(w_n18316_0[1]),.dinb(w_asqrt61_12[0]),.dout(n18317),.clk(gclk));
	jxor g18018(.dina(w_n17665_0[0]),.dinb(w_n290_15[1]),.dout(n18318),.clk(gclk));
	jand g18019(.dina(n18318),.dinb(w_asqrt6_13[0]),.dout(n18319),.clk(gclk));
	jxor g18020(.dina(n18319),.dinb(w_n17675_0[0]),.dout(n18320),.clk(gclk));
	jnot g18021(.din(n18320),.dout(n18321),.clk(gclk));
	jor g18022(.dina(w_n18316_0[0]),.dinb(w_asqrt61_11[2]),.dout(n18322),.clk(gclk));
	jand g18023(.dina(w_n18322_0[1]),.dinb(w_n18321_0[1]),.dout(n18323),.clk(gclk));
	jor g18024(.dina(w_n18323_0[2]),.dinb(w_n18317_0[2]),.dout(n18324),.clk(gclk));
	jand g18025(.dina(n18324),.dinb(w_asqrt62_12[0]),.dout(n18325),.clk(gclk));
	jnot g18026(.din(w_n17680_0[0]),.dout(n18326),.clk(gclk));
	jand g18027(.dina(n18326),.dinb(w_n17678_0[0]),.dout(n18327),.clk(gclk));
	jand g18028(.dina(n18327),.dinb(w_asqrt6_12[2]),.dout(n18328),.clk(gclk));
	jxor g18029(.dina(n18328),.dinb(w_n17688_0[0]),.dout(n18329),.clk(gclk));
	jnot g18030(.din(n18329),.dout(n18330),.clk(gclk));
	jor g18031(.dina(w_n18317_0[1]),.dinb(w_asqrt62_11[2]),.dout(n18331),.clk(gclk));
	jor g18032(.dina(n18331),.dinb(w_n18323_0[1]),.dout(n18332),.clk(gclk));
	jand g18033(.dina(w_n18332_0[1]),.dinb(w_n18330_0[1]),.dout(n18333),.clk(gclk));
	jor g18034(.dina(w_n18333_0[1]),.dinb(w_n18325_0[1]),.dout(n18334),.clk(gclk));
	jxor g18035(.dina(w_n17690_0[0]),.dinb(w_n199_17[2]),.dout(n18335),.clk(gclk));
	jand g18036(.dina(n18335),.dinb(w_asqrt6_12[1]),.dout(n18336),.clk(gclk));
	jxor g18037(.dina(n18336),.dinb(w_n17695_0[0]),.dout(n18337),.clk(gclk));
	jnot g18038(.din(w_n17697_0[0]),.dout(n18338),.clk(gclk));
	jnot g18039(.din(w_n17701_0[0]),.dout(n18339),.clk(gclk));
	jand g18040(.dina(w_asqrt6_12[0]),.dinb(w_n18339_0[1]),.dout(n18340),.clk(gclk));
	jand g18041(.dina(w_n18340_0[1]),.dinb(w_n18338_0[2]),.dout(n18341),.clk(gclk));
	jor g18042(.dina(n18341),.dinb(w_n17708_0[0]),.dout(n18342),.clk(gclk));
	jor g18043(.dina(n18342),.dinb(w_n18337_0[1]),.dout(n18343),.clk(gclk));
	jnot g18044(.din(n18343),.dout(n18344),.clk(gclk));
	jand g18045(.dina(n18344),.dinb(w_n18334_1[2]),.dout(n18345),.clk(gclk));
	jor g18046(.dina(n18345),.dinb(w_asqrt63_6[2]),.dout(n18346),.clk(gclk));
	jnot g18047(.din(w_n18337_0[0]),.dout(n18347),.clk(gclk));
	jor g18048(.dina(w_n18347_0[2]),.dinb(w_n18334_1[1]),.dout(n18348),.clk(gclk));
	jor g18049(.dina(w_n18340_0[0]),.dinb(w_n18338_0[1]),.dout(n18349),.clk(gclk));
	jand g18050(.dina(w_n18339_0[0]),.dinb(w_n18338_0[0]),.dout(n18350),.clk(gclk));
	jor g18051(.dina(n18350),.dinb(w_n194_16[2]),.dout(n18351),.clk(gclk));
	jnot g18052(.din(n18351),.dout(n18352),.clk(gclk));
	jand g18053(.dina(n18352),.dinb(n18349),.dout(n18353),.clk(gclk));
	jnot g18054(.din(n18353),.dout(n18354),.clk(gclk));
	jand g18055(.dina(n18354),.dinb(w_n18348_0[1]),.dout(n18355),.clk(gclk));
	jand g18056(.dina(n18355),.dinb(n18346),.dout(n18356),.clk(gclk));
	jxor g18057(.dina(w_n18270_0[0]),.dinb(w_n430_15[0]),.dout(n18357),.clk(gclk));
	jor g18058(.dina(n18357),.dinb(w_n18356_19[1]),.dout(n18358),.clk(gclk));
	jxor g18059(.dina(n18358),.dinb(w_n17720_0[0]),.dout(n18359),.clk(gclk));
	jnot g18060(.din(w_asqrt6_11[2]),.dout(n18360),.clk(gclk));
	jor g18061(.dina(w_n18356_19[0]),.dinb(w_n17722_1[0]),.dout(n18361),.clk(gclk));
	jnot g18062(.din(w_a8_0[1]),.dout(n18362),.clk(gclk));
	jnot g18063(.din(a[9]),.dout(n18363),.clk(gclk));
	jand g18064(.dina(w_n17722_0[2]),.dinb(w_n18363_0[2]),.dout(n18364),.clk(gclk));
	jand g18065(.dina(n18364),.dinb(w_n18362_1[1]),.dout(n18365),.clk(gclk));
	jnot g18066(.din(n18365),.dout(n18366),.clk(gclk));
	jand g18067(.dina(n18366),.dinb(n18361),.dout(n18367),.clk(gclk));
	jor g18068(.dina(w_n18367_0[2]),.dinb(w_n18360_3[2]),.dout(n18368),.clk(gclk));
	jor g18069(.dina(w_n18356_18[2]),.dinb(w_a10_0[0]),.dout(n18369),.clk(gclk));
	jxor g18070(.dina(w_n18369_0[1]),.dinb(w_n17723_0[0]),.dout(n18370),.clk(gclk));
	jand g18071(.dina(w_n18367_0[1]),.dinb(w_n18360_3[1]),.dout(n18371),.clk(gclk));
	jor g18072(.dina(n18371),.dinb(w_n18370_0[1]),.dout(n18372),.clk(gclk));
	jand g18073(.dina(w_n18372_0[1]),.dinb(w_n18368_0[1]),.dout(n18373),.clk(gclk));
	jor g18074(.dina(n18373),.dinb(w_n17140_9[1]),.dout(n18374),.clk(gclk));
	jand g18075(.dina(w_n18368_0[0]),.dinb(w_n17140_9[0]),.dout(n18375),.clk(gclk));
	jand g18076(.dina(n18375),.dinb(w_n18372_0[0]),.dout(n18376),.clk(gclk));
	jor g18077(.dina(w_n18369_0[0]),.dinb(w_a11_0[0]),.dout(n18377),.clk(gclk));
	jnot g18078(.din(w_n18356_18[1]),.dout(asqrt_fa_6),.clk(gclk));
	jor g18079(.dina(w_asqrt5_15[1]),.dinb(w_n18360_3[0]),.dout(n18379),.clk(gclk));
	jand g18080(.dina(n18379),.dinb(n18377),.dout(n18380),.clk(gclk));
	jxor g18081(.dina(n18380),.dinb(w_n17145_0[1]),.dout(n18381),.clk(gclk));
	jor g18082(.dina(w_n18381_0[1]),.dinb(w_n18376_0[1]),.dout(n18382),.clk(gclk));
	jand g18083(.dina(n18382),.dinb(w_n18374_0[1]),.dout(n18383),.clk(gclk));
	jor g18084(.dina(w_n18383_0[2]),.dinb(w_n17135_4[0]),.dout(n18384),.clk(gclk));
	jand g18085(.dina(w_n18383_0[1]),.dinb(w_n17135_3[2]),.dout(n18385),.clk(gclk));
	jxor g18086(.dina(w_n17726_0[0]),.dinb(w_n17140_8[2]),.dout(n18386),.clk(gclk));
	jor g18087(.dina(n18386),.dinb(w_n18356_18[0]),.dout(n18387),.clk(gclk));
	jxor g18088(.dina(n18387),.dinb(w_n17729_0[0]),.dout(n18388),.clk(gclk));
	jor g18089(.dina(w_n18388_0[1]),.dinb(n18385),.dout(n18389),.clk(gclk));
	jand g18090(.dina(w_n18389_0[1]),.dinb(w_n18384_0[1]),.dout(n18390),.clk(gclk));
	jor g18091(.dina(n18390),.dinb(w_n15955_9[2]),.dout(n18391),.clk(gclk));
	jnot g18092(.din(w_n17735_0[0]),.dout(n18392),.clk(gclk));
	jor g18093(.dina(n18392),.dinb(w_n17733_0[0]),.dout(n18393),.clk(gclk));
	jor g18094(.dina(n18393),.dinb(w_n18356_17[2]),.dout(n18394),.clk(gclk));
	jxor g18095(.dina(n18394),.dinb(w_n17744_0[0]),.dout(n18395),.clk(gclk));
	jand g18096(.dina(w_n18384_0[0]),.dinb(w_n15955_9[1]),.dout(n18396),.clk(gclk));
	jand g18097(.dina(n18396),.dinb(w_n18389_0[0]),.dout(n18397),.clk(gclk));
	jor g18098(.dina(w_n18397_0[1]),.dinb(w_n18395_0[1]),.dout(n18398),.clk(gclk));
	jand g18099(.dina(w_n18398_0[1]),.dinb(w_n18391_0[1]),.dout(n18399),.clk(gclk));
	jor g18100(.dina(w_n18399_0[2]),.dinb(w_n15950_4[1]),.dout(n18400),.clk(gclk));
	jand g18101(.dina(w_n18399_0[1]),.dinb(w_n15950_4[0]),.dout(n18401),.clk(gclk));
	jxor g18102(.dina(w_n17746_0[0]),.dinb(w_n15955_9[0]),.dout(n18402),.clk(gclk));
	jor g18103(.dina(n18402),.dinb(w_n18356_17[1]),.dout(n18403),.clk(gclk));
	jxor g18104(.dina(n18403),.dinb(w_n17751_0[0]),.dout(n18404),.clk(gclk));
	jnot g18105(.din(w_n18404_0[1]),.dout(n18405),.clk(gclk));
	jor g18106(.dina(n18405),.dinb(n18401),.dout(n18406),.clk(gclk));
	jand g18107(.dina(w_n18406_0[1]),.dinb(w_n18400_0[1]),.dout(n18407),.clk(gclk));
	jor g18108(.dina(n18407),.dinb(w_n14821_10[0]),.dout(n18408),.clk(gclk));
	jand g18109(.dina(w_n18400_0[0]),.dinb(w_n14821_9[2]),.dout(n18409),.clk(gclk));
	jand g18110(.dina(n18409),.dinb(w_n18406_0[0]),.dout(n18410),.clk(gclk));
	jnot g18111(.din(w_n17755_0[0]),.dout(n18411),.clk(gclk));
	jand g18112(.dina(w_asqrt5_15[0]),.dinb(n18411),.dout(n18412),.clk(gclk));
	jand g18113(.dina(w_n18412_0[1]),.dinb(w_n17762_0[0]),.dout(n18413),.clk(gclk));
	jor g18114(.dina(n18413),.dinb(w_n17760_0[0]),.dout(n18414),.clk(gclk));
	jand g18115(.dina(w_n18412_0[0]),.dinb(w_n17763_0[0]),.dout(n18415),.clk(gclk));
	jnot g18116(.din(n18415),.dout(n18416),.clk(gclk));
	jand g18117(.dina(n18416),.dinb(n18414),.dout(n18417),.clk(gclk));
	jnot g18118(.din(n18417),.dout(n18418),.clk(gclk));
	jor g18119(.dina(w_n18418_0[1]),.dinb(w_n18410_0[1]),.dout(n18419),.clk(gclk));
	jand g18120(.dina(n18419),.dinb(w_n18408_0[1]),.dout(n18420),.clk(gclk));
	jor g18121(.dina(w_n18420_0[2]),.dinb(w_n14816_5[0]),.dout(n18421),.clk(gclk));
	jand g18122(.dina(w_n18420_0[1]),.dinb(w_n14816_4[2]),.dout(n18422),.clk(gclk));
	jnot g18123(.din(w_n17770_0[0]),.dout(n18423),.clk(gclk));
	jxor g18124(.dina(w_n17764_0[0]),.dinb(w_n14821_9[1]),.dout(n18424),.clk(gclk));
	jor g18125(.dina(n18424),.dinb(w_n18356_17[0]),.dout(n18425),.clk(gclk));
	jxor g18126(.dina(n18425),.dinb(n18423),.dout(n18426),.clk(gclk));
	jnot g18127(.din(w_n18426_0[1]),.dout(n18427),.clk(gclk));
	jor g18128(.dina(n18427),.dinb(n18422),.dout(n18428),.clk(gclk));
	jand g18129(.dina(w_n18428_0[1]),.dinb(w_n18421_0[1]),.dout(n18429),.clk(gclk));
	jor g18130(.dina(n18429),.dinb(w_n13723_9[2]),.dout(n18430),.clk(gclk));
	jnot g18131(.din(w_n17775_0[0]),.dout(n18431),.clk(gclk));
	jor g18132(.dina(n18431),.dinb(w_n17773_0[0]),.dout(n18432),.clk(gclk));
	jor g18133(.dina(n18432),.dinb(w_n18356_16[2]),.dout(n18433),.clk(gclk));
	jxor g18134(.dina(n18433),.dinb(w_n17784_0[0]),.dout(n18434),.clk(gclk));
	jand g18135(.dina(w_n18421_0[0]),.dinb(w_n13723_9[1]),.dout(n18435),.clk(gclk));
	jand g18136(.dina(n18435),.dinb(w_n18428_0[0]),.dout(n18436),.clk(gclk));
	jor g18137(.dina(w_n18436_0[1]),.dinb(w_n18434_0[1]),.dout(n18437),.clk(gclk));
	jand g18138(.dina(w_n18437_0[1]),.dinb(w_n18430_0[1]),.dout(n18438),.clk(gclk));
	jor g18139(.dina(w_n18438_0[2]),.dinb(w_n13718_5[0]),.dout(n18439),.clk(gclk));
	jand g18140(.dina(w_n18438_0[1]),.dinb(w_n13718_4[2]),.dout(n18440),.clk(gclk));
	jnot g18141(.din(w_n17791_0[0]),.dout(n18441),.clk(gclk));
	jxor g18142(.dina(w_n17786_0[0]),.dinb(w_n13723_9[0]),.dout(n18442),.clk(gclk));
	jor g18143(.dina(n18442),.dinb(w_n18356_16[1]),.dout(n18443),.clk(gclk));
	jxor g18144(.dina(n18443),.dinb(n18441),.dout(n18444),.clk(gclk));
	jnot g18145(.din(n18444),.dout(n18445),.clk(gclk));
	jor g18146(.dina(w_n18445_0[1]),.dinb(n18440),.dout(n18446),.clk(gclk));
	jand g18147(.dina(w_n18446_0[1]),.dinb(w_n18439_0[1]),.dout(n18447),.clk(gclk));
	jor g18148(.dina(n18447),.dinb(w_n12675_10[1]),.dout(n18448),.clk(gclk));
	jand g18149(.dina(w_n18439_0[0]),.dinb(w_n12675_10[0]),.dout(n18449),.clk(gclk));
	jand g18150(.dina(n18449),.dinb(w_n18446_0[0]),.dout(n18450),.clk(gclk));
	jnot g18151(.din(w_n17794_0[0]),.dout(n18451),.clk(gclk));
	jand g18152(.dina(w_asqrt5_14[2]),.dinb(n18451),.dout(n18452),.clk(gclk));
	jand g18153(.dina(w_n18452_0[1]),.dinb(w_n17801_0[0]),.dout(n18453),.clk(gclk));
	jor g18154(.dina(n18453),.dinb(w_n17799_0[0]),.dout(n18454),.clk(gclk));
	jand g18155(.dina(w_n18452_0[0]),.dinb(w_n17802_0[0]),.dout(n18455),.clk(gclk));
	jnot g18156(.din(n18455),.dout(n18456),.clk(gclk));
	jand g18157(.dina(n18456),.dinb(n18454),.dout(n18457),.clk(gclk));
	jnot g18158(.din(n18457),.dout(n18458),.clk(gclk));
	jor g18159(.dina(w_n18458_0[1]),.dinb(w_n18450_0[1]),.dout(n18459),.clk(gclk));
	jand g18160(.dina(n18459),.dinb(w_n18448_0[1]),.dout(n18460),.clk(gclk));
	jor g18161(.dina(w_n18460_0[1]),.dinb(w_n12670_5[1]),.dout(n18461),.clk(gclk));
	jxor g18162(.dina(w_n17803_0[0]),.dinb(w_n12675_9[2]),.dout(n18462),.clk(gclk));
	jor g18163(.dina(n18462),.dinb(w_n18356_16[0]),.dout(n18463),.clk(gclk));
	jxor g18164(.dina(n18463),.dinb(w_n17808_0[0]),.dout(n18464),.clk(gclk));
	jand g18165(.dina(w_n18460_0[0]),.dinb(w_n12670_5[0]),.dout(n18465),.clk(gclk));
	jor g18166(.dina(w_n18465_0[1]),.dinb(w_n18464_0[1]),.dout(n18466),.clk(gclk));
	jand g18167(.dina(w_n18466_0[2]),.dinb(w_n18461_0[2]),.dout(n18467),.clk(gclk));
	jor g18168(.dina(n18467),.dinb(w_n11662_10[0]),.dout(n18468),.clk(gclk));
	jnot g18169(.din(w_n17813_0[0]),.dout(n18469),.clk(gclk));
	jor g18170(.dina(n18469),.dinb(w_n17811_0[0]),.dout(n18470),.clk(gclk));
	jor g18171(.dina(n18470),.dinb(w_n18356_15[2]),.dout(n18471),.clk(gclk));
	jxor g18172(.dina(n18471),.dinb(w_n17822_0[0]),.dout(n18472),.clk(gclk));
	jand g18173(.dina(w_n18461_0[1]),.dinb(w_n11662_9[2]),.dout(n18473),.clk(gclk));
	jand g18174(.dina(n18473),.dinb(w_n18466_0[1]),.dout(n18474),.clk(gclk));
	jor g18175(.dina(w_n18474_0[1]),.dinb(w_n18472_0[1]),.dout(n18475),.clk(gclk));
	jand g18176(.dina(w_n18475_0[1]),.dinb(w_n18468_0[1]),.dout(n18476),.clk(gclk));
	jor g18177(.dina(w_n18476_0[2]),.dinb(w_n11657_5[2]),.dout(n18477),.clk(gclk));
	jand g18178(.dina(w_n18476_0[1]),.dinb(w_n11657_5[1]),.dout(n18478),.clk(gclk));
	jnot g18179(.din(w_n17825_0[0]),.dout(n18479),.clk(gclk));
	jand g18180(.dina(w_asqrt5_14[1]),.dinb(n18479),.dout(n18480),.clk(gclk));
	jand g18181(.dina(w_n18480_0[1]),.dinb(w_n17830_0[0]),.dout(n18481),.clk(gclk));
	jor g18182(.dina(n18481),.dinb(w_n17829_0[0]),.dout(n18482),.clk(gclk));
	jand g18183(.dina(w_n18480_0[0]),.dinb(w_n17831_0[0]),.dout(n18483),.clk(gclk));
	jnot g18184(.din(n18483),.dout(n18484),.clk(gclk));
	jand g18185(.dina(n18484),.dinb(n18482),.dout(n18485),.clk(gclk));
	jnot g18186(.din(n18485),.dout(n18486),.clk(gclk));
	jor g18187(.dina(w_n18486_0[1]),.dinb(n18478),.dout(n18487),.clk(gclk));
	jand g18188(.dina(w_n18487_0[1]),.dinb(w_n18477_0[1]),.dout(n18488),.clk(gclk));
	jor g18189(.dina(n18488),.dinb(w_n10701_10[2]),.dout(n18489),.clk(gclk));
	jand g18190(.dina(w_n18477_0[0]),.dinb(w_n10701_10[1]),.dout(n18490),.clk(gclk));
	jand g18191(.dina(n18490),.dinb(w_n18487_0[0]),.dout(n18491),.clk(gclk));
	jnot g18192(.din(w_n17833_0[0]),.dout(n18492),.clk(gclk));
	jand g18193(.dina(w_asqrt5_14[0]),.dinb(n18492),.dout(n18493),.clk(gclk));
	jand g18194(.dina(w_n18493_0[1]),.dinb(w_n17840_0[0]),.dout(n18494),.clk(gclk));
	jor g18195(.dina(n18494),.dinb(w_n17838_0[0]),.dout(n18495),.clk(gclk));
	jand g18196(.dina(w_n18493_0[0]),.dinb(w_n17841_0[0]),.dout(n18496),.clk(gclk));
	jnot g18197(.din(n18496),.dout(n18497),.clk(gclk));
	jand g18198(.dina(n18497),.dinb(n18495),.dout(n18498),.clk(gclk));
	jnot g18199(.din(n18498),.dout(n18499),.clk(gclk));
	jor g18200(.dina(w_n18499_0[1]),.dinb(w_n18491_0[1]),.dout(n18500),.clk(gclk));
	jand g18201(.dina(n18500),.dinb(w_n18489_0[1]),.dout(n18501),.clk(gclk));
	jor g18202(.dina(w_n18501_0[1]),.dinb(w_n10696_6[1]),.dout(n18502),.clk(gclk));
	jxor g18203(.dina(w_n17842_0[0]),.dinb(w_n10701_10[0]),.dout(n18503),.clk(gclk));
	jor g18204(.dina(n18503),.dinb(w_n18356_15[1]),.dout(n18504),.clk(gclk));
	jxor g18205(.dina(n18504),.dinb(w_n17853_0[0]),.dout(n18505),.clk(gclk));
	jand g18206(.dina(w_n18501_0[0]),.dinb(w_n10696_6[0]),.dout(n18506),.clk(gclk));
	jor g18207(.dina(w_n18506_0[1]),.dinb(w_n18505_0[1]),.dout(n18507),.clk(gclk));
	jand g18208(.dina(w_n18507_0[2]),.dinb(w_n18502_0[2]),.dout(n18508),.clk(gclk));
	jor g18209(.dina(n18508),.dinb(w_n9774_10[1]),.dout(n18509),.clk(gclk));
	jnot g18210(.din(w_n17858_0[0]),.dout(n18510),.clk(gclk));
	jor g18211(.dina(n18510),.dinb(w_n17856_0[0]),.dout(n18511),.clk(gclk));
	jor g18212(.dina(n18511),.dinb(w_n18356_15[0]),.dout(n18512),.clk(gclk));
	jxor g18213(.dina(n18512),.dinb(w_n17867_0[0]),.dout(n18513),.clk(gclk));
	jand g18214(.dina(w_n18502_0[1]),.dinb(w_n9774_10[0]),.dout(n18514),.clk(gclk));
	jand g18215(.dina(n18514),.dinb(w_n18507_0[1]),.dout(n18515),.clk(gclk));
	jor g18216(.dina(w_n18515_0[1]),.dinb(w_n18513_0[1]),.dout(n18516),.clk(gclk));
	jand g18217(.dina(w_n18516_0[1]),.dinb(w_n18509_0[1]),.dout(n18517),.clk(gclk));
	jor g18218(.dina(w_n18517_0[2]),.dinb(w_n9769_6[2]),.dout(n18518),.clk(gclk));
	jand g18219(.dina(w_n18517_0[1]),.dinb(w_n9769_6[1]),.dout(n18519),.clk(gclk));
	jnot g18220(.din(w_n17870_0[0]),.dout(n18520),.clk(gclk));
	jand g18221(.dina(w_asqrt5_13[2]),.dinb(n18520),.dout(n18521),.clk(gclk));
	jand g18222(.dina(w_n18521_0[1]),.dinb(w_n17875_0[0]),.dout(n18522),.clk(gclk));
	jor g18223(.dina(n18522),.dinb(w_n17874_0[0]),.dout(n18523),.clk(gclk));
	jand g18224(.dina(w_n18521_0[0]),.dinb(w_n17876_0[0]),.dout(n18524),.clk(gclk));
	jnot g18225(.din(n18524),.dout(n18525),.clk(gclk));
	jand g18226(.dina(n18525),.dinb(n18523),.dout(n18526),.clk(gclk));
	jnot g18227(.din(n18526),.dout(n18527),.clk(gclk));
	jor g18228(.dina(w_n18527_0[1]),.dinb(n18519),.dout(n18528),.clk(gclk));
	jand g18229(.dina(w_n18528_0[1]),.dinb(w_n18518_0[1]),.dout(n18529),.clk(gclk));
	jor g18230(.dina(n18529),.dinb(w_n8898_11[1]),.dout(n18530),.clk(gclk));
	jand g18231(.dina(w_n18518_0[0]),.dinb(w_n8898_11[0]),.dout(n18531),.clk(gclk));
	jand g18232(.dina(n18531),.dinb(w_n18528_0[0]),.dout(n18532),.clk(gclk));
	jnot g18233(.din(w_n17878_0[0]),.dout(n18533),.clk(gclk));
	jand g18234(.dina(w_asqrt5_13[1]),.dinb(n18533),.dout(n18534),.clk(gclk));
	jand g18235(.dina(w_n18534_0[1]),.dinb(w_n17885_0[0]),.dout(n18535),.clk(gclk));
	jor g18236(.dina(n18535),.dinb(w_n17883_0[0]),.dout(n18536),.clk(gclk));
	jand g18237(.dina(w_n18534_0[0]),.dinb(w_n17886_0[0]),.dout(n18537),.clk(gclk));
	jnot g18238(.din(n18537),.dout(n18538),.clk(gclk));
	jand g18239(.dina(n18538),.dinb(n18536),.dout(n18539),.clk(gclk));
	jnot g18240(.din(n18539),.dout(n18540),.clk(gclk));
	jor g18241(.dina(w_n18540_0[1]),.dinb(w_n18532_0[1]),.dout(n18541),.clk(gclk));
	jand g18242(.dina(n18541),.dinb(w_n18530_0[1]),.dout(n18542),.clk(gclk));
	jor g18243(.dina(w_n18542_0[1]),.dinb(w_n8893_7[0]),.dout(n18543),.clk(gclk));
	jxor g18244(.dina(w_n17887_0[0]),.dinb(w_n8898_10[2]),.dout(n18544),.clk(gclk));
	jor g18245(.dina(n18544),.dinb(w_n18356_14[2]),.dout(n18545),.clk(gclk));
	jxor g18246(.dina(n18545),.dinb(w_n17898_0[0]),.dout(n18546),.clk(gclk));
	jand g18247(.dina(w_n18542_0[0]),.dinb(w_n8893_6[2]),.dout(n18547),.clk(gclk));
	jor g18248(.dina(w_n18547_0[1]),.dinb(w_n18546_0[1]),.dout(n18548),.clk(gclk));
	jand g18249(.dina(w_n18548_0[2]),.dinb(w_n18543_0[2]),.dout(n18549),.clk(gclk));
	jor g18250(.dina(n18549),.dinb(w_n8058_11[0]),.dout(n18550),.clk(gclk));
	jnot g18251(.din(w_n17903_0[0]),.dout(n18551),.clk(gclk));
	jor g18252(.dina(n18551),.dinb(w_n17901_0[0]),.dout(n18552),.clk(gclk));
	jor g18253(.dina(n18552),.dinb(w_n18356_14[1]),.dout(n18553),.clk(gclk));
	jxor g18254(.dina(n18553),.dinb(w_n17912_0[0]),.dout(n18554),.clk(gclk));
	jand g18255(.dina(w_n18543_0[1]),.dinb(w_n8058_10[2]),.dout(n18555),.clk(gclk));
	jand g18256(.dina(n18555),.dinb(w_n18548_0[1]),.dout(n18556),.clk(gclk));
	jor g18257(.dina(w_n18556_0[1]),.dinb(w_n18554_0[1]),.dout(n18557),.clk(gclk));
	jand g18258(.dina(w_n18557_0[1]),.dinb(w_n18550_0[1]),.dout(n18558),.clk(gclk));
	jor g18259(.dina(w_n18558_0[2]),.dinb(w_n8053_7[1]),.dout(n18559),.clk(gclk));
	jand g18260(.dina(w_n18558_0[1]),.dinb(w_n8053_7[0]),.dout(n18560),.clk(gclk));
	jnot g18261(.din(w_n17915_0[0]),.dout(n18561),.clk(gclk));
	jand g18262(.dina(w_asqrt5_13[0]),.dinb(n18561),.dout(n18562),.clk(gclk));
	jand g18263(.dina(w_n18562_0[1]),.dinb(w_n17920_0[0]),.dout(n18563),.clk(gclk));
	jor g18264(.dina(n18563),.dinb(w_n17919_0[0]),.dout(n18564),.clk(gclk));
	jand g18265(.dina(w_n18562_0[0]),.dinb(w_n17921_0[0]),.dout(n18565),.clk(gclk));
	jnot g18266(.din(n18565),.dout(n18566),.clk(gclk));
	jand g18267(.dina(n18566),.dinb(n18564),.dout(n18567),.clk(gclk));
	jnot g18268(.din(n18567),.dout(n18568),.clk(gclk));
	jor g18269(.dina(w_n18568_0[1]),.dinb(n18560),.dout(n18569),.clk(gclk));
	jand g18270(.dina(w_n18569_0[1]),.dinb(w_n18559_0[1]),.dout(n18570),.clk(gclk));
	jor g18271(.dina(n18570),.dinb(w_n7265_11[2]),.dout(n18571),.clk(gclk));
	jand g18272(.dina(w_n18559_0[0]),.dinb(w_n7265_11[1]),.dout(n18572),.clk(gclk));
	jand g18273(.dina(n18572),.dinb(w_n18569_0[0]),.dout(n18573),.clk(gclk));
	jnot g18274(.din(w_n17923_0[0]),.dout(n18574),.clk(gclk));
	jand g18275(.dina(w_asqrt5_12[2]),.dinb(n18574),.dout(n18575),.clk(gclk));
	jand g18276(.dina(w_n18575_0[1]),.dinb(w_n17930_0[0]),.dout(n18576),.clk(gclk));
	jor g18277(.dina(n18576),.dinb(w_n17928_0[0]),.dout(n18577),.clk(gclk));
	jand g18278(.dina(w_n18575_0[0]),.dinb(w_n17931_0[0]),.dout(n18578),.clk(gclk));
	jnot g18279(.din(n18578),.dout(n18579),.clk(gclk));
	jand g18280(.dina(n18579),.dinb(n18577),.dout(n18580),.clk(gclk));
	jnot g18281(.din(n18580),.dout(n18581),.clk(gclk));
	jor g18282(.dina(w_n18581_0[1]),.dinb(w_n18573_0[1]),.dout(n18582),.clk(gclk));
	jand g18283(.dina(n18582),.dinb(w_n18571_0[1]),.dout(n18583),.clk(gclk));
	jor g18284(.dina(w_n18583_0[1]),.dinb(w_n7260_8[0]),.dout(n18584),.clk(gclk));
	jxor g18285(.dina(w_n17932_0[0]),.dinb(w_n7265_11[0]),.dout(n18585),.clk(gclk));
	jor g18286(.dina(n18585),.dinb(w_n18356_14[0]),.dout(n18586),.clk(gclk));
	jxor g18287(.dina(n18586),.dinb(w_n17943_0[0]),.dout(n18587),.clk(gclk));
	jand g18288(.dina(w_n18583_0[0]),.dinb(w_n7260_7[2]),.dout(n18588),.clk(gclk));
	jor g18289(.dina(w_n18588_0[1]),.dinb(w_n18587_0[1]),.dout(n18589),.clk(gclk));
	jand g18290(.dina(w_n18589_0[2]),.dinb(w_n18584_0[2]),.dout(n18590),.clk(gclk));
	jor g18291(.dina(n18590),.dinb(w_n6505_11[1]),.dout(n18591),.clk(gclk));
	jnot g18292(.din(w_n17948_0[0]),.dout(n18592),.clk(gclk));
	jor g18293(.dina(n18592),.dinb(w_n17946_0[0]),.dout(n18593),.clk(gclk));
	jor g18294(.dina(n18593),.dinb(w_n18356_13[2]),.dout(n18594),.clk(gclk));
	jxor g18295(.dina(n18594),.dinb(w_n17957_0[0]),.dout(n18595),.clk(gclk));
	jand g18296(.dina(w_n18584_0[1]),.dinb(w_n6505_11[0]),.dout(n18596),.clk(gclk));
	jand g18297(.dina(n18596),.dinb(w_n18589_0[1]),.dout(n18597),.clk(gclk));
	jor g18298(.dina(w_n18597_0[1]),.dinb(w_n18595_0[1]),.dout(n18598),.clk(gclk));
	jand g18299(.dina(w_n18598_0[1]),.dinb(w_n18591_0[1]),.dout(n18599),.clk(gclk));
	jor g18300(.dina(w_n18599_0[2]),.dinb(w_n6500_8[1]),.dout(n18600),.clk(gclk));
	jand g18301(.dina(w_n18599_0[1]),.dinb(w_n6500_8[0]),.dout(n18601),.clk(gclk));
	jnot g18302(.din(w_n17960_0[0]),.dout(n18602),.clk(gclk));
	jand g18303(.dina(w_asqrt5_12[1]),.dinb(n18602),.dout(n18603),.clk(gclk));
	jand g18304(.dina(w_n18603_0[1]),.dinb(w_n17965_0[0]),.dout(n18604),.clk(gclk));
	jor g18305(.dina(n18604),.dinb(w_n17964_0[0]),.dout(n18605),.clk(gclk));
	jand g18306(.dina(w_n18603_0[0]),.dinb(w_n17966_0[0]),.dout(n18606),.clk(gclk));
	jnot g18307(.din(n18606),.dout(n18607),.clk(gclk));
	jand g18308(.dina(n18607),.dinb(n18605),.dout(n18608),.clk(gclk));
	jnot g18309(.din(n18608),.dout(n18609),.clk(gclk));
	jor g18310(.dina(w_n18609_0[1]),.dinb(n18601),.dout(n18610),.clk(gclk));
	jand g18311(.dina(w_n18610_0[1]),.dinb(w_n18600_0[1]),.dout(n18611),.clk(gclk));
	jor g18312(.dina(n18611),.dinb(w_n5793_12[0]),.dout(n18612),.clk(gclk));
	jand g18313(.dina(w_n18600_0[0]),.dinb(w_n5793_11[2]),.dout(n18613),.clk(gclk));
	jand g18314(.dina(n18613),.dinb(w_n18610_0[0]),.dout(n18614),.clk(gclk));
	jnot g18315(.din(w_n17968_0[0]),.dout(n18615),.clk(gclk));
	jand g18316(.dina(w_asqrt5_12[0]),.dinb(n18615),.dout(n18616),.clk(gclk));
	jand g18317(.dina(w_n18616_0[1]),.dinb(w_n17975_0[0]),.dout(n18617),.clk(gclk));
	jor g18318(.dina(n18617),.dinb(w_n17973_0[0]),.dout(n18618),.clk(gclk));
	jand g18319(.dina(w_n18616_0[0]),.dinb(w_n17976_0[0]),.dout(n18619),.clk(gclk));
	jnot g18320(.din(n18619),.dout(n18620),.clk(gclk));
	jand g18321(.dina(n18620),.dinb(n18618),.dout(n18621),.clk(gclk));
	jnot g18322(.din(n18621),.dout(n18622),.clk(gclk));
	jor g18323(.dina(w_n18622_0[1]),.dinb(w_n18614_0[1]),.dout(n18623),.clk(gclk));
	jand g18324(.dina(n18623),.dinb(w_n18612_0[1]),.dout(n18624),.clk(gclk));
	jor g18325(.dina(w_n18624_0[1]),.dinb(w_n5788_8[2]),.dout(n18625),.clk(gclk));
	jxor g18326(.dina(w_n17977_0[0]),.dinb(w_n5793_11[1]),.dout(n18626),.clk(gclk));
	jor g18327(.dina(n18626),.dinb(w_n18356_13[1]),.dout(n18627),.clk(gclk));
	jxor g18328(.dina(n18627),.dinb(w_n17988_0[0]),.dout(n18628),.clk(gclk));
	jand g18329(.dina(w_n18624_0[0]),.dinb(w_n5788_8[1]),.dout(n18629),.clk(gclk));
	jor g18330(.dina(w_n18629_0[1]),.dinb(w_n18628_0[1]),.dout(n18630),.clk(gclk));
	jand g18331(.dina(w_n18630_0[2]),.dinb(w_n18625_0[2]),.dout(n18631),.clk(gclk));
	jor g18332(.dina(n18631),.dinb(w_n5121_11[2]),.dout(n18632),.clk(gclk));
	jnot g18333(.din(w_n17993_0[0]),.dout(n18633),.clk(gclk));
	jor g18334(.dina(n18633),.dinb(w_n17991_0[0]),.dout(n18634),.clk(gclk));
	jor g18335(.dina(n18634),.dinb(w_n18356_13[0]),.dout(n18635),.clk(gclk));
	jxor g18336(.dina(n18635),.dinb(w_n18002_0[0]),.dout(n18636),.clk(gclk));
	jand g18337(.dina(w_n18625_0[1]),.dinb(w_n5121_11[1]),.dout(n18637),.clk(gclk));
	jand g18338(.dina(n18637),.dinb(w_n18630_0[1]),.dout(n18638),.clk(gclk));
	jor g18339(.dina(w_n18638_0[1]),.dinb(w_n18636_0[1]),.dout(n18639),.clk(gclk));
	jand g18340(.dina(w_n18639_0[1]),.dinb(w_n18632_0[1]),.dout(n18640),.clk(gclk));
	jor g18341(.dina(w_n18640_0[2]),.dinb(w_n5116_9[0]),.dout(n18641),.clk(gclk));
	jand g18342(.dina(w_n18640_0[1]),.dinb(w_n5116_8[2]),.dout(n18642),.clk(gclk));
	jnot g18343(.din(w_n18005_0[0]),.dout(n18643),.clk(gclk));
	jand g18344(.dina(w_asqrt5_11[2]),.dinb(n18643),.dout(n18644),.clk(gclk));
	jand g18345(.dina(w_n18644_0[1]),.dinb(w_n18010_0[0]),.dout(n18645),.clk(gclk));
	jor g18346(.dina(n18645),.dinb(w_n18009_0[0]),.dout(n18646),.clk(gclk));
	jand g18347(.dina(w_n18644_0[0]),.dinb(w_n18011_0[0]),.dout(n18647),.clk(gclk));
	jnot g18348(.din(n18647),.dout(n18648),.clk(gclk));
	jand g18349(.dina(n18648),.dinb(n18646),.dout(n18649),.clk(gclk));
	jnot g18350(.din(n18649),.dout(n18650),.clk(gclk));
	jor g18351(.dina(w_n18650_0[1]),.dinb(n18642),.dout(n18651),.clk(gclk));
	jand g18352(.dina(w_n18651_0[1]),.dinb(w_n18641_0[1]),.dout(n18652),.clk(gclk));
	jor g18353(.dina(n18652),.dinb(w_n4499_12[2]),.dout(n18653),.clk(gclk));
	jand g18354(.dina(w_n18641_0[0]),.dinb(w_n4499_12[1]),.dout(n18654),.clk(gclk));
	jand g18355(.dina(n18654),.dinb(w_n18651_0[0]),.dout(n18655),.clk(gclk));
	jnot g18356(.din(w_n18013_0[0]),.dout(n18656),.clk(gclk));
	jand g18357(.dina(w_asqrt5_11[1]),.dinb(n18656),.dout(n18657),.clk(gclk));
	jand g18358(.dina(w_n18657_0[1]),.dinb(w_n18020_0[0]),.dout(n18658),.clk(gclk));
	jor g18359(.dina(n18658),.dinb(w_n18018_0[0]),.dout(n18659),.clk(gclk));
	jand g18360(.dina(w_n18657_0[0]),.dinb(w_n18021_0[0]),.dout(n18660),.clk(gclk));
	jnot g18361(.din(n18660),.dout(n18661),.clk(gclk));
	jand g18362(.dina(n18661),.dinb(n18659),.dout(n18662),.clk(gclk));
	jnot g18363(.din(n18662),.dout(n18663),.clk(gclk));
	jor g18364(.dina(w_n18663_0[1]),.dinb(w_n18655_0[1]),.dout(n18664),.clk(gclk));
	jand g18365(.dina(n18664),.dinb(w_n18653_0[1]),.dout(n18665),.clk(gclk));
	jor g18366(.dina(w_n18665_0[1]),.dinb(w_n4494_9[2]),.dout(n18666),.clk(gclk));
	jxor g18367(.dina(w_n18022_0[0]),.dinb(w_n4499_12[0]),.dout(n18667),.clk(gclk));
	jor g18368(.dina(n18667),.dinb(w_n18356_12[2]),.dout(n18668),.clk(gclk));
	jxor g18369(.dina(n18668),.dinb(w_n18033_0[0]),.dout(n18669),.clk(gclk));
	jand g18370(.dina(w_n18665_0[0]),.dinb(w_n4494_9[1]),.dout(n18670),.clk(gclk));
	jor g18371(.dina(w_n18670_0[1]),.dinb(w_n18669_0[1]),.dout(n18671),.clk(gclk));
	jand g18372(.dina(w_n18671_0[2]),.dinb(w_n18666_0[2]),.dout(n18672),.clk(gclk));
	jor g18373(.dina(n18672),.dinb(w_n3912_12[1]),.dout(n18673),.clk(gclk));
	jnot g18374(.din(w_n18038_0[0]),.dout(n18674),.clk(gclk));
	jor g18375(.dina(n18674),.dinb(w_n18036_0[0]),.dout(n18675),.clk(gclk));
	jor g18376(.dina(n18675),.dinb(w_n18356_12[1]),.dout(n18676),.clk(gclk));
	jxor g18377(.dina(n18676),.dinb(w_n18047_0[0]),.dout(n18677),.clk(gclk));
	jand g18378(.dina(w_n18666_0[1]),.dinb(w_n3912_12[0]),.dout(n18678),.clk(gclk));
	jand g18379(.dina(n18678),.dinb(w_n18671_0[1]),.dout(n18679),.clk(gclk));
	jor g18380(.dina(w_n18679_0[1]),.dinb(w_n18677_0[1]),.dout(n18680),.clk(gclk));
	jand g18381(.dina(w_n18680_0[1]),.dinb(w_n18673_0[1]),.dout(n18681),.clk(gclk));
	jor g18382(.dina(w_n18681_0[2]),.dinb(w_n3907_10[0]),.dout(n18682),.clk(gclk));
	jand g18383(.dina(w_n18681_0[1]),.dinb(w_n3907_9[2]),.dout(n18683),.clk(gclk));
	jnot g18384(.din(w_n18050_0[0]),.dout(n18684),.clk(gclk));
	jand g18385(.dina(w_asqrt5_11[0]),.dinb(n18684),.dout(n18685),.clk(gclk));
	jand g18386(.dina(w_n18685_0[1]),.dinb(w_n18055_0[0]),.dout(n18686),.clk(gclk));
	jor g18387(.dina(n18686),.dinb(w_n18054_0[0]),.dout(n18687),.clk(gclk));
	jand g18388(.dina(w_n18685_0[0]),.dinb(w_n18056_0[0]),.dout(n18688),.clk(gclk));
	jnot g18389(.din(n18688),.dout(n18689),.clk(gclk));
	jand g18390(.dina(n18689),.dinb(n18687),.dout(n18690),.clk(gclk));
	jnot g18391(.din(n18690),.dout(n18691),.clk(gclk));
	jor g18392(.dina(w_n18691_0[1]),.dinb(n18683),.dout(n18692),.clk(gclk));
	jand g18393(.dina(w_n18692_0[1]),.dinb(w_n18682_0[1]),.dout(n18693),.clk(gclk));
	jor g18394(.dina(n18693),.dinb(w_n3376_13[1]),.dout(n18694),.clk(gclk));
	jand g18395(.dina(w_n18682_0[0]),.dinb(w_n3376_13[0]),.dout(n18695),.clk(gclk));
	jand g18396(.dina(n18695),.dinb(w_n18692_0[0]),.dout(n18696),.clk(gclk));
	jnot g18397(.din(w_n18058_0[0]),.dout(n18697),.clk(gclk));
	jand g18398(.dina(w_asqrt5_10[2]),.dinb(n18697),.dout(n18698),.clk(gclk));
	jand g18399(.dina(w_n18698_0[1]),.dinb(w_n18065_0[0]),.dout(n18699),.clk(gclk));
	jor g18400(.dina(n18699),.dinb(w_n18063_0[0]),.dout(n18700),.clk(gclk));
	jand g18401(.dina(w_n18698_0[0]),.dinb(w_n18066_0[0]),.dout(n18701),.clk(gclk));
	jnot g18402(.din(n18701),.dout(n18702),.clk(gclk));
	jand g18403(.dina(n18702),.dinb(n18700),.dout(n18703),.clk(gclk));
	jnot g18404(.din(n18703),.dout(n18704),.clk(gclk));
	jor g18405(.dina(w_n18704_0[1]),.dinb(w_n18696_0[1]),.dout(n18705),.clk(gclk));
	jand g18406(.dina(n18705),.dinb(w_n18694_0[1]),.dout(n18706),.clk(gclk));
	jor g18407(.dina(w_n18706_0[1]),.dinb(w_n3371_10[1]),.dout(n18707),.clk(gclk));
	jxor g18408(.dina(w_n18067_0[0]),.dinb(w_n3376_12[2]),.dout(n18708),.clk(gclk));
	jor g18409(.dina(n18708),.dinb(w_n18356_12[0]),.dout(n18709),.clk(gclk));
	jxor g18410(.dina(n18709),.dinb(w_n18078_0[0]),.dout(n18710),.clk(gclk));
	jand g18411(.dina(w_n18706_0[0]),.dinb(w_n3371_10[0]),.dout(n18711),.clk(gclk));
	jor g18412(.dina(w_n18711_0[1]),.dinb(w_n18710_0[1]),.dout(n18712),.clk(gclk));
	jand g18413(.dina(w_n18712_0[2]),.dinb(w_n18707_0[2]),.dout(n18713),.clk(gclk));
	jor g18414(.dina(n18713),.dinb(w_n2875_13[0]),.dout(n18714),.clk(gclk));
	jnot g18415(.din(w_n18083_0[0]),.dout(n18715),.clk(gclk));
	jor g18416(.dina(n18715),.dinb(w_n18081_0[0]),.dout(n18716),.clk(gclk));
	jor g18417(.dina(n18716),.dinb(w_n18356_11[2]),.dout(n18717),.clk(gclk));
	jxor g18418(.dina(n18717),.dinb(w_n18092_0[0]),.dout(n18718),.clk(gclk));
	jand g18419(.dina(w_n18707_0[1]),.dinb(w_n2875_12[2]),.dout(n18719),.clk(gclk));
	jand g18420(.dina(n18719),.dinb(w_n18712_0[1]),.dout(n18720),.clk(gclk));
	jor g18421(.dina(w_n18720_0[1]),.dinb(w_n18718_0[1]),.dout(n18721),.clk(gclk));
	jand g18422(.dina(w_n18721_0[1]),.dinb(w_n18714_0[1]),.dout(n18722),.clk(gclk));
	jor g18423(.dina(w_n18722_0[2]),.dinb(w_n2870_10[2]),.dout(n18723),.clk(gclk));
	jand g18424(.dina(w_n18722_0[1]),.dinb(w_n2870_10[1]),.dout(n18724),.clk(gclk));
	jnot g18425(.din(w_n18095_0[0]),.dout(n18725),.clk(gclk));
	jand g18426(.dina(w_asqrt5_10[1]),.dinb(n18725),.dout(n18726),.clk(gclk));
	jand g18427(.dina(w_n18726_0[1]),.dinb(w_n18100_0[0]),.dout(n18727),.clk(gclk));
	jor g18428(.dina(n18727),.dinb(w_n18099_0[0]),.dout(n18728),.clk(gclk));
	jand g18429(.dina(w_n18726_0[0]),.dinb(w_n18101_0[0]),.dout(n18729),.clk(gclk));
	jnot g18430(.din(n18729),.dout(n18730),.clk(gclk));
	jand g18431(.dina(n18730),.dinb(n18728),.dout(n18731),.clk(gclk));
	jnot g18432(.din(n18731),.dout(n18732),.clk(gclk));
	jor g18433(.dina(w_n18732_0[1]),.dinb(n18724),.dout(n18733),.clk(gclk));
	jand g18434(.dina(w_n18733_0[1]),.dinb(w_n18723_0[1]),.dout(n18734),.clk(gclk));
	jor g18435(.dina(n18734),.dinb(w_n2425_13[2]),.dout(n18735),.clk(gclk));
	jand g18436(.dina(w_n18723_0[0]),.dinb(w_n2425_13[1]),.dout(n18736),.clk(gclk));
	jand g18437(.dina(n18736),.dinb(w_n18733_0[0]),.dout(n18737),.clk(gclk));
	jnot g18438(.din(w_n18103_0[0]),.dout(n18738),.clk(gclk));
	jand g18439(.dina(w_asqrt5_10[0]),.dinb(n18738),.dout(n18739),.clk(gclk));
	jand g18440(.dina(w_n18739_0[1]),.dinb(w_n18110_0[0]),.dout(n18740),.clk(gclk));
	jor g18441(.dina(n18740),.dinb(w_n18108_0[0]),.dout(n18741),.clk(gclk));
	jand g18442(.dina(w_n18739_0[0]),.dinb(w_n18111_0[0]),.dout(n18742),.clk(gclk));
	jnot g18443(.din(n18742),.dout(n18743),.clk(gclk));
	jand g18444(.dina(n18743),.dinb(n18741),.dout(n18744),.clk(gclk));
	jnot g18445(.din(n18744),.dout(n18745),.clk(gclk));
	jor g18446(.dina(w_n18745_0[1]),.dinb(w_n18737_0[1]),.dout(n18746),.clk(gclk));
	jand g18447(.dina(n18746),.dinb(w_n18735_0[1]),.dout(n18747),.clk(gclk));
	jor g18448(.dina(w_n18747_0[1]),.dinb(w_n2420_11[1]),.dout(n18748),.clk(gclk));
	jxor g18449(.dina(w_n18112_0[0]),.dinb(w_n2425_13[0]),.dout(n18749),.clk(gclk));
	jor g18450(.dina(n18749),.dinb(w_n18356_11[1]),.dout(n18750),.clk(gclk));
	jxor g18451(.dina(n18750),.dinb(w_n18123_0[0]),.dout(n18751),.clk(gclk));
	jand g18452(.dina(w_n18747_0[0]),.dinb(w_n2420_11[0]),.dout(n18752),.clk(gclk));
	jor g18453(.dina(w_n18752_0[1]),.dinb(w_n18751_0[1]),.dout(n18753),.clk(gclk));
	jand g18454(.dina(w_n18753_0[2]),.dinb(w_n18748_0[2]),.dout(n18754),.clk(gclk));
	jor g18455(.dina(n18754),.dinb(w_n2010_13[1]),.dout(n18755),.clk(gclk));
	jnot g18456(.din(w_n18128_0[0]),.dout(n18756),.clk(gclk));
	jor g18457(.dina(n18756),.dinb(w_n18126_0[0]),.dout(n18757),.clk(gclk));
	jor g18458(.dina(n18757),.dinb(w_n18356_11[0]),.dout(n18758),.clk(gclk));
	jxor g18459(.dina(n18758),.dinb(w_n18137_0[0]),.dout(n18759),.clk(gclk));
	jand g18460(.dina(w_n18748_0[1]),.dinb(w_n2010_13[0]),.dout(n18760),.clk(gclk));
	jand g18461(.dina(n18760),.dinb(w_n18753_0[1]),.dout(n18761),.clk(gclk));
	jor g18462(.dina(w_n18761_0[1]),.dinb(w_n18759_0[1]),.dout(n18762),.clk(gclk));
	jand g18463(.dina(w_n18762_0[1]),.dinb(w_n18755_0[1]),.dout(n18763),.clk(gclk));
	jor g18464(.dina(w_n18763_0[2]),.dinb(w_n2005_11[2]),.dout(n18764),.clk(gclk));
	jand g18465(.dina(w_n18763_0[1]),.dinb(w_n2005_11[1]),.dout(n18765),.clk(gclk));
	jnot g18466(.din(w_n18140_0[0]),.dout(n18766),.clk(gclk));
	jand g18467(.dina(w_asqrt5_9[2]),.dinb(n18766),.dout(n18767),.clk(gclk));
	jand g18468(.dina(w_n18767_0[1]),.dinb(w_n18145_0[0]),.dout(n18768),.clk(gclk));
	jor g18469(.dina(n18768),.dinb(w_n18144_0[0]),.dout(n18769),.clk(gclk));
	jand g18470(.dina(w_n18767_0[0]),.dinb(w_n18146_0[0]),.dout(n18770),.clk(gclk));
	jnot g18471(.din(n18770),.dout(n18771),.clk(gclk));
	jand g18472(.dina(n18771),.dinb(n18769),.dout(n18772),.clk(gclk));
	jnot g18473(.din(n18772),.dout(n18773),.clk(gclk));
	jor g18474(.dina(w_n18773_0[1]),.dinb(n18765),.dout(n18774),.clk(gclk));
	jand g18475(.dina(w_n18774_0[1]),.dinb(w_n18764_0[1]),.dout(n18775),.clk(gclk));
	jor g18476(.dina(n18775),.dinb(w_n1646_14[1]),.dout(n18776),.clk(gclk));
	jand g18477(.dina(w_n18764_0[0]),.dinb(w_n1646_14[0]),.dout(n18777),.clk(gclk));
	jand g18478(.dina(n18777),.dinb(w_n18774_0[0]),.dout(n18778),.clk(gclk));
	jnot g18479(.din(w_n18148_0[0]),.dout(n18779),.clk(gclk));
	jand g18480(.dina(w_asqrt5_9[1]),.dinb(n18779),.dout(n18780),.clk(gclk));
	jand g18481(.dina(w_n18780_0[1]),.dinb(w_n18155_0[0]),.dout(n18781),.clk(gclk));
	jor g18482(.dina(n18781),.dinb(w_n18153_0[0]),.dout(n18782),.clk(gclk));
	jand g18483(.dina(w_n18780_0[0]),.dinb(w_n18156_0[0]),.dout(n18783),.clk(gclk));
	jnot g18484(.din(n18783),.dout(n18784),.clk(gclk));
	jand g18485(.dina(n18784),.dinb(n18782),.dout(n18785),.clk(gclk));
	jnot g18486(.din(n18785),.dout(n18786),.clk(gclk));
	jor g18487(.dina(w_n18786_0[1]),.dinb(w_n18778_0[1]),.dout(n18787),.clk(gclk));
	jand g18488(.dina(n18787),.dinb(w_n18776_0[1]),.dout(n18788),.clk(gclk));
	jor g18489(.dina(w_n18788_0[1]),.dinb(w_n1641_12[0]),.dout(n18789),.clk(gclk));
	jxor g18490(.dina(w_n18157_0[0]),.dinb(w_n1646_13[2]),.dout(n18790),.clk(gclk));
	jor g18491(.dina(n18790),.dinb(w_n18356_10[2]),.dout(n18791),.clk(gclk));
	jxor g18492(.dina(n18791),.dinb(w_n18168_0[0]),.dout(n18792),.clk(gclk));
	jand g18493(.dina(w_n18788_0[0]),.dinb(w_n1641_11[2]),.dout(n18793),.clk(gclk));
	jor g18494(.dina(w_n18793_0[1]),.dinb(w_n18792_0[1]),.dout(n18794),.clk(gclk));
	jand g18495(.dina(w_n18794_0[2]),.dinb(w_n18789_0[2]),.dout(n18795),.clk(gclk));
	jor g18496(.dina(n18795),.dinb(w_n1317_14[0]),.dout(n18796),.clk(gclk));
	jnot g18497(.din(w_n18173_0[0]),.dout(n18797),.clk(gclk));
	jor g18498(.dina(n18797),.dinb(w_n18171_0[0]),.dout(n18798),.clk(gclk));
	jor g18499(.dina(n18798),.dinb(w_n18356_10[1]),.dout(n18799),.clk(gclk));
	jxor g18500(.dina(n18799),.dinb(w_n18182_0[0]),.dout(n18800),.clk(gclk));
	jand g18501(.dina(w_n18789_0[1]),.dinb(w_n1317_13[2]),.dout(n18801),.clk(gclk));
	jand g18502(.dina(n18801),.dinb(w_n18794_0[1]),.dout(n18802),.clk(gclk));
	jor g18503(.dina(w_n18802_0[1]),.dinb(w_n18800_0[1]),.dout(n18803),.clk(gclk));
	jand g18504(.dina(w_n18803_0[1]),.dinb(w_n18796_0[1]),.dout(n18804),.clk(gclk));
	jor g18505(.dina(w_n18804_0[2]),.dinb(w_n1312_12[1]),.dout(n18805),.clk(gclk));
	jand g18506(.dina(w_n18804_0[1]),.dinb(w_n1312_12[0]),.dout(n18806),.clk(gclk));
	jnot g18507(.din(w_n18185_0[0]),.dout(n18807),.clk(gclk));
	jand g18508(.dina(w_asqrt5_9[0]),.dinb(n18807),.dout(n18808),.clk(gclk));
	jand g18509(.dina(w_n18808_0[1]),.dinb(w_n18190_0[0]),.dout(n18809),.clk(gclk));
	jor g18510(.dina(n18809),.dinb(w_n18189_0[0]),.dout(n18810),.clk(gclk));
	jand g18511(.dina(w_n18808_0[0]),.dinb(w_n18191_0[0]),.dout(n18811),.clk(gclk));
	jnot g18512(.din(n18811),.dout(n18812),.clk(gclk));
	jand g18513(.dina(n18812),.dinb(n18810),.dout(n18813),.clk(gclk));
	jnot g18514(.din(n18813),.dout(n18814),.clk(gclk));
	jor g18515(.dina(w_n18814_0[1]),.dinb(n18806),.dout(n18815),.clk(gclk));
	jand g18516(.dina(w_n18815_0[1]),.dinb(w_n18805_0[1]),.dout(n18816),.clk(gclk));
	jor g18517(.dina(n18816),.dinb(w_n1039_14[2]),.dout(n18817),.clk(gclk));
	jand g18518(.dina(w_n18805_0[0]),.dinb(w_n1039_14[1]),.dout(n18818),.clk(gclk));
	jand g18519(.dina(n18818),.dinb(w_n18815_0[0]),.dout(n18819),.clk(gclk));
	jnot g18520(.din(w_n18193_0[0]),.dout(n18820),.clk(gclk));
	jand g18521(.dina(w_asqrt5_8[2]),.dinb(n18820),.dout(n18821),.clk(gclk));
	jand g18522(.dina(w_n18821_0[1]),.dinb(w_n18200_0[0]),.dout(n18822),.clk(gclk));
	jor g18523(.dina(n18822),.dinb(w_n18198_0[0]),.dout(n18823),.clk(gclk));
	jand g18524(.dina(w_n18821_0[0]),.dinb(w_n18201_0[0]),.dout(n18824),.clk(gclk));
	jnot g18525(.din(n18824),.dout(n18825),.clk(gclk));
	jand g18526(.dina(n18825),.dinb(n18823),.dout(n18826),.clk(gclk));
	jnot g18527(.din(n18826),.dout(n18827),.clk(gclk));
	jor g18528(.dina(w_n18827_0[1]),.dinb(w_n18819_0[1]),.dout(n18828),.clk(gclk));
	jand g18529(.dina(n18828),.dinb(w_n18817_0[1]),.dout(n18829),.clk(gclk));
	jor g18530(.dina(w_n18829_0[1]),.dinb(w_n1034_13[0]),.dout(n18830),.clk(gclk));
	jxor g18531(.dina(w_n18202_0[0]),.dinb(w_n1039_14[0]),.dout(n18831),.clk(gclk));
	jor g18532(.dina(n18831),.dinb(w_n18356_10[0]),.dout(n18832),.clk(gclk));
	jxor g18533(.dina(n18832),.dinb(w_n18213_0[0]),.dout(n18833),.clk(gclk));
	jand g18534(.dina(w_n18829_0[0]),.dinb(w_n1034_12[2]),.dout(n18834),.clk(gclk));
	jor g18535(.dina(w_n18834_0[1]),.dinb(w_n18833_0[1]),.dout(n18835),.clk(gclk));
	jand g18536(.dina(w_n18835_0[2]),.dinb(w_n18830_0[2]),.dout(n18836),.clk(gclk));
	jor g18537(.dina(n18836),.dinb(w_n796_14[1]),.dout(n18837),.clk(gclk));
	jnot g18538(.din(w_n18218_0[0]),.dout(n18838),.clk(gclk));
	jor g18539(.dina(n18838),.dinb(w_n18216_0[0]),.dout(n18839),.clk(gclk));
	jor g18540(.dina(n18839),.dinb(w_n18356_9[2]),.dout(n18840),.clk(gclk));
	jxor g18541(.dina(n18840),.dinb(w_n18227_0[0]),.dout(n18841),.clk(gclk));
	jand g18542(.dina(w_n18830_0[1]),.dinb(w_n796_14[0]),.dout(n18842),.clk(gclk));
	jand g18543(.dina(n18842),.dinb(w_n18835_0[1]),.dout(n18843),.clk(gclk));
	jor g18544(.dina(w_n18843_0[1]),.dinb(w_n18841_0[1]),.dout(n18844),.clk(gclk));
	jand g18545(.dina(w_n18844_0[1]),.dinb(w_n18837_0[1]),.dout(n18845),.clk(gclk));
	jor g18546(.dina(w_n18845_0[2]),.dinb(w_n791_13[1]),.dout(n18846),.clk(gclk));
	jand g18547(.dina(w_n18845_0[1]),.dinb(w_n791_13[0]),.dout(n18847),.clk(gclk));
	jnot g18548(.din(w_n18230_0[0]),.dout(n18848),.clk(gclk));
	jand g18549(.dina(w_asqrt5_8[1]),.dinb(n18848),.dout(n18849),.clk(gclk));
	jand g18550(.dina(w_n18849_0[1]),.dinb(w_n18235_0[0]),.dout(n18850),.clk(gclk));
	jor g18551(.dina(n18850),.dinb(w_n18234_0[0]),.dout(n18851),.clk(gclk));
	jand g18552(.dina(w_n18849_0[0]),.dinb(w_n18236_0[0]),.dout(n18852),.clk(gclk));
	jnot g18553(.din(n18852),.dout(n18853),.clk(gclk));
	jand g18554(.dina(n18853),.dinb(n18851),.dout(n18854),.clk(gclk));
	jnot g18555(.din(n18854),.dout(n18855),.clk(gclk));
	jor g18556(.dina(w_n18855_0[1]),.dinb(n18847),.dout(n18856),.clk(gclk));
	jand g18557(.dina(w_n18856_0[1]),.dinb(w_n18846_0[1]),.dout(n18857),.clk(gclk));
	jor g18558(.dina(n18857),.dinb(w_n595_15[0]),.dout(n18858),.clk(gclk));
	jand g18559(.dina(w_n18846_0[0]),.dinb(w_n595_14[2]),.dout(n18859),.clk(gclk));
	jand g18560(.dina(n18859),.dinb(w_n18856_0[0]),.dout(n18860),.clk(gclk));
	jnot g18561(.din(w_n18238_0[0]),.dout(n18861),.clk(gclk));
	jand g18562(.dina(w_asqrt5_8[0]),.dinb(n18861),.dout(n18862),.clk(gclk));
	jand g18563(.dina(w_n18862_0[1]),.dinb(w_n18245_0[0]),.dout(n18863),.clk(gclk));
	jor g18564(.dina(n18863),.dinb(w_n18243_0[0]),.dout(n18864),.clk(gclk));
	jand g18565(.dina(w_n18862_0[0]),.dinb(w_n18246_0[0]),.dout(n18865),.clk(gclk));
	jnot g18566(.din(n18865),.dout(n18866),.clk(gclk));
	jand g18567(.dina(n18866),.dinb(n18864),.dout(n18867),.clk(gclk));
	jnot g18568(.din(n18867),.dout(n18868),.clk(gclk));
	jor g18569(.dina(w_n18868_0[1]),.dinb(w_n18860_0[1]),.dout(n18869),.clk(gclk));
	jand g18570(.dina(n18869),.dinb(w_n18858_0[1]),.dout(n18870),.clk(gclk));
	jor g18571(.dina(w_n18870_0[1]),.dinb(w_n590_13[2]),.dout(n18871),.clk(gclk));
	jxor g18572(.dina(w_n18247_0[0]),.dinb(w_n595_14[1]),.dout(n18872),.clk(gclk));
	jor g18573(.dina(n18872),.dinb(w_n18356_9[1]),.dout(n18873),.clk(gclk));
	jxor g18574(.dina(n18873),.dinb(w_n18258_0[0]),.dout(n18874),.clk(gclk));
	jand g18575(.dina(w_n18870_0[0]),.dinb(w_n590_13[1]),.dout(n18875),.clk(gclk));
	jor g18576(.dina(w_n18875_0[1]),.dinb(w_n18874_0[1]),.dout(n18876),.clk(gclk));
	jand g18577(.dina(w_n18876_0[2]),.dinb(w_n18871_0[2]),.dout(n18877),.clk(gclk));
	jor g18578(.dina(n18877),.dinb(w_n430_14[2]),.dout(n18878),.clk(gclk));
	jand g18579(.dina(w_n18871_0[1]),.dinb(w_n430_14[1]),.dout(n18879),.clk(gclk));
	jand g18580(.dina(n18879),.dinb(w_n18876_0[1]),.dout(n18880),.clk(gclk));
	jnot g18581(.din(w_n18261_0[0]),.dout(n18881),.clk(gclk));
	jand g18582(.dina(w_asqrt5_7[2]),.dinb(n18881),.dout(n18882),.clk(gclk));
	jand g18583(.dina(w_n18882_0[1]),.dinb(w_n18268_0[0]),.dout(n18883),.clk(gclk));
	jor g18584(.dina(n18883),.dinb(w_n18266_0[0]),.dout(n18884),.clk(gclk));
	jand g18585(.dina(w_n18882_0[0]),.dinb(w_n18269_0[0]),.dout(n18885),.clk(gclk));
	jnot g18586(.din(n18885),.dout(n18886),.clk(gclk));
	jand g18587(.dina(n18886),.dinb(n18884),.dout(n18887),.clk(gclk));
	jnot g18588(.din(n18887),.dout(n18888),.clk(gclk));
	jor g18589(.dina(w_n18888_0[1]),.dinb(w_n18880_0[1]),.dout(n18889),.clk(gclk));
	jand g18590(.dina(n18889),.dinb(w_n18878_0[1]),.dout(n18890),.clk(gclk));
	jor g18591(.dina(w_n18890_0[2]),.dinb(w_n425_14[0]),.dout(n18891),.clk(gclk));
	jnot g18592(.din(w_n18359_0[1]),.dout(n18892),.clk(gclk));
	jand g18593(.dina(w_n18890_0[1]),.dinb(w_n425_13[2]),.dout(n18893),.clk(gclk));
	jor g18594(.dina(n18893),.dinb(n18892),.dout(n18894),.clk(gclk));
	jand g18595(.dina(w_n18894_0[1]),.dinb(w_n18891_0[1]),.dout(n18895),.clk(gclk));
	jor g18596(.dina(n18895),.dinb(w_n305_15[2]),.dout(n18896),.clk(gclk));
	jnot g18597(.din(w_n18278_0[0]),.dout(n18897),.clk(gclk));
	jor g18598(.dina(n18897),.dinb(w_n18276_0[0]),.dout(n18898),.clk(gclk));
	jor g18599(.dina(n18898),.dinb(w_n18356_9[0]),.dout(n18899),.clk(gclk));
	jxor g18600(.dina(n18899),.dinb(w_n18287_0[0]),.dout(n18900),.clk(gclk));
	jand g18601(.dina(w_n18891_0[0]),.dinb(w_n305_15[1]),.dout(n18901),.clk(gclk));
	jand g18602(.dina(n18901),.dinb(w_n18894_0[0]),.dout(n18902),.clk(gclk));
	jor g18603(.dina(w_n18902_0[1]),.dinb(w_n18900_0[1]),.dout(n18903),.clk(gclk));
	jand g18604(.dina(w_n18903_0[1]),.dinb(w_n18896_0[1]),.dout(n18904),.clk(gclk));
	jor g18605(.dina(w_n18904_0[1]),.dinb(w_n290_15[0]),.dout(n18905),.clk(gclk));
	jxor g18606(.dina(w_n18289_0[0]),.dinb(w_n305_15[0]),.dout(n18906),.clk(gclk));
	jor g18607(.dina(n18906),.dinb(w_n18356_8[2]),.dout(n18907),.clk(gclk));
	jxor g18608(.dina(n18907),.dinb(w_n18300_0[0]),.dout(n18908),.clk(gclk));
	jand g18609(.dina(w_n18904_0[0]),.dinb(w_n290_14[2]),.dout(n18909),.clk(gclk));
	jor g18610(.dina(w_n18909_0[1]),.dinb(w_n18908_0[1]),.dout(n18910),.clk(gclk));
	jand g18611(.dina(w_n18910_0[2]),.dinb(w_n18905_0[2]),.dout(n18911),.clk(gclk));
	jor g18612(.dina(n18911),.dinb(w_n223_15[1]),.dout(n18912),.clk(gclk));
	jnot g18613(.din(w_n18305_0[0]),.dout(n18913),.clk(gclk));
	jor g18614(.dina(n18913),.dinb(w_n18303_0[0]),.dout(n18914),.clk(gclk));
	jor g18615(.dina(n18914),.dinb(w_n18356_8[1]),.dout(n18915),.clk(gclk));
	jxor g18616(.dina(n18915),.dinb(w_n18314_0[0]),.dout(n18916),.clk(gclk));
	jand g18617(.dina(w_n18905_0[1]),.dinb(w_n223_15[0]),.dout(n18917),.clk(gclk));
	jand g18618(.dina(n18917),.dinb(w_n18910_0[1]),.dout(n18918),.clk(gclk));
	jor g18619(.dina(w_n18918_0[1]),.dinb(w_n18916_0[1]),.dout(n18919),.clk(gclk));
	jand g18620(.dina(w_n18919_0[1]),.dinb(w_n18912_0[1]),.dout(n18920),.clk(gclk));
	jor g18621(.dina(w_n18920_0[2]),.dinb(w_n199_17[1]),.dout(n18921),.clk(gclk));
	jand g18622(.dina(w_n18920_0[1]),.dinb(w_n199_17[0]),.dout(n18922),.clk(gclk));
	jnot g18623(.din(w_n18317_0[0]),.dout(n18923),.clk(gclk));
	jand g18624(.dina(w_asqrt5_7[1]),.dinb(n18923),.dout(n18924),.clk(gclk));
	jand g18625(.dina(w_n18924_0[1]),.dinb(w_n18322_0[0]),.dout(n18925),.clk(gclk));
	jor g18626(.dina(n18925),.dinb(w_n18321_0[0]),.dout(n18926),.clk(gclk));
	jand g18627(.dina(w_n18924_0[0]),.dinb(w_n18323_0[0]),.dout(n18927),.clk(gclk));
	jnot g18628(.din(n18927),.dout(n18928),.clk(gclk));
	jand g18629(.dina(n18928),.dinb(n18926),.dout(n18929),.clk(gclk));
	jnot g18630(.din(n18929),.dout(n18930),.clk(gclk));
	jor g18631(.dina(w_n18930_0[1]),.dinb(n18922),.dout(n18931),.clk(gclk));
	jand g18632(.dina(n18931),.dinb(n18921),.dout(n18932),.clk(gclk));
	jnot g18633(.din(w_n18325_0[0]),.dout(n18933),.clk(gclk));
	jand g18634(.dina(w_asqrt5_7[0]),.dinb(n18933),.dout(n18934),.clk(gclk));
	jand g18635(.dina(w_n18934_0[1]),.dinb(w_n18332_0[0]),.dout(n18935),.clk(gclk));
	jor g18636(.dina(n18935),.dinb(w_n18330_0[0]),.dout(n18936),.clk(gclk));
	jand g18637(.dina(w_n18934_0[0]),.dinb(w_n18333_0[0]),.dout(n18937),.clk(gclk));
	jnot g18638(.din(n18937),.dout(n18938),.clk(gclk));
	jand g18639(.dina(n18938),.dinb(n18936),.dout(n18939),.clk(gclk));
	jnot g18640(.din(w_n18939_0[2]),.dout(n18940),.clk(gclk));
	jnot g18641(.din(w_n18348_0[0]),.dout(n18941),.clk(gclk));
	jand g18642(.dina(w_asqrt5_6[2]),.dinb(w_n18347_0[1]),.dout(n18942),.clk(gclk));
	jand g18643(.dina(w_n18942_0[1]),.dinb(w_n18334_1[0]),.dout(n18943),.clk(gclk));
	jor g18644(.dina(n18943),.dinb(n18941),.dout(n18944),.clk(gclk));
	jor g18645(.dina(n18944),.dinb(w_n18940_0[1]),.dout(n18945),.clk(gclk));
	jor g18646(.dina(n18945),.dinb(w_n18932_0[2]),.dout(n18946),.clk(gclk));
	jand g18647(.dina(n18946),.dinb(w_n194_16[1]),.dout(n18947),.clk(gclk));
	jand g18648(.dina(w_n18940_0[0]),.dinb(w_n18932_0[1]),.dout(n18948),.clk(gclk));
	jor g18649(.dina(w_n18942_0[0]),.dinb(w_n18334_0[2]),.dout(n18949),.clk(gclk));
	jand g18650(.dina(w_n18347_0[0]),.dinb(w_n18334_0[1]),.dout(n18950),.clk(gclk));
	jor g18651(.dina(n18950),.dinb(w_n194_16[0]),.dout(n18951),.clk(gclk));
	jnot g18652(.din(n18951),.dout(n18952),.clk(gclk));
	jand g18653(.dina(n18952),.dinb(n18949),.dout(n18953),.clk(gclk));
	jor g18654(.dina(n18953),.dinb(w_n18948_0[1]),.dout(n18954),.clk(gclk));
	jor g18655(.dina(n18954),.dinb(n18947),.dout(asqrt_fa_5),.clk(gclk));
	jxor g18656(.dina(w_n18890_0[0]),.dinb(w_n425_13[1]),.dout(n18956),.clk(gclk));
	jand g18657(.dina(n18956),.dinb(w_asqrt4_31),.dout(n18957),.clk(gclk));
	jxor g18658(.dina(n18957),.dinb(w_n18359_0[0]),.dout(n18958),.clk(gclk));
	jnot g18659(.din(w_n18958_0[1]),.dout(n18959),.clk(gclk));
	jand g18660(.dina(w_asqrt4_30[2]),.dinb(w_a8_0[0]),.dout(n18960),.clk(gclk));
	jnot g18661(.din(w_a6_0[1]),.dout(n18961),.clk(gclk));
	jnot g18662(.din(w_a7_0[1]),.dout(n18962),.clk(gclk));
	jand g18663(.dina(w_n18362_1[0]),.dinb(w_n18962_0[1]),.dout(n18963),.clk(gclk));
	jand g18664(.dina(n18963),.dinb(w_n18961_1[1]),.dout(n18964),.clk(gclk));
	jor g18665(.dina(n18964),.dinb(n18960),.dout(n18965),.clk(gclk));
	jand g18666(.dina(w_n18965_0[2]),.dinb(w_asqrt5_6[1]),.dout(n18966),.clk(gclk));
	jand g18667(.dina(w_asqrt4_30[1]),.dinb(w_n18362_0[2]),.dout(n18967),.clk(gclk));
	jxor g18668(.dina(w_n18967_0[1]),.dinb(w_n18363_0[1]),.dout(n18968),.clk(gclk));
	jor g18669(.dina(w_n18965_0[1]),.dinb(w_asqrt5_6[0]),.dout(n18969),.clk(gclk));
	jand g18670(.dina(n18969),.dinb(w_n18968_0[1]),.dout(n18970),.clk(gclk));
	jor g18671(.dina(w_n18970_0[1]),.dinb(w_n18966_0[1]),.dout(n18971),.clk(gclk));
	jand g18672(.dina(n18971),.dinb(w_asqrt6_11[1]),.dout(n18972),.clk(gclk));
	jor g18673(.dina(w_n18966_0[0]),.dinb(w_asqrt6_11[0]),.dout(n18973),.clk(gclk));
	jor g18674(.dina(n18973),.dinb(w_n18970_0[0]),.dout(n18974),.clk(gclk));
	jand g18675(.dina(w_n18967_0[0]),.dinb(w_n18363_0[0]),.dout(n18975),.clk(gclk));
	jnot g18676(.din(w_asqrt4_30[0]),.dout(n18976),.clk(gclk));
	jand g18677(.dina(w_n18976_2[2]),.dinb(w_asqrt5_5[2]),.dout(n18977),.clk(gclk));
	jor g18678(.dina(n18977),.dinb(n18975),.dout(n18978),.clk(gclk));
	jxor g18679(.dina(n18978),.dinb(w_n17722_0[1]),.dout(n18979),.clk(gclk));
	jand g18680(.dina(w_n18979_0[1]),.dinb(w_n18974_0[1]),.dout(n18980),.clk(gclk));
	jor g18681(.dina(n18980),.dinb(w_n18972_0[1]),.dout(n18981),.clk(gclk));
	jand g18682(.dina(w_n18981_0[2]),.dinb(w_asqrt7_6[0]),.dout(n18982),.clk(gclk));
	jor g18683(.dina(w_n18981_0[1]),.dinb(w_asqrt7_5[2]),.dout(n18983),.clk(gclk));
	jxor g18684(.dina(w_n18367_0[0]),.dinb(w_n18360_2[2]),.dout(n18984),.clk(gclk));
	jand g18685(.dina(n18984),.dinb(w_asqrt4_29[2]),.dout(n18985),.clk(gclk));
	jxor g18686(.dina(n18985),.dinb(w_n18370_0[0]),.dout(n18986),.clk(gclk));
	jnot g18687(.din(w_n18986_0[1]),.dout(n18987),.clk(gclk));
	jand g18688(.dina(n18987),.dinb(n18983),.dout(n18988),.clk(gclk));
	jor g18689(.dina(w_n18988_0[1]),.dinb(w_n18982_0[1]),.dout(n18989),.clk(gclk));
	jand g18690(.dina(n18989),.dinb(w_asqrt8_11[1]),.dout(n18990),.clk(gclk));
	jnot g18691(.din(w_n18376_0[0]),.dout(n18991),.clk(gclk));
	jand g18692(.dina(n18991),.dinb(w_n18374_0[0]),.dout(n18992),.clk(gclk));
	jand g18693(.dina(n18992),.dinb(w_asqrt4_29[1]),.dout(n18993),.clk(gclk));
	jxor g18694(.dina(n18993),.dinb(w_n18381_0[0]),.dout(n18994),.clk(gclk));
	jnot g18695(.din(n18994),.dout(n18995),.clk(gclk));
	jor g18696(.dina(w_n18982_0[0]),.dinb(w_asqrt8_11[0]),.dout(n18996),.clk(gclk));
	jor g18697(.dina(n18996),.dinb(w_n18988_0[0]),.dout(n18997),.clk(gclk));
	jand g18698(.dina(w_n18997_0[1]),.dinb(w_n18995_0[1]),.dout(n18998),.clk(gclk));
	jor g18699(.dina(w_n18998_0[1]),.dinb(w_n18990_0[1]),.dout(n18999),.clk(gclk));
	jand g18700(.dina(w_n18999_0[2]),.dinb(w_asqrt9_6[1]),.dout(n19000),.clk(gclk));
	jor g18701(.dina(w_n18999_0[1]),.dinb(w_asqrt9_6[0]),.dout(n19001),.clk(gclk));
	jnot g18702(.din(w_n18388_0[0]),.dout(n19002),.clk(gclk));
	jxor g18703(.dina(w_n18383_0[0]),.dinb(w_n17135_3[1]),.dout(n19003),.clk(gclk));
	jand g18704(.dina(n19003),.dinb(w_asqrt4_29[0]),.dout(n19004),.clk(gclk));
	jxor g18705(.dina(n19004),.dinb(n19002),.dout(n19005),.clk(gclk));
	jand g18706(.dina(w_n19005_0[1]),.dinb(n19001),.dout(n19006),.clk(gclk));
	jor g18707(.dina(w_n19006_0[1]),.dinb(w_n19000_0[1]),.dout(n19007),.clk(gclk));
	jand g18708(.dina(n19007),.dinb(w_asqrt10_11[1]),.dout(n19008),.clk(gclk));
	jor g18709(.dina(w_n19000_0[0]),.dinb(w_asqrt10_11[0]),.dout(n19009),.clk(gclk));
	jor g18710(.dina(n19009),.dinb(w_n19006_0[0]),.dout(n19010),.clk(gclk));
	jnot g18711(.din(w_n18395_0[0]),.dout(n19011),.clk(gclk));
	jnot g18712(.din(w_n18397_0[0]),.dout(n19012),.clk(gclk));
	jand g18713(.dina(w_asqrt4_28[2]),.dinb(w_n18391_0[0]),.dout(n19013),.clk(gclk));
	jand g18714(.dina(w_n19013_0[1]),.dinb(n19012),.dout(n19014),.clk(gclk));
	jor g18715(.dina(n19014),.dinb(n19011),.dout(n19015),.clk(gclk));
	jnot g18716(.din(w_n18398_0[0]),.dout(n19016),.clk(gclk));
	jand g18717(.dina(w_n19013_0[0]),.dinb(n19016),.dout(n19017),.clk(gclk));
	jnot g18718(.din(n19017),.dout(n19018),.clk(gclk));
	jand g18719(.dina(n19018),.dinb(n19015),.dout(n19019),.clk(gclk));
	jand g18720(.dina(w_n19019_0[1]),.dinb(w_n19010_0[1]),.dout(n19020),.clk(gclk));
	jor g18721(.dina(n19020),.dinb(w_n19008_0[1]),.dout(n19021),.clk(gclk));
	jand g18722(.dina(w_n19021_0[2]),.dinb(w_asqrt11_6[1]),.dout(n19022),.clk(gclk));
	jor g18723(.dina(w_n19021_0[1]),.dinb(w_asqrt11_6[0]),.dout(n19023),.clk(gclk));
	jxor g18724(.dina(w_n18399_0[0]),.dinb(w_n15950_3[2]),.dout(n19024),.clk(gclk));
	jand g18725(.dina(n19024),.dinb(w_asqrt4_28[1]),.dout(n19025),.clk(gclk));
	jxor g18726(.dina(n19025),.dinb(w_n18404_0[0]),.dout(n19026),.clk(gclk));
	jand g18727(.dina(w_n19026_0[1]),.dinb(n19023),.dout(n19027),.clk(gclk));
	jor g18728(.dina(w_n19027_0[1]),.dinb(w_n19022_0[1]),.dout(n19028),.clk(gclk));
	jand g18729(.dina(n19028),.dinb(w_asqrt12_11[1]),.dout(n19029),.clk(gclk));
	jnot g18730(.din(w_n18410_0[0]),.dout(n19030),.clk(gclk));
	jand g18731(.dina(n19030),.dinb(w_n18408_0[0]),.dout(n19031),.clk(gclk));
	jand g18732(.dina(n19031),.dinb(w_asqrt4_28[0]),.dout(n19032),.clk(gclk));
	jxor g18733(.dina(n19032),.dinb(w_n18418_0[0]),.dout(n19033),.clk(gclk));
	jnot g18734(.din(n19033),.dout(n19034),.clk(gclk));
	jor g18735(.dina(w_n19022_0[0]),.dinb(w_asqrt12_11[0]),.dout(n19035),.clk(gclk));
	jor g18736(.dina(n19035),.dinb(w_n19027_0[0]),.dout(n19036),.clk(gclk));
	jand g18737(.dina(w_n19036_0[1]),.dinb(w_n19034_0[1]),.dout(n19037),.clk(gclk));
	jor g18738(.dina(w_n19037_0[1]),.dinb(w_n19029_0[1]),.dout(n19038),.clk(gclk));
	jand g18739(.dina(w_n19038_0[2]),.dinb(w_asqrt13_6[2]),.dout(n19039),.clk(gclk));
	jor g18740(.dina(w_n19038_0[1]),.dinb(w_asqrt13_6[1]),.dout(n19040),.clk(gclk));
	jxor g18741(.dina(w_n18420_0[0]),.dinb(w_n14816_4[1]),.dout(n19041),.clk(gclk));
	jand g18742(.dina(n19041),.dinb(w_asqrt4_27[2]),.dout(n19042),.clk(gclk));
	jxor g18743(.dina(n19042),.dinb(w_n18426_0[0]),.dout(n19043),.clk(gclk));
	jand g18744(.dina(w_n19043_0[1]),.dinb(n19040),.dout(n19044),.clk(gclk));
	jor g18745(.dina(w_n19044_0[1]),.dinb(w_n19039_0[1]),.dout(n19045),.clk(gclk));
	jand g18746(.dina(n19045),.dinb(w_asqrt14_11[1]),.dout(n19046),.clk(gclk));
	jor g18747(.dina(w_n19039_0[0]),.dinb(w_asqrt14_11[0]),.dout(n19047),.clk(gclk));
	jor g18748(.dina(n19047),.dinb(w_n19044_0[0]),.dout(n19048),.clk(gclk));
	jnot g18749(.din(w_n18434_0[0]),.dout(n19049),.clk(gclk));
	jnot g18750(.din(w_n18436_0[0]),.dout(n19050),.clk(gclk));
	jand g18751(.dina(w_asqrt4_27[1]),.dinb(w_n18430_0[0]),.dout(n19051),.clk(gclk));
	jand g18752(.dina(w_n19051_0[1]),.dinb(n19050),.dout(n19052),.clk(gclk));
	jor g18753(.dina(n19052),.dinb(n19049),.dout(n19053),.clk(gclk));
	jnot g18754(.din(w_n18437_0[0]),.dout(n19054),.clk(gclk));
	jand g18755(.dina(w_n19051_0[0]),.dinb(n19054),.dout(n19055),.clk(gclk));
	jnot g18756(.din(n19055),.dout(n19056),.clk(gclk));
	jand g18757(.dina(n19056),.dinb(n19053),.dout(n19057),.clk(gclk));
	jand g18758(.dina(w_n19057_0[1]),.dinb(w_n19048_0[1]),.dout(n19058),.clk(gclk));
	jor g18759(.dina(n19058),.dinb(w_n19046_0[1]),.dout(n19059),.clk(gclk));
	jand g18760(.dina(w_n19059_0[1]),.dinb(w_asqrt15_6[2]),.dout(n19060),.clk(gclk));
	jxor g18761(.dina(w_n18438_0[0]),.dinb(w_n13718_4[1]),.dout(n19061),.clk(gclk));
	jand g18762(.dina(n19061),.dinb(w_asqrt4_27[0]),.dout(n19062),.clk(gclk));
	jxor g18763(.dina(n19062),.dinb(w_n18445_0[0]),.dout(n19063),.clk(gclk));
	jnot g18764(.din(n19063),.dout(n19064),.clk(gclk));
	jor g18765(.dina(w_n19059_0[0]),.dinb(w_asqrt15_6[1]),.dout(n19065),.clk(gclk));
	jand g18766(.dina(w_n19065_0[1]),.dinb(w_n19064_0[1]),.dout(n19066),.clk(gclk));
	jor g18767(.dina(w_n19066_0[2]),.dinb(w_n19060_0[2]),.dout(n19067),.clk(gclk));
	jand g18768(.dina(n19067),.dinb(w_asqrt16_11[1]),.dout(n19068),.clk(gclk));
	jnot g18769(.din(w_n18450_0[0]),.dout(n19069),.clk(gclk));
	jand g18770(.dina(n19069),.dinb(w_n18448_0[0]),.dout(n19070),.clk(gclk));
	jand g18771(.dina(n19070),.dinb(w_asqrt4_26[2]),.dout(n19071),.clk(gclk));
	jxor g18772(.dina(n19071),.dinb(w_n18458_0[0]),.dout(n19072),.clk(gclk));
	jnot g18773(.din(n19072),.dout(n19073),.clk(gclk));
	jor g18774(.dina(w_n19060_0[1]),.dinb(w_asqrt16_11[0]),.dout(n19074),.clk(gclk));
	jor g18775(.dina(n19074),.dinb(w_n19066_0[1]),.dout(n19075),.clk(gclk));
	jand g18776(.dina(w_n19075_0[1]),.dinb(w_n19073_0[1]),.dout(n19076),.clk(gclk));
	jor g18777(.dina(w_n19076_0[1]),.dinb(w_n19068_0[1]),.dout(n19077),.clk(gclk));
	jand g18778(.dina(w_n19077_0[2]),.dinb(w_asqrt17_7[0]),.dout(n19078),.clk(gclk));
	jor g18779(.dina(w_n19077_0[1]),.dinb(w_asqrt17_6[2]),.dout(n19079),.clk(gclk));
	jnot g18780(.din(w_n18464_0[0]),.dout(n19080),.clk(gclk));
	jnot g18781(.din(w_n18465_0[0]),.dout(n19081),.clk(gclk));
	jand g18782(.dina(w_asqrt4_26[1]),.dinb(w_n18461_0[0]),.dout(n19082),.clk(gclk));
	jand g18783(.dina(w_n19082_0[1]),.dinb(n19081),.dout(n19083),.clk(gclk));
	jor g18784(.dina(n19083),.dinb(n19080),.dout(n19084),.clk(gclk));
	jnot g18785(.din(w_n18466_0[0]),.dout(n19085),.clk(gclk));
	jand g18786(.dina(w_n19082_0[0]),.dinb(n19085),.dout(n19086),.clk(gclk));
	jnot g18787(.din(n19086),.dout(n19087),.clk(gclk));
	jand g18788(.dina(n19087),.dinb(n19084),.dout(n19088),.clk(gclk));
	jand g18789(.dina(w_n19088_0[1]),.dinb(n19079),.dout(n19089),.clk(gclk));
	jor g18790(.dina(w_n19089_0[1]),.dinb(w_n19078_0[1]),.dout(n19090),.clk(gclk));
	jand g18791(.dina(n19090),.dinb(w_asqrt18_11[1]),.dout(n19091),.clk(gclk));
	jor g18792(.dina(w_n19078_0[0]),.dinb(w_asqrt18_11[0]),.dout(n19092),.clk(gclk));
	jor g18793(.dina(n19092),.dinb(w_n19089_0[0]),.dout(n19093),.clk(gclk));
	jnot g18794(.din(w_n18472_0[0]),.dout(n19094),.clk(gclk));
	jnot g18795(.din(w_n18474_0[0]),.dout(n19095),.clk(gclk));
	jand g18796(.dina(w_asqrt4_26[0]),.dinb(w_n18468_0[0]),.dout(n19096),.clk(gclk));
	jand g18797(.dina(w_n19096_0[1]),.dinb(n19095),.dout(n19097),.clk(gclk));
	jor g18798(.dina(n19097),.dinb(n19094),.dout(n19098),.clk(gclk));
	jnot g18799(.din(w_n18475_0[0]),.dout(n19099),.clk(gclk));
	jand g18800(.dina(w_n19096_0[0]),.dinb(n19099),.dout(n19100),.clk(gclk));
	jnot g18801(.din(n19100),.dout(n19101),.clk(gclk));
	jand g18802(.dina(n19101),.dinb(n19098),.dout(n19102),.clk(gclk));
	jand g18803(.dina(w_n19102_0[1]),.dinb(w_n19093_0[1]),.dout(n19103),.clk(gclk));
	jor g18804(.dina(n19103),.dinb(w_n19091_0[1]),.dout(n19104),.clk(gclk));
	jand g18805(.dina(w_n19104_0[1]),.dinb(w_asqrt19_7[0]),.dout(n19105),.clk(gclk));
	jxor g18806(.dina(w_n18476_0[0]),.dinb(w_n11657_5[0]),.dout(n19106),.clk(gclk));
	jand g18807(.dina(n19106),.dinb(w_asqrt4_25[2]),.dout(n19107),.clk(gclk));
	jxor g18808(.dina(n19107),.dinb(w_n18486_0[0]),.dout(n19108),.clk(gclk));
	jnot g18809(.din(n19108),.dout(n19109),.clk(gclk));
	jor g18810(.dina(w_n19104_0[0]),.dinb(w_asqrt19_6[2]),.dout(n19110),.clk(gclk));
	jand g18811(.dina(w_n19110_0[1]),.dinb(w_n19109_0[1]),.dout(n19111),.clk(gclk));
	jor g18812(.dina(w_n19111_0[2]),.dinb(w_n19105_0[2]),.dout(n19112),.clk(gclk));
	jand g18813(.dina(n19112),.dinb(w_asqrt20_11[1]),.dout(n19113),.clk(gclk));
	jnot g18814(.din(w_n18491_0[0]),.dout(n19114),.clk(gclk));
	jand g18815(.dina(n19114),.dinb(w_n18489_0[0]),.dout(n19115),.clk(gclk));
	jand g18816(.dina(n19115),.dinb(w_asqrt4_25[1]),.dout(n19116),.clk(gclk));
	jxor g18817(.dina(n19116),.dinb(w_n18499_0[0]),.dout(n19117),.clk(gclk));
	jnot g18818(.din(n19117),.dout(n19118),.clk(gclk));
	jor g18819(.dina(w_n19105_0[1]),.dinb(w_asqrt20_11[0]),.dout(n19119),.clk(gclk));
	jor g18820(.dina(n19119),.dinb(w_n19111_0[1]),.dout(n19120),.clk(gclk));
	jand g18821(.dina(w_n19120_0[1]),.dinb(w_n19118_0[1]),.dout(n19121),.clk(gclk));
	jor g18822(.dina(w_n19121_0[1]),.dinb(w_n19113_0[1]),.dout(n19122),.clk(gclk));
	jand g18823(.dina(w_n19122_0[2]),.dinb(w_asqrt21_7[1]),.dout(n19123),.clk(gclk));
	jor g18824(.dina(w_n19122_0[1]),.dinb(w_asqrt21_7[0]),.dout(n19124),.clk(gclk));
	jnot g18825(.din(w_n18505_0[0]),.dout(n19125),.clk(gclk));
	jnot g18826(.din(w_n18506_0[0]),.dout(n19126),.clk(gclk));
	jand g18827(.dina(w_asqrt4_25[0]),.dinb(w_n18502_0[0]),.dout(n19127),.clk(gclk));
	jand g18828(.dina(w_n19127_0[1]),.dinb(n19126),.dout(n19128),.clk(gclk));
	jor g18829(.dina(n19128),.dinb(n19125),.dout(n19129),.clk(gclk));
	jnot g18830(.din(w_n18507_0[0]),.dout(n19130),.clk(gclk));
	jand g18831(.dina(w_n19127_0[0]),.dinb(n19130),.dout(n19131),.clk(gclk));
	jnot g18832(.din(n19131),.dout(n19132),.clk(gclk));
	jand g18833(.dina(n19132),.dinb(n19129),.dout(n19133),.clk(gclk));
	jand g18834(.dina(w_n19133_0[1]),.dinb(n19124),.dout(n19134),.clk(gclk));
	jor g18835(.dina(w_n19134_0[1]),.dinb(w_n19123_0[1]),.dout(n19135),.clk(gclk));
	jand g18836(.dina(n19135),.dinb(w_asqrt22_11[1]),.dout(n19136),.clk(gclk));
	jor g18837(.dina(w_n19123_0[0]),.dinb(w_asqrt22_11[0]),.dout(n19137),.clk(gclk));
	jor g18838(.dina(n19137),.dinb(w_n19134_0[0]),.dout(n19138),.clk(gclk));
	jnot g18839(.din(w_n18513_0[0]),.dout(n19139),.clk(gclk));
	jnot g18840(.din(w_n18515_0[0]),.dout(n19140),.clk(gclk));
	jand g18841(.dina(w_asqrt4_24[2]),.dinb(w_n18509_0[0]),.dout(n19141),.clk(gclk));
	jand g18842(.dina(w_n19141_0[1]),.dinb(n19140),.dout(n19142),.clk(gclk));
	jor g18843(.dina(n19142),.dinb(n19139),.dout(n19143),.clk(gclk));
	jnot g18844(.din(w_n18516_0[0]),.dout(n19144),.clk(gclk));
	jand g18845(.dina(w_n19141_0[0]),.dinb(n19144),.dout(n19145),.clk(gclk));
	jnot g18846(.din(n19145),.dout(n19146),.clk(gclk));
	jand g18847(.dina(n19146),.dinb(n19143),.dout(n19147),.clk(gclk));
	jand g18848(.dina(w_n19147_0[1]),.dinb(w_n19138_0[1]),.dout(n19148),.clk(gclk));
	jor g18849(.dina(n19148),.dinb(w_n19136_0[1]),.dout(n19149),.clk(gclk));
	jand g18850(.dina(w_n19149_0[1]),.dinb(w_asqrt23_7[1]),.dout(n19150),.clk(gclk));
	jxor g18851(.dina(w_n18517_0[0]),.dinb(w_n9769_6[0]),.dout(n19151),.clk(gclk));
	jand g18852(.dina(n19151),.dinb(w_asqrt4_24[1]),.dout(n19152),.clk(gclk));
	jxor g18853(.dina(n19152),.dinb(w_n18527_0[0]),.dout(n19153),.clk(gclk));
	jnot g18854(.din(n19153),.dout(n19154),.clk(gclk));
	jor g18855(.dina(w_n19149_0[0]),.dinb(w_asqrt23_7[0]),.dout(n19155),.clk(gclk));
	jand g18856(.dina(w_n19155_0[1]),.dinb(w_n19154_0[1]),.dout(n19156),.clk(gclk));
	jor g18857(.dina(w_n19156_0[2]),.dinb(w_n19150_0[2]),.dout(n19157),.clk(gclk));
	jand g18858(.dina(n19157),.dinb(w_asqrt24_11[1]),.dout(n19158),.clk(gclk));
	jnot g18859(.din(w_n18532_0[0]),.dout(n19159),.clk(gclk));
	jand g18860(.dina(n19159),.dinb(w_n18530_0[0]),.dout(n19160),.clk(gclk));
	jand g18861(.dina(n19160),.dinb(w_asqrt4_24[0]),.dout(n19161),.clk(gclk));
	jxor g18862(.dina(n19161),.dinb(w_n18540_0[0]),.dout(n19162),.clk(gclk));
	jnot g18863(.din(n19162),.dout(n19163),.clk(gclk));
	jor g18864(.dina(w_n19150_0[1]),.dinb(w_asqrt24_11[0]),.dout(n19164),.clk(gclk));
	jor g18865(.dina(n19164),.dinb(w_n19156_0[1]),.dout(n19165),.clk(gclk));
	jand g18866(.dina(w_n19165_0[1]),.dinb(w_n19163_0[1]),.dout(n19166),.clk(gclk));
	jor g18867(.dina(w_n19166_0[1]),.dinb(w_n19158_0[1]),.dout(n19167),.clk(gclk));
	jand g18868(.dina(w_n19167_0[2]),.dinb(w_asqrt25_7[2]),.dout(n19168),.clk(gclk));
	jor g18869(.dina(w_n19167_0[1]),.dinb(w_asqrt25_7[1]),.dout(n19169),.clk(gclk));
	jnot g18870(.din(w_n18546_0[0]),.dout(n19170),.clk(gclk));
	jnot g18871(.din(w_n18547_0[0]),.dout(n19171),.clk(gclk));
	jand g18872(.dina(w_asqrt4_23[2]),.dinb(w_n18543_0[0]),.dout(n19172),.clk(gclk));
	jand g18873(.dina(w_n19172_0[1]),.dinb(n19171),.dout(n19173),.clk(gclk));
	jor g18874(.dina(n19173),.dinb(n19170),.dout(n19174),.clk(gclk));
	jnot g18875(.din(w_n18548_0[0]),.dout(n19175),.clk(gclk));
	jand g18876(.dina(w_n19172_0[0]),.dinb(n19175),.dout(n19176),.clk(gclk));
	jnot g18877(.din(n19176),.dout(n19177),.clk(gclk));
	jand g18878(.dina(n19177),.dinb(n19174),.dout(n19178),.clk(gclk));
	jand g18879(.dina(w_n19178_0[1]),.dinb(n19169),.dout(n19179),.clk(gclk));
	jor g18880(.dina(w_n19179_0[1]),.dinb(w_n19168_0[1]),.dout(n19180),.clk(gclk));
	jand g18881(.dina(n19180),.dinb(w_asqrt26_11[1]),.dout(n19181),.clk(gclk));
	jor g18882(.dina(w_n19168_0[0]),.dinb(w_asqrt26_11[0]),.dout(n19182),.clk(gclk));
	jor g18883(.dina(n19182),.dinb(w_n19179_0[0]),.dout(n19183),.clk(gclk));
	jnot g18884(.din(w_n18554_0[0]),.dout(n19184),.clk(gclk));
	jnot g18885(.din(w_n18556_0[0]),.dout(n19185),.clk(gclk));
	jand g18886(.dina(w_asqrt4_23[1]),.dinb(w_n18550_0[0]),.dout(n19186),.clk(gclk));
	jand g18887(.dina(w_n19186_0[1]),.dinb(n19185),.dout(n19187),.clk(gclk));
	jor g18888(.dina(n19187),.dinb(n19184),.dout(n19188),.clk(gclk));
	jnot g18889(.din(w_n18557_0[0]),.dout(n19189),.clk(gclk));
	jand g18890(.dina(w_n19186_0[0]),.dinb(n19189),.dout(n19190),.clk(gclk));
	jnot g18891(.din(n19190),.dout(n19191),.clk(gclk));
	jand g18892(.dina(n19191),.dinb(n19188),.dout(n19192),.clk(gclk));
	jand g18893(.dina(w_n19192_0[1]),.dinb(w_n19183_0[1]),.dout(n19193),.clk(gclk));
	jor g18894(.dina(n19193),.dinb(w_n19181_0[1]),.dout(n19194),.clk(gclk));
	jand g18895(.dina(w_n19194_0[1]),.dinb(w_asqrt27_7[2]),.dout(n19195),.clk(gclk));
	jxor g18896(.dina(w_n18558_0[0]),.dinb(w_n8053_6[2]),.dout(n19196),.clk(gclk));
	jand g18897(.dina(n19196),.dinb(w_asqrt4_23[0]),.dout(n19197),.clk(gclk));
	jxor g18898(.dina(n19197),.dinb(w_n18568_0[0]),.dout(n19198),.clk(gclk));
	jnot g18899(.din(n19198),.dout(n19199),.clk(gclk));
	jor g18900(.dina(w_n19194_0[0]),.dinb(w_asqrt27_7[1]),.dout(n19200),.clk(gclk));
	jand g18901(.dina(w_n19200_0[1]),.dinb(w_n19199_0[1]),.dout(n19201),.clk(gclk));
	jor g18902(.dina(w_n19201_0[2]),.dinb(w_n19195_0[2]),.dout(n19202),.clk(gclk));
	jand g18903(.dina(n19202),.dinb(w_asqrt28_11[1]),.dout(n19203),.clk(gclk));
	jnot g18904(.din(w_n18573_0[0]),.dout(n19204),.clk(gclk));
	jand g18905(.dina(n19204),.dinb(w_n18571_0[0]),.dout(n19205),.clk(gclk));
	jand g18906(.dina(n19205),.dinb(w_asqrt4_22[2]),.dout(n19206),.clk(gclk));
	jxor g18907(.dina(n19206),.dinb(w_n18581_0[0]),.dout(n19207),.clk(gclk));
	jnot g18908(.din(n19207),.dout(n19208),.clk(gclk));
	jor g18909(.dina(w_n19195_0[1]),.dinb(w_asqrt28_11[0]),.dout(n19209),.clk(gclk));
	jor g18910(.dina(n19209),.dinb(w_n19201_0[1]),.dout(n19210),.clk(gclk));
	jand g18911(.dina(w_n19210_0[1]),.dinb(w_n19208_0[1]),.dout(n19211),.clk(gclk));
	jor g18912(.dina(w_n19211_0[1]),.dinb(w_n19203_0[1]),.dout(n19212),.clk(gclk));
	jand g18913(.dina(w_n19212_0[2]),.dinb(w_asqrt29_8[0]),.dout(n19213),.clk(gclk));
	jor g18914(.dina(w_n19212_0[1]),.dinb(w_asqrt29_7[2]),.dout(n19214),.clk(gclk));
	jnot g18915(.din(w_n18587_0[0]),.dout(n19215),.clk(gclk));
	jnot g18916(.din(w_n18588_0[0]),.dout(n19216),.clk(gclk));
	jand g18917(.dina(w_asqrt4_22[1]),.dinb(w_n18584_0[0]),.dout(n19217),.clk(gclk));
	jand g18918(.dina(w_n19217_0[1]),.dinb(n19216),.dout(n19218),.clk(gclk));
	jor g18919(.dina(n19218),.dinb(n19215),.dout(n19219),.clk(gclk));
	jnot g18920(.din(w_n18589_0[0]),.dout(n19220),.clk(gclk));
	jand g18921(.dina(w_n19217_0[0]),.dinb(n19220),.dout(n19221),.clk(gclk));
	jnot g18922(.din(n19221),.dout(n19222),.clk(gclk));
	jand g18923(.dina(n19222),.dinb(n19219),.dout(n19223),.clk(gclk));
	jand g18924(.dina(w_n19223_0[1]),.dinb(n19214),.dout(n19224),.clk(gclk));
	jor g18925(.dina(w_n19224_0[1]),.dinb(w_n19213_0[1]),.dout(n19225),.clk(gclk));
	jand g18926(.dina(n19225),.dinb(w_asqrt30_11[1]),.dout(n19226),.clk(gclk));
	jor g18927(.dina(w_n19213_0[0]),.dinb(w_asqrt30_11[0]),.dout(n19227),.clk(gclk));
	jor g18928(.dina(n19227),.dinb(w_n19224_0[0]),.dout(n19228),.clk(gclk));
	jnot g18929(.din(w_n18595_0[0]),.dout(n19229),.clk(gclk));
	jnot g18930(.din(w_n18597_0[0]),.dout(n19230),.clk(gclk));
	jand g18931(.dina(w_asqrt4_22[0]),.dinb(w_n18591_0[0]),.dout(n19231),.clk(gclk));
	jand g18932(.dina(w_n19231_0[1]),.dinb(n19230),.dout(n19232),.clk(gclk));
	jor g18933(.dina(n19232),.dinb(n19229),.dout(n19233),.clk(gclk));
	jnot g18934(.din(w_n18598_0[0]),.dout(n19234),.clk(gclk));
	jand g18935(.dina(w_n19231_0[0]),.dinb(n19234),.dout(n19235),.clk(gclk));
	jnot g18936(.din(n19235),.dout(n19236),.clk(gclk));
	jand g18937(.dina(n19236),.dinb(n19233),.dout(n19237),.clk(gclk));
	jand g18938(.dina(w_n19237_0[1]),.dinb(w_n19228_0[1]),.dout(n19238),.clk(gclk));
	jor g18939(.dina(n19238),.dinb(w_n19226_0[1]),.dout(n19239),.clk(gclk));
	jand g18940(.dina(w_n19239_0[1]),.dinb(w_asqrt31_8[0]),.dout(n19240),.clk(gclk));
	jxor g18941(.dina(w_n18599_0[0]),.dinb(w_n6500_7[2]),.dout(n19241),.clk(gclk));
	jand g18942(.dina(n19241),.dinb(w_asqrt4_21[2]),.dout(n19242),.clk(gclk));
	jxor g18943(.dina(n19242),.dinb(w_n18609_0[0]),.dout(n19243),.clk(gclk));
	jnot g18944(.din(n19243),.dout(n19244),.clk(gclk));
	jor g18945(.dina(w_n19239_0[0]),.dinb(w_asqrt31_7[2]),.dout(n19245),.clk(gclk));
	jand g18946(.dina(w_n19245_0[1]),.dinb(w_n19244_0[1]),.dout(n19246),.clk(gclk));
	jor g18947(.dina(w_n19246_0[2]),.dinb(w_n19240_0[2]),.dout(n19247),.clk(gclk));
	jand g18948(.dina(n19247),.dinb(w_asqrt32_11[1]),.dout(n19248),.clk(gclk));
	jnot g18949(.din(w_n18614_0[0]),.dout(n19249),.clk(gclk));
	jand g18950(.dina(n19249),.dinb(w_n18612_0[0]),.dout(n19250),.clk(gclk));
	jand g18951(.dina(n19250),.dinb(w_asqrt4_21[1]),.dout(n19251),.clk(gclk));
	jxor g18952(.dina(n19251),.dinb(w_n18622_0[0]),.dout(n19252),.clk(gclk));
	jnot g18953(.din(n19252),.dout(n19253),.clk(gclk));
	jor g18954(.dina(w_n19240_0[1]),.dinb(w_asqrt32_11[0]),.dout(n19254),.clk(gclk));
	jor g18955(.dina(n19254),.dinb(w_n19246_0[1]),.dout(n19255),.clk(gclk));
	jand g18956(.dina(w_n19255_0[1]),.dinb(w_n19253_0[1]),.dout(n19256),.clk(gclk));
	jor g18957(.dina(w_n19256_0[1]),.dinb(w_n19248_0[1]),.dout(n19257),.clk(gclk));
	jand g18958(.dina(w_n19257_0[2]),.dinb(w_asqrt33_8[1]),.dout(n19258),.clk(gclk));
	jor g18959(.dina(w_n19257_0[1]),.dinb(w_asqrt33_8[0]),.dout(n19259),.clk(gclk));
	jnot g18960(.din(w_n18628_0[0]),.dout(n19260),.clk(gclk));
	jnot g18961(.din(w_n18629_0[0]),.dout(n19261),.clk(gclk));
	jand g18962(.dina(w_asqrt4_21[0]),.dinb(w_n18625_0[0]),.dout(n19262),.clk(gclk));
	jand g18963(.dina(w_n19262_0[1]),.dinb(n19261),.dout(n19263),.clk(gclk));
	jor g18964(.dina(n19263),.dinb(n19260),.dout(n19264),.clk(gclk));
	jnot g18965(.din(w_n18630_0[0]),.dout(n19265),.clk(gclk));
	jand g18966(.dina(w_n19262_0[0]),.dinb(n19265),.dout(n19266),.clk(gclk));
	jnot g18967(.din(n19266),.dout(n19267),.clk(gclk));
	jand g18968(.dina(n19267),.dinb(n19264),.dout(n19268),.clk(gclk));
	jand g18969(.dina(w_n19268_0[1]),.dinb(n19259),.dout(n19269),.clk(gclk));
	jor g18970(.dina(w_n19269_0[1]),.dinb(w_n19258_0[1]),.dout(n19270),.clk(gclk));
	jand g18971(.dina(n19270),.dinb(w_asqrt34_11[1]),.dout(n19271),.clk(gclk));
	jor g18972(.dina(w_n19258_0[0]),.dinb(w_asqrt34_11[0]),.dout(n19272),.clk(gclk));
	jor g18973(.dina(n19272),.dinb(w_n19269_0[0]),.dout(n19273),.clk(gclk));
	jnot g18974(.din(w_n18636_0[0]),.dout(n19274),.clk(gclk));
	jnot g18975(.din(w_n18638_0[0]),.dout(n19275),.clk(gclk));
	jand g18976(.dina(w_asqrt4_20[2]),.dinb(w_n18632_0[0]),.dout(n19276),.clk(gclk));
	jand g18977(.dina(w_n19276_0[1]),.dinb(n19275),.dout(n19277),.clk(gclk));
	jor g18978(.dina(n19277),.dinb(n19274),.dout(n19278),.clk(gclk));
	jnot g18979(.din(w_n18639_0[0]),.dout(n19279),.clk(gclk));
	jand g18980(.dina(w_n19276_0[0]),.dinb(n19279),.dout(n19280),.clk(gclk));
	jnot g18981(.din(n19280),.dout(n19281),.clk(gclk));
	jand g18982(.dina(n19281),.dinb(n19278),.dout(n19282),.clk(gclk));
	jand g18983(.dina(w_n19282_0[1]),.dinb(w_n19273_0[1]),.dout(n19283),.clk(gclk));
	jor g18984(.dina(n19283),.dinb(w_n19271_0[1]),.dout(n19284),.clk(gclk));
	jand g18985(.dina(w_n19284_0[1]),.dinb(w_asqrt35_8[1]),.dout(n19285),.clk(gclk));
	jxor g18986(.dina(w_n18640_0[0]),.dinb(w_n5116_8[1]),.dout(n19286),.clk(gclk));
	jand g18987(.dina(n19286),.dinb(w_asqrt4_20[1]),.dout(n19287),.clk(gclk));
	jxor g18988(.dina(n19287),.dinb(w_n18650_0[0]),.dout(n19288),.clk(gclk));
	jnot g18989(.din(n19288),.dout(n19289),.clk(gclk));
	jor g18990(.dina(w_n19284_0[0]),.dinb(w_asqrt35_8[0]),.dout(n19290),.clk(gclk));
	jand g18991(.dina(w_n19290_0[1]),.dinb(w_n19289_0[1]),.dout(n19291),.clk(gclk));
	jor g18992(.dina(w_n19291_0[2]),.dinb(w_n19285_0[2]),.dout(n19292),.clk(gclk));
	jand g18993(.dina(n19292),.dinb(w_asqrt36_11[1]),.dout(n19293),.clk(gclk));
	jnot g18994(.din(w_n18655_0[0]),.dout(n19294),.clk(gclk));
	jand g18995(.dina(n19294),.dinb(w_n18653_0[0]),.dout(n19295),.clk(gclk));
	jand g18996(.dina(n19295),.dinb(w_asqrt4_20[0]),.dout(n19296),.clk(gclk));
	jxor g18997(.dina(n19296),.dinb(w_n18663_0[0]),.dout(n19297),.clk(gclk));
	jnot g18998(.din(n19297),.dout(n19298),.clk(gclk));
	jor g18999(.dina(w_n19285_0[1]),.dinb(w_asqrt36_11[0]),.dout(n19299),.clk(gclk));
	jor g19000(.dina(n19299),.dinb(w_n19291_0[1]),.dout(n19300),.clk(gclk));
	jand g19001(.dina(w_n19300_0[1]),.dinb(w_n19298_0[1]),.dout(n19301),.clk(gclk));
	jor g19002(.dina(w_n19301_0[1]),.dinb(w_n19293_0[1]),.dout(n19302),.clk(gclk));
	jand g19003(.dina(w_n19302_0[2]),.dinb(w_asqrt37_8[2]),.dout(n19303),.clk(gclk));
	jor g19004(.dina(w_n19302_0[1]),.dinb(w_asqrt37_8[1]),.dout(n19304),.clk(gclk));
	jnot g19005(.din(w_n18669_0[0]),.dout(n19305),.clk(gclk));
	jnot g19006(.din(w_n18670_0[0]),.dout(n19306),.clk(gclk));
	jand g19007(.dina(w_asqrt4_19[2]),.dinb(w_n18666_0[0]),.dout(n19307),.clk(gclk));
	jand g19008(.dina(w_n19307_0[1]),.dinb(n19306),.dout(n19308),.clk(gclk));
	jor g19009(.dina(n19308),.dinb(n19305),.dout(n19309),.clk(gclk));
	jnot g19010(.din(w_n18671_0[0]),.dout(n19310),.clk(gclk));
	jand g19011(.dina(w_n19307_0[0]),.dinb(n19310),.dout(n19311),.clk(gclk));
	jnot g19012(.din(n19311),.dout(n19312),.clk(gclk));
	jand g19013(.dina(n19312),.dinb(n19309),.dout(n19313),.clk(gclk));
	jand g19014(.dina(w_n19313_0[1]),.dinb(n19304),.dout(n19314),.clk(gclk));
	jor g19015(.dina(w_n19314_0[1]),.dinb(w_n19303_0[1]),.dout(n19315),.clk(gclk));
	jand g19016(.dina(n19315),.dinb(w_asqrt38_11[1]),.dout(n19316),.clk(gclk));
	jor g19017(.dina(w_n19303_0[0]),.dinb(w_asqrt38_11[0]),.dout(n19317),.clk(gclk));
	jor g19018(.dina(n19317),.dinb(w_n19314_0[0]),.dout(n19318),.clk(gclk));
	jnot g19019(.din(w_n18677_0[0]),.dout(n19319),.clk(gclk));
	jnot g19020(.din(w_n18679_0[0]),.dout(n19320),.clk(gclk));
	jand g19021(.dina(w_asqrt4_19[1]),.dinb(w_n18673_0[0]),.dout(n19321),.clk(gclk));
	jand g19022(.dina(w_n19321_0[1]),.dinb(n19320),.dout(n19322),.clk(gclk));
	jor g19023(.dina(n19322),.dinb(n19319),.dout(n19323),.clk(gclk));
	jnot g19024(.din(w_n18680_0[0]),.dout(n19324),.clk(gclk));
	jand g19025(.dina(w_n19321_0[0]),.dinb(n19324),.dout(n19325),.clk(gclk));
	jnot g19026(.din(n19325),.dout(n19326),.clk(gclk));
	jand g19027(.dina(n19326),.dinb(n19323),.dout(n19327),.clk(gclk));
	jand g19028(.dina(w_n19327_0[1]),.dinb(w_n19318_0[1]),.dout(n19328),.clk(gclk));
	jor g19029(.dina(n19328),.dinb(w_n19316_0[1]),.dout(n19329),.clk(gclk));
	jand g19030(.dina(w_n19329_0[1]),.dinb(w_asqrt39_8[2]),.dout(n19330),.clk(gclk));
	jxor g19031(.dina(w_n18681_0[0]),.dinb(w_n3907_9[1]),.dout(n19331),.clk(gclk));
	jand g19032(.dina(n19331),.dinb(w_asqrt4_19[0]),.dout(n19332),.clk(gclk));
	jxor g19033(.dina(n19332),.dinb(w_n18691_0[0]),.dout(n19333),.clk(gclk));
	jnot g19034(.din(n19333),.dout(n19334),.clk(gclk));
	jor g19035(.dina(w_n19329_0[0]),.dinb(w_asqrt39_8[1]),.dout(n19335),.clk(gclk));
	jand g19036(.dina(w_n19335_0[1]),.dinb(w_n19334_0[1]),.dout(n19336),.clk(gclk));
	jor g19037(.dina(w_n19336_0[2]),.dinb(w_n19330_0[2]),.dout(n19337),.clk(gclk));
	jand g19038(.dina(n19337),.dinb(w_asqrt40_11[1]),.dout(n19338),.clk(gclk));
	jnot g19039(.din(w_n18696_0[0]),.dout(n19339),.clk(gclk));
	jand g19040(.dina(n19339),.dinb(w_n18694_0[0]),.dout(n19340),.clk(gclk));
	jand g19041(.dina(n19340),.dinb(w_asqrt4_18[2]),.dout(n19341),.clk(gclk));
	jxor g19042(.dina(n19341),.dinb(w_n18704_0[0]),.dout(n19342),.clk(gclk));
	jnot g19043(.din(n19342),.dout(n19343),.clk(gclk));
	jor g19044(.dina(w_n19330_0[1]),.dinb(w_asqrt40_11[0]),.dout(n19344),.clk(gclk));
	jor g19045(.dina(n19344),.dinb(w_n19336_0[1]),.dout(n19345),.clk(gclk));
	jand g19046(.dina(w_n19345_0[1]),.dinb(w_n19343_0[1]),.dout(n19346),.clk(gclk));
	jor g19047(.dina(w_n19346_0[1]),.dinb(w_n19338_0[1]),.dout(n19347),.clk(gclk));
	jand g19048(.dina(w_n19347_0[2]),.dinb(w_asqrt41_9[0]),.dout(n19348),.clk(gclk));
	jor g19049(.dina(w_n19347_0[1]),.dinb(w_asqrt41_8[2]),.dout(n19349),.clk(gclk));
	jnot g19050(.din(w_n18710_0[0]),.dout(n19350),.clk(gclk));
	jnot g19051(.din(w_n18711_0[0]),.dout(n19351),.clk(gclk));
	jand g19052(.dina(w_asqrt4_18[1]),.dinb(w_n18707_0[0]),.dout(n19352),.clk(gclk));
	jand g19053(.dina(w_n19352_0[1]),.dinb(n19351),.dout(n19353),.clk(gclk));
	jor g19054(.dina(n19353),.dinb(n19350),.dout(n19354),.clk(gclk));
	jnot g19055(.din(w_n18712_0[0]),.dout(n19355),.clk(gclk));
	jand g19056(.dina(w_n19352_0[0]),.dinb(n19355),.dout(n19356),.clk(gclk));
	jnot g19057(.din(n19356),.dout(n19357),.clk(gclk));
	jand g19058(.dina(n19357),.dinb(n19354),.dout(n19358),.clk(gclk));
	jand g19059(.dina(w_n19358_0[1]),.dinb(n19349),.dout(n19359),.clk(gclk));
	jor g19060(.dina(w_n19359_0[1]),.dinb(w_n19348_0[1]),.dout(n19360),.clk(gclk));
	jand g19061(.dina(n19360),.dinb(w_asqrt42_11[1]),.dout(n19361),.clk(gclk));
	jor g19062(.dina(w_n19348_0[0]),.dinb(w_asqrt42_11[0]),.dout(n19362),.clk(gclk));
	jor g19063(.dina(n19362),.dinb(w_n19359_0[0]),.dout(n19363),.clk(gclk));
	jnot g19064(.din(w_n18718_0[0]),.dout(n19364),.clk(gclk));
	jnot g19065(.din(w_n18720_0[0]),.dout(n19365),.clk(gclk));
	jand g19066(.dina(w_asqrt4_18[0]),.dinb(w_n18714_0[0]),.dout(n19366),.clk(gclk));
	jand g19067(.dina(w_n19366_0[1]),.dinb(n19365),.dout(n19367),.clk(gclk));
	jor g19068(.dina(n19367),.dinb(n19364),.dout(n19368),.clk(gclk));
	jnot g19069(.din(w_n18721_0[0]),.dout(n19369),.clk(gclk));
	jand g19070(.dina(w_n19366_0[0]),.dinb(n19369),.dout(n19370),.clk(gclk));
	jnot g19071(.din(n19370),.dout(n19371),.clk(gclk));
	jand g19072(.dina(n19371),.dinb(n19368),.dout(n19372),.clk(gclk));
	jand g19073(.dina(w_n19372_0[1]),.dinb(w_n19363_0[1]),.dout(n19373),.clk(gclk));
	jor g19074(.dina(n19373),.dinb(w_n19361_0[1]),.dout(n19374),.clk(gclk));
	jand g19075(.dina(w_n19374_0[1]),.dinb(w_asqrt43_9[0]),.dout(n19375),.clk(gclk));
	jxor g19076(.dina(w_n18722_0[0]),.dinb(w_n2870_10[0]),.dout(n19376),.clk(gclk));
	jand g19077(.dina(n19376),.dinb(w_asqrt4_17[2]),.dout(n19377),.clk(gclk));
	jxor g19078(.dina(n19377),.dinb(w_n18732_0[0]),.dout(n19378),.clk(gclk));
	jnot g19079(.din(n19378),.dout(n19379),.clk(gclk));
	jor g19080(.dina(w_n19374_0[0]),.dinb(w_asqrt43_8[2]),.dout(n19380),.clk(gclk));
	jand g19081(.dina(w_n19380_0[1]),.dinb(w_n19379_0[1]),.dout(n19381),.clk(gclk));
	jor g19082(.dina(w_n19381_0[2]),.dinb(w_n19375_0[2]),.dout(n19382),.clk(gclk));
	jand g19083(.dina(n19382),.dinb(w_asqrt44_11[1]),.dout(n19383),.clk(gclk));
	jnot g19084(.din(w_n18737_0[0]),.dout(n19384),.clk(gclk));
	jand g19085(.dina(n19384),.dinb(w_n18735_0[0]),.dout(n19385),.clk(gclk));
	jand g19086(.dina(n19385),.dinb(w_asqrt4_17[1]),.dout(n19386),.clk(gclk));
	jxor g19087(.dina(n19386),.dinb(w_n18745_0[0]),.dout(n19387),.clk(gclk));
	jnot g19088(.din(n19387),.dout(n19388),.clk(gclk));
	jor g19089(.dina(w_n19375_0[1]),.dinb(w_asqrt44_11[0]),.dout(n19389),.clk(gclk));
	jor g19090(.dina(n19389),.dinb(w_n19381_0[1]),.dout(n19390),.clk(gclk));
	jand g19091(.dina(w_n19390_0[1]),.dinb(w_n19388_0[1]),.dout(n19391),.clk(gclk));
	jor g19092(.dina(w_n19391_0[1]),.dinb(w_n19383_0[1]),.dout(n19392),.clk(gclk));
	jand g19093(.dina(w_n19392_0[2]),.dinb(w_asqrt45_9[1]),.dout(n19393),.clk(gclk));
	jor g19094(.dina(w_n19392_0[1]),.dinb(w_asqrt45_9[0]),.dout(n19394),.clk(gclk));
	jnot g19095(.din(w_n18751_0[0]),.dout(n19395),.clk(gclk));
	jnot g19096(.din(w_n18752_0[0]),.dout(n19396),.clk(gclk));
	jand g19097(.dina(w_asqrt4_17[0]),.dinb(w_n18748_0[0]),.dout(n19397),.clk(gclk));
	jand g19098(.dina(w_n19397_0[1]),.dinb(n19396),.dout(n19398),.clk(gclk));
	jor g19099(.dina(n19398),.dinb(n19395),.dout(n19399),.clk(gclk));
	jnot g19100(.din(w_n18753_0[0]),.dout(n19400),.clk(gclk));
	jand g19101(.dina(w_n19397_0[0]),.dinb(n19400),.dout(n19401),.clk(gclk));
	jnot g19102(.din(n19401),.dout(n19402),.clk(gclk));
	jand g19103(.dina(n19402),.dinb(n19399),.dout(n19403),.clk(gclk));
	jand g19104(.dina(w_n19403_0[1]),.dinb(n19394),.dout(n19404),.clk(gclk));
	jor g19105(.dina(w_n19404_0[1]),.dinb(w_n19393_0[1]),.dout(n19405),.clk(gclk));
	jand g19106(.dina(n19405),.dinb(w_asqrt46_11[1]),.dout(n19406),.clk(gclk));
	jor g19107(.dina(w_n19393_0[0]),.dinb(w_asqrt46_11[0]),.dout(n19407),.clk(gclk));
	jor g19108(.dina(n19407),.dinb(w_n19404_0[0]),.dout(n19408),.clk(gclk));
	jnot g19109(.din(w_n18759_0[0]),.dout(n19409),.clk(gclk));
	jnot g19110(.din(w_n18761_0[0]),.dout(n19410),.clk(gclk));
	jand g19111(.dina(w_asqrt4_16[2]),.dinb(w_n18755_0[0]),.dout(n19411),.clk(gclk));
	jand g19112(.dina(w_n19411_0[1]),.dinb(n19410),.dout(n19412),.clk(gclk));
	jor g19113(.dina(n19412),.dinb(n19409),.dout(n19413),.clk(gclk));
	jnot g19114(.din(w_n18762_0[0]),.dout(n19414),.clk(gclk));
	jand g19115(.dina(w_n19411_0[0]),.dinb(n19414),.dout(n19415),.clk(gclk));
	jnot g19116(.din(n19415),.dout(n19416),.clk(gclk));
	jand g19117(.dina(n19416),.dinb(n19413),.dout(n19417),.clk(gclk));
	jand g19118(.dina(w_n19417_0[1]),.dinb(w_n19408_0[1]),.dout(n19418),.clk(gclk));
	jor g19119(.dina(n19418),.dinb(w_n19406_0[1]),.dout(n19419),.clk(gclk));
	jand g19120(.dina(w_n19419_0[1]),.dinb(w_asqrt47_9[1]),.dout(n19420),.clk(gclk));
	jxor g19121(.dina(w_n18763_0[0]),.dinb(w_n2005_11[0]),.dout(n19421),.clk(gclk));
	jand g19122(.dina(n19421),.dinb(w_asqrt4_16[1]),.dout(n19422),.clk(gclk));
	jxor g19123(.dina(n19422),.dinb(w_n18773_0[0]),.dout(n19423),.clk(gclk));
	jnot g19124(.din(n19423),.dout(n19424),.clk(gclk));
	jor g19125(.dina(w_n19419_0[0]),.dinb(w_asqrt47_9[0]),.dout(n19425),.clk(gclk));
	jand g19126(.dina(w_n19425_0[1]),.dinb(w_n19424_0[1]),.dout(n19426),.clk(gclk));
	jor g19127(.dina(w_n19426_0[2]),.dinb(w_n19420_0[2]),.dout(n19427),.clk(gclk));
	jand g19128(.dina(n19427),.dinb(w_asqrt48_11[1]),.dout(n19428),.clk(gclk));
	jnot g19129(.din(w_n18778_0[0]),.dout(n19429),.clk(gclk));
	jand g19130(.dina(n19429),.dinb(w_n18776_0[0]),.dout(n19430),.clk(gclk));
	jand g19131(.dina(n19430),.dinb(w_asqrt4_16[0]),.dout(n19431),.clk(gclk));
	jxor g19132(.dina(n19431),.dinb(w_n18786_0[0]),.dout(n19432),.clk(gclk));
	jnot g19133(.din(n19432),.dout(n19433),.clk(gclk));
	jor g19134(.dina(w_n19420_0[1]),.dinb(w_asqrt48_11[0]),.dout(n19434),.clk(gclk));
	jor g19135(.dina(n19434),.dinb(w_n19426_0[1]),.dout(n19435),.clk(gclk));
	jand g19136(.dina(w_n19435_0[1]),.dinb(w_n19433_0[1]),.dout(n19436),.clk(gclk));
	jor g19137(.dina(w_n19436_0[1]),.dinb(w_n19428_0[1]),.dout(n19437),.clk(gclk));
	jand g19138(.dina(w_n19437_0[2]),.dinb(w_asqrt49_9[2]),.dout(n19438),.clk(gclk));
	jor g19139(.dina(w_n19437_0[1]),.dinb(w_asqrt49_9[1]),.dout(n19439),.clk(gclk));
	jnot g19140(.din(w_n18792_0[0]),.dout(n19440),.clk(gclk));
	jnot g19141(.din(w_n18793_0[0]),.dout(n19441),.clk(gclk));
	jand g19142(.dina(w_asqrt4_15[2]),.dinb(w_n18789_0[0]),.dout(n19442),.clk(gclk));
	jand g19143(.dina(w_n19442_0[1]),.dinb(n19441),.dout(n19443),.clk(gclk));
	jor g19144(.dina(n19443),.dinb(n19440),.dout(n19444),.clk(gclk));
	jnot g19145(.din(w_n18794_0[0]),.dout(n19445),.clk(gclk));
	jand g19146(.dina(w_n19442_0[0]),.dinb(n19445),.dout(n19446),.clk(gclk));
	jnot g19147(.din(n19446),.dout(n19447),.clk(gclk));
	jand g19148(.dina(n19447),.dinb(n19444),.dout(n19448),.clk(gclk));
	jand g19149(.dina(w_n19448_0[1]),.dinb(n19439),.dout(n19449),.clk(gclk));
	jor g19150(.dina(w_n19449_0[1]),.dinb(w_n19438_0[1]),.dout(n19450),.clk(gclk));
	jand g19151(.dina(n19450),.dinb(w_asqrt50_11[1]),.dout(n19451),.clk(gclk));
	jor g19152(.dina(w_n19438_0[0]),.dinb(w_asqrt50_11[0]),.dout(n19452),.clk(gclk));
	jor g19153(.dina(n19452),.dinb(w_n19449_0[0]),.dout(n19453),.clk(gclk));
	jnot g19154(.din(w_n18800_0[0]),.dout(n19454),.clk(gclk));
	jnot g19155(.din(w_n18802_0[0]),.dout(n19455),.clk(gclk));
	jand g19156(.dina(w_asqrt4_15[1]),.dinb(w_n18796_0[0]),.dout(n19456),.clk(gclk));
	jand g19157(.dina(w_n19456_0[1]),.dinb(n19455),.dout(n19457),.clk(gclk));
	jor g19158(.dina(n19457),.dinb(n19454),.dout(n19458),.clk(gclk));
	jnot g19159(.din(w_n18803_0[0]),.dout(n19459),.clk(gclk));
	jand g19160(.dina(w_n19456_0[0]),.dinb(n19459),.dout(n19460),.clk(gclk));
	jnot g19161(.din(n19460),.dout(n19461),.clk(gclk));
	jand g19162(.dina(n19461),.dinb(n19458),.dout(n19462),.clk(gclk));
	jand g19163(.dina(w_n19462_0[1]),.dinb(w_n19453_0[1]),.dout(n19463),.clk(gclk));
	jor g19164(.dina(n19463),.dinb(w_n19451_0[1]),.dout(n19464),.clk(gclk));
	jand g19165(.dina(w_n19464_0[1]),.dinb(w_asqrt51_9[2]),.dout(n19465),.clk(gclk));
	jxor g19166(.dina(w_n18804_0[0]),.dinb(w_n1312_11[2]),.dout(n19466),.clk(gclk));
	jand g19167(.dina(n19466),.dinb(w_asqrt4_15[0]),.dout(n19467),.clk(gclk));
	jxor g19168(.dina(n19467),.dinb(w_n18814_0[0]),.dout(n19468),.clk(gclk));
	jnot g19169(.din(n19468),.dout(n19469),.clk(gclk));
	jor g19170(.dina(w_n19464_0[0]),.dinb(w_asqrt51_9[1]),.dout(n19470),.clk(gclk));
	jand g19171(.dina(w_n19470_0[1]),.dinb(w_n19469_0[1]),.dout(n19471),.clk(gclk));
	jor g19172(.dina(w_n19471_0[2]),.dinb(w_n19465_0[2]),.dout(n19472),.clk(gclk));
	jand g19173(.dina(n19472),.dinb(w_asqrt52_11[1]),.dout(n19473),.clk(gclk));
	jnot g19174(.din(w_n18819_0[0]),.dout(n19474),.clk(gclk));
	jand g19175(.dina(n19474),.dinb(w_n18817_0[0]),.dout(n19475),.clk(gclk));
	jand g19176(.dina(n19475),.dinb(w_asqrt4_14[2]),.dout(n19476),.clk(gclk));
	jxor g19177(.dina(n19476),.dinb(w_n18827_0[0]),.dout(n19477),.clk(gclk));
	jnot g19178(.din(n19477),.dout(n19478),.clk(gclk));
	jor g19179(.dina(w_n19465_0[1]),.dinb(w_asqrt52_11[0]),.dout(n19479),.clk(gclk));
	jor g19180(.dina(n19479),.dinb(w_n19471_0[1]),.dout(n19480),.clk(gclk));
	jand g19181(.dina(w_n19480_0[1]),.dinb(w_n19478_0[1]),.dout(n19481),.clk(gclk));
	jor g19182(.dina(w_n19481_0[1]),.dinb(w_n19473_0[1]),.dout(n19482),.clk(gclk));
	jand g19183(.dina(w_n19482_0[2]),.dinb(w_asqrt53_10[0]),.dout(n19483),.clk(gclk));
	jor g19184(.dina(w_n19482_0[1]),.dinb(w_asqrt53_9[2]),.dout(n19484),.clk(gclk));
	jnot g19185(.din(w_n18833_0[0]),.dout(n19485),.clk(gclk));
	jnot g19186(.din(w_n18834_0[0]),.dout(n19486),.clk(gclk));
	jand g19187(.dina(w_asqrt4_14[1]),.dinb(w_n18830_0[0]),.dout(n19487),.clk(gclk));
	jand g19188(.dina(w_n19487_0[1]),.dinb(n19486),.dout(n19488),.clk(gclk));
	jor g19189(.dina(n19488),.dinb(n19485),.dout(n19489),.clk(gclk));
	jnot g19190(.din(w_n18835_0[0]),.dout(n19490),.clk(gclk));
	jand g19191(.dina(w_n19487_0[0]),.dinb(n19490),.dout(n19491),.clk(gclk));
	jnot g19192(.din(n19491),.dout(n19492),.clk(gclk));
	jand g19193(.dina(n19492),.dinb(n19489),.dout(n19493),.clk(gclk));
	jand g19194(.dina(w_n19493_0[1]),.dinb(n19484),.dout(n19494),.clk(gclk));
	jor g19195(.dina(w_n19494_0[1]),.dinb(w_n19483_0[1]),.dout(n19495),.clk(gclk));
	jand g19196(.dina(n19495),.dinb(w_asqrt54_11[1]),.dout(n19496),.clk(gclk));
	jor g19197(.dina(w_n19483_0[0]),.dinb(w_asqrt54_11[0]),.dout(n19497),.clk(gclk));
	jor g19198(.dina(n19497),.dinb(w_n19494_0[0]),.dout(n19498),.clk(gclk));
	jnot g19199(.din(w_n18841_0[0]),.dout(n19499),.clk(gclk));
	jnot g19200(.din(w_n18843_0[0]),.dout(n19500),.clk(gclk));
	jand g19201(.dina(w_asqrt4_14[0]),.dinb(w_n18837_0[0]),.dout(n19501),.clk(gclk));
	jand g19202(.dina(w_n19501_0[1]),.dinb(n19500),.dout(n19502),.clk(gclk));
	jor g19203(.dina(n19502),.dinb(n19499),.dout(n19503),.clk(gclk));
	jnot g19204(.din(w_n18844_0[0]),.dout(n19504),.clk(gclk));
	jand g19205(.dina(w_n19501_0[0]),.dinb(n19504),.dout(n19505),.clk(gclk));
	jnot g19206(.din(n19505),.dout(n19506),.clk(gclk));
	jand g19207(.dina(n19506),.dinb(n19503),.dout(n19507),.clk(gclk));
	jand g19208(.dina(w_n19507_0[1]),.dinb(w_n19498_0[1]),.dout(n19508),.clk(gclk));
	jor g19209(.dina(n19508),.dinb(w_n19496_0[1]),.dout(n19509),.clk(gclk));
	jand g19210(.dina(w_n19509_0[1]),.dinb(w_asqrt55_10[1]),.dout(n19510),.clk(gclk));
	jxor g19211(.dina(w_n18845_0[0]),.dinb(w_n791_12[2]),.dout(n19511),.clk(gclk));
	jand g19212(.dina(n19511),.dinb(w_asqrt4_13[2]),.dout(n19512),.clk(gclk));
	jxor g19213(.dina(n19512),.dinb(w_n18855_0[0]),.dout(n19513),.clk(gclk));
	jnot g19214(.din(n19513),.dout(n19514),.clk(gclk));
	jor g19215(.dina(w_n19509_0[0]),.dinb(w_asqrt55_10[0]),.dout(n19515),.clk(gclk));
	jand g19216(.dina(w_n19515_0[1]),.dinb(w_n19514_0[1]),.dout(n19516),.clk(gclk));
	jor g19217(.dina(w_n19516_0[2]),.dinb(w_n19510_0[2]),.dout(n19517),.clk(gclk));
	jand g19218(.dina(n19517),.dinb(w_asqrt56_11[1]),.dout(n19518),.clk(gclk));
	jnot g19219(.din(w_n18860_0[0]),.dout(n19519),.clk(gclk));
	jand g19220(.dina(n19519),.dinb(w_n18858_0[0]),.dout(n19520),.clk(gclk));
	jand g19221(.dina(n19520),.dinb(w_asqrt4_13[1]),.dout(n19521),.clk(gclk));
	jxor g19222(.dina(n19521),.dinb(w_n18868_0[0]),.dout(n19522),.clk(gclk));
	jnot g19223(.din(n19522),.dout(n19523),.clk(gclk));
	jor g19224(.dina(w_n19510_0[1]),.dinb(w_asqrt56_11[0]),.dout(n19524),.clk(gclk));
	jor g19225(.dina(n19524),.dinb(w_n19516_0[1]),.dout(n19525),.clk(gclk));
	jand g19226(.dina(w_n19525_0[1]),.dinb(w_n19523_0[1]),.dout(n19526),.clk(gclk));
	jor g19227(.dina(w_n19526_0[1]),.dinb(w_n19518_0[1]),.dout(n19527),.clk(gclk));
	jand g19228(.dina(w_n19527_0[2]),.dinb(w_asqrt57_10[2]),.dout(n19528),.clk(gclk));
	jor g19229(.dina(w_n19527_0[1]),.dinb(w_asqrt57_10[1]),.dout(n19529),.clk(gclk));
	jnot g19230(.din(w_n18874_0[0]),.dout(n19530),.clk(gclk));
	jnot g19231(.din(w_n18875_0[0]),.dout(n19531),.clk(gclk));
	jand g19232(.dina(w_asqrt4_13[0]),.dinb(w_n18871_0[0]),.dout(n19532),.clk(gclk));
	jand g19233(.dina(w_n19532_0[1]),.dinb(n19531),.dout(n19533),.clk(gclk));
	jor g19234(.dina(n19533),.dinb(n19530),.dout(n19534),.clk(gclk));
	jnot g19235(.din(w_n18876_0[0]),.dout(n19535),.clk(gclk));
	jand g19236(.dina(w_n19532_0[0]),.dinb(n19535),.dout(n19536),.clk(gclk));
	jnot g19237(.din(n19536),.dout(n19537),.clk(gclk));
	jand g19238(.dina(n19537),.dinb(n19534),.dout(n19538),.clk(gclk));
	jand g19239(.dina(w_n19538_0[1]),.dinb(n19529),.dout(n19539),.clk(gclk));
	jor g19240(.dina(w_n19539_0[1]),.dinb(w_n19528_0[1]),.dout(n19540),.clk(gclk));
	jand g19241(.dina(n19540),.dinb(w_asqrt58_11[1]),.dout(n19541),.clk(gclk));
	jnot g19242(.din(w_n18880_0[0]),.dout(n19542),.clk(gclk));
	jand g19243(.dina(n19542),.dinb(w_n18878_0[0]),.dout(n19543),.clk(gclk));
	jand g19244(.dina(n19543),.dinb(w_asqrt4_12[2]),.dout(n19544),.clk(gclk));
	jxor g19245(.dina(n19544),.dinb(w_n18888_0[0]),.dout(n19545),.clk(gclk));
	jnot g19246(.din(n19545),.dout(n19546),.clk(gclk));
	jor g19247(.dina(w_n19528_0[0]),.dinb(w_asqrt58_11[0]),.dout(n19547),.clk(gclk));
	jor g19248(.dina(n19547),.dinb(w_n19539_0[0]),.dout(n19548),.clk(gclk));
	jand g19249(.dina(w_n19548_0[1]),.dinb(w_n19546_0[1]),.dout(n19549),.clk(gclk));
	jor g19250(.dina(w_n19549_0[1]),.dinb(w_n19541_0[1]),.dout(n19550),.clk(gclk));
	jand g19251(.dina(w_n19550_0[2]),.dinb(w_asqrt59_11[0]),.dout(n19551),.clk(gclk));
	jor g19252(.dina(w_n19550_0[1]),.dinb(w_asqrt59_10[2]),.dout(n19552),.clk(gclk));
	jand g19253(.dina(n19552),.dinb(w_n18958_0[0]),.dout(n19553),.clk(gclk));
	jor g19254(.dina(w_n19553_0[1]),.dinb(w_n19551_0[1]),.dout(n19554),.clk(gclk));
	jand g19255(.dina(n19554),.dinb(w_asqrt60_11[0]),.dout(n19555),.clk(gclk));
	jor g19256(.dina(w_n19551_0[0]),.dinb(w_asqrt60_10[2]),.dout(n19556),.clk(gclk));
	jor g19257(.dina(n19556),.dinb(w_n19553_0[0]),.dout(n19557),.clk(gclk));
	jnot g19258(.din(w_n18900_0[0]),.dout(n19558),.clk(gclk));
	jnot g19259(.din(w_n18902_0[0]),.dout(n19559),.clk(gclk));
	jand g19260(.dina(w_asqrt4_12[1]),.dinb(w_n18896_0[0]),.dout(n19560),.clk(gclk));
	jand g19261(.dina(w_n19560_0[1]),.dinb(n19559),.dout(n19561),.clk(gclk));
	jor g19262(.dina(n19561),.dinb(n19558),.dout(n19562),.clk(gclk));
	jnot g19263(.din(w_n18903_0[0]),.dout(n19563),.clk(gclk));
	jand g19264(.dina(w_n19560_0[0]),.dinb(n19563),.dout(n19564),.clk(gclk));
	jnot g19265(.din(n19564),.dout(n19565),.clk(gclk));
	jand g19266(.dina(n19565),.dinb(n19562),.dout(n19566),.clk(gclk));
	jand g19267(.dina(w_n19566_0[1]),.dinb(w_n19557_0[1]),.dout(n19567),.clk(gclk));
	jor g19268(.dina(n19567),.dinb(w_n19555_0[1]),.dout(n19568),.clk(gclk));
	jand g19269(.dina(w_n19568_0[2]),.dinb(w_asqrt61_11[1]),.dout(n19569),.clk(gclk));
	jor g19270(.dina(w_n19568_0[1]),.dinb(w_asqrt61_11[0]),.dout(n19570),.clk(gclk));
	jnot g19271(.din(w_n18908_0[0]),.dout(n19571),.clk(gclk));
	jnot g19272(.din(w_n18909_0[0]),.dout(n19572),.clk(gclk));
	jand g19273(.dina(w_asqrt4_12[0]),.dinb(w_n18905_0[0]),.dout(n19573),.clk(gclk));
	jand g19274(.dina(w_n19573_0[1]),.dinb(n19572),.dout(n19574),.clk(gclk));
	jor g19275(.dina(n19574),.dinb(n19571),.dout(n19575),.clk(gclk));
	jnot g19276(.din(w_n18910_0[0]),.dout(n19576),.clk(gclk));
	jand g19277(.dina(w_n19573_0[0]),.dinb(n19576),.dout(n19577),.clk(gclk));
	jnot g19278(.din(n19577),.dout(n19578),.clk(gclk));
	jand g19279(.dina(n19578),.dinb(n19575),.dout(n19579),.clk(gclk));
	jand g19280(.dina(w_n19579_0[1]),.dinb(n19570),.dout(n19580),.clk(gclk));
	jor g19281(.dina(w_n19580_0[1]),.dinb(w_n19569_0[1]),.dout(n19581),.clk(gclk));
	jand g19282(.dina(n19581),.dinb(w_asqrt62_11[1]),.dout(n19582),.clk(gclk));
	jor g19283(.dina(w_n19569_0[0]),.dinb(w_asqrt62_11[0]),.dout(n19583),.clk(gclk));
	jor g19284(.dina(n19583),.dinb(w_n19580_0[0]),.dout(n19584),.clk(gclk));
	jnot g19285(.din(w_n18916_0[0]),.dout(n19585),.clk(gclk));
	jnot g19286(.din(w_n18918_0[0]),.dout(n19586),.clk(gclk));
	jand g19287(.dina(w_asqrt4_11[2]),.dinb(w_n18912_0[0]),.dout(n19587),.clk(gclk));
	jand g19288(.dina(w_n19587_0[1]),.dinb(n19586),.dout(n19588),.clk(gclk));
	jor g19289(.dina(n19588),.dinb(n19585),.dout(n19589),.clk(gclk));
	jnot g19290(.din(w_n18919_0[0]),.dout(n19590),.clk(gclk));
	jand g19291(.dina(w_n19587_0[0]),.dinb(n19590),.dout(n19591),.clk(gclk));
	jnot g19292(.din(n19591),.dout(n19592),.clk(gclk));
	jand g19293(.dina(n19592),.dinb(n19589),.dout(n19593),.clk(gclk));
	jand g19294(.dina(w_n19593_0[1]),.dinb(w_n19584_0[1]),.dout(n19594),.clk(gclk));
	jor g19295(.dina(n19594),.dinb(w_n19582_0[1]),.dout(n19595),.clk(gclk));
	jxor g19296(.dina(w_n18920_0[0]),.dinb(w_n199_16[2]),.dout(n19596),.clk(gclk));
	jand g19297(.dina(n19596),.dinb(w_asqrt4_11[1]),.dout(n19597),.clk(gclk));
	jxor g19298(.dina(n19597),.dinb(w_n18930_0[0]),.dout(n19598),.clk(gclk));
	jnot g19299(.din(w_n18932_0[0]),.dout(n19599),.clk(gclk));
	jand g19300(.dina(w_asqrt4_11[0]),.dinb(w_n18939_0[1]),.dout(n19600),.clk(gclk));
	jand g19301(.dina(w_n19600_0[1]),.dinb(w_n19599_0[2]),.dout(n19601),.clk(gclk));
	jor g19302(.dina(n19601),.dinb(w_n18948_0[0]),.dout(n19602),.clk(gclk));
	jor g19303(.dina(n19602),.dinb(w_n19598_0[1]),.dout(n19603),.clk(gclk));
	jnot g19304(.din(n19603),.dout(n19604),.clk(gclk));
	jand g19305(.dina(n19604),.dinb(w_n19595_1[2]),.dout(n19605),.clk(gclk));
	jor g19306(.dina(n19605),.dinb(w_asqrt63_6[1]),.dout(n19606),.clk(gclk));
	jnot g19307(.din(w_n19598_0[0]),.dout(n19607),.clk(gclk));
	jor g19308(.dina(w_n19607_0[2]),.dinb(w_n19595_1[1]),.dout(n19608),.clk(gclk));
	jor g19309(.dina(w_n19600_0[0]),.dinb(w_n19599_0[1]),.dout(n19609),.clk(gclk));
	jand g19310(.dina(w_n18939_0[0]),.dinb(w_n19599_0[0]),.dout(n19610),.clk(gclk));
	jor g19311(.dina(n19610),.dinb(w_n194_15[2]),.dout(n19611),.clk(gclk));
	jnot g19312(.din(n19611),.dout(n19612),.clk(gclk));
	jand g19313(.dina(n19612),.dinb(n19609),.dout(n19613),.clk(gclk));
	jnot g19314(.din(n19613),.dout(n19614),.clk(gclk));
	jand g19315(.dina(n19614),.dinb(w_n19608_0[1]),.dout(n19615),.clk(gclk));
	jand g19316(.dina(n19615),.dinb(n19606),.dout(n19616),.clk(gclk));
	jxor g19317(.dina(w_n19550_0[0]),.dinb(w_n305_14[2]),.dout(n19617),.clk(gclk));
	jor g19318(.dina(n19617),.dinb(w_n19616_18[2]),.dout(n19618),.clk(gclk));
	jxor g19319(.dina(n19618),.dinb(n18959),.dout(n19619),.clk(gclk));
	jnot g19320(.din(n19619),.dout(n19620),.clk(gclk));
	jor g19321(.dina(w_n19616_18[1]),.dinb(w_n18961_1[0]),.dout(n19621),.clk(gclk));
	jnot g19322(.din(w_a4_0[1]),.dout(n19622),.clk(gclk));
	jnot g19323(.din(a[5]),.dout(n19623),.clk(gclk));
	jand g19324(.dina(w_n18961_0[2]),.dinb(w_n19623_0[2]),.dout(n19624),.clk(gclk));
	jand g19325(.dina(n19624),.dinb(w_n19622_1[1]),.dout(n19625),.clk(gclk));
	jnot g19326(.din(n19625),.dout(n19626),.clk(gclk));
	jand g19327(.dina(n19626),.dinb(n19621),.dout(n19627),.clk(gclk));
	jor g19328(.dina(w_n19627_0[2]),.dinb(w_n18976_2[1]),.dout(n19628),.clk(gclk));
	jor g19329(.dina(w_n19616_18[0]),.dinb(w_a6_0[0]),.dout(n19629),.clk(gclk));
	jxor g19330(.dina(w_n19629_0[1]),.dinb(w_n18962_0[0]),.dout(n19630),.clk(gclk));
	jand g19331(.dina(w_n19627_0[1]),.dinb(w_n18976_2[0]),.dout(n19631),.clk(gclk));
	jor g19332(.dina(n19631),.dinb(w_n19630_0[1]),.dout(n19632),.clk(gclk));
	jand g19333(.dina(w_n19632_0[1]),.dinb(w_n19628_0[1]),.dout(n19633),.clk(gclk));
	jor g19334(.dina(n19633),.dinb(w_n18356_8[0]),.dout(n19634),.clk(gclk));
	jand g19335(.dina(w_n19628_0[0]),.dinb(w_n18356_7[2]),.dout(n19635),.clk(gclk));
	jand g19336(.dina(n19635),.dinb(w_n19632_0[0]),.dout(n19636),.clk(gclk));
	jor g19337(.dina(w_n19629_0[0]),.dinb(w_a7_0[0]),.dout(n19637),.clk(gclk));
	jnot g19338(.din(w_n19616_17[2]),.dout(asqrt_fa_4),.clk(gclk));
	jor g19339(.dina(w_asqrt3_14[1]),.dinb(w_n18976_1[2]),.dout(n19639),.clk(gclk));
	jand g19340(.dina(n19639),.dinb(n19637),.dout(n19640),.clk(gclk));
	jxor g19341(.dina(n19640),.dinb(w_n18362_0[1]),.dout(n19641),.clk(gclk));
	jor g19342(.dina(w_n19641_0[1]),.dinb(w_n19636_0[1]),.dout(n19642),.clk(gclk));
	jand g19343(.dina(n19642),.dinb(w_n19634_0[1]),.dout(n19643),.clk(gclk));
	jor g19344(.dina(w_n19643_0[2]),.dinb(w_n18360_2[1]),.dout(n19644),.clk(gclk));
	jand g19345(.dina(w_n19643_0[1]),.dinb(w_n18360_2[0]),.dout(n19645),.clk(gclk));
	jxor g19346(.dina(w_n18965_0[0]),.dinb(w_n18356_7[1]),.dout(n19646),.clk(gclk));
	jor g19347(.dina(n19646),.dinb(w_n19616_17[1]),.dout(n19647),.clk(gclk));
	jxor g19348(.dina(n19647),.dinb(w_n18968_0[0]),.dout(n19648),.clk(gclk));
	jor g19349(.dina(w_n19648_0[1]),.dinb(n19645),.dout(n19649),.clk(gclk));
	jand g19350(.dina(w_n19649_0[1]),.dinb(w_n19644_0[1]),.dout(n19650),.clk(gclk));
	jor g19351(.dina(n19650),.dinb(w_n17140_8[1]),.dout(n19651),.clk(gclk));
	jnot g19352(.din(w_n18974_0[0]),.dout(n19652),.clk(gclk));
	jor g19353(.dina(n19652),.dinb(w_n18972_0[0]),.dout(n19653),.clk(gclk));
	jor g19354(.dina(n19653),.dinb(w_n19616_17[0]),.dout(n19654),.clk(gclk));
	jxor g19355(.dina(n19654),.dinb(w_n18979_0[0]),.dout(n19655),.clk(gclk));
	jand g19356(.dina(w_n19644_0[0]),.dinb(w_n17140_8[0]),.dout(n19656),.clk(gclk));
	jand g19357(.dina(n19656),.dinb(w_n19649_0[0]),.dout(n19657),.clk(gclk));
	jor g19358(.dina(w_n19657_0[1]),.dinb(w_n19655_0[1]),.dout(n19658),.clk(gclk));
	jand g19359(.dina(w_n19658_0[1]),.dinb(w_n19651_0[1]),.dout(n19659),.clk(gclk));
	jor g19360(.dina(w_n19659_0[2]),.dinb(w_n17135_3[0]),.dout(n19660),.clk(gclk));
	jand g19361(.dina(w_n19659_0[1]),.dinb(w_n17135_2[2]),.dout(n19661),.clk(gclk));
	jxor g19362(.dina(w_n18981_0[0]),.dinb(w_n17140_7[2]),.dout(n19662),.clk(gclk));
	jor g19363(.dina(n19662),.dinb(w_n19616_16[2]),.dout(n19663),.clk(gclk));
	jxor g19364(.dina(n19663),.dinb(w_n18986_0[0]),.dout(n19664),.clk(gclk));
	jnot g19365(.din(w_n19664_0[1]),.dout(n19665),.clk(gclk));
	jor g19366(.dina(n19665),.dinb(n19661),.dout(n19666),.clk(gclk));
	jand g19367(.dina(w_n19666_0[1]),.dinb(w_n19660_0[1]),.dout(n19667),.clk(gclk));
	jor g19368(.dina(n19667),.dinb(w_n15955_8[2]),.dout(n19668),.clk(gclk));
	jand g19369(.dina(w_n19660_0[0]),.dinb(w_n15955_8[1]),.dout(n19669),.clk(gclk));
	jand g19370(.dina(n19669),.dinb(w_n19666_0[0]),.dout(n19670),.clk(gclk));
	jnot g19371(.din(w_n18990_0[0]),.dout(n19671),.clk(gclk));
	jand g19372(.dina(w_asqrt3_14[0]),.dinb(n19671),.dout(n19672),.clk(gclk));
	jand g19373(.dina(w_n19672_0[1]),.dinb(w_n18997_0[0]),.dout(n19673),.clk(gclk));
	jor g19374(.dina(n19673),.dinb(w_n18995_0[0]),.dout(n19674),.clk(gclk));
	jand g19375(.dina(w_n19672_0[0]),.dinb(w_n18998_0[0]),.dout(n19675),.clk(gclk));
	jnot g19376(.din(n19675),.dout(n19676),.clk(gclk));
	jand g19377(.dina(n19676),.dinb(n19674),.dout(n19677),.clk(gclk));
	jnot g19378(.din(n19677),.dout(n19678),.clk(gclk));
	jor g19379(.dina(w_n19678_0[1]),.dinb(w_n19670_0[1]),.dout(n19679),.clk(gclk));
	jand g19380(.dina(n19679),.dinb(w_n19668_0[1]),.dout(n19680),.clk(gclk));
	jor g19381(.dina(w_n19680_0[2]),.dinb(w_n15950_3[1]),.dout(n19681),.clk(gclk));
	jand g19382(.dina(w_n19680_0[1]),.dinb(w_n15950_3[0]),.dout(n19682),.clk(gclk));
	jnot g19383(.din(w_n19005_0[0]),.dout(n19683),.clk(gclk));
	jxor g19384(.dina(w_n18999_0[0]),.dinb(w_n15955_8[0]),.dout(n19684),.clk(gclk));
	jor g19385(.dina(n19684),.dinb(w_n19616_16[1]),.dout(n19685),.clk(gclk));
	jxor g19386(.dina(n19685),.dinb(n19683),.dout(n19686),.clk(gclk));
	jnot g19387(.din(w_n19686_0[1]),.dout(n19687),.clk(gclk));
	jor g19388(.dina(n19687),.dinb(n19682),.dout(n19688),.clk(gclk));
	jand g19389(.dina(w_n19688_0[1]),.dinb(w_n19681_0[1]),.dout(n19689),.clk(gclk));
	jor g19390(.dina(n19689),.dinb(w_n14821_9[0]),.dout(n19690),.clk(gclk));
	jnot g19391(.din(w_n19010_0[0]),.dout(n19691),.clk(gclk));
	jor g19392(.dina(n19691),.dinb(w_n19008_0[0]),.dout(n19692),.clk(gclk));
	jor g19393(.dina(n19692),.dinb(w_n19616_16[0]),.dout(n19693),.clk(gclk));
	jxor g19394(.dina(n19693),.dinb(w_n19019_0[0]),.dout(n19694),.clk(gclk));
	jand g19395(.dina(w_n19681_0[0]),.dinb(w_n14821_8[2]),.dout(n19695),.clk(gclk));
	jand g19396(.dina(n19695),.dinb(w_n19688_0[0]),.dout(n19696),.clk(gclk));
	jor g19397(.dina(w_n19696_0[1]),.dinb(w_n19694_0[1]),.dout(n19697),.clk(gclk));
	jand g19398(.dina(w_n19697_0[1]),.dinb(w_n19690_0[1]),.dout(n19698),.clk(gclk));
	jor g19399(.dina(w_n19698_0[2]),.dinb(w_n14816_4[0]),.dout(n19699),.clk(gclk));
	jand g19400(.dina(w_n19698_0[1]),.dinb(w_n14816_3[2]),.dout(n19700),.clk(gclk));
	jnot g19401(.din(w_n19026_0[0]),.dout(n19701),.clk(gclk));
	jxor g19402(.dina(w_n19021_0[0]),.dinb(w_n14821_8[1]),.dout(n19702),.clk(gclk));
	jor g19403(.dina(n19702),.dinb(w_n19616_15[2]),.dout(n19703),.clk(gclk));
	jxor g19404(.dina(n19703),.dinb(n19701),.dout(n19704),.clk(gclk));
	jnot g19405(.din(n19704),.dout(n19705),.clk(gclk));
	jor g19406(.dina(w_n19705_0[1]),.dinb(n19700),.dout(n19706),.clk(gclk));
	jand g19407(.dina(w_n19706_0[1]),.dinb(w_n19699_0[1]),.dout(n19707),.clk(gclk));
	jor g19408(.dina(n19707),.dinb(w_n13723_8[2]),.dout(n19708),.clk(gclk));
	jand g19409(.dina(w_n19699_0[0]),.dinb(w_n13723_8[1]),.dout(n19709),.clk(gclk));
	jand g19410(.dina(n19709),.dinb(w_n19706_0[0]),.dout(n19710),.clk(gclk));
	jnot g19411(.din(w_n19029_0[0]),.dout(n19711),.clk(gclk));
	jand g19412(.dina(w_asqrt3_13[2]),.dinb(n19711),.dout(n19712),.clk(gclk));
	jand g19413(.dina(w_n19712_0[1]),.dinb(w_n19036_0[0]),.dout(n19713),.clk(gclk));
	jor g19414(.dina(n19713),.dinb(w_n19034_0[0]),.dout(n19714),.clk(gclk));
	jand g19415(.dina(w_n19712_0[0]),.dinb(w_n19037_0[0]),.dout(n19715),.clk(gclk));
	jnot g19416(.din(n19715),.dout(n19716),.clk(gclk));
	jand g19417(.dina(n19716),.dinb(n19714),.dout(n19717),.clk(gclk));
	jnot g19418(.din(n19717),.dout(n19718),.clk(gclk));
	jor g19419(.dina(w_n19718_0[1]),.dinb(w_n19710_0[1]),.dout(n19719),.clk(gclk));
	jand g19420(.dina(n19719),.dinb(w_n19708_0[1]),.dout(n19720),.clk(gclk));
	jor g19421(.dina(w_n19720_0[1]),.dinb(w_n13718_4[0]),.dout(n19721),.clk(gclk));
	jxor g19422(.dina(w_n19038_0[0]),.dinb(w_n13723_8[0]),.dout(n19722),.clk(gclk));
	jor g19423(.dina(n19722),.dinb(w_n19616_15[1]),.dout(n19723),.clk(gclk));
	jxor g19424(.dina(n19723),.dinb(w_n19043_0[0]),.dout(n19724),.clk(gclk));
	jand g19425(.dina(w_n19720_0[0]),.dinb(w_n13718_3[2]),.dout(n19725),.clk(gclk));
	jor g19426(.dina(w_n19725_0[1]),.dinb(w_n19724_0[1]),.dout(n19726),.clk(gclk));
	jand g19427(.dina(w_n19726_0[2]),.dinb(w_n19721_0[2]),.dout(n19727),.clk(gclk));
	jor g19428(.dina(n19727),.dinb(w_n12675_9[1]),.dout(n19728),.clk(gclk));
	jnot g19429(.din(w_n19048_0[0]),.dout(n19729),.clk(gclk));
	jor g19430(.dina(n19729),.dinb(w_n19046_0[0]),.dout(n19730),.clk(gclk));
	jor g19431(.dina(n19730),.dinb(w_n19616_15[0]),.dout(n19731),.clk(gclk));
	jxor g19432(.dina(n19731),.dinb(w_n19057_0[0]),.dout(n19732),.clk(gclk));
	jand g19433(.dina(w_n19721_0[1]),.dinb(w_n12675_9[0]),.dout(n19733),.clk(gclk));
	jand g19434(.dina(n19733),.dinb(w_n19726_0[1]),.dout(n19734),.clk(gclk));
	jor g19435(.dina(w_n19734_0[1]),.dinb(w_n19732_0[1]),.dout(n19735),.clk(gclk));
	jand g19436(.dina(w_n19735_0[1]),.dinb(w_n19728_0[1]),.dout(n19736),.clk(gclk));
	jor g19437(.dina(w_n19736_0[2]),.dinb(w_n12670_4[2]),.dout(n19737),.clk(gclk));
	jand g19438(.dina(w_n19736_0[1]),.dinb(w_n12670_4[1]),.dout(n19738),.clk(gclk));
	jnot g19439(.din(w_n19060_0[0]),.dout(n19739),.clk(gclk));
	jand g19440(.dina(w_asqrt3_13[1]),.dinb(n19739),.dout(n19740),.clk(gclk));
	jand g19441(.dina(w_n19740_0[1]),.dinb(w_n19065_0[0]),.dout(n19741),.clk(gclk));
	jor g19442(.dina(n19741),.dinb(w_n19064_0[0]),.dout(n19742),.clk(gclk));
	jand g19443(.dina(w_n19740_0[0]),.dinb(w_n19066_0[0]),.dout(n19743),.clk(gclk));
	jnot g19444(.din(n19743),.dout(n19744),.clk(gclk));
	jand g19445(.dina(n19744),.dinb(n19742),.dout(n19745),.clk(gclk));
	jnot g19446(.din(n19745),.dout(n19746),.clk(gclk));
	jor g19447(.dina(w_n19746_0[1]),.dinb(n19738),.dout(n19747),.clk(gclk));
	jand g19448(.dina(w_n19747_0[1]),.dinb(w_n19737_0[1]),.dout(n19748),.clk(gclk));
	jor g19449(.dina(n19748),.dinb(w_n11662_9[1]),.dout(n19749),.clk(gclk));
	jand g19450(.dina(w_n19737_0[0]),.dinb(w_n11662_9[0]),.dout(n19750),.clk(gclk));
	jand g19451(.dina(n19750),.dinb(w_n19747_0[0]),.dout(n19751),.clk(gclk));
	jnot g19452(.din(w_n19068_0[0]),.dout(n19752),.clk(gclk));
	jand g19453(.dina(w_asqrt3_13[0]),.dinb(n19752),.dout(n19753),.clk(gclk));
	jand g19454(.dina(w_n19753_0[1]),.dinb(w_n19075_0[0]),.dout(n19754),.clk(gclk));
	jor g19455(.dina(n19754),.dinb(w_n19073_0[0]),.dout(n19755),.clk(gclk));
	jand g19456(.dina(w_n19753_0[0]),.dinb(w_n19076_0[0]),.dout(n19756),.clk(gclk));
	jnot g19457(.din(n19756),.dout(n19757),.clk(gclk));
	jand g19458(.dina(n19757),.dinb(n19755),.dout(n19758),.clk(gclk));
	jnot g19459(.din(n19758),.dout(n19759),.clk(gclk));
	jor g19460(.dina(w_n19759_0[1]),.dinb(w_n19751_0[1]),.dout(n19760),.clk(gclk));
	jand g19461(.dina(n19760),.dinb(w_n19749_0[1]),.dout(n19761),.clk(gclk));
	jor g19462(.dina(w_n19761_0[1]),.dinb(w_n11657_4[2]),.dout(n19762),.clk(gclk));
	jxor g19463(.dina(w_n19077_0[0]),.dinb(w_n11662_8[2]),.dout(n19763),.clk(gclk));
	jor g19464(.dina(n19763),.dinb(w_n19616_14[2]),.dout(n19764),.clk(gclk));
	jxor g19465(.dina(n19764),.dinb(w_n19088_0[0]),.dout(n19765),.clk(gclk));
	jand g19466(.dina(w_n19761_0[0]),.dinb(w_n11657_4[1]),.dout(n19766),.clk(gclk));
	jor g19467(.dina(w_n19766_0[1]),.dinb(w_n19765_0[1]),.dout(n19767),.clk(gclk));
	jand g19468(.dina(w_n19767_0[2]),.dinb(w_n19762_0[2]),.dout(n19768),.clk(gclk));
	jor g19469(.dina(n19768),.dinb(w_n10701_9[2]),.dout(n19769),.clk(gclk));
	jnot g19470(.din(w_n19093_0[0]),.dout(n19770),.clk(gclk));
	jor g19471(.dina(n19770),.dinb(w_n19091_0[0]),.dout(n19771),.clk(gclk));
	jor g19472(.dina(n19771),.dinb(w_n19616_14[1]),.dout(n19772),.clk(gclk));
	jxor g19473(.dina(n19772),.dinb(w_n19102_0[0]),.dout(n19773),.clk(gclk));
	jand g19474(.dina(w_n19762_0[1]),.dinb(w_n10701_9[1]),.dout(n19774),.clk(gclk));
	jand g19475(.dina(n19774),.dinb(w_n19767_0[1]),.dout(n19775),.clk(gclk));
	jor g19476(.dina(w_n19775_0[1]),.dinb(w_n19773_0[1]),.dout(n19776),.clk(gclk));
	jand g19477(.dina(w_n19776_0[1]),.dinb(w_n19769_0[1]),.dout(n19777),.clk(gclk));
	jor g19478(.dina(w_n19777_0[2]),.dinb(w_n10696_5[2]),.dout(n19778),.clk(gclk));
	jand g19479(.dina(w_n19777_0[1]),.dinb(w_n10696_5[1]),.dout(n19779),.clk(gclk));
	jnot g19480(.din(w_n19105_0[0]),.dout(n19780),.clk(gclk));
	jand g19481(.dina(w_asqrt3_12[2]),.dinb(n19780),.dout(n19781),.clk(gclk));
	jand g19482(.dina(w_n19781_0[1]),.dinb(w_n19110_0[0]),.dout(n19782),.clk(gclk));
	jor g19483(.dina(n19782),.dinb(w_n19109_0[0]),.dout(n19783),.clk(gclk));
	jand g19484(.dina(w_n19781_0[0]),.dinb(w_n19111_0[0]),.dout(n19784),.clk(gclk));
	jnot g19485(.din(n19784),.dout(n19785),.clk(gclk));
	jand g19486(.dina(n19785),.dinb(n19783),.dout(n19786),.clk(gclk));
	jnot g19487(.din(n19786),.dout(n19787),.clk(gclk));
	jor g19488(.dina(w_n19787_0[1]),.dinb(n19779),.dout(n19788),.clk(gclk));
	jand g19489(.dina(w_n19788_0[1]),.dinb(w_n19778_0[1]),.dout(n19789),.clk(gclk));
	jor g19490(.dina(n19789),.dinb(w_n9774_9[2]),.dout(n19790),.clk(gclk));
	jand g19491(.dina(w_n19778_0[0]),.dinb(w_n9774_9[1]),.dout(n19791),.clk(gclk));
	jand g19492(.dina(n19791),.dinb(w_n19788_0[0]),.dout(n19792),.clk(gclk));
	jnot g19493(.din(w_n19113_0[0]),.dout(n19793),.clk(gclk));
	jand g19494(.dina(w_asqrt3_12[1]),.dinb(n19793),.dout(n19794),.clk(gclk));
	jand g19495(.dina(w_n19794_0[1]),.dinb(w_n19120_0[0]),.dout(n19795),.clk(gclk));
	jor g19496(.dina(n19795),.dinb(w_n19118_0[0]),.dout(n19796),.clk(gclk));
	jand g19497(.dina(w_n19794_0[0]),.dinb(w_n19121_0[0]),.dout(n19797),.clk(gclk));
	jnot g19498(.din(n19797),.dout(n19798),.clk(gclk));
	jand g19499(.dina(n19798),.dinb(n19796),.dout(n19799),.clk(gclk));
	jnot g19500(.din(n19799),.dout(n19800),.clk(gclk));
	jor g19501(.dina(w_n19800_0[1]),.dinb(w_n19792_0[1]),.dout(n19801),.clk(gclk));
	jand g19502(.dina(n19801),.dinb(w_n19790_0[1]),.dout(n19802),.clk(gclk));
	jor g19503(.dina(w_n19802_0[1]),.dinb(w_n9769_5[2]),.dout(n19803),.clk(gclk));
	jxor g19504(.dina(w_n19122_0[0]),.dinb(w_n9774_9[0]),.dout(n19804),.clk(gclk));
	jor g19505(.dina(n19804),.dinb(w_n19616_14[0]),.dout(n19805),.clk(gclk));
	jxor g19506(.dina(n19805),.dinb(w_n19133_0[0]),.dout(n19806),.clk(gclk));
	jand g19507(.dina(w_n19802_0[0]),.dinb(w_n9769_5[1]),.dout(n19807),.clk(gclk));
	jor g19508(.dina(w_n19807_0[1]),.dinb(w_n19806_0[1]),.dout(n19808),.clk(gclk));
	jand g19509(.dina(w_n19808_0[2]),.dinb(w_n19803_0[2]),.dout(n19809),.clk(gclk));
	jor g19510(.dina(n19809),.dinb(w_n8898_10[1]),.dout(n19810),.clk(gclk));
	jnot g19511(.din(w_n19138_0[0]),.dout(n19811),.clk(gclk));
	jor g19512(.dina(n19811),.dinb(w_n19136_0[0]),.dout(n19812),.clk(gclk));
	jor g19513(.dina(n19812),.dinb(w_n19616_13[2]),.dout(n19813),.clk(gclk));
	jxor g19514(.dina(n19813),.dinb(w_n19147_0[0]),.dout(n19814),.clk(gclk));
	jand g19515(.dina(w_n19803_0[1]),.dinb(w_n8898_10[0]),.dout(n19815),.clk(gclk));
	jand g19516(.dina(n19815),.dinb(w_n19808_0[1]),.dout(n19816),.clk(gclk));
	jor g19517(.dina(w_n19816_0[1]),.dinb(w_n19814_0[1]),.dout(n19817),.clk(gclk));
	jand g19518(.dina(w_n19817_0[1]),.dinb(w_n19810_0[1]),.dout(n19818),.clk(gclk));
	jor g19519(.dina(w_n19818_0[2]),.dinb(w_n8893_6[1]),.dout(n19819),.clk(gclk));
	jand g19520(.dina(w_n19818_0[1]),.dinb(w_n8893_6[0]),.dout(n19820),.clk(gclk));
	jnot g19521(.din(w_n19150_0[0]),.dout(n19821),.clk(gclk));
	jand g19522(.dina(w_asqrt3_12[0]),.dinb(n19821),.dout(n19822),.clk(gclk));
	jand g19523(.dina(w_n19822_0[1]),.dinb(w_n19155_0[0]),.dout(n19823),.clk(gclk));
	jor g19524(.dina(n19823),.dinb(w_n19154_0[0]),.dout(n19824),.clk(gclk));
	jand g19525(.dina(w_n19822_0[0]),.dinb(w_n19156_0[0]),.dout(n19825),.clk(gclk));
	jnot g19526(.din(n19825),.dout(n19826),.clk(gclk));
	jand g19527(.dina(n19826),.dinb(n19824),.dout(n19827),.clk(gclk));
	jnot g19528(.din(n19827),.dout(n19828),.clk(gclk));
	jor g19529(.dina(w_n19828_0[1]),.dinb(n19820),.dout(n19829),.clk(gclk));
	jand g19530(.dina(w_n19829_0[1]),.dinb(w_n19819_0[1]),.dout(n19830),.clk(gclk));
	jor g19531(.dina(n19830),.dinb(w_n8058_10[1]),.dout(n19831),.clk(gclk));
	jand g19532(.dina(w_n19819_0[0]),.dinb(w_n8058_10[0]),.dout(n19832),.clk(gclk));
	jand g19533(.dina(n19832),.dinb(w_n19829_0[0]),.dout(n19833),.clk(gclk));
	jnot g19534(.din(w_n19158_0[0]),.dout(n19834),.clk(gclk));
	jand g19535(.dina(w_asqrt3_11[2]),.dinb(n19834),.dout(n19835),.clk(gclk));
	jand g19536(.dina(w_n19835_0[1]),.dinb(w_n19165_0[0]),.dout(n19836),.clk(gclk));
	jor g19537(.dina(n19836),.dinb(w_n19163_0[0]),.dout(n19837),.clk(gclk));
	jand g19538(.dina(w_n19835_0[0]),.dinb(w_n19166_0[0]),.dout(n19838),.clk(gclk));
	jnot g19539(.din(n19838),.dout(n19839),.clk(gclk));
	jand g19540(.dina(n19839),.dinb(n19837),.dout(n19840),.clk(gclk));
	jnot g19541(.din(n19840),.dout(n19841),.clk(gclk));
	jor g19542(.dina(w_n19841_0[1]),.dinb(w_n19833_0[1]),.dout(n19842),.clk(gclk));
	jand g19543(.dina(n19842),.dinb(w_n19831_0[1]),.dout(n19843),.clk(gclk));
	jor g19544(.dina(w_n19843_0[1]),.dinb(w_n8053_6[1]),.dout(n19844),.clk(gclk));
	jxor g19545(.dina(w_n19167_0[0]),.dinb(w_n8058_9[2]),.dout(n19845),.clk(gclk));
	jor g19546(.dina(n19845),.dinb(w_n19616_13[1]),.dout(n19846),.clk(gclk));
	jxor g19547(.dina(n19846),.dinb(w_n19178_0[0]),.dout(n19847),.clk(gclk));
	jand g19548(.dina(w_n19843_0[0]),.dinb(w_n8053_6[0]),.dout(n19848),.clk(gclk));
	jor g19549(.dina(w_n19848_0[1]),.dinb(w_n19847_0[1]),.dout(n19849),.clk(gclk));
	jand g19550(.dina(w_n19849_0[2]),.dinb(w_n19844_0[2]),.dout(n19850),.clk(gclk));
	jor g19551(.dina(n19850),.dinb(w_n7265_10[2]),.dout(n19851),.clk(gclk));
	jnot g19552(.din(w_n19183_0[0]),.dout(n19852),.clk(gclk));
	jor g19553(.dina(n19852),.dinb(w_n19181_0[0]),.dout(n19853),.clk(gclk));
	jor g19554(.dina(n19853),.dinb(w_n19616_13[0]),.dout(n19854),.clk(gclk));
	jxor g19555(.dina(n19854),.dinb(w_n19192_0[0]),.dout(n19855),.clk(gclk));
	jand g19556(.dina(w_n19844_0[1]),.dinb(w_n7265_10[1]),.dout(n19856),.clk(gclk));
	jand g19557(.dina(n19856),.dinb(w_n19849_0[1]),.dout(n19857),.clk(gclk));
	jor g19558(.dina(w_n19857_0[1]),.dinb(w_n19855_0[1]),.dout(n19858),.clk(gclk));
	jand g19559(.dina(w_n19858_0[1]),.dinb(w_n19851_0[1]),.dout(n19859),.clk(gclk));
	jor g19560(.dina(w_n19859_0[2]),.dinb(w_n7260_7[1]),.dout(n19860),.clk(gclk));
	jand g19561(.dina(w_n19859_0[1]),.dinb(w_n7260_7[0]),.dout(n19861),.clk(gclk));
	jnot g19562(.din(w_n19195_0[0]),.dout(n19862),.clk(gclk));
	jand g19563(.dina(w_asqrt3_11[1]),.dinb(n19862),.dout(n19863),.clk(gclk));
	jand g19564(.dina(w_n19863_0[1]),.dinb(w_n19200_0[0]),.dout(n19864),.clk(gclk));
	jor g19565(.dina(n19864),.dinb(w_n19199_0[0]),.dout(n19865),.clk(gclk));
	jand g19566(.dina(w_n19863_0[0]),.dinb(w_n19201_0[0]),.dout(n19866),.clk(gclk));
	jnot g19567(.din(n19866),.dout(n19867),.clk(gclk));
	jand g19568(.dina(n19867),.dinb(n19865),.dout(n19868),.clk(gclk));
	jnot g19569(.din(n19868),.dout(n19869),.clk(gclk));
	jor g19570(.dina(w_n19869_0[1]),.dinb(n19861),.dout(n19870),.clk(gclk));
	jand g19571(.dina(w_n19870_0[1]),.dinb(w_n19860_0[1]),.dout(n19871),.clk(gclk));
	jor g19572(.dina(n19871),.dinb(w_n6505_10[2]),.dout(n19872),.clk(gclk));
	jand g19573(.dina(w_n19860_0[0]),.dinb(w_n6505_10[1]),.dout(n19873),.clk(gclk));
	jand g19574(.dina(n19873),.dinb(w_n19870_0[0]),.dout(n19874),.clk(gclk));
	jnot g19575(.din(w_n19203_0[0]),.dout(n19875),.clk(gclk));
	jand g19576(.dina(w_asqrt3_11[0]),.dinb(n19875),.dout(n19876),.clk(gclk));
	jand g19577(.dina(w_n19876_0[1]),.dinb(w_n19210_0[0]),.dout(n19877),.clk(gclk));
	jor g19578(.dina(n19877),.dinb(w_n19208_0[0]),.dout(n19878),.clk(gclk));
	jand g19579(.dina(w_n19876_0[0]),.dinb(w_n19211_0[0]),.dout(n19879),.clk(gclk));
	jnot g19580(.din(n19879),.dout(n19880),.clk(gclk));
	jand g19581(.dina(n19880),.dinb(n19878),.dout(n19881),.clk(gclk));
	jnot g19582(.din(n19881),.dout(n19882),.clk(gclk));
	jor g19583(.dina(w_n19882_0[1]),.dinb(w_n19874_0[1]),.dout(n19883),.clk(gclk));
	jand g19584(.dina(n19883),.dinb(w_n19872_0[1]),.dout(n19884),.clk(gclk));
	jor g19585(.dina(w_n19884_0[1]),.dinb(w_n6500_7[1]),.dout(n19885),.clk(gclk));
	jxor g19586(.dina(w_n19212_0[0]),.dinb(w_n6505_10[0]),.dout(n19886),.clk(gclk));
	jor g19587(.dina(n19886),.dinb(w_n19616_12[2]),.dout(n19887),.clk(gclk));
	jxor g19588(.dina(n19887),.dinb(w_n19223_0[0]),.dout(n19888),.clk(gclk));
	jand g19589(.dina(w_n19884_0[0]),.dinb(w_n6500_7[0]),.dout(n19889),.clk(gclk));
	jor g19590(.dina(w_n19889_0[1]),.dinb(w_n19888_0[1]),.dout(n19890),.clk(gclk));
	jand g19591(.dina(w_n19890_0[2]),.dinb(w_n19885_0[2]),.dout(n19891),.clk(gclk));
	jor g19592(.dina(n19891),.dinb(w_n5793_11[0]),.dout(n19892),.clk(gclk));
	jnot g19593(.din(w_n19228_0[0]),.dout(n19893),.clk(gclk));
	jor g19594(.dina(n19893),.dinb(w_n19226_0[0]),.dout(n19894),.clk(gclk));
	jor g19595(.dina(n19894),.dinb(w_n19616_12[1]),.dout(n19895),.clk(gclk));
	jxor g19596(.dina(n19895),.dinb(w_n19237_0[0]),.dout(n19896),.clk(gclk));
	jand g19597(.dina(w_n19885_0[1]),.dinb(w_n5793_10[2]),.dout(n19897),.clk(gclk));
	jand g19598(.dina(n19897),.dinb(w_n19890_0[1]),.dout(n19898),.clk(gclk));
	jor g19599(.dina(w_n19898_0[1]),.dinb(w_n19896_0[1]),.dout(n19899),.clk(gclk));
	jand g19600(.dina(w_n19899_0[1]),.dinb(w_n19892_0[1]),.dout(n19900),.clk(gclk));
	jor g19601(.dina(w_n19900_0[2]),.dinb(w_n5788_8[0]),.dout(n19901),.clk(gclk));
	jand g19602(.dina(w_n19900_0[1]),.dinb(w_n5788_7[2]),.dout(n19902),.clk(gclk));
	jnot g19603(.din(w_n19240_0[0]),.dout(n19903),.clk(gclk));
	jand g19604(.dina(w_asqrt3_10[2]),.dinb(n19903),.dout(n19904),.clk(gclk));
	jand g19605(.dina(w_n19904_0[1]),.dinb(w_n19245_0[0]),.dout(n19905),.clk(gclk));
	jor g19606(.dina(n19905),.dinb(w_n19244_0[0]),.dout(n19906),.clk(gclk));
	jand g19607(.dina(w_n19904_0[0]),.dinb(w_n19246_0[0]),.dout(n19907),.clk(gclk));
	jnot g19608(.din(n19907),.dout(n19908),.clk(gclk));
	jand g19609(.dina(n19908),.dinb(n19906),.dout(n19909),.clk(gclk));
	jnot g19610(.din(n19909),.dout(n19910),.clk(gclk));
	jor g19611(.dina(w_n19910_0[1]),.dinb(n19902),.dout(n19911),.clk(gclk));
	jand g19612(.dina(w_n19911_0[1]),.dinb(w_n19901_0[1]),.dout(n19912),.clk(gclk));
	jor g19613(.dina(n19912),.dinb(w_n5121_11[0]),.dout(n19913),.clk(gclk));
	jand g19614(.dina(w_n19901_0[0]),.dinb(w_n5121_10[2]),.dout(n19914),.clk(gclk));
	jand g19615(.dina(n19914),.dinb(w_n19911_0[0]),.dout(n19915),.clk(gclk));
	jnot g19616(.din(w_n19248_0[0]),.dout(n19916),.clk(gclk));
	jand g19617(.dina(w_asqrt3_10[1]),.dinb(n19916),.dout(n19917),.clk(gclk));
	jand g19618(.dina(w_n19917_0[1]),.dinb(w_n19255_0[0]),.dout(n19918),.clk(gclk));
	jor g19619(.dina(n19918),.dinb(w_n19253_0[0]),.dout(n19919),.clk(gclk));
	jand g19620(.dina(w_n19917_0[0]),.dinb(w_n19256_0[0]),.dout(n19920),.clk(gclk));
	jnot g19621(.din(n19920),.dout(n19921),.clk(gclk));
	jand g19622(.dina(n19921),.dinb(n19919),.dout(n19922),.clk(gclk));
	jnot g19623(.din(n19922),.dout(n19923),.clk(gclk));
	jor g19624(.dina(w_n19923_0[1]),.dinb(w_n19915_0[1]),.dout(n19924),.clk(gclk));
	jand g19625(.dina(n19924),.dinb(w_n19913_0[1]),.dout(n19925),.clk(gclk));
	jor g19626(.dina(w_n19925_0[1]),.dinb(w_n5116_8[0]),.dout(n19926),.clk(gclk));
	jxor g19627(.dina(w_n19257_0[0]),.dinb(w_n5121_10[1]),.dout(n19927),.clk(gclk));
	jor g19628(.dina(n19927),.dinb(w_n19616_12[0]),.dout(n19928),.clk(gclk));
	jxor g19629(.dina(n19928),.dinb(w_n19268_0[0]),.dout(n19929),.clk(gclk));
	jand g19630(.dina(w_n19925_0[0]),.dinb(w_n5116_7[2]),.dout(n19930),.clk(gclk));
	jor g19631(.dina(w_n19930_0[1]),.dinb(w_n19929_0[1]),.dout(n19931),.clk(gclk));
	jand g19632(.dina(w_n19931_0[2]),.dinb(w_n19926_0[2]),.dout(n19932),.clk(gclk));
	jor g19633(.dina(n19932),.dinb(w_n4499_11[2]),.dout(n19933),.clk(gclk));
	jnot g19634(.din(w_n19273_0[0]),.dout(n19934),.clk(gclk));
	jor g19635(.dina(n19934),.dinb(w_n19271_0[0]),.dout(n19935),.clk(gclk));
	jor g19636(.dina(n19935),.dinb(w_n19616_11[2]),.dout(n19936),.clk(gclk));
	jxor g19637(.dina(n19936),.dinb(w_n19282_0[0]),.dout(n19937),.clk(gclk));
	jand g19638(.dina(w_n19926_0[1]),.dinb(w_n4499_11[1]),.dout(n19938),.clk(gclk));
	jand g19639(.dina(n19938),.dinb(w_n19931_0[1]),.dout(n19939),.clk(gclk));
	jor g19640(.dina(w_n19939_0[1]),.dinb(w_n19937_0[1]),.dout(n19940),.clk(gclk));
	jand g19641(.dina(w_n19940_0[1]),.dinb(w_n19933_0[1]),.dout(n19941),.clk(gclk));
	jor g19642(.dina(w_n19941_0[2]),.dinb(w_n4494_9[0]),.dout(n19942),.clk(gclk));
	jand g19643(.dina(w_n19941_0[1]),.dinb(w_n4494_8[2]),.dout(n19943),.clk(gclk));
	jnot g19644(.din(w_n19285_0[0]),.dout(n19944),.clk(gclk));
	jand g19645(.dina(w_asqrt3_10[0]),.dinb(n19944),.dout(n19945),.clk(gclk));
	jand g19646(.dina(w_n19945_0[1]),.dinb(w_n19290_0[0]),.dout(n19946),.clk(gclk));
	jor g19647(.dina(n19946),.dinb(w_n19289_0[0]),.dout(n19947),.clk(gclk));
	jand g19648(.dina(w_n19945_0[0]),.dinb(w_n19291_0[0]),.dout(n19948),.clk(gclk));
	jnot g19649(.din(n19948),.dout(n19949),.clk(gclk));
	jand g19650(.dina(n19949),.dinb(n19947),.dout(n19950),.clk(gclk));
	jnot g19651(.din(n19950),.dout(n19951),.clk(gclk));
	jor g19652(.dina(w_n19951_0[1]),.dinb(n19943),.dout(n19952),.clk(gclk));
	jand g19653(.dina(w_n19952_0[1]),.dinb(w_n19942_0[1]),.dout(n19953),.clk(gclk));
	jor g19654(.dina(n19953),.dinb(w_n3912_11[2]),.dout(n19954),.clk(gclk));
	jand g19655(.dina(w_n19942_0[0]),.dinb(w_n3912_11[1]),.dout(n19955),.clk(gclk));
	jand g19656(.dina(n19955),.dinb(w_n19952_0[0]),.dout(n19956),.clk(gclk));
	jnot g19657(.din(w_n19293_0[0]),.dout(n19957),.clk(gclk));
	jand g19658(.dina(w_asqrt3_9[2]),.dinb(n19957),.dout(n19958),.clk(gclk));
	jand g19659(.dina(w_n19958_0[1]),.dinb(w_n19300_0[0]),.dout(n19959),.clk(gclk));
	jor g19660(.dina(n19959),.dinb(w_n19298_0[0]),.dout(n19960),.clk(gclk));
	jand g19661(.dina(w_n19958_0[0]),.dinb(w_n19301_0[0]),.dout(n19961),.clk(gclk));
	jnot g19662(.din(n19961),.dout(n19962),.clk(gclk));
	jand g19663(.dina(n19962),.dinb(n19960),.dout(n19963),.clk(gclk));
	jnot g19664(.din(n19963),.dout(n19964),.clk(gclk));
	jor g19665(.dina(w_n19964_0[1]),.dinb(w_n19956_0[1]),.dout(n19965),.clk(gclk));
	jand g19666(.dina(n19965),.dinb(w_n19954_0[1]),.dout(n19966),.clk(gclk));
	jor g19667(.dina(w_n19966_0[1]),.dinb(w_n3907_9[0]),.dout(n19967),.clk(gclk));
	jxor g19668(.dina(w_n19302_0[0]),.dinb(w_n3912_11[0]),.dout(n19968),.clk(gclk));
	jor g19669(.dina(n19968),.dinb(w_n19616_11[1]),.dout(n19969),.clk(gclk));
	jxor g19670(.dina(n19969),.dinb(w_n19313_0[0]),.dout(n19970),.clk(gclk));
	jand g19671(.dina(w_n19966_0[0]),.dinb(w_n3907_8[2]),.dout(n19971),.clk(gclk));
	jor g19672(.dina(w_n19971_0[1]),.dinb(w_n19970_0[1]),.dout(n19972),.clk(gclk));
	jand g19673(.dina(w_n19972_0[2]),.dinb(w_n19967_0[2]),.dout(n19973),.clk(gclk));
	jor g19674(.dina(n19973),.dinb(w_n3376_12[1]),.dout(n19974),.clk(gclk));
	jnot g19675(.din(w_n19318_0[0]),.dout(n19975),.clk(gclk));
	jor g19676(.dina(n19975),.dinb(w_n19316_0[0]),.dout(n19976),.clk(gclk));
	jor g19677(.dina(n19976),.dinb(w_n19616_11[0]),.dout(n19977),.clk(gclk));
	jxor g19678(.dina(n19977),.dinb(w_n19327_0[0]),.dout(n19978),.clk(gclk));
	jand g19679(.dina(w_n19967_0[1]),.dinb(w_n3376_12[0]),.dout(n19979),.clk(gclk));
	jand g19680(.dina(n19979),.dinb(w_n19972_0[1]),.dout(n19980),.clk(gclk));
	jor g19681(.dina(w_n19980_0[1]),.dinb(w_n19978_0[1]),.dout(n19981),.clk(gclk));
	jand g19682(.dina(w_n19981_0[1]),.dinb(w_n19974_0[1]),.dout(n19982),.clk(gclk));
	jor g19683(.dina(w_n19982_0[2]),.dinb(w_n3371_9[2]),.dout(n19983),.clk(gclk));
	jand g19684(.dina(w_n19982_0[1]),.dinb(w_n3371_9[1]),.dout(n19984),.clk(gclk));
	jnot g19685(.din(w_n19330_0[0]),.dout(n19985),.clk(gclk));
	jand g19686(.dina(w_asqrt3_9[1]),.dinb(n19985),.dout(n19986),.clk(gclk));
	jand g19687(.dina(w_n19986_0[1]),.dinb(w_n19335_0[0]),.dout(n19987),.clk(gclk));
	jor g19688(.dina(n19987),.dinb(w_n19334_0[0]),.dout(n19988),.clk(gclk));
	jand g19689(.dina(w_n19986_0[0]),.dinb(w_n19336_0[0]),.dout(n19989),.clk(gclk));
	jnot g19690(.din(n19989),.dout(n19990),.clk(gclk));
	jand g19691(.dina(n19990),.dinb(n19988),.dout(n19991),.clk(gclk));
	jnot g19692(.din(n19991),.dout(n19992),.clk(gclk));
	jor g19693(.dina(w_n19992_0[1]),.dinb(n19984),.dout(n19993),.clk(gclk));
	jand g19694(.dina(w_n19993_0[1]),.dinb(w_n19983_0[1]),.dout(n19994),.clk(gclk));
	jor g19695(.dina(n19994),.dinb(w_n2875_12[1]),.dout(n19995),.clk(gclk));
	jand g19696(.dina(w_n19983_0[0]),.dinb(w_n2875_12[0]),.dout(n19996),.clk(gclk));
	jand g19697(.dina(n19996),.dinb(w_n19993_0[0]),.dout(n19997),.clk(gclk));
	jnot g19698(.din(w_n19338_0[0]),.dout(n19998),.clk(gclk));
	jand g19699(.dina(w_asqrt3_9[0]),.dinb(n19998),.dout(n19999),.clk(gclk));
	jand g19700(.dina(w_n19999_0[1]),.dinb(w_n19345_0[0]),.dout(n20000),.clk(gclk));
	jor g19701(.dina(n20000),.dinb(w_n19343_0[0]),.dout(n20001),.clk(gclk));
	jand g19702(.dina(w_n19999_0[0]),.dinb(w_n19346_0[0]),.dout(n20002),.clk(gclk));
	jnot g19703(.din(n20002),.dout(n20003),.clk(gclk));
	jand g19704(.dina(n20003),.dinb(n20001),.dout(n20004),.clk(gclk));
	jnot g19705(.din(n20004),.dout(n20005),.clk(gclk));
	jor g19706(.dina(w_n20005_0[1]),.dinb(w_n19997_0[1]),.dout(n20006),.clk(gclk));
	jand g19707(.dina(n20006),.dinb(w_n19995_0[1]),.dout(n20007),.clk(gclk));
	jor g19708(.dina(w_n20007_0[1]),.dinb(w_n2870_9[2]),.dout(n20008),.clk(gclk));
	jxor g19709(.dina(w_n19347_0[0]),.dinb(w_n2875_11[2]),.dout(n20009),.clk(gclk));
	jor g19710(.dina(n20009),.dinb(w_n19616_10[2]),.dout(n20010),.clk(gclk));
	jxor g19711(.dina(n20010),.dinb(w_n19358_0[0]),.dout(n20011),.clk(gclk));
	jand g19712(.dina(w_n20007_0[0]),.dinb(w_n2870_9[1]),.dout(n20012),.clk(gclk));
	jor g19713(.dina(w_n20012_0[1]),.dinb(w_n20011_0[1]),.dout(n20013),.clk(gclk));
	jand g19714(.dina(w_n20013_0[2]),.dinb(w_n20008_0[2]),.dout(n20014),.clk(gclk));
	jor g19715(.dina(n20014),.dinb(w_n2425_12[2]),.dout(n20015),.clk(gclk));
	jnot g19716(.din(w_n19363_0[0]),.dout(n20016),.clk(gclk));
	jor g19717(.dina(n20016),.dinb(w_n19361_0[0]),.dout(n20017),.clk(gclk));
	jor g19718(.dina(n20017),.dinb(w_n19616_10[1]),.dout(n20018),.clk(gclk));
	jxor g19719(.dina(n20018),.dinb(w_n19372_0[0]),.dout(n20019),.clk(gclk));
	jand g19720(.dina(w_n20008_0[1]),.dinb(w_n2425_12[1]),.dout(n20020),.clk(gclk));
	jand g19721(.dina(n20020),.dinb(w_n20013_0[1]),.dout(n20021),.clk(gclk));
	jor g19722(.dina(w_n20021_0[1]),.dinb(w_n20019_0[1]),.dout(n20022),.clk(gclk));
	jand g19723(.dina(w_n20022_0[1]),.dinb(w_n20015_0[1]),.dout(n20023),.clk(gclk));
	jor g19724(.dina(w_n20023_0[2]),.dinb(w_n2420_10[2]),.dout(n20024),.clk(gclk));
	jand g19725(.dina(w_n20023_0[1]),.dinb(w_n2420_10[1]),.dout(n20025),.clk(gclk));
	jnot g19726(.din(w_n19375_0[0]),.dout(n20026),.clk(gclk));
	jand g19727(.dina(w_asqrt3_8[2]),.dinb(n20026),.dout(n20027),.clk(gclk));
	jand g19728(.dina(w_n20027_0[1]),.dinb(w_n19380_0[0]),.dout(n20028),.clk(gclk));
	jor g19729(.dina(n20028),.dinb(w_n19379_0[0]),.dout(n20029),.clk(gclk));
	jand g19730(.dina(w_n20027_0[0]),.dinb(w_n19381_0[0]),.dout(n20030),.clk(gclk));
	jnot g19731(.din(n20030),.dout(n20031),.clk(gclk));
	jand g19732(.dina(n20031),.dinb(n20029),.dout(n20032),.clk(gclk));
	jnot g19733(.din(n20032),.dout(n20033),.clk(gclk));
	jor g19734(.dina(w_n20033_0[1]),.dinb(n20025),.dout(n20034),.clk(gclk));
	jand g19735(.dina(w_n20034_0[1]),.dinb(w_n20024_0[1]),.dout(n20035),.clk(gclk));
	jor g19736(.dina(n20035),.dinb(w_n2010_12[2]),.dout(n20036),.clk(gclk));
	jand g19737(.dina(w_n20024_0[0]),.dinb(w_n2010_12[1]),.dout(n20037),.clk(gclk));
	jand g19738(.dina(n20037),.dinb(w_n20034_0[0]),.dout(n20038),.clk(gclk));
	jnot g19739(.din(w_n19383_0[0]),.dout(n20039),.clk(gclk));
	jand g19740(.dina(w_asqrt3_8[1]),.dinb(n20039),.dout(n20040),.clk(gclk));
	jand g19741(.dina(w_n20040_0[1]),.dinb(w_n19390_0[0]),.dout(n20041),.clk(gclk));
	jor g19742(.dina(n20041),.dinb(w_n19388_0[0]),.dout(n20042),.clk(gclk));
	jand g19743(.dina(w_n20040_0[0]),.dinb(w_n19391_0[0]),.dout(n20043),.clk(gclk));
	jnot g19744(.din(n20043),.dout(n20044),.clk(gclk));
	jand g19745(.dina(n20044),.dinb(n20042),.dout(n20045),.clk(gclk));
	jnot g19746(.din(n20045),.dout(n20046),.clk(gclk));
	jor g19747(.dina(w_n20046_0[1]),.dinb(w_n20038_0[1]),.dout(n20047),.clk(gclk));
	jand g19748(.dina(n20047),.dinb(w_n20036_0[1]),.dout(n20048),.clk(gclk));
	jor g19749(.dina(w_n20048_0[1]),.dinb(w_n2005_10[2]),.dout(n20049),.clk(gclk));
	jxor g19750(.dina(w_n19392_0[0]),.dinb(w_n2010_12[0]),.dout(n20050),.clk(gclk));
	jor g19751(.dina(n20050),.dinb(w_n19616_10[0]),.dout(n20051),.clk(gclk));
	jxor g19752(.dina(n20051),.dinb(w_n19403_0[0]),.dout(n20052),.clk(gclk));
	jand g19753(.dina(w_n20048_0[0]),.dinb(w_n2005_10[1]),.dout(n20053),.clk(gclk));
	jor g19754(.dina(w_n20053_0[1]),.dinb(w_n20052_0[1]),.dout(n20054),.clk(gclk));
	jand g19755(.dina(w_n20054_0[2]),.dinb(w_n20049_0[2]),.dout(n20055),.clk(gclk));
	jor g19756(.dina(n20055),.dinb(w_n1646_13[1]),.dout(n20056),.clk(gclk));
	jnot g19757(.din(w_n19408_0[0]),.dout(n20057),.clk(gclk));
	jor g19758(.dina(n20057),.dinb(w_n19406_0[0]),.dout(n20058),.clk(gclk));
	jor g19759(.dina(n20058),.dinb(w_n19616_9[2]),.dout(n20059),.clk(gclk));
	jxor g19760(.dina(n20059),.dinb(w_n19417_0[0]),.dout(n20060),.clk(gclk));
	jand g19761(.dina(w_n20049_0[1]),.dinb(w_n1646_13[0]),.dout(n20061),.clk(gclk));
	jand g19762(.dina(n20061),.dinb(w_n20054_0[1]),.dout(n20062),.clk(gclk));
	jor g19763(.dina(w_n20062_0[1]),.dinb(w_n20060_0[1]),.dout(n20063),.clk(gclk));
	jand g19764(.dina(w_n20063_0[1]),.dinb(w_n20056_0[1]),.dout(n20064),.clk(gclk));
	jor g19765(.dina(w_n20064_0[2]),.dinb(w_n1641_11[1]),.dout(n20065),.clk(gclk));
	jand g19766(.dina(w_n20064_0[1]),.dinb(w_n1641_11[0]),.dout(n20066),.clk(gclk));
	jnot g19767(.din(w_n19420_0[0]),.dout(n20067),.clk(gclk));
	jand g19768(.dina(w_asqrt3_8[0]),.dinb(n20067),.dout(n20068),.clk(gclk));
	jand g19769(.dina(w_n20068_0[1]),.dinb(w_n19425_0[0]),.dout(n20069),.clk(gclk));
	jor g19770(.dina(n20069),.dinb(w_n19424_0[0]),.dout(n20070),.clk(gclk));
	jand g19771(.dina(w_n20068_0[0]),.dinb(w_n19426_0[0]),.dout(n20071),.clk(gclk));
	jnot g19772(.din(n20071),.dout(n20072),.clk(gclk));
	jand g19773(.dina(n20072),.dinb(n20070),.dout(n20073),.clk(gclk));
	jnot g19774(.din(n20073),.dout(n20074),.clk(gclk));
	jor g19775(.dina(w_n20074_0[1]),.dinb(n20066),.dout(n20075),.clk(gclk));
	jand g19776(.dina(w_n20075_0[1]),.dinb(w_n20065_0[1]),.dout(n20076),.clk(gclk));
	jor g19777(.dina(n20076),.dinb(w_n1317_13[1]),.dout(n20077),.clk(gclk));
	jand g19778(.dina(w_n20065_0[0]),.dinb(w_n1317_13[0]),.dout(n20078),.clk(gclk));
	jand g19779(.dina(n20078),.dinb(w_n20075_0[0]),.dout(n20079),.clk(gclk));
	jnot g19780(.din(w_n19428_0[0]),.dout(n20080),.clk(gclk));
	jand g19781(.dina(w_asqrt3_7[2]),.dinb(n20080),.dout(n20081),.clk(gclk));
	jand g19782(.dina(w_n20081_0[1]),.dinb(w_n19435_0[0]),.dout(n20082),.clk(gclk));
	jor g19783(.dina(n20082),.dinb(w_n19433_0[0]),.dout(n20083),.clk(gclk));
	jand g19784(.dina(w_n20081_0[0]),.dinb(w_n19436_0[0]),.dout(n20084),.clk(gclk));
	jnot g19785(.din(n20084),.dout(n20085),.clk(gclk));
	jand g19786(.dina(n20085),.dinb(n20083),.dout(n20086),.clk(gclk));
	jnot g19787(.din(n20086),.dout(n20087),.clk(gclk));
	jor g19788(.dina(w_n20087_0[1]),.dinb(w_n20079_0[1]),.dout(n20088),.clk(gclk));
	jand g19789(.dina(n20088),.dinb(w_n20077_0[1]),.dout(n20089),.clk(gclk));
	jor g19790(.dina(w_n20089_0[1]),.dinb(w_n1312_11[1]),.dout(n20090),.clk(gclk));
	jxor g19791(.dina(w_n19437_0[0]),.dinb(w_n1317_12[2]),.dout(n20091),.clk(gclk));
	jor g19792(.dina(n20091),.dinb(w_n19616_9[1]),.dout(n20092),.clk(gclk));
	jxor g19793(.dina(n20092),.dinb(w_n19448_0[0]),.dout(n20093),.clk(gclk));
	jand g19794(.dina(w_n20089_0[0]),.dinb(w_n1312_11[0]),.dout(n20094),.clk(gclk));
	jor g19795(.dina(w_n20094_0[1]),.dinb(w_n20093_0[1]),.dout(n20095),.clk(gclk));
	jand g19796(.dina(w_n20095_0[2]),.dinb(w_n20090_0[2]),.dout(n20096),.clk(gclk));
	jor g19797(.dina(n20096),.dinb(w_n1039_13[2]),.dout(n20097),.clk(gclk));
	jnot g19798(.din(w_n19453_0[0]),.dout(n20098),.clk(gclk));
	jor g19799(.dina(n20098),.dinb(w_n19451_0[0]),.dout(n20099),.clk(gclk));
	jor g19800(.dina(n20099),.dinb(w_n19616_9[0]),.dout(n20100),.clk(gclk));
	jxor g19801(.dina(n20100),.dinb(w_n19462_0[0]),.dout(n20101),.clk(gclk));
	jand g19802(.dina(w_n20090_0[1]),.dinb(w_n1039_13[1]),.dout(n20102),.clk(gclk));
	jand g19803(.dina(n20102),.dinb(w_n20095_0[1]),.dout(n20103),.clk(gclk));
	jor g19804(.dina(w_n20103_0[1]),.dinb(w_n20101_0[1]),.dout(n20104),.clk(gclk));
	jand g19805(.dina(w_n20104_0[1]),.dinb(w_n20097_0[1]),.dout(n20105),.clk(gclk));
	jor g19806(.dina(w_n20105_0[2]),.dinb(w_n1034_12[1]),.dout(n20106),.clk(gclk));
	jand g19807(.dina(w_n20105_0[1]),.dinb(w_n1034_12[0]),.dout(n20107),.clk(gclk));
	jnot g19808(.din(w_n19465_0[0]),.dout(n20108),.clk(gclk));
	jand g19809(.dina(w_asqrt3_7[1]),.dinb(n20108),.dout(n20109),.clk(gclk));
	jand g19810(.dina(w_n20109_0[1]),.dinb(w_n19470_0[0]),.dout(n20110),.clk(gclk));
	jor g19811(.dina(n20110),.dinb(w_n19469_0[0]),.dout(n20111),.clk(gclk));
	jand g19812(.dina(w_n20109_0[0]),.dinb(w_n19471_0[0]),.dout(n20112),.clk(gclk));
	jnot g19813(.din(n20112),.dout(n20113),.clk(gclk));
	jand g19814(.dina(n20113),.dinb(n20111),.dout(n20114),.clk(gclk));
	jnot g19815(.din(n20114),.dout(n20115),.clk(gclk));
	jor g19816(.dina(w_n20115_0[1]),.dinb(n20107),.dout(n20116),.clk(gclk));
	jand g19817(.dina(w_n20116_0[1]),.dinb(w_n20106_0[1]),.dout(n20117),.clk(gclk));
	jor g19818(.dina(n20117),.dinb(w_n796_13[2]),.dout(n20118),.clk(gclk));
	jand g19819(.dina(w_n20106_0[0]),.dinb(w_n796_13[1]),.dout(n20119),.clk(gclk));
	jand g19820(.dina(n20119),.dinb(w_n20116_0[0]),.dout(n20120),.clk(gclk));
	jnot g19821(.din(w_n19473_0[0]),.dout(n20121),.clk(gclk));
	jand g19822(.dina(w_asqrt3_7[0]),.dinb(n20121),.dout(n20122),.clk(gclk));
	jand g19823(.dina(w_n20122_0[1]),.dinb(w_n19480_0[0]),.dout(n20123),.clk(gclk));
	jor g19824(.dina(n20123),.dinb(w_n19478_0[0]),.dout(n20124),.clk(gclk));
	jand g19825(.dina(w_n20122_0[0]),.dinb(w_n19481_0[0]),.dout(n20125),.clk(gclk));
	jnot g19826(.din(n20125),.dout(n20126),.clk(gclk));
	jand g19827(.dina(n20126),.dinb(n20124),.dout(n20127),.clk(gclk));
	jnot g19828(.din(n20127),.dout(n20128),.clk(gclk));
	jor g19829(.dina(w_n20128_0[1]),.dinb(w_n20120_0[1]),.dout(n20129),.clk(gclk));
	jand g19830(.dina(n20129),.dinb(w_n20118_0[1]),.dout(n20130),.clk(gclk));
	jor g19831(.dina(w_n20130_0[1]),.dinb(w_n791_12[1]),.dout(n20131),.clk(gclk));
	jxor g19832(.dina(w_n19482_0[0]),.dinb(w_n796_13[0]),.dout(n20132),.clk(gclk));
	jor g19833(.dina(n20132),.dinb(w_n19616_8[2]),.dout(n20133),.clk(gclk));
	jxor g19834(.dina(n20133),.dinb(w_n19493_0[0]),.dout(n20134),.clk(gclk));
	jand g19835(.dina(w_n20130_0[0]),.dinb(w_n791_12[0]),.dout(n20135),.clk(gclk));
	jor g19836(.dina(w_n20135_0[1]),.dinb(w_n20134_0[1]),.dout(n20136),.clk(gclk));
	jand g19837(.dina(w_n20136_0[2]),.dinb(w_n20131_0[2]),.dout(n20137),.clk(gclk));
	jor g19838(.dina(n20137),.dinb(w_n595_14[0]),.dout(n20138),.clk(gclk));
	jnot g19839(.din(w_n19498_0[0]),.dout(n20139),.clk(gclk));
	jor g19840(.dina(n20139),.dinb(w_n19496_0[0]),.dout(n20140),.clk(gclk));
	jor g19841(.dina(n20140),.dinb(w_n19616_8[1]),.dout(n20141),.clk(gclk));
	jxor g19842(.dina(n20141),.dinb(w_n19507_0[0]),.dout(n20142),.clk(gclk));
	jand g19843(.dina(w_n20131_0[1]),.dinb(w_n595_13[2]),.dout(n20143),.clk(gclk));
	jand g19844(.dina(n20143),.dinb(w_n20136_0[1]),.dout(n20144),.clk(gclk));
	jor g19845(.dina(w_n20144_0[1]),.dinb(w_n20142_0[1]),.dout(n20145),.clk(gclk));
	jand g19846(.dina(w_n20145_0[1]),.dinb(w_n20138_0[1]),.dout(n20146),.clk(gclk));
	jor g19847(.dina(w_n20146_0[2]),.dinb(w_n590_13[0]),.dout(n20147),.clk(gclk));
	jand g19848(.dina(w_n20146_0[1]),.dinb(w_n590_12[2]),.dout(n20148),.clk(gclk));
	jnot g19849(.din(w_n19510_0[0]),.dout(n20149),.clk(gclk));
	jand g19850(.dina(w_asqrt3_6[2]),.dinb(n20149),.dout(n20150),.clk(gclk));
	jand g19851(.dina(w_n20150_0[1]),.dinb(w_n19515_0[0]),.dout(n20151),.clk(gclk));
	jor g19852(.dina(n20151),.dinb(w_n19514_0[0]),.dout(n20152),.clk(gclk));
	jand g19853(.dina(w_n20150_0[0]),.dinb(w_n19516_0[0]),.dout(n20153),.clk(gclk));
	jnot g19854(.din(n20153),.dout(n20154),.clk(gclk));
	jand g19855(.dina(n20154),.dinb(n20152),.dout(n20155),.clk(gclk));
	jnot g19856(.din(n20155),.dout(n20156),.clk(gclk));
	jor g19857(.dina(w_n20156_0[1]),.dinb(n20148),.dout(n20157),.clk(gclk));
	jand g19858(.dina(w_n20157_0[1]),.dinb(w_n20147_0[1]),.dout(n20158),.clk(gclk));
	jor g19859(.dina(n20158),.dinb(w_n430_14[0]),.dout(n20159),.clk(gclk));
	jand g19860(.dina(w_n20147_0[0]),.dinb(w_n430_13[2]),.dout(n20160),.clk(gclk));
	jand g19861(.dina(n20160),.dinb(w_n20157_0[0]),.dout(n20161),.clk(gclk));
	jnot g19862(.din(w_n19518_0[0]),.dout(n20162),.clk(gclk));
	jand g19863(.dina(w_asqrt3_6[1]),.dinb(n20162),.dout(n20163),.clk(gclk));
	jand g19864(.dina(w_n20163_0[1]),.dinb(w_n19525_0[0]),.dout(n20164),.clk(gclk));
	jor g19865(.dina(n20164),.dinb(w_n19523_0[0]),.dout(n20165),.clk(gclk));
	jand g19866(.dina(w_n20163_0[0]),.dinb(w_n19526_0[0]),.dout(n20166),.clk(gclk));
	jnot g19867(.din(n20166),.dout(n20167),.clk(gclk));
	jand g19868(.dina(n20167),.dinb(n20165),.dout(n20168),.clk(gclk));
	jnot g19869(.din(n20168),.dout(n20169),.clk(gclk));
	jor g19870(.dina(w_n20169_0[1]),.dinb(w_n20161_0[1]),.dout(n20170),.clk(gclk));
	jand g19871(.dina(n20170),.dinb(w_n20159_0[1]),.dout(n20171),.clk(gclk));
	jor g19872(.dina(w_n20171_0[1]),.dinb(w_n425_13[0]),.dout(n20172),.clk(gclk));
	jxor g19873(.dina(w_n19527_0[0]),.dinb(w_n430_13[1]),.dout(n20173),.clk(gclk));
	jor g19874(.dina(n20173),.dinb(w_n19616_8[0]),.dout(n20174),.clk(gclk));
	jxor g19875(.dina(n20174),.dinb(w_n19538_0[0]),.dout(n20175),.clk(gclk));
	jand g19876(.dina(w_n20171_0[0]),.dinb(w_n425_12[2]),.dout(n20176),.clk(gclk));
	jor g19877(.dina(w_n20176_0[1]),.dinb(w_n20175_0[1]),.dout(n20177),.clk(gclk));
	jand g19878(.dina(w_n20177_0[2]),.dinb(w_n20172_0[2]),.dout(n20178),.clk(gclk));
	jor g19879(.dina(n20178),.dinb(w_n305_14[1]),.dout(n20179),.clk(gclk));
	jand g19880(.dina(w_n20172_0[1]),.dinb(w_n305_14[0]),.dout(n20180),.clk(gclk));
	jand g19881(.dina(n20180),.dinb(w_n20177_0[1]),.dout(n20181),.clk(gclk));
	jnot g19882(.din(w_n19541_0[0]),.dout(n20182),.clk(gclk));
	jand g19883(.dina(w_asqrt3_6[0]),.dinb(n20182),.dout(n20183),.clk(gclk));
	jand g19884(.dina(w_n20183_0[1]),.dinb(w_n19548_0[0]),.dout(n20184),.clk(gclk));
	jor g19885(.dina(n20184),.dinb(w_n19546_0[0]),.dout(n20185),.clk(gclk));
	jand g19886(.dina(w_n20183_0[0]),.dinb(w_n19549_0[0]),.dout(n20186),.clk(gclk));
	jnot g19887(.din(n20186),.dout(n20187),.clk(gclk));
	jand g19888(.dina(n20187),.dinb(n20185),.dout(n20188),.clk(gclk));
	jnot g19889(.din(n20188),.dout(n20189),.clk(gclk));
	jor g19890(.dina(w_n20189_0[1]),.dinb(w_n20181_0[1]),.dout(n20190),.clk(gclk));
	jand g19891(.dina(n20190),.dinb(w_n20179_0[1]),.dout(n20191),.clk(gclk));
	jor g19892(.dina(w_n20191_0[2]),.dinb(w_n290_14[1]),.dout(n20192),.clk(gclk));
	jand g19893(.dina(w_n20191_0[1]),.dinb(w_n290_14[0]),.dout(n20193),.clk(gclk));
	jor g19894(.dina(n20193),.dinb(w_n19620_0[1]),.dout(n20194),.clk(gclk));
	jand g19895(.dina(w_n20194_0[1]),.dinb(w_n20192_0[1]),.dout(n20195),.clk(gclk));
	jor g19896(.dina(n20195),.dinb(w_n223_14[2]),.dout(n20196),.clk(gclk));
	jnot g19897(.din(w_n19557_0[0]),.dout(n20197),.clk(gclk));
	jor g19898(.dina(n20197),.dinb(w_n19555_0[0]),.dout(n20198),.clk(gclk));
	jor g19899(.dina(n20198),.dinb(w_n19616_7[2]),.dout(n20199),.clk(gclk));
	jxor g19900(.dina(n20199),.dinb(w_n19566_0[0]),.dout(n20200),.clk(gclk));
	jand g19901(.dina(w_n20192_0[0]),.dinb(w_n223_14[1]),.dout(n20201),.clk(gclk));
	jand g19902(.dina(n20201),.dinb(w_n20194_0[0]),.dout(n20202),.clk(gclk));
	jor g19903(.dina(w_n20202_0[1]),.dinb(w_n20200_0[1]),.dout(n20203),.clk(gclk));
	jand g19904(.dina(w_n20203_0[1]),.dinb(w_n20196_0[1]),.dout(n20204),.clk(gclk));
	jor g19905(.dina(w_n20204_0[2]),.dinb(w_n199_16[1]),.dout(n20205),.clk(gclk));
	jand g19906(.dina(w_n20204_0[1]),.dinb(w_n199_16[0]),.dout(n20206),.clk(gclk));
	jxor g19907(.dina(w_n19568_0[0]),.dinb(w_n223_14[0]),.dout(n20207),.clk(gclk));
	jor g19908(.dina(n20207),.dinb(w_n19616_7[1]),.dout(n20208),.clk(gclk));
	jxor g19909(.dina(n20208),.dinb(w_n19579_0[0]),.dout(n20209),.clk(gclk));
	jor g19910(.dina(w_n20209_0[1]),.dinb(n20206),.dout(n20210),.clk(gclk));
	jand g19911(.dina(n20210),.dinb(n20205),.dout(n20211),.clk(gclk));
	jnot g19912(.din(w_n19584_0[0]),.dout(n20212),.clk(gclk));
	jor g19913(.dina(n20212),.dinb(w_n19582_0[0]),.dout(n20213),.clk(gclk));
	jor g19914(.dina(n20213),.dinb(w_n19616_7[0]),.dout(n20214),.clk(gclk));
	jxor g19915(.dina(n20214),.dinb(w_n19593_0[0]),.dout(n20215),.clk(gclk));
	jnot g19916(.din(w_n19608_0[0]),.dout(n20216),.clk(gclk));
	jand g19917(.dina(w_asqrt3_5[2]),.dinb(w_n19607_0[1]),.dout(n20217),.clk(gclk));
	jand g19918(.dina(w_n20217_0[1]),.dinb(w_n19595_1[0]),.dout(n20218),.clk(gclk));
	jor g19919(.dina(n20218),.dinb(n20216),.dout(n20219),.clk(gclk));
	jor g19920(.dina(n20219),.dinb(w_n20215_0[2]),.dout(n20220),.clk(gclk));
	jor g19921(.dina(n20220),.dinb(w_n20211_0[2]),.dout(n20221),.clk(gclk));
	jand g19922(.dina(n20221),.dinb(w_n194_15[1]),.dout(n20222),.clk(gclk));
	jand g19923(.dina(w_n20215_0[1]),.dinb(w_n20211_0[1]),.dout(n20223),.clk(gclk));
	jor g19924(.dina(w_n20217_0[0]),.dinb(w_n19595_0[2]),.dout(n20224),.clk(gclk));
	jand g19925(.dina(w_n19607_0[0]),.dinb(w_n19595_0[1]),.dout(n20225),.clk(gclk));
	jor g19926(.dina(n20225),.dinb(w_n194_15[0]),.dout(n20226),.clk(gclk));
	jnot g19927(.din(n20226),.dout(n20227),.clk(gclk));
	jand g19928(.dina(n20227),.dinb(n20224),.dout(n20228),.clk(gclk));
	jor g19929(.dina(n20228),.dinb(w_n20223_0[1]),.dout(n20229),.clk(gclk));
	jor g19930(.dina(n20229),.dinb(n20222),.dout(asqrt_fa_3),.clk(gclk));
	jxor g19931(.dina(w_n20191_0[0]),.dinb(w_n290_13[2]),.dout(n20231),.clk(gclk));
	jand g19932(.dina(n20231),.dinb(w_asqrt2_31),.dout(n20232),.clk(gclk));
	jxor g19933(.dina(n20232),.dinb(w_n19620_0[0]),.dout(n20233),.clk(gclk));
	jnot g19934(.din(n20233),.dout(n20234),.clk(gclk));
	jand g19935(.dina(w_asqrt2_30[2]),.dinb(w_a4_0[0]),.dout(n20235),.clk(gclk));
	jnot g19936(.din(w_a2_0[2]),.dout(n20236),.clk(gclk));
	jnot g19937(.din(w_a3_0[1]),.dout(n20237),.clk(gclk));
	jand g19938(.dina(w_n19622_1[0]),.dinb(w_n20237_0[1]),.dout(n20238),.clk(gclk));
	jand g19939(.dina(n20238),.dinb(w_n20236_0[1]),.dout(n20239),.clk(gclk));
	jor g19940(.dina(n20239),.dinb(n20235),.dout(n20240),.clk(gclk));
	jand g19941(.dina(w_n20240_0[2]),.dinb(w_asqrt3_5[1]),.dout(n20241),.clk(gclk));
	jand g19942(.dina(w_asqrt2_30[1]),.dinb(w_n19622_0[2]),.dout(n20242),.clk(gclk));
	jxor g19943(.dina(w_n20242_0[1]),.dinb(w_n19623_0[1]),.dout(n20243),.clk(gclk));
	jor g19944(.dina(w_n20240_0[1]),.dinb(w_asqrt3_5[0]),.dout(n20244),.clk(gclk));
	jand g19945(.dina(n20244),.dinb(w_n20243_0[1]),.dout(n20245),.clk(gclk));
	jor g19946(.dina(w_n20245_0[1]),.dinb(w_n20241_0[1]),.dout(n20246),.clk(gclk));
	jand g19947(.dina(n20246),.dinb(w_asqrt4_10[2]),.dout(n20247),.clk(gclk));
	jor g19948(.dina(w_n20241_0[0]),.dinb(w_asqrt4_10[1]),.dout(n20248),.clk(gclk));
	jor g19949(.dina(n20248),.dinb(w_n20245_0[0]),.dout(n20249),.clk(gclk));
	jand g19950(.dina(w_n20242_0[0]),.dinb(w_n19623_0[0]),.dout(n20250),.clk(gclk));
	jnot g19951(.din(w_asqrt2_30[0]),.dout(n20251),.clk(gclk));
	jand g19952(.dina(w_n20251_1[1]),.dinb(w_asqrt3_4[2]),.dout(n20252),.clk(gclk));
	jor g19953(.dina(n20252),.dinb(n20250),.dout(n20253),.clk(gclk));
	jxor g19954(.dina(n20253),.dinb(w_n18961_0[1]),.dout(n20254),.clk(gclk));
	jand g19955(.dina(w_n20254_0[1]),.dinb(w_n20249_0[1]),.dout(n20255),.clk(gclk));
	jor g19956(.dina(n20255),.dinb(w_n20247_0[1]),.dout(n20256),.clk(gclk));
	jand g19957(.dina(w_n20256_0[2]),.dinb(w_asqrt5_5[1]),.dout(n20257),.clk(gclk));
	jor g19958(.dina(w_n20256_0[1]),.dinb(w_asqrt5_5[0]),.dout(n20258),.clk(gclk));
	jxor g19959(.dina(w_n19627_0[0]),.dinb(w_n18976_1[1]),.dout(n20259),.clk(gclk));
	jand g19960(.dina(n20259),.dinb(w_asqrt2_29[2]),.dout(n20260),.clk(gclk));
	jxor g19961(.dina(n20260),.dinb(w_n19630_0[0]),.dout(n20261),.clk(gclk));
	jnot g19962(.din(n20261),.dout(n20262),.clk(gclk));
	jand g19963(.dina(w_n20262_0[1]),.dinb(n20258),.dout(n20263),.clk(gclk));
	jor g19964(.dina(w_n20263_0[1]),.dinb(w_n20257_0[1]),.dout(n20264),.clk(gclk));
	jand g19965(.dina(n20264),.dinb(w_asqrt6_10[2]),.dout(n20265),.clk(gclk));
	jnot g19966(.din(w_n19636_0[0]),.dout(n20266),.clk(gclk));
	jand g19967(.dina(n20266),.dinb(w_n19634_0[0]),.dout(n20267),.clk(gclk));
	jand g19968(.dina(n20267),.dinb(w_asqrt2_29[1]),.dout(n20268),.clk(gclk));
	jxor g19969(.dina(n20268),.dinb(w_n19641_0[0]),.dout(n20269),.clk(gclk));
	jnot g19970(.din(w_n20269_0[1]),.dout(n20270),.clk(gclk));
	jor g19971(.dina(w_n20257_0[0]),.dinb(w_asqrt6_10[1]),.dout(n20271),.clk(gclk));
	jor g19972(.dina(n20271),.dinb(w_n20263_0[0]),.dout(n20272),.clk(gclk));
	jand g19973(.dina(w_n20272_0[1]),.dinb(n20270),.dout(n20273),.clk(gclk));
	jor g19974(.dina(w_n20273_0[1]),.dinb(w_n20265_0[1]),.dout(n20274),.clk(gclk));
	jand g19975(.dina(w_n20274_0[2]),.dinb(w_asqrt7_5[1]),.dout(n20275),.clk(gclk));
	jor g19976(.dina(w_n20274_0[1]),.dinb(w_asqrt7_5[0]),.dout(n20276),.clk(gclk));
	jnot g19977(.din(w_n19648_0[0]),.dout(n20277),.clk(gclk));
	jxor g19978(.dina(w_n19643_0[0]),.dinb(w_n18360_1[2]),.dout(n20278),.clk(gclk));
	jand g19979(.dina(n20278),.dinb(w_asqrt2_29[0]),.dout(n20279),.clk(gclk));
	jxor g19980(.dina(n20279),.dinb(n20277),.dout(n20280),.clk(gclk));
	jand g19981(.dina(w_n20280_0[1]),.dinb(n20276),.dout(n20281),.clk(gclk));
	jor g19982(.dina(w_n20281_0[1]),.dinb(w_n20275_0[1]),.dout(n20282),.clk(gclk));
	jand g19983(.dina(n20282),.dinb(w_asqrt8_10[2]),.dout(n20283),.clk(gclk));
	jor g19984(.dina(w_n20275_0[0]),.dinb(w_asqrt8_10[1]),.dout(n20284),.clk(gclk));
	jor g19985(.dina(n20284),.dinb(w_n20281_0[0]),.dout(n20285),.clk(gclk));
	jnot g19986(.din(w_n19655_0[0]),.dout(n20286),.clk(gclk));
	jnot g19987(.din(w_n19657_0[0]),.dout(n20287),.clk(gclk));
	jand g19988(.dina(w_asqrt2_28[2]),.dinb(w_n19651_0[0]),.dout(n20288),.clk(gclk));
	jand g19989(.dina(w_n20288_0[1]),.dinb(n20287),.dout(n20289),.clk(gclk));
	jor g19990(.dina(n20289),.dinb(n20286),.dout(n20290),.clk(gclk));
	jnot g19991(.din(w_n19658_0[0]),.dout(n20291),.clk(gclk));
	jand g19992(.dina(w_n20288_0[0]),.dinb(n20291),.dout(n20292),.clk(gclk));
	jnot g19993(.din(n20292),.dout(n20293),.clk(gclk));
	jand g19994(.dina(n20293),.dinb(n20290),.dout(n20294),.clk(gclk));
	jand g19995(.dina(w_n20294_0[1]),.dinb(w_n20285_0[1]),.dout(n20295),.clk(gclk));
	jor g19996(.dina(n20295),.dinb(w_n20283_0[1]),.dout(n20296),.clk(gclk));
	jand g19997(.dina(w_n20296_0[2]),.dinb(w_asqrt9_5[2]),.dout(n20297),.clk(gclk));
	jor g19998(.dina(w_n20296_0[1]),.dinb(w_asqrt9_5[1]),.dout(n20298),.clk(gclk));
	jxor g19999(.dina(w_n19659_0[0]),.dinb(w_n17135_2[1]),.dout(n20299),.clk(gclk));
	jand g20000(.dina(n20299),.dinb(w_asqrt2_28[1]),.dout(n20300),.clk(gclk));
	jxor g20001(.dina(n20300),.dinb(w_n19664_0[0]),.dout(n20301),.clk(gclk));
	jand g20002(.dina(w_n20301_0[1]),.dinb(n20298),.dout(n20302),.clk(gclk));
	jor g20003(.dina(w_n20302_0[1]),.dinb(w_n20297_0[1]),.dout(n20303),.clk(gclk));
	jand g20004(.dina(n20303),.dinb(w_asqrt10_10[2]),.dout(n20304),.clk(gclk));
	jnot g20005(.din(w_n19670_0[0]),.dout(n20305),.clk(gclk));
	jand g20006(.dina(n20305),.dinb(w_n19668_0[0]),.dout(n20306),.clk(gclk));
	jand g20007(.dina(n20306),.dinb(w_asqrt2_28[0]),.dout(n20307),.clk(gclk));
	jxor g20008(.dina(n20307),.dinb(w_n19678_0[0]),.dout(n20308),.clk(gclk));
	jnot g20009(.din(w_n20308_0[1]),.dout(n20309),.clk(gclk));
	jor g20010(.dina(w_n20297_0[0]),.dinb(w_asqrt10_10[1]),.dout(n20310),.clk(gclk));
	jor g20011(.dina(n20310),.dinb(w_n20302_0[0]),.dout(n20311),.clk(gclk));
	jand g20012(.dina(w_n20311_0[1]),.dinb(n20309),.dout(n20312),.clk(gclk));
	jor g20013(.dina(w_n20312_0[1]),.dinb(w_n20304_0[1]),.dout(n20313),.clk(gclk));
	jand g20014(.dina(w_n20313_0[2]),.dinb(w_asqrt11_5[2]),.dout(n20314),.clk(gclk));
	jor g20015(.dina(w_n20313_0[1]),.dinb(w_asqrt11_5[1]),.dout(n20315),.clk(gclk));
	jxor g20016(.dina(w_n19680_0[0]),.dinb(w_n15950_2[2]),.dout(n20316),.clk(gclk));
	jand g20017(.dina(n20316),.dinb(w_asqrt2_27[2]),.dout(n20317),.clk(gclk));
	jxor g20018(.dina(n20317),.dinb(w_n19686_0[0]),.dout(n20318),.clk(gclk));
	jand g20019(.dina(w_n20318_0[1]),.dinb(n20315),.dout(n20319),.clk(gclk));
	jor g20020(.dina(w_n20319_0[1]),.dinb(w_n20314_0[1]),.dout(n20320),.clk(gclk));
	jand g20021(.dina(n20320),.dinb(w_asqrt12_10[2]),.dout(n20321),.clk(gclk));
	jor g20022(.dina(w_n20314_0[0]),.dinb(w_asqrt12_10[1]),.dout(n20322),.clk(gclk));
	jor g20023(.dina(n20322),.dinb(w_n20319_0[0]),.dout(n20323),.clk(gclk));
	jnot g20024(.din(w_n19694_0[0]),.dout(n20324),.clk(gclk));
	jnot g20025(.din(w_n19696_0[0]),.dout(n20325),.clk(gclk));
	jand g20026(.dina(w_asqrt2_27[1]),.dinb(w_n19690_0[0]),.dout(n20326),.clk(gclk));
	jand g20027(.dina(w_n20326_0[1]),.dinb(n20325),.dout(n20327),.clk(gclk));
	jor g20028(.dina(n20327),.dinb(n20324),.dout(n20328),.clk(gclk));
	jnot g20029(.din(w_n19697_0[0]),.dout(n20329),.clk(gclk));
	jand g20030(.dina(w_n20326_0[0]),.dinb(n20329),.dout(n20330),.clk(gclk));
	jnot g20031(.din(n20330),.dout(n20331),.clk(gclk));
	jand g20032(.dina(n20331),.dinb(n20328),.dout(n20332),.clk(gclk));
	jand g20033(.dina(w_n20332_0[1]),.dinb(w_n20323_0[1]),.dout(n20333),.clk(gclk));
	jor g20034(.dina(n20333),.dinb(w_n20321_0[1]),.dout(n20334),.clk(gclk));
	jand g20035(.dina(w_n20334_0[1]),.dinb(w_asqrt13_6[0]),.dout(n20335),.clk(gclk));
	jxor g20036(.dina(w_n19698_0[0]),.dinb(w_n14816_3[1]),.dout(n20336),.clk(gclk));
	jand g20037(.dina(n20336),.dinb(w_asqrt2_27[0]),.dout(n20337),.clk(gclk));
	jxor g20038(.dina(n20337),.dinb(w_n19705_0[0]),.dout(n20338),.clk(gclk));
	jnot g20039(.din(w_n20338_0[1]),.dout(n20339),.clk(gclk));
	jor g20040(.dina(w_n20334_0[0]),.dinb(w_asqrt13_5[2]),.dout(n20340),.clk(gclk));
	jand g20041(.dina(w_n20340_0[1]),.dinb(n20339),.dout(n20341),.clk(gclk));
	jor g20042(.dina(w_n20341_0[2]),.dinb(w_n20335_0[2]),.dout(n20342),.clk(gclk));
	jand g20043(.dina(n20342),.dinb(w_asqrt14_10[2]),.dout(n20343),.clk(gclk));
	jnot g20044(.din(w_n19710_0[0]),.dout(n20344),.clk(gclk));
	jand g20045(.dina(n20344),.dinb(w_n19708_0[0]),.dout(n20345),.clk(gclk));
	jand g20046(.dina(n20345),.dinb(w_asqrt2_26[2]),.dout(n20346),.clk(gclk));
	jxor g20047(.dina(n20346),.dinb(w_n19718_0[0]),.dout(n20347),.clk(gclk));
	jnot g20048(.din(w_n20347_0[1]),.dout(n20348),.clk(gclk));
	jor g20049(.dina(w_n20335_0[1]),.dinb(w_asqrt14_10[1]),.dout(n20349),.clk(gclk));
	jor g20050(.dina(n20349),.dinb(w_n20341_0[1]),.dout(n20350),.clk(gclk));
	jand g20051(.dina(w_n20350_0[1]),.dinb(n20348),.dout(n20351),.clk(gclk));
	jor g20052(.dina(w_n20351_0[1]),.dinb(w_n20343_0[1]),.dout(n20352),.clk(gclk));
	jand g20053(.dina(w_n20352_0[2]),.dinb(w_asqrt15_6[0]),.dout(n20353),.clk(gclk));
	jor g20054(.dina(w_n20352_0[1]),.dinb(w_asqrt15_5[2]),.dout(n20354),.clk(gclk));
	jnot g20055(.din(w_n19724_0[0]),.dout(n20355),.clk(gclk));
	jnot g20056(.din(w_n19725_0[0]),.dout(n20356),.clk(gclk));
	jand g20057(.dina(w_asqrt2_26[1]),.dinb(w_n19721_0[0]),.dout(n20357),.clk(gclk));
	jand g20058(.dina(w_n20357_0[1]),.dinb(n20356),.dout(n20358),.clk(gclk));
	jor g20059(.dina(n20358),.dinb(n20355),.dout(n20359),.clk(gclk));
	jnot g20060(.din(w_n19726_0[0]),.dout(n20360),.clk(gclk));
	jand g20061(.dina(w_n20357_0[0]),.dinb(n20360),.dout(n20361),.clk(gclk));
	jnot g20062(.din(n20361),.dout(n20362),.clk(gclk));
	jand g20063(.dina(n20362),.dinb(n20359),.dout(n20363),.clk(gclk));
	jand g20064(.dina(w_n20363_0[1]),.dinb(n20354),.dout(n20364),.clk(gclk));
	jor g20065(.dina(w_n20364_0[1]),.dinb(w_n20353_0[1]),.dout(n20365),.clk(gclk));
	jand g20066(.dina(n20365),.dinb(w_asqrt16_10[2]),.dout(n20366),.clk(gclk));
	jor g20067(.dina(w_n20353_0[0]),.dinb(w_asqrt16_10[1]),.dout(n20367),.clk(gclk));
	jor g20068(.dina(n20367),.dinb(w_n20364_0[0]),.dout(n20368),.clk(gclk));
	jnot g20069(.din(w_n19732_0[0]),.dout(n20369),.clk(gclk));
	jnot g20070(.din(w_n19734_0[0]),.dout(n20370),.clk(gclk));
	jand g20071(.dina(w_asqrt2_26[0]),.dinb(w_n19728_0[0]),.dout(n20371),.clk(gclk));
	jand g20072(.dina(w_n20371_0[1]),.dinb(n20370),.dout(n20372),.clk(gclk));
	jor g20073(.dina(n20372),.dinb(n20369),.dout(n20373),.clk(gclk));
	jnot g20074(.din(w_n19735_0[0]),.dout(n20374),.clk(gclk));
	jand g20075(.dina(w_n20371_0[0]),.dinb(n20374),.dout(n20375),.clk(gclk));
	jnot g20076(.din(n20375),.dout(n20376),.clk(gclk));
	jand g20077(.dina(n20376),.dinb(n20373),.dout(n20377),.clk(gclk));
	jand g20078(.dina(w_n20377_0[1]),.dinb(w_n20368_0[1]),.dout(n20378),.clk(gclk));
	jor g20079(.dina(n20378),.dinb(w_n20366_0[1]),.dout(n20379),.clk(gclk));
	jand g20080(.dina(w_n20379_0[1]),.dinb(w_asqrt17_6[1]),.dout(n20380),.clk(gclk));
	jxor g20081(.dina(w_n19736_0[0]),.dinb(w_n12670_4[0]),.dout(n20381),.clk(gclk));
	jand g20082(.dina(n20381),.dinb(w_asqrt2_25[2]),.dout(n20382),.clk(gclk));
	jxor g20083(.dina(n20382),.dinb(w_n19746_0[0]),.dout(n20383),.clk(gclk));
	jnot g20084(.din(w_n20383_0[1]),.dout(n20384),.clk(gclk));
	jor g20085(.dina(w_n20379_0[0]),.dinb(w_asqrt17_6[0]),.dout(n20385),.clk(gclk));
	jand g20086(.dina(w_n20385_0[1]),.dinb(n20384),.dout(n20386),.clk(gclk));
	jor g20087(.dina(w_n20386_0[2]),.dinb(w_n20380_0[2]),.dout(n20387),.clk(gclk));
	jand g20088(.dina(n20387),.dinb(w_asqrt18_10[2]),.dout(n20388),.clk(gclk));
	jnot g20089(.din(w_n19751_0[0]),.dout(n20389),.clk(gclk));
	jand g20090(.dina(n20389),.dinb(w_n19749_0[0]),.dout(n20390),.clk(gclk));
	jand g20091(.dina(n20390),.dinb(w_asqrt2_25[1]),.dout(n20391),.clk(gclk));
	jxor g20092(.dina(n20391),.dinb(w_n19759_0[0]),.dout(n20392),.clk(gclk));
	jnot g20093(.din(w_n20392_0[1]),.dout(n20393),.clk(gclk));
	jor g20094(.dina(w_n20380_0[1]),.dinb(w_asqrt18_10[1]),.dout(n20394),.clk(gclk));
	jor g20095(.dina(n20394),.dinb(w_n20386_0[1]),.dout(n20395),.clk(gclk));
	jand g20096(.dina(w_n20395_0[1]),.dinb(n20393),.dout(n20396),.clk(gclk));
	jor g20097(.dina(w_n20396_0[1]),.dinb(w_n20388_0[1]),.dout(n20397),.clk(gclk));
	jand g20098(.dina(w_n20397_0[2]),.dinb(w_asqrt19_6[1]),.dout(n20398),.clk(gclk));
	jor g20099(.dina(w_n20397_0[1]),.dinb(w_asqrt19_6[0]),.dout(n20399),.clk(gclk));
	jnot g20100(.din(w_n19765_0[0]),.dout(n20400),.clk(gclk));
	jnot g20101(.din(w_n19766_0[0]),.dout(n20401),.clk(gclk));
	jand g20102(.dina(w_asqrt2_25[0]),.dinb(w_n19762_0[0]),.dout(n20402),.clk(gclk));
	jand g20103(.dina(w_n20402_0[1]),.dinb(n20401),.dout(n20403),.clk(gclk));
	jor g20104(.dina(n20403),.dinb(n20400),.dout(n20404),.clk(gclk));
	jnot g20105(.din(w_n19767_0[0]),.dout(n20405),.clk(gclk));
	jand g20106(.dina(w_n20402_0[0]),.dinb(n20405),.dout(n20406),.clk(gclk));
	jnot g20107(.din(n20406),.dout(n20407),.clk(gclk));
	jand g20108(.dina(n20407),.dinb(n20404),.dout(n20408),.clk(gclk));
	jand g20109(.dina(w_n20408_0[1]),.dinb(n20399),.dout(n20409),.clk(gclk));
	jor g20110(.dina(w_n20409_0[1]),.dinb(w_n20398_0[1]),.dout(n20410),.clk(gclk));
	jand g20111(.dina(n20410),.dinb(w_asqrt20_10[2]),.dout(n20411),.clk(gclk));
	jor g20112(.dina(w_n20398_0[0]),.dinb(w_asqrt20_10[1]),.dout(n20412),.clk(gclk));
	jor g20113(.dina(n20412),.dinb(w_n20409_0[0]),.dout(n20413),.clk(gclk));
	jnot g20114(.din(w_n19773_0[0]),.dout(n20414),.clk(gclk));
	jnot g20115(.din(w_n19775_0[0]),.dout(n20415),.clk(gclk));
	jand g20116(.dina(w_asqrt2_24[2]),.dinb(w_n19769_0[0]),.dout(n20416),.clk(gclk));
	jand g20117(.dina(w_n20416_0[1]),.dinb(n20415),.dout(n20417),.clk(gclk));
	jor g20118(.dina(n20417),.dinb(n20414),.dout(n20418),.clk(gclk));
	jnot g20119(.din(w_n19776_0[0]),.dout(n20419),.clk(gclk));
	jand g20120(.dina(w_n20416_0[0]),.dinb(n20419),.dout(n20420),.clk(gclk));
	jnot g20121(.din(n20420),.dout(n20421),.clk(gclk));
	jand g20122(.dina(n20421),.dinb(n20418),.dout(n20422),.clk(gclk));
	jand g20123(.dina(w_n20422_0[1]),.dinb(w_n20413_0[1]),.dout(n20423),.clk(gclk));
	jor g20124(.dina(n20423),.dinb(w_n20411_0[1]),.dout(n20424),.clk(gclk));
	jand g20125(.dina(w_n20424_0[1]),.dinb(w_asqrt21_6[2]),.dout(n20425),.clk(gclk));
	jxor g20126(.dina(w_n19777_0[0]),.dinb(w_n10696_5[0]),.dout(n20426),.clk(gclk));
	jand g20127(.dina(n20426),.dinb(w_asqrt2_24[1]),.dout(n20427),.clk(gclk));
	jxor g20128(.dina(n20427),.dinb(w_n19787_0[0]),.dout(n20428),.clk(gclk));
	jnot g20129(.din(w_n20428_0[1]),.dout(n20429),.clk(gclk));
	jor g20130(.dina(w_n20424_0[0]),.dinb(w_asqrt21_6[1]),.dout(n20430),.clk(gclk));
	jand g20131(.dina(w_n20430_0[1]),.dinb(n20429),.dout(n20431),.clk(gclk));
	jor g20132(.dina(w_n20431_0[2]),.dinb(w_n20425_0[2]),.dout(n20432),.clk(gclk));
	jand g20133(.dina(n20432),.dinb(w_asqrt22_10[2]),.dout(n20433),.clk(gclk));
	jnot g20134(.din(w_n19792_0[0]),.dout(n20434),.clk(gclk));
	jand g20135(.dina(n20434),.dinb(w_n19790_0[0]),.dout(n20435),.clk(gclk));
	jand g20136(.dina(n20435),.dinb(w_asqrt2_24[0]),.dout(n20436),.clk(gclk));
	jxor g20137(.dina(n20436),.dinb(w_n19800_0[0]),.dout(n20437),.clk(gclk));
	jnot g20138(.din(w_n20437_0[1]),.dout(n20438),.clk(gclk));
	jor g20139(.dina(w_n20425_0[1]),.dinb(w_asqrt22_10[1]),.dout(n20439),.clk(gclk));
	jor g20140(.dina(n20439),.dinb(w_n20431_0[1]),.dout(n20440),.clk(gclk));
	jand g20141(.dina(w_n20440_0[1]),.dinb(n20438),.dout(n20441),.clk(gclk));
	jor g20142(.dina(w_n20441_0[1]),.dinb(w_n20433_0[1]),.dout(n20442),.clk(gclk));
	jand g20143(.dina(w_n20442_0[2]),.dinb(w_asqrt23_6[2]),.dout(n20443),.clk(gclk));
	jor g20144(.dina(w_n20442_0[1]),.dinb(w_asqrt23_6[1]),.dout(n20444),.clk(gclk));
	jnot g20145(.din(w_n19806_0[0]),.dout(n20445),.clk(gclk));
	jnot g20146(.din(w_n19807_0[0]),.dout(n20446),.clk(gclk));
	jand g20147(.dina(w_asqrt2_23[2]),.dinb(w_n19803_0[0]),.dout(n20447),.clk(gclk));
	jand g20148(.dina(w_n20447_0[1]),.dinb(n20446),.dout(n20448),.clk(gclk));
	jor g20149(.dina(n20448),.dinb(n20445),.dout(n20449),.clk(gclk));
	jnot g20150(.din(w_n19808_0[0]),.dout(n20450),.clk(gclk));
	jand g20151(.dina(w_n20447_0[0]),.dinb(n20450),.dout(n20451),.clk(gclk));
	jnot g20152(.din(n20451),.dout(n20452),.clk(gclk));
	jand g20153(.dina(n20452),.dinb(n20449),.dout(n20453),.clk(gclk));
	jand g20154(.dina(w_n20453_0[1]),.dinb(n20444),.dout(n20454),.clk(gclk));
	jor g20155(.dina(w_n20454_0[1]),.dinb(w_n20443_0[1]),.dout(n20455),.clk(gclk));
	jand g20156(.dina(n20455),.dinb(w_asqrt24_10[2]),.dout(n20456),.clk(gclk));
	jor g20157(.dina(w_n20443_0[0]),.dinb(w_asqrt24_10[1]),.dout(n20457),.clk(gclk));
	jor g20158(.dina(n20457),.dinb(w_n20454_0[0]),.dout(n20458),.clk(gclk));
	jnot g20159(.din(w_n19814_0[0]),.dout(n20459),.clk(gclk));
	jnot g20160(.din(w_n19816_0[0]),.dout(n20460),.clk(gclk));
	jand g20161(.dina(w_asqrt2_23[1]),.dinb(w_n19810_0[0]),.dout(n20461),.clk(gclk));
	jand g20162(.dina(w_n20461_0[1]),.dinb(n20460),.dout(n20462),.clk(gclk));
	jor g20163(.dina(n20462),.dinb(n20459),.dout(n20463),.clk(gclk));
	jnot g20164(.din(w_n19817_0[0]),.dout(n20464),.clk(gclk));
	jand g20165(.dina(w_n20461_0[0]),.dinb(n20464),.dout(n20465),.clk(gclk));
	jnot g20166(.din(n20465),.dout(n20466),.clk(gclk));
	jand g20167(.dina(n20466),.dinb(n20463),.dout(n20467),.clk(gclk));
	jand g20168(.dina(w_n20467_0[1]),.dinb(w_n20458_0[1]),.dout(n20468),.clk(gclk));
	jor g20169(.dina(n20468),.dinb(w_n20456_0[1]),.dout(n20469),.clk(gclk));
	jand g20170(.dina(w_n20469_0[1]),.dinb(w_asqrt25_7[0]),.dout(n20470),.clk(gclk));
	jxor g20171(.dina(w_n19818_0[0]),.dinb(w_n8893_5[2]),.dout(n20471),.clk(gclk));
	jand g20172(.dina(n20471),.dinb(w_asqrt2_23[0]),.dout(n20472),.clk(gclk));
	jxor g20173(.dina(n20472),.dinb(w_n19828_0[0]),.dout(n20473),.clk(gclk));
	jnot g20174(.din(w_n20473_0[1]),.dout(n20474),.clk(gclk));
	jor g20175(.dina(w_n20469_0[0]),.dinb(w_asqrt25_6[2]),.dout(n20475),.clk(gclk));
	jand g20176(.dina(w_n20475_0[1]),.dinb(n20474),.dout(n20476),.clk(gclk));
	jor g20177(.dina(w_n20476_0[2]),.dinb(w_n20470_0[2]),.dout(n20477),.clk(gclk));
	jand g20178(.dina(n20477),.dinb(w_asqrt26_10[2]),.dout(n20478),.clk(gclk));
	jnot g20179(.din(w_n19833_0[0]),.dout(n20479),.clk(gclk));
	jand g20180(.dina(n20479),.dinb(w_n19831_0[0]),.dout(n20480),.clk(gclk));
	jand g20181(.dina(n20480),.dinb(w_asqrt2_22[2]),.dout(n20481),.clk(gclk));
	jxor g20182(.dina(n20481),.dinb(w_n19841_0[0]),.dout(n20482),.clk(gclk));
	jnot g20183(.din(w_n20482_0[1]),.dout(n20483),.clk(gclk));
	jor g20184(.dina(w_n20470_0[1]),.dinb(w_asqrt26_10[1]),.dout(n20484),.clk(gclk));
	jor g20185(.dina(n20484),.dinb(w_n20476_0[1]),.dout(n20485),.clk(gclk));
	jand g20186(.dina(w_n20485_0[1]),.dinb(n20483),.dout(n20486),.clk(gclk));
	jor g20187(.dina(w_n20486_0[1]),.dinb(w_n20478_0[1]),.dout(n20487),.clk(gclk));
	jand g20188(.dina(w_n20487_0[2]),.dinb(w_asqrt27_7[0]),.dout(n20488),.clk(gclk));
	jor g20189(.dina(w_n20487_0[1]),.dinb(w_asqrt27_6[2]),.dout(n20489),.clk(gclk));
	jnot g20190(.din(w_n19847_0[0]),.dout(n20490),.clk(gclk));
	jnot g20191(.din(w_n19848_0[0]),.dout(n20491),.clk(gclk));
	jand g20192(.dina(w_asqrt2_22[1]),.dinb(w_n19844_0[0]),.dout(n20492),.clk(gclk));
	jand g20193(.dina(w_n20492_0[1]),.dinb(n20491),.dout(n20493),.clk(gclk));
	jor g20194(.dina(n20493),.dinb(n20490),.dout(n20494),.clk(gclk));
	jnot g20195(.din(w_n19849_0[0]),.dout(n20495),.clk(gclk));
	jand g20196(.dina(w_n20492_0[0]),.dinb(n20495),.dout(n20496),.clk(gclk));
	jnot g20197(.din(n20496),.dout(n20497),.clk(gclk));
	jand g20198(.dina(n20497),.dinb(n20494),.dout(n20498),.clk(gclk));
	jand g20199(.dina(w_n20498_0[1]),.dinb(n20489),.dout(n20499),.clk(gclk));
	jor g20200(.dina(w_n20499_0[1]),.dinb(w_n20488_0[1]),.dout(n20500),.clk(gclk));
	jand g20201(.dina(n20500),.dinb(w_asqrt28_10[2]),.dout(n20501),.clk(gclk));
	jor g20202(.dina(w_n20488_0[0]),.dinb(w_asqrt28_10[1]),.dout(n20502),.clk(gclk));
	jor g20203(.dina(n20502),.dinb(w_n20499_0[0]),.dout(n20503),.clk(gclk));
	jnot g20204(.din(w_n19855_0[0]),.dout(n20504),.clk(gclk));
	jnot g20205(.din(w_n19857_0[0]),.dout(n20505),.clk(gclk));
	jand g20206(.dina(w_asqrt2_22[0]),.dinb(w_n19851_0[0]),.dout(n20506),.clk(gclk));
	jand g20207(.dina(w_n20506_0[1]),.dinb(n20505),.dout(n20507),.clk(gclk));
	jor g20208(.dina(n20507),.dinb(n20504),.dout(n20508),.clk(gclk));
	jnot g20209(.din(w_n19858_0[0]),.dout(n20509),.clk(gclk));
	jand g20210(.dina(w_n20506_0[0]),.dinb(n20509),.dout(n20510),.clk(gclk));
	jnot g20211(.din(n20510),.dout(n20511),.clk(gclk));
	jand g20212(.dina(n20511),.dinb(n20508),.dout(n20512),.clk(gclk));
	jand g20213(.dina(w_n20512_0[1]),.dinb(w_n20503_0[1]),.dout(n20513),.clk(gclk));
	jor g20214(.dina(n20513),.dinb(w_n20501_0[1]),.dout(n20514),.clk(gclk));
	jand g20215(.dina(w_n20514_0[1]),.dinb(w_asqrt29_7[1]),.dout(n20515),.clk(gclk));
	jxor g20216(.dina(w_n19859_0[0]),.dinb(w_n7260_6[2]),.dout(n20516),.clk(gclk));
	jand g20217(.dina(n20516),.dinb(w_asqrt2_21[2]),.dout(n20517),.clk(gclk));
	jxor g20218(.dina(n20517),.dinb(w_n19869_0[0]),.dout(n20518),.clk(gclk));
	jnot g20219(.din(w_n20518_0[1]),.dout(n20519),.clk(gclk));
	jor g20220(.dina(w_n20514_0[0]),.dinb(w_asqrt29_7[0]),.dout(n20520),.clk(gclk));
	jand g20221(.dina(w_n20520_0[1]),.dinb(n20519),.dout(n20521),.clk(gclk));
	jor g20222(.dina(w_n20521_0[2]),.dinb(w_n20515_0[2]),.dout(n20522),.clk(gclk));
	jand g20223(.dina(n20522),.dinb(w_asqrt30_10[2]),.dout(n20523),.clk(gclk));
	jnot g20224(.din(w_n19874_0[0]),.dout(n20524),.clk(gclk));
	jand g20225(.dina(n20524),.dinb(w_n19872_0[0]),.dout(n20525),.clk(gclk));
	jand g20226(.dina(n20525),.dinb(w_asqrt2_21[1]),.dout(n20526),.clk(gclk));
	jxor g20227(.dina(n20526),.dinb(w_n19882_0[0]),.dout(n20527),.clk(gclk));
	jnot g20228(.din(w_n20527_0[1]),.dout(n20528),.clk(gclk));
	jor g20229(.dina(w_n20515_0[1]),.dinb(w_asqrt30_10[1]),.dout(n20529),.clk(gclk));
	jor g20230(.dina(n20529),.dinb(w_n20521_0[1]),.dout(n20530),.clk(gclk));
	jand g20231(.dina(w_n20530_0[1]),.dinb(n20528),.dout(n20531),.clk(gclk));
	jor g20232(.dina(w_n20531_0[1]),.dinb(w_n20523_0[1]),.dout(n20532),.clk(gclk));
	jand g20233(.dina(w_n20532_0[2]),.dinb(w_asqrt31_7[1]),.dout(n20533),.clk(gclk));
	jor g20234(.dina(w_n20532_0[1]),.dinb(w_asqrt31_7[0]),.dout(n20534),.clk(gclk));
	jnot g20235(.din(w_n19888_0[0]),.dout(n20535),.clk(gclk));
	jnot g20236(.din(w_n19889_0[0]),.dout(n20536),.clk(gclk));
	jand g20237(.dina(w_asqrt2_21[0]),.dinb(w_n19885_0[0]),.dout(n20537),.clk(gclk));
	jand g20238(.dina(w_n20537_0[1]),.dinb(n20536),.dout(n20538),.clk(gclk));
	jor g20239(.dina(n20538),.dinb(n20535),.dout(n20539),.clk(gclk));
	jnot g20240(.din(w_n19890_0[0]),.dout(n20540),.clk(gclk));
	jand g20241(.dina(w_n20537_0[0]),.dinb(n20540),.dout(n20541),.clk(gclk));
	jnot g20242(.din(n20541),.dout(n20542),.clk(gclk));
	jand g20243(.dina(n20542),.dinb(n20539),.dout(n20543),.clk(gclk));
	jand g20244(.dina(w_n20543_0[1]),.dinb(n20534),.dout(n20544),.clk(gclk));
	jor g20245(.dina(w_n20544_0[1]),.dinb(w_n20533_0[1]),.dout(n20545),.clk(gclk));
	jand g20246(.dina(n20545),.dinb(w_asqrt32_10[2]),.dout(n20546),.clk(gclk));
	jor g20247(.dina(w_n20533_0[0]),.dinb(w_asqrt32_10[1]),.dout(n20547),.clk(gclk));
	jor g20248(.dina(n20547),.dinb(w_n20544_0[0]),.dout(n20548),.clk(gclk));
	jnot g20249(.din(w_n19896_0[0]),.dout(n20549),.clk(gclk));
	jnot g20250(.din(w_n19898_0[0]),.dout(n20550),.clk(gclk));
	jand g20251(.dina(w_asqrt2_20[2]),.dinb(w_n19892_0[0]),.dout(n20551),.clk(gclk));
	jand g20252(.dina(w_n20551_0[1]),.dinb(n20550),.dout(n20552),.clk(gclk));
	jor g20253(.dina(n20552),.dinb(n20549),.dout(n20553),.clk(gclk));
	jnot g20254(.din(w_n19899_0[0]),.dout(n20554),.clk(gclk));
	jand g20255(.dina(w_n20551_0[0]),.dinb(n20554),.dout(n20555),.clk(gclk));
	jnot g20256(.din(n20555),.dout(n20556),.clk(gclk));
	jand g20257(.dina(n20556),.dinb(n20553),.dout(n20557),.clk(gclk));
	jand g20258(.dina(w_n20557_0[1]),.dinb(w_n20548_0[1]),.dout(n20558),.clk(gclk));
	jor g20259(.dina(n20558),.dinb(w_n20546_0[1]),.dout(n20559),.clk(gclk));
	jand g20260(.dina(w_n20559_0[1]),.dinb(w_asqrt33_7[2]),.dout(n20560),.clk(gclk));
	jxor g20261(.dina(w_n19900_0[0]),.dinb(w_n5788_7[1]),.dout(n20561),.clk(gclk));
	jand g20262(.dina(n20561),.dinb(w_asqrt2_20[1]),.dout(n20562),.clk(gclk));
	jxor g20263(.dina(n20562),.dinb(w_n19910_0[0]),.dout(n20563),.clk(gclk));
	jnot g20264(.din(w_n20563_0[1]),.dout(n20564),.clk(gclk));
	jor g20265(.dina(w_n20559_0[0]),.dinb(w_asqrt33_7[1]),.dout(n20565),.clk(gclk));
	jand g20266(.dina(w_n20565_0[1]),.dinb(n20564),.dout(n20566),.clk(gclk));
	jor g20267(.dina(w_n20566_0[2]),.dinb(w_n20560_0[2]),.dout(n20567),.clk(gclk));
	jand g20268(.dina(n20567),.dinb(w_asqrt34_10[2]),.dout(n20568),.clk(gclk));
	jnot g20269(.din(w_n19915_0[0]),.dout(n20569),.clk(gclk));
	jand g20270(.dina(n20569),.dinb(w_n19913_0[0]),.dout(n20570),.clk(gclk));
	jand g20271(.dina(n20570),.dinb(w_asqrt2_20[0]),.dout(n20571),.clk(gclk));
	jxor g20272(.dina(n20571),.dinb(w_n19923_0[0]),.dout(n20572),.clk(gclk));
	jnot g20273(.din(w_n20572_0[1]),.dout(n20573),.clk(gclk));
	jor g20274(.dina(w_n20560_0[1]),.dinb(w_asqrt34_10[1]),.dout(n20574),.clk(gclk));
	jor g20275(.dina(n20574),.dinb(w_n20566_0[1]),.dout(n20575),.clk(gclk));
	jand g20276(.dina(w_n20575_0[1]),.dinb(n20573),.dout(n20576),.clk(gclk));
	jor g20277(.dina(w_n20576_0[1]),.dinb(w_n20568_0[1]),.dout(n20577),.clk(gclk));
	jand g20278(.dina(w_n20577_0[2]),.dinb(w_asqrt35_7[2]),.dout(n20578),.clk(gclk));
	jor g20279(.dina(w_n20577_0[1]),.dinb(w_asqrt35_7[1]),.dout(n20579),.clk(gclk));
	jnot g20280(.din(w_n19929_0[0]),.dout(n20580),.clk(gclk));
	jnot g20281(.din(w_n19930_0[0]),.dout(n20581),.clk(gclk));
	jand g20282(.dina(w_asqrt2_19[2]),.dinb(w_n19926_0[0]),.dout(n20582),.clk(gclk));
	jand g20283(.dina(w_n20582_0[1]),.dinb(n20581),.dout(n20583),.clk(gclk));
	jor g20284(.dina(n20583),.dinb(n20580),.dout(n20584),.clk(gclk));
	jnot g20285(.din(w_n19931_0[0]),.dout(n20585),.clk(gclk));
	jand g20286(.dina(w_n20582_0[0]),.dinb(n20585),.dout(n20586),.clk(gclk));
	jnot g20287(.din(n20586),.dout(n20587),.clk(gclk));
	jand g20288(.dina(n20587),.dinb(n20584),.dout(n20588),.clk(gclk));
	jand g20289(.dina(w_n20588_0[1]),.dinb(n20579),.dout(n20589),.clk(gclk));
	jor g20290(.dina(w_n20589_0[1]),.dinb(w_n20578_0[1]),.dout(n20590),.clk(gclk));
	jand g20291(.dina(n20590),.dinb(w_asqrt36_10[2]),.dout(n20591),.clk(gclk));
	jor g20292(.dina(w_n20578_0[0]),.dinb(w_asqrt36_10[1]),.dout(n20592),.clk(gclk));
	jor g20293(.dina(n20592),.dinb(w_n20589_0[0]),.dout(n20593),.clk(gclk));
	jnot g20294(.din(w_n19937_0[0]),.dout(n20594),.clk(gclk));
	jnot g20295(.din(w_n19939_0[0]),.dout(n20595),.clk(gclk));
	jand g20296(.dina(w_asqrt2_19[1]),.dinb(w_n19933_0[0]),.dout(n20596),.clk(gclk));
	jand g20297(.dina(w_n20596_0[1]),.dinb(n20595),.dout(n20597),.clk(gclk));
	jor g20298(.dina(n20597),.dinb(n20594),.dout(n20598),.clk(gclk));
	jnot g20299(.din(w_n19940_0[0]),.dout(n20599),.clk(gclk));
	jand g20300(.dina(w_n20596_0[0]),.dinb(n20599),.dout(n20600),.clk(gclk));
	jnot g20301(.din(n20600),.dout(n20601),.clk(gclk));
	jand g20302(.dina(n20601),.dinb(n20598),.dout(n20602),.clk(gclk));
	jand g20303(.dina(w_n20602_0[1]),.dinb(w_n20593_0[1]),.dout(n20603),.clk(gclk));
	jor g20304(.dina(n20603),.dinb(w_n20591_0[1]),.dout(n20604),.clk(gclk));
	jand g20305(.dina(w_n20604_0[1]),.dinb(w_asqrt37_8[0]),.dout(n20605),.clk(gclk));
	jxor g20306(.dina(w_n19941_0[0]),.dinb(w_n4494_8[1]),.dout(n20606),.clk(gclk));
	jand g20307(.dina(n20606),.dinb(w_asqrt2_19[0]),.dout(n20607),.clk(gclk));
	jxor g20308(.dina(n20607),.dinb(w_n19951_0[0]),.dout(n20608),.clk(gclk));
	jnot g20309(.din(w_n20608_0[1]),.dout(n20609),.clk(gclk));
	jor g20310(.dina(w_n20604_0[0]),.dinb(w_asqrt37_7[2]),.dout(n20610),.clk(gclk));
	jand g20311(.dina(w_n20610_0[1]),.dinb(n20609),.dout(n20611),.clk(gclk));
	jor g20312(.dina(w_n20611_0[2]),.dinb(w_n20605_0[2]),.dout(n20612),.clk(gclk));
	jand g20313(.dina(n20612),.dinb(w_asqrt38_10[2]),.dout(n20613),.clk(gclk));
	jnot g20314(.din(w_n19956_0[0]),.dout(n20614),.clk(gclk));
	jand g20315(.dina(n20614),.dinb(w_n19954_0[0]),.dout(n20615),.clk(gclk));
	jand g20316(.dina(n20615),.dinb(w_asqrt2_18[2]),.dout(n20616),.clk(gclk));
	jxor g20317(.dina(n20616),.dinb(w_n19964_0[0]),.dout(n20617),.clk(gclk));
	jnot g20318(.din(w_n20617_0[1]),.dout(n20618),.clk(gclk));
	jor g20319(.dina(w_n20605_0[1]),.dinb(w_asqrt38_10[1]),.dout(n20619),.clk(gclk));
	jor g20320(.dina(n20619),.dinb(w_n20611_0[1]),.dout(n20620),.clk(gclk));
	jand g20321(.dina(w_n20620_0[1]),.dinb(n20618),.dout(n20621),.clk(gclk));
	jor g20322(.dina(w_n20621_0[1]),.dinb(w_n20613_0[1]),.dout(n20622),.clk(gclk));
	jand g20323(.dina(w_n20622_0[2]),.dinb(w_asqrt39_8[0]),.dout(n20623),.clk(gclk));
	jor g20324(.dina(w_n20622_0[1]),.dinb(w_asqrt39_7[2]),.dout(n20624),.clk(gclk));
	jnot g20325(.din(w_n19970_0[0]),.dout(n20625),.clk(gclk));
	jnot g20326(.din(w_n19971_0[0]),.dout(n20626),.clk(gclk));
	jand g20327(.dina(w_asqrt2_18[1]),.dinb(w_n19967_0[0]),.dout(n20627),.clk(gclk));
	jand g20328(.dina(w_n20627_0[1]),.dinb(n20626),.dout(n20628),.clk(gclk));
	jor g20329(.dina(n20628),.dinb(n20625),.dout(n20629),.clk(gclk));
	jnot g20330(.din(w_n19972_0[0]),.dout(n20630),.clk(gclk));
	jand g20331(.dina(w_n20627_0[0]),.dinb(n20630),.dout(n20631),.clk(gclk));
	jnot g20332(.din(n20631),.dout(n20632),.clk(gclk));
	jand g20333(.dina(n20632),.dinb(n20629),.dout(n20633),.clk(gclk));
	jand g20334(.dina(w_n20633_0[1]),.dinb(n20624),.dout(n20634),.clk(gclk));
	jor g20335(.dina(w_n20634_0[1]),.dinb(w_n20623_0[1]),.dout(n20635),.clk(gclk));
	jand g20336(.dina(n20635),.dinb(w_asqrt40_10[2]),.dout(n20636),.clk(gclk));
	jor g20337(.dina(w_n20623_0[0]),.dinb(w_asqrt40_10[1]),.dout(n20637),.clk(gclk));
	jor g20338(.dina(n20637),.dinb(w_n20634_0[0]),.dout(n20638),.clk(gclk));
	jnot g20339(.din(w_n19978_0[0]),.dout(n20639),.clk(gclk));
	jnot g20340(.din(w_n19980_0[0]),.dout(n20640),.clk(gclk));
	jand g20341(.dina(w_asqrt2_18[0]),.dinb(w_n19974_0[0]),.dout(n20641),.clk(gclk));
	jand g20342(.dina(w_n20641_0[1]),.dinb(n20640),.dout(n20642),.clk(gclk));
	jor g20343(.dina(n20642),.dinb(n20639),.dout(n20643),.clk(gclk));
	jnot g20344(.din(w_n19981_0[0]),.dout(n20644),.clk(gclk));
	jand g20345(.dina(w_n20641_0[0]),.dinb(n20644),.dout(n20645),.clk(gclk));
	jnot g20346(.din(n20645),.dout(n20646),.clk(gclk));
	jand g20347(.dina(n20646),.dinb(n20643),.dout(n20647),.clk(gclk));
	jand g20348(.dina(w_n20647_0[1]),.dinb(w_n20638_0[1]),.dout(n20648),.clk(gclk));
	jor g20349(.dina(n20648),.dinb(w_n20636_0[1]),.dout(n20649),.clk(gclk));
	jand g20350(.dina(w_n20649_0[1]),.dinb(w_asqrt41_8[1]),.dout(n20650),.clk(gclk));
	jxor g20351(.dina(w_n19982_0[0]),.dinb(w_n3371_9[0]),.dout(n20651),.clk(gclk));
	jand g20352(.dina(n20651),.dinb(w_asqrt2_17[2]),.dout(n20652),.clk(gclk));
	jxor g20353(.dina(n20652),.dinb(w_n19992_0[0]),.dout(n20653),.clk(gclk));
	jnot g20354(.din(w_n20653_0[1]),.dout(n20654),.clk(gclk));
	jor g20355(.dina(w_n20649_0[0]),.dinb(w_asqrt41_8[0]),.dout(n20655),.clk(gclk));
	jand g20356(.dina(w_n20655_0[1]),.dinb(n20654),.dout(n20656),.clk(gclk));
	jor g20357(.dina(w_n20656_0[2]),.dinb(w_n20650_0[2]),.dout(n20657),.clk(gclk));
	jand g20358(.dina(n20657),.dinb(w_asqrt42_10[2]),.dout(n20658),.clk(gclk));
	jnot g20359(.din(w_n19997_0[0]),.dout(n20659),.clk(gclk));
	jand g20360(.dina(n20659),.dinb(w_n19995_0[0]),.dout(n20660),.clk(gclk));
	jand g20361(.dina(n20660),.dinb(w_asqrt2_17[1]),.dout(n20661),.clk(gclk));
	jxor g20362(.dina(n20661),.dinb(w_n20005_0[0]),.dout(n20662),.clk(gclk));
	jnot g20363(.din(w_n20662_0[1]),.dout(n20663),.clk(gclk));
	jor g20364(.dina(w_n20650_0[1]),.dinb(w_asqrt42_10[1]),.dout(n20664),.clk(gclk));
	jor g20365(.dina(n20664),.dinb(w_n20656_0[1]),.dout(n20665),.clk(gclk));
	jand g20366(.dina(w_n20665_0[1]),.dinb(n20663),.dout(n20666),.clk(gclk));
	jor g20367(.dina(w_n20666_0[1]),.dinb(w_n20658_0[1]),.dout(n20667),.clk(gclk));
	jand g20368(.dina(w_n20667_0[2]),.dinb(w_asqrt43_8[1]),.dout(n20668),.clk(gclk));
	jor g20369(.dina(w_n20667_0[1]),.dinb(w_asqrt43_8[0]),.dout(n20669),.clk(gclk));
	jnot g20370(.din(w_n20011_0[0]),.dout(n20670),.clk(gclk));
	jnot g20371(.din(w_n20012_0[0]),.dout(n20671),.clk(gclk));
	jand g20372(.dina(w_asqrt2_17[0]),.dinb(w_n20008_0[0]),.dout(n20672),.clk(gclk));
	jand g20373(.dina(w_n20672_0[1]),.dinb(n20671),.dout(n20673),.clk(gclk));
	jor g20374(.dina(n20673),.dinb(n20670),.dout(n20674),.clk(gclk));
	jnot g20375(.din(w_n20013_0[0]),.dout(n20675),.clk(gclk));
	jand g20376(.dina(w_n20672_0[0]),.dinb(n20675),.dout(n20676),.clk(gclk));
	jnot g20377(.din(n20676),.dout(n20677),.clk(gclk));
	jand g20378(.dina(n20677),.dinb(n20674),.dout(n20678),.clk(gclk));
	jand g20379(.dina(w_n20678_0[1]),.dinb(n20669),.dout(n20679),.clk(gclk));
	jor g20380(.dina(w_n20679_0[1]),.dinb(w_n20668_0[1]),.dout(n20680),.clk(gclk));
	jand g20381(.dina(n20680),.dinb(w_asqrt44_10[2]),.dout(n20681),.clk(gclk));
	jor g20382(.dina(w_n20668_0[0]),.dinb(w_asqrt44_10[1]),.dout(n20682),.clk(gclk));
	jor g20383(.dina(n20682),.dinb(w_n20679_0[0]),.dout(n20683),.clk(gclk));
	jnot g20384(.din(w_n20019_0[0]),.dout(n20684),.clk(gclk));
	jnot g20385(.din(w_n20021_0[0]),.dout(n20685),.clk(gclk));
	jand g20386(.dina(w_asqrt2_16[2]),.dinb(w_n20015_0[0]),.dout(n20686),.clk(gclk));
	jand g20387(.dina(w_n20686_0[1]),.dinb(n20685),.dout(n20687),.clk(gclk));
	jor g20388(.dina(n20687),.dinb(n20684),.dout(n20688),.clk(gclk));
	jnot g20389(.din(w_n20022_0[0]),.dout(n20689),.clk(gclk));
	jand g20390(.dina(w_n20686_0[0]),.dinb(n20689),.dout(n20690),.clk(gclk));
	jnot g20391(.din(n20690),.dout(n20691),.clk(gclk));
	jand g20392(.dina(n20691),.dinb(n20688),.dout(n20692),.clk(gclk));
	jand g20393(.dina(w_n20692_0[1]),.dinb(w_n20683_0[1]),.dout(n20693),.clk(gclk));
	jor g20394(.dina(n20693),.dinb(w_n20681_0[1]),.dout(n20694),.clk(gclk));
	jand g20395(.dina(w_n20694_0[1]),.dinb(w_asqrt45_8[2]),.dout(n20695),.clk(gclk));
	jxor g20396(.dina(w_n20023_0[0]),.dinb(w_n2420_10[0]),.dout(n20696),.clk(gclk));
	jand g20397(.dina(n20696),.dinb(w_asqrt2_16[1]),.dout(n20697),.clk(gclk));
	jxor g20398(.dina(n20697),.dinb(w_n20033_0[0]),.dout(n20698),.clk(gclk));
	jnot g20399(.din(w_n20698_0[1]),.dout(n20699),.clk(gclk));
	jor g20400(.dina(w_n20694_0[0]),.dinb(w_asqrt45_8[1]),.dout(n20700),.clk(gclk));
	jand g20401(.dina(w_n20700_0[1]),.dinb(n20699),.dout(n20701),.clk(gclk));
	jor g20402(.dina(w_n20701_0[2]),.dinb(w_n20695_0[2]),.dout(n20702),.clk(gclk));
	jand g20403(.dina(n20702),.dinb(w_asqrt46_10[2]),.dout(n20703),.clk(gclk));
	jnot g20404(.din(w_n20038_0[0]),.dout(n20704),.clk(gclk));
	jand g20405(.dina(n20704),.dinb(w_n20036_0[0]),.dout(n20705),.clk(gclk));
	jand g20406(.dina(n20705),.dinb(w_asqrt2_16[0]),.dout(n20706),.clk(gclk));
	jxor g20407(.dina(n20706),.dinb(w_n20046_0[0]),.dout(n20707),.clk(gclk));
	jnot g20408(.din(w_n20707_0[1]),.dout(n20708),.clk(gclk));
	jor g20409(.dina(w_n20695_0[1]),.dinb(w_asqrt46_10[1]),.dout(n20709),.clk(gclk));
	jor g20410(.dina(n20709),.dinb(w_n20701_0[1]),.dout(n20710),.clk(gclk));
	jand g20411(.dina(w_n20710_0[1]),.dinb(n20708),.dout(n20711),.clk(gclk));
	jor g20412(.dina(w_n20711_0[1]),.dinb(w_n20703_0[1]),.dout(n20712),.clk(gclk));
	jand g20413(.dina(w_n20712_0[2]),.dinb(w_asqrt47_8[2]),.dout(n20713),.clk(gclk));
	jor g20414(.dina(w_n20712_0[1]),.dinb(w_asqrt47_8[1]),.dout(n20714),.clk(gclk));
	jnot g20415(.din(w_n20052_0[0]),.dout(n20715),.clk(gclk));
	jnot g20416(.din(w_n20053_0[0]),.dout(n20716),.clk(gclk));
	jand g20417(.dina(w_asqrt2_15[2]),.dinb(w_n20049_0[0]),.dout(n20717),.clk(gclk));
	jand g20418(.dina(w_n20717_0[1]),.dinb(n20716),.dout(n20718),.clk(gclk));
	jor g20419(.dina(n20718),.dinb(n20715),.dout(n20719),.clk(gclk));
	jnot g20420(.din(w_n20054_0[0]),.dout(n20720),.clk(gclk));
	jand g20421(.dina(w_n20717_0[0]),.dinb(n20720),.dout(n20721),.clk(gclk));
	jnot g20422(.din(n20721),.dout(n20722),.clk(gclk));
	jand g20423(.dina(n20722),.dinb(n20719),.dout(n20723),.clk(gclk));
	jand g20424(.dina(w_n20723_0[1]),.dinb(n20714),.dout(n20724),.clk(gclk));
	jor g20425(.dina(w_n20724_0[1]),.dinb(w_n20713_0[1]),.dout(n20725),.clk(gclk));
	jand g20426(.dina(n20725),.dinb(w_asqrt48_10[2]),.dout(n20726),.clk(gclk));
	jor g20427(.dina(w_n20713_0[0]),.dinb(w_asqrt48_10[1]),.dout(n20727),.clk(gclk));
	jor g20428(.dina(n20727),.dinb(w_n20724_0[0]),.dout(n20728),.clk(gclk));
	jnot g20429(.din(w_n20060_0[0]),.dout(n20729),.clk(gclk));
	jnot g20430(.din(w_n20062_0[0]),.dout(n20730),.clk(gclk));
	jand g20431(.dina(w_asqrt2_15[1]),.dinb(w_n20056_0[0]),.dout(n20731),.clk(gclk));
	jand g20432(.dina(w_n20731_0[1]),.dinb(n20730),.dout(n20732),.clk(gclk));
	jor g20433(.dina(n20732),.dinb(n20729),.dout(n20733),.clk(gclk));
	jnot g20434(.din(w_n20063_0[0]),.dout(n20734),.clk(gclk));
	jand g20435(.dina(w_n20731_0[0]),.dinb(n20734),.dout(n20735),.clk(gclk));
	jnot g20436(.din(n20735),.dout(n20736),.clk(gclk));
	jand g20437(.dina(n20736),.dinb(n20733),.dout(n20737),.clk(gclk));
	jand g20438(.dina(w_n20737_0[1]),.dinb(w_n20728_0[1]),.dout(n20738),.clk(gclk));
	jor g20439(.dina(n20738),.dinb(w_n20726_0[1]),.dout(n20739),.clk(gclk));
	jand g20440(.dina(w_n20739_0[1]),.dinb(w_asqrt49_9[0]),.dout(n20740),.clk(gclk));
	jxor g20441(.dina(w_n20064_0[0]),.dinb(w_n1641_10[2]),.dout(n20741),.clk(gclk));
	jand g20442(.dina(n20741),.dinb(w_asqrt2_15[0]),.dout(n20742),.clk(gclk));
	jxor g20443(.dina(n20742),.dinb(w_n20074_0[0]),.dout(n20743),.clk(gclk));
	jnot g20444(.din(w_n20743_0[1]),.dout(n20744),.clk(gclk));
	jor g20445(.dina(w_n20739_0[0]),.dinb(w_asqrt49_8[2]),.dout(n20745),.clk(gclk));
	jand g20446(.dina(w_n20745_0[1]),.dinb(n20744),.dout(n20746),.clk(gclk));
	jor g20447(.dina(w_n20746_0[2]),.dinb(w_n20740_0[2]),.dout(n20747),.clk(gclk));
	jand g20448(.dina(n20747),.dinb(w_asqrt50_10[2]),.dout(n20748),.clk(gclk));
	jnot g20449(.din(w_n20079_0[0]),.dout(n20749),.clk(gclk));
	jand g20450(.dina(n20749),.dinb(w_n20077_0[0]),.dout(n20750),.clk(gclk));
	jand g20451(.dina(n20750),.dinb(w_asqrt2_14[2]),.dout(n20751),.clk(gclk));
	jxor g20452(.dina(n20751),.dinb(w_n20087_0[0]),.dout(n20752),.clk(gclk));
	jnot g20453(.din(w_n20752_0[1]),.dout(n20753),.clk(gclk));
	jor g20454(.dina(w_n20740_0[1]),.dinb(w_asqrt50_10[1]),.dout(n20754),.clk(gclk));
	jor g20455(.dina(n20754),.dinb(w_n20746_0[1]),.dout(n20755),.clk(gclk));
	jand g20456(.dina(w_n20755_0[1]),.dinb(n20753),.dout(n20756),.clk(gclk));
	jor g20457(.dina(w_n20756_0[1]),.dinb(w_n20748_0[1]),.dout(n20757),.clk(gclk));
	jand g20458(.dina(w_n20757_0[2]),.dinb(w_asqrt51_9[0]),.dout(n20758),.clk(gclk));
	jor g20459(.dina(w_n20757_0[1]),.dinb(w_asqrt51_8[2]),.dout(n20759),.clk(gclk));
	jnot g20460(.din(w_n20093_0[0]),.dout(n20760),.clk(gclk));
	jnot g20461(.din(w_n20094_0[0]),.dout(n20761),.clk(gclk));
	jand g20462(.dina(w_asqrt2_14[1]),.dinb(w_n20090_0[0]),.dout(n20762),.clk(gclk));
	jand g20463(.dina(w_n20762_0[1]),.dinb(n20761),.dout(n20763),.clk(gclk));
	jor g20464(.dina(n20763),.dinb(n20760),.dout(n20764),.clk(gclk));
	jnot g20465(.din(w_n20095_0[0]),.dout(n20765),.clk(gclk));
	jand g20466(.dina(w_n20762_0[0]),.dinb(n20765),.dout(n20766),.clk(gclk));
	jnot g20467(.din(n20766),.dout(n20767),.clk(gclk));
	jand g20468(.dina(n20767),.dinb(n20764),.dout(n20768),.clk(gclk));
	jand g20469(.dina(w_n20768_0[1]),.dinb(n20759),.dout(n20769),.clk(gclk));
	jor g20470(.dina(w_n20769_0[1]),.dinb(w_n20758_0[1]),.dout(n20770),.clk(gclk));
	jand g20471(.dina(n20770),.dinb(w_asqrt52_10[2]),.dout(n20771),.clk(gclk));
	jor g20472(.dina(w_n20758_0[0]),.dinb(w_asqrt52_10[1]),.dout(n20772),.clk(gclk));
	jor g20473(.dina(n20772),.dinb(w_n20769_0[0]),.dout(n20773),.clk(gclk));
	jnot g20474(.din(w_n20101_0[0]),.dout(n20774),.clk(gclk));
	jnot g20475(.din(w_n20103_0[0]),.dout(n20775),.clk(gclk));
	jand g20476(.dina(w_asqrt2_14[0]),.dinb(w_n20097_0[0]),.dout(n20776),.clk(gclk));
	jand g20477(.dina(w_n20776_0[1]),.dinb(n20775),.dout(n20777),.clk(gclk));
	jor g20478(.dina(n20777),.dinb(n20774),.dout(n20778),.clk(gclk));
	jnot g20479(.din(w_n20104_0[0]),.dout(n20779),.clk(gclk));
	jand g20480(.dina(w_n20776_0[0]),.dinb(n20779),.dout(n20780),.clk(gclk));
	jnot g20481(.din(n20780),.dout(n20781),.clk(gclk));
	jand g20482(.dina(n20781),.dinb(n20778),.dout(n20782),.clk(gclk));
	jand g20483(.dina(w_n20782_0[1]),.dinb(w_n20773_0[1]),.dout(n20783),.clk(gclk));
	jor g20484(.dina(n20783),.dinb(w_n20771_0[1]),.dout(n20784),.clk(gclk));
	jand g20485(.dina(w_n20784_0[1]),.dinb(w_asqrt53_9[1]),.dout(n20785),.clk(gclk));
	jxor g20486(.dina(w_n20105_0[0]),.dinb(w_n1034_11[2]),.dout(n20786),.clk(gclk));
	jand g20487(.dina(n20786),.dinb(w_asqrt2_13[2]),.dout(n20787),.clk(gclk));
	jxor g20488(.dina(n20787),.dinb(w_n20115_0[0]),.dout(n20788),.clk(gclk));
	jnot g20489(.din(w_n20788_0[1]),.dout(n20789),.clk(gclk));
	jor g20490(.dina(w_n20784_0[0]),.dinb(w_asqrt53_9[0]),.dout(n20790),.clk(gclk));
	jand g20491(.dina(w_n20790_0[1]),.dinb(n20789),.dout(n20791),.clk(gclk));
	jor g20492(.dina(w_n20791_0[2]),.dinb(w_n20785_0[2]),.dout(n20792),.clk(gclk));
	jand g20493(.dina(n20792),.dinb(w_asqrt54_10[2]),.dout(n20793),.clk(gclk));
	jnot g20494(.din(w_n20120_0[0]),.dout(n20794),.clk(gclk));
	jand g20495(.dina(n20794),.dinb(w_n20118_0[0]),.dout(n20795),.clk(gclk));
	jand g20496(.dina(n20795),.dinb(w_asqrt2_13[1]),.dout(n20796),.clk(gclk));
	jxor g20497(.dina(n20796),.dinb(w_n20128_0[0]),.dout(n20797),.clk(gclk));
	jnot g20498(.din(w_n20797_0[1]),.dout(n20798),.clk(gclk));
	jor g20499(.dina(w_n20785_0[1]),.dinb(w_asqrt54_10[1]),.dout(n20799),.clk(gclk));
	jor g20500(.dina(n20799),.dinb(w_n20791_0[1]),.dout(n20800),.clk(gclk));
	jand g20501(.dina(w_n20800_0[1]),.dinb(n20798),.dout(n20801),.clk(gclk));
	jor g20502(.dina(w_n20801_0[1]),.dinb(w_n20793_0[1]),.dout(n20802),.clk(gclk));
	jand g20503(.dina(w_n20802_0[2]),.dinb(w_asqrt55_9[2]),.dout(n20803),.clk(gclk));
	jor g20504(.dina(w_n20802_0[1]),.dinb(w_asqrt55_9[1]),.dout(n20804),.clk(gclk));
	jnot g20505(.din(w_n20134_0[0]),.dout(n20805),.clk(gclk));
	jnot g20506(.din(w_n20135_0[0]),.dout(n20806),.clk(gclk));
	jand g20507(.dina(w_asqrt2_13[0]),.dinb(w_n20131_0[0]),.dout(n20807),.clk(gclk));
	jand g20508(.dina(w_n20807_0[1]),.dinb(n20806),.dout(n20808),.clk(gclk));
	jor g20509(.dina(n20808),.dinb(n20805),.dout(n20809),.clk(gclk));
	jnot g20510(.din(w_n20136_0[0]),.dout(n20810),.clk(gclk));
	jand g20511(.dina(w_n20807_0[0]),.dinb(n20810),.dout(n20811),.clk(gclk));
	jnot g20512(.din(n20811),.dout(n20812),.clk(gclk));
	jand g20513(.dina(n20812),.dinb(n20809),.dout(n20813),.clk(gclk));
	jand g20514(.dina(w_n20813_0[1]),.dinb(n20804),.dout(n20814),.clk(gclk));
	jor g20515(.dina(w_n20814_0[1]),.dinb(w_n20803_0[1]),.dout(n20815),.clk(gclk));
	jand g20516(.dina(n20815),.dinb(w_asqrt56_10[2]),.dout(n20816),.clk(gclk));
	jor g20517(.dina(w_n20803_0[0]),.dinb(w_asqrt56_10[1]),.dout(n20817),.clk(gclk));
	jor g20518(.dina(n20817),.dinb(w_n20814_0[0]),.dout(n20818),.clk(gclk));
	jnot g20519(.din(w_n20142_0[0]),.dout(n20819),.clk(gclk));
	jnot g20520(.din(w_n20144_0[0]),.dout(n20820),.clk(gclk));
	jand g20521(.dina(w_asqrt2_12[2]),.dinb(w_n20138_0[0]),.dout(n20821),.clk(gclk));
	jand g20522(.dina(w_n20821_0[1]),.dinb(n20820),.dout(n20822),.clk(gclk));
	jor g20523(.dina(n20822),.dinb(n20819),.dout(n20823),.clk(gclk));
	jnot g20524(.din(w_n20145_0[0]),.dout(n20824),.clk(gclk));
	jand g20525(.dina(w_n20821_0[0]),.dinb(n20824),.dout(n20825),.clk(gclk));
	jnot g20526(.din(n20825),.dout(n20826),.clk(gclk));
	jand g20527(.dina(n20826),.dinb(n20823),.dout(n20827),.clk(gclk));
	jand g20528(.dina(w_n20827_0[1]),.dinb(w_n20818_0[1]),.dout(n20828),.clk(gclk));
	jor g20529(.dina(n20828),.dinb(w_n20816_0[1]),.dout(n20829),.clk(gclk));
	jand g20530(.dina(w_n20829_0[1]),.dinb(w_asqrt57_10[0]),.dout(n20830),.clk(gclk));
	jxor g20531(.dina(w_n20146_0[0]),.dinb(w_n590_12[1]),.dout(n20831),.clk(gclk));
	jand g20532(.dina(n20831),.dinb(w_asqrt2_12[1]),.dout(n20832),.clk(gclk));
	jxor g20533(.dina(n20832),.dinb(w_n20156_0[0]),.dout(n20833),.clk(gclk));
	jnot g20534(.din(w_n20833_0[1]),.dout(n20834),.clk(gclk));
	jor g20535(.dina(w_n20829_0[0]),.dinb(w_asqrt57_9[2]),.dout(n20835),.clk(gclk));
	jand g20536(.dina(w_n20835_0[1]),.dinb(n20834),.dout(n20836),.clk(gclk));
	jor g20537(.dina(w_n20836_0[2]),.dinb(w_n20830_0[2]),.dout(n20837),.clk(gclk));
	jand g20538(.dina(n20837),.dinb(w_asqrt58_10[2]),.dout(n20838),.clk(gclk));
	jnot g20539(.din(w_n20161_0[0]),.dout(n20839),.clk(gclk));
	jand g20540(.dina(n20839),.dinb(w_n20159_0[0]),.dout(n20840),.clk(gclk));
	jand g20541(.dina(n20840),.dinb(w_asqrt2_12[0]),.dout(n20841),.clk(gclk));
	jxor g20542(.dina(n20841),.dinb(w_n20169_0[0]),.dout(n20842),.clk(gclk));
	jnot g20543(.din(w_n20842_0[1]),.dout(n20843),.clk(gclk));
	jor g20544(.dina(w_n20830_0[1]),.dinb(w_asqrt58_10[1]),.dout(n20844),.clk(gclk));
	jor g20545(.dina(n20844),.dinb(w_n20836_0[1]),.dout(n20845),.clk(gclk));
	jand g20546(.dina(w_n20845_0[1]),.dinb(n20843),.dout(n20846),.clk(gclk));
	jor g20547(.dina(w_n20846_0[1]),.dinb(w_n20838_0[1]),.dout(n20847),.clk(gclk));
	jand g20548(.dina(w_n20847_0[2]),.dinb(w_asqrt59_10[1]),.dout(n20848),.clk(gclk));
	jor g20549(.dina(w_n20847_0[1]),.dinb(w_asqrt59_10[0]),.dout(n20849),.clk(gclk));
	jnot g20550(.din(w_n20175_0[0]),.dout(n20850),.clk(gclk));
	jnot g20551(.din(w_n20176_0[0]),.dout(n20851),.clk(gclk));
	jand g20552(.dina(w_asqrt2_11[2]),.dinb(w_n20172_0[0]),.dout(n20852),.clk(gclk));
	jand g20553(.dina(w_n20852_0[1]),.dinb(n20851),.dout(n20853),.clk(gclk));
	jor g20554(.dina(n20853),.dinb(n20850),.dout(n20854),.clk(gclk));
	jnot g20555(.din(w_n20177_0[0]),.dout(n20855),.clk(gclk));
	jand g20556(.dina(w_n20852_0[0]),.dinb(n20855),.dout(n20856),.clk(gclk));
	jnot g20557(.din(n20856),.dout(n20857),.clk(gclk));
	jand g20558(.dina(n20857),.dinb(n20854),.dout(n20858),.clk(gclk));
	jand g20559(.dina(w_n20858_0[1]),.dinb(n20849),.dout(n20859),.clk(gclk));
	jor g20560(.dina(w_n20859_0[1]),.dinb(w_n20848_0[1]),.dout(n20860),.clk(gclk));
	jand g20561(.dina(n20860),.dinb(w_asqrt60_10[1]),.dout(n20861),.clk(gclk));
	jnot g20562(.din(w_n20181_0[0]),.dout(n20862),.clk(gclk));
	jand g20563(.dina(n20862),.dinb(w_n20179_0[0]),.dout(n20863),.clk(gclk));
	jand g20564(.dina(n20863),.dinb(w_asqrt2_11[1]),.dout(n20864),.clk(gclk));
	jxor g20565(.dina(n20864),.dinb(w_n20189_0[0]),.dout(n20865),.clk(gclk));
	jnot g20566(.din(w_n20865_0[1]),.dout(n20866),.clk(gclk));
	jor g20567(.dina(w_n20848_0[0]),.dinb(w_asqrt60_10[0]),.dout(n20867),.clk(gclk));
	jor g20568(.dina(n20867),.dinb(w_n20859_0[0]),.dout(n20868),.clk(gclk));
	jand g20569(.dina(w_n20868_0[1]),.dinb(n20866),.dout(n20869),.clk(gclk));
	jor g20570(.dina(w_n20869_0[1]),.dinb(w_n20861_0[1]),.dout(n20870),.clk(gclk));
	jand g20571(.dina(w_n20870_0[2]),.dinb(w_asqrt61_10[2]),.dout(n20871),.clk(gclk));
	jor g20572(.dina(w_n20870_0[1]),.dinb(w_asqrt61_10[1]),.dout(n20872),.clk(gclk));
	jand g20573(.dina(n20872),.dinb(w_n20234_0[1]),.dout(n20873),.clk(gclk));
	jor g20574(.dina(w_n20873_0[1]),.dinb(w_n20871_0[1]),.dout(n20874),.clk(gclk));
	jand g20575(.dina(n20874),.dinb(w_asqrt62_10[2]),.dout(n20875),.clk(gclk));
	jor g20576(.dina(w_n20871_0[0]),.dinb(w_asqrt62_10[1]),.dout(n20876),.clk(gclk));
	jor g20577(.dina(n20876),.dinb(w_n20873_0[0]),.dout(n20877),.clk(gclk));
	jnot g20578(.din(w_n20200_0[0]),.dout(n20878),.clk(gclk));
	jnot g20579(.din(w_n20202_0[0]),.dout(n20879),.clk(gclk));
	jand g20580(.dina(w_asqrt2_11[0]),.dinb(w_n20196_0[0]),.dout(n20880),.clk(gclk));
	jand g20581(.dina(w_n20880_0[1]),.dinb(n20879),.dout(n20881),.clk(gclk));
	jor g20582(.dina(n20881),.dinb(n20878),.dout(n20882),.clk(gclk));
	jnot g20583(.din(w_n20203_0[0]),.dout(n20883),.clk(gclk));
	jand g20584(.dina(w_n20880_0[0]),.dinb(n20883),.dout(n20884),.clk(gclk));
	jnot g20585(.din(n20884),.dout(n20885),.clk(gclk));
	jand g20586(.dina(n20885),.dinb(n20882),.dout(n20886),.clk(gclk));
	jand g20587(.dina(w_n20886_0[1]),.dinb(w_n20877_0[1]),.dout(n20887),.clk(gclk));
	jor g20588(.dina(n20887),.dinb(w_n20875_0[1]),.dout(n20888),.clk(gclk));
	jxor g20589(.dina(w_n20204_0[0]),.dinb(w_n199_15[2]),.dout(n20889),.clk(gclk));
	jand g20590(.dina(n20889),.dinb(w_asqrt2_10[2]),.dout(n20890),.clk(gclk));
	jxor g20591(.dina(n20890),.dinb(w_n20209_0[0]),.dout(n20891),.clk(gclk));
	jnot g20592(.din(w_n20211_0[0]),.dout(n20892),.clk(gclk));
	jnot g20593(.din(w_n20215_0[0]),.dout(n20893),.clk(gclk));
	jand g20594(.dina(w_asqrt2_10[1]),.dinb(w_n20893_0[1]),.dout(n20894),.clk(gclk));
	jand g20595(.dina(w_n20894_0[1]),.dinb(w_n20892_0[2]),.dout(n20895),.clk(gclk));
	jor g20596(.dina(n20895),.dinb(w_n20223_0[0]),.dout(n20896),.clk(gclk));
	jor g20597(.dina(n20896),.dinb(w_n20891_0[2]),.dout(n20897),.clk(gclk));
	jnot g20598(.din(n20897),.dout(n20898),.clk(gclk));
	jand g20599(.dina(n20898),.dinb(w_n20888_1[2]),.dout(n20899),.clk(gclk));
	jor g20600(.dina(n20899),.dinb(w_asqrt63_6[0]),.dout(n20900),.clk(gclk));
	jnot g20601(.din(w_n20891_0[1]),.dout(n20901),.clk(gclk));
	jor g20602(.dina(w_n20901_0[1]),.dinb(w_n20888_1[1]),.dout(n20902),.clk(gclk));
	jor g20603(.dina(w_n20894_0[0]),.dinb(w_n20892_0[1]),.dout(n20903),.clk(gclk));
	jand g20604(.dina(w_n20893_0[0]),.dinb(w_n20892_0[0]),.dout(n20904),.clk(gclk));
	jor g20605(.dina(n20904),.dinb(w_n194_14[2]),.dout(n20905),.clk(gclk));
	jnot g20606(.din(n20905),.dout(n20906),.clk(gclk));
	jand g20607(.dina(n20906),.dinb(n20903),.dout(n20907),.clk(gclk));
	jnot g20608(.din(n20907),.dout(n20908),.clk(gclk));
	jand g20609(.dina(n20908),.dinb(w_n20902_0[1]),.dout(n20909),.clk(gclk));
	jand g20610(.dina(n20909),.dinb(n20900),.dout(n20910),.clk(gclk));
	jxor g20611(.dina(w_n20870_0[0]),.dinb(w_n223_13[2]),.dout(n20911),.clk(gclk));
	jor g20612(.dina(n20911),.dinb(w_n20910_17[2]),.dout(n20912),.clk(gclk));
	jxor g20613(.dina(n20912),.dinb(w_n20234_0[0]),.dout(n20913),.clk(gclk));
	jor g20614(.dina(w_n20913_0[1]),.dinb(w_n199_15[1]),.dout(n20914),.clk(gclk));
	jor g20615(.dina(a[1]),.dinb(a[0]),.dout(n20915),.clk(gclk));
	jand g20616(.dina(n20915),.dinb(w_n20236_0[0]),.dout(n20916),.clk(gclk));
	jand g20617(.dina(w_n20910_17[1]),.dinb(w_a2_0[1]),.dout(n20917),.clk(gclk));
	jor g20618(.dina(n20917),.dinb(n20916),.dout(n20918),.clk(gclk));
	jand g20619(.dina(w_n20918_0[1]),.dinb(w_n20251_1[0]),.dout(n20919),.clk(gclk));
	jor g20620(.dina(w_n20918_0[0]),.dinb(w_n20251_0[2]),.dout(n20920),.clk(gclk));
	jor g20621(.dina(w_n20910_17[0]),.dinb(w_a2_0[0]),.dout(n20921),.clk(gclk));
	jxor g20622(.dina(w_n20921_0[1]),.dinb(w_n20237_0[0]),.dout(n20922),.clk(gclk));
	jand g20623(.dina(n20922),.dinb(n20920),.dout(n20923),.clk(gclk));
	jor g20624(.dina(n20923),.dinb(n20919),.dout(n20924),.clk(gclk));
	jor g20625(.dina(w_n20924_0[1]),.dinb(w_n19616_6[2]),.dout(n20925),.clk(gclk));
	jor g20626(.dina(w_n20921_0[0]),.dinb(w_a3_0[0]),.dout(n20926),.clk(gclk));
	jnot g20627(.din(w_n20910_16[2]),.dout(asqrt_fa_2),.clk(gclk));
	jor g20628(.dina(w_asqrt1_13[1]),.dinb(w_n20251_0[1]),.dout(n20928),.clk(gclk));
	jand g20629(.dina(n20928),.dinb(n20926),.dout(n20929),.clk(gclk));
	jxor g20630(.dina(n20929),.dinb(w_n19622_0[1]),.dout(n20930),.clk(gclk));
	jand g20631(.dina(n20930),.dinb(n20925),.dout(n20931),.clk(gclk));
	jxor g20632(.dina(w_n20240_0[0]),.dinb(w_n19616_6[1]),.dout(n20932),.clk(gclk));
	jor g20633(.dina(n20932),.dinb(w_n20910_16[1]),.dout(n20933),.clk(gclk));
	jxor g20634(.dina(n20933),.dinb(w_n20243_0[0]),.dout(n20934),.clk(gclk));
	jand g20635(.dina(w_n20934_0[1]),.dinb(w_n18976_1[0]),.dout(n20935),.clk(gclk));
	jand g20636(.dina(w_n20924_0[0]),.dinb(w_n19616_6[0]),.dout(n20936),.clk(gclk));
	jor g20637(.dina(n20936),.dinb(n20935),.dout(n20937),.clk(gclk));
	jor g20638(.dina(n20937),.dinb(n20931),.dout(n20938),.clk(gclk));
	jnot g20639(.din(w_n20249_0[0]),.dout(n20939),.clk(gclk));
	jor g20640(.dina(n20939),.dinb(w_n20247_0[0]),.dout(n20940),.clk(gclk));
	jor g20641(.dina(n20940),.dinb(w_n20910_16[0]),.dout(n20941),.clk(gclk));
	jxor g20642(.dina(n20941),.dinb(w_n20254_0[0]),.dout(n20942),.clk(gclk));
	jor g20643(.dina(w_n20942_0[1]),.dinb(w_n18356_7[0]),.dout(n20943),.clk(gclk));
	jor g20644(.dina(w_n20934_0[0]),.dinb(w_n18976_0[2]),.dout(n20944),.clk(gclk));
	jand g20645(.dina(n20944),.dinb(n20943),.dout(n20945),.clk(gclk));
	jand g20646(.dina(n20945),.dinb(n20938),.dout(n20946),.clk(gclk));
	jand g20647(.dina(w_n20942_0[0]),.dinb(w_n18356_6[2]),.dout(n20947),.clk(gclk));
	jxor g20648(.dina(w_n20256_0[0]),.dinb(w_n18356_6[1]),.dout(n20948),.clk(gclk));
	jor g20649(.dina(n20948),.dinb(w_n20910_15[2]),.dout(n20949),.clk(gclk));
	jxor g20650(.dina(n20949),.dinb(w_n20262_0[0]),.dout(n20950),.clk(gclk));
	jand g20651(.dina(w_n20950_0[1]),.dinb(w_n18360_1[1]),.dout(n20951),.clk(gclk));
	jor g20652(.dina(n20951),.dinb(n20947),.dout(n20952),.clk(gclk));
	jor g20653(.dina(n20952),.dinb(n20946),.dout(n20953),.clk(gclk));
	jnot g20654(.din(w_n20272_0[0]),.dout(n20954),.clk(gclk));
	jor g20655(.dina(w_n20910_15[1]),.dinb(w_n20265_0[0]),.dout(n20955),.clk(gclk));
	jor g20656(.dina(w_n20955_0[1]),.dinb(n20954),.dout(n20956),.clk(gclk));
	jand g20657(.dina(n20956),.dinb(w_n20269_0[0]),.dout(n20957),.clk(gclk));
	jnot g20658(.din(w_n20955_0[0]),.dout(n20958),.clk(gclk));
	jand g20659(.dina(n20958),.dinb(w_n20273_0[0]),.dout(n20959),.clk(gclk));
	jor g20660(.dina(n20959),.dinb(n20957),.dout(n20960),.clk(gclk));
	jor g20661(.dina(w_n20960_0[1]),.dinb(w_n17140_7[1]),.dout(n20961),.clk(gclk));
	jor g20662(.dina(w_n20950_0[0]),.dinb(w_n18360_1[0]),.dout(n20962),.clk(gclk));
	jand g20663(.dina(n20962),.dinb(n20961),.dout(n20963),.clk(gclk));
	jand g20664(.dina(n20963),.dinb(n20953),.dout(n20964),.clk(gclk));
	jxor g20665(.dina(w_n20274_0[0]),.dinb(w_n17140_7[0]),.dout(n20965),.clk(gclk));
	jor g20666(.dina(n20965),.dinb(w_n20910_15[0]),.dout(n20966),.clk(gclk));
	jxor g20667(.dina(n20966),.dinb(w_n20280_0[0]),.dout(n20967),.clk(gclk));
	jand g20668(.dina(w_n20967_0[1]),.dinb(w_n17135_2[0]),.dout(n20968),.clk(gclk));
	jand g20669(.dina(w_n20960_0[0]),.dinb(w_n17140_6[2]),.dout(n20969),.clk(gclk));
	jor g20670(.dina(n20969),.dinb(n20968),.dout(n20970),.clk(gclk));
	jor g20671(.dina(n20970),.dinb(n20964),.dout(n20971),.clk(gclk));
	jnot g20672(.din(w_n20285_0[0]),.dout(n20972),.clk(gclk));
	jor g20673(.dina(n20972),.dinb(w_n20283_0[0]),.dout(n20973),.clk(gclk));
	jor g20674(.dina(n20973),.dinb(w_n20910_14[2]),.dout(n20974),.clk(gclk));
	jxor g20675(.dina(n20974),.dinb(w_n20294_0[0]),.dout(n20975),.clk(gclk));
	jor g20676(.dina(w_n20975_0[1]),.dinb(w_n15955_7[2]),.dout(n20976),.clk(gclk));
	jor g20677(.dina(w_n20967_0[0]),.dinb(w_n17135_1[2]),.dout(n20977),.clk(gclk));
	jand g20678(.dina(n20977),.dinb(n20976),.dout(n20978),.clk(gclk));
	jand g20679(.dina(n20978),.dinb(n20971),.dout(n20979),.clk(gclk));
	jxor g20680(.dina(w_n20296_0[0]),.dinb(w_n15955_7[1]),.dout(n20980),.clk(gclk));
	jor g20681(.dina(n20980),.dinb(w_n20910_14[1]),.dout(n20981),.clk(gclk));
	jxor g20682(.dina(n20981),.dinb(w_n20301_0[0]),.dout(n20982),.clk(gclk));
	jand g20683(.dina(w_n20982_0[1]),.dinb(w_n15950_2[1]),.dout(n20983),.clk(gclk));
	jand g20684(.dina(w_n20975_0[0]),.dinb(w_n15955_7[0]),.dout(n20984),.clk(gclk));
	jor g20685(.dina(n20984),.dinb(n20983),.dout(n20985),.clk(gclk));
	jor g20686(.dina(n20985),.dinb(n20979),.dout(n20986),.clk(gclk));
	jnot g20687(.din(w_n20311_0[0]),.dout(n20987),.clk(gclk));
	jnot g20688(.din(w_n20304_0[0]),.dout(n20988),.clk(gclk));
	jand g20689(.dina(w_asqrt1_13[0]),.dinb(n20988),.dout(n20989),.clk(gclk));
	jnot g20690(.din(w_n20989_0[1]),.dout(n20990),.clk(gclk));
	jor g20691(.dina(n20990),.dinb(n20987),.dout(n20991),.clk(gclk));
	jand g20692(.dina(n20991),.dinb(w_n20308_0[0]),.dout(n20992),.clk(gclk));
	jand g20693(.dina(w_n20989_0[0]),.dinb(w_n20312_0[0]),.dout(n20993),.clk(gclk));
	jor g20694(.dina(n20993),.dinb(n20992),.dout(n20994),.clk(gclk));
	jor g20695(.dina(w_n20994_0[1]),.dinb(w_n14821_8[0]),.dout(n20995),.clk(gclk));
	jor g20696(.dina(w_n20982_0[0]),.dinb(w_n15950_2[0]),.dout(n20996),.clk(gclk));
	jand g20697(.dina(n20996),.dinb(n20995),.dout(n20997),.clk(gclk));
	jand g20698(.dina(n20997),.dinb(n20986),.dout(n20998),.clk(gclk));
	jxor g20699(.dina(w_n20313_0[0]),.dinb(w_n14821_7[2]),.dout(n20999),.clk(gclk));
	jor g20700(.dina(n20999),.dinb(w_n20910_14[0]),.dout(n21000),.clk(gclk));
	jxor g20701(.dina(n21000),.dinb(w_n20318_0[0]),.dout(n21001),.clk(gclk));
	jand g20702(.dina(w_n21001_0[1]),.dinb(w_n14816_3[0]),.dout(n21002),.clk(gclk));
	jand g20703(.dina(w_n20994_0[0]),.dinb(w_n14821_7[1]),.dout(n21003),.clk(gclk));
	jor g20704(.dina(n21003),.dinb(n21002),.dout(n21004),.clk(gclk));
	jor g20705(.dina(n21004),.dinb(n20998),.dout(n21005),.clk(gclk));
	jnot g20706(.din(w_n20323_0[0]),.dout(n21006),.clk(gclk));
	jor g20707(.dina(n21006),.dinb(w_n20321_0[0]),.dout(n21007),.clk(gclk));
	jor g20708(.dina(n21007),.dinb(w_n20910_13[2]),.dout(n21008),.clk(gclk));
	jxor g20709(.dina(n21008),.dinb(w_n20332_0[0]),.dout(n21009),.clk(gclk));
	jor g20710(.dina(w_n21009_0[1]),.dinb(w_n13723_7[2]),.dout(n21010),.clk(gclk));
	jor g20711(.dina(w_n21001_0[0]),.dinb(w_n14816_2[2]),.dout(n21011),.clk(gclk));
	jand g20712(.dina(n21011),.dinb(n21010),.dout(n21012),.clk(gclk));
	jand g20713(.dina(n21012),.dinb(n21005),.dout(n21013),.clk(gclk));
	jnot g20714(.din(w_n20340_0[0]),.dout(n21014),.clk(gclk));
	jnot g20715(.din(w_n20335_0[0]),.dout(n21015),.clk(gclk));
	jand g20716(.dina(w_asqrt1_12[2]),.dinb(n21015),.dout(n21016),.clk(gclk));
	jnot g20717(.din(w_n21016_0[1]),.dout(n21017),.clk(gclk));
	jor g20718(.dina(n21017),.dinb(n21014),.dout(n21018),.clk(gclk));
	jand g20719(.dina(n21018),.dinb(w_n20338_0[0]),.dout(n21019),.clk(gclk));
	jand g20720(.dina(w_n21016_0[0]),.dinb(w_n20341_0[0]),.dout(n21020),.clk(gclk));
	jor g20721(.dina(n21020),.dinb(n21019),.dout(n21021),.clk(gclk));
	jand g20722(.dina(w_n21021_0[1]),.dinb(w_n13718_3[1]),.dout(n21022),.clk(gclk));
	jand g20723(.dina(w_n21009_0[0]),.dinb(w_n13723_7[1]),.dout(n21023),.clk(gclk));
	jor g20724(.dina(n21023),.dinb(n21022),.dout(n21024),.clk(gclk));
	jor g20725(.dina(n21024),.dinb(n21013),.dout(n21025),.clk(gclk));
	jnot g20726(.din(w_n20350_0[0]),.dout(n21026),.clk(gclk));
	jnot g20727(.din(w_n20343_0[0]),.dout(n21027),.clk(gclk));
	jand g20728(.dina(w_asqrt1_12[1]),.dinb(n21027),.dout(n21028),.clk(gclk));
	jnot g20729(.din(w_n21028_0[1]),.dout(n21029),.clk(gclk));
	jor g20730(.dina(n21029),.dinb(n21026),.dout(n21030),.clk(gclk));
	jand g20731(.dina(n21030),.dinb(w_n20347_0[0]),.dout(n21031),.clk(gclk));
	jand g20732(.dina(w_n21028_0[0]),.dinb(w_n20351_0[0]),.dout(n21032),.clk(gclk));
	jor g20733(.dina(n21032),.dinb(n21031),.dout(n21033),.clk(gclk));
	jor g20734(.dina(w_n21033_0[1]),.dinb(w_n12675_8[2]),.dout(n21034),.clk(gclk));
	jor g20735(.dina(w_n21021_0[0]),.dinb(w_n13718_3[0]),.dout(n21035),.clk(gclk));
	jand g20736(.dina(n21035),.dinb(n21034),.dout(n21036),.clk(gclk));
	jand g20737(.dina(n21036),.dinb(n21025),.dout(n21037),.clk(gclk));
	jxor g20738(.dina(w_n20352_0[0]),.dinb(w_n12675_8[1]),.dout(n21038),.clk(gclk));
	jor g20739(.dina(n21038),.dinb(w_n20910_13[1]),.dout(n21039),.clk(gclk));
	jxor g20740(.dina(n21039),.dinb(w_n20363_0[0]),.dout(n21040),.clk(gclk));
	jand g20741(.dina(w_n21040_0[1]),.dinb(w_n12670_3[2]),.dout(n21041),.clk(gclk));
	jand g20742(.dina(w_n21033_0[0]),.dinb(w_n12675_8[0]),.dout(n21042),.clk(gclk));
	jor g20743(.dina(n21042),.dinb(n21041),.dout(n21043),.clk(gclk));
	jor g20744(.dina(n21043),.dinb(n21037),.dout(n21044),.clk(gclk));
	jnot g20745(.din(w_n20368_0[0]),.dout(n21045),.clk(gclk));
	jor g20746(.dina(n21045),.dinb(w_n20366_0[0]),.dout(n21046),.clk(gclk));
	jor g20747(.dina(n21046),.dinb(w_n20910_13[0]),.dout(n21047),.clk(gclk));
	jxor g20748(.dina(n21047),.dinb(w_n20377_0[0]),.dout(n21048),.clk(gclk));
	jor g20749(.dina(w_n21048_0[1]),.dinb(w_n11662_8[1]),.dout(n21049),.clk(gclk));
	jor g20750(.dina(w_n21040_0[0]),.dinb(w_n12670_3[1]),.dout(n21050),.clk(gclk));
	jand g20751(.dina(n21050),.dinb(n21049),.dout(n21051),.clk(gclk));
	jand g20752(.dina(n21051),.dinb(n21044),.dout(n21052),.clk(gclk));
	jnot g20753(.din(w_n20385_0[0]),.dout(n21053),.clk(gclk));
	jnot g20754(.din(w_n20380_0[0]),.dout(n21054),.clk(gclk));
	jand g20755(.dina(w_asqrt1_12[0]),.dinb(n21054),.dout(n21055),.clk(gclk));
	jnot g20756(.din(w_n21055_0[1]),.dout(n21056),.clk(gclk));
	jor g20757(.dina(n21056),.dinb(n21053),.dout(n21057),.clk(gclk));
	jand g20758(.dina(n21057),.dinb(w_n20383_0[0]),.dout(n21058),.clk(gclk));
	jand g20759(.dina(w_n21055_0[0]),.dinb(w_n20386_0[0]),.dout(n21059),.clk(gclk));
	jor g20760(.dina(n21059),.dinb(n21058),.dout(n21060),.clk(gclk));
	jand g20761(.dina(w_n21060_0[1]),.dinb(w_n11657_4[0]),.dout(n21061),.clk(gclk));
	jand g20762(.dina(w_n21048_0[0]),.dinb(w_n11662_8[0]),.dout(n21062),.clk(gclk));
	jor g20763(.dina(n21062),.dinb(n21061),.dout(n21063),.clk(gclk));
	jor g20764(.dina(n21063),.dinb(n21052),.dout(n21064),.clk(gclk));
	jnot g20765(.din(w_n20395_0[0]),.dout(n21065),.clk(gclk));
	jnot g20766(.din(w_n20388_0[0]),.dout(n21066),.clk(gclk));
	jand g20767(.dina(w_asqrt1_11[2]),.dinb(n21066),.dout(n21067),.clk(gclk));
	jnot g20768(.din(w_n21067_0[1]),.dout(n21068),.clk(gclk));
	jor g20769(.dina(n21068),.dinb(n21065),.dout(n21069),.clk(gclk));
	jand g20770(.dina(n21069),.dinb(w_n20392_0[0]),.dout(n21070),.clk(gclk));
	jand g20771(.dina(w_n21067_0[0]),.dinb(w_n20396_0[0]),.dout(n21071),.clk(gclk));
	jor g20772(.dina(n21071),.dinb(n21070),.dout(n21072),.clk(gclk));
	jor g20773(.dina(w_n21072_0[1]),.dinb(w_n10701_9[0]),.dout(n21073),.clk(gclk));
	jor g20774(.dina(w_n21060_0[0]),.dinb(w_n11657_3[2]),.dout(n21074),.clk(gclk));
	jand g20775(.dina(n21074),.dinb(n21073),.dout(n21075),.clk(gclk));
	jand g20776(.dina(n21075),.dinb(n21064),.dout(n21076),.clk(gclk));
	jxor g20777(.dina(w_n20397_0[0]),.dinb(w_n10701_8[2]),.dout(n21077),.clk(gclk));
	jor g20778(.dina(n21077),.dinb(w_n20910_12[2]),.dout(n21078),.clk(gclk));
	jxor g20779(.dina(n21078),.dinb(w_n20408_0[0]),.dout(n21079),.clk(gclk));
	jand g20780(.dina(w_n21079_0[1]),.dinb(w_n10696_4[2]),.dout(n21080),.clk(gclk));
	jand g20781(.dina(w_n21072_0[0]),.dinb(w_n10701_8[1]),.dout(n21081),.clk(gclk));
	jor g20782(.dina(n21081),.dinb(n21080),.dout(n21082),.clk(gclk));
	jor g20783(.dina(n21082),.dinb(n21076),.dout(n21083),.clk(gclk));
	jnot g20784(.din(w_n20413_0[0]),.dout(n21084),.clk(gclk));
	jor g20785(.dina(n21084),.dinb(w_n20411_0[0]),.dout(n21085),.clk(gclk));
	jor g20786(.dina(n21085),.dinb(w_n20910_12[1]),.dout(n21086),.clk(gclk));
	jxor g20787(.dina(n21086),.dinb(w_n20422_0[0]),.dout(n21087),.clk(gclk));
	jor g20788(.dina(w_n21087_0[1]),.dinb(w_n9774_8[2]),.dout(n21088),.clk(gclk));
	jor g20789(.dina(w_n21079_0[0]),.dinb(w_n10696_4[1]),.dout(n21089),.clk(gclk));
	jand g20790(.dina(n21089),.dinb(n21088),.dout(n21090),.clk(gclk));
	jand g20791(.dina(n21090),.dinb(n21083),.dout(n21091),.clk(gclk));
	jnot g20792(.din(w_n20430_0[0]),.dout(n21092),.clk(gclk));
	jnot g20793(.din(w_n20425_0[0]),.dout(n21093),.clk(gclk));
	jand g20794(.dina(w_asqrt1_11[1]),.dinb(n21093),.dout(n21094),.clk(gclk));
	jnot g20795(.din(w_n21094_0[1]),.dout(n21095),.clk(gclk));
	jor g20796(.dina(n21095),.dinb(n21092),.dout(n21096),.clk(gclk));
	jand g20797(.dina(n21096),.dinb(w_n20428_0[0]),.dout(n21097),.clk(gclk));
	jand g20798(.dina(w_n21094_0[0]),.dinb(w_n20431_0[0]),.dout(n21098),.clk(gclk));
	jor g20799(.dina(n21098),.dinb(n21097),.dout(n21099),.clk(gclk));
	jand g20800(.dina(w_n21099_0[1]),.dinb(w_n9769_5[0]),.dout(n21100),.clk(gclk));
	jand g20801(.dina(w_n21087_0[0]),.dinb(w_n9774_8[1]),.dout(n21101),.clk(gclk));
	jor g20802(.dina(n21101),.dinb(n21100),.dout(n21102),.clk(gclk));
	jor g20803(.dina(n21102),.dinb(n21091),.dout(n21103),.clk(gclk));
	jnot g20804(.din(w_n20440_0[0]),.dout(n21104),.clk(gclk));
	jnot g20805(.din(w_n20433_0[0]),.dout(n21105),.clk(gclk));
	jand g20806(.dina(w_asqrt1_11[0]),.dinb(n21105),.dout(n21106),.clk(gclk));
	jnot g20807(.din(w_n21106_0[1]),.dout(n21107),.clk(gclk));
	jor g20808(.dina(n21107),.dinb(n21104),.dout(n21108),.clk(gclk));
	jand g20809(.dina(n21108),.dinb(w_n20437_0[0]),.dout(n21109),.clk(gclk));
	jand g20810(.dina(w_n21106_0[0]),.dinb(w_n20441_0[0]),.dout(n21110),.clk(gclk));
	jor g20811(.dina(n21110),.dinb(n21109),.dout(n21111),.clk(gclk));
	jor g20812(.dina(w_n21111_0[1]),.dinb(w_n8898_9[2]),.dout(n21112),.clk(gclk));
	jor g20813(.dina(w_n21099_0[0]),.dinb(w_n9769_4[2]),.dout(n21113),.clk(gclk));
	jand g20814(.dina(n21113),.dinb(n21112),.dout(n21114),.clk(gclk));
	jand g20815(.dina(n21114),.dinb(n21103),.dout(n21115),.clk(gclk));
	jxor g20816(.dina(w_n20442_0[0]),.dinb(w_n8898_9[1]),.dout(n21116),.clk(gclk));
	jor g20817(.dina(n21116),.dinb(w_n20910_12[0]),.dout(n21117),.clk(gclk));
	jxor g20818(.dina(n21117),.dinb(w_n20453_0[0]),.dout(n21118),.clk(gclk));
	jand g20819(.dina(w_n21118_0[1]),.dinb(w_n8893_5[1]),.dout(n21119),.clk(gclk));
	jand g20820(.dina(w_n21111_0[0]),.dinb(w_n8898_9[0]),.dout(n21120),.clk(gclk));
	jor g20821(.dina(n21120),.dinb(n21119),.dout(n21121),.clk(gclk));
	jor g20822(.dina(n21121),.dinb(n21115),.dout(n21122),.clk(gclk));
	jnot g20823(.din(w_n20458_0[0]),.dout(n21123),.clk(gclk));
	jor g20824(.dina(n21123),.dinb(w_n20456_0[0]),.dout(n21124),.clk(gclk));
	jor g20825(.dina(n21124),.dinb(w_n20910_11[2]),.dout(n21125),.clk(gclk));
	jxor g20826(.dina(n21125),.dinb(w_n20467_0[0]),.dout(n21126),.clk(gclk));
	jor g20827(.dina(w_n21126_0[1]),.dinb(w_n8058_9[1]),.dout(n21127),.clk(gclk));
	jor g20828(.dina(w_n21118_0[0]),.dinb(w_n8893_5[0]),.dout(n21128),.clk(gclk));
	jand g20829(.dina(n21128),.dinb(n21127),.dout(n21129),.clk(gclk));
	jand g20830(.dina(n21129),.dinb(n21122),.dout(n21130),.clk(gclk));
	jnot g20831(.din(w_n20475_0[0]),.dout(n21131),.clk(gclk));
	jnot g20832(.din(w_n20470_0[0]),.dout(n21132),.clk(gclk));
	jand g20833(.dina(w_asqrt1_10[2]),.dinb(n21132),.dout(n21133),.clk(gclk));
	jnot g20834(.din(w_n21133_0[1]),.dout(n21134),.clk(gclk));
	jor g20835(.dina(n21134),.dinb(n21131),.dout(n21135),.clk(gclk));
	jand g20836(.dina(n21135),.dinb(w_n20473_0[0]),.dout(n21136),.clk(gclk));
	jand g20837(.dina(w_n21133_0[0]),.dinb(w_n20476_0[0]),.dout(n21137),.clk(gclk));
	jor g20838(.dina(n21137),.dinb(n21136),.dout(n21138),.clk(gclk));
	jand g20839(.dina(w_n21138_0[1]),.dinb(w_n8053_5[2]),.dout(n21139),.clk(gclk));
	jand g20840(.dina(w_n21126_0[0]),.dinb(w_n8058_9[0]),.dout(n21140),.clk(gclk));
	jor g20841(.dina(n21140),.dinb(n21139),.dout(n21141),.clk(gclk));
	jor g20842(.dina(n21141),.dinb(n21130),.dout(n21142),.clk(gclk));
	jnot g20843(.din(w_n20485_0[0]),.dout(n21143),.clk(gclk));
	jnot g20844(.din(w_n20478_0[0]),.dout(n21144),.clk(gclk));
	jand g20845(.dina(w_asqrt1_10[1]),.dinb(n21144),.dout(n21145),.clk(gclk));
	jnot g20846(.din(w_n21145_0[1]),.dout(n21146),.clk(gclk));
	jor g20847(.dina(n21146),.dinb(n21143),.dout(n21147),.clk(gclk));
	jand g20848(.dina(n21147),.dinb(w_n20482_0[0]),.dout(n21148),.clk(gclk));
	jand g20849(.dina(w_n21145_0[0]),.dinb(w_n20486_0[0]),.dout(n21149),.clk(gclk));
	jor g20850(.dina(n21149),.dinb(n21148),.dout(n21150),.clk(gclk));
	jor g20851(.dina(w_n21150_0[1]),.dinb(w_n7265_10[0]),.dout(n21151),.clk(gclk));
	jor g20852(.dina(w_n21138_0[0]),.dinb(w_n8053_5[1]),.dout(n21152),.clk(gclk));
	jand g20853(.dina(n21152),.dinb(n21151),.dout(n21153),.clk(gclk));
	jand g20854(.dina(n21153),.dinb(n21142),.dout(n21154),.clk(gclk));
	jxor g20855(.dina(w_n20487_0[0]),.dinb(w_n7265_9[2]),.dout(n21155),.clk(gclk));
	jor g20856(.dina(n21155),.dinb(w_n20910_11[1]),.dout(n21156),.clk(gclk));
	jxor g20857(.dina(n21156),.dinb(w_n20498_0[0]),.dout(n21157),.clk(gclk));
	jand g20858(.dina(w_n21157_0[1]),.dinb(w_n7260_6[1]),.dout(n21158),.clk(gclk));
	jand g20859(.dina(w_n21150_0[0]),.dinb(w_n7265_9[1]),.dout(n21159),.clk(gclk));
	jor g20860(.dina(n21159),.dinb(n21158),.dout(n21160),.clk(gclk));
	jor g20861(.dina(n21160),.dinb(n21154),.dout(n21161),.clk(gclk));
	jnot g20862(.din(w_n20503_0[0]),.dout(n21162),.clk(gclk));
	jor g20863(.dina(n21162),.dinb(w_n20501_0[0]),.dout(n21163),.clk(gclk));
	jor g20864(.dina(n21163),.dinb(w_n20910_11[0]),.dout(n21164),.clk(gclk));
	jxor g20865(.dina(n21164),.dinb(w_n20512_0[0]),.dout(n21165),.clk(gclk));
	jor g20866(.dina(w_n21165_0[1]),.dinb(w_n6505_9[2]),.dout(n21166),.clk(gclk));
	jor g20867(.dina(w_n21157_0[0]),.dinb(w_n7260_6[0]),.dout(n21167),.clk(gclk));
	jand g20868(.dina(n21167),.dinb(n21166),.dout(n21168),.clk(gclk));
	jand g20869(.dina(n21168),.dinb(n21161),.dout(n21169),.clk(gclk));
	jnot g20870(.din(w_n20520_0[0]),.dout(n21170),.clk(gclk));
	jnot g20871(.din(w_n20515_0[0]),.dout(n21171),.clk(gclk));
	jand g20872(.dina(w_asqrt1_10[0]),.dinb(n21171),.dout(n21172),.clk(gclk));
	jnot g20873(.din(w_n21172_0[1]),.dout(n21173),.clk(gclk));
	jor g20874(.dina(n21173),.dinb(n21170),.dout(n21174),.clk(gclk));
	jand g20875(.dina(n21174),.dinb(w_n20518_0[0]),.dout(n21175),.clk(gclk));
	jand g20876(.dina(w_n21172_0[0]),.dinb(w_n20521_0[0]),.dout(n21176),.clk(gclk));
	jor g20877(.dina(n21176),.dinb(n21175),.dout(n21177),.clk(gclk));
	jand g20878(.dina(w_n21177_0[1]),.dinb(w_n6500_6[2]),.dout(n21178),.clk(gclk));
	jand g20879(.dina(w_n21165_0[0]),.dinb(w_n6505_9[1]),.dout(n21179),.clk(gclk));
	jor g20880(.dina(n21179),.dinb(n21178),.dout(n21180),.clk(gclk));
	jor g20881(.dina(n21180),.dinb(n21169),.dout(n21181),.clk(gclk));
	jnot g20882(.din(w_n20530_0[0]),.dout(n21182),.clk(gclk));
	jnot g20883(.din(w_n20523_0[0]),.dout(n21183),.clk(gclk));
	jand g20884(.dina(w_asqrt1_9[2]),.dinb(n21183),.dout(n21184),.clk(gclk));
	jnot g20885(.din(w_n21184_0[1]),.dout(n21185),.clk(gclk));
	jor g20886(.dina(n21185),.dinb(n21182),.dout(n21186),.clk(gclk));
	jand g20887(.dina(n21186),.dinb(w_n20527_0[0]),.dout(n21187),.clk(gclk));
	jand g20888(.dina(w_n21184_0[0]),.dinb(w_n20531_0[0]),.dout(n21188),.clk(gclk));
	jor g20889(.dina(n21188),.dinb(n21187),.dout(n21189),.clk(gclk));
	jor g20890(.dina(w_n21189_0[1]),.dinb(w_n5793_10[1]),.dout(n21190),.clk(gclk));
	jor g20891(.dina(w_n21177_0[0]),.dinb(w_n6500_6[1]),.dout(n21191),.clk(gclk));
	jand g20892(.dina(n21191),.dinb(n21190),.dout(n21192),.clk(gclk));
	jand g20893(.dina(n21192),.dinb(n21181),.dout(n21193),.clk(gclk));
	jxor g20894(.dina(w_n20532_0[0]),.dinb(w_n5793_10[0]),.dout(n21194),.clk(gclk));
	jor g20895(.dina(n21194),.dinb(w_n20910_10[2]),.dout(n21195),.clk(gclk));
	jxor g20896(.dina(n21195),.dinb(w_n20543_0[0]),.dout(n21196),.clk(gclk));
	jand g20897(.dina(w_n21196_0[1]),.dinb(w_n5788_7[0]),.dout(n21197),.clk(gclk));
	jand g20898(.dina(w_n21189_0[0]),.dinb(w_n5793_9[2]),.dout(n21198),.clk(gclk));
	jor g20899(.dina(n21198),.dinb(n21197),.dout(n21199),.clk(gclk));
	jor g20900(.dina(n21199),.dinb(n21193),.dout(n21200),.clk(gclk));
	jnot g20901(.din(w_n20548_0[0]),.dout(n21201),.clk(gclk));
	jor g20902(.dina(n21201),.dinb(w_n20546_0[0]),.dout(n21202),.clk(gclk));
	jor g20903(.dina(n21202),.dinb(w_n20910_10[1]),.dout(n21203),.clk(gclk));
	jxor g20904(.dina(n21203),.dinb(w_n20557_0[0]),.dout(n21204),.clk(gclk));
	jor g20905(.dina(w_n21204_0[1]),.dinb(w_n5121_10[0]),.dout(n21205),.clk(gclk));
	jor g20906(.dina(w_n21196_0[0]),.dinb(w_n5788_6[2]),.dout(n21206),.clk(gclk));
	jand g20907(.dina(n21206),.dinb(n21205),.dout(n21207),.clk(gclk));
	jand g20908(.dina(n21207),.dinb(n21200),.dout(n21208),.clk(gclk));
	jnot g20909(.din(w_n20565_0[0]),.dout(n21209),.clk(gclk));
	jnot g20910(.din(w_n20560_0[0]),.dout(n21210),.clk(gclk));
	jand g20911(.dina(w_asqrt1_9[1]),.dinb(n21210),.dout(n21211),.clk(gclk));
	jnot g20912(.din(w_n21211_0[1]),.dout(n21212),.clk(gclk));
	jor g20913(.dina(n21212),.dinb(n21209),.dout(n21213),.clk(gclk));
	jand g20914(.dina(n21213),.dinb(w_n20563_0[0]),.dout(n21214),.clk(gclk));
	jand g20915(.dina(w_n21211_0[0]),.dinb(w_n20566_0[0]),.dout(n21215),.clk(gclk));
	jor g20916(.dina(n21215),.dinb(n21214),.dout(n21216),.clk(gclk));
	jand g20917(.dina(w_n21216_0[1]),.dinb(w_n5116_7[1]),.dout(n21217),.clk(gclk));
	jand g20918(.dina(w_n21204_0[0]),.dinb(w_n5121_9[2]),.dout(n21218),.clk(gclk));
	jor g20919(.dina(n21218),.dinb(n21217),.dout(n21219),.clk(gclk));
	jor g20920(.dina(n21219),.dinb(n21208),.dout(n21220),.clk(gclk));
	jnot g20921(.din(w_n20575_0[0]),.dout(n21221),.clk(gclk));
	jnot g20922(.din(w_n20568_0[0]),.dout(n21222),.clk(gclk));
	jand g20923(.dina(w_asqrt1_9[0]),.dinb(n21222),.dout(n21223),.clk(gclk));
	jnot g20924(.din(w_n21223_0[1]),.dout(n21224),.clk(gclk));
	jor g20925(.dina(n21224),.dinb(n21221),.dout(n21225),.clk(gclk));
	jand g20926(.dina(n21225),.dinb(w_n20572_0[0]),.dout(n21226),.clk(gclk));
	jand g20927(.dina(w_n21223_0[0]),.dinb(w_n20576_0[0]),.dout(n21227),.clk(gclk));
	jor g20928(.dina(n21227),.dinb(n21226),.dout(n21228),.clk(gclk));
	jor g20929(.dina(w_n21228_0[1]),.dinb(w_n4499_11[0]),.dout(n21229),.clk(gclk));
	jor g20930(.dina(w_n21216_0[0]),.dinb(w_n5116_7[0]),.dout(n21230),.clk(gclk));
	jand g20931(.dina(n21230),.dinb(n21229),.dout(n21231),.clk(gclk));
	jand g20932(.dina(n21231),.dinb(n21220),.dout(n21232),.clk(gclk));
	jxor g20933(.dina(w_n20577_0[0]),.dinb(w_n4499_10[2]),.dout(n21233),.clk(gclk));
	jor g20934(.dina(n21233),.dinb(w_n20910_10[0]),.dout(n21234),.clk(gclk));
	jxor g20935(.dina(n21234),.dinb(w_n20588_0[0]),.dout(n21235),.clk(gclk));
	jand g20936(.dina(w_n21235_0[1]),.dinb(w_n4494_8[0]),.dout(n21236),.clk(gclk));
	jand g20937(.dina(w_n21228_0[0]),.dinb(w_n4499_10[1]),.dout(n21237),.clk(gclk));
	jor g20938(.dina(n21237),.dinb(n21236),.dout(n21238),.clk(gclk));
	jor g20939(.dina(n21238),.dinb(n21232),.dout(n21239),.clk(gclk));
	jnot g20940(.din(w_n20593_0[0]),.dout(n21240),.clk(gclk));
	jor g20941(.dina(n21240),.dinb(w_n20591_0[0]),.dout(n21241),.clk(gclk));
	jor g20942(.dina(n21241),.dinb(w_n20910_9[2]),.dout(n21242),.clk(gclk));
	jxor g20943(.dina(n21242),.dinb(w_n20602_0[0]),.dout(n21243),.clk(gclk));
	jor g20944(.dina(w_n21243_0[1]),.dinb(w_n3912_10[2]),.dout(n21244),.clk(gclk));
	jor g20945(.dina(w_n21235_0[0]),.dinb(w_n4494_7[2]),.dout(n21245),.clk(gclk));
	jand g20946(.dina(n21245),.dinb(n21244),.dout(n21246),.clk(gclk));
	jand g20947(.dina(n21246),.dinb(n21239),.dout(n21247),.clk(gclk));
	jnot g20948(.din(w_n20610_0[0]),.dout(n21248),.clk(gclk));
	jnot g20949(.din(w_n20605_0[0]),.dout(n21249),.clk(gclk));
	jand g20950(.dina(w_asqrt1_8[2]),.dinb(n21249),.dout(n21250),.clk(gclk));
	jnot g20951(.din(w_n21250_0[1]),.dout(n21251),.clk(gclk));
	jor g20952(.dina(n21251),.dinb(n21248),.dout(n21252),.clk(gclk));
	jand g20953(.dina(n21252),.dinb(w_n20608_0[0]),.dout(n21253),.clk(gclk));
	jand g20954(.dina(w_n21250_0[0]),.dinb(w_n20611_0[0]),.dout(n21254),.clk(gclk));
	jor g20955(.dina(n21254),.dinb(n21253),.dout(n21255),.clk(gclk));
	jand g20956(.dina(w_n21255_0[1]),.dinb(w_n3907_8[1]),.dout(n21256),.clk(gclk));
	jand g20957(.dina(w_n21243_0[0]),.dinb(w_n3912_10[1]),.dout(n21257),.clk(gclk));
	jor g20958(.dina(n21257),.dinb(n21256),.dout(n21258),.clk(gclk));
	jor g20959(.dina(n21258),.dinb(n21247),.dout(n21259),.clk(gclk));
	jnot g20960(.din(w_n20620_0[0]),.dout(n21260),.clk(gclk));
	jnot g20961(.din(w_n20613_0[0]),.dout(n21261),.clk(gclk));
	jand g20962(.dina(w_asqrt1_8[1]),.dinb(n21261),.dout(n21262),.clk(gclk));
	jnot g20963(.din(w_n21262_0[1]),.dout(n21263),.clk(gclk));
	jor g20964(.dina(n21263),.dinb(n21260),.dout(n21264),.clk(gclk));
	jand g20965(.dina(n21264),.dinb(w_n20617_0[0]),.dout(n21265),.clk(gclk));
	jand g20966(.dina(w_n21262_0[0]),.dinb(w_n20621_0[0]),.dout(n21266),.clk(gclk));
	jor g20967(.dina(n21266),.dinb(n21265),.dout(n21267),.clk(gclk));
	jor g20968(.dina(w_n21267_0[1]),.dinb(w_n3376_11[2]),.dout(n21268),.clk(gclk));
	jor g20969(.dina(w_n21255_0[0]),.dinb(w_n3907_8[0]),.dout(n21269),.clk(gclk));
	jand g20970(.dina(n21269),.dinb(n21268),.dout(n21270),.clk(gclk));
	jand g20971(.dina(n21270),.dinb(n21259),.dout(n21271),.clk(gclk));
	jxor g20972(.dina(w_n20622_0[0]),.dinb(w_n3376_11[1]),.dout(n21272),.clk(gclk));
	jor g20973(.dina(n21272),.dinb(w_n20910_9[1]),.dout(n21273),.clk(gclk));
	jxor g20974(.dina(n21273),.dinb(w_n20633_0[0]),.dout(n21274),.clk(gclk));
	jand g20975(.dina(w_n21274_0[1]),.dinb(w_n3371_8[2]),.dout(n21275),.clk(gclk));
	jand g20976(.dina(w_n21267_0[0]),.dinb(w_n3376_11[0]),.dout(n21276),.clk(gclk));
	jor g20977(.dina(n21276),.dinb(n21275),.dout(n21277),.clk(gclk));
	jor g20978(.dina(n21277),.dinb(n21271),.dout(n21278),.clk(gclk));
	jnot g20979(.din(w_n20638_0[0]),.dout(n21279),.clk(gclk));
	jor g20980(.dina(n21279),.dinb(w_n20636_0[0]),.dout(n21280),.clk(gclk));
	jor g20981(.dina(n21280),.dinb(w_n20910_9[0]),.dout(n21281),.clk(gclk));
	jxor g20982(.dina(n21281),.dinb(w_n20647_0[0]),.dout(n21282),.clk(gclk));
	jor g20983(.dina(w_n21282_0[1]),.dinb(w_n2875_11[1]),.dout(n21283),.clk(gclk));
	jor g20984(.dina(w_n21274_0[0]),.dinb(w_n3371_8[1]),.dout(n21284),.clk(gclk));
	jand g20985(.dina(n21284),.dinb(n21283),.dout(n21285),.clk(gclk));
	jand g20986(.dina(n21285),.dinb(n21278),.dout(n21286),.clk(gclk));
	jnot g20987(.din(w_n20655_0[0]),.dout(n21287),.clk(gclk));
	jnot g20988(.din(w_n20650_0[0]),.dout(n21288),.clk(gclk));
	jand g20989(.dina(w_asqrt1_8[0]),.dinb(n21288),.dout(n21289),.clk(gclk));
	jnot g20990(.din(w_n21289_0[1]),.dout(n21290),.clk(gclk));
	jor g20991(.dina(n21290),.dinb(n21287),.dout(n21291),.clk(gclk));
	jand g20992(.dina(n21291),.dinb(w_n20653_0[0]),.dout(n21292),.clk(gclk));
	jand g20993(.dina(w_n21289_0[0]),.dinb(w_n20656_0[0]),.dout(n21293),.clk(gclk));
	jor g20994(.dina(n21293),.dinb(n21292),.dout(n21294),.clk(gclk));
	jand g20995(.dina(w_n21294_0[1]),.dinb(w_n2870_9[0]),.dout(n21295),.clk(gclk));
	jand g20996(.dina(w_n21282_0[0]),.dinb(w_n2875_11[0]),.dout(n21296),.clk(gclk));
	jor g20997(.dina(n21296),.dinb(n21295),.dout(n21297),.clk(gclk));
	jor g20998(.dina(n21297),.dinb(n21286),.dout(n21298),.clk(gclk));
	jnot g20999(.din(w_n20665_0[0]),.dout(n21299),.clk(gclk));
	jnot g21000(.din(w_n20658_0[0]),.dout(n21300),.clk(gclk));
	jand g21001(.dina(w_asqrt1_7[2]),.dinb(n21300),.dout(n21301),.clk(gclk));
	jnot g21002(.din(w_n21301_0[1]),.dout(n21302),.clk(gclk));
	jor g21003(.dina(n21302),.dinb(n21299),.dout(n21303),.clk(gclk));
	jand g21004(.dina(n21303),.dinb(w_n20662_0[0]),.dout(n21304),.clk(gclk));
	jand g21005(.dina(w_n21301_0[0]),.dinb(w_n20666_0[0]),.dout(n21305),.clk(gclk));
	jor g21006(.dina(n21305),.dinb(n21304),.dout(n21306),.clk(gclk));
	jor g21007(.dina(w_n21306_0[1]),.dinb(w_n2425_12[0]),.dout(n21307),.clk(gclk));
	jor g21008(.dina(w_n21294_0[0]),.dinb(w_n2870_8[2]),.dout(n21308),.clk(gclk));
	jand g21009(.dina(n21308),.dinb(n21307),.dout(n21309),.clk(gclk));
	jand g21010(.dina(n21309),.dinb(n21298),.dout(n21310),.clk(gclk));
	jxor g21011(.dina(w_n20667_0[0]),.dinb(w_n2425_11[2]),.dout(n21311),.clk(gclk));
	jor g21012(.dina(n21311),.dinb(w_n20910_8[2]),.dout(n21312),.clk(gclk));
	jxor g21013(.dina(n21312),.dinb(w_n20678_0[0]),.dout(n21313),.clk(gclk));
	jand g21014(.dina(w_n21313_0[1]),.dinb(w_n2420_9[2]),.dout(n21314),.clk(gclk));
	jand g21015(.dina(w_n21306_0[0]),.dinb(w_n2425_11[1]),.dout(n21315),.clk(gclk));
	jor g21016(.dina(n21315),.dinb(n21314),.dout(n21316),.clk(gclk));
	jor g21017(.dina(n21316),.dinb(n21310),.dout(n21317),.clk(gclk));
	jnot g21018(.din(w_n20683_0[0]),.dout(n21318),.clk(gclk));
	jor g21019(.dina(n21318),.dinb(w_n20681_0[0]),.dout(n21319),.clk(gclk));
	jor g21020(.dina(n21319),.dinb(w_n20910_8[1]),.dout(n21320),.clk(gclk));
	jxor g21021(.dina(n21320),.dinb(w_n20692_0[0]),.dout(n21321),.clk(gclk));
	jor g21022(.dina(w_n21321_0[1]),.dinb(w_n2010_11[2]),.dout(n21322),.clk(gclk));
	jor g21023(.dina(w_n21313_0[0]),.dinb(w_n2420_9[1]),.dout(n21323),.clk(gclk));
	jand g21024(.dina(n21323),.dinb(n21322),.dout(n21324),.clk(gclk));
	jand g21025(.dina(n21324),.dinb(n21317),.dout(n21325),.clk(gclk));
	jnot g21026(.din(w_n20700_0[0]),.dout(n21326),.clk(gclk));
	jnot g21027(.din(w_n20695_0[0]),.dout(n21327),.clk(gclk));
	jand g21028(.dina(w_asqrt1_7[1]),.dinb(n21327),.dout(n21328),.clk(gclk));
	jnot g21029(.din(w_n21328_0[1]),.dout(n21329),.clk(gclk));
	jor g21030(.dina(n21329),.dinb(n21326),.dout(n21330),.clk(gclk));
	jand g21031(.dina(n21330),.dinb(w_n20698_0[0]),.dout(n21331),.clk(gclk));
	jand g21032(.dina(w_n21328_0[0]),.dinb(w_n20701_0[0]),.dout(n21332),.clk(gclk));
	jor g21033(.dina(n21332),.dinb(n21331),.dout(n21333),.clk(gclk));
	jand g21034(.dina(w_n21333_0[1]),.dinb(w_n2005_10[0]),.dout(n21334),.clk(gclk));
	jand g21035(.dina(w_n21321_0[0]),.dinb(w_n2010_11[1]),.dout(n21335),.clk(gclk));
	jor g21036(.dina(n21335),.dinb(n21334),.dout(n21336),.clk(gclk));
	jor g21037(.dina(n21336),.dinb(n21325),.dout(n21337),.clk(gclk));
	jnot g21038(.din(w_n20710_0[0]),.dout(n21338),.clk(gclk));
	jnot g21039(.din(w_n20703_0[0]),.dout(n21339),.clk(gclk));
	jand g21040(.dina(w_asqrt1_7[0]),.dinb(n21339),.dout(n21340),.clk(gclk));
	jnot g21041(.din(w_n21340_0[1]),.dout(n21341),.clk(gclk));
	jor g21042(.dina(n21341),.dinb(n21338),.dout(n21342),.clk(gclk));
	jand g21043(.dina(n21342),.dinb(w_n20707_0[0]),.dout(n21343),.clk(gclk));
	jand g21044(.dina(w_n21340_0[0]),.dinb(w_n20711_0[0]),.dout(n21344),.clk(gclk));
	jor g21045(.dina(n21344),.dinb(n21343),.dout(n21345),.clk(gclk));
	jor g21046(.dina(w_n21345_0[1]),.dinb(w_n1646_12[2]),.dout(n21346),.clk(gclk));
	jor g21047(.dina(w_n21333_0[0]),.dinb(w_n2005_9[2]),.dout(n21347),.clk(gclk));
	jand g21048(.dina(n21347),.dinb(n21346),.dout(n21348),.clk(gclk));
	jand g21049(.dina(n21348),.dinb(n21337),.dout(n21349),.clk(gclk));
	jxor g21050(.dina(w_n20712_0[0]),.dinb(w_n1646_12[1]),.dout(n21350),.clk(gclk));
	jor g21051(.dina(n21350),.dinb(w_n20910_8[0]),.dout(n21351),.clk(gclk));
	jxor g21052(.dina(n21351),.dinb(w_n20723_0[0]),.dout(n21352),.clk(gclk));
	jand g21053(.dina(w_n21352_0[1]),.dinb(w_n1641_10[1]),.dout(n21353),.clk(gclk));
	jand g21054(.dina(w_n21345_0[0]),.dinb(w_n1646_12[0]),.dout(n21354),.clk(gclk));
	jor g21055(.dina(n21354),.dinb(n21353),.dout(n21355),.clk(gclk));
	jor g21056(.dina(n21355),.dinb(n21349),.dout(n21356),.clk(gclk));
	jnot g21057(.din(w_n20728_0[0]),.dout(n21357),.clk(gclk));
	jor g21058(.dina(n21357),.dinb(w_n20726_0[0]),.dout(n21358),.clk(gclk));
	jor g21059(.dina(n21358),.dinb(w_n20910_7[2]),.dout(n21359),.clk(gclk));
	jxor g21060(.dina(n21359),.dinb(w_n20737_0[0]),.dout(n21360),.clk(gclk));
	jor g21061(.dina(w_n21360_0[1]),.dinb(w_n1317_12[1]),.dout(n21361),.clk(gclk));
	jor g21062(.dina(w_n21352_0[0]),.dinb(w_n1641_10[0]),.dout(n21362),.clk(gclk));
	jand g21063(.dina(n21362),.dinb(n21361),.dout(n21363),.clk(gclk));
	jand g21064(.dina(n21363),.dinb(n21356),.dout(n21364),.clk(gclk));
	jnot g21065(.din(w_n20745_0[0]),.dout(n21365),.clk(gclk));
	jnot g21066(.din(w_n20740_0[0]),.dout(n21366),.clk(gclk));
	jand g21067(.dina(w_asqrt1_6[2]),.dinb(n21366),.dout(n21367),.clk(gclk));
	jnot g21068(.din(w_n21367_0[1]),.dout(n21368),.clk(gclk));
	jor g21069(.dina(n21368),.dinb(n21365),.dout(n21369),.clk(gclk));
	jand g21070(.dina(n21369),.dinb(w_n20743_0[0]),.dout(n21370),.clk(gclk));
	jand g21071(.dina(w_n21367_0[0]),.dinb(w_n20746_0[0]),.dout(n21371),.clk(gclk));
	jor g21072(.dina(n21371),.dinb(n21370),.dout(n21372),.clk(gclk));
	jand g21073(.dina(w_n21372_0[1]),.dinb(w_n1312_10[2]),.dout(n21373),.clk(gclk));
	jand g21074(.dina(w_n21360_0[0]),.dinb(w_n1317_12[0]),.dout(n21374),.clk(gclk));
	jor g21075(.dina(n21374),.dinb(n21373),.dout(n21375),.clk(gclk));
	jor g21076(.dina(n21375),.dinb(n21364),.dout(n21376),.clk(gclk));
	jnot g21077(.din(w_n20755_0[0]),.dout(n21377),.clk(gclk));
	jnot g21078(.din(w_n20748_0[0]),.dout(n21378),.clk(gclk));
	jand g21079(.dina(w_asqrt1_6[1]),.dinb(n21378),.dout(n21379),.clk(gclk));
	jnot g21080(.din(w_n21379_0[1]),.dout(n21380),.clk(gclk));
	jor g21081(.dina(n21380),.dinb(n21377),.dout(n21381),.clk(gclk));
	jand g21082(.dina(n21381),.dinb(w_n20752_0[0]),.dout(n21382),.clk(gclk));
	jand g21083(.dina(w_n21379_0[0]),.dinb(w_n20756_0[0]),.dout(n21383),.clk(gclk));
	jor g21084(.dina(n21383),.dinb(n21382),.dout(n21384),.clk(gclk));
	jor g21085(.dina(w_n21384_0[1]),.dinb(w_n1039_13[0]),.dout(n21385),.clk(gclk));
	jor g21086(.dina(w_n21372_0[0]),.dinb(w_n1312_10[1]),.dout(n21386),.clk(gclk));
	jand g21087(.dina(n21386),.dinb(n21385),.dout(n21387),.clk(gclk));
	jand g21088(.dina(n21387),.dinb(n21376),.dout(n21388),.clk(gclk));
	jxor g21089(.dina(w_n20757_0[0]),.dinb(w_n1039_12[2]),.dout(n21389),.clk(gclk));
	jor g21090(.dina(n21389),.dinb(w_n20910_7[1]),.dout(n21390),.clk(gclk));
	jxor g21091(.dina(n21390),.dinb(w_n20768_0[0]),.dout(n21391),.clk(gclk));
	jand g21092(.dina(w_n21391_0[1]),.dinb(w_n1034_11[1]),.dout(n21392),.clk(gclk));
	jand g21093(.dina(w_n21384_0[0]),.dinb(w_n1039_12[1]),.dout(n21393),.clk(gclk));
	jor g21094(.dina(n21393),.dinb(n21392),.dout(n21394),.clk(gclk));
	jor g21095(.dina(n21394),.dinb(n21388),.dout(n21395),.clk(gclk));
	jnot g21096(.din(w_n20773_0[0]),.dout(n21396),.clk(gclk));
	jor g21097(.dina(n21396),.dinb(w_n20771_0[0]),.dout(n21397),.clk(gclk));
	jor g21098(.dina(n21397),.dinb(w_n20910_7[0]),.dout(n21398),.clk(gclk));
	jxor g21099(.dina(n21398),.dinb(w_n20782_0[0]),.dout(n21399),.clk(gclk));
	jor g21100(.dina(w_n21399_0[1]),.dinb(w_n796_12[2]),.dout(n21400),.clk(gclk));
	jor g21101(.dina(w_n21391_0[0]),.dinb(w_n1034_11[0]),.dout(n21401),.clk(gclk));
	jand g21102(.dina(n21401),.dinb(n21400),.dout(n21402),.clk(gclk));
	jand g21103(.dina(n21402),.dinb(n21395),.dout(n21403),.clk(gclk));
	jnot g21104(.din(w_n20790_0[0]),.dout(n21404),.clk(gclk));
	jnot g21105(.din(w_n20785_0[0]),.dout(n21405),.clk(gclk));
	jand g21106(.dina(w_asqrt1_6[0]),.dinb(n21405),.dout(n21406),.clk(gclk));
	jnot g21107(.din(w_n21406_0[1]),.dout(n21407),.clk(gclk));
	jor g21108(.dina(n21407),.dinb(n21404),.dout(n21408),.clk(gclk));
	jand g21109(.dina(n21408),.dinb(w_n20788_0[0]),.dout(n21409),.clk(gclk));
	jand g21110(.dina(w_n21406_0[0]),.dinb(w_n20791_0[0]),.dout(n21410),.clk(gclk));
	jor g21111(.dina(n21410),.dinb(n21409),.dout(n21411),.clk(gclk));
	jand g21112(.dina(w_n21411_0[1]),.dinb(w_n791_11[2]),.dout(n21412),.clk(gclk));
	jand g21113(.dina(w_n21399_0[0]),.dinb(w_n796_12[1]),.dout(n21413),.clk(gclk));
	jor g21114(.dina(n21413),.dinb(n21412),.dout(n21414),.clk(gclk));
	jor g21115(.dina(n21414),.dinb(n21403),.dout(n21415),.clk(gclk));
	jnot g21116(.din(w_n20800_0[0]),.dout(n21416),.clk(gclk));
	jnot g21117(.din(w_n20793_0[0]),.dout(n21417),.clk(gclk));
	jand g21118(.dina(w_asqrt1_5[2]),.dinb(n21417),.dout(n21418),.clk(gclk));
	jnot g21119(.din(w_n21418_0[1]),.dout(n21419),.clk(gclk));
	jor g21120(.dina(n21419),.dinb(n21416),.dout(n21420),.clk(gclk));
	jand g21121(.dina(n21420),.dinb(w_n20797_0[0]),.dout(n21421),.clk(gclk));
	jand g21122(.dina(w_n21418_0[0]),.dinb(w_n20801_0[0]),.dout(n21422),.clk(gclk));
	jor g21123(.dina(n21422),.dinb(n21421),.dout(n21423),.clk(gclk));
	jor g21124(.dina(w_n21423_0[1]),.dinb(w_n595_13[1]),.dout(n21424),.clk(gclk));
	jor g21125(.dina(w_n21411_0[0]),.dinb(w_n791_11[1]),.dout(n21425),.clk(gclk));
	jand g21126(.dina(n21425),.dinb(n21424),.dout(n21426),.clk(gclk));
	jand g21127(.dina(n21426),.dinb(n21415),.dout(n21427),.clk(gclk));
	jxor g21128(.dina(w_n20802_0[0]),.dinb(w_n595_13[0]),.dout(n21428),.clk(gclk));
	jor g21129(.dina(n21428),.dinb(w_n20910_6[2]),.dout(n21429),.clk(gclk));
	jxor g21130(.dina(n21429),.dinb(w_n20813_0[0]),.dout(n21430),.clk(gclk));
	jand g21131(.dina(w_n21430_0[1]),.dinb(w_n590_12[0]),.dout(n21431),.clk(gclk));
	jand g21132(.dina(w_n21423_0[0]),.dinb(w_n595_12[2]),.dout(n21432),.clk(gclk));
	jor g21133(.dina(n21432),.dinb(n21431),.dout(n21433),.clk(gclk));
	jor g21134(.dina(n21433),.dinb(n21427),.dout(n21434),.clk(gclk));
	jnot g21135(.din(w_n20818_0[0]),.dout(n21435),.clk(gclk));
	jor g21136(.dina(n21435),.dinb(w_n20816_0[0]),.dout(n21436),.clk(gclk));
	jor g21137(.dina(n21436),.dinb(w_n20910_6[1]),.dout(n21437),.clk(gclk));
	jxor g21138(.dina(n21437),.dinb(w_n20827_0[0]),.dout(n21438),.clk(gclk));
	jor g21139(.dina(w_n21438_0[1]),.dinb(w_n430_13[0]),.dout(n21439),.clk(gclk));
	jor g21140(.dina(w_n21430_0[0]),.dinb(w_n590_11[2]),.dout(n21440),.clk(gclk));
	jand g21141(.dina(n21440),.dinb(n21439),.dout(n21441),.clk(gclk));
	jand g21142(.dina(n21441),.dinb(n21434),.dout(n21442),.clk(gclk));
	jnot g21143(.din(w_n20835_0[0]),.dout(n21443),.clk(gclk));
	jnot g21144(.din(w_n20830_0[0]),.dout(n21444),.clk(gclk));
	jand g21145(.dina(w_asqrt1_5[1]),.dinb(n21444),.dout(n21445),.clk(gclk));
	jnot g21146(.din(w_n21445_0[1]),.dout(n21446),.clk(gclk));
	jor g21147(.dina(n21446),.dinb(n21443),.dout(n21447),.clk(gclk));
	jand g21148(.dina(n21447),.dinb(w_n20833_0[0]),.dout(n21448),.clk(gclk));
	jand g21149(.dina(w_n21445_0[0]),.dinb(w_n20836_0[0]),.dout(n21449),.clk(gclk));
	jor g21150(.dina(n21449),.dinb(n21448),.dout(n21450),.clk(gclk));
	jand g21151(.dina(w_n21450_0[1]),.dinb(w_n425_12[1]),.dout(n21451),.clk(gclk));
	jand g21152(.dina(w_n21438_0[0]),.dinb(w_n430_12[2]),.dout(n21452),.clk(gclk));
	jor g21153(.dina(n21452),.dinb(n21451),.dout(n21453),.clk(gclk));
	jor g21154(.dina(n21453),.dinb(n21442),.dout(n21454),.clk(gclk));
	jnot g21155(.din(w_n20845_0[0]),.dout(n21455),.clk(gclk));
	jnot g21156(.din(w_n20838_0[0]),.dout(n21456),.clk(gclk));
	jand g21157(.dina(w_asqrt1_5[0]),.dinb(n21456),.dout(n21457),.clk(gclk));
	jnot g21158(.din(w_n21457_0[1]),.dout(n21458),.clk(gclk));
	jor g21159(.dina(n21458),.dinb(n21455),.dout(n21459),.clk(gclk));
	jand g21160(.dina(n21459),.dinb(w_n20842_0[0]),.dout(n21460),.clk(gclk));
	jand g21161(.dina(w_n21457_0[0]),.dinb(w_n20846_0[0]),.dout(n21461),.clk(gclk));
	jor g21162(.dina(n21461),.dinb(n21460),.dout(n21462),.clk(gclk));
	jor g21163(.dina(w_n21462_0[1]),.dinb(w_n305_13[2]),.dout(n21463),.clk(gclk));
	jor g21164(.dina(w_n21450_0[0]),.dinb(w_n425_12[0]),.dout(n21464),.clk(gclk));
	jand g21165(.dina(n21464),.dinb(n21463),.dout(n21465),.clk(gclk));
	jand g21166(.dina(n21465),.dinb(n21454),.dout(n21466),.clk(gclk));
	jxor g21167(.dina(w_n20847_0[0]),.dinb(w_n305_13[1]),.dout(n21467),.clk(gclk));
	jor g21168(.dina(n21467),.dinb(w_n20910_6[0]),.dout(n21468),.clk(gclk));
	jxor g21169(.dina(n21468),.dinb(w_n20858_0[0]),.dout(n21469),.clk(gclk));
	jand g21170(.dina(w_n21469_0[1]),.dinb(w_n290_13[1]),.dout(n21470),.clk(gclk));
	jand g21171(.dina(w_n21462_0[0]),.dinb(w_n305_13[0]),.dout(n21471),.clk(gclk));
	jor g21172(.dina(n21471),.dinb(n21470),.dout(n21472),.clk(gclk));
	jor g21173(.dina(n21472),.dinb(n21466),.dout(n21473),.clk(gclk));
	jnot g21174(.din(w_n20868_0[0]),.dout(n21474),.clk(gclk));
	jnot g21175(.din(w_n20861_0[0]),.dout(n21475),.clk(gclk));
	jand g21176(.dina(w_asqrt1_4[2]),.dinb(n21475),.dout(n21476),.clk(gclk));
	jnot g21177(.din(w_n21476_0[1]),.dout(n21477),.clk(gclk));
	jor g21178(.dina(n21477),.dinb(n21474),.dout(n21478),.clk(gclk));
	jand g21179(.dina(n21478),.dinb(w_n20865_0[0]),.dout(n21479),.clk(gclk));
	jand g21180(.dina(w_n21476_0[0]),.dinb(w_n20869_0[0]),.dout(n21480),.clk(gclk));
	jor g21181(.dina(n21480),.dinb(n21479),.dout(n21481),.clk(gclk));
	jor g21182(.dina(w_n21481_0[1]),.dinb(w_n223_13[1]),.dout(n21482),.clk(gclk));
	jor g21183(.dina(w_n21469_0[0]),.dinb(w_n290_13[0]),.dout(n21483),.clk(gclk));
	jand g21184(.dina(n21483),.dinb(n21482),.dout(n21484),.clk(gclk));
	jand g21185(.dina(n21484),.dinb(n21473),.dout(n21485),.clk(gclk));
	jand g21186(.dina(w_n20913_0[0]),.dinb(w_n199_15[0]),.dout(n21486),.clk(gclk));
	jand g21187(.dina(w_n21481_0[0]),.dinb(w_n223_13[0]),.dout(n21487),.clk(gclk));
	jor g21188(.dina(n21487),.dinb(n21486),.dout(n21488),.clk(gclk));
	jor g21189(.dina(n21488),.dinb(n21485),.dout(n21489),.clk(gclk));
	jand g21190(.dina(n21489),.dinb(n20914),.dout(n21490),.clk(gclk));
	jnot g21191(.din(w_n20877_0[0]),.dout(n21491),.clk(gclk));
	jor g21192(.dina(n21491),.dinb(w_n20875_0[0]),.dout(n21492),.clk(gclk));
	jor g21193(.dina(n21492),.dinb(w_n20910_5[2]),.dout(n21493),.clk(gclk));
	jxor g21194(.dina(n21493),.dinb(w_n20886_0[0]),.dout(n21494),.clk(gclk));
	jnot g21195(.din(w_n20902_0[0]),.dout(n21495),.clk(gclk));
	jand g21196(.dina(w_asqrt1_4[1]),.dinb(w_n20901_0[0]),.dout(n21496),.clk(gclk));
	jand g21197(.dina(w_n21496_0[1]),.dinb(w_n20888_1[0]),.dout(n21497),.clk(gclk));
	jor g21198(.dina(n21497),.dinb(n21495),.dout(n21498),.clk(gclk));
	jor g21199(.dina(n21498),.dinb(w_n21494_0[1]),.dout(n21499),.clk(gclk));
	jor g21200(.dina(n21499),.dinb(w_n21490_0[1]),.dout(n21500),.clk(gclk));
	jand g21201(.dina(n21500),.dinb(w_n194_14[1]),.dout(n21501),.clk(gclk));
	jand g21202(.dina(w_n21494_0[0]),.dinb(w_n21490_0[0]),.dout(n21502),.clk(gclk));
	jor g21203(.dina(w_n21496_0[0]),.dinb(w_n20888_0[2]),.dout(n21503),.clk(gclk));
	jnot g21204(.din(w_n20888_0[1]),.dout(n21504),.clk(gclk));
	jor g21205(.dina(w_n20891_0[0]),.dinb(n21504),.dout(n21505),.clk(gclk));
	jand g21206(.dina(n21505),.dinb(w_asqrt63_5[2]),.dout(n21506),.clk(gclk));
	jand g21207(.dina(n21506),.dinb(n21503),.dout(n21507),.clk(gclk));
	jor g21208(.dina(n21507),.dinb(n21502),.dout(n21508),.clk(gclk));
	jor g21209(.dina(n21508),.dinb(n21501),.dout(asqrt_fa_1),.clk(gclk));
	jspl3 jspl3_w_a2_0(.douta(w_a2_0[0]),.doutb(w_a2_0[1]),.doutc(w_a2_0[2]),.din(a[2]));
	jspl jspl_w_a3_0(.douta(w_a3_0[0]),.doutb(w_a3_0[1]),.din(a[3]));
	jspl jspl_w_a4_0(.douta(w_a4_0[0]),.doutb(w_a4_0[1]),.din(a[4]));
	jspl jspl_w_a6_0(.douta(w_a6_0[0]),.doutb(w_a6_0[1]),.din(a[6]));
	jspl jspl_w_a7_0(.douta(w_a7_0[0]),.doutb(w_a7_0[1]),.din(a[7]));
	jspl jspl_w_a8_0(.douta(w_a8_0[0]),.doutb(w_a8_0[1]),.din(a[8]));
	jspl jspl_w_a10_0(.douta(w_a10_0[0]),.doutb(w_a10_0[1]),.din(a[10]));
	jspl jspl_w_a11_0(.douta(w_a11_0[0]),.doutb(w_a11_0[1]),.din(a[11]));
	jspl jspl_w_a12_0(.douta(w_a12_0[0]),.doutb(w_a12_0[1]),.din(a[12]));
	jspl jspl_w_a14_0(.douta(w_a14_0[0]),.doutb(w_a14_0[1]),.din(a[14]));
	jspl jspl_w_a15_0(.douta(w_a15_0[0]),.doutb(w_a15_0[1]),.din(a[15]));
	jspl jspl_w_a16_0(.douta(w_a16_0[0]),.doutb(w_a16_0[1]),.din(a[16]));
	jspl jspl_w_a18_0(.douta(w_a18_0[0]),.doutb(w_a18_0[1]),.din(a[18]));
	jspl jspl_w_a19_0(.douta(w_a19_0[0]),.doutb(w_a19_0[1]),.din(a[19]));
	jspl jspl_w_a20_0(.douta(w_a20_0[0]),.doutb(w_a20_0[1]),.din(a[20]));
	jspl jspl_w_a22_0(.douta(w_a22_0[0]),.doutb(w_a22_0[1]),.din(a[22]));
	jspl jspl_w_a23_0(.douta(w_a23_0[0]),.doutb(w_a23_0[1]),.din(a[23]));
	jspl jspl_w_a24_0(.douta(w_a24_0[0]),.doutb(w_a24_0[1]),.din(a[24]));
	jspl jspl_w_a26_0(.douta(w_a26_0[0]),.doutb(w_a26_0[1]),.din(a[26]));
	jspl jspl_w_a27_0(.douta(w_a27_0[0]),.doutb(w_a27_0[1]),.din(a[27]));
	jspl jspl_w_a28_0(.douta(w_a28_0[0]),.doutb(w_a28_0[1]),.din(a[28]));
	jspl jspl_w_a30_0(.douta(w_a30_0[0]),.doutb(w_a30_0[1]),.din(a[30]));
	jspl jspl_w_a31_0(.douta(w_a31_0[0]),.doutb(w_a31_0[1]),.din(a[31]));
	jspl jspl_w_a32_0(.douta(w_a32_0[0]),.doutb(w_a32_0[1]),.din(a[32]));
	jspl jspl_w_a34_0(.douta(w_a34_0[0]),.doutb(w_a34_0[1]),.din(a[34]));
	jspl jspl_w_a35_0(.douta(w_a35_0[0]),.doutb(w_a35_0[1]),.din(a[35]));
	jspl jspl_w_a36_0(.douta(w_a36_0[0]),.doutb(w_a36_0[1]),.din(a[36]));
	jspl jspl_w_a38_0(.douta(w_a38_0[0]),.doutb(w_a38_0[1]),.din(a[38]));
	jspl jspl_w_a39_0(.douta(w_a39_0[0]),.doutb(w_a39_0[1]),.din(a[39]));
	jspl jspl_w_a40_0(.douta(w_a40_0[0]),.doutb(w_a40_0[1]),.din(a[40]));
	jspl jspl_w_a42_0(.douta(w_a42_0[0]),.doutb(w_a42_0[1]),.din(a[42]));
	jspl jspl_w_a43_0(.douta(w_a43_0[0]),.doutb(w_a43_0[1]),.din(a[43]));
	jspl jspl_w_a44_0(.douta(w_a44_0[0]),.doutb(w_a44_0[1]),.din(a[44]));
	jspl jspl_w_a46_0(.douta(w_a46_0[0]),.doutb(w_a46_0[1]),.din(a[46]));
	jspl jspl_w_a47_0(.douta(w_a47_0[0]),.doutb(w_a47_0[1]),.din(a[47]));
	jspl jspl_w_a48_0(.douta(w_a48_0[0]),.doutb(w_a48_0[1]),.din(a[48]));
	jspl jspl_w_a50_0(.douta(w_a50_0[0]),.doutb(w_a50_0[1]),.din(a[50]));
	jspl jspl_w_a51_0(.douta(w_a51_0[0]),.doutb(w_a51_0[1]),.din(a[51]));
	jspl jspl_w_a52_0(.douta(w_a52_0[0]),.doutb(w_a52_0[1]),.din(a[52]));
	jspl jspl_w_a54_0(.douta(w_a54_0[0]),.doutb(w_a54_0[1]),.din(a[54]));
	jspl jspl_w_a55_0(.douta(w_a55_0[0]),.doutb(w_a55_0[1]),.din(a[55]));
	jspl jspl_w_a56_0(.douta(w_a56_0[0]),.doutb(w_a56_0[1]),.din(a[56]));
	jspl jspl_w_a58_0(.douta(w_a58_0[0]),.doutb(w_a58_0[1]),.din(a[58]));
	jspl jspl_w_a59_0(.douta(w_a59_0[0]),.doutb(w_a59_0[1]),.din(a[59]));
	jspl jspl_w_a60_0(.douta(w_a60_0[0]),.doutb(w_a60_0[1]),.din(a[60]));
	jspl jspl_w_a62_0(.douta(w_a62_0[0]),.doutb(w_a62_0[1]),.din(a[62]));
	jspl jspl_w_a63_0(.douta(w_a63_0[0]),.doutb(w_a63_0[1]),.din(a[63]));
	jspl jspl_w_a64_0(.douta(w_a64_0[0]),.doutb(w_a64_0[1]),.din(a[64]));
	jspl jspl_w_a66_0(.douta(w_a66_0[0]),.doutb(w_a66_0[1]),.din(a[66]));
	jspl jspl_w_a67_0(.douta(w_a67_0[0]),.doutb(w_a67_0[1]),.din(a[67]));
	jspl jspl_w_a68_0(.douta(w_a68_0[0]),.doutb(w_a68_0[1]),.din(a[68]));
	jspl jspl_w_a70_0(.douta(w_a70_0[0]),.doutb(w_a70_0[1]),.din(a[70]));
	jspl jspl_w_a71_0(.douta(w_a71_0[0]),.doutb(w_a71_0[1]),.din(a[71]));
	jspl jspl_w_a72_0(.douta(w_a72_0[0]),.doutb(w_a72_0[1]),.din(a[72]));
	jspl jspl_w_a74_0(.douta(w_a74_0[0]),.doutb(w_a74_0[1]),.din(a[74]));
	jspl jspl_w_a75_0(.douta(w_a75_0[0]),.doutb(w_a75_0[1]),.din(a[75]));
	jspl jspl_w_a76_0(.douta(w_a76_0[0]),.doutb(w_a76_0[1]),.din(a[76]));
	jspl jspl_w_a78_0(.douta(w_a78_0[0]),.doutb(w_a78_0[1]),.din(a[78]));
	jspl jspl_w_a79_0(.douta(w_a79_0[0]),.doutb(w_a79_0[1]),.din(a[79]));
	jspl jspl_w_a80_0(.douta(w_a80_0[0]),.doutb(w_a80_0[1]),.din(a[80]));
	jspl jspl_w_a82_0(.douta(w_a82_0[0]),.doutb(w_a82_0[1]),.din(a[82]));
	jspl jspl_w_a83_0(.douta(w_a83_0[0]),.doutb(w_a83_0[1]),.din(a[83]));
	jspl jspl_w_a84_0(.douta(w_a84_0[0]),.doutb(w_a84_0[1]),.din(a[84]));
	jspl jspl_w_a86_0(.douta(w_a86_0[0]),.doutb(w_a86_0[1]),.din(a[86]));
	jspl jspl_w_a87_0(.douta(w_a87_0[0]),.doutb(w_a87_0[1]),.din(a[87]));
	jspl jspl_w_a88_0(.douta(w_a88_0[0]),.doutb(w_a88_0[1]),.din(a[88]));
	jspl jspl_w_a90_0(.douta(w_a90_0[0]),.doutb(w_a90_0[1]),.din(a[90]));
	jspl jspl_w_a91_0(.douta(w_a91_0[0]),.doutb(w_a91_0[1]),.din(a[91]));
	jspl jspl_w_a92_0(.douta(w_a92_0[0]),.doutb(w_a92_0[1]),.din(a[92]));
	jspl jspl_w_a94_0(.douta(w_a94_0[0]),.doutb(w_a94_0[1]),.din(a[94]));
	jspl jspl_w_a95_0(.douta(w_a95_0[0]),.doutb(w_a95_0[1]),.din(a[95]));
	jspl jspl_w_a96_0(.douta(w_a96_0[0]),.doutb(w_a96_0[1]),.din(a[96]));
	jspl jspl_w_a98_0(.douta(w_a98_0[0]),.doutb(w_a98_0[1]),.din(a[98]));
	jspl jspl_w_a99_0(.douta(w_a99_0[0]),.doutb(w_a99_0[1]),.din(a[99]));
	jspl jspl_w_a100_0(.douta(w_a100_0[0]),.doutb(w_a100_0[1]),.din(a[100]));
	jspl jspl_w_a102_0(.douta(w_a102_0[0]),.doutb(w_a102_0[1]),.din(a[102]));
	jspl jspl_w_a103_0(.douta(w_a103_0[0]),.doutb(w_a103_0[1]),.din(a[103]));
	jspl jspl_w_a104_0(.douta(w_a104_0[0]),.doutb(w_a104_0[1]),.din(a[104]));
	jspl jspl_w_a106_0(.douta(w_a106_0[0]),.doutb(w_a106_0[1]),.din(a[106]));
	jspl jspl_w_a107_0(.douta(w_a107_0[0]),.doutb(w_a107_0[1]),.din(a[107]));
	jspl jspl_w_a108_0(.douta(w_a108_0[0]),.doutb(w_a108_0[1]),.din(a[108]));
	jspl jspl_w_a110_0(.douta(w_a110_0[0]),.doutb(w_a110_0[1]),.din(a[110]));
	jspl jspl_w_a111_0(.douta(w_a111_0[0]),.doutb(w_a111_0[1]),.din(a[111]));
	jspl jspl_w_a112_0(.douta(w_a112_0[0]),.doutb(w_a112_0[1]),.din(a[112]));
	jspl jspl_w_a114_0(.douta(w_a114_0[0]),.doutb(w_a114_0[1]),.din(a[114]));
	jspl jspl_w_a115_0(.douta(w_a115_0[0]),.doutb(w_a115_0[1]),.din(a[115]));
	jspl jspl_w_a116_0(.douta(w_a116_0[0]),.doutb(w_a116_0[1]),.din(a[116]));
	jspl jspl_w_a118_0(.douta(w_a118_0[0]),.doutb(w_a118_0[1]),.din(a[118]));
	jspl jspl_w_a119_0(.douta(w_a119_0[0]),.doutb(w_a119_0[1]),.din(a[119]));
	jspl jspl_w_a120_0(.douta(w_a120_0[0]),.doutb(w_a120_0[1]),.din(a[120]));
	jspl jspl_w_a122_0(.douta(w_a122_0[0]),.doutb(w_a122_0[1]),.din(a[122]));
	jspl jspl_w_a123_0(.douta(w_a123_0[0]),.doutb(w_a123_0[1]),.din(a[123]));
	jspl3 jspl3_w_a124_0(.douta(w_a124_0[0]),.doutb(w_a124_0[1]),.doutc(w_a124_0[2]),.din(a[124]));
	jspl jspl_w_a125_0(.douta(w_a125_0[0]),.doutb(w_a125_0[1]),.din(a[125]));
	jspl3 jspl3_w_a126_0(.douta(w_a126_0[0]),.doutb(w_a126_0[1]),.doutc(w_a126_0[2]),.din(a[126]));
	jspl jspl_w_a127_0(.douta(w_a127_0[0]),.doutb(w_a127_0[1]),.din(a[127]));
	jspl3 jspl3_w_asqrt1_0(.douta(w_asqrt1_0[0]),.doutb(w_asqrt1_0[1]),.doutc(w_asqrt1_0[2]),.din(asqrt_fa_1));
	jspl3 jspl3_w_asqrt1_1(.douta(w_asqrt1_1[0]),.doutb(w_asqrt1_1[1]),.doutc(w_asqrt1_1[2]),.din(w_asqrt1_0[0]));
	jspl3 jspl3_w_asqrt1_2(.douta(w_asqrt1_2[0]),.doutb(w_asqrt1_2[1]),.doutc(w_asqrt1_2[2]),.din(w_asqrt1_0[1]));
	jspl3 jspl3_w_asqrt1_3(.douta(w_asqrt1_3[0]),.doutb(w_asqrt1_3[1]),.doutc(w_asqrt1_3[2]),.din(w_asqrt1_0[2]));
	jspl3 jspl3_w_asqrt1_4(.douta(w_asqrt1_4[0]),.doutb(w_asqrt1_4[1]),.doutc(w_asqrt1_4[2]),.din(w_asqrt1_1[0]));
	jspl3 jspl3_w_asqrt1_5(.douta(w_asqrt1_5[0]),.doutb(w_asqrt1_5[1]),.doutc(w_asqrt1_5[2]),.din(w_asqrt1_1[1]));
	jspl3 jspl3_w_asqrt1_6(.douta(w_asqrt1_6[0]),.doutb(w_asqrt1_6[1]),.doutc(w_asqrt1_6[2]),.din(w_asqrt1_1[2]));
	jspl3 jspl3_w_asqrt1_7(.douta(w_asqrt1_7[0]),.doutb(w_asqrt1_7[1]),.doutc(w_asqrt1_7[2]),.din(w_asqrt1_2[0]));
	jspl3 jspl3_w_asqrt1_8(.douta(w_asqrt1_8[0]),.doutb(w_asqrt1_8[1]),.doutc(w_asqrt1_8[2]),.din(w_asqrt1_2[1]));
	jspl3 jspl3_w_asqrt1_9(.douta(w_asqrt1_9[0]),.doutb(w_asqrt1_9[1]),.doutc(w_asqrt1_9[2]),.din(w_asqrt1_2[2]));
	jspl3 jspl3_w_asqrt1_10(.douta(w_asqrt1_10[0]),.doutb(w_asqrt1_10[1]),.doutc(w_asqrt1_10[2]),.din(w_asqrt1_3[0]));
	jspl3 jspl3_w_asqrt1_11(.douta(w_asqrt1_11[0]),.doutb(w_asqrt1_11[1]),.doutc(w_asqrt1_11[2]),.din(w_asqrt1_3[1]));
	jspl3 jspl3_w_asqrt1_12(.douta(w_asqrt1_12[0]),.doutb(w_asqrt1_12[1]),.doutc(w_asqrt1_12[2]),.din(w_asqrt1_3[2]));
	jspl3 jspl3_w_asqrt1_13(.douta(w_asqrt1_13[0]),.doutb(w_asqrt1_13[1]),.doutc(asqrt[0]),.din(w_asqrt1_4[0]));
	jspl3 jspl3_w_asqrt2_0(.douta(w_asqrt2_0[0]),.doutb(w_asqrt2_0[1]),.doutc(w_asqrt2_0[2]),.din(asqrt_fa_2));
	jspl3 jspl3_w_asqrt2_1(.douta(w_asqrt2_1[0]),.doutb(w_asqrt2_1[1]),.doutc(w_asqrt2_1[2]),.din(w_asqrt2_0[0]));
	jspl3 jspl3_w_asqrt2_2(.douta(w_asqrt2_2[0]),.doutb(w_asqrt2_2[1]),.doutc(w_asqrt2_2[2]),.din(w_asqrt2_0[1]));
	jspl3 jspl3_w_asqrt2_3(.douta(w_asqrt2_3[0]),.doutb(w_asqrt2_3[1]),.doutc(w_asqrt2_3[2]),.din(w_asqrt2_0[2]));
	jspl3 jspl3_w_asqrt2_4(.douta(w_asqrt2_4[0]),.doutb(w_asqrt2_4[1]),.doutc(w_asqrt2_4[2]),.din(w_asqrt2_1[0]));
	jspl3 jspl3_w_asqrt2_5(.douta(w_asqrt2_5[0]),.doutb(w_asqrt2_5[1]),.doutc(w_asqrt2_5[2]),.din(w_asqrt2_1[1]));
	jspl3 jspl3_w_asqrt2_6(.douta(w_asqrt2_6[0]),.doutb(w_asqrt2_6[1]),.doutc(w_asqrt2_6[2]),.din(w_asqrt2_1[2]));
	jspl3 jspl3_w_asqrt2_7(.douta(w_asqrt2_7[0]),.doutb(w_asqrt2_7[1]),.doutc(w_asqrt2_7[2]),.din(w_asqrt2_2[0]));
	jspl3 jspl3_w_asqrt2_8(.douta(w_asqrt2_8[0]),.doutb(w_asqrt2_8[1]),.doutc(w_asqrt2_8[2]),.din(w_asqrt2_2[1]));
	jspl3 jspl3_w_asqrt2_9(.douta(w_asqrt2_9[0]),.doutb(w_asqrt2_9[1]),.doutc(w_asqrt2_9[2]),.din(w_asqrt2_2[2]));
	jspl3 jspl3_w_asqrt2_10(.douta(w_asqrt2_10[0]),.doutb(w_asqrt2_10[1]),.doutc(w_asqrt2_10[2]),.din(w_asqrt2_3[0]));
	jspl3 jspl3_w_asqrt2_11(.douta(w_asqrt2_11[0]),.doutb(w_asqrt2_11[1]),.doutc(w_asqrt2_11[2]),.din(w_asqrt2_3[1]));
	jspl3 jspl3_w_asqrt2_12(.douta(w_asqrt2_12[0]),.doutb(w_asqrt2_12[1]),.doutc(w_asqrt2_12[2]),.din(w_asqrt2_3[2]));
	jspl3 jspl3_w_asqrt2_13(.douta(w_asqrt2_13[0]),.doutb(w_asqrt2_13[1]),.doutc(w_asqrt2_13[2]),.din(w_asqrt2_4[0]));
	jspl3 jspl3_w_asqrt2_14(.douta(w_asqrt2_14[0]),.doutb(w_asqrt2_14[1]),.doutc(w_asqrt2_14[2]),.din(w_asqrt2_4[1]));
	jspl3 jspl3_w_asqrt2_15(.douta(w_asqrt2_15[0]),.doutb(w_asqrt2_15[1]),.doutc(w_asqrt2_15[2]),.din(w_asqrt2_4[2]));
	jspl3 jspl3_w_asqrt2_16(.douta(w_asqrt2_16[0]),.doutb(w_asqrt2_16[1]),.doutc(w_asqrt2_16[2]),.din(w_asqrt2_5[0]));
	jspl3 jspl3_w_asqrt2_17(.douta(w_asqrt2_17[0]),.doutb(w_asqrt2_17[1]),.doutc(w_asqrt2_17[2]),.din(w_asqrt2_5[1]));
	jspl3 jspl3_w_asqrt2_18(.douta(w_asqrt2_18[0]),.doutb(w_asqrt2_18[1]),.doutc(w_asqrt2_18[2]),.din(w_asqrt2_5[2]));
	jspl3 jspl3_w_asqrt2_19(.douta(w_asqrt2_19[0]),.doutb(w_asqrt2_19[1]),.doutc(w_asqrt2_19[2]),.din(w_asqrt2_6[0]));
	jspl3 jspl3_w_asqrt2_20(.douta(w_asqrt2_20[0]),.doutb(w_asqrt2_20[1]),.doutc(w_asqrt2_20[2]),.din(w_asqrt2_6[1]));
	jspl3 jspl3_w_asqrt2_21(.douta(w_asqrt2_21[0]),.doutb(w_asqrt2_21[1]),.doutc(w_asqrt2_21[2]),.din(w_asqrt2_6[2]));
	jspl3 jspl3_w_asqrt2_22(.douta(w_asqrt2_22[0]),.doutb(w_asqrt2_22[1]),.doutc(w_asqrt2_22[2]),.din(w_asqrt2_7[0]));
	jspl3 jspl3_w_asqrt2_23(.douta(w_asqrt2_23[0]),.doutb(w_asqrt2_23[1]),.doutc(w_asqrt2_23[2]),.din(w_asqrt2_7[1]));
	jspl3 jspl3_w_asqrt2_24(.douta(w_asqrt2_24[0]),.doutb(w_asqrt2_24[1]),.doutc(w_asqrt2_24[2]),.din(w_asqrt2_7[2]));
	jspl3 jspl3_w_asqrt2_25(.douta(w_asqrt2_25[0]),.doutb(w_asqrt2_25[1]),.doutc(w_asqrt2_25[2]),.din(w_asqrt2_8[0]));
	jspl3 jspl3_w_asqrt2_26(.douta(w_asqrt2_26[0]),.doutb(w_asqrt2_26[1]),.doutc(w_asqrt2_26[2]),.din(w_asqrt2_8[1]));
	jspl3 jspl3_w_asqrt2_27(.douta(w_asqrt2_27[0]),.doutb(w_asqrt2_27[1]),.doutc(w_asqrt2_27[2]),.din(w_asqrt2_8[2]));
	jspl3 jspl3_w_asqrt2_28(.douta(w_asqrt2_28[0]),.doutb(w_asqrt2_28[1]),.doutc(w_asqrt2_28[2]),.din(w_asqrt2_9[0]));
	jspl3 jspl3_w_asqrt2_29(.douta(w_asqrt2_29[0]),.doutb(w_asqrt2_29[1]),.doutc(w_asqrt2_29[2]),.din(w_asqrt2_9[1]));
	jspl3 jspl3_w_asqrt2_30(.douta(w_asqrt2_30[0]),.doutb(w_asqrt2_30[1]),.doutc(w_asqrt2_30[2]),.din(w_asqrt2_9[2]));
	jspl jspl_w_asqrt2_31(.douta(w_asqrt2_31),.doutb(asqrt[1]),.din(w_asqrt2_10[0]));
	jspl3 jspl3_w_asqrt3_0(.douta(w_asqrt3_0[0]),.doutb(w_asqrt3_0[1]),.doutc(w_asqrt3_0[2]),.din(asqrt_fa_3));
	jspl3 jspl3_w_asqrt3_1(.douta(w_asqrt3_1[0]),.doutb(w_asqrt3_1[1]),.doutc(w_asqrt3_1[2]),.din(w_asqrt3_0[0]));
	jspl3 jspl3_w_asqrt3_2(.douta(w_asqrt3_2[0]),.doutb(w_asqrt3_2[1]),.doutc(w_asqrt3_2[2]),.din(w_asqrt3_0[1]));
	jspl3 jspl3_w_asqrt3_3(.douta(w_asqrt3_3[0]),.doutb(w_asqrt3_3[1]),.doutc(w_asqrt3_3[2]),.din(w_asqrt3_0[2]));
	jspl3 jspl3_w_asqrt3_4(.douta(w_asqrt3_4[0]),.doutb(w_asqrt3_4[1]),.doutc(w_asqrt3_4[2]),.din(w_asqrt3_1[0]));
	jspl3 jspl3_w_asqrt3_5(.douta(w_asqrt3_5[0]),.doutb(w_asqrt3_5[1]),.doutc(w_asqrt3_5[2]),.din(w_asqrt3_1[1]));
	jspl3 jspl3_w_asqrt3_6(.douta(w_asqrt3_6[0]),.doutb(w_asqrt3_6[1]),.doutc(w_asqrt3_6[2]),.din(w_asqrt3_1[2]));
	jspl3 jspl3_w_asqrt3_7(.douta(w_asqrt3_7[0]),.doutb(w_asqrt3_7[1]),.doutc(w_asqrt3_7[2]),.din(w_asqrt3_2[0]));
	jspl3 jspl3_w_asqrt3_8(.douta(w_asqrt3_8[0]),.doutb(w_asqrt3_8[1]),.doutc(w_asqrt3_8[2]),.din(w_asqrt3_2[1]));
	jspl3 jspl3_w_asqrt3_9(.douta(w_asqrt3_9[0]),.doutb(w_asqrt3_9[1]),.doutc(w_asqrt3_9[2]),.din(w_asqrt3_2[2]));
	jspl3 jspl3_w_asqrt3_10(.douta(w_asqrt3_10[0]),.doutb(w_asqrt3_10[1]),.doutc(w_asqrt3_10[2]),.din(w_asqrt3_3[0]));
	jspl3 jspl3_w_asqrt3_11(.douta(w_asqrt3_11[0]),.doutb(w_asqrt3_11[1]),.doutc(w_asqrt3_11[2]),.din(w_asqrt3_3[1]));
	jspl3 jspl3_w_asqrt3_12(.douta(w_asqrt3_12[0]),.doutb(w_asqrt3_12[1]),.doutc(w_asqrt3_12[2]),.din(w_asqrt3_3[2]));
	jspl3 jspl3_w_asqrt3_13(.douta(w_asqrt3_13[0]),.doutb(w_asqrt3_13[1]),.doutc(w_asqrt3_13[2]),.din(w_asqrt3_4[0]));
	jspl3 jspl3_w_asqrt3_14(.douta(w_asqrt3_14[0]),.doutb(w_asqrt3_14[1]),.doutc(asqrt[2]),.din(w_asqrt3_4[1]));
	jspl3 jspl3_w_asqrt4_0(.douta(w_asqrt4_0[0]),.doutb(w_asqrt4_0[1]),.doutc(w_asqrt4_0[2]),.din(asqrt_fa_4));
	jspl3 jspl3_w_asqrt4_1(.douta(w_asqrt4_1[0]),.doutb(w_asqrt4_1[1]),.doutc(w_asqrt4_1[2]),.din(w_asqrt4_0[0]));
	jspl3 jspl3_w_asqrt4_2(.douta(w_asqrt4_2[0]),.doutb(w_asqrt4_2[1]),.doutc(w_asqrt4_2[2]),.din(w_asqrt4_0[1]));
	jspl3 jspl3_w_asqrt4_3(.douta(w_asqrt4_3[0]),.doutb(w_asqrt4_3[1]),.doutc(w_asqrt4_3[2]),.din(w_asqrt4_0[2]));
	jspl3 jspl3_w_asqrt4_4(.douta(w_asqrt4_4[0]),.doutb(w_asqrt4_4[1]),.doutc(w_asqrt4_4[2]),.din(w_asqrt4_1[0]));
	jspl3 jspl3_w_asqrt4_5(.douta(w_asqrt4_5[0]),.doutb(w_asqrt4_5[1]),.doutc(w_asqrt4_5[2]),.din(w_asqrt4_1[1]));
	jspl3 jspl3_w_asqrt4_6(.douta(w_asqrt4_6[0]),.doutb(w_asqrt4_6[1]),.doutc(w_asqrt4_6[2]),.din(w_asqrt4_1[2]));
	jspl3 jspl3_w_asqrt4_7(.douta(w_asqrt4_7[0]),.doutb(w_asqrt4_7[1]),.doutc(w_asqrt4_7[2]),.din(w_asqrt4_2[0]));
	jspl3 jspl3_w_asqrt4_8(.douta(w_asqrt4_8[0]),.doutb(w_asqrt4_8[1]),.doutc(w_asqrt4_8[2]),.din(w_asqrt4_2[1]));
	jspl3 jspl3_w_asqrt4_9(.douta(w_asqrt4_9[0]),.doutb(w_asqrt4_9[1]),.doutc(w_asqrt4_9[2]),.din(w_asqrt4_2[2]));
	jspl3 jspl3_w_asqrt4_10(.douta(w_asqrt4_10[0]),.doutb(w_asqrt4_10[1]),.doutc(w_asqrt4_10[2]),.din(w_asqrt4_3[0]));
	jspl3 jspl3_w_asqrt4_11(.douta(w_asqrt4_11[0]),.doutb(w_asqrt4_11[1]),.doutc(w_asqrt4_11[2]),.din(w_asqrt4_3[1]));
	jspl3 jspl3_w_asqrt4_12(.douta(w_asqrt4_12[0]),.doutb(w_asqrt4_12[1]),.doutc(w_asqrt4_12[2]),.din(w_asqrt4_3[2]));
	jspl3 jspl3_w_asqrt4_13(.douta(w_asqrt4_13[0]),.doutb(w_asqrt4_13[1]),.doutc(w_asqrt4_13[2]),.din(w_asqrt4_4[0]));
	jspl3 jspl3_w_asqrt4_14(.douta(w_asqrt4_14[0]),.doutb(w_asqrt4_14[1]),.doutc(w_asqrt4_14[2]),.din(w_asqrt4_4[1]));
	jspl3 jspl3_w_asqrt4_15(.douta(w_asqrt4_15[0]),.doutb(w_asqrt4_15[1]),.doutc(w_asqrt4_15[2]),.din(w_asqrt4_4[2]));
	jspl3 jspl3_w_asqrt4_16(.douta(w_asqrt4_16[0]),.doutb(w_asqrt4_16[1]),.doutc(w_asqrt4_16[2]),.din(w_asqrt4_5[0]));
	jspl3 jspl3_w_asqrt4_17(.douta(w_asqrt4_17[0]),.doutb(w_asqrt4_17[1]),.doutc(w_asqrt4_17[2]),.din(w_asqrt4_5[1]));
	jspl3 jspl3_w_asqrt4_18(.douta(w_asqrt4_18[0]),.doutb(w_asqrt4_18[1]),.doutc(w_asqrt4_18[2]),.din(w_asqrt4_5[2]));
	jspl3 jspl3_w_asqrt4_19(.douta(w_asqrt4_19[0]),.doutb(w_asqrt4_19[1]),.doutc(w_asqrt4_19[2]),.din(w_asqrt4_6[0]));
	jspl3 jspl3_w_asqrt4_20(.douta(w_asqrt4_20[0]),.doutb(w_asqrt4_20[1]),.doutc(w_asqrt4_20[2]),.din(w_asqrt4_6[1]));
	jspl3 jspl3_w_asqrt4_21(.douta(w_asqrt4_21[0]),.doutb(w_asqrt4_21[1]),.doutc(w_asqrt4_21[2]),.din(w_asqrt4_6[2]));
	jspl3 jspl3_w_asqrt4_22(.douta(w_asqrt4_22[0]),.doutb(w_asqrt4_22[1]),.doutc(w_asqrt4_22[2]),.din(w_asqrt4_7[0]));
	jspl3 jspl3_w_asqrt4_23(.douta(w_asqrt4_23[0]),.doutb(w_asqrt4_23[1]),.doutc(w_asqrt4_23[2]),.din(w_asqrt4_7[1]));
	jspl3 jspl3_w_asqrt4_24(.douta(w_asqrt4_24[0]),.doutb(w_asqrt4_24[1]),.doutc(w_asqrt4_24[2]),.din(w_asqrt4_7[2]));
	jspl3 jspl3_w_asqrt4_25(.douta(w_asqrt4_25[0]),.doutb(w_asqrt4_25[1]),.doutc(w_asqrt4_25[2]),.din(w_asqrt4_8[0]));
	jspl3 jspl3_w_asqrt4_26(.douta(w_asqrt4_26[0]),.doutb(w_asqrt4_26[1]),.doutc(w_asqrt4_26[2]),.din(w_asqrt4_8[1]));
	jspl3 jspl3_w_asqrt4_27(.douta(w_asqrt4_27[0]),.doutb(w_asqrt4_27[1]),.doutc(w_asqrt4_27[2]),.din(w_asqrt4_8[2]));
	jspl3 jspl3_w_asqrt4_28(.douta(w_asqrt4_28[0]),.doutb(w_asqrt4_28[1]),.doutc(w_asqrt4_28[2]),.din(w_asqrt4_9[0]));
	jspl3 jspl3_w_asqrt4_29(.douta(w_asqrt4_29[0]),.doutb(w_asqrt4_29[1]),.doutc(w_asqrt4_29[2]),.din(w_asqrt4_9[1]));
	jspl3 jspl3_w_asqrt4_30(.douta(w_asqrt4_30[0]),.doutb(w_asqrt4_30[1]),.doutc(w_asqrt4_30[2]),.din(w_asqrt4_9[2]));
	jspl jspl_w_asqrt4_31(.douta(w_asqrt4_31),.doutb(asqrt[3]),.din(w_asqrt4_10[0]));
	jspl3 jspl3_w_asqrt5_0(.douta(w_asqrt5_0[0]),.doutb(w_asqrt5_0[1]),.doutc(w_asqrt5_0[2]),.din(asqrt_fa_5));
	jspl3 jspl3_w_asqrt5_1(.douta(w_asqrt5_1[0]),.doutb(w_asqrt5_1[1]),.doutc(w_asqrt5_1[2]),.din(w_asqrt5_0[0]));
	jspl3 jspl3_w_asqrt5_2(.douta(w_asqrt5_2[0]),.doutb(w_asqrt5_2[1]),.doutc(w_asqrt5_2[2]),.din(w_asqrt5_0[1]));
	jspl3 jspl3_w_asqrt5_3(.douta(w_asqrt5_3[0]),.doutb(w_asqrt5_3[1]),.doutc(w_asqrt5_3[2]),.din(w_asqrt5_0[2]));
	jspl3 jspl3_w_asqrt5_4(.douta(w_asqrt5_4[0]),.doutb(w_asqrt5_4[1]),.doutc(w_asqrt5_4[2]),.din(w_asqrt5_1[0]));
	jspl3 jspl3_w_asqrt5_5(.douta(w_asqrt5_5[0]),.doutb(w_asqrt5_5[1]),.doutc(w_asqrt5_5[2]),.din(w_asqrt5_1[1]));
	jspl3 jspl3_w_asqrt5_6(.douta(w_asqrt5_6[0]),.doutb(w_asqrt5_6[1]),.doutc(w_asqrt5_6[2]),.din(w_asqrt5_1[2]));
	jspl3 jspl3_w_asqrt5_7(.douta(w_asqrt5_7[0]),.doutb(w_asqrt5_7[1]),.doutc(w_asqrt5_7[2]),.din(w_asqrt5_2[0]));
	jspl3 jspl3_w_asqrt5_8(.douta(w_asqrt5_8[0]),.doutb(w_asqrt5_8[1]),.doutc(w_asqrt5_8[2]),.din(w_asqrt5_2[1]));
	jspl3 jspl3_w_asqrt5_9(.douta(w_asqrt5_9[0]),.doutb(w_asqrt5_9[1]),.doutc(w_asqrt5_9[2]),.din(w_asqrt5_2[2]));
	jspl3 jspl3_w_asqrt5_10(.douta(w_asqrt5_10[0]),.doutb(w_asqrt5_10[1]),.doutc(w_asqrt5_10[2]),.din(w_asqrt5_3[0]));
	jspl3 jspl3_w_asqrt5_11(.douta(w_asqrt5_11[0]),.doutb(w_asqrt5_11[1]),.doutc(w_asqrt5_11[2]),.din(w_asqrt5_3[1]));
	jspl3 jspl3_w_asqrt5_12(.douta(w_asqrt5_12[0]),.doutb(w_asqrt5_12[1]),.doutc(w_asqrt5_12[2]),.din(w_asqrt5_3[2]));
	jspl3 jspl3_w_asqrt5_13(.douta(w_asqrt5_13[0]),.doutb(w_asqrt5_13[1]),.doutc(w_asqrt5_13[2]),.din(w_asqrt5_4[0]));
	jspl3 jspl3_w_asqrt5_14(.douta(w_asqrt5_14[0]),.doutb(w_asqrt5_14[1]),.doutc(w_asqrt5_14[2]),.din(w_asqrt5_4[1]));
	jspl3 jspl3_w_asqrt5_15(.douta(w_asqrt5_15[0]),.doutb(w_asqrt5_15[1]),.doutc(asqrt[4]),.din(w_asqrt5_4[2]));
	jspl3 jspl3_w_asqrt6_0(.douta(w_asqrt6_0[0]),.doutb(w_asqrt6_0[1]),.doutc(w_asqrt6_0[2]),.din(asqrt_fa_6));
	jspl3 jspl3_w_asqrt6_1(.douta(w_asqrt6_1[0]),.doutb(w_asqrt6_1[1]),.doutc(w_asqrt6_1[2]),.din(w_asqrt6_0[0]));
	jspl3 jspl3_w_asqrt6_2(.douta(w_asqrt6_2[0]),.doutb(w_asqrt6_2[1]),.doutc(w_asqrt6_2[2]),.din(w_asqrt6_0[1]));
	jspl3 jspl3_w_asqrt6_3(.douta(w_asqrt6_3[0]),.doutb(w_asqrt6_3[1]),.doutc(w_asqrt6_3[2]),.din(w_asqrt6_0[2]));
	jspl3 jspl3_w_asqrt6_4(.douta(w_asqrt6_4[0]),.doutb(w_asqrt6_4[1]),.doutc(w_asqrt6_4[2]),.din(w_asqrt6_1[0]));
	jspl3 jspl3_w_asqrt6_5(.douta(w_asqrt6_5[0]),.doutb(w_asqrt6_5[1]),.doutc(w_asqrt6_5[2]),.din(w_asqrt6_1[1]));
	jspl3 jspl3_w_asqrt6_6(.douta(w_asqrt6_6[0]),.doutb(w_asqrt6_6[1]),.doutc(w_asqrt6_6[2]),.din(w_asqrt6_1[2]));
	jspl3 jspl3_w_asqrt6_7(.douta(w_asqrt6_7[0]),.doutb(w_asqrt6_7[1]),.doutc(w_asqrt6_7[2]),.din(w_asqrt6_2[0]));
	jspl3 jspl3_w_asqrt6_8(.douta(w_asqrt6_8[0]),.doutb(w_asqrt6_8[1]),.doutc(w_asqrt6_8[2]),.din(w_asqrt6_2[1]));
	jspl3 jspl3_w_asqrt6_9(.douta(w_asqrt6_9[0]),.doutb(w_asqrt6_9[1]),.doutc(w_asqrt6_9[2]),.din(w_asqrt6_2[2]));
	jspl3 jspl3_w_asqrt6_10(.douta(w_asqrt6_10[0]),.doutb(w_asqrt6_10[1]),.doutc(w_asqrt6_10[2]),.din(w_asqrt6_3[0]));
	jspl3 jspl3_w_asqrt6_11(.douta(w_asqrt6_11[0]),.doutb(w_asqrt6_11[1]),.doutc(w_asqrt6_11[2]),.din(w_asqrt6_3[1]));
	jspl3 jspl3_w_asqrt6_12(.douta(w_asqrt6_12[0]),.doutb(w_asqrt6_12[1]),.doutc(w_asqrt6_12[2]),.din(w_asqrt6_3[2]));
	jspl3 jspl3_w_asqrt6_13(.douta(w_asqrt6_13[0]),.doutb(w_asqrt6_13[1]),.doutc(w_asqrt6_13[2]),.din(w_asqrt6_4[0]));
	jspl3 jspl3_w_asqrt6_14(.douta(w_asqrt6_14[0]),.doutb(w_asqrt6_14[1]),.doutc(w_asqrt6_14[2]),.din(w_asqrt6_4[1]));
	jspl3 jspl3_w_asqrt6_15(.douta(w_asqrt6_15[0]),.doutb(w_asqrt6_15[1]),.doutc(w_asqrt6_15[2]),.din(w_asqrt6_4[2]));
	jspl3 jspl3_w_asqrt6_16(.douta(w_asqrt6_16[0]),.doutb(w_asqrt6_16[1]),.doutc(w_asqrt6_16[2]),.din(w_asqrt6_5[0]));
	jspl3 jspl3_w_asqrt6_17(.douta(w_asqrt6_17[0]),.doutb(w_asqrt6_17[1]),.doutc(w_asqrt6_17[2]),.din(w_asqrt6_5[1]));
	jspl3 jspl3_w_asqrt6_18(.douta(w_asqrt6_18[0]),.doutb(w_asqrt6_18[1]),.doutc(w_asqrt6_18[2]),.din(w_asqrt6_5[2]));
	jspl3 jspl3_w_asqrt6_19(.douta(w_asqrt6_19[0]),.doutb(w_asqrt6_19[1]),.doutc(w_asqrt6_19[2]),.din(w_asqrt6_6[0]));
	jspl3 jspl3_w_asqrt6_20(.douta(w_asqrt6_20[0]),.doutb(w_asqrt6_20[1]),.doutc(w_asqrt6_20[2]),.din(w_asqrt6_6[1]));
	jspl3 jspl3_w_asqrt6_21(.douta(w_asqrt6_21[0]),.doutb(w_asqrt6_21[1]),.doutc(w_asqrt6_21[2]),.din(w_asqrt6_6[2]));
	jspl3 jspl3_w_asqrt6_22(.douta(w_asqrt6_22[0]),.doutb(w_asqrt6_22[1]),.doutc(w_asqrt6_22[2]),.din(w_asqrt6_7[0]));
	jspl3 jspl3_w_asqrt6_23(.douta(w_asqrt6_23[0]),.doutb(w_asqrt6_23[1]),.doutc(w_asqrt6_23[2]),.din(w_asqrt6_7[1]));
	jspl3 jspl3_w_asqrt6_24(.douta(w_asqrt6_24[0]),.doutb(w_asqrt6_24[1]),.doutc(w_asqrt6_24[2]),.din(w_asqrt6_7[2]));
	jspl3 jspl3_w_asqrt6_25(.douta(w_asqrt6_25[0]),.doutb(w_asqrt6_25[1]),.doutc(w_asqrt6_25[2]),.din(w_asqrt6_8[0]));
	jspl3 jspl3_w_asqrt6_26(.douta(w_asqrt6_26[0]),.doutb(w_asqrt6_26[1]),.doutc(w_asqrt6_26[2]),.din(w_asqrt6_8[1]));
	jspl3 jspl3_w_asqrt6_27(.douta(w_asqrt6_27[0]),.doutb(w_asqrt6_27[1]),.doutc(w_asqrt6_27[2]),.din(w_asqrt6_8[2]));
	jspl3 jspl3_w_asqrt6_28(.douta(w_asqrt6_28[0]),.doutb(w_asqrt6_28[1]),.doutc(w_asqrt6_28[2]),.din(w_asqrt6_9[0]));
	jspl3 jspl3_w_asqrt6_29(.douta(w_asqrt6_29[0]),.doutb(w_asqrt6_29[1]),.doutc(w_asqrt6_29[2]),.din(w_asqrt6_9[1]));
	jspl3 jspl3_w_asqrt6_30(.douta(w_asqrt6_30[0]),.doutb(w_asqrt6_30[1]),.doutc(w_asqrt6_30[2]),.din(w_asqrt6_9[2]));
	jspl jspl_w_asqrt6_31(.douta(w_asqrt6_31),.doutb(asqrt[5]),.din(w_asqrt6_10[0]));
	jspl3 jspl3_w_asqrt7_0(.douta(w_asqrt7_0[0]),.doutb(w_asqrt7_0[1]),.doutc(w_asqrt7_0[2]),.din(asqrt_fa_7));
	jspl3 jspl3_w_asqrt7_1(.douta(w_asqrt7_1[0]),.doutb(w_asqrt7_1[1]),.doutc(w_asqrt7_1[2]),.din(w_asqrt7_0[0]));
	jspl3 jspl3_w_asqrt7_2(.douta(w_asqrt7_2[0]),.doutb(w_asqrt7_2[1]),.doutc(w_asqrt7_2[2]),.din(w_asqrt7_0[1]));
	jspl3 jspl3_w_asqrt7_3(.douta(w_asqrt7_3[0]),.doutb(w_asqrt7_3[1]),.doutc(w_asqrt7_3[2]),.din(w_asqrt7_0[2]));
	jspl3 jspl3_w_asqrt7_4(.douta(w_asqrt7_4[0]),.doutb(w_asqrt7_4[1]),.doutc(w_asqrt7_4[2]),.din(w_asqrt7_1[0]));
	jspl3 jspl3_w_asqrt7_5(.douta(w_asqrt7_5[0]),.doutb(w_asqrt7_5[1]),.doutc(w_asqrt7_5[2]),.din(w_asqrt7_1[1]));
	jspl3 jspl3_w_asqrt7_6(.douta(w_asqrt7_6[0]),.doutb(w_asqrt7_6[1]),.doutc(w_asqrt7_6[2]),.din(w_asqrt7_1[2]));
	jspl3 jspl3_w_asqrt7_7(.douta(w_asqrt7_7[0]),.doutb(w_asqrt7_7[1]),.doutc(w_asqrt7_7[2]),.din(w_asqrt7_2[0]));
	jspl3 jspl3_w_asqrt7_8(.douta(w_asqrt7_8[0]),.doutb(w_asqrt7_8[1]),.doutc(w_asqrt7_8[2]),.din(w_asqrt7_2[1]));
	jspl3 jspl3_w_asqrt7_9(.douta(w_asqrt7_9[0]),.doutb(w_asqrt7_9[1]),.doutc(w_asqrt7_9[2]),.din(w_asqrt7_2[2]));
	jspl3 jspl3_w_asqrt7_10(.douta(w_asqrt7_10[0]),.doutb(w_asqrt7_10[1]),.doutc(w_asqrt7_10[2]),.din(w_asqrt7_3[0]));
	jspl3 jspl3_w_asqrt7_11(.douta(w_asqrt7_11[0]),.doutb(w_asqrt7_11[1]),.doutc(w_asqrt7_11[2]),.din(w_asqrt7_3[1]));
	jspl3 jspl3_w_asqrt7_12(.douta(w_asqrt7_12[0]),.doutb(w_asqrt7_12[1]),.doutc(w_asqrt7_12[2]),.din(w_asqrt7_3[2]));
	jspl3 jspl3_w_asqrt7_13(.douta(w_asqrt7_13[0]),.doutb(w_asqrt7_13[1]),.doutc(w_asqrt7_13[2]),.din(w_asqrt7_4[0]));
	jspl3 jspl3_w_asqrt7_14(.douta(w_asqrt7_14[0]),.doutb(w_asqrt7_14[1]),.doutc(w_asqrt7_14[2]),.din(w_asqrt7_4[1]));
	jspl jspl_w_asqrt7_15(.douta(w_asqrt7_15),.doutb(asqrt[6]),.din(w_asqrt7_4[2]));
	jspl3 jspl3_w_asqrt8_0(.douta(w_asqrt8_0[0]),.doutb(w_asqrt8_0[1]),.doutc(w_asqrt8_0[2]),.din(asqrt_fa_8));
	jspl3 jspl3_w_asqrt8_1(.douta(w_asqrt8_1[0]),.doutb(w_asqrt8_1[1]),.doutc(w_asqrt8_1[2]),.din(w_asqrt8_0[0]));
	jspl3 jspl3_w_asqrt8_2(.douta(w_asqrt8_2[0]),.doutb(w_asqrt8_2[1]),.doutc(w_asqrt8_2[2]),.din(w_asqrt8_0[1]));
	jspl3 jspl3_w_asqrt8_3(.douta(w_asqrt8_3[0]),.doutb(w_asqrt8_3[1]),.doutc(w_asqrt8_3[2]),.din(w_asqrt8_0[2]));
	jspl3 jspl3_w_asqrt8_4(.douta(w_asqrt8_4[0]),.doutb(w_asqrt8_4[1]),.doutc(w_asqrt8_4[2]),.din(w_asqrt8_1[0]));
	jspl3 jspl3_w_asqrt8_5(.douta(w_asqrt8_5[0]),.doutb(w_asqrt8_5[1]),.doutc(w_asqrt8_5[2]),.din(w_asqrt8_1[1]));
	jspl3 jspl3_w_asqrt8_6(.douta(w_asqrt8_6[0]),.doutb(w_asqrt8_6[1]),.doutc(w_asqrt8_6[2]),.din(w_asqrt8_1[2]));
	jspl3 jspl3_w_asqrt8_7(.douta(w_asqrt8_7[0]),.doutb(w_asqrt8_7[1]),.doutc(w_asqrt8_7[2]),.din(w_asqrt8_2[0]));
	jspl3 jspl3_w_asqrt8_8(.douta(w_asqrt8_8[0]),.doutb(w_asqrt8_8[1]),.doutc(w_asqrt8_8[2]),.din(w_asqrt8_2[1]));
	jspl3 jspl3_w_asqrt8_9(.douta(w_asqrt8_9[0]),.doutb(w_asqrt8_9[1]),.doutc(w_asqrt8_9[2]),.din(w_asqrt8_2[2]));
	jspl3 jspl3_w_asqrt8_10(.douta(w_asqrt8_10[0]),.doutb(w_asqrt8_10[1]),.doutc(w_asqrt8_10[2]),.din(w_asqrt8_3[0]));
	jspl3 jspl3_w_asqrt8_11(.douta(w_asqrt8_11[0]),.doutb(w_asqrt8_11[1]),.doutc(w_asqrt8_11[2]),.din(w_asqrt8_3[1]));
	jspl3 jspl3_w_asqrt8_12(.douta(w_asqrt8_12[0]),.doutb(w_asqrt8_12[1]),.doutc(w_asqrt8_12[2]),.din(w_asqrt8_3[2]));
	jspl3 jspl3_w_asqrt8_13(.douta(w_asqrt8_13[0]),.doutb(w_asqrt8_13[1]),.doutc(w_asqrt8_13[2]),.din(w_asqrt8_4[0]));
	jspl3 jspl3_w_asqrt8_14(.douta(w_asqrt8_14[0]),.doutb(w_asqrt8_14[1]),.doutc(w_asqrt8_14[2]),.din(w_asqrt8_4[1]));
	jspl3 jspl3_w_asqrt8_15(.douta(w_asqrt8_15[0]),.doutb(w_asqrt8_15[1]),.doutc(w_asqrt8_15[2]),.din(w_asqrt8_4[2]));
	jspl3 jspl3_w_asqrt8_16(.douta(w_asqrt8_16[0]),.doutb(w_asqrt8_16[1]),.doutc(w_asqrt8_16[2]),.din(w_asqrt8_5[0]));
	jspl3 jspl3_w_asqrt8_17(.douta(w_asqrt8_17[0]),.doutb(w_asqrt8_17[1]),.doutc(w_asqrt8_17[2]),.din(w_asqrt8_5[1]));
	jspl3 jspl3_w_asqrt8_18(.douta(w_asqrt8_18[0]),.doutb(w_asqrt8_18[1]),.doutc(w_asqrt8_18[2]),.din(w_asqrt8_5[2]));
	jspl3 jspl3_w_asqrt8_19(.douta(w_asqrt8_19[0]),.doutb(w_asqrt8_19[1]),.doutc(w_asqrt8_19[2]),.din(w_asqrt8_6[0]));
	jspl3 jspl3_w_asqrt8_20(.douta(w_asqrt8_20[0]),.doutb(w_asqrt8_20[1]),.doutc(w_asqrt8_20[2]),.din(w_asqrt8_6[1]));
	jspl3 jspl3_w_asqrt8_21(.douta(w_asqrt8_21[0]),.doutb(w_asqrt8_21[1]),.doutc(w_asqrt8_21[2]),.din(w_asqrt8_6[2]));
	jspl3 jspl3_w_asqrt8_22(.douta(w_asqrt8_22[0]),.doutb(w_asqrt8_22[1]),.doutc(w_asqrt8_22[2]),.din(w_asqrt8_7[0]));
	jspl3 jspl3_w_asqrt8_23(.douta(w_asqrt8_23[0]),.doutb(w_asqrt8_23[1]),.doutc(w_asqrt8_23[2]),.din(w_asqrt8_7[1]));
	jspl3 jspl3_w_asqrt8_24(.douta(w_asqrt8_24[0]),.doutb(w_asqrt8_24[1]),.doutc(w_asqrt8_24[2]),.din(w_asqrt8_7[2]));
	jspl3 jspl3_w_asqrt8_25(.douta(w_asqrt8_25[0]),.doutb(w_asqrt8_25[1]),.doutc(w_asqrt8_25[2]),.din(w_asqrt8_8[0]));
	jspl3 jspl3_w_asqrt8_26(.douta(w_asqrt8_26[0]),.doutb(w_asqrt8_26[1]),.doutc(w_asqrt8_26[2]),.din(w_asqrt8_8[1]));
	jspl3 jspl3_w_asqrt8_27(.douta(w_asqrt8_27[0]),.doutb(w_asqrt8_27[1]),.doutc(w_asqrt8_27[2]),.din(w_asqrt8_8[2]));
	jspl3 jspl3_w_asqrt8_28(.douta(w_asqrt8_28[0]),.doutb(w_asqrt8_28[1]),.doutc(w_asqrt8_28[2]),.din(w_asqrt8_9[0]));
	jspl3 jspl3_w_asqrt8_29(.douta(w_asqrt8_29[0]),.doutb(w_asqrt8_29[1]),.doutc(w_asqrt8_29[2]),.din(w_asqrt8_9[1]));
	jspl3 jspl3_w_asqrt8_30(.douta(w_asqrt8_30[0]),.doutb(w_asqrt8_30[1]),.doutc(w_asqrt8_30[2]),.din(w_asqrt8_9[2]));
	jspl jspl_w_asqrt8_31(.douta(w_asqrt8_31),.doutb(asqrt[7]),.din(w_asqrt8_10[0]));
	jspl3 jspl3_w_asqrt9_0(.douta(w_asqrt9_0[0]),.doutb(w_asqrt9_0[1]),.doutc(w_asqrt9_0[2]),.din(asqrt_fa_9));
	jspl3 jspl3_w_asqrt9_1(.douta(w_asqrt9_1[0]),.doutb(w_asqrt9_1[1]),.doutc(w_asqrt9_1[2]),.din(w_asqrt9_0[0]));
	jspl3 jspl3_w_asqrt9_2(.douta(w_asqrt9_2[0]),.doutb(w_asqrt9_2[1]),.doutc(w_asqrt9_2[2]),.din(w_asqrt9_0[1]));
	jspl3 jspl3_w_asqrt9_3(.douta(w_asqrt9_3[0]),.doutb(w_asqrt9_3[1]),.doutc(w_asqrt9_3[2]),.din(w_asqrt9_0[2]));
	jspl3 jspl3_w_asqrt9_4(.douta(w_asqrt9_4[0]),.doutb(w_asqrt9_4[1]),.doutc(w_asqrt9_4[2]),.din(w_asqrt9_1[0]));
	jspl3 jspl3_w_asqrt9_5(.douta(w_asqrt9_5[0]),.doutb(w_asqrt9_5[1]),.doutc(w_asqrt9_5[2]),.din(w_asqrt9_1[1]));
	jspl3 jspl3_w_asqrt9_6(.douta(w_asqrt9_6[0]),.doutb(w_asqrt9_6[1]),.doutc(w_asqrt9_6[2]),.din(w_asqrt9_1[2]));
	jspl3 jspl3_w_asqrt9_7(.douta(w_asqrt9_7[0]),.doutb(w_asqrt9_7[1]),.doutc(w_asqrt9_7[2]),.din(w_asqrt9_2[0]));
	jspl3 jspl3_w_asqrt9_8(.douta(w_asqrt9_8[0]),.doutb(w_asqrt9_8[1]),.doutc(w_asqrt9_8[2]),.din(w_asqrt9_2[1]));
	jspl3 jspl3_w_asqrt9_9(.douta(w_asqrt9_9[0]),.doutb(w_asqrt9_9[1]),.doutc(w_asqrt9_9[2]),.din(w_asqrt9_2[2]));
	jspl3 jspl3_w_asqrt9_10(.douta(w_asqrt9_10[0]),.doutb(w_asqrt9_10[1]),.doutc(w_asqrt9_10[2]),.din(w_asqrt9_3[0]));
	jspl3 jspl3_w_asqrt9_11(.douta(w_asqrt9_11[0]),.doutb(w_asqrt9_11[1]),.doutc(w_asqrt9_11[2]),.din(w_asqrt9_3[1]));
	jspl3 jspl3_w_asqrt9_12(.douta(w_asqrt9_12[0]),.doutb(w_asqrt9_12[1]),.doutc(w_asqrt9_12[2]),.din(w_asqrt9_3[2]));
	jspl3 jspl3_w_asqrt9_13(.douta(w_asqrt9_13[0]),.doutb(w_asqrt9_13[1]),.doutc(w_asqrt9_13[2]),.din(w_asqrt9_4[0]));
	jspl3 jspl3_w_asqrt9_14(.douta(w_asqrt9_14[0]),.doutb(w_asqrt9_14[1]),.doutc(w_asqrt9_14[2]),.din(w_asqrt9_4[1]));
	jspl3 jspl3_w_asqrt9_15(.douta(w_asqrt9_15[0]),.doutb(w_asqrt9_15[1]),.doutc(w_asqrt9_15[2]),.din(w_asqrt9_4[2]));
	jspl jspl_w_asqrt9_16(.douta(w_asqrt9_16),.doutb(asqrt[8]),.din(w_asqrt9_5[0]));
	jspl3 jspl3_w_asqrt10_0(.douta(w_asqrt10_0[0]),.doutb(w_asqrt10_0[1]),.doutc(w_asqrt10_0[2]),.din(asqrt_fa_10));
	jspl3 jspl3_w_asqrt10_1(.douta(w_asqrt10_1[0]),.doutb(w_asqrt10_1[1]),.doutc(w_asqrt10_1[2]),.din(w_asqrt10_0[0]));
	jspl3 jspl3_w_asqrt10_2(.douta(w_asqrt10_2[0]),.doutb(w_asqrt10_2[1]),.doutc(w_asqrt10_2[2]),.din(w_asqrt10_0[1]));
	jspl3 jspl3_w_asqrt10_3(.douta(w_asqrt10_3[0]),.doutb(w_asqrt10_3[1]),.doutc(w_asqrt10_3[2]),.din(w_asqrt10_0[2]));
	jspl3 jspl3_w_asqrt10_4(.douta(w_asqrt10_4[0]),.doutb(w_asqrt10_4[1]),.doutc(w_asqrt10_4[2]),.din(w_asqrt10_1[0]));
	jspl3 jspl3_w_asqrt10_5(.douta(w_asqrt10_5[0]),.doutb(w_asqrt10_5[1]),.doutc(w_asqrt10_5[2]),.din(w_asqrt10_1[1]));
	jspl3 jspl3_w_asqrt10_6(.douta(w_asqrt10_6[0]),.doutb(w_asqrt10_6[1]),.doutc(w_asqrt10_6[2]),.din(w_asqrt10_1[2]));
	jspl3 jspl3_w_asqrt10_7(.douta(w_asqrt10_7[0]),.doutb(w_asqrt10_7[1]),.doutc(w_asqrt10_7[2]),.din(w_asqrt10_2[0]));
	jspl3 jspl3_w_asqrt10_8(.douta(w_asqrt10_8[0]),.doutb(w_asqrt10_8[1]),.doutc(w_asqrt10_8[2]),.din(w_asqrt10_2[1]));
	jspl3 jspl3_w_asqrt10_9(.douta(w_asqrt10_9[0]),.doutb(w_asqrt10_9[1]),.doutc(w_asqrt10_9[2]),.din(w_asqrt10_2[2]));
	jspl3 jspl3_w_asqrt10_10(.douta(w_asqrt10_10[0]),.doutb(w_asqrt10_10[1]),.doutc(w_asqrt10_10[2]),.din(w_asqrt10_3[0]));
	jspl3 jspl3_w_asqrt10_11(.douta(w_asqrt10_11[0]),.doutb(w_asqrt10_11[1]),.doutc(w_asqrt10_11[2]),.din(w_asqrt10_3[1]));
	jspl3 jspl3_w_asqrt10_12(.douta(w_asqrt10_12[0]),.doutb(w_asqrt10_12[1]),.doutc(w_asqrt10_12[2]),.din(w_asqrt10_3[2]));
	jspl3 jspl3_w_asqrt10_13(.douta(w_asqrt10_13[0]),.doutb(w_asqrt10_13[1]),.doutc(w_asqrt10_13[2]),.din(w_asqrt10_4[0]));
	jspl3 jspl3_w_asqrt10_14(.douta(w_asqrt10_14[0]),.doutb(w_asqrt10_14[1]),.doutc(w_asqrt10_14[2]),.din(w_asqrt10_4[1]));
	jspl3 jspl3_w_asqrt10_15(.douta(w_asqrt10_15[0]),.doutb(w_asqrt10_15[1]),.doutc(w_asqrt10_15[2]),.din(w_asqrt10_4[2]));
	jspl3 jspl3_w_asqrt10_16(.douta(w_asqrt10_16[0]),.doutb(w_asqrt10_16[1]),.doutc(w_asqrt10_16[2]),.din(w_asqrt10_5[0]));
	jspl3 jspl3_w_asqrt10_17(.douta(w_asqrt10_17[0]),.doutb(w_asqrt10_17[1]),.doutc(w_asqrt10_17[2]),.din(w_asqrt10_5[1]));
	jspl3 jspl3_w_asqrt10_18(.douta(w_asqrt10_18[0]),.doutb(w_asqrt10_18[1]),.doutc(w_asqrt10_18[2]),.din(w_asqrt10_5[2]));
	jspl3 jspl3_w_asqrt10_19(.douta(w_asqrt10_19[0]),.doutb(w_asqrt10_19[1]),.doutc(w_asqrt10_19[2]),.din(w_asqrt10_6[0]));
	jspl3 jspl3_w_asqrt10_20(.douta(w_asqrt10_20[0]),.doutb(w_asqrt10_20[1]),.doutc(w_asqrt10_20[2]),.din(w_asqrt10_6[1]));
	jspl3 jspl3_w_asqrt10_21(.douta(w_asqrt10_21[0]),.doutb(w_asqrt10_21[1]),.doutc(w_asqrt10_21[2]),.din(w_asqrt10_6[2]));
	jspl3 jspl3_w_asqrt10_22(.douta(w_asqrt10_22[0]),.doutb(w_asqrt10_22[1]),.doutc(w_asqrt10_22[2]),.din(w_asqrt10_7[0]));
	jspl3 jspl3_w_asqrt10_23(.douta(w_asqrt10_23[0]),.doutb(w_asqrt10_23[1]),.doutc(w_asqrt10_23[2]),.din(w_asqrt10_7[1]));
	jspl3 jspl3_w_asqrt10_24(.douta(w_asqrt10_24[0]),.doutb(w_asqrt10_24[1]),.doutc(w_asqrt10_24[2]),.din(w_asqrt10_7[2]));
	jspl3 jspl3_w_asqrt10_25(.douta(w_asqrt10_25[0]),.doutb(w_asqrt10_25[1]),.doutc(w_asqrt10_25[2]),.din(w_asqrt10_8[0]));
	jspl3 jspl3_w_asqrt10_26(.douta(w_asqrt10_26[0]),.doutb(w_asqrt10_26[1]),.doutc(w_asqrt10_26[2]),.din(w_asqrt10_8[1]));
	jspl3 jspl3_w_asqrt10_27(.douta(w_asqrt10_27[0]),.doutb(w_asqrt10_27[1]),.doutc(w_asqrt10_27[2]),.din(w_asqrt10_8[2]));
	jspl3 jspl3_w_asqrt10_28(.douta(w_asqrt10_28[0]),.doutb(w_asqrt10_28[1]),.doutc(w_asqrt10_28[2]),.din(w_asqrt10_9[0]));
	jspl3 jspl3_w_asqrt10_29(.douta(w_asqrt10_29[0]),.doutb(w_asqrt10_29[1]),.doutc(w_asqrt10_29[2]),.din(w_asqrt10_9[1]));
	jspl3 jspl3_w_asqrt10_30(.douta(w_asqrt10_30[0]),.doutb(w_asqrt10_30[1]),.doutc(w_asqrt10_30[2]),.din(w_asqrt10_9[2]));
	jspl jspl_w_asqrt10_31(.douta(w_asqrt10_31),.doutb(asqrt[9]),.din(w_asqrt10_10[0]));
	jspl3 jspl3_w_asqrt11_0(.douta(w_asqrt11_0[0]),.doutb(w_asqrt11_0[1]),.doutc(w_asqrt11_0[2]),.din(asqrt_fa_11));
	jspl3 jspl3_w_asqrt11_1(.douta(w_asqrt11_1[0]),.doutb(w_asqrt11_1[1]),.doutc(w_asqrt11_1[2]),.din(w_asqrt11_0[0]));
	jspl3 jspl3_w_asqrt11_2(.douta(w_asqrt11_2[0]),.doutb(w_asqrt11_2[1]),.doutc(w_asqrt11_2[2]),.din(w_asqrt11_0[1]));
	jspl3 jspl3_w_asqrt11_3(.douta(w_asqrt11_3[0]),.doutb(w_asqrt11_3[1]),.doutc(w_asqrt11_3[2]),.din(w_asqrt11_0[2]));
	jspl3 jspl3_w_asqrt11_4(.douta(w_asqrt11_4[0]),.doutb(w_asqrt11_4[1]),.doutc(w_asqrt11_4[2]),.din(w_asqrt11_1[0]));
	jspl3 jspl3_w_asqrt11_5(.douta(w_asqrt11_5[0]),.doutb(w_asqrt11_5[1]),.doutc(w_asqrt11_5[2]),.din(w_asqrt11_1[1]));
	jspl3 jspl3_w_asqrt11_6(.douta(w_asqrt11_6[0]),.doutb(w_asqrt11_6[1]),.doutc(w_asqrt11_6[2]),.din(w_asqrt11_1[2]));
	jspl3 jspl3_w_asqrt11_7(.douta(w_asqrt11_7[0]),.doutb(w_asqrt11_7[1]),.doutc(w_asqrt11_7[2]),.din(w_asqrt11_2[0]));
	jspl3 jspl3_w_asqrt11_8(.douta(w_asqrt11_8[0]),.doutb(w_asqrt11_8[1]),.doutc(w_asqrt11_8[2]),.din(w_asqrt11_2[1]));
	jspl3 jspl3_w_asqrt11_9(.douta(w_asqrt11_9[0]),.doutb(w_asqrt11_9[1]),.doutc(w_asqrt11_9[2]),.din(w_asqrt11_2[2]));
	jspl3 jspl3_w_asqrt11_10(.douta(w_asqrt11_10[0]),.doutb(w_asqrt11_10[1]),.doutc(w_asqrt11_10[2]),.din(w_asqrt11_3[0]));
	jspl3 jspl3_w_asqrt11_11(.douta(w_asqrt11_11[0]),.doutb(w_asqrt11_11[1]),.doutc(w_asqrt11_11[2]),.din(w_asqrt11_3[1]));
	jspl3 jspl3_w_asqrt11_12(.douta(w_asqrt11_12[0]),.doutb(w_asqrt11_12[1]),.doutc(w_asqrt11_12[2]),.din(w_asqrt11_3[2]));
	jspl3 jspl3_w_asqrt11_13(.douta(w_asqrt11_13[0]),.doutb(w_asqrt11_13[1]),.doutc(w_asqrt11_13[2]),.din(w_asqrt11_4[0]));
	jspl3 jspl3_w_asqrt11_14(.douta(w_asqrt11_14[0]),.doutb(w_asqrt11_14[1]),.doutc(w_asqrt11_14[2]),.din(w_asqrt11_4[1]));
	jspl3 jspl3_w_asqrt11_15(.douta(w_asqrt11_15[0]),.doutb(w_asqrt11_15[1]),.doutc(w_asqrt11_15[2]),.din(w_asqrt11_4[2]));
	jspl jspl_w_asqrt11_16(.douta(w_asqrt11_16),.doutb(asqrt[10]),.din(w_asqrt11_5[0]));
	jspl3 jspl3_w_asqrt12_0(.douta(w_asqrt12_0[0]),.doutb(w_asqrt12_0[1]),.doutc(w_asqrt12_0[2]),.din(asqrt_fa_12));
	jspl3 jspl3_w_asqrt12_1(.douta(w_asqrt12_1[0]),.doutb(w_asqrt12_1[1]),.doutc(w_asqrt12_1[2]),.din(w_asqrt12_0[0]));
	jspl3 jspl3_w_asqrt12_2(.douta(w_asqrt12_2[0]),.doutb(w_asqrt12_2[1]),.doutc(w_asqrt12_2[2]),.din(w_asqrt12_0[1]));
	jspl3 jspl3_w_asqrt12_3(.douta(w_asqrt12_3[0]),.doutb(w_asqrt12_3[1]),.doutc(w_asqrt12_3[2]),.din(w_asqrt12_0[2]));
	jspl3 jspl3_w_asqrt12_4(.douta(w_asqrt12_4[0]),.doutb(w_asqrt12_4[1]),.doutc(w_asqrt12_4[2]),.din(w_asqrt12_1[0]));
	jspl3 jspl3_w_asqrt12_5(.douta(w_asqrt12_5[0]),.doutb(w_asqrt12_5[1]),.doutc(w_asqrt12_5[2]),.din(w_asqrt12_1[1]));
	jspl3 jspl3_w_asqrt12_6(.douta(w_asqrt12_6[0]),.doutb(w_asqrt12_6[1]),.doutc(w_asqrt12_6[2]),.din(w_asqrt12_1[2]));
	jspl3 jspl3_w_asqrt12_7(.douta(w_asqrt12_7[0]),.doutb(w_asqrt12_7[1]),.doutc(w_asqrt12_7[2]),.din(w_asqrt12_2[0]));
	jspl3 jspl3_w_asqrt12_8(.douta(w_asqrt12_8[0]),.doutb(w_asqrt12_8[1]),.doutc(w_asqrt12_8[2]),.din(w_asqrt12_2[1]));
	jspl3 jspl3_w_asqrt12_9(.douta(w_asqrt12_9[0]),.doutb(w_asqrt12_9[1]),.doutc(w_asqrt12_9[2]),.din(w_asqrt12_2[2]));
	jspl3 jspl3_w_asqrt12_10(.douta(w_asqrt12_10[0]),.doutb(w_asqrt12_10[1]),.doutc(w_asqrt12_10[2]),.din(w_asqrt12_3[0]));
	jspl3 jspl3_w_asqrt12_11(.douta(w_asqrt12_11[0]),.doutb(w_asqrt12_11[1]),.doutc(w_asqrt12_11[2]),.din(w_asqrt12_3[1]));
	jspl3 jspl3_w_asqrt12_12(.douta(w_asqrt12_12[0]),.doutb(w_asqrt12_12[1]),.doutc(w_asqrt12_12[2]),.din(w_asqrt12_3[2]));
	jspl3 jspl3_w_asqrt12_13(.douta(w_asqrt12_13[0]),.doutb(w_asqrt12_13[1]),.doutc(w_asqrt12_13[2]),.din(w_asqrt12_4[0]));
	jspl3 jspl3_w_asqrt12_14(.douta(w_asqrt12_14[0]),.doutb(w_asqrt12_14[1]),.doutc(w_asqrt12_14[2]),.din(w_asqrt12_4[1]));
	jspl3 jspl3_w_asqrt12_15(.douta(w_asqrt12_15[0]),.doutb(w_asqrt12_15[1]),.doutc(w_asqrt12_15[2]),.din(w_asqrt12_4[2]));
	jspl3 jspl3_w_asqrt12_16(.douta(w_asqrt12_16[0]),.doutb(w_asqrt12_16[1]),.doutc(w_asqrt12_16[2]),.din(w_asqrt12_5[0]));
	jspl3 jspl3_w_asqrt12_17(.douta(w_asqrt12_17[0]),.doutb(w_asqrt12_17[1]),.doutc(w_asqrt12_17[2]),.din(w_asqrt12_5[1]));
	jspl3 jspl3_w_asqrt12_18(.douta(w_asqrt12_18[0]),.doutb(w_asqrt12_18[1]),.doutc(w_asqrt12_18[2]),.din(w_asqrt12_5[2]));
	jspl3 jspl3_w_asqrt12_19(.douta(w_asqrt12_19[0]),.doutb(w_asqrt12_19[1]),.doutc(w_asqrt12_19[2]),.din(w_asqrt12_6[0]));
	jspl3 jspl3_w_asqrt12_20(.douta(w_asqrt12_20[0]),.doutb(w_asqrt12_20[1]),.doutc(w_asqrt12_20[2]),.din(w_asqrt12_6[1]));
	jspl3 jspl3_w_asqrt12_21(.douta(w_asqrt12_21[0]),.doutb(w_asqrt12_21[1]),.doutc(w_asqrt12_21[2]),.din(w_asqrt12_6[2]));
	jspl3 jspl3_w_asqrt12_22(.douta(w_asqrt12_22[0]),.doutb(w_asqrt12_22[1]),.doutc(w_asqrt12_22[2]),.din(w_asqrt12_7[0]));
	jspl3 jspl3_w_asqrt12_23(.douta(w_asqrt12_23[0]),.doutb(w_asqrt12_23[1]),.doutc(w_asqrt12_23[2]),.din(w_asqrt12_7[1]));
	jspl3 jspl3_w_asqrt12_24(.douta(w_asqrt12_24[0]),.doutb(w_asqrt12_24[1]),.doutc(w_asqrt12_24[2]),.din(w_asqrt12_7[2]));
	jspl3 jspl3_w_asqrt12_25(.douta(w_asqrt12_25[0]),.doutb(w_asqrt12_25[1]),.doutc(w_asqrt12_25[2]),.din(w_asqrt12_8[0]));
	jspl3 jspl3_w_asqrt12_26(.douta(w_asqrt12_26[0]),.doutb(w_asqrt12_26[1]),.doutc(w_asqrt12_26[2]),.din(w_asqrt12_8[1]));
	jspl3 jspl3_w_asqrt12_27(.douta(w_asqrt12_27[0]),.doutb(w_asqrt12_27[1]),.doutc(w_asqrt12_27[2]),.din(w_asqrt12_8[2]));
	jspl3 jspl3_w_asqrt12_28(.douta(w_asqrt12_28[0]),.doutb(w_asqrt12_28[1]),.doutc(w_asqrt12_28[2]),.din(w_asqrt12_9[0]));
	jspl3 jspl3_w_asqrt12_29(.douta(w_asqrt12_29[0]),.doutb(w_asqrt12_29[1]),.doutc(w_asqrt12_29[2]),.din(w_asqrt12_9[1]));
	jspl3 jspl3_w_asqrt12_30(.douta(w_asqrt12_30[0]),.doutb(w_asqrt12_30[1]),.doutc(w_asqrt12_30[2]),.din(w_asqrt12_9[2]));
	jspl jspl_w_asqrt12_31(.douta(w_asqrt12_31),.doutb(asqrt[11]),.din(w_asqrt12_10[0]));
	jspl3 jspl3_w_asqrt13_0(.douta(w_asqrt13_0[0]),.doutb(w_asqrt13_0[1]),.doutc(w_asqrt13_0[2]),.din(asqrt_fa_13));
	jspl3 jspl3_w_asqrt13_1(.douta(w_asqrt13_1[0]),.doutb(w_asqrt13_1[1]),.doutc(w_asqrt13_1[2]),.din(w_asqrt13_0[0]));
	jspl3 jspl3_w_asqrt13_2(.douta(w_asqrt13_2[0]),.doutb(w_asqrt13_2[1]),.doutc(w_asqrt13_2[2]),.din(w_asqrt13_0[1]));
	jspl3 jspl3_w_asqrt13_3(.douta(w_asqrt13_3[0]),.doutb(w_asqrt13_3[1]),.doutc(w_asqrt13_3[2]),.din(w_asqrt13_0[2]));
	jspl3 jspl3_w_asqrt13_4(.douta(w_asqrt13_4[0]),.doutb(w_asqrt13_4[1]),.doutc(w_asqrt13_4[2]),.din(w_asqrt13_1[0]));
	jspl3 jspl3_w_asqrt13_5(.douta(w_asqrt13_5[0]),.doutb(w_asqrt13_5[1]),.doutc(w_asqrt13_5[2]),.din(w_asqrt13_1[1]));
	jspl3 jspl3_w_asqrt13_6(.douta(w_asqrt13_6[0]),.doutb(w_asqrt13_6[1]),.doutc(w_asqrt13_6[2]),.din(w_asqrt13_1[2]));
	jspl3 jspl3_w_asqrt13_7(.douta(w_asqrt13_7[0]),.doutb(w_asqrt13_7[1]),.doutc(w_asqrt13_7[2]),.din(w_asqrt13_2[0]));
	jspl3 jspl3_w_asqrt13_8(.douta(w_asqrt13_8[0]),.doutb(w_asqrt13_8[1]),.doutc(w_asqrt13_8[2]),.din(w_asqrt13_2[1]));
	jspl3 jspl3_w_asqrt13_9(.douta(w_asqrt13_9[0]),.doutb(w_asqrt13_9[1]),.doutc(w_asqrt13_9[2]),.din(w_asqrt13_2[2]));
	jspl3 jspl3_w_asqrt13_10(.douta(w_asqrt13_10[0]),.doutb(w_asqrt13_10[1]),.doutc(w_asqrt13_10[2]),.din(w_asqrt13_3[0]));
	jspl3 jspl3_w_asqrt13_11(.douta(w_asqrt13_11[0]),.doutb(w_asqrt13_11[1]),.doutc(w_asqrt13_11[2]),.din(w_asqrt13_3[1]));
	jspl3 jspl3_w_asqrt13_12(.douta(w_asqrt13_12[0]),.doutb(w_asqrt13_12[1]),.doutc(w_asqrt13_12[2]),.din(w_asqrt13_3[2]));
	jspl3 jspl3_w_asqrt13_13(.douta(w_asqrt13_13[0]),.doutb(w_asqrt13_13[1]),.doutc(w_asqrt13_13[2]),.din(w_asqrt13_4[0]));
	jspl3 jspl3_w_asqrt13_14(.douta(w_asqrt13_14[0]),.doutb(w_asqrt13_14[1]),.doutc(w_asqrt13_14[2]),.din(w_asqrt13_4[1]));
	jspl3 jspl3_w_asqrt13_15(.douta(w_asqrt13_15[0]),.doutb(w_asqrt13_15[1]),.doutc(w_asqrt13_15[2]),.din(w_asqrt13_4[2]));
	jspl3 jspl3_w_asqrt13_16(.douta(w_asqrt13_16[0]),.doutb(w_asqrt13_16[1]),.doutc(w_asqrt13_16[2]),.din(w_asqrt13_5[0]));
	jspl jspl_w_asqrt13_17(.douta(w_asqrt13_17),.doutb(asqrt[12]),.din(w_asqrt13_5[1]));
	jspl3 jspl3_w_asqrt14_0(.douta(w_asqrt14_0[0]),.doutb(w_asqrt14_0[1]),.doutc(w_asqrt14_0[2]),.din(asqrt_fa_14));
	jspl3 jspl3_w_asqrt14_1(.douta(w_asqrt14_1[0]),.doutb(w_asqrt14_1[1]),.doutc(w_asqrt14_1[2]),.din(w_asqrt14_0[0]));
	jspl3 jspl3_w_asqrt14_2(.douta(w_asqrt14_2[0]),.doutb(w_asqrt14_2[1]),.doutc(w_asqrt14_2[2]),.din(w_asqrt14_0[1]));
	jspl3 jspl3_w_asqrt14_3(.douta(w_asqrt14_3[0]),.doutb(w_asqrt14_3[1]),.doutc(w_asqrt14_3[2]),.din(w_asqrt14_0[2]));
	jspl3 jspl3_w_asqrt14_4(.douta(w_asqrt14_4[0]),.doutb(w_asqrt14_4[1]),.doutc(w_asqrt14_4[2]),.din(w_asqrt14_1[0]));
	jspl3 jspl3_w_asqrt14_5(.douta(w_asqrt14_5[0]),.doutb(w_asqrt14_5[1]),.doutc(w_asqrt14_5[2]),.din(w_asqrt14_1[1]));
	jspl3 jspl3_w_asqrt14_6(.douta(w_asqrt14_6[0]),.doutb(w_asqrt14_6[1]),.doutc(w_asqrt14_6[2]),.din(w_asqrt14_1[2]));
	jspl3 jspl3_w_asqrt14_7(.douta(w_asqrt14_7[0]),.doutb(w_asqrt14_7[1]),.doutc(w_asqrt14_7[2]),.din(w_asqrt14_2[0]));
	jspl3 jspl3_w_asqrt14_8(.douta(w_asqrt14_8[0]),.doutb(w_asqrt14_8[1]),.doutc(w_asqrt14_8[2]),.din(w_asqrt14_2[1]));
	jspl3 jspl3_w_asqrt14_9(.douta(w_asqrt14_9[0]),.doutb(w_asqrt14_9[1]),.doutc(w_asqrt14_9[2]),.din(w_asqrt14_2[2]));
	jspl3 jspl3_w_asqrt14_10(.douta(w_asqrt14_10[0]),.doutb(w_asqrt14_10[1]),.doutc(w_asqrt14_10[2]),.din(w_asqrt14_3[0]));
	jspl3 jspl3_w_asqrt14_11(.douta(w_asqrt14_11[0]),.doutb(w_asqrt14_11[1]),.doutc(w_asqrt14_11[2]),.din(w_asqrt14_3[1]));
	jspl3 jspl3_w_asqrt14_12(.douta(w_asqrt14_12[0]),.doutb(w_asqrt14_12[1]),.doutc(w_asqrt14_12[2]),.din(w_asqrt14_3[2]));
	jspl3 jspl3_w_asqrt14_13(.douta(w_asqrt14_13[0]),.doutb(w_asqrt14_13[1]),.doutc(w_asqrt14_13[2]),.din(w_asqrt14_4[0]));
	jspl3 jspl3_w_asqrt14_14(.douta(w_asqrt14_14[0]),.doutb(w_asqrt14_14[1]),.doutc(w_asqrt14_14[2]),.din(w_asqrt14_4[1]));
	jspl3 jspl3_w_asqrt14_15(.douta(w_asqrt14_15[0]),.doutb(w_asqrt14_15[1]),.doutc(w_asqrt14_15[2]),.din(w_asqrt14_4[2]));
	jspl3 jspl3_w_asqrt14_16(.douta(w_asqrt14_16[0]),.doutb(w_asqrt14_16[1]),.doutc(w_asqrt14_16[2]),.din(w_asqrt14_5[0]));
	jspl3 jspl3_w_asqrt14_17(.douta(w_asqrt14_17[0]),.doutb(w_asqrt14_17[1]),.doutc(w_asqrt14_17[2]),.din(w_asqrt14_5[1]));
	jspl3 jspl3_w_asqrt14_18(.douta(w_asqrt14_18[0]),.doutb(w_asqrt14_18[1]),.doutc(w_asqrt14_18[2]),.din(w_asqrt14_5[2]));
	jspl3 jspl3_w_asqrt14_19(.douta(w_asqrt14_19[0]),.doutb(w_asqrt14_19[1]),.doutc(w_asqrt14_19[2]),.din(w_asqrt14_6[0]));
	jspl3 jspl3_w_asqrt14_20(.douta(w_asqrt14_20[0]),.doutb(w_asqrt14_20[1]),.doutc(w_asqrt14_20[2]),.din(w_asqrt14_6[1]));
	jspl3 jspl3_w_asqrt14_21(.douta(w_asqrt14_21[0]),.doutb(w_asqrt14_21[1]),.doutc(w_asqrt14_21[2]),.din(w_asqrt14_6[2]));
	jspl3 jspl3_w_asqrt14_22(.douta(w_asqrt14_22[0]),.doutb(w_asqrt14_22[1]),.doutc(w_asqrt14_22[2]),.din(w_asqrt14_7[0]));
	jspl3 jspl3_w_asqrt14_23(.douta(w_asqrt14_23[0]),.doutb(w_asqrt14_23[1]),.doutc(w_asqrt14_23[2]),.din(w_asqrt14_7[1]));
	jspl3 jspl3_w_asqrt14_24(.douta(w_asqrt14_24[0]),.doutb(w_asqrt14_24[1]),.doutc(w_asqrt14_24[2]),.din(w_asqrt14_7[2]));
	jspl3 jspl3_w_asqrt14_25(.douta(w_asqrt14_25[0]),.doutb(w_asqrt14_25[1]),.doutc(w_asqrt14_25[2]),.din(w_asqrt14_8[0]));
	jspl3 jspl3_w_asqrt14_26(.douta(w_asqrt14_26[0]),.doutb(w_asqrt14_26[1]),.doutc(w_asqrt14_26[2]),.din(w_asqrt14_8[1]));
	jspl3 jspl3_w_asqrt14_27(.douta(w_asqrt14_27[0]),.doutb(w_asqrt14_27[1]),.doutc(w_asqrt14_27[2]),.din(w_asqrt14_8[2]));
	jspl3 jspl3_w_asqrt14_28(.douta(w_asqrt14_28[0]),.doutb(w_asqrt14_28[1]),.doutc(w_asqrt14_28[2]),.din(w_asqrt14_9[0]));
	jspl3 jspl3_w_asqrt14_29(.douta(w_asqrt14_29[0]),.doutb(w_asqrt14_29[1]),.doutc(w_asqrt14_29[2]),.din(w_asqrt14_9[1]));
	jspl3 jspl3_w_asqrt14_30(.douta(w_asqrt14_30[0]),.doutb(w_asqrt14_30[1]),.doutc(w_asqrt14_30[2]),.din(w_asqrt14_9[2]));
	jspl jspl_w_asqrt14_31(.douta(w_asqrt14_31),.doutb(asqrt[13]),.din(w_asqrt14_10[0]));
	jspl3 jspl3_w_asqrt15_0(.douta(w_asqrt15_0[0]),.doutb(w_asqrt15_0[1]),.doutc(w_asqrt15_0[2]),.din(asqrt_fa_15));
	jspl3 jspl3_w_asqrt15_1(.douta(w_asqrt15_1[0]),.doutb(w_asqrt15_1[1]),.doutc(w_asqrt15_1[2]),.din(w_asqrt15_0[0]));
	jspl3 jspl3_w_asqrt15_2(.douta(w_asqrt15_2[0]),.doutb(w_asqrt15_2[1]),.doutc(w_asqrt15_2[2]),.din(w_asqrt15_0[1]));
	jspl3 jspl3_w_asqrt15_3(.douta(w_asqrt15_3[0]),.doutb(w_asqrt15_3[1]),.doutc(w_asqrt15_3[2]),.din(w_asqrt15_0[2]));
	jspl3 jspl3_w_asqrt15_4(.douta(w_asqrt15_4[0]),.doutb(w_asqrt15_4[1]),.doutc(w_asqrt15_4[2]),.din(w_asqrt15_1[0]));
	jspl3 jspl3_w_asqrt15_5(.douta(w_asqrt15_5[0]),.doutb(w_asqrt15_5[1]),.doutc(w_asqrt15_5[2]),.din(w_asqrt15_1[1]));
	jspl3 jspl3_w_asqrt15_6(.douta(w_asqrt15_6[0]),.doutb(w_asqrt15_6[1]),.doutc(w_asqrt15_6[2]),.din(w_asqrt15_1[2]));
	jspl3 jspl3_w_asqrt15_7(.douta(w_asqrt15_7[0]),.doutb(w_asqrt15_7[1]),.doutc(w_asqrt15_7[2]),.din(w_asqrt15_2[0]));
	jspl3 jspl3_w_asqrt15_8(.douta(w_asqrt15_8[0]),.doutb(w_asqrt15_8[1]),.doutc(w_asqrt15_8[2]),.din(w_asqrt15_2[1]));
	jspl3 jspl3_w_asqrt15_9(.douta(w_asqrt15_9[0]),.doutb(w_asqrt15_9[1]),.doutc(w_asqrt15_9[2]),.din(w_asqrt15_2[2]));
	jspl3 jspl3_w_asqrt15_10(.douta(w_asqrt15_10[0]),.doutb(w_asqrt15_10[1]),.doutc(w_asqrt15_10[2]),.din(w_asqrt15_3[0]));
	jspl3 jspl3_w_asqrt15_11(.douta(w_asqrt15_11[0]),.doutb(w_asqrt15_11[1]),.doutc(w_asqrt15_11[2]),.din(w_asqrt15_3[1]));
	jspl3 jspl3_w_asqrt15_12(.douta(w_asqrt15_12[0]),.doutb(w_asqrt15_12[1]),.doutc(w_asqrt15_12[2]),.din(w_asqrt15_3[2]));
	jspl3 jspl3_w_asqrt15_13(.douta(w_asqrt15_13[0]),.doutb(w_asqrt15_13[1]),.doutc(w_asqrt15_13[2]),.din(w_asqrt15_4[0]));
	jspl3 jspl3_w_asqrt15_14(.douta(w_asqrt15_14[0]),.doutb(w_asqrt15_14[1]),.doutc(w_asqrt15_14[2]),.din(w_asqrt15_4[1]));
	jspl3 jspl3_w_asqrt15_15(.douta(w_asqrt15_15[0]),.doutb(w_asqrt15_15[1]),.doutc(w_asqrt15_15[2]),.din(w_asqrt15_4[2]));
	jspl3 jspl3_w_asqrt15_16(.douta(w_asqrt15_16[0]),.doutb(w_asqrt15_16[1]),.doutc(w_asqrt15_16[2]),.din(w_asqrt15_5[0]));
	jspl jspl_w_asqrt15_17(.douta(w_asqrt15_17),.doutb(asqrt[14]),.din(w_asqrt15_5[1]));
	jspl3 jspl3_w_asqrt16_0(.douta(w_asqrt16_0[0]),.doutb(w_asqrt16_0[1]),.doutc(w_asqrt16_0[2]),.din(asqrt_fa_16));
	jspl3 jspl3_w_asqrt16_1(.douta(w_asqrt16_1[0]),.doutb(w_asqrt16_1[1]),.doutc(w_asqrt16_1[2]),.din(w_asqrt16_0[0]));
	jspl3 jspl3_w_asqrt16_2(.douta(w_asqrt16_2[0]),.doutb(w_asqrt16_2[1]),.doutc(w_asqrt16_2[2]),.din(w_asqrt16_0[1]));
	jspl3 jspl3_w_asqrt16_3(.douta(w_asqrt16_3[0]),.doutb(w_asqrt16_3[1]),.doutc(w_asqrt16_3[2]),.din(w_asqrt16_0[2]));
	jspl3 jspl3_w_asqrt16_4(.douta(w_asqrt16_4[0]),.doutb(w_asqrt16_4[1]),.doutc(w_asqrt16_4[2]),.din(w_asqrt16_1[0]));
	jspl3 jspl3_w_asqrt16_5(.douta(w_asqrt16_5[0]),.doutb(w_asqrt16_5[1]),.doutc(w_asqrt16_5[2]),.din(w_asqrt16_1[1]));
	jspl3 jspl3_w_asqrt16_6(.douta(w_asqrt16_6[0]),.doutb(w_asqrt16_6[1]),.doutc(w_asqrt16_6[2]),.din(w_asqrt16_1[2]));
	jspl3 jspl3_w_asqrt16_7(.douta(w_asqrt16_7[0]),.doutb(w_asqrt16_7[1]),.doutc(w_asqrt16_7[2]),.din(w_asqrt16_2[0]));
	jspl3 jspl3_w_asqrt16_8(.douta(w_asqrt16_8[0]),.doutb(w_asqrt16_8[1]),.doutc(w_asqrt16_8[2]),.din(w_asqrt16_2[1]));
	jspl3 jspl3_w_asqrt16_9(.douta(w_asqrt16_9[0]),.doutb(w_asqrt16_9[1]),.doutc(w_asqrt16_9[2]),.din(w_asqrt16_2[2]));
	jspl3 jspl3_w_asqrt16_10(.douta(w_asqrt16_10[0]),.doutb(w_asqrt16_10[1]),.doutc(w_asqrt16_10[2]),.din(w_asqrt16_3[0]));
	jspl3 jspl3_w_asqrt16_11(.douta(w_asqrt16_11[0]),.doutb(w_asqrt16_11[1]),.doutc(w_asqrt16_11[2]),.din(w_asqrt16_3[1]));
	jspl3 jspl3_w_asqrt16_12(.douta(w_asqrt16_12[0]),.doutb(w_asqrt16_12[1]),.doutc(w_asqrt16_12[2]),.din(w_asqrt16_3[2]));
	jspl3 jspl3_w_asqrt16_13(.douta(w_asqrt16_13[0]),.doutb(w_asqrt16_13[1]),.doutc(w_asqrt16_13[2]),.din(w_asqrt16_4[0]));
	jspl3 jspl3_w_asqrt16_14(.douta(w_asqrt16_14[0]),.doutb(w_asqrt16_14[1]),.doutc(w_asqrt16_14[2]),.din(w_asqrt16_4[1]));
	jspl3 jspl3_w_asqrt16_15(.douta(w_asqrt16_15[0]),.doutb(w_asqrt16_15[1]),.doutc(w_asqrt16_15[2]),.din(w_asqrt16_4[2]));
	jspl3 jspl3_w_asqrt16_16(.douta(w_asqrt16_16[0]),.doutb(w_asqrt16_16[1]),.doutc(w_asqrt16_16[2]),.din(w_asqrt16_5[0]));
	jspl3 jspl3_w_asqrt16_17(.douta(w_asqrt16_17[0]),.doutb(w_asqrt16_17[1]),.doutc(w_asqrt16_17[2]),.din(w_asqrt16_5[1]));
	jspl3 jspl3_w_asqrt16_18(.douta(w_asqrt16_18[0]),.doutb(w_asqrt16_18[1]),.doutc(w_asqrt16_18[2]),.din(w_asqrt16_5[2]));
	jspl3 jspl3_w_asqrt16_19(.douta(w_asqrt16_19[0]),.doutb(w_asqrt16_19[1]),.doutc(w_asqrt16_19[2]),.din(w_asqrt16_6[0]));
	jspl3 jspl3_w_asqrt16_20(.douta(w_asqrt16_20[0]),.doutb(w_asqrt16_20[1]),.doutc(w_asqrt16_20[2]),.din(w_asqrt16_6[1]));
	jspl3 jspl3_w_asqrt16_21(.douta(w_asqrt16_21[0]),.doutb(w_asqrt16_21[1]),.doutc(w_asqrt16_21[2]),.din(w_asqrt16_6[2]));
	jspl3 jspl3_w_asqrt16_22(.douta(w_asqrt16_22[0]),.doutb(w_asqrt16_22[1]),.doutc(w_asqrt16_22[2]),.din(w_asqrt16_7[0]));
	jspl3 jspl3_w_asqrt16_23(.douta(w_asqrt16_23[0]),.doutb(w_asqrt16_23[1]),.doutc(w_asqrt16_23[2]),.din(w_asqrt16_7[1]));
	jspl3 jspl3_w_asqrt16_24(.douta(w_asqrt16_24[0]),.doutb(w_asqrt16_24[1]),.doutc(w_asqrt16_24[2]),.din(w_asqrt16_7[2]));
	jspl3 jspl3_w_asqrt16_25(.douta(w_asqrt16_25[0]),.doutb(w_asqrt16_25[1]),.doutc(w_asqrt16_25[2]),.din(w_asqrt16_8[0]));
	jspl3 jspl3_w_asqrt16_26(.douta(w_asqrt16_26[0]),.doutb(w_asqrt16_26[1]),.doutc(w_asqrt16_26[2]),.din(w_asqrt16_8[1]));
	jspl3 jspl3_w_asqrt16_27(.douta(w_asqrt16_27[0]),.doutb(w_asqrt16_27[1]),.doutc(w_asqrt16_27[2]),.din(w_asqrt16_8[2]));
	jspl3 jspl3_w_asqrt16_28(.douta(w_asqrt16_28[0]),.doutb(w_asqrt16_28[1]),.doutc(w_asqrt16_28[2]),.din(w_asqrt16_9[0]));
	jspl3 jspl3_w_asqrt16_29(.douta(w_asqrt16_29[0]),.doutb(w_asqrt16_29[1]),.doutc(w_asqrt16_29[2]),.din(w_asqrt16_9[1]));
	jspl3 jspl3_w_asqrt16_30(.douta(w_asqrt16_30[0]),.doutb(w_asqrt16_30[1]),.doutc(w_asqrt16_30[2]),.din(w_asqrt16_9[2]));
	jspl jspl_w_asqrt16_31(.douta(w_asqrt16_31),.doutb(asqrt[15]),.din(w_asqrt16_10[0]));
	jspl3 jspl3_w_asqrt17_0(.douta(w_asqrt17_0[0]),.doutb(w_asqrt17_0[1]),.doutc(w_asqrt17_0[2]),.din(asqrt_fa_17));
	jspl3 jspl3_w_asqrt17_1(.douta(w_asqrt17_1[0]),.doutb(w_asqrt17_1[1]),.doutc(w_asqrt17_1[2]),.din(w_asqrt17_0[0]));
	jspl3 jspl3_w_asqrt17_2(.douta(w_asqrt17_2[0]),.doutb(w_asqrt17_2[1]),.doutc(w_asqrt17_2[2]),.din(w_asqrt17_0[1]));
	jspl3 jspl3_w_asqrt17_3(.douta(w_asqrt17_3[0]),.doutb(w_asqrt17_3[1]),.doutc(w_asqrt17_3[2]),.din(w_asqrt17_0[2]));
	jspl3 jspl3_w_asqrt17_4(.douta(w_asqrt17_4[0]),.doutb(w_asqrt17_4[1]),.doutc(w_asqrt17_4[2]),.din(w_asqrt17_1[0]));
	jspl3 jspl3_w_asqrt17_5(.douta(w_asqrt17_5[0]),.doutb(w_asqrt17_5[1]),.doutc(w_asqrt17_5[2]),.din(w_asqrt17_1[1]));
	jspl3 jspl3_w_asqrt17_6(.douta(w_asqrt17_6[0]),.doutb(w_asqrt17_6[1]),.doutc(w_asqrt17_6[2]),.din(w_asqrt17_1[2]));
	jspl3 jspl3_w_asqrt17_7(.douta(w_asqrt17_7[0]),.doutb(w_asqrt17_7[1]),.doutc(w_asqrt17_7[2]),.din(w_asqrt17_2[0]));
	jspl3 jspl3_w_asqrt17_8(.douta(w_asqrt17_8[0]),.doutb(w_asqrt17_8[1]),.doutc(w_asqrt17_8[2]),.din(w_asqrt17_2[1]));
	jspl3 jspl3_w_asqrt17_9(.douta(w_asqrt17_9[0]),.doutb(w_asqrt17_9[1]),.doutc(w_asqrt17_9[2]),.din(w_asqrt17_2[2]));
	jspl3 jspl3_w_asqrt17_10(.douta(w_asqrt17_10[0]),.doutb(w_asqrt17_10[1]),.doutc(w_asqrt17_10[2]),.din(w_asqrt17_3[0]));
	jspl3 jspl3_w_asqrt17_11(.douta(w_asqrt17_11[0]),.doutb(w_asqrt17_11[1]),.doutc(w_asqrt17_11[2]),.din(w_asqrt17_3[1]));
	jspl3 jspl3_w_asqrt17_12(.douta(w_asqrt17_12[0]),.doutb(w_asqrt17_12[1]),.doutc(w_asqrt17_12[2]),.din(w_asqrt17_3[2]));
	jspl3 jspl3_w_asqrt17_13(.douta(w_asqrt17_13[0]),.doutb(w_asqrt17_13[1]),.doutc(w_asqrt17_13[2]),.din(w_asqrt17_4[0]));
	jspl3 jspl3_w_asqrt17_14(.douta(w_asqrt17_14[0]),.doutb(w_asqrt17_14[1]),.doutc(w_asqrt17_14[2]),.din(w_asqrt17_4[1]));
	jspl3 jspl3_w_asqrt17_15(.douta(w_asqrt17_15[0]),.doutb(w_asqrt17_15[1]),.doutc(w_asqrt17_15[2]),.din(w_asqrt17_4[2]));
	jspl3 jspl3_w_asqrt17_16(.douta(w_asqrt17_16[0]),.doutb(w_asqrt17_16[1]),.doutc(w_asqrt17_16[2]),.din(w_asqrt17_5[0]));
	jspl3 jspl3_w_asqrt17_17(.douta(w_asqrt17_17[0]),.doutb(w_asqrt17_17[1]),.doutc(w_asqrt17_17[2]),.din(w_asqrt17_5[1]));
	jspl jspl_w_asqrt17_18(.douta(w_asqrt17_18),.doutb(asqrt[16]),.din(w_asqrt17_5[2]));
	jspl3 jspl3_w_asqrt18_0(.douta(w_asqrt18_0[0]),.doutb(w_asqrt18_0[1]),.doutc(w_asqrt18_0[2]),.din(asqrt_fa_18));
	jspl3 jspl3_w_asqrt18_1(.douta(w_asqrt18_1[0]),.doutb(w_asqrt18_1[1]),.doutc(w_asqrt18_1[2]),.din(w_asqrt18_0[0]));
	jspl3 jspl3_w_asqrt18_2(.douta(w_asqrt18_2[0]),.doutb(w_asqrt18_2[1]),.doutc(w_asqrt18_2[2]),.din(w_asqrt18_0[1]));
	jspl3 jspl3_w_asqrt18_3(.douta(w_asqrt18_3[0]),.doutb(w_asqrt18_3[1]),.doutc(w_asqrt18_3[2]),.din(w_asqrt18_0[2]));
	jspl3 jspl3_w_asqrt18_4(.douta(w_asqrt18_4[0]),.doutb(w_asqrt18_4[1]),.doutc(w_asqrt18_4[2]),.din(w_asqrt18_1[0]));
	jspl3 jspl3_w_asqrt18_5(.douta(w_asqrt18_5[0]),.doutb(w_asqrt18_5[1]),.doutc(w_asqrt18_5[2]),.din(w_asqrt18_1[1]));
	jspl3 jspl3_w_asqrt18_6(.douta(w_asqrt18_6[0]),.doutb(w_asqrt18_6[1]),.doutc(w_asqrt18_6[2]),.din(w_asqrt18_1[2]));
	jspl3 jspl3_w_asqrt18_7(.douta(w_asqrt18_7[0]),.doutb(w_asqrt18_7[1]),.doutc(w_asqrt18_7[2]),.din(w_asqrt18_2[0]));
	jspl3 jspl3_w_asqrt18_8(.douta(w_asqrt18_8[0]),.doutb(w_asqrt18_8[1]),.doutc(w_asqrt18_8[2]),.din(w_asqrt18_2[1]));
	jspl3 jspl3_w_asqrt18_9(.douta(w_asqrt18_9[0]),.doutb(w_asqrt18_9[1]),.doutc(w_asqrt18_9[2]),.din(w_asqrt18_2[2]));
	jspl3 jspl3_w_asqrt18_10(.douta(w_asqrt18_10[0]),.doutb(w_asqrt18_10[1]),.doutc(w_asqrt18_10[2]),.din(w_asqrt18_3[0]));
	jspl3 jspl3_w_asqrt18_11(.douta(w_asqrt18_11[0]),.doutb(w_asqrt18_11[1]),.doutc(w_asqrt18_11[2]),.din(w_asqrt18_3[1]));
	jspl3 jspl3_w_asqrt18_12(.douta(w_asqrt18_12[0]),.doutb(w_asqrt18_12[1]),.doutc(w_asqrt18_12[2]),.din(w_asqrt18_3[2]));
	jspl3 jspl3_w_asqrt18_13(.douta(w_asqrt18_13[0]),.doutb(w_asqrt18_13[1]),.doutc(w_asqrt18_13[2]),.din(w_asqrt18_4[0]));
	jspl3 jspl3_w_asqrt18_14(.douta(w_asqrt18_14[0]),.doutb(w_asqrt18_14[1]),.doutc(w_asqrt18_14[2]),.din(w_asqrt18_4[1]));
	jspl3 jspl3_w_asqrt18_15(.douta(w_asqrt18_15[0]),.doutb(w_asqrt18_15[1]),.doutc(w_asqrt18_15[2]),.din(w_asqrt18_4[2]));
	jspl3 jspl3_w_asqrt18_16(.douta(w_asqrt18_16[0]),.doutb(w_asqrt18_16[1]),.doutc(w_asqrt18_16[2]),.din(w_asqrt18_5[0]));
	jspl3 jspl3_w_asqrt18_17(.douta(w_asqrt18_17[0]),.doutb(w_asqrt18_17[1]),.doutc(w_asqrt18_17[2]),.din(w_asqrt18_5[1]));
	jspl3 jspl3_w_asqrt18_18(.douta(w_asqrt18_18[0]),.doutb(w_asqrt18_18[1]),.doutc(w_asqrt18_18[2]),.din(w_asqrt18_5[2]));
	jspl3 jspl3_w_asqrt18_19(.douta(w_asqrt18_19[0]),.doutb(w_asqrt18_19[1]),.doutc(w_asqrt18_19[2]),.din(w_asqrt18_6[0]));
	jspl3 jspl3_w_asqrt18_20(.douta(w_asqrt18_20[0]),.doutb(w_asqrt18_20[1]),.doutc(w_asqrt18_20[2]),.din(w_asqrt18_6[1]));
	jspl3 jspl3_w_asqrt18_21(.douta(w_asqrt18_21[0]),.doutb(w_asqrt18_21[1]),.doutc(w_asqrt18_21[2]),.din(w_asqrt18_6[2]));
	jspl3 jspl3_w_asqrt18_22(.douta(w_asqrt18_22[0]),.doutb(w_asqrt18_22[1]),.doutc(w_asqrt18_22[2]),.din(w_asqrt18_7[0]));
	jspl3 jspl3_w_asqrt18_23(.douta(w_asqrt18_23[0]),.doutb(w_asqrt18_23[1]),.doutc(w_asqrt18_23[2]),.din(w_asqrt18_7[1]));
	jspl3 jspl3_w_asqrt18_24(.douta(w_asqrt18_24[0]),.doutb(w_asqrt18_24[1]),.doutc(w_asqrt18_24[2]),.din(w_asqrt18_7[2]));
	jspl3 jspl3_w_asqrt18_25(.douta(w_asqrt18_25[0]),.doutb(w_asqrt18_25[1]),.doutc(w_asqrt18_25[2]),.din(w_asqrt18_8[0]));
	jspl3 jspl3_w_asqrt18_26(.douta(w_asqrt18_26[0]),.doutb(w_asqrt18_26[1]),.doutc(w_asqrt18_26[2]),.din(w_asqrt18_8[1]));
	jspl3 jspl3_w_asqrt18_27(.douta(w_asqrt18_27[0]),.doutb(w_asqrt18_27[1]),.doutc(w_asqrt18_27[2]),.din(w_asqrt18_8[2]));
	jspl3 jspl3_w_asqrt18_28(.douta(w_asqrt18_28[0]),.doutb(w_asqrt18_28[1]),.doutc(w_asqrt18_28[2]),.din(w_asqrt18_9[0]));
	jspl3 jspl3_w_asqrt18_29(.douta(w_asqrt18_29[0]),.doutb(w_asqrt18_29[1]),.doutc(w_asqrt18_29[2]),.din(w_asqrt18_9[1]));
	jspl3 jspl3_w_asqrt18_30(.douta(w_asqrt18_30[0]),.doutb(w_asqrt18_30[1]),.doutc(w_asqrt18_30[2]),.din(w_asqrt18_9[2]));
	jspl jspl_w_asqrt18_31(.douta(w_asqrt18_31),.doutb(asqrt[17]),.din(w_asqrt18_10[0]));
	jspl3 jspl3_w_asqrt19_0(.douta(w_asqrt19_0[0]),.doutb(w_asqrt19_0[1]),.doutc(w_asqrt19_0[2]),.din(asqrt_fa_19));
	jspl3 jspl3_w_asqrt19_1(.douta(w_asqrt19_1[0]),.doutb(w_asqrt19_1[1]),.doutc(w_asqrt19_1[2]),.din(w_asqrt19_0[0]));
	jspl3 jspl3_w_asqrt19_2(.douta(w_asqrt19_2[0]),.doutb(w_asqrt19_2[1]),.doutc(w_asqrt19_2[2]),.din(w_asqrt19_0[1]));
	jspl3 jspl3_w_asqrt19_3(.douta(w_asqrt19_3[0]),.doutb(w_asqrt19_3[1]),.doutc(w_asqrt19_3[2]),.din(w_asqrt19_0[2]));
	jspl3 jspl3_w_asqrt19_4(.douta(w_asqrt19_4[0]),.doutb(w_asqrt19_4[1]),.doutc(w_asqrt19_4[2]),.din(w_asqrt19_1[0]));
	jspl3 jspl3_w_asqrt19_5(.douta(w_asqrt19_5[0]),.doutb(w_asqrt19_5[1]),.doutc(w_asqrt19_5[2]),.din(w_asqrt19_1[1]));
	jspl3 jspl3_w_asqrt19_6(.douta(w_asqrt19_6[0]),.doutb(w_asqrt19_6[1]),.doutc(w_asqrt19_6[2]),.din(w_asqrt19_1[2]));
	jspl3 jspl3_w_asqrt19_7(.douta(w_asqrt19_7[0]),.doutb(w_asqrt19_7[1]),.doutc(w_asqrt19_7[2]),.din(w_asqrt19_2[0]));
	jspl3 jspl3_w_asqrt19_8(.douta(w_asqrt19_8[0]),.doutb(w_asqrt19_8[1]),.doutc(w_asqrt19_8[2]),.din(w_asqrt19_2[1]));
	jspl3 jspl3_w_asqrt19_9(.douta(w_asqrt19_9[0]),.doutb(w_asqrt19_9[1]),.doutc(w_asqrt19_9[2]),.din(w_asqrt19_2[2]));
	jspl3 jspl3_w_asqrt19_10(.douta(w_asqrt19_10[0]),.doutb(w_asqrt19_10[1]),.doutc(w_asqrt19_10[2]),.din(w_asqrt19_3[0]));
	jspl3 jspl3_w_asqrt19_11(.douta(w_asqrt19_11[0]),.doutb(w_asqrt19_11[1]),.doutc(w_asqrt19_11[2]),.din(w_asqrt19_3[1]));
	jspl3 jspl3_w_asqrt19_12(.douta(w_asqrt19_12[0]),.doutb(w_asqrt19_12[1]),.doutc(w_asqrt19_12[2]),.din(w_asqrt19_3[2]));
	jspl3 jspl3_w_asqrt19_13(.douta(w_asqrt19_13[0]),.doutb(w_asqrt19_13[1]),.doutc(w_asqrt19_13[2]),.din(w_asqrt19_4[0]));
	jspl3 jspl3_w_asqrt19_14(.douta(w_asqrt19_14[0]),.doutb(w_asqrt19_14[1]),.doutc(w_asqrt19_14[2]),.din(w_asqrt19_4[1]));
	jspl3 jspl3_w_asqrt19_15(.douta(w_asqrt19_15[0]),.doutb(w_asqrt19_15[1]),.doutc(w_asqrt19_15[2]),.din(w_asqrt19_4[2]));
	jspl3 jspl3_w_asqrt19_16(.douta(w_asqrt19_16[0]),.doutb(w_asqrt19_16[1]),.doutc(w_asqrt19_16[2]),.din(w_asqrt19_5[0]));
	jspl3 jspl3_w_asqrt19_17(.douta(w_asqrt19_17[0]),.doutb(w_asqrt19_17[1]),.doutc(w_asqrt19_17[2]),.din(w_asqrt19_5[1]));
	jspl jspl_w_asqrt19_18(.douta(w_asqrt19_18),.doutb(asqrt[18]),.din(w_asqrt19_5[2]));
	jspl3 jspl3_w_asqrt20_0(.douta(w_asqrt20_0[0]),.doutb(w_asqrt20_0[1]),.doutc(w_asqrt20_0[2]),.din(asqrt_fa_20));
	jspl3 jspl3_w_asqrt20_1(.douta(w_asqrt20_1[0]),.doutb(w_asqrt20_1[1]),.doutc(w_asqrt20_1[2]),.din(w_asqrt20_0[0]));
	jspl3 jspl3_w_asqrt20_2(.douta(w_asqrt20_2[0]),.doutb(w_asqrt20_2[1]),.doutc(w_asqrt20_2[2]),.din(w_asqrt20_0[1]));
	jspl3 jspl3_w_asqrt20_3(.douta(w_asqrt20_3[0]),.doutb(w_asqrt20_3[1]),.doutc(w_asqrt20_3[2]),.din(w_asqrt20_0[2]));
	jspl3 jspl3_w_asqrt20_4(.douta(w_asqrt20_4[0]),.doutb(w_asqrt20_4[1]),.doutc(w_asqrt20_4[2]),.din(w_asqrt20_1[0]));
	jspl3 jspl3_w_asqrt20_5(.douta(w_asqrt20_5[0]),.doutb(w_asqrt20_5[1]),.doutc(w_asqrt20_5[2]),.din(w_asqrt20_1[1]));
	jspl3 jspl3_w_asqrt20_6(.douta(w_asqrt20_6[0]),.doutb(w_asqrt20_6[1]),.doutc(w_asqrt20_6[2]),.din(w_asqrt20_1[2]));
	jspl3 jspl3_w_asqrt20_7(.douta(w_asqrt20_7[0]),.doutb(w_asqrt20_7[1]),.doutc(w_asqrt20_7[2]),.din(w_asqrt20_2[0]));
	jspl3 jspl3_w_asqrt20_8(.douta(w_asqrt20_8[0]),.doutb(w_asqrt20_8[1]),.doutc(w_asqrt20_8[2]),.din(w_asqrt20_2[1]));
	jspl3 jspl3_w_asqrt20_9(.douta(w_asqrt20_9[0]),.doutb(w_asqrt20_9[1]),.doutc(w_asqrt20_9[2]),.din(w_asqrt20_2[2]));
	jspl3 jspl3_w_asqrt20_10(.douta(w_asqrt20_10[0]),.doutb(w_asqrt20_10[1]),.doutc(w_asqrt20_10[2]),.din(w_asqrt20_3[0]));
	jspl3 jspl3_w_asqrt20_11(.douta(w_asqrt20_11[0]),.doutb(w_asqrt20_11[1]),.doutc(w_asqrt20_11[2]),.din(w_asqrt20_3[1]));
	jspl3 jspl3_w_asqrt20_12(.douta(w_asqrt20_12[0]),.doutb(w_asqrt20_12[1]),.doutc(w_asqrt20_12[2]),.din(w_asqrt20_3[2]));
	jspl3 jspl3_w_asqrt20_13(.douta(w_asqrt20_13[0]),.doutb(w_asqrt20_13[1]),.doutc(w_asqrt20_13[2]),.din(w_asqrt20_4[0]));
	jspl3 jspl3_w_asqrt20_14(.douta(w_asqrt20_14[0]),.doutb(w_asqrt20_14[1]),.doutc(w_asqrt20_14[2]),.din(w_asqrt20_4[1]));
	jspl3 jspl3_w_asqrt20_15(.douta(w_asqrt20_15[0]),.doutb(w_asqrt20_15[1]),.doutc(w_asqrt20_15[2]),.din(w_asqrt20_4[2]));
	jspl3 jspl3_w_asqrt20_16(.douta(w_asqrt20_16[0]),.doutb(w_asqrt20_16[1]),.doutc(w_asqrt20_16[2]),.din(w_asqrt20_5[0]));
	jspl3 jspl3_w_asqrt20_17(.douta(w_asqrt20_17[0]),.doutb(w_asqrt20_17[1]),.doutc(w_asqrt20_17[2]),.din(w_asqrt20_5[1]));
	jspl3 jspl3_w_asqrt20_18(.douta(w_asqrt20_18[0]),.doutb(w_asqrt20_18[1]),.doutc(w_asqrt20_18[2]),.din(w_asqrt20_5[2]));
	jspl3 jspl3_w_asqrt20_19(.douta(w_asqrt20_19[0]),.doutb(w_asqrt20_19[1]),.doutc(w_asqrt20_19[2]),.din(w_asqrt20_6[0]));
	jspl3 jspl3_w_asqrt20_20(.douta(w_asqrt20_20[0]),.doutb(w_asqrt20_20[1]),.doutc(w_asqrt20_20[2]),.din(w_asqrt20_6[1]));
	jspl3 jspl3_w_asqrt20_21(.douta(w_asqrt20_21[0]),.doutb(w_asqrt20_21[1]),.doutc(w_asqrt20_21[2]),.din(w_asqrt20_6[2]));
	jspl3 jspl3_w_asqrt20_22(.douta(w_asqrt20_22[0]),.doutb(w_asqrt20_22[1]),.doutc(w_asqrt20_22[2]),.din(w_asqrt20_7[0]));
	jspl3 jspl3_w_asqrt20_23(.douta(w_asqrt20_23[0]),.doutb(w_asqrt20_23[1]),.doutc(w_asqrt20_23[2]),.din(w_asqrt20_7[1]));
	jspl3 jspl3_w_asqrt20_24(.douta(w_asqrt20_24[0]),.doutb(w_asqrt20_24[1]),.doutc(w_asqrt20_24[2]),.din(w_asqrt20_7[2]));
	jspl3 jspl3_w_asqrt20_25(.douta(w_asqrt20_25[0]),.doutb(w_asqrt20_25[1]),.doutc(w_asqrt20_25[2]),.din(w_asqrt20_8[0]));
	jspl3 jspl3_w_asqrt20_26(.douta(w_asqrt20_26[0]),.doutb(w_asqrt20_26[1]),.doutc(w_asqrt20_26[2]),.din(w_asqrt20_8[1]));
	jspl3 jspl3_w_asqrt20_27(.douta(w_asqrt20_27[0]),.doutb(w_asqrt20_27[1]),.doutc(w_asqrt20_27[2]),.din(w_asqrt20_8[2]));
	jspl3 jspl3_w_asqrt20_28(.douta(w_asqrt20_28[0]),.doutb(w_asqrt20_28[1]),.doutc(w_asqrt20_28[2]),.din(w_asqrt20_9[0]));
	jspl3 jspl3_w_asqrt20_29(.douta(w_asqrt20_29[0]),.doutb(w_asqrt20_29[1]),.doutc(w_asqrt20_29[2]),.din(w_asqrt20_9[1]));
	jspl3 jspl3_w_asqrt20_30(.douta(w_asqrt20_30[0]),.doutb(w_asqrt20_30[1]),.doutc(w_asqrt20_30[2]),.din(w_asqrt20_9[2]));
	jspl jspl_w_asqrt20_31(.douta(w_asqrt20_31),.doutb(asqrt[19]),.din(w_asqrt20_10[0]));
	jspl3 jspl3_w_asqrt21_0(.douta(w_asqrt21_0[0]),.doutb(w_asqrt21_0[1]),.doutc(w_asqrt21_0[2]),.din(asqrt_fa_21));
	jspl3 jspl3_w_asqrt21_1(.douta(w_asqrt21_1[0]),.doutb(w_asqrt21_1[1]),.doutc(w_asqrt21_1[2]),.din(w_asqrt21_0[0]));
	jspl3 jspl3_w_asqrt21_2(.douta(w_asqrt21_2[0]),.doutb(w_asqrt21_2[1]),.doutc(w_asqrt21_2[2]),.din(w_asqrt21_0[1]));
	jspl3 jspl3_w_asqrt21_3(.douta(w_asqrt21_3[0]),.doutb(w_asqrt21_3[1]),.doutc(w_asqrt21_3[2]),.din(w_asqrt21_0[2]));
	jspl3 jspl3_w_asqrt21_4(.douta(w_asqrt21_4[0]),.doutb(w_asqrt21_4[1]),.doutc(w_asqrt21_4[2]),.din(w_asqrt21_1[0]));
	jspl3 jspl3_w_asqrt21_5(.douta(w_asqrt21_5[0]),.doutb(w_asqrt21_5[1]),.doutc(w_asqrt21_5[2]),.din(w_asqrt21_1[1]));
	jspl3 jspl3_w_asqrt21_6(.douta(w_asqrt21_6[0]),.doutb(w_asqrt21_6[1]),.doutc(w_asqrt21_6[2]),.din(w_asqrt21_1[2]));
	jspl3 jspl3_w_asqrt21_7(.douta(w_asqrt21_7[0]),.doutb(w_asqrt21_7[1]),.doutc(w_asqrt21_7[2]),.din(w_asqrt21_2[0]));
	jspl3 jspl3_w_asqrt21_8(.douta(w_asqrt21_8[0]),.doutb(w_asqrt21_8[1]),.doutc(w_asqrt21_8[2]),.din(w_asqrt21_2[1]));
	jspl3 jspl3_w_asqrt21_9(.douta(w_asqrt21_9[0]),.doutb(w_asqrt21_9[1]),.doutc(w_asqrt21_9[2]),.din(w_asqrt21_2[2]));
	jspl3 jspl3_w_asqrt21_10(.douta(w_asqrt21_10[0]),.doutb(w_asqrt21_10[1]),.doutc(w_asqrt21_10[2]),.din(w_asqrt21_3[0]));
	jspl3 jspl3_w_asqrt21_11(.douta(w_asqrt21_11[0]),.doutb(w_asqrt21_11[1]),.doutc(w_asqrt21_11[2]),.din(w_asqrt21_3[1]));
	jspl3 jspl3_w_asqrt21_12(.douta(w_asqrt21_12[0]),.doutb(w_asqrt21_12[1]),.doutc(w_asqrt21_12[2]),.din(w_asqrt21_3[2]));
	jspl3 jspl3_w_asqrt21_13(.douta(w_asqrt21_13[0]),.doutb(w_asqrt21_13[1]),.doutc(w_asqrt21_13[2]),.din(w_asqrt21_4[0]));
	jspl3 jspl3_w_asqrt21_14(.douta(w_asqrt21_14[0]),.doutb(w_asqrt21_14[1]),.doutc(w_asqrt21_14[2]),.din(w_asqrt21_4[1]));
	jspl3 jspl3_w_asqrt21_15(.douta(w_asqrt21_15[0]),.doutb(w_asqrt21_15[1]),.doutc(w_asqrt21_15[2]),.din(w_asqrt21_4[2]));
	jspl3 jspl3_w_asqrt21_16(.douta(w_asqrt21_16[0]),.doutb(w_asqrt21_16[1]),.doutc(w_asqrt21_16[2]),.din(w_asqrt21_5[0]));
	jspl3 jspl3_w_asqrt21_17(.douta(w_asqrt21_17[0]),.doutb(w_asqrt21_17[1]),.doutc(w_asqrt21_17[2]),.din(w_asqrt21_5[1]));
	jspl3 jspl3_w_asqrt21_18(.douta(w_asqrt21_18[0]),.doutb(w_asqrt21_18[1]),.doutc(w_asqrt21_18[2]),.din(w_asqrt21_5[2]));
	jspl jspl_w_asqrt21_19(.douta(w_asqrt21_19),.doutb(asqrt[20]),.din(w_asqrt21_6[0]));
	jspl3 jspl3_w_asqrt22_0(.douta(w_asqrt22_0[0]),.doutb(w_asqrt22_0[1]),.doutc(w_asqrt22_0[2]),.din(asqrt_fa_22));
	jspl3 jspl3_w_asqrt22_1(.douta(w_asqrt22_1[0]),.doutb(w_asqrt22_1[1]),.doutc(w_asqrt22_1[2]),.din(w_asqrt22_0[0]));
	jspl3 jspl3_w_asqrt22_2(.douta(w_asqrt22_2[0]),.doutb(w_asqrt22_2[1]),.doutc(w_asqrt22_2[2]),.din(w_asqrt22_0[1]));
	jspl3 jspl3_w_asqrt22_3(.douta(w_asqrt22_3[0]),.doutb(w_asqrt22_3[1]),.doutc(w_asqrt22_3[2]),.din(w_asqrt22_0[2]));
	jspl3 jspl3_w_asqrt22_4(.douta(w_asqrt22_4[0]),.doutb(w_asqrt22_4[1]),.doutc(w_asqrt22_4[2]),.din(w_asqrt22_1[0]));
	jspl3 jspl3_w_asqrt22_5(.douta(w_asqrt22_5[0]),.doutb(w_asqrt22_5[1]),.doutc(w_asqrt22_5[2]),.din(w_asqrt22_1[1]));
	jspl3 jspl3_w_asqrt22_6(.douta(w_asqrt22_6[0]),.doutb(w_asqrt22_6[1]),.doutc(w_asqrt22_6[2]),.din(w_asqrt22_1[2]));
	jspl3 jspl3_w_asqrt22_7(.douta(w_asqrt22_7[0]),.doutb(w_asqrt22_7[1]),.doutc(w_asqrt22_7[2]),.din(w_asqrt22_2[0]));
	jspl3 jspl3_w_asqrt22_8(.douta(w_asqrt22_8[0]),.doutb(w_asqrt22_8[1]),.doutc(w_asqrt22_8[2]),.din(w_asqrt22_2[1]));
	jspl3 jspl3_w_asqrt22_9(.douta(w_asqrt22_9[0]),.doutb(w_asqrt22_9[1]),.doutc(w_asqrt22_9[2]),.din(w_asqrt22_2[2]));
	jspl3 jspl3_w_asqrt22_10(.douta(w_asqrt22_10[0]),.doutb(w_asqrt22_10[1]),.doutc(w_asqrt22_10[2]),.din(w_asqrt22_3[0]));
	jspl3 jspl3_w_asqrt22_11(.douta(w_asqrt22_11[0]),.doutb(w_asqrt22_11[1]),.doutc(w_asqrt22_11[2]),.din(w_asqrt22_3[1]));
	jspl3 jspl3_w_asqrt22_12(.douta(w_asqrt22_12[0]),.doutb(w_asqrt22_12[1]),.doutc(w_asqrt22_12[2]),.din(w_asqrt22_3[2]));
	jspl3 jspl3_w_asqrt22_13(.douta(w_asqrt22_13[0]),.doutb(w_asqrt22_13[1]),.doutc(w_asqrt22_13[2]),.din(w_asqrt22_4[0]));
	jspl3 jspl3_w_asqrt22_14(.douta(w_asqrt22_14[0]),.doutb(w_asqrt22_14[1]),.doutc(w_asqrt22_14[2]),.din(w_asqrt22_4[1]));
	jspl3 jspl3_w_asqrt22_15(.douta(w_asqrt22_15[0]),.doutb(w_asqrt22_15[1]),.doutc(w_asqrt22_15[2]),.din(w_asqrt22_4[2]));
	jspl3 jspl3_w_asqrt22_16(.douta(w_asqrt22_16[0]),.doutb(w_asqrt22_16[1]),.doutc(w_asqrt22_16[2]),.din(w_asqrt22_5[0]));
	jspl3 jspl3_w_asqrt22_17(.douta(w_asqrt22_17[0]),.doutb(w_asqrt22_17[1]),.doutc(w_asqrt22_17[2]),.din(w_asqrt22_5[1]));
	jspl3 jspl3_w_asqrt22_18(.douta(w_asqrt22_18[0]),.doutb(w_asqrt22_18[1]),.doutc(w_asqrt22_18[2]),.din(w_asqrt22_5[2]));
	jspl3 jspl3_w_asqrt22_19(.douta(w_asqrt22_19[0]),.doutb(w_asqrt22_19[1]),.doutc(w_asqrt22_19[2]),.din(w_asqrt22_6[0]));
	jspl3 jspl3_w_asqrt22_20(.douta(w_asqrt22_20[0]),.doutb(w_asqrt22_20[1]),.doutc(w_asqrt22_20[2]),.din(w_asqrt22_6[1]));
	jspl3 jspl3_w_asqrt22_21(.douta(w_asqrt22_21[0]),.doutb(w_asqrt22_21[1]),.doutc(w_asqrt22_21[2]),.din(w_asqrt22_6[2]));
	jspl3 jspl3_w_asqrt22_22(.douta(w_asqrt22_22[0]),.doutb(w_asqrt22_22[1]),.doutc(w_asqrt22_22[2]),.din(w_asqrt22_7[0]));
	jspl3 jspl3_w_asqrt22_23(.douta(w_asqrt22_23[0]),.doutb(w_asqrt22_23[1]),.doutc(w_asqrt22_23[2]),.din(w_asqrt22_7[1]));
	jspl3 jspl3_w_asqrt22_24(.douta(w_asqrt22_24[0]),.doutb(w_asqrt22_24[1]),.doutc(w_asqrt22_24[2]),.din(w_asqrt22_7[2]));
	jspl3 jspl3_w_asqrt22_25(.douta(w_asqrt22_25[0]),.doutb(w_asqrt22_25[1]),.doutc(w_asqrt22_25[2]),.din(w_asqrt22_8[0]));
	jspl3 jspl3_w_asqrt22_26(.douta(w_asqrt22_26[0]),.doutb(w_asqrt22_26[1]),.doutc(w_asqrt22_26[2]),.din(w_asqrt22_8[1]));
	jspl3 jspl3_w_asqrt22_27(.douta(w_asqrt22_27[0]),.doutb(w_asqrt22_27[1]),.doutc(w_asqrt22_27[2]),.din(w_asqrt22_8[2]));
	jspl3 jspl3_w_asqrt22_28(.douta(w_asqrt22_28[0]),.doutb(w_asqrt22_28[1]),.doutc(w_asqrt22_28[2]),.din(w_asqrt22_9[0]));
	jspl3 jspl3_w_asqrt22_29(.douta(w_asqrt22_29[0]),.doutb(w_asqrt22_29[1]),.doutc(w_asqrt22_29[2]),.din(w_asqrt22_9[1]));
	jspl3 jspl3_w_asqrt22_30(.douta(w_asqrt22_30[0]),.doutb(w_asqrt22_30[1]),.doutc(w_asqrt22_30[2]),.din(w_asqrt22_9[2]));
	jspl jspl_w_asqrt22_31(.douta(w_asqrt22_31),.doutb(asqrt[21]),.din(w_asqrt22_10[0]));
	jspl3 jspl3_w_asqrt23_0(.douta(w_asqrt23_0[0]),.doutb(w_asqrt23_0[1]),.doutc(w_asqrt23_0[2]),.din(asqrt_fa_23));
	jspl3 jspl3_w_asqrt23_1(.douta(w_asqrt23_1[0]),.doutb(w_asqrt23_1[1]),.doutc(w_asqrt23_1[2]),.din(w_asqrt23_0[0]));
	jspl3 jspl3_w_asqrt23_2(.douta(w_asqrt23_2[0]),.doutb(w_asqrt23_2[1]),.doutc(w_asqrt23_2[2]),.din(w_asqrt23_0[1]));
	jspl3 jspl3_w_asqrt23_3(.douta(w_asqrt23_3[0]),.doutb(w_asqrt23_3[1]),.doutc(w_asqrt23_3[2]),.din(w_asqrt23_0[2]));
	jspl3 jspl3_w_asqrt23_4(.douta(w_asqrt23_4[0]),.doutb(w_asqrt23_4[1]),.doutc(w_asqrt23_4[2]),.din(w_asqrt23_1[0]));
	jspl3 jspl3_w_asqrt23_5(.douta(w_asqrt23_5[0]),.doutb(w_asqrt23_5[1]),.doutc(w_asqrt23_5[2]),.din(w_asqrt23_1[1]));
	jspl3 jspl3_w_asqrt23_6(.douta(w_asqrt23_6[0]),.doutb(w_asqrt23_6[1]),.doutc(w_asqrt23_6[2]),.din(w_asqrt23_1[2]));
	jspl3 jspl3_w_asqrt23_7(.douta(w_asqrt23_7[0]),.doutb(w_asqrt23_7[1]),.doutc(w_asqrt23_7[2]),.din(w_asqrt23_2[0]));
	jspl3 jspl3_w_asqrt23_8(.douta(w_asqrt23_8[0]),.doutb(w_asqrt23_8[1]),.doutc(w_asqrt23_8[2]),.din(w_asqrt23_2[1]));
	jspl3 jspl3_w_asqrt23_9(.douta(w_asqrt23_9[0]),.doutb(w_asqrt23_9[1]),.doutc(w_asqrt23_9[2]),.din(w_asqrt23_2[2]));
	jspl3 jspl3_w_asqrt23_10(.douta(w_asqrt23_10[0]),.doutb(w_asqrt23_10[1]),.doutc(w_asqrt23_10[2]),.din(w_asqrt23_3[0]));
	jspl3 jspl3_w_asqrt23_11(.douta(w_asqrt23_11[0]),.doutb(w_asqrt23_11[1]),.doutc(w_asqrt23_11[2]),.din(w_asqrt23_3[1]));
	jspl3 jspl3_w_asqrt23_12(.douta(w_asqrt23_12[0]),.doutb(w_asqrt23_12[1]),.doutc(w_asqrt23_12[2]),.din(w_asqrt23_3[2]));
	jspl3 jspl3_w_asqrt23_13(.douta(w_asqrt23_13[0]),.doutb(w_asqrt23_13[1]),.doutc(w_asqrt23_13[2]),.din(w_asqrt23_4[0]));
	jspl3 jspl3_w_asqrt23_14(.douta(w_asqrt23_14[0]),.doutb(w_asqrt23_14[1]),.doutc(w_asqrt23_14[2]),.din(w_asqrt23_4[1]));
	jspl3 jspl3_w_asqrt23_15(.douta(w_asqrt23_15[0]),.doutb(w_asqrt23_15[1]),.doutc(w_asqrt23_15[2]),.din(w_asqrt23_4[2]));
	jspl3 jspl3_w_asqrt23_16(.douta(w_asqrt23_16[0]),.doutb(w_asqrt23_16[1]),.doutc(w_asqrt23_16[2]),.din(w_asqrt23_5[0]));
	jspl3 jspl3_w_asqrt23_17(.douta(w_asqrt23_17[0]),.doutb(w_asqrt23_17[1]),.doutc(w_asqrt23_17[2]),.din(w_asqrt23_5[1]));
	jspl3 jspl3_w_asqrt23_18(.douta(w_asqrt23_18[0]),.doutb(w_asqrt23_18[1]),.doutc(w_asqrt23_18[2]),.din(w_asqrt23_5[2]));
	jspl jspl_w_asqrt23_19(.douta(w_asqrt23_19),.doutb(asqrt[22]),.din(w_asqrt23_6[0]));
	jspl3 jspl3_w_asqrt24_0(.douta(w_asqrt24_0[0]),.doutb(w_asqrt24_0[1]),.doutc(w_asqrt24_0[2]),.din(asqrt_fa_24));
	jspl3 jspl3_w_asqrt24_1(.douta(w_asqrt24_1[0]),.doutb(w_asqrt24_1[1]),.doutc(w_asqrt24_1[2]),.din(w_asqrt24_0[0]));
	jspl3 jspl3_w_asqrt24_2(.douta(w_asqrt24_2[0]),.doutb(w_asqrt24_2[1]),.doutc(w_asqrt24_2[2]),.din(w_asqrt24_0[1]));
	jspl3 jspl3_w_asqrt24_3(.douta(w_asqrt24_3[0]),.doutb(w_asqrt24_3[1]),.doutc(w_asqrt24_3[2]),.din(w_asqrt24_0[2]));
	jspl3 jspl3_w_asqrt24_4(.douta(w_asqrt24_4[0]),.doutb(w_asqrt24_4[1]),.doutc(w_asqrt24_4[2]),.din(w_asqrt24_1[0]));
	jspl3 jspl3_w_asqrt24_5(.douta(w_asqrt24_5[0]),.doutb(w_asqrt24_5[1]),.doutc(w_asqrt24_5[2]),.din(w_asqrt24_1[1]));
	jspl3 jspl3_w_asqrt24_6(.douta(w_asqrt24_6[0]),.doutb(w_asqrt24_6[1]),.doutc(w_asqrt24_6[2]),.din(w_asqrt24_1[2]));
	jspl3 jspl3_w_asqrt24_7(.douta(w_asqrt24_7[0]),.doutb(w_asqrt24_7[1]),.doutc(w_asqrt24_7[2]),.din(w_asqrt24_2[0]));
	jspl3 jspl3_w_asqrt24_8(.douta(w_asqrt24_8[0]),.doutb(w_asqrt24_8[1]),.doutc(w_asqrt24_8[2]),.din(w_asqrt24_2[1]));
	jspl3 jspl3_w_asqrt24_9(.douta(w_asqrt24_9[0]),.doutb(w_asqrt24_9[1]),.doutc(w_asqrt24_9[2]),.din(w_asqrt24_2[2]));
	jspl3 jspl3_w_asqrt24_10(.douta(w_asqrt24_10[0]),.doutb(w_asqrt24_10[1]),.doutc(w_asqrt24_10[2]),.din(w_asqrt24_3[0]));
	jspl3 jspl3_w_asqrt24_11(.douta(w_asqrt24_11[0]),.doutb(w_asqrt24_11[1]),.doutc(w_asqrt24_11[2]),.din(w_asqrt24_3[1]));
	jspl3 jspl3_w_asqrt24_12(.douta(w_asqrt24_12[0]),.doutb(w_asqrt24_12[1]),.doutc(w_asqrt24_12[2]),.din(w_asqrt24_3[2]));
	jspl3 jspl3_w_asqrt24_13(.douta(w_asqrt24_13[0]),.doutb(w_asqrt24_13[1]),.doutc(w_asqrt24_13[2]),.din(w_asqrt24_4[0]));
	jspl3 jspl3_w_asqrt24_14(.douta(w_asqrt24_14[0]),.doutb(w_asqrt24_14[1]),.doutc(w_asqrt24_14[2]),.din(w_asqrt24_4[1]));
	jspl3 jspl3_w_asqrt24_15(.douta(w_asqrt24_15[0]),.doutb(w_asqrt24_15[1]),.doutc(w_asqrt24_15[2]),.din(w_asqrt24_4[2]));
	jspl3 jspl3_w_asqrt24_16(.douta(w_asqrt24_16[0]),.doutb(w_asqrt24_16[1]),.doutc(w_asqrt24_16[2]),.din(w_asqrt24_5[0]));
	jspl3 jspl3_w_asqrt24_17(.douta(w_asqrt24_17[0]),.doutb(w_asqrt24_17[1]),.doutc(w_asqrt24_17[2]),.din(w_asqrt24_5[1]));
	jspl3 jspl3_w_asqrt24_18(.douta(w_asqrt24_18[0]),.doutb(w_asqrt24_18[1]),.doutc(w_asqrt24_18[2]),.din(w_asqrt24_5[2]));
	jspl3 jspl3_w_asqrt24_19(.douta(w_asqrt24_19[0]),.doutb(w_asqrt24_19[1]),.doutc(w_asqrt24_19[2]),.din(w_asqrt24_6[0]));
	jspl3 jspl3_w_asqrt24_20(.douta(w_asqrt24_20[0]),.doutb(w_asqrt24_20[1]),.doutc(w_asqrt24_20[2]),.din(w_asqrt24_6[1]));
	jspl3 jspl3_w_asqrt24_21(.douta(w_asqrt24_21[0]),.doutb(w_asqrt24_21[1]),.doutc(w_asqrt24_21[2]),.din(w_asqrt24_6[2]));
	jspl3 jspl3_w_asqrt24_22(.douta(w_asqrt24_22[0]),.doutb(w_asqrt24_22[1]),.doutc(w_asqrt24_22[2]),.din(w_asqrt24_7[0]));
	jspl3 jspl3_w_asqrt24_23(.douta(w_asqrt24_23[0]),.doutb(w_asqrt24_23[1]),.doutc(w_asqrt24_23[2]),.din(w_asqrt24_7[1]));
	jspl3 jspl3_w_asqrt24_24(.douta(w_asqrt24_24[0]),.doutb(w_asqrt24_24[1]),.doutc(w_asqrt24_24[2]),.din(w_asqrt24_7[2]));
	jspl3 jspl3_w_asqrt24_25(.douta(w_asqrt24_25[0]),.doutb(w_asqrt24_25[1]),.doutc(w_asqrt24_25[2]),.din(w_asqrt24_8[0]));
	jspl3 jspl3_w_asqrt24_26(.douta(w_asqrt24_26[0]),.doutb(w_asqrt24_26[1]),.doutc(w_asqrt24_26[2]),.din(w_asqrt24_8[1]));
	jspl3 jspl3_w_asqrt24_27(.douta(w_asqrt24_27[0]),.doutb(w_asqrt24_27[1]),.doutc(w_asqrt24_27[2]),.din(w_asqrt24_8[2]));
	jspl3 jspl3_w_asqrt24_28(.douta(w_asqrt24_28[0]),.doutb(w_asqrt24_28[1]),.doutc(w_asqrt24_28[2]),.din(w_asqrt24_9[0]));
	jspl3 jspl3_w_asqrt24_29(.douta(w_asqrt24_29[0]),.doutb(w_asqrt24_29[1]),.doutc(w_asqrt24_29[2]),.din(w_asqrt24_9[1]));
	jspl3 jspl3_w_asqrt24_30(.douta(w_asqrt24_30[0]),.doutb(w_asqrt24_30[1]),.doutc(w_asqrt24_30[2]),.din(w_asqrt24_9[2]));
	jspl jspl_w_asqrt24_31(.douta(w_asqrt24_31),.doutb(asqrt[23]),.din(w_asqrt24_10[0]));
	jspl3 jspl3_w_asqrt25_0(.douta(w_asqrt25_0[0]),.doutb(w_asqrt25_0[1]),.doutc(w_asqrt25_0[2]),.din(asqrt_fa_25));
	jspl3 jspl3_w_asqrt25_1(.douta(w_asqrt25_1[0]),.doutb(w_asqrt25_1[1]),.doutc(w_asqrt25_1[2]),.din(w_asqrt25_0[0]));
	jspl3 jspl3_w_asqrt25_2(.douta(w_asqrt25_2[0]),.doutb(w_asqrt25_2[1]),.doutc(w_asqrt25_2[2]),.din(w_asqrt25_0[1]));
	jspl3 jspl3_w_asqrt25_3(.douta(w_asqrt25_3[0]),.doutb(w_asqrt25_3[1]),.doutc(w_asqrt25_3[2]),.din(w_asqrt25_0[2]));
	jspl3 jspl3_w_asqrt25_4(.douta(w_asqrt25_4[0]),.doutb(w_asqrt25_4[1]),.doutc(w_asqrt25_4[2]),.din(w_asqrt25_1[0]));
	jspl3 jspl3_w_asqrt25_5(.douta(w_asqrt25_5[0]),.doutb(w_asqrt25_5[1]),.doutc(w_asqrt25_5[2]),.din(w_asqrt25_1[1]));
	jspl3 jspl3_w_asqrt25_6(.douta(w_asqrt25_6[0]),.doutb(w_asqrt25_6[1]),.doutc(w_asqrt25_6[2]),.din(w_asqrt25_1[2]));
	jspl3 jspl3_w_asqrt25_7(.douta(w_asqrt25_7[0]),.doutb(w_asqrt25_7[1]),.doutc(w_asqrt25_7[2]),.din(w_asqrt25_2[0]));
	jspl3 jspl3_w_asqrt25_8(.douta(w_asqrt25_8[0]),.doutb(w_asqrt25_8[1]),.doutc(w_asqrt25_8[2]),.din(w_asqrt25_2[1]));
	jspl3 jspl3_w_asqrt25_9(.douta(w_asqrt25_9[0]),.doutb(w_asqrt25_9[1]),.doutc(w_asqrt25_9[2]),.din(w_asqrt25_2[2]));
	jspl3 jspl3_w_asqrt25_10(.douta(w_asqrt25_10[0]),.doutb(w_asqrt25_10[1]),.doutc(w_asqrt25_10[2]),.din(w_asqrt25_3[0]));
	jspl3 jspl3_w_asqrt25_11(.douta(w_asqrt25_11[0]),.doutb(w_asqrt25_11[1]),.doutc(w_asqrt25_11[2]),.din(w_asqrt25_3[1]));
	jspl3 jspl3_w_asqrt25_12(.douta(w_asqrt25_12[0]),.doutb(w_asqrt25_12[1]),.doutc(w_asqrt25_12[2]),.din(w_asqrt25_3[2]));
	jspl3 jspl3_w_asqrt25_13(.douta(w_asqrt25_13[0]),.doutb(w_asqrt25_13[1]),.doutc(w_asqrt25_13[2]),.din(w_asqrt25_4[0]));
	jspl3 jspl3_w_asqrt25_14(.douta(w_asqrt25_14[0]),.doutb(w_asqrt25_14[1]),.doutc(w_asqrt25_14[2]),.din(w_asqrt25_4[1]));
	jspl3 jspl3_w_asqrt25_15(.douta(w_asqrt25_15[0]),.doutb(w_asqrt25_15[1]),.doutc(w_asqrt25_15[2]),.din(w_asqrt25_4[2]));
	jspl3 jspl3_w_asqrt25_16(.douta(w_asqrt25_16[0]),.doutb(w_asqrt25_16[1]),.doutc(w_asqrt25_16[2]),.din(w_asqrt25_5[0]));
	jspl3 jspl3_w_asqrt25_17(.douta(w_asqrt25_17[0]),.doutb(w_asqrt25_17[1]),.doutc(w_asqrt25_17[2]),.din(w_asqrt25_5[1]));
	jspl3 jspl3_w_asqrt25_18(.douta(w_asqrt25_18[0]),.doutb(w_asqrt25_18[1]),.doutc(w_asqrt25_18[2]),.din(w_asqrt25_5[2]));
	jspl3 jspl3_w_asqrt25_19(.douta(w_asqrt25_19[0]),.doutb(w_asqrt25_19[1]),.doutc(w_asqrt25_19[2]),.din(w_asqrt25_6[0]));
	jspl jspl_w_asqrt25_20(.douta(w_asqrt25_20),.doutb(asqrt[24]),.din(w_asqrt25_6[1]));
	jspl3 jspl3_w_asqrt26_0(.douta(w_asqrt26_0[0]),.doutb(w_asqrt26_0[1]),.doutc(w_asqrt26_0[2]),.din(asqrt_fa_26));
	jspl3 jspl3_w_asqrt26_1(.douta(w_asqrt26_1[0]),.doutb(w_asqrt26_1[1]),.doutc(w_asqrt26_1[2]),.din(w_asqrt26_0[0]));
	jspl3 jspl3_w_asqrt26_2(.douta(w_asqrt26_2[0]),.doutb(w_asqrt26_2[1]),.doutc(w_asqrt26_2[2]),.din(w_asqrt26_0[1]));
	jspl3 jspl3_w_asqrt26_3(.douta(w_asqrt26_3[0]),.doutb(w_asqrt26_3[1]),.doutc(w_asqrt26_3[2]),.din(w_asqrt26_0[2]));
	jspl3 jspl3_w_asqrt26_4(.douta(w_asqrt26_4[0]),.doutb(w_asqrt26_4[1]),.doutc(w_asqrt26_4[2]),.din(w_asqrt26_1[0]));
	jspl3 jspl3_w_asqrt26_5(.douta(w_asqrt26_5[0]),.doutb(w_asqrt26_5[1]),.doutc(w_asqrt26_5[2]),.din(w_asqrt26_1[1]));
	jspl3 jspl3_w_asqrt26_6(.douta(w_asqrt26_6[0]),.doutb(w_asqrt26_6[1]),.doutc(w_asqrt26_6[2]),.din(w_asqrt26_1[2]));
	jspl3 jspl3_w_asqrt26_7(.douta(w_asqrt26_7[0]),.doutb(w_asqrt26_7[1]),.doutc(w_asqrt26_7[2]),.din(w_asqrt26_2[0]));
	jspl3 jspl3_w_asqrt26_8(.douta(w_asqrt26_8[0]),.doutb(w_asqrt26_8[1]),.doutc(w_asqrt26_8[2]),.din(w_asqrt26_2[1]));
	jspl3 jspl3_w_asqrt26_9(.douta(w_asqrt26_9[0]),.doutb(w_asqrt26_9[1]),.doutc(w_asqrt26_9[2]),.din(w_asqrt26_2[2]));
	jspl3 jspl3_w_asqrt26_10(.douta(w_asqrt26_10[0]),.doutb(w_asqrt26_10[1]),.doutc(w_asqrt26_10[2]),.din(w_asqrt26_3[0]));
	jspl3 jspl3_w_asqrt26_11(.douta(w_asqrt26_11[0]),.doutb(w_asqrt26_11[1]),.doutc(w_asqrt26_11[2]),.din(w_asqrt26_3[1]));
	jspl3 jspl3_w_asqrt26_12(.douta(w_asqrt26_12[0]),.doutb(w_asqrt26_12[1]),.doutc(w_asqrt26_12[2]),.din(w_asqrt26_3[2]));
	jspl3 jspl3_w_asqrt26_13(.douta(w_asqrt26_13[0]),.doutb(w_asqrt26_13[1]),.doutc(w_asqrt26_13[2]),.din(w_asqrt26_4[0]));
	jspl3 jspl3_w_asqrt26_14(.douta(w_asqrt26_14[0]),.doutb(w_asqrt26_14[1]),.doutc(w_asqrt26_14[2]),.din(w_asqrt26_4[1]));
	jspl3 jspl3_w_asqrt26_15(.douta(w_asqrt26_15[0]),.doutb(w_asqrt26_15[1]),.doutc(w_asqrt26_15[2]),.din(w_asqrt26_4[2]));
	jspl3 jspl3_w_asqrt26_16(.douta(w_asqrt26_16[0]),.doutb(w_asqrt26_16[1]),.doutc(w_asqrt26_16[2]),.din(w_asqrt26_5[0]));
	jspl3 jspl3_w_asqrt26_17(.douta(w_asqrt26_17[0]),.doutb(w_asqrt26_17[1]),.doutc(w_asqrt26_17[2]),.din(w_asqrt26_5[1]));
	jspl3 jspl3_w_asqrt26_18(.douta(w_asqrt26_18[0]),.doutb(w_asqrt26_18[1]),.doutc(w_asqrt26_18[2]),.din(w_asqrt26_5[2]));
	jspl3 jspl3_w_asqrt26_19(.douta(w_asqrt26_19[0]),.doutb(w_asqrt26_19[1]),.doutc(w_asqrt26_19[2]),.din(w_asqrt26_6[0]));
	jspl3 jspl3_w_asqrt26_20(.douta(w_asqrt26_20[0]),.doutb(w_asqrt26_20[1]),.doutc(w_asqrt26_20[2]),.din(w_asqrt26_6[1]));
	jspl3 jspl3_w_asqrt26_21(.douta(w_asqrt26_21[0]),.doutb(w_asqrt26_21[1]),.doutc(w_asqrt26_21[2]),.din(w_asqrt26_6[2]));
	jspl3 jspl3_w_asqrt26_22(.douta(w_asqrt26_22[0]),.doutb(w_asqrt26_22[1]),.doutc(w_asqrt26_22[2]),.din(w_asqrt26_7[0]));
	jspl3 jspl3_w_asqrt26_23(.douta(w_asqrt26_23[0]),.doutb(w_asqrt26_23[1]),.doutc(w_asqrt26_23[2]),.din(w_asqrt26_7[1]));
	jspl3 jspl3_w_asqrt26_24(.douta(w_asqrt26_24[0]),.doutb(w_asqrt26_24[1]),.doutc(w_asqrt26_24[2]),.din(w_asqrt26_7[2]));
	jspl3 jspl3_w_asqrt26_25(.douta(w_asqrt26_25[0]),.doutb(w_asqrt26_25[1]),.doutc(w_asqrt26_25[2]),.din(w_asqrt26_8[0]));
	jspl3 jspl3_w_asqrt26_26(.douta(w_asqrt26_26[0]),.doutb(w_asqrt26_26[1]),.doutc(w_asqrt26_26[2]),.din(w_asqrt26_8[1]));
	jspl3 jspl3_w_asqrt26_27(.douta(w_asqrt26_27[0]),.doutb(w_asqrt26_27[1]),.doutc(w_asqrt26_27[2]),.din(w_asqrt26_8[2]));
	jspl3 jspl3_w_asqrt26_28(.douta(w_asqrt26_28[0]),.doutb(w_asqrt26_28[1]),.doutc(w_asqrt26_28[2]),.din(w_asqrt26_9[0]));
	jspl3 jspl3_w_asqrt26_29(.douta(w_asqrt26_29[0]),.doutb(w_asqrt26_29[1]),.doutc(w_asqrt26_29[2]),.din(w_asqrt26_9[1]));
	jspl3 jspl3_w_asqrt26_30(.douta(w_asqrt26_30[0]),.doutb(w_asqrt26_30[1]),.doutc(w_asqrt26_30[2]),.din(w_asqrt26_9[2]));
	jspl jspl_w_asqrt26_31(.douta(w_asqrt26_31),.doutb(asqrt[25]),.din(w_asqrt26_10[0]));
	jspl3 jspl3_w_asqrt27_0(.douta(w_asqrt27_0[0]),.doutb(w_asqrt27_0[1]),.doutc(w_asqrt27_0[2]),.din(asqrt_fa_27));
	jspl3 jspl3_w_asqrt27_1(.douta(w_asqrt27_1[0]),.doutb(w_asqrt27_1[1]),.doutc(w_asqrt27_1[2]),.din(w_asqrt27_0[0]));
	jspl3 jspl3_w_asqrt27_2(.douta(w_asqrt27_2[0]),.doutb(w_asqrt27_2[1]),.doutc(w_asqrt27_2[2]),.din(w_asqrt27_0[1]));
	jspl3 jspl3_w_asqrt27_3(.douta(w_asqrt27_3[0]),.doutb(w_asqrt27_3[1]),.doutc(w_asqrt27_3[2]),.din(w_asqrt27_0[2]));
	jspl3 jspl3_w_asqrt27_4(.douta(w_asqrt27_4[0]),.doutb(w_asqrt27_4[1]),.doutc(w_asqrt27_4[2]),.din(w_asqrt27_1[0]));
	jspl3 jspl3_w_asqrt27_5(.douta(w_asqrt27_5[0]),.doutb(w_asqrt27_5[1]),.doutc(w_asqrt27_5[2]),.din(w_asqrt27_1[1]));
	jspl3 jspl3_w_asqrt27_6(.douta(w_asqrt27_6[0]),.doutb(w_asqrt27_6[1]),.doutc(w_asqrt27_6[2]),.din(w_asqrt27_1[2]));
	jspl3 jspl3_w_asqrt27_7(.douta(w_asqrt27_7[0]),.doutb(w_asqrt27_7[1]),.doutc(w_asqrt27_7[2]),.din(w_asqrt27_2[0]));
	jspl3 jspl3_w_asqrt27_8(.douta(w_asqrt27_8[0]),.doutb(w_asqrt27_8[1]),.doutc(w_asqrt27_8[2]),.din(w_asqrt27_2[1]));
	jspl3 jspl3_w_asqrt27_9(.douta(w_asqrt27_9[0]),.doutb(w_asqrt27_9[1]),.doutc(w_asqrt27_9[2]),.din(w_asqrt27_2[2]));
	jspl3 jspl3_w_asqrt27_10(.douta(w_asqrt27_10[0]),.doutb(w_asqrt27_10[1]),.doutc(w_asqrt27_10[2]),.din(w_asqrt27_3[0]));
	jspl3 jspl3_w_asqrt27_11(.douta(w_asqrt27_11[0]),.doutb(w_asqrt27_11[1]),.doutc(w_asqrt27_11[2]),.din(w_asqrt27_3[1]));
	jspl3 jspl3_w_asqrt27_12(.douta(w_asqrt27_12[0]),.doutb(w_asqrt27_12[1]),.doutc(w_asqrt27_12[2]),.din(w_asqrt27_3[2]));
	jspl3 jspl3_w_asqrt27_13(.douta(w_asqrt27_13[0]),.doutb(w_asqrt27_13[1]),.doutc(w_asqrt27_13[2]),.din(w_asqrt27_4[0]));
	jspl3 jspl3_w_asqrt27_14(.douta(w_asqrt27_14[0]),.doutb(w_asqrt27_14[1]),.doutc(w_asqrt27_14[2]),.din(w_asqrt27_4[1]));
	jspl3 jspl3_w_asqrt27_15(.douta(w_asqrt27_15[0]),.doutb(w_asqrt27_15[1]),.doutc(w_asqrt27_15[2]),.din(w_asqrt27_4[2]));
	jspl3 jspl3_w_asqrt27_16(.douta(w_asqrt27_16[0]),.doutb(w_asqrt27_16[1]),.doutc(w_asqrt27_16[2]),.din(w_asqrt27_5[0]));
	jspl3 jspl3_w_asqrt27_17(.douta(w_asqrt27_17[0]),.doutb(w_asqrt27_17[1]),.doutc(w_asqrt27_17[2]),.din(w_asqrt27_5[1]));
	jspl3 jspl3_w_asqrt27_18(.douta(w_asqrt27_18[0]),.doutb(w_asqrt27_18[1]),.doutc(w_asqrt27_18[2]),.din(w_asqrt27_5[2]));
	jspl3 jspl3_w_asqrt27_19(.douta(w_asqrt27_19[0]),.doutb(w_asqrt27_19[1]),.doutc(w_asqrt27_19[2]),.din(w_asqrt27_6[0]));
	jspl3 jspl3_w_asqrt27_20(.douta(w_asqrt27_20[0]),.doutb(w_asqrt27_20[1]),.doutc(asqrt[26]),.din(w_asqrt27_6[1]));
	jspl3 jspl3_w_asqrt28_0(.douta(w_asqrt28_0[0]),.doutb(w_asqrt28_0[1]),.doutc(w_asqrt28_0[2]),.din(asqrt_fa_28));
	jspl3 jspl3_w_asqrt28_1(.douta(w_asqrt28_1[0]),.doutb(w_asqrt28_1[1]),.doutc(w_asqrt28_1[2]),.din(w_asqrt28_0[0]));
	jspl3 jspl3_w_asqrt28_2(.douta(w_asqrt28_2[0]),.doutb(w_asqrt28_2[1]),.doutc(w_asqrt28_2[2]),.din(w_asqrt28_0[1]));
	jspl3 jspl3_w_asqrt28_3(.douta(w_asqrt28_3[0]),.doutb(w_asqrt28_3[1]),.doutc(w_asqrt28_3[2]),.din(w_asqrt28_0[2]));
	jspl3 jspl3_w_asqrt28_4(.douta(w_asqrt28_4[0]),.doutb(w_asqrt28_4[1]),.doutc(w_asqrt28_4[2]),.din(w_asqrt28_1[0]));
	jspl3 jspl3_w_asqrt28_5(.douta(w_asqrt28_5[0]),.doutb(w_asqrt28_5[1]),.doutc(w_asqrt28_5[2]),.din(w_asqrt28_1[1]));
	jspl3 jspl3_w_asqrt28_6(.douta(w_asqrt28_6[0]),.doutb(w_asqrt28_6[1]),.doutc(w_asqrt28_6[2]),.din(w_asqrt28_1[2]));
	jspl3 jspl3_w_asqrt28_7(.douta(w_asqrt28_7[0]),.doutb(w_asqrt28_7[1]),.doutc(w_asqrt28_7[2]),.din(w_asqrt28_2[0]));
	jspl3 jspl3_w_asqrt28_8(.douta(w_asqrt28_8[0]),.doutb(w_asqrt28_8[1]),.doutc(w_asqrt28_8[2]),.din(w_asqrt28_2[1]));
	jspl3 jspl3_w_asqrt28_9(.douta(w_asqrt28_9[0]),.doutb(w_asqrt28_9[1]),.doutc(w_asqrt28_9[2]),.din(w_asqrt28_2[2]));
	jspl3 jspl3_w_asqrt28_10(.douta(w_asqrt28_10[0]),.doutb(w_asqrt28_10[1]),.doutc(w_asqrt28_10[2]),.din(w_asqrt28_3[0]));
	jspl3 jspl3_w_asqrt28_11(.douta(w_asqrt28_11[0]),.doutb(w_asqrt28_11[1]),.doutc(w_asqrt28_11[2]),.din(w_asqrt28_3[1]));
	jspl3 jspl3_w_asqrt28_12(.douta(w_asqrt28_12[0]),.doutb(w_asqrt28_12[1]),.doutc(w_asqrt28_12[2]),.din(w_asqrt28_3[2]));
	jspl3 jspl3_w_asqrt28_13(.douta(w_asqrt28_13[0]),.doutb(w_asqrt28_13[1]),.doutc(w_asqrt28_13[2]),.din(w_asqrt28_4[0]));
	jspl3 jspl3_w_asqrt28_14(.douta(w_asqrt28_14[0]),.doutb(w_asqrt28_14[1]),.doutc(w_asqrt28_14[2]),.din(w_asqrt28_4[1]));
	jspl3 jspl3_w_asqrt28_15(.douta(w_asqrt28_15[0]),.doutb(w_asqrt28_15[1]),.doutc(w_asqrt28_15[2]),.din(w_asqrt28_4[2]));
	jspl3 jspl3_w_asqrt28_16(.douta(w_asqrt28_16[0]),.doutb(w_asqrt28_16[1]),.doutc(w_asqrt28_16[2]),.din(w_asqrt28_5[0]));
	jspl3 jspl3_w_asqrt28_17(.douta(w_asqrt28_17[0]),.doutb(w_asqrt28_17[1]),.doutc(w_asqrt28_17[2]),.din(w_asqrt28_5[1]));
	jspl3 jspl3_w_asqrt28_18(.douta(w_asqrt28_18[0]),.doutb(w_asqrt28_18[1]),.doutc(w_asqrt28_18[2]),.din(w_asqrt28_5[2]));
	jspl3 jspl3_w_asqrt28_19(.douta(w_asqrt28_19[0]),.doutb(w_asqrt28_19[1]),.doutc(w_asqrt28_19[2]),.din(w_asqrt28_6[0]));
	jspl3 jspl3_w_asqrt28_20(.douta(w_asqrt28_20[0]),.doutb(w_asqrt28_20[1]),.doutc(w_asqrt28_20[2]),.din(w_asqrt28_6[1]));
	jspl3 jspl3_w_asqrt28_21(.douta(w_asqrt28_21[0]),.doutb(w_asqrt28_21[1]),.doutc(w_asqrt28_21[2]),.din(w_asqrt28_6[2]));
	jspl3 jspl3_w_asqrt28_22(.douta(w_asqrt28_22[0]),.doutb(w_asqrt28_22[1]),.doutc(w_asqrt28_22[2]),.din(w_asqrt28_7[0]));
	jspl3 jspl3_w_asqrt28_23(.douta(w_asqrt28_23[0]),.doutb(w_asqrt28_23[1]),.doutc(w_asqrt28_23[2]),.din(w_asqrt28_7[1]));
	jspl3 jspl3_w_asqrt28_24(.douta(w_asqrt28_24[0]),.doutb(w_asqrt28_24[1]),.doutc(w_asqrt28_24[2]),.din(w_asqrt28_7[2]));
	jspl3 jspl3_w_asqrt28_25(.douta(w_asqrt28_25[0]),.doutb(w_asqrt28_25[1]),.doutc(w_asqrt28_25[2]),.din(w_asqrt28_8[0]));
	jspl3 jspl3_w_asqrt28_26(.douta(w_asqrt28_26[0]),.doutb(w_asqrt28_26[1]),.doutc(w_asqrt28_26[2]),.din(w_asqrt28_8[1]));
	jspl3 jspl3_w_asqrt28_27(.douta(w_asqrt28_27[0]),.doutb(w_asqrt28_27[1]),.doutc(w_asqrt28_27[2]),.din(w_asqrt28_8[2]));
	jspl3 jspl3_w_asqrt28_28(.douta(w_asqrt28_28[0]),.doutb(w_asqrt28_28[1]),.doutc(w_asqrt28_28[2]),.din(w_asqrt28_9[0]));
	jspl3 jspl3_w_asqrt28_29(.douta(w_asqrt28_29[0]),.doutb(w_asqrt28_29[1]),.doutc(w_asqrt28_29[2]),.din(w_asqrt28_9[1]));
	jspl3 jspl3_w_asqrt28_30(.douta(w_asqrt28_30[0]),.doutb(w_asqrt28_30[1]),.doutc(w_asqrt28_30[2]),.din(w_asqrt28_9[2]));
	jspl jspl_w_asqrt28_31(.douta(w_asqrt28_31),.doutb(asqrt[27]),.din(w_asqrt28_10[0]));
	jspl3 jspl3_w_asqrt29_0(.douta(w_asqrt29_0[0]),.doutb(w_asqrt29_0[1]),.doutc(w_asqrt29_0[2]),.din(asqrt_fa_29));
	jspl3 jspl3_w_asqrt29_1(.douta(w_asqrt29_1[0]),.doutb(w_asqrt29_1[1]),.doutc(w_asqrt29_1[2]),.din(w_asqrt29_0[0]));
	jspl3 jspl3_w_asqrt29_2(.douta(w_asqrt29_2[0]),.doutb(w_asqrt29_2[1]),.doutc(w_asqrt29_2[2]),.din(w_asqrt29_0[1]));
	jspl3 jspl3_w_asqrt29_3(.douta(w_asqrt29_3[0]),.doutb(w_asqrt29_3[1]),.doutc(w_asqrt29_3[2]),.din(w_asqrt29_0[2]));
	jspl3 jspl3_w_asqrt29_4(.douta(w_asqrt29_4[0]),.doutb(w_asqrt29_4[1]),.doutc(w_asqrt29_4[2]),.din(w_asqrt29_1[0]));
	jspl3 jspl3_w_asqrt29_5(.douta(w_asqrt29_5[0]),.doutb(w_asqrt29_5[1]),.doutc(w_asqrt29_5[2]),.din(w_asqrt29_1[1]));
	jspl3 jspl3_w_asqrt29_6(.douta(w_asqrt29_6[0]),.doutb(w_asqrt29_6[1]),.doutc(w_asqrt29_6[2]),.din(w_asqrt29_1[2]));
	jspl3 jspl3_w_asqrt29_7(.douta(w_asqrt29_7[0]),.doutb(w_asqrt29_7[1]),.doutc(w_asqrt29_7[2]),.din(w_asqrt29_2[0]));
	jspl3 jspl3_w_asqrt29_8(.douta(w_asqrt29_8[0]),.doutb(w_asqrt29_8[1]),.doutc(w_asqrt29_8[2]),.din(w_asqrt29_2[1]));
	jspl3 jspl3_w_asqrt29_9(.douta(w_asqrt29_9[0]),.doutb(w_asqrt29_9[1]),.doutc(w_asqrt29_9[2]),.din(w_asqrt29_2[2]));
	jspl3 jspl3_w_asqrt29_10(.douta(w_asqrt29_10[0]),.doutb(w_asqrt29_10[1]),.doutc(w_asqrt29_10[2]),.din(w_asqrt29_3[0]));
	jspl3 jspl3_w_asqrt29_11(.douta(w_asqrt29_11[0]),.doutb(w_asqrt29_11[1]),.doutc(w_asqrt29_11[2]),.din(w_asqrt29_3[1]));
	jspl3 jspl3_w_asqrt29_12(.douta(w_asqrt29_12[0]),.doutb(w_asqrt29_12[1]),.doutc(w_asqrt29_12[2]),.din(w_asqrt29_3[2]));
	jspl3 jspl3_w_asqrt29_13(.douta(w_asqrt29_13[0]),.doutb(w_asqrt29_13[1]),.doutc(w_asqrt29_13[2]),.din(w_asqrt29_4[0]));
	jspl3 jspl3_w_asqrt29_14(.douta(w_asqrt29_14[0]),.doutb(w_asqrt29_14[1]),.doutc(w_asqrt29_14[2]),.din(w_asqrt29_4[1]));
	jspl3 jspl3_w_asqrt29_15(.douta(w_asqrt29_15[0]),.doutb(w_asqrt29_15[1]),.doutc(w_asqrt29_15[2]),.din(w_asqrt29_4[2]));
	jspl3 jspl3_w_asqrt29_16(.douta(w_asqrt29_16[0]),.doutb(w_asqrt29_16[1]),.doutc(w_asqrt29_16[2]),.din(w_asqrt29_5[0]));
	jspl3 jspl3_w_asqrt29_17(.douta(w_asqrt29_17[0]),.doutb(w_asqrt29_17[1]),.doutc(w_asqrt29_17[2]),.din(w_asqrt29_5[1]));
	jspl3 jspl3_w_asqrt29_18(.douta(w_asqrt29_18[0]),.doutb(w_asqrt29_18[1]),.doutc(w_asqrt29_18[2]),.din(w_asqrt29_5[2]));
	jspl3 jspl3_w_asqrt29_19(.douta(w_asqrt29_19[0]),.doutb(w_asqrt29_19[1]),.doutc(w_asqrt29_19[2]),.din(w_asqrt29_6[0]));
	jspl3 jspl3_w_asqrt29_20(.douta(w_asqrt29_20[0]),.doutb(w_asqrt29_20[1]),.doutc(w_asqrt29_20[2]),.din(w_asqrt29_6[1]));
	jspl3 jspl3_w_asqrt29_21(.douta(w_asqrt29_21[0]),.doutb(w_asqrt29_21[1]),.doutc(asqrt[28]),.din(w_asqrt29_6[2]));
	jspl3 jspl3_w_asqrt30_0(.douta(w_asqrt30_0[0]),.doutb(w_asqrt30_0[1]),.doutc(w_asqrt30_0[2]),.din(asqrt_fa_30));
	jspl3 jspl3_w_asqrt30_1(.douta(w_asqrt30_1[0]),.doutb(w_asqrt30_1[1]),.doutc(w_asqrt30_1[2]),.din(w_asqrt30_0[0]));
	jspl3 jspl3_w_asqrt30_2(.douta(w_asqrt30_2[0]),.doutb(w_asqrt30_2[1]),.doutc(w_asqrt30_2[2]),.din(w_asqrt30_0[1]));
	jspl3 jspl3_w_asqrt30_3(.douta(w_asqrt30_3[0]),.doutb(w_asqrt30_3[1]),.doutc(w_asqrt30_3[2]),.din(w_asqrt30_0[2]));
	jspl3 jspl3_w_asqrt30_4(.douta(w_asqrt30_4[0]),.doutb(w_asqrt30_4[1]),.doutc(w_asqrt30_4[2]),.din(w_asqrt30_1[0]));
	jspl3 jspl3_w_asqrt30_5(.douta(w_asqrt30_5[0]),.doutb(w_asqrt30_5[1]),.doutc(w_asqrt30_5[2]),.din(w_asqrt30_1[1]));
	jspl3 jspl3_w_asqrt30_6(.douta(w_asqrt30_6[0]),.doutb(w_asqrt30_6[1]),.doutc(w_asqrt30_6[2]),.din(w_asqrt30_1[2]));
	jspl3 jspl3_w_asqrt30_7(.douta(w_asqrt30_7[0]),.doutb(w_asqrt30_7[1]),.doutc(w_asqrt30_7[2]),.din(w_asqrt30_2[0]));
	jspl3 jspl3_w_asqrt30_8(.douta(w_asqrt30_8[0]),.doutb(w_asqrt30_8[1]),.doutc(w_asqrt30_8[2]),.din(w_asqrt30_2[1]));
	jspl3 jspl3_w_asqrt30_9(.douta(w_asqrt30_9[0]),.doutb(w_asqrt30_9[1]),.doutc(w_asqrt30_9[2]),.din(w_asqrt30_2[2]));
	jspl3 jspl3_w_asqrt30_10(.douta(w_asqrt30_10[0]),.doutb(w_asqrt30_10[1]),.doutc(w_asqrt30_10[2]),.din(w_asqrt30_3[0]));
	jspl3 jspl3_w_asqrt30_11(.douta(w_asqrt30_11[0]),.doutb(w_asqrt30_11[1]),.doutc(w_asqrt30_11[2]),.din(w_asqrt30_3[1]));
	jspl3 jspl3_w_asqrt30_12(.douta(w_asqrt30_12[0]),.doutb(w_asqrt30_12[1]),.doutc(w_asqrt30_12[2]),.din(w_asqrt30_3[2]));
	jspl3 jspl3_w_asqrt30_13(.douta(w_asqrt30_13[0]),.doutb(w_asqrt30_13[1]),.doutc(w_asqrt30_13[2]),.din(w_asqrt30_4[0]));
	jspl3 jspl3_w_asqrt30_14(.douta(w_asqrt30_14[0]),.doutb(w_asqrt30_14[1]),.doutc(w_asqrt30_14[2]),.din(w_asqrt30_4[1]));
	jspl3 jspl3_w_asqrt30_15(.douta(w_asqrt30_15[0]),.doutb(w_asqrt30_15[1]),.doutc(w_asqrt30_15[2]),.din(w_asqrt30_4[2]));
	jspl3 jspl3_w_asqrt30_16(.douta(w_asqrt30_16[0]),.doutb(w_asqrt30_16[1]),.doutc(w_asqrt30_16[2]),.din(w_asqrt30_5[0]));
	jspl3 jspl3_w_asqrt30_17(.douta(w_asqrt30_17[0]),.doutb(w_asqrt30_17[1]),.doutc(w_asqrt30_17[2]),.din(w_asqrt30_5[1]));
	jspl3 jspl3_w_asqrt30_18(.douta(w_asqrt30_18[0]),.doutb(w_asqrt30_18[1]),.doutc(w_asqrt30_18[2]),.din(w_asqrt30_5[2]));
	jspl3 jspl3_w_asqrt30_19(.douta(w_asqrt30_19[0]),.doutb(w_asqrt30_19[1]),.doutc(w_asqrt30_19[2]),.din(w_asqrt30_6[0]));
	jspl3 jspl3_w_asqrt30_20(.douta(w_asqrt30_20[0]),.doutb(w_asqrt30_20[1]),.doutc(w_asqrt30_20[2]),.din(w_asqrt30_6[1]));
	jspl3 jspl3_w_asqrt30_21(.douta(w_asqrt30_21[0]),.doutb(w_asqrt30_21[1]),.doutc(w_asqrt30_21[2]),.din(w_asqrt30_6[2]));
	jspl3 jspl3_w_asqrt30_22(.douta(w_asqrt30_22[0]),.doutb(w_asqrt30_22[1]),.doutc(w_asqrt30_22[2]),.din(w_asqrt30_7[0]));
	jspl3 jspl3_w_asqrt30_23(.douta(w_asqrt30_23[0]),.doutb(w_asqrt30_23[1]),.doutc(w_asqrt30_23[2]),.din(w_asqrt30_7[1]));
	jspl3 jspl3_w_asqrt30_24(.douta(w_asqrt30_24[0]),.doutb(w_asqrt30_24[1]),.doutc(w_asqrt30_24[2]),.din(w_asqrt30_7[2]));
	jspl3 jspl3_w_asqrt30_25(.douta(w_asqrt30_25[0]),.doutb(w_asqrt30_25[1]),.doutc(w_asqrt30_25[2]),.din(w_asqrt30_8[0]));
	jspl3 jspl3_w_asqrt30_26(.douta(w_asqrt30_26[0]),.doutb(w_asqrt30_26[1]),.doutc(w_asqrt30_26[2]),.din(w_asqrt30_8[1]));
	jspl3 jspl3_w_asqrt30_27(.douta(w_asqrt30_27[0]),.doutb(w_asqrt30_27[1]),.doutc(w_asqrt30_27[2]),.din(w_asqrt30_8[2]));
	jspl3 jspl3_w_asqrt30_28(.douta(w_asqrt30_28[0]),.doutb(w_asqrt30_28[1]),.doutc(w_asqrt30_28[2]),.din(w_asqrt30_9[0]));
	jspl3 jspl3_w_asqrt30_29(.douta(w_asqrt30_29[0]),.doutb(w_asqrt30_29[1]),.doutc(w_asqrt30_29[2]),.din(w_asqrt30_9[1]));
	jspl3 jspl3_w_asqrt30_30(.douta(w_asqrt30_30[0]),.doutb(w_asqrt30_30[1]),.doutc(w_asqrt30_30[2]),.din(w_asqrt30_9[2]));
	jspl jspl_w_asqrt30_31(.douta(w_asqrt30_31),.doutb(asqrt[29]),.din(w_asqrt30_10[0]));
	jspl3 jspl3_w_asqrt31_0(.douta(w_asqrt31_0[0]),.doutb(w_asqrt31_0[1]),.doutc(w_asqrt31_0[2]),.din(asqrt_fa_31));
	jspl3 jspl3_w_asqrt31_1(.douta(w_asqrt31_1[0]),.doutb(w_asqrt31_1[1]),.doutc(w_asqrt31_1[2]),.din(w_asqrt31_0[0]));
	jspl3 jspl3_w_asqrt31_2(.douta(w_asqrt31_2[0]),.doutb(w_asqrt31_2[1]),.doutc(w_asqrt31_2[2]),.din(w_asqrt31_0[1]));
	jspl3 jspl3_w_asqrt31_3(.douta(w_asqrt31_3[0]),.doutb(w_asqrt31_3[1]),.doutc(w_asqrt31_3[2]),.din(w_asqrt31_0[2]));
	jspl3 jspl3_w_asqrt31_4(.douta(w_asqrt31_4[0]),.doutb(w_asqrt31_4[1]),.doutc(w_asqrt31_4[2]),.din(w_asqrt31_1[0]));
	jspl3 jspl3_w_asqrt31_5(.douta(w_asqrt31_5[0]),.doutb(w_asqrt31_5[1]),.doutc(w_asqrt31_5[2]),.din(w_asqrt31_1[1]));
	jspl3 jspl3_w_asqrt31_6(.douta(w_asqrt31_6[0]),.doutb(w_asqrt31_6[1]),.doutc(w_asqrt31_6[2]),.din(w_asqrt31_1[2]));
	jspl3 jspl3_w_asqrt31_7(.douta(w_asqrt31_7[0]),.doutb(w_asqrt31_7[1]),.doutc(w_asqrt31_7[2]),.din(w_asqrt31_2[0]));
	jspl3 jspl3_w_asqrt31_8(.douta(w_asqrt31_8[0]),.doutb(w_asqrt31_8[1]),.doutc(w_asqrt31_8[2]),.din(w_asqrt31_2[1]));
	jspl3 jspl3_w_asqrt31_9(.douta(w_asqrt31_9[0]),.doutb(w_asqrt31_9[1]),.doutc(w_asqrt31_9[2]),.din(w_asqrt31_2[2]));
	jspl3 jspl3_w_asqrt31_10(.douta(w_asqrt31_10[0]),.doutb(w_asqrt31_10[1]),.doutc(w_asqrt31_10[2]),.din(w_asqrt31_3[0]));
	jspl3 jspl3_w_asqrt31_11(.douta(w_asqrt31_11[0]),.doutb(w_asqrt31_11[1]),.doutc(w_asqrt31_11[2]),.din(w_asqrt31_3[1]));
	jspl3 jspl3_w_asqrt31_12(.douta(w_asqrt31_12[0]),.doutb(w_asqrt31_12[1]),.doutc(w_asqrt31_12[2]),.din(w_asqrt31_3[2]));
	jspl3 jspl3_w_asqrt31_13(.douta(w_asqrt31_13[0]),.doutb(w_asqrt31_13[1]),.doutc(w_asqrt31_13[2]),.din(w_asqrt31_4[0]));
	jspl3 jspl3_w_asqrt31_14(.douta(w_asqrt31_14[0]),.doutb(w_asqrt31_14[1]),.doutc(w_asqrt31_14[2]),.din(w_asqrt31_4[1]));
	jspl3 jspl3_w_asqrt31_15(.douta(w_asqrt31_15[0]),.doutb(w_asqrt31_15[1]),.doutc(w_asqrt31_15[2]),.din(w_asqrt31_4[2]));
	jspl3 jspl3_w_asqrt31_16(.douta(w_asqrt31_16[0]),.doutb(w_asqrt31_16[1]),.doutc(w_asqrt31_16[2]),.din(w_asqrt31_5[0]));
	jspl3 jspl3_w_asqrt31_17(.douta(w_asqrt31_17[0]),.doutb(w_asqrt31_17[1]),.doutc(w_asqrt31_17[2]),.din(w_asqrt31_5[1]));
	jspl3 jspl3_w_asqrt31_18(.douta(w_asqrt31_18[0]),.doutb(w_asqrt31_18[1]),.doutc(w_asqrt31_18[2]),.din(w_asqrt31_5[2]));
	jspl3 jspl3_w_asqrt31_19(.douta(w_asqrt31_19[0]),.doutb(w_asqrt31_19[1]),.doutc(w_asqrt31_19[2]),.din(w_asqrt31_6[0]));
	jspl3 jspl3_w_asqrt31_20(.douta(w_asqrt31_20[0]),.doutb(w_asqrt31_20[1]),.doutc(w_asqrt31_20[2]),.din(w_asqrt31_6[1]));
	jspl3 jspl3_w_asqrt31_21(.douta(w_asqrt31_21[0]),.doutb(w_asqrt31_21[1]),.doutc(asqrt[30]),.din(w_asqrt31_6[2]));
	jspl3 jspl3_w_asqrt32_0(.douta(w_asqrt32_0[0]),.doutb(w_asqrt32_0[1]),.doutc(w_asqrt32_0[2]),.din(asqrt_fa_32));
	jspl3 jspl3_w_asqrt32_1(.douta(w_asqrt32_1[0]),.doutb(w_asqrt32_1[1]),.doutc(w_asqrt32_1[2]),.din(w_asqrt32_0[0]));
	jspl3 jspl3_w_asqrt32_2(.douta(w_asqrt32_2[0]),.doutb(w_asqrt32_2[1]),.doutc(w_asqrt32_2[2]),.din(w_asqrt32_0[1]));
	jspl3 jspl3_w_asqrt32_3(.douta(w_asqrt32_3[0]),.doutb(w_asqrt32_3[1]),.doutc(w_asqrt32_3[2]),.din(w_asqrt32_0[2]));
	jspl3 jspl3_w_asqrt32_4(.douta(w_asqrt32_4[0]),.doutb(w_asqrt32_4[1]),.doutc(w_asqrt32_4[2]),.din(w_asqrt32_1[0]));
	jspl3 jspl3_w_asqrt32_5(.douta(w_asqrt32_5[0]),.doutb(w_asqrt32_5[1]),.doutc(w_asqrt32_5[2]),.din(w_asqrt32_1[1]));
	jspl3 jspl3_w_asqrt32_6(.douta(w_asqrt32_6[0]),.doutb(w_asqrt32_6[1]),.doutc(w_asqrt32_6[2]),.din(w_asqrt32_1[2]));
	jspl3 jspl3_w_asqrt32_7(.douta(w_asqrt32_7[0]),.doutb(w_asqrt32_7[1]),.doutc(w_asqrt32_7[2]),.din(w_asqrt32_2[0]));
	jspl3 jspl3_w_asqrt32_8(.douta(w_asqrt32_8[0]),.doutb(w_asqrt32_8[1]),.doutc(w_asqrt32_8[2]),.din(w_asqrt32_2[1]));
	jspl3 jspl3_w_asqrt32_9(.douta(w_asqrt32_9[0]),.doutb(w_asqrt32_9[1]),.doutc(w_asqrt32_9[2]),.din(w_asqrt32_2[2]));
	jspl3 jspl3_w_asqrt32_10(.douta(w_asqrt32_10[0]),.doutb(w_asqrt32_10[1]),.doutc(w_asqrt32_10[2]),.din(w_asqrt32_3[0]));
	jspl3 jspl3_w_asqrt32_11(.douta(w_asqrt32_11[0]),.doutb(w_asqrt32_11[1]),.doutc(w_asqrt32_11[2]),.din(w_asqrt32_3[1]));
	jspl3 jspl3_w_asqrt32_12(.douta(w_asqrt32_12[0]),.doutb(w_asqrt32_12[1]),.doutc(w_asqrt32_12[2]),.din(w_asqrt32_3[2]));
	jspl3 jspl3_w_asqrt32_13(.douta(w_asqrt32_13[0]),.doutb(w_asqrt32_13[1]),.doutc(w_asqrt32_13[2]),.din(w_asqrt32_4[0]));
	jspl3 jspl3_w_asqrt32_14(.douta(w_asqrt32_14[0]),.doutb(w_asqrt32_14[1]),.doutc(w_asqrt32_14[2]),.din(w_asqrt32_4[1]));
	jspl3 jspl3_w_asqrt32_15(.douta(w_asqrt32_15[0]),.doutb(w_asqrt32_15[1]),.doutc(w_asqrt32_15[2]),.din(w_asqrt32_4[2]));
	jspl3 jspl3_w_asqrt32_16(.douta(w_asqrt32_16[0]),.doutb(w_asqrt32_16[1]),.doutc(w_asqrt32_16[2]),.din(w_asqrt32_5[0]));
	jspl3 jspl3_w_asqrt32_17(.douta(w_asqrt32_17[0]),.doutb(w_asqrt32_17[1]),.doutc(w_asqrt32_17[2]),.din(w_asqrt32_5[1]));
	jspl3 jspl3_w_asqrt32_18(.douta(w_asqrt32_18[0]),.doutb(w_asqrt32_18[1]),.doutc(w_asqrt32_18[2]),.din(w_asqrt32_5[2]));
	jspl3 jspl3_w_asqrt32_19(.douta(w_asqrt32_19[0]),.doutb(w_asqrt32_19[1]),.doutc(w_asqrt32_19[2]),.din(w_asqrt32_6[0]));
	jspl3 jspl3_w_asqrt32_20(.douta(w_asqrt32_20[0]),.doutb(w_asqrt32_20[1]),.doutc(w_asqrt32_20[2]),.din(w_asqrt32_6[1]));
	jspl3 jspl3_w_asqrt32_21(.douta(w_asqrt32_21[0]),.doutb(w_asqrt32_21[1]),.doutc(w_asqrt32_21[2]),.din(w_asqrt32_6[2]));
	jspl3 jspl3_w_asqrt32_22(.douta(w_asqrt32_22[0]),.doutb(w_asqrt32_22[1]),.doutc(w_asqrt32_22[2]),.din(w_asqrt32_7[0]));
	jspl3 jspl3_w_asqrt32_23(.douta(w_asqrt32_23[0]),.doutb(w_asqrt32_23[1]),.doutc(w_asqrt32_23[2]),.din(w_asqrt32_7[1]));
	jspl3 jspl3_w_asqrt32_24(.douta(w_asqrt32_24[0]),.doutb(w_asqrt32_24[1]),.doutc(w_asqrt32_24[2]),.din(w_asqrt32_7[2]));
	jspl3 jspl3_w_asqrt32_25(.douta(w_asqrt32_25[0]),.doutb(w_asqrt32_25[1]),.doutc(w_asqrt32_25[2]),.din(w_asqrt32_8[0]));
	jspl3 jspl3_w_asqrt32_26(.douta(w_asqrt32_26[0]),.doutb(w_asqrt32_26[1]),.doutc(w_asqrt32_26[2]),.din(w_asqrt32_8[1]));
	jspl3 jspl3_w_asqrt32_27(.douta(w_asqrt32_27[0]),.doutb(w_asqrt32_27[1]),.doutc(w_asqrt32_27[2]),.din(w_asqrt32_8[2]));
	jspl3 jspl3_w_asqrt32_28(.douta(w_asqrt32_28[0]),.doutb(w_asqrt32_28[1]),.doutc(w_asqrt32_28[2]),.din(w_asqrt32_9[0]));
	jspl3 jspl3_w_asqrt32_29(.douta(w_asqrt32_29[0]),.doutb(w_asqrt32_29[1]),.doutc(w_asqrt32_29[2]),.din(w_asqrt32_9[1]));
	jspl3 jspl3_w_asqrt32_30(.douta(w_asqrt32_30[0]),.doutb(w_asqrt32_30[1]),.doutc(w_asqrt32_30[2]),.din(w_asqrt32_9[2]));
	jspl jspl_w_asqrt32_31(.douta(w_asqrt32_31),.doutb(asqrt[31]),.din(w_asqrt32_10[0]));
	jspl3 jspl3_w_asqrt33_0(.douta(w_asqrt33_0[0]),.doutb(w_asqrt33_0[1]),.doutc(w_asqrt33_0[2]),.din(asqrt_fa_33));
	jspl3 jspl3_w_asqrt33_1(.douta(w_asqrt33_1[0]),.doutb(w_asqrt33_1[1]),.doutc(w_asqrt33_1[2]),.din(w_asqrt33_0[0]));
	jspl3 jspl3_w_asqrt33_2(.douta(w_asqrt33_2[0]),.doutb(w_asqrt33_2[1]),.doutc(w_asqrt33_2[2]),.din(w_asqrt33_0[1]));
	jspl3 jspl3_w_asqrt33_3(.douta(w_asqrt33_3[0]),.doutb(w_asqrt33_3[1]),.doutc(w_asqrt33_3[2]),.din(w_asqrt33_0[2]));
	jspl3 jspl3_w_asqrt33_4(.douta(w_asqrt33_4[0]),.doutb(w_asqrt33_4[1]),.doutc(w_asqrt33_4[2]),.din(w_asqrt33_1[0]));
	jspl3 jspl3_w_asqrt33_5(.douta(w_asqrt33_5[0]),.doutb(w_asqrt33_5[1]),.doutc(w_asqrt33_5[2]),.din(w_asqrt33_1[1]));
	jspl3 jspl3_w_asqrt33_6(.douta(w_asqrt33_6[0]),.doutb(w_asqrt33_6[1]),.doutc(w_asqrt33_6[2]),.din(w_asqrt33_1[2]));
	jspl3 jspl3_w_asqrt33_7(.douta(w_asqrt33_7[0]),.doutb(w_asqrt33_7[1]),.doutc(w_asqrt33_7[2]),.din(w_asqrt33_2[0]));
	jspl3 jspl3_w_asqrt33_8(.douta(w_asqrt33_8[0]),.doutb(w_asqrt33_8[1]),.doutc(w_asqrt33_8[2]),.din(w_asqrt33_2[1]));
	jspl3 jspl3_w_asqrt33_9(.douta(w_asqrt33_9[0]),.doutb(w_asqrt33_9[1]),.doutc(w_asqrt33_9[2]),.din(w_asqrt33_2[2]));
	jspl3 jspl3_w_asqrt33_10(.douta(w_asqrt33_10[0]),.doutb(w_asqrt33_10[1]),.doutc(w_asqrt33_10[2]),.din(w_asqrt33_3[0]));
	jspl3 jspl3_w_asqrt33_11(.douta(w_asqrt33_11[0]),.doutb(w_asqrt33_11[1]),.doutc(w_asqrt33_11[2]),.din(w_asqrt33_3[1]));
	jspl3 jspl3_w_asqrt33_12(.douta(w_asqrt33_12[0]),.doutb(w_asqrt33_12[1]),.doutc(w_asqrt33_12[2]),.din(w_asqrt33_3[2]));
	jspl3 jspl3_w_asqrt33_13(.douta(w_asqrt33_13[0]),.doutb(w_asqrt33_13[1]),.doutc(w_asqrt33_13[2]),.din(w_asqrt33_4[0]));
	jspl3 jspl3_w_asqrt33_14(.douta(w_asqrt33_14[0]),.doutb(w_asqrt33_14[1]),.doutc(w_asqrt33_14[2]),.din(w_asqrt33_4[1]));
	jspl3 jspl3_w_asqrt33_15(.douta(w_asqrt33_15[0]),.doutb(w_asqrt33_15[1]),.doutc(w_asqrt33_15[2]),.din(w_asqrt33_4[2]));
	jspl3 jspl3_w_asqrt33_16(.douta(w_asqrt33_16[0]),.doutb(w_asqrt33_16[1]),.doutc(w_asqrt33_16[2]),.din(w_asqrt33_5[0]));
	jspl3 jspl3_w_asqrt33_17(.douta(w_asqrt33_17[0]),.doutb(w_asqrt33_17[1]),.doutc(w_asqrt33_17[2]),.din(w_asqrt33_5[1]));
	jspl3 jspl3_w_asqrt33_18(.douta(w_asqrt33_18[0]),.doutb(w_asqrt33_18[1]),.doutc(w_asqrt33_18[2]),.din(w_asqrt33_5[2]));
	jspl3 jspl3_w_asqrt33_19(.douta(w_asqrt33_19[0]),.doutb(w_asqrt33_19[1]),.doutc(w_asqrt33_19[2]),.din(w_asqrt33_6[0]));
	jspl3 jspl3_w_asqrt33_20(.douta(w_asqrt33_20[0]),.doutb(w_asqrt33_20[1]),.doutc(w_asqrt33_20[2]),.din(w_asqrt33_6[1]));
	jspl3 jspl3_w_asqrt33_21(.douta(w_asqrt33_21[0]),.doutb(w_asqrt33_21[1]),.doutc(w_asqrt33_21[2]),.din(w_asqrt33_6[2]));
	jspl3 jspl3_w_asqrt33_22(.douta(w_asqrt33_22[0]),.doutb(w_asqrt33_22[1]),.doutc(asqrt[32]),.din(w_asqrt33_7[0]));
	jspl3 jspl3_w_asqrt34_0(.douta(w_asqrt34_0[0]),.doutb(w_asqrt34_0[1]),.doutc(w_asqrt34_0[2]),.din(asqrt_fa_34));
	jspl3 jspl3_w_asqrt34_1(.douta(w_asqrt34_1[0]),.doutb(w_asqrt34_1[1]),.doutc(w_asqrt34_1[2]),.din(w_asqrt34_0[0]));
	jspl3 jspl3_w_asqrt34_2(.douta(w_asqrt34_2[0]),.doutb(w_asqrt34_2[1]),.doutc(w_asqrt34_2[2]),.din(w_asqrt34_0[1]));
	jspl3 jspl3_w_asqrt34_3(.douta(w_asqrt34_3[0]),.doutb(w_asqrt34_3[1]),.doutc(w_asqrt34_3[2]),.din(w_asqrt34_0[2]));
	jspl3 jspl3_w_asqrt34_4(.douta(w_asqrt34_4[0]),.doutb(w_asqrt34_4[1]),.doutc(w_asqrt34_4[2]),.din(w_asqrt34_1[0]));
	jspl3 jspl3_w_asqrt34_5(.douta(w_asqrt34_5[0]),.doutb(w_asqrt34_5[1]),.doutc(w_asqrt34_5[2]),.din(w_asqrt34_1[1]));
	jspl3 jspl3_w_asqrt34_6(.douta(w_asqrt34_6[0]),.doutb(w_asqrt34_6[1]),.doutc(w_asqrt34_6[2]),.din(w_asqrt34_1[2]));
	jspl3 jspl3_w_asqrt34_7(.douta(w_asqrt34_7[0]),.doutb(w_asqrt34_7[1]),.doutc(w_asqrt34_7[2]),.din(w_asqrt34_2[0]));
	jspl3 jspl3_w_asqrt34_8(.douta(w_asqrt34_8[0]),.doutb(w_asqrt34_8[1]),.doutc(w_asqrt34_8[2]),.din(w_asqrt34_2[1]));
	jspl3 jspl3_w_asqrt34_9(.douta(w_asqrt34_9[0]),.doutb(w_asqrt34_9[1]),.doutc(w_asqrt34_9[2]),.din(w_asqrt34_2[2]));
	jspl3 jspl3_w_asqrt34_10(.douta(w_asqrt34_10[0]),.doutb(w_asqrt34_10[1]),.doutc(w_asqrt34_10[2]),.din(w_asqrt34_3[0]));
	jspl3 jspl3_w_asqrt34_11(.douta(w_asqrt34_11[0]),.doutb(w_asqrt34_11[1]),.doutc(w_asqrt34_11[2]),.din(w_asqrt34_3[1]));
	jspl3 jspl3_w_asqrt34_12(.douta(w_asqrt34_12[0]),.doutb(w_asqrt34_12[1]),.doutc(w_asqrt34_12[2]),.din(w_asqrt34_3[2]));
	jspl3 jspl3_w_asqrt34_13(.douta(w_asqrt34_13[0]),.doutb(w_asqrt34_13[1]),.doutc(w_asqrt34_13[2]),.din(w_asqrt34_4[0]));
	jspl3 jspl3_w_asqrt34_14(.douta(w_asqrt34_14[0]),.doutb(w_asqrt34_14[1]),.doutc(w_asqrt34_14[2]),.din(w_asqrt34_4[1]));
	jspl3 jspl3_w_asqrt34_15(.douta(w_asqrt34_15[0]),.doutb(w_asqrt34_15[1]),.doutc(w_asqrt34_15[2]),.din(w_asqrt34_4[2]));
	jspl3 jspl3_w_asqrt34_16(.douta(w_asqrt34_16[0]),.doutb(w_asqrt34_16[1]),.doutc(w_asqrt34_16[2]),.din(w_asqrt34_5[0]));
	jspl3 jspl3_w_asqrt34_17(.douta(w_asqrt34_17[0]),.doutb(w_asqrt34_17[1]),.doutc(w_asqrt34_17[2]),.din(w_asqrt34_5[1]));
	jspl3 jspl3_w_asqrt34_18(.douta(w_asqrt34_18[0]),.doutb(w_asqrt34_18[1]),.doutc(w_asqrt34_18[2]),.din(w_asqrt34_5[2]));
	jspl3 jspl3_w_asqrt34_19(.douta(w_asqrt34_19[0]),.doutb(w_asqrt34_19[1]),.doutc(w_asqrt34_19[2]),.din(w_asqrt34_6[0]));
	jspl3 jspl3_w_asqrt34_20(.douta(w_asqrt34_20[0]),.doutb(w_asqrt34_20[1]),.doutc(w_asqrt34_20[2]),.din(w_asqrt34_6[1]));
	jspl3 jspl3_w_asqrt34_21(.douta(w_asqrt34_21[0]),.doutb(w_asqrt34_21[1]),.doutc(w_asqrt34_21[2]),.din(w_asqrt34_6[2]));
	jspl3 jspl3_w_asqrt34_22(.douta(w_asqrt34_22[0]),.doutb(w_asqrt34_22[1]),.doutc(w_asqrt34_22[2]),.din(w_asqrt34_7[0]));
	jspl3 jspl3_w_asqrt34_23(.douta(w_asqrt34_23[0]),.doutb(w_asqrt34_23[1]),.doutc(w_asqrt34_23[2]),.din(w_asqrt34_7[1]));
	jspl3 jspl3_w_asqrt34_24(.douta(w_asqrt34_24[0]),.doutb(w_asqrt34_24[1]),.doutc(w_asqrt34_24[2]),.din(w_asqrt34_7[2]));
	jspl3 jspl3_w_asqrt34_25(.douta(w_asqrt34_25[0]),.doutb(w_asqrt34_25[1]),.doutc(w_asqrt34_25[2]),.din(w_asqrt34_8[0]));
	jspl3 jspl3_w_asqrt34_26(.douta(w_asqrt34_26[0]),.doutb(w_asqrt34_26[1]),.doutc(w_asqrt34_26[2]),.din(w_asqrt34_8[1]));
	jspl3 jspl3_w_asqrt34_27(.douta(w_asqrt34_27[0]),.doutb(w_asqrt34_27[1]),.doutc(w_asqrt34_27[2]),.din(w_asqrt34_8[2]));
	jspl3 jspl3_w_asqrt34_28(.douta(w_asqrt34_28[0]),.doutb(w_asqrt34_28[1]),.doutc(w_asqrt34_28[2]),.din(w_asqrt34_9[0]));
	jspl3 jspl3_w_asqrt34_29(.douta(w_asqrt34_29[0]),.doutb(w_asqrt34_29[1]),.doutc(w_asqrt34_29[2]),.din(w_asqrt34_9[1]));
	jspl3 jspl3_w_asqrt34_30(.douta(w_asqrt34_30[0]),.doutb(w_asqrt34_30[1]),.doutc(w_asqrt34_30[2]),.din(w_asqrt34_9[2]));
	jspl jspl_w_asqrt34_31(.douta(w_asqrt34_31),.doutb(asqrt[33]),.din(w_asqrt34_10[0]));
	jspl3 jspl3_w_asqrt35_0(.douta(w_asqrt35_0[0]),.doutb(w_asqrt35_0[1]),.doutc(w_asqrt35_0[2]),.din(asqrt_fa_35));
	jspl3 jspl3_w_asqrt35_1(.douta(w_asqrt35_1[0]),.doutb(w_asqrt35_1[1]),.doutc(w_asqrt35_1[2]),.din(w_asqrt35_0[0]));
	jspl3 jspl3_w_asqrt35_2(.douta(w_asqrt35_2[0]),.doutb(w_asqrt35_2[1]),.doutc(w_asqrt35_2[2]),.din(w_asqrt35_0[1]));
	jspl3 jspl3_w_asqrt35_3(.douta(w_asqrt35_3[0]),.doutb(w_asqrt35_3[1]),.doutc(w_asqrt35_3[2]),.din(w_asqrt35_0[2]));
	jspl3 jspl3_w_asqrt35_4(.douta(w_asqrt35_4[0]),.doutb(w_asqrt35_4[1]),.doutc(w_asqrt35_4[2]),.din(w_asqrt35_1[0]));
	jspl3 jspl3_w_asqrt35_5(.douta(w_asqrt35_5[0]),.doutb(w_asqrt35_5[1]),.doutc(w_asqrt35_5[2]),.din(w_asqrt35_1[1]));
	jspl3 jspl3_w_asqrt35_6(.douta(w_asqrt35_6[0]),.doutb(w_asqrt35_6[1]),.doutc(w_asqrt35_6[2]),.din(w_asqrt35_1[2]));
	jspl3 jspl3_w_asqrt35_7(.douta(w_asqrt35_7[0]),.doutb(w_asqrt35_7[1]),.doutc(w_asqrt35_7[2]),.din(w_asqrt35_2[0]));
	jspl3 jspl3_w_asqrt35_8(.douta(w_asqrt35_8[0]),.doutb(w_asqrt35_8[1]),.doutc(w_asqrt35_8[2]),.din(w_asqrt35_2[1]));
	jspl3 jspl3_w_asqrt35_9(.douta(w_asqrt35_9[0]),.doutb(w_asqrt35_9[1]),.doutc(w_asqrt35_9[2]),.din(w_asqrt35_2[2]));
	jspl3 jspl3_w_asqrt35_10(.douta(w_asqrt35_10[0]),.doutb(w_asqrt35_10[1]),.doutc(w_asqrt35_10[2]),.din(w_asqrt35_3[0]));
	jspl3 jspl3_w_asqrt35_11(.douta(w_asqrt35_11[0]),.doutb(w_asqrt35_11[1]),.doutc(w_asqrt35_11[2]),.din(w_asqrt35_3[1]));
	jspl3 jspl3_w_asqrt35_12(.douta(w_asqrt35_12[0]),.doutb(w_asqrt35_12[1]),.doutc(w_asqrt35_12[2]),.din(w_asqrt35_3[2]));
	jspl3 jspl3_w_asqrt35_13(.douta(w_asqrt35_13[0]),.doutb(w_asqrt35_13[1]),.doutc(w_asqrt35_13[2]),.din(w_asqrt35_4[0]));
	jspl3 jspl3_w_asqrt35_14(.douta(w_asqrt35_14[0]),.doutb(w_asqrt35_14[1]),.doutc(w_asqrt35_14[2]),.din(w_asqrt35_4[1]));
	jspl3 jspl3_w_asqrt35_15(.douta(w_asqrt35_15[0]),.doutb(w_asqrt35_15[1]),.doutc(w_asqrt35_15[2]),.din(w_asqrt35_4[2]));
	jspl3 jspl3_w_asqrt35_16(.douta(w_asqrt35_16[0]),.doutb(w_asqrt35_16[1]),.doutc(w_asqrt35_16[2]),.din(w_asqrt35_5[0]));
	jspl3 jspl3_w_asqrt35_17(.douta(w_asqrt35_17[0]),.doutb(w_asqrt35_17[1]),.doutc(w_asqrt35_17[2]),.din(w_asqrt35_5[1]));
	jspl3 jspl3_w_asqrt35_18(.douta(w_asqrt35_18[0]),.doutb(w_asqrt35_18[1]),.doutc(w_asqrt35_18[2]),.din(w_asqrt35_5[2]));
	jspl3 jspl3_w_asqrt35_19(.douta(w_asqrt35_19[0]),.doutb(w_asqrt35_19[1]),.doutc(w_asqrt35_19[2]),.din(w_asqrt35_6[0]));
	jspl3 jspl3_w_asqrt35_20(.douta(w_asqrt35_20[0]),.doutb(w_asqrt35_20[1]),.doutc(w_asqrt35_20[2]),.din(w_asqrt35_6[1]));
	jspl3 jspl3_w_asqrt35_21(.douta(w_asqrt35_21[0]),.doutb(w_asqrt35_21[1]),.doutc(w_asqrt35_21[2]),.din(w_asqrt35_6[2]));
	jspl3 jspl3_w_asqrt35_22(.douta(w_asqrt35_22[0]),.doutb(w_asqrt35_22[1]),.doutc(asqrt[34]),.din(w_asqrt35_7[0]));
	jspl3 jspl3_w_asqrt36_0(.douta(w_asqrt36_0[0]),.doutb(w_asqrt36_0[1]),.doutc(w_asqrt36_0[2]),.din(asqrt_fa_36));
	jspl3 jspl3_w_asqrt36_1(.douta(w_asqrt36_1[0]),.doutb(w_asqrt36_1[1]),.doutc(w_asqrt36_1[2]),.din(w_asqrt36_0[0]));
	jspl3 jspl3_w_asqrt36_2(.douta(w_asqrt36_2[0]),.doutb(w_asqrt36_2[1]),.doutc(w_asqrt36_2[2]),.din(w_asqrt36_0[1]));
	jspl3 jspl3_w_asqrt36_3(.douta(w_asqrt36_3[0]),.doutb(w_asqrt36_3[1]),.doutc(w_asqrt36_3[2]),.din(w_asqrt36_0[2]));
	jspl3 jspl3_w_asqrt36_4(.douta(w_asqrt36_4[0]),.doutb(w_asqrt36_4[1]),.doutc(w_asqrt36_4[2]),.din(w_asqrt36_1[0]));
	jspl3 jspl3_w_asqrt36_5(.douta(w_asqrt36_5[0]),.doutb(w_asqrt36_5[1]),.doutc(w_asqrt36_5[2]),.din(w_asqrt36_1[1]));
	jspl3 jspl3_w_asqrt36_6(.douta(w_asqrt36_6[0]),.doutb(w_asqrt36_6[1]),.doutc(w_asqrt36_6[2]),.din(w_asqrt36_1[2]));
	jspl3 jspl3_w_asqrt36_7(.douta(w_asqrt36_7[0]),.doutb(w_asqrt36_7[1]),.doutc(w_asqrt36_7[2]),.din(w_asqrt36_2[0]));
	jspl3 jspl3_w_asqrt36_8(.douta(w_asqrt36_8[0]),.doutb(w_asqrt36_8[1]),.doutc(w_asqrt36_8[2]),.din(w_asqrt36_2[1]));
	jspl3 jspl3_w_asqrt36_9(.douta(w_asqrt36_9[0]),.doutb(w_asqrt36_9[1]),.doutc(w_asqrt36_9[2]),.din(w_asqrt36_2[2]));
	jspl3 jspl3_w_asqrt36_10(.douta(w_asqrt36_10[0]),.doutb(w_asqrt36_10[1]),.doutc(w_asqrt36_10[2]),.din(w_asqrt36_3[0]));
	jspl3 jspl3_w_asqrt36_11(.douta(w_asqrt36_11[0]),.doutb(w_asqrt36_11[1]),.doutc(w_asqrt36_11[2]),.din(w_asqrt36_3[1]));
	jspl3 jspl3_w_asqrt36_12(.douta(w_asqrt36_12[0]),.doutb(w_asqrt36_12[1]),.doutc(w_asqrt36_12[2]),.din(w_asqrt36_3[2]));
	jspl3 jspl3_w_asqrt36_13(.douta(w_asqrt36_13[0]),.doutb(w_asqrt36_13[1]),.doutc(w_asqrt36_13[2]),.din(w_asqrt36_4[0]));
	jspl3 jspl3_w_asqrt36_14(.douta(w_asqrt36_14[0]),.doutb(w_asqrt36_14[1]),.doutc(w_asqrt36_14[2]),.din(w_asqrt36_4[1]));
	jspl3 jspl3_w_asqrt36_15(.douta(w_asqrt36_15[0]),.doutb(w_asqrt36_15[1]),.doutc(w_asqrt36_15[2]),.din(w_asqrt36_4[2]));
	jspl3 jspl3_w_asqrt36_16(.douta(w_asqrt36_16[0]),.doutb(w_asqrt36_16[1]),.doutc(w_asqrt36_16[2]),.din(w_asqrt36_5[0]));
	jspl3 jspl3_w_asqrt36_17(.douta(w_asqrt36_17[0]),.doutb(w_asqrt36_17[1]),.doutc(w_asqrt36_17[2]),.din(w_asqrt36_5[1]));
	jspl3 jspl3_w_asqrt36_18(.douta(w_asqrt36_18[0]),.doutb(w_asqrt36_18[1]),.doutc(w_asqrt36_18[2]),.din(w_asqrt36_5[2]));
	jspl3 jspl3_w_asqrt36_19(.douta(w_asqrt36_19[0]),.doutb(w_asqrt36_19[1]),.doutc(w_asqrt36_19[2]),.din(w_asqrt36_6[0]));
	jspl3 jspl3_w_asqrt36_20(.douta(w_asqrt36_20[0]),.doutb(w_asqrt36_20[1]),.doutc(w_asqrt36_20[2]),.din(w_asqrt36_6[1]));
	jspl3 jspl3_w_asqrt36_21(.douta(w_asqrt36_21[0]),.doutb(w_asqrt36_21[1]),.doutc(w_asqrt36_21[2]),.din(w_asqrt36_6[2]));
	jspl3 jspl3_w_asqrt36_22(.douta(w_asqrt36_22[0]),.doutb(w_asqrt36_22[1]),.doutc(w_asqrt36_22[2]),.din(w_asqrt36_7[0]));
	jspl3 jspl3_w_asqrt36_23(.douta(w_asqrt36_23[0]),.doutb(w_asqrt36_23[1]),.doutc(w_asqrt36_23[2]),.din(w_asqrt36_7[1]));
	jspl3 jspl3_w_asqrt36_24(.douta(w_asqrt36_24[0]),.doutb(w_asqrt36_24[1]),.doutc(w_asqrt36_24[2]),.din(w_asqrt36_7[2]));
	jspl3 jspl3_w_asqrt36_25(.douta(w_asqrt36_25[0]),.doutb(w_asqrt36_25[1]),.doutc(w_asqrt36_25[2]),.din(w_asqrt36_8[0]));
	jspl3 jspl3_w_asqrt36_26(.douta(w_asqrt36_26[0]),.doutb(w_asqrt36_26[1]),.doutc(w_asqrt36_26[2]),.din(w_asqrt36_8[1]));
	jspl3 jspl3_w_asqrt36_27(.douta(w_asqrt36_27[0]),.doutb(w_asqrt36_27[1]),.doutc(w_asqrt36_27[2]),.din(w_asqrt36_8[2]));
	jspl3 jspl3_w_asqrt36_28(.douta(w_asqrt36_28[0]),.doutb(w_asqrt36_28[1]),.doutc(w_asqrt36_28[2]),.din(w_asqrt36_9[0]));
	jspl3 jspl3_w_asqrt36_29(.douta(w_asqrt36_29[0]),.doutb(w_asqrt36_29[1]),.doutc(w_asqrt36_29[2]),.din(w_asqrt36_9[1]));
	jspl3 jspl3_w_asqrt36_30(.douta(w_asqrt36_30[0]),.doutb(w_asqrt36_30[1]),.doutc(w_asqrt36_30[2]),.din(w_asqrt36_9[2]));
	jspl jspl_w_asqrt36_31(.douta(w_asqrt36_31),.doutb(asqrt[35]),.din(w_asqrt36_10[0]));
	jspl3 jspl3_w_asqrt37_0(.douta(w_asqrt37_0[0]),.doutb(w_asqrt37_0[1]),.doutc(w_asqrt37_0[2]),.din(asqrt_fa_37));
	jspl3 jspl3_w_asqrt37_1(.douta(w_asqrt37_1[0]),.doutb(w_asqrt37_1[1]),.doutc(w_asqrt37_1[2]),.din(w_asqrt37_0[0]));
	jspl3 jspl3_w_asqrt37_2(.douta(w_asqrt37_2[0]),.doutb(w_asqrt37_2[1]),.doutc(w_asqrt37_2[2]),.din(w_asqrt37_0[1]));
	jspl3 jspl3_w_asqrt37_3(.douta(w_asqrt37_3[0]),.doutb(w_asqrt37_3[1]),.doutc(w_asqrt37_3[2]),.din(w_asqrt37_0[2]));
	jspl3 jspl3_w_asqrt37_4(.douta(w_asqrt37_4[0]),.doutb(w_asqrt37_4[1]),.doutc(w_asqrt37_4[2]),.din(w_asqrt37_1[0]));
	jspl3 jspl3_w_asqrt37_5(.douta(w_asqrt37_5[0]),.doutb(w_asqrt37_5[1]),.doutc(w_asqrt37_5[2]),.din(w_asqrt37_1[1]));
	jspl3 jspl3_w_asqrt37_6(.douta(w_asqrt37_6[0]),.doutb(w_asqrt37_6[1]),.doutc(w_asqrt37_6[2]),.din(w_asqrt37_1[2]));
	jspl3 jspl3_w_asqrt37_7(.douta(w_asqrt37_7[0]),.doutb(w_asqrt37_7[1]),.doutc(w_asqrt37_7[2]),.din(w_asqrt37_2[0]));
	jspl3 jspl3_w_asqrt37_8(.douta(w_asqrt37_8[0]),.doutb(w_asqrt37_8[1]),.doutc(w_asqrt37_8[2]),.din(w_asqrt37_2[1]));
	jspl3 jspl3_w_asqrt37_9(.douta(w_asqrt37_9[0]),.doutb(w_asqrt37_9[1]),.doutc(w_asqrt37_9[2]),.din(w_asqrt37_2[2]));
	jspl3 jspl3_w_asqrt37_10(.douta(w_asqrt37_10[0]),.doutb(w_asqrt37_10[1]),.doutc(w_asqrt37_10[2]),.din(w_asqrt37_3[0]));
	jspl3 jspl3_w_asqrt37_11(.douta(w_asqrt37_11[0]),.doutb(w_asqrt37_11[1]),.doutc(w_asqrt37_11[2]),.din(w_asqrt37_3[1]));
	jspl3 jspl3_w_asqrt37_12(.douta(w_asqrt37_12[0]),.doutb(w_asqrt37_12[1]),.doutc(w_asqrt37_12[2]),.din(w_asqrt37_3[2]));
	jspl3 jspl3_w_asqrt37_13(.douta(w_asqrt37_13[0]),.doutb(w_asqrt37_13[1]),.doutc(w_asqrt37_13[2]),.din(w_asqrt37_4[0]));
	jspl3 jspl3_w_asqrt37_14(.douta(w_asqrt37_14[0]),.doutb(w_asqrt37_14[1]),.doutc(w_asqrt37_14[2]),.din(w_asqrt37_4[1]));
	jspl3 jspl3_w_asqrt37_15(.douta(w_asqrt37_15[0]),.doutb(w_asqrt37_15[1]),.doutc(w_asqrt37_15[2]),.din(w_asqrt37_4[2]));
	jspl3 jspl3_w_asqrt37_16(.douta(w_asqrt37_16[0]),.doutb(w_asqrt37_16[1]),.doutc(w_asqrt37_16[2]),.din(w_asqrt37_5[0]));
	jspl3 jspl3_w_asqrt37_17(.douta(w_asqrt37_17[0]),.doutb(w_asqrt37_17[1]),.doutc(w_asqrt37_17[2]),.din(w_asqrt37_5[1]));
	jspl3 jspl3_w_asqrt37_18(.douta(w_asqrt37_18[0]),.doutb(w_asqrt37_18[1]),.doutc(w_asqrt37_18[2]),.din(w_asqrt37_5[2]));
	jspl3 jspl3_w_asqrt37_19(.douta(w_asqrt37_19[0]),.doutb(w_asqrt37_19[1]),.doutc(w_asqrt37_19[2]),.din(w_asqrt37_6[0]));
	jspl3 jspl3_w_asqrt37_20(.douta(w_asqrt37_20[0]),.doutb(w_asqrt37_20[1]),.doutc(w_asqrt37_20[2]),.din(w_asqrt37_6[1]));
	jspl3 jspl3_w_asqrt37_21(.douta(w_asqrt37_21[0]),.doutb(w_asqrt37_21[1]),.doutc(w_asqrt37_21[2]),.din(w_asqrt37_6[2]));
	jspl3 jspl3_w_asqrt37_22(.douta(w_asqrt37_22[0]),.doutb(w_asqrt37_22[1]),.doutc(w_asqrt37_22[2]),.din(w_asqrt37_7[0]));
	jspl3 jspl3_w_asqrt37_23(.douta(w_asqrt37_23[0]),.doutb(w_asqrt37_23[1]),.doutc(asqrt[36]),.din(w_asqrt37_7[1]));
	jspl3 jspl3_w_asqrt38_0(.douta(w_asqrt38_0[0]),.doutb(w_asqrt38_0[1]),.doutc(w_asqrt38_0[2]),.din(asqrt_fa_38));
	jspl3 jspl3_w_asqrt38_1(.douta(w_asqrt38_1[0]),.doutb(w_asqrt38_1[1]),.doutc(w_asqrt38_1[2]),.din(w_asqrt38_0[0]));
	jspl3 jspl3_w_asqrt38_2(.douta(w_asqrt38_2[0]),.doutb(w_asqrt38_2[1]),.doutc(w_asqrt38_2[2]),.din(w_asqrt38_0[1]));
	jspl3 jspl3_w_asqrt38_3(.douta(w_asqrt38_3[0]),.doutb(w_asqrt38_3[1]),.doutc(w_asqrt38_3[2]),.din(w_asqrt38_0[2]));
	jspl3 jspl3_w_asqrt38_4(.douta(w_asqrt38_4[0]),.doutb(w_asqrt38_4[1]),.doutc(w_asqrt38_4[2]),.din(w_asqrt38_1[0]));
	jspl3 jspl3_w_asqrt38_5(.douta(w_asqrt38_5[0]),.doutb(w_asqrt38_5[1]),.doutc(w_asqrt38_5[2]),.din(w_asqrt38_1[1]));
	jspl3 jspl3_w_asqrt38_6(.douta(w_asqrt38_6[0]),.doutb(w_asqrt38_6[1]),.doutc(w_asqrt38_6[2]),.din(w_asqrt38_1[2]));
	jspl3 jspl3_w_asqrt38_7(.douta(w_asqrt38_7[0]),.doutb(w_asqrt38_7[1]),.doutc(w_asqrt38_7[2]),.din(w_asqrt38_2[0]));
	jspl3 jspl3_w_asqrt38_8(.douta(w_asqrt38_8[0]),.doutb(w_asqrt38_8[1]),.doutc(w_asqrt38_8[2]),.din(w_asqrt38_2[1]));
	jspl3 jspl3_w_asqrt38_9(.douta(w_asqrt38_9[0]),.doutb(w_asqrt38_9[1]),.doutc(w_asqrt38_9[2]),.din(w_asqrt38_2[2]));
	jspl3 jspl3_w_asqrt38_10(.douta(w_asqrt38_10[0]),.doutb(w_asqrt38_10[1]),.doutc(w_asqrt38_10[2]),.din(w_asqrt38_3[0]));
	jspl3 jspl3_w_asqrt38_11(.douta(w_asqrt38_11[0]),.doutb(w_asqrt38_11[1]),.doutc(w_asqrt38_11[2]),.din(w_asqrt38_3[1]));
	jspl3 jspl3_w_asqrt38_12(.douta(w_asqrt38_12[0]),.doutb(w_asqrt38_12[1]),.doutc(w_asqrt38_12[2]),.din(w_asqrt38_3[2]));
	jspl3 jspl3_w_asqrt38_13(.douta(w_asqrt38_13[0]),.doutb(w_asqrt38_13[1]),.doutc(w_asqrt38_13[2]),.din(w_asqrt38_4[0]));
	jspl3 jspl3_w_asqrt38_14(.douta(w_asqrt38_14[0]),.doutb(w_asqrt38_14[1]),.doutc(w_asqrt38_14[2]),.din(w_asqrt38_4[1]));
	jspl3 jspl3_w_asqrt38_15(.douta(w_asqrt38_15[0]),.doutb(w_asqrt38_15[1]),.doutc(w_asqrt38_15[2]),.din(w_asqrt38_4[2]));
	jspl3 jspl3_w_asqrt38_16(.douta(w_asqrt38_16[0]),.doutb(w_asqrt38_16[1]),.doutc(w_asqrt38_16[2]),.din(w_asqrt38_5[0]));
	jspl3 jspl3_w_asqrt38_17(.douta(w_asqrt38_17[0]),.doutb(w_asqrt38_17[1]),.doutc(w_asqrt38_17[2]),.din(w_asqrt38_5[1]));
	jspl3 jspl3_w_asqrt38_18(.douta(w_asqrt38_18[0]),.doutb(w_asqrt38_18[1]),.doutc(w_asqrt38_18[2]),.din(w_asqrt38_5[2]));
	jspl3 jspl3_w_asqrt38_19(.douta(w_asqrt38_19[0]),.doutb(w_asqrt38_19[1]),.doutc(w_asqrt38_19[2]),.din(w_asqrt38_6[0]));
	jspl3 jspl3_w_asqrt38_20(.douta(w_asqrt38_20[0]),.doutb(w_asqrt38_20[1]),.doutc(w_asqrt38_20[2]),.din(w_asqrt38_6[1]));
	jspl3 jspl3_w_asqrt38_21(.douta(w_asqrt38_21[0]),.doutb(w_asqrt38_21[1]),.doutc(w_asqrt38_21[2]),.din(w_asqrt38_6[2]));
	jspl3 jspl3_w_asqrt38_22(.douta(w_asqrt38_22[0]),.doutb(w_asqrt38_22[1]),.doutc(w_asqrt38_22[2]),.din(w_asqrt38_7[0]));
	jspl3 jspl3_w_asqrt38_23(.douta(w_asqrt38_23[0]),.doutb(w_asqrt38_23[1]),.doutc(w_asqrt38_23[2]),.din(w_asqrt38_7[1]));
	jspl3 jspl3_w_asqrt38_24(.douta(w_asqrt38_24[0]),.doutb(w_asqrt38_24[1]),.doutc(w_asqrt38_24[2]),.din(w_asqrt38_7[2]));
	jspl3 jspl3_w_asqrt38_25(.douta(w_asqrt38_25[0]),.doutb(w_asqrt38_25[1]),.doutc(w_asqrt38_25[2]),.din(w_asqrt38_8[0]));
	jspl3 jspl3_w_asqrt38_26(.douta(w_asqrt38_26[0]),.doutb(w_asqrt38_26[1]),.doutc(w_asqrt38_26[2]),.din(w_asqrt38_8[1]));
	jspl3 jspl3_w_asqrt38_27(.douta(w_asqrt38_27[0]),.doutb(w_asqrt38_27[1]),.doutc(w_asqrt38_27[2]),.din(w_asqrt38_8[2]));
	jspl3 jspl3_w_asqrt38_28(.douta(w_asqrt38_28[0]),.doutb(w_asqrt38_28[1]),.doutc(w_asqrt38_28[2]),.din(w_asqrt38_9[0]));
	jspl3 jspl3_w_asqrt38_29(.douta(w_asqrt38_29[0]),.doutb(w_asqrt38_29[1]),.doutc(w_asqrt38_29[2]),.din(w_asqrt38_9[1]));
	jspl3 jspl3_w_asqrt38_30(.douta(w_asqrt38_30[0]),.doutb(w_asqrt38_30[1]),.doutc(w_asqrt38_30[2]),.din(w_asqrt38_9[2]));
	jspl jspl_w_asqrt38_31(.douta(w_asqrt38_31),.doutb(asqrt[37]),.din(w_asqrt38_10[0]));
	jspl3 jspl3_w_asqrt39_0(.douta(w_asqrt39_0[0]),.doutb(w_asqrt39_0[1]),.doutc(w_asqrt39_0[2]),.din(asqrt_fa_39));
	jspl3 jspl3_w_asqrt39_1(.douta(w_asqrt39_1[0]),.doutb(w_asqrt39_1[1]),.doutc(w_asqrt39_1[2]),.din(w_asqrt39_0[0]));
	jspl3 jspl3_w_asqrt39_2(.douta(w_asqrt39_2[0]),.doutb(w_asqrt39_2[1]),.doutc(w_asqrt39_2[2]),.din(w_asqrt39_0[1]));
	jspl3 jspl3_w_asqrt39_3(.douta(w_asqrt39_3[0]),.doutb(w_asqrt39_3[1]),.doutc(w_asqrt39_3[2]),.din(w_asqrt39_0[2]));
	jspl3 jspl3_w_asqrt39_4(.douta(w_asqrt39_4[0]),.doutb(w_asqrt39_4[1]),.doutc(w_asqrt39_4[2]),.din(w_asqrt39_1[0]));
	jspl3 jspl3_w_asqrt39_5(.douta(w_asqrt39_5[0]),.doutb(w_asqrt39_5[1]),.doutc(w_asqrt39_5[2]),.din(w_asqrt39_1[1]));
	jspl3 jspl3_w_asqrt39_6(.douta(w_asqrt39_6[0]),.doutb(w_asqrt39_6[1]),.doutc(w_asqrt39_6[2]),.din(w_asqrt39_1[2]));
	jspl3 jspl3_w_asqrt39_7(.douta(w_asqrt39_7[0]),.doutb(w_asqrt39_7[1]),.doutc(w_asqrt39_7[2]),.din(w_asqrt39_2[0]));
	jspl3 jspl3_w_asqrt39_8(.douta(w_asqrt39_8[0]),.doutb(w_asqrt39_8[1]),.doutc(w_asqrt39_8[2]),.din(w_asqrt39_2[1]));
	jspl3 jspl3_w_asqrt39_9(.douta(w_asqrt39_9[0]),.doutb(w_asqrt39_9[1]),.doutc(w_asqrt39_9[2]),.din(w_asqrt39_2[2]));
	jspl3 jspl3_w_asqrt39_10(.douta(w_asqrt39_10[0]),.doutb(w_asqrt39_10[1]),.doutc(w_asqrt39_10[2]),.din(w_asqrt39_3[0]));
	jspl3 jspl3_w_asqrt39_11(.douta(w_asqrt39_11[0]),.doutb(w_asqrt39_11[1]),.doutc(w_asqrt39_11[2]),.din(w_asqrt39_3[1]));
	jspl3 jspl3_w_asqrt39_12(.douta(w_asqrt39_12[0]),.doutb(w_asqrt39_12[1]),.doutc(w_asqrt39_12[2]),.din(w_asqrt39_3[2]));
	jspl3 jspl3_w_asqrt39_13(.douta(w_asqrt39_13[0]),.doutb(w_asqrt39_13[1]),.doutc(w_asqrt39_13[2]),.din(w_asqrt39_4[0]));
	jspl3 jspl3_w_asqrt39_14(.douta(w_asqrt39_14[0]),.doutb(w_asqrt39_14[1]),.doutc(w_asqrt39_14[2]),.din(w_asqrt39_4[1]));
	jspl3 jspl3_w_asqrt39_15(.douta(w_asqrt39_15[0]),.doutb(w_asqrt39_15[1]),.doutc(w_asqrt39_15[2]),.din(w_asqrt39_4[2]));
	jspl3 jspl3_w_asqrt39_16(.douta(w_asqrt39_16[0]),.doutb(w_asqrt39_16[1]),.doutc(w_asqrt39_16[2]),.din(w_asqrt39_5[0]));
	jspl3 jspl3_w_asqrt39_17(.douta(w_asqrt39_17[0]),.doutb(w_asqrt39_17[1]),.doutc(w_asqrt39_17[2]),.din(w_asqrt39_5[1]));
	jspl3 jspl3_w_asqrt39_18(.douta(w_asqrt39_18[0]),.doutb(w_asqrt39_18[1]),.doutc(w_asqrt39_18[2]),.din(w_asqrt39_5[2]));
	jspl3 jspl3_w_asqrt39_19(.douta(w_asqrt39_19[0]),.doutb(w_asqrt39_19[1]),.doutc(w_asqrt39_19[2]),.din(w_asqrt39_6[0]));
	jspl3 jspl3_w_asqrt39_20(.douta(w_asqrt39_20[0]),.doutb(w_asqrt39_20[1]),.doutc(w_asqrt39_20[2]),.din(w_asqrt39_6[1]));
	jspl3 jspl3_w_asqrt39_21(.douta(w_asqrt39_21[0]),.doutb(w_asqrt39_21[1]),.doutc(w_asqrt39_21[2]),.din(w_asqrt39_6[2]));
	jspl3 jspl3_w_asqrt39_22(.douta(w_asqrt39_22[0]),.doutb(w_asqrt39_22[1]),.doutc(w_asqrt39_22[2]),.din(w_asqrt39_7[0]));
	jspl3 jspl3_w_asqrt39_23(.douta(w_asqrt39_23[0]),.doutb(w_asqrt39_23[1]),.doutc(asqrt[38]),.din(w_asqrt39_7[1]));
	jspl3 jspl3_w_asqrt40_0(.douta(w_asqrt40_0[0]),.doutb(w_asqrt40_0[1]),.doutc(w_asqrt40_0[2]),.din(asqrt_fa_40));
	jspl3 jspl3_w_asqrt40_1(.douta(w_asqrt40_1[0]),.doutb(w_asqrt40_1[1]),.doutc(w_asqrt40_1[2]),.din(w_asqrt40_0[0]));
	jspl3 jspl3_w_asqrt40_2(.douta(w_asqrt40_2[0]),.doutb(w_asqrt40_2[1]),.doutc(w_asqrt40_2[2]),.din(w_asqrt40_0[1]));
	jspl3 jspl3_w_asqrt40_3(.douta(w_asqrt40_3[0]),.doutb(w_asqrt40_3[1]),.doutc(w_asqrt40_3[2]),.din(w_asqrt40_0[2]));
	jspl3 jspl3_w_asqrt40_4(.douta(w_asqrt40_4[0]),.doutb(w_asqrt40_4[1]),.doutc(w_asqrt40_4[2]),.din(w_asqrt40_1[0]));
	jspl3 jspl3_w_asqrt40_5(.douta(w_asqrt40_5[0]),.doutb(w_asqrt40_5[1]),.doutc(w_asqrt40_5[2]),.din(w_asqrt40_1[1]));
	jspl3 jspl3_w_asqrt40_6(.douta(w_asqrt40_6[0]),.doutb(w_asqrt40_6[1]),.doutc(w_asqrt40_6[2]),.din(w_asqrt40_1[2]));
	jspl3 jspl3_w_asqrt40_7(.douta(w_asqrt40_7[0]),.doutb(w_asqrt40_7[1]),.doutc(w_asqrt40_7[2]),.din(w_asqrt40_2[0]));
	jspl3 jspl3_w_asqrt40_8(.douta(w_asqrt40_8[0]),.doutb(w_asqrt40_8[1]),.doutc(w_asqrt40_8[2]),.din(w_asqrt40_2[1]));
	jspl3 jspl3_w_asqrt40_9(.douta(w_asqrt40_9[0]),.doutb(w_asqrt40_9[1]),.doutc(w_asqrt40_9[2]),.din(w_asqrt40_2[2]));
	jspl3 jspl3_w_asqrt40_10(.douta(w_asqrt40_10[0]),.doutb(w_asqrt40_10[1]),.doutc(w_asqrt40_10[2]),.din(w_asqrt40_3[0]));
	jspl3 jspl3_w_asqrt40_11(.douta(w_asqrt40_11[0]),.doutb(w_asqrt40_11[1]),.doutc(w_asqrt40_11[2]),.din(w_asqrt40_3[1]));
	jspl3 jspl3_w_asqrt40_12(.douta(w_asqrt40_12[0]),.doutb(w_asqrt40_12[1]),.doutc(w_asqrt40_12[2]),.din(w_asqrt40_3[2]));
	jspl3 jspl3_w_asqrt40_13(.douta(w_asqrt40_13[0]),.doutb(w_asqrt40_13[1]),.doutc(w_asqrt40_13[2]),.din(w_asqrt40_4[0]));
	jspl3 jspl3_w_asqrt40_14(.douta(w_asqrt40_14[0]),.doutb(w_asqrt40_14[1]),.doutc(w_asqrt40_14[2]),.din(w_asqrt40_4[1]));
	jspl3 jspl3_w_asqrt40_15(.douta(w_asqrt40_15[0]),.doutb(w_asqrt40_15[1]),.doutc(w_asqrt40_15[2]),.din(w_asqrt40_4[2]));
	jspl3 jspl3_w_asqrt40_16(.douta(w_asqrt40_16[0]),.doutb(w_asqrt40_16[1]),.doutc(w_asqrt40_16[2]),.din(w_asqrt40_5[0]));
	jspl3 jspl3_w_asqrt40_17(.douta(w_asqrt40_17[0]),.doutb(w_asqrt40_17[1]),.doutc(w_asqrt40_17[2]),.din(w_asqrt40_5[1]));
	jspl3 jspl3_w_asqrt40_18(.douta(w_asqrt40_18[0]),.doutb(w_asqrt40_18[1]),.doutc(w_asqrt40_18[2]),.din(w_asqrt40_5[2]));
	jspl3 jspl3_w_asqrt40_19(.douta(w_asqrt40_19[0]),.doutb(w_asqrt40_19[1]),.doutc(w_asqrt40_19[2]),.din(w_asqrt40_6[0]));
	jspl3 jspl3_w_asqrt40_20(.douta(w_asqrt40_20[0]),.doutb(w_asqrt40_20[1]),.doutc(w_asqrt40_20[2]),.din(w_asqrt40_6[1]));
	jspl3 jspl3_w_asqrt40_21(.douta(w_asqrt40_21[0]),.doutb(w_asqrt40_21[1]),.doutc(w_asqrt40_21[2]),.din(w_asqrt40_6[2]));
	jspl3 jspl3_w_asqrt40_22(.douta(w_asqrt40_22[0]),.doutb(w_asqrt40_22[1]),.doutc(w_asqrt40_22[2]),.din(w_asqrt40_7[0]));
	jspl3 jspl3_w_asqrt40_23(.douta(w_asqrt40_23[0]),.doutb(w_asqrt40_23[1]),.doutc(w_asqrt40_23[2]),.din(w_asqrt40_7[1]));
	jspl3 jspl3_w_asqrt40_24(.douta(w_asqrt40_24[0]),.doutb(w_asqrt40_24[1]),.doutc(w_asqrt40_24[2]),.din(w_asqrt40_7[2]));
	jspl3 jspl3_w_asqrt40_25(.douta(w_asqrt40_25[0]),.doutb(w_asqrt40_25[1]),.doutc(w_asqrt40_25[2]),.din(w_asqrt40_8[0]));
	jspl3 jspl3_w_asqrt40_26(.douta(w_asqrt40_26[0]),.doutb(w_asqrt40_26[1]),.doutc(w_asqrt40_26[2]),.din(w_asqrt40_8[1]));
	jspl3 jspl3_w_asqrt40_27(.douta(w_asqrt40_27[0]),.doutb(w_asqrt40_27[1]),.doutc(w_asqrt40_27[2]),.din(w_asqrt40_8[2]));
	jspl3 jspl3_w_asqrt40_28(.douta(w_asqrt40_28[0]),.doutb(w_asqrt40_28[1]),.doutc(w_asqrt40_28[2]),.din(w_asqrt40_9[0]));
	jspl3 jspl3_w_asqrt40_29(.douta(w_asqrt40_29[0]),.doutb(w_asqrt40_29[1]),.doutc(w_asqrt40_29[2]),.din(w_asqrt40_9[1]));
	jspl3 jspl3_w_asqrt40_30(.douta(w_asqrt40_30[0]),.doutb(w_asqrt40_30[1]),.doutc(w_asqrt40_30[2]),.din(w_asqrt40_9[2]));
	jspl jspl_w_asqrt40_31(.douta(w_asqrt40_31),.doutb(asqrt[39]),.din(w_asqrt40_10[0]));
	jspl3 jspl3_w_asqrt41_0(.douta(w_asqrt41_0[0]),.doutb(w_asqrt41_0[1]),.doutc(w_asqrt41_0[2]),.din(asqrt_fa_41));
	jspl3 jspl3_w_asqrt41_1(.douta(w_asqrt41_1[0]),.doutb(w_asqrt41_1[1]),.doutc(w_asqrt41_1[2]),.din(w_asqrt41_0[0]));
	jspl3 jspl3_w_asqrt41_2(.douta(w_asqrt41_2[0]),.doutb(w_asqrt41_2[1]),.doutc(w_asqrt41_2[2]),.din(w_asqrt41_0[1]));
	jspl3 jspl3_w_asqrt41_3(.douta(w_asqrt41_3[0]),.doutb(w_asqrt41_3[1]),.doutc(w_asqrt41_3[2]),.din(w_asqrt41_0[2]));
	jspl3 jspl3_w_asqrt41_4(.douta(w_asqrt41_4[0]),.doutb(w_asqrt41_4[1]),.doutc(w_asqrt41_4[2]),.din(w_asqrt41_1[0]));
	jspl3 jspl3_w_asqrt41_5(.douta(w_asqrt41_5[0]),.doutb(w_asqrt41_5[1]),.doutc(w_asqrt41_5[2]),.din(w_asqrt41_1[1]));
	jspl3 jspl3_w_asqrt41_6(.douta(w_asqrt41_6[0]),.doutb(w_asqrt41_6[1]),.doutc(w_asqrt41_6[2]),.din(w_asqrt41_1[2]));
	jspl3 jspl3_w_asqrt41_7(.douta(w_asqrt41_7[0]),.doutb(w_asqrt41_7[1]),.doutc(w_asqrt41_7[2]),.din(w_asqrt41_2[0]));
	jspl3 jspl3_w_asqrt41_8(.douta(w_asqrt41_8[0]),.doutb(w_asqrt41_8[1]),.doutc(w_asqrt41_8[2]),.din(w_asqrt41_2[1]));
	jspl3 jspl3_w_asqrt41_9(.douta(w_asqrt41_9[0]),.doutb(w_asqrt41_9[1]),.doutc(w_asqrt41_9[2]),.din(w_asqrt41_2[2]));
	jspl3 jspl3_w_asqrt41_10(.douta(w_asqrt41_10[0]),.doutb(w_asqrt41_10[1]),.doutc(w_asqrt41_10[2]),.din(w_asqrt41_3[0]));
	jspl3 jspl3_w_asqrt41_11(.douta(w_asqrt41_11[0]),.doutb(w_asqrt41_11[1]),.doutc(w_asqrt41_11[2]),.din(w_asqrt41_3[1]));
	jspl3 jspl3_w_asqrt41_12(.douta(w_asqrt41_12[0]),.doutb(w_asqrt41_12[1]),.doutc(w_asqrt41_12[2]),.din(w_asqrt41_3[2]));
	jspl3 jspl3_w_asqrt41_13(.douta(w_asqrt41_13[0]),.doutb(w_asqrt41_13[1]),.doutc(w_asqrt41_13[2]),.din(w_asqrt41_4[0]));
	jspl3 jspl3_w_asqrt41_14(.douta(w_asqrt41_14[0]),.doutb(w_asqrt41_14[1]),.doutc(w_asqrt41_14[2]),.din(w_asqrt41_4[1]));
	jspl3 jspl3_w_asqrt41_15(.douta(w_asqrt41_15[0]),.doutb(w_asqrt41_15[1]),.doutc(w_asqrt41_15[2]),.din(w_asqrt41_4[2]));
	jspl3 jspl3_w_asqrt41_16(.douta(w_asqrt41_16[0]),.doutb(w_asqrt41_16[1]),.doutc(w_asqrt41_16[2]),.din(w_asqrt41_5[0]));
	jspl3 jspl3_w_asqrt41_17(.douta(w_asqrt41_17[0]),.doutb(w_asqrt41_17[1]),.doutc(w_asqrt41_17[2]),.din(w_asqrt41_5[1]));
	jspl3 jspl3_w_asqrt41_18(.douta(w_asqrt41_18[0]),.doutb(w_asqrt41_18[1]),.doutc(w_asqrt41_18[2]),.din(w_asqrt41_5[2]));
	jspl3 jspl3_w_asqrt41_19(.douta(w_asqrt41_19[0]),.doutb(w_asqrt41_19[1]),.doutc(w_asqrt41_19[2]),.din(w_asqrt41_6[0]));
	jspl3 jspl3_w_asqrt41_20(.douta(w_asqrt41_20[0]),.doutb(w_asqrt41_20[1]),.doutc(w_asqrt41_20[2]),.din(w_asqrt41_6[1]));
	jspl3 jspl3_w_asqrt41_21(.douta(w_asqrt41_21[0]),.doutb(w_asqrt41_21[1]),.doutc(w_asqrt41_21[2]),.din(w_asqrt41_6[2]));
	jspl3 jspl3_w_asqrt41_22(.douta(w_asqrt41_22[0]),.doutb(w_asqrt41_22[1]),.doutc(w_asqrt41_22[2]),.din(w_asqrt41_7[0]));
	jspl3 jspl3_w_asqrt41_23(.douta(w_asqrt41_23[0]),.doutb(w_asqrt41_23[1]),.doutc(w_asqrt41_23[2]),.din(w_asqrt41_7[1]));
	jspl3 jspl3_w_asqrt41_24(.douta(w_asqrt41_24[0]),.doutb(w_asqrt41_24[1]),.doutc(asqrt[40]),.din(w_asqrt41_7[2]));
	jspl3 jspl3_w_asqrt42_0(.douta(w_asqrt42_0[0]),.doutb(w_asqrt42_0[1]),.doutc(w_asqrt42_0[2]),.din(asqrt_fa_42));
	jspl3 jspl3_w_asqrt42_1(.douta(w_asqrt42_1[0]),.doutb(w_asqrt42_1[1]),.doutc(w_asqrt42_1[2]),.din(w_asqrt42_0[0]));
	jspl3 jspl3_w_asqrt42_2(.douta(w_asqrt42_2[0]),.doutb(w_asqrt42_2[1]),.doutc(w_asqrt42_2[2]),.din(w_asqrt42_0[1]));
	jspl3 jspl3_w_asqrt42_3(.douta(w_asqrt42_3[0]),.doutb(w_asqrt42_3[1]),.doutc(w_asqrt42_3[2]),.din(w_asqrt42_0[2]));
	jspl3 jspl3_w_asqrt42_4(.douta(w_asqrt42_4[0]),.doutb(w_asqrt42_4[1]),.doutc(w_asqrt42_4[2]),.din(w_asqrt42_1[0]));
	jspl3 jspl3_w_asqrt42_5(.douta(w_asqrt42_5[0]),.doutb(w_asqrt42_5[1]),.doutc(w_asqrt42_5[2]),.din(w_asqrt42_1[1]));
	jspl3 jspl3_w_asqrt42_6(.douta(w_asqrt42_6[0]),.doutb(w_asqrt42_6[1]),.doutc(w_asqrt42_6[2]),.din(w_asqrt42_1[2]));
	jspl3 jspl3_w_asqrt42_7(.douta(w_asqrt42_7[0]),.doutb(w_asqrt42_7[1]),.doutc(w_asqrt42_7[2]),.din(w_asqrt42_2[0]));
	jspl3 jspl3_w_asqrt42_8(.douta(w_asqrt42_8[0]),.doutb(w_asqrt42_8[1]),.doutc(w_asqrt42_8[2]),.din(w_asqrt42_2[1]));
	jspl3 jspl3_w_asqrt42_9(.douta(w_asqrt42_9[0]),.doutb(w_asqrt42_9[1]),.doutc(w_asqrt42_9[2]),.din(w_asqrt42_2[2]));
	jspl3 jspl3_w_asqrt42_10(.douta(w_asqrt42_10[0]),.doutb(w_asqrt42_10[1]),.doutc(w_asqrt42_10[2]),.din(w_asqrt42_3[0]));
	jspl3 jspl3_w_asqrt42_11(.douta(w_asqrt42_11[0]),.doutb(w_asqrt42_11[1]),.doutc(w_asqrt42_11[2]),.din(w_asqrt42_3[1]));
	jspl3 jspl3_w_asqrt42_12(.douta(w_asqrt42_12[0]),.doutb(w_asqrt42_12[1]),.doutc(w_asqrt42_12[2]),.din(w_asqrt42_3[2]));
	jspl3 jspl3_w_asqrt42_13(.douta(w_asqrt42_13[0]),.doutb(w_asqrt42_13[1]),.doutc(w_asqrt42_13[2]),.din(w_asqrt42_4[0]));
	jspl3 jspl3_w_asqrt42_14(.douta(w_asqrt42_14[0]),.doutb(w_asqrt42_14[1]),.doutc(w_asqrt42_14[2]),.din(w_asqrt42_4[1]));
	jspl3 jspl3_w_asqrt42_15(.douta(w_asqrt42_15[0]),.doutb(w_asqrt42_15[1]),.doutc(w_asqrt42_15[2]),.din(w_asqrt42_4[2]));
	jspl3 jspl3_w_asqrt42_16(.douta(w_asqrt42_16[0]),.doutb(w_asqrt42_16[1]),.doutc(w_asqrt42_16[2]),.din(w_asqrt42_5[0]));
	jspl3 jspl3_w_asqrt42_17(.douta(w_asqrt42_17[0]),.doutb(w_asqrt42_17[1]),.doutc(w_asqrt42_17[2]),.din(w_asqrt42_5[1]));
	jspl3 jspl3_w_asqrt42_18(.douta(w_asqrt42_18[0]),.doutb(w_asqrt42_18[1]),.doutc(w_asqrt42_18[2]),.din(w_asqrt42_5[2]));
	jspl3 jspl3_w_asqrt42_19(.douta(w_asqrt42_19[0]),.doutb(w_asqrt42_19[1]),.doutc(w_asqrt42_19[2]),.din(w_asqrt42_6[0]));
	jspl3 jspl3_w_asqrt42_20(.douta(w_asqrt42_20[0]),.doutb(w_asqrt42_20[1]),.doutc(w_asqrt42_20[2]),.din(w_asqrt42_6[1]));
	jspl3 jspl3_w_asqrt42_21(.douta(w_asqrt42_21[0]),.doutb(w_asqrt42_21[1]),.doutc(w_asqrt42_21[2]),.din(w_asqrt42_6[2]));
	jspl3 jspl3_w_asqrt42_22(.douta(w_asqrt42_22[0]),.doutb(w_asqrt42_22[1]),.doutc(w_asqrt42_22[2]),.din(w_asqrt42_7[0]));
	jspl3 jspl3_w_asqrt42_23(.douta(w_asqrt42_23[0]),.doutb(w_asqrt42_23[1]),.doutc(w_asqrt42_23[2]),.din(w_asqrt42_7[1]));
	jspl3 jspl3_w_asqrt42_24(.douta(w_asqrt42_24[0]),.doutb(w_asqrt42_24[1]),.doutc(w_asqrt42_24[2]),.din(w_asqrt42_7[2]));
	jspl3 jspl3_w_asqrt42_25(.douta(w_asqrt42_25[0]),.doutb(w_asqrt42_25[1]),.doutc(w_asqrt42_25[2]),.din(w_asqrt42_8[0]));
	jspl3 jspl3_w_asqrt42_26(.douta(w_asqrt42_26[0]),.doutb(w_asqrt42_26[1]),.doutc(w_asqrt42_26[2]),.din(w_asqrt42_8[1]));
	jspl3 jspl3_w_asqrt42_27(.douta(w_asqrt42_27[0]),.doutb(w_asqrt42_27[1]),.doutc(w_asqrt42_27[2]),.din(w_asqrt42_8[2]));
	jspl3 jspl3_w_asqrt42_28(.douta(w_asqrt42_28[0]),.doutb(w_asqrt42_28[1]),.doutc(w_asqrt42_28[2]),.din(w_asqrt42_9[0]));
	jspl3 jspl3_w_asqrt42_29(.douta(w_asqrt42_29[0]),.doutb(w_asqrt42_29[1]),.doutc(w_asqrt42_29[2]),.din(w_asqrt42_9[1]));
	jspl3 jspl3_w_asqrt42_30(.douta(w_asqrt42_30[0]),.doutb(w_asqrt42_30[1]),.doutc(w_asqrt42_30[2]),.din(w_asqrt42_9[2]));
	jspl jspl_w_asqrt42_31(.douta(w_asqrt42_31),.doutb(asqrt[41]),.din(w_asqrt42_10[0]));
	jspl3 jspl3_w_asqrt43_0(.douta(w_asqrt43_0[0]),.doutb(w_asqrt43_0[1]),.doutc(w_asqrt43_0[2]),.din(asqrt_fa_43));
	jspl3 jspl3_w_asqrt43_1(.douta(w_asqrt43_1[0]),.doutb(w_asqrt43_1[1]),.doutc(w_asqrt43_1[2]),.din(w_asqrt43_0[0]));
	jspl3 jspl3_w_asqrt43_2(.douta(w_asqrt43_2[0]),.doutb(w_asqrt43_2[1]),.doutc(w_asqrt43_2[2]),.din(w_asqrt43_0[1]));
	jspl3 jspl3_w_asqrt43_3(.douta(w_asqrt43_3[0]),.doutb(w_asqrt43_3[1]),.doutc(w_asqrt43_3[2]),.din(w_asqrt43_0[2]));
	jspl3 jspl3_w_asqrt43_4(.douta(w_asqrt43_4[0]),.doutb(w_asqrt43_4[1]),.doutc(w_asqrt43_4[2]),.din(w_asqrt43_1[0]));
	jspl3 jspl3_w_asqrt43_5(.douta(w_asqrt43_5[0]),.doutb(w_asqrt43_5[1]),.doutc(w_asqrt43_5[2]),.din(w_asqrt43_1[1]));
	jspl3 jspl3_w_asqrt43_6(.douta(w_asqrt43_6[0]),.doutb(w_asqrt43_6[1]),.doutc(w_asqrt43_6[2]),.din(w_asqrt43_1[2]));
	jspl3 jspl3_w_asqrt43_7(.douta(w_asqrt43_7[0]),.doutb(w_asqrt43_7[1]),.doutc(w_asqrt43_7[2]),.din(w_asqrt43_2[0]));
	jspl3 jspl3_w_asqrt43_8(.douta(w_asqrt43_8[0]),.doutb(w_asqrt43_8[1]),.doutc(w_asqrt43_8[2]),.din(w_asqrt43_2[1]));
	jspl3 jspl3_w_asqrt43_9(.douta(w_asqrt43_9[0]),.doutb(w_asqrt43_9[1]),.doutc(w_asqrt43_9[2]),.din(w_asqrt43_2[2]));
	jspl3 jspl3_w_asqrt43_10(.douta(w_asqrt43_10[0]),.doutb(w_asqrt43_10[1]),.doutc(w_asqrt43_10[2]),.din(w_asqrt43_3[0]));
	jspl3 jspl3_w_asqrt43_11(.douta(w_asqrt43_11[0]),.doutb(w_asqrt43_11[1]),.doutc(w_asqrt43_11[2]),.din(w_asqrt43_3[1]));
	jspl3 jspl3_w_asqrt43_12(.douta(w_asqrt43_12[0]),.doutb(w_asqrt43_12[1]),.doutc(w_asqrt43_12[2]),.din(w_asqrt43_3[2]));
	jspl3 jspl3_w_asqrt43_13(.douta(w_asqrt43_13[0]),.doutb(w_asqrt43_13[1]),.doutc(w_asqrt43_13[2]),.din(w_asqrt43_4[0]));
	jspl3 jspl3_w_asqrt43_14(.douta(w_asqrt43_14[0]),.doutb(w_asqrt43_14[1]),.doutc(w_asqrt43_14[2]),.din(w_asqrt43_4[1]));
	jspl3 jspl3_w_asqrt43_15(.douta(w_asqrt43_15[0]),.doutb(w_asqrt43_15[1]),.doutc(w_asqrt43_15[2]),.din(w_asqrt43_4[2]));
	jspl3 jspl3_w_asqrt43_16(.douta(w_asqrt43_16[0]),.doutb(w_asqrt43_16[1]),.doutc(w_asqrt43_16[2]),.din(w_asqrt43_5[0]));
	jspl3 jspl3_w_asqrt43_17(.douta(w_asqrt43_17[0]),.doutb(w_asqrt43_17[1]),.doutc(w_asqrt43_17[2]),.din(w_asqrt43_5[1]));
	jspl3 jspl3_w_asqrt43_18(.douta(w_asqrt43_18[0]),.doutb(w_asqrt43_18[1]),.doutc(w_asqrt43_18[2]),.din(w_asqrt43_5[2]));
	jspl3 jspl3_w_asqrt43_19(.douta(w_asqrt43_19[0]),.doutb(w_asqrt43_19[1]),.doutc(w_asqrt43_19[2]),.din(w_asqrt43_6[0]));
	jspl3 jspl3_w_asqrt43_20(.douta(w_asqrt43_20[0]),.doutb(w_asqrt43_20[1]),.doutc(w_asqrt43_20[2]),.din(w_asqrt43_6[1]));
	jspl3 jspl3_w_asqrt43_21(.douta(w_asqrt43_21[0]),.doutb(w_asqrt43_21[1]),.doutc(w_asqrt43_21[2]),.din(w_asqrt43_6[2]));
	jspl3 jspl3_w_asqrt43_22(.douta(w_asqrt43_22[0]),.doutb(w_asqrt43_22[1]),.doutc(w_asqrt43_22[2]),.din(w_asqrt43_7[0]));
	jspl3 jspl3_w_asqrt43_23(.douta(w_asqrt43_23[0]),.doutb(w_asqrt43_23[1]),.doutc(w_asqrt43_23[2]),.din(w_asqrt43_7[1]));
	jspl3 jspl3_w_asqrt43_24(.douta(w_asqrt43_24[0]),.doutb(w_asqrt43_24[1]),.doutc(asqrt[42]),.din(w_asqrt43_7[2]));
	jspl3 jspl3_w_asqrt44_0(.douta(w_asqrt44_0[0]),.doutb(w_asqrt44_0[1]),.doutc(w_asqrt44_0[2]),.din(asqrt_fa_44));
	jspl3 jspl3_w_asqrt44_1(.douta(w_asqrt44_1[0]),.doutb(w_asqrt44_1[1]),.doutc(w_asqrt44_1[2]),.din(w_asqrt44_0[0]));
	jspl3 jspl3_w_asqrt44_2(.douta(w_asqrt44_2[0]),.doutb(w_asqrt44_2[1]),.doutc(w_asqrt44_2[2]),.din(w_asqrt44_0[1]));
	jspl3 jspl3_w_asqrt44_3(.douta(w_asqrt44_3[0]),.doutb(w_asqrt44_3[1]),.doutc(w_asqrt44_3[2]),.din(w_asqrt44_0[2]));
	jspl3 jspl3_w_asqrt44_4(.douta(w_asqrt44_4[0]),.doutb(w_asqrt44_4[1]),.doutc(w_asqrt44_4[2]),.din(w_asqrt44_1[0]));
	jspl3 jspl3_w_asqrt44_5(.douta(w_asqrt44_5[0]),.doutb(w_asqrt44_5[1]),.doutc(w_asqrt44_5[2]),.din(w_asqrt44_1[1]));
	jspl3 jspl3_w_asqrt44_6(.douta(w_asqrt44_6[0]),.doutb(w_asqrt44_6[1]),.doutc(w_asqrt44_6[2]),.din(w_asqrt44_1[2]));
	jspl3 jspl3_w_asqrt44_7(.douta(w_asqrt44_7[0]),.doutb(w_asqrt44_7[1]),.doutc(w_asqrt44_7[2]),.din(w_asqrt44_2[0]));
	jspl3 jspl3_w_asqrt44_8(.douta(w_asqrt44_8[0]),.doutb(w_asqrt44_8[1]),.doutc(w_asqrt44_8[2]),.din(w_asqrt44_2[1]));
	jspl3 jspl3_w_asqrt44_9(.douta(w_asqrt44_9[0]),.doutb(w_asqrt44_9[1]),.doutc(w_asqrt44_9[2]),.din(w_asqrt44_2[2]));
	jspl3 jspl3_w_asqrt44_10(.douta(w_asqrt44_10[0]),.doutb(w_asqrt44_10[1]),.doutc(w_asqrt44_10[2]),.din(w_asqrt44_3[0]));
	jspl3 jspl3_w_asqrt44_11(.douta(w_asqrt44_11[0]),.doutb(w_asqrt44_11[1]),.doutc(w_asqrt44_11[2]),.din(w_asqrt44_3[1]));
	jspl3 jspl3_w_asqrt44_12(.douta(w_asqrt44_12[0]),.doutb(w_asqrt44_12[1]),.doutc(w_asqrt44_12[2]),.din(w_asqrt44_3[2]));
	jspl3 jspl3_w_asqrt44_13(.douta(w_asqrt44_13[0]),.doutb(w_asqrt44_13[1]),.doutc(w_asqrt44_13[2]),.din(w_asqrt44_4[0]));
	jspl3 jspl3_w_asqrt44_14(.douta(w_asqrt44_14[0]),.doutb(w_asqrt44_14[1]),.doutc(w_asqrt44_14[2]),.din(w_asqrt44_4[1]));
	jspl3 jspl3_w_asqrt44_15(.douta(w_asqrt44_15[0]),.doutb(w_asqrt44_15[1]),.doutc(w_asqrt44_15[2]),.din(w_asqrt44_4[2]));
	jspl3 jspl3_w_asqrt44_16(.douta(w_asqrt44_16[0]),.doutb(w_asqrt44_16[1]),.doutc(w_asqrt44_16[2]),.din(w_asqrt44_5[0]));
	jspl3 jspl3_w_asqrt44_17(.douta(w_asqrt44_17[0]),.doutb(w_asqrt44_17[1]),.doutc(w_asqrt44_17[2]),.din(w_asqrt44_5[1]));
	jspl3 jspl3_w_asqrt44_18(.douta(w_asqrt44_18[0]),.doutb(w_asqrt44_18[1]),.doutc(w_asqrt44_18[2]),.din(w_asqrt44_5[2]));
	jspl3 jspl3_w_asqrt44_19(.douta(w_asqrt44_19[0]),.doutb(w_asqrt44_19[1]),.doutc(w_asqrt44_19[2]),.din(w_asqrt44_6[0]));
	jspl3 jspl3_w_asqrt44_20(.douta(w_asqrt44_20[0]),.doutb(w_asqrt44_20[1]),.doutc(w_asqrt44_20[2]),.din(w_asqrt44_6[1]));
	jspl3 jspl3_w_asqrt44_21(.douta(w_asqrt44_21[0]),.doutb(w_asqrt44_21[1]),.doutc(w_asqrt44_21[2]),.din(w_asqrt44_6[2]));
	jspl3 jspl3_w_asqrt44_22(.douta(w_asqrt44_22[0]),.doutb(w_asqrt44_22[1]),.doutc(w_asqrt44_22[2]),.din(w_asqrt44_7[0]));
	jspl3 jspl3_w_asqrt44_23(.douta(w_asqrt44_23[0]),.doutb(w_asqrt44_23[1]),.doutc(w_asqrt44_23[2]),.din(w_asqrt44_7[1]));
	jspl3 jspl3_w_asqrt44_24(.douta(w_asqrt44_24[0]),.doutb(w_asqrt44_24[1]),.doutc(w_asqrt44_24[2]),.din(w_asqrt44_7[2]));
	jspl3 jspl3_w_asqrt44_25(.douta(w_asqrt44_25[0]),.doutb(w_asqrt44_25[1]),.doutc(w_asqrt44_25[2]),.din(w_asqrt44_8[0]));
	jspl3 jspl3_w_asqrt44_26(.douta(w_asqrt44_26[0]),.doutb(w_asqrt44_26[1]),.doutc(w_asqrt44_26[2]),.din(w_asqrt44_8[1]));
	jspl3 jspl3_w_asqrt44_27(.douta(w_asqrt44_27[0]),.doutb(w_asqrt44_27[1]),.doutc(w_asqrt44_27[2]),.din(w_asqrt44_8[2]));
	jspl3 jspl3_w_asqrt44_28(.douta(w_asqrt44_28[0]),.doutb(w_asqrt44_28[1]),.doutc(w_asqrt44_28[2]),.din(w_asqrt44_9[0]));
	jspl3 jspl3_w_asqrt44_29(.douta(w_asqrt44_29[0]),.doutb(w_asqrt44_29[1]),.doutc(w_asqrt44_29[2]),.din(w_asqrt44_9[1]));
	jspl3 jspl3_w_asqrt44_30(.douta(w_asqrt44_30[0]),.doutb(w_asqrt44_30[1]),.doutc(w_asqrt44_30[2]),.din(w_asqrt44_9[2]));
	jspl jspl_w_asqrt44_31(.douta(w_asqrt44_31),.doutb(asqrt[43]),.din(w_asqrt44_10[0]));
	jspl3 jspl3_w_asqrt45_0(.douta(w_asqrt45_0[0]),.doutb(w_asqrt45_0[1]),.doutc(w_asqrt45_0[2]),.din(asqrt_fa_45));
	jspl3 jspl3_w_asqrt45_1(.douta(w_asqrt45_1[0]),.doutb(w_asqrt45_1[1]),.doutc(w_asqrt45_1[2]),.din(w_asqrt45_0[0]));
	jspl3 jspl3_w_asqrt45_2(.douta(w_asqrt45_2[0]),.doutb(w_asqrt45_2[1]),.doutc(w_asqrt45_2[2]),.din(w_asqrt45_0[1]));
	jspl3 jspl3_w_asqrt45_3(.douta(w_asqrt45_3[0]),.doutb(w_asqrt45_3[1]),.doutc(w_asqrt45_3[2]),.din(w_asqrt45_0[2]));
	jspl3 jspl3_w_asqrt45_4(.douta(w_asqrt45_4[0]),.doutb(w_asqrt45_4[1]),.doutc(w_asqrt45_4[2]),.din(w_asqrt45_1[0]));
	jspl3 jspl3_w_asqrt45_5(.douta(w_asqrt45_5[0]),.doutb(w_asqrt45_5[1]),.doutc(w_asqrt45_5[2]),.din(w_asqrt45_1[1]));
	jspl3 jspl3_w_asqrt45_6(.douta(w_asqrt45_6[0]),.doutb(w_asqrt45_6[1]),.doutc(w_asqrt45_6[2]),.din(w_asqrt45_1[2]));
	jspl3 jspl3_w_asqrt45_7(.douta(w_asqrt45_7[0]),.doutb(w_asqrt45_7[1]),.doutc(w_asqrt45_7[2]),.din(w_asqrt45_2[0]));
	jspl3 jspl3_w_asqrt45_8(.douta(w_asqrt45_8[0]),.doutb(w_asqrt45_8[1]),.doutc(w_asqrt45_8[2]),.din(w_asqrt45_2[1]));
	jspl3 jspl3_w_asqrt45_9(.douta(w_asqrt45_9[0]),.doutb(w_asqrt45_9[1]),.doutc(w_asqrt45_9[2]),.din(w_asqrt45_2[2]));
	jspl3 jspl3_w_asqrt45_10(.douta(w_asqrt45_10[0]),.doutb(w_asqrt45_10[1]),.doutc(w_asqrt45_10[2]),.din(w_asqrt45_3[0]));
	jspl3 jspl3_w_asqrt45_11(.douta(w_asqrt45_11[0]),.doutb(w_asqrt45_11[1]),.doutc(w_asqrt45_11[2]),.din(w_asqrt45_3[1]));
	jspl3 jspl3_w_asqrt45_12(.douta(w_asqrt45_12[0]),.doutb(w_asqrt45_12[1]),.doutc(w_asqrt45_12[2]),.din(w_asqrt45_3[2]));
	jspl3 jspl3_w_asqrt45_13(.douta(w_asqrt45_13[0]),.doutb(w_asqrt45_13[1]),.doutc(w_asqrt45_13[2]),.din(w_asqrt45_4[0]));
	jspl3 jspl3_w_asqrt45_14(.douta(w_asqrt45_14[0]),.doutb(w_asqrt45_14[1]),.doutc(w_asqrt45_14[2]),.din(w_asqrt45_4[1]));
	jspl3 jspl3_w_asqrt45_15(.douta(w_asqrt45_15[0]),.doutb(w_asqrt45_15[1]),.doutc(w_asqrt45_15[2]),.din(w_asqrt45_4[2]));
	jspl3 jspl3_w_asqrt45_16(.douta(w_asqrt45_16[0]),.doutb(w_asqrt45_16[1]),.doutc(w_asqrt45_16[2]),.din(w_asqrt45_5[0]));
	jspl3 jspl3_w_asqrt45_17(.douta(w_asqrt45_17[0]),.doutb(w_asqrt45_17[1]),.doutc(w_asqrt45_17[2]),.din(w_asqrt45_5[1]));
	jspl3 jspl3_w_asqrt45_18(.douta(w_asqrt45_18[0]),.doutb(w_asqrt45_18[1]),.doutc(w_asqrt45_18[2]),.din(w_asqrt45_5[2]));
	jspl3 jspl3_w_asqrt45_19(.douta(w_asqrt45_19[0]),.doutb(w_asqrt45_19[1]),.doutc(w_asqrt45_19[2]),.din(w_asqrt45_6[0]));
	jspl3 jspl3_w_asqrt45_20(.douta(w_asqrt45_20[0]),.doutb(w_asqrt45_20[1]),.doutc(w_asqrt45_20[2]),.din(w_asqrt45_6[1]));
	jspl3 jspl3_w_asqrt45_21(.douta(w_asqrt45_21[0]),.doutb(w_asqrt45_21[1]),.doutc(w_asqrt45_21[2]),.din(w_asqrt45_6[2]));
	jspl3 jspl3_w_asqrt45_22(.douta(w_asqrt45_22[0]),.doutb(w_asqrt45_22[1]),.doutc(w_asqrt45_22[2]),.din(w_asqrt45_7[0]));
	jspl3 jspl3_w_asqrt45_23(.douta(w_asqrt45_23[0]),.doutb(w_asqrt45_23[1]),.doutc(w_asqrt45_23[2]),.din(w_asqrt45_7[1]));
	jspl3 jspl3_w_asqrt45_24(.douta(w_asqrt45_24[0]),.doutb(w_asqrt45_24[1]),.doutc(w_asqrt45_24[2]),.din(w_asqrt45_7[2]));
	jspl3 jspl3_w_asqrt45_25(.douta(w_asqrt45_25[0]),.doutb(w_asqrt45_25[1]),.doutc(asqrt[44]),.din(w_asqrt45_8[0]));
	jspl3 jspl3_w_asqrt46_0(.douta(w_asqrt46_0[0]),.doutb(w_asqrt46_0[1]),.doutc(w_asqrt46_0[2]),.din(asqrt_fa_46));
	jspl3 jspl3_w_asqrt46_1(.douta(w_asqrt46_1[0]),.doutb(w_asqrt46_1[1]),.doutc(w_asqrt46_1[2]),.din(w_asqrt46_0[0]));
	jspl3 jspl3_w_asqrt46_2(.douta(w_asqrt46_2[0]),.doutb(w_asqrt46_2[1]),.doutc(w_asqrt46_2[2]),.din(w_asqrt46_0[1]));
	jspl3 jspl3_w_asqrt46_3(.douta(w_asqrt46_3[0]),.doutb(w_asqrt46_3[1]),.doutc(w_asqrt46_3[2]),.din(w_asqrt46_0[2]));
	jspl3 jspl3_w_asqrt46_4(.douta(w_asqrt46_4[0]),.doutb(w_asqrt46_4[1]),.doutc(w_asqrt46_4[2]),.din(w_asqrt46_1[0]));
	jspl3 jspl3_w_asqrt46_5(.douta(w_asqrt46_5[0]),.doutb(w_asqrt46_5[1]),.doutc(w_asqrt46_5[2]),.din(w_asqrt46_1[1]));
	jspl3 jspl3_w_asqrt46_6(.douta(w_asqrt46_6[0]),.doutb(w_asqrt46_6[1]),.doutc(w_asqrt46_6[2]),.din(w_asqrt46_1[2]));
	jspl3 jspl3_w_asqrt46_7(.douta(w_asqrt46_7[0]),.doutb(w_asqrt46_7[1]),.doutc(w_asqrt46_7[2]),.din(w_asqrt46_2[0]));
	jspl3 jspl3_w_asqrt46_8(.douta(w_asqrt46_8[0]),.doutb(w_asqrt46_8[1]),.doutc(w_asqrt46_8[2]),.din(w_asqrt46_2[1]));
	jspl3 jspl3_w_asqrt46_9(.douta(w_asqrt46_9[0]),.doutb(w_asqrt46_9[1]),.doutc(w_asqrt46_9[2]),.din(w_asqrt46_2[2]));
	jspl3 jspl3_w_asqrt46_10(.douta(w_asqrt46_10[0]),.doutb(w_asqrt46_10[1]),.doutc(w_asqrt46_10[2]),.din(w_asqrt46_3[0]));
	jspl3 jspl3_w_asqrt46_11(.douta(w_asqrt46_11[0]),.doutb(w_asqrt46_11[1]),.doutc(w_asqrt46_11[2]),.din(w_asqrt46_3[1]));
	jspl3 jspl3_w_asqrt46_12(.douta(w_asqrt46_12[0]),.doutb(w_asqrt46_12[1]),.doutc(w_asqrt46_12[2]),.din(w_asqrt46_3[2]));
	jspl3 jspl3_w_asqrt46_13(.douta(w_asqrt46_13[0]),.doutb(w_asqrt46_13[1]),.doutc(w_asqrt46_13[2]),.din(w_asqrt46_4[0]));
	jspl3 jspl3_w_asqrt46_14(.douta(w_asqrt46_14[0]),.doutb(w_asqrt46_14[1]),.doutc(w_asqrt46_14[2]),.din(w_asqrt46_4[1]));
	jspl3 jspl3_w_asqrt46_15(.douta(w_asqrt46_15[0]),.doutb(w_asqrt46_15[1]),.doutc(w_asqrt46_15[2]),.din(w_asqrt46_4[2]));
	jspl3 jspl3_w_asqrt46_16(.douta(w_asqrt46_16[0]),.doutb(w_asqrt46_16[1]),.doutc(w_asqrt46_16[2]),.din(w_asqrt46_5[0]));
	jspl3 jspl3_w_asqrt46_17(.douta(w_asqrt46_17[0]),.doutb(w_asqrt46_17[1]),.doutc(w_asqrt46_17[2]),.din(w_asqrt46_5[1]));
	jspl3 jspl3_w_asqrt46_18(.douta(w_asqrt46_18[0]),.doutb(w_asqrt46_18[1]),.doutc(w_asqrt46_18[2]),.din(w_asqrt46_5[2]));
	jspl3 jspl3_w_asqrt46_19(.douta(w_asqrt46_19[0]),.doutb(w_asqrt46_19[1]),.doutc(w_asqrt46_19[2]),.din(w_asqrt46_6[0]));
	jspl3 jspl3_w_asqrt46_20(.douta(w_asqrt46_20[0]),.doutb(w_asqrt46_20[1]),.doutc(w_asqrt46_20[2]),.din(w_asqrt46_6[1]));
	jspl3 jspl3_w_asqrt46_21(.douta(w_asqrt46_21[0]),.doutb(w_asqrt46_21[1]),.doutc(w_asqrt46_21[2]),.din(w_asqrt46_6[2]));
	jspl3 jspl3_w_asqrt46_22(.douta(w_asqrt46_22[0]),.doutb(w_asqrt46_22[1]),.doutc(w_asqrt46_22[2]),.din(w_asqrt46_7[0]));
	jspl3 jspl3_w_asqrt46_23(.douta(w_asqrt46_23[0]),.doutb(w_asqrt46_23[1]),.doutc(w_asqrt46_23[2]),.din(w_asqrt46_7[1]));
	jspl3 jspl3_w_asqrt46_24(.douta(w_asqrt46_24[0]),.doutb(w_asqrt46_24[1]),.doutc(w_asqrt46_24[2]),.din(w_asqrt46_7[2]));
	jspl3 jspl3_w_asqrt46_25(.douta(w_asqrt46_25[0]),.doutb(w_asqrt46_25[1]),.doutc(w_asqrt46_25[2]),.din(w_asqrt46_8[0]));
	jspl3 jspl3_w_asqrt46_26(.douta(w_asqrt46_26[0]),.doutb(w_asqrt46_26[1]),.doutc(w_asqrt46_26[2]),.din(w_asqrt46_8[1]));
	jspl3 jspl3_w_asqrt46_27(.douta(w_asqrt46_27[0]),.doutb(w_asqrt46_27[1]),.doutc(w_asqrt46_27[2]),.din(w_asqrt46_8[2]));
	jspl3 jspl3_w_asqrt46_28(.douta(w_asqrt46_28[0]),.doutb(w_asqrt46_28[1]),.doutc(w_asqrt46_28[2]),.din(w_asqrt46_9[0]));
	jspl3 jspl3_w_asqrt46_29(.douta(w_asqrt46_29[0]),.doutb(w_asqrt46_29[1]),.doutc(w_asqrt46_29[2]),.din(w_asqrt46_9[1]));
	jspl3 jspl3_w_asqrt46_30(.douta(w_asqrt46_30[0]),.doutb(w_asqrt46_30[1]),.doutc(w_asqrt46_30[2]),.din(w_asqrt46_9[2]));
	jspl jspl_w_asqrt46_31(.douta(w_asqrt46_31),.doutb(asqrt[45]),.din(w_asqrt46_10[0]));
	jspl3 jspl3_w_asqrt47_0(.douta(w_asqrt47_0[0]),.doutb(w_asqrt47_0[1]),.doutc(w_asqrt47_0[2]),.din(asqrt_fa_47));
	jspl3 jspl3_w_asqrt47_1(.douta(w_asqrt47_1[0]),.doutb(w_asqrt47_1[1]),.doutc(w_asqrt47_1[2]),.din(w_asqrt47_0[0]));
	jspl3 jspl3_w_asqrt47_2(.douta(w_asqrt47_2[0]),.doutb(w_asqrt47_2[1]),.doutc(w_asqrt47_2[2]),.din(w_asqrt47_0[1]));
	jspl3 jspl3_w_asqrt47_3(.douta(w_asqrt47_3[0]),.doutb(w_asqrt47_3[1]),.doutc(w_asqrt47_3[2]),.din(w_asqrt47_0[2]));
	jspl3 jspl3_w_asqrt47_4(.douta(w_asqrt47_4[0]),.doutb(w_asqrt47_4[1]),.doutc(w_asqrt47_4[2]),.din(w_asqrt47_1[0]));
	jspl3 jspl3_w_asqrt47_5(.douta(w_asqrt47_5[0]),.doutb(w_asqrt47_5[1]),.doutc(w_asqrt47_5[2]),.din(w_asqrt47_1[1]));
	jspl3 jspl3_w_asqrt47_6(.douta(w_asqrt47_6[0]),.doutb(w_asqrt47_6[1]),.doutc(w_asqrt47_6[2]),.din(w_asqrt47_1[2]));
	jspl3 jspl3_w_asqrt47_7(.douta(w_asqrt47_7[0]),.doutb(w_asqrt47_7[1]),.doutc(w_asqrt47_7[2]),.din(w_asqrt47_2[0]));
	jspl3 jspl3_w_asqrt47_8(.douta(w_asqrt47_8[0]),.doutb(w_asqrt47_8[1]),.doutc(w_asqrt47_8[2]),.din(w_asqrt47_2[1]));
	jspl3 jspl3_w_asqrt47_9(.douta(w_asqrt47_9[0]),.doutb(w_asqrt47_9[1]),.doutc(w_asqrt47_9[2]),.din(w_asqrt47_2[2]));
	jspl3 jspl3_w_asqrt47_10(.douta(w_asqrt47_10[0]),.doutb(w_asqrt47_10[1]),.doutc(w_asqrt47_10[2]),.din(w_asqrt47_3[0]));
	jspl3 jspl3_w_asqrt47_11(.douta(w_asqrt47_11[0]),.doutb(w_asqrt47_11[1]),.doutc(w_asqrt47_11[2]),.din(w_asqrt47_3[1]));
	jspl3 jspl3_w_asqrt47_12(.douta(w_asqrt47_12[0]),.doutb(w_asqrt47_12[1]),.doutc(w_asqrt47_12[2]),.din(w_asqrt47_3[2]));
	jspl3 jspl3_w_asqrt47_13(.douta(w_asqrt47_13[0]),.doutb(w_asqrt47_13[1]),.doutc(w_asqrt47_13[2]),.din(w_asqrt47_4[0]));
	jspl3 jspl3_w_asqrt47_14(.douta(w_asqrt47_14[0]),.doutb(w_asqrt47_14[1]),.doutc(w_asqrt47_14[2]),.din(w_asqrt47_4[1]));
	jspl3 jspl3_w_asqrt47_15(.douta(w_asqrt47_15[0]),.doutb(w_asqrt47_15[1]),.doutc(w_asqrt47_15[2]),.din(w_asqrt47_4[2]));
	jspl3 jspl3_w_asqrt47_16(.douta(w_asqrt47_16[0]),.doutb(w_asqrt47_16[1]),.doutc(w_asqrt47_16[2]),.din(w_asqrt47_5[0]));
	jspl3 jspl3_w_asqrt47_17(.douta(w_asqrt47_17[0]),.doutb(w_asqrt47_17[1]),.doutc(w_asqrt47_17[2]),.din(w_asqrt47_5[1]));
	jspl3 jspl3_w_asqrt47_18(.douta(w_asqrt47_18[0]),.doutb(w_asqrt47_18[1]),.doutc(w_asqrt47_18[2]),.din(w_asqrt47_5[2]));
	jspl3 jspl3_w_asqrt47_19(.douta(w_asqrt47_19[0]),.doutb(w_asqrt47_19[1]),.doutc(w_asqrt47_19[2]),.din(w_asqrt47_6[0]));
	jspl3 jspl3_w_asqrt47_20(.douta(w_asqrt47_20[0]),.doutb(w_asqrt47_20[1]),.doutc(w_asqrt47_20[2]),.din(w_asqrt47_6[1]));
	jspl3 jspl3_w_asqrt47_21(.douta(w_asqrt47_21[0]),.doutb(w_asqrt47_21[1]),.doutc(w_asqrt47_21[2]),.din(w_asqrt47_6[2]));
	jspl3 jspl3_w_asqrt47_22(.douta(w_asqrt47_22[0]),.doutb(w_asqrt47_22[1]),.doutc(w_asqrt47_22[2]),.din(w_asqrt47_7[0]));
	jspl3 jspl3_w_asqrt47_23(.douta(w_asqrt47_23[0]),.doutb(w_asqrt47_23[1]),.doutc(w_asqrt47_23[2]),.din(w_asqrt47_7[1]));
	jspl3 jspl3_w_asqrt47_24(.douta(w_asqrt47_24[0]),.doutb(w_asqrt47_24[1]),.doutc(w_asqrt47_24[2]),.din(w_asqrt47_7[2]));
	jspl3 jspl3_w_asqrt47_25(.douta(w_asqrt47_25[0]),.doutb(w_asqrt47_25[1]),.doutc(asqrt[46]),.din(w_asqrt47_8[0]));
	jspl3 jspl3_w_asqrt48_0(.douta(w_asqrt48_0[0]),.doutb(w_asqrt48_0[1]),.doutc(w_asqrt48_0[2]),.din(asqrt_fa_48));
	jspl3 jspl3_w_asqrt48_1(.douta(w_asqrt48_1[0]),.doutb(w_asqrt48_1[1]),.doutc(w_asqrt48_1[2]),.din(w_asqrt48_0[0]));
	jspl3 jspl3_w_asqrt48_2(.douta(w_asqrt48_2[0]),.doutb(w_asqrt48_2[1]),.doutc(w_asqrt48_2[2]),.din(w_asqrt48_0[1]));
	jspl3 jspl3_w_asqrt48_3(.douta(w_asqrt48_3[0]),.doutb(w_asqrt48_3[1]),.doutc(w_asqrt48_3[2]),.din(w_asqrt48_0[2]));
	jspl3 jspl3_w_asqrt48_4(.douta(w_asqrt48_4[0]),.doutb(w_asqrt48_4[1]),.doutc(w_asqrt48_4[2]),.din(w_asqrt48_1[0]));
	jspl3 jspl3_w_asqrt48_5(.douta(w_asqrt48_5[0]),.doutb(w_asqrt48_5[1]),.doutc(w_asqrt48_5[2]),.din(w_asqrt48_1[1]));
	jspl3 jspl3_w_asqrt48_6(.douta(w_asqrt48_6[0]),.doutb(w_asqrt48_6[1]),.doutc(w_asqrt48_6[2]),.din(w_asqrt48_1[2]));
	jspl3 jspl3_w_asqrt48_7(.douta(w_asqrt48_7[0]),.doutb(w_asqrt48_7[1]),.doutc(w_asqrt48_7[2]),.din(w_asqrt48_2[0]));
	jspl3 jspl3_w_asqrt48_8(.douta(w_asqrt48_8[0]),.doutb(w_asqrt48_8[1]),.doutc(w_asqrt48_8[2]),.din(w_asqrt48_2[1]));
	jspl3 jspl3_w_asqrt48_9(.douta(w_asqrt48_9[0]),.doutb(w_asqrt48_9[1]),.doutc(w_asqrt48_9[2]),.din(w_asqrt48_2[2]));
	jspl3 jspl3_w_asqrt48_10(.douta(w_asqrt48_10[0]),.doutb(w_asqrt48_10[1]),.doutc(w_asqrt48_10[2]),.din(w_asqrt48_3[0]));
	jspl3 jspl3_w_asqrt48_11(.douta(w_asqrt48_11[0]),.doutb(w_asqrt48_11[1]),.doutc(w_asqrt48_11[2]),.din(w_asqrt48_3[1]));
	jspl3 jspl3_w_asqrt48_12(.douta(w_asqrt48_12[0]),.doutb(w_asqrt48_12[1]),.doutc(w_asqrt48_12[2]),.din(w_asqrt48_3[2]));
	jspl3 jspl3_w_asqrt48_13(.douta(w_asqrt48_13[0]),.doutb(w_asqrt48_13[1]),.doutc(w_asqrt48_13[2]),.din(w_asqrt48_4[0]));
	jspl3 jspl3_w_asqrt48_14(.douta(w_asqrt48_14[0]),.doutb(w_asqrt48_14[1]),.doutc(w_asqrt48_14[2]),.din(w_asqrt48_4[1]));
	jspl3 jspl3_w_asqrt48_15(.douta(w_asqrt48_15[0]),.doutb(w_asqrt48_15[1]),.doutc(w_asqrt48_15[2]),.din(w_asqrt48_4[2]));
	jspl3 jspl3_w_asqrt48_16(.douta(w_asqrt48_16[0]),.doutb(w_asqrt48_16[1]),.doutc(w_asqrt48_16[2]),.din(w_asqrt48_5[0]));
	jspl3 jspl3_w_asqrt48_17(.douta(w_asqrt48_17[0]),.doutb(w_asqrt48_17[1]),.doutc(w_asqrt48_17[2]),.din(w_asqrt48_5[1]));
	jspl3 jspl3_w_asqrt48_18(.douta(w_asqrt48_18[0]),.doutb(w_asqrt48_18[1]),.doutc(w_asqrt48_18[2]),.din(w_asqrt48_5[2]));
	jspl3 jspl3_w_asqrt48_19(.douta(w_asqrt48_19[0]),.doutb(w_asqrt48_19[1]),.doutc(w_asqrt48_19[2]),.din(w_asqrt48_6[0]));
	jspl3 jspl3_w_asqrt48_20(.douta(w_asqrt48_20[0]),.doutb(w_asqrt48_20[1]),.doutc(w_asqrt48_20[2]),.din(w_asqrt48_6[1]));
	jspl3 jspl3_w_asqrt48_21(.douta(w_asqrt48_21[0]),.doutb(w_asqrt48_21[1]),.doutc(w_asqrt48_21[2]),.din(w_asqrt48_6[2]));
	jspl3 jspl3_w_asqrt48_22(.douta(w_asqrt48_22[0]),.doutb(w_asqrt48_22[1]),.doutc(w_asqrt48_22[2]),.din(w_asqrt48_7[0]));
	jspl3 jspl3_w_asqrt48_23(.douta(w_asqrt48_23[0]),.doutb(w_asqrt48_23[1]),.doutc(w_asqrt48_23[2]),.din(w_asqrt48_7[1]));
	jspl3 jspl3_w_asqrt48_24(.douta(w_asqrt48_24[0]),.doutb(w_asqrt48_24[1]),.doutc(w_asqrt48_24[2]),.din(w_asqrt48_7[2]));
	jspl3 jspl3_w_asqrt48_25(.douta(w_asqrt48_25[0]),.doutb(w_asqrt48_25[1]),.doutc(w_asqrt48_25[2]),.din(w_asqrt48_8[0]));
	jspl3 jspl3_w_asqrt48_26(.douta(w_asqrt48_26[0]),.doutb(w_asqrt48_26[1]),.doutc(w_asqrt48_26[2]),.din(w_asqrt48_8[1]));
	jspl3 jspl3_w_asqrt48_27(.douta(w_asqrt48_27[0]),.doutb(w_asqrt48_27[1]),.doutc(w_asqrt48_27[2]),.din(w_asqrt48_8[2]));
	jspl3 jspl3_w_asqrt48_28(.douta(w_asqrt48_28[0]),.doutb(w_asqrt48_28[1]),.doutc(w_asqrt48_28[2]),.din(w_asqrt48_9[0]));
	jspl3 jspl3_w_asqrt48_29(.douta(w_asqrt48_29[0]),.doutb(w_asqrt48_29[1]),.doutc(w_asqrt48_29[2]),.din(w_asqrt48_9[1]));
	jspl3 jspl3_w_asqrt48_30(.douta(w_asqrt48_30[0]),.doutb(w_asqrt48_30[1]),.doutc(w_asqrt48_30[2]),.din(w_asqrt48_9[2]));
	jspl jspl_w_asqrt48_31(.douta(w_asqrt48_31),.doutb(asqrt[47]),.din(w_asqrt48_10[0]));
	jspl3 jspl3_w_asqrt49_0(.douta(w_asqrt49_0[0]),.doutb(w_asqrt49_0[1]),.doutc(w_asqrt49_0[2]),.din(asqrt_fa_49));
	jspl3 jspl3_w_asqrt49_1(.douta(w_asqrt49_1[0]),.doutb(w_asqrt49_1[1]),.doutc(w_asqrt49_1[2]),.din(w_asqrt49_0[0]));
	jspl3 jspl3_w_asqrt49_2(.douta(w_asqrt49_2[0]),.doutb(w_asqrt49_2[1]),.doutc(w_asqrt49_2[2]),.din(w_asqrt49_0[1]));
	jspl3 jspl3_w_asqrt49_3(.douta(w_asqrt49_3[0]),.doutb(w_asqrt49_3[1]),.doutc(w_asqrt49_3[2]),.din(w_asqrt49_0[2]));
	jspl3 jspl3_w_asqrt49_4(.douta(w_asqrt49_4[0]),.doutb(w_asqrt49_4[1]),.doutc(w_asqrt49_4[2]),.din(w_asqrt49_1[0]));
	jspl3 jspl3_w_asqrt49_5(.douta(w_asqrt49_5[0]),.doutb(w_asqrt49_5[1]),.doutc(w_asqrt49_5[2]),.din(w_asqrt49_1[1]));
	jspl3 jspl3_w_asqrt49_6(.douta(w_asqrt49_6[0]),.doutb(w_asqrt49_6[1]),.doutc(w_asqrt49_6[2]),.din(w_asqrt49_1[2]));
	jspl3 jspl3_w_asqrt49_7(.douta(w_asqrt49_7[0]),.doutb(w_asqrt49_7[1]),.doutc(w_asqrt49_7[2]),.din(w_asqrt49_2[0]));
	jspl3 jspl3_w_asqrt49_8(.douta(w_asqrt49_8[0]),.doutb(w_asqrt49_8[1]),.doutc(w_asqrt49_8[2]),.din(w_asqrt49_2[1]));
	jspl3 jspl3_w_asqrt49_9(.douta(w_asqrt49_9[0]),.doutb(w_asqrt49_9[1]),.doutc(w_asqrt49_9[2]),.din(w_asqrt49_2[2]));
	jspl3 jspl3_w_asqrt49_10(.douta(w_asqrt49_10[0]),.doutb(w_asqrt49_10[1]),.doutc(w_asqrt49_10[2]),.din(w_asqrt49_3[0]));
	jspl3 jspl3_w_asqrt49_11(.douta(w_asqrt49_11[0]),.doutb(w_asqrt49_11[1]),.doutc(w_asqrt49_11[2]),.din(w_asqrt49_3[1]));
	jspl3 jspl3_w_asqrt49_12(.douta(w_asqrt49_12[0]),.doutb(w_asqrt49_12[1]),.doutc(w_asqrt49_12[2]),.din(w_asqrt49_3[2]));
	jspl3 jspl3_w_asqrt49_13(.douta(w_asqrt49_13[0]),.doutb(w_asqrt49_13[1]),.doutc(w_asqrt49_13[2]),.din(w_asqrt49_4[0]));
	jspl3 jspl3_w_asqrt49_14(.douta(w_asqrt49_14[0]),.doutb(w_asqrt49_14[1]),.doutc(w_asqrt49_14[2]),.din(w_asqrt49_4[1]));
	jspl3 jspl3_w_asqrt49_15(.douta(w_asqrt49_15[0]),.doutb(w_asqrt49_15[1]),.doutc(w_asqrt49_15[2]),.din(w_asqrt49_4[2]));
	jspl3 jspl3_w_asqrt49_16(.douta(w_asqrt49_16[0]),.doutb(w_asqrt49_16[1]),.doutc(w_asqrt49_16[2]),.din(w_asqrt49_5[0]));
	jspl3 jspl3_w_asqrt49_17(.douta(w_asqrt49_17[0]),.doutb(w_asqrt49_17[1]),.doutc(w_asqrt49_17[2]),.din(w_asqrt49_5[1]));
	jspl3 jspl3_w_asqrt49_18(.douta(w_asqrt49_18[0]),.doutb(w_asqrt49_18[1]),.doutc(w_asqrt49_18[2]),.din(w_asqrt49_5[2]));
	jspl3 jspl3_w_asqrt49_19(.douta(w_asqrt49_19[0]),.doutb(w_asqrt49_19[1]),.doutc(w_asqrt49_19[2]),.din(w_asqrt49_6[0]));
	jspl3 jspl3_w_asqrt49_20(.douta(w_asqrt49_20[0]),.doutb(w_asqrt49_20[1]),.doutc(w_asqrt49_20[2]),.din(w_asqrt49_6[1]));
	jspl3 jspl3_w_asqrt49_21(.douta(w_asqrt49_21[0]),.doutb(w_asqrt49_21[1]),.doutc(w_asqrt49_21[2]),.din(w_asqrt49_6[2]));
	jspl3 jspl3_w_asqrt49_22(.douta(w_asqrt49_22[0]),.doutb(w_asqrt49_22[1]),.doutc(w_asqrt49_22[2]),.din(w_asqrt49_7[0]));
	jspl3 jspl3_w_asqrt49_23(.douta(w_asqrt49_23[0]),.doutb(w_asqrt49_23[1]),.doutc(w_asqrt49_23[2]),.din(w_asqrt49_7[1]));
	jspl3 jspl3_w_asqrt49_24(.douta(w_asqrt49_24[0]),.doutb(w_asqrt49_24[1]),.doutc(w_asqrt49_24[2]),.din(w_asqrt49_7[2]));
	jspl3 jspl3_w_asqrt49_25(.douta(w_asqrt49_25[0]),.doutb(w_asqrt49_25[1]),.doutc(w_asqrt49_25[2]),.din(w_asqrt49_8[0]));
	jspl3 jspl3_w_asqrt49_26(.douta(w_asqrt49_26[0]),.doutb(w_asqrt49_26[1]),.doutc(asqrt[48]),.din(w_asqrt49_8[1]));
	jspl3 jspl3_w_asqrt50_0(.douta(w_asqrt50_0[0]),.doutb(w_asqrt50_0[1]),.doutc(w_asqrt50_0[2]),.din(asqrt_fa_50));
	jspl3 jspl3_w_asqrt50_1(.douta(w_asqrt50_1[0]),.doutb(w_asqrt50_1[1]),.doutc(w_asqrt50_1[2]),.din(w_asqrt50_0[0]));
	jspl3 jspl3_w_asqrt50_2(.douta(w_asqrt50_2[0]),.doutb(w_asqrt50_2[1]),.doutc(w_asqrt50_2[2]),.din(w_asqrt50_0[1]));
	jspl3 jspl3_w_asqrt50_3(.douta(w_asqrt50_3[0]),.doutb(w_asqrt50_3[1]),.doutc(w_asqrt50_3[2]),.din(w_asqrt50_0[2]));
	jspl3 jspl3_w_asqrt50_4(.douta(w_asqrt50_4[0]),.doutb(w_asqrt50_4[1]),.doutc(w_asqrt50_4[2]),.din(w_asqrt50_1[0]));
	jspl3 jspl3_w_asqrt50_5(.douta(w_asqrt50_5[0]),.doutb(w_asqrt50_5[1]),.doutc(w_asqrt50_5[2]),.din(w_asqrt50_1[1]));
	jspl3 jspl3_w_asqrt50_6(.douta(w_asqrt50_6[0]),.doutb(w_asqrt50_6[1]),.doutc(w_asqrt50_6[2]),.din(w_asqrt50_1[2]));
	jspl3 jspl3_w_asqrt50_7(.douta(w_asqrt50_7[0]),.doutb(w_asqrt50_7[1]),.doutc(w_asqrt50_7[2]),.din(w_asqrt50_2[0]));
	jspl3 jspl3_w_asqrt50_8(.douta(w_asqrt50_8[0]),.doutb(w_asqrt50_8[1]),.doutc(w_asqrt50_8[2]),.din(w_asqrt50_2[1]));
	jspl3 jspl3_w_asqrt50_9(.douta(w_asqrt50_9[0]),.doutb(w_asqrt50_9[1]),.doutc(w_asqrt50_9[2]),.din(w_asqrt50_2[2]));
	jspl3 jspl3_w_asqrt50_10(.douta(w_asqrt50_10[0]),.doutb(w_asqrt50_10[1]),.doutc(w_asqrt50_10[2]),.din(w_asqrt50_3[0]));
	jspl3 jspl3_w_asqrt50_11(.douta(w_asqrt50_11[0]),.doutb(w_asqrt50_11[1]),.doutc(w_asqrt50_11[2]),.din(w_asqrt50_3[1]));
	jspl3 jspl3_w_asqrt50_12(.douta(w_asqrt50_12[0]),.doutb(w_asqrt50_12[1]),.doutc(w_asqrt50_12[2]),.din(w_asqrt50_3[2]));
	jspl3 jspl3_w_asqrt50_13(.douta(w_asqrt50_13[0]),.doutb(w_asqrt50_13[1]),.doutc(w_asqrt50_13[2]),.din(w_asqrt50_4[0]));
	jspl3 jspl3_w_asqrt50_14(.douta(w_asqrt50_14[0]),.doutb(w_asqrt50_14[1]),.doutc(w_asqrt50_14[2]),.din(w_asqrt50_4[1]));
	jspl3 jspl3_w_asqrt50_15(.douta(w_asqrt50_15[0]),.doutb(w_asqrt50_15[1]),.doutc(w_asqrt50_15[2]),.din(w_asqrt50_4[2]));
	jspl3 jspl3_w_asqrt50_16(.douta(w_asqrt50_16[0]),.doutb(w_asqrt50_16[1]),.doutc(w_asqrt50_16[2]),.din(w_asqrt50_5[0]));
	jspl3 jspl3_w_asqrt50_17(.douta(w_asqrt50_17[0]),.doutb(w_asqrt50_17[1]),.doutc(w_asqrt50_17[2]),.din(w_asqrt50_5[1]));
	jspl3 jspl3_w_asqrt50_18(.douta(w_asqrt50_18[0]),.doutb(w_asqrt50_18[1]),.doutc(w_asqrt50_18[2]),.din(w_asqrt50_5[2]));
	jspl3 jspl3_w_asqrt50_19(.douta(w_asqrt50_19[0]),.doutb(w_asqrt50_19[1]),.doutc(w_asqrt50_19[2]),.din(w_asqrt50_6[0]));
	jspl3 jspl3_w_asqrt50_20(.douta(w_asqrt50_20[0]),.doutb(w_asqrt50_20[1]),.doutc(w_asqrt50_20[2]),.din(w_asqrt50_6[1]));
	jspl3 jspl3_w_asqrt50_21(.douta(w_asqrt50_21[0]),.doutb(w_asqrt50_21[1]),.doutc(w_asqrt50_21[2]),.din(w_asqrt50_6[2]));
	jspl3 jspl3_w_asqrt50_22(.douta(w_asqrt50_22[0]),.doutb(w_asqrt50_22[1]),.doutc(w_asqrt50_22[2]),.din(w_asqrt50_7[0]));
	jspl3 jspl3_w_asqrt50_23(.douta(w_asqrt50_23[0]),.doutb(w_asqrt50_23[1]),.doutc(w_asqrt50_23[2]),.din(w_asqrt50_7[1]));
	jspl3 jspl3_w_asqrt50_24(.douta(w_asqrt50_24[0]),.doutb(w_asqrt50_24[1]),.doutc(w_asqrt50_24[2]),.din(w_asqrt50_7[2]));
	jspl3 jspl3_w_asqrt50_25(.douta(w_asqrt50_25[0]),.doutb(w_asqrt50_25[1]),.doutc(w_asqrt50_25[2]),.din(w_asqrt50_8[0]));
	jspl3 jspl3_w_asqrt50_26(.douta(w_asqrt50_26[0]),.doutb(w_asqrt50_26[1]),.doutc(w_asqrt50_26[2]),.din(w_asqrt50_8[1]));
	jspl3 jspl3_w_asqrt50_27(.douta(w_asqrt50_27[0]),.doutb(w_asqrt50_27[1]),.doutc(w_asqrt50_27[2]),.din(w_asqrt50_8[2]));
	jspl3 jspl3_w_asqrt50_28(.douta(w_asqrt50_28[0]),.doutb(w_asqrt50_28[1]),.doutc(w_asqrt50_28[2]),.din(w_asqrt50_9[0]));
	jspl3 jspl3_w_asqrt50_29(.douta(w_asqrt50_29[0]),.doutb(w_asqrt50_29[1]),.doutc(w_asqrt50_29[2]),.din(w_asqrt50_9[1]));
	jspl3 jspl3_w_asqrt50_30(.douta(w_asqrt50_30[0]),.doutb(w_asqrt50_30[1]),.doutc(w_asqrt50_30[2]),.din(w_asqrt50_9[2]));
	jspl jspl_w_asqrt50_31(.douta(w_asqrt50_31),.doutb(asqrt[49]),.din(w_asqrt50_10[0]));
	jspl3 jspl3_w_asqrt51_0(.douta(w_asqrt51_0[0]),.doutb(w_asqrt51_0[1]),.doutc(w_asqrt51_0[2]),.din(asqrt_fa_51));
	jspl3 jspl3_w_asqrt51_1(.douta(w_asqrt51_1[0]),.doutb(w_asqrt51_1[1]),.doutc(w_asqrt51_1[2]),.din(w_asqrt51_0[0]));
	jspl3 jspl3_w_asqrt51_2(.douta(w_asqrt51_2[0]),.doutb(w_asqrt51_2[1]),.doutc(w_asqrt51_2[2]),.din(w_asqrt51_0[1]));
	jspl3 jspl3_w_asqrt51_3(.douta(w_asqrt51_3[0]),.doutb(w_asqrt51_3[1]),.doutc(w_asqrt51_3[2]),.din(w_asqrt51_0[2]));
	jspl3 jspl3_w_asqrt51_4(.douta(w_asqrt51_4[0]),.doutb(w_asqrt51_4[1]),.doutc(w_asqrt51_4[2]),.din(w_asqrt51_1[0]));
	jspl3 jspl3_w_asqrt51_5(.douta(w_asqrt51_5[0]),.doutb(w_asqrt51_5[1]),.doutc(w_asqrt51_5[2]),.din(w_asqrt51_1[1]));
	jspl3 jspl3_w_asqrt51_6(.douta(w_asqrt51_6[0]),.doutb(w_asqrt51_6[1]),.doutc(w_asqrt51_6[2]),.din(w_asqrt51_1[2]));
	jspl3 jspl3_w_asqrt51_7(.douta(w_asqrt51_7[0]),.doutb(w_asqrt51_7[1]),.doutc(w_asqrt51_7[2]),.din(w_asqrt51_2[0]));
	jspl3 jspl3_w_asqrt51_8(.douta(w_asqrt51_8[0]),.doutb(w_asqrt51_8[1]),.doutc(w_asqrt51_8[2]),.din(w_asqrt51_2[1]));
	jspl3 jspl3_w_asqrt51_9(.douta(w_asqrt51_9[0]),.doutb(w_asqrt51_9[1]),.doutc(w_asqrt51_9[2]),.din(w_asqrt51_2[2]));
	jspl3 jspl3_w_asqrt51_10(.douta(w_asqrt51_10[0]),.doutb(w_asqrt51_10[1]),.doutc(w_asqrt51_10[2]),.din(w_asqrt51_3[0]));
	jspl3 jspl3_w_asqrt51_11(.douta(w_asqrt51_11[0]),.doutb(w_asqrt51_11[1]),.doutc(w_asqrt51_11[2]),.din(w_asqrt51_3[1]));
	jspl3 jspl3_w_asqrt51_12(.douta(w_asqrt51_12[0]),.doutb(w_asqrt51_12[1]),.doutc(w_asqrt51_12[2]),.din(w_asqrt51_3[2]));
	jspl3 jspl3_w_asqrt51_13(.douta(w_asqrt51_13[0]),.doutb(w_asqrt51_13[1]),.doutc(w_asqrt51_13[2]),.din(w_asqrt51_4[0]));
	jspl3 jspl3_w_asqrt51_14(.douta(w_asqrt51_14[0]),.doutb(w_asqrt51_14[1]),.doutc(w_asqrt51_14[2]),.din(w_asqrt51_4[1]));
	jspl3 jspl3_w_asqrt51_15(.douta(w_asqrt51_15[0]),.doutb(w_asqrt51_15[1]),.doutc(w_asqrt51_15[2]),.din(w_asqrt51_4[2]));
	jspl3 jspl3_w_asqrt51_16(.douta(w_asqrt51_16[0]),.doutb(w_asqrt51_16[1]),.doutc(w_asqrt51_16[2]),.din(w_asqrt51_5[0]));
	jspl3 jspl3_w_asqrt51_17(.douta(w_asqrt51_17[0]),.doutb(w_asqrt51_17[1]),.doutc(w_asqrt51_17[2]),.din(w_asqrt51_5[1]));
	jspl3 jspl3_w_asqrt51_18(.douta(w_asqrt51_18[0]),.doutb(w_asqrt51_18[1]),.doutc(w_asqrt51_18[2]),.din(w_asqrt51_5[2]));
	jspl3 jspl3_w_asqrt51_19(.douta(w_asqrt51_19[0]),.doutb(w_asqrt51_19[1]),.doutc(w_asqrt51_19[2]),.din(w_asqrt51_6[0]));
	jspl3 jspl3_w_asqrt51_20(.douta(w_asqrt51_20[0]),.doutb(w_asqrt51_20[1]),.doutc(w_asqrt51_20[2]),.din(w_asqrt51_6[1]));
	jspl3 jspl3_w_asqrt51_21(.douta(w_asqrt51_21[0]),.doutb(w_asqrt51_21[1]),.doutc(w_asqrt51_21[2]),.din(w_asqrt51_6[2]));
	jspl3 jspl3_w_asqrt51_22(.douta(w_asqrt51_22[0]),.doutb(w_asqrt51_22[1]),.doutc(w_asqrt51_22[2]),.din(w_asqrt51_7[0]));
	jspl3 jspl3_w_asqrt51_23(.douta(w_asqrt51_23[0]),.doutb(w_asqrt51_23[1]),.doutc(w_asqrt51_23[2]),.din(w_asqrt51_7[1]));
	jspl3 jspl3_w_asqrt51_24(.douta(w_asqrt51_24[0]),.doutb(w_asqrt51_24[1]),.doutc(w_asqrt51_24[2]),.din(w_asqrt51_7[2]));
	jspl3 jspl3_w_asqrt51_25(.douta(w_asqrt51_25[0]),.doutb(w_asqrt51_25[1]),.doutc(w_asqrt51_25[2]),.din(w_asqrt51_8[0]));
	jspl3 jspl3_w_asqrt51_26(.douta(w_asqrt51_26[0]),.doutb(w_asqrt51_26[1]),.doutc(asqrt[50]),.din(w_asqrt51_8[1]));
	jspl3 jspl3_w_asqrt52_0(.douta(w_asqrt52_0[0]),.doutb(w_asqrt52_0[1]),.doutc(w_asqrt52_0[2]),.din(asqrt_fa_52));
	jspl3 jspl3_w_asqrt52_1(.douta(w_asqrt52_1[0]),.doutb(w_asqrt52_1[1]),.doutc(w_asqrt52_1[2]),.din(w_asqrt52_0[0]));
	jspl3 jspl3_w_asqrt52_2(.douta(w_asqrt52_2[0]),.doutb(w_asqrt52_2[1]),.doutc(w_asqrt52_2[2]),.din(w_asqrt52_0[1]));
	jspl3 jspl3_w_asqrt52_3(.douta(w_asqrt52_3[0]),.doutb(w_asqrt52_3[1]),.doutc(w_asqrt52_3[2]),.din(w_asqrt52_0[2]));
	jspl3 jspl3_w_asqrt52_4(.douta(w_asqrt52_4[0]),.doutb(w_asqrt52_4[1]),.doutc(w_asqrt52_4[2]),.din(w_asqrt52_1[0]));
	jspl3 jspl3_w_asqrt52_5(.douta(w_asqrt52_5[0]),.doutb(w_asqrt52_5[1]),.doutc(w_asqrt52_5[2]),.din(w_asqrt52_1[1]));
	jspl3 jspl3_w_asqrt52_6(.douta(w_asqrt52_6[0]),.doutb(w_asqrt52_6[1]),.doutc(w_asqrt52_6[2]),.din(w_asqrt52_1[2]));
	jspl3 jspl3_w_asqrt52_7(.douta(w_asqrt52_7[0]),.doutb(w_asqrt52_7[1]),.doutc(w_asqrt52_7[2]),.din(w_asqrt52_2[0]));
	jspl3 jspl3_w_asqrt52_8(.douta(w_asqrt52_8[0]),.doutb(w_asqrt52_8[1]),.doutc(w_asqrt52_8[2]),.din(w_asqrt52_2[1]));
	jspl3 jspl3_w_asqrt52_9(.douta(w_asqrt52_9[0]),.doutb(w_asqrt52_9[1]),.doutc(w_asqrt52_9[2]),.din(w_asqrt52_2[2]));
	jspl3 jspl3_w_asqrt52_10(.douta(w_asqrt52_10[0]),.doutb(w_asqrt52_10[1]),.doutc(w_asqrt52_10[2]),.din(w_asqrt52_3[0]));
	jspl3 jspl3_w_asqrt52_11(.douta(w_asqrt52_11[0]),.doutb(w_asqrt52_11[1]),.doutc(w_asqrt52_11[2]),.din(w_asqrt52_3[1]));
	jspl3 jspl3_w_asqrt52_12(.douta(w_asqrt52_12[0]),.doutb(w_asqrt52_12[1]),.doutc(w_asqrt52_12[2]),.din(w_asqrt52_3[2]));
	jspl3 jspl3_w_asqrt52_13(.douta(w_asqrt52_13[0]),.doutb(w_asqrt52_13[1]),.doutc(w_asqrt52_13[2]),.din(w_asqrt52_4[0]));
	jspl3 jspl3_w_asqrt52_14(.douta(w_asqrt52_14[0]),.doutb(w_asqrt52_14[1]),.doutc(w_asqrt52_14[2]),.din(w_asqrt52_4[1]));
	jspl3 jspl3_w_asqrt52_15(.douta(w_asqrt52_15[0]),.doutb(w_asqrt52_15[1]),.doutc(w_asqrt52_15[2]),.din(w_asqrt52_4[2]));
	jspl3 jspl3_w_asqrt52_16(.douta(w_asqrt52_16[0]),.doutb(w_asqrt52_16[1]),.doutc(w_asqrt52_16[2]),.din(w_asqrt52_5[0]));
	jspl3 jspl3_w_asqrt52_17(.douta(w_asqrt52_17[0]),.doutb(w_asqrt52_17[1]),.doutc(w_asqrt52_17[2]),.din(w_asqrt52_5[1]));
	jspl3 jspl3_w_asqrt52_18(.douta(w_asqrt52_18[0]),.doutb(w_asqrt52_18[1]),.doutc(w_asqrt52_18[2]),.din(w_asqrt52_5[2]));
	jspl3 jspl3_w_asqrt52_19(.douta(w_asqrt52_19[0]),.doutb(w_asqrt52_19[1]),.doutc(w_asqrt52_19[2]),.din(w_asqrt52_6[0]));
	jspl3 jspl3_w_asqrt52_20(.douta(w_asqrt52_20[0]),.doutb(w_asqrt52_20[1]),.doutc(w_asqrt52_20[2]),.din(w_asqrt52_6[1]));
	jspl3 jspl3_w_asqrt52_21(.douta(w_asqrt52_21[0]),.doutb(w_asqrt52_21[1]),.doutc(w_asqrt52_21[2]),.din(w_asqrt52_6[2]));
	jspl3 jspl3_w_asqrt52_22(.douta(w_asqrt52_22[0]),.doutb(w_asqrt52_22[1]),.doutc(w_asqrt52_22[2]),.din(w_asqrt52_7[0]));
	jspl3 jspl3_w_asqrt52_23(.douta(w_asqrt52_23[0]),.doutb(w_asqrt52_23[1]),.doutc(w_asqrt52_23[2]),.din(w_asqrt52_7[1]));
	jspl3 jspl3_w_asqrt52_24(.douta(w_asqrt52_24[0]),.doutb(w_asqrt52_24[1]),.doutc(w_asqrt52_24[2]),.din(w_asqrt52_7[2]));
	jspl3 jspl3_w_asqrt52_25(.douta(w_asqrt52_25[0]),.doutb(w_asqrt52_25[1]),.doutc(w_asqrt52_25[2]),.din(w_asqrt52_8[0]));
	jspl3 jspl3_w_asqrt52_26(.douta(w_asqrt52_26[0]),.doutb(w_asqrt52_26[1]),.doutc(w_asqrt52_26[2]),.din(w_asqrt52_8[1]));
	jspl3 jspl3_w_asqrt52_27(.douta(w_asqrt52_27[0]),.doutb(w_asqrt52_27[1]),.doutc(w_asqrt52_27[2]),.din(w_asqrt52_8[2]));
	jspl3 jspl3_w_asqrt52_28(.douta(w_asqrt52_28[0]),.doutb(w_asqrt52_28[1]),.doutc(w_asqrt52_28[2]),.din(w_asqrt52_9[0]));
	jspl3 jspl3_w_asqrt52_29(.douta(w_asqrt52_29[0]),.doutb(w_asqrt52_29[1]),.doutc(w_asqrt52_29[2]),.din(w_asqrt52_9[1]));
	jspl3 jspl3_w_asqrt52_30(.douta(w_asqrt52_30[0]),.doutb(w_asqrt52_30[1]),.doutc(w_asqrt52_30[2]),.din(w_asqrt52_9[2]));
	jspl jspl_w_asqrt52_31(.douta(w_asqrt52_31),.doutb(asqrt[51]),.din(w_asqrt52_10[0]));
	jspl3 jspl3_w_asqrt53_0(.douta(w_asqrt53_0[0]),.doutb(w_asqrt53_0[1]),.doutc(w_asqrt53_0[2]),.din(asqrt_fa_53));
	jspl3 jspl3_w_asqrt53_1(.douta(w_asqrt53_1[0]),.doutb(w_asqrt53_1[1]),.doutc(w_asqrt53_1[2]),.din(w_asqrt53_0[0]));
	jspl3 jspl3_w_asqrt53_2(.douta(w_asqrt53_2[0]),.doutb(w_asqrt53_2[1]),.doutc(w_asqrt53_2[2]),.din(w_asqrt53_0[1]));
	jspl3 jspl3_w_asqrt53_3(.douta(w_asqrt53_3[0]),.doutb(w_asqrt53_3[1]),.doutc(w_asqrt53_3[2]),.din(w_asqrt53_0[2]));
	jspl3 jspl3_w_asqrt53_4(.douta(w_asqrt53_4[0]),.doutb(w_asqrt53_4[1]),.doutc(w_asqrt53_4[2]),.din(w_asqrt53_1[0]));
	jspl3 jspl3_w_asqrt53_5(.douta(w_asqrt53_5[0]),.doutb(w_asqrt53_5[1]),.doutc(w_asqrt53_5[2]),.din(w_asqrt53_1[1]));
	jspl3 jspl3_w_asqrt53_6(.douta(w_asqrt53_6[0]),.doutb(w_asqrt53_6[1]),.doutc(w_asqrt53_6[2]),.din(w_asqrt53_1[2]));
	jspl3 jspl3_w_asqrt53_7(.douta(w_asqrt53_7[0]),.doutb(w_asqrt53_7[1]),.doutc(w_asqrt53_7[2]),.din(w_asqrt53_2[0]));
	jspl3 jspl3_w_asqrt53_8(.douta(w_asqrt53_8[0]),.doutb(w_asqrt53_8[1]),.doutc(w_asqrt53_8[2]),.din(w_asqrt53_2[1]));
	jspl3 jspl3_w_asqrt53_9(.douta(w_asqrt53_9[0]),.doutb(w_asqrt53_9[1]),.doutc(w_asqrt53_9[2]),.din(w_asqrt53_2[2]));
	jspl3 jspl3_w_asqrt53_10(.douta(w_asqrt53_10[0]),.doutb(w_asqrt53_10[1]),.doutc(w_asqrt53_10[2]),.din(w_asqrt53_3[0]));
	jspl3 jspl3_w_asqrt53_11(.douta(w_asqrt53_11[0]),.doutb(w_asqrt53_11[1]),.doutc(w_asqrt53_11[2]),.din(w_asqrt53_3[1]));
	jspl3 jspl3_w_asqrt53_12(.douta(w_asqrt53_12[0]),.doutb(w_asqrt53_12[1]),.doutc(w_asqrt53_12[2]),.din(w_asqrt53_3[2]));
	jspl3 jspl3_w_asqrt53_13(.douta(w_asqrt53_13[0]),.doutb(w_asqrt53_13[1]),.doutc(w_asqrt53_13[2]),.din(w_asqrt53_4[0]));
	jspl3 jspl3_w_asqrt53_14(.douta(w_asqrt53_14[0]),.doutb(w_asqrt53_14[1]),.doutc(w_asqrt53_14[2]),.din(w_asqrt53_4[1]));
	jspl3 jspl3_w_asqrt53_15(.douta(w_asqrt53_15[0]),.doutb(w_asqrt53_15[1]),.doutc(w_asqrt53_15[2]),.din(w_asqrt53_4[2]));
	jspl3 jspl3_w_asqrt53_16(.douta(w_asqrt53_16[0]),.doutb(w_asqrt53_16[1]),.doutc(w_asqrt53_16[2]),.din(w_asqrt53_5[0]));
	jspl3 jspl3_w_asqrt53_17(.douta(w_asqrt53_17[0]),.doutb(w_asqrt53_17[1]),.doutc(w_asqrt53_17[2]),.din(w_asqrt53_5[1]));
	jspl3 jspl3_w_asqrt53_18(.douta(w_asqrt53_18[0]),.doutb(w_asqrt53_18[1]),.doutc(w_asqrt53_18[2]),.din(w_asqrt53_5[2]));
	jspl3 jspl3_w_asqrt53_19(.douta(w_asqrt53_19[0]),.doutb(w_asqrt53_19[1]),.doutc(w_asqrt53_19[2]),.din(w_asqrt53_6[0]));
	jspl3 jspl3_w_asqrt53_20(.douta(w_asqrt53_20[0]),.doutb(w_asqrt53_20[1]),.doutc(w_asqrt53_20[2]),.din(w_asqrt53_6[1]));
	jspl3 jspl3_w_asqrt53_21(.douta(w_asqrt53_21[0]),.doutb(w_asqrt53_21[1]),.doutc(w_asqrt53_21[2]),.din(w_asqrt53_6[2]));
	jspl3 jspl3_w_asqrt53_22(.douta(w_asqrt53_22[0]),.doutb(w_asqrt53_22[1]),.doutc(w_asqrt53_22[2]),.din(w_asqrt53_7[0]));
	jspl3 jspl3_w_asqrt53_23(.douta(w_asqrt53_23[0]),.doutb(w_asqrt53_23[1]),.doutc(w_asqrt53_23[2]),.din(w_asqrt53_7[1]));
	jspl3 jspl3_w_asqrt53_24(.douta(w_asqrt53_24[0]),.doutb(w_asqrt53_24[1]),.doutc(w_asqrt53_24[2]),.din(w_asqrt53_7[2]));
	jspl3 jspl3_w_asqrt53_25(.douta(w_asqrt53_25[0]),.doutb(w_asqrt53_25[1]),.doutc(w_asqrt53_25[2]),.din(w_asqrt53_8[0]));
	jspl3 jspl3_w_asqrt53_26(.douta(w_asqrt53_26[0]),.doutb(w_asqrt53_26[1]),.doutc(w_asqrt53_26[2]),.din(w_asqrt53_8[1]));
	jspl3 jspl3_w_asqrt53_27(.douta(w_asqrt53_27[0]),.doutb(w_asqrt53_27[1]),.doutc(asqrt[52]),.din(w_asqrt53_8[2]));
	jspl3 jspl3_w_asqrt54_0(.douta(w_asqrt54_0[0]),.doutb(w_asqrt54_0[1]),.doutc(w_asqrt54_0[2]),.din(asqrt_fa_54));
	jspl3 jspl3_w_asqrt54_1(.douta(w_asqrt54_1[0]),.doutb(w_asqrt54_1[1]),.doutc(w_asqrt54_1[2]),.din(w_asqrt54_0[0]));
	jspl3 jspl3_w_asqrt54_2(.douta(w_asqrt54_2[0]),.doutb(w_asqrt54_2[1]),.doutc(w_asqrt54_2[2]),.din(w_asqrt54_0[1]));
	jspl3 jspl3_w_asqrt54_3(.douta(w_asqrt54_3[0]),.doutb(w_asqrt54_3[1]),.doutc(w_asqrt54_3[2]),.din(w_asqrt54_0[2]));
	jspl3 jspl3_w_asqrt54_4(.douta(w_asqrt54_4[0]),.doutb(w_asqrt54_4[1]),.doutc(w_asqrt54_4[2]),.din(w_asqrt54_1[0]));
	jspl3 jspl3_w_asqrt54_5(.douta(w_asqrt54_5[0]),.doutb(w_asqrt54_5[1]),.doutc(w_asqrt54_5[2]),.din(w_asqrt54_1[1]));
	jspl3 jspl3_w_asqrt54_6(.douta(w_asqrt54_6[0]),.doutb(w_asqrt54_6[1]),.doutc(w_asqrt54_6[2]),.din(w_asqrt54_1[2]));
	jspl3 jspl3_w_asqrt54_7(.douta(w_asqrt54_7[0]),.doutb(w_asqrt54_7[1]),.doutc(w_asqrt54_7[2]),.din(w_asqrt54_2[0]));
	jspl3 jspl3_w_asqrt54_8(.douta(w_asqrt54_8[0]),.doutb(w_asqrt54_8[1]),.doutc(w_asqrt54_8[2]),.din(w_asqrt54_2[1]));
	jspl3 jspl3_w_asqrt54_9(.douta(w_asqrt54_9[0]),.doutb(w_asqrt54_9[1]),.doutc(w_asqrt54_9[2]),.din(w_asqrt54_2[2]));
	jspl3 jspl3_w_asqrt54_10(.douta(w_asqrt54_10[0]),.doutb(w_asqrt54_10[1]),.doutc(w_asqrt54_10[2]),.din(w_asqrt54_3[0]));
	jspl3 jspl3_w_asqrt54_11(.douta(w_asqrt54_11[0]),.doutb(w_asqrt54_11[1]),.doutc(w_asqrt54_11[2]),.din(w_asqrt54_3[1]));
	jspl3 jspl3_w_asqrt54_12(.douta(w_asqrt54_12[0]),.doutb(w_asqrt54_12[1]),.doutc(w_asqrt54_12[2]),.din(w_asqrt54_3[2]));
	jspl3 jspl3_w_asqrt54_13(.douta(w_asqrt54_13[0]),.doutb(w_asqrt54_13[1]),.doutc(w_asqrt54_13[2]),.din(w_asqrt54_4[0]));
	jspl3 jspl3_w_asqrt54_14(.douta(w_asqrt54_14[0]),.doutb(w_asqrt54_14[1]),.doutc(w_asqrt54_14[2]),.din(w_asqrt54_4[1]));
	jspl3 jspl3_w_asqrt54_15(.douta(w_asqrt54_15[0]),.doutb(w_asqrt54_15[1]),.doutc(w_asqrt54_15[2]),.din(w_asqrt54_4[2]));
	jspl3 jspl3_w_asqrt54_16(.douta(w_asqrt54_16[0]),.doutb(w_asqrt54_16[1]),.doutc(w_asqrt54_16[2]),.din(w_asqrt54_5[0]));
	jspl3 jspl3_w_asqrt54_17(.douta(w_asqrt54_17[0]),.doutb(w_asqrt54_17[1]),.doutc(w_asqrt54_17[2]),.din(w_asqrt54_5[1]));
	jspl3 jspl3_w_asqrt54_18(.douta(w_asqrt54_18[0]),.doutb(w_asqrt54_18[1]),.doutc(w_asqrt54_18[2]),.din(w_asqrt54_5[2]));
	jspl3 jspl3_w_asqrt54_19(.douta(w_asqrt54_19[0]),.doutb(w_asqrt54_19[1]),.doutc(w_asqrt54_19[2]),.din(w_asqrt54_6[0]));
	jspl3 jspl3_w_asqrt54_20(.douta(w_asqrt54_20[0]),.doutb(w_asqrt54_20[1]),.doutc(w_asqrt54_20[2]),.din(w_asqrt54_6[1]));
	jspl3 jspl3_w_asqrt54_21(.douta(w_asqrt54_21[0]),.doutb(w_asqrt54_21[1]),.doutc(w_asqrt54_21[2]),.din(w_asqrt54_6[2]));
	jspl3 jspl3_w_asqrt54_22(.douta(w_asqrt54_22[0]),.doutb(w_asqrt54_22[1]),.doutc(w_asqrt54_22[2]),.din(w_asqrt54_7[0]));
	jspl3 jspl3_w_asqrt54_23(.douta(w_asqrt54_23[0]),.doutb(w_asqrt54_23[1]),.doutc(w_asqrt54_23[2]),.din(w_asqrt54_7[1]));
	jspl3 jspl3_w_asqrt54_24(.douta(w_asqrt54_24[0]),.doutb(w_asqrt54_24[1]),.doutc(w_asqrt54_24[2]),.din(w_asqrt54_7[2]));
	jspl3 jspl3_w_asqrt54_25(.douta(w_asqrt54_25[0]),.doutb(w_asqrt54_25[1]),.doutc(w_asqrt54_25[2]),.din(w_asqrt54_8[0]));
	jspl3 jspl3_w_asqrt54_26(.douta(w_asqrt54_26[0]),.doutb(w_asqrt54_26[1]),.doutc(w_asqrt54_26[2]),.din(w_asqrt54_8[1]));
	jspl3 jspl3_w_asqrt54_27(.douta(w_asqrt54_27[0]),.doutb(w_asqrt54_27[1]),.doutc(w_asqrt54_27[2]),.din(w_asqrt54_8[2]));
	jspl3 jspl3_w_asqrt54_28(.douta(w_asqrt54_28[0]),.doutb(w_asqrt54_28[1]),.doutc(w_asqrt54_28[2]),.din(w_asqrt54_9[0]));
	jspl3 jspl3_w_asqrt54_29(.douta(w_asqrt54_29[0]),.doutb(w_asqrt54_29[1]),.doutc(w_asqrt54_29[2]),.din(w_asqrt54_9[1]));
	jspl3 jspl3_w_asqrt54_30(.douta(w_asqrt54_30[0]),.doutb(w_asqrt54_30[1]),.doutc(w_asqrt54_30[2]),.din(w_asqrt54_9[2]));
	jspl jspl_w_asqrt54_31(.douta(w_asqrt54_31),.doutb(asqrt[53]),.din(w_asqrt54_10[0]));
	jspl3 jspl3_w_asqrt55_0(.douta(w_asqrt55_0[0]),.doutb(w_asqrt55_0[1]),.doutc(w_asqrt55_0[2]),.din(asqrt_fa_55));
	jspl3 jspl3_w_asqrt55_1(.douta(w_asqrt55_1[0]),.doutb(w_asqrt55_1[1]),.doutc(w_asqrt55_1[2]),.din(w_asqrt55_0[0]));
	jspl3 jspl3_w_asqrt55_2(.douta(w_asqrt55_2[0]),.doutb(w_asqrt55_2[1]),.doutc(w_asqrt55_2[2]),.din(w_asqrt55_0[1]));
	jspl3 jspl3_w_asqrt55_3(.douta(w_asqrt55_3[0]),.doutb(w_asqrt55_3[1]),.doutc(w_asqrt55_3[2]),.din(w_asqrt55_0[2]));
	jspl3 jspl3_w_asqrt55_4(.douta(w_asqrt55_4[0]),.doutb(w_asqrt55_4[1]),.doutc(w_asqrt55_4[2]),.din(w_asqrt55_1[0]));
	jspl3 jspl3_w_asqrt55_5(.douta(w_asqrt55_5[0]),.doutb(w_asqrt55_5[1]),.doutc(w_asqrt55_5[2]),.din(w_asqrt55_1[1]));
	jspl3 jspl3_w_asqrt55_6(.douta(w_asqrt55_6[0]),.doutb(w_asqrt55_6[1]),.doutc(w_asqrt55_6[2]),.din(w_asqrt55_1[2]));
	jspl3 jspl3_w_asqrt55_7(.douta(w_asqrt55_7[0]),.doutb(w_asqrt55_7[1]),.doutc(w_asqrt55_7[2]),.din(w_asqrt55_2[0]));
	jspl3 jspl3_w_asqrt55_8(.douta(w_asqrt55_8[0]),.doutb(w_asqrt55_8[1]),.doutc(w_asqrt55_8[2]),.din(w_asqrt55_2[1]));
	jspl3 jspl3_w_asqrt55_9(.douta(w_asqrt55_9[0]),.doutb(w_asqrt55_9[1]),.doutc(w_asqrt55_9[2]),.din(w_asqrt55_2[2]));
	jspl3 jspl3_w_asqrt55_10(.douta(w_asqrt55_10[0]),.doutb(w_asqrt55_10[1]),.doutc(w_asqrt55_10[2]),.din(w_asqrt55_3[0]));
	jspl3 jspl3_w_asqrt55_11(.douta(w_asqrt55_11[0]),.doutb(w_asqrt55_11[1]),.doutc(w_asqrt55_11[2]),.din(w_asqrt55_3[1]));
	jspl3 jspl3_w_asqrt55_12(.douta(w_asqrt55_12[0]),.doutb(w_asqrt55_12[1]),.doutc(w_asqrt55_12[2]),.din(w_asqrt55_3[2]));
	jspl3 jspl3_w_asqrt55_13(.douta(w_asqrt55_13[0]),.doutb(w_asqrt55_13[1]),.doutc(w_asqrt55_13[2]),.din(w_asqrt55_4[0]));
	jspl3 jspl3_w_asqrt55_14(.douta(w_asqrt55_14[0]),.doutb(w_asqrt55_14[1]),.doutc(w_asqrt55_14[2]),.din(w_asqrt55_4[1]));
	jspl3 jspl3_w_asqrt55_15(.douta(w_asqrt55_15[0]),.doutb(w_asqrt55_15[1]),.doutc(w_asqrt55_15[2]),.din(w_asqrt55_4[2]));
	jspl3 jspl3_w_asqrt55_16(.douta(w_asqrt55_16[0]),.doutb(w_asqrt55_16[1]),.doutc(w_asqrt55_16[2]),.din(w_asqrt55_5[0]));
	jspl3 jspl3_w_asqrt55_17(.douta(w_asqrt55_17[0]),.doutb(w_asqrt55_17[1]),.doutc(w_asqrt55_17[2]),.din(w_asqrt55_5[1]));
	jspl3 jspl3_w_asqrt55_18(.douta(w_asqrt55_18[0]),.doutb(w_asqrt55_18[1]),.doutc(w_asqrt55_18[2]),.din(w_asqrt55_5[2]));
	jspl3 jspl3_w_asqrt55_19(.douta(w_asqrt55_19[0]),.doutb(w_asqrt55_19[1]),.doutc(w_asqrt55_19[2]),.din(w_asqrt55_6[0]));
	jspl3 jspl3_w_asqrt55_20(.douta(w_asqrt55_20[0]),.doutb(w_asqrt55_20[1]),.doutc(w_asqrt55_20[2]),.din(w_asqrt55_6[1]));
	jspl3 jspl3_w_asqrt55_21(.douta(w_asqrt55_21[0]),.doutb(w_asqrt55_21[1]),.doutc(w_asqrt55_21[2]),.din(w_asqrt55_6[2]));
	jspl3 jspl3_w_asqrt55_22(.douta(w_asqrt55_22[0]),.doutb(w_asqrt55_22[1]),.doutc(w_asqrt55_22[2]),.din(w_asqrt55_7[0]));
	jspl3 jspl3_w_asqrt55_23(.douta(w_asqrt55_23[0]),.doutb(w_asqrt55_23[1]),.doutc(w_asqrt55_23[2]),.din(w_asqrt55_7[1]));
	jspl3 jspl3_w_asqrt55_24(.douta(w_asqrt55_24[0]),.doutb(w_asqrt55_24[1]),.doutc(w_asqrt55_24[2]),.din(w_asqrt55_7[2]));
	jspl3 jspl3_w_asqrt55_25(.douta(w_asqrt55_25[0]),.doutb(w_asqrt55_25[1]),.doutc(w_asqrt55_25[2]),.din(w_asqrt55_8[0]));
	jspl3 jspl3_w_asqrt55_26(.douta(w_asqrt55_26[0]),.doutb(w_asqrt55_26[1]),.doutc(w_asqrt55_26[2]),.din(w_asqrt55_8[1]));
	jspl3 jspl3_w_asqrt55_27(.douta(w_asqrt55_27[0]),.doutb(w_asqrt55_27[1]),.doutc(w_asqrt55_27[2]),.din(w_asqrt55_8[2]));
	jspl jspl_w_asqrt55_28(.douta(w_asqrt55_28),.doutb(asqrt[54]),.din(w_asqrt55_9[0]));
	jspl3 jspl3_w_asqrt56_0(.douta(w_asqrt56_0[0]),.doutb(w_asqrt56_0[1]),.doutc(w_asqrt56_0[2]),.din(asqrt_fa_56));
	jspl3 jspl3_w_asqrt56_1(.douta(w_asqrt56_1[0]),.doutb(w_asqrt56_1[1]),.doutc(w_asqrt56_1[2]),.din(w_asqrt56_0[0]));
	jspl3 jspl3_w_asqrt56_2(.douta(w_asqrt56_2[0]),.doutb(w_asqrt56_2[1]),.doutc(w_asqrt56_2[2]),.din(w_asqrt56_0[1]));
	jspl3 jspl3_w_asqrt56_3(.douta(w_asqrt56_3[0]),.doutb(w_asqrt56_3[1]),.doutc(w_asqrt56_3[2]),.din(w_asqrt56_0[2]));
	jspl3 jspl3_w_asqrt56_4(.douta(w_asqrt56_4[0]),.doutb(w_asqrt56_4[1]),.doutc(w_asqrt56_4[2]),.din(w_asqrt56_1[0]));
	jspl3 jspl3_w_asqrt56_5(.douta(w_asqrt56_5[0]),.doutb(w_asqrt56_5[1]),.doutc(w_asqrt56_5[2]),.din(w_asqrt56_1[1]));
	jspl3 jspl3_w_asqrt56_6(.douta(w_asqrt56_6[0]),.doutb(w_asqrt56_6[1]),.doutc(w_asqrt56_6[2]),.din(w_asqrt56_1[2]));
	jspl3 jspl3_w_asqrt56_7(.douta(w_asqrt56_7[0]),.doutb(w_asqrt56_7[1]),.doutc(w_asqrt56_7[2]),.din(w_asqrt56_2[0]));
	jspl3 jspl3_w_asqrt56_8(.douta(w_asqrt56_8[0]),.doutb(w_asqrt56_8[1]),.doutc(w_asqrt56_8[2]),.din(w_asqrt56_2[1]));
	jspl3 jspl3_w_asqrt56_9(.douta(w_asqrt56_9[0]),.doutb(w_asqrt56_9[1]),.doutc(w_asqrt56_9[2]),.din(w_asqrt56_2[2]));
	jspl3 jspl3_w_asqrt56_10(.douta(w_asqrt56_10[0]),.doutb(w_asqrt56_10[1]),.doutc(w_asqrt56_10[2]),.din(w_asqrt56_3[0]));
	jspl3 jspl3_w_asqrt56_11(.douta(w_asqrt56_11[0]),.doutb(w_asqrt56_11[1]),.doutc(w_asqrt56_11[2]),.din(w_asqrt56_3[1]));
	jspl3 jspl3_w_asqrt56_12(.douta(w_asqrt56_12[0]),.doutb(w_asqrt56_12[1]),.doutc(w_asqrt56_12[2]),.din(w_asqrt56_3[2]));
	jspl3 jspl3_w_asqrt56_13(.douta(w_asqrt56_13[0]),.doutb(w_asqrt56_13[1]),.doutc(w_asqrt56_13[2]),.din(w_asqrt56_4[0]));
	jspl3 jspl3_w_asqrt56_14(.douta(w_asqrt56_14[0]),.doutb(w_asqrt56_14[1]),.doutc(w_asqrt56_14[2]),.din(w_asqrt56_4[1]));
	jspl3 jspl3_w_asqrt56_15(.douta(w_asqrt56_15[0]),.doutb(w_asqrt56_15[1]),.doutc(w_asqrt56_15[2]),.din(w_asqrt56_4[2]));
	jspl3 jspl3_w_asqrt56_16(.douta(w_asqrt56_16[0]),.doutb(w_asqrt56_16[1]),.doutc(w_asqrt56_16[2]),.din(w_asqrt56_5[0]));
	jspl3 jspl3_w_asqrt56_17(.douta(w_asqrt56_17[0]),.doutb(w_asqrt56_17[1]),.doutc(w_asqrt56_17[2]),.din(w_asqrt56_5[1]));
	jspl3 jspl3_w_asqrt56_18(.douta(w_asqrt56_18[0]),.doutb(w_asqrt56_18[1]),.doutc(w_asqrt56_18[2]),.din(w_asqrt56_5[2]));
	jspl3 jspl3_w_asqrt56_19(.douta(w_asqrt56_19[0]),.doutb(w_asqrt56_19[1]),.doutc(w_asqrt56_19[2]),.din(w_asqrt56_6[0]));
	jspl3 jspl3_w_asqrt56_20(.douta(w_asqrt56_20[0]),.doutb(w_asqrt56_20[1]),.doutc(w_asqrt56_20[2]),.din(w_asqrt56_6[1]));
	jspl3 jspl3_w_asqrt56_21(.douta(w_asqrt56_21[0]),.doutb(w_asqrt56_21[1]),.doutc(w_asqrt56_21[2]),.din(w_asqrt56_6[2]));
	jspl3 jspl3_w_asqrt56_22(.douta(w_asqrt56_22[0]),.doutb(w_asqrt56_22[1]),.doutc(w_asqrt56_22[2]),.din(w_asqrt56_7[0]));
	jspl3 jspl3_w_asqrt56_23(.douta(w_asqrt56_23[0]),.doutb(w_asqrt56_23[1]),.doutc(w_asqrt56_23[2]),.din(w_asqrt56_7[1]));
	jspl3 jspl3_w_asqrt56_24(.douta(w_asqrt56_24[0]),.doutb(w_asqrt56_24[1]),.doutc(w_asqrt56_24[2]),.din(w_asqrt56_7[2]));
	jspl3 jspl3_w_asqrt56_25(.douta(w_asqrt56_25[0]),.doutb(w_asqrt56_25[1]),.doutc(w_asqrt56_25[2]),.din(w_asqrt56_8[0]));
	jspl3 jspl3_w_asqrt56_26(.douta(w_asqrt56_26[0]),.doutb(w_asqrt56_26[1]),.doutc(w_asqrt56_26[2]),.din(w_asqrt56_8[1]));
	jspl3 jspl3_w_asqrt56_27(.douta(w_asqrt56_27[0]),.doutb(w_asqrt56_27[1]),.doutc(w_asqrt56_27[2]),.din(w_asqrt56_8[2]));
	jspl3 jspl3_w_asqrt56_28(.douta(w_asqrt56_28[0]),.doutb(w_asqrt56_28[1]),.doutc(w_asqrt56_28[2]),.din(w_asqrt56_9[0]));
	jspl3 jspl3_w_asqrt56_29(.douta(w_asqrt56_29[0]),.doutb(w_asqrt56_29[1]),.doutc(w_asqrt56_29[2]),.din(w_asqrt56_9[1]));
	jspl3 jspl3_w_asqrt56_30(.douta(w_asqrt56_30[0]),.doutb(w_asqrt56_30[1]),.doutc(w_asqrt56_30[2]),.din(w_asqrt56_9[2]));
	jspl jspl_w_asqrt56_31(.douta(w_asqrt56_31),.doutb(asqrt[55]),.din(w_asqrt56_10[0]));
	jspl3 jspl3_w_asqrt57_0(.douta(w_asqrt57_0[0]),.doutb(w_asqrt57_0[1]),.doutc(w_asqrt57_0[2]),.din(asqrt_fa_57));
	jspl3 jspl3_w_asqrt57_1(.douta(w_asqrt57_1[0]),.doutb(w_asqrt57_1[1]),.doutc(w_asqrt57_1[2]),.din(w_asqrt57_0[0]));
	jspl3 jspl3_w_asqrt57_2(.douta(w_asqrt57_2[0]),.doutb(w_asqrt57_2[1]),.doutc(w_asqrt57_2[2]),.din(w_asqrt57_0[1]));
	jspl3 jspl3_w_asqrt57_3(.douta(w_asqrt57_3[0]),.doutb(w_asqrt57_3[1]),.doutc(w_asqrt57_3[2]),.din(w_asqrt57_0[2]));
	jspl3 jspl3_w_asqrt57_4(.douta(w_asqrt57_4[0]),.doutb(w_asqrt57_4[1]),.doutc(w_asqrt57_4[2]),.din(w_asqrt57_1[0]));
	jspl3 jspl3_w_asqrt57_5(.douta(w_asqrt57_5[0]),.doutb(w_asqrt57_5[1]),.doutc(w_asqrt57_5[2]),.din(w_asqrt57_1[1]));
	jspl3 jspl3_w_asqrt57_6(.douta(w_asqrt57_6[0]),.doutb(w_asqrt57_6[1]),.doutc(w_asqrt57_6[2]),.din(w_asqrt57_1[2]));
	jspl3 jspl3_w_asqrt57_7(.douta(w_asqrt57_7[0]),.doutb(w_asqrt57_7[1]),.doutc(w_asqrt57_7[2]),.din(w_asqrt57_2[0]));
	jspl3 jspl3_w_asqrt57_8(.douta(w_asqrt57_8[0]),.doutb(w_asqrt57_8[1]),.doutc(w_asqrt57_8[2]),.din(w_asqrt57_2[1]));
	jspl3 jspl3_w_asqrt57_9(.douta(w_asqrt57_9[0]),.doutb(w_asqrt57_9[1]),.doutc(w_asqrt57_9[2]),.din(w_asqrt57_2[2]));
	jspl3 jspl3_w_asqrt57_10(.douta(w_asqrt57_10[0]),.doutb(w_asqrt57_10[1]),.doutc(w_asqrt57_10[2]),.din(w_asqrt57_3[0]));
	jspl3 jspl3_w_asqrt57_11(.douta(w_asqrt57_11[0]),.doutb(w_asqrt57_11[1]),.doutc(w_asqrt57_11[2]),.din(w_asqrt57_3[1]));
	jspl3 jspl3_w_asqrt57_12(.douta(w_asqrt57_12[0]),.doutb(w_asqrt57_12[1]),.doutc(w_asqrt57_12[2]),.din(w_asqrt57_3[2]));
	jspl3 jspl3_w_asqrt57_13(.douta(w_asqrt57_13[0]),.doutb(w_asqrt57_13[1]),.doutc(w_asqrt57_13[2]),.din(w_asqrt57_4[0]));
	jspl3 jspl3_w_asqrt57_14(.douta(w_asqrt57_14[0]),.doutb(w_asqrt57_14[1]),.doutc(w_asqrt57_14[2]),.din(w_asqrt57_4[1]));
	jspl3 jspl3_w_asqrt57_15(.douta(w_asqrt57_15[0]),.doutb(w_asqrt57_15[1]),.doutc(w_asqrt57_15[2]),.din(w_asqrt57_4[2]));
	jspl3 jspl3_w_asqrt57_16(.douta(w_asqrt57_16[0]),.doutb(w_asqrt57_16[1]),.doutc(w_asqrt57_16[2]),.din(w_asqrt57_5[0]));
	jspl3 jspl3_w_asqrt57_17(.douta(w_asqrt57_17[0]),.doutb(w_asqrt57_17[1]),.doutc(w_asqrt57_17[2]),.din(w_asqrt57_5[1]));
	jspl3 jspl3_w_asqrt57_18(.douta(w_asqrt57_18[0]),.doutb(w_asqrt57_18[1]),.doutc(w_asqrt57_18[2]),.din(w_asqrt57_5[2]));
	jspl3 jspl3_w_asqrt57_19(.douta(w_asqrt57_19[0]),.doutb(w_asqrt57_19[1]),.doutc(w_asqrt57_19[2]),.din(w_asqrt57_6[0]));
	jspl3 jspl3_w_asqrt57_20(.douta(w_asqrt57_20[0]),.doutb(w_asqrt57_20[1]),.doutc(w_asqrt57_20[2]),.din(w_asqrt57_6[1]));
	jspl3 jspl3_w_asqrt57_21(.douta(w_asqrt57_21[0]),.doutb(w_asqrt57_21[1]),.doutc(w_asqrt57_21[2]),.din(w_asqrt57_6[2]));
	jspl3 jspl3_w_asqrt57_22(.douta(w_asqrt57_22[0]),.doutb(w_asqrt57_22[1]),.doutc(w_asqrt57_22[2]),.din(w_asqrt57_7[0]));
	jspl3 jspl3_w_asqrt57_23(.douta(w_asqrt57_23[0]),.doutb(w_asqrt57_23[1]),.doutc(w_asqrt57_23[2]),.din(w_asqrt57_7[1]));
	jspl3 jspl3_w_asqrt57_24(.douta(w_asqrt57_24[0]),.doutb(w_asqrt57_24[1]),.doutc(w_asqrt57_24[2]),.din(w_asqrt57_7[2]));
	jspl3 jspl3_w_asqrt57_25(.douta(w_asqrt57_25[0]),.doutb(w_asqrt57_25[1]),.doutc(w_asqrt57_25[2]),.din(w_asqrt57_8[0]));
	jspl3 jspl3_w_asqrt57_26(.douta(w_asqrt57_26[0]),.doutb(w_asqrt57_26[1]),.doutc(w_asqrt57_26[2]),.din(w_asqrt57_8[1]));
	jspl3 jspl3_w_asqrt57_27(.douta(w_asqrt57_27[0]),.doutb(w_asqrt57_27[1]),.doutc(w_asqrt57_27[2]),.din(w_asqrt57_8[2]));
	jspl3 jspl3_w_asqrt57_28(.douta(w_asqrt57_28[0]),.doutb(w_asqrt57_28[1]),.doutc(w_asqrt57_28[2]),.din(w_asqrt57_9[0]));
	jspl jspl_w_asqrt57_29(.douta(w_asqrt57_29),.doutb(asqrt[56]),.din(w_asqrt57_9[1]));
	jspl3 jspl3_w_asqrt58_0(.douta(w_asqrt58_0[0]),.doutb(w_asqrt58_0[1]),.doutc(w_asqrt58_0[2]),.din(asqrt_fa_58));
	jspl3 jspl3_w_asqrt58_1(.douta(w_asqrt58_1[0]),.doutb(w_asqrt58_1[1]),.doutc(w_asqrt58_1[2]),.din(w_asqrt58_0[0]));
	jspl3 jspl3_w_asqrt58_2(.douta(w_asqrt58_2[0]),.doutb(w_asqrt58_2[1]),.doutc(w_asqrt58_2[2]),.din(w_asqrt58_0[1]));
	jspl3 jspl3_w_asqrt58_3(.douta(w_asqrt58_3[0]),.doutb(w_asqrt58_3[1]),.doutc(w_asqrt58_3[2]),.din(w_asqrt58_0[2]));
	jspl3 jspl3_w_asqrt58_4(.douta(w_asqrt58_4[0]),.doutb(w_asqrt58_4[1]),.doutc(w_asqrt58_4[2]),.din(w_asqrt58_1[0]));
	jspl3 jspl3_w_asqrt58_5(.douta(w_asqrt58_5[0]),.doutb(w_asqrt58_5[1]),.doutc(w_asqrt58_5[2]),.din(w_asqrt58_1[1]));
	jspl3 jspl3_w_asqrt58_6(.douta(w_asqrt58_6[0]),.doutb(w_asqrt58_6[1]),.doutc(w_asqrt58_6[2]),.din(w_asqrt58_1[2]));
	jspl3 jspl3_w_asqrt58_7(.douta(w_asqrt58_7[0]),.doutb(w_asqrt58_7[1]),.doutc(w_asqrt58_7[2]),.din(w_asqrt58_2[0]));
	jspl3 jspl3_w_asqrt58_8(.douta(w_asqrt58_8[0]),.doutb(w_asqrt58_8[1]),.doutc(w_asqrt58_8[2]),.din(w_asqrt58_2[1]));
	jspl3 jspl3_w_asqrt58_9(.douta(w_asqrt58_9[0]),.doutb(w_asqrt58_9[1]),.doutc(w_asqrt58_9[2]),.din(w_asqrt58_2[2]));
	jspl3 jspl3_w_asqrt58_10(.douta(w_asqrt58_10[0]),.doutb(w_asqrt58_10[1]),.doutc(w_asqrt58_10[2]),.din(w_asqrt58_3[0]));
	jspl3 jspl3_w_asqrt58_11(.douta(w_asqrt58_11[0]),.doutb(w_asqrt58_11[1]),.doutc(w_asqrt58_11[2]),.din(w_asqrt58_3[1]));
	jspl3 jspl3_w_asqrt58_12(.douta(w_asqrt58_12[0]),.doutb(w_asqrt58_12[1]),.doutc(w_asqrt58_12[2]),.din(w_asqrt58_3[2]));
	jspl3 jspl3_w_asqrt58_13(.douta(w_asqrt58_13[0]),.doutb(w_asqrt58_13[1]),.doutc(w_asqrt58_13[2]),.din(w_asqrt58_4[0]));
	jspl3 jspl3_w_asqrt58_14(.douta(w_asqrt58_14[0]),.doutb(w_asqrt58_14[1]),.doutc(w_asqrt58_14[2]),.din(w_asqrt58_4[1]));
	jspl3 jspl3_w_asqrt58_15(.douta(w_asqrt58_15[0]),.doutb(w_asqrt58_15[1]),.doutc(w_asqrt58_15[2]),.din(w_asqrt58_4[2]));
	jspl3 jspl3_w_asqrt58_16(.douta(w_asqrt58_16[0]),.doutb(w_asqrt58_16[1]),.doutc(w_asqrt58_16[2]),.din(w_asqrt58_5[0]));
	jspl3 jspl3_w_asqrt58_17(.douta(w_asqrt58_17[0]),.doutb(w_asqrt58_17[1]),.doutc(w_asqrt58_17[2]),.din(w_asqrt58_5[1]));
	jspl3 jspl3_w_asqrt58_18(.douta(w_asqrt58_18[0]),.doutb(w_asqrt58_18[1]),.doutc(w_asqrt58_18[2]),.din(w_asqrt58_5[2]));
	jspl3 jspl3_w_asqrt58_19(.douta(w_asqrt58_19[0]),.doutb(w_asqrt58_19[1]),.doutc(w_asqrt58_19[2]),.din(w_asqrt58_6[0]));
	jspl3 jspl3_w_asqrt58_20(.douta(w_asqrt58_20[0]),.doutb(w_asqrt58_20[1]),.doutc(w_asqrt58_20[2]),.din(w_asqrt58_6[1]));
	jspl3 jspl3_w_asqrt58_21(.douta(w_asqrt58_21[0]),.doutb(w_asqrt58_21[1]),.doutc(w_asqrt58_21[2]),.din(w_asqrt58_6[2]));
	jspl3 jspl3_w_asqrt58_22(.douta(w_asqrt58_22[0]),.doutb(w_asqrt58_22[1]),.doutc(w_asqrt58_22[2]),.din(w_asqrt58_7[0]));
	jspl3 jspl3_w_asqrt58_23(.douta(w_asqrt58_23[0]),.doutb(w_asqrt58_23[1]),.doutc(w_asqrt58_23[2]),.din(w_asqrt58_7[1]));
	jspl3 jspl3_w_asqrt58_24(.douta(w_asqrt58_24[0]),.doutb(w_asqrt58_24[1]),.doutc(w_asqrt58_24[2]),.din(w_asqrt58_7[2]));
	jspl3 jspl3_w_asqrt58_25(.douta(w_asqrt58_25[0]),.doutb(w_asqrt58_25[1]),.doutc(w_asqrt58_25[2]),.din(w_asqrt58_8[0]));
	jspl3 jspl3_w_asqrt58_26(.douta(w_asqrt58_26[0]),.doutb(w_asqrt58_26[1]),.doutc(w_asqrt58_26[2]),.din(w_asqrt58_8[1]));
	jspl3 jspl3_w_asqrt58_27(.douta(w_asqrt58_27[0]),.doutb(w_asqrt58_27[1]),.doutc(w_asqrt58_27[2]),.din(w_asqrt58_8[2]));
	jspl3 jspl3_w_asqrt58_28(.douta(w_asqrt58_28[0]),.doutb(w_asqrt58_28[1]),.doutc(w_asqrt58_28[2]),.din(w_asqrt58_9[0]));
	jspl3 jspl3_w_asqrt58_29(.douta(w_asqrt58_29[0]),.doutb(w_asqrt58_29[1]),.doutc(w_asqrt58_29[2]),.din(w_asqrt58_9[1]));
	jspl3 jspl3_w_asqrt58_30(.douta(w_asqrt58_30[0]),.doutb(w_asqrt58_30[1]),.doutc(w_asqrt58_30[2]),.din(w_asqrt58_9[2]));
	jspl jspl_w_asqrt58_31(.douta(w_asqrt58_31),.doutb(asqrt[57]),.din(w_asqrt58_10[0]));
	jspl3 jspl3_w_asqrt59_0(.douta(w_asqrt59_0[0]),.doutb(w_asqrt59_0[1]),.doutc(w_asqrt59_0[2]),.din(asqrt_fa_59));
	jspl3 jspl3_w_asqrt59_1(.douta(w_asqrt59_1[0]),.doutb(w_asqrt59_1[1]),.doutc(w_asqrt59_1[2]),.din(w_asqrt59_0[0]));
	jspl3 jspl3_w_asqrt59_2(.douta(w_asqrt59_2[0]),.doutb(w_asqrt59_2[1]),.doutc(w_asqrt59_2[2]),.din(w_asqrt59_0[1]));
	jspl3 jspl3_w_asqrt59_3(.douta(w_asqrt59_3[0]),.doutb(w_asqrt59_3[1]),.doutc(w_asqrt59_3[2]),.din(w_asqrt59_0[2]));
	jspl3 jspl3_w_asqrt59_4(.douta(w_asqrt59_4[0]),.doutb(w_asqrt59_4[1]),.doutc(w_asqrt59_4[2]),.din(w_asqrt59_1[0]));
	jspl3 jspl3_w_asqrt59_5(.douta(w_asqrt59_5[0]),.doutb(w_asqrt59_5[1]),.doutc(w_asqrt59_5[2]),.din(w_asqrt59_1[1]));
	jspl3 jspl3_w_asqrt59_6(.douta(w_asqrt59_6[0]),.doutb(w_asqrt59_6[1]),.doutc(w_asqrt59_6[2]),.din(w_asqrt59_1[2]));
	jspl3 jspl3_w_asqrt59_7(.douta(w_asqrt59_7[0]),.doutb(w_asqrt59_7[1]),.doutc(w_asqrt59_7[2]),.din(w_asqrt59_2[0]));
	jspl3 jspl3_w_asqrt59_8(.douta(w_asqrt59_8[0]),.doutb(w_asqrt59_8[1]),.doutc(w_asqrt59_8[2]),.din(w_asqrt59_2[1]));
	jspl3 jspl3_w_asqrt59_9(.douta(w_asqrt59_9[0]),.doutb(w_asqrt59_9[1]),.doutc(w_asqrt59_9[2]),.din(w_asqrt59_2[2]));
	jspl3 jspl3_w_asqrt59_10(.douta(w_asqrt59_10[0]),.doutb(w_asqrt59_10[1]),.doutc(w_asqrt59_10[2]),.din(w_asqrt59_3[0]));
	jspl3 jspl3_w_asqrt59_11(.douta(w_asqrt59_11[0]),.doutb(w_asqrt59_11[1]),.doutc(w_asqrt59_11[2]),.din(w_asqrt59_3[1]));
	jspl3 jspl3_w_asqrt59_12(.douta(w_asqrt59_12[0]),.doutb(w_asqrt59_12[1]),.doutc(w_asqrt59_12[2]),.din(w_asqrt59_3[2]));
	jspl3 jspl3_w_asqrt59_13(.douta(w_asqrt59_13[0]),.doutb(w_asqrt59_13[1]),.doutc(w_asqrt59_13[2]),.din(w_asqrt59_4[0]));
	jspl3 jspl3_w_asqrt59_14(.douta(w_asqrt59_14[0]),.doutb(w_asqrt59_14[1]),.doutc(w_asqrt59_14[2]),.din(w_asqrt59_4[1]));
	jspl3 jspl3_w_asqrt59_15(.douta(w_asqrt59_15[0]),.doutb(w_asqrt59_15[1]),.doutc(w_asqrt59_15[2]),.din(w_asqrt59_4[2]));
	jspl3 jspl3_w_asqrt59_16(.douta(w_asqrt59_16[0]),.doutb(w_asqrt59_16[1]),.doutc(w_asqrt59_16[2]),.din(w_asqrt59_5[0]));
	jspl3 jspl3_w_asqrt59_17(.douta(w_asqrt59_17[0]),.doutb(w_asqrt59_17[1]),.doutc(w_asqrt59_17[2]),.din(w_asqrt59_5[1]));
	jspl3 jspl3_w_asqrt59_18(.douta(w_asqrt59_18[0]),.doutb(w_asqrt59_18[1]),.doutc(w_asqrt59_18[2]),.din(w_asqrt59_5[2]));
	jspl3 jspl3_w_asqrt59_19(.douta(w_asqrt59_19[0]),.doutb(w_asqrt59_19[1]),.doutc(w_asqrt59_19[2]),.din(w_asqrt59_6[0]));
	jspl3 jspl3_w_asqrt59_20(.douta(w_asqrt59_20[0]),.doutb(w_asqrt59_20[1]),.doutc(w_asqrt59_20[2]),.din(w_asqrt59_6[1]));
	jspl3 jspl3_w_asqrt59_21(.douta(w_asqrt59_21[0]),.doutb(w_asqrt59_21[1]),.doutc(w_asqrt59_21[2]),.din(w_asqrt59_6[2]));
	jspl3 jspl3_w_asqrt59_22(.douta(w_asqrt59_22[0]),.doutb(w_asqrt59_22[1]),.doutc(w_asqrt59_22[2]),.din(w_asqrt59_7[0]));
	jspl3 jspl3_w_asqrt59_23(.douta(w_asqrt59_23[0]),.doutb(w_asqrt59_23[1]),.doutc(w_asqrt59_23[2]),.din(w_asqrt59_7[1]));
	jspl3 jspl3_w_asqrt59_24(.douta(w_asqrt59_24[0]),.doutb(w_asqrt59_24[1]),.doutc(w_asqrt59_24[2]),.din(w_asqrt59_7[2]));
	jspl3 jspl3_w_asqrt59_25(.douta(w_asqrt59_25[0]),.doutb(w_asqrt59_25[1]),.doutc(w_asqrt59_25[2]),.din(w_asqrt59_8[0]));
	jspl3 jspl3_w_asqrt59_26(.douta(w_asqrt59_26[0]),.doutb(w_asqrt59_26[1]),.doutc(w_asqrt59_26[2]),.din(w_asqrt59_8[1]));
	jspl3 jspl3_w_asqrt59_27(.douta(w_asqrt59_27[0]),.doutb(w_asqrt59_27[1]),.doutc(w_asqrt59_27[2]),.din(w_asqrt59_8[2]));
	jspl3 jspl3_w_asqrt59_28(.douta(w_asqrt59_28[0]),.doutb(w_asqrt59_28[1]),.doutc(w_asqrt59_28[2]),.din(w_asqrt59_9[0]));
	jspl3 jspl3_w_asqrt59_29(.douta(w_asqrt59_29[0]),.doutb(w_asqrt59_29[1]),.doutc(w_asqrt59_29[2]),.din(w_asqrt59_9[1]));
	jspl3 jspl3_w_asqrt59_30(.douta(w_asqrt59_30[0]),.doutb(w_asqrt59_30[1]),.doutc(asqrt[58]),.din(w_asqrt59_9[2]));
	jspl3 jspl3_w_asqrt60_0(.douta(w_asqrt60_0[0]),.doutb(w_asqrt60_0[1]),.doutc(w_asqrt60_0[2]),.din(asqrt_fa_60));
	jspl3 jspl3_w_asqrt60_1(.douta(w_asqrt60_1[0]),.doutb(w_asqrt60_1[1]),.doutc(w_asqrt60_1[2]),.din(w_asqrt60_0[0]));
	jspl3 jspl3_w_asqrt60_2(.douta(w_asqrt60_2[0]),.doutb(w_asqrt60_2[1]),.doutc(w_asqrt60_2[2]),.din(w_asqrt60_0[1]));
	jspl3 jspl3_w_asqrt60_3(.douta(w_asqrt60_3[0]),.doutb(w_asqrt60_3[1]),.doutc(w_asqrt60_3[2]),.din(w_asqrt60_0[2]));
	jspl3 jspl3_w_asqrt60_4(.douta(w_asqrt60_4[0]),.doutb(w_asqrt60_4[1]),.doutc(w_asqrt60_4[2]),.din(w_asqrt60_1[0]));
	jspl3 jspl3_w_asqrt60_5(.douta(w_asqrt60_5[0]),.doutb(w_asqrt60_5[1]),.doutc(w_asqrt60_5[2]),.din(w_asqrt60_1[1]));
	jspl3 jspl3_w_asqrt60_6(.douta(w_asqrt60_6[0]),.doutb(w_asqrt60_6[1]),.doutc(w_asqrt60_6[2]),.din(w_asqrt60_1[2]));
	jspl3 jspl3_w_asqrt60_7(.douta(w_asqrt60_7[0]),.doutb(w_asqrt60_7[1]),.doutc(w_asqrt60_7[2]),.din(w_asqrt60_2[0]));
	jspl3 jspl3_w_asqrt60_8(.douta(w_asqrt60_8[0]),.doutb(w_asqrt60_8[1]),.doutc(w_asqrt60_8[2]),.din(w_asqrt60_2[1]));
	jspl3 jspl3_w_asqrt60_9(.douta(w_asqrt60_9[0]),.doutb(w_asqrt60_9[1]),.doutc(w_asqrt60_9[2]),.din(w_asqrt60_2[2]));
	jspl3 jspl3_w_asqrt60_10(.douta(w_asqrt60_10[0]),.doutb(w_asqrt60_10[1]),.doutc(w_asqrt60_10[2]),.din(w_asqrt60_3[0]));
	jspl3 jspl3_w_asqrt60_11(.douta(w_asqrt60_11[0]),.doutb(w_asqrt60_11[1]),.doutc(w_asqrt60_11[2]),.din(w_asqrt60_3[1]));
	jspl3 jspl3_w_asqrt60_12(.douta(w_asqrt60_12[0]),.doutb(w_asqrt60_12[1]),.doutc(w_asqrt60_12[2]),.din(w_asqrt60_3[2]));
	jspl3 jspl3_w_asqrt60_13(.douta(w_asqrt60_13[0]),.doutb(w_asqrt60_13[1]),.doutc(w_asqrt60_13[2]),.din(w_asqrt60_4[0]));
	jspl3 jspl3_w_asqrt60_14(.douta(w_asqrt60_14[0]),.doutb(w_asqrt60_14[1]),.doutc(w_asqrt60_14[2]),.din(w_asqrt60_4[1]));
	jspl3 jspl3_w_asqrt60_15(.douta(w_asqrt60_15[0]),.doutb(w_asqrt60_15[1]),.doutc(w_asqrt60_15[2]),.din(w_asqrt60_4[2]));
	jspl3 jspl3_w_asqrt60_16(.douta(w_asqrt60_16[0]),.doutb(w_asqrt60_16[1]),.doutc(w_asqrt60_16[2]),.din(w_asqrt60_5[0]));
	jspl3 jspl3_w_asqrt60_17(.douta(w_asqrt60_17[0]),.doutb(w_asqrt60_17[1]),.doutc(w_asqrt60_17[2]),.din(w_asqrt60_5[1]));
	jspl3 jspl3_w_asqrt60_18(.douta(w_asqrt60_18[0]),.doutb(w_asqrt60_18[1]),.doutc(w_asqrt60_18[2]),.din(w_asqrt60_5[2]));
	jspl3 jspl3_w_asqrt60_19(.douta(w_asqrt60_19[0]),.doutb(w_asqrt60_19[1]),.doutc(w_asqrt60_19[2]),.din(w_asqrt60_6[0]));
	jspl3 jspl3_w_asqrt60_20(.douta(w_asqrt60_20[0]),.doutb(w_asqrt60_20[1]),.doutc(w_asqrt60_20[2]),.din(w_asqrt60_6[1]));
	jspl3 jspl3_w_asqrt60_21(.douta(w_asqrt60_21[0]),.doutb(w_asqrt60_21[1]),.doutc(w_asqrt60_21[2]),.din(w_asqrt60_6[2]));
	jspl3 jspl3_w_asqrt60_22(.douta(w_asqrt60_22[0]),.doutb(w_asqrt60_22[1]),.doutc(w_asqrt60_22[2]),.din(w_asqrt60_7[0]));
	jspl3 jspl3_w_asqrt60_23(.douta(w_asqrt60_23[0]),.doutb(w_asqrt60_23[1]),.doutc(w_asqrt60_23[2]),.din(w_asqrt60_7[1]));
	jspl3 jspl3_w_asqrt60_24(.douta(w_asqrt60_24[0]),.doutb(w_asqrt60_24[1]),.doutc(w_asqrt60_24[2]),.din(w_asqrt60_7[2]));
	jspl3 jspl3_w_asqrt60_25(.douta(w_asqrt60_25[0]),.doutb(w_asqrt60_25[1]),.doutc(w_asqrt60_25[2]),.din(w_asqrt60_8[0]));
	jspl3 jspl3_w_asqrt60_26(.douta(w_asqrt60_26[0]),.doutb(w_asqrt60_26[1]),.doutc(w_asqrt60_26[2]),.din(w_asqrt60_8[1]));
	jspl3 jspl3_w_asqrt60_27(.douta(w_asqrt60_27[0]),.doutb(w_asqrt60_27[1]),.doutc(w_asqrt60_27[2]),.din(w_asqrt60_8[2]));
	jspl3 jspl3_w_asqrt60_28(.douta(w_asqrt60_28[0]),.doutb(w_asqrt60_28[1]),.doutc(w_asqrt60_28[2]),.din(w_asqrt60_9[0]));
	jspl3 jspl3_w_asqrt60_29(.douta(w_asqrt60_29[0]),.doutb(w_asqrt60_29[1]),.doutc(w_asqrt60_29[2]),.din(w_asqrt60_9[1]));
	jspl3 jspl3_w_asqrt60_30(.douta(w_asqrt60_30[0]),.doutb(w_asqrt60_30[1]),.doutc(asqrt[59]),.din(w_asqrt60_9[2]));
	jspl3 jspl3_w_asqrt61_0(.douta(w_asqrt61_0[0]),.doutb(w_asqrt61_0[1]),.doutc(w_asqrt61_0[2]),.din(asqrt_fa_61));
	jspl3 jspl3_w_asqrt61_1(.douta(w_asqrt61_1[0]),.doutb(w_asqrt61_1[1]),.doutc(w_asqrt61_1[2]),.din(w_asqrt61_0[0]));
	jspl3 jspl3_w_asqrt61_2(.douta(w_asqrt61_2[0]),.doutb(w_asqrt61_2[1]),.doutc(w_asqrt61_2[2]),.din(w_asqrt61_0[1]));
	jspl3 jspl3_w_asqrt61_3(.douta(w_asqrt61_3[0]),.doutb(w_asqrt61_3[1]),.doutc(w_asqrt61_3[2]),.din(w_asqrt61_0[2]));
	jspl3 jspl3_w_asqrt61_4(.douta(w_asqrt61_4[0]),.doutb(w_asqrt61_4[1]),.doutc(w_asqrt61_4[2]),.din(w_asqrt61_1[0]));
	jspl3 jspl3_w_asqrt61_5(.douta(w_asqrt61_5[0]),.doutb(w_asqrt61_5[1]),.doutc(w_asqrt61_5[2]),.din(w_asqrt61_1[1]));
	jspl3 jspl3_w_asqrt61_6(.douta(w_asqrt61_6[0]),.doutb(w_asqrt61_6[1]),.doutc(w_asqrt61_6[2]),.din(w_asqrt61_1[2]));
	jspl3 jspl3_w_asqrt61_7(.douta(w_asqrt61_7[0]),.doutb(w_asqrt61_7[1]),.doutc(w_asqrt61_7[2]),.din(w_asqrt61_2[0]));
	jspl3 jspl3_w_asqrt61_8(.douta(w_asqrt61_8[0]),.doutb(w_asqrt61_8[1]),.doutc(w_asqrt61_8[2]),.din(w_asqrt61_2[1]));
	jspl3 jspl3_w_asqrt61_9(.douta(w_asqrt61_9[0]),.doutb(w_asqrt61_9[1]),.doutc(w_asqrt61_9[2]),.din(w_asqrt61_2[2]));
	jspl3 jspl3_w_asqrt61_10(.douta(w_asqrt61_10[0]),.doutb(w_asqrt61_10[1]),.doutc(w_asqrt61_10[2]),.din(w_asqrt61_3[0]));
	jspl3 jspl3_w_asqrt61_11(.douta(w_asqrt61_11[0]),.doutb(w_asqrt61_11[1]),.doutc(w_asqrt61_11[2]),.din(w_asqrt61_3[1]));
	jspl3 jspl3_w_asqrt61_12(.douta(w_asqrt61_12[0]),.doutb(w_asqrt61_12[1]),.doutc(w_asqrt61_12[2]),.din(w_asqrt61_3[2]));
	jspl3 jspl3_w_asqrt61_13(.douta(w_asqrt61_13[0]),.doutb(w_asqrt61_13[1]),.doutc(w_asqrt61_13[2]),.din(w_asqrt61_4[0]));
	jspl3 jspl3_w_asqrt61_14(.douta(w_asqrt61_14[0]),.doutb(w_asqrt61_14[1]),.doutc(w_asqrt61_14[2]),.din(w_asqrt61_4[1]));
	jspl3 jspl3_w_asqrt61_15(.douta(w_asqrt61_15[0]),.doutb(w_asqrt61_15[1]),.doutc(w_asqrt61_15[2]),.din(w_asqrt61_4[2]));
	jspl3 jspl3_w_asqrt61_16(.douta(w_asqrt61_16[0]),.doutb(w_asqrt61_16[1]),.doutc(w_asqrt61_16[2]),.din(w_asqrt61_5[0]));
	jspl3 jspl3_w_asqrt61_17(.douta(w_asqrt61_17[0]),.doutb(w_asqrt61_17[1]),.doutc(w_asqrt61_17[2]),.din(w_asqrt61_5[1]));
	jspl3 jspl3_w_asqrt61_18(.douta(w_asqrt61_18[0]),.doutb(w_asqrt61_18[1]),.doutc(w_asqrt61_18[2]),.din(w_asqrt61_5[2]));
	jspl3 jspl3_w_asqrt61_19(.douta(w_asqrt61_19[0]),.doutb(w_asqrt61_19[1]),.doutc(w_asqrt61_19[2]),.din(w_asqrt61_6[0]));
	jspl3 jspl3_w_asqrt61_20(.douta(w_asqrt61_20[0]),.doutb(w_asqrt61_20[1]),.doutc(w_asqrt61_20[2]),.din(w_asqrt61_6[1]));
	jspl3 jspl3_w_asqrt61_21(.douta(w_asqrt61_21[0]),.doutb(w_asqrt61_21[1]),.doutc(w_asqrt61_21[2]),.din(w_asqrt61_6[2]));
	jspl3 jspl3_w_asqrt61_22(.douta(w_asqrt61_22[0]),.doutb(w_asqrt61_22[1]),.doutc(w_asqrt61_22[2]),.din(w_asqrt61_7[0]));
	jspl3 jspl3_w_asqrt61_23(.douta(w_asqrt61_23[0]),.doutb(w_asqrt61_23[1]),.doutc(w_asqrt61_23[2]),.din(w_asqrt61_7[1]));
	jspl3 jspl3_w_asqrt61_24(.douta(w_asqrt61_24[0]),.doutb(w_asqrt61_24[1]),.doutc(w_asqrt61_24[2]),.din(w_asqrt61_7[2]));
	jspl3 jspl3_w_asqrt61_25(.douta(w_asqrt61_25[0]),.doutb(w_asqrt61_25[1]),.doutc(w_asqrt61_25[2]),.din(w_asqrt61_8[0]));
	jspl3 jspl3_w_asqrt61_26(.douta(w_asqrt61_26[0]),.doutb(w_asqrt61_26[1]),.doutc(w_asqrt61_26[2]),.din(w_asqrt61_8[1]));
	jspl3 jspl3_w_asqrt61_27(.douta(w_asqrt61_27[0]),.doutb(w_asqrt61_27[1]),.doutc(w_asqrt61_27[2]),.din(w_asqrt61_8[2]));
	jspl3 jspl3_w_asqrt61_28(.douta(w_asqrt61_28[0]),.doutb(w_asqrt61_28[1]),.doutc(w_asqrt61_28[2]),.din(w_asqrt61_9[0]));
	jspl3 jspl3_w_asqrt61_29(.douta(w_asqrt61_29[0]),.doutb(w_asqrt61_29[1]),.doutc(w_asqrt61_29[2]),.din(w_asqrt61_9[1]));
	jspl3 jspl3_w_asqrt61_30(.douta(w_asqrt61_30[0]),.doutb(w_asqrt61_30[1]),.doutc(w_asqrt61_30[2]),.din(w_asqrt61_9[2]));
	jspl jspl_w_asqrt61_31(.douta(w_asqrt61_31),.doutb(asqrt[60]),.din(w_asqrt61_10[0]));
	jspl3 jspl3_w_asqrt62_0(.douta(w_asqrt62_0[0]),.doutb(w_asqrt62_0[1]),.doutc(w_asqrt62_0[2]),.din(asqrt_fa_62));
	jspl3 jspl3_w_asqrt62_1(.douta(w_asqrt62_1[0]),.doutb(w_asqrt62_1[1]),.doutc(w_asqrt62_1[2]),.din(w_asqrt62_0[0]));
	jspl3 jspl3_w_asqrt62_2(.douta(w_asqrt62_2[0]),.doutb(w_asqrt62_2[1]),.doutc(w_asqrt62_2[2]),.din(w_asqrt62_0[1]));
	jspl3 jspl3_w_asqrt62_3(.douta(w_asqrt62_3[0]),.doutb(w_asqrt62_3[1]),.doutc(w_asqrt62_3[2]),.din(w_asqrt62_0[2]));
	jspl3 jspl3_w_asqrt62_4(.douta(w_asqrt62_4[0]),.doutb(w_asqrt62_4[1]),.doutc(w_asqrt62_4[2]),.din(w_asqrt62_1[0]));
	jspl3 jspl3_w_asqrt62_5(.douta(w_asqrt62_5[0]),.doutb(w_asqrt62_5[1]),.doutc(w_asqrt62_5[2]),.din(w_asqrt62_1[1]));
	jspl3 jspl3_w_asqrt62_6(.douta(w_asqrt62_6[0]),.doutb(w_asqrt62_6[1]),.doutc(w_asqrt62_6[2]),.din(w_asqrt62_1[2]));
	jspl3 jspl3_w_asqrt62_7(.douta(w_asqrt62_7[0]),.doutb(w_asqrt62_7[1]),.doutc(w_asqrt62_7[2]),.din(w_asqrt62_2[0]));
	jspl3 jspl3_w_asqrt62_8(.douta(w_asqrt62_8[0]),.doutb(w_asqrt62_8[1]),.doutc(w_asqrt62_8[2]),.din(w_asqrt62_2[1]));
	jspl3 jspl3_w_asqrt62_9(.douta(w_asqrt62_9[0]),.doutb(w_asqrt62_9[1]),.doutc(w_asqrt62_9[2]),.din(w_asqrt62_2[2]));
	jspl3 jspl3_w_asqrt62_10(.douta(w_asqrt62_10[0]),.doutb(w_asqrt62_10[1]),.doutc(w_asqrt62_10[2]),.din(w_asqrt62_3[0]));
	jspl3 jspl3_w_asqrt62_11(.douta(w_asqrt62_11[0]),.doutb(w_asqrt62_11[1]),.doutc(w_asqrt62_11[2]),.din(w_asqrt62_3[1]));
	jspl3 jspl3_w_asqrt62_12(.douta(w_asqrt62_12[0]),.doutb(w_asqrt62_12[1]),.doutc(w_asqrt62_12[2]),.din(w_asqrt62_3[2]));
	jspl3 jspl3_w_asqrt62_13(.douta(w_asqrt62_13[0]),.doutb(w_asqrt62_13[1]),.doutc(w_asqrt62_13[2]),.din(w_asqrt62_4[0]));
	jspl3 jspl3_w_asqrt62_14(.douta(w_asqrt62_14[0]),.doutb(w_asqrt62_14[1]),.doutc(w_asqrt62_14[2]),.din(w_asqrt62_4[1]));
	jspl3 jspl3_w_asqrt62_15(.douta(w_asqrt62_15[0]),.doutb(w_asqrt62_15[1]),.doutc(w_asqrt62_15[2]),.din(w_asqrt62_4[2]));
	jspl3 jspl3_w_asqrt62_16(.douta(w_asqrt62_16[0]),.doutb(w_asqrt62_16[1]),.doutc(w_asqrt62_16[2]),.din(w_asqrt62_5[0]));
	jspl3 jspl3_w_asqrt62_17(.douta(w_asqrt62_17[0]),.doutb(w_asqrt62_17[1]),.doutc(w_asqrt62_17[2]),.din(w_asqrt62_5[1]));
	jspl3 jspl3_w_asqrt62_18(.douta(w_asqrt62_18[0]),.doutb(w_asqrt62_18[1]),.doutc(w_asqrt62_18[2]),.din(w_asqrt62_5[2]));
	jspl3 jspl3_w_asqrt62_19(.douta(w_asqrt62_19[0]),.doutb(w_asqrt62_19[1]),.doutc(w_asqrt62_19[2]),.din(w_asqrt62_6[0]));
	jspl3 jspl3_w_asqrt62_20(.douta(w_asqrt62_20[0]),.doutb(w_asqrt62_20[1]),.doutc(w_asqrt62_20[2]),.din(w_asqrt62_6[1]));
	jspl3 jspl3_w_asqrt62_21(.douta(w_asqrt62_21[0]),.doutb(w_asqrt62_21[1]),.doutc(w_asqrt62_21[2]),.din(w_asqrt62_6[2]));
	jspl3 jspl3_w_asqrt62_22(.douta(w_asqrt62_22[0]),.doutb(w_asqrt62_22[1]),.doutc(w_asqrt62_22[2]),.din(w_asqrt62_7[0]));
	jspl3 jspl3_w_asqrt62_23(.douta(w_asqrt62_23[0]),.doutb(w_asqrt62_23[1]),.doutc(w_asqrt62_23[2]),.din(w_asqrt62_7[1]));
	jspl3 jspl3_w_asqrt62_24(.douta(w_asqrt62_24[0]),.doutb(w_asqrt62_24[1]),.doutc(w_asqrt62_24[2]),.din(w_asqrt62_7[2]));
	jspl3 jspl3_w_asqrt62_25(.douta(w_asqrt62_25[0]),.doutb(w_asqrt62_25[1]),.doutc(w_asqrt62_25[2]),.din(w_asqrt62_8[0]));
	jspl3 jspl3_w_asqrt62_26(.douta(w_asqrt62_26[0]),.doutb(w_asqrt62_26[1]),.doutc(w_asqrt62_26[2]),.din(w_asqrt62_8[1]));
	jspl3 jspl3_w_asqrt62_27(.douta(w_asqrt62_27[0]),.doutb(w_asqrt62_27[1]),.doutc(w_asqrt62_27[2]),.din(w_asqrt62_8[2]));
	jspl3 jspl3_w_asqrt62_28(.douta(w_asqrt62_28[0]),.doutb(w_asqrt62_28[1]),.doutc(w_asqrt62_28[2]),.din(w_asqrt62_9[0]));
	jspl3 jspl3_w_asqrt62_29(.douta(w_asqrt62_29[0]),.doutb(w_asqrt62_29[1]),.doutc(w_asqrt62_29[2]),.din(w_asqrt62_9[1]));
	jspl3 jspl3_w_asqrt62_30(.douta(w_asqrt62_30[0]),.doutb(w_asqrt62_30[1]),.doutc(w_asqrt62_30[2]),.din(w_asqrt62_9[2]));
	jspl jspl_w_asqrt62_31(.douta(w_asqrt62_31),.doutb(asqrt[61]),.din(w_asqrt62_10[0]));
	jspl3 jspl3_w_asqrt63_0(.douta(w_asqrt63_0[0]),.doutb(w_asqrt63_0[1]),.doutc(w_asqrt63_0[2]),.din(asqrt_fa_63));
	jspl3 jspl3_w_asqrt63_1(.douta(w_asqrt63_1[0]),.doutb(w_asqrt63_1[1]),.doutc(w_asqrt63_1[2]),.din(w_asqrt63_0[0]));
	jspl3 jspl3_w_asqrt63_2(.douta(w_asqrt63_2[0]),.doutb(w_asqrt63_2[1]),.doutc(w_asqrt63_2[2]),.din(w_asqrt63_0[1]));
	jspl3 jspl3_w_asqrt63_3(.douta(w_asqrt63_3[0]),.doutb(w_asqrt63_3[1]),.doutc(w_asqrt63_3[2]),.din(w_asqrt63_0[2]));
	jspl3 jspl3_w_asqrt63_4(.douta(w_asqrt63_4[0]),.doutb(w_asqrt63_4[1]),.doutc(w_asqrt63_4[2]),.din(w_asqrt63_1[0]));
	jspl3 jspl3_w_asqrt63_5(.douta(w_asqrt63_5[0]),.doutb(w_asqrt63_5[1]),.doutc(w_asqrt63_5[2]),.din(w_asqrt63_1[1]));
	jspl3 jspl3_w_asqrt63_6(.douta(w_asqrt63_6[0]),.doutb(w_asqrt63_6[1]),.doutc(w_asqrt63_6[2]),.din(w_asqrt63_1[2]));
	jspl3 jspl3_w_asqrt63_7(.douta(w_asqrt63_7[0]),.doutb(w_asqrt63_7[1]),.doutc(w_asqrt63_7[2]),.din(w_asqrt63_2[0]));
	jspl3 jspl3_w_asqrt63_8(.douta(w_asqrt63_8[0]),.doutb(w_asqrt63_8[1]),.doutc(w_asqrt63_8[2]),.din(w_asqrt63_2[1]));
	jspl3 jspl3_w_asqrt63_9(.douta(w_asqrt63_9[0]),.doutb(w_asqrt63_9[1]),.doutc(w_asqrt63_9[2]),.din(w_asqrt63_2[2]));
	jspl3 jspl3_w_asqrt63_10(.douta(w_asqrt63_10[0]),.doutb(w_asqrt63_10[1]),.doutc(w_asqrt63_10[2]),.din(w_asqrt63_3[0]));
	jspl3 jspl3_w_asqrt63_11(.douta(w_asqrt63_11[0]),.doutb(w_asqrt63_11[1]),.doutc(w_asqrt63_11[2]),.din(w_asqrt63_3[1]));
	jspl3 jspl3_w_asqrt63_12(.douta(w_asqrt63_12[0]),.doutb(w_asqrt63_12[1]),.doutc(w_asqrt63_12[2]),.din(w_asqrt63_3[2]));
	jspl3 jspl3_w_asqrt63_13(.douta(w_asqrt63_13[0]),.doutb(w_asqrt63_13[1]),.doutc(w_asqrt63_13[2]),.din(w_asqrt63_4[0]));
	jspl3 jspl3_w_asqrt63_14(.douta(w_asqrt63_14[0]),.doutb(w_asqrt63_14[1]),.doutc(w_asqrt63_14[2]),.din(w_asqrt63_4[1]));
	jspl3 jspl3_w_asqrt63_15(.douta(w_asqrt63_15[0]),.doutb(w_asqrt63_15[1]),.doutc(w_asqrt63_15[2]),.din(w_asqrt63_4[2]));
	jspl3 jspl3_w_asqrt63_16(.douta(w_asqrt63_16[0]),.doutb(w_asqrt63_16[1]),.doutc(w_asqrt63_16[2]),.din(w_asqrt63_5[0]));
	jspl jspl_w_asqrt63_17(.douta(w_asqrt63_17),.doutb(asqrt[62]),.din(w_asqrt63_5[1]));
	jspl jspl_w_n192_0(.douta(w_n192_0[0]),.doutb(w_n192_0[1]),.din(n192));
	jspl jspl_w_n193_0(.douta(w_n193_0[0]),.doutb(w_n193_0[1]),.din(n193));
	jspl3 jspl3_w_n194_0(.douta(w_n194_0[0]),.doutb(w_n194_0[1]),.doutc(w_n194_0[2]),.din(n194));
	jspl3 jspl3_w_n194_1(.douta(w_n194_1[0]),.doutb(w_n194_1[1]),.doutc(w_n194_1[2]),.din(w_n194_0[0]));
	jspl3 jspl3_w_n194_2(.douta(w_n194_2[0]),.doutb(w_n194_2[1]),.doutc(w_n194_2[2]),.din(w_n194_0[1]));
	jspl3 jspl3_w_n194_3(.douta(w_n194_3[0]),.doutb(w_n194_3[1]),.doutc(w_n194_3[2]),.din(w_n194_0[2]));
	jspl3 jspl3_w_n194_4(.douta(w_n194_4[0]),.doutb(w_n194_4[1]),.doutc(w_n194_4[2]),.din(w_n194_1[0]));
	jspl3 jspl3_w_n194_5(.douta(w_n194_5[0]),.doutb(w_n194_5[1]),.doutc(w_n194_5[2]),.din(w_n194_1[1]));
	jspl3 jspl3_w_n194_6(.douta(w_n194_6[0]),.doutb(w_n194_6[1]),.doutc(w_n194_6[2]),.din(w_n194_1[2]));
	jspl3 jspl3_w_n194_7(.douta(w_n194_7[0]),.doutb(w_n194_7[1]),.doutc(w_n194_7[2]),.din(w_n194_2[0]));
	jspl3 jspl3_w_n194_8(.douta(w_n194_8[0]),.doutb(w_n194_8[1]),.doutc(w_n194_8[2]),.din(w_n194_2[1]));
	jspl3 jspl3_w_n194_9(.douta(w_n194_9[0]),.doutb(w_n194_9[1]),.doutc(w_n194_9[2]),.din(w_n194_2[2]));
	jspl3 jspl3_w_n194_10(.douta(w_n194_10[0]),.doutb(w_n194_10[1]),.doutc(w_n194_10[2]),.din(w_n194_3[0]));
	jspl3 jspl3_w_n194_11(.douta(w_n194_11[0]),.doutb(w_n194_11[1]),.doutc(w_n194_11[2]),.din(w_n194_3[1]));
	jspl3 jspl3_w_n194_12(.douta(w_n194_12[0]),.doutb(w_n194_12[1]),.doutc(w_n194_12[2]),.din(w_n194_3[2]));
	jspl3 jspl3_w_n194_13(.douta(w_n194_13[0]),.doutb(w_n194_13[1]),.doutc(w_n194_13[2]),.din(w_n194_4[0]));
	jspl3 jspl3_w_n194_14(.douta(w_n194_14[0]),.doutb(w_n194_14[1]),.doutc(w_n194_14[2]),.din(w_n194_4[1]));
	jspl3 jspl3_w_n194_15(.douta(w_n194_15[0]),.doutb(w_n194_15[1]),.doutc(w_n194_15[2]),.din(w_n194_4[2]));
	jspl3 jspl3_w_n194_16(.douta(w_n194_16[0]),.doutb(w_n194_16[1]),.doutc(w_n194_16[2]),.din(w_n194_5[0]));
	jspl3 jspl3_w_n194_17(.douta(w_n194_17[0]),.doutb(w_n194_17[1]),.doutc(w_n194_17[2]),.din(w_n194_5[1]));
	jspl3 jspl3_w_n194_18(.douta(w_n194_18[0]),.doutb(w_n194_18[1]),.doutc(w_n194_18[2]),.din(w_n194_5[2]));
	jspl3 jspl3_w_n194_19(.douta(w_n194_19[0]),.doutb(w_n194_19[1]),.doutc(w_n194_19[2]),.din(w_n194_6[0]));
	jspl3 jspl3_w_n194_20(.douta(w_n194_20[0]),.doutb(w_n194_20[1]),.doutc(w_n194_20[2]),.din(w_n194_6[1]));
	jspl3 jspl3_w_n194_21(.douta(w_n194_21[0]),.doutb(w_n194_21[1]),.doutc(w_n194_21[2]),.din(w_n194_6[2]));
	jspl3 jspl3_w_n194_22(.douta(w_n194_22[0]),.doutb(w_n194_22[1]),.doutc(w_n194_22[2]),.din(w_n194_7[0]));
	jspl3 jspl3_w_n194_23(.douta(w_n194_23[0]),.doutb(w_n194_23[1]),.doutc(w_n194_23[2]),.din(w_n194_7[1]));
	jspl3 jspl3_w_n194_24(.douta(w_n194_24[0]),.doutb(w_n194_24[1]),.doutc(w_n194_24[2]),.din(w_n194_7[2]));
	jspl3 jspl3_w_n194_25(.douta(w_n194_25[0]),.doutb(w_n194_25[1]),.doutc(w_n194_25[2]),.din(w_n194_8[0]));
	jspl3 jspl3_w_n194_26(.douta(w_n194_26[0]),.doutb(w_n194_26[1]),.doutc(w_n194_26[2]),.din(w_n194_8[1]));
	jspl3 jspl3_w_n194_27(.douta(w_n194_27[0]),.doutb(w_n194_27[1]),.doutc(w_n194_27[2]),.din(w_n194_8[2]));
	jspl3 jspl3_w_n194_28(.douta(w_n194_28[0]),.doutb(w_n194_28[1]),.doutc(w_n194_28[2]),.din(w_n194_9[0]));
	jspl3 jspl3_w_n194_29(.douta(w_n194_29[0]),.doutb(w_n194_29[1]),.doutc(w_n194_29[2]),.din(w_n194_9[1]));
	jspl3 jspl3_w_n194_30(.douta(w_n194_30[0]),.doutb(w_n194_30[1]),.doutc(w_n194_30[2]),.din(w_n194_9[2]));
	jspl3 jspl3_w_n194_31(.douta(w_n194_31[0]),.doutb(w_n194_31[1]),.doutc(w_n194_31[2]),.din(w_n194_10[0]));
	jspl3 jspl3_w_n194_32(.douta(w_n194_32[0]),.doutb(w_n194_32[1]),.doutc(w_n194_32[2]),.din(w_n194_10[1]));
	jspl3 jspl3_w_n194_33(.douta(w_n194_33[0]),.doutb(w_n194_33[1]),.doutc(w_n194_33[2]),.din(w_n194_10[2]));
	jspl3 jspl3_w_n194_34(.douta(w_n194_34[0]),.doutb(w_n194_34[1]),.doutc(w_n194_34[2]),.din(w_n194_11[0]));
	jspl3 jspl3_w_n194_35(.douta(w_n194_35[0]),.doutb(w_n194_35[1]),.doutc(w_n194_35[2]),.din(w_n194_11[1]));
	jspl3 jspl3_w_n194_36(.douta(w_n194_36[0]),.doutb(w_n194_36[1]),.doutc(w_n194_36[2]),.din(w_n194_11[2]));
	jspl3 jspl3_w_n194_37(.douta(w_n194_37[0]),.doutb(w_n194_37[1]),.doutc(w_n194_37[2]),.din(w_n194_12[0]));
	jspl3 jspl3_w_n194_38(.douta(w_n194_38[0]),.doutb(w_n194_38[1]),.doutc(w_n194_38[2]),.din(w_n194_12[1]));
	jspl3 jspl3_w_n194_39(.douta(w_n194_39[0]),.doutb(w_n194_39[1]),.doutc(w_n194_39[2]),.din(w_n194_12[2]));
	jspl3 jspl3_w_n194_40(.douta(w_n194_40[0]),.doutb(w_n194_40[1]),.doutc(w_n194_40[2]),.din(w_n194_13[0]));
	jspl3 jspl3_w_n194_41(.douta(w_n194_41[0]),.doutb(w_n194_41[1]),.doutc(w_n194_41[2]),.din(w_n194_13[1]));
	jspl3 jspl3_w_n194_42(.douta(w_n194_42[0]),.doutb(w_n194_42[1]),.doutc(w_n194_42[2]),.din(w_n194_13[2]));
	jspl3 jspl3_w_n194_43(.douta(w_n194_43[0]),.doutb(w_n194_43[1]),.doutc(w_n194_43[2]),.din(w_n194_14[0]));
	jspl jspl_w_n195_0(.douta(w_n195_0[0]),.doutb(w_n195_0[1]),.din(n195));
	jspl jspl_w_n196_0(.douta(w_n196_0[0]),.doutb(w_n196_0[1]),.din(n196));
	jspl jspl_w_n197_0(.douta(w_n197_0[0]),.doutb(w_n197_0[1]),.din(n197));
	jspl3 jspl3_w_n199_0(.douta(w_n199_0[0]),.doutb(w_n199_0[1]),.doutc(w_n199_0[2]),.din(n199));
	jspl3 jspl3_w_n199_1(.douta(w_n199_1[0]),.doutb(w_n199_1[1]),.doutc(w_n199_1[2]),.din(w_n199_0[0]));
	jspl3 jspl3_w_n199_2(.douta(w_n199_2[0]),.doutb(w_n199_2[1]),.doutc(w_n199_2[2]),.din(w_n199_0[1]));
	jspl3 jspl3_w_n199_3(.douta(w_n199_3[0]),.doutb(w_n199_3[1]),.doutc(w_n199_3[2]),.din(w_n199_0[2]));
	jspl3 jspl3_w_n199_4(.douta(w_n199_4[0]),.doutb(w_n199_4[1]),.doutc(w_n199_4[2]),.din(w_n199_1[0]));
	jspl3 jspl3_w_n199_5(.douta(w_n199_5[0]),.doutb(w_n199_5[1]),.doutc(w_n199_5[2]),.din(w_n199_1[1]));
	jspl3 jspl3_w_n199_6(.douta(w_n199_6[0]),.doutb(w_n199_6[1]),.doutc(w_n199_6[2]),.din(w_n199_1[2]));
	jspl3 jspl3_w_n199_7(.douta(w_n199_7[0]),.doutb(w_n199_7[1]),.doutc(w_n199_7[2]),.din(w_n199_2[0]));
	jspl3 jspl3_w_n199_8(.douta(w_n199_8[0]),.doutb(w_n199_8[1]),.doutc(w_n199_8[2]),.din(w_n199_2[1]));
	jspl3 jspl3_w_n199_9(.douta(w_n199_9[0]),.doutb(w_n199_9[1]),.doutc(w_n199_9[2]),.din(w_n199_2[2]));
	jspl3 jspl3_w_n199_10(.douta(w_n199_10[0]),.doutb(w_n199_10[1]),.doutc(w_n199_10[2]),.din(w_n199_3[0]));
	jspl3 jspl3_w_n199_11(.douta(w_n199_11[0]),.doutb(w_n199_11[1]),.doutc(w_n199_11[2]),.din(w_n199_3[1]));
	jspl3 jspl3_w_n199_12(.douta(w_n199_12[0]),.doutb(w_n199_12[1]),.doutc(w_n199_12[2]),.din(w_n199_3[2]));
	jspl3 jspl3_w_n199_13(.douta(w_n199_13[0]),.doutb(w_n199_13[1]),.doutc(w_n199_13[2]),.din(w_n199_4[0]));
	jspl3 jspl3_w_n199_14(.douta(w_n199_14[0]),.doutb(w_n199_14[1]),.doutc(w_n199_14[2]),.din(w_n199_4[1]));
	jspl3 jspl3_w_n199_15(.douta(w_n199_15[0]),.doutb(w_n199_15[1]),.doutc(w_n199_15[2]),.din(w_n199_4[2]));
	jspl3 jspl3_w_n199_16(.douta(w_n199_16[0]),.doutb(w_n199_16[1]),.doutc(w_n199_16[2]),.din(w_n199_5[0]));
	jspl3 jspl3_w_n199_17(.douta(w_n199_17[0]),.doutb(w_n199_17[1]),.doutc(w_n199_17[2]),.din(w_n199_5[1]));
	jspl3 jspl3_w_n199_18(.douta(w_n199_18[0]),.doutb(w_n199_18[1]),.doutc(w_n199_18[2]),.din(w_n199_5[2]));
	jspl3 jspl3_w_n199_19(.douta(w_n199_19[0]),.doutb(w_n199_19[1]),.doutc(w_n199_19[2]),.din(w_n199_6[0]));
	jspl3 jspl3_w_n199_20(.douta(w_n199_20[0]),.doutb(w_n199_20[1]),.doutc(w_n199_20[2]),.din(w_n199_6[1]));
	jspl3 jspl3_w_n199_21(.douta(w_n199_21[0]),.doutb(w_n199_21[1]),.doutc(w_n199_21[2]),.din(w_n199_6[2]));
	jspl3 jspl3_w_n199_22(.douta(w_n199_22[0]),.doutb(w_n199_22[1]),.doutc(w_n199_22[2]),.din(w_n199_7[0]));
	jspl3 jspl3_w_n199_23(.douta(w_n199_23[0]),.doutb(w_n199_23[1]),.doutc(w_n199_23[2]),.din(w_n199_7[1]));
	jspl3 jspl3_w_n199_24(.douta(w_n199_24[0]),.doutb(w_n199_24[1]),.doutc(w_n199_24[2]),.din(w_n199_7[2]));
	jspl3 jspl3_w_n199_25(.douta(w_n199_25[0]),.doutb(w_n199_25[1]),.doutc(w_n199_25[2]),.din(w_n199_8[0]));
	jspl3 jspl3_w_n199_26(.douta(w_n199_26[0]),.doutb(w_n199_26[1]),.doutc(w_n199_26[2]),.din(w_n199_8[1]));
	jspl3 jspl3_w_n199_27(.douta(w_n199_27[0]),.doutb(w_n199_27[1]),.doutc(w_n199_27[2]),.din(w_n199_8[2]));
	jspl3 jspl3_w_n199_28(.douta(w_n199_28[0]),.doutb(w_n199_28[1]),.doutc(w_n199_28[2]),.din(w_n199_9[0]));
	jspl3 jspl3_w_n199_29(.douta(w_n199_29[0]),.doutb(w_n199_29[1]),.doutc(w_n199_29[2]),.din(w_n199_9[1]));
	jspl3 jspl3_w_n199_30(.douta(w_n199_30[0]),.doutb(w_n199_30[1]),.doutc(w_n199_30[2]),.din(w_n199_9[2]));
	jspl3 jspl3_w_n199_31(.douta(w_n199_31[0]),.doutb(w_n199_31[1]),.doutc(w_n199_31[2]),.din(w_n199_10[0]));
	jspl3 jspl3_w_n199_32(.douta(w_n199_32[0]),.doutb(w_n199_32[1]),.doutc(w_n199_32[2]),.din(w_n199_10[1]));
	jspl3 jspl3_w_n199_33(.douta(w_n199_33[0]),.doutb(w_n199_33[1]),.doutc(w_n199_33[2]),.din(w_n199_10[2]));
	jspl3 jspl3_w_n199_34(.douta(w_n199_34[0]),.doutb(w_n199_34[1]),.doutc(w_n199_34[2]),.din(w_n199_11[0]));
	jspl3 jspl3_w_n199_35(.douta(w_n199_35[0]),.doutb(w_n199_35[1]),.doutc(w_n199_35[2]),.din(w_n199_11[1]));
	jspl3 jspl3_w_n199_36(.douta(w_n199_36[0]),.doutb(w_n199_36[1]),.doutc(w_n199_36[2]),.din(w_n199_11[2]));
	jspl3 jspl3_w_n199_37(.douta(w_n199_37[0]),.doutb(w_n199_37[1]),.doutc(w_n199_37[2]),.din(w_n199_12[0]));
	jspl3 jspl3_w_n199_38(.douta(w_n199_38[0]),.doutb(w_n199_38[1]),.doutc(w_n199_38[2]),.din(w_n199_12[1]));
	jspl3 jspl3_w_n199_39(.douta(w_n199_39[0]),.doutb(w_n199_39[1]),.doutc(w_n199_39[2]),.din(w_n199_12[2]));
	jspl3 jspl3_w_n199_40(.douta(w_n199_40[0]),.doutb(w_n199_40[1]),.doutc(w_n199_40[2]),.din(w_n199_13[0]));
	jspl3 jspl3_w_n199_41(.douta(w_n199_41[0]),.doutb(w_n199_41[1]),.doutc(w_n199_41[2]),.din(w_n199_13[1]));
	jspl3 jspl3_w_n199_42(.douta(w_n199_42[0]),.doutb(w_n199_42[1]),.doutc(w_n199_42[2]),.din(w_n199_13[2]));
	jspl3 jspl3_w_n199_43(.douta(w_n199_43[0]),.doutb(w_n199_43[1]),.doutc(w_n199_43[2]),.din(w_n199_14[0]));
	jspl3 jspl3_w_n199_44(.douta(w_n199_44[0]),.doutb(w_n199_44[1]),.doutc(w_n199_44[2]),.din(w_n199_14[1]));
	jspl3 jspl3_w_n199_45(.douta(w_n199_45[0]),.doutb(w_n199_45[1]),.doutc(w_n199_45[2]),.din(w_n199_14[2]));
	jspl jspl_w_n200_0(.douta(w_n200_0[0]),.doutb(w_n200_0[1]),.din(n200));
	jspl3 jspl3_w_n203_0(.douta(w_n203_0[0]),.doutb(w_n203_0[1]),.doutc(w_n203_0[2]),.din(n203));
	jspl jspl_w_n206_0(.douta(w_n206_0[0]),.doutb(w_n206_0[1]),.din(n206));
	jspl3 jspl3_w_n209_0(.douta(w_n209_0[0]),.doutb(w_n209_0[1]),.doutc(w_n209_0[2]),.din(n209));
	jspl3 jspl3_w_n211_0(.douta(w_n211_0[0]),.doutb(w_n211_0[1]),.doutc(w_n211_0[2]),.din(n211));
	jspl jspl_w_n211_1(.douta(w_n211_1[0]),.doutb(w_n211_1[1]),.din(w_n211_0[0]));
	jspl jspl_w_n212_0(.douta(w_n212_0[0]),.doutb(w_n212_0[1]),.din(n212));
	jspl3 jspl3_w_n215_0(.douta(w_n215_0[0]),.doutb(w_n215_0[1]),.doutc(w_n215_0[2]),.din(n215));
	jspl3 jspl3_w_n216_0(.douta(w_n216_0[0]),.doutb(w_n216_0[1]),.doutc(w_n216_0[2]),.din(n216));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.din(n218));
	jspl jspl_w_n221_0(.douta(w_n221_0[0]),.doutb(w_n221_0[1]),.din(n221));
	jspl3 jspl3_w_n223_0(.douta(w_n223_0[0]),.doutb(w_n223_0[1]),.doutc(w_n223_0[2]),.din(n223));
	jspl3 jspl3_w_n223_1(.douta(w_n223_1[0]),.doutb(w_n223_1[1]),.doutc(w_n223_1[2]),.din(w_n223_0[0]));
	jspl3 jspl3_w_n223_2(.douta(w_n223_2[0]),.doutb(w_n223_2[1]),.doutc(w_n223_2[2]),.din(w_n223_0[1]));
	jspl3 jspl3_w_n223_3(.douta(w_n223_3[0]),.doutb(w_n223_3[1]),.doutc(w_n223_3[2]),.din(w_n223_0[2]));
	jspl3 jspl3_w_n223_4(.douta(w_n223_4[0]),.doutb(w_n223_4[1]),.doutc(w_n223_4[2]),.din(w_n223_1[0]));
	jspl3 jspl3_w_n223_5(.douta(w_n223_5[0]),.doutb(w_n223_5[1]),.doutc(w_n223_5[2]),.din(w_n223_1[1]));
	jspl3 jspl3_w_n223_6(.douta(w_n223_6[0]),.doutb(w_n223_6[1]),.doutc(w_n223_6[2]),.din(w_n223_1[2]));
	jspl3 jspl3_w_n223_7(.douta(w_n223_7[0]),.doutb(w_n223_7[1]),.doutc(w_n223_7[2]),.din(w_n223_2[0]));
	jspl3 jspl3_w_n223_8(.douta(w_n223_8[0]),.doutb(w_n223_8[1]),.doutc(w_n223_8[2]),.din(w_n223_2[1]));
	jspl3 jspl3_w_n223_9(.douta(w_n223_9[0]),.doutb(w_n223_9[1]),.doutc(w_n223_9[2]),.din(w_n223_2[2]));
	jspl3 jspl3_w_n223_10(.douta(w_n223_10[0]),.doutb(w_n223_10[1]),.doutc(w_n223_10[2]),.din(w_n223_3[0]));
	jspl3 jspl3_w_n223_11(.douta(w_n223_11[0]),.doutb(w_n223_11[1]),.doutc(w_n223_11[2]),.din(w_n223_3[1]));
	jspl3 jspl3_w_n223_12(.douta(w_n223_12[0]),.doutb(w_n223_12[1]),.doutc(w_n223_12[2]),.din(w_n223_3[2]));
	jspl3 jspl3_w_n223_13(.douta(w_n223_13[0]),.doutb(w_n223_13[1]),.doutc(w_n223_13[2]),.din(w_n223_4[0]));
	jspl3 jspl3_w_n223_14(.douta(w_n223_14[0]),.doutb(w_n223_14[1]),.doutc(w_n223_14[2]),.din(w_n223_4[1]));
	jspl3 jspl3_w_n223_15(.douta(w_n223_15[0]),.doutb(w_n223_15[1]),.doutc(w_n223_15[2]),.din(w_n223_4[2]));
	jspl3 jspl3_w_n223_16(.douta(w_n223_16[0]),.doutb(w_n223_16[1]),.doutc(w_n223_16[2]),.din(w_n223_5[0]));
	jspl3 jspl3_w_n223_17(.douta(w_n223_17[0]),.doutb(w_n223_17[1]),.doutc(w_n223_17[2]),.din(w_n223_5[1]));
	jspl3 jspl3_w_n223_18(.douta(w_n223_18[0]),.doutb(w_n223_18[1]),.doutc(w_n223_18[2]),.din(w_n223_5[2]));
	jspl3 jspl3_w_n223_19(.douta(w_n223_19[0]),.doutb(w_n223_19[1]),.doutc(w_n223_19[2]),.din(w_n223_6[0]));
	jspl3 jspl3_w_n223_20(.douta(w_n223_20[0]),.doutb(w_n223_20[1]),.doutc(w_n223_20[2]),.din(w_n223_6[1]));
	jspl3 jspl3_w_n223_21(.douta(w_n223_21[0]),.doutb(w_n223_21[1]),.doutc(w_n223_21[2]),.din(w_n223_6[2]));
	jspl3 jspl3_w_n223_22(.douta(w_n223_22[0]),.doutb(w_n223_22[1]),.doutc(w_n223_22[2]),.din(w_n223_7[0]));
	jspl3 jspl3_w_n223_23(.douta(w_n223_23[0]),.doutb(w_n223_23[1]),.doutc(w_n223_23[2]),.din(w_n223_7[1]));
	jspl3 jspl3_w_n223_24(.douta(w_n223_24[0]),.doutb(w_n223_24[1]),.doutc(w_n223_24[2]),.din(w_n223_7[2]));
	jspl3 jspl3_w_n223_25(.douta(w_n223_25[0]),.doutb(w_n223_25[1]),.doutc(w_n223_25[2]),.din(w_n223_8[0]));
	jspl3 jspl3_w_n223_26(.douta(w_n223_26[0]),.doutb(w_n223_26[1]),.doutc(w_n223_26[2]),.din(w_n223_8[1]));
	jspl3 jspl3_w_n223_27(.douta(w_n223_27[0]),.doutb(w_n223_27[1]),.doutc(w_n223_27[2]),.din(w_n223_8[2]));
	jspl3 jspl3_w_n223_28(.douta(w_n223_28[0]),.doutb(w_n223_28[1]),.doutc(w_n223_28[2]),.din(w_n223_9[0]));
	jspl3 jspl3_w_n223_29(.douta(w_n223_29[0]),.doutb(w_n223_29[1]),.doutc(w_n223_29[2]),.din(w_n223_9[1]));
	jspl3 jspl3_w_n223_30(.douta(w_n223_30[0]),.doutb(w_n223_30[1]),.doutc(w_n223_30[2]),.din(w_n223_9[2]));
	jspl3 jspl3_w_n223_31(.douta(w_n223_31[0]),.doutb(w_n223_31[1]),.doutc(w_n223_31[2]),.din(w_n223_10[0]));
	jspl3 jspl3_w_n223_32(.douta(w_n223_32[0]),.doutb(w_n223_32[1]),.doutc(w_n223_32[2]),.din(w_n223_10[1]));
	jspl3 jspl3_w_n223_33(.douta(w_n223_33[0]),.doutb(w_n223_33[1]),.doutc(w_n223_33[2]),.din(w_n223_10[2]));
	jspl3 jspl3_w_n223_34(.douta(w_n223_34[0]),.doutb(w_n223_34[1]),.doutc(w_n223_34[2]),.din(w_n223_11[0]));
	jspl3 jspl3_w_n223_35(.douta(w_n223_35[0]),.doutb(w_n223_35[1]),.doutc(w_n223_35[2]),.din(w_n223_11[1]));
	jspl3 jspl3_w_n223_36(.douta(w_n223_36[0]),.doutb(w_n223_36[1]),.doutc(w_n223_36[2]),.din(w_n223_11[2]));
	jspl3 jspl3_w_n223_37(.douta(w_n223_37[0]),.doutb(w_n223_37[1]),.doutc(w_n223_37[2]),.din(w_n223_12[0]));
	jspl3 jspl3_w_n223_38(.douta(w_n223_38[0]),.doutb(w_n223_38[1]),.doutc(w_n223_38[2]),.din(w_n223_12[1]));
	jspl3 jspl3_w_n223_39(.douta(w_n223_39[0]),.doutb(w_n223_39[1]),.doutc(w_n223_39[2]),.din(w_n223_12[2]));
	jspl jspl_w_n226_0(.douta(w_n226_0[0]),.doutb(w_n226_0[1]),.din(n226));
	jspl3 jspl3_w_n229_0(.douta(w_n229_0[0]),.doutb(w_n229_0[1]),.doutc(w_n229_0[2]),.din(n229));
	jspl3 jspl3_w_n231_0(.douta(w_n231_0[0]),.doutb(w_n231_0[1]),.doutc(w_n231_0[2]),.din(n231));
	jspl jspl_w_n231_1(.douta(w_n231_1[0]),.doutb(w_n231_1[1]),.din(w_n231_0[0]));
	jspl3 jspl3_w_n232_0(.douta(w_n232_0[0]),.doutb(w_n232_0[1]),.doutc(w_n232_0[2]),.din(n232));
	jspl3 jspl3_w_n236_0(.douta(w_n236_0[0]),.doutb(w_n236_0[1]),.doutc(w_n236_0[2]),.din(n236));
	jspl jspl_w_n239_0(.douta(w_n239_0[0]),.doutb(w_n239_0[1]),.din(n239));
	jspl jspl_w_n241_0(.douta(w_n241_0[0]),.doutb(w_n241_0[1]),.din(n241));
	jspl3 jspl3_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.doutc(w_n242_0[2]),.din(n242));
	jspl jspl_w_n248_0(.douta(w_n248_0[0]),.doutb(w_n248_0[1]),.din(n248));
	jspl jspl_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.din(n249));
	jspl jspl_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.din(n254));
	jspl3 jspl3_w_n261_0(.douta(w_n261_0[0]),.doutb(w_n261_0[1]),.doutc(w_n261_0[2]),.din(n261));
	jspl jspl_w_n261_1(.douta(w_n261_1[0]),.doutb(w_n261_1[1]),.din(w_n261_0[0]));
	jspl jspl_w_n262_0(.douta(w_n262_0[0]),.doutb(w_n262_0[1]),.din(n262));
	jspl3 jspl3_w_n265_0(.douta(w_n265_0[0]),.doutb(w_n265_0[1]),.doutc(w_n265_0[2]),.din(n265));
	jspl jspl_w_n266_0(.douta(w_n266_0[0]),.doutb(w_n266_0[1]),.din(n266));
	jspl jspl_w_n267_0(.douta(w_n267_0[0]),.doutb(w_n267_0[1]),.din(n267));
	jspl jspl_w_n268_0(.douta(w_n268_0[0]),.doutb(w_n268_0[1]),.din(n268));
	jspl jspl_w_n270_0(.douta(w_n270_0[0]),.doutb(w_n270_0[1]),.din(n270));
	jspl jspl_w_n272_0(.douta(w_n272_0[0]),.doutb(w_n272_0[1]),.din(n272));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_n274_0[1]),.din(n274));
	jspl3 jspl3_w_n277_0(.douta(w_n277_0[0]),.doutb(w_n277_0[1]),.doutc(w_n277_0[2]),.din(n277));
	jspl jspl_w_n283_0(.douta(w_n283_0[0]),.doutb(w_n283_0[1]),.din(n283));
	jspl3 jspl3_w_n285_0(.douta(w_n285_0[0]),.doutb(w_n285_0[1]),.doutc(w_n285_0[2]),.din(n285));
	jspl jspl_w_n285_1(.douta(w_n285_1[0]),.doutb(w_n285_1[1]),.din(w_n285_0[0]));
	jspl3 jspl3_w_n289_0(.douta(w_n289_0[0]),.doutb(w_n289_0[1]),.doutc(w_n289_0[2]),.din(n289));
	jspl jspl_w_n289_1(.douta(w_n289_1[0]),.doutb(w_n289_1[1]),.din(w_n289_0[0]));
	jspl3 jspl3_w_n290_0(.douta(w_n290_0[0]),.doutb(w_n290_0[1]),.doutc(w_n290_0[2]),.din(n290));
	jspl3 jspl3_w_n290_1(.douta(w_n290_1[0]),.doutb(w_n290_1[1]),.doutc(w_n290_1[2]),.din(w_n290_0[0]));
	jspl3 jspl3_w_n290_2(.douta(w_n290_2[0]),.doutb(w_n290_2[1]),.doutc(w_n290_2[2]),.din(w_n290_0[1]));
	jspl3 jspl3_w_n290_3(.douta(w_n290_3[0]),.doutb(w_n290_3[1]),.doutc(w_n290_3[2]),.din(w_n290_0[2]));
	jspl3 jspl3_w_n290_4(.douta(w_n290_4[0]),.doutb(w_n290_4[1]),.doutc(w_n290_4[2]),.din(w_n290_1[0]));
	jspl3 jspl3_w_n290_5(.douta(w_n290_5[0]),.doutb(w_n290_5[1]),.doutc(w_n290_5[2]),.din(w_n290_1[1]));
	jspl3 jspl3_w_n290_6(.douta(w_n290_6[0]),.doutb(w_n290_6[1]),.doutc(w_n290_6[2]),.din(w_n290_1[2]));
	jspl3 jspl3_w_n290_7(.douta(w_n290_7[0]),.doutb(w_n290_7[1]),.doutc(w_n290_7[2]),.din(w_n290_2[0]));
	jspl3 jspl3_w_n290_8(.douta(w_n290_8[0]),.doutb(w_n290_8[1]),.doutc(w_n290_8[2]),.din(w_n290_2[1]));
	jspl3 jspl3_w_n290_9(.douta(w_n290_9[0]),.doutb(w_n290_9[1]),.doutc(w_n290_9[2]),.din(w_n290_2[2]));
	jspl3 jspl3_w_n290_10(.douta(w_n290_10[0]),.doutb(w_n290_10[1]),.doutc(w_n290_10[2]),.din(w_n290_3[0]));
	jspl3 jspl3_w_n290_11(.douta(w_n290_11[0]),.doutb(w_n290_11[1]),.doutc(w_n290_11[2]),.din(w_n290_3[1]));
	jspl3 jspl3_w_n290_12(.douta(w_n290_12[0]),.doutb(w_n290_12[1]),.doutc(w_n290_12[2]),.din(w_n290_3[2]));
	jspl3 jspl3_w_n290_13(.douta(w_n290_13[0]),.doutb(w_n290_13[1]),.doutc(w_n290_13[2]),.din(w_n290_4[0]));
	jspl3 jspl3_w_n290_14(.douta(w_n290_14[0]),.doutb(w_n290_14[1]),.doutc(w_n290_14[2]),.din(w_n290_4[1]));
	jspl3 jspl3_w_n290_15(.douta(w_n290_15[0]),.doutb(w_n290_15[1]),.doutc(w_n290_15[2]),.din(w_n290_4[2]));
	jspl3 jspl3_w_n290_16(.douta(w_n290_16[0]),.doutb(w_n290_16[1]),.doutc(w_n290_16[2]),.din(w_n290_5[0]));
	jspl3 jspl3_w_n290_17(.douta(w_n290_17[0]),.doutb(w_n290_17[1]),.doutc(w_n290_17[2]),.din(w_n290_5[1]));
	jspl3 jspl3_w_n290_18(.douta(w_n290_18[0]),.doutb(w_n290_18[1]),.doutc(w_n290_18[2]),.din(w_n290_5[2]));
	jspl3 jspl3_w_n290_19(.douta(w_n290_19[0]),.doutb(w_n290_19[1]),.doutc(w_n290_19[2]),.din(w_n290_6[0]));
	jspl3 jspl3_w_n290_20(.douta(w_n290_20[0]),.doutb(w_n290_20[1]),.doutc(w_n290_20[2]),.din(w_n290_6[1]));
	jspl3 jspl3_w_n290_21(.douta(w_n290_21[0]),.doutb(w_n290_21[1]),.doutc(w_n290_21[2]),.din(w_n290_6[2]));
	jspl3 jspl3_w_n290_22(.douta(w_n290_22[0]),.doutb(w_n290_22[1]),.doutc(w_n290_22[2]),.din(w_n290_7[0]));
	jspl3 jspl3_w_n290_23(.douta(w_n290_23[0]),.doutb(w_n290_23[1]),.doutc(w_n290_23[2]),.din(w_n290_7[1]));
	jspl3 jspl3_w_n290_24(.douta(w_n290_24[0]),.doutb(w_n290_24[1]),.doutc(w_n290_24[2]),.din(w_n290_7[2]));
	jspl3 jspl3_w_n290_25(.douta(w_n290_25[0]),.doutb(w_n290_25[1]),.doutc(w_n290_25[2]),.din(w_n290_8[0]));
	jspl3 jspl3_w_n290_26(.douta(w_n290_26[0]),.doutb(w_n290_26[1]),.doutc(w_n290_26[2]),.din(w_n290_8[1]));
	jspl3 jspl3_w_n290_27(.douta(w_n290_27[0]),.doutb(w_n290_27[1]),.doutc(w_n290_27[2]),.din(w_n290_8[2]));
	jspl3 jspl3_w_n290_28(.douta(w_n290_28[0]),.doutb(w_n290_28[1]),.doutc(w_n290_28[2]),.din(w_n290_9[0]));
	jspl3 jspl3_w_n290_29(.douta(w_n290_29[0]),.doutb(w_n290_29[1]),.doutc(w_n290_29[2]),.din(w_n290_9[1]));
	jspl3 jspl3_w_n290_30(.douta(w_n290_30[0]),.doutb(w_n290_30[1]),.doutc(w_n290_30[2]),.din(w_n290_9[2]));
	jspl3 jspl3_w_n290_31(.douta(w_n290_31[0]),.doutb(w_n290_31[1]),.doutc(w_n290_31[2]),.din(w_n290_10[0]));
	jspl3 jspl3_w_n290_32(.douta(w_n290_32[0]),.doutb(w_n290_32[1]),.doutc(w_n290_32[2]),.din(w_n290_10[1]));
	jspl3 jspl3_w_n290_33(.douta(w_n290_33[0]),.doutb(w_n290_33[1]),.doutc(w_n290_33[2]),.din(w_n290_10[2]));
	jspl3 jspl3_w_n290_34(.douta(w_n290_34[0]),.doutb(w_n290_34[1]),.doutc(w_n290_34[2]),.din(w_n290_11[0]));
	jspl3 jspl3_w_n290_35(.douta(w_n290_35[0]),.doutb(w_n290_35[1]),.doutc(w_n290_35[2]),.din(w_n290_11[1]));
	jspl3 jspl3_w_n290_36(.douta(w_n290_36[0]),.doutb(w_n290_36[1]),.doutc(w_n290_36[2]),.din(w_n290_11[2]));
	jspl3 jspl3_w_n290_37(.douta(w_n290_37[0]),.doutb(w_n290_37[1]),.doutc(w_n290_37[2]),.din(w_n290_12[0]));
	jspl3 jspl3_w_n290_38(.douta(w_n290_38[0]),.doutb(w_n290_38[1]),.doutc(w_n290_38[2]),.din(w_n290_12[1]));
	jspl jspl_w_n290_39(.douta(w_n290_39[0]),.doutb(w_n290_39[1]),.din(w_n290_12[2]));
	jspl jspl_w_n295_0(.douta(w_n295_0[0]),.doutb(w_n295_0[1]),.din(n295));
	jspl3 jspl3_w_n296_0(.douta(w_n296_0[0]),.doutb(w_n296_0[1]),.doutc(w_n296_0[2]),.din(n296));
	jspl jspl_w_n301_0(.douta(w_n301_0[0]),.doutb(w_n301_0[1]),.din(n301));
	jspl3 jspl3_w_n305_0(.douta(w_n305_0[0]),.doutb(w_n305_0[1]),.doutc(w_n305_0[2]),.din(n305));
	jspl3 jspl3_w_n305_1(.douta(w_n305_1[0]),.doutb(w_n305_1[1]),.doutc(w_n305_1[2]),.din(w_n305_0[0]));
	jspl3 jspl3_w_n305_2(.douta(w_n305_2[0]),.doutb(w_n305_2[1]),.doutc(w_n305_2[2]),.din(w_n305_0[1]));
	jspl3 jspl3_w_n305_3(.douta(w_n305_3[0]),.doutb(w_n305_3[1]),.doutc(w_n305_3[2]),.din(w_n305_0[2]));
	jspl3 jspl3_w_n305_4(.douta(w_n305_4[0]),.doutb(w_n305_4[1]),.doutc(w_n305_4[2]),.din(w_n305_1[0]));
	jspl3 jspl3_w_n305_5(.douta(w_n305_5[0]),.doutb(w_n305_5[1]),.doutc(w_n305_5[2]),.din(w_n305_1[1]));
	jspl3 jspl3_w_n305_6(.douta(w_n305_6[0]),.doutb(w_n305_6[1]),.doutc(w_n305_6[2]),.din(w_n305_1[2]));
	jspl3 jspl3_w_n305_7(.douta(w_n305_7[0]),.doutb(w_n305_7[1]),.doutc(w_n305_7[2]),.din(w_n305_2[0]));
	jspl3 jspl3_w_n305_8(.douta(w_n305_8[0]),.doutb(w_n305_8[1]),.doutc(w_n305_8[2]),.din(w_n305_2[1]));
	jspl3 jspl3_w_n305_9(.douta(w_n305_9[0]),.doutb(w_n305_9[1]),.doutc(w_n305_9[2]),.din(w_n305_2[2]));
	jspl3 jspl3_w_n305_10(.douta(w_n305_10[0]),.doutb(w_n305_10[1]),.doutc(w_n305_10[2]),.din(w_n305_3[0]));
	jspl3 jspl3_w_n305_11(.douta(w_n305_11[0]),.doutb(w_n305_11[1]),.doutc(w_n305_11[2]),.din(w_n305_3[1]));
	jspl3 jspl3_w_n305_12(.douta(w_n305_12[0]),.doutb(w_n305_12[1]),.doutc(w_n305_12[2]),.din(w_n305_3[2]));
	jspl3 jspl3_w_n305_13(.douta(w_n305_13[0]),.doutb(w_n305_13[1]),.doutc(w_n305_13[2]),.din(w_n305_4[0]));
	jspl3 jspl3_w_n305_14(.douta(w_n305_14[0]),.doutb(w_n305_14[1]),.doutc(w_n305_14[2]),.din(w_n305_4[1]));
	jspl3 jspl3_w_n305_15(.douta(w_n305_15[0]),.doutb(w_n305_15[1]),.doutc(w_n305_15[2]),.din(w_n305_4[2]));
	jspl3 jspl3_w_n305_16(.douta(w_n305_16[0]),.doutb(w_n305_16[1]),.doutc(w_n305_16[2]),.din(w_n305_5[0]));
	jspl3 jspl3_w_n305_17(.douta(w_n305_17[0]),.doutb(w_n305_17[1]),.doutc(w_n305_17[2]),.din(w_n305_5[1]));
	jspl3 jspl3_w_n305_18(.douta(w_n305_18[0]),.doutb(w_n305_18[1]),.doutc(w_n305_18[2]),.din(w_n305_5[2]));
	jspl3 jspl3_w_n305_19(.douta(w_n305_19[0]),.doutb(w_n305_19[1]),.doutc(w_n305_19[2]),.din(w_n305_6[0]));
	jspl3 jspl3_w_n305_20(.douta(w_n305_20[0]),.doutb(w_n305_20[1]),.doutc(w_n305_20[2]),.din(w_n305_6[1]));
	jspl3 jspl3_w_n305_21(.douta(w_n305_21[0]),.doutb(w_n305_21[1]),.doutc(w_n305_21[2]),.din(w_n305_6[2]));
	jspl3 jspl3_w_n305_22(.douta(w_n305_22[0]),.doutb(w_n305_22[1]),.doutc(w_n305_22[2]),.din(w_n305_7[0]));
	jspl3 jspl3_w_n305_23(.douta(w_n305_23[0]),.doutb(w_n305_23[1]),.doutc(w_n305_23[2]),.din(w_n305_7[1]));
	jspl3 jspl3_w_n305_24(.douta(w_n305_24[0]),.doutb(w_n305_24[1]),.doutc(w_n305_24[2]),.din(w_n305_7[2]));
	jspl3 jspl3_w_n305_25(.douta(w_n305_25[0]),.doutb(w_n305_25[1]),.doutc(w_n305_25[2]),.din(w_n305_8[0]));
	jspl3 jspl3_w_n305_26(.douta(w_n305_26[0]),.doutb(w_n305_26[1]),.doutc(w_n305_26[2]),.din(w_n305_8[1]));
	jspl3 jspl3_w_n305_27(.douta(w_n305_27[0]),.doutb(w_n305_27[1]),.doutc(w_n305_27[2]),.din(w_n305_8[2]));
	jspl3 jspl3_w_n305_28(.douta(w_n305_28[0]),.doutb(w_n305_28[1]),.doutc(w_n305_28[2]),.din(w_n305_9[0]));
	jspl3 jspl3_w_n305_29(.douta(w_n305_29[0]),.doutb(w_n305_29[1]),.doutc(w_n305_29[2]),.din(w_n305_9[1]));
	jspl3 jspl3_w_n305_30(.douta(w_n305_30[0]),.doutb(w_n305_30[1]),.doutc(w_n305_30[2]),.din(w_n305_9[2]));
	jspl3 jspl3_w_n305_31(.douta(w_n305_31[0]),.doutb(w_n305_31[1]),.doutc(w_n305_31[2]),.din(w_n305_10[0]));
	jspl3 jspl3_w_n305_32(.douta(w_n305_32[0]),.doutb(w_n305_32[1]),.doutc(w_n305_32[2]),.din(w_n305_10[1]));
	jspl3 jspl3_w_n305_33(.douta(w_n305_33[0]),.doutb(w_n305_33[1]),.doutc(w_n305_33[2]),.din(w_n305_10[2]));
	jspl3 jspl3_w_n305_34(.douta(w_n305_34[0]),.doutb(w_n305_34[1]),.doutc(w_n305_34[2]),.din(w_n305_11[0]));
	jspl3 jspl3_w_n305_35(.douta(w_n305_35[0]),.doutb(w_n305_35[1]),.doutc(w_n305_35[2]),.din(w_n305_11[1]));
	jspl3 jspl3_w_n305_36(.douta(w_n305_36[0]),.doutb(w_n305_36[1]),.doutc(w_n305_36[2]),.din(w_n305_11[2]));
	jspl3 jspl3_w_n305_37(.douta(w_n305_37[0]),.doutb(w_n305_37[1]),.doutc(w_n305_37[2]),.din(w_n305_12[0]));
	jspl3 jspl3_w_n305_38(.douta(w_n305_38[0]),.doutb(w_n305_38[1]),.doutc(w_n305_38[2]),.din(w_n305_12[1]));
	jspl3 jspl3_w_n305_39(.douta(w_n305_39[0]),.doutb(w_n305_39[1]),.doutc(w_n305_39[2]),.din(w_n305_12[2]));
	jspl3 jspl3_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.doutc(w_n308_0[2]),.din(n308));
	jspl jspl_w_n308_1(.douta(w_n308_1[0]),.doutb(w_n308_1[1]),.din(w_n308_0[0]));
	jspl3 jspl3_w_n309_0(.douta(w_n309_0[0]),.doutb(w_n309_0[1]),.doutc(w_n309_0[2]),.din(n309));
	jspl3 jspl3_w_n313_0(.douta(w_n313_0[0]),.doutb(w_n313_0[1]),.doutc(w_n313_0[2]),.din(n313));
	jspl jspl_w_n314_0(.douta(w_n314_0[0]),.doutb(w_n314_0[1]),.din(n314));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl jspl_w_n316_0(.douta(w_n316_0[0]),.doutb(w_n316_0[1]),.din(n316));
	jspl jspl_w_n318_0(.douta(w_n318_0[0]),.doutb(w_n318_0[1]),.din(n318));
	jspl jspl_w_n320_0(.douta(w_n320_0[0]),.doutb(w_n320_0[1]),.din(n320));
	jspl jspl_w_n322_0(.douta(w_n322_0[0]),.doutb(w_n322_0[1]),.din(n322));
	jspl jspl_w_n325_0(.douta(w_n325_0[0]),.doutb(w_n325_0[1]),.din(n325));
	jspl jspl_w_n329_0(.douta(w_n329_0[0]),.doutb(w_n329_0[1]),.din(n329));
	jspl3 jspl3_w_n331_0(.douta(w_n331_0[0]),.doutb(w_n331_0[1]),.doutc(w_n331_0[2]),.din(n331));
	jspl jspl_w_n336_0(.douta(w_n336_0[0]),.doutb(w_n336_0[1]),.din(n336));
	jspl3 jspl3_w_n338_0(.douta(w_n338_0[0]),.doutb(w_n338_0[1]),.doutc(w_n338_0[2]),.din(n338));
	jspl3 jspl3_w_n342_0(.douta(w_n342_0[0]),.doutb(w_n342_0[1]),.doutc(w_n342_0[2]),.din(n342));
	jspl jspl_w_n348_0(.douta(w_n348_0[0]),.doutb(w_n348_0[1]),.din(n348));
	jspl3 jspl3_w_n349_0(.douta(w_n349_0[0]),.doutb(w_n349_0[1]),.doutc(w_n349_0[2]),.din(n349));
	jspl jspl_w_n358_0(.douta(w_n358_0[0]),.doutb(w_n358_0[1]),.din(n358));
	jspl3 jspl3_w_n363_0(.douta(w_n363_0[0]),.doutb(w_n363_0[1]),.doutc(w_n363_0[2]),.din(n363));
	jspl jspl_w_n363_1(.douta(w_n363_1[0]),.doutb(w_n363_1[1]),.din(w_n363_0[0]));
	jspl jspl_w_n364_0(.douta(w_n364_0[0]),.doutb(w_n364_0[1]),.din(n364));
	jspl3 jspl3_w_n367_0(.douta(w_n367_0[0]),.doutb(w_n367_0[1]),.doutc(w_n367_0[2]),.din(n367));
	jspl jspl_w_n368_0(.douta(w_n368_0[0]),.doutb(w_n368_0[1]),.din(n368));
	jspl jspl_w_n369_0(.douta(w_n369_0[0]),.doutb(w_n369_0[1]),.din(n369));
	jspl jspl_w_n370_0(.douta(w_n370_0[0]),.doutb(w_n370_0[1]),.din(n370));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.din(n372));
	jspl jspl_w_n374_0(.douta(w_n374_0[0]),.doutb(w_n374_0[1]),.din(n374));
	jspl jspl_w_n376_0(.douta(w_n376_0[0]),.doutb(w_n376_0[1]),.din(n376));
	jspl jspl_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.din(n385));
	jspl3 jspl3_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.doutc(w_n387_0[2]),.din(n387));
	jspl jspl_w_n388_0(.douta(w_n388_0[0]),.doutb(w_n388_0[1]),.din(n388));
	jspl jspl_w_n392_0(.douta(w_n392_0[0]),.doutb(w_n392_0[1]),.din(n392));
	jspl jspl_w_n394_0(.douta(w_n394_0[0]),.doutb(w_n394_0[1]),.din(n394));
	jspl jspl_w_n396_0(.douta(w_n396_0[0]),.doutb(w_n396_0[1]),.din(n396));
	jspl jspl_w_n401_0(.douta(w_n401_0[0]),.doutb(w_n401_0[1]),.din(n401));
	jspl jspl_w_n403_0(.douta(w_n403_0[0]),.doutb(w_n403_0[1]),.din(n403));
	jspl jspl_w_n404_0(.douta(w_n404_0[0]),.doutb(w_n404_0[1]),.din(n404));
	jspl3 jspl3_w_n405_0(.douta(w_n405_0[0]),.doutb(w_n405_0[1]),.doutc(w_n405_0[2]),.din(n405));
	jspl3 jspl3_w_n405_1(.douta(w_n405_1[0]),.doutb(w_n405_1[1]),.doutc(w_n405_1[2]),.din(w_n405_0[0]));
	jspl jspl_w_n408_0(.douta(w_n408_0[0]),.doutb(w_n408_0[1]),.din(n408));
	jspl3 jspl3_w_n409_0(.douta(w_n409_0[0]),.doutb(w_n409_0[1]),.doutc(w_n409_0[2]),.din(n409));
	jspl jspl_w_n410_0(.douta(w_n410_0[0]),.doutb(w_n410_0[1]),.din(n410));
	jspl jspl_w_n411_0(.douta(w_n411_0[0]),.doutb(w_n411_0[1]),.din(n411));
	jspl jspl_w_n417_0(.douta(w_n417_0[0]),.doutb(w_n417_0[1]),.din(n417));
	jspl3 jspl3_w_n418_0(.douta(w_n418_0[0]),.doutb(w_n418_0[1]),.doutc(w_n418_0[2]),.din(n418));
	jspl jspl_w_n419_0(.douta(w_n419_0[0]),.doutb(w_n419_0[1]),.din(n419));
	jspl jspl_w_n424_0(.douta(w_n424_0[0]),.doutb(w_n424_0[1]),.din(n424));
	jspl3 jspl3_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.doutc(w_n425_0[2]),.din(n425));
	jspl3 jspl3_w_n425_1(.douta(w_n425_1[0]),.doutb(w_n425_1[1]),.doutc(w_n425_1[2]),.din(w_n425_0[0]));
	jspl3 jspl3_w_n425_2(.douta(w_n425_2[0]),.doutb(w_n425_2[1]),.doutc(w_n425_2[2]),.din(w_n425_0[1]));
	jspl3 jspl3_w_n425_3(.douta(w_n425_3[0]),.doutb(w_n425_3[1]),.doutc(w_n425_3[2]),.din(w_n425_0[2]));
	jspl3 jspl3_w_n425_4(.douta(w_n425_4[0]),.doutb(w_n425_4[1]),.doutc(w_n425_4[2]),.din(w_n425_1[0]));
	jspl3 jspl3_w_n425_5(.douta(w_n425_5[0]),.doutb(w_n425_5[1]),.doutc(w_n425_5[2]),.din(w_n425_1[1]));
	jspl3 jspl3_w_n425_6(.douta(w_n425_6[0]),.doutb(w_n425_6[1]),.doutc(w_n425_6[2]),.din(w_n425_1[2]));
	jspl3 jspl3_w_n425_7(.douta(w_n425_7[0]),.doutb(w_n425_7[1]),.doutc(w_n425_7[2]),.din(w_n425_2[0]));
	jspl3 jspl3_w_n425_8(.douta(w_n425_8[0]),.doutb(w_n425_8[1]),.doutc(w_n425_8[2]),.din(w_n425_2[1]));
	jspl3 jspl3_w_n425_9(.douta(w_n425_9[0]),.doutb(w_n425_9[1]),.doutc(w_n425_9[2]),.din(w_n425_2[2]));
	jspl3 jspl3_w_n425_10(.douta(w_n425_10[0]),.doutb(w_n425_10[1]),.doutc(w_n425_10[2]),.din(w_n425_3[0]));
	jspl3 jspl3_w_n425_11(.douta(w_n425_11[0]),.doutb(w_n425_11[1]),.doutc(w_n425_11[2]),.din(w_n425_3[1]));
	jspl3 jspl3_w_n425_12(.douta(w_n425_12[0]),.doutb(w_n425_12[1]),.doutc(w_n425_12[2]),.din(w_n425_3[2]));
	jspl3 jspl3_w_n425_13(.douta(w_n425_13[0]),.doutb(w_n425_13[1]),.doutc(w_n425_13[2]),.din(w_n425_4[0]));
	jspl3 jspl3_w_n425_14(.douta(w_n425_14[0]),.doutb(w_n425_14[1]),.doutc(w_n425_14[2]),.din(w_n425_4[1]));
	jspl3 jspl3_w_n425_15(.douta(w_n425_15[0]),.doutb(w_n425_15[1]),.doutc(w_n425_15[2]),.din(w_n425_4[2]));
	jspl3 jspl3_w_n425_16(.douta(w_n425_16[0]),.doutb(w_n425_16[1]),.doutc(w_n425_16[2]),.din(w_n425_5[0]));
	jspl3 jspl3_w_n425_17(.douta(w_n425_17[0]),.doutb(w_n425_17[1]),.doutc(w_n425_17[2]),.din(w_n425_5[1]));
	jspl3 jspl3_w_n425_18(.douta(w_n425_18[0]),.doutb(w_n425_18[1]),.doutc(w_n425_18[2]),.din(w_n425_5[2]));
	jspl3 jspl3_w_n425_19(.douta(w_n425_19[0]),.doutb(w_n425_19[1]),.doutc(w_n425_19[2]),.din(w_n425_6[0]));
	jspl3 jspl3_w_n425_20(.douta(w_n425_20[0]),.doutb(w_n425_20[1]),.doutc(w_n425_20[2]),.din(w_n425_6[1]));
	jspl3 jspl3_w_n425_21(.douta(w_n425_21[0]),.doutb(w_n425_21[1]),.doutc(w_n425_21[2]),.din(w_n425_6[2]));
	jspl3 jspl3_w_n425_22(.douta(w_n425_22[0]),.doutb(w_n425_22[1]),.doutc(w_n425_22[2]),.din(w_n425_7[0]));
	jspl3 jspl3_w_n425_23(.douta(w_n425_23[0]),.doutb(w_n425_23[1]),.doutc(w_n425_23[2]),.din(w_n425_7[1]));
	jspl3 jspl3_w_n425_24(.douta(w_n425_24[0]),.doutb(w_n425_24[1]),.doutc(w_n425_24[2]),.din(w_n425_7[2]));
	jspl3 jspl3_w_n425_25(.douta(w_n425_25[0]),.doutb(w_n425_25[1]),.doutc(w_n425_25[2]),.din(w_n425_8[0]));
	jspl3 jspl3_w_n425_26(.douta(w_n425_26[0]),.doutb(w_n425_26[1]),.doutc(w_n425_26[2]),.din(w_n425_8[1]));
	jspl3 jspl3_w_n425_27(.douta(w_n425_27[0]),.doutb(w_n425_27[1]),.doutc(w_n425_27[2]),.din(w_n425_8[2]));
	jspl3 jspl3_w_n425_28(.douta(w_n425_28[0]),.doutb(w_n425_28[1]),.doutc(w_n425_28[2]),.din(w_n425_9[0]));
	jspl3 jspl3_w_n425_29(.douta(w_n425_29[0]),.doutb(w_n425_29[1]),.doutc(w_n425_29[2]),.din(w_n425_9[1]));
	jspl3 jspl3_w_n425_30(.douta(w_n425_30[0]),.doutb(w_n425_30[1]),.doutc(w_n425_30[2]),.din(w_n425_9[2]));
	jspl3 jspl3_w_n425_31(.douta(w_n425_31[0]),.doutb(w_n425_31[1]),.doutc(w_n425_31[2]),.din(w_n425_10[0]));
	jspl3 jspl3_w_n425_32(.douta(w_n425_32[0]),.doutb(w_n425_32[1]),.doutc(w_n425_32[2]),.din(w_n425_10[1]));
	jspl3 jspl3_w_n425_33(.douta(w_n425_33[0]),.doutb(w_n425_33[1]),.doutc(w_n425_33[2]),.din(w_n425_10[2]));
	jspl3 jspl3_w_n425_34(.douta(w_n425_34[0]),.doutb(w_n425_34[1]),.doutc(w_n425_34[2]),.din(w_n425_11[0]));
	jspl3 jspl3_w_n425_35(.douta(w_n425_35[0]),.doutb(w_n425_35[1]),.doutc(w_n425_35[2]),.din(w_n425_11[1]));
	jspl3 jspl3_w_n425_36(.douta(w_n425_36[0]),.doutb(w_n425_36[1]),.doutc(w_n425_36[2]),.din(w_n425_11[2]));
	jspl3 jspl3_w_n430_0(.douta(w_n430_0[0]),.doutb(w_n430_0[1]),.doutc(w_n430_0[2]),.din(n430));
	jspl3 jspl3_w_n430_1(.douta(w_n430_1[0]),.doutb(w_n430_1[1]),.doutc(w_n430_1[2]),.din(w_n430_0[0]));
	jspl3 jspl3_w_n430_2(.douta(w_n430_2[0]),.doutb(w_n430_2[1]),.doutc(w_n430_2[2]),.din(w_n430_0[1]));
	jspl3 jspl3_w_n430_3(.douta(w_n430_3[0]),.doutb(w_n430_3[1]),.doutc(w_n430_3[2]),.din(w_n430_0[2]));
	jspl3 jspl3_w_n430_4(.douta(w_n430_4[0]),.doutb(w_n430_4[1]),.doutc(w_n430_4[2]),.din(w_n430_1[0]));
	jspl3 jspl3_w_n430_5(.douta(w_n430_5[0]),.doutb(w_n430_5[1]),.doutc(w_n430_5[2]),.din(w_n430_1[1]));
	jspl3 jspl3_w_n430_6(.douta(w_n430_6[0]),.doutb(w_n430_6[1]),.doutc(w_n430_6[2]),.din(w_n430_1[2]));
	jspl3 jspl3_w_n430_7(.douta(w_n430_7[0]),.doutb(w_n430_7[1]),.doutc(w_n430_7[2]),.din(w_n430_2[0]));
	jspl3 jspl3_w_n430_8(.douta(w_n430_8[0]),.doutb(w_n430_8[1]),.doutc(w_n430_8[2]),.din(w_n430_2[1]));
	jspl3 jspl3_w_n430_9(.douta(w_n430_9[0]),.doutb(w_n430_9[1]),.doutc(w_n430_9[2]),.din(w_n430_2[2]));
	jspl3 jspl3_w_n430_10(.douta(w_n430_10[0]),.doutb(w_n430_10[1]),.doutc(w_n430_10[2]),.din(w_n430_3[0]));
	jspl3 jspl3_w_n430_11(.douta(w_n430_11[0]),.doutb(w_n430_11[1]),.doutc(w_n430_11[2]),.din(w_n430_3[1]));
	jspl3 jspl3_w_n430_12(.douta(w_n430_12[0]),.doutb(w_n430_12[1]),.doutc(w_n430_12[2]),.din(w_n430_3[2]));
	jspl3 jspl3_w_n430_13(.douta(w_n430_13[0]),.doutb(w_n430_13[1]),.doutc(w_n430_13[2]),.din(w_n430_4[0]));
	jspl3 jspl3_w_n430_14(.douta(w_n430_14[0]),.doutb(w_n430_14[1]),.doutc(w_n430_14[2]),.din(w_n430_4[1]));
	jspl3 jspl3_w_n430_15(.douta(w_n430_15[0]),.doutb(w_n430_15[1]),.doutc(w_n430_15[2]),.din(w_n430_4[2]));
	jspl3 jspl3_w_n430_16(.douta(w_n430_16[0]),.doutb(w_n430_16[1]),.doutc(w_n430_16[2]),.din(w_n430_5[0]));
	jspl3 jspl3_w_n430_17(.douta(w_n430_17[0]),.doutb(w_n430_17[1]),.doutc(w_n430_17[2]),.din(w_n430_5[1]));
	jspl3 jspl3_w_n430_18(.douta(w_n430_18[0]),.doutb(w_n430_18[1]),.doutc(w_n430_18[2]),.din(w_n430_5[2]));
	jspl3 jspl3_w_n430_19(.douta(w_n430_19[0]),.doutb(w_n430_19[1]),.doutc(w_n430_19[2]),.din(w_n430_6[0]));
	jspl3 jspl3_w_n430_20(.douta(w_n430_20[0]),.doutb(w_n430_20[1]),.doutc(w_n430_20[2]),.din(w_n430_6[1]));
	jspl3 jspl3_w_n430_21(.douta(w_n430_21[0]),.doutb(w_n430_21[1]),.doutc(w_n430_21[2]),.din(w_n430_6[2]));
	jspl3 jspl3_w_n430_22(.douta(w_n430_22[0]),.doutb(w_n430_22[1]),.doutc(w_n430_22[2]),.din(w_n430_7[0]));
	jspl3 jspl3_w_n430_23(.douta(w_n430_23[0]),.doutb(w_n430_23[1]),.doutc(w_n430_23[2]),.din(w_n430_7[1]));
	jspl3 jspl3_w_n430_24(.douta(w_n430_24[0]),.doutb(w_n430_24[1]),.doutc(w_n430_24[2]),.din(w_n430_7[2]));
	jspl3 jspl3_w_n430_25(.douta(w_n430_25[0]),.doutb(w_n430_25[1]),.doutc(w_n430_25[2]),.din(w_n430_8[0]));
	jspl3 jspl3_w_n430_26(.douta(w_n430_26[0]),.doutb(w_n430_26[1]),.doutc(w_n430_26[2]),.din(w_n430_8[1]));
	jspl3 jspl3_w_n430_27(.douta(w_n430_27[0]),.doutb(w_n430_27[1]),.doutc(w_n430_27[2]),.din(w_n430_8[2]));
	jspl3 jspl3_w_n430_28(.douta(w_n430_28[0]),.doutb(w_n430_28[1]),.doutc(w_n430_28[2]),.din(w_n430_9[0]));
	jspl3 jspl3_w_n430_29(.douta(w_n430_29[0]),.doutb(w_n430_29[1]),.doutc(w_n430_29[2]),.din(w_n430_9[1]));
	jspl3 jspl3_w_n430_30(.douta(w_n430_30[0]),.doutb(w_n430_30[1]),.doutc(w_n430_30[2]),.din(w_n430_9[2]));
	jspl3 jspl3_w_n430_31(.douta(w_n430_31[0]),.doutb(w_n430_31[1]),.doutc(w_n430_31[2]),.din(w_n430_10[0]));
	jspl3 jspl3_w_n430_32(.douta(w_n430_32[0]),.doutb(w_n430_32[1]),.doutc(w_n430_32[2]),.din(w_n430_10[1]));
	jspl3 jspl3_w_n430_33(.douta(w_n430_33[0]),.doutb(w_n430_33[1]),.doutc(w_n430_33[2]),.din(w_n430_10[2]));
	jspl3 jspl3_w_n430_34(.douta(w_n430_34[0]),.doutb(w_n430_34[1]),.doutc(w_n430_34[2]),.din(w_n430_11[0]));
	jspl3 jspl3_w_n430_35(.douta(w_n430_35[0]),.doutb(w_n430_35[1]),.doutc(w_n430_35[2]),.din(w_n430_11[1]));
	jspl3 jspl3_w_n430_36(.douta(w_n430_36[0]),.doutb(w_n430_36[1]),.doutc(w_n430_36[2]),.din(w_n430_11[2]));
	jspl3 jspl3_w_n430_37(.douta(w_n430_37[0]),.doutb(w_n430_37[1]),.doutc(w_n430_37[2]),.din(w_n430_12[0]));
	jspl3 jspl3_w_n430_38(.douta(w_n430_38[0]),.doutb(w_n430_38[1]),.doutc(w_n430_38[2]),.din(w_n430_12[1]));
	jspl3 jspl3_w_n433_0(.douta(w_n433_0[0]),.doutb(w_n433_0[1]),.doutc(w_n433_0[2]),.din(n433));
	jspl jspl_w_n433_1(.douta(w_n433_1[0]),.doutb(w_n433_1[1]),.din(w_n433_0[0]));
	jspl3 jspl3_w_n434_0(.douta(w_n434_0[0]),.doutb(w_n434_0[1]),.doutc(w_n434_0[2]),.din(n434));
	jspl3 jspl3_w_n438_0(.douta(w_n438_0[0]),.doutb(w_n438_0[1]),.doutc(w_n438_0[2]),.din(n438));
	jspl jspl_w_n439_0(.douta(w_n439_0[0]),.doutb(w_n439_0[1]),.din(n439));
	jspl jspl_w_n440_0(.douta(w_n440_0[0]),.doutb(w_n440_0[1]),.din(n440));
	jspl jspl_w_n441_0(.douta(w_n441_0[0]),.doutb(w_n441_0[1]),.din(n441));
	jspl jspl_w_n443_0(.douta(w_n443_0[0]),.doutb(w_n443_0[1]),.din(n443));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl jspl_w_n447_0(.douta(w_n447_0[0]),.doutb(w_n447_0[1]),.din(n447));
	jspl jspl_w_n450_0(.douta(w_n450_0[0]),.doutb(w_n450_0[1]),.din(n450));
	jspl jspl_w_n455_0(.douta(w_n455_0[0]),.doutb(w_n455_0[1]),.din(n455));
	jspl3 jspl3_w_n457_0(.douta(w_n457_0[0]),.doutb(w_n457_0[1]),.doutc(w_n457_0[2]),.din(n457));
	jspl jspl_w_n458_0(.douta(w_n458_0[0]),.doutb(w_n458_0[1]),.din(n458));
	jspl jspl_w_n462_0(.douta(w_n462_0[0]),.doutb(w_n462_0[1]),.din(n462));
	jspl jspl_w_n463_0(.douta(w_n463_0[0]),.doutb(w_n463_0[1]),.din(n463));
	jspl jspl_w_n465_0(.douta(w_n465_0[0]),.doutb(w_n465_0[1]),.din(n465));
	jspl jspl_w_n469_0(.douta(w_n469_0[0]),.doutb(w_n469_0[1]),.din(n469));
	jspl jspl_w_n471_0(.douta(w_n471_0[0]),.doutb(w_n471_0[1]),.din(n471));
	jspl jspl_w_n472_0(.douta(w_n472_0[0]),.doutb(w_n472_0[1]),.din(n472));
	jspl3 jspl3_w_n473_0(.douta(w_n473_0[0]),.doutb(w_n473_0[1]),.doutc(w_n473_0[2]),.din(n473));
	jspl jspl_w_n478_0(.douta(w_n478_0[0]),.doutb(w_n478_0[1]),.din(n478));
	jspl3 jspl3_w_n481_0(.douta(w_n481_0[0]),.doutb(w_n481_0[1]),.doutc(w_n481_0[2]),.din(n481));
	jspl jspl_w_n483_0(.douta(w_n483_0[0]),.doutb(w_n483_0[1]),.din(n483));
	jspl3 jspl3_w_n488_0(.douta(w_n488_0[0]),.doutb(w_n488_0[1]),.doutc(w_n488_0[2]),.din(n488));
	jspl jspl_w_n489_0(.douta(w_n489_0[0]),.doutb(w_n489_0[1]),.din(n489));
	jspl jspl_w_n490_0(.douta(w_n490_0[0]),.doutb(w_n490_0[1]),.din(n490));
	jspl jspl_w_n495_0(.douta(w_n495_0[0]),.doutb(w_n495_0[1]),.din(n495));
	jspl3 jspl3_w_n496_0(.douta(w_n496_0[0]),.doutb(w_n496_0[1]),.doutc(w_n496_0[2]),.din(n496));
	jspl jspl_w_n501_0(.douta(w_n501_0[0]),.doutb(w_n501_0[1]),.din(n501));
	jspl3 jspl3_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.doutc(w_n507_0[2]),.din(n507));
	jspl jspl_w_n507_1(.douta(w_n507_1[0]),.doutb(w_n507_1[1]),.din(w_n507_0[0]));
	jspl jspl_w_n508_0(.douta(w_n508_0[0]),.doutb(w_n508_0[1]),.din(n508));
	jspl3 jspl3_w_n511_0(.douta(w_n511_0[0]),.doutb(w_n511_0[1]),.doutc(w_n511_0[2]),.din(n511));
	jspl jspl_w_n512_0(.douta(w_n512_0[0]),.doutb(w_n512_0[1]),.din(n512));
	jspl jspl_w_n513_0(.douta(w_n513_0[0]),.doutb(w_n513_0[1]),.din(n513));
	jspl jspl_w_n514_0(.douta(w_n514_0[0]),.doutb(w_n514_0[1]),.din(n514));
	jspl jspl_w_n516_0(.douta(w_n516_0[0]),.doutb(w_n516_0[1]),.din(n516));
	jspl jspl_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.din(n518));
	jspl jspl_w_n520_0(.douta(w_n520_0[0]),.doutb(w_n520_0[1]),.din(n520));
	jspl jspl_w_n529_0(.douta(w_n529_0[0]),.doutb(w_n529_0[1]),.din(n529));
	jspl3 jspl3_w_n531_0(.douta(w_n531_0[0]),.doutb(w_n531_0[1]),.doutc(w_n531_0[2]),.din(n531));
	jspl jspl_w_n532_0(.douta(w_n532_0[0]),.doutb(w_n532_0[1]),.din(n532));
	jspl jspl_w_n536_0(.douta(w_n536_0[0]),.doutb(w_n536_0[1]),.din(n536));
	jspl jspl_w_n538_0(.douta(w_n538_0[0]),.doutb(w_n538_0[1]),.din(n538));
	jspl jspl_w_n540_0(.douta(w_n540_0[0]),.doutb(w_n540_0[1]),.din(n540));
	jspl jspl_w_n545_0(.douta(w_n545_0[0]),.doutb(w_n545_0[1]),.din(n545));
	jspl jspl_w_n547_0(.douta(w_n547_0[0]),.doutb(w_n547_0[1]),.din(n547));
	jspl jspl_w_n548_0(.douta(w_n548_0[0]),.doutb(w_n548_0[1]),.din(n548));
	jspl3 jspl3_w_n549_0(.douta(w_n549_0[0]),.doutb(w_n549_0[1]),.doutc(w_n549_0[2]),.din(n549));
	jspl jspl_w_n550_0(.douta(w_n550_0[0]),.doutb(w_n550_0[1]),.din(n550));
	jspl jspl_w_n555_0(.douta(w_n555_0[0]),.doutb(w_n555_0[1]),.din(n555));
	jspl jspl_w_n556_0(.douta(w_n556_0[0]),.doutb(w_n556_0[1]),.din(n556));
	jspl jspl_w_n558_0(.douta(w_n558_0[0]),.doutb(w_n558_0[1]),.din(n558));
	jspl jspl_w_n560_0(.douta(w_n560_0[0]),.doutb(w_n560_0[1]),.din(n560));
	jspl jspl_w_n563_0(.douta(w_n563_0[0]),.doutb(w_n563_0[1]),.din(n563));
	jspl jspl_w_n569_0(.douta(w_n569_0[0]),.doutb(w_n569_0[1]),.din(n569));
	jspl3 jspl3_w_n571_0(.douta(w_n571_0[0]),.doutb(w_n571_0[1]),.doutc(w_n571_0[2]),.din(n571));
	jspl3 jspl3_w_n571_1(.douta(w_n571_1[0]),.doutb(w_n571_1[1]),.doutc(w_n571_1[2]),.din(w_n571_0[0]));
	jspl3 jspl3_w_n574_0(.douta(w_n574_0[0]),.doutb(w_n574_0[1]),.doutc(w_n574_0[2]),.din(n574));
	jspl jspl_w_n574_1(.douta(w_n574_1[0]),.doutb(w_n574_1[1]),.din(w_n574_0[0]));
	jspl3 jspl3_w_n576_0(.douta(w_n576_0[0]),.doutb(w_n576_0[1]),.doutc(w_n576_0[2]),.din(n576));
	jspl jspl_w_n577_0(.douta(w_n577_0[0]),.doutb(w_n577_0[1]),.din(n577));
	jspl jspl_w_n583_0(.douta(w_n583_0[0]),.doutb(w_n583_0[1]),.din(n583));
	jspl jspl_w_n584_0(.douta(w_n584_0[0]),.doutb(w_n584_0[1]),.din(n584));
	jspl jspl_w_n589_0(.douta(w_n589_0[0]),.doutb(w_n589_0[1]),.din(n589));
	jspl3 jspl3_w_n590_0(.douta(w_n590_0[0]),.doutb(w_n590_0[1]),.doutc(w_n590_0[2]),.din(n590));
	jspl3 jspl3_w_n590_1(.douta(w_n590_1[0]),.doutb(w_n590_1[1]),.doutc(w_n590_1[2]),.din(w_n590_0[0]));
	jspl3 jspl3_w_n590_2(.douta(w_n590_2[0]),.doutb(w_n590_2[1]),.doutc(w_n590_2[2]),.din(w_n590_0[1]));
	jspl3 jspl3_w_n590_3(.douta(w_n590_3[0]),.doutb(w_n590_3[1]),.doutc(w_n590_3[2]),.din(w_n590_0[2]));
	jspl3 jspl3_w_n590_4(.douta(w_n590_4[0]),.doutb(w_n590_4[1]),.doutc(w_n590_4[2]),.din(w_n590_1[0]));
	jspl3 jspl3_w_n590_5(.douta(w_n590_5[0]),.doutb(w_n590_5[1]),.doutc(w_n590_5[2]),.din(w_n590_1[1]));
	jspl3 jspl3_w_n590_6(.douta(w_n590_6[0]),.doutb(w_n590_6[1]),.doutc(w_n590_6[2]),.din(w_n590_1[2]));
	jspl3 jspl3_w_n590_7(.douta(w_n590_7[0]),.doutb(w_n590_7[1]),.doutc(w_n590_7[2]),.din(w_n590_2[0]));
	jspl3 jspl3_w_n590_8(.douta(w_n590_8[0]),.doutb(w_n590_8[1]),.doutc(w_n590_8[2]),.din(w_n590_2[1]));
	jspl3 jspl3_w_n590_9(.douta(w_n590_9[0]),.doutb(w_n590_9[1]),.doutc(w_n590_9[2]),.din(w_n590_2[2]));
	jspl3 jspl3_w_n590_10(.douta(w_n590_10[0]),.doutb(w_n590_10[1]),.doutc(w_n590_10[2]),.din(w_n590_3[0]));
	jspl3 jspl3_w_n590_11(.douta(w_n590_11[0]),.doutb(w_n590_11[1]),.doutc(w_n590_11[2]),.din(w_n590_3[1]));
	jspl3 jspl3_w_n590_12(.douta(w_n590_12[0]),.doutb(w_n590_12[1]),.doutc(w_n590_12[2]),.din(w_n590_3[2]));
	jspl3 jspl3_w_n590_13(.douta(w_n590_13[0]),.doutb(w_n590_13[1]),.doutc(w_n590_13[2]),.din(w_n590_4[0]));
	jspl3 jspl3_w_n590_14(.douta(w_n590_14[0]),.doutb(w_n590_14[1]),.doutc(w_n590_14[2]),.din(w_n590_4[1]));
	jspl3 jspl3_w_n590_15(.douta(w_n590_15[0]),.doutb(w_n590_15[1]),.doutc(w_n590_15[2]),.din(w_n590_4[2]));
	jspl3 jspl3_w_n590_16(.douta(w_n590_16[0]),.doutb(w_n590_16[1]),.doutc(w_n590_16[2]),.din(w_n590_5[0]));
	jspl3 jspl3_w_n590_17(.douta(w_n590_17[0]),.doutb(w_n590_17[1]),.doutc(w_n590_17[2]),.din(w_n590_5[1]));
	jspl3 jspl3_w_n590_18(.douta(w_n590_18[0]),.doutb(w_n590_18[1]),.doutc(w_n590_18[2]),.din(w_n590_5[2]));
	jspl3 jspl3_w_n590_19(.douta(w_n590_19[0]),.doutb(w_n590_19[1]),.doutc(w_n590_19[2]),.din(w_n590_6[0]));
	jspl3 jspl3_w_n590_20(.douta(w_n590_20[0]),.doutb(w_n590_20[1]),.doutc(w_n590_20[2]),.din(w_n590_6[1]));
	jspl3 jspl3_w_n590_21(.douta(w_n590_21[0]),.doutb(w_n590_21[1]),.doutc(w_n590_21[2]),.din(w_n590_6[2]));
	jspl3 jspl3_w_n590_22(.douta(w_n590_22[0]),.doutb(w_n590_22[1]),.doutc(w_n590_22[2]),.din(w_n590_7[0]));
	jspl3 jspl3_w_n590_23(.douta(w_n590_23[0]),.doutb(w_n590_23[1]),.doutc(w_n590_23[2]),.din(w_n590_7[1]));
	jspl3 jspl3_w_n590_24(.douta(w_n590_24[0]),.doutb(w_n590_24[1]),.doutc(w_n590_24[2]),.din(w_n590_7[2]));
	jspl3 jspl3_w_n590_25(.douta(w_n590_25[0]),.doutb(w_n590_25[1]),.doutc(w_n590_25[2]),.din(w_n590_8[0]));
	jspl3 jspl3_w_n590_26(.douta(w_n590_26[0]),.doutb(w_n590_26[1]),.doutc(w_n590_26[2]),.din(w_n590_8[1]));
	jspl3 jspl3_w_n590_27(.douta(w_n590_27[0]),.doutb(w_n590_27[1]),.doutc(w_n590_27[2]),.din(w_n590_8[2]));
	jspl3 jspl3_w_n590_28(.douta(w_n590_28[0]),.doutb(w_n590_28[1]),.doutc(w_n590_28[2]),.din(w_n590_9[0]));
	jspl3 jspl3_w_n590_29(.douta(w_n590_29[0]),.doutb(w_n590_29[1]),.doutc(w_n590_29[2]),.din(w_n590_9[1]));
	jspl3 jspl3_w_n590_30(.douta(w_n590_30[0]),.doutb(w_n590_30[1]),.doutc(w_n590_30[2]),.din(w_n590_9[2]));
	jspl3 jspl3_w_n590_31(.douta(w_n590_31[0]),.doutb(w_n590_31[1]),.doutc(w_n590_31[2]),.din(w_n590_10[0]));
	jspl3 jspl3_w_n590_32(.douta(w_n590_32[0]),.doutb(w_n590_32[1]),.doutc(w_n590_32[2]),.din(w_n590_10[1]));
	jspl3 jspl3_w_n590_33(.douta(w_n590_33[0]),.doutb(w_n590_33[1]),.doutc(w_n590_33[2]),.din(w_n590_10[2]));
	jspl3 jspl3_w_n590_34(.douta(w_n590_34[0]),.doutb(w_n590_34[1]),.doutc(w_n590_34[2]),.din(w_n590_11[0]));
	jspl3 jspl3_w_n590_35(.douta(w_n590_35[0]),.doutb(w_n590_35[1]),.doutc(w_n590_35[2]),.din(w_n590_11[1]));
	jspl3 jspl3_w_n595_0(.douta(w_n595_0[0]),.doutb(w_n595_0[1]),.doutc(w_n595_0[2]),.din(n595));
	jspl3 jspl3_w_n595_1(.douta(w_n595_1[0]),.doutb(w_n595_1[1]),.doutc(w_n595_1[2]),.din(w_n595_0[0]));
	jspl3 jspl3_w_n595_2(.douta(w_n595_2[0]),.doutb(w_n595_2[1]),.doutc(w_n595_2[2]),.din(w_n595_0[1]));
	jspl3 jspl3_w_n595_3(.douta(w_n595_3[0]),.doutb(w_n595_3[1]),.doutc(w_n595_3[2]),.din(w_n595_0[2]));
	jspl3 jspl3_w_n595_4(.douta(w_n595_4[0]),.doutb(w_n595_4[1]),.doutc(w_n595_4[2]),.din(w_n595_1[0]));
	jspl3 jspl3_w_n595_5(.douta(w_n595_5[0]),.doutb(w_n595_5[1]),.doutc(w_n595_5[2]),.din(w_n595_1[1]));
	jspl3 jspl3_w_n595_6(.douta(w_n595_6[0]),.doutb(w_n595_6[1]),.doutc(w_n595_6[2]),.din(w_n595_1[2]));
	jspl3 jspl3_w_n595_7(.douta(w_n595_7[0]),.doutb(w_n595_7[1]),.doutc(w_n595_7[2]),.din(w_n595_2[0]));
	jspl3 jspl3_w_n595_8(.douta(w_n595_8[0]),.doutb(w_n595_8[1]),.doutc(w_n595_8[2]),.din(w_n595_2[1]));
	jspl3 jspl3_w_n595_9(.douta(w_n595_9[0]),.doutb(w_n595_9[1]),.doutc(w_n595_9[2]),.din(w_n595_2[2]));
	jspl3 jspl3_w_n595_10(.douta(w_n595_10[0]),.doutb(w_n595_10[1]),.doutc(w_n595_10[2]),.din(w_n595_3[0]));
	jspl3 jspl3_w_n595_11(.douta(w_n595_11[0]),.doutb(w_n595_11[1]),.doutc(w_n595_11[2]),.din(w_n595_3[1]));
	jspl3 jspl3_w_n595_12(.douta(w_n595_12[0]),.doutb(w_n595_12[1]),.doutc(w_n595_12[2]),.din(w_n595_3[2]));
	jspl3 jspl3_w_n595_13(.douta(w_n595_13[0]),.doutb(w_n595_13[1]),.doutc(w_n595_13[2]),.din(w_n595_4[0]));
	jspl3 jspl3_w_n595_14(.douta(w_n595_14[0]),.doutb(w_n595_14[1]),.doutc(w_n595_14[2]),.din(w_n595_4[1]));
	jspl3 jspl3_w_n595_15(.douta(w_n595_15[0]),.doutb(w_n595_15[1]),.doutc(w_n595_15[2]),.din(w_n595_4[2]));
	jspl3 jspl3_w_n595_16(.douta(w_n595_16[0]),.doutb(w_n595_16[1]),.doutc(w_n595_16[2]),.din(w_n595_5[0]));
	jspl3 jspl3_w_n595_17(.douta(w_n595_17[0]),.doutb(w_n595_17[1]),.doutc(w_n595_17[2]),.din(w_n595_5[1]));
	jspl3 jspl3_w_n595_18(.douta(w_n595_18[0]),.doutb(w_n595_18[1]),.doutc(w_n595_18[2]),.din(w_n595_5[2]));
	jspl3 jspl3_w_n595_19(.douta(w_n595_19[0]),.doutb(w_n595_19[1]),.doutc(w_n595_19[2]),.din(w_n595_6[0]));
	jspl3 jspl3_w_n595_20(.douta(w_n595_20[0]),.doutb(w_n595_20[1]),.doutc(w_n595_20[2]),.din(w_n595_6[1]));
	jspl3 jspl3_w_n595_21(.douta(w_n595_21[0]),.doutb(w_n595_21[1]),.doutc(w_n595_21[2]),.din(w_n595_6[2]));
	jspl3 jspl3_w_n595_22(.douta(w_n595_22[0]),.doutb(w_n595_22[1]),.doutc(w_n595_22[2]),.din(w_n595_7[0]));
	jspl3 jspl3_w_n595_23(.douta(w_n595_23[0]),.doutb(w_n595_23[1]),.doutc(w_n595_23[2]),.din(w_n595_7[1]));
	jspl3 jspl3_w_n595_24(.douta(w_n595_24[0]),.doutb(w_n595_24[1]),.doutc(w_n595_24[2]),.din(w_n595_7[2]));
	jspl3 jspl3_w_n595_25(.douta(w_n595_25[0]),.doutb(w_n595_25[1]),.doutc(w_n595_25[2]),.din(w_n595_8[0]));
	jspl3 jspl3_w_n595_26(.douta(w_n595_26[0]),.doutb(w_n595_26[1]),.doutc(w_n595_26[2]),.din(w_n595_8[1]));
	jspl3 jspl3_w_n595_27(.douta(w_n595_27[0]),.doutb(w_n595_27[1]),.doutc(w_n595_27[2]),.din(w_n595_8[2]));
	jspl3 jspl3_w_n595_28(.douta(w_n595_28[0]),.doutb(w_n595_28[1]),.doutc(w_n595_28[2]),.din(w_n595_9[0]));
	jspl3 jspl3_w_n595_29(.douta(w_n595_29[0]),.doutb(w_n595_29[1]),.doutc(w_n595_29[2]),.din(w_n595_9[1]));
	jspl3 jspl3_w_n595_30(.douta(w_n595_30[0]),.doutb(w_n595_30[1]),.doutc(w_n595_30[2]),.din(w_n595_9[2]));
	jspl3 jspl3_w_n595_31(.douta(w_n595_31[0]),.doutb(w_n595_31[1]),.doutc(w_n595_31[2]),.din(w_n595_10[0]));
	jspl3 jspl3_w_n595_32(.douta(w_n595_32[0]),.doutb(w_n595_32[1]),.doutc(w_n595_32[2]),.din(w_n595_10[1]));
	jspl3 jspl3_w_n595_33(.douta(w_n595_33[0]),.doutb(w_n595_33[1]),.doutc(w_n595_33[2]),.din(w_n595_10[2]));
	jspl3 jspl3_w_n595_34(.douta(w_n595_34[0]),.doutb(w_n595_34[1]),.doutc(w_n595_34[2]),.din(w_n595_11[0]));
	jspl3 jspl3_w_n595_35(.douta(w_n595_35[0]),.doutb(w_n595_35[1]),.doutc(w_n595_35[2]),.din(w_n595_11[1]));
	jspl3 jspl3_w_n595_36(.douta(w_n595_36[0]),.doutb(w_n595_36[1]),.doutc(w_n595_36[2]),.din(w_n595_11[2]));
	jspl3 jspl3_w_n595_37(.douta(w_n595_37[0]),.doutb(w_n595_37[1]),.doutc(w_n595_37[2]),.din(w_n595_12[0]));
	jspl3 jspl3_w_n595_38(.douta(w_n595_38[0]),.doutb(w_n595_38[1]),.doutc(w_n595_38[2]),.din(w_n595_12[1]));
	jspl3 jspl3_w_n598_0(.douta(w_n598_0[0]),.doutb(w_n598_0[1]),.doutc(w_n598_0[2]),.din(n598));
	jspl jspl_w_n598_1(.douta(w_n598_1[0]),.doutb(w_n598_1[1]),.din(w_n598_0[0]));
	jspl3 jspl3_w_n599_0(.douta(w_n599_0[0]),.doutb(w_n599_0[1]),.doutc(w_n599_0[2]),.din(n599));
	jspl3 jspl3_w_n603_0(.douta(w_n603_0[0]),.doutb(w_n603_0[1]),.doutc(w_n603_0[2]),.din(n603));
	jspl jspl_w_n604_0(.douta(w_n604_0[0]),.doutb(w_n604_0[1]),.din(n604));
	jspl jspl_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.din(n605));
	jspl jspl_w_n606_0(.douta(w_n606_0[0]),.doutb(w_n606_0[1]),.din(n606));
	jspl jspl_w_n608_0(.douta(w_n608_0[0]),.doutb(w_n608_0[1]),.din(n608));
	jspl jspl_w_n610_0(.douta(w_n610_0[0]),.doutb(w_n610_0[1]),.din(n610));
	jspl jspl_w_n612_0(.douta(w_n612_0[0]),.doutb(w_n612_0[1]),.din(n612));
	jspl jspl_w_n615_0(.douta(w_n615_0[0]),.doutb(w_n615_0[1]),.din(n615));
	jspl jspl_w_n620_0(.douta(w_n620_0[0]),.doutb(w_n620_0[1]),.din(n620));
	jspl3 jspl3_w_n622_0(.douta(w_n622_0[0]),.doutb(w_n622_0[1]),.doutc(w_n622_0[2]),.din(n622));
	jspl jspl_w_n623_0(.douta(w_n623_0[0]),.doutb(w_n623_0[1]),.din(n623));
	jspl jspl_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.din(n627));
	jspl jspl_w_n628_0(.douta(w_n628_0[0]),.doutb(w_n628_0[1]),.din(n628));
	jspl jspl_w_n630_0(.douta(w_n630_0[0]),.doutb(w_n630_0[1]),.din(n630));
	jspl jspl_w_n634_0(.douta(w_n634_0[0]),.doutb(w_n634_0[1]),.din(n634));
	jspl jspl_w_n636_0(.douta(w_n636_0[0]),.doutb(w_n636_0[1]),.din(n636));
	jspl jspl_w_n637_0(.douta(w_n637_0[0]),.doutb(w_n637_0[1]),.din(n637));
	jspl3 jspl3_w_n638_0(.douta(w_n638_0[0]),.doutb(w_n638_0[1]),.doutc(w_n638_0[2]),.din(n638));
	jspl jspl_w_n639_0(.douta(w_n639_0[0]),.doutb(w_n639_0[1]),.din(n639));
	jspl jspl_w_n643_0(.douta(w_n643_0[0]),.doutb(w_n643_0[1]),.din(n643));
	jspl jspl_w_n645_0(.douta(w_n645_0[0]),.doutb(w_n645_0[1]),.din(n645));
	jspl jspl_w_n647_0(.douta(w_n647_0[0]),.doutb(w_n647_0[1]),.din(n647));
	jspl jspl_w_n649_0(.douta(w_n649_0[0]),.doutb(w_n649_0[1]),.din(n649));
	jspl jspl_w_n651_0(.douta(w_n651_0[0]),.doutb(w_n651_0[1]),.din(n651));
	jspl jspl_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.din(n657));
	jspl3 jspl3_w_n659_0(.douta(w_n659_0[0]),.doutb(w_n659_0[1]),.doutc(w_n659_0[2]),.din(n659));
	jspl jspl_w_n665_0(.douta(w_n665_0[0]),.doutb(w_n665_0[1]),.din(n665));
	jspl3 jspl3_w_n668_0(.douta(w_n668_0[0]),.doutb(w_n668_0[1]),.doutc(w_n668_0[2]),.din(n668));
	jspl3 jspl3_w_n672_0(.douta(w_n672_0[0]),.doutb(w_n672_0[1]),.doutc(w_n672_0[2]),.din(n672));
	jspl jspl_w_n673_0(.douta(w_n673_0[0]),.doutb(w_n673_0[1]),.din(n673));
	jspl jspl_w_n678_0(.douta(w_n678_0[0]),.doutb(w_n678_0[1]),.din(n678));
	jspl3 jspl3_w_n679_0(.douta(w_n679_0[0]),.doutb(w_n679_0[1]),.doutc(w_n679_0[2]),.din(n679));
	jspl jspl_w_n684_0(.douta(w_n684_0[0]),.doutb(w_n684_0[1]),.din(n684));
	jspl3 jspl3_w_n690_0(.douta(w_n690_0[0]),.doutb(w_n690_0[1]),.doutc(w_n690_0[2]),.din(n690));
	jspl jspl_w_n690_1(.douta(w_n690_1[0]),.doutb(w_n690_1[1]),.din(w_n690_0[0]));
	jspl jspl_w_n691_0(.douta(w_n691_0[0]),.doutb(w_n691_0[1]),.din(n691));
	jspl3 jspl3_w_n694_0(.douta(w_n694_0[0]),.doutb(w_n694_0[1]),.doutc(w_n694_0[2]),.din(n694));
	jspl jspl_w_n695_0(.douta(w_n695_0[0]),.doutb(w_n695_0[1]),.din(n695));
	jspl jspl_w_n696_0(.douta(w_n696_0[0]),.doutb(w_n696_0[1]),.din(n696));
	jspl jspl_w_n697_0(.douta(w_n697_0[0]),.doutb(w_n697_0[1]),.din(n697));
	jspl jspl_w_n699_0(.douta(w_n699_0[0]),.doutb(w_n699_0[1]),.din(n699));
	jspl jspl_w_n701_0(.douta(w_n701_0[0]),.doutb(w_n701_0[1]),.din(n701));
	jspl jspl_w_n703_0(.douta(w_n703_0[0]),.doutb(w_n703_0[1]),.din(n703));
	jspl jspl_w_n712_0(.douta(w_n712_0[0]),.doutb(w_n712_0[1]),.din(n712));
	jspl3 jspl3_w_n714_0(.douta(w_n714_0[0]),.doutb(w_n714_0[1]),.doutc(w_n714_0[2]),.din(n714));
	jspl jspl_w_n715_0(.douta(w_n715_0[0]),.doutb(w_n715_0[1]),.din(n715));
	jspl jspl_w_n719_0(.douta(w_n719_0[0]),.doutb(w_n719_0[1]),.din(n719));
	jspl jspl_w_n721_0(.douta(w_n721_0[0]),.doutb(w_n721_0[1]),.din(n721));
	jspl jspl_w_n723_0(.douta(w_n723_0[0]),.doutb(w_n723_0[1]),.din(n723));
	jspl jspl_w_n728_0(.douta(w_n728_0[0]),.doutb(w_n728_0[1]),.din(n728));
	jspl jspl_w_n730_0(.douta(w_n730_0[0]),.doutb(w_n730_0[1]),.din(n730));
	jspl jspl_w_n731_0(.douta(w_n731_0[0]),.doutb(w_n731_0[1]),.din(n731));
	jspl3 jspl3_w_n732_0(.douta(w_n732_0[0]),.doutb(w_n732_0[1]),.doutc(w_n732_0[2]),.din(n732));
	jspl jspl_w_n733_0(.douta(w_n733_0[0]),.doutb(w_n733_0[1]),.din(n733));
	jspl jspl_w_n738_0(.douta(w_n738_0[0]),.doutb(w_n738_0[1]),.din(n738));
	jspl jspl_w_n739_0(.douta(w_n739_0[0]),.doutb(w_n739_0[1]),.din(n739));
	jspl jspl_w_n741_0(.douta(w_n741_0[0]),.doutb(w_n741_0[1]),.din(n741));
	jspl jspl_w_n743_0(.douta(w_n743_0[0]),.doutb(w_n743_0[1]),.din(n743));
	jspl jspl_w_n746_0(.douta(w_n746_0[0]),.doutb(w_n746_0[1]),.din(n746));
	jspl jspl_w_n752_0(.douta(w_n752_0[0]),.doutb(w_n752_0[1]),.din(n752));
	jspl3 jspl3_w_n754_0(.douta(w_n754_0[0]),.doutb(w_n754_0[1]),.doutc(w_n754_0[2]),.din(n754));
	jspl jspl_w_n755_0(.douta(w_n755_0[0]),.doutb(w_n755_0[1]),.din(n755));
	jspl jspl_w_n759_0(.douta(w_n759_0[0]),.doutb(w_n759_0[1]),.din(n759));
	jspl jspl_w_n760_0(.douta(w_n760_0[0]),.doutb(w_n760_0[1]),.din(n760));
	jspl jspl_w_n762_0(.douta(w_n762_0[0]),.doutb(w_n762_0[1]),.din(n762));
	jspl jspl_w_n767_0(.douta(w_n767_0[0]),.doutb(w_n767_0[1]),.din(n767));
	jspl jspl_w_n769_0(.douta(w_n769_0[0]),.doutb(w_n769_0[1]),.din(n769));
	jspl jspl_w_n770_0(.douta(w_n770_0[0]),.doutb(w_n770_0[1]),.din(n770));
	jspl3 jspl3_w_n771_0(.douta(w_n771_0[0]),.doutb(w_n771_0[1]),.doutc(w_n771_0[2]),.din(n771));
	jspl3 jspl3_w_n771_1(.douta(w_n771_1[0]),.doutb(w_n771_1[1]),.doutc(w_n771_1[2]),.din(w_n771_0[0]));
	jspl3 jspl3_w_n774_0(.douta(w_n774_0[0]),.doutb(w_n774_0[1]),.doutc(w_n774_0[2]),.din(n774));
	jspl jspl_w_n774_1(.douta(w_n774_1[0]),.doutb(w_n774_1[1]),.din(w_n774_0[0]));
	jspl3 jspl3_w_n776_0(.douta(w_n776_0[0]),.doutb(w_n776_0[1]),.doutc(w_n776_0[2]),.din(n776));
	jspl jspl_w_n777_0(.douta(w_n777_0[0]),.doutb(w_n777_0[1]),.din(n777));
	jspl jspl_w_n778_0(.douta(w_n778_0[0]),.doutb(w_n778_0[1]),.din(n778));
	jspl jspl_w_n784_0(.douta(w_n784_0[0]),.doutb(w_n784_0[1]),.din(n784));
	jspl jspl_w_n785_0(.douta(w_n785_0[0]),.doutb(w_n785_0[1]),.din(n785));
	jspl jspl_w_n790_0(.douta(w_n790_0[0]),.doutb(w_n790_0[1]),.din(n790));
	jspl3 jspl3_w_n791_0(.douta(w_n791_0[0]),.doutb(w_n791_0[1]),.doutc(w_n791_0[2]),.din(n791));
	jspl3 jspl3_w_n791_1(.douta(w_n791_1[0]),.doutb(w_n791_1[1]),.doutc(w_n791_1[2]),.din(w_n791_0[0]));
	jspl3 jspl3_w_n791_2(.douta(w_n791_2[0]),.doutb(w_n791_2[1]),.doutc(w_n791_2[2]),.din(w_n791_0[1]));
	jspl3 jspl3_w_n791_3(.douta(w_n791_3[0]),.doutb(w_n791_3[1]),.doutc(w_n791_3[2]),.din(w_n791_0[2]));
	jspl3 jspl3_w_n791_4(.douta(w_n791_4[0]),.doutb(w_n791_4[1]),.doutc(w_n791_4[2]),.din(w_n791_1[0]));
	jspl3 jspl3_w_n791_5(.douta(w_n791_5[0]),.doutb(w_n791_5[1]),.doutc(w_n791_5[2]),.din(w_n791_1[1]));
	jspl3 jspl3_w_n791_6(.douta(w_n791_6[0]),.doutb(w_n791_6[1]),.doutc(w_n791_6[2]),.din(w_n791_1[2]));
	jspl3 jspl3_w_n791_7(.douta(w_n791_7[0]),.doutb(w_n791_7[1]),.doutc(w_n791_7[2]),.din(w_n791_2[0]));
	jspl3 jspl3_w_n791_8(.douta(w_n791_8[0]),.doutb(w_n791_8[1]),.doutc(w_n791_8[2]),.din(w_n791_2[1]));
	jspl3 jspl3_w_n791_9(.douta(w_n791_9[0]),.doutb(w_n791_9[1]),.doutc(w_n791_9[2]),.din(w_n791_2[2]));
	jspl3 jspl3_w_n791_10(.douta(w_n791_10[0]),.doutb(w_n791_10[1]),.doutc(w_n791_10[2]),.din(w_n791_3[0]));
	jspl3 jspl3_w_n791_11(.douta(w_n791_11[0]),.doutb(w_n791_11[1]),.doutc(w_n791_11[2]),.din(w_n791_3[1]));
	jspl3 jspl3_w_n791_12(.douta(w_n791_12[0]),.doutb(w_n791_12[1]),.doutc(w_n791_12[2]),.din(w_n791_3[2]));
	jspl3 jspl3_w_n791_13(.douta(w_n791_13[0]),.doutb(w_n791_13[1]),.doutc(w_n791_13[2]),.din(w_n791_4[0]));
	jspl3 jspl3_w_n791_14(.douta(w_n791_14[0]),.doutb(w_n791_14[1]),.doutc(w_n791_14[2]),.din(w_n791_4[1]));
	jspl3 jspl3_w_n791_15(.douta(w_n791_15[0]),.doutb(w_n791_15[1]),.doutc(w_n791_15[2]),.din(w_n791_4[2]));
	jspl3 jspl3_w_n791_16(.douta(w_n791_16[0]),.doutb(w_n791_16[1]),.doutc(w_n791_16[2]),.din(w_n791_5[0]));
	jspl3 jspl3_w_n791_17(.douta(w_n791_17[0]),.doutb(w_n791_17[1]),.doutc(w_n791_17[2]),.din(w_n791_5[1]));
	jspl3 jspl3_w_n791_18(.douta(w_n791_18[0]),.doutb(w_n791_18[1]),.doutc(w_n791_18[2]),.din(w_n791_5[2]));
	jspl3 jspl3_w_n791_19(.douta(w_n791_19[0]),.doutb(w_n791_19[1]),.doutc(w_n791_19[2]),.din(w_n791_6[0]));
	jspl3 jspl3_w_n791_20(.douta(w_n791_20[0]),.doutb(w_n791_20[1]),.doutc(w_n791_20[2]),.din(w_n791_6[1]));
	jspl3 jspl3_w_n791_21(.douta(w_n791_21[0]),.doutb(w_n791_21[1]),.doutc(w_n791_21[2]),.din(w_n791_6[2]));
	jspl3 jspl3_w_n791_22(.douta(w_n791_22[0]),.doutb(w_n791_22[1]),.doutc(w_n791_22[2]),.din(w_n791_7[0]));
	jspl3 jspl3_w_n791_23(.douta(w_n791_23[0]),.doutb(w_n791_23[1]),.doutc(w_n791_23[2]),.din(w_n791_7[1]));
	jspl3 jspl3_w_n791_24(.douta(w_n791_24[0]),.doutb(w_n791_24[1]),.doutc(w_n791_24[2]),.din(w_n791_7[2]));
	jspl3 jspl3_w_n791_25(.douta(w_n791_25[0]),.doutb(w_n791_25[1]),.doutc(w_n791_25[2]),.din(w_n791_8[0]));
	jspl3 jspl3_w_n791_26(.douta(w_n791_26[0]),.doutb(w_n791_26[1]),.doutc(w_n791_26[2]),.din(w_n791_8[1]));
	jspl3 jspl3_w_n791_27(.douta(w_n791_27[0]),.doutb(w_n791_27[1]),.doutc(w_n791_27[2]),.din(w_n791_8[2]));
	jspl3 jspl3_w_n791_28(.douta(w_n791_28[0]),.doutb(w_n791_28[1]),.doutc(w_n791_28[2]),.din(w_n791_9[0]));
	jspl3 jspl3_w_n791_29(.douta(w_n791_29[0]),.doutb(w_n791_29[1]),.doutc(w_n791_29[2]),.din(w_n791_9[1]));
	jspl3 jspl3_w_n791_30(.douta(w_n791_30[0]),.doutb(w_n791_30[1]),.doutc(w_n791_30[2]),.din(w_n791_9[2]));
	jspl3 jspl3_w_n791_31(.douta(w_n791_31[0]),.doutb(w_n791_31[1]),.doutc(w_n791_31[2]),.din(w_n791_10[0]));
	jspl3 jspl3_w_n791_32(.douta(w_n791_32[0]),.doutb(w_n791_32[1]),.doutc(w_n791_32[2]),.din(w_n791_10[1]));
	jspl3 jspl3_w_n791_33(.douta(w_n791_33[0]),.doutb(w_n791_33[1]),.doutc(w_n791_33[2]),.din(w_n791_10[2]));
	jspl jspl_w_n791_34(.douta(w_n791_34[0]),.doutb(w_n791_34[1]),.din(w_n791_11[0]));
	jspl3 jspl3_w_n796_0(.douta(w_n796_0[0]),.doutb(w_n796_0[1]),.doutc(w_n796_0[2]),.din(n796));
	jspl3 jspl3_w_n796_1(.douta(w_n796_1[0]),.doutb(w_n796_1[1]),.doutc(w_n796_1[2]),.din(w_n796_0[0]));
	jspl3 jspl3_w_n796_2(.douta(w_n796_2[0]),.doutb(w_n796_2[1]),.doutc(w_n796_2[2]),.din(w_n796_0[1]));
	jspl3 jspl3_w_n796_3(.douta(w_n796_3[0]),.doutb(w_n796_3[1]),.doutc(w_n796_3[2]),.din(w_n796_0[2]));
	jspl3 jspl3_w_n796_4(.douta(w_n796_4[0]),.doutb(w_n796_4[1]),.doutc(w_n796_4[2]),.din(w_n796_1[0]));
	jspl3 jspl3_w_n796_5(.douta(w_n796_5[0]),.doutb(w_n796_5[1]),.doutc(w_n796_5[2]),.din(w_n796_1[1]));
	jspl3 jspl3_w_n796_6(.douta(w_n796_6[0]),.doutb(w_n796_6[1]),.doutc(w_n796_6[2]),.din(w_n796_1[2]));
	jspl3 jspl3_w_n796_7(.douta(w_n796_7[0]),.doutb(w_n796_7[1]),.doutc(w_n796_7[2]),.din(w_n796_2[0]));
	jspl3 jspl3_w_n796_8(.douta(w_n796_8[0]),.doutb(w_n796_8[1]),.doutc(w_n796_8[2]),.din(w_n796_2[1]));
	jspl3 jspl3_w_n796_9(.douta(w_n796_9[0]),.doutb(w_n796_9[1]),.doutc(w_n796_9[2]),.din(w_n796_2[2]));
	jspl3 jspl3_w_n796_10(.douta(w_n796_10[0]),.doutb(w_n796_10[1]),.doutc(w_n796_10[2]),.din(w_n796_3[0]));
	jspl3 jspl3_w_n796_11(.douta(w_n796_11[0]),.doutb(w_n796_11[1]),.doutc(w_n796_11[2]),.din(w_n796_3[1]));
	jspl3 jspl3_w_n796_12(.douta(w_n796_12[0]),.doutb(w_n796_12[1]),.doutc(w_n796_12[2]),.din(w_n796_3[2]));
	jspl3 jspl3_w_n796_13(.douta(w_n796_13[0]),.doutb(w_n796_13[1]),.doutc(w_n796_13[2]),.din(w_n796_4[0]));
	jspl3 jspl3_w_n796_14(.douta(w_n796_14[0]),.doutb(w_n796_14[1]),.doutc(w_n796_14[2]),.din(w_n796_4[1]));
	jspl3 jspl3_w_n796_15(.douta(w_n796_15[0]),.doutb(w_n796_15[1]),.doutc(w_n796_15[2]),.din(w_n796_4[2]));
	jspl3 jspl3_w_n796_16(.douta(w_n796_16[0]),.doutb(w_n796_16[1]),.doutc(w_n796_16[2]),.din(w_n796_5[0]));
	jspl3 jspl3_w_n796_17(.douta(w_n796_17[0]),.doutb(w_n796_17[1]),.doutc(w_n796_17[2]),.din(w_n796_5[1]));
	jspl3 jspl3_w_n796_18(.douta(w_n796_18[0]),.doutb(w_n796_18[1]),.doutc(w_n796_18[2]),.din(w_n796_5[2]));
	jspl3 jspl3_w_n796_19(.douta(w_n796_19[0]),.doutb(w_n796_19[1]),.doutc(w_n796_19[2]),.din(w_n796_6[0]));
	jspl3 jspl3_w_n796_20(.douta(w_n796_20[0]),.doutb(w_n796_20[1]),.doutc(w_n796_20[2]),.din(w_n796_6[1]));
	jspl3 jspl3_w_n796_21(.douta(w_n796_21[0]),.doutb(w_n796_21[1]),.doutc(w_n796_21[2]),.din(w_n796_6[2]));
	jspl3 jspl3_w_n796_22(.douta(w_n796_22[0]),.doutb(w_n796_22[1]),.doutc(w_n796_22[2]),.din(w_n796_7[0]));
	jspl3 jspl3_w_n796_23(.douta(w_n796_23[0]),.doutb(w_n796_23[1]),.doutc(w_n796_23[2]),.din(w_n796_7[1]));
	jspl3 jspl3_w_n796_24(.douta(w_n796_24[0]),.doutb(w_n796_24[1]),.doutc(w_n796_24[2]),.din(w_n796_7[2]));
	jspl3 jspl3_w_n796_25(.douta(w_n796_25[0]),.doutb(w_n796_25[1]),.doutc(w_n796_25[2]),.din(w_n796_8[0]));
	jspl3 jspl3_w_n796_26(.douta(w_n796_26[0]),.doutb(w_n796_26[1]),.doutc(w_n796_26[2]),.din(w_n796_8[1]));
	jspl3 jspl3_w_n796_27(.douta(w_n796_27[0]),.doutb(w_n796_27[1]),.doutc(w_n796_27[2]),.din(w_n796_8[2]));
	jspl3 jspl3_w_n796_28(.douta(w_n796_28[0]),.doutb(w_n796_28[1]),.doutc(w_n796_28[2]),.din(w_n796_9[0]));
	jspl3 jspl3_w_n796_29(.douta(w_n796_29[0]),.doutb(w_n796_29[1]),.doutc(w_n796_29[2]),.din(w_n796_9[1]));
	jspl3 jspl3_w_n796_30(.douta(w_n796_30[0]),.doutb(w_n796_30[1]),.doutc(w_n796_30[2]),.din(w_n796_9[2]));
	jspl3 jspl3_w_n796_31(.douta(w_n796_31[0]),.doutb(w_n796_31[1]),.doutc(w_n796_31[2]),.din(w_n796_10[0]));
	jspl3 jspl3_w_n796_32(.douta(w_n796_32[0]),.doutb(w_n796_32[1]),.doutc(w_n796_32[2]),.din(w_n796_10[1]));
	jspl3 jspl3_w_n796_33(.douta(w_n796_33[0]),.doutb(w_n796_33[1]),.doutc(w_n796_33[2]),.din(w_n796_10[2]));
	jspl3 jspl3_w_n796_34(.douta(w_n796_34[0]),.doutb(w_n796_34[1]),.doutc(w_n796_34[2]),.din(w_n796_11[0]));
	jspl3 jspl3_w_n796_35(.douta(w_n796_35[0]),.doutb(w_n796_35[1]),.doutc(w_n796_35[2]),.din(w_n796_11[1]));
	jspl3 jspl3_w_n796_36(.douta(w_n796_36[0]),.doutb(w_n796_36[1]),.doutc(w_n796_36[2]),.din(w_n796_11[2]));
	jspl3 jspl3_w_n796_37(.douta(w_n796_37[0]),.doutb(w_n796_37[1]),.doutc(w_n796_37[2]),.din(w_n796_12[0]));
	jspl3 jspl3_w_n799_0(.douta(w_n799_0[0]),.doutb(w_n799_0[1]),.doutc(w_n799_0[2]),.din(n799));
	jspl jspl_w_n799_1(.douta(w_n799_1[0]),.doutb(w_n799_1[1]),.din(w_n799_0[0]));
	jspl3 jspl3_w_n800_0(.douta(w_n800_0[0]),.doutb(w_n800_0[1]),.doutc(w_n800_0[2]),.din(n800));
	jspl3 jspl3_w_n804_0(.douta(w_n804_0[0]),.doutb(w_n804_0[1]),.doutc(w_n804_0[2]),.din(n804));
	jspl jspl_w_n805_0(.douta(w_n805_0[0]),.doutb(w_n805_0[1]),.din(n805));
	jspl jspl_w_n806_0(.douta(w_n806_0[0]),.doutb(w_n806_0[1]),.din(n806));
	jspl jspl_w_n807_0(.douta(w_n807_0[0]),.doutb(w_n807_0[1]),.din(n807));
	jspl jspl_w_n809_0(.douta(w_n809_0[0]),.doutb(w_n809_0[1]),.din(n809));
	jspl jspl_w_n811_0(.douta(w_n811_0[0]),.doutb(w_n811_0[1]),.din(n811));
	jspl jspl_w_n813_0(.douta(w_n813_0[0]),.doutb(w_n813_0[1]),.din(n813));
	jspl jspl_w_n816_0(.douta(w_n816_0[0]),.doutb(w_n816_0[1]),.din(n816));
	jspl jspl_w_n821_0(.douta(w_n821_0[0]),.doutb(w_n821_0[1]),.din(n821));
	jspl3 jspl3_w_n823_0(.douta(w_n823_0[0]),.doutb(w_n823_0[1]),.doutc(w_n823_0[2]),.din(n823));
	jspl jspl_w_n824_0(.douta(w_n824_0[0]),.doutb(w_n824_0[1]),.din(n824));
	jspl jspl_w_n828_0(.douta(w_n828_0[0]),.doutb(w_n828_0[1]),.din(n828));
	jspl jspl_w_n829_0(.douta(w_n829_0[0]),.doutb(w_n829_0[1]),.din(n829));
	jspl jspl_w_n831_0(.douta(w_n831_0[0]),.doutb(w_n831_0[1]),.din(n831));
	jspl jspl_w_n835_0(.douta(w_n835_0[0]),.doutb(w_n835_0[1]),.din(n835));
	jspl jspl_w_n837_0(.douta(w_n837_0[0]),.doutb(w_n837_0[1]),.din(n837));
	jspl jspl_w_n838_0(.douta(w_n838_0[0]),.doutb(w_n838_0[1]),.din(n838));
	jspl3 jspl3_w_n839_0(.douta(w_n839_0[0]),.doutb(w_n839_0[1]),.doutc(w_n839_0[2]),.din(n839));
	jspl jspl_w_n840_0(.douta(w_n840_0[0]),.doutb(w_n840_0[1]),.din(n840));
	jspl jspl_w_n844_0(.douta(w_n844_0[0]),.doutb(w_n844_0[1]),.din(n844));
	jspl jspl_w_n846_0(.douta(w_n846_0[0]),.doutb(w_n846_0[1]),.din(n846));
	jspl jspl_w_n848_0(.douta(w_n848_0[0]),.doutb(w_n848_0[1]),.din(n848));
	jspl jspl_w_n850_0(.douta(w_n850_0[0]),.doutb(w_n850_0[1]),.din(n850));
	jspl jspl_w_n852_0(.douta(w_n852_0[0]),.doutb(w_n852_0[1]),.din(n852));
	jspl jspl_w_n858_0(.douta(w_n858_0[0]),.doutb(w_n858_0[1]),.din(n858));
	jspl3 jspl3_w_n860_0(.douta(w_n860_0[0]),.doutb(w_n860_0[1]),.doutc(w_n860_0[2]),.din(n860));
	jspl jspl_w_n861_0(.douta(w_n861_0[0]),.doutb(w_n861_0[1]),.din(n861));
	jspl jspl_w_n866_0(.douta(w_n866_0[0]),.doutb(w_n866_0[1]),.din(n866));
	jspl jspl_w_n868_0(.douta(w_n868_0[0]),.doutb(w_n868_0[1]),.din(n868));
	jspl jspl_w_n870_0(.douta(w_n870_0[0]),.doutb(w_n870_0[1]),.din(n870));
	jspl jspl_w_n874_0(.douta(w_n874_0[0]),.doutb(w_n874_0[1]),.din(n874));
	jspl jspl_w_n876_0(.douta(w_n876_0[0]),.doutb(w_n876_0[1]),.din(n876));
	jspl jspl_w_n877_0(.douta(w_n877_0[0]),.doutb(w_n877_0[1]),.din(n877));
	jspl3 jspl3_w_n878_0(.douta(w_n878_0[0]),.doutb(w_n878_0[1]),.doutc(w_n878_0[2]),.din(n878));
	jspl jspl_w_n885_0(.douta(w_n885_0[0]),.doutb(w_n885_0[1]),.din(n885));
	jspl3 jspl3_w_n887_0(.douta(w_n887_0[0]),.doutb(w_n887_0[1]),.doutc(w_n887_0[2]),.din(n887));
	jspl jspl_w_n889_0(.douta(w_n889_0[0]),.doutb(w_n889_0[1]),.din(n889));
	jspl3 jspl3_w_n894_0(.douta(w_n894_0[0]),.doutb(w_n894_0[1]),.doutc(w_n894_0[2]),.din(n894));
	jspl jspl_w_n895_0(.douta(w_n895_0[0]),.doutb(w_n895_0[1]),.din(n895));
	jspl jspl_w_n896_0(.douta(w_n896_0[0]),.doutb(w_n896_0[1]),.din(n896));
	jspl jspl_w_n901_0(.douta(w_n901_0[0]),.doutb(w_n901_0[1]),.din(n901));
	jspl3 jspl3_w_n902_0(.douta(w_n902_0[0]),.doutb(w_n902_0[1]),.doutc(w_n902_0[2]),.din(n902));
	jspl jspl_w_n907_0(.douta(w_n907_0[0]),.doutb(w_n907_0[1]),.din(n907));
	jspl3 jspl3_w_n913_0(.douta(w_n913_0[0]),.doutb(w_n913_0[1]),.doutc(w_n913_0[2]),.din(n913));
	jspl jspl_w_n913_1(.douta(w_n913_1[0]),.doutb(w_n913_1[1]),.din(w_n913_0[0]));
	jspl jspl_w_n914_0(.douta(w_n914_0[0]),.doutb(w_n914_0[1]),.din(n914));
	jspl3 jspl3_w_n917_0(.douta(w_n917_0[0]),.doutb(w_n917_0[1]),.doutc(w_n917_0[2]),.din(n917));
	jspl jspl_w_n918_0(.douta(w_n918_0[0]),.doutb(w_n918_0[1]),.din(n918));
	jspl jspl_w_n919_0(.douta(w_n919_0[0]),.doutb(w_n919_0[1]),.din(n919));
	jspl jspl_w_n920_0(.douta(w_n920_0[0]),.doutb(w_n920_0[1]),.din(n920));
	jspl jspl_w_n922_0(.douta(w_n922_0[0]),.doutb(w_n922_0[1]),.din(n922));
	jspl jspl_w_n924_0(.douta(w_n924_0[0]),.doutb(w_n924_0[1]),.din(n924));
	jspl jspl_w_n926_0(.douta(w_n926_0[0]),.doutb(w_n926_0[1]),.din(n926));
	jspl jspl_w_n935_0(.douta(w_n935_0[0]),.doutb(w_n935_0[1]),.din(n935));
	jspl3 jspl3_w_n937_0(.douta(w_n937_0[0]),.doutb(w_n937_0[1]),.doutc(w_n937_0[2]),.din(n937));
	jspl jspl_w_n938_0(.douta(w_n938_0[0]),.doutb(w_n938_0[1]),.din(n938));
	jspl jspl_w_n942_0(.douta(w_n942_0[0]),.doutb(w_n942_0[1]),.din(n942));
	jspl jspl_w_n944_0(.douta(w_n944_0[0]),.doutb(w_n944_0[1]),.din(n944));
	jspl jspl_w_n946_0(.douta(w_n946_0[0]),.doutb(w_n946_0[1]),.din(n946));
	jspl jspl_w_n951_0(.douta(w_n951_0[0]),.doutb(w_n951_0[1]),.din(n951));
	jspl jspl_w_n953_0(.douta(w_n953_0[0]),.doutb(w_n953_0[1]),.din(n953));
	jspl jspl_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.din(n954));
	jspl3 jspl3_w_n955_0(.douta(w_n955_0[0]),.doutb(w_n955_0[1]),.doutc(w_n955_0[2]),.din(n955));
	jspl jspl_w_n956_0(.douta(w_n956_0[0]),.doutb(w_n956_0[1]),.din(n956));
	jspl jspl_w_n961_0(.douta(w_n961_0[0]),.doutb(w_n961_0[1]),.din(n961));
	jspl jspl_w_n962_0(.douta(w_n962_0[0]),.doutb(w_n962_0[1]),.din(n962));
	jspl jspl_w_n964_0(.douta(w_n964_0[0]),.doutb(w_n964_0[1]),.din(n964));
	jspl jspl_w_n966_0(.douta(w_n966_0[0]),.doutb(w_n966_0[1]),.din(n966));
	jspl jspl_w_n969_0(.douta(w_n969_0[0]),.doutb(w_n969_0[1]),.din(n969));
	jspl jspl_w_n975_0(.douta(w_n975_0[0]),.doutb(w_n975_0[1]),.din(n975));
	jspl3 jspl3_w_n977_0(.douta(w_n977_0[0]),.doutb(w_n977_0[1]),.doutc(w_n977_0[2]),.din(n977));
	jspl jspl_w_n978_0(.douta(w_n978_0[0]),.doutb(w_n978_0[1]),.din(n978));
	jspl jspl_w_n982_0(.douta(w_n982_0[0]),.doutb(w_n982_0[1]),.din(n982));
	jspl jspl_w_n983_0(.douta(w_n983_0[0]),.doutb(w_n983_0[1]),.din(n983));
	jspl jspl_w_n985_0(.douta(w_n985_0[0]),.doutb(w_n985_0[1]),.din(n985));
	jspl jspl_w_n990_0(.douta(w_n990_0[0]),.doutb(w_n990_0[1]),.din(n990));
	jspl jspl_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.din(n992));
	jspl jspl_w_n993_0(.douta(w_n993_0[0]),.doutb(w_n993_0[1]),.din(n993));
	jspl3 jspl3_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.doutc(w_n994_0[2]),.din(n994));
	jspl jspl_w_n995_0(.douta(w_n995_0[0]),.doutb(w_n995_0[1]),.din(n995));
	jspl jspl_w_n999_0(.douta(w_n999_0[0]),.doutb(w_n999_0[1]),.din(n999));
	jspl jspl_w_n1000_0(.douta(w_n1000_0[0]),.doutb(w_n1000_0[1]),.din(n1000));
	jspl jspl_w_n1002_0(.douta(w_n1002_0[0]),.doutb(w_n1002_0[1]),.din(n1002));
	jspl jspl_w_n1004_0(.douta(w_n1004_0[0]),.doutb(w_n1004_0[1]),.din(n1004));
	jspl jspl_w_n1007_0(.douta(w_n1007_0[0]),.doutb(w_n1007_0[1]),.din(n1007));
	jspl jspl_w_n1013_0(.douta(w_n1013_0[0]),.doutb(w_n1013_0[1]),.din(n1013));
	jspl3 jspl3_w_n1015_0(.douta(w_n1015_0[0]),.doutb(w_n1015_0[1]),.doutc(w_n1015_0[2]),.din(n1015));
	jspl3 jspl3_w_n1015_1(.douta(w_n1015_1[0]),.doutb(w_n1015_1[1]),.doutc(w_n1015_1[2]),.din(w_n1015_0[0]));
	jspl jspl_w_n1018_0(.douta(w_n1018_0[0]),.doutb(w_n1018_0[1]),.din(n1018));
	jspl3 jspl3_w_n1019_0(.douta(w_n1019_0[0]),.doutb(w_n1019_0[1]),.doutc(w_n1019_0[2]),.din(n1019));
	jspl jspl_w_n1020_0(.douta(w_n1020_0[0]),.doutb(w_n1020_0[1]),.din(n1020));
	jspl jspl_w_n1026_0(.douta(w_n1026_0[0]),.doutb(w_n1026_0[1]),.din(n1026));
	jspl3 jspl3_w_n1027_0(.douta(w_n1027_0[0]),.doutb(w_n1027_0[1]),.doutc(w_n1027_0[2]),.din(n1027));
	jspl jspl_w_n1028_0(.douta(w_n1028_0[0]),.doutb(w_n1028_0[1]),.din(n1028));
	jspl jspl_w_n1033_0(.douta(w_n1033_0[0]),.doutb(w_n1033_0[1]),.din(n1033));
	jspl3 jspl3_w_n1034_0(.douta(w_n1034_0[0]),.doutb(w_n1034_0[1]),.doutc(w_n1034_0[2]),.din(n1034));
	jspl3 jspl3_w_n1034_1(.douta(w_n1034_1[0]),.doutb(w_n1034_1[1]),.doutc(w_n1034_1[2]),.din(w_n1034_0[0]));
	jspl3 jspl3_w_n1034_2(.douta(w_n1034_2[0]),.doutb(w_n1034_2[1]),.doutc(w_n1034_2[2]),.din(w_n1034_0[1]));
	jspl3 jspl3_w_n1034_3(.douta(w_n1034_3[0]),.doutb(w_n1034_3[1]),.doutc(w_n1034_3[2]),.din(w_n1034_0[2]));
	jspl3 jspl3_w_n1034_4(.douta(w_n1034_4[0]),.doutb(w_n1034_4[1]),.doutc(w_n1034_4[2]),.din(w_n1034_1[0]));
	jspl3 jspl3_w_n1034_5(.douta(w_n1034_5[0]),.doutb(w_n1034_5[1]),.doutc(w_n1034_5[2]),.din(w_n1034_1[1]));
	jspl3 jspl3_w_n1034_6(.douta(w_n1034_6[0]),.doutb(w_n1034_6[1]),.doutc(w_n1034_6[2]),.din(w_n1034_1[2]));
	jspl3 jspl3_w_n1034_7(.douta(w_n1034_7[0]),.doutb(w_n1034_7[1]),.doutc(w_n1034_7[2]),.din(w_n1034_2[0]));
	jspl3 jspl3_w_n1034_8(.douta(w_n1034_8[0]),.doutb(w_n1034_8[1]),.doutc(w_n1034_8[2]),.din(w_n1034_2[1]));
	jspl3 jspl3_w_n1034_9(.douta(w_n1034_9[0]),.doutb(w_n1034_9[1]),.doutc(w_n1034_9[2]),.din(w_n1034_2[2]));
	jspl3 jspl3_w_n1034_10(.douta(w_n1034_10[0]),.doutb(w_n1034_10[1]),.doutc(w_n1034_10[2]),.din(w_n1034_3[0]));
	jspl3 jspl3_w_n1034_11(.douta(w_n1034_11[0]),.doutb(w_n1034_11[1]),.doutc(w_n1034_11[2]),.din(w_n1034_3[1]));
	jspl3 jspl3_w_n1034_12(.douta(w_n1034_12[0]),.doutb(w_n1034_12[1]),.doutc(w_n1034_12[2]),.din(w_n1034_3[2]));
	jspl3 jspl3_w_n1034_13(.douta(w_n1034_13[0]),.doutb(w_n1034_13[1]),.doutc(w_n1034_13[2]),.din(w_n1034_4[0]));
	jspl3 jspl3_w_n1034_14(.douta(w_n1034_14[0]),.doutb(w_n1034_14[1]),.doutc(w_n1034_14[2]),.din(w_n1034_4[1]));
	jspl3 jspl3_w_n1034_15(.douta(w_n1034_15[0]),.doutb(w_n1034_15[1]),.doutc(w_n1034_15[2]),.din(w_n1034_4[2]));
	jspl3 jspl3_w_n1034_16(.douta(w_n1034_16[0]),.doutb(w_n1034_16[1]),.doutc(w_n1034_16[2]),.din(w_n1034_5[0]));
	jspl3 jspl3_w_n1034_17(.douta(w_n1034_17[0]),.doutb(w_n1034_17[1]),.doutc(w_n1034_17[2]),.din(w_n1034_5[1]));
	jspl3 jspl3_w_n1034_18(.douta(w_n1034_18[0]),.doutb(w_n1034_18[1]),.doutc(w_n1034_18[2]),.din(w_n1034_5[2]));
	jspl3 jspl3_w_n1034_19(.douta(w_n1034_19[0]),.doutb(w_n1034_19[1]),.doutc(w_n1034_19[2]),.din(w_n1034_6[0]));
	jspl3 jspl3_w_n1034_20(.douta(w_n1034_20[0]),.doutb(w_n1034_20[1]),.doutc(w_n1034_20[2]),.din(w_n1034_6[1]));
	jspl3 jspl3_w_n1034_21(.douta(w_n1034_21[0]),.doutb(w_n1034_21[1]),.doutc(w_n1034_21[2]),.din(w_n1034_6[2]));
	jspl3 jspl3_w_n1034_22(.douta(w_n1034_22[0]),.doutb(w_n1034_22[1]),.doutc(w_n1034_22[2]),.din(w_n1034_7[0]));
	jspl3 jspl3_w_n1034_23(.douta(w_n1034_23[0]),.doutb(w_n1034_23[1]),.doutc(w_n1034_23[2]),.din(w_n1034_7[1]));
	jspl3 jspl3_w_n1034_24(.douta(w_n1034_24[0]),.doutb(w_n1034_24[1]),.doutc(w_n1034_24[2]),.din(w_n1034_7[2]));
	jspl3 jspl3_w_n1034_25(.douta(w_n1034_25[0]),.doutb(w_n1034_25[1]),.doutc(w_n1034_25[2]),.din(w_n1034_8[0]));
	jspl3 jspl3_w_n1034_26(.douta(w_n1034_26[0]),.doutb(w_n1034_26[1]),.doutc(w_n1034_26[2]),.din(w_n1034_8[1]));
	jspl3 jspl3_w_n1034_27(.douta(w_n1034_27[0]),.doutb(w_n1034_27[1]),.doutc(w_n1034_27[2]),.din(w_n1034_8[2]));
	jspl3 jspl3_w_n1034_28(.douta(w_n1034_28[0]),.doutb(w_n1034_28[1]),.doutc(w_n1034_28[2]),.din(w_n1034_9[0]));
	jspl3 jspl3_w_n1034_29(.douta(w_n1034_29[0]),.doutb(w_n1034_29[1]),.doutc(w_n1034_29[2]),.din(w_n1034_9[1]));
	jspl3 jspl3_w_n1034_30(.douta(w_n1034_30[0]),.doutb(w_n1034_30[1]),.doutc(w_n1034_30[2]),.din(w_n1034_9[2]));
	jspl3 jspl3_w_n1034_31(.douta(w_n1034_31[0]),.doutb(w_n1034_31[1]),.doutc(w_n1034_31[2]),.din(w_n1034_10[0]));
	jspl3 jspl3_w_n1034_32(.douta(w_n1034_32[0]),.doutb(w_n1034_32[1]),.doutc(w_n1034_32[2]),.din(w_n1034_10[1]));
	jspl jspl_w_n1034_33(.douta(w_n1034_33[0]),.doutb(w_n1034_33[1]),.din(w_n1034_10[2]));
	jspl3 jspl3_w_n1039_0(.douta(w_n1039_0[0]),.doutb(w_n1039_0[1]),.doutc(w_n1039_0[2]),.din(n1039));
	jspl3 jspl3_w_n1039_1(.douta(w_n1039_1[0]),.doutb(w_n1039_1[1]),.doutc(w_n1039_1[2]),.din(w_n1039_0[0]));
	jspl3 jspl3_w_n1039_2(.douta(w_n1039_2[0]),.doutb(w_n1039_2[1]),.doutc(w_n1039_2[2]),.din(w_n1039_0[1]));
	jspl3 jspl3_w_n1039_3(.douta(w_n1039_3[0]),.doutb(w_n1039_3[1]),.doutc(w_n1039_3[2]),.din(w_n1039_0[2]));
	jspl3 jspl3_w_n1039_4(.douta(w_n1039_4[0]),.doutb(w_n1039_4[1]),.doutc(w_n1039_4[2]),.din(w_n1039_1[0]));
	jspl3 jspl3_w_n1039_5(.douta(w_n1039_5[0]),.doutb(w_n1039_5[1]),.doutc(w_n1039_5[2]),.din(w_n1039_1[1]));
	jspl3 jspl3_w_n1039_6(.douta(w_n1039_6[0]),.doutb(w_n1039_6[1]),.doutc(w_n1039_6[2]),.din(w_n1039_1[2]));
	jspl3 jspl3_w_n1039_7(.douta(w_n1039_7[0]),.doutb(w_n1039_7[1]),.doutc(w_n1039_7[2]),.din(w_n1039_2[0]));
	jspl3 jspl3_w_n1039_8(.douta(w_n1039_8[0]),.doutb(w_n1039_8[1]),.doutc(w_n1039_8[2]),.din(w_n1039_2[1]));
	jspl3 jspl3_w_n1039_9(.douta(w_n1039_9[0]),.doutb(w_n1039_9[1]),.doutc(w_n1039_9[2]),.din(w_n1039_2[2]));
	jspl3 jspl3_w_n1039_10(.douta(w_n1039_10[0]),.doutb(w_n1039_10[1]),.doutc(w_n1039_10[2]),.din(w_n1039_3[0]));
	jspl3 jspl3_w_n1039_11(.douta(w_n1039_11[0]),.doutb(w_n1039_11[1]),.doutc(w_n1039_11[2]),.din(w_n1039_3[1]));
	jspl3 jspl3_w_n1039_12(.douta(w_n1039_12[0]),.doutb(w_n1039_12[1]),.doutc(w_n1039_12[2]),.din(w_n1039_3[2]));
	jspl3 jspl3_w_n1039_13(.douta(w_n1039_13[0]),.doutb(w_n1039_13[1]),.doutc(w_n1039_13[2]),.din(w_n1039_4[0]));
	jspl3 jspl3_w_n1039_14(.douta(w_n1039_14[0]),.doutb(w_n1039_14[1]),.doutc(w_n1039_14[2]),.din(w_n1039_4[1]));
	jspl3 jspl3_w_n1039_15(.douta(w_n1039_15[0]),.doutb(w_n1039_15[1]),.doutc(w_n1039_15[2]),.din(w_n1039_4[2]));
	jspl3 jspl3_w_n1039_16(.douta(w_n1039_16[0]),.doutb(w_n1039_16[1]),.doutc(w_n1039_16[2]),.din(w_n1039_5[0]));
	jspl3 jspl3_w_n1039_17(.douta(w_n1039_17[0]),.doutb(w_n1039_17[1]),.doutc(w_n1039_17[2]),.din(w_n1039_5[1]));
	jspl3 jspl3_w_n1039_18(.douta(w_n1039_18[0]),.doutb(w_n1039_18[1]),.doutc(w_n1039_18[2]),.din(w_n1039_5[2]));
	jspl3 jspl3_w_n1039_19(.douta(w_n1039_19[0]),.doutb(w_n1039_19[1]),.doutc(w_n1039_19[2]),.din(w_n1039_6[0]));
	jspl3 jspl3_w_n1039_20(.douta(w_n1039_20[0]),.doutb(w_n1039_20[1]),.doutc(w_n1039_20[2]),.din(w_n1039_6[1]));
	jspl3 jspl3_w_n1039_21(.douta(w_n1039_21[0]),.doutb(w_n1039_21[1]),.doutc(w_n1039_21[2]),.din(w_n1039_6[2]));
	jspl3 jspl3_w_n1039_22(.douta(w_n1039_22[0]),.doutb(w_n1039_22[1]),.doutc(w_n1039_22[2]),.din(w_n1039_7[0]));
	jspl3 jspl3_w_n1039_23(.douta(w_n1039_23[0]),.doutb(w_n1039_23[1]),.doutc(w_n1039_23[2]),.din(w_n1039_7[1]));
	jspl3 jspl3_w_n1039_24(.douta(w_n1039_24[0]),.doutb(w_n1039_24[1]),.doutc(w_n1039_24[2]),.din(w_n1039_7[2]));
	jspl3 jspl3_w_n1039_25(.douta(w_n1039_25[0]),.doutb(w_n1039_25[1]),.doutc(w_n1039_25[2]),.din(w_n1039_8[0]));
	jspl3 jspl3_w_n1039_26(.douta(w_n1039_26[0]),.doutb(w_n1039_26[1]),.doutc(w_n1039_26[2]),.din(w_n1039_8[1]));
	jspl3 jspl3_w_n1039_27(.douta(w_n1039_27[0]),.doutb(w_n1039_27[1]),.doutc(w_n1039_27[2]),.din(w_n1039_8[2]));
	jspl3 jspl3_w_n1039_28(.douta(w_n1039_28[0]),.doutb(w_n1039_28[1]),.doutc(w_n1039_28[2]),.din(w_n1039_9[0]));
	jspl3 jspl3_w_n1039_29(.douta(w_n1039_29[0]),.doutb(w_n1039_29[1]),.doutc(w_n1039_29[2]),.din(w_n1039_9[1]));
	jspl3 jspl3_w_n1039_30(.douta(w_n1039_30[0]),.doutb(w_n1039_30[1]),.doutc(w_n1039_30[2]),.din(w_n1039_9[2]));
	jspl3 jspl3_w_n1039_31(.douta(w_n1039_31[0]),.doutb(w_n1039_31[1]),.doutc(w_n1039_31[2]),.din(w_n1039_10[0]));
	jspl3 jspl3_w_n1039_32(.douta(w_n1039_32[0]),.doutb(w_n1039_32[1]),.doutc(w_n1039_32[2]),.din(w_n1039_10[1]));
	jspl3 jspl3_w_n1039_33(.douta(w_n1039_33[0]),.doutb(w_n1039_33[1]),.doutc(w_n1039_33[2]),.din(w_n1039_10[2]));
	jspl3 jspl3_w_n1039_34(.douta(w_n1039_34[0]),.doutb(w_n1039_34[1]),.doutc(w_n1039_34[2]),.din(w_n1039_11[0]));
	jspl3 jspl3_w_n1039_35(.douta(w_n1039_35[0]),.doutb(w_n1039_35[1]),.doutc(w_n1039_35[2]),.din(w_n1039_11[1]));
	jspl3 jspl3_w_n1039_36(.douta(w_n1039_36[0]),.doutb(w_n1039_36[1]),.doutc(w_n1039_36[2]),.din(w_n1039_11[2]));
	jspl3 jspl3_w_n1039_37(.douta(w_n1039_37[0]),.doutb(w_n1039_37[1]),.doutc(w_n1039_37[2]),.din(w_n1039_12[0]));
	jspl3 jspl3_w_n1042_0(.douta(w_n1042_0[0]),.doutb(w_n1042_0[1]),.doutc(w_n1042_0[2]),.din(n1042));
	jspl jspl_w_n1042_1(.douta(w_n1042_1[0]),.doutb(w_n1042_1[1]),.din(w_n1042_0[0]));
	jspl3 jspl3_w_n1043_0(.douta(w_n1043_0[0]),.doutb(w_n1043_0[1]),.doutc(w_n1043_0[2]),.din(n1043));
	jspl3 jspl3_w_n1047_0(.douta(w_n1047_0[0]),.doutb(w_n1047_0[1]),.doutc(w_n1047_0[2]),.din(n1047));
	jspl jspl_w_n1048_0(.douta(w_n1048_0[0]),.doutb(w_n1048_0[1]),.din(n1048));
	jspl jspl_w_n1049_0(.douta(w_n1049_0[0]),.doutb(w_n1049_0[1]),.din(n1049));
	jspl jspl_w_n1050_0(.douta(w_n1050_0[0]),.doutb(w_n1050_0[1]),.din(n1050));
	jspl jspl_w_n1052_0(.douta(w_n1052_0[0]),.doutb(w_n1052_0[1]),.din(n1052));
	jspl jspl_w_n1054_0(.douta(w_n1054_0[0]),.doutb(w_n1054_0[1]),.din(n1054));
	jspl jspl_w_n1056_0(.douta(w_n1056_0[0]),.doutb(w_n1056_0[1]),.din(n1056));
	jspl jspl_w_n1059_0(.douta(w_n1059_0[0]),.doutb(w_n1059_0[1]),.din(n1059));
	jspl jspl_w_n1064_0(.douta(w_n1064_0[0]),.doutb(w_n1064_0[1]),.din(n1064));
	jspl3 jspl3_w_n1066_0(.douta(w_n1066_0[0]),.doutb(w_n1066_0[1]),.doutc(w_n1066_0[2]),.din(n1066));
	jspl jspl_w_n1067_0(.douta(w_n1067_0[0]),.doutb(w_n1067_0[1]),.din(n1067));
	jspl jspl_w_n1071_0(.douta(w_n1071_0[0]),.doutb(w_n1071_0[1]),.din(n1071));
	jspl jspl_w_n1072_0(.douta(w_n1072_0[0]),.doutb(w_n1072_0[1]),.din(n1072));
	jspl jspl_w_n1074_0(.douta(w_n1074_0[0]),.doutb(w_n1074_0[1]),.din(n1074));
	jspl jspl_w_n1078_0(.douta(w_n1078_0[0]),.doutb(w_n1078_0[1]),.din(n1078));
	jspl jspl_w_n1080_0(.douta(w_n1080_0[0]),.doutb(w_n1080_0[1]),.din(n1080));
	jspl jspl_w_n1081_0(.douta(w_n1081_0[0]),.doutb(w_n1081_0[1]),.din(n1081));
	jspl3 jspl3_w_n1082_0(.douta(w_n1082_0[0]),.doutb(w_n1082_0[1]),.doutc(w_n1082_0[2]),.din(n1082));
	jspl jspl_w_n1083_0(.douta(w_n1083_0[0]),.doutb(w_n1083_0[1]),.din(n1083));
	jspl jspl_w_n1087_0(.douta(w_n1087_0[0]),.doutb(w_n1087_0[1]),.din(n1087));
	jspl jspl_w_n1089_0(.douta(w_n1089_0[0]),.doutb(w_n1089_0[1]),.din(n1089));
	jspl jspl_w_n1091_0(.douta(w_n1091_0[0]),.doutb(w_n1091_0[1]),.din(n1091));
	jspl jspl_w_n1093_0(.douta(w_n1093_0[0]),.doutb(w_n1093_0[1]),.din(n1093));
	jspl jspl_w_n1095_0(.douta(w_n1095_0[0]),.doutb(w_n1095_0[1]),.din(n1095));
	jspl jspl_w_n1101_0(.douta(w_n1101_0[0]),.doutb(w_n1101_0[1]),.din(n1101));
	jspl3 jspl3_w_n1103_0(.douta(w_n1103_0[0]),.doutb(w_n1103_0[1]),.doutc(w_n1103_0[2]),.din(n1103));
	jspl jspl_w_n1104_0(.douta(w_n1104_0[0]),.doutb(w_n1104_0[1]),.din(n1104));
	jspl jspl_w_n1109_0(.douta(w_n1109_0[0]),.doutb(w_n1109_0[1]),.din(n1109));
	jspl jspl_w_n1111_0(.douta(w_n1111_0[0]),.doutb(w_n1111_0[1]),.din(n1111));
	jspl jspl_w_n1113_0(.douta(w_n1113_0[0]),.doutb(w_n1113_0[1]),.din(n1113));
	jspl jspl_w_n1117_0(.douta(w_n1117_0[0]),.doutb(w_n1117_0[1]),.din(n1117));
	jspl jspl_w_n1119_0(.douta(w_n1119_0[0]),.doutb(w_n1119_0[1]),.din(n1119));
	jspl jspl_w_n1120_0(.douta(w_n1120_0[0]),.doutb(w_n1120_0[1]),.din(n1120));
	jspl3 jspl3_w_n1121_0(.douta(w_n1121_0[0]),.doutb(w_n1121_0[1]),.doutc(w_n1121_0[2]),.din(n1121));
	jspl jspl_w_n1122_0(.douta(w_n1122_0[0]),.doutb(w_n1122_0[1]),.din(n1122));
	jspl jspl_w_n1128_0(.douta(w_n1128_0[0]),.doutb(w_n1128_0[1]),.din(n1128));
	jspl jspl_w_n1129_0(.douta(w_n1129_0[0]),.doutb(w_n1129_0[1]),.din(n1129));
	jspl jspl_w_n1131_0(.douta(w_n1131_0[0]),.doutb(w_n1131_0[1]),.din(n1131));
	jspl jspl_w_n1133_0(.douta(w_n1133_0[0]),.doutb(w_n1133_0[1]),.din(n1133));
	jspl jspl_w_n1135_0(.douta(w_n1135_0[0]),.doutb(w_n1135_0[1]),.din(n1135));
	jspl jspl_w_n1141_0(.douta(w_n1141_0[0]),.doutb(w_n1141_0[1]),.din(n1141));
	jspl3 jspl3_w_n1143_0(.douta(w_n1143_0[0]),.doutb(w_n1143_0[1]),.doutc(w_n1143_0[2]),.din(n1143));
	jspl jspl_w_n1148_0(.douta(w_n1148_0[0]),.doutb(w_n1148_0[1]),.din(n1148));
	jspl3 jspl3_w_n1150_0(.douta(w_n1150_0[0]),.doutb(w_n1150_0[1]),.doutc(w_n1150_0[2]),.din(n1150));
	jspl3 jspl3_w_n1154_0(.douta(w_n1154_0[0]),.doutb(w_n1154_0[1]),.doutc(w_n1154_0[2]),.din(n1154));
	jspl jspl_w_n1155_0(.douta(w_n1155_0[0]),.doutb(w_n1155_0[1]),.din(n1155));
	jspl jspl_w_n1160_0(.douta(w_n1160_0[0]),.doutb(w_n1160_0[1]),.din(n1160));
	jspl3 jspl3_w_n1161_0(.douta(w_n1161_0[0]),.doutb(w_n1161_0[1]),.doutc(w_n1161_0[2]),.din(n1161));
	jspl jspl_w_n1166_0(.douta(w_n1166_0[0]),.doutb(w_n1166_0[1]),.din(n1166));
	jspl3 jspl3_w_n1172_0(.douta(w_n1172_0[0]),.doutb(w_n1172_0[1]),.doutc(w_n1172_0[2]),.din(n1172));
	jspl jspl_w_n1172_1(.douta(w_n1172_1[0]),.doutb(w_n1172_1[1]),.din(w_n1172_0[0]));
	jspl jspl_w_n1173_0(.douta(w_n1173_0[0]),.doutb(w_n1173_0[1]),.din(n1173));
	jspl3 jspl3_w_n1176_0(.douta(w_n1176_0[0]),.doutb(w_n1176_0[1]),.doutc(w_n1176_0[2]),.din(n1176));
	jspl jspl_w_n1177_0(.douta(w_n1177_0[0]),.doutb(w_n1177_0[1]),.din(n1177));
	jspl jspl_w_n1178_0(.douta(w_n1178_0[0]),.doutb(w_n1178_0[1]),.din(n1178));
	jspl jspl_w_n1179_0(.douta(w_n1179_0[0]),.doutb(w_n1179_0[1]),.din(n1179));
	jspl jspl_w_n1181_0(.douta(w_n1181_0[0]),.doutb(w_n1181_0[1]),.din(n1181));
	jspl jspl_w_n1183_0(.douta(w_n1183_0[0]),.doutb(w_n1183_0[1]),.din(n1183));
	jspl jspl_w_n1185_0(.douta(w_n1185_0[0]),.doutb(w_n1185_0[1]),.din(n1185));
	jspl jspl_w_n1194_0(.douta(w_n1194_0[0]),.doutb(w_n1194_0[1]),.din(n1194));
	jspl3 jspl3_w_n1196_0(.douta(w_n1196_0[0]),.doutb(w_n1196_0[1]),.doutc(w_n1196_0[2]),.din(n1196));
	jspl jspl_w_n1197_0(.douta(w_n1197_0[0]),.doutb(w_n1197_0[1]),.din(n1197));
	jspl jspl_w_n1201_0(.douta(w_n1201_0[0]),.doutb(w_n1201_0[1]),.din(n1201));
	jspl jspl_w_n1203_0(.douta(w_n1203_0[0]),.doutb(w_n1203_0[1]),.din(n1203));
	jspl jspl_w_n1205_0(.douta(w_n1205_0[0]),.doutb(w_n1205_0[1]),.din(n1205));
	jspl jspl_w_n1210_0(.douta(w_n1210_0[0]),.doutb(w_n1210_0[1]),.din(n1210));
	jspl jspl_w_n1212_0(.douta(w_n1212_0[0]),.doutb(w_n1212_0[1]),.din(n1212));
	jspl jspl_w_n1213_0(.douta(w_n1213_0[0]),.doutb(w_n1213_0[1]),.din(n1213));
	jspl3 jspl3_w_n1214_0(.douta(w_n1214_0[0]),.doutb(w_n1214_0[1]),.doutc(w_n1214_0[2]),.din(n1214));
	jspl jspl_w_n1215_0(.douta(w_n1215_0[0]),.doutb(w_n1215_0[1]),.din(n1215));
	jspl jspl_w_n1220_0(.douta(w_n1220_0[0]),.doutb(w_n1220_0[1]),.din(n1220));
	jspl jspl_w_n1221_0(.douta(w_n1221_0[0]),.doutb(w_n1221_0[1]),.din(n1221));
	jspl jspl_w_n1223_0(.douta(w_n1223_0[0]),.doutb(w_n1223_0[1]),.din(n1223));
	jspl jspl_w_n1225_0(.douta(w_n1225_0[0]),.doutb(w_n1225_0[1]),.din(n1225));
	jspl jspl_w_n1228_0(.douta(w_n1228_0[0]),.doutb(w_n1228_0[1]),.din(n1228));
	jspl jspl_w_n1234_0(.douta(w_n1234_0[0]),.doutb(w_n1234_0[1]),.din(n1234));
	jspl3 jspl3_w_n1236_0(.douta(w_n1236_0[0]),.doutb(w_n1236_0[1]),.doutc(w_n1236_0[2]),.din(n1236));
	jspl jspl_w_n1237_0(.douta(w_n1237_0[0]),.doutb(w_n1237_0[1]),.din(n1237));
	jspl jspl_w_n1241_0(.douta(w_n1241_0[0]),.doutb(w_n1241_0[1]),.din(n1241));
	jspl jspl_w_n1242_0(.douta(w_n1242_0[0]),.doutb(w_n1242_0[1]),.din(n1242));
	jspl jspl_w_n1244_0(.douta(w_n1244_0[0]),.doutb(w_n1244_0[1]),.din(n1244));
	jspl jspl_w_n1249_0(.douta(w_n1249_0[0]),.doutb(w_n1249_0[1]),.din(n1249));
	jspl jspl_w_n1251_0(.douta(w_n1251_0[0]),.doutb(w_n1251_0[1]),.din(n1251));
	jspl jspl_w_n1252_0(.douta(w_n1252_0[0]),.doutb(w_n1252_0[1]),.din(n1252));
	jspl3 jspl3_w_n1253_0(.douta(w_n1253_0[0]),.doutb(w_n1253_0[1]),.doutc(w_n1253_0[2]),.din(n1253));
	jspl jspl_w_n1254_0(.douta(w_n1254_0[0]),.doutb(w_n1254_0[1]),.din(n1254));
	jspl jspl_w_n1258_0(.douta(w_n1258_0[0]),.doutb(w_n1258_0[1]),.din(n1258));
	jspl jspl_w_n1259_0(.douta(w_n1259_0[0]),.doutb(w_n1259_0[1]),.din(n1259));
	jspl jspl_w_n1261_0(.douta(w_n1261_0[0]),.doutb(w_n1261_0[1]),.din(n1261));
	jspl jspl_w_n1263_0(.douta(w_n1263_0[0]),.doutb(w_n1263_0[1]),.din(n1263));
	jspl jspl_w_n1266_0(.douta(w_n1266_0[0]),.doutb(w_n1266_0[1]),.din(n1266));
	jspl jspl_w_n1272_0(.douta(w_n1272_0[0]),.doutb(w_n1272_0[1]),.din(n1272));
	jspl jspl_w_n1274_0(.douta(w_n1274_0[0]),.doutb(w_n1274_0[1]),.din(n1274));
	jspl3 jspl3_w_n1275_0(.douta(w_n1275_0[0]),.doutb(w_n1275_0[1]),.doutc(w_n1275_0[2]),.din(n1275));
	jspl jspl_w_n1279_0(.douta(w_n1279_0[0]),.doutb(w_n1279_0[1]),.din(n1279));
	jspl jspl_w_n1280_0(.douta(w_n1280_0[0]),.doutb(w_n1280_0[1]),.din(n1280));
	jspl3 jspl3_w_n1281_0(.douta(w_n1281_0[0]),.doutb(w_n1281_0[1]),.doutc(w_n1281_0[2]),.din(n1281));
	jspl jspl_w_n1283_0(.douta(w_n1283_0[0]),.doutb(w_n1283_0[1]),.din(n1283));
	jspl jspl_w_n1288_0(.douta(w_n1288_0[0]),.doutb(w_n1288_0[1]),.din(n1288));
	jspl jspl_w_n1290_0(.douta(w_n1290_0[0]),.doutb(w_n1290_0[1]),.din(n1290));
	jspl jspl_w_n1291_0(.douta(w_n1291_0[0]),.doutb(w_n1291_0[1]),.din(n1291));
	jspl3 jspl3_w_n1292_0(.douta(w_n1292_0[0]),.doutb(w_n1292_0[1]),.doutc(w_n1292_0[2]),.din(n1292));
	jspl3 jspl3_w_n1292_1(.douta(w_n1292_1[0]),.doutb(w_n1292_1[1]),.doutc(w_n1292_1[2]),.din(w_n1292_0[0]));
	jspl jspl_w_n1295_0(.douta(w_n1295_0[0]),.doutb(w_n1295_0[1]),.din(n1295));
	jspl3 jspl3_w_n1296_0(.douta(w_n1296_0[0]),.doutb(w_n1296_0[1]),.doutc(w_n1296_0[2]),.din(n1296));
	jspl jspl_w_n1297_0(.douta(w_n1297_0[0]),.doutb(w_n1297_0[1]),.din(n1297));
	jspl jspl_w_n1298_0(.douta(w_n1298_0[0]),.doutb(w_n1298_0[1]),.din(n1298));
	jspl jspl_w_n1304_0(.douta(w_n1304_0[0]),.doutb(w_n1304_0[1]),.din(n1304));
	jspl3 jspl3_w_n1305_0(.douta(w_n1305_0[0]),.doutb(w_n1305_0[1]),.doutc(w_n1305_0[2]),.din(n1305));
	jspl jspl_w_n1306_0(.douta(w_n1306_0[0]),.doutb(w_n1306_0[1]),.din(n1306));
	jspl jspl_w_n1311_0(.douta(w_n1311_0[0]),.doutb(w_n1311_0[1]),.din(n1311));
	jspl3 jspl3_w_n1312_0(.douta(w_n1312_0[0]),.doutb(w_n1312_0[1]),.doutc(w_n1312_0[2]),.din(n1312));
	jspl3 jspl3_w_n1312_1(.douta(w_n1312_1[0]),.doutb(w_n1312_1[1]),.doutc(w_n1312_1[2]),.din(w_n1312_0[0]));
	jspl3 jspl3_w_n1312_2(.douta(w_n1312_2[0]),.doutb(w_n1312_2[1]),.doutc(w_n1312_2[2]),.din(w_n1312_0[1]));
	jspl3 jspl3_w_n1312_3(.douta(w_n1312_3[0]),.doutb(w_n1312_3[1]),.doutc(w_n1312_3[2]),.din(w_n1312_0[2]));
	jspl3 jspl3_w_n1312_4(.douta(w_n1312_4[0]),.doutb(w_n1312_4[1]),.doutc(w_n1312_4[2]),.din(w_n1312_1[0]));
	jspl3 jspl3_w_n1312_5(.douta(w_n1312_5[0]),.doutb(w_n1312_5[1]),.doutc(w_n1312_5[2]),.din(w_n1312_1[1]));
	jspl3 jspl3_w_n1312_6(.douta(w_n1312_6[0]),.doutb(w_n1312_6[1]),.doutc(w_n1312_6[2]),.din(w_n1312_1[2]));
	jspl3 jspl3_w_n1312_7(.douta(w_n1312_7[0]),.doutb(w_n1312_7[1]),.doutc(w_n1312_7[2]),.din(w_n1312_2[0]));
	jspl3 jspl3_w_n1312_8(.douta(w_n1312_8[0]),.doutb(w_n1312_8[1]),.doutc(w_n1312_8[2]),.din(w_n1312_2[1]));
	jspl3 jspl3_w_n1312_9(.douta(w_n1312_9[0]),.doutb(w_n1312_9[1]),.doutc(w_n1312_9[2]),.din(w_n1312_2[2]));
	jspl3 jspl3_w_n1312_10(.douta(w_n1312_10[0]),.doutb(w_n1312_10[1]),.doutc(w_n1312_10[2]),.din(w_n1312_3[0]));
	jspl3 jspl3_w_n1312_11(.douta(w_n1312_11[0]),.doutb(w_n1312_11[1]),.doutc(w_n1312_11[2]),.din(w_n1312_3[1]));
	jspl3 jspl3_w_n1312_12(.douta(w_n1312_12[0]),.doutb(w_n1312_12[1]),.doutc(w_n1312_12[2]),.din(w_n1312_3[2]));
	jspl3 jspl3_w_n1312_13(.douta(w_n1312_13[0]),.doutb(w_n1312_13[1]),.doutc(w_n1312_13[2]),.din(w_n1312_4[0]));
	jspl3 jspl3_w_n1312_14(.douta(w_n1312_14[0]),.doutb(w_n1312_14[1]),.doutc(w_n1312_14[2]),.din(w_n1312_4[1]));
	jspl3 jspl3_w_n1312_15(.douta(w_n1312_15[0]),.doutb(w_n1312_15[1]),.doutc(w_n1312_15[2]),.din(w_n1312_4[2]));
	jspl3 jspl3_w_n1312_16(.douta(w_n1312_16[0]),.doutb(w_n1312_16[1]),.doutc(w_n1312_16[2]),.din(w_n1312_5[0]));
	jspl3 jspl3_w_n1312_17(.douta(w_n1312_17[0]),.doutb(w_n1312_17[1]),.doutc(w_n1312_17[2]),.din(w_n1312_5[1]));
	jspl3 jspl3_w_n1312_18(.douta(w_n1312_18[0]),.doutb(w_n1312_18[1]),.doutc(w_n1312_18[2]),.din(w_n1312_5[2]));
	jspl3 jspl3_w_n1312_19(.douta(w_n1312_19[0]),.doutb(w_n1312_19[1]),.doutc(w_n1312_19[2]),.din(w_n1312_6[0]));
	jspl3 jspl3_w_n1312_20(.douta(w_n1312_20[0]),.doutb(w_n1312_20[1]),.doutc(w_n1312_20[2]),.din(w_n1312_6[1]));
	jspl3 jspl3_w_n1312_21(.douta(w_n1312_21[0]),.doutb(w_n1312_21[1]),.doutc(w_n1312_21[2]),.din(w_n1312_6[2]));
	jspl3 jspl3_w_n1312_22(.douta(w_n1312_22[0]),.doutb(w_n1312_22[1]),.doutc(w_n1312_22[2]),.din(w_n1312_7[0]));
	jspl3 jspl3_w_n1312_23(.douta(w_n1312_23[0]),.doutb(w_n1312_23[1]),.doutc(w_n1312_23[2]),.din(w_n1312_7[1]));
	jspl3 jspl3_w_n1312_24(.douta(w_n1312_24[0]),.doutb(w_n1312_24[1]),.doutc(w_n1312_24[2]),.din(w_n1312_7[2]));
	jspl3 jspl3_w_n1312_25(.douta(w_n1312_25[0]),.doutb(w_n1312_25[1]),.doutc(w_n1312_25[2]),.din(w_n1312_8[0]));
	jspl3 jspl3_w_n1312_26(.douta(w_n1312_26[0]),.doutb(w_n1312_26[1]),.doutc(w_n1312_26[2]),.din(w_n1312_8[1]));
	jspl3 jspl3_w_n1312_27(.douta(w_n1312_27[0]),.doutb(w_n1312_27[1]),.doutc(w_n1312_27[2]),.din(w_n1312_8[2]));
	jspl3 jspl3_w_n1312_28(.douta(w_n1312_28[0]),.doutb(w_n1312_28[1]),.doutc(w_n1312_28[2]),.din(w_n1312_9[0]));
	jspl3 jspl3_w_n1312_29(.douta(w_n1312_29[0]),.doutb(w_n1312_29[1]),.doutc(w_n1312_29[2]),.din(w_n1312_9[1]));
	jspl3 jspl3_w_n1312_30(.douta(w_n1312_30[0]),.doutb(w_n1312_30[1]),.doutc(w_n1312_30[2]),.din(w_n1312_9[2]));
	jspl3 jspl3_w_n1312_31(.douta(w_n1312_31[0]),.doutb(w_n1312_31[1]),.doutc(w_n1312_31[2]),.din(w_n1312_10[0]));
	jspl3 jspl3_w_n1317_0(.douta(w_n1317_0[0]),.doutb(w_n1317_0[1]),.doutc(w_n1317_0[2]),.din(n1317));
	jspl3 jspl3_w_n1317_1(.douta(w_n1317_1[0]),.doutb(w_n1317_1[1]),.doutc(w_n1317_1[2]),.din(w_n1317_0[0]));
	jspl3 jspl3_w_n1317_2(.douta(w_n1317_2[0]),.doutb(w_n1317_2[1]),.doutc(w_n1317_2[2]),.din(w_n1317_0[1]));
	jspl3 jspl3_w_n1317_3(.douta(w_n1317_3[0]),.doutb(w_n1317_3[1]),.doutc(w_n1317_3[2]),.din(w_n1317_0[2]));
	jspl3 jspl3_w_n1317_4(.douta(w_n1317_4[0]),.doutb(w_n1317_4[1]),.doutc(w_n1317_4[2]),.din(w_n1317_1[0]));
	jspl3 jspl3_w_n1317_5(.douta(w_n1317_5[0]),.doutb(w_n1317_5[1]),.doutc(w_n1317_5[2]),.din(w_n1317_1[1]));
	jspl3 jspl3_w_n1317_6(.douta(w_n1317_6[0]),.doutb(w_n1317_6[1]),.doutc(w_n1317_6[2]),.din(w_n1317_1[2]));
	jspl3 jspl3_w_n1317_7(.douta(w_n1317_7[0]),.doutb(w_n1317_7[1]),.doutc(w_n1317_7[2]),.din(w_n1317_2[0]));
	jspl3 jspl3_w_n1317_8(.douta(w_n1317_8[0]),.doutb(w_n1317_8[1]),.doutc(w_n1317_8[2]),.din(w_n1317_2[1]));
	jspl3 jspl3_w_n1317_9(.douta(w_n1317_9[0]),.doutb(w_n1317_9[1]),.doutc(w_n1317_9[2]),.din(w_n1317_2[2]));
	jspl3 jspl3_w_n1317_10(.douta(w_n1317_10[0]),.doutb(w_n1317_10[1]),.doutc(w_n1317_10[2]),.din(w_n1317_3[0]));
	jspl3 jspl3_w_n1317_11(.douta(w_n1317_11[0]),.doutb(w_n1317_11[1]),.doutc(w_n1317_11[2]),.din(w_n1317_3[1]));
	jspl3 jspl3_w_n1317_12(.douta(w_n1317_12[0]),.doutb(w_n1317_12[1]),.doutc(w_n1317_12[2]),.din(w_n1317_3[2]));
	jspl3 jspl3_w_n1317_13(.douta(w_n1317_13[0]),.doutb(w_n1317_13[1]),.doutc(w_n1317_13[2]),.din(w_n1317_4[0]));
	jspl3 jspl3_w_n1317_14(.douta(w_n1317_14[0]),.doutb(w_n1317_14[1]),.doutc(w_n1317_14[2]),.din(w_n1317_4[1]));
	jspl3 jspl3_w_n1317_15(.douta(w_n1317_15[0]),.doutb(w_n1317_15[1]),.doutc(w_n1317_15[2]),.din(w_n1317_4[2]));
	jspl3 jspl3_w_n1317_16(.douta(w_n1317_16[0]),.doutb(w_n1317_16[1]),.doutc(w_n1317_16[2]),.din(w_n1317_5[0]));
	jspl3 jspl3_w_n1317_17(.douta(w_n1317_17[0]),.doutb(w_n1317_17[1]),.doutc(w_n1317_17[2]),.din(w_n1317_5[1]));
	jspl3 jspl3_w_n1317_18(.douta(w_n1317_18[0]),.doutb(w_n1317_18[1]),.doutc(w_n1317_18[2]),.din(w_n1317_5[2]));
	jspl3 jspl3_w_n1317_19(.douta(w_n1317_19[0]),.doutb(w_n1317_19[1]),.doutc(w_n1317_19[2]),.din(w_n1317_6[0]));
	jspl3 jspl3_w_n1317_20(.douta(w_n1317_20[0]),.doutb(w_n1317_20[1]),.doutc(w_n1317_20[2]),.din(w_n1317_6[1]));
	jspl3 jspl3_w_n1317_21(.douta(w_n1317_21[0]),.doutb(w_n1317_21[1]),.doutc(w_n1317_21[2]),.din(w_n1317_6[2]));
	jspl3 jspl3_w_n1317_22(.douta(w_n1317_22[0]),.doutb(w_n1317_22[1]),.doutc(w_n1317_22[2]),.din(w_n1317_7[0]));
	jspl3 jspl3_w_n1317_23(.douta(w_n1317_23[0]),.doutb(w_n1317_23[1]),.doutc(w_n1317_23[2]),.din(w_n1317_7[1]));
	jspl3 jspl3_w_n1317_24(.douta(w_n1317_24[0]),.doutb(w_n1317_24[1]),.doutc(w_n1317_24[2]),.din(w_n1317_7[2]));
	jspl3 jspl3_w_n1317_25(.douta(w_n1317_25[0]),.doutb(w_n1317_25[1]),.doutc(w_n1317_25[2]),.din(w_n1317_8[0]));
	jspl3 jspl3_w_n1317_26(.douta(w_n1317_26[0]),.doutb(w_n1317_26[1]),.doutc(w_n1317_26[2]),.din(w_n1317_8[1]));
	jspl3 jspl3_w_n1317_27(.douta(w_n1317_27[0]),.doutb(w_n1317_27[1]),.doutc(w_n1317_27[2]),.din(w_n1317_8[2]));
	jspl3 jspl3_w_n1317_28(.douta(w_n1317_28[0]),.doutb(w_n1317_28[1]),.doutc(w_n1317_28[2]),.din(w_n1317_9[0]));
	jspl3 jspl3_w_n1317_29(.douta(w_n1317_29[0]),.doutb(w_n1317_29[1]),.doutc(w_n1317_29[2]),.din(w_n1317_9[1]));
	jspl3 jspl3_w_n1317_30(.douta(w_n1317_30[0]),.doutb(w_n1317_30[1]),.doutc(w_n1317_30[2]),.din(w_n1317_9[2]));
	jspl3 jspl3_w_n1317_31(.douta(w_n1317_31[0]),.doutb(w_n1317_31[1]),.doutc(w_n1317_31[2]),.din(w_n1317_10[0]));
	jspl3 jspl3_w_n1317_32(.douta(w_n1317_32[0]),.doutb(w_n1317_32[1]),.doutc(w_n1317_32[2]),.din(w_n1317_10[1]));
	jspl3 jspl3_w_n1317_33(.douta(w_n1317_33[0]),.doutb(w_n1317_33[1]),.doutc(w_n1317_33[2]),.din(w_n1317_10[2]));
	jspl3 jspl3_w_n1317_34(.douta(w_n1317_34[0]),.doutb(w_n1317_34[1]),.doutc(w_n1317_34[2]),.din(w_n1317_11[0]));
	jspl3 jspl3_w_n1317_35(.douta(w_n1317_35[0]),.doutb(w_n1317_35[1]),.doutc(w_n1317_35[2]),.din(w_n1317_11[1]));
	jspl jspl_w_n1317_36(.douta(w_n1317_36[0]),.doutb(w_n1317_36[1]),.din(w_n1317_11[2]));
	jspl3 jspl3_w_n1320_0(.douta(w_n1320_0[0]),.doutb(w_n1320_0[1]),.doutc(w_n1320_0[2]),.din(n1320));
	jspl jspl_w_n1320_1(.douta(w_n1320_1[0]),.doutb(w_n1320_1[1]),.din(w_n1320_0[0]));
	jspl3 jspl3_w_n1321_0(.douta(w_n1321_0[0]),.doutb(w_n1321_0[1]),.doutc(w_n1321_0[2]),.din(n1321));
	jspl3 jspl3_w_n1325_0(.douta(w_n1325_0[0]),.doutb(w_n1325_0[1]),.doutc(w_n1325_0[2]),.din(n1325));
	jspl jspl_w_n1326_0(.douta(w_n1326_0[0]),.doutb(w_n1326_0[1]),.din(n1326));
	jspl jspl_w_n1327_0(.douta(w_n1327_0[0]),.doutb(w_n1327_0[1]),.din(n1327));
	jspl jspl_w_n1328_0(.douta(w_n1328_0[0]),.doutb(w_n1328_0[1]),.din(n1328));
	jspl jspl_w_n1330_0(.douta(w_n1330_0[0]),.doutb(w_n1330_0[1]),.din(n1330));
	jspl jspl_w_n1332_0(.douta(w_n1332_0[0]),.doutb(w_n1332_0[1]),.din(n1332));
	jspl jspl_w_n1334_0(.douta(w_n1334_0[0]),.doutb(w_n1334_0[1]),.din(n1334));
	jspl jspl_w_n1337_0(.douta(w_n1337_0[0]),.doutb(w_n1337_0[1]),.din(n1337));
	jspl jspl_w_n1342_0(.douta(w_n1342_0[0]),.doutb(w_n1342_0[1]),.din(n1342));
	jspl3 jspl3_w_n1344_0(.douta(w_n1344_0[0]),.doutb(w_n1344_0[1]),.doutc(w_n1344_0[2]),.din(n1344));
	jspl jspl_w_n1345_0(.douta(w_n1345_0[0]),.doutb(w_n1345_0[1]),.din(n1345));
	jspl jspl_w_n1349_0(.douta(w_n1349_0[0]),.doutb(w_n1349_0[1]),.din(n1349));
	jspl jspl_w_n1350_0(.douta(w_n1350_0[0]),.doutb(w_n1350_0[1]),.din(n1350));
	jspl jspl_w_n1352_0(.douta(w_n1352_0[0]),.doutb(w_n1352_0[1]),.din(n1352));
	jspl jspl_w_n1356_0(.douta(w_n1356_0[0]),.doutb(w_n1356_0[1]),.din(n1356));
	jspl jspl_w_n1358_0(.douta(w_n1358_0[0]),.doutb(w_n1358_0[1]),.din(n1358));
	jspl jspl_w_n1359_0(.douta(w_n1359_0[0]),.doutb(w_n1359_0[1]),.din(n1359));
	jspl3 jspl3_w_n1360_0(.douta(w_n1360_0[0]),.doutb(w_n1360_0[1]),.doutc(w_n1360_0[2]),.din(n1360));
	jspl jspl_w_n1361_0(.douta(w_n1361_0[0]),.doutb(w_n1361_0[1]),.din(n1361));
	jspl jspl_w_n1365_0(.douta(w_n1365_0[0]),.doutb(w_n1365_0[1]),.din(n1365));
	jspl jspl_w_n1367_0(.douta(w_n1367_0[0]),.doutb(w_n1367_0[1]),.din(n1367));
	jspl jspl_w_n1369_0(.douta(w_n1369_0[0]),.doutb(w_n1369_0[1]),.din(n1369));
	jspl jspl_w_n1371_0(.douta(w_n1371_0[0]),.doutb(w_n1371_0[1]),.din(n1371));
	jspl jspl_w_n1373_0(.douta(w_n1373_0[0]),.doutb(w_n1373_0[1]),.din(n1373));
	jspl jspl_w_n1379_0(.douta(w_n1379_0[0]),.doutb(w_n1379_0[1]),.din(n1379));
	jspl3 jspl3_w_n1381_0(.douta(w_n1381_0[0]),.doutb(w_n1381_0[1]),.doutc(w_n1381_0[2]),.din(n1381));
	jspl jspl_w_n1382_0(.douta(w_n1382_0[0]),.doutb(w_n1382_0[1]),.din(n1382));
	jspl jspl_w_n1387_0(.douta(w_n1387_0[0]),.doutb(w_n1387_0[1]),.din(n1387));
	jspl jspl_w_n1389_0(.douta(w_n1389_0[0]),.doutb(w_n1389_0[1]),.din(n1389));
	jspl jspl_w_n1391_0(.douta(w_n1391_0[0]),.doutb(w_n1391_0[1]),.din(n1391));
	jspl jspl_w_n1395_0(.douta(w_n1395_0[0]),.doutb(w_n1395_0[1]),.din(n1395));
	jspl jspl_w_n1397_0(.douta(w_n1397_0[0]),.doutb(w_n1397_0[1]),.din(n1397));
	jspl jspl_w_n1398_0(.douta(w_n1398_0[0]),.doutb(w_n1398_0[1]),.din(n1398));
	jspl3 jspl3_w_n1399_0(.douta(w_n1399_0[0]),.doutb(w_n1399_0[1]),.doutc(w_n1399_0[2]),.din(n1399));
	jspl jspl_w_n1400_0(.douta(w_n1400_0[0]),.doutb(w_n1400_0[1]),.din(n1400));
	jspl jspl_w_n1406_0(.douta(w_n1406_0[0]),.doutb(w_n1406_0[1]),.din(n1406));
	jspl jspl_w_n1407_0(.douta(w_n1407_0[0]),.doutb(w_n1407_0[1]),.din(n1407));
	jspl jspl_w_n1409_0(.douta(w_n1409_0[0]),.doutb(w_n1409_0[1]),.din(n1409));
	jspl jspl_w_n1411_0(.douta(w_n1411_0[0]),.doutb(w_n1411_0[1]),.din(n1411));
	jspl jspl_w_n1413_0(.douta(w_n1413_0[0]),.doutb(w_n1413_0[1]),.din(n1413));
	jspl jspl_w_n1419_0(.douta(w_n1419_0[0]),.doutb(w_n1419_0[1]),.din(n1419));
	jspl jspl_w_n1421_0(.douta(w_n1421_0[0]),.doutb(w_n1421_0[1]),.din(n1421));
	jspl3 jspl3_w_n1422_0(.douta(w_n1422_0[0]),.doutb(w_n1422_0[1]),.doutc(w_n1422_0[2]),.din(n1422));
	jspl jspl_w_n1425_0(.douta(w_n1425_0[0]),.doutb(w_n1425_0[1]),.din(n1425));
	jspl jspl_w_n1426_0(.douta(w_n1426_0[0]),.doutb(w_n1426_0[1]),.din(n1426));
	jspl3 jspl3_w_n1427_0(.douta(w_n1427_0[0]),.doutb(w_n1427_0[1]),.doutc(w_n1427_0[2]),.din(n1427));
	jspl jspl_w_n1429_0(.douta(w_n1429_0[0]),.doutb(w_n1429_0[1]),.din(n1429));
	jspl jspl_w_n1433_0(.douta(w_n1433_0[0]),.doutb(w_n1433_0[1]),.din(n1433));
	jspl jspl_w_n1435_0(.douta(w_n1435_0[0]),.doutb(w_n1435_0[1]),.din(n1435));
	jspl jspl_w_n1436_0(.douta(w_n1436_0[0]),.doutb(w_n1436_0[1]),.din(n1436));
	jspl3 jspl3_w_n1437_0(.douta(w_n1437_0[0]),.doutb(w_n1437_0[1]),.doutc(w_n1437_0[2]),.din(n1437));
	jspl jspl_w_n1441_0(.douta(w_n1441_0[0]),.doutb(w_n1441_0[1]),.din(n1441));
	jspl jspl_w_n1447_0(.douta(w_n1447_0[0]),.doutb(w_n1447_0[1]),.din(n1447));
	jspl3 jspl3_w_n1449_0(.douta(w_n1449_0[0]),.doutb(w_n1449_0[1]),.doutc(w_n1449_0[2]),.din(n1449));
	jspl jspl_w_n1451_0(.douta(w_n1451_0[0]),.doutb(w_n1451_0[1]),.din(n1451));
	jspl3 jspl3_w_n1456_0(.douta(w_n1456_0[0]),.doutb(w_n1456_0[1]),.doutc(w_n1456_0[2]),.din(n1456));
	jspl jspl_w_n1457_0(.douta(w_n1457_0[0]),.doutb(w_n1457_0[1]),.din(n1457));
	jspl jspl_w_n1458_0(.douta(w_n1458_0[0]),.doutb(w_n1458_0[1]),.din(n1458));
	jspl jspl_w_n1463_0(.douta(w_n1463_0[0]),.doutb(w_n1463_0[1]),.din(n1463));
	jspl3 jspl3_w_n1464_0(.douta(w_n1464_0[0]),.doutb(w_n1464_0[1]),.doutc(w_n1464_0[2]),.din(n1464));
	jspl jspl_w_n1469_0(.douta(w_n1469_0[0]),.doutb(w_n1469_0[1]),.din(n1469));
	jspl3 jspl3_w_n1475_0(.douta(w_n1475_0[0]),.doutb(w_n1475_0[1]),.doutc(w_n1475_0[2]),.din(n1475));
	jspl jspl_w_n1475_1(.douta(w_n1475_1[0]),.doutb(w_n1475_1[1]),.din(w_n1475_0[0]));
	jspl jspl_w_n1476_0(.douta(w_n1476_0[0]),.doutb(w_n1476_0[1]),.din(n1476));
	jspl3 jspl3_w_n1479_0(.douta(w_n1479_0[0]),.doutb(w_n1479_0[1]),.doutc(w_n1479_0[2]),.din(n1479));
	jspl jspl_w_n1480_0(.douta(w_n1480_0[0]),.doutb(w_n1480_0[1]),.din(n1480));
	jspl jspl_w_n1481_0(.douta(w_n1481_0[0]),.doutb(w_n1481_0[1]),.din(n1481));
	jspl jspl_w_n1482_0(.douta(w_n1482_0[0]),.doutb(w_n1482_0[1]),.din(n1482));
	jspl jspl_w_n1484_0(.douta(w_n1484_0[0]),.doutb(w_n1484_0[1]),.din(n1484));
	jspl jspl_w_n1486_0(.douta(w_n1486_0[0]),.doutb(w_n1486_0[1]),.din(n1486));
	jspl jspl_w_n1488_0(.douta(w_n1488_0[0]),.doutb(w_n1488_0[1]),.din(n1488));
	jspl jspl_w_n1497_0(.douta(w_n1497_0[0]),.doutb(w_n1497_0[1]),.din(n1497));
	jspl3 jspl3_w_n1499_0(.douta(w_n1499_0[0]),.doutb(w_n1499_0[1]),.doutc(w_n1499_0[2]),.din(n1499));
	jspl jspl_w_n1500_0(.douta(w_n1500_0[0]),.doutb(w_n1500_0[1]),.din(n1500));
	jspl jspl_w_n1504_0(.douta(w_n1504_0[0]),.doutb(w_n1504_0[1]),.din(n1504));
	jspl jspl_w_n1506_0(.douta(w_n1506_0[0]),.doutb(w_n1506_0[1]),.din(n1506));
	jspl jspl_w_n1508_0(.douta(w_n1508_0[0]),.doutb(w_n1508_0[1]),.din(n1508));
	jspl jspl_w_n1513_0(.douta(w_n1513_0[0]),.doutb(w_n1513_0[1]),.din(n1513));
	jspl jspl_w_n1515_0(.douta(w_n1515_0[0]),.doutb(w_n1515_0[1]),.din(n1515));
	jspl jspl_w_n1516_0(.douta(w_n1516_0[0]),.doutb(w_n1516_0[1]),.din(n1516));
	jspl3 jspl3_w_n1517_0(.douta(w_n1517_0[0]),.doutb(w_n1517_0[1]),.doutc(w_n1517_0[2]),.din(n1517));
	jspl jspl_w_n1518_0(.douta(w_n1518_0[0]),.doutb(w_n1518_0[1]),.din(n1518));
	jspl jspl_w_n1523_0(.douta(w_n1523_0[0]),.doutb(w_n1523_0[1]),.din(n1523));
	jspl jspl_w_n1524_0(.douta(w_n1524_0[0]),.doutb(w_n1524_0[1]),.din(n1524));
	jspl jspl_w_n1526_0(.douta(w_n1526_0[0]),.doutb(w_n1526_0[1]),.din(n1526));
	jspl jspl_w_n1528_0(.douta(w_n1528_0[0]),.doutb(w_n1528_0[1]),.din(n1528));
	jspl jspl_w_n1531_0(.douta(w_n1531_0[0]),.doutb(w_n1531_0[1]),.din(n1531));
	jspl jspl_w_n1537_0(.douta(w_n1537_0[0]),.doutb(w_n1537_0[1]),.din(n1537));
	jspl3 jspl3_w_n1539_0(.douta(w_n1539_0[0]),.doutb(w_n1539_0[1]),.doutc(w_n1539_0[2]),.din(n1539));
	jspl jspl_w_n1540_0(.douta(w_n1540_0[0]),.doutb(w_n1540_0[1]),.din(n1540));
	jspl jspl_w_n1544_0(.douta(w_n1544_0[0]),.doutb(w_n1544_0[1]),.din(n1544));
	jspl jspl_w_n1545_0(.douta(w_n1545_0[0]),.doutb(w_n1545_0[1]),.din(n1545));
	jspl jspl_w_n1547_0(.douta(w_n1547_0[0]),.doutb(w_n1547_0[1]),.din(n1547));
	jspl jspl_w_n1552_0(.douta(w_n1552_0[0]),.doutb(w_n1552_0[1]),.din(n1552));
	jspl jspl_w_n1554_0(.douta(w_n1554_0[0]),.doutb(w_n1554_0[1]),.din(n1554));
	jspl jspl_w_n1555_0(.douta(w_n1555_0[0]),.doutb(w_n1555_0[1]),.din(n1555));
	jspl3 jspl3_w_n1556_0(.douta(w_n1556_0[0]),.doutb(w_n1556_0[1]),.doutc(w_n1556_0[2]),.din(n1556));
	jspl jspl_w_n1557_0(.douta(w_n1557_0[0]),.doutb(w_n1557_0[1]),.din(n1557));
	jspl jspl_w_n1561_0(.douta(w_n1561_0[0]),.doutb(w_n1561_0[1]),.din(n1561));
	jspl jspl_w_n1562_0(.douta(w_n1562_0[0]),.doutb(w_n1562_0[1]),.din(n1562));
	jspl jspl_w_n1564_0(.douta(w_n1564_0[0]),.doutb(w_n1564_0[1]),.din(n1564));
	jspl jspl_w_n1566_0(.douta(w_n1566_0[0]),.doutb(w_n1566_0[1]),.din(n1566));
	jspl jspl_w_n1569_0(.douta(w_n1569_0[0]),.doutb(w_n1569_0[1]),.din(n1569));
	jspl jspl_w_n1575_0(.douta(w_n1575_0[0]),.doutb(w_n1575_0[1]),.din(n1575));
	jspl jspl_w_n1577_0(.douta(w_n1577_0[0]),.doutb(w_n1577_0[1]),.din(n1577));
	jspl3 jspl3_w_n1578_0(.douta(w_n1578_0[0]),.doutb(w_n1578_0[1]),.doutc(w_n1578_0[2]),.din(n1578));
	jspl jspl_w_n1582_0(.douta(w_n1582_0[0]),.doutb(w_n1582_0[1]),.din(n1582));
	jspl jspl_w_n1583_0(.douta(w_n1583_0[0]),.doutb(w_n1583_0[1]),.din(n1583));
	jspl3 jspl3_w_n1584_0(.douta(w_n1584_0[0]),.doutb(w_n1584_0[1]),.doutc(w_n1584_0[2]),.din(n1584));
	jspl jspl_w_n1586_0(.douta(w_n1586_0[0]),.doutb(w_n1586_0[1]),.din(n1586));
	jspl jspl_w_n1591_0(.douta(w_n1591_0[0]),.doutb(w_n1591_0[1]),.din(n1591));
	jspl jspl_w_n1593_0(.douta(w_n1593_0[0]),.doutb(w_n1593_0[1]),.din(n1593));
	jspl jspl_w_n1594_0(.douta(w_n1594_0[0]),.doutb(w_n1594_0[1]),.din(n1594));
	jspl3 jspl3_w_n1595_0(.douta(w_n1595_0[0]),.doutb(w_n1595_0[1]),.doutc(w_n1595_0[2]),.din(n1595));
	jspl jspl_w_n1596_0(.douta(w_n1596_0[0]),.doutb(w_n1596_0[1]),.din(n1596));
	jspl jspl_w_n1600_0(.douta(w_n1600_0[0]),.doutb(w_n1600_0[1]),.din(n1600));
	jspl jspl_w_n1606_0(.douta(w_n1606_0[0]),.doutb(w_n1606_0[1]),.din(n1606));
	jspl jspl_w_n1607_0(.douta(w_n1607_0[0]),.doutb(w_n1607_0[1]),.din(n1607));
	jspl jspl_w_n1609_0(.douta(w_n1609_0[0]),.doutb(w_n1609_0[1]),.din(n1609));
	jspl jspl_w_n1611_0(.douta(w_n1611_0[0]),.doutb(w_n1611_0[1]),.din(n1611));
	jspl jspl_w_n1614_0(.douta(w_n1614_0[0]),.doutb(w_n1614_0[1]),.din(n1614));
	jspl jspl_w_n1620_0(.douta(w_n1620_0[0]),.doutb(w_n1620_0[1]),.din(n1620));
	jspl3 jspl3_w_n1622_0(.douta(w_n1622_0[0]),.doutb(w_n1622_0[1]),.doutc(w_n1622_0[2]),.din(n1622));
	jspl3 jspl3_w_n1622_1(.douta(w_n1622_1[0]),.doutb(w_n1622_1[1]),.doutc(w_n1622_1[2]),.din(w_n1622_0[0]));
	jspl jspl_w_n1625_0(.douta(w_n1625_0[0]),.doutb(w_n1625_0[1]),.din(n1625));
	jspl3 jspl3_w_n1626_0(.douta(w_n1626_0[0]),.doutb(w_n1626_0[1]),.doutc(w_n1626_0[2]),.din(n1626));
	jspl jspl_w_n1627_0(.douta(w_n1627_0[0]),.doutb(w_n1627_0[1]),.din(n1627));
	jspl jspl_w_n1633_0(.douta(w_n1633_0[0]),.doutb(w_n1633_0[1]),.din(n1633));
	jspl3 jspl3_w_n1634_0(.douta(w_n1634_0[0]),.doutb(w_n1634_0[1]),.doutc(w_n1634_0[2]),.din(n1634));
	jspl jspl_w_n1635_0(.douta(w_n1635_0[0]),.doutb(w_n1635_0[1]),.din(n1635));
	jspl jspl_w_n1640_0(.douta(w_n1640_0[0]),.doutb(w_n1640_0[1]),.din(n1640));
	jspl3 jspl3_w_n1641_0(.douta(w_n1641_0[0]),.doutb(w_n1641_0[1]),.doutc(w_n1641_0[2]),.din(n1641));
	jspl3 jspl3_w_n1641_1(.douta(w_n1641_1[0]),.doutb(w_n1641_1[1]),.doutc(w_n1641_1[2]),.din(w_n1641_0[0]));
	jspl3 jspl3_w_n1641_2(.douta(w_n1641_2[0]),.doutb(w_n1641_2[1]),.doutc(w_n1641_2[2]),.din(w_n1641_0[1]));
	jspl3 jspl3_w_n1641_3(.douta(w_n1641_3[0]),.doutb(w_n1641_3[1]),.doutc(w_n1641_3[2]),.din(w_n1641_0[2]));
	jspl3 jspl3_w_n1641_4(.douta(w_n1641_4[0]),.doutb(w_n1641_4[1]),.doutc(w_n1641_4[2]),.din(w_n1641_1[0]));
	jspl3 jspl3_w_n1641_5(.douta(w_n1641_5[0]),.doutb(w_n1641_5[1]),.doutc(w_n1641_5[2]),.din(w_n1641_1[1]));
	jspl3 jspl3_w_n1641_6(.douta(w_n1641_6[0]),.doutb(w_n1641_6[1]),.doutc(w_n1641_6[2]),.din(w_n1641_1[2]));
	jspl3 jspl3_w_n1641_7(.douta(w_n1641_7[0]),.doutb(w_n1641_7[1]),.doutc(w_n1641_7[2]),.din(w_n1641_2[0]));
	jspl3 jspl3_w_n1641_8(.douta(w_n1641_8[0]),.doutb(w_n1641_8[1]),.doutc(w_n1641_8[2]),.din(w_n1641_2[1]));
	jspl3 jspl3_w_n1641_9(.douta(w_n1641_9[0]),.doutb(w_n1641_9[1]),.doutc(w_n1641_9[2]),.din(w_n1641_2[2]));
	jspl3 jspl3_w_n1641_10(.douta(w_n1641_10[0]),.doutb(w_n1641_10[1]),.doutc(w_n1641_10[2]),.din(w_n1641_3[0]));
	jspl3 jspl3_w_n1641_11(.douta(w_n1641_11[0]),.doutb(w_n1641_11[1]),.doutc(w_n1641_11[2]),.din(w_n1641_3[1]));
	jspl3 jspl3_w_n1641_12(.douta(w_n1641_12[0]),.doutb(w_n1641_12[1]),.doutc(w_n1641_12[2]),.din(w_n1641_3[2]));
	jspl3 jspl3_w_n1641_13(.douta(w_n1641_13[0]),.doutb(w_n1641_13[1]),.doutc(w_n1641_13[2]),.din(w_n1641_4[0]));
	jspl3 jspl3_w_n1641_14(.douta(w_n1641_14[0]),.doutb(w_n1641_14[1]),.doutc(w_n1641_14[2]),.din(w_n1641_4[1]));
	jspl3 jspl3_w_n1641_15(.douta(w_n1641_15[0]),.doutb(w_n1641_15[1]),.doutc(w_n1641_15[2]),.din(w_n1641_4[2]));
	jspl3 jspl3_w_n1641_16(.douta(w_n1641_16[0]),.doutb(w_n1641_16[1]),.doutc(w_n1641_16[2]),.din(w_n1641_5[0]));
	jspl3 jspl3_w_n1641_17(.douta(w_n1641_17[0]),.doutb(w_n1641_17[1]),.doutc(w_n1641_17[2]),.din(w_n1641_5[1]));
	jspl3 jspl3_w_n1641_18(.douta(w_n1641_18[0]),.doutb(w_n1641_18[1]),.doutc(w_n1641_18[2]),.din(w_n1641_5[2]));
	jspl3 jspl3_w_n1641_19(.douta(w_n1641_19[0]),.doutb(w_n1641_19[1]),.doutc(w_n1641_19[2]),.din(w_n1641_6[0]));
	jspl3 jspl3_w_n1641_20(.douta(w_n1641_20[0]),.doutb(w_n1641_20[1]),.doutc(w_n1641_20[2]),.din(w_n1641_6[1]));
	jspl3 jspl3_w_n1641_21(.douta(w_n1641_21[0]),.doutb(w_n1641_21[1]),.doutc(w_n1641_21[2]),.din(w_n1641_6[2]));
	jspl3 jspl3_w_n1641_22(.douta(w_n1641_22[0]),.doutb(w_n1641_22[1]),.doutc(w_n1641_22[2]),.din(w_n1641_7[0]));
	jspl3 jspl3_w_n1641_23(.douta(w_n1641_23[0]),.doutb(w_n1641_23[1]),.doutc(w_n1641_23[2]),.din(w_n1641_7[1]));
	jspl3 jspl3_w_n1641_24(.douta(w_n1641_24[0]),.doutb(w_n1641_24[1]),.doutc(w_n1641_24[2]),.din(w_n1641_7[2]));
	jspl3 jspl3_w_n1641_25(.douta(w_n1641_25[0]),.doutb(w_n1641_25[1]),.doutc(w_n1641_25[2]),.din(w_n1641_8[0]));
	jspl3 jspl3_w_n1641_26(.douta(w_n1641_26[0]),.doutb(w_n1641_26[1]),.doutc(w_n1641_26[2]),.din(w_n1641_8[1]));
	jspl3 jspl3_w_n1641_27(.douta(w_n1641_27[0]),.doutb(w_n1641_27[1]),.doutc(w_n1641_27[2]),.din(w_n1641_8[2]));
	jspl3 jspl3_w_n1641_28(.douta(w_n1641_28[0]),.doutb(w_n1641_28[1]),.doutc(w_n1641_28[2]),.din(w_n1641_9[0]));
	jspl3 jspl3_w_n1641_29(.douta(w_n1641_29[0]),.doutb(w_n1641_29[1]),.doutc(w_n1641_29[2]),.din(w_n1641_9[1]));
	jspl3 jspl3_w_n1641_30(.douta(w_n1641_30[0]),.doutb(w_n1641_30[1]),.doutc(w_n1641_30[2]),.din(w_n1641_9[2]));
	jspl3 jspl3_w_n1646_0(.douta(w_n1646_0[0]),.doutb(w_n1646_0[1]),.doutc(w_n1646_0[2]),.din(n1646));
	jspl3 jspl3_w_n1646_1(.douta(w_n1646_1[0]),.doutb(w_n1646_1[1]),.doutc(w_n1646_1[2]),.din(w_n1646_0[0]));
	jspl3 jspl3_w_n1646_2(.douta(w_n1646_2[0]),.doutb(w_n1646_2[1]),.doutc(w_n1646_2[2]),.din(w_n1646_0[1]));
	jspl3 jspl3_w_n1646_3(.douta(w_n1646_3[0]),.doutb(w_n1646_3[1]),.doutc(w_n1646_3[2]),.din(w_n1646_0[2]));
	jspl3 jspl3_w_n1646_4(.douta(w_n1646_4[0]),.doutb(w_n1646_4[1]),.doutc(w_n1646_4[2]),.din(w_n1646_1[0]));
	jspl3 jspl3_w_n1646_5(.douta(w_n1646_5[0]),.doutb(w_n1646_5[1]),.doutc(w_n1646_5[2]),.din(w_n1646_1[1]));
	jspl3 jspl3_w_n1646_6(.douta(w_n1646_6[0]),.doutb(w_n1646_6[1]),.doutc(w_n1646_6[2]),.din(w_n1646_1[2]));
	jspl3 jspl3_w_n1646_7(.douta(w_n1646_7[0]),.doutb(w_n1646_7[1]),.doutc(w_n1646_7[2]),.din(w_n1646_2[0]));
	jspl3 jspl3_w_n1646_8(.douta(w_n1646_8[0]),.doutb(w_n1646_8[1]),.doutc(w_n1646_8[2]),.din(w_n1646_2[1]));
	jspl3 jspl3_w_n1646_9(.douta(w_n1646_9[0]),.doutb(w_n1646_9[1]),.doutc(w_n1646_9[2]),.din(w_n1646_2[2]));
	jspl3 jspl3_w_n1646_10(.douta(w_n1646_10[0]),.doutb(w_n1646_10[1]),.doutc(w_n1646_10[2]),.din(w_n1646_3[0]));
	jspl3 jspl3_w_n1646_11(.douta(w_n1646_11[0]),.doutb(w_n1646_11[1]),.doutc(w_n1646_11[2]),.din(w_n1646_3[1]));
	jspl3 jspl3_w_n1646_12(.douta(w_n1646_12[0]),.doutb(w_n1646_12[1]),.doutc(w_n1646_12[2]),.din(w_n1646_3[2]));
	jspl3 jspl3_w_n1646_13(.douta(w_n1646_13[0]),.doutb(w_n1646_13[1]),.doutc(w_n1646_13[2]),.din(w_n1646_4[0]));
	jspl3 jspl3_w_n1646_14(.douta(w_n1646_14[0]),.doutb(w_n1646_14[1]),.doutc(w_n1646_14[2]),.din(w_n1646_4[1]));
	jspl3 jspl3_w_n1646_15(.douta(w_n1646_15[0]),.doutb(w_n1646_15[1]),.doutc(w_n1646_15[2]),.din(w_n1646_4[2]));
	jspl3 jspl3_w_n1646_16(.douta(w_n1646_16[0]),.doutb(w_n1646_16[1]),.doutc(w_n1646_16[2]),.din(w_n1646_5[0]));
	jspl3 jspl3_w_n1646_17(.douta(w_n1646_17[0]),.doutb(w_n1646_17[1]),.doutc(w_n1646_17[2]),.din(w_n1646_5[1]));
	jspl3 jspl3_w_n1646_18(.douta(w_n1646_18[0]),.doutb(w_n1646_18[1]),.doutc(w_n1646_18[2]),.din(w_n1646_5[2]));
	jspl3 jspl3_w_n1646_19(.douta(w_n1646_19[0]),.doutb(w_n1646_19[1]),.doutc(w_n1646_19[2]),.din(w_n1646_6[0]));
	jspl3 jspl3_w_n1646_20(.douta(w_n1646_20[0]),.doutb(w_n1646_20[1]),.doutc(w_n1646_20[2]),.din(w_n1646_6[1]));
	jspl3 jspl3_w_n1646_21(.douta(w_n1646_21[0]),.doutb(w_n1646_21[1]),.doutc(w_n1646_21[2]),.din(w_n1646_6[2]));
	jspl3 jspl3_w_n1646_22(.douta(w_n1646_22[0]),.doutb(w_n1646_22[1]),.doutc(w_n1646_22[2]),.din(w_n1646_7[0]));
	jspl3 jspl3_w_n1646_23(.douta(w_n1646_23[0]),.doutb(w_n1646_23[1]),.doutc(w_n1646_23[2]),.din(w_n1646_7[1]));
	jspl3 jspl3_w_n1646_24(.douta(w_n1646_24[0]),.doutb(w_n1646_24[1]),.doutc(w_n1646_24[2]),.din(w_n1646_7[2]));
	jspl3 jspl3_w_n1646_25(.douta(w_n1646_25[0]),.doutb(w_n1646_25[1]),.doutc(w_n1646_25[2]),.din(w_n1646_8[0]));
	jspl3 jspl3_w_n1646_26(.douta(w_n1646_26[0]),.doutb(w_n1646_26[1]),.doutc(w_n1646_26[2]),.din(w_n1646_8[1]));
	jspl3 jspl3_w_n1646_27(.douta(w_n1646_27[0]),.doutb(w_n1646_27[1]),.doutc(w_n1646_27[2]),.din(w_n1646_8[2]));
	jspl3 jspl3_w_n1646_28(.douta(w_n1646_28[0]),.doutb(w_n1646_28[1]),.doutc(w_n1646_28[2]),.din(w_n1646_9[0]));
	jspl3 jspl3_w_n1646_29(.douta(w_n1646_29[0]),.doutb(w_n1646_29[1]),.doutc(w_n1646_29[2]),.din(w_n1646_9[1]));
	jspl3 jspl3_w_n1646_30(.douta(w_n1646_30[0]),.doutb(w_n1646_30[1]),.doutc(w_n1646_30[2]),.din(w_n1646_9[2]));
	jspl3 jspl3_w_n1646_31(.douta(w_n1646_31[0]),.doutb(w_n1646_31[1]),.doutc(w_n1646_31[2]),.din(w_n1646_10[0]));
	jspl3 jspl3_w_n1646_32(.douta(w_n1646_32[0]),.doutb(w_n1646_32[1]),.doutc(w_n1646_32[2]),.din(w_n1646_10[1]));
	jspl3 jspl3_w_n1646_33(.douta(w_n1646_33[0]),.doutb(w_n1646_33[1]),.doutc(w_n1646_33[2]),.din(w_n1646_10[2]));
	jspl3 jspl3_w_n1646_34(.douta(w_n1646_34[0]),.doutb(w_n1646_34[1]),.doutc(w_n1646_34[2]),.din(w_n1646_11[0]));
	jspl3 jspl3_w_n1646_35(.douta(w_n1646_35[0]),.doutb(w_n1646_35[1]),.doutc(w_n1646_35[2]),.din(w_n1646_11[1]));
	jspl jspl_w_n1646_36(.douta(w_n1646_36[0]),.doutb(w_n1646_36[1]),.din(w_n1646_11[2]));
	jspl3 jspl3_w_n1649_0(.douta(w_n1649_0[0]),.doutb(w_n1649_0[1]),.doutc(w_n1649_0[2]),.din(n1649));
	jspl jspl_w_n1649_1(.douta(w_n1649_1[0]),.doutb(w_n1649_1[1]),.din(w_n1649_0[0]));
	jspl3 jspl3_w_n1650_0(.douta(w_n1650_0[0]),.doutb(w_n1650_0[1]),.doutc(w_n1650_0[2]),.din(n1650));
	jspl3 jspl3_w_n1654_0(.douta(w_n1654_0[0]),.doutb(w_n1654_0[1]),.doutc(w_n1654_0[2]),.din(n1654));
	jspl jspl_w_n1655_0(.douta(w_n1655_0[0]),.doutb(w_n1655_0[1]),.din(n1655));
	jspl jspl_w_n1656_0(.douta(w_n1656_0[0]),.doutb(w_n1656_0[1]),.din(n1656));
	jspl jspl_w_n1657_0(.douta(w_n1657_0[0]),.doutb(w_n1657_0[1]),.din(n1657));
	jspl jspl_w_n1659_0(.douta(w_n1659_0[0]),.doutb(w_n1659_0[1]),.din(n1659));
	jspl jspl_w_n1661_0(.douta(w_n1661_0[0]),.doutb(w_n1661_0[1]),.din(n1661));
	jspl jspl_w_n1663_0(.douta(w_n1663_0[0]),.doutb(w_n1663_0[1]),.din(n1663));
	jspl jspl_w_n1666_0(.douta(w_n1666_0[0]),.doutb(w_n1666_0[1]),.din(n1666));
	jspl jspl_w_n1671_0(.douta(w_n1671_0[0]),.doutb(w_n1671_0[1]),.din(n1671));
	jspl3 jspl3_w_n1673_0(.douta(w_n1673_0[0]),.doutb(w_n1673_0[1]),.doutc(w_n1673_0[2]),.din(n1673));
	jspl jspl_w_n1674_0(.douta(w_n1674_0[0]),.doutb(w_n1674_0[1]),.din(n1674));
	jspl jspl_w_n1678_0(.douta(w_n1678_0[0]),.doutb(w_n1678_0[1]),.din(n1678));
	jspl jspl_w_n1679_0(.douta(w_n1679_0[0]),.doutb(w_n1679_0[1]),.din(n1679));
	jspl jspl_w_n1681_0(.douta(w_n1681_0[0]),.doutb(w_n1681_0[1]),.din(n1681));
	jspl jspl_w_n1685_0(.douta(w_n1685_0[0]),.doutb(w_n1685_0[1]),.din(n1685));
	jspl jspl_w_n1687_0(.douta(w_n1687_0[0]),.doutb(w_n1687_0[1]),.din(n1687));
	jspl jspl_w_n1688_0(.douta(w_n1688_0[0]),.doutb(w_n1688_0[1]),.din(n1688));
	jspl3 jspl3_w_n1689_0(.douta(w_n1689_0[0]),.doutb(w_n1689_0[1]),.doutc(w_n1689_0[2]),.din(n1689));
	jspl jspl_w_n1690_0(.douta(w_n1690_0[0]),.doutb(w_n1690_0[1]),.din(n1690));
	jspl jspl_w_n1694_0(.douta(w_n1694_0[0]),.doutb(w_n1694_0[1]),.din(n1694));
	jspl jspl_w_n1696_0(.douta(w_n1696_0[0]),.doutb(w_n1696_0[1]),.din(n1696));
	jspl jspl_w_n1698_0(.douta(w_n1698_0[0]),.doutb(w_n1698_0[1]),.din(n1698));
	jspl jspl_w_n1700_0(.douta(w_n1700_0[0]),.doutb(w_n1700_0[1]),.din(n1700));
	jspl jspl_w_n1702_0(.douta(w_n1702_0[0]),.doutb(w_n1702_0[1]),.din(n1702));
	jspl jspl_w_n1708_0(.douta(w_n1708_0[0]),.doutb(w_n1708_0[1]),.din(n1708));
	jspl3 jspl3_w_n1710_0(.douta(w_n1710_0[0]),.doutb(w_n1710_0[1]),.doutc(w_n1710_0[2]),.din(n1710));
	jspl jspl_w_n1711_0(.douta(w_n1711_0[0]),.doutb(w_n1711_0[1]),.din(n1711));
	jspl jspl_w_n1716_0(.douta(w_n1716_0[0]),.doutb(w_n1716_0[1]),.din(n1716));
	jspl jspl_w_n1718_0(.douta(w_n1718_0[0]),.doutb(w_n1718_0[1]),.din(n1718));
	jspl jspl_w_n1720_0(.douta(w_n1720_0[0]),.doutb(w_n1720_0[1]),.din(n1720));
	jspl jspl_w_n1724_0(.douta(w_n1724_0[0]),.doutb(w_n1724_0[1]),.din(n1724));
	jspl jspl_w_n1726_0(.douta(w_n1726_0[0]),.doutb(w_n1726_0[1]),.din(n1726));
	jspl jspl_w_n1727_0(.douta(w_n1727_0[0]),.doutb(w_n1727_0[1]),.din(n1727));
	jspl3 jspl3_w_n1728_0(.douta(w_n1728_0[0]),.doutb(w_n1728_0[1]),.doutc(w_n1728_0[2]),.din(n1728));
	jspl jspl_w_n1729_0(.douta(w_n1729_0[0]),.doutb(w_n1729_0[1]),.din(n1729));
	jspl jspl_w_n1735_0(.douta(w_n1735_0[0]),.doutb(w_n1735_0[1]),.din(n1735));
	jspl jspl_w_n1736_0(.douta(w_n1736_0[0]),.doutb(w_n1736_0[1]),.din(n1736));
	jspl jspl_w_n1738_0(.douta(w_n1738_0[0]),.doutb(w_n1738_0[1]),.din(n1738));
	jspl jspl_w_n1740_0(.douta(w_n1740_0[0]),.doutb(w_n1740_0[1]),.din(n1740));
	jspl jspl_w_n1742_0(.douta(w_n1742_0[0]),.doutb(w_n1742_0[1]),.din(n1742));
	jspl jspl_w_n1748_0(.douta(w_n1748_0[0]),.doutb(w_n1748_0[1]),.din(n1748));
	jspl jspl_w_n1750_0(.douta(w_n1750_0[0]),.doutb(w_n1750_0[1]),.din(n1750));
	jspl3 jspl3_w_n1751_0(.douta(w_n1751_0[0]),.doutb(w_n1751_0[1]),.doutc(w_n1751_0[2]),.din(n1751));
	jspl jspl_w_n1754_0(.douta(w_n1754_0[0]),.doutb(w_n1754_0[1]),.din(n1754));
	jspl jspl_w_n1755_0(.douta(w_n1755_0[0]),.doutb(w_n1755_0[1]),.din(n1755));
	jspl3 jspl3_w_n1756_0(.douta(w_n1756_0[0]),.doutb(w_n1756_0[1]),.doutc(w_n1756_0[2]),.din(n1756));
	jspl jspl_w_n1758_0(.douta(w_n1758_0[0]),.doutb(w_n1758_0[1]),.din(n1758));
	jspl jspl_w_n1762_0(.douta(w_n1762_0[0]),.doutb(w_n1762_0[1]),.din(n1762));
	jspl jspl_w_n1764_0(.douta(w_n1764_0[0]),.doutb(w_n1764_0[1]),.din(n1764));
	jspl jspl_w_n1765_0(.douta(w_n1765_0[0]),.doutb(w_n1765_0[1]),.din(n1765));
	jspl3 jspl3_w_n1766_0(.douta(w_n1766_0[0]),.doutb(w_n1766_0[1]),.doutc(w_n1766_0[2]),.din(n1766));
	jspl jspl_w_n1767_0(.douta(w_n1767_0[0]),.doutb(w_n1767_0[1]),.din(n1767));
	jspl jspl_w_n1770_0(.douta(w_n1770_0[0]),.doutb(w_n1770_0[1]),.din(n1770));
	jspl jspl_w_n1776_0(.douta(w_n1776_0[0]),.doutb(w_n1776_0[1]),.din(n1776));
	jspl jspl_w_n1777_0(.douta(w_n1777_0[0]),.doutb(w_n1777_0[1]),.din(n1777));
	jspl jspl_w_n1779_0(.douta(w_n1779_0[0]),.doutb(w_n1779_0[1]),.din(n1779));
	jspl jspl_w_n1781_0(.douta(w_n1781_0[0]),.doutb(w_n1781_0[1]),.din(n1781));
	jspl jspl_w_n1783_0(.douta(w_n1783_0[0]),.doutb(w_n1783_0[1]),.din(n1783));
	jspl jspl_w_n1789_0(.douta(w_n1789_0[0]),.doutb(w_n1789_0[1]),.din(n1789));
	jspl3 jspl3_w_n1791_0(.douta(w_n1791_0[0]),.doutb(w_n1791_0[1]),.doutc(w_n1791_0[2]),.din(n1791));
	jspl jspl_w_n1796_0(.douta(w_n1796_0[0]),.doutb(w_n1796_0[1]),.din(n1796));
	jspl3 jspl3_w_n1798_0(.douta(w_n1798_0[0]),.doutb(w_n1798_0[1]),.doutc(w_n1798_0[2]),.din(n1798));
	jspl3 jspl3_w_n1802_0(.douta(w_n1802_0[0]),.doutb(w_n1802_0[1]),.doutc(w_n1802_0[2]),.din(n1802));
	jspl jspl_w_n1803_0(.douta(w_n1803_0[0]),.doutb(w_n1803_0[1]),.din(n1803));
	jspl jspl_w_n1808_0(.douta(w_n1808_0[0]),.doutb(w_n1808_0[1]),.din(n1808));
	jspl3 jspl3_w_n1809_0(.douta(w_n1809_0[0]),.doutb(w_n1809_0[1]),.doutc(w_n1809_0[2]),.din(n1809));
	jspl jspl_w_n1814_0(.douta(w_n1814_0[0]),.doutb(w_n1814_0[1]),.din(n1814));
	jspl3 jspl3_w_n1820_0(.douta(w_n1820_0[0]),.doutb(w_n1820_0[1]),.doutc(w_n1820_0[2]),.din(n1820));
	jspl jspl_w_n1820_1(.douta(w_n1820_1[0]),.doutb(w_n1820_1[1]),.din(w_n1820_0[0]));
	jspl jspl_w_n1821_0(.douta(w_n1821_0[0]),.doutb(w_n1821_0[1]),.din(n1821));
	jspl3 jspl3_w_n1824_0(.douta(w_n1824_0[0]),.doutb(w_n1824_0[1]),.doutc(w_n1824_0[2]),.din(n1824));
	jspl jspl_w_n1825_0(.douta(w_n1825_0[0]),.doutb(w_n1825_0[1]),.din(n1825));
	jspl jspl_w_n1826_0(.douta(w_n1826_0[0]),.doutb(w_n1826_0[1]),.din(n1826));
	jspl jspl_w_n1827_0(.douta(w_n1827_0[0]),.doutb(w_n1827_0[1]),.din(n1827));
	jspl jspl_w_n1829_0(.douta(w_n1829_0[0]),.doutb(w_n1829_0[1]),.din(n1829));
	jspl jspl_w_n1831_0(.douta(w_n1831_0[0]),.doutb(w_n1831_0[1]),.din(n1831));
	jspl jspl_w_n1833_0(.douta(w_n1833_0[0]),.doutb(w_n1833_0[1]),.din(n1833));
	jspl jspl_w_n1842_0(.douta(w_n1842_0[0]),.doutb(w_n1842_0[1]),.din(n1842));
	jspl3 jspl3_w_n1844_0(.douta(w_n1844_0[0]),.doutb(w_n1844_0[1]),.doutc(w_n1844_0[2]),.din(n1844));
	jspl jspl_w_n1845_0(.douta(w_n1845_0[0]),.doutb(w_n1845_0[1]),.din(n1845));
	jspl jspl_w_n1849_0(.douta(w_n1849_0[0]),.doutb(w_n1849_0[1]),.din(n1849));
	jspl jspl_w_n1851_0(.douta(w_n1851_0[0]),.doutb(w_n1851_0[1]),.din(n1851));
	jspl jspl_w_n1853_0(.douta(w_n1853_0[0]),.doutb(w_n1853_0[1]),.din(n1853));
	jspl jspl_w_n1858_0(.douta(w_n1858_0[0]),.doutb(w_n1858_0[1]),.din(n1858));
	jspl jspl_w_n1860_0(.douta(w_n1860_0[0]),.doutb(w_n1860_0[1]),.din(n1860));
	jspl jspl_w_n1861_0(.douta(w_n1861_0[0]),.doutb(w_n1861_0[1]),.din(n1861));
	jspl3 jspl3_w_n1862_0(.douta(w_n1862_0[0]),.doutb(w_n1862_0[1]),.doutc(w_n1862_0[2]),.din(n1862));
	jspl jspl_w_n1863_0(.douta(w_n1863_0[0]),.doutb(w_n1863_0[1]),.din(n1863));
	jspl jspl_w_n1868_0(.douta(w_n1868_0[0]),.doutb(w_n1868_0[1]),.din(n1868));
	jspl jspl_w_n1869_0(.douta(w_n1869_0[0]),.doutb(w_n1869_0[1]),.din(n1869));
	jspl jspl_w_n1871_0(.douta(w_n1871_0[0]),.doutb(w_n1871_0[1]),.din(n1871));
	jspl jspl_w_n1873_0(.douta(w_n1873_0[0]),.doutb(w_n1873_0[1]),.din(n1873));
	jspl jspl_w_n1876_0(.douta(w_n1876_0[0]),.doutb(w_n1876_0[1]),.din(n1876));
	jspl jspl_w_n1882_0(.douta(w_n1882_0[0]),.doutb(w_n1882_0[1]),.din(n1882));
	jspl3 jspl3_w_n1884_0(.douta(w_n1884_0[0]),.doutb(w_n1884_0[1]),.doutc(w_n1884_0[2]),.din(n1884));
	jspl jspl_w_n1885_0(.douta(w_n1885_0[0]),.doutb(w_n1885_0[1]),.din(n1885));
	jspl jspl_w_n1889_0(.douta(w_n1889_0[0]),.doutb(w_n1889_0[1]),.din(n1889));
	jspl jspl_w_n1890_0(.douta(w_n1890_0[0]),.doutb(w_n1890_0[1]),.din(n1890));
	jspl jspl_w_n1892_0(.douta(w_n1892_0[0]),.doutb(w_n1892_0[1]),.din(n1892));
	jspl jspl_w_n1897_0(.douta(w_n1897_0[0]),.doutb(w_n1897_0[1]),.din(n1897));
	jspl jspl_w_n1899_0(.douta(w_n1899_0[0]),.doutb(w_n1899_0[1]),.din(n1899));
	jspl jspl_w_n1900_0(.douta(w_n1900_0[0]),.doutb(w_n1900_0[1]),.din(n1900));
	jspl3 jspl3_w_n1901_0(.douta(w_n1901_0[0]),.doutb(w_n1901_0[1]),.doutc(w_n1901_0[2]),.din(n1901));
	jspl jspl_w_n1902_0(.douta(w_n1902_0[0]),.doutb(w_n1902_0[1]),.din(n1902));
	jspl jspl_w_n1906_0(.douta(w_n1906_0[0]),.doutb(w_n1906_0[1]),.din(n1906));
	jspl jspl_w_n1907_0(.douta(w_n1907_0[0]),.doutb(w_n1907_0[1]),.din(n1907));
	jspl jspl_w_n1909_0(.douta(w_n1909_0[0]),.doutb(w_n1909_0[1]),.din(n1909));
	jspl jspl_w_n1911_0(.douta(w_n1911_0[0]),.doutb(w_n1911_0[1]),.din(n1911));
	jspl jspl_w_n1914_0(.douta(w_n1914_0[0]),.doutb(w_n1914_0[1]),.din(n1914));
	jspl jspl_w_n1920_0(.douta(w_n1920_0[0]),.doutb(w_n1920_0[1]),.din(n1920));
	jspl jspl_w_n1922_0(.douta(w_n1922_0[0]),.doutb(w_n1922_0[1]),.din(n1922));
	jspl3 jspl3_w_n1923_0(.douta(w_n1923_0[0]),.doutb(w_n1923_0[1]),.doutc(w_n1923_0[2]),.din(n1923));
	jspl jspl_w_n1927_0(.douta(w_n1927_0[0]),.doutb(w_n1927_0[1]),.din(n1927));
	jspl jspl_w_n1928_0(.douta(w_n1928_0[0]),.doutb(w_n1928_0[1]),.din(n1928));
	jspl3 jspl3_w_n1929_0(.douta(w_n1929_0[0]),.doutb(w_n1929_0[1]),.doutc(w_n1929_0[2]),.din(n1929));
	jspl jspl_w_n1931_0(.douta(w_n1931_0[0]),.doutb(w_n1931_0[1]),.din(n1931));
	jspl jspl_w_n1936_0(.douta(w_n1936_0[0]),.doutb(w_n1936_0[1]),.din(n1936));
	jspl jspl_w_n1938_0(.douta(w_n1938_0[0]),.doutb(w_n1938_0[1]),.din(n1938));
	jspl jspl_w_n1939_0(.douta(w_n1939_0[0]),.doutb(w_n1939_0[1]),.din(n1939));
	jspl3 jspl3_w_n1940_0(.douta(w_n1940_0[0]),.doutb(w_n1940_0[1]),.doutc(w_n1940_0[2]),.din(n1940));
	jspl jspl_w_n1941_0(.douta(w_n1941_0[0]),.doutb(w_n1941_0[1]),.din(n1941));
	jspl jspl_w_n1945_0(.douta(w_n1945_0[0]),.doutb(w_n1945_0[1]),.din(n1945));
	jspl jspl_w_n1951_0(.douta(w_n1951_0[0]),.doutb(w_n1951_0[1]),.din(n1951));
	jspl jspl_w_n1952_0(.douta(w_n1952_0[0]),.doutb(w_n1952_0[1]),.din(n1952));
	jspl jspl_w_n1954_0(.douta(w_n1954_0[0]),.doutb(w_n1954_0[1]),.din(n1954));
	jspl jspl_w_n1956_0(.douta(w_n1956_0[0]),.doutb(w_n1956_0[1]),.din(n1956));
	jspl jspl_w_n1959_0(.douta(w_n1959_0[0]),.doutb(w_n1959_0[1]),.din(n1959));
	jspl jspl_w_n1965_0(.douta(w_n1965_0[0]),.doutb(w_n1965_0[1]),.din(n1965));
	jspl jspl_w_n1967_0(.douta(w_n1967_0[0]),.doutb(w_n1967_0[1]),.din(n1967));
	jspl3 jspl3_w_n1968_0(.douta(w_n1968_0[0]),.doutb(w_n1968_0[1]),.doutc(w_n1968_0[2]),.din(n1968));
	jspl jspl_w_n1972_0(.douta(w_n1972_0[0]),.doutb(w_n1972_0[1]),.din(n1972));
	jspl jspl_w_n1973_0(.douta(w_n1973_0[0]),.doutb(w_n1973_0[1]),.din(n1973));
	jspl3 jspl3_w_n1974_0(.douta(w_n1974_0[0]),.doutb(w_n1974_0[1]),.doutc(w_n1974_0[2]),.din(n1974));
	jspl jspl_w_n1976_0(.douta(w_n1976_0[0]),.doutb(w_n1976_0[1]),.din(n1976));
	jspl jspl_w_n1981_0(.douta(w_n1981_0[0]),.doutb(w_n1981_0[1]),.din(n1981));
	jspl jspl_w_n1983_0(.douta(w_n1983_0[0]),.doutb(w_n1983_0[1]),.din(n1983));
	jspl jspl_w_n1984_0(.douta(w_n1984_0[0]),.doutb(w_n1984_0[1]),.din(n1984));
	jspl3 jspl3_w_n1985_0(.douta(w_n1985_0[0]),.doutb(w_n1985_0[1]),.doutc(w_n1985_0[2]),.din(n1985));
	jspl3 jspl3_w_n1985_1(.douta(w_n1985_1[0]),.doutb(w_n1985_1[1]),.doutc(w_n1985_1[2]),.din(w_n1985_0[0]));
	jspl jspl_w_n1988_0(.douta(w_n1988_0[0]),.doutb(w_n1988_0[1]),.din(n1988));
	jspl3 jspl3_w_n1989_0(.douta(w_n1989_0[0]),.doutb(w_n1989_0[1]),.doutc(w_n1989_0[2]),.din(n1989));
	jspl jspl_w_n1990_0(.douta(w_n1990_0[0]),.doutb(w_n1990_0[1]),.din(n1990));
	jspl jspl_w_n1991_0(.douta(w_n1991_0[0]),.doutb(w_n1991_0[1]),.din(n1991));
	jspl jspl_w_n1997_0(.douta(w_n1997_0[0]),.doutb(w_n1997_0[1]),.din(n1997));
	jspl3 jspl3_w_n1998_0(.douta(w_n1998_0[0]),.doutb(w_n1998_0[1]),.doutc(w_n1998_0[2]),.din(n1998));
	jspl jspl_w_n1999_0(.douta(w_n1999_0[0]),.doutb(w_n1999_0[1]),.din(n1999));
	jspl jspl_w_n2004_0(.douta(w_n2004_0[0]),.doutb(w_n2004_0[1]),.din(n2004));
	jspl3 jspl3_w_n2005_0(.douta(w_n2005_0[0]),.doutb(w_n2005_0[1]),.doutc(w_n2005_0[2]),.din(n2005));
	jspl3 jspl3_w_n2005_1(.douta(w_n2005_1[0]),.doutb(w_n2005_1[1]),.doutc(w_n2005_1[2]),.din(w_n2005_0[0]));
	jspl3 jspl3_w_n2005_2(.douta(w_n2005_2[0]),.doutb(w_n2005_2[1]),.doutc(w_n2005_2[2]),.din(w_n2005_0[1]));
	jspl3 jspl3_w_n2005_3(.douta(w_n2005_3[0]),.doutb(w_n2005_3[1]),.doutc(w_n2005_3[2]),.din(w_n2005_0[2]));
	jspl3 jspl3_w_n2005_4(.douta(w_n2005_4[0]),.doutb(w_n2005_4[1]),.doutc(w_n2005_4[2]),.din(w_n2005_1[0]));
	jspl3 jspl3_w_n2005_5(.douta(w_n2005_5[0]),.doutb(w_n2005_5[1]),.doutc(w_n2005_5[2]),.din(w_n2005_1[1]));
	jspl3 jspl3_w_n2005_6(.douta(w_n2005_6[0]),.doutb(w_n2005_6[1]),.doutc(w_n2005_6[2]),.din(w_n2005_1[2]));
	jspl3 jspl3_w_n2005_7(.douta(w_n2005_7[0]),.doutb(w_n2005_7[1]),.doutc(w_n2005_7[2]),.din(w_n2005_2[0]));
	jspl3 jspl3_w_n2005_8(.douta(w_n2005_8[0]),.doutb(w_n2005_8[1]),.doutc(w_n2005_8[2]),.din(w_n2005_2[1]));
	jspl3 jspl3_w_n2005_9(.douta(w_n2005_9[0]),.doutb(w_n2005_9[1]),.doutc(w_n2005_9[2]),.din(w_n2005_2[2]));
	jspl3 jspl3_w_n2005_10(.douta(w_n2005_10[0]),.doutb(w_n2005_10[1]),.doutc(w_n2005_10[2]),.din(w_n2005_3[0]));
	jspl3 jspl3_w_n2005_11(.douta(w_n2005_11[0]),.doutb(w_n2005_11[1]),.doutc(w_n2005_11[2]),.din(w_n2005_3[1]));
	jspl3 jspl3_w_n2005_12(.douta(w_n2005_12[0]),.doutb(w_n2005_12[1]),.doutc(w_n2005_12[2]),.din(w_n2005_3[2]));
	jspl3 jspl3_w_n2005_13(.douta(w_n2005_13[0]),.doutb(w_n2005_13[1]),.doutc(w_n2005_13[2]),.din(w_n2005_4[0]));
	jspl3 jspl3_w_n2005_14(.douta(w_n2005_14[0]),.doutb(w_n2005_14[1]),.doutc(w_n2005_14[2]),.din(w_n2005_4[1]));
	jspl3 jspl3_w_n2005_15(.douta(w_n2005_15[0]),.doutb(w_n2005_15[1]),.doutc(w_n2005_15[2]),.din(w_n2005_4[2]));
	jspl3 jspl3_w_n2005_16(.douta(w_n2005_16[0]),.doutb(w_n2005_16[1]),.doutc(w_n2005_16[2]),.din(w_n2005_5[0]));
	jspl3 jspl3_w_n2005_17(.douta(w_n2005_17[0]),.doutb(w_n2005_17[1]),.doutc(w_n2005_17[2]),.din(w_n2005_5[1]));
	jspl3 jspl3_w_n2005_18(.douta(w_n2005_18[0]),.doutb(w_n2005_18[1]),.doutc(w_n2005_18[2]),.din(w_n2005_5[2]));
	jspl3 jspl3_w_n2005_19(.douta(w_n2005_19[0]),.doutb(w_n2005_19[1]),.doutc(w_n2005_19[2]),.din(w_n2005_6[0]));
	jspl3 jspl3_w_n2005_20(.douta(w_n2005_20[0]),.doutb(w_n2005_20[1]),.doutc(w_n2005_20[2]),.din(w_n2005_6[1]));
	jspl3 jspl3_w_n2005_21(.douta(w_n2005_21[0]),.doutb(w_n2005_21[1]),.doutc(w_n2005_21[2]),.din(w_n2005_6[2]));
	jspl3 jspl3_w_n2005_22(.douta(w_n2005_22[0]),.doutb(w_n2005_22[1]),.doutc(w_n2005_22[2]),.din(w_n2005_7[0]));
	jspl3 jspl3_w_n2005_23(.douta(w_n2005_23[0]),.doutb(w_n2005_23[1]),.doutc(w_n2005_23[2]),.din(w_n2005_7[1]));
	jspl3 jspl3_w_n2005_24(.douta(w_n2005_24[0]),.doutb(w_n2005_24[1]),.doutc(w_n2005_24[2]),.din(w_n2005_7[2]));
	jspl3 jspl3_w_n2005_25(.douta(w_n2005_25[0]),.doutb(w_n2005_25[1]),.doutc(w_n2005_25[2]),.din(w_n2005_8[0]));
	jspl3 jspl3_w_n2005_26(.douta(w_n2005_26[0]),.doutb(w_n2005_26[1]),.doutc(w_n2005_26[2]),.din(w_n2005_8[1]));
	jspl3 jspl3_w_n2005_27(.douta(w_n2005_27[0]),.doutb(w_n2005_27[1]),.doutc(w_n2005_27[2]),.din(w_n2005_8[2]));
	jspl3 jspl3_w_n2005_28(.douta(w_n2005_28[0]),.doutb(w_n2005_28[1]),.doutc(w_n2005_28[2]),.din(w_n2005_9[0]));
	jspl jspl_w_n2005_29(.douta(w_n2005_29[0]),.doutb(w_n2005_29[1]),.din(w_n2005_9[1]));
	jspl3 jspl3_w_n2010_0(.douta(w_n2010_0[0]),.doutb(w_n2010_0[1]),.doutc(w_n2010_0[2]),.din(n2010));
	jspl3 jspl3_w_n2010_1(.douta(w_n2010_1[0]),.doutb(w_n2010_1[1]),.doutc(w_n2010_1[2]),.din(w_n2010_0[0]));
	jspl3 jspl3_w_n2010_2(.douta(w_n2010_2[0]),.doutb(w_n2010_2[1]),.doutc(w_n2010_2[2]),.din(w_n2010_0[1]));
	jspl3 jspl3_w_n2010_3(.douta(w_n2010_3[0]),.doutb(w_n2010_3[1]),.doutc(w_n2010_3[2]),.din(w_n2010_0[2]));
	jspl3 jspl3_w_n2010_4(.douta(w_n2010_4[0]),.doutb(w_n2010_4[1]),.doutc(w_n2010_4[2]),.din(w_n2010_1[0]));
	jspl3 jspl3_w_n2010_5(.douta(w_n2010_5[0]),.doutb(w_n2010_5[1]),.doutc(w_n2010_5[2]),.din(w_n2010_1[1]));
	jspl3 jspl3_w_n2010_6(.douta(w_n2010_6[0]),.doutb(w_n2010_6[1]),.doutc(w_n2010_6[2]),.din(w_n2010_1[2]));
	jspl3 jspl3_w_n2010_7(.douta(w_n2010_7[0]),.doutb(w_n2010_7[1]),.doutc(w_n2010_7[2]),.din(w_n2010_2[0]));
	jspl3 jspl3_w_n2010_8(.douta(w_n2010_8[0]),.doutb(w_n2010_8[1]),.doutc(w_n2010_8[2]),.din(w_n2010_2[1]));
	jspl3 jspl3_w_n2010_9(.douta(w_n2010_9[0]),.doutb(w_n2010_9[1]),.doutc(w_n2010_9[2]),.din(w_n2010_2[2]));
	jspl3 jspl3_w_n2010_10(.douta(w_n2010_10[0]),.doutb(w_n2010_10[1]),.doutc(w_n2010_10[2]),.din(w_n2010_3[0]));
	jspl3 jspl3_w_n2010_11(.douta(w_n2010_11[0]),.doutb(w_n2010_11[1]),.doutc(w_n2010_11[2]),.din(w_n2010_3[1]));
	jspl3 jspl3_w_n2010_12(.douta(w_n2010_12[0]),.doutb(w_n2010_12[1]),.doutc(w_n2010_12[2]),.din(w_n2010_3[2]));
	jspl3 jspl3_w_n2010_13(.douta(w_n2010_13[0]),.doutb(w_n2010_13[1]),.doutc(w_n2010_13[2]),.din(w_n2010_4[0]));
	jspl3 jspl3_w_n2010_14(.douta(w_n2010_14[0]),.doutb(w_n2010_14[1]),.doutc(w_n2010_14[2]),.din(w_n2010_4[1]));
	jspl3 jspl3_w_n2010_15(.douta(w_n2010_15[0]),.doutb(w_n2010_15[1]),.doutc(w_n2010_15[2]),.din(w_n2010_4[2]));
	jspl3 jspl3_w_n2010_16(.douta(w_n2010_16[0]),.doutb(w_n2010_16[1]),.doutc(w_n2010_16[2]),.din(w_n2010_5[0]));
	jspl3 jspl3_w_n2010_17(.douta(w_n2010_17[0]),.doutb(w_n2010_17[1]),.doutc(w_n2010_17[2]),.din(w_n2010_5[1]));
	jspl3 jspl3_w_n2010_18(.douta(w_n2010_18[0]),.doutb(w_n2010_18[1]),.doutc(w_n2010_18[2]),.din(w_n2010_5[2]));
	jspl3 jspl3_w_n2010_19(.douta(w_n2010_19[0]),.doutb(w_n2010_19[1]),.doutc(w_n2010_19[2]),.din(w_n2010_6[0]));
	jspl3 jspl3_w_n2010_20(.douta(w_n2010_20[0]),.doutb(w_n2010_20[1]),.doutc(w_n2010_20[2]),.din(w_n2010_6[1]));
	jspl3 jspl3_w_n2010_21(.douta(w_n2010_21[0]),.doutb(w_n2010_21[1]),.doutc(w_n2010_21[2]),.din(w_n2010_6[2]));
	jspl3 jspl3_w_n2010_22(.douta(w_n2010_22[0]),.doutb(w_n2010_22[1]),.doutc(w_n2010_22[2]),.din(w_n2010_7[0]));
	jspl3 jspl3_w_n2010_23(.douta(w_n2010_23[0]),.doutb(w_n2010_23[1]),.doutc(w_n2010_23[2]),.din(w_n2010_7[1]));
	jspl3 jspl3_w_n2010_24(.douta(w_n2010_24[0]),.doutb(w_n2010_24[1]),.doutc(w_n2010_24[2]),.din(w_n2010_7[2]));
	jspl3 jspl3_w_n2010_25(.douta(w_n2010_25[0]),.doutb(w_n2010_25[1]),.doutc(w_n2010_25[2]),.din(w_n2010_8[0]));
	jspl3 jspl3_w_n2010_26(.douta(w_n2010_26[0]),.doutb(w_n2010_26[1]),.doutc(w_n2010_26[2]),.din(w_n2010_8[1]));
	jspl3 jspl3_w_n2010_27(.douta(w_n2010_27[0]),.doutb(w_n2010_27[1]),.doutc(w_n2010_27[2]),.din(w_n2010_8[2]));
	jspl3 jspl3_w_n2010_28(.douta(w_n2010_28[0]),.doutb(w_n2010_28[1]),.doutc(w_n2010_28[2]),.din(w_n2010_9[0]));
	jspl3 jspl3_w_n2010_29(.douta(w_n2010_29[0]),.doutb(w_n2010_29[1]),.doutc(w_n2010_29[2]),.din(w_n2010_9[1]));
	jspl3 jspl3_w_n2010_30(.douta(w_n2010_30[0]),.doutb(w_n2010_30[1]),.doutc(w_n2010_30[2]),.din(w_n2010_9[2]));
	jspl3 jspl3_w_n2010_31(.douta(w_n2010_31[0]),.doutb(w_n2010_31[1]),.doutc(w_n2010_31[2]),.din(w_n2010_10[0]));
	jspl3 jspl3_w_n2010_32(.douta(w_n2010_32[0]),.doutb(w_n2010_32[1]),.doutc(w_n2010_32[2]),.din(w_n2010_10[1]));
	jspl3 jspl3_w_n2010_33(.douta(w_n2010_33[0]),.doutb(w_n2010_33[1]),.doutc(w_n2010_33[2]),.din(w_n2010_10[2]));
	jspl3 jspl3_w_n2010_34(.douta(w_n2010_34[0]),.doutb(w_n2010_34[1]),.doutc(w_n2010_34[2]),.din(w_n2010_11[0]));
	jspl3 jspl3_w_n2013_0(.douta(w_n2013_0[0]),.doutb(w_n2013_0[1]),.doutc(w_n2013_0[2]),.din(n2013));
	jspl jspl_w_n2013_1(.douta(w_n2013_1[0]),.doutb(w_n2013_1[1]),.din(w_n2013_0[0]));
	jspl3 jspl3_w_n2014_0(.douta(w_n2014_0[0]),.doutb(w_n2014_0[1]),.doutc(w_n2014_0[2]),.din(n2014));
	jspl3 jspl3_w_n2018_0(.douta(w_n2018_0[0]),.doutb(w_n2018_0[1]),.doutc(w_n2018_0[2]),.din(n2018));
	jspl jspl_w_n2019_0(.douta(w_n2019_0[0]),.doutb(w_n2019_0[1]),.din(n2019));
	jspl jspl_w_n2020_0(.douta(w_n2020_0[0]),.doutb(w_n2020_0[1]),.din(n2020));
	jspl jspl_w_n2021_0(.douta(w_n2021_0[0]),.doutb(w_n2021_0[1]),.din(n2021));
	jspl jspl_w_n2023_0(.douta(w_n2023_0[0]),.doutb(w_n2023_0[1]),.din(n2023));
	jspl jspl_w_n2025_0(.douta(w_n2025_0[0]),.doutb(w_n2025_0[1]),.din(n2025));
	jspl jspl_w_n2027_0(.douta(w_n2027_0[0]),.doutb(w_n2027_0[1]),.din(n2027));
	jspl jspl_w_n2030_0(.douta(w_n2030_0[0]),.doutb(w_n2030_0[1]),.din(n2030));
	jspl jspl_w_n2035_0(.douta(w_n2035_0[0]),.doutb(w_n2035_0[1]),.din(n2035));
	jspl3 jspl3_w_n2037_0(.douta(w_n2037_0[0]),.doutb(w_n2037_0[1]),.doutc(w_n2037_0[2]),.din(n2037));
	jspl jspl_w_n2038_0(.douta(w_n2038_0[0]),.doutb(w_n2038_0[1]),.din(n2038));
	jspl jspl_w_n2042_0(.douta(w_n2042_0[0]),.doutb(w_n2042_0[1]),.din(n2042));
	jspl jspl_w_n2043_0(.douta(w_n2043_0[0]),.doutb(w_n2043_0[1]),.din(n2043));
	jspl jspl_w_n2045_0(.douta(w_n2045_0[0]),.doutb(w_n2045_0[1]),.din(n2045));
	jspl jspl_w_n2049_0(.douta(w_n2049_0[0]),.doutb(w_n2049_0[1]),.din(n2049));
	jspl jspl_w_n2051_0(.douta(w_n2051_0[0]),.doutb(w_n2051_0[1]),.din(n2051));
	jspl jspl_w_n2052_0(.douta(w_n2052_0[0]),.doutb(w_n2052_0[1]),.din(n2052));
	jspl3 jspl3_w_n2053_0(.douta(w_n2053_0[0]),.doutb(w_n2053_0[1]),.doutc(w_n2053_0[2]),.din(n2053));
	jspl jspl_w_n2054_0(.douta(w_n2054_0[0]),.doutb(w_n2054_0[1]),.din(n2054));
	jspl jspl_w_n2058_0(.douta(w_n2058_0[0]),.doutb(w_n2058_0[1]),.din(n2058));
	jspl jspl_w_n2060_0(.douta(w_n2060_0[0]),.doutb(w_n2060_0[1]),.din(n2060));
	jspl jspl_w_n2062_0(.douta(w_n2062_0[0]),.doutb(w_n2062_0[1]),.din(n2062));
	jspl jspl_w_n2064_0(.douta(w_n2064_0[0]),.doutb(w_n2064_0[1]),.din(n2064));
	jspl jspl_w_n2066_0(.douta(w_n2066_0[0]),.doutb(w_n2066_0[1]),.din(n2066));
	jspl jspl_w_n2072_0(.douta(w_n2072_0[0]),.doutb(w_n2072_0[1]),.din(n2072));
	jspl3 jspl3_w_n2074_0(.douta(w_n2074_0[0]),.doutb(w_n2074_0[1]),.doutc(w_n2074_0[2]),.din(n2074));
	jspl jspl_w_n2075_0(.douta(w_n2075_0[0]),.doutb(w_n2075_0[1]),.din(n2075));
	jspl jspl_w_n2080_0(.douta(w_n2080_0[0]),.doutb(w_n2080_0[1]),.din(n2080));
	jspl jspl_w_n2082_0(.douta(w_n2082_0[0]),.doutb(w_n2082_0[1]),.din(n2082));
	jspl jspl_w_n2084_0(.douta(w_n2084_0[0]),.doutb(w_n2084_0[1]),.din(n2084));
	jspl jspl_w_n2088_0(.douta(w_n2088_0[0]),.doutb(w_n2088_0[1]),.din(n2088));
	jspl jspl_w_n2090_0(.douta(w_n2090_0[0]),.doutb(w_n2090_0[1]),.din(n2090));
	jspl jspl_w_n2091_0(.douta(w_n2091_0[0]),.doutb(w_n2091_0[1]),.din(n2091));
	jspl3 jspl3_w_n2092_0(.douta(w_n2092_0[0]),.doutb(w_n2092_0[1]),.doutc(w_n2092_0[2]),.din(n2092));
	jspl jspl_w_n2093_0(.douta(w_n2093_0[0]),.doutb(w_n2093_0[1]),.din(n2093));
	jspl jspl_w_n2099_0(.douta(w_n2099_0[0]),.doutb(w_n2099_0[1]),.din(n2099));
	jspl jspl_w_n2100_0(.douta(w_n2100_0[0]),.doutb(w_n2100_0[1]),.din(n2100));
	jspl jspl_w_n2102_0(.douta(w_n2102_0[0]),.doutb(w_n2102_0[1]),.din(n2102));
	jspl jspl_w_n2104_0(.douta(w_n2104_0[0]),.doutb(w_n2104_0[1]),.din(n2104));
	jspl jspl_w_n2106_0(.douta(w_n2106_0[0]),.doutb(w_n2106_0[1]),.din(n2106));
	jspl jspl_w_n2112_0(.douta(w_n2112_0[0]),.doutb(w_n2112_0[1]),.din(n2112));
	jspl jspl_w_n2114_0(.douta(w_n2114_0[0]),.doutb(w_n2114_0[1]),.din(n2114));
	jspl3 jspl3_w_n2115_0(.douta(w_n2115_0[0]),.doutb(w_n2115_0[1]),.doutc(w_n2115_0[2]),.din(n2115));
	jspl jspl_w_n2118_0(.douta(w_n2118_0[0]),.doutb(w_n2118_0[1]),.din(n2118));
	jspl jspl_w_n2119_0(.douta(w_n2119_0[0]),.doutb(w_n2119_0[1]),.din(n2119));
	jspl3 jspl3_w_n2120_0(.douta(w_n2120_0[0]),.doutb(w_n2120_0[1]),.doutc(w_n2120_0[2]),.din(n2120));
	jspl jspl_w_n2122_0(.douta(w_n2122_0[0]),.doutb(w_n2122_0[1]),.din(n2122));
	jspl jspl_w_n2126_0(.douta(w_n2126_0[0]),.doutb(w_n2126_0[1]),.din(n2126));
	jspl jspl_w_n2128_0(.douta(w_n2128_0[0]),.doutb(w_n2128_0[1]),.din(n2128));
	jspl jspl_w_n2129_0(.douta(w_n2129_0[0]),.doutb(w_n2129_0[1]),.din(n2129));
	jspl3 jspl3_w_n2130_0(.douta(w_n2130_0[0]),.doutb(w_n2130_0[1]),.doutc(w_n2130_0[2]),.din(n2130));
	jspl jspl_w_n2131_0(.douta(w_n2131_0[0]),.doutb(w_n2131_0[1]),.din(n2131));
	jspl jspl_w_n2134_0(.douta(w_n2134_0[0]),.doutb(w_n2134_0[1]),.din(n2134));
	jspl jspl_w_n2140_0(.douta(w_n2140_0[0]),.doutb(w_n2140_0[1]),.din(n2140));
	jspl jspl_w_n2141_0(.douta(w_n2141_0[0]),.doutb(w_n2141_0[1]),.din(n2141));
	jspl jspl_w_n2143_0(.douta(w_n2143_0[0]),.doutb(w_n2143_0[1]),.din(n2143));
	jspl jspl_w_n2145_0(.douta(w_n2145_0[0]),.doutb(w_n2145_0[1]),.din(n2145));
	jspl jspl_w_n2147_0(.douta(w_n2147_0[0]),.doutb(w_n2147_0[1]),.din(n2147));
	jspl jspl_w_n2153_0(.douta(w_n2153_0[0]),.doutb(w_n2153_0[1]),.din(n2153));
	jspl jspl_w_n2155_0(.douta(w_n2155_0[0]),.doutb(w_n2155_0[1]),.din(n2155));
	jspl3 jspl3_w_n2156_0(.douta(w_n2156_0[0]),.doutb(w_n2156_0[1]),.doutc(w_n2156_0[2]),.din(n2156));
	jspl jspl_w_n2159_0(.douta(w_n2159_0[0]),.doutb(w_n2159_0[1]),.din(n2159));
	jspl jspl_w_n2160_0(.douta(w_n2160_0[0]),.doutb(w_n2160_0[1]),.din(n2160));
	jspl3 jspl3_w_n2161_0(.douta(w_n2161_0[0]),.doutb(w_n2161_0[1]),.doutc(w_n2161_0[2]),.din(n2161));
	jspl jspl_w_n2163_0(.douta(w_n2163_0[0]),.doutb(w_n2163_0[1]),.din(n2163));
	jspl jspl_w_n2167_0(.douta(w_n2167_0[0]),.doutb(w_n2167_0[1]),.din(n2167));
	jspl jspl_w_n2169_0(.douta(w_n2169_0[0]),.doutb(w_n2169_0[1]),.din(n2169));
	jspl jspl_w_n2170_0(.douta(w_n2170_0[0]),.doutb(w_n2170_0[1]),.din(n2170));
	jspl3 jspl3_w_n2171_0(.douta(w_n2171_0[0]),.doutb(w_n2171_0[1]),.doutc(w_n2171_0[2]),.din(n2171));
	jspl jspl_w_n2175_0(.douta(w_n2175_0[0]),.doutb(w_n2175_0[1]),.din(n2175));
	jspl jspl_w_n2181_0(.douta(w_n2181_0[0]),.doutb(w_n2181_0[1]),.din(n2181));
	jspl3 jspl3_w_n2183_0(.douta(w_n2183_0[0]),.doutb(w_n2183_0[1]),.doutc(w_n2183_0[2]),.din(n2183));
	jspl jspl_w_n2185_0(.douta(w_n2185_0[0]),.doutb(w_n2185_0[1]),.din(n2185));
	jspl3 jspl3_w_n2190_0(.douta(w_n2190_0[0]),.doutb(w_n2190_0[1]),.doutc(w_n2190_0[2]),.din(n2190));
	jspl jspl_w_n2191_0(.douta(w_n2191_0[0]),.doutb(w_n2191_0[1]),.din(n2191));
	jspl jspl_w_n2192_0(.douta(w_n2192_0[0]),.doutb(w_n2192_0[1]),.din(n2192));
	jspl jspl_w_n2197_0(.douta(w_n2197_0[0]),.doutb(w_n2197_0[1]),.din(n2197));
	jspl3 jspl3_w_n2198_0(.douta(w_n2198_0[0]),.doutb(w_n2198_0[1]),.doutc(w_n2198_0[2]),.din(n2198));
	jspl jspl_w_n2203_0(.douta(w_n2203_0[0]),.doutb(w_n2203_0[1]),.din(n2203));
	jspl3 jspl3_w_n2209_0(.douta(w_n2209_0[0]),.doutb(w_n2209_0[1]),.doutc(w_n2209_0[2]),.din(n2209));
	jspl jspl_w_n2209_1(.douta(w_n2209_1[0]),.doutb(w_n2209_1[1]),.din(w_n2209_0[0]));
	jspl jspl_w_n2210_0(.douta(w_n2210_0[0]),.doutb(w_n2210_0[1]),.din(n2210));
	jspl3 jspl3_w_n2213_0(.douta(w_n2213_0[0]),.doutb(w_n2213_0[1]),.doutc(w_n2213_0[2]),.din(n2213));
	jspl jspl_w_n2214_0(.douta(w_n2214_0[0]),.doutb(w_n2214_0[1]),.din(n2214));
	jspl jspl_w_n2215_0(.douta(w_n2215_0[0]),.doutb(w_n2215_0[1]),.din(n2215));
	jspl jspl_w_n2216_0(.douta(w_n2216_0[0]),.doutb(w_n2216_0[1]),.din(n2216));
	jspl jspl_w_n2218_0(.douta(w_n2218_0[0]),.doutb(w_n2218_0[1]),.din(n2218));
	jspl jspl_w_n2220_0(.douta(w_n2220_0[0]),.doutb(w_n2220_0[1]),.din(n2220));
	jspl jspl_w_n2222_0(.douta(w_n2222_0[0]),.doutb(w_n2222_0[1]),.din(n2222));
	jspl jspl_w_n2231_0(.douta(w_n2231_0[0]),.doutb(w_n2231_0[1]),.din(n2231));
	jspl3 jspl3_w_n2233_0(.douta(w_n2233_0[0]),.doutb(w_n2233_0[1]),.doutc(w_n2233_0[2]),.din(n2233));
	jspl jspl_w_n2234_0(.douta(w_n2234_0[0]),.doutb(w_n2234_0[1]),.din(n2234));
	jspl jspl_w_n2238_0(.douta(w_n2238_0[0]),.doutb(w_n2238_0[1]),.din(n2238));
	jspl jspl_w_n2240_0(.douta(w_n2240_0[0]),.doutb(w_n2240_0[1]),.din(n2240));
	jspl jspl_w_n2242_0(.douta(w_n2242_0[0]),.doutb(w_n2242_0[1]),.din(n2242));
	jspl jspl_w_n2247_0(.douta(w_n2247_0[0]),.doutb(w_n2247_0[1]),.din(n2247));
	jspl jspl_w_n2249_0(.douta(w_n2249_0[0]),.doutb(w_n2249_0[1]),.din(n2249));
	jspl jspl_w_n2250_0(.douta(w_n2250_0[0]),.doutb(w_n2250_0[1]),.din(n2250));
	jspl3 jspl3_w_n2251_0(.douta(w_n2251_0[0]),.doutb(w_n2251_0[1]),.doutc(w_n2251_0[2]),.din(n2251));
	jspl jspl_w_n2252_0(.douta(w_n2252_0[0]),.doutb(w_n2252_0[1]),.din(n2252));
	jspl jspl_w_n2257_0(.douta(w_n2257_0[0]),.doutb(w_n2257_0[1]),.din(n2257));
	jspl jspl_w_n2258_0(.douta(w_n2258_0[0]),.doutb(w_n2258_0[1]),.din(n2258));
	jspl jspl_w_n2260_0(.douta(w_n2260_0[0]),.doutb(w_n2260_0[1]),.din(n2260));
	jspl jspl_w_n2262_0(.douta(w_n2262_0[0]),.doutb(w_n2262_0[1]),.din(n2262));
	jspl jspl_w_n2265_0(.douta(w_n2265_0[0]),.doutb(w_n2265_0[1]),.din(n2265));
	jspl jspl_w_n2271_0(.douta(w_n2271_0[0]),.doutb(w_n2271_0[1]),.din(n2271));
	jspl3 jspl3_w_n2273_0(.douta(w_n2273_0[0]),.doutb(w_n2273_0[1]),.doutc(w_n2273_0[2]),.din(n2273));
	jspl jspl_w_n2274_0(.douta(w_n2274_0[0]),.doutb(w_n2274_0[1]),.din(n2274));
	jspl jspl_w_n2278_0(.douta(w_n2278_0[0]),.doutb(w_n2278_0[1]),.din(n2278));
	jspl jspl_w_n2279_0(.douta(w_n2279_0[0]),.doutb(w_n2279_0[1]),.din(n2279));
	jspl jspl_w_n2281_0(.douta(w_n2281_0[0]),.doutb(w_n2281_0[1]),.din(n2281));
	jspl jspl_w_n2286_0(.douta(w_n2286_0[0]),.doutb(w_n2286_0[1]),.din(n2286));
	jspl jspl_w_n2288_0(.douta(w_n2288_0[0]),.doutb(w_n2288_0[1]),.din(n2288));
	jspl jspl_w_n2289_0(.douta(w_n2289_0[0]),.doutb(w_n2289_0[1]),.din(n2289));
	jspl3 jspl3_w_n2290_0(.douta(w_n2290_0[0]),.doutb(w_n2290_0[1]),.doutc(w_n2290_0[2]),.din(n2290));
	jspl jspl_w_n2291_0(.douta(w_n2291_0[0]),.doutb(w_n2291_0[1]),.din(n2291));
	jspl jspl_w_n2295_0(.douta(w_n2295_0[0]),.doutb(w_n2295_0[1]),.din(n2295));
	jspl jspl_w_n2296_0(.douta(w_n2296_0[0]),.doutb(w_n2296_0[1]),.din(n2296));
	jspl jspl_w_n2298_0(.douta(w_n2298_0[0]),.doutb(w_n2298_0[1]),.din(n2298));
	jspl jspl_w_n2300_0(.douta(w_n2300_0[0]),.doutb(w_n2300_0[1]),.din(n2300));
	jspl jspl_w_n2303_0(.douta(w_n2303_0[0]),.doutb(w_n2303_0[1]),.din(n2303));
	jspl jspl_w_n2309_0(.douta(w_n2309_0[0]),.doutb(w_n2309_0[1]),.din(n2309));
	jspl jspl_w_n2311_0(.douta(w_n2311_0[0]),.doutb(w_n2311_0[1]),.din(n2311));
	jspl3 jspl3_w_n2312_0(.douta(w_n2312_0[0]),.doutb(w_n2312_0[1]),.doutc(w_n2312_0[2]),.din(n2312));
	jspl jspl_w_n2316_0(.douta(w_n2316_0[0]),.doutb(w_n2316_0[1]),.din(n2316));
	jspl jspl_w_n2317_0(.douta(w_n2317_0[0]),.doutb(w_n2317_0[1]),.din(n2317));
	jspl3 jspl3_w_n2318_0(.douta(w_n2318_0[0]),.doutb(w_n2318_0[1]),.doutc(w_n2318_0[2]),.din(n2318));
	jspl jspl_w_n2320_0(.douta(w_n2320_0[0]),.doutb(w_n2320_0[1]),.din(n2320));
	jspl jspl_w_n2325_0(.douta(w_n2325_0[0]),.doutb(w_n2325_0[1]),.din(n2325));
	jspl jspl_w_n2327_0(.douta(w_n2327_0[0]),.doutb(w_n2327_0[1]),.din(n2327));
	jspl jspl_w_n2328_0(.douta(w_n2328_0[0]),.doutb(w_n2328_0[1]),.din(n2328));
	jspl3 jspl3_w_n2329_0(.douta(w_n2329_0[0]),.doutb(w_n2329_0[1]),.doutc(w_n2329_0[2]),.din(n2329));
	jspl jspl_w_n2330_0(.douta(w_n2330_0[0]),.doutb(w_n2330_0[1]),.din(n2330));
	jspl jspl_w_n2334_0(.douta(w_n2334_0[0]),.doutb(w_n2334_0[1]),.din(n2334));
	jspl jspl_w_n2340_0(.douta(w_n2340_0[0]),.doutb(w_n2340_0[1]),.din(n2340));
	jspl jspl_w_n2341_0(.douta(w_n2341_0[0]),.doutb(w_n2341_0[1]),.din(n2341));
	jspl jspl_w_n2343_0(.douta(w_n2343_0[0]),.doutb(w_n2343_0[1]),.din(n2343));
	jspl jspl_w_n2345_0(.douta(w_n2345_0[0]),.doutb(w_n2345_0[1]),.din(n2345));
	jspl jspl_w_n2348_0(.douta(w_n2348_0[0]),.doutb(w_n2348_0[1]),.din(n2348));
	jspl jspl_w_n2354_0(.douta(w_n2354_0[0]),.doutb(w_n2354_0[1]),.din(n2354));
	jspl jspl_w_n2356_0(.douta(w_n2356_0[0]),.doutb(w_n2356_0[1]),.din(n2356));
	jspl3 jspl3_w_n2357_0(.douta(w_n2357_0[0]),.doutb(w_n2357_0[1]),.doutc(w_n2357_0[2]),.din(n2357));
	jspl jspl_w_n2361_0(.douta(w_n2361_0[0]),.doutb(w_n2361_0[1]),.din(n2361));
	jspl jspl_w_n2362_0(.douta(w_n2362_0[0]),.doutb(w_n2362_0[1]),.din(n2362));
	jspl3 jspl3_w_n2363_0(.douta(w_n2363_0[0]),.doutb(w_n2363_0[1]),.doutc(w_n2363_0[2]),.din(n2363));
	jspl jspl_w_n2365_0(.douta(w_n2365_0[0]),.doutb(w_n2365_0[1]),.din(n2365));
	jspl jspl_w_n2370_0(.douta(w_n2370_0[0]),.doutb(w_n2370_0[1]),.din(n2370));
	jspl jspl_w_n2372_0(.douta(w_n2372_0[0]),.doutb(w_n2372_0[1]),.din(n2372));
	jspl jspl_w_n2373_0(.douta(w_n2373_0[0]),.doutb(w_n2373_0[1]),.din(n2373));
	jspl3 jspl3_w_n2374_0(.douta(w_n2374_0[0]),.doutb(w_n2374_0[1]),.doutc(w_n2374_0[2]),.din(n2374));
	jspl jspl_w_n2375_0(.douta(w_n2375_0[0]),.doutb(w_n2375_0[1]),.din(n2375));
	jspl jspl_w_n2379_0(.douta(w_n2379_0[0]),.doutb(w_n2379_0[1]),.din(n2379));
	jspl jspl_w_n2385_0(.douta(w_n2385_0[0]),.doutb(w_n2385_0[1]),.din(n2385));
	jspl jspl_w_n2386_0(.douta(w_n2386_0[0]),.doutb(w_n2386_0[1]),.din(n2386));
	jspl jspl_w_n2388_0(.douta(w_n2388_0[0]),.doutb(w_n2388_0[1]),.din(n2388));
	jspl jspl_w_n2390_0(.douta(w_n2390_0[0]),.doutb(w_n2390_0[1]),.din(n2390));
	jspl jspl_w_n2393_0(.douta(w_n2393_0[0]),.doutb(w_n2393_0[1]),.din(n2393));
	jspl jspl_w_n2399_0(.douta(w_n2399_0[0]),.doutb(w_n2399_0[1]),.din(n2399));
	jspl3 jspl3_w_n2401_0(.douta(w_n2401_0[0]),.doutb(w_n2401_0[1]),.doutc(w_n2401_0[2]),.din(n2401));
	jspl3 jspl3_w_n2401_1(.douta(w_n2401_1[0]),.doutb(w_n2401_1[1]),.doutc(w_n2401_1[2]),.din(w_n2401_0[0]));
	jspl jspl_w_n2404_0(.douta(w_n2404_0[0]),.doutb(w_n2404_0[1]),.din(n2404));
	jspl3 jspl3_w_n2405_0(.douta(w_n2405_0[0]),.doutb(w_n2405_0[1]),.doutc(w_n2405_0[2]),.din(n2405));
	jspl jspl_w_n2406_0(.douta(w_n2406_0[0]),.doutb(w_n2406_0[1]),.din(n2406));
	jspl jspl_w_n2412_0(.douta(w_n2412_0[0]),.doutb(w_n2412_0[1]),.din(n2412));
	jspl3 jspl3_w_n2413_0(.douta(w_n2413_0[0]),.doutb(w_n2413_0[1]),.doutc(w_n2413_0[2]),.din(n2413));
	jspl jspl_w_n2414_0(.douta(w_n2414_0[0]),.doutb(w_n2414_0[1]),.din(n2414));
	jspl jspl_w_n2419_0(.douta(w_n2419_0[0]),.doutb(w_n2419_0[1]),.din(n2419));
	jspl3 jspl3_w_n2420_0(.douta(w_n2420_0[0]),.doutb(w_n2420_0[1]),.doutc(w_n2420_0[2]),.din(n2420));
	jspl3 jspl3_w_n2420_1(.douta(w_n2420_1[0]),.doutb(w_n2420_1[1]),.doutc(w_n2420_1[2]),.din(w_n2420_0[0]));
	jspl3 jspl3_w_n2420_2(.douta(w_n2420_2[0]),.doutb(w_n2420_2[1]),.doutc(w_n2420_2[2]),.din(w_n2420_0[1]));
	jspl3 jspl3_w_n2420_3(.douta(w_n2420_3[0]),.doutb(w_n2420_3[1]),.doutc(w_n2420_3[2]),.din(w_n2420_0[2]));
	jspl3 jspl3_w_n2420_4(.douta(w_n2420_4[0]),.doutb(w_n2420_4[1]),.doutc(w_n2420_4[2]),.din(w_n2420_1[0]));
	jspl3 jspl3_w_n2420_5(.douta(w_n2420_5[0]),.doutb(w_n2420_5[1]),.doutc(w_n2420_5[2]),.din(w_n2420_1[1]));
	jspl3 jspl3_w_n2420_6(.douta(w_n2420_6[0]),.doutb(w_n2420_6[1]),.doutc(w_n2420_6[2]),.din(w_n2420_1[2]));
	jspl3 jspl3_w_n2420_7(.douta(w_n2420_7[0]),.doutb(w_n2420_7[1]),.doutc(w_n2420_7[2]),.din(w_n2420_2[0]));
	jspl3 jspl3_w_n2420_8(.douta(w_n2420_8[0]),.doutb(w_n2420_8[1]),.doutc(w_n2420_8[2]),.din(w_n2420_2[1]));
	jspl3 jspl3_w_n2420_9(.douta(w_n2420_9[0]),.doutb(w_n2420_9[1]),.doutc(w_n2420_9[2]),.din(w_n2420_2[2]));
	jspl3 jspl3_w_n2420_10(.douta(w_n2420_10[0]),.doutb(w_n2420_10[1]),.doutc(w_n2420_10[2]),.din(w_n2420_3[0]));
	jspl3 jspl3_w_n2420_11(.douta(w_n2420_11[0]),.doutb(w_n2420_11[1]),.doutc(w_n2420_11[2]),.din(w_n2420_3[1]));
	jspl3 jspl3_w_n2420_12(.douta(w_n2420_12[0]),.doutb(w_n2420_12[1]),.doutc(w_n2420_12[2]),.din(w_n2420_3[2]));
	jspl3 jspl3_w_n2420_13(.douta(w_n2420_13[0]),.doutb(w_n2420_13[1]),.doutc(w_n2420_13[2]),.din(w_n2420_4[0]));
	jspl3 jspl3_w_n2420_14(.douta(w_n2420_14[0]),.doutb(w_n2420_14[1]),.doutc(w_n2420_14[2]),.din(w_n2420_4[1]));
	jspl3 jspl3_w_n2420_15(.douta(w_n2420_15[0]),.doutb(w_n2420_15[1]),.doutc(w_n2420_15[2]),.din(w_n2420_4[2]));
	jspl3 jspl3_w_n2420_16(.douta(w_n2420_16[0]),.doutb(w_n2420_16[1]),.doutc(w_n2420_16[2]),.din(w_n2420_5[0]));
	jspl3 jspl3_w_n2420_17(.douta(w_n2420_17[0]),.doutb(w_n2420_17[1]),.doutc(w_n2420_17[2]),.din(w_n2420_5[1]));
	jspl3 jspl3_w_n2420_18(.douta(w_n2420_18[0]),.doutb(w_n2420_18[1]),.doutc(w_n2420_18[2]),.din(w_n2420_5[2]));
	jspl3 jspl3_w_n2420_19(.douta(w_n2420_19[0]),.doutb(w_n2420_19[1]),.doutc(w_n2420_19[2]),.din(w_n2420_6[0]));
	jspl3 jspl3_w_n2420_20(.douta(w_n2420_20[0]),.doutb(w_n2420_20[1]),.doutc(w_n2420_20[2]),.din(w_n2420_6[1]));
	jspl3 jspl3_w_n2420_21(.douta(w_n2420_21[0]),.doutb(w_n2420_21[1]),.doutc(w_n2420_21[2]),.din(w_n2420_6[2]));
	jspl3 jspl3_w_n2420_22(.douta(w_n2420_22[0]),.doutb(w_n2420_22[1]),.doutc(w_n2420_22[2]),.din(w_n2420_7[0]));
	jspl3 jspl3_w_n2420_23(.douta(w_n2420_23[0]),.doutb(w_n2420_23[1]),.doutc(w_n2420_23[2]),.din(w_n2420_7[1]));
	jspl3 jspl3_w_n2420_24(.douta(w_n2420_24[0]),.doutb(w_n2420_24[1]),.doutc(w_n2420_24[2]),.din(w_n2420_7[2]));
	jspl3 jspl3_w_n2420_25(.douta(w_n2420_25[0]),.doutb(w_n2420_25[1]),.doutc(w_n2420_25[2]),.din(w_n2420_8[0]));
	jspl3 jspl3_w_n2420_26(.douta(w_n2420_26[0]),.doutb(w_n2420_26[1]),.doutc(w_n2420_26[2]),.din(w_n2420_8[1]));
	jspl3 jspl3_w_n2420_27(.douta(w_n2420_27[0]),.doutb(w_n2420_27[1]),.doutc(w_n2420_27[2]),.din(w_n2420_8[2]));
	jspl jspl_w_n2420_28(.douta(w_n2420_28[0]),.doutb(w_n2420_28[1]),.din(w_n2420_9[0]));
	jspl3 jspl3_w_n2425_0(.douta(w_n2425_0[0]),.doutb(w_n2425_0[1]),.doutc(w_n2425_0[2]),.din(n2425));
	jspl3 jspl3_w_n2425_1(.douta(w_n2425_1[0]),.doutb(w_n2425_1[1]),.doutc(w_n2425_1[2]),.din(w_n2425_0[0]));
	jspl3 jspl3_w_n2425_2(.douta(w_n2425_2[0]),.doutb(w_n2425_2[1]),.doutc(w_n2425_2[2]),.din(w_n2425_0[1]));
	jspl3 jspl3_w_n2425_3(.douta(w_n2425_3[0]),.doutb(w_n2425_3[1]),.doutc(w_n2425_3[2]),.din(w_n2425_0[2]));
	jspl3 jspl3_w_n2425_4(.douta(w_n2425_4[0]),.doutb(w_n2425_4[1]),.doutc(w_n2425_4[2]),.din(w_n2425_1[0]));
	jspl3 jspl3_w_n2425_5(.douta(w_n2425_5[0]),.doutb(w_n2425_5[1]),.doutc(w_n2425_5[2]),.din(w_n2425_1[1]));
	jspl3 jspl3_w_n2425_6(.douta(w_n2425_6[0]),.doutb(w_n2425_6[1]),.doutc(w_n2425_6[2]),.din(w_n2425_1[2]));
	jspl3 jspl3_w_n2425_7(.douta(w_n2425_7[0]),.doutb(w_n2425_7[1]),.doutc(w_n2425_7[2]),.din(w_n2425_2[0]));
	jspl3 jspl3_w_n2425_8(.douta(w_n2425_8[0]),.doutb(w_n2425_8[1]),.doutc(w_n2425_8[2]),.din(w_n2425_2[1]));
	jspl3 jspl3_w_n2425_9(.douta(w_n2425_9[0]),.doutb(w_n2425_9[1]),.doutc(w_n2425_9[2]),.din(w_n2425_2[2]));
	jspl3 jspl3_w_n2425_10(.douta(w_n2425_10[0]),.doutb(w_n2425_10[1]),.doutc(w_n2425_10[2]),.din(w_n2425_3[0]));
	jspl3 jspl3_w_n2425_11(.douta(w_n2425_11[0]),.doutb(w_n2425_11[1]),.doutc(w_n2425_11[2]),.din(w_n2425_3[1]));
	jspl3 jspl3_w_n2425_12(.douta(w_n2425_12[0]),.doutb(w_n2425_12[1]),.doutc(w_n2425_12[2]),.din(w_n2425_3[2]));
	jspl3 jspl3_w_n2425_13(.douta(w_n2425_13[0]),.doutb(w_n2425_13[1]),.doutc(w_n2425_13[2]),.din(w_n2425_4[0]));
	jspl3 jspl3_w_n2425_14(.douta(w_n2425_14[0]),.doutb(w_n2425_14[1]),.doutc(w_n2425_14[2]),.din(w_n2425_4[1]));
	jspl3 jspl3_w_n2425_15(.douta(w_n2425_15[0]),.doutb(w_n2425_15[1]),.doutc(w_n2425_15[2]),.din(w_n2425_4[2]));
	jspl3 jspl3_w_n2425_16(.douta(w_n2425_16[0]),.doutb(w_n2425_16[1]),.doutc(w_n2425_16[2]),.din(w_n2425_5[0]));
	jspl3 jspl3_w_n2425_17(.douta(w_n2425_17[0]),.doutb(w_n2425_17[1]),.doutc(w_n2425_17[2]),.din(w_n2425_5[1]));
	jspl3 jspl3_w_n2425_18(.douta(w_n2425_18[0]),.doutb(w_n2425_18[1]),.doutc(w_n2425_18[2]),.din(w_n2425_5[2]));
	jspl3 jspl3_w_n2425_19(.douta(w_n2425_19[0]),.doutb(w_n2425_19[1]),.doutc(w_n2425_19[2]),.din(w_n2425_6[0]));
	jspl3 jspl3_w_n2425_20(.douta(w_n2425_20[0]),.doutb(w_n2425_20[1]),.doutc(w_n2425_20[2]),.din(w_n2425_6[1]));
	jspl3 jspl3_w_n2425_21(.douta(w_n2425_21[0]),.doutb(w_n2425_21[1]),.doutc(w_n2425_21[2]),.din(w_n2425_6[2]));
	jspl3 jspl3_w_n2425_22(.douta(w_n2425_22[0]),.doutb(w_n2425_22[1]),.doutc(w_n2425_22[2]),.din(w_n2425_7[0]));
	jspl3 jspl3_w_n2425_23(.douta(w_n2425_23[0]),.doutb(w_n2425_23[1]),.doutc(w_n2425_23[2]),.din(w_n2425_7[1]));
	jspl3 jspl3_w_n2425_24(.douta(w_n2425_24[0]),.doutb(w_n2425_24[1]),.doutc(w_n2425_24[2]),.din(w_n2425_7[2]));
	jspl3 jspl3_w_n2425_25(.douta(w_n2425_25[0]),.doutb(w_n2425_25[1]),.doutc(w_n2425_25[2]),.din(w_n2425_8[0]));
	jspl3 jspl3_w_n2425_26(.douta(w_n2425_26[0]),.doutb(w_n2425_26[1]),.doutc(w_n2425_26[2]),.din(w_n2425_8[1]));
	jspl3 jspl3_w_n2425_27(.douta(w_n2425_27[0]),.doutb(w_n2425_27[1]),.doutc(w_n2425_27[2]),.din(w_n2425_8[2]));
	jspl3 jspl3_w_n2425_28(.douta(w_n2425_28[0]),.doutb(w_n2425_28[1]),.doutc(w_n2425_28[2]),.din(w_n2425_9[0]));
	jspl3 jspl3_w_n2425_29(.douta(w_n2425_29[0]),.doutb(w_n2425_29[1]),.doutc(w_n2425_29[2]),.din(w_n2425_9[1]));
	jspl3 jspl3_w_n2425_30(.douta(w_n2425_30[0]),.doutb(w_n2425_30[1]),.doutc(w_n2425_30[2]),.din(w_n2425_9[2]));
	jspl3 jspl3_w_n2425_31(.douta(w_n2425_31[0]),.doutb(w_n2425_31[1]),.doutc(w_n2425_31[2]),.din(w_n2425_10[0]));
	jspl3 jspl3_w_n2425_32(.douta(w_n2425_32[0]),.doutb(w_n2425_32[1]),.doutc(w_n2425_32[2]),.din(w_n2425_10[1]));
	jspl3 jspl3_w_n2425_33(.douta(w_n2425_33[0]),.doutb(w_n2425_33[1]),.doutc(w_n2425_33[2]),.din(w_n2425_10[2]));
	jspl3 jspl3_w_n2425_34(.douta(w_n2425_34[0]),.doutb(w_n2425_34[1]),.doutc(w_n2425_34[2]),.din(w_n2425_11[0]));
	jspl3 jspl3_w_n2428_0(.douta(w_n2428_0[0]),.doutb(w_n2428_0[1]),.doutc(w_n2428_0[2]),.din(n2428));
	jspl jspl_w_n2428_1(.douta(w_n2428_1[0]),.doutb(w_n2428_1[1]),.din(w_n2428_0[0]));
	jspl3 jspl3_w_n2429_0(.douta(w_n2429_0[0]),.doutb(w_n2429_0[1]),.doutc(w_n2429_0[2]),.din(n2429));
	jspl3 jspl3_w_n2433_0(.douta(w_n2433_0[0]),.doutb(w_n2433_0[1]),.doutc(w_n2433_0[2]),.din(n2433));
	jspl jspl_w_n2434_0(.douta(w_n2434_0[0]),.doutb(w_n2434_0[1]),.din(n2434));
	jspl jspl_w_n2435_0(.douta(w_n2435_0[0]),.doutb(w_n2435_0[1]),.din(n2435));
	jspl jspl_w_n2436_0(.douta(w_n2436_0[0]),.doutb(w_n2436_0[1]),.din(n2436));
	jspl jspl_w_n2438_0(.douta(w_n2438_0[0]),.doutb(w_n2438_0[1]),.din(n2438));
	jspl jspl_w_n2440_0(.douta(w_n2440_0[0]),.doutb(w_n2440_0[1]),.din(n2440));
	jspl jspl_w_n2442_0(.douta(w_n2442_0[0]),.doutb(w_n2442_0[1]),.din(n2442));
	jspl jspl_w_n2445_0(.douta(w_n2445_0[0]),.doutb(w_n2445_0[1]),.din(n2445));
	jspl jspl_w_n2450_0(.douta(w_n2450_0[0]),.doutb(w_n2450_0[1]),.din(n2450));
	jspl3 jspl3_w_n2452_0(.douta(w_n2452_0[0]),.doutb(w_n2452_0[1]),.doutc(w_n2452_0[2]),.din(n2452));
	jspl jspl_w_n2453_0(.douta(w_n2453_0[0]),.doutb(w_n2453_0[1]),.din(n2453));
	jspl jspl_w_n2457_0(.douta(w_n2457_0[0]),.doutb(w_n2457_0[1]),.din(n2457));
	jspl jspl_w_n2458_0(.douta(w_n2458_0[0]),.doutb(w_n2458_0[1]),.din(n2458));
	jspl jspl_w_n2460_0(.douta(w_n2460_0[0]),.doutb(w_n2460_0[1]),.din(n2460));
	jspl jspl_w_n2464_0(.douta(w_n2464_0[0]),.doutb(w_n2464_0[1]),.din(n2464));
	jspl jspl_w_n2466_0(.douta(w_n2466_0[0]),.doutb(w_n2466_0[1]),.din(n2466));
	jspl jspl_w_n2467_0(.douta(w_n2467_0[0]),.doutb(w_n2467_0[1]),.din(n2467));
	jspl3 jspl3_w_n2468_0(.douta(w_n2468_0[0]),.doutb(w_n2468_0[1]),.doutc(w_n2468_0[2]),.din(n2468));
	jspl jspl_w_n2469_0(.douta(w_n2469_0[0]),.doutb(w_n2469_0[1]),.din(n2469));
	jspl jspl_w_n2473_0(.douta(w_n2473_0[0]),.doutb(w_n2473_0[1]),.din(n2473));
	jspl jspl_w_n2475_0(.douta(w_n2475_0[0]),.doutb(w_n2475_0[1]),.din(n2475));
	jspl jspl_w_n2477_0(.douta(w_n2477_0[0]),.doutb(w_n2477_0[1]),.din(n2477));
	jspl jspl_w_n2479_0(.douta(w_n2479_0[0]),.doutb(w_n2479_0[1]),.din(n2479));
	jspl jspl_w_n2481_0(.douta(w_n2481_0[0]),.doutb(w_n2481_0[1]),.din(n2481));
	jspl jspl_w_n2487_0(.douta(w_n2487_0[0]),.doutb(w_n2487_0[1]),.din(n2487));
	jspl3 jspl3_w_n2489_0(.douta(w_n2489_0[0]),.doutb(w_n2489_0[1]),.doutc(w_n2489_0[2]),.din(n2489));
	jspl jspl_w_n2490_0(.douta(w_n2490_0[0]),.doutb(w_n2490_0[1]),.din(n2490));
	jspl jspl_w_n2495_0(.douta(w_n2495_0[0]),.doutb(w_n2495_0[1]),.din(n2495));
	jspl jspl_w_n2497_0(.douta(w_n2497_0[0]),.doutb(w_n2497_0[1]),.din(n2497));
	jspl jspl_w_n2499_0(.douta(w_n2499_0[0]),.doutb(w_n2499_0[1]),.din(n2499));
	jspl jspl_w_n2503_0(.douta(w_n2503_0[0]),.doutb(w_n2503_0[1]),.din(n2503));
	jspl jspl_w_n2505_0(.douta(w_n2505_0[0]),.doutb(w_n2505_0[1]),.din(n2505));
	jspl jspl_w_n2506_0(.douta(w_n2506_0[0]),.doutb(w_n2506_0[1]),.din(n2506));
	jspl3 jspl3_w_n2507_0(.douta(w_n2507_0[0]),.doutb(w_n2507_0[1]),.doutc(w_n2507_0[2]),.din(n2507));
	jspl jspl_w_n2508_0(.douta(w_n2508_0[0]),.doutb(w_n2508_0[1]),.din(n2508));
	jspl jspl_w_n2514_0(.douta(w_n2514_0[0]),.doutb(w_n2514_0[1]),.din(n2514));
	jspl jspl_w_n2515_0(.douta(w_n2515_0[0]),.doutb(w_n2515_0[1]),.din(n2515));
	jspl jspl_w_n2517_0(.douta(w_n2517_0[0]),.doutb(w_n2517_0[1]),.din(n2517));
	jspl jspl_w_n2519_0(.douta(w_n2519_0[0]),.doutb(w_n2519_0[1]),.din(n2519));
	jspl jspl_w_n2521_0(.douta(w_n2521_0[0]),.doutb(w_n2521_0[1]),.din(n2521));
	jspl jspl_w_n2527_0(.douta(w_n2527_0[0]),.doutb(w_n2527_0[1]),.din(n2527));
	jspl jspl_w_n2529_0(.douta(w_n2529_0[0]),.doutb(w_n2529_0[1]),.din(n2529));
	jspl3 jspl3_w_n2530_0(.douta(w_n2530_0[0]),.doutb(w_n2530_0[1]),.doutc(w_n2530_0[2]),.din(n2530));
	jspl jspl_w_n2533_0(.douta(w_n2533_0[0]),.doutb(w_n2533_0[1]),.din(n2533));
	jspl jspl_w_n2534_0(.douta(w_n2534_0[0]),.doutb(w_n2534_0[1]),.din(n2534));
	jspl3 jspl3_w_n2535_0(.douta(w_n2535_0[0]),.doutb(w_n2535_0[1]),.doutc(w_n2535_0[2]),.din(n2535));
	jspl jspl_w_n2537_0(.douta(w_n2537_0[0]),.doutb(w_n2537_0[1]),.din(n2537));
	jspl jspl_w_n2541_0(.douta(w_n2541_0[0]),.doutb(w_n2541_0[1]),.din(n2541));
	jspl jspl_w_n2543_0(.douta(w_n2543_0[0]),.doutb(w_n2543_0[1]),.din(n2543));
	jspl jspl_w_n2544_0(.douta(w_n2544_0[0]),.doutb(w_n2544_0[1]),.din(n2544));
	jspl3 jspl3_w_n2545_0(.douta(w_n2545_0[0]),.doutb(w_n2545_0[1]),.doutc(w_n2545_0[2]),.din(n2545));
	jspl jspl_w_n2546_0(.douta(w_n2546_0[0]),.doutb(w_n2546_0[1]),.din(n2546));
	jspl jspl_w_n2549_0(.douta(w_n2549_0[0]),.doutb(w_n2549_0[1]),.din(n2549));
	jspl jspl_w_n2555_0(.douta(w_n2555_0[0]),.doutb(w_n2555_0[1]),.din(n2555));
	jspl jspl_w_n2556_0(.douta(w_n2556_0[0]),.doutb(w_n2556_0[1]),.din(n2556));
	jspl jspl_w_n2558_0(.douta(w_n2558_0[0]),.doutb(w_n2558_0[1]),.din(n2558));
	jspl jspl_w_n2560_0(.douta(w_n2560_0[0]),.doutb(w_n2560_0[1]),.din(n2560));
	jspl jspl_w_n2562_0(.douta(w_n2562_0[0]),.doutb(w_n2562_0[1]),.din(n2562));
	jspl jspl_w_n2568_0(.douta(w_n2568_0[0]),.doutb(w_n2568_0[1]),.din(n2568));
	jspl jspl_w_n2570_0(.douta(w_n2570_0[0]),.doutb(w_n2570_0[1]),.din(n2570));
	jspl3 jspl3_w_n2571_0(.douta(w_n2571_0[0]),.doutb(w_n2571_0[1]),.doutc(w_n2571_0[2]),.din(n2571));
	jspl jspl_w_n2574_0(.douta(w_n2574_0[0]),.doutb(w_n2574_0[1]),.din(n2574));
	jspl jspl_w_n2575_0(.douta(w_n2575_0[0]),.doutb(w_n2575_0[1]),.din(n2575));
	jspl3 jspl3_w_n2576_0(.douta(w_n2576_0[0]),.doutb(w_n2576_0[1]),.doutc(w_n2576_0[2]),.din(n2576));
	jspl jspl_w_n2578_0(.douta(w_n2578_0[0]),.doutb(w_n2578_0[1]),.din(n2578));
	jspl jspl_w_n2582_0(.douta(w_n2582_0[0]),.doutb(w_n2582_0[1]),.din(n2582));
	jspl jspl_w_n2584_0(.douta(w_n2584_0[0]),.doutb(w_n2584_0[1]),.din(n2584));
	jspl jspl_w_n2585_0(.douta(w_n2585_0[0]),.doutb(w_n2585_0[1]),.din(n2585));
	jspl3 jspl3_w_n2586_0(.douta(w_n2586_0[0]),.doutb(w_n2586_0[1]),.doutc(w_n2586_0[2]),.din(n2586));
	jspl jspl_w_n2587_0(.douta(w_n2587_0[0]),.doutb(w_n2587_0[1]),.din(n2587));
	jspl jspl_w_n2590_0(.douta(w_n2590_0[0]),.doutb(w_n2590_0[1]),.din(n2590));
	jspl jspl_w_n2596_0(.douta(w_n2596_0[0]),.doutb(w_n2596_0[1]),.din(n2596));
	jspl jspl_w_n2597_0(.douta(w_n2597_0[0]),.doutb(w_n2597_0[1]),.din(n2597));
	jspl jspl_w_n2599_0(.douta(w_n2599_0[0]),.doutb(w_n2599_0[1]),.din(n2599));
	jspl jspl_w_n2601_0(.douta(w_n2601_0[0]),.doutb(w_n2601_0[1]),.din(n2601));
	jspl jspl_w_n2603_0(.douta(w_n2603_0[0]),.doutb(w_n2603_0[1]),.din(n2603));
	jspl jspl_w_n2609_0(.douta(w_n2609_0[0]),.doutb(w_n2609_0[1]),.din(n2609));
	jspl3 jspl3_w_n2611_0(.douta(w_n2611_0[0]),.doutb(w_n2611_0[1]),.doutc(w_n2611_0[2]),.din(n2611));
	jspl jspl_w_n2616_0(.douta(w_n2616_0[0]),.doutb(w_n2616_0[1]),.din(n2616));
	jspl3 jspl3_w_n2618_0(.douta(w_n2618_0[0]),.doutb(w_n2618_0[1]),.doutc(w_n2618_0[2]),.din(n2618));
	jspl3 jspl3_w_n2622_0(.douta(w_n2622_0[0]),.doutb(w_n2622_0[1]),.doutc(w_n2622_0[2]),.din(n2622));
	jspl jspl_w_n2623_0(.douta(w_n2623_0[0]),.doutb(w_n2623_0[1]),.din(n2623));
	jspl jspl_w_n2628_0(.douta(w_n2628_0[0]),.doutb(w_n2628_0[1]),.din(n2628));
	jspl3 jspl3_w_n2629_0(.douta(w_n2629_0[0]),.doutb(w_n2629_0[1]),.doutc(w_n2629_0[2]),.din(n2629));
	jspl jspl_w_n2634_0(.douta(w_n2634_0[0]),.doutb(w_n2634_0[1]),.din(n2634));
	jspl3 jspl3_w_n2640_0(.douta(w_n2640_0[0]),.doutb(w_n2640_0[1]),.doutc(w_n2640_0[2]),.din(n2640));
	jspl jspl_w_n2640_1(.douta(w_n2640_1[0]),.doutb(w_n2640_1[1]),.din(w_n2640_0[0]));
	jspl jspl_w_n2641_0(.douta(w_n2641_0[0]),.doutb(w_n2641_0[1]),.din(n2641));
	jspl3 jspl3_w_n2644_0(.douta(w_n2644_0[0]),.doutb(w_n2644_0[1]),.doutc(w_n2644_0[2]),.din(n2644));
	jspl jspl_w_n2645_0(.douta(w_n2645_0[0]),.doutb(w_n2645_0[1]),.din(n2645));
	jspl jspl_w_n2646_0(.douta(w_n2646_0[0]),.doutb(w_n2646_0[1]),.din(n2646));
	jspl jspl_w_n2647_0(.douta(w_n2647_0[0]),.doutb(w_n2647_0[1]),.din(n2647));
	jspl jspl_w_n2649_0(.douta(w_n2649_0[0]),.doutb(w_n2649_0[1]),.din(n2649));
	jspl jspl_w_n2651_0(.douta(w_n2651_0[0]),.doutb(w_n2651_0[1]),.din(n2651));
	jspl jspl_w_n2653_0(.douta(w_n2653_0[0]),.doutb(w_n2653_0[1]),.din(n2653));
	jspl jspl_w_n2662_0(.douta(w_n2662_0[0]),.doutb(w_n2662_0[1]),.din(n2662));
	jspl3 jspl3_w_n2664_0(.douta(w_n2664_0[0]),.doutb(w_n2664_0[1]),.doutc(w_n2664_0[2]),.din(n2664));
	jspl jspl_w_n2665_0(.douta(w_n2665_0[0]),.doutb(w_n2665_0[1]),.din(n2665));
	jspl jspl_w_n2669_0(.douta(w_n2669_0[0]),.doutb(w_n2669_0[1]),.din(n2669));
	jspl jspl_w_n2671_0(.douta(w_n2671_0[0]),.doutb(w_n2671_0[1]),.din(n2671));
	jspl jspl_w_n2673_0(.douta(w_n2673_0[0]),.doutb(w_n2673_0[1]),.din(n2673));
	jspl jspl_w_n2678_0(.douta(w_n2678_0[0]),.doutb(w_n2678_0[1]),.din(n2678));
	jspl jspl_w_n2680_0(.douta(w_n2680_0[0]),.doutb(w_n2680_0[1]),.din(n2680));
	jspl jspl_w_n2681_0(.douta(w_n2681_0[0]),.doutb(w_n2681_0[1]),.din(n2681));
	jspl3 jspl3_w_n2682_0(.douta(w_n2682_0[0]),.doutb(w_n2682_0[1]),.doutc(w_n2682_0[2]),.din(n2682));
	jspl jspl_w_n2683_0(.douta(w_n2683_0[0]),.doutb(w_n2683_0[1]),.din(n2683));
	jspl jspl_w_n2688_0(.douta(w_n2688_0[0]),.doutb(w_n2688_0[1]),.din(n2688));
	jspl jspl_w_n2689_0(.douta(w_n2689_0[0]),.doutb(w_n2689_0[1]),.din(n2689));
	jspl jspl_w_n2691_0(.douta(w_n2691_0[0]),.doutb(w_n2691_0[1]),.din(n2691));
	jspl jspl_w_n2693_0(.douta(w_n2693_0[0]),.doutb(w_n2693_0[1]),.din(n2693));
	jspl jspl_w_n2696_0(.douta(w_n2696_0[0]),.doutb(w_n2696_0[1]),.din(n2696));
	jspl jspl_w_n2702_0(.douta(w_n2702_0[0]),.doutb(w_n2702_0[1]),.din(n2702));
	jspl3 jspl3_w_n2704_0(.douta(w_n2704_0[0]),.doutb(w_n2704_0[1]),.doutc(w_n2704_0[2]),.din(n2704));
	jspl jspl_w_n2705_0(.douta(w_n2705_0[0]),.doutb(w_n2705_0[1]),.din(n2705));
	jspl jspl_w_n2709_0(.douta(w_n2709_0[0]),.doutb(w_n2709_0[1]),.din(n2709));
	jspl jspl_w_n2710_0(.douta(w_n2710_0[0]),.doutb(w_n2710_0[1]),.din(n2710));
	jspl jspl_w_n2712_0(.douta(w_n2712_0[0]),.doutb(w_n2712_0[1]),.din(n2712));
	jspl jspl_w_n2717_0(.douta(w_n2717_0[0]),.doutb(w_n2717_0[1]),.din(n2717));
	jspl jspl_w_n2719_0(.douta(w_n2719_0[0]),.doutb(w_n2719_0[1]),.din(n2719));
	jspl jspl_w_n2720_0(.douta(w_n2720_0[0]),.doutb(w_n2720_0[1]),.din(n2720));
	jspl3 jspl3_w_n2721_0(.douta(w_n2721_0[0]),.doutb(w_n2721_0[1]),.doutc(w_n2721_0[2]),.din(n2721));
	jspl jspl_w_n2722_0(.douta(w_n2722_0[0]),.doutb(w_n2722_0[1]),.din(n2722));
	jspl jspl_w_n2726_0(.douta(w_n2726_0[0]),.doutb(w_n2726_0[1]),.din(n2726));
	jspl jspl_w_n2727_0(.douta(w_n2727_0[0]),.doutb(w_n2727_0[1]),.din(n2727));
	jspl jspl_w_n2729_0(.douta(w_n2729_0[0]),.doutb(w_n2729_0[1]),.din(n2729));
	jspl jspl_w_n2731_0(.douta(w_n2731_0[0]),.doutb(w_n2731_0[1]),.din(n2731));
	jspl jspl_w_n2734_0(.douta(w_n2734_0[0]),.doutb(w_n2734_0[1]),.din(n2734));
	jspl jspl_w_n2740_0(.douta(w_n2740_0[0]),.doutb(w_n2740_0[1]),.din(n2740));
	jspl jspl_w_n2742_0(.douta(w_n2742_0[0]),.doutb(w_n2742_0[1]),.din(n2742));
	jspl3 jspl3_w_n2743_0(.douta(w_n2743_0[0]),.doutb(w_n2743_0[1]),.doutc(w_n2743_0[2]),.din(n2743));
	jspl jspl_w_n2747_0(.douta(w_n2747_0[0]),.doutb(w_n2747_0[1]),.din(n2747));
	jspl jspl_w_n2748_0(.douta(w_n2748_0[0]),.doutb(w_n2748_0[1]),.din(n2748));
	jspl3 jspl3_w_n2749_0(.douta(w_n2749_0[0]),.doutb(w_n2749_0[1]),.doutc(w_n2749_0[2]),.din(n2749));
	jspl jspl_w_n2751_0(.douta(w_n2751_0[0]),.doutb(w_n2751_0[1]),.din(n2751));
	jspl jspl_w_n2756_0(.douta(w_n2756_0[0]),.doutb(w_n2756_0[1]),.din(n2756));
	jspl jspl_w_n2758_0(.douta(w_n2758_0[0]),.doutb(w_n2758_0[1]),.din(n2758));
	jspl jspl_w_n2759_0(.douta(w_n2759_0[0]),.doutb(w_n2759_0[1]),.din(n2759));
	jspl3 jspl3_w_n2760_0(.douta(w_n2760_0[0]),.doutb(w_n2760_0[1]),.doutc(w_n2760_0[2]),.din(n2760));
	jspl jspl_w_n2761_0(.douta(w_n2761_0[0]),.doutb(w_n2761_0[1]),.din(n2761));
	jspl jspl_w_n2765_0(.douta(w_n2765_0[0]),.doutb(w_n2765_0[1]),.din(n2765));
	jspl jspl_w_n2771_0(.douta(w_n2771_0[0]),.doutb(w_n2771_0[1]),.din(n2771));
	jspl jspl_w_n2772_0(.douta(w_n2772_0[0]),.doutb(w_n2772_0[1]),.din(n2772));
	jspl jspl_w_n2774_0(.douta(w_n2774_0[0]),.doutb(w_n2774_0[1]),.din(n2774));
	jspl jspl_w_n2776_0(.douta(w_n2776_0[0]),.doutb(w_n2776_0[1]),.din(n2776));
	jspl jspl_w_n2779_0(.douta(w_n2779_0[0]),.doutb(w_n2779_0[1]),.din(n2779));
	jspl jspl_w_n2785_0(.douta(w_n2785_0[0]),.doutb(w_n2785_0[1]),.din(n2785));
	jspl jspl_w_n2787_0(.douta(w_n2787_0[0]),.doutb(w_n2787_0[1]),.din(n2787));
	jspl3 jspl3_w_n2788_0(.douta(w_n2788_0[0]),.doutb(w_n2788_0[1]),.doutc(w_n2788_0[2]),.din(n2788));
	jspl jspl_w_n2792_0(.douta(w_n2792_0[0]),.doutb(w_n2792_0[1]),.din(n2792));
	jspl jspl_w_n2793_0(.douta(w_n2793_0[0]),.doutb(w_n2793_0[1]),.din(n2793));
	jspl3 jspl3_w_n2794_0(.douta(w_n2794_0[0]),.doutb(w_n2794_0[1]),.doutc(w_n2794_0[2]),.din(n2794));
	jspl jspl_w_n2796_0(.douta(w_n2796_0[0]),.doutb(w_n2796_0[1]),.din(n2796));
	jspl jspl_w_n2801_0(.douta(w_n2801_0[0]),.doutb(w_n2801_0[1]),.din(n2801));
	jspl jspl_w_n2803_0(.douta(w_n2803_0[0]),.doutb(w_n2803_0[1]),.din(n2803));
	jspl jspl_w_n2804_0(.douta(w_n2804_0[0]),.doutb(w_n2804_0[1]),.din(n2804));
	jspl3 jspl3_w_n2805_0(.douta(w_n2805_0[0]),.doutb(w_n2805_0[1]),.doutc(w_n2805_0[2]),.din(n2805));
	jspl jspl_w_n2806_0(.douta(w_n2806_0[0]),.doutb(w_n2806_0[1]),.din(n2806));
	jspl jspl_w_n2810_0(.douta(w_n2810_0[0]),.doutb(w_n2810_0[1]),.din(n2810));
	jspl jspl_w_n2816_0(.douta(w_n2816_0[0]),.doutb(w_n2816_0[1]),.din(n2816));
	jspl jspl_w_n2817_0(.douta(w_n2817_0[0]),.doutb(w_n2817_0[1]),.din(n2817));
	jspl jspl_w_n2819_0(.douta(w_n2819_0[0]),.doutb(w_n2819_0[1]),.din(n2819));
	jspl jspl_w_n2821_0(.douta(w_n2821_0[0]),.doutb(w_n2821_0[1]),.din(n2821));
	jspl jspl_w_n2824_0(.douta(w_n2824_0[0]),.doutb(w_n2824_0[1]),.din(n2824));
	jspl jspl_w_n2830_0(.douta(w_n2830_0[0]),.doutb(w_n2830_0[1]),.din(n2830));
	jspl jspl_w_n2832_0(.douta(w_n2832_0[0]),.doutb(w_n2832_0[1]),.din(n2832));
	jspl3 jspl3_w_n2833_0(.douta(w_n2833_0[0]),.doutb(w_n2833_0[1]),.doutc(w_n2833_0[2]),.din(n2833));
	jspl jspl_w_n2837_0(.douta(w_n2837_0[0]),.doutb(w_n2837_0[1]),.din(n2837));
	jspl jspl_w_n2838_0(.douta(w_n2838_0[0]),.doutb(w_n2838_0[1]),.din(n2838));
	jspl3 jspl3_w_n2839_0(.douta(w_n2839_0[0]),.doutb(w_n2839_0[1]),.doutc(w_n2839_0[2]),.din(n2839));
	jspl jspl_w_n2841_0(.douta(w_n2841_0[0]),.doutb(w_n2841_0[1]),.din(n2841));
	jspl jspl_w_n2846_0(.douta(w_n2846_0[0]),.doutb(w_n2846_0[1]),.din(n2846));
	jspl jspl_w_n2848_0(.douta(w_n2848_0[0]),.doutb(w_n2848_0[1]),.din(n2848));
	jspl jspl_w_n2849_0(.douta(w_n2849_0[0]),.doutb(w_n2849_0[1]),.din(n2849));
	jspl3 jspl3_w_n2850_0(.douta(w_n2850_0[0]),.doutb(w_n2850_0[1]),.doutc(w_n2850_0[2]),.din(n2850));
	jspl3 jspl3_w_n2850_1(.douta(w_n2850_1[0]),.doutb(w_n2850_1[1]),.doutc(w_n2850_1[2]),.din(w_n2850_0[0]));
	jspl jspl_w_n2853_0(.douta(w_n2853_0[0]),.doutb(w_n2853_0[1]),.din(n2853));
	jspl3 jspl3_w_n2854_0(.douta(w_n2854_0[0]),.doutb(w_n2854_0[1]),.doutc(w_n2854_0[2]),.din(n2854));
	jspl jspl_w_n2855_0(.douta(w_n2855_0[0]),.doutb(w_n2855_0[1]),.din(n2855));
	jspl jspl_w_n2856_0(.douta(w_n2856_0[0]),.doutb(w_n2856_0[1]),.din(n2856));
	jspl jspl_w_n2862_0(.douta(w_n2862_0[0]),.doutb(w_n2862_0[1]),.din(n2862));
	jspl3 jspl3_w_n2863_0(.douta(w_n2863_0[0]),.doutb(w_n2863_0[1]),.doutc(w_n2863_0[2]),.din(n2863));
	jspl jspl_w_n2864_0(.douta(w_n2864_0[0]),.doutb(w_n2864_0[1]),.din(n2864));
	jspl jspl_w_n2869_0(.douta(w_n2869_0[0]),.doutb(w_n2869_0[1]),.din(n2869));
	jspl3 jspl3_w_n2870_0(.douta(w_n2870_0[0]),.doutb(w_n2870_0[1]),.doutc(w_n2870_0[2]),.din(n2870));
	jspl3 jspl3_w_n2870_1(.douta(w_n2870_1[0]),.doutb(w_n2870_1[1]),.doutc(w_n2870_1[2]),.din(w_n2870_0[0]));
	jspl3 jspl3_w_n2870_2(.douta(w_n2870_2[0]),.doutb(w_n2870_2[1]),.doutc(w_n2870_2[2]),.din(w_n2870_0[1]));
	jspl3 jspl3_w_n2870_3(.douta(w_n2870_3[0]),.doutb(w_n2870_3[1]),.doutc(w_n2870_3[2]),.din(w_n2870_0[2]));
	jspl3 jspl3_w_n2870_4(.douta(w_n2870_4[0]),.doutb(w_n2870_4[1]),.doutc(w_n2870_4[2]),.din(w_n2870_1[0]));
	jspl3 jspl3_w_n2870_5(.douta(w_n2870_5[0]),.doutb(w_n2870_5[1]),.doutc(w_n2870_5[2]),.din(w_n2870_1[1]));
	jspl3 jspl3_w_n2870_6(.douta(w_n2870_6[0]),.doutb(w_n2870_6[1]),.doutc(w_n2870_6[2]),.din(w_n2870_1[2]));
	jspl3 jspl3_w_n2870_7(.douta(w_n2870_7[0]),.doutb(w_n2870_7[1]),.doutc(w_n2870_7[2]),.din(w_n2870_2[0]));
	jspl3 jspl3_w_n2870_8(.douta(w_n2870_8[0]),.doutb(w_n2870_8[1]),.doutc(w_n2870_8[2]),.din(w_n2870_2[1]));
	jspl3 jspl3_w_n2870_9(.douta(w_n2870_9[0]),.doutb(w_n2870_9[1]),.doutc(w_n2870_9[2]),.din(w_n2870_2[2]));
	jspl3 jspl3_w_n2870_10(.douta(w_n2870_10[0]),.doutb(w_n2870_10[1]),.doutc(w_n2870_10[2]),.din(w_n2870_3[0]));
	jspl3 jspl3_w_n2870_11(.douta(w_n2870_11[0]),.doutb(w_n2870_11[1]),.doutc(w_n2870_11[2]),.din(w_n2870_3[1]));
	jspl3 jspl3_w_n2870_12(.douta(w_n2870_12[0]),.doutb(w_n2870_12[1]),.doutc(w_n2870_12[2]),.din(w_n2870_3[2]));
	jspl3 jspl3_w_n2870_13(.douta(w_n2870_13[0]),.doutb(w_n2870_13[1]),.doutc(w_n2870_13[2]),.din(w_n2870_4[0]));
	jspl3 jspl3_w_n2870_14(.douta(w_n2870_14[0]),.doutb(w_n2870_14[1]),.doutc(w_n2870_14[2]),.din(w_n2870_4[1]));
	jspl3 jspl3_w_n2870_15(.douta(w_n2870_15[0]),.doutb(w_n2870_15[1]),.doutc(w_n2870_15[2]),.din(w_n2870_4[2]));
	jspl3 jspl3_w_n2870_16(.douta(w_n2870_16[0]),.doutb(w_n2870_16[1]),.doutc(w_n2870_16[2]),.din(w_n2870_5[0]));
	jspl3 jspl3_w_n2870_17(.douta(w_n2870_17[0]),.doutb(w_n2870_17[1]),.doutc(w_n2870_17[2]),.din(w_n2870_5[1]));
	jspl3 jspl3_w_n2870_18(.douta(w_n2870_18[0]),.doutb(w_n2870_18[1]),.doutc(w_n2870_18[2]),.din(w_n2870_5[2]));
	jspl3 jspl3_w_n2870_19(.douta(w_n2870_19[0]),.doutb(w_n2870_19[1]),.doutc(w_n2870_19[2]),.din(w_n2870_6[0]));
	jspl3 jspl3_w_n2870_20(.douta(w_n2870_20[0]),.doutb(w_n2870_20[1]),.doutc(w_n2870_20[2]),.din(w_n2870_6[1]));
	jspl3 jspl3_w_n2870_21(.douta(w_n2870_21[0]),.doutb(w_n2870_21[1]),.doutc(w_n2870_21[2]),.din(w_n2870_6[2]));
	jspl3 jspl3_w_n2870_22(.douta(w_n2870_22[0]),.doutb(w_n2870_22[1]),.doutc(w_n2870_22[2]),.din(w_n2870_7[0]));
	jspl3 jspl3_w_n2870_23(.douta(w_n2870_23[0]),.doutb(w_n2870_23[1]),.doutc(w_n2870_23[2]),.din(w_n2870_7[1]));
	jspl3 jspl3_w_n2870_24(.douta(w_n2870_24[0]),.doutb(w_n2870_24[1]),.doutc(w_n2870_24[2]),.din(w_n2870_7[2]));
	jspl3 jspl3_w_n2870_25(.douta(w_n2870_25[0]),.doutb(w_n2870_25[1]),.doutc(w_n2870_25[2]),.din(w_n2870_8[0]));
	jspl3 jspl3_w_n2870_26(.douta(w_n2870_26[0]),.doutb(w_n2870_26[1]),.doutc(w_n2870_26[2]),.din(w_n2870_8[1]));
	jspl3 jspl3_w_n2875_0(.douta(w_n2875_0[0]),.doutb(w_n2875_0[1]),.doutc(w_n2875_0[2]),.din(n2875));
	jspl3 jspl3_w_n2875_1(.douta(w_n2875_1[0]),.doutb(w_n2875_1[1]),.doutc(w_n2875_1[2]),.din(w_n2875_0[0]));
	jspl3 jspl3_w_n2875_2(.douta(w_n2875_2[0]),.doutb(w_n2875_2[1]),.doutc(w_n2875_2[2]),.din(w_n2875_0[1]));
	jspl3 jspl3_w_n2875_3(.douta(w_n2875_3[0]),.doutb(w_n2875_3[1]),.doutc(w_n2875_3[2]),.din(w_n2875_0[2]));
	jspl3 jspl3_w_n2875_4(.douta(w_n2875_4[0]),.doutb(w_n2875_4[1]),.doutc(w_n2875_4[2]),.din(w_n2875_1[0]));
	jspl3 jspl3_w_n2875_5(.douta(w_n2875_5[0]),.doutb(w_n2875_5[1]),.doutc(w_n2875_5[2]),.din(w_n2875_1[1]));
	jspl3 jspl3_w_n2875_6(.douta(w_n2875_6[0]),.doutb(w_n2875_6[1]),.doutc(w_n2875_6[2]),.din(w_n2875_1[2]));
	jspl3 jspl3_w_n2875_7(.douta(w_n2875_7[0]),.doutb(w_n2875_7[1]),.doutc(w_n2875_7[2]),.din(w_n2875_2[0]));
	jspl3 jspl3_w_n2875_8(.douta(w_n2875_8[0]),.doutb(w_n2875_8[1]),.doutc(w_n2875_8[2]),.din(w_n2875_2[1]));
	jspl3 jspl3_w_n2875_9(.douta(w_n2875_9[0]),.doutb(w_n2875_9[1]),.doutc(w_n2875_9[2]),.din(w_n2875_2[2]));
	jspl3 jspl3_w_n2875_10(.douta(w_n2875_10[0]),.doutb(w_n2875_10[1]),.doutc(w_n2875_10[2]),.din(w_n2875_3[0]));
	jspl3 jspl3_w_n2875_11(.douta(w_n2875_11[0]),.doutb(w_n2875_11[1]),.doutc(w_n2875_11[2]),.din(w_n2875_3[1]));
	jspl3 jspl3_w_n2875_12(.douta(w_n2875_12[0]),.doutb(w_n2875_12[1]),.doutc(w_n2875_12[2]),.din(w_n2875_3[2]));
	jspl3 jspl3_w_n2875_13(.douta(w_n2875_13[0]),.doutb(w_n2875_13[1]),.doutc(w_n2875_13[2]),.din(w_n2875_4[0]));
	jspl3 jspl3_w_n2875_14(.douta(w_n2875_14[0]),.doutb(w_n2875_14[1]),.doutc(w_n2875_14[2]),.din(w_n2875_4[1]));
	jspl3 jspl3_w_n2875_15(.douta(w_n2875_15[0]),.doutb(w_n2875_15[1]),.doutc(w_n2875_15[2]),.din(w_n2875_4[2]));
	jspl3 jspl3_w_n2875_16(.douta(w_n2875_16[0]),.doutb(w_n2875_16[1]),.doutc(w_n2875_16[2]),.din(w_n2875_5[0]));
	jspl3 jspl3_w_n2875_17(.douta(w_n2875_17[0]),.doutb(w_n2875_17[1]),.doutc(w_n2875_17[2]),.din(w_n2875_5[1]));
	jspl3 jspl3_w_n2875_18(.douta(w_n2875_18[0]),.doutb(w_n2875_18[1]),.doutc(w_n2875_18[2]),.din(w_n2875_5[2]));
	jspl3 jspl3_w_n2875_19(.douta(w_n2875_19[0]),.doutb(w_n2875_19[1]),.doutc(w_n2875_19[2]),.din(w_n2875_6[0]));
	jspl3 jspl3_w_n2875_20(.douta(w_n2875_20[0]),.doutb(w_n2875_20[1]),.doutc(w_n2875_20[2]),.din(w_n2875_6[1]));
	jspl3 jspl3_w_n2875_21(.douta(w_n2875_21[0]),.doutb(w_n2875_21[1]),.doutc(w_n2875_21[2]),.din(w_n2875_6[2]));
	jspl3 jspl3_w_n2875_22(.douta(w_n2875_22[0]),.doutb(w_n2875_22[1]),.doutc(w_n2875_22[2]),.din(w_n2875_7[0]));
	jspl3 jspl3_w_n2875_23(.douta(w_n2875_23[0]),.doutb(w_n2875_23[1]),.doutc(w_n2875_23[2]),.din(w_n2875_7[1]));
	jspl3 jspl3_w_n2875_24(.douta(w_n2875_24[0]),.doutb(w_n2875_24[1]),.doutc(w_n2875_24[2]),.din(w_n2875_7[2]));
	jspl3 jspl3_w_n2875_25(.douta(w_n2875_25[0]),.doutb(w_n2875_25[1]),.doutc(w_n2875_25[2]),.din(w_n2875_8[0]));
	jspl3 jspl3_w_n2875_26(.douta(w_n2875_26[0]),.doutb(w_n2875_26[1]),.doutc(w_n2875_26[2]),.din(w_n2875_8[1]));
	jspl3 jspl3_w_n2875_27(.douta(w_n2875_27[0]),.doutb(w_n2875_27[1]),.doutc(w_n2875_27[2]),.din(w_n2875_8[2]));
	jspl3 jspl3_w_n2875_28(.douta(w_n2875_28[0]),.doutb(w_n2875_28[1]),.doutc(w_n2875_28[2]),.din(w_n2875_9[0]));
	jspl3 jspl3_w_n2875_29(.douta(w_n2875_29[0]),.doutb(w_n2875_29[1]),.doutc(w_n2875_29[2]),.din(w_n2875_9[1]));
	jspl3 jspl3_w_n2875_30(.douta(w_n2875_30[0]),.doutb(w_n2875_30[1]),.doutc(w_n2875_30[2]),.din(w_n2875_9[2]));
	jspl3 jspl3_w_n2875_31(.douta(w_n2875_31[0]),.doutb(w_n2875_31[1]),.doutc(w_n2875_31[2]),.din(w_n2875_10[0]));
	jspl3 jspl3_w_n2875_32(.douta(w_n2875_32[0]),.doutb(w_n2875_32[1]),.doutc(w_n2875_32[2]),.din(w_n2875_10[1]));
	jspl jspl_w_n2875_33(.douta(w_n2875_33[0]),.doutb(w_n2875_33[1]),.din(w_n2875_10[2]));
	jspl3 jspl3_w_n2878_0(.douta(w_n2878_0[0]),.doutb(w_n2878_0[1]),.doutc(w_n2878_0[2]),.din(n2878));
	jspl jspl_w_n2878_1(.douta(w_n2878_1[0]),.doutb(w_n2878_1[1]),.din(w_n2878_0[0]));
	jspl3 jspl3_w_n2879_0(.douta(w_n2879_0[0]),.doutb(w_n2879_0[1]),.doutc(w_n2879_0[2]),.din(n2879));
	jspl3 jspl3_w_n2883_0(.douta(w_n2883_0[0]),.doutb(w_n2883_0[1]),.doutc(w_n2883_0[2]),.din(n2883));
	jspl jspl_w_n2884_0(.douta(w_n2884_0[0]),.doutb(w_n2884_0[1]),.din(n2884));
	jspl jspl_w_n2885_0(.douta(w_n2885_0[0]),.doutb(w_n2885_0[1]),.din(n2885));
	jspl jspl_w_n2886_0(.douta(w_n2886_0[0]),.doutb(w_n2886_0[1]),.din(n2886));
	jspl jspl_w_n2888_0(.douta(w_n2888_0[0]),.doutb(w_n2888_0[1]),.din(n2888));
	jspl jspl_w_n2890_0(.douta(w_n2890_0[0]),.doutb(w_n2890_0[1]),.din(n2890));
	jspl jspl_w_n2892_0(.douta(w_n2892_0[0]),.doutb(w_n2892_0[1]),.din(n2892));
	jspl jspl_w_n2895_0(.douta(w_n2895_0[0]),.doutb(w_n2895_0[1]),.din(n2895));
	jspl jspl_w_n2900_0(.douta(w_n2900_0[0]),.doutb(w_n2900_0[1]),.din(n2900));
	jspl3 jspl3_w_n2902_0(.douta(w_n2902_0[0]),.doutb(w_n2902_0[1]),.doutc(w_n2902_0[2]),.din(n2902));
	jspl jspl_w_n2903_0(.douta(w_n2903_0[0]),.doutb(w_n2903_0[1]),.din(n2903));
	jspl jspl_w_n2907_0(.douta(w_n2907_0[0]),.doutb(w_n2907_0[1]),.din(n2907));
	jspl jspl_w_n2908_0(.douta(w_n2908_0[0]),.doutb(w_n2908_0[1]),.din(n2908));
	jspl jspl_w_n2910_0(.douta(w_n2910_0[0]),.doutb(w_n2910_0[1]),.din(n2910));
	jspl jspl_w_n2914_0(.douta(w_n2914_0[0]),.doutb(w_n2914_0[1]),.din(n2914));
	jspl jspl_w_n2916_0(.douta(w_n2916_0[0]),.doutb(w_n2916_0[1]),.din(n2916));
	jspl jspl_w_n2917_0(.douta(w_n2917_0[0]),.doutb(w_n2917_0[1]),.din(n2917));
	jspl3 jspl3_w_n2918_0(.douta(w_n2918_0[0]),.doutb(w_n2918_0[1]),.doutc(w_n2918_0[2]),.din(n2918));
	jspl jspl_w_n2919_0(.douta(w_n2919_0[0]),.doutb(w_n2919_0[1]),.din(n2919));
	jspl jspl_w_n2923_0(.douta(w_n2923_0[0]),.doutb(w_n2923_0[1]),.din(n2923));
	jspl jspl_w_n2925_0(.douta(w_n2925_0[0]),.doutb(w_n2925_0[1]),.din(n2925));
	jspl jspl_w_n2927_0(.douta(w_n2927_0[0]),.doutb(w_n2927_0[1]),.din(n2927));
	jspl jspl_w_n2929_0(.douta(w_n2929_0[0]),.doutb(w_n2929_0[1]),.din(n2929));
	jspl jspl_w_n2931_0(.douta(w_n2931_0[0]),.doutb(w_n2931_0[1]),.din(n2931));
	jspl jspl_w_n2937_0(.douta(w_n2937_0[0]),.doutb(w_n2937_0[1]),.din(n2937));
	jspl3 jspl3_w_n2939_0(.douta(w_n2939_0[0]),.doutb(w_n2939_0[1]),.doutc(w_n2939_0[2]),.din(n2939));
	jspl jspl_w_n2940_0(.douta(w_n2940_0[0]),.doutb(w_n2940_0[1]),.din(n2940));
	jspl jspl_w_n2945_0(.douta(w_n2945_0[0]),.doutb(w_n2945_0[1]),.din(n2945));
	jspl jspl_w_n2947_0(.douta(w_n2947_0[0]),.doutb(w_n2947_0[1]),.din(n2947));
	jspl jspl_w_n2949_0(.douta(w_n2949_0[0]),.doutb(w_n2949_0[1]),.din(n2949));
	jspl jspl_w_n2953_0(.douta(w_n2953_0[0]),.doutb(w_n2953_0[1]),.din(n2953));
	jspl jspl_w_n2955_0(.douta(w_n2955_0[0]),.doutb(w_n2955_0[1]),.din(n2955));
	jspl jspl_w_n2956_0(.douta(w_n2956_0[0]),.doutb(w_n2956_0[1]),.din(n2956));
	jspl3 jspl3_w_n2957_0(.douta(w_n2957_0[0]),.doutb(w_n2957_0[1]),.doutc(w_n2957_0[2]),.din(n2957));
	jspl jspl_w_n2958_0(.douta(w_n2958_0[0]),.doutb(w_n2958_0[1]),.din(n2958));
	jspl jspl_w_n2964_0(.douta(w_n2964_0[0]),.doutb(w_n2964_0[1]),.din(n2964));
	jspl jspl_w_n2965_0(.douta(w_n2965_0[0]),.doutb(w_n2965_0[1]),.din(n2965));
	jspl jspl_w_n2967_0(.douta(w_n2967_0[0]),.doutb(w_n2967_0[1]),.din(n2967));
	jspl jspl_w_n2969_0(.douta(w_n2969_0[0]),.doutb(w_n2969_0[1]),.din(n2969));
	jspl jspl_w_n2971_0(.douta(w_n2971_0[0]),.doutb(w_n2971_0[1]),.din(n2971));
	jspl jspl_w_n2977_0(.douta(w_n2977_0[0]),.doutb(w_n2977_0[1]),.din(n2977));
	jspl jspl_w_n2979_0(.douta(w_n2979_0[0]),.doutb(w_n2979_0[1]),.din(n2979));
	jspl3 jspl3_w_n2980_0(.douta(w_n2980_0[0]),.doutb(w_n2980_0[1]),.doutc(w_n2980_0[2]),.din(n2980));
	jspl jspl_w_n2983_0(.douta(w_n2983_0[0]),.doutb(w_n2983_0[1]),.din(n2983));
	jspl jspl_w_n2984_0(.douta(w_n2984_0[0]),.doutb(w_n2984_0[1]),.din(n2984));
	jspl3 jspl3_w_n2985_0(.douta(w_n2985_0[0]),.doutb(w_n2985_0[1]),.doutc(w_n2985_0[2]),.din(n2985));
	jspl jspl_w_n2987_0(.douta(w_n2987_0[0]),.doutb(w_n2987_0[1]),.din(n2987));
	jspl jspl_w_n2991_0(.douta(w_n2991_0[0]),.doutb(w_n2991_0[1]),.din(n2991));
	jspl jspl_w_n2993_0(.douta(w_n2993_0[0]),.doutb(w_n2993_0[1]),.din(n2993));
	jspl jspl_w_n2994_0(.douta(w_n2994_0[0]),.doutb(w_n2994_0[1]),.din(n2994));
	jspl3 jspl3_w_n2995_0(.douta(w_n2995_0[0]),.doutb(w_n2995_0[1]),.doutc(w_n2995_0[2]),.din(n2995));
	jspl jspl_w_n2996_0(.douta(w_n2996_0[0]),.doutb(w_n2996_0[1]),.din(n2996));
	jspl jspl_w_n2999_0(.douta(w_n2999_0[0]),.doutb(w_n2999_0[1]),.din(n2999));
	jspl jspl_w_n3005_0(.douta(w_n3005_0[0]),.doutb(w_n3005_0[1]),.din(n3005));
	jspl jspl_w_n3006_0(.douta(w_n3006_0[0]),.doutb(w_n3006_0[1]),.din(n3006));
	jspl jspl_w_n3008_0(.douta(w_n3008_0[0]),.doutb(w_n3008_0[1]),.din(n3008));
	jspl jspl_w_n3010_0(.douta(w_n3010_0[0]),.doutb(w_n3010_0[1]),.din(n3010));
	jspl jspl_w_n3012_0(.douta(w_n3012_0[0]),.doutb(w_n3012_0[1]),.din(n3012));
	jspl jspl_w_n3018_0(.douta(w_n3018_0[0]),.doutb(w_n3018_0[1]),.din(n3018));
	jspl jspl_w_n3020_0(.douta(w_n3020_0[0]),.doutb(w_n3020_0[1]),.din(n3020));
	jspl3 jspl3_w_n3021_0(.douta(w_n3021_0[0]),.doutb(w_n3021_0[1]),.doutc(w_n3021_0[2]),.din(n3021));
	jspl jspl_w_n3024_0(.douta(w_n3024_0[0]),.doutb(w_n3024_0[1]),.din(n3024));
	jspl jspl_w_n3025_0(.douta(w_n3025_0[0]),.doutb(w_n3025_0[1]),.din(n3025));
	jspl3 jspl3_w_n3026_0(.douta(w_n3026_0[0]),.doutb(w_n3026_0[1]),.doutc(w_n3026_0[2]),.din(n3026));
	jspl jspl_w_n3028_0(.douta(w_n3028_0[0]),.doutb(w_n3028_0[1]),.din(n3028));
	jspl jspl_w_n3032_0(.douta(w_n3032_0[0]),.doutb(w_n3032_0[1]),.din(n3032));
	jspl jspl_w_n3034_0(.douta(w_n3034_0[0]),.doutb(w_n3034_0[1]),.din(n3034));
	jspl jspl_w_n3035_0(.douta(w_n3035_0[0]),.doutb(w_n3035_0[1]),.din(n3035));
	jspl3 jspl3_w_n3036_0(.douta(w_n3036_0[0]),.doutb(w_n3036_0[1]),.doutc(w_n3036_0[2]),.din(n3036));
	jspl jspl_w_n3037_0(.douta(w_n3037_0[0]),.doutb(w_n3037_0[1]),.din(n3037));
	jspl jspl_w_n3040_0(.douta(w_n3040_0[0]),.doutb(w_n3040_0[1]),.din(n3040));
	jspl jspl_w_n3046_0(.douta(w_n3046_0[0]),.doutb(w_n3046_0[1]),.din(n3046));
	jspl jspl_w_n3047_0(.douta(w_n3047_0[0]),.doutb(w_n3047_0[1]),.din(n3047));
	jspl jspl_w_n3049_0(.douta(w_n3049_0[0]),.doutb(w_n3049_0[1]),.din(n3049));
	jspl jspl_w_n3051_0(.douta(w_n3051_0[0]),.doutb(w_n3051_0[1]),.din(n3051));
	jspl jspl_w_n3053_0(.douta(w_n3053_0[0]),.doutb(w_n3053_0[1]),.din(n3053));
	jspl jspl_w_n3059_0(.douta(w_n3059_0[0]),.doutb(w_n3059_0[1]),.din(n3059));
	jspl jspl_w_n3061_0(.douta(w_n3061_0[0]),.doutb(w_n3061_0[1]),.din(n3061));
	jspl3 jspl3_w_n3062_0(.douta(w_n3062_0[0]),.doutb(w_n3062_0[1]),.doutc(w_n3062_0[2]),.din(n3062));
	jspl jspl_w_n3065_0(.douta(w_n3065_0[0]),.doutb(w_n3065_0[1]),.din(n3065));
	jspl jspl_w_n3066_0(.douta(w_n3066_0[0]),.doutb(w_n3066_0[1]),.din(n3066));
	jspl3 jspl3_w_n3067_0(.douta(w_n3067_0[0]),.doutb(w_n3067_0[1]),.doutc(w_n3067_0[2]),.din(n3067));
	jspl jspl_w_n3069_0(.douta(w_n3069_0[0]),.doutb(w_n3069_0[1]),.din(n3069));
	jspl jspl_w_n3073_0(.douta(w_n3073_0[0]),.doutb(w_n3073_0[1]),.din(n3073));
	jspl jspl_w_n3075_0(.douta(w_n3075_0[0]),.doutb(w_n3075_0[1]),.din(n3075));
	jspl jspl_w_n3076_0(.douta(w_n3076_0[0]),.doutb(w_n3076_0[1]),.din(n3076));
	jspl3 jspl3_w_n3077_0(.douta(w_n3077_0[0]),.doutb(w_n3077_0[1]),.doutc(w_n3077_0[2]),.din(n3077));
	jspl jspl_w_n3081_0(.douta(w_n3081_0[0]),.doutb(w_n3081_0[1]),.din(n3081));
	jspl jspl_w_n3087_0(.douta(w_n3087_0[0]),.doutb(w_n3087_0[1]),.din(n3087));
	jspl3 jspl3_w_n3089_0(.douta(w_n3089_0[0]),.doutb(w_n3089_0[1]),.doutc(w_n3089_0[2]),.din(n3089));
	jspl jspl_w_n3091_0(.douta(w_n3091_0[0]),.doutb(w_n3091_0[1]),.din(n3091));
	jspl3 jspl3_w_n3096_0(.douta(w_n3096_0[0]),.doutb(w_n3096_0[1]),.doutc(w_n3096_0[2]),.din(n3096));
	jspl jspl_w_n3097_0(.douta(w_n3097_0[0]),.doutb(w_n3097_0[1]),.din(n3097));
	jspl jspl_w_n3098_0(.douta(w_n3098_0[0]),.doutb(w_n3098_0[1]),.din(n3098));
	jspl jspl_w_n3103_0(.douta(w_n3103_0[0]),.doutb(w_n3103_0[1]),.din(n3103));
	jspl3 jspl3_w_n3104_0(.douta(w_n3104_0[0]),.doutb(w_n3104_0[1]),.doutc(w_n3104_0[2]),.din(n3104));
	jspl jspl_w_n3109_0(.douta(w_n3109_0[0]),.doutb(w_n3109_0[1]),.din(n3109));
	jspl3 jspl3_w_n3115_0(.douta(w_n3115_0[0]),.doutb(w_n3115_0[1]),.doutc(w_n3115_0[2]),.din(n3115));
	jspl jspl_w_n3115_1(.douta(w_n3115_1[0]),.doutb(w_n3115_1[1]),.din(w_n3115_0[0]));
	jspl jspl_w_n3116_0(.douta(w_n3116_0[0]),.doutb(w_n3116_0[1]),.din(n3116));
	jspl3 jspl3_w_n3119_0(.douta(w_n3119_0[0]),.doutb(w_n3119_0[1]),.doutc(w_n3119_0[2]),.din(n3119));
	jspl jspl_w_n3120_0(.douta(w_n3120_0[0]),.doutb(w_n3120_0[1]),.din(n3120));
	jspl jspl_w_n3121_0(.douta(w_n3121_0[0]),.doutb(w_n3121_0[1]),.din(n3121));
	jspl jspl_w_n3122_0(.douta(w_n3122_0[0]),.doutb(w_n3122_0[1]),.din(n3122));
	jspl jspl_w_n3124_0(.douta(w_n3124_0[0]),.doutb(w_n3124_0[1]),.din(n3124));
	jspl jspl_w_n3126_0(.douta(w_n3126_0[0]),.doutb(w_n3126_0[1]),.din(n3126));
	jspl jspl_w_n3128_0(.douta(w_n3128_0[0]),.doutb(w_n3128_0[1]),.din(n3128));
	jspl jspl_w_n3137_0(.douta(w_n3137_0[0]),.doutb(w_n3137_0[1]),.din(n3137));
	jspl3 jspl3_w_n3139_0(.douta(w_n3139_0[0]),.doutb(w_n3139_0[1]),.doutc(w_n3139_0[2]),.din(n3139));
	jspl jspl_w_n3140_0(.douta(w_n3140_0[0]),.doutb(w_n3140_0[1]),.din(n3140));
	jspl jspl_w_n3144_0(.douta(w_n3144_0[0]),.doutb(w_n3144_0[1]),.din(n3144));
	jspl jspl_w_n3146_0(.douta(w_n3146_0[0]),.doutb(w_n3146_0[1]),.din(n3146));
	jspl jspl_w_n3148_0(.douta(w_n3148_0[0]),.doutb(w_n3148_0[1]),.din(n3148));
	jspl jspl_w_n3153_0(.douta(w_n3153_0[0]),.doutb(w_n3153_0[1]),.din(n3153));
	jspl jspl_w_n3155_0(.douta(w_n3155_0[0]),.doutb(w_n3155_0[1]),.din(n3155));
	jspl jspl_w_n3156_0(.douta(w_n3156_0[0]),.doutb(w_n3156_0[1]),.din(n3156));
	jspl3 jspl3_w_n3157_0(.douta(w_n3157_0[0]),.doutb(w_n3157_0[1]),.doutc(w_n3157_0[2]),.din(n3157));
	jspl jspl_w_n3158_0(.douta(w_n3158_0[0]),.doutb(w_n3158_0[1]),.din(n3158));
	jspl jspl_w_n3163_0(.douta(w_n3163_0[0]),.doutb(w_n3163_0[1]),.din(n3163));
	jspl jspl_w_n3164_0(.douta(w_n3164_0[0]),.doutb(w_n3164_0[1]),.din(n3164));
	jspl jspl_w_n3166_0(.douta(w_n3166_0[0]),.doutb(w_n3166_0[1]),.din(n3166));
	jspl jspl_w_n3168_0(.douta(w_n3168_0[0]),.doutb(w_n3168_0[1]),.din(n3168));
	jspl jspl_w_n3171_0(.douta(w_n3171_0[0]),.doutb(w_n3171_0[1]),.din(n3171));
	jspl jspl_w_n3177_0(.douta(w_n3177_0[0]),.doutb(w_n3177_0[1]),.din(n3177));
	jspl3 jspl3_w_n3179_0(.douta(w_n3179_0[0]),.doutb(w_n3179_0[1]),.doutc(w_n3179_0[2]),.din(n3179));
	jspl jspl_w_n3180_0(.douta(w_n3180_0[0]),.doutb(w_n3180_0[1]),.din(n3180));
	jspl jspl_w_n3184_0(.douta(w_n3184_0[0]),.doutb(w_n3184_0[1]),.din(n3184));
	jspl jspl_w_n3185_0(.douta(w_n3185_0[0]),.doutb(w_n3185_0[1]),.din(n3185));
	jspl jspl_w_n3187_0(.douta(w_n3187_0[0]),.doutb(w_n3187_0[1]),.din(n3187));
	jspl jspl_w_n3192_0(.douta(w_n3192_0[0]),.doutb(w_n3192_0[1]),.din(n3192));
	jspl jspl_w_n3194_0(.douta(w_n3194_0[0]),.doutb(w_n3194_0[1]),.din(n3194));
	jspl jspl_w_n3195_0(.douta(w_n3195_0[0]),.doutb(w_n3195_0[1]),.din(n3195));
	jspl3 jspl3_w_n3196_0(.douta(w_n3196_0[0]),.doutb(w_n3196_0[1]),.doutc(w_n3196_0[2]),.din(n3196));
	jspl jspl_w_n3197_0(.douta(w_n3197_0[0]),.doutb(w_n3197_0[1]),.din(n3197));
	jspl jspl_w_n3201_0(.douta(w_n3201_0[0]),.doutb(w_n3201_0[1]),.din(n3201));
	jspl jspl_w_n3202_0(.douta(w_n3202_0[0]),.doutb(w_n3202_0[1]),.din(n3202));
	jspl jspl_w_n3204_0(.douta(w_n3204_0[0]),.doutb(w_n3204_0[1]),.din(n3204));
	jspl jspl_w_n3206_0(.douta(w_n3206_0[0]),.doutb(w_n3206_0[1]),.din(n3206));
	jspl jspl_w_n3209_0(.douta(w_n3209_0[0]),.doutb(w_n3209_0[1]),.din(n3209));
	jspl jspl_w_n3215_0(.douta(w_n3215_0[0]),.doutb(w_n3215_0[1]),.din(n3215));
	jspl jspl_w_n3217_0(.douta(w_n3217_0[0]),.doutb(w_n3217_0[1]),.din(n3217));
	jspl3 jspl3_w_n3218_0(.douta(w_n3218_0[0]),.doutb(w_n3218_0[1]),.doutc(w_n3218_0[2]),.din(n3218));
	jspl jspl_w_n3222_0(.douta(w_n3222_0[0]),.doutb(w_n3222_0[1]),.din(n3222));
	jspl jspl_w_n3223_0(.douta(w_n3223_0[0]),.doutb(w_n3223_0[1]),.din(n3223));
	jspl3 jspl3_w_n3224_0(.douta(w_n3224_0[0]),.doutb(w_n3224_0[1]),.doutc(w_n3224_0[2]),.din(n3224));
	jspl jspl_w_n3226_0(.douta(w_n3226_0[0]),.doutb(w_n3226_0[1]),.din(n3226));
	jspl jspl_w_n3231_0(.douta(w_n3231_0[0]),.doutb(w_n3231_0[1]),.din(n3231));
	jspl jspl_w_n3233_0(.douta(w_n3233_0[0]),.doutb(w_n3233_0[1]),.din(n3233));
	jspl jspl_w_n3234_0(.douta(w_n3234_0[0]),.doutb(w_n3234_0[1]),.din(n3234));
	jspl3 jspl3_w_n3235_0(.douta(w_n3235_0[0]),.doutb(w_n3235_0[1]),.doutc(w_n3235_0[2]),.din(n3235));
	jspl jspl_w_n3236_0(.douta(w_n3236_0[0]),.doutb(w_n3236_0[1]),.din(n3236));
	jspl jspl_w_n3240_0(.douta(w_n3240_0[0]),.doutb(w_n3240_0[1]),.din(n3240));
	jspl jspl_w_n3246_0(.douta(w_n3246_0[0]),.doutb(w_n3246_0[1]),.din(n3246));
	jspl jspl_w_n3247_0(.douta(w_n3247_0[0]),.doutb(w_n3247_0[1]),.din(n3247));
	jspl jspl_w_n3249_0(.douta(w_n3249_0[0]),.doutb(w_n3249_0[1]),.din(n3249));
	jspl jspl_w_n3251_0(.douta(w_n3251_0[0]),.doutb(w_n3251_0[1]),.din(n3251));
	jspl jspl_w_n3254_0(.douta(w_n3254_0[0]),.doutb(w_n3254_0[1]),.din(n3254));
	jspl jspl_w_n3260_0(.douta(w_n3260_0[0]),.doutb(w_n3260_0[1]),.din(n3260));
	jspl jspl_w_n3262_0(.douta(w_n3262_0[0]),.doutb(w_n3262_0[1]),.din(n3262));
	jspl3 jspl3_w_n3263_0(.douta(w_n3263_0[0]),.doutb(w_n3263_0[1]),.doutc(w_n3263_0[2]),.din(n3263));
	jspl jspl_w_n3267_0(.douta(w_n3267_0[0]),.doutb(w_n3267_0[1]),.din(n3267));
	jspl jspl_w_n3268_0(.douta(w_n3268_0[0]),.doutb(w_n3268_0[1]),.din(n3268));
	jspl3 jspl3_w_n3269_0(.douta(w_n3269_0[0]),.doutb(w_n3269_0[1]),.doutc(w_n3269_0[2]),.din(n3269));
	jspl jspl_w_n3271_0(.douta(w_n3271_0[0]),.doutb(w_n3271_0[1]),.din(n3271));
	jspl jspl_w_n3276_0(.douta(w_n3276_0[0]),.doutb(w_n3276_0[1]),.din(n3276));
	jspl jspl_w_n3278_0(.douta(w_n3278_0[0]),.doutb(w_n3278_0[1]),.din(n3278));
	jspl jspl_w_n3279_0(.douta(w_n3279_0[0]),.doutb(w_n3279_0[1]),.din(n3279));
	jspl3 jspl3_w_n3280_0(.douta(w_n3280_0[0]),.doutb(w_n3280_0[1]),.doutc(w_n3280_0[2]),.din(n3280));
	jspl jspl_w_n3281_0(.douta(w_n3281_0[0]),.doutb(w_n3281_0[1]),.din(n3281));
	jspl jspl_w_n3285_0(.douta(w_n3285_0[0]),.doutb(w_n3285_0[1]),.din(n3285));
	jspl jspl_w_n3291_0(.douta(w_n3291_0[0]),.doutb(w_n3291_0[1]),.din(n3291));
	jspl jspl_w_n3292_0(.douta(w_n3292_0[0]),.doutb(w_n3292_0[1]),.din(n3292));
	jspl jspl_w_n3294_0(.douta(w_n3294_0[0]),.doutb(w_n3294_0[1]),.din(n3294));
	jspl jspl_w_n3296_0(.douta(w_n3296_0[0]),.doutb(w_n3296_0[1]),.din(n3296));
	jspl jspl_w_n3299_0(.douta(w_n3299_0[0]),.doutb(w_n3299_0[1]),.din(n3299));
	jspl jspl_w_n3305_0(.douta(w_n3305_0[0]),.doutb(w_n3305_0[1]),.din(n3305));
	jspl jspl_w_n3307_0(.douta(w_n3307_0[0]),.doutb(w_n3307_0[1]),.din(n3307));
	jspl3 jspl3_w_n3308_0(.douta(w_n3308_0[0]),.doutb(w_n3308_0[1]),.doutc(w_n3308_0[2]),.din(n3308));
	jspl jspl_w_n3312_0(.douta(w_n3312_0[0]),.doutb(w_n3312_0[1]),.din(n3312));
	jspl jspl_w_n3313_0(.douta(w_n3313_0[0]),.doutb(w_n3313_0[1]),.din(n3313));
	jspl3 jspl3_w_n3314_0(.douta(w_n3314_0[0]),.doutb(w_n3314_0[1]),.doutc(w_n3314_0[2]),.din(n3314));
	jspl jspl_w_n3316_0(.douta(w_n3316_0[0]),.doutb(w_n3316_0[1]),.din(n3316));
	jspl jspl_w_n3321_0(.douta(w_n3321_0[0]),.doutb(w_n3321_0[1]),.din(n3321));
	jspl jspl_w_n3323_0(.douta(w_n3323_0[0]),.doutb(w_n3323_0[1]),.din(n3323));
	jspl jspl_w_n3324_0(.douta(w_n3324_0[0]),.doutb(w_n3324_0[1]),.din(n3324));
	jspl3 jspl3_w_n3325_0(.douta(w_n3325_0[0]),.doutb(w_n3325_0[1]),.doutc(w_n3325_0[2]),.din(n3325));
	jspl jspl_w_n3326_0(.douta(w_n3326_0[0]),.doutb(w_n3326_0[1]),.din(n3326));
	jspl jspl_w_n3330_0(.douta(w_n3330_0[0]),.doutb(w_n3330_0[1]),.din(n3330));
	jspl jspl_w_n3336_0(.douta(w_n3336_0[0]),.doutb(w_n3336_0[1]),.din(n3336));
	jspl jspl_w_n3337_0(.douta(w_n3337_0[0]),.doutb(w_n3337_0[1]),.din(n3337));
	jspl jspl_w_n3339_0(.douta(w_n3339_0[0]),.doutb(w_n3339_0[1]),.din(n3339));
	jspl jspl_w_n3341_0(.douta(w_n3341_0[0]),.doutb(w_n3341_0[1]),.din(n3341));
	jspl jspl_w_n3344_0(.douta(w_n3344_0[0]),.doutb(w_n3344_0[1]),.din(n3344));
	jspl jspl_w_n3350_0(.douta(w_n3350_0[0]),.doutb(w_n3350_0[1]),.din(n3350));
	jspl3 jspl3_w_n3352_0(.douta(w_n3352_0[0]),.doutb(w_n3352_0[1]),.doutc(w_n3352_0[2]),.din(n3352));
	jspl3 jspl3_w_n3352_1(.douta(w_n3352_1[0]),.doutb(w_n3352_1[1]),.doutc(w_n3352_1[2]),.din(w_n3352_0[0]));
	jspl jspl_w_n3355_0(.douta(w_n3355_0[0]),.doutb(w_n3355_0[1]),.din(n3355));
	jspl3 jspl3_w_n3356_0(.douta(w_n3356_0[0]),.doutb(w_n3356_0[1]),.doutc(w_n3356_0[2]),.din(n3356));
	jspl jspl_w_n3357_0(.douta(w_n3357_0[0]),.doutb(w_n3357_0[1]),.din(n3357));
	jspl jspl_w_n3363_0(.douta(w_n3363_0[0]),.doutb(w_n3363_0[1]),.din(n3363));
	jspl3 jspl3_w_n3364_0(.douta(w_n3364_0[0]),.doutb(w_n3364_0[1]),.doutc(w_n3364_0[2]),.din(n3364));
	jspl jspl_w_n3365_0(.douta(w_n3365_0[0]),.doutb(w_n3365_0[1]),.din(n3365));
	jspl jspl_w_n3370_0(.douta(w_n3370_0[0]),.doutb(w_n3370_0[1]),.din(n3370));
	jspl3 jspl3_w_n3371_0(.douta(w_n3371_0[0]),.doutb(w_n3371_0[1]),.doutc(w_n3371_0[2]),.din(n3371));
	jspl3 jspl3_w_n3371_1(.douta(w_n3371_1[0]),.doutb(w_n3371_1[1]),.doutc(w_n3371_1[2]),.din(w_n3371_0[0]));
	jspl3 jspl3_w_n3371_2(.douta(w_n3371_2[0]),.doutb(w_n3371_2[1]),.doutc(w_n3371_2[2]),.din(w_n3371_0[1]));
	jspl3 jspl3_w_n3371_3(.douta(w_n3371_3[0]),.doutb(w_n3371_3[1]),.doutc(w_n3371_3[2]),.din(w_n3371_0[2]));
	jspl3 jspl3_w_n3371_4(.douta(w_n3371_4[0]),.doutb(w_n3371_4[1]),.doutc(w_n3371_4[2]),.din(w_n3371_1[0]));
	jspl3 jspl3_w_n3371_5(.douta(w_n3371_5[0]),.doutb(w_n3371_5[1]),.doutc(w_n3371_5[2]),.din(w_n3371_1[1]));
	jspl3 jspl3_w_n3371_6(.douta(w_n3371_6[0]),.doutb(w_n3371_6[1]),.doutc(w_n3371_6[2]),.din(w_n3371_1[2]));
	jspl3 jspl3_w_n3371_7(.douta(w_n3371_7[0]),.doutb(w_n3371_7[1]),.doutc(w_n3371_7[2]),.din(w_n3371_2[0]));
	jspl3 jspl3_w_n3371_8(.douta(w_n3371_8[0]),.doutb(w_n3371_8[1]),.doutc(w_n3371_8[2]),.din(w_n3371_2[1]));
	jspl3 jspl3_w_n3371_9(.douta(w_n3371_9[0]),.doutb(w_n3371_9[1]),.doutc(w_n3371_9[2]),.din(w_n3371_2[2]));
	jspl3 jspl3_w_n3371_10(.douta(w_n3371_10[0]),.doutb(w_n3371_10[1]),.doutc(w_n3371_10[2]),.din(w_n3371_3[0]));
	jspl3 jspl3_w_n3371_11(.douta(w_n3371_11[0]),.doutb(w_n3371_11[1]),.doutc(w_n3371_11[2]),.din(w_n3371_3[1]));
	jspl3 jspl3_w_n3371_12(.douta(w_n3371_12[0]),.doutb(w_n3371_12[1]),.doutc(w_n3371_12[2]),.din(w_n3371_3[2]));
	jspl3 jspl3_w_n3371_13(.douta(w_n3371_13[0]),.doutb(w_n3371_13[1]),.doutc(w_n3371_13[2]),.din(w_n3371_4[0]));
	jspl3 jspl3_w_n3371_14(.douta(w_n3371_14[0]),.doutb(w_n3371_14[1]),.doutc(w_n3371_14[2]),.din(w_n3371_4[1]));
	jspl3 jspl3_w_n3371_15(.douta(w_n3371_15[0]),.doutb(w_n3371_15[1]),.doutc(w_n3371_15[2]),.din(w_n3371_4[2]));
	jspl3 jspl3_w_n3371_16(.douta(w_n3371_16[0]),.doutb(w_n3371_16[1]),.doutc(w_n3371_16[2]),.din(w_n3371_5[0]));
	jspl3 jspl3_w_n3371_17(.douta(w_n3371_17[0]),.doutb(w_n3371_17[1]),.doutc(w_n3371_17[2]),.din(w_n3371_5[1]));
	jspl3 jspl3_w_n3371_18(.douta(w_n3371_18[0]),.doutb(w_n3371_18[1]),.doutc(w_n3371_18[2]),.din(w_n3371_5[2]));
	jspl3 jspl3_w_n3371_19(.douta(w_n3371_19[0]),.doutb(w_n3371_19[1]),.doutc(w_n3371_19[2]),.din(w_n3371_6[0]));
	jspl3 jspl3_w_n3371_20(.douta(w_n3371_20[0]),.doutb(w_n3371_20[1]),.doutc(w_n3371_20[2]),.din(w_n3371_6[1]));
	jspl3 jspl3_w_n3371_21(.douta(w_n3371_21[0]),.doutb(w_n3371_21[1]),.doutc(w_n3371_21[2]),.din(w_n3371_6[2]));
	jspl3 jspl3_w_n3371_22(.douta(w_n3371_22[0]),.doutb(w_n3371_22[1]),.doutc(w_n3371_22[2]),.din(w_n3371_7[0]));
	jspl3 jspl3_w_n3371_23(.douta(w_n3371_23[0]),.doutb(w_n3371_23[1]),.doutc(w_n3371_23[2]),.din(w_n3371_7[1]));
	jspl3 jspl3_w_n3371_24(.douta(w_n3371_24[0]),.doutb(w_n3371_24[1]),.doutc(w_n3371_24[2]),.din(w_n3371_7[2]));
	jspl3 jspl3_w_n3371_25(.douta(w_n3371_25[0]),.doutb(w_n3371_25[1]),.doutc(w_n3371_25[2]),.din(w_n3371_8[0]));
	jspl3 jspl3_w_n3376_0(.douta(w_n3376_0[0]),.doutb(w_n3376_0[1]),.doutc(w_n3376_0[2]),.din(n3376));
	jspl3 jspl3_w_n3376_1(.douta(w_n3376_1[0]),.doutb(w_n3376_1[1]),.doutc(w_n3376_1[2]),.din(w_n3376_0[0]));
	jspl3 jspl3_w_n3376_2(.douta(w_n3376_2[0]),.doutb(w_n3376_2[1]),.doutc(w_n3376_2[2]),.din(w_n3376_0[1]));
	jspl3 jspl3_w_n3376_3(.douta(w_n3376_3[0]),.doutb(w_n3376_3[1]),.doutc(w_n3376_3[2]),.din(w_n3376_0[2]));
	jspl3 jspl3_w_n3376_4(.douta(w_n3376_4[0]),.doutb(w_n3376_4[1]),.doutc(w_n3376_4[2]),.din(w_n3376_1[0]));
	jspl3 jspl3_w_n3376_5(.douta(w_n3376_5[0]),.doutb(w_n3376_5[1]),.doutc(w_n3376_5[2]),.din(w_n3376_1[1]));
	jspl3 jspl3_w_n3376_6(.douta(w_n3376_6[0]),.doutb(w_n3376_6[1]),.doutc(w_n3376_6[2]),.din(w_n3376_1[2]));
	jspl3 jspl3_w_n3376_7(.douta(w_n3376_7[0]),.doutb(w_n3376_7[1]),.doutc(w_n3376_7[2]),.din(w_n3376_2[0]));
	jspl3 jspl3_w_n3376_8(.douta(w_n3376_8[0]),.doutb(w_n3376_8[1]),.doutc(w_n3376_8[2]),.din(w_n3376_2[1]));
	jspl3 jspl3_w_n3376_9(.douta(w_n3376_9[0]),.doutb(w_n3376_9[1]),.doutc(w_n3376_9[2]),.din(w_n3376_2[2]));
	jspl3 jspl3_w_n3376_10(.douta(w_n3376_10[0]),.doutb(w_n3376_10[1]),.doutc(w_n3376_10[2]),.din(w_n3376_3[0]));
	jspl3 jspl3_w_n3376_11(.douta(w_n3376_11[0]),.doutb(w_n3376_11[1]),.doutc(w_n3376_11[2]),.din(w_n3376_3[1]));
	jspl3 jspl3_w_n3376_12(.douta(w_n3376_12[0]),.doutb(w_n3376_12[1]),.doutc(w_n3376_12[2]),.din(w_n3376_3[2]));
	jspl3 jspl3_w_n3376_13(.douta(w_n3376_13[0]),.doutb(w_n3376_13[1]),.doutc(w_n3376_13[2]),.din(w_n3376_4[0]));
	jspl3 jspl3_w_n3376_14(.douta(w_n3376_14[0]),.doutb(w_n3376_14[1]),.doutc(w_n3376_14[2]),.din(w_n3376_4[1]));
	jspl3 jspl3_w_n3376_15(.douta(w_n3376_15[0]),.doutb(w_n3376_15[1]),.doutc(w_n3376_15[2]),.din(w_n3376_4[2]));
	jspl3 jspl3_w_n3376_16(.douta(w_n3376_16[0]),.doutb(w_n3376_16[1]),.doutc(w_n3376_16[2]),.din(w_n3376_5[0]));
	jspl3 jspl3_w_n3376_17(.douta(w_n3376_17[0]),.doutb(w_n3376_17[1]),.doutc(w_n3376_17[2]),.din(w_n3376_5[1]));
	jspl3 jspl3_w_n3376_18(.douta(w_n3376_18[0]),.doutb(w_n3376_18[1]),.doutc(w_n3376_18[2]),.din(w_n3376_5[2]));
	jspl3 jspl3_w_n3376_19(.douta(w_n3376_19[0]),.doutb(w_n3376_19[1]),.doutc(w_n3376_19[2]),.din(w_n3376_6[0]));
	jspl3 jspl3_w_n3376_20(.douta(w_n3376_20[0]),.doutb(w_n3376_20[1]),.doutc(w_n3376_20[2]),.din(w_n3376_6[1]));
	jspl3 jspl3_w_n3376_21(.douta(w_n3376_21[0]),.doutb(w_n3376_21[1]),.doutc(w_n3376_21[2]),.din(w_n3376_6[2]));
	jspl3 jspl3_w_n3376_22(.douta(w_n3376_22[0]),.doutb(w_n3376_22[1]),.doutc(w_n3376_22[2]),.din(w_n3376_7[0]));
	jspl3 jspl3_w_n3376_23(.douta(w_n3376_23[0]),.doutb(w_n3376_23[1]),.doutc(w_n3376_23[2]),.din(w_n3376_7[1]));
	jspl3 jspl3_w_n3376_24(.douta(w_n3376_24[0]),.doutb(w_n3376_24[1]),.doutc(w_n3376_24[2]),.din(w_n3376_7[2]));
	jspl3 jspl3_w_n3376_25(.douta(w_n3376_25[0]),.doutb(w_n3376_25[1]),.doutc(w_n3376_25[2]),.din(w_n3376_8[0]));
	jspl3 jspl3_w_n3376_26(.douta(w_n3376_26[0]),.doutb(w_n3376_26[1]),.doutc(w_n3376_26[2]),.din(w_n3376_8[1]));
	jspl3 jspl3_w_n3376_27(.douta(w_n3376_27[0]),.doutb(w_n3376_27[1]),.doutc(w_n3376_27[2]),.din(w_n3376_8[2]));
	jspl3 jspl3_w_n3376_28(.douta(w_n3376_28[0]),.doutb(w_n3376_28[1]),.doutc(w_n3376_28[2]),.din(w_n3376_9[0]));
	jspl3 jspl3_w_n3376_29(.douta(w_n3376_29[0]),.doutb(w_n3376_29[1]),.doutc(w_n3376_29[2]),.din(w_n3376_9[1]));
	jspl3 jspl3_w_n3376_30(.douta(w_n3376_30[0]),.doutb(w_n3376_30[1]),.doutc(w_n3376_30[2]),.din(w_n3376_9[2]));
	jspl3 jspl3_w_n3376_31(.douta(w_n3376_31[0]),.doutb(w_n3376_31[1]),.doutc(w_n3376_31[2]),.din(w_n3376_10[0]));
	jspl3 jspl3_w_n3376_32(.douta(w_n3376_32[0]),.doutb(w_n3376_32[1]),.doutc(w_n3376_32[2]),.din(w_n3376_10[1]));
	jspl jspl_w_n3376_33(.douta(w_n3376_33[0]),.doutb(w_n3376_33[1]),.din(w_n3376_10[2]));
	jspl3 jspl3_w_n3379_0(.douta(w_n3379_0[0]),.doutb(w_n3379_0[1]),.doutc(w_n3379_0[2]),.din(n3379));
	jspl jspl_w_n3379_1(.douta(w_n3379_1[0]),.doutb(w_n3379_1[1]),.din(w_n3379_0[0]));
	jspl3 jspl3_w_n3380_0(.douta(w_n3380_0[0]),.doutb(w_n3380_0[1]),.doutc(w_n3380_0[2]),.din(n3380));
	jspl3 jspl3_w_n3384_0(.douta(w_n3384_0[0]),.doutb(w_n3384_0[1]),.doutc(w_n3384_0[2]),.din(n3384));
	jspl jspl_w_n3385_0(.douta(w_n3385_0[0]),.doutb(w_n3385_0[1]),.din(n3385));
	jspl jspl_w_n3386_0(.douta(w_n3386_0[0]),.doutb(w_n3386_0[1]),.din(n3386));
	jspl jspl_w_n3387_0(.douta(w_n3387_0[0]),.doutb(w_n3387_0[1]),.din(n3387));
	jspl jspl_w_n3389_0(.douta(w_n3389_0[0]),.doutb(w_n3389_0[1]),.din(n3389));
	jspl jspl_w_n3391_0(.douta(w_n3391_0[0]),.doutb(w_n3391_0[1]),.din(n3391));
	jspl jspl_w_n3393_0(.douta(w_n3393_0[0]),.doutb(w_n3393_0[1]),.din(n3393));
	jspl jspl_w_n3396_0(.douta(w_n3396_0[0]),.doutb(w_n3396_0[1]),.din(n3396));
	jspl jspl_w_n3401_0(.douta(w_n3401_0[0]),.doutb(w_n3401_0[1]),.din(n3401));
	jspl3 jspl3_w_n3403_0(.douta(w_n3403_0[0]),.doutb(w_n3403_0[1]),.doutc(w_n3403_0[2]),.din(n3403));
	jspl jspl_w_n3404_0(.douta(w_n3404_0[0]),.doutb(w_n3404_0[1]),.din(n3404));
	jspl jspl_w_n3408_0(.douta(w_n3408_0[0]),.doutb(w_n3408_0[1]),.din(n3408));
	jspl jspl_w_n3409_0(.douta(w_n3409_0[0]),.doutb(w_n3409_0[1]),.din(n3409));
	jspl jspl_w_n3411_0(.douta(w_n3411_0[0]),.doutb(w_n3411_0[1]),.din(n3411));
	jspl jspl_w_n3415_0(.douta(w_n3415_0[0]),.doutb(w_n3415_0[1]),.din(n3415));
	jspl jspl_w_n3417_0(.douta(w_n3417_0[0]),.doutb(w_n3417_0[1]),.din(n3417));
	jspl jspl_w_n3418_0(.douta(w_n3418_0[0]),.doutb(w_n3418_0[1]),.din(n3418));
	jspl3 jspl3_w_n3419_0(.douta(w_n3419_0[0]),.doutb(w_n3419_0[1]),.doutc(w_n3419_0[2]),.din(n3419));
	jspl jspl_w_n3420_0(.douta(w_n3420_0[0]),.doutb(w_n3420_0[1]),.din(n3420));
	jspl jspl_w_n3424_0(.douta(w_n3424_0[0]),.doutb(w_n3424_0[1]),.din(n3424));
	jspl jspl_w_n3426_0(.douta(w_n3426_0[0]),.doutb(w_n3426_0[1]),.din(n3426));
	jspl jspl_w_n3428_0(.douta(w_n3428_0[0]),.doutb(w_n3428_0[1]),.din(n3428));
	jspl jspl_w_n3430_0(.douta(w_n3430_0[0]),.doutb(w_n3430_0[1]),.din(n3430));
	jspl jspl_w_n3432_0(.douta(w_n3432_0[0]),.doutb(w_n3432_0[1]),.din(n3432));
	jspl jspl_w_n3438_0(.douta(w_n3438_0[0]),.doutb(w_n3438_0[1]),.din(n3438));
	jspl3 jspl3_w_n3440_0(.douta(w_n3440_0[0]),.doutb(w_n3440_0[1]),.doutc(w_n3440_0[2]),.din(n3440));
	jspl jspl_w_n3441_0(.douta(w_n3441_0[0]),.doutb(w_n3441_0[1]),.din(n3441));
	jspl jspl_w_n3446_0(.douta(w_n3446_0[0]),.doutb(w_n3446_0[1]),.din(n3446));
	jspl jspl_w_n3448_0(.douta(w_n3448_0[0]),.doutb(w_n3448_0[1]),.din(n3448));
	jspl jspl_w_n3450_0(.douta(w_n3450_0[0]),.doutb(w_n3450_0[1]),.din(n3450));
	jspl jspl_w_n3454_0(.douta(w_n3454_0[0]),.doutb(w_n3454_0[1]),.din(n3454));
	jspl jspl_w_n3456_0(.douta(w_n3456_0[0]),.doutb(w_n3456_0[1]),.din(n3456));
	jspl jspl_w_n3457_0(.douta(w_n3457_0[0]),.doutb(w_n3457_0[1]),.din(n3457));
	jspl3 jspl3_w_n3458_0(.douta(w_n3458_0[0]),.doutb(w_n3458_0[1]),.doutc(w_n3458_0[2]),.din(n3458));
	jspl jspl_w_n3459_0(.douta(w_n3459_0[0]),.doutb(w_n3459_0[1]),.din(n3459));
	jspl jspl_w_n3465_0(.douta(w_n3465_0[0]),.doutb(w_n3465_0[1]),.din(n3465));
	jspl jspl_w_n3466_0(.douta(w_n3466_0[0]),.doutb(w_n3466_0[1]),.din(n3466));
	jspl jspl_w_n3468_0(.douta(w_n3468_0[0]),.doutb(w_n3468_0[1]),.din(n3468));
	jspl jspl_w_n3470_0(.douta(w_n3470_0[0]),.doutb(w_n3470_0[1]),.din(n3470));
	jspl jspl_w_n3472_0(.douta(w_n3472_0[0]),.doutb(w_n3472_0[1]),.din(n3472));
	jspl jspl_w_n3478_0(.douta(w_n3478_0[0]),.doutb(w_n3478_0[1]),.din(n3478));
	jspl jspl_w_n3480_0(.douta(w_n3480_0[0]),.doutb(w_n3480_0[1]),.din(n3480));
	jspl3 jspl3_w_n3481_0(.douta(w_n3481_0[0]),.doutb(w_n3481_0[1]),.doutc(w_n3481_0[2]),.din(n3481));
	jspl jspl_w_n3484_0(.douta(w_n3484_0[0]),.doutb(w_n3484_0[1]),.din(n3484));
	jspl jspl_w_n3485_0(.douta(w_n3485_0[0]),.doutb(w_n3485_0[1]),.din(n3485));
	jspl3 jspl3_w_n3486_0(.douta(w_n3486_0[0]),.doutb(w_n3486_0[1]),.doutc(w_n3486_0[2]),.din(n3486));
	jspl jspl_w_n3488_0(.douta(w_n3488_0[0]),.doutb(w_n3488_0[1]),.din(n3488));
	jspl jspl_w_n3492_0(.douta(w_n3492_0[0]),.doutb(w_n3492_0[1]),.din(n3492));
	jspl jspl_w_n3494_0(.douta(w_n3494_0[0]),.doutb(w_n3494_0[1]),.din(n3494));
	jspl jspl_w_n3495_0(.douta(w_n3495_0[0]),.doutb(w_n3495_0[1]),.din(n3495));
	jspl3 jspl3_w_n3496_0(.douta(w_n3496_0[0]),.doutb(w_n3496_0[1]),.doutc(w_n3496_0[2]),.din(n3496));
	jspl jspl_w_n3497_0(.douta(w_n3497_0[0]),.doutb(w_n3497_0[1]),.din(n3497));
	jspl jspl_w_n3500_0(.douta(w_n3500_0[0]),.doutb(w_n3500_0[1]),.din(n3500));
	jspl jspl_w_n3506_0(.douta(w_n3506_0[0]),.doutb(w_n3506_0[1]),.din(n3506));
	jspl jspl_w_n3507_0(.douta(w_n3507_0[0]),.doutb(w_n3507_0[1]),.din(n3507));
	jspl jspl_w_n3509_0(.douta(w_n3509_0[0]),.doutb(w_n3509_0[1]),.din(n3509));
	jspl jspl_w_n3511_0(.douta(w_n3511_0[0]),.doutb(w_n3511_0[1]),.din(n3511));
	jspl jspl_w_n3513_0(.douta(w_n3513_0[0]),.doutb(w_n3513_0[1]),.din(n3513));
	jspl jspl_w_n3519_0(.douta(w_n3519_0[0]),.doutb(w_n3519_0[1]),.din(n3519));
	jspl jspl_w_n3521_0(.douta(w_n3521_0[0]),.doutb(w_n3521_0[1]),.din(n3521));
	jspl3 jspl3_w_n3522_0(.douta(w_n3522_0[0]),.doutb(w_n3522_0[1]),.doutc(w_n3522_0[2]),.din(n3522));
	jspl jspl_w_n3525_0(.douta(w_n3525_0[0]),.doutb(w_n3525_0[1]),.din(n3525));
	jspl jspl_w_n3526_0(.douta(w_n3526_0[0]),.doutb(w_n3526_0[1]),.din(n3526));
	jspl3 jspl3_w_n3527_0(.douta(w_n3527_0[0]),.doutb(w_n3527_0[1]),.doutc(w_n3527_0[2]),.din(n3527));
	jspl jspl_w_n3529_0(.douta(w_n3529_0[0]),.doutb(w_n3529_0[1]),.din(n3529));
	jspl jspl_w_n3533_0(.douta(w_n3533_0[0]),.doutb(w_n3533_0[1]),.din(n3533));
	jspl jspl_w_n3535_0(.douta(w_n3535_0[0]),.doutb(w_n3535_0[1]),.din(n3535));
	jspl jspl_w_n3536_0(.douta(w_n3536_0[0]),.doutb(w_n3536_0[1]),.din(n3536));
	jspl3 jspl3_w_n3537_0(.douta(w_n3537_0[0]),.doutb(w_n3537_0[1]),.doutc(w_n3537_0[2]),.din(n3537));
	jspl jspl_w_n3538_0(.douta(w_n3538_0[0]),.doutb(w_n3538_0[1]),.din(n3538));
	jspl jspl_w_n3541_0(.douta(w_n3541_0[0]),.doutb(w_n3541_0[1]),.din(n3541));
	jspl jspl_w_n3547_0(.douta(w_n3547_0[0]),.doutb(w_n3547_0[1]),.din(n3547));
	jspl jspl_w_n3548_0(.douta(w_n3548_0[0]),.doutb(w_n3548_0[1]),.din(n3548));
	jspl jspl_w_n3550_0(.douta(w_n3550_0[0]),.doutb(w_n3550_0[1]),.din(n3550));
	jspl jspl_w_n3552_0(.douta(w_n3552_0[0]),.doutb(w_n3552_0[1]),.din(n3552));
	jspl jspl_w_n3554_0(.douta(w_n3554_0[0]),.doutb(w_n3554_0[1]),.din(n3554));
	jspl jspl_w_n3560_0(.douta(w_n3560_0[0]),.doutb(w_n3560_0[1]),.din(n3560));
	jspl jspl_w_n3562_0(.douta(w_n3562_0[0]),.doutb(w_n3562_0[1]),.din(n3562));
	jspl3 jspl3_w_n3563_0(.douta(w_n3563_0[0]),.doutb(w_n3563_0[1]),.doutc(w_n3563_0[2]),.din(n3563));
	jspl jspl_w_n3566_0(.douta(w_n3566_0[0]),.doutb(w_n3566_0[1]),.din(n3566));
	jspl jspl_w_n3567_0(.douta(w_n3567_0[0]),.doutb(w_n3567_0[1]),.din(n3567));
	jspl3 jspl3_w_n3568_0(.douta(w_n3568_0[0]),.doutb(w_n3568_0[1]),.doutc(w_n3568_0[2]),.din(n3568));
	jspl jspl_w_n3570_0(.douta(w_n3570_0[0]),.doutb(w_n3570_0[1]),.din(n3570));
	jspl jspl_w_n3574_0(.douta(w_n3574_0[0]),.doutb(w_n3574_0[1]),.din(n3574));
	jspl jspl_w_n3576_0(.douta(w_n3576_0[0]),.doutb(w_n3576_0[1]),.din(n3576));
	jspl jspl_w_n3577_0(.douta(w_n3577_0[0]),.doutb(w_n3577_0[1]),.din(n3577));
	jspl3 jspl3_w_n3578_0(.douta(w_n3578_0[0]),.doutb(w_n3578_0[1]),.doutc(w_n3578_0[2]),.din(n3578));
	jspl jspl_w_n3579_0(.douta(w_n3579_0[0]),.doutb(w_n3579_0[1]),.din(n3579));
	jspl jspl_w_n3582_0(.douta(w_n3582_0[0]),.doutb(w_n3582_0[1]),.din(n3582));
	jspl jspl_w_n3588_0(.douta(w_n3588_0[0]),.doutb(w_n3588_0[1]),.din(n3588));
	jspl jspl_w_n3589_0(.douta(w_n3589_0[0]),.doutb(w_n3589_0[1]),.din(n3589));
	jspl jspl_w_n3591_0(.douta(w_n3591_0[0]),.doutb(w_n3591_0[1]),.din(n3591));
	jspl jspl_w_n3593_0(.douta(w_n3593_0[0]),.doutb(w_n3593_0[1]),.din(n3593));
	jspl jspl_w_n3595_0(.douta(w_n3595_0[0]),.doutb(w_n3595_0[1]),.din(n3595));
	jspl jspl_w_n3601_0(.douta(w_n3601_0[0]),.doutb(w_n3601_0[1]),.din(n3601));
	jspl3 jspl3_w_n3603_0(.douta(w_n3603_0[0]),.doutb(w_n3603_0[1]),.doutc(w_n3603_0[2]),.din(n3603));
	jspl jspl_w_n3608_0(.douta(w_n3608_0[0]),.doutb(w_n3608_0[1]),.din(n3608));
	jspl3 jspl3_w_n3610_0(.douta(w_n3610_0[0]),.doutb(w_n3610_0[1]),.doutc(w_n3610_0[2]),.din(n3610));
	jspl3 jspl3_w_n3614_0(.douta(w_n3614_0[0]),.doutb(w_n3614_0[1]),.doutc(w_n3614_0[2]),.din(n3614));
	jspl jspl_w_n3615_0(.douta(w_n3615_0[0]),.doutb(w_n3615_0[1]),.din(n3615));
	jspl jspl_w_n3620_0(.douta(w_n3620_0[0]),.doutb(w_n3620_0[1]),.din(n3620));
	jspl3 jspl3_w_n3621_0(.douta(w_n3621_0[0]),.doutb(w_n3621_0[1]),.doutc(w_n3621_0[2]),.din(n3621));
	jspl jspl_w_n3626_0(.douta(w_n3626_0[0]),.doutb(w_n3626_0[1]),.din(n3626));
	jspl3 jspl3_w_n3632_0(.douta(w_n3632_0[0]),.doutb(w_n3632_0[1]),.doutc(w_n3632_0[2]),.din(n3632));
	jspl jspl_w_n3632_1(.douta(w_n3632_1[0]),.doutb(w_n3632_1[1]),.din(w_n3632_0[0]));
	jspl jspl_w_n3633_0(.douta(w_n3633_0[0]),.doutb(w_n3633_0[1]),.din(n3633));
	jspl3 jspl3_w_n3636_0(.douta(w_n3636_0[0]),.doutb(w_n3636_0[1]),.doutc(w_n3636_0[2]),.din(n3636));
	jspl jspl_w_n3637_0(.douta(w_n3637_0[0]),.doutb(w_n3637_0[1]),.din(n3637));
	jspl jspl_w_n3638_0(.douta(w_n3638_0[0]),.doutb(w_n3638_0[1]),.din(n3638));
	jspl jspl_w_n3639_0(.douta(w_n3639_0[0]),.doutb(w_n3639_0[1]),.din(n3639));
	jspl jspl_w_n3641_0(.douta(w_n3641_0[0]),.doutb(w_n3641_0[1]),.din(n3641));
	jspl jspl_w_n3643_0(.douta(w_n3643_0[0]),.doutb(w_n3643_0[1]),.din(n3643));
	jspl jspl_w_n3645_0(.douta(w_n3645_0[0]),.doutb(w_n3645_0[1]),.din(n3645));
	jspl jspl_w_n3654_0(.douta(w_n3654_0[0]),.doutb(w_n3654_0[1]),.din(n3654));
	jspl3 jspl3_w_n3656_0(.douta(w_n3656_0[0]),.doutb(w_n3656_0[1]),.doutc(w_n3656_0[2]),.din(n3656));
	jspl jspl_w_n3657_0(.douta(w_n3657_0[0]),.doutb(w_n3657_0[1]),.din(n3657));
	jspl jspl_w_n3661_0(.douta(w_n3661_0[0]),.doutb(w_n3661_0[1]),.din(n3661));
	jspl jspl_w_n3663_0(.douta(w_n3663_0[0]),.doutb(w_n3663_0[1]),.din(n3663));
	jspl jspl_w_n3665_0(.douta(w_n3665_0[0]),.doutb(w_n3665_0[1]),.din(n3665));
	jspl jspl_w_n3670_0(.douta(w_n3670_0[0]),.doutb(w_n3670_0[1]),.din(n3670));
	jspl jspl_w_n3672_0(.douta(w_n3672_0[0]),.doutb(w_n3672_0[1]),.din(n3672));
	jspl jspl_w_n3673_0(.douta(w_n3673_0[0]),.doutb(w_n3673_0[1]),.din(n3673));
	jspl3 jspl3_w_n3674_0(.douta(w_n3674_0[0]),.doutb(w_n3674_0[1]),.doutc(w_n3674_0[2]),.din(n3674));
	jspl jspl_w_n3675_0(.douta(w_n3675_0[0]),.doutb(w_n3675_0[1]),.din(n3675));
	jspl jspl_w_n3680_0(.douta(w_n3680_0[0]),.doutb(w_n3680_0[1]),.din(n3680));
	jspl jspl_w_n3681_0(.douta(w_n3681_0[0]),.doutb(w_n3681_0[1]),.din(n3681));
	jspl jspl_w_n3683_0(.douta(w_n3683_0[0]),.doutb(w_n3683_0[1]),.din(n3683));
	jspl jspl_w_n3685_0(.douta(w_n3685_0[0]),.doutb(w_n3685_0[1]),.din(n3685));
	jspl jspl_w_n3688_0(.douta(w_n3688_0[0]),.doutb(w_n3688_0[1]),.din(n3688));
	jspl jspl_w_n3694_0(.douta(w_n3694_0[0]),.doutb(w_n3694_0[1]),.din(n3694));
	jspl3 jspl3_w_n3696_0(.douta(w_n3696_0[0]),.doutb(w_n3696_0[1]),.doutc(w_n3696_0[2]),.din(n3696));
	jspl jspl_w_n3697_0(.douta(w_n3697_0[0]),.doutb(w_n3697_0[1]),.din(n3697));
	jspl jspl_w_n3701_0(.douta(w_n3701_0[0]),.doutb(w_n3701_0[1]),.din(n3701));
	jspl jspl_w_n3702_0(.douta(w_n3702_0[0]),.doutb(w_n3702_0[1]),.din(n3702));
	jspl jspl_w_n3704_0(.douta(w_n3704_0[0]),.doutb(w_n3704_0[1]),.din(n3704));
	jspl jspl_w_n3709_0(.douta(w_n3709_0[0]),.doutb(w_n3709_0[1]),.din(n3709));
	jspl jspl_w_n3711_0(.douta(w_n3711_0[0]),.doutb(w_n3711_0[1]),.din(n3711));
	jspl jspl_w_n3712_0(.douta(w_n3712_0[0]),.doutb(w_n3712_0[1]),.din(n3712));
	jspl3 jspl3_w_n3713_0(.douta(w_n3713_0[0]),.doutb(w_n3713_0[1]),.doutc(w_n3713_0[2]),.din(n3713));
	jspl jspl_w_n3714_0(.douta(w_n3714_0[0]),.doutb(w_n3714_0[1]),.din(n3714));
	jspl jspl_w_n3718_0(.douta(w_n3718_0[0]),.doutb(w_n3718_0[1]),.din(n3718));
	jspl jspl_w_n3719_0(.douta(w_n3719_0[0]),.doutb(w_n3719_0[1]),.din(n3719));
	jspl jspl_w_n3721_0(.douta(w_n3721_0[0]),.doutb(w_n3721_0[1]),.din(n3721));
	jspl jspl_w_n3723_0(.douta(w_n3723_0[0]),.doutb(w_n3723_0[1]),.din(n3723));
	jspl jspl_w_n3726_0(.douta(w_n3726_0[0]),.doutb(w_n3726_0[1]),.din(n3726));
	jspl jspl_w_n3732_0(.douta(w_n3732_0[0]),.doutb(w_n3732_0[1]),.din(n3732));
	jspl jspl_w_n3734_0(.douta(w_n3734_0[0]),.doutb(w_n3734_0[1]),.din(n3734));
	jspl3 jspl3_w_n3735_0(.douta(w_n3735_0[0]),.doutb(w_n3735_0[1]),.doutc(w_n3735_0[2]),.din(n3735));
	jspl jspl_w_n3739_0(.douta(w_n3739_0[0]),.doutb(w_n3739_0[1]),.din(n3739));
	jspl jspl_w_n3740_0(.douta(w_n3740_0[0]),.doutb(w_n3740_0[1]),.din(n3740));
	jspl3 jspl3_w_n3741_0(.douta(w_n3741_0[0]),.doutb(w_n3741_0[1]),.doutc(w_n3741_0[2]),.din(n3741));
	jspl jspl_w_n3743_0(.douta(w_n3743_0[0]),.doutb(w_n3743_0[1]),.din(n3743));
	jspl jspl_w_n3748_0(.douta(w_n3748_0[0]),.doutb(w_n3748_0[1]),.din(n3748));
	jspl jspl_w_n3750_0(.douta(w_n3750_0[0]),.doutb(w_n3750_0[1]),.din(n3750));
	jspl jspl_w_n3751_0(.douta(w_n3751_0[0]),.doutb(w_n3751_0[1]),.din(n3751));
	jspl3 jspl3_w_n3752_0(.douta(w_n3752_0[0]),.doutb(w_n3752_0[1]),.doutc(w_n3752_0[2]),.din(n3752));
	jspl jspl_w_n3753_0(.douta(w_n3753_0[0]),.doutb(w_n3753_0[1]),.din(n3753));
	jspl jspl_w_n3757_0(.douta(w_n3757_0[0]),.doutb(w_n3757_0[1]),.din(n3757));
	jspl jspl_w_n3763_0(.douta(w_n3763_0[0]),.doutb(w_n3763_0[1]),.din(n3763));
	jspl jspl_w_n3764_0(.douta(w_n3764_0[0]),.doutb(w_n3764_0[1]),.din(n3764));
	jspl jspl_w_n3766_0(.douta(w_n3766_0[0]),.doutb(w_n3766_0[1]),.din(n3766));
	jspl jspl_w_n3768_0(.douta(w_n3768_0[0]),.doutb(w_n3768_0[1]),.din(n3768));
	jspl jspl_w_n3771_0(.douta(w_n3771_0[0]),.doutb(w_n3771_0[1]),.din(n3771));
	jspl jspl_w_n3777_0(.douta(w_n3777_0[0]),.doutb(w_n3777_0[1]),.din(n3777));
	jspl jspl_w_n3779_0(.douta(w_n3779_0[0]),.doutb(w_n3779_0[1]),.din(n3779));
	jspl3 jspl3_w_n3780_0(.douta(w_n3780_0[0]),.doutb(w_n3780_0[1]),.doutc(w_n3780_0[2]),.din(n3780));
	jspl jspl_w_n3784_0(.douta(w_n3784_0[0]),.doutb(w_n3784_0[1]),.din(n3784));
	jspl jspl_w_n3785_0(.douta(w_n3785_0[0]),.doutb(w_n3785_0[1]),.din(n3785));
	jspl3 jspl3_w_n3786_0(.douta(w_n3786_0[0]),.doutb(w_n3786_0[1]),.doutc(w_n3786_0[2]),.din(n3786));
	jspl jspl_w_n3788_0(.douta(w_n3788_0[0]),.doutb(w_n3788_0[1]),.din(n3788));
	jspl jspl_w_n3793_0(.douta(w_n3793_0[0]),.doutb(w_n3793_0[1]),.din(n3793));
	jspl jspl_w_n3795_0(.douta(w_n3795_0[0]),.doutb(w_n3795_0[1]),.din(n3795));
	jspl jspl_w_n3796_0(.douta(w_n3796_0[0]),.doutb(w_n3796_0[1]),.din(n3796));
	jspl3 jspl3_w_n3797_0(.douta(w_n3797_0[0]),.doutb(w_n3797_0[1]),.doutc(w_n3797_0[2]),.din(n3797));
	jspl jspl_w_n3798_0(.douta(w_n3798_0[0]),.doutb(w_n3798_0[1]),.din(n3798));
	jspl jspl_w_n3802_0(.douta(w_n3802_0[0]),.doutb(w_n3802_0[1]),.din(n3802));
	jspl jspl_w_n3808_0(.douta(w_n3808_0[0]),.doutb(w_n3808_0[1]),.din(n3808));
	jspl jspl_w_n3809_0(.douta(w_n3809_0[0]),.doutb(w_n3809_0[1]),.din(n3809));
	jspl jspl_w_n3811_0(.douta(w_n3811_0[0]),.doutb(w_n3811_0[1]),.din(n3811));
	jspl jspl_w_n3813_0(.douta(w_n3813_0[0]),.doutb(w_n3813_0[1]),.din(n3813));
	jspl jspl_w_n3816_0(.douta(w_n3816_0[0]),.doutb(w_n3816_0[1]),.din(n3816));
	jspl jspl_w_n3822_0(.douta(w_n3822_0[0]),.doutb(w_n3822_0[1]),.din(n3822));
	jspl jspl_w_n3824_0(.douta(w_n3824_0[0]),.doutb(w_n3824_0[1]),.din(n3824));
	jspl3 jspl3_w_n3825_0(.douta(w_n3825_0[0]),.doutb(w_n3825_0[1]),.doutc(w_n3825_0[2]),.din(n3825));
	jspl jspl_w_n3829_0(.douta(w_n3829_0[0]),.doutb(w_n3829_0[1]),.din(n3829));
	jspl jspl_w_n3830_0(.douta(w_n3830_0[0]),.doutb(w_n3830_0[1]),.din(n3830));
	jspl3 jspl3_w_n3831_0(.douta(w_n3831_0[0]),.doutb(w_n3831_0[1]),.doutc(w_n3831_0[2]),.din(n3831));
	jspl jspl_w_n3833_0(.douta(w_n3833_0[0]),.doutb(w_n3833_0[1]),.din(n3833));
	jspl jspl_w_n3838_0(.douta(w_n3838_0[0]),.doutb(w_n3838_0[1]),.din(n3838));
	jspl jspl_w_n3840_0(.douta(w_n3840_0[0]),.doutb(w_n3840_0[1]),.din(n3840));
	jspl jspl_w_n3841_0(.douta(w_n3841_0[0]),.doutb(w_n3841_0[1]),.din(n3841));
	jspl3 jspl3_w_n3842_0(.douta(w_n3842_0[0]),.doutb(w_n3842_0[1]),.doutc(w_n3842_0[2]),.din(n3842));
	jspl jspl_w_n3843_0(.douta(w_n3843_0[0]),.doutb(w_n3843_0[1]),.din(n3843));
	jspl jspl_w_n3847_0(.douta(w_n3847_0[0]),.doutb(w_n3847_0[1]),.din(n3847));
	jspl jspl_w_n3853_0(.douta(w_n3853_0[0]),.doutb(w_n3853_0[1]),.din(n3853));
	jspl jspl_w_n3854_0(.douta(w_n3854_0[0]),.doutb(w_n3854_0[1]),.din(n3854));
	jspl jspl_w_n3856_0(.douta(w_n3856_0[0]),.doutb(w_n3856_0[1]),.din(n3856));
	jspl jspl_w_n3858_0(.douta(w_n3858_0[0]),.doutb(w_n3858_0[1]),.din(n3858));
	jspl jspl_w_n3861_0(.douta(w_n3861_0[0]),.doutb(w_n3861_0[1]),.din(n3861));
	jspl jspl_w_n3867_0(.douta(w_n3867_0[0]),.doutb(w_n3867_0[1]),.din(n3867));
	jspl jspl_w_n3869_0(.douta(w_n3869_0[0]),.doutb(w_n3869_0[1]),.din(n3869));
	jspl3 jspl3_w_n3870_0(.douta(w_n3870_0[0]),.doutb(w_n3870_0[1]),.doutc(w_n3870_0[2]),.din(n3870));
	jspl jspl_w_n3874_0(.douta(w_n3874_0[0]),.doutb(w_n3874_0[1]),.din(n3874));
	jspl jspl_w_n3875_0(.douta(w_n3875_0[0]),.doutb(w_n3875_0[1]),.din(n3875));
	jspl3 jspl3_w_n3876_0(.douta(w_n3876_0[0]),.doutb(w_n3876_0[1]),.doutc(w_n3876_0[2]),.din(n3876));
	jspl jspl_w_n3878_0(.douta(w_n3878_0[0]),.doutb(w_n3878_0[1]),.din(n3878));
	jspl jspl_w_n3883_0(.douta(w_n3883_0[0]),.doutb(w_n3883_0[1]),.din(n3883));
	jspl jspl_w_n3885_0(.douta(w_n3885_0[0]),.doutb(w_n3885_0[1]),.din(n3885));
	jspl jspl_w_n3886_0(.douta(w_n3886_0[0]),.doutb(w_n3886_0[1]),.din(n3886));
	jspl3 jspl3_w_n3887_0(.douta(w_n3887_0[0]),.doutb(w_n3887_0[1]),.doutc(w_n3887_0[2]),.din(n3887));
	jspl3 jspl3_w_n3887_1(.douta(w_n3887_1[0]),.doutb(w_n3887_1[1]),.doutc(w_n3887_1[2]),.din(w_n3887_0[0]));
	jspl jspl_w_n3890_0(.douta(w_n3890_0[0]),.doutb(w_n3890_0[1]),.din(n3890));
	jspl3 jspl3_w_n3891_0(.douta(w_n3891_0[0]),.doutb(w_n3891_0[1]),.doutc(w_n3891_0[2]),.din(n3891));
	jspl jspl_w_n3892_0(.douta(w_n3892_0[0]),.doutb(w_n3892_0[1]),.din(n3892));
	jspl jspl_w_n3893_0(.douta(w_n3893_0[0]),.doutb(w_n3893_0[1]),.din(n3893));
	jspl jspl_w_n3899_0(.douta(w_n3899_0[0]),.doutb(w_n3899_0[1]),.din(n3899));
	jspl3 jspl3_w_n3900_0(.douta(w_n3900_0[0]),.doutb(w_n3900_0[1]),.doutc(w_n3900_0[2]),.din(n3900));
	jspl jspl_w_n3901_0(.douta(w_n3901_0[0]),.doutb(w_n3901_0[1]),.din(n3901));
	jspl jspl_w_n3906_0(.douta(w_n3906_0[0]),.doutb(w_n3906_0[1]),.din(n3906));
	jspl3 jspl3_w_n3907_0(.douta(w_n3907_0[0]),.doutb(w_n3907_0[1]),.doutc(w_n3907_0[2]),.din(n3907));
	jspl3 jspl3_w_n3907_1(.douta(w_n3907_1[0]),.doutb(w_n3907_1[1]),.doutc(w_n3907_1[2]),.din(w_n3907_0[0]));
	jspl3 jspl3_w_n3907_2(.douta(w_n3907_2[0]),.doutb(w_n3907_2[1]),.doutc(w_n3907_2[2]),.din(w_n3907_0[1]));
	jspl3 jspl3_w_n3907_3(.douta(w_n3907_3[0]),.doutb(w_n3907_3[1]),.doutc(w_n3907_3[2]),.din(w_n3907_0[2]));
	jspl3 jspl3_w_n3907_4(.douta(w_n3907_4[0]),.doutb(w_n3907_4[1]),.doutc(w_n3907_4[2]),.din(w_n3907_1[0]));
	jspl3 jspl3_w_n3907_5(.douta(w_n3907_5[0]),.doutb(w_n3907_5[1]),.doutc(w_n3907_5[2]),.din(w_n3907_1[1]));
	jspl3 jspl3_w_n3907_6(.douta(w_n3907_6[0]),.doutb(w_n3907_6[1]),.doutc(w_n3907_6[2]),.din(w_n3907_1[2]));
	jspl3 jspl3_w_n3907_7(.douta(w_n3907_7[0]),.doutb(w_n3907_7[1]),.doutc(w_n3907_7[2]),.din(w_n3907_2[0]));
	jspl3 jspl3_w_n3907_8(.douta(w_n3907_8[0]),.doutb(w_n3907_8[1]),.doutc(w_n3907_8[2]),.din(w_n3907_2[1]));
	jspl3 jspl3_w_n3907_9(.douta(w_n3907_9[0]),.doutb(w_n3907_9[1]),.doutc(w_n3907_9[2]),.din(w_n3907_2[2]));
	jspl3 jspl3_w_n3907_10(.douta(w_n3907_10[0]),.doutb(w_n3907_10[1]),.doutc(w_n3907_10[2]),.din(w_n3907_3[0]));
	jspl3 jspl3_w_n3907_11(.douta(w_n3907_11[0]),.doutb(w_n3907_11[1]),.doutc(w_n3907_11[2]),.din(w_n3907_3[1]));
	jspl3 jspl3_w_n3907_12(.douta(w_n3907_12[0]),.doutb(w_n3907_12[1]),.doutc(w_n3907_12[2]),.din(w_n3907_3[2]));
	jspl3 jspl3_w_n3907_13(.douta(w_n3907_13[0]),.doutb(w_n3907_13[1]),.doutc(w_n3907_13[2]),.din(w_n3907_4[0]));
	jspl3 jspl3_w_n3907_14(.douta(w_n3907_14[0]),.doutb(w_n3907_14[1]),.doutc(w_n3907_14[2]),.din(w_n3907_4[1]));
	jspl3 jspl3_w_n3907_15(.douta(w_n3907_15[0]),.doutb(w_n3907_15[1]),.doutc(w_n3907_15[2]),.din(w_n3907_4[2]));
	jspl3 jspl3_w_n3907_16(.douta(w_n3907_16[0]),.doutb(w_n3907_16[1]),.doutc(w_n3907_16[2]),.din(w_n3907_5[0]));
	jspl3 jspl3_w_n3907_17(.douta(w_n3907_17[0]),.doutb(w_n3907_17[1]),.doutc(w_n3907_17[2]),.din(w_n3907_5[1]));
	jspl3 jspl3_w_n3907_18(.douta(w_n3907_18[0]),.doutb(w_n3907_18[1]),.doutc(w_n3907_18[2]),.din(w_n3907_5[2]));
	jspl3 jspl3_w_n3907_19(.douta(w_n3907_19[0]),.doutb(w_n3907_19[1]),.doutc(w_n3907_19[2]),.din(w_n3907_6[0]));
	jspl3 jspl3_w_n3907_20(.douta(w_n3907_20[0]),.doutb(w_n3907_20[1]),.doutc(w_n3907_20[2]),.din(w_n3907_6[1]));
	jspl3 jspl3_w_n3907_21(.douta(w_n3907_21[0]),.doutb(w_n3907_21[1]),.doutc(w_n3907_21[2]),.din(w_n3907_6[2]));
	jspl3 jspl3_w_n3907_22(.douta(w_n3907_22[0]),.doutb(w_n3907_22[1]),.doutc(w_n3907_22[2]),.din(w_n3907_7[0]));
	jspl3 jspl3_w_n3907_23(.douta(w_n3907_23[0]),.doutb(w_n3907_23[1]),.doutc(w_n3907_23[2]),.din(w_n3907_7[1]));
	jspl jspl_w_n3907_24(.douta(w_n3907_24[0]),.doutb(w_n3907_24[1]),.din(w_n3907_7[2]));
	jspl3 jspl3_w_n3912_0(.douta(w_n3912_0[0]),.doutb(w_n3912_0[1]),.doutc(w_n3912_0[2]),.din(n3912));
	jspl3 jspl3_w_n3912_1(.douta(w_n3912_1[0]),.doutb(w_n3912_1[1]),.doutc(w_n3912_1[2]),.din(w_n3912_0[0]));
	jspl3 jspl3_w_n3912_2(.douta(w_n3912_2[0]),.doutb(w_n3912_2[1]),.doutc(w_n3912_2[2]),.din(w_n3912_0[1]));
	jspl3 jspl3_w_n3912_3(.douta(w_n3912_3[0]),.doutb(w_n3912_3[1]),.doutc(w_n3912_3[2]),.din(w_n3912_0[2]));
	jspl3 jspl3_w_n3912_4(.douta(w_n3912_4[0]),.doutb(w_n3912_4[1]),.doutc(w_n3912_4[2]),.din(w_n3912_1[0]));
	jspl3 jspl3_w_n3912_5(.douta(w_n3912_5[0]),.doutb(w_n3912_5[1]),.doutc(w_n3912_5[2]),.din(w_n3912_1[1]));
	jspl3 jspl3_w_n3912_6(.douta(w_n3912_6[0]),.doutb(w_n3912_6[1]),.doutc(w_n3912_6[2]),.din(w_n3912_1[2]));
	jspl3 jspl3_w_n3912_7(.douta(w_n3912_7[0]),.doutb(w_n3912_7[1]),.doutc(w_n3912_7[2]),.din(w_n3912_2[0]));
	jspl3 jspl3_w_n3912_8(.douta(w_n3912_8[0]),.doutb(w_n3912_8[1]),.doutc(w_n3912_8[2]),.din(w_n3912_2[1]));
	jspl3 jspl3_w_n3912_9(.douta(w_n3912_9[0]),.doutb(w_n3912_9[1]),.doutc(w_n3912_9[2]),.din(w_n3912_2[2]));
	jspl3 jspl3_w_n3912_10(.douta(w_n3912_10[0]),.doutb(w_n3912_10[1]),.doutc(w_n3912_10[2]),.din(w_n3912_3[0]));
	jspl3 jspl3_w_n3912_11(.douta(w_n3912_11[0]),.doutb(w_n3912_11[1]),.doutc(w_n3912_11[2]),.din(w_n3912_3[1]));
	jspl3 jspl3_w_n3912_12(.douta(w_n3912_12[0]),.doutb(w_n3912_12[1]),.doutc(w_n3912_12[2]),.din(w_n3912_3[2]));
	jspl3 jspl3_w_n3912_13(.douta(w_n3912_13[0]),.doutb(w_n3912_13[1]),.doutc(w_n3912_13[2]),.din(w_n3912_4[0]));
	jspl3 jspl3_w_n3912_14(.douta(w_n3912_14[0]),.doutb(w_n3912_14[1]),.doutc(w_n3912_14[2]),.din(w_n3912_4[1]));
	jspl3 jspl3_w_n3912_15(.douta(w_n3912_15[0]),.doutb(w_n3912_15[1]),.doutc(w_n3912_15[2]),.din(w_n3912_4[2]));
	jspl3 jspl3_w_n3912_16(.douta(w_n3912_16[0]),.doutb(w_n3912_16[1]),.doutc(w_n3912_16[2]),.din(w_n3912_5[0]));
	jspl3 jspl3_w_n3912_17(.douta(w_n3912_17[0]),.doutb(w_n3912_17[1]),.doutc(w_n3912_17[2]),.din(w_n3912_5[1]));
	jspl3 jspl3_w_n3912_18(.douta(w_n3912_18[0]),.doutb(w_n3912_18[1]),.doutc(w_n3912_18[2]),.din(w_n3912_5[2]));
	jspl3 jspl3_w_n3912_19(.douta(w_n3912_19[0]),.doutb(w_n3912_19[1]),.doutc(w_n3912_19[2]),.din(w_n3912_6[0]));
	jspl3 jspl3_w_n3912_20(.douta(w_n3912_20[0]),.doutb(w_n3912_20[1]),.doutc(w_n3912_20[2]),.din(w_n3912_6[1]));
	jspl3 jspl3_w_n3912_21(.douta(w_n3912_21[0]),.doutb(w_n3912_21[1]),.doutc(w_n3912_21[2]),.din(w_n3912_6[2]));
	jspl3 jspl3_w_n3912_22(.douta(w_n3912_22[0]),.doutb(w_n3912_22[1]),.doutc(w_n3912_22[2]),.din(w_n3912_7[0]));
	jspl3 jspl3_w_n3912_23(.douta(w_n3912_23[0]),.doutb(w_n3912_23[1]),.doutc(w_n3912_23[2]),.din(w_n3912_7[1]));
	jspl3 jspl3_w_n3912_24(.douta(w_n3912_24[0]),.doutb(w_n3912_24[1]),.doutc(w_n3912_24[2]),.din(w_n3912_7[2]));
	jspl3 jspl3_w_n3912_25(.douta(w_n3912_25[0]),.doutb(w_n3912_25[1]),.doutc(w_n3912_25[2]),.din(w_n3912_8[0]));
	jspl3 jspl3_w_n3912_26(.douta(w_n3912_26[0]),.doutb(w_n3912_26[1]),.doutc(w_n3912_26[2]),.din(w_n3912_8[1]));
	jspl3 jspl3_w_n3912_27(.douta(w_n3912_27[0]),.doutb(w_n3912_27[1]),.doutc(w_n3912_27[2]),.din(w_n3912_8[2]));
	jspl3 jspl3_w_n3912_28(.douta(w_n3912_28[0]),.doutb(w_n3912_28[1]),.doutc(w_n3912_28[2]),.din(w_n3912_9[0]));
	jspl3 jspl3_w_n3912_29(.douta(w_n3912_29[0]),.doutb(w_n3912_29[1]),.doutc(w_n3912_29[2]),.din(w_n3912_9[1]));
	jspl3 jspl3_w_n3912_30(.douta(w_n3912_30[0]),.doutb(w_n3912_30[1]),.doutc(w_n3912_30[2]),.din(w_n3912_9[2]));
	jspl3 jspl3_w_n3912_31(.douta(w_n3912_31[0]),.doutb(w_n3912_31[1]),.doutc(w_n3912_31[2]),.din(w_n3912_10[0]));
	jspl3 jspl3_w_n3915_0(.douta(w_n3915_0[0]),.doutb(w_n3915_0[1]),.doutc(w_n3915_0[2]),.din(n3915));
	jspl jspl_w_n3915_1(.douta(w_n3915_1[0]),.doutb(w_n3915_1[1]),.din(w_n3915_0[0]));
	jspl3 jspl3_w_n3916_0(.douta(w_n3916_0[0]),.doutb(w_n3916_0[1]),.doutc(w_n3916_0[2]),.din(n3916));
	jspl3 jspl3_w_n3920_0(.douta(w_n3920_0[0]),.doutb(w_n3920_0[1]),.doutc(w_n3920_0[2]),.din(n3920));
	jspl jspl_w_n3921_0(.douta(w_n3921_0[0]),.doutb(w_n3921_0[1]),.din(n3921));
	jspl jspl_w_n3922_0(.douta(w_n3922_0[0]),.doutb(w_n3922_0[1]),.din(n3922));
	jspl jspl_w_n3923_0(.douta(w_n3923_0[0]),.doutb(w_n3923_0[1]),.din(n3923));
	jspl jspl_w_n3925_0(.douta(w_n3925_0[0]),.doutb(w_n3925_0[1]),.din(n3925));
	jspl jspl_w_n3927_0(.douta(w_n3927_0[0]),.doutb(w_n3927_0[1]),.din(n3927));
	jspl jspl_w_n3929_0(.douta(w_n3929_0[0]),.doutb(w_n3929_0[1]),.din(n3929));
	jspl jspl_w_n3932_0(.douta(w_n3932_0[0]),.doutb(w_n3932_0[1]),.din(n3932));
	jspl jspl_w_n3937_0(.douta(w_n3937_0[0]),.doutb(w_n3937_0[1]),.din(n3937));
	jspl3 jspl3_w_n3939_0(.douta(w_n3939_0[0]),.doutb(w_n3939_0[1]),.doutc(w_n3939_0[2]),.din(n3939));
	jspl jspl_w_n3940_0(.douta(w_n3940_0[0]),.doutb(w_n3940_0[1]),.din(n3940));
	jspl jspl_w_n3944_0(.douta(w_n3944_0[0]),.doutb(w_n3944_0[1]),.din(n3944));
	jspl jspl_w_n3945_0(.douta(w_n3945_0[0]),.doutb(w_n3945_0[1]),.din(n3945));
	jspl jspl_w_n3947_0(.douta(w_n3947_0[0]),.doutb(w_n3947_0[1]),.din(n3947));
	jspl jspl_w_n3951_0(.douta(w_n3951_0[0]),.doutb(w_n3951_0[1]),.din(n3951));
	jspl jspl_w_n3953_0(.douta(w_n3953_0[0]),.doutb(w_n3953_0[1]),.din(n3953));
	jspl jspl_w_n3954_0(.douta(w_n3954_0[0]),.doutb(w_n3954_0[1]),.din(n3954));
	jspl3 jspl3_w_n3955_0(.douta(w_n3955_0[0]),.doutb(w_n3955_0[1]),.doutc(w_n3955_0[2]),.din(n3955));
	jspl jspl_w_n3956_0(.douta(w_n3956_0[0]),.doutb(w_n3956_0[1]),.din(n3956));
	jspl jspl_w_n3960_0(.douta(w_n3960_0[0]),.doutb(w_n3960_0[1]),.din(n3960));
	jspl jspl_w_n3962_0(.douta(w_n3962_0[0]),.doutb(w_n3962_0[1]),.din(n3962));
	jspl jspl_w_n3964_0(.douta(w_n3964_0[0]),.doutb(w_n3964_0[1]),.din(n3964));
	jspl jspl_w_n3966_0(.douta(w_n3966_0[0]),.doutb(w_n3966_0[1]),.din(n3966));
	jspl jspl_w_n3968_0(.douta(w_n3968_0[0]),.doutb(w_n3968_0[1]),.din(n3968));
	jspl jspl_w_n3974_0(.douta(w_n3974_0[0]),.doutb(w_n3974_0[1]),.din(n3974));
	jspl3 jspl3_w_n3976_0(.douta(w_n3976_0[0]),.doutb(w_n3976_0[1]),.doutc(w_n3976_0[2]),.din(n3976));
	jspl jspl_w_n3977_0(.douta(w_n3977_0[0]),.doutb(w_n3977_0[1]),.din(n3977));
	jspl jspl_w_n3982_0(.douta(w_n3982_0[0]),.doutb(w_n3982_0[1]),.din(n3982));
	jspl jspl_w_n3984_0(.douta(w_n3984_0[0]),.doutb(w_n3984_0[1]),.din(n3984));
	jspl jspl_w_n3986_0(.douta(w_n3986_0[0]),.doutb(w_n3986_0[1]),.din(n3986));
	jspl jspl_w_n3990_0(.douta(w_n3990_0[0]),.doutb(w_n3990_0[1]),.din(n3990));
	jspl jspl_w_n3992_0(.douta(w_n3992_0[0]),.doutb(w_n3992_0[1]),.din(n3992));
	jspl jspl_w_n3993_0(.douta(w_n3993_0[0]),.doutb(w_n3993_0[1]),.din(n3993));
	jspl3 jspl3_w_n3994_0(.douta(w_n3994_0[0]),.doutb(w_n3994_0[1]),.doutc(w_n3994_0[2]),.din(n3994));
	jspl jspl_w_n3995_0(.douta(w_n3995_0[0]),.doutb(w_n3995_0[1]),.din(n3995));
	jspl jspl_w_n4001_0(.douta(w_n4001_0[0]),.doutb(w_n4001_0[1]),.din(n4001));
	jspl jspl_w_n4002_0(.douta(w_n4002_0[0]),.doutb(w_n4002_0[1]),.din(n4002));
	jspl jspl_w_n4004_0(.douta(w_n4004_0[0]),.doutb(w_n4004_0[1]),.din(n4004));
	jspl jspl_w_n4006_0(.douta(w_n4006_0[0]),.doutb(w_n4006_0[1]),.din(n4006));
	jspl jspl_w_n4008_0(.douta(w_n4008_0[0]),.doutb(w_n4008_0[1]),.din(n4008));
	jspl jspl_w_n4014_0(.douta(w_n4014_0[0]),.doutb(w_n4014_0[1]),.din(n4014));
	jspl jspl_w_n4016_0(.douta(w_n4016_0[0]),.doutb(w_n4016_0[1]),.din(n4016));
	jspl3 jspl3_w_n4017_0(.douta(w_n4017_0[0]),.doutb(w_n4017_0[1]),.doutc(w_n4017_0[2]),.din(n4017));
	jspl jspl_w_n4020_0(.douta(w_n4020_0[0]),.doutb(w_n4020_0[1]),.din(n4020));
	jspl jspl_w_n4021_0(.douta(w_n4021_0[0]),.doutb(w_n4021_0[1]),.din(n4021));
	jspl3 jspl3_w_n4022_0(.douta(w_n4022_0[0]),.doutb(w_n4022_0[1]),.doutc(w_n4022_0[2]),.din(n4022));
	jspl jspl_w_n4024_0(.douta(w_n4024_0[0]),.doutb(w_n4024_0[1]),.din(n4024));
	jspl jspl_w_n4028_0(.douta(w_n4028_0[0]),.doutb(w_n4028_0[1]),.din(n4028));
	jspl jspl_w_n4030_0(.douta(w_n4030_0[0]),.doutb(w_n4030_0[1]),.din(n4030));
	jspl jspl_w_n4031_0(.douta(w_n4031_0[0]),.doutb(w_n4031_0[1]),.din(n4031));
	jspl3 jspl3_w_n4032_0(.douta(w_n4032_0[0]),.doutb(w_n4032_0[1]),.doutc(w_n4032_0[2]),.din(n4032));
	jspl jspl_w_n4033_0(.douta(w_n4033_0[0]),.doutb(w_n4033_0[1]),.din(n4033));
	jspl jspl_w_n4036_0(.douta(w_n4036_0[0]),.doutb(w_n4036_0[1]),.din(n4036));
	jspl jspl_w_n4042_0(.douta(w_n4042_0[0]),.doutb(w_n4042_0[1]),.din(n4042));
	jspl jspl_w_n4043_0(.douta(w_n4043_0[0]),.doutb(w_n4043_0[1]),.din(n4043));
	jspl jspl_w_n4045_0(.douta(w_n4045_0[0]),.doutb(w_n4045_0[1]),.din(n4045));
	jspl jspl_w_n4047_0(.douta(w_n4047_0[0]),.doutb(w_n4047_0[1]),.din(n4047));
	jspl jspl_w_n4049_0(.douta(w_n4049_0[0]),.doutb(w_n4049_0[1]),.din(n4049));
	jspl jspl_w_n4055_0(.douta(w_n4055_0[0]),.doutb(w_n4055_0[1]),.din(n4055));
	jspl jspl_w_n4057_0(.douta(w_n4057_0[0]),.doutb(w_n4057_0[1]),.din(n4057));
	jspl3 jspl3_w_n4058_0(.douta(w_n4058_0[0]),.doutb(w_n4058_0[1]),.doutc(w_n4058_0[2]),.din(n4058));
	jspl jspl_w_n4061_0(.douta(w_n4061_0[0]),.doutb(w_n4061_0[1]),.din(n4061));
	jspl jspl_w_n4062_0(.douta(w_n4062_0[0]),.doutb(w_n4062_0[1]),.din(n4062));
	jspl3 jspl3_w_n4063_0(.douta(w_n4063_0[0]),.doutb(w_n4063_0[1]),.doutc(w_n4063_0[2]),.din(n4063));
	jspl jspl_w_n4065_0(.douta(w_n4065_0[0]),.doutb(w_n4065_0[1]),.din(n4065));
	jspl jspl_w_n4069_0(.douta(w_n4069_0[0]),.doutb(w_n4069_0[1]),.din(n4069));
	jspl jspl_w_n4071_0(.douta(w_n4071_0[0]),.doutb(w_n4071_0[1]),.din(n4071));
	jspl jspl_w_n4072_0(.douta(w_n4072_0[0]),.doutb(w_n4072_0[1]),.din(n4072));
	jspl3 jspl3_w_n4073_0(.douta(w_n4073_0[0]),.doutb(w_n4073_0[1]),.doutc(w_n4073_0[2]),.din(n4073));
	jspl jspl_w_n4074_0(.douta(w_n4074_0[0]),.doutb(w_n4074_0[1]),.din(n4074));
	jspl jspl_w_n4077_0(.douta(w_n4077_0[0]),.doutb(w_n4077_0[1]),.din(n4077));
	jspl jspl_w_n4083_0(.douta(w_n4083_0[0]),.doutb(w_n4083_0[1]),.din(n4083));
	jspl jspl_w_n4084_0(.douta(w_n4084_0[0]),.doutb(w_n4084_0[1]),.din(n4084));
	jspl jspl_w_n4086_0(.douta(w_n4086_0[0]),.doutb(w_n4086_0[1]),.din(n4086));
	jspl jspl_w_n4088_0(.douta(w_n4088_0[0]),.doutb(w_n4088_0[1]),.din(n4088));
	jspl jspl_w_n4090_0(.douta(w_n4090_0[0]),.doutb(w_n4090_0[1]),.din(n4090));
	jspl jspl_w_n4096_0(.douta(w_n4096_0[0]),.doutb(w_n4096_0[1]),.din(n4096));
	jspl jspl_w_n4098_0(.douta(w_n4098_0[0]),.doutb(w_n4098_0[1]),.din(n4098));
	jspl3 jspl3_w_n4099_0(.douta(w_n4099_0[0]),.doutb(w_n4099_0[1]),.doutc(w_n4099_0[2]),.din(n4099));
	jspl jspl_w_n4102_0(.douta(w_n4102_0[0]),.doutb(w_n4102_0[1]),.din(n4102));
	jspl jspl_w_n4103_0(.douta(w_n4103_0[0]),.doutb(w_n4103_0[1]),.din(n4103));
	jspl3 jspl3_w_n4104_0(.douta(w_n4104_0[0]),.doutb(w_n4104_0[1]),.doutc(w_n4104_0[2]),.din(n4104));
	jspl jspl_w_n4106_0(.douta(w_n4106_0[0]),.doutb(w_n4106_0[1]),.din(n4106));
	jspl jspl_w_n4110_0(.douta(w_n4110_0[0]),.doutb(w_n4110_0[1]),.din(n4110));
	jspl jspl_w_n4112_0(.douta(w_n4112_0[0]),.doutb(w_n4112_0[1]),.din(n4112));
	jspl jspl_w_n4113_0(.douta(w_n4113_0[0]),.doutb(w_n4113_0[1]),.din(n4113));
	jspl3 jspl3_w_n4114_0(.douta(w_n4114_0[0]),.doutb(w_n4114_0[1]),.doutc(w_n4114_0[2]),.din(n4114));
	jspl jspl_w_n4115_0(.douta(w_n4115_0[0]),.doutb(w_n4115_0[1]),.din(n4115));
	jspl jspl_w_n4118_0(.douta(w_n4118_0[0]),.doutb(w_n4118_0[1]),.din(n4118));
	jspl jspl_w_n4124_0(.douta(w_n4124_0[0]),.doutb(w_n4124_0[1]),.din(n4124));
	jspl jspl_w_n4125_0(.douta(w_n4125_0[0]),.doutb(w_n4125_0[1]),.din(n4125));
	jspl jspl_w_n4127_0(.douta(w_n4127_0[0]),.doutb(w_n4127_0[1]),.din(n4127));
	jspl jspl_w_n4129_0(.douta(w_n4129_0[0]),.doutb(w_n4129_0[1]),.din(n4129));
	jspl jspl_w_n4131_0(.douta(w_n4131_0[0]),.doutb(w_n4131_0[1]),.din(n4131));
	jspl jspl_w_n4137_0(.douta(w_n4137_0[0]),.doutb(w_n4137_0[1]),.din(n4137));
	jspl jspl_w_n4139_0(.douta(w_n4139_0[0]),.doutb(w_n4139_0[1]),.din(n4139));
	jspl3 jspl3_w_n4140_0(.douta(w_n4140_0[0]),.doutb(w_n4140_0[1]),.doutc(w_n4140_0[2]),.din(n4140));
	jspl jspl_w_n4143_0(.douta(w_n4143_0[0]),.doutb(w_n4143_0[1]),.din(n4143));
	jspl jspl_w_n4144_0(.douta(w_n4144_0[0]),.doutb(w_n4144_0[1]),.din(n4144));
	jspl3 jspl3_w_n4145_0(.douta(w_n4145_0[0]),.doutb(w_n4145_0[1]),.doutc(w_n4145_0[2]),.din(n4145));
	jspl jspl_w_n4147_0(.douta(w_n4147_0[0]),.doutb(w_n4147_0[1]),.din(n4147));
	jspl jspl_w_n4151_0(.douta(w_n4151_0[0]),.doutb(w_n4151_0[1]),.din(n4151));
	jspl jspl_w_n4153_0(.douta(w_n4153_0[0]),.doutb(w_n4153_0[1]),.din(n4153));
	jspl jspl_w_n4154_0(.douta(w_n4154_0[0]),.doutb(w_n4154_0[1]),.din(n4154));
	jspl3 jspl3_w_n4155_0(.douta(w_n4155_0[0]),.doutb(w_n4155_0[1]),.doutc(w_n4155_0[2]),.din(n4155));
	jspl jspl_w_n4159_0(.douta(w_n4159_0[0]),.doutb(w_n4159_0[1]),.din(n4159));
	jspl jspl_w_n4165_0(.douta(w_n4165_0[0]),.doutb(w_n4165_0[1]),.din(n4165));
	jspl3 jspl3_w_n4167_0(.douta(w_n4167_0[0]),.doutb(w_n4167_0[1]),.doutc(w_n4167_0[2]),.din(n4167));
	jspl jspl_w_n4169_0(.douta(w_n4169_0[0]),.doutb(w_n4169_0[1]),.din(n4169));
	jspl3 jspl3_w_n4174_0(.douta(w_n4174_0[0]),.doutb(w_n4174_0[1]),.doutc(w_n4174_0[2]),.din(n4174));
	jspl jspl_w_n4175_0(.douta(w_n4175_0[0]),.doutb(w_n4175_0[1]),.din(n4175));
	jspl jspl_w_n4176_0(.douta(w_n4176_0[0]),.doutb(w_n4176_0[1]),.din(n4176));
	jspl jspl_w_n4181_0(.douta(w_n4181_0[0]),.doutb(w_n4181_0[1]),.din(n4181));
	jspl3 jspl3_w_n4182_0(.douta(w_n4182_0[0]),.doutb(w_n4182_0[1]),.doutc(w_n4182_0[2]),.din(n4182));
	jspl jspl_w_n4187_0(.douta(w_n4187_0[0]),.doutb(w_n4187_0[1]),.din(n4187));
	jspl3 jspl3_w_n4193_0(.douta(w_n4193_0[0]),.doutb(w_n4193_0[1]),.doutc(w_n4193_0[2]),.din(n4193));
	jspl jspl_w_n4193_1(.douta(w_n4193_1[0]),.doutb(w_n4193_1[1]),.din(w_n4193_0[0]));
	jspl jspl_w_n4194_0(.douta(w_n4194_0[0]),.doutb(w_n4194_0[1]),.din(n4194));
	jspl3 jspl3_w_n4197_0(.douta(w_n4197_0[0]),.doutb(w_n4197_0[1]),.doutc(w_n4197_0[2]),.din(n4197));
	jspl jspl_w_n4198_0(.douta(w_n4198_0[0]),.doutb(w_n4198_0[1]),.din(n4198));
	jspl jspl_w_n4199_0(.douta(w_n4199_0[0]),.doutb(w_n4199_0[1]),.din(n4199));
	jspl jspl_w_n4200_0(.douta(w_n4200_0[0]),.doutb(w_n4200_0[1]),.din(n4200));
	jspl jspl_w_n4202_0(.douta(w_n4202_0[0]),.doutb(w_n4202_0[1]),.din(n4202));
	jspl jspl_w_n4204_0(.douta(w_n4204_0[0]),.doutb(w_n4204_0[1]),.din(n4204));
	jspl jspl_w_n4206_0(.douta(w_n4206_0[0]),.doutb(w_n4206_0[1]),.din(n4206));
	jspl jspl_w_n4215_0(.douta(w_n4215_0[0]),.doutb(w_n4215_0[1]),.din(n4215));
	jspl3 jspl3_w_n4217_0(.douta(w_n4217_0[0]),.doutb(w_n4217_0[1]),.doutc(w_n4217_0[2]),.din(n4217));
	jspl jspl_w_n4218_0(.douta(w_n4218_0[0]),.doutb(w_n4218_0[1]),.din(n4218));
	jspl jspl_w_n4222_0(.douta(w_n4222_0[0]),.doutb(w_n4222_0[1]),.din(n4222));
	jspl jspl_w_n4224_0(.douta(w_n4224_0[0]),.doutb(w_n4224_0[1]),.din(n4224));
	jspl jspl_w_n4226_0(.douta(w_n4226_0[0]),.doutb(w_n4226_0[1]),.din(n4226));
	jspl jspl_w_n4231_0(.douta(w_n4231_0[0]),.doutb(w_n4231_0[1]),.din(n4231));
	jspl jspl_w_n4233_0(.douta(w_n4233_0[0]),.doutb(w_n4233_0[1]),.din(n4233));
	jspl jspl_w_n4234_0(.douta(w_n4234_0[0]),.doutb(w_n4234_0[1]),.din(n4234));
	jspl3 jspl3_w_n4235_0(.douta(w_n4235_0[0]),.doutb(w_n4235_0[1]),.doutc(w_n4235_0[2]),.din(n4235));
	jspl jspl_w_n4236_0(.douta(w_n4236_0[0]),.doutb(w_n4236_0[1]),.din(n4236));
	jspl jspl_w_n4241_0(.douta(w_n4241_0[0]),.doutb(w_n4241_0[1]),.din(n4241));
	jspl jspl_w_n4242_0(.douta(w_n4242_0[0]),.doutb(w_n4242_0[1]),.din(n4242));
	jspl jspl_w_n4244_0(.douta(w_n4244_0[0]),.doutb(w_n4244_0[1]),.din(n4244));
	jspl jspl_w_n4246_0(.douta(w_n4246_0[0]),.doutb(w_n4246_0[1]),.din(n4246));
	jspl jspl_w_n4249_0(.douta(w_n4249_0[0]),.doutb(w_n4249_0[1]),.din(n4249));
	jspl jspl_w_n4255_0(.douta(w_n4255_0[0]),.doutb(w_n4255_0[1]),.din(n4255));
	jspl3 jspl3_w_n4257_0(.douta(w_n4257_0[0]),.doutb(w_n4257_0[1]),.doutc(w_n4257_0[2]),.din(n4257));
	jspl jspl_w_n4258_0(.douta(w_n4258_0[0]),.doutb(w_n4258_0[1]),.din(n4258));
	jspl jspl_w_n4262_0(.douta(w_n4262_0[0]),.doutb(w_n4262_0[1]),.din(n4262));
	jspl jspl_w_n4263_0(.douta(w_n4263_0[0]),.doutb(w_n4263_0[1]),.din(n4263));
	jspl jspl_w_n4265_0(.douta(w_n4265_0[0]),.doutb(w_n4265_0[1]),.din(n4265));
	jspl jspl_w_n4270_0(.douta(w_n4270_0[0]),.doutb(w_n4270_0[1]),.din(n4270));
	jspl jspl_w_n4272_0(.douta(w_n4272_0[0]),.doutb(w_n4272_0[1]),.din(n4272));
	jspl jspl_w_n4273_0(.douta(w_n4273_0[0]),.doutb(w_n4273_0[1]),.din(n4273));
	jspl3 jspl3_w_n4274_0(.douta(w_n4274_0[0]),.doutb(w_n4274_0[1]),.doutc(w_n4274_0[2]),.din(n4274));
	jspl jspl_w_n4275_0(.douta(w_n4275_0[0]),.doutb(w_n4275_0[1]),.din(n4275));
	jspl jspl_w_n4279_0(.douta(w_n4279_0[0]),.doutb(w_n4279_0[1]),.din(n4279));
	jspl jspl_w_n4280_0(.douta(w_n4280_0[0]),.doutb(w_n4280_0[1]),.din(n4280));
	jspl jspl_w_n4282_0(.douta(w_n4282_0[0]),.doutb(w_n4282_0[1]),.din(n4282));
	jspl jspl_w_n4284_0(.douta(w_n4284_0[0]),.doutb(w_n4284_0[1]),.din(n4284));
	jspl jspl_w_n4287_0(.douta(w_n4287_0[0]),.doutb(w_n4287_0[1]),.din(n4287));
	jspl jspl_w_n4293_0(.douta(w_n4293_0[0]),.doutb(w_n4293_0[1]),.din(n4293));
	jspl jspl_w_n4295_0(.douta(w_n4295_0[0]),.doutb(w_n4295_0[1]),.din(n4295));
	jspl3 jspl3_w_n4296_0(.douta(w_n4296_0[0]),.doutb(w_n4296_0[1]),.doutc(w_n4296_0[2]),.din(n4296));
	jspl jspl_w_n4300_0(.douta(w_n4300_0[0]),.doutb(w_n4300_0[1]),.din(n4300));
	jspl jspl_w_n4301_0(.douta(w_n4301_0[0]),.doutb(w_n4301_0[1]),.din(n4301));
	jspl3 jspl3_w_n4302_0(.douta(w_n4302_0[0]),.doutb(w_n4302_0[1]),.doutc(w_n4302_0[2]),.din(n4302));
	jspl jspl_w_n4304_0(.douta(w_n4304_0[0]),.doutb(w_n4304_0[1]),.din(n4304));
	jspl jspl_w_n4309_0(.douta(w_n4309_0[0]),.doutb(w_n4309_0[1]),.din(n4309));
	jspl jspl_w_n4311_0(.douta(w_n4311_0[0]),.doutb(w_n4311_0[1]),.din(n4311));
	jspl jspl_w_n4312_0(.douta(w_n4312_0[0]),.doutb(w_n4312_0[1]),.din(n4312));
	jspl3 jspl3_w_n4313_0(.douta(w_n4313_0[0]),.doutb(w_n4313_0[1]),.doutc(w_n4313_0[2]),.din(n4313));
	jspl jspl_w_n4314_0(.douta(w_n4314_0[0]),.doutb(w_n4314_0[1]),.din(n4314));
	jspl jspl_w_n4318_0(.douta(w_n4318_0[0]),.doutb(w_n4318_0[1]),.din(n4318));
	jspl jspl_w_n4324_0(.douta(w_n4324_0[0]),.doutb(w_n4324_0[1]),.din(n4324));
	jspl jspl_w_n4325_0(.douta(w_n4325_0[0]),.doutb(w_n4325_0[1]),.din(n4325));
	jspl jspl_w_n4327_0(.douta(w_n4327_0[0]),.doutb(w_n4327_0[1]),.din(n4327));
	jspl jspl_w_n4329_0(.douta(w_n4329_0[0]),.doutb(w_n4329_0[1]),.din(n4329));
	jspl jspl_w_n4332_0(.douta(w_n4332_0[0]),.doutb(w_n4332_0[1]),.din(n4332));
	jspl jspl_w_n4338_0(.douta(w_n4338_0[0]),.doutb(w_n4338_0[1]),.din(n4338));
	jspl jspl_w_n4340_0(.douta(w_n4340_0[0]),.doutb(w_n4340_0[1]),.din(n4340));
	jspl3 jspl3_w_n4341_0(.douta(w_n4341_0[0]),.doutb(w_n4341_0[1]),.doutc(w_n4341_0[2]),.din(n4341));
	jspl jspl_w_n4345_0(.douta(w_n4345_0[0]),.doutb(w_n4345_0[1]),.din(n4345));
	jspl jspl_w_n4346_0(.douta(w_n4346_0[0]),.doutb(w_n4346_0[1]),.din(n4346));
	jspl3 jspl3_w_n4347_0(.douta(w_n4347_0[0]),.doutb(w_n4347_0[1]),.doutc(w_n4347_0[2]),.din(n4347));
	jspl jspl_w_n4349_0(.douta(w_n4349_0[0]),.doutb(w_n4349_0[1]),.din(n4349));
	jspl jspl_w_n4354_0(.douta(w_n4354_0[0]),.doutb(w_n4354_0[1]),.din(n4354));
	jspl jspl_w_n4356_0(.douta(w_n4356_0[0]),.doutb(w_n4356_0[1]),.din(n4356));
	jspl jspl_w_n4357_0(.douta(w_n4357_0[0]),.doutb(w_n4357_0[1]),.din(n4357));
	jspl3 jspl3_w_n4358_0(.douta(w_n4358_0[0]),.doutb(w_n4358_0[1]),.doutc(w_n4358_0[2]),.din(n4358));
	jspl jspl_w_n4359_0(.douta(w_n4359_0[0]),.doutb(w_n4359_0[1]),.din(n4359));
	jspl jspl_w_n4363_0(.douta(w_n4363_0[0]),.doutb(w_n4363_0[1]),.din(n4363));
	jspl jspl_w_n4369_0(.douta(w_n4369_0[0]),.doutb(w_n4369_0[1]),.din(n4369));
	jspl jspl_w_n4370_0(.douta(w_n4370_0[0]),.doutb(w_n4370_0[1]),.din(n4370));
	jspl jspl_w_n4372_0(.douta(w_n4372_0[0]),.doutb(w_n4372_0[1]),.din(n4372));
	jspl jspl_w_n4374_0(.douta(w_n4374_0[0]),.doutb(w_n4374_0[1]),.din(n4374));
	jspl jspl_w_n4377_0(.douta(w_n4377_0[0]),.doutb(w_n4377_0[1]),.din(n4377));
	jspl jspl_w_n4383_0(.douta(w_n4383_0[0]),.doutb(w_n4383_0[1]),.din(n4383));
	jspl jspl_w_n4385_0(.douta(w_n4385_0[0]),.doutb(w_n4385_0[1]),.din(n4385));
	jspl3 jspl3_w_n4386_0(.douta(w_n4386_0[0]),.doutb(w_n4386_0[1]),.doutc(w_n4386_0[2]),.din(n4386));
	jspl jspl_w_n4390_0(.douta(w_n4390_0[0]),.doutb(w_n4390_0[1]),.din(n4390));
	jspl jspl_w_n4391_0(.douta(w_n4391_0[0]),.doutb(w_n4391_0[1]),.din(n4391));
	jspl3 jspl3_w_n4392_0(.douta(w_n4392_0[0]),.doutb(w_n4392_0[1]),.doutc(w_n4392_0[2]),.din(n4392));
	jspl jspl_w_n4394_0(.douta(w_n4394_0[0]),.doutb(w_n4394_0[1]),.din(n4394));
	jspl jspl_w_n4399_0(.douta(w_n4399_0[0]),.doutb(w_n4399_0[1]),.din(n4399));
	jspl jspl_w_n4401_0(.douta(w_n4401_0[0]),.doutb(w_n4401_0[1]),.din(n4401));
	jspl jspl_w_n4402_0(.douta(w_n4402_0[0]),.doutb(w_n4402_0[1]),.din(n4402));
	jspl3 jspl3_w_n4403_0(.douta(w_n4403_0[0]),.doutb(w_n4403_0[1]),.doutc(w_n4403_0[2]),.din(n4403));
	jspl jspl_w_n4404_0(.douta(w_n4404_0[0]),.doutb(w_n4404_0[1]),.din(n4404));
	jspl jspl_w_n4408_0(.douta(w_n4408_0[0]),.doutb(w_n4408_0[1]),.din(n4408));
	jspl jspl_w_n4414_0(.douta(w_n4414_0[0]),.doutb(w_n4414_0[1]),.din(n4414));
	jspl jspl_w_n4415_0(.douta(w_n4415_0[0]),.doutb(w_n4415_0[1]),.din(n4415));
	jspl jspl_w_n4417_0(.douta(w_n4417_0[0]),.doutb(w_n4417_0[1]),.din(n4417));
	jspl jspl_w_n4419_0(.douta(w_n4419_0[0]),.doutb(w_n4419_0[1]),.din(n4419));
	jspl jspl_w_n4422_0(.douta(w_n4422_0[0]),.doutb(w_n4422_0[1]),.din(n4422));
	jspl jspl_w_n4428_0(.douta(w_n4428_0[0]),.doutb(w_n4428_0[1]),.din(n4428));
	jspl jspl_w_n4430_0(.douta(w_n4430_0[0]),.doutb(w_n4430_0[1]),.din(n4430));
	jspl3 jspl3_w_n4431_0(.douta(w_n4431_0[0]),.doutb(w_n4431_0[1]),.doutc(w_n4431_0[2]),.din(n4431));
	jspl jspl_w_n4435_0(.douta(w_n4435_0[0]),.doutb(w_n4435_0[1]),.din(n4435));
	jspl jspl_w_n4436_0(.douta(w_n4436_0[0]),.doutb(w_n4436_0[1]),.din(n4436));
	jspl3 jspl3_w_n4437_0(.douta(w_n4437_0[0]),.doutb(w_n4437_0[1]),.doutc(w_n4437_0[2]),.din(n4437));
	jspl jspl_w_n4439_0(.douta(w_n4439_0[0]),.doutb(w_n4439_0[1]),.din(n4439));
	jspl jspl_w_n4444_0(.douta(w_n4444_0[0]),.doutb(w_n4444_0[1]),.din(n4444));
	jspl jspl_w_n4446_0(.douta(w_n4446_0[0]),.doutb(w_n4446_0[1]),.din(n4446));
	jspl jspl_w_n4447_0(.douta(w_n4447_0[0]),.doutb(w_n4447_0[1]),.din(n4447));
	jspl3 jspl3_w_n4448_0(.douta(w_n4448_0[0]),.doutb(w_n4448_0[1]),.doutc(w_n4448_0[2]),.din(n4448));
	jspl jspl_w_n4449_0(.douta(w_n4449_0[0]),.doutb(w_n4449_0[1]),.din(n4449));
	jspl jspl_w_n4453_0(.douta(w_n4453_0[0]),.doutb(w_n4453_0[1]),.din(n4453));
	jspl jspl_w_n4459_0(.douta(w_n4459_0[0]),.doutb(w_n4459_0[1]),.din(n4459));
	jspl jspl_w_n4460_0(.douta(w_n4460_0[0]),.doutb(w_n4460_0[1]),.din(n4460));
	jspl jspl_w_n4462_0(.douta(w_n4462_0[0]),.doutb(w_n4462_0[1]),.din(n4462));
	jspl jspl_w_n4464_0(.douta(w_n4464_0[0]),.doutb(w_n4464_0[1]),.din(n4464));
	jspl jspl_w_n4467_0(.douta(w_n4467_0[0]),.doutb(w_n4467_0[1]),.din(n4467));
	jspl jspl_w_n4473_0(.douta(w_n4473_0[0]),.doutb(w_n4473_0[1]),.din(n4473));
	jspl3 jspl3_w_n4475_0(.douta(w_n4475_0[0]),.doutb(w_n4475_0[1]),.doutc(w_n4475_0[2]),.din(n4475));
	jspl3 jspl3_w_n4475_1(.douta(w_n4475_1[0]),.doutb(w_n4475_1[1]),.doutc(w_n4475_1[2]),.din(w_n4475_0[0]));
	jspl jspl_w_n4478_0(.douta(w_n4478_0[0]),.doutb(w_n4478_0[1]),.din(n4478));
	jspl3 jspl3_w_n4479_0(.douta(w_n4479_0[0]),.doutb(w_n4479_0[1]),.doutc(w_n4479_0[2]),.din(n4479));
	jspl jspl_w_n4480_0(.douta(w_n4480_0[0]),.doutb(w_n4480_0[1]),.din(n4480));
	jspl jspl_w_n4486_0(.douta(w_n4486_0[0]),.doutb(w_n4486_0[1]),.din(n4486));
	jspl3 jspl3_w_n4487_0(.douta(w_n4487_0[0]),.doutb(w_n4487_0[1]),.doutc(w_n4487_0[2]),.din(n4487));
	jspl jspl_w_n4488_0(.douta(w_n4488_0[0]),.doutb(w_n4488_0[1]),.din(n4488));
	jspl jspl_w_n4493_0(.douta(w_n4493_0[0]),.doutb(w_n4493_0[1]),.din(n4493));
	jspl3 jspl3_w_n4494_0(.douta(w_n4494_0[0]),.doutb(w_n4494_0[1]),.doutc(w_n4494_0[2]),.din(n4494));
	jspl3 jspl3_w_n4494_1(.douta(w_n4494_1[0]),.doutb(w_n4494_1[1]),.doutc(w_n4494_1[2]),.din(w_n4494_0[0]));
	jspl3 jspl3_w_n4494_2(.douta(w_n4494_2[0]),.doutb(w_n4494_2[1]),.doutc(w_n4494_2[2]),.din(w_n4494_0[1]));
	jspl3 jspl3_w_n4494_3(.douta(w_n4494_3[0]),.doutb(w_n4494_3[1]),.doutc(w_n4494_3[2]),.din(w_n4494_0[2]));
	jspl3 jspl3_w_n4494_4(.douta(w_n4494_4[0]),.doutb(w_n4494_4[1]),.doutc(w_n4494_4[2]),.din(w_n4494_1[0]));
	jspl3 jspl3_w_n4494_5(.douta(w_n4494_5[0]),.doutb(w_n4494_5[1]),.doutc(w_n4494_5[2]),.din(w_n4494_1[1]));
	jspl3 jspl3_w_n4494_6(.douta(w_n4494_6[0]),.doutb(w_n4494_6[1]),.doutc(w_n4494_6[2]),.din(w_n4494_1[2]));
	jspl3 jspl3_w_n4494_7(.douta(w_n4494_7[0]),.doutb(w_n4494_7[1]),.doutc(w_n4494_7[2]),.din(w_n4494_2[0]));
	jspl3 jspl3_w_n4494_8(.douta(w_n4494_8[0]),.doutb(w_n4494_8[1]),.doutc(w_n4494_8[2]),.din(w_n4494_2[1]));
	jspl3 jspl3_w_n4494_9(.douta(w_n4494_9[0]),.doutb(w_n4494_9[1]),.doutc(w_n4494_9[2]),.din(w_n4494_2[2]));
	jspl3 jspl3_w_n4494_10(.douta(w_n4494_10[0]),.doutb(w_n4494_10[1]),.doutc(w_n4494_10[2]),.din(w_n4494_3[0]));
	jspl3 jspl3_w_n4494_11(.douta(w_n4494_11[0]),.doutb(w_n4494_11[1]),.doutc(w_n4494_11[2]),.din(w_n4494_3[1]));
	jspl3 jspl3_w_n4494_12(.douta(w_n4494_12[0]),.doutb(w_n4494_12[1]),.doutc(w_n4494_12[2]),.din(w_n4494_3[2]));
	jspl3 jspl3_w_n4494_13(.douta(w_n4494_13[0]),.doutb(w_n4494_13[1]),.doutc(w_n4494_13[2]),.din(w_n4494_4[0]));
	jspl3 jspl3_w_n4494_14(.douta(w_n4494_14[0]),.doutb(w_n4494_14[1]),.doutc(w_n4494_14[2]),.din(w_n4494_4[1]));
	jspl3 jspl3_w_n4494_15(.douta(w_n4494_15[0]),.doutb(w_n4494_15[1]),.doutc(w_n4494_15[2]),.din(w_n4494_4[2]));
	jspl3 jspl3_w_n4494_16(.douta(w_n4494_16[0]),.doutb(w_n4494_16[1]),.doutc(w_n4494_16[2]),.din(w_n4494_5[0]));
	jspl3 jspl3_w_n4494_17(.douta(w_n4494_17[0]),.doutb(w_n4494_17[1]),.doutc(w_n4494_17[2]),.din(w_n4494_5[1]));
	jspl3 jspl3_w_n4494_18(.douta(w_n4494_18[0]),.doutb(w_n4494_18[1]),.doutc(w_n4494_18[2]),.din(w_n4494_5[2]));
	jspl3 jspl3_w_n4494_19(.douta(w_n4494_19[0]),.doutb(w_n4494_19[1]),.doutc(w_n4494_19[2]),.din(w_n4494_6[0]));
	jspl3 jspl3_w_n4494_20(.douta(w_n4494_20[0]),.doutb(w_n4494_20[1]),.doutc(w_n4494_20[2]),.din(w_n4494_6[1]));
	jspl3 jspl3_w_n4494_21(.douta(w_n4494_21[0]),.doutb(w_n4494_21[1]),.doutc(w_n4494_21[2]),.din(w_n4494_6[2]));
	jspl3 jspl3_w_n4494_22(.douta(w_n4494_22[0]),.doutb(w_n4494_22[1]),.doutc(w_n4494_22[2]),.din(w_n4494_7[0]));
	jspl jspl_w_n4494_23(.douta(w_n4494_23[0]),.doutb(w_n4494_23[1]),.din(w_n4494_7[1]));
	jspl3 jspl3_w_n4499_0(.douta(w_n4499_0[0]),.doutb(w_n4499_0[1]),.doutc(w_n4499_0[2]),.din(n4499));
	jspl3 jspl3_w_n4499_1(.douta(w_n4499_1[0]),.doutb(w_n4499_1[1]),.doutc(w_n4499_1[2]),.din(w_n4499_0[0]));
	jspl3 jspl3_w_n4499_2(.douta(w_n4499_2[0]),.doutb(w_n4499_2[1]),.doutc(w_n4499_2[2]),.din(w_n4499_0[1]));
	jspl3 jspl3_w_n4499_3(.douta(w_n4499_3[0]),.doutb(w_n4499_3[1]),.doutc(w_n4499_3[2]),.din(w_n4499_0[2]));
	jspl3 jspl3_w_n4499_4(.douta(w_n4499_4[0]),.doutb(w_n4499_4[1]),.doutc(w_n4499_4[2]),.din(w_n4499_1[0]));
	jspl3 jspl3_w_n4499_5(.douta(w_n4499_5[0]),.doutb(w_n4499_5[1]),.doutc(w_n4499_5[2]),.din(w_n4499_1[1]));
	jspl3 jspl3_w_n4499_6(.douta(w_n4499_6[0]),.doutb(w_n4499_6[1]),.doutc(w_n4499_6[2]),.din(w_n4499_1[2]));
	jspl3 jspl3_w_n4499_7(.douta(w_n4499_7[0]),.doutb(w_n4499_7[1]),.doutc(w_n4499_7[2]),.din(w_n4499_2[0]));
	jspl3 jspl3_w_n4499_8(.douta(w_n4499_8[0]),.doutb(w_n4499_8[1]),.doutc(w_n4499_8[2]),.din(w_n4499_2[1]));
	jspl3 jspl3_w_n4499_9(.douta(w_n4499_9[0]),.doutb(w_n4499_9[1]),.doutc(w_n4499_9[2]),.din(w_n4499_2[2]));
	jspl3 jspl3_w_n4499_10(.douta(w_n4499_10[0]),.doutb(w_n4499_10[1]),.doutc(w_n4499_10[2]),.din(w_n4499_3[0]));
	jspl3 jspl3_w_n4499_11(.douta(w_n4499_11[0]),.doutb(w_n4499_11[1]),.doutc(w_n4499_11[2]),.din(w_n4499_3[1]));
	jspl3 jspl3_w_n4499_12(.douta(w_n4499_12[0]),.doutb(w_n4499_12[1]),.doutc(w_n4499_12[2]),.din(w_n4499_3[2]));
	jspl3 jspl3_w_n4499_13(.douta(w_n4499_13[0]),.doutb(w_n4499_13[1]),.doutc(w_n4499_13[2]),.din(w_n4499_4[0]));
	jspl3 jspl3_w_n4499_14(.douta(w_n4499_14[0]),.doutb(w_n4499_14[1]),.doutc(w_n4499_14[2]),.din(w_n4499_4[1]));
	jspl3 jspl3_w_n4499_15(.douta(w_n4499_15[0]),.doutb(w_n4499_15[1]),.doutc(w_n4499_15[2]),.din(w_n4499_4[2]));
	jspl3 jspl3_w_n4499_16(.douta(w_n4499_16[0]),.doutb(w_n4499_16[1]),.doutc(w_n4499_16[2]),.din(w_n4499_5[0]));
	jspl3 jspl3_w_n4499_17(.douta(w_n4499_17[0]),.doutb(w_n4499_17[1]),.doutc(w_n4499_17[2]),.din(w_n4499_5[1]));
	jspl3 jspl3_w_n4499_18(.douta(w_n4499_18[0]),.doutb(w_n4499_18[1]),.doutc(w_n4499_18[2]),.din(w_n4499_5[2]));
	jspl3 jspl3_w_n4499_19(.douta(w_n4499_19[0]),.doutb(w_n4499_19[1]),.doutc(w_n4499_19[2]),.din(w_n4499_6[0]));
	jspl3 jspl3_w_n4499_20(.douta(w_n4499_20[0]),.doutb(w_n4499_20[1]),.doutc(w_n4499_20[2]),.din(w_n4499_6[1]));
	jspl3 jspl3_w_n4499_21(.douta(w_n4499_21[0]),.doutb(w_n4499_21[1]),.doutc(w_n4499_21[2]),.din(w_n4499_6[2]));
	jspl3 jspl3_w_n4499_22(.douta(w_n4499_22[0]),.doutb(w_n4499_22[1]),.doutc(w_n4499_22[2]),.din(w_n4499_7[0]));
	jspl3 jspl3_w_n4499_23(.douta(w_n4499_23[0]),.doutb(w_n4499_23[1]),.doutc(w_n4499_23[2]),.din(w_n4499_7[1]));
	jspl3 jspl3_w_n4499_24(.douta(w_n4499_24[0]),.doutb(w_n4499_24[1]),.doutc(w_n4499_24[2]),.din(w_n4499_7[2]));
	jspl3 jspl3_w_n4499_25(.douta(w_n4499_25[0]),.doutb(w_n4499_25[1]),.doutc(w_n4499_25[2]),.din(w_n4499_8[0]));
	jspl3 jspl3_w_n4499_26(.douta(w_n4499_26[0]),.doutb(w_n4499_26[1]),.doutc(w_n4499_26[2]),.din(w_n4499_8[1]));
	jspl3 jspl3_w_n4499_27(.douta(w_n4499_27[0]),.doutb(w_n4499_27[1]),.doutc(w_n4499_27[2]),.din(w_n4499_8[2]));
	jspl3 jspl3_w_n4499_28(.douta(w_n4499_28[0]),.doutb(w_n4499_28[1]),.doutc(w_n4499_28[2]),.din(w_n4499_9[0]));
	jspl3 jspl3_w_n4499_29(.douta(w_n4499_29[0]),.doutb(w_n4499_29[1]),.doutc(w_n4499_29[2]),.din(w_n4499_9[1]));
	jspl3 jspl3_w_n4499_30(.douta(w_n4499_30[0]),.doutb(w_n4499_30[1]),.doutc(w_n4499_30[2]),.din(w_n4499_9[2]));
	jspl jspl_w_n4499_31(.douta(w_n4499_31[0]),.doutb(w_n4499_31[1]),.din(w_n4499_10[0]));
	jspl3 jspl3_w_n4502_0(.douta(w_n4502_0[0]),.doutb(w_n4502_0[1]),.doutc(w_n4502_0[2]),.din(n4502));
	jspl jspl_w_n4502_1(.douta(w_n4502_1[0]),.doutb(w_n4502_1[1]),.din(w_n4502_0[0]));
	jspl3 jspl3_w_n4503_0(.douta(w_n4503_0[0]),.doutb(w_n4503_0[1]),.doutc(w_n4503_0[2]),.din(n4503));
	jspl3 jspl3_w_n4507_0(.douta(w_n4507_0[0]),.doutb(w_n4507_0[1]),.doutc(w_n4507_0[2]),.din(n4507));
	jspl jspl_w_n4508_0(.douta(w_n4508_0[0]),.doutb(w_n4508_0[1]),.din(n4508));
	jspl jspl_w_n4509_0(.douta(w_n4509_0[0]),.doutb(w_n4509_0[1]),.din(n4509));
	jspl jspl_w_n4510_0(.douta(w_n4510_0[0]),.doutb(w_n4510_0[1]),.din(n4510));
	jspl jspl_w_n4512_0(.douta(w_n4512_0[0]),.doutb(w_n4512_0[1]),.din(n4512));
	jspl jspl_w_n4514_0(.douta(w_n4514_0[0]),.doutb(w_n4514_0[1]),.din(n4514));
	jspl jspl_w_n4516_0(.douta(w_n4516_0[0]),.doutb(w_n4516_0[1]),.din(n4516));
	jspl jspl_w_n4519_0(.douta(w_n4519_0[0]),.doutb(w_n4519_0[1]),.din(n4519));
	jspl jspl_w_n4524_0(.douta(w_n4524_0[0]),.doutb(w_n4524_0[1]),.din(n4524));
	jspl3 jspl3_w_n4526_0(.douta(w_n4526_0[0]),.doutb(w_n4526_0[1]),.doutc(w_n4526_0[2]),.din(n4526));
	jspl jspl_w_n4527_0(.douta(w_n4527_0[0]),.doutb(w_n4527_0[1]),.din(n4527));
	jspl jspl_w_n4531_0(.douta(w_n4531_0[0]),.doutb(w_n4531_0[1]),.din(n4531));
	jspl jspl_w_n4532_0(.douta(w_n4532_0[0]),.doutb(w_n4532_0[1]),.din(n4532));
	jspl jspl_w_n4534_0(.douta(w_n4534_0[0]),.doutb(w_n4534_0[1]),.din(n4534));
	jspl jspl_w_n4538_0(.douta(w_n4538_0[0]),.doutb(w_n4538_0[1]),.din(n4538));
	jspl jspl_w_n4540_0(.douta(w_n4540_0[0]),.doutb(w_n4540_0[1]),.din(n4540));
	jspl jspl_w_n4541_0(.douta(w_n4541_0[0]),.doutb(w_n4541_0[1]),.din(n4541));
	jspl3 jspl3_w_n4542_0(.douta(w_n4542_0[0]),.doutb(w_n4542_0[1]),.doutc(w_n4542_0[2]),.din(n4542));
	jspl jspl_w_n4543_0(.douta(w_n4543_0[0]),.doutb(w_n4543_0[1]),.din(n4543));
	jspl jspl_w_n4547_0(.douta(w_n4547_0[0]),.doutb(w_n4547_0[1]),.din(n4547));
	jspl jspl_w_n4549_0(.douta(w_n4549_0[0]),.doutb(w_n4549_0[1]),.din(n4549));
	jspl jspl_w_n4551_0(.douta(w_n4551_0[0]),.doutb(w_n4551_0[1]),.din(n4551));
	jspl jspl_w_n4553_0(.douta(w_n4553_0[0]),.doutb(w_n4553_0[1]),.din(n4553));
	jspl jspl_w_n4555_0(.douta(w_n4555_0[0]),.doutb(w_n4555_0[1]),.din(n4555));
	jspl jspl_w_n4561_0(.douta(w_n4561_0[0]),.doutb(w_n4561_0[1]),.din(n4561));
	jspl3 jspl3_w_n4563_0(.douta(w_n4563_0[0]),.doutb(w_n4563_0[1]),.doutc(w_n4563_0[2]),.din(n4563));
	jspl jspl_w_n4564_0(.douta(w_n4564_0[0]),.doutb(w_n4564_0[1]),.din(n4564));
	jspl jspl_w_n4569_0(.douta(w_n4569_0[0]),.doutb(w_n4569_0[1]),.din(n4569));
	jspl jspl_w_n4571_0(.douta(w_n4571_0[0]),.doutb(w_n4571_0[1]),.din(n4571));
	jspl jspl_w_n4573_0(.douta(w_n4573_0[0]),.doutb(w_n4573_0[1]),.din(n4573));
	jspl jspl_w_n4577_0(.douta(w_n4577_0[0]),.doutb(w_n4577_0[1]),.din(n4577));
	jspl jspl_w_n4579_0(.douta(w_n4579_0[0]),.doutb(w_n4579_0[1]),.din(n4579));
	jspl jspl_w_n4580_0(.douta(w_n4580_0[0]),.doutb(w_n4580_0[1]),.din(n4580));
	jspl3 jspl3_w_n4581_0(.douta(w_n4581_0[0]),.doutb(w_n4581_0[1]),.doutc(w_n4581_0[2]),.din(n4581));
	jspl jspl_w_n4582_0(.douta(w_n4582_0[0]),.doutb(w_n4582_0[1]),.din(n4582));
	jspl jspl_w_n4588_0(.douta(w_n4588_0[0]),.doutb(w_n4588_0[1]),.din(n4588));
	jspl jspl_w_n4589_0(.douta(w_n4589_0[0]),.doutb(w_n4589_0[1]),.din(n4589));
	jspl jspl_w_n4591_0(.douta(w_n4591_0[0]),.doutb(w_n4591_0[1]),.din(n4591));
	jspl jspl_w_n4593_0(.douta(w_n4593_0[0]),.doutb(w_n4593_0[1]),.din(n4593));
	jspl jspl_w_n4595_0(.douta(w_n4595_0[0]),.doutb(w_n4595_0[1]),.din(n4595));
	jspl jspl_w_n4601_0(.douta(w_n4601_0[0]),.doutb(w_n4601_0[1]),.din(n4601));
	jspl jspl_w_n4603_0(.douta(w_n4603_0[0]),.doutb(w_n4603_0[1]),.din(n4603));
	jspl3 jspl3_w_n4604_0(.douta(w_n4604_0[0]),.doutb(w_n4604_0[1]),.doutc(w_n4604_0[2]),.din(n4604));
	jspl jspl_w_n4607_0(.douta(w_n4607_0[0]),.doutb(w_n4607_0[1]),.din(n4607));
	jspl jspl_w_n4608_0(.douta(w_n4608_0[0]),.doutb(w_n4608_0[1]),.din(n4608));
	jspl3 jspl3_w_n4609_0(.douta(w_n4609_0[0]),.doutb(w_n4609_0[1]),.doutc(w_n4609_0[2]),.din(n4609));
	jspl jspl_w_n4611_0(.douta(w_n4611_0[0]),.doutb(w_n4611_0[1]),.din(n4611));
	jspl jspl_w_n4615_0(.douta(w_n4615_0[0]),.doutb(w_n4615_0[1]),.din(n4615));
	jspl jspl_w_n4617_0(.douta(w_n4617_0[0]),.doutb(w_n4617_0[1]),.din(n4617));
	jspl jspl_w_n4618_0(.douta(w_n4618_0[0]),.doutb(w_n4618_0[1]),.din(n4618));
	jspl3 jspl3_w_n4619_0(.douta(w_n4619_0[0]),.doutb(w_n4619_0[1]),.doutc(w_n4619_0[2]),.din(n4619));
	jspl jspl_w_n4620_0(.douta(w_n4620_0[0]),.doutb(w_n4620_0[1]),.din(n4620));
	jspl jspl_w_n4623_0(.douta(w_n4623_0[0]),.doutb(w_n4623_0[1]),.din(n4623));
	jspl jspl_w_n4629_0(.douta(w_n4629_0[0]),.doutb(w_n4629_0[1]),.din(n4629));
	jspl jspl_w_n4630_0(.douta(w_n4630_0[0]),.doutb(w_n4630_0[1]),.din(n4630));
	jspl jspl_w_n4632_0(.douta(w_n4632_0[0]),.doutb(w_n4632_0[1]),.din(n4632));
	jspl jspl_w_n4634_0(.douta(w_n4634_0[0]),.doutb(w_n4634_0[1]),.din(n4634));
	jspl jspl_w_n4636_0(.douta(w_n4636_0[0]),.doutb(w_n4636_0[1]),.din(n4636));
	jspl jspl_w_n4642_0(.douta(w_n4642_0[0]),.doutb(w_n4642_0[1]),.din(n4642));
	jspl jspl_w_n4644_0(.douta(w_n4644_0[0]),.doutb(w_n4644_0[1]),.din(n4644));
	jspl3 jspl3_w_n4645_0(.douta(w_n4645_0[0]),.doutb(w_n4645_0[1]),.doutc(w_n4645_0[2]),.din(n4645));
	jspl jspl_w_n4648_0(.douta(w_n4648_0[0]),.doutb(w_n4648_0[1]),.din(n4648));
	jspl jspl_w_n4649_0(.douta(w_n4649_0[0]),.doutb(w_n4649_0[1]),.din(n4649));
	jspl3 jspl3_w_n4650_0(.douta(w_n4650_0[0]),.doutb(w_n4650_0[1]),.doutc(w_n4650_0[2]),.din(n4650));
	jspl jspl_w_n4652_0(.douta(w_n4652_0[0]),.doutb(w_n4652_0[1]),.din(n4652));
	jspl jspl_w_n4656_0(.douta(w_n4656_0[0]),.doutb(w_n4656_0[1]),.din(n4656));
	jspl jspl_w_n4658_0(.douta(w_n4658_0[0]),.doutb(w_n4658_0[1]),.din(n4658));
	jspl jspl_w_n4659_0(.douta(w_n4659_0[0]),.doutb(w_n4659_0[1]),.din(n4659));
	jspl3 jspl3_w_n4660_0(.douta(w_n4660_0[0]),.doutb(w_n4660_0[1]),.doutc(w_n4660_0[2]),.din(n4660));
	jspl jspl_w_n4661_0(.douta(w_n4661_0[0]),.doutb(w_n4661_0[1]),.din(n4661));
	jspl jspl_w_n4664_0(.douta(w_n4664_0[0]),.doutb(w_n4664_0[1]),.din(n4664));
	jspl jspl_w_n4670_0(.douta(w_n4670_0[0]),.doutb(w_n4670_0[1]),.din(n4670));
	jspl jspl_w_n4671_0(.douta(w_n4671_0[0]),.doutb(w_n4671_0[1]),.din(n4671));
	jspl jspl_w_n4673_0(.douta(w_n4673_0[0]),.doutb(w_n4673_0[1]),.din(n4673));
	jspl jspl_w_n4675_0(.douta(w_n4675_0[0]),.doutb(w_n4675_0[1]),.din(n4675));
	jspl jspl_w_n4677_0(.douta(w_n4677_0[0]),.doutb(w_n4677_0[1]),.din(n4677));
	jspl jspl_w_n4683_0(.douta(w_n4683_0[0]),.doutb(w_n4683_0[1]),.din(n4683));
	jspl jspl_w_n4685_0(.douta(w_n4685_0[0]),.doutb(w_n4685_0[1]),.din(n4685));
	jspl3 jspl3_w_n4686_0(.douta(w_n4686_0[0]),.doutb(w_n4686_0[1]),.doutc(w_n4686_0[2]),.din(n4686));
	jspl jspl_w_n4689_0(.douta(w_n4689_0[0]),.doutb(w_n4689_0[1]),.din(n4689));
	jspl jspl_w_n4690_0(.douta(w_n4690_0[0]),.doutb(w_n4690_0[1]),.din(n4690));
	jspl3 jspl3_w_n4691_0(.douta(w_n4691_0[0]),.doutb(w_n4691_0[1]),.doutc(w_n4691_0[2]),.din(n4691));
	jspl jspl_w_n4693_0(.douta(w_n4693_0[0]),.doutb(w_n4693_0[1]),.din(n4693));
	jspl jspl_w_n4697_0(.douta(w_n4697_0[0]),.doutb(w_n4697_0[1]),.din(n4697));
	jspl jspl_w_n4699_0(.douta(w_n4699_0[0]),.doutb(w_n4699_0[1]),.din(n4699));
	jspl jspl_w_n4700_0(.douta(w_n4700_0[0]),.doutb(w_n4700_0[1]),.din(n4700));
	jspl3 jspl3_w_n4701_0(.douta(w_n4701_0[0]),.doutb(w_n4701_0[1]),.doutc(w_n4701_0[2]),.din(n4701));
	jspl jspl_w_n4702_0(.douta(w_n4702_0[0]),.doutb(w_n4702_0[1]),.din(n4702));
	jspl jspl_w_n4705_0(.douta(w_n4705_0[0]),.doutb(w_n4705_0[1]),.din(n4705));
	jspl jspl_w_n4711_0(.douta(w_n4711_0[0]),.doutb(w_n4711_0[1]),.din(n4711));
	jspl jspl_w_n4712_0(.douta(w_n4712_0[0]),.doutb(w_n4712_0[1]),.din(n4712));
	jspl jspl_w_n4714_0(.douta(w_n4714_0[0]),.doutb(w_n4714_0[1]),.din(n4714));
	jspl jspl_w_n4716_0(.douta(w_n4716_0[0]),.doutb(w_n4716_0[1]),.din(n4716));
	jspl jspl_w_n4718_0(.douta(w_n4718_0[0]),.doutb(w_n4718_0[1]),.din(n4718));
	jspl jspl_w_n4724_0(.douta(w_n4724_0[0]),.doutb(w_n4724_0[1]),.din(n4724));
	jspl jspl_w_n4726_0(.douta(w_n4726_0[0]),.doutb(w_n4726_0[1]),.din(n4726));
	jspl3 jspl3_w_n4727_0(.douta(w_n4727_0[0]),.doutb(w_n4727_0[1]),.doutc(w_n4727_0[2]),.din(n4727));
	jspl jspl_w_n4730_0(.douta(w_n4730_0[0]),.doutb(w_n4730_0[1]),.din(n4730));
	jspl jspl_w_n4731_0(.douta(w_n4731_0[0]),.doutb(w_n4731_0[1]),.din(n4731));
	jspl3 jspl3_w_n4732_0(.douta(w_n4732_0[0]),.doutb(w_n4732_0[1]),.doutc(w_n4732_0[2]),.din(n4732));
	jspl jspl_w_n4734_0(.douta(w_n4734_0[0]),.doutb(w_n4734_0[1]),.din(n4734));
	jspl jspl_w_n4738_0(.douta(w_n4738_0[0]),.doutb(w_n4738_0[1]),.din(n4738));
	jspl jspl_w_n4740_0(.douta(w_n4740_0[0]),.doutb(w_n4740_0[1]),.din(n4740));
	jspl jspl_w_n4741_0(.douta(w_n4741_0[0]),.doutb(w_n4741_0[1]),.din(n4741));
	jspl3 jspl3_w_n4742_0(.douta(w_n4742_0[0]),.doutb(w_n4742_0[1]),.doutc(w_n4742_0[2]),.din(n4742));
	jspl jspl_w_n4743_0(.douta(w_n4743_0[0]),.doutb(w_n4743_0[1]),.din(n4743));
	jspl jspl_w_n4746_0(.douta(w_n4746_0[0]),.doutb(w_n4746_0[1]),.din(n4746));
	jspl jspl_w_n4752_0(.douta(w_n4752_0[0]),.doutb(w_n4752_0[1]),.din(n4752));
	jspl jspl_w_n4753_0(.douta(w_n4753_0[0]),.doutb(w_n4753_0[1]),.din(n4753));
	jspl jspl_w_n4755_0(.douta(w_n4755_0[0]),.doutb(w_n4755_0[1]),.din(n4755));
	jspl jspl_w_n4757_0(.douta(w_n4757_0[0]),.doutb(w_n4757_0[1]),.din(n4757));
	jspl jspl_w_n4759_0(.douta(w_n4759_0[0]),.doutb(w_n4759_0[1]),.din(n4759));
	jspl jspl_w_n4765_0(.douta(w_n4765_0[0]),.doutb(w_n4765_0[1]),.din(n4765));
	jspl3 jspl3_w_n4767_0(.douta(w_n4767_0[0]),.doutb(w_n4767_0[1]),.doutc(w_n4767_0[2]),.din(n4767));
	jspl jspl_w_n4772_0(.douta(w_n4772_0[0]),.doutb(w_n4772_0[1]),.din(n4772));
	jspl3 jspl3_w_n4774_0(.douta(w_n4774_0[0]),.doutb(w_n4774_0[1]),.doutc(w_n4774_0[2]),.din(n4774));
	jspl3 jspl3_w_n4778_0(.douta(w_n4778_0[0]),.doutb(w_n4778_0[1]),.doutc(w_n4778_0[2]),.din(n4778));
	jspl jspl_w_n4779_0(.douta(w_n4779_0[0]),.doutb(w_n4779_0[1]),.din(n4779));
	jspl jspl_w_n4784_0(.douta(w_n4784_0[0]),.doutb(w_n4784_0[1]),.din(n4784));
	jspl3 jspl3_w_n4785_0(.douta(w_n4785_0[0]),.doutb(w_n4785_0[1]),.doutc(w_n4785_0[2]),.din(n4785));
	jspl jspl_w_n4790_0(.douta(w_n4790_0[0]),.doutb(w_n4790_0[1]),.din(n4790));
	jspl3 jspl3_w_n4796_0(.douta(w_n4796_0[0]),.doutb(w_n4796_0[1]),.doutc(w_n4796_0[2]),.din(n4796));
	jspl jspl_w_n4796_1(.douta(w_n4796_1[0]),.doutb(w_n4796_1[1]),.din(w_n4796_0[0]));
	jspl jspl_w_n4797_0(.douta(w_n4797_0[0]),.doutb(w_n4797_0[1]),.din(n4797));
	jspl3 jspl3_w_n4800_0(.douta(w_n4800_0[0]),.doutb(w_n4800_0[1]),.doutc(w_n4800_0[2]),.din(n4800));
	jspl jspl_w_n4801_0(.douta(w_n4801_0[0]),.doutb(w_n4801_0[1]),.din(n4801));
	jspl jspl_w_n4802_0(.douta(w_n4802_0[0]),.doutb(w_n4802_0[1]),.din(n4802));
	jspl jspl_w_n4803_0(.douta(w_n4803_0[0]),.doutb(w_n4803_0[1]),.din(n4803));
	jspl jspl_w_n4805_0(.douta(w_n4805_0[0]),.doutb(w_n4805_0[1]),.din(n4805));
	jspl jspl_w_n4807_0(.douta(w_n4807_0[0]),.doutb(w_n4807_0[1]),.din(n4807));
	jspl jspl_w_n4809_0(.douta(w_n4809_0[0]),.doutb(w_n4809_0[1]),.din(n4809));
	jspl jspl_w_n4818_0(.douta(w_n4818_0[0]),.doutb(w_n4818_0[1]),.din(n4818));
	jspl3 jspl3_w_n4820_0(.douta(w_n4820_0[0]),.doutb(w_n4820_0[1]),.doutc(w_n4820_0[2]),.din(n4820));
	jspl jspl_w_n4821_0(.douta(w_n4821_0[0]),.doutb(w_n4821_0[1]),.din(n4821));
	jspl jspl_w_n4825_0(.douta(w_n4825_0[0]),.doutb(w_n4825_0[1]),.din(n4825));
	jspl jspl_w_n4827_0(.douta(w_n4827_0[0]),.doutb(w_n4827_0[1]),.din(n4827));
	jspl jspl_w_n4829_0(.douta(w_n4829_0[0]),.doutb(w_n4829_0[1]),.din(n4829));
	jspl jspl_w_n4834_0(.douta(w_n4834_0[0]),.doutb(w_n4834_0[1]),.din(n4834));
	jspl jspl_w_n4836_0(.douta(w_n4836_0[0]),.doutb(w_n4836_0[1]),.din(n4836));
	jspl jspl_w_n4837_0(.douta(w_n4837_0[0]),.doutb(w_n4837_0[1]),.din(n4837));
	jspl3 jspl3_w_n4838_0(.douta(w_n4838_0[0]),.doutb(w_n4838_0[1]),.doutc(w_n4838_0[2]),.din(n4838));
	jspl jspl_w_n4839_0(.douta(w_n4839_0[0]),.doutb(w_n4839_0[1]),.din(n4839));
	jspl jspl_w_n4844_0(.douta(w_n4844_0[0]),.doutb(w_n4844_0[1]),.din(n4844));
	jspl jspl_w_n4845_0(.douta(w_n4845_0[0]),.doutb(w_n4845_0[1]),.din(n4845));
	jspl jspl_w_n4847_0(.douta(w_n4847_0[0]),.doutb(w_n4847_0[1]),.din(n4847));
	jspl jspl_w_n4849_0(.douta(w_n4849_0[0]),.doutb(w_n4849_0[1]),.din(n4849));
	jspl jspl_w_n4852_0(.douta(w_n4852_0[0]),.doutb(w_n4852_0[1]),.din(n4852));
	jspl jspl_w_n4858_0(.douta(w_n4858_0[0]),.doutb(w_n4858_0[1]),.din(n4858));
	jspl3 jspl3_w_n4860_0(.douta(w_n4860_0[0]),.doutb(w_n4860_0[1]),.doutc(w_n4860_0[2]),.din(n4860));
	jspl jspl_w_n4861_0(.douta(w_n4861_0[0]),.doutb(w_n4861_0[1]),.din(n4861));
	jspl jspl_w_n4865_0(.douta(w_n4865_0[0]),.doutb(w_n4865_0[1]),.din(n4865));
	jspl jspl_w_n4866_0(.douta(w_n4866_0[0]),.doutb(w_n4866_0[1]),.din(n4866));
	jspl jspl_w_n4868_0(.douta(w_n4868_0[0]),.doutb(w_n4868_0[1]),.din(n4868));
	jspl jspl_w_n4873_0(.douta(w_n4873_0[0]),.doutb(w_n4873_0[1]),.din(n4873));
	jspl jspl_w_n4875_0(.douta(w_n4875_0[0]),.doutb(w_n4875_0[1]),.din(n4875));
	jspl jspl_w_n4876_0(.douta(w_n4876_0[0]),.doutb(w_n4876_0[1]),.din(n4876));
	jspl3 jspl3_w_n4877_0(.douta(w_n4877_0[0]),.doutb(w_n4877_0[1]),.doutc(w_n4877_0[2]),.din(n4877));
	jspl jspl_w_n4878_0(.douta(w_n4878_0[0]),.doutb(w_n4878_0[1]),.din(n4878));
	jspl jspl_w_n4882_0(.douta(w_n4882_0[0]),.doutb(w_n4882_0[1]),.din(n4882));
	jspl jspl_w_n4883_0(.douta(w_n4883_0[0]),.doutb(w_n4883_0[1]),.din(n4883));
	jspl jspl_w_n4885_0(.douta(w_n4885_0[0]),.doutb(w_n4885_0[1]),.din(n4885));
	jspl jspl_w_n4887_0(.douta(w_n4887_0[0]),.doutb(w_n4887_0[1]),.din(n4887));
	jspl jspl_w_n4890_0(.douta(w_n4890_0[0]),.doutb(w_n4890_0[1]),.din(n4890));
	jspl jspl_w_n4896_0(.douta(w_n4896_0[0]),.doutb(w_n4896_0[1]),.din(n4896));
	jspl jspl_w_n4898_0(.douta(w_n4898_0[0]),.doutb(w_n4898_0[1]),.din(n4898));
	jspl3 jspl3_w_n4899_0(.douta(w_n4899_0[0]),.doutb(w_n4899_0[1]),.doutc(w_n4899_0[2]),.din(n4899));
	jspl jspl_w_n4903_0(.douta(w_n4903_0[0]),.doutb(w_n4903_0[1]),.din(n4903));
	jspl jspl_w_n4904_0(.douta(w_n4904_0[0]),.doutb(w_n4904_0[1]),.din(n4904));
	jspl3 jspl3_w_n4905_0(.douta(w_n4905_0[0]),.doutb(w_n4905_0[1]),.doutc(w_n4905_0[2]),.din(n4905));
	jspl jspl_w_n4907_0(.douta(w_n4907_0[0]),.doutb(w_n4907_0[1]),.din(n4907));
	jspl jspl_w_n4912_0(.douta(w_n4912_0[0]),.doutb(w_n4912_0[1]),.din(n4912));
	jspl jspl_w_n4914_0(.douta(w_n4914_0[0]),.doutb(w_n4914_0[1]),.din(n4914));
	jspl jspl_w_n4915_0(.douta(w_n4915_0[0]),.doutb(w_n4915_0[1]),.din(n4915));
	jspl3 jspl3_w_n4916_0(.douta(w_n4916_0[0]),.doutb(w_n4916_0[1]),.doutc(w_n4916_0[2]),.din(n4916));
	jspl jspl_w_n4917_0(.douta(w_n4917_0[0]),.doutb(w_n4917_0[1]),.din(n4917));
	jspl jspl_w_n4921_0(.douta(w_n4921_0[0]),.doutb(w_n4921_0[1]),.din(n4921));
	jspl jspl_w_n4927_0(.douta(w_n4927_0[0]),.doutb(w_n4927_0[1]),.din(n4927));
	jspl jspl_w_n4928_0(.douta(w_n4928_0[0]),.doutb(w_n4928_0[1]),.din(n4928));
	jspl jspl_w_n4930_0(.douta(w_n4930_0[0]),.doutb(w_n4930_0[1]),.din(n4930));
	jspl jspl_w_n4932_0(.douta(w_n4932_0[0]),.doutb(w_n4932_0[1]),.din(n4932));
	jspl jspl_w_n4935_0(.douta(w_n4935_0[0]),.doutb(w_n4935_0[1]),.din(n4935));
	jspl jspl_w_n4941_0(.douta(w_n4941_0[0]),.doutb(w_n4941_0[1]),.din(n4941));
	jspl jspl_w_n4943_0(.douta(w_n4943_0[0]),.doutb(w_n4943_0[1]),.din(n4943));
	jspl3 jspl3_w_n4944_0(.douta(w_n4944_0[0]),.doutb(w_n4944_0[1]),.doutc(w_n4944_0[2]),.din(n4944));
	jspl jspl_w_n4948_0(.douta(w_n4948_0[0]),.doutb(w_n4948_0[1]),.din(n4948));
	jspl jspl_w_n4949_0(.douta(w_n4949_0[0]),.doutb(w_n4949_0[1]),.din(n4949));
	jspl3 jspl3_w_n4950_0(.douta(w_n4950_0[0]),.doutb(w_n4950_0[1]),.doutc(w_n4950_0[2]),.din(n4950));
	jspl jspl_w_n4952_0(.douta(w_n4952_0[0]),.doutb(w_n4952_0[1]),.din(n4952));
	jspl jspl_w_n4957_0(.douta(w_n4957_0[0]),.doutb(w_n4957_0[1]),.din(n4957));
	jspl jspl_w_n4959_0(.douta(w_n4959_0[0]),.doutb(w_n4959_0[1]),.din(n4959));
	jspl jspl_w_n4960_0(.douta(w_n4960_0[0]),.doutb(w_n4960_0[1]),.din(n4960));
	jspl3 jspl3_w_n4961_0(.douta(w_n4961_0[0]),.doutb(w_n4961_0[1]),.doutc(w_n4961_0[2]),.din(n4961));
	jspl jspl_w_n4962_0(.douta(w_n4962_0[0]),.doutb(w_n4962_0[1]),.din(n4962));
	jspl jspl_w_n4966_0(.douta(w_n4966_0[0]),.doutb(w_n4966_0[1]),.din(n4966));
	jspl jspl_w_n4972_0(.douta(w_n4972_0[0]),.doutb(w_n4972_0[1]),.din(n4972));
	jspl jspl_w_n4973_0(.douta(w_n4973_0[0]),.doutb(w_n4973_0[1]),.din(n4973));
	jspl jspl_w_n4975_0(.douta(w_n4975_0[0]),.doutb(w_n4975_0[1]),.din(n4975));
	jspl jspl_w_n4977_0(.douta(w_n4977_0[0]),.doutb(w_n4977_0[1]),.din(n4977));
	jspl jspl_w_n4980_0(.douta(w_n4980_0[0]),.doutb(w_n4980_0[1]),.din(n4980));
	jspl jspl_w_n4986_0(.douta(w_n4986_0[0]),.doutb(w_n4986_0[1]),.din(n4986));
	jspl jspl_w_n4988_0(.douta(w_n4988_0[0]),.doutb(w_n4988_0[1]),.din(n4988));
	jspl3 jspl3_w_n4989_0(.douta(w_n4989_0[0]),.doutb(w_n4989_0[1]),.doutc(w_n4989_0[2]),.din(n4989));
	jspl jspl_w_n4993_0(.douta(w_n4993_0[0]),.doutb(w_n4993_0[1]),.din(n4993));
	jspl jspl_w_n4994_0(.douta(w_n4994_0[0]),.doutb(w_n4994_0[1]),.din(n4994));
	jspl3 jspl3_w_n4995_0(.douta(w_n4995_0[0]),.doutb(w_n4995_0[1]),.doutc(w_n4995_0[2]),.din(n4995));
	jspl jspl_w_n4997_0(.douta(w_n4997_0[0]),.doutb(w_n4997_0[1]),.din(n4997));
	jspl jspl_w_n5002_0(.douta(w_n5002_0[0]),.doutb(w_n5002_0[1]),.din(n5002));
	jspl jspl_w_n5004_0(.douta(w_n5004_0[0]),.doutb(w_n5004_0[1]),.din(n5004));
	jspl jspl_w_n5005_0(.douta(w_n5005_0[0]),.doutb(w_n5005_0[1]),.din(n5005));
	jspl3 jspl3_w_n5006_0(.douta(w_n5006_0[0]),.doutb(w_n5006_0[1]),.doutc(w_n5006_0[2]),.din(n5006));
	jspl jspl_w_n5007_0(.douta(w_n5007_0[0]),.doutb(w_n5007_0[1]),.din(n5007));
	jspl jspl_w_n5011_0(.douta(w_n5011_0[0]),.doutb(w_n5011_0[1]),.din(n5011));
	jspl jspl_w_n5017_0(.douta(w_n5017_0[0]),.doutb(w_n5017_0[1]),.din(n5017));
	jspl jspl_w_n5018_0(.douta(w_n5018_0[0]),.doutb(w_n5018_0[1]),.din(n5018));
	jspl jspl_w_n5020_0(.douta(w_n5020_0[0]),.doutb(w_n5020_0[1]),.din(n5020));
	jspl jspl_w_n5022_0(.douta(w_n5022_0[0]),.doutb(w_n5022_0[1]),.din(n5022));
	jspl jspl_w_n5025_0(.douta(w_n5025_0[0]),.doutb(w_n5025_0[1]),.din(n5025));
	jspl jspl_w_n5031_0(.douta(w_n5031_0[0]),.doutb(w_n5031_0[1]),.din(n5031));
	jspl jspl_w_n5033_0(.douta(w_n5033_0[0]),.doutb(w_n5033_0[1]),.din(n5033));
	jspl3 jspl3_w_n5034_0(.douta(w_n5034_0[0]),.doutb(w_n5034_0[1]),.doutc(w_n5034_0[2]),.din(n5034));
	jspl jspl_w_n5038_0(.douta(w_n5038_0[0]),.doutb(w_n5038_0[1]),.din(n5038));
	jspl jspl_w_n5039_0(.douta(w_n5039_0[0]),.doutb(w_n5039_0[1]),.din(n5039));
	jspl3 jspl3_w_n5040_0(.douta(w_n5040_0[0]),.doutb(w_n5040_0[1]),.doutc(w_n5040_0[2]),.din(n5040));
	jspl jspl_w_n5042_0(.douta(w_n5042_0[0]),.doutb(w_n5042_0[1]),.din(n5042));
	jspl jspl_w_n5047_0(.douta(w_n5047_0[0]),.doutb(w_n5047_0[1]),.din(n5047));
	jspl jspl_w_n5049_0(.douta(w_n5049_0[0]),.doutb(w_n5049_0[1]),.din(n5049));
	jspl jspl_w_n5050_0(.douta(w_n5050_0[0]),.doutb(w_n5050_0[1]),.din(n5050));
	jspl3 jspl3_w_n5051_0(.douta(w_n5051_0[0]),.doutb(w_n5051_0[1]),.doutc(w_n5051_0[2]),.din(n5051));
	jspl jspl_w_n5052_0(.douta(w_n5052_0[0]),.doutb(w_n5052_0[1]),.din(n5052));
	jspl jspl_w_n5056_0(.douta(w_n5056_0[0]),.doutb(w_n5056_0[1]),.din(n5056));
	jspl jspl_w_n5062_0(.douta(w_n5062_0[0]),.doutb(w_n5062_0[1]),.din(n5062));
	jspl jspl_w_n5063_0(.douta(w_n5063_0[0]),.doutb(w_n5063_0[1]),.din(n5063));
	jspl jspl_w_n5065_0(.douta(w_n5065_0[0]),.doutb(w_n5065_0[1]),.din(n5065));
	jspl jspl_w_n5067_0(.douta(w_n5067_0[0]),.doutb(w_n5067_0[1]),.din(n5067));
	jspl jspl_w_n5070_0(.douta(w_n5070_0[0]),.doutb(w_n5070_0[1]),.din(n5070));
	jspl jspl_w_n5076_0(.douta(w_n5076_0[0]),.doutb(w_n5076_0[1]),.din(n5076));
	jspl jspl_w_n5078_0(.douta(w_n5078_0[0]),.doutb(w_n5078_0[1]),.din(n5078));
	jspl3 jspl3_w_n5079_0(.douta(w_n5079_0[0]),.doutb(w_n5079_0[1]),.doutc(w_n5079_0[2]),.din(n5079));
	jspl jspl_w_n5083_0(.douta(w_n5083_0[0]),.doutb(w_n5083_0[1]),.din(n5083));
	jspl jspl_w_n5084_0(.douta(w_n5084_0[0]),.doutb(w_n5084_0[1]),.din(n5084));
	jspl3 jspl3_w_n5085_0(.douta(w_n5085_0[0]),.doutb(w_n5085_0[1]),.doutc(w_n5085_0[2]),.din(n5085));
	jspl jspl_w_n5087_0(.douta(w_n5087_0[0]),.doutb(w_n5087_0[1]),.din(n5087));
	jspl jspl_w_n5092_0(.douta(w_n5092_0[0]),.doutb(w_n5092_0[1]),.din(n5092));
	jspl jspl_w_n5094_0(.douta(w_n5094_0[0]),.doutb(w_n5094_0[1]),.din(n5094));
	jspl jspl_w_n5095_0(.douta(w_n5095_0[0]),.doutb(w_n5095_0[1]),.din(n5095));
	jspl3 jspl3_w_n5096_0(.douta(w_n5096_0[0]),.doutb(w_n5096_0[1]),.doutc(w_n5096_0[2]),.din(n5096));
	jspl3 jspl3_w_n5096_1(.douta(w_n5096_1[0]),.doutb(w_n5096_1[1]),.doutc(w_n5096_1[2]),.din(w_n5096_0[0]));
	jspl jspl_w_n5099_0(.douta(w_n5099_0[0]),.doutb(w_n5099_0[1]),.din(n5099));
	jspl3 jspl3_w_n5100_0(.douta(w_n5100_0[0]),.doutb(w_n5100_0[1]),.doutc(w_n5100_0[2]),.din(n5100));
	jspl jspl_w_n5101_0(.douta(w_n5101_0[0]),.doutb(w_n5101_0[1]),.din(n5101));
	jspl jspl_w_n5102_0(.douta(w_n5102_0[0]),.doutb(w_n5102_0[1]),.din(n5102));
	jspl jspl_w_n5108_0(.douta(w_n5108_0[0]),.doutb(w_n5108_0[1]),.din(n5108));
	jspl3 jspl3_w_n5109_0(.douta(w_n5109_0[0]),.doutb(w_n5109_0[1]),.doutc(w_n5109_0[2]),.din(n5109));
	jspl jspl_w_n5110_0(.douta(w_n5110_0[0]),.doutb(w_n5110_0[1]),.din(n5110));
	jspl jspl_w_n5115_0(.douta(w_n5115_0[0]),.doutb(w_n5115_0[1]),.din(n5115));
	jspl3 jspl3_w_n5116_0(.douta(w_n5116_0[0]),.doutb(w_n5116_0[1]),.doutc(w_n5116_0[2]),.din(n5116));
	jspl3 jspl3_w_n5116_1(.douta(w_n5116_1[0]),.doutb(w_n5116_1[1]),.doutc(w_n5116_1[2]),.din(w_n5116_0[0]));
	jspl3 jspl3_w_n5116_2(.douta(w_n5116_2[0]),.doutb(w_n5116_2[1]),.doutc(w_n5116_2[2]),.din(w_n5116_0[1]));
	jspl3 jspl3_w_n5116_3(.douta(w_n5116_3[0]),.doutb(w_n5116_3[1]),.doutc(w_n5116_3[2]),.din(w_n5116_0[2]));
	jspl3 jspl3_w_n5116_4(.douta(w_n5116_4[0]),.doutb(w_n5116_4[1]),.doutc(w_n5116_4[2]),.din(w_n5116_1[0]));
	jspl3 jspl3_w_n5116_5(.douta(w_n5116_5[0]),.doutb(w_n5116_5[1]),.doutc(w_n5116_5[2]),.din(w_n5116_1[1]));
	jspl3 jspl3_w_n5116_6(.douta(w_n5116_6[0]),.doutb(w_n5116_6[1]),.doutc(w_n5116_6[2]),.din(w_n5116_1[2]));
	jspl3 jspl3_w_n5116_7(.douta(w_n5116_7[0]),.doutb(w_n5116_7[1]),.doutc(w_n5116_7[2]),.din(w_n5116_2[0]));
	jspl3 jspl3_w_n5116_8(.douta(w_n5116_8[0]),.doutb(w_n5116_8[1]),.doutc(w_n5116_8[2]),.din(w_n5116_2[1]));
	jspl3 jspl3_w_n5116_9(.douta(w_n5116_9[0]),.doutb(w_n5116_9[1]),.doutc(w_n5116_9[2]),.din(w_n5116_2[2]));
	jspl3 jspl3_w_n5116_10(.douta(w_n5116_10[0]),.doutb(w_n5116_10[1]),.doutc(w_n5116_10[2]),.din(w_n5116_3[0]));
	jspl3 jspl3_w_n5116_11(.douta(w_n5116_11[0]),.doutb(w_n5116_11[1]),.doutc(w_n5116_11[2]),.din(w_n5116_3[1]));
	jspl3 jspl3_w_n5116_12(.douta(w_n5116_12[0]),.doutb(w_n5116_12[1]),.doutc(w_n5116_12[2]),.din(w_n5116_3[2]));
	jspl3 jspl3_w_n5116_13(.douta(w_n5116_13[0]),.doutb(w_n5116_13[1]),.doutc(w_n5116_13[2]),.din(w_n5116_4[0]));
	jspl3 jspl3_w_n5116_14(.douta(w_n5116_14[0]),.doutb(w_n5116_14[1]),.doutc(w_n5116_14[2]),.din(w_n5116_4[1]));
	jspl3 jspl3_w_n5116_15(.douta(w_n5116_15[0]),.doutb(w_n5116_15[1]),.doutc(w_n5116_15[2]),.din(w_n5116_4[2]));
	jspl3 jspl3_w_n5116_16(.douta(w_n5116_16[0]),.doutb(w_n5116_16[1]),.doutc(w_n5116_16[2]),.din(w_n5116_5[0]));
	jspl3 jspl3_w_n5116_17(.douta(w_n5116_17[0]),.doutb(w_n5116_17[1]),.doutc(w_n5116_17[2]),.din(w_n5116_5[1]));
	jspl3 jspl3_w_n5116_18(.douta(w_n5116_18[0]),.doutb(w_n5116_18[1]),.doutc(w_n5116_18[2]),.din(w_n5116_5[2]));
	jspl3 jspl3_w_n5116_19(.douta(w_n5116_19[0]),.doutb(w_n5116_19[1]),.doutc(w_n5116_19[2]),.din(w_n5116_6[0]));
	jspl3 jspl3_w_n5116_20(.douta(w_n5116_20[0]),.doutb(w_n5116_20[1]),.doutc(w_n5116_20[2]),.din(w_n5116_6[1]));
	jspl3 jspl3_w_n5116_21(.douta(w_n5116_21[0]),.doutb(w_n5116_21[1]),.doutc(w_n5116_21[2]),.din(w_n5116_6[2]));
	jspl3 jspl3_w_n5121_0(.douta(w_n5121_0[0]),.doutb(w_n5121_0[1]),.doutc(w_n5121_0[2]),.din(n5121));
	jspl3 jspl3_w_n5121_1(.douta(w_n5121_1[0]),.doutb(w_n5121_1[1]),.doutc(w_n5121_1[2]),.din(w_n5121_0[0]));
	jspl3 jspl3_w_n5121_2(.douta(w_n5121_2[0]),.doutb(w_n5121_2[1]),.doutc(w_n5121_2[2]),.din(w_n5121_0[1]));
	jspl3 jspl3_w_n5121_3(.douta(w_n5121_3[0]),.doutb(w_n5121_3[1]),.doutc(w_n5121_3[2]),.din(w_n5121_0[2]));
	jspl3 jspl3_w_n5121_4(.douta(w_n5121_4[0]),.doutb(w_n5121_4[1]),.doutc(w_n5121_4[2]),.din(w_n5121_1[0]));
	jspl3 jspl3_w_n5121_5(.douta(w_n5121_5[0]),.doutb(w_n5121_5[1]),.doutc(w_n5121_5[2]),.din(w_n5121_1[1]));
	jspl3 jspl3_w_n5121_6(.douta(w_n5121_6[0]),.doutb(w_n5121_6[1]),.doutc(w_n5121_6[2]),.din(w_n5121_1[2]));
	jspl3 jspl3_w_n5121_7(.douta(w_n5121_7[0]),.doutb(w_n5121_7[1]),.doutc(w_n5121_7[2]),.din(w_n5121_2[0]));
	jspl3 jspl3_w_n5121_8(.douta(w_n5121_8[0]),.doutb(w_n5121_8[1]),.doutc(w_n5121_8[2]),.din(w_n5121_2[1]));
	jspl3 jspl3_w_n5121_9(.douta(w_n5121_9[0]),.doutb(w_n5121_9[1]),.doutc(w_n5121_9[2]),.din(w_n5121_2[2]));
	jspl3 jspl3_w_n5121_10(.douta(w_n5121_10[0]),.doutb(w_n5121_10[1]),.doutc(w_n5121_10[2]),.din(w_n5121_3[0]));
	jspl3 jspl3_w_n5121_11(.douta(w_n5121_11[0]),.doutb(w_n5121_11[1]),.doutc(w_n5121_11[2]),.din(w_n5121_3[1]));
	jspl3 jspl3_w_n5121_12(.douta(w_n5121_12[0]),.doutb(w_n5121_12[1]),.doutc(w_n5121_12[2]),.din(w_n5121_3[2]));
	jspl3 jspl3_w_n5121_13(.douta(w_n5121_13[0]),.doutb(w_n5121_13[1]),.doutc(w_n5121_13[2]),.din(w_n5121_4[0]));
	jspl3 jspl3_w_n5121_14(.douta(w_n5121_14[0]),.doutb(w_n5121_14[1]),.doutc(w_n5121_14[2]),.din(w_n5121_4[1]));
	jspl3 jspl3_w_n5121_15(.douta(w_n5121_15[0]),.doutb(w_n5121_15[1]),.doutc(w_n5121_15[2]),.din(w_n5121_4[2]));
	jspl3 jspl3_w_n5121_16(.douta(w_n5121_16[0]),.doutb(w_n5121_16[1]),.doutc(w_n5121_16[2]),.din(w_n5121_5[0]));
	jspl3 jspl3_w_n5121_17(.douta(w_n5121_17[0]),.doutb(w_n5121_17[1]),.doutc(w_n5121_17[2]),.din(w_n5121_5[1]));
	jspl3 jspl3_w_n5121_18(.douta(w_n5121_18[0]),.doutb(w_n5121_18[1]),.doutc(w_n5121_18[2]),.din(w_n5121_5[2]));
	jspl3 jspl3_w_n5121_19(.douta(w_n5121_19[0]),.doutb(w_n5121_19[1]),.doutc(w_n5121_19[2]),.din(w_n5121_6[0]));
	jspl3 jspl3_w_n5121_20(.douta(w_n5121_20[0]),.doutb(w_n5121_20[1]),.doutc(w_n5121_20[2]),.din(w_n5121_6[1]));
	jspl3 jspl3_w_n5121_21(.douta(w_n5121_21[0]),.doutb(w_n5121_21[1]),.doutc(w_n5121_21[2]),.din(w_n5121_6[2]));
	jspl3 jspl3_w_n5121_22(.douta(w_n5121_22[0]),.doutb(w_n5121_22[1]),.doutc(w_n5121_22[2]),.din(w_n5121_7[0]));
	jspl3 jspl3_w_n5121_23(.douta(w_n5121_23[0]),.doutb(w_n5121_23[1]),.doutc(w_n5121_23[2]),.din(w_n5121_7[1]));
	jspl3 jspl3_w_n5121_24(.douta(w_n5121_24[0]),.doutb(w_n5121_24[1]),.doutc(w_n5121_24[2]),.din(w_n5121_7[2]));
	jspl3 jspl3_w_n5121_25(.douta(w_n5121_25[0]),.doutb(w_n5121_25[1]),.doutc(w_n5121_25[2]),.din(w_n5121_8[0]));
	jspl3 jspl3_w_n5121_26(.douta(w_n5121_26[0]),.doutb(w_n5121_26[1]),.doutc(w_n5121_26[2]),.din(w_n5121_8[1]));
	jspl3 jspl3_w_n5121_27(.douta(w_n5121_27[0]),.doutb(w_n5121_27[1]),.doutc(w_n5121_27[2]),.din(w_n5121_8[2]));
	jspl3 jspl3_w_n5121_28(.douta(w_n5121_28[0]),.doutb(w_n5121_28[1]),.doutc(w_n5121_28[2]),.din(w_n5121_9[0]));
	jspl3 jspl3_w_n5121_29(.douta(w_n5121_29[0]),.doutb(w_n5121_29[1]),.doutc(w_n5121_29[2]),.din(w_n5121_9[1]));
	jspl3 jspl3_w_n5124_0(.douta(w_n5124_0[0]),.doutb(w_n5124_0[1]),.doutc(w_n5124_0[2]),.din(n5124));
	jspl jspl_w_n5124_1(.douta(w_n5124_1[0]),.doutb(w_n5124_1[1]),.din(w_n5124_0[0]));
	jspl3 jspl3_w_n5125_0(.douta(w_n5125_0[0]),.doutb(w_n5125_0[1]),.doutc(w_n5125_0[2]),.din(n5125));
	jspl3 jspl3_w_n5129_0(.douta(w_n5129_0[0]),.doutb(w_n5129_0[1]),.doutc(w_n5129_0[2]),.din(n5129));
	jspl jspl_w_n5130_0(.douta(w_n5130_0[0]),.doutb(w_n5130_0[1]),.din(n5130));
	jspl jspl_w_n5131_0(.douta(w_n5131_0[0]),.doutb(w_n5131_0[1]),.din(n5131));
	jspl jspl_w_n5132_0(.douta(w_n5132_0[0]),.doutb(w_n5132_0[1]),.din(n5132));
	jspl jspl_w_n5134_0(.douta(w_n5134_0[0]),.doutb(w_n5134_0[1]),.din(n5134));
	jspl jspl_w_n5136_0(.douta(w_n5136_0[0]),.doutb(w_n5136_0[1]),.din(n5136));
	jspl jspl_w_n5138_0(.douta(w_n5138_0[0]),.doutb(w_n5138_0[1]),.din(n5138));
	jspl jspl_w_n5141_0(.douta(w_n5141_0[0]),.doutb(w_n5141_0[1]),.din(n5141));
	jspl jspl_w_n5146_0(.douta(w_n5146_0[0]),.doutb(w_n5146_0[1]),.din(n5146));
	jspl3 jspl3_w_n5148_0(.douta(w_n5148_0[0]),.doutb(w_n5148_0[1]),.doutc(w_n5148_0[2]),.din(n5148));
	jspl jspl_w_n5149_0(.douta(w_n5149_0[0]),.doutb(w_n5149_0[1]),.din(n5149));
	jspl jspl_w_n5153_0(.douta(w_n5153_0[0]),.doutb(w_n5153_0[1]),.din(n5153));
	jspl jspl_w_n5154_0(.douta(w_n5154_0[0]),.doutb(w_n5154_0[1]),.din(n5154));
	jspl jspl_w_n5156_0(.douta(w_n5156_0[0]),.doutb(w_n5156_0[1]),.din(n5156));
	jspl jspl_w_n5160_0(.douta(w_n5160_0[0]),.doutb(w_n5160_0[1]),.din(n5160));
	jspl jspl_w_n5162_0(.douta(w_n5162_0[0]),.doutb(w_n5162_0[1]),.din(n5162));
	jspl jspl_w_n5163_0(.douta(w_n5163_0[0]),.doutb(w_n5163_0[1]),.din(n5163));
	jspl3 jspl3_w_n5164_0(.douta(w_n5164_0[0]),.doutb(w_n5164_0[1]),.doutc(w_n5164_0[2]),.din(n5164));
	jspl jspl_w_n5165_0(.douta(w_n5165_0[0]),.doutb(w_n5165_0[1]),.din(n5165));
	jspl jspl_w_n5169_0(.douta(w_n5169_0[0]),.doutb(w_n5169_0[1]),.din(n5169));
	jspl jspl_w_n5171_0(.douta(w_n5171_0[0]),.doutb(w_n5171_0[1]),.din(n5171));
	jspl jspl_w_n5173_0(.douta(w_n5173_0[0]),.doutb(w_n5173_0[1]),.din(n5173));
	jspl jspl_w_n5175_0(.douta(w_n5175_0[0]),.doutb(w_n5175_0[1]),.din(n5175));
	jspl jspl_w_n5177_0(.douta(w_n5177_0[0]),.doutb(w_n5177_0[1]),.din(n5177));
	jspl jspl_w_n5183_0(.douta(w_n5183_0[0]),.doutb(w_n5183_0[1]),.din(n5183));
	jspl3 jspl3_w_n5185_0(.douta(w_n5185_0[0]),.doutb(w_n5185_0[1]),.doutc(w_n5185_0[2]),.din(n5185));
	jspl jspl_w_n5186_0(.douta(w_n5186_0[0]),.doutb(w_n5186_0[1]),.din(n5186));
	jspl jspl_w_n5191_0(.douta(w_n5191_0[0]),.doutb(w_n5191_0[1]),.din(n5191));
	jspl jspl_w_n5193_0(.douta(w_n5193_0[0]),.doutb(w_n5193_0[1]),.din(n5193));
	jspl jspl_w_n5195_0(.douta(w_n5195_0[0]),.doutb(w_n5195_0[1]),.din(n5195));
	jspl jspl_w_n5199_0(.douta(w_n5199_0[0]),.doutb(w_n5199_0[1]),.din(n5199));
	jspl jspl_w_n5201_0(.douta(w_n5201_0[0]),.doutb(w_n5201_0[1]),.din(n5201));
	jspl jspl_w_n5202_0(.douta(w_n5202_0[0]),.doutb(w_n5202_0[1]),.din(n5202));
	jspl3 jspl3_w_n5203_0(.douta(w_n5203_0[0]),.doutb(w_n5203_0[1]),.doutc(w_n5203_0[2]),.din(n5203));
	jspl jspl_w_n5204_0(.douta(w_n5204_0[0]),.doutb(w_n5204_0[1]),.din(n5204));
	jspl jspl_w_n5210_0(.douta(w_n5210_0[0]),.doutb(w_n5210_0[1]),.din(n5210));
	jspl jspl_w_n5211_0(.douta(w_n5211_0[0]),.doutb(w_n5211_0[1]),.din(n5211));
	jspl jspl_w_n5213_0(.douta(w_n5213_0[0]),.doutb(w_n5213_0[1]),.din(n5213));
	jspl jspl_w_n5215_0(.douta(w_n5215_0[0]),.doutb(w_n5215_0[1]),.din(n5215));
	jspl jspl_w_n5217_0(.douta(w_n5217_0[0]),.doutb(w_n5217_0[1]),.din(n5217));
	jspl jspl_w_n5223_0(.douta(w_n5223_0[0]),.doutb(w_n5223_0[1]),.din(n5223));
	jspl jspl_w_n5225_0(.douta(w_n5225_0[0]),.doutb(w_n5225_0[1]),.din(n5225));
	jspl3 jspl3_w_n5226_0(.douta(w_n5226_0[0]),.doutb(w_n5226_0[1]),.doutc(w_n5226_0[2]),.din(n5226));
	jspl jspl_w_n5229_0(.douta(w_n5229_0[0]),.doutb(w_n5229_0[1]),.din(n5229));
	jspl jspl_w_n5230_0(.douta(w_n5230_0[0]),.doutb(w_n5230_0[1]),.din(n5230));
	jspl3 jspl3_w_n5231_0(.douta(w_n5231_0[0]),.doutb(w_n5231_0[1]),.doutc(w_n5231_0[2]),.din(n5231));
	jspl jspl_w_n5233_0(.douta(w_n5233_0[0]),.doutb(w_n5233_0[1]),.din(n5233));
	jspl jspl_w_n5237_0(.douta(w_n5237_0[0]),.doutb(w_n5237_0[1]),.din(n5237));
	jspl jspl_w_n5239_0(.douta(w_n5239_0[0]),.doutb(w_n5239_0[1]),.din(n5239));
	jspl jspl_w_n5240_0(.douta(w_n5240_0[0]),.doutb(w_n5240_0[1]),.din(n5240));
	jspl3 jspl3_w_n5241_0(.douta(w_n5241_0[0]),.doutb(w_n5241_0[1]),.doutc(w_n5241_0[2]),.din(n5241));
	jspl jspl_w_n5242_0(.douta(w_n5242_0[0]),.doutb(w_n5242_0[1]),.din(n5242));
	jspl jspl_w_n5245_0(.douta(w_n5245_0[0]),.doutb(w_n5245_0[1]),.din(n5245));
	jspl jspl_w_n5251_0(.douta(w_n5251_0[0]),.doutb(w_n5251_0[1]),.din(n5251));
	jspl jspl_w_n5252_0(.douta(w_n5252_0[0]),.doutb(w_n5252_0[1]),.din(n5252));
	jspl jspl_w_n5254_0(.douta(w_n5254_0[0]),.doutb(w_n5254_0[1]),.din(n5254));
	jspl jspl_w_n5256_0(.douta(w_n5256_0[0]),.doutb(w_n5256_0[1]),.din(n5256));
	jspl jspl_w_n5258_0(.douta(w_n5258_0[0]),.doutb(w_n5258_0[1]),.din(n5258));
	jspl jspl_w_n5264_0(.douta(w_n5264_0[0]),.doutb(w_n5264_0[1]),.din(n5264));
	jspl jspl_w_n5266_0(.douta(w_n5266_0[0]),.doutb(w_n5266_0[1]),.din(n5266));
	jspl3 jspl3_w_n5267_0(.douta(w_n5267_0[0]),.doutb(w_n5267_0[1]),.doutc(w_n5267_0[2]),.din(n5267));
	jspl jspl_w_n5270_0(.douta(w_n5270_0[0]),.doutb(w_n5270_0[1]),.din(n5270));
	jspl jspl_w_n5271_0(.douta(w_n5271_0[0]),.doutb(w_n5271_0[1]),.din(n5271));
	jspl3 jspl3_w_n5272_0(.douta(w_n5272_0[0]),.doutb(w_n5272_0[1]),.doutc(w_n5272_0[2]),.din(n5272));
	jspl jspl_w_n5274_0(.douta(w_n5274_0[0]),.doutb(w_n5274_0[1]),.din(n5274));
	jspl jspl_w_n5278_0(.douta(w_n5278_0[0]),.doutb(w_n5278_0[1]),.din(n5278));
	jspl jspl_w_n5280_0(.douta(w_n5280_0[0]),.doutb(w_n5280_0[1]),.din(n5280));
	jspl jspl_w_n5281_0(.douta(w_n5281_0[0]),.doutb(w_n5281_0[1]),.din(n5281));
	jspl3 jspl3_w_n5282_0(.douta(w_n5282_0[0]),.doutb(w_n5282_0[1]),.doutc(w_n5282_0[2]),.din(n5282));
	jspl jspl_w_n5283_0(.douta(w_n5283_0[0]),.doutb(w_n5283_0[1]),.din(n5283));
	jspl jspl_w_n5286_0(.douta(w_n5286_0[0]),.doutb(w_n5286_0[1]),.din(n5286));
	jspl jspl_w_n5292_0(.douta(w_n5292_0[0]),.doutb(w_n5292_0[1]),.din(n5292));
	jspl jspl_w_n5293_0(.douta(w_n5293_0[0]),.doutb(w_n5293_0[1]),.din(n5293));
	jspl jspl_w_n5295_0(.douta(w_n5295_0[0]),.doutb(w_n5295_0[1]),.din(n5295));
	jspl jspl_w_n5297_0(.douta(w_n5297_0[0]),.doutb(w_n5297_0[1]),.din(n5297));
	jspl jspl_w_n5299_0(.douta(w_n5299_0[0]),.doutb(w_n5299_0[1]),.din(n5299));
	jspl jspl_w_n5305_0(.douta(w_n5305_0[0]),.doutb(w_n5305_0[1]),.din(n5305));
	jspl jspl_w_n5307_0(.douta(w_n5307_0[0]),.doutb(w_n5307_0[1]),.din(n5307));
	jspl3 jspl3_w_n5308_0(.douta(w_n5308_0[0]),.doutb(w_n5308_0[1]),.doutc(w_n5308_0[2]),.din(n5308));
	jspl jspl_w_n5311_0(.douta(w_n5311_0[0]),.doutb(w_n5311_0[1]),.din(n5311));
	jspl jspl_w_n5312_0(.douta(w_n5312_0[0]),.doutb(w_n5312_0[1]),.din(n5312));
	jspl3 jspl3_w_n5313_0(.douta(w_n5313_0[0]),.doutb(w_n5313_0[1]),.doutc(w_n5313_0[2]),.din(n5313));
	jspl jspl_w_n5315_0(.douta(w_n5315_0[0]),.doutb(w_n5315_0[1]),.din(n5315));
	jspl jspl_w_n5319_0(.douta(w_n5319_0[0]),.doutb(w_n5319_0[1]),.din(n5319));
	jspl jspl_w_n5321_0(.douta(w_n5321_0[0]),.doutb(w_n5321_0[1]),.din(n5321));
	jspl jspl_w_n5322_0(.douta(w_n5322_0[0]),.doutb(w_n5322_0[1]),.din(n5322));
	jspl3 jspl3_w_n5323_0(.douta(w_n5323_0[0]),.doutb(w_n5323_0[1]),.doutc(w_n5323_0[2]),.din(n5323));
	jspl jspl_w_n5324_0(.douta(w_n5324_0[0]),.doutb(w_n5324_0[1]),.din(n5324));
	jspl jspl_w_n5327_0(.douta(w_n5327_0[0]),.doutb(w_n5327_0[1]),.din(n5327));
	jspl jspl_w_n5333_0(.douta(w_n5333_0[0]),.doutb(w_n5333_0[1]),.din(n5333));
	jspl jspl_w_n5334_0(.douta(w_n5334_0[0]),.doutb(w_n5334_0[1]),.din(n5334));
	jspl jspl_w_n5336_0(.douta(w_n5336_0[0]),.doutb(w_n5336_0[1]),.din(n5336));
	jspl jspl_w_n5338_0(.douta(w_n5338_0[0]),.doutb(w_n5338_0[1]),.din(n5338));
	jspl jspl_w_n5340_0(.douta(w_n5340_0[0]),.doutb(w_n5340_0[1]),.din(n5340));
	jspl jspl_w_n5346_0(.douta(w_n5346_0[0]),.doutb(w_n5346_0[1]),.din(n5346));
	jspl jspl_w_n5348_0(.douta(w_n5348_0[0]),.doutb(w_n5348_0[1]),.din(n5348));
	jspl3 jspl3_w_n5349_0(.douta(w_n5349_0[0]),.doutb(w_n5349_0[1]),.doutc(w_n5349_0[2]),.din(n5349));
	jspl jspl_w_n5352_0(.douta(w_n5352_0[0]),.doutb(w_n5352_0[1]),.din(n5352));
	jspl jspl_w_n5353_0(.douta(w_n5353_0[0]),.doutb(w_n5353_0[1]),.din(n5353));
	jspl3 jspl3_w_n5354_0(.douta(w_n5354_0[0]),.doutb(w_n5354_0[1]),.doutc(w_n5354_0[2]),.din(n5354));
	jspl jspl_w_n5356_0(.douta(w_n5356_0[0]),.doutb(w_n5356_0[1]),.din(n5356));
	jspl jspl_w_n5360_0(.douta(w_n5360_0[0]),.doutb(w_n5360_0[1]),.din(n5360));
	jspl jspl_w_n5362_0(.douta(w_n5362_0[0]),.doutb(w_n5362_0[1]),.din(n5362));
	jspl jspl_w_n5363_0(.douta(w_n5363_0[0]),.doutb(w_n5363_0[1]),.din(n5363));
	jspl3 jspl3_w_n5364_0(.douta(w_n5364_0[0]),.doutb(w_n5364_0[1]),.doutc(w_n5364_0[2]),.din(n5364));
	jspl jspl_w_n5365_0(.douta(w_n5365_0[0]),.doutb(w_n5365_0[1]),.din(n5365));
	jspl jspl_w_n5368_0(.douta(w_n5368_0[0]),.doutb(w_n5368_0[1]),.din(n5368));
	jspl jspl_w_n5374_0(.douta(w_n5374_0[0]),.doutb(w_n5374_0[1]),.din(n5374));
	jspl jspl_w_n5375_0(.douta(w_n5375_0[0]),.doutb(w_n5375_0[1]),.din(n5375));
	jspl jspl_w_n5377_0(.douta(w_n5377_0[0]),.doutb(w_n5377_0[1]),.din(n5377));
	jspl jspl_w_n5379_0(.douta(w_n5379_0[0]),.doutb(w_n5379_0[1]),.din(n5379));
	jspl jspl_w_n5381_0(.douta(w_n5381_0[0]),.doutb(w_n5381_0[1]),.din(n5381));
	jspl jspl_w_n5387_0(.douta(w_n5387_0[0]),.doutb(w_n5387_0[1]),.din(n5387));
	jspl jspl_w_n5389_0(.douta(w_n5389_0[0]),.doutb(w_n5389_0[1]),.din(n5389));
	jspl3 jspl3_w_n5390_0(.douta(w_n5390_0[0]),.doutb(w_n5390_0[1]),.doutc(w_n5390_0[2]),.din(n5390));
	jspl jspl_w_n5393_0(.douta(w_n5393_0[0]),.doutb(w_n5393_0[1]),.din(n5393));
	jspl jspl_w_n5394_0(.douta(w_n5394_0[0]),.doutb(w_n5394_0[1]),.din(n5394));
	jspl3 jspl3_w_n5395_0(.douta(w_n5395_0[0]),.doutb(w_n5395_0[1]),.doutc(w_n5395_0[2]),.din(n5395));
	jspl jspl_w_n5397_0(.douta(w_n5397_0[0]),.doutb(w_n5397_0[1]),.din(n5397));
	jspl jspl_w_n5401_0(.douta(w_n5401_0[0]),.doutb(w_n5401_0[1]),.din(n5401));
	jspl jspl_w_n5403_0(.douta(w_n5403_0[0]),.doutb(w_n5403_0[1]),.din(n5403));
	jspl jspl_w_n5404_0(.douta(w_n5404_0[0]),.doutb(w_n5404_0[1]),.din(n5404));
	jspl3 jspl3_w_n5405_0(.douta(w_n5405_0[0]),.doutb(w_n5405_0[1]),.doutc(w_n5405_0[2]),.din(n5405));
	jspl jspl_w_n5409_0(.douta(w_n5409_0[0]),.doutb(w_n5409_0[1]),.din(n5409));
	jspl jspl_w_n5415_0(.douta(w_n5415_0[0]),.doutb(w_n5415_0[1]),.din(n5415));
	jspl3 jspl3_w_n5417_0(.douta(w_n5417_0[0]),.doutb(w_n5417_0[1]),.doutc(w_n5417_0[2]),.din(n5417));
	jspl jspl_w_n5419_0(.douta(w_n5419_0[0]),.doutb(w_n5419_0[1]),.din(n5419));
	jspl3 jspl3_w_n5424_0(.douta(w_n5424_0[0]),.doutb(w_n5424_0[1]),.doutc(w_n5424_0[2]),.din(n5424));
	jspl jspl_w_n5425_0(.douta(w_n5425_0[0]),.doutb(w_n5425_0[1]),.din(n5425));
	jspl jspl_w_n5426_0(.douta(w_n5426_0[0]),.doutb(w_n5426_0[1]),.din(n5426));
	jspl jspl_w_n5431_0(.douta(w_n5431_0[0]),.doutb(w_n5431_0[1]),.din(n5431));
	jspl3 jspl3_w_n5432_0(.douta(w_n5432_0[0]),.doutb(w_n5432_0[1]),.doutc(w_n5432_0[2]),.din(n5432));
	jspl jspl_w_n5437_0(.douta(w_n5437_0[0]),.doutb(w_n5437_0[1]),.din(n5437));
	jspl3 jspl3_w_n5443_0(.douta(w_n5443_0[0]),.doutb(w_n5443_0[1]),.doutc(w_n5443_0[2]),.din(n5443));
	jspl jspl_w_n5443_1(.douta(w_n5443_1[0]),.doutb(w_n5443_1[1]),.din(w_n5443_0[0]));
	jspl3 jspl3_w_n5446_0(.douta(w_n5446_0[0]),.doutb(w_n5446_0[1]),.doutc(w_n5446_0[2]),.din(n5446));
	jspl jspl_w_n5447_0(.douta(w_n5447_0[0]),.doutb(w_n5447_0[1]),.din(n5447));
	jspl jspl_w_n5448_0(.douta(w_n5448_0[0]),.doutb(w_n5448_0[1]),.din(n5448));
	jspl jspl_w_n5449_0(.douta(w_n5449_0[0]),.doutb(w_n5449_0[1]),.din(n5449));
	jspl jspl_w_n5451_0(.douta(w_n5451_0[0]),.doutb(w_n5451_0[1]),.din(n5451));
	jspl jspl_w_n5453_0(.douta(w_n5453_0[0]),.doutb(w_n5453_0[1]),.din(n5453));
	jspl jspl_w_n5455_0(.douta(w_n5455_0[0]),.doutb(w_n5455_0[1]),.din(n5455));
	jspl jspl_w_n5464_0(.douta(w_n5464_0[0]),.doutb(w_n5464_0[1]),.din(n5464));
	jspl3 jspl3_w_n5466_0(.douta(w_n5466_0[0]),.doutb(w_n5466_0[1]),.doutc(w_n5466_0[2]),.din(n5466));
	jspl jspl_w_n5467_0(.douta(w_n5467_0[0]),.doutb(w_n5467_0[1]),.din(n5467));
	jspl jspl_w_n5471_0(.douta(w_n5471_0[0]),.doutb(w_n5471_0[1]),.din(n5471));
	jspl jspl_w_n5473_0(.douta(w_n5473_0[0]),.doutb(w_n5473_0[1]),.din(n5473));
	jspl jspl_w_n5475_0(.douta(w_n5475_0[0]),.doutb(w_n5475_0[1]),.din(n5475));
	jspl jspl_w_n5480_0(.douta(w_n5480_0[0]),.doutb(w_n5480_0[1]),.din(n5480));
	jspl jspl_w_n5482_0(.douta(w_n5482_0[0]),.doutb(w_n5482_0[1]),.din(n5482));
	jspl jspl_w_n5483_0(.douta(w_n5483_0[0]),.doutb(w_n5483_0[1]),.din(n5483));
	jspl3 jspl3_w_n5484_0(.douta(w_n5484_0[0]),.doutb(w_n5484_0[1]),.doutc(w_n5484_0[2]),.din(n5484));
	jspl jspl_w_n5485_0(.douta(w_n5485_0[0]),.doutb(w_n5485_0[1]),.din(n5485));
	jspl jspl_w_n5490_0(.douta(w_n5490_0[0]),.doutb(w_n5490_0[1]),.din(n5490));
	jspl jspl_w_n5491_0(.douta(w_n5491_0[0]),.doutb(w_n5491_0[1]),.din(n5491));
	jspl jspl_w_n5493_0(.douta(w_n5493_0[0]),.doutb(w_n5493_0[1]),.din(n5493));
	jspl jspl_w_n5495_0(.douta(w_n5495_0[0]),.doutb(w_n5495_0[1]),.din(n5495));
	jspl jspl_w_n5498_0(.douta(w_n5498_0[0]),.doutb(w_n5498_0[1]),.din(n5498));
	jspl jspl_w_n5504_0(.douta(w_n5504_0[0]),.doutb(w_n5504_0[1]),.din(n5504));
	jspl3 jspl3_w_n5506_0(.douta(w_n5506_0[0]),.doutb(w_n5506_0[1]),.doutc(w_n5506_0[2]),.din(n5506));
	jspl jspl_w_n5507_0(.douta(w_n5507_0[0]),.doutb(w_n5507_0[1]),.din(n5507));
	jspl jspl_w_n5511_0(.douta(w_n5511_0[0]),.doutb(w_n5511_0[1]),.din(n5511));
	jspl jspl_w_n5512_0(.douta(w_n5512_0[0]),.doutb(w_n5512_0[1]),.din(n5512));
	jspl jspl_w_n5514_0(.douta(w_n5514_0[0]),.doutb(w_n5514_0[1]),.din(n5514));
	jspl jspl_w_n5519_0(.douta(w_n5519_0[0]),.doutb(w_n5519_0[1]),.din(n5519));
	jspl jspl_w_n5521_0(.douta(w_n5521_0[0]),.doutb(w_n5521_0[1]),.din(n5521));
	jspl jspl_w_n5522_0(.douta(w_n5522_0[0]),.doutb(w_n5522_0[1]),.din(n5522));
	jspl3 jspl3_w_n5523_0(.douta(w_n5523_0[0]),.doutb(w_n5523_0[1]),.doutc(w_n5523_0[2]),.din(n5523));
	jspl jspl_w_n5524_0(.douta(w_n5524_0[0]),.doutb(w_n5524_0[1]),.din(n5524));
	jspl jspl_w_n5528_0(.douta(w_n5528_0[0]),.doutb(w_n5528_0[1]),.din(n5528));
	jspl jspl_w_n5529_0(.douta(w_n5529_0[0]),.doutb(w_n5529_0[1]),.din(n5529));
	jspl jspl_w_n5531_0(.douta(w_n5531_0[0]),.doutb(w_n5531_0[1]),.din(n5531));
	jspl jspl_w_n5533_0(.douta(w_n5533_0[0]),.doutb(w_n5533_0[1]),.din(n5533));
	jspl jspl_w_n5536_0(.douta(w_n5536_0[0]),.doutb(w_n5536_0[1]),.din(n5536));
	jspl jspl_w_n5542_0(.douta(w_n5542_0[0]),.doutb(w_n5542_0[1]),.din(n5542));
	jspl jspl_w_n5544_0(.douta(w_n5544_0[0]),.doutb(w_n5544_0[1]),.din(n5544));
	jspl3 jspl3_w_n5545_0(.douta(w_n5545_0[0]),.doutb(w_n5545_0[1]),.doutc(w_n5545_0[2]),.din(n5545));
	jspl jspl_w_n5549_0(.douta(w_n5549_0[0]),.doutb(w_n5549_0[1]),.din(n5549));
	jspl jspl_w_n5550_0(.douta(w_n5550_0[0]),.doutb(w_n5550_0[1]),.din(n5550));
	jspl3 jspl3_w_n5551_0(.douta(w_n5551_0[0]),.doutb(w_n5551_0[1]),.doutc(w_n5551_0[2]),.din(n5551));
	jspl jspl_w_n5553_0(.douta(w_n5553_0[0]),.doutb(w_n5553_0[1]),.din(n5553));
	jspl jspl_w_n5558_0(.douta(w_n5558_0[0]),.doutb(w_n5558_0[1]),.din(n5558));
	jspl jspl_w_n5560_0(.douta(w_n5560_0[0]),.doutb(w_n5560_0[1]),.din(n5560));
	jspl jspl_w_n5561_0(.douta(w_n5561_0[0]),.doutb(w_n5561_0[1]),.din(n5561));
	jspl3 jspl3_w_n5562_0(.douta(w_n5562_0[0]),.doutb(w_n5562_0[1]),.doutc(w_n5562_0[2]),.din(n5562));
	jspl jspl_w_n5563_0(.douta(w_n5563_0[0]),.doutb(w_n5563_0[1]),.din(n5563));
	jspl jspl_w_n5567_0(.douta(w_n5567_0[0]),.doutb(w_n5567_0[1]),.din(n5567));
	jspl jspl_w_n5573_0(.douta(w_n5573_0[0]),.doutb(w_n5573_0[1]),.din(n5573));
	jspl jspl_w_n5574_0(.douta(w_n5574_0[0]),.doutb(w_n5574_0[1]),.din(n5574));
	jspl jspl_w_n5576_0(.douta(w_n5576_0[0]),.doutb(w_n5576_0[1]),.din(n5576));
	jspl jspl_w_n5578_0(.douta(w_n5578_0[0]),.doutb(w_n5578_0[1]),.din(n5578));
	jspl jspl_w_n5581_0(.douta(w_n5581_0[0]),.doutb(w_n5581_0[1]),.din(n5581));
	jspl jspl_w_n5587_0(.douta(w_n5587_0[0]),.doutb(w_n5587_0[1]),.din(n5587));
	jspl jspl_w_n5589_0(.douta(w_n5589_0[0]),.doutb(w_n5589_0[1]),.din(n5589));
	jspl3 jspl3_w_n5590_0(.douta(w_n5590_0[0]),.doutb(w_n5590_0[1]),.doutc(w_n5590_0[2]),.din(n5590));
	jspl jspl_w_n5594_0(.douta(w_n5594_0[0]),.doutb(w_n5594_0[1]),.din(n5594));
	jspl jspl_w_n5595_0(.douta(w_n5595_0[0]),.doutb(w_n5595_0[1]),.din(n5595));
	jspl3 jspl3_w_n5596_0(.douta(w_n5596_0[0]),.doutb(w_n5596_0[1]),.doutc(w_n5596_0[2]),.din(n5596));
	jspl jspl_w_n5598_0(.douta(w_n5598_0[0]),.doutb(w_n5598_0[1]),.din(n5598));
	jspl jspl_w_n5603_0(.douta(w_n5603_0[0]),.doutb(w_n5603_0[1]),.din(n5603));
	jspl jspl_w_n5605_0(.douta(w_n5605_0[0]),.doutb(w_n5605_0[1]),.din(n5605));
	jspl jspl_w_n5606_0(.douta(w_n5606_0[0]),.doutb(w_n5606_0[1]),.din(n5606));
	jspl3 jspl3_w_n5607_0(.douta(w_n5607_0[0]),.doutb(w_n5607_0[1]),.doutc(w_n5607_0[2]),.din(n5607));
	jspl jspl_w_n5608_0(.douta(w_n5608_0[0]),.doutb(w_n5608_0[1]),.din(n5608));
	jspl jspl_w_n5612_0(.douta(w_n5612_0[0]),.doutb(w_n5612_0[1]),.din(n5612));
	jspl jspl_w_n5618_0(.douta(w_n5618_0[0]),.doutb(w_n5618_0[1]),.din(n5618));
	jspl jspl_w_n5619_0(.douta(w_n5619_0[0]),.doutb(w_n5619_0[1]),.din(n5619));
	jspl jspl_w_n5621_0(.douta(w_n5621_0[0]),.doutb(w_n5621_0[1]),.din(n5621));
	jspl jspl_w_n5623_0(.douta(w_n5623_0[0]),.doutb(w_n5623_0[1]),.din(n5623));
	jspl jspl_w_n5626_0(.douta(w_n5626_0[0]),.doutb(w_n5626_0[1]),.din(n5626));
	jspl jspl_w_n5632_0(.douta(w_n5632_0[0]),.doutb(w_n5632_0[1]),.din(n5632));
	jspl jspl_w_n5634_0(.douta(w_n5634_0[0]),.doutb(w_n5634_0[1]),.din(n5634));
	jspl3 jspl3_w_n5635_0(.douta(w_n5635_0[0]),.doutb(w_n5635_0[1]),.doutc(w_n5635_0[2]),.din(n5635));
	jspl jspl_w_n5639_0(.douta(w_n5639_0[0]),.doutb(w_n5639_0[1]),.din(n5639));
	jspl jspl_w_n5640_0(.douta(w_n5640_0[0]),.doutb(w_n5640_0[1]),.din(n5640));
	jspl3 jspl3_w_n5641_0(.douta(w_n5641_0[0]),.doutb(w_n5641_0[1]),.doutc(w_n5641_0[2]),.din(n5641));
	jspl jspl_w_n5643_0(.douta(w_n5643_0[0]),.doutb(w_n5643_0[1]),.din(n5643));
	jspl jspl_w_n5648_0(.douta(w_n5648_0[0]),.doutb(w_n5648_0[1]),.din(n5648));
	jspl jspl_w_n5650_0(.douta(w_n5650_0[0]),.doutb(w_n5650_0[1]),.din(n5650));
	jspl jspl_w_n5651_0(.douta(w_n5651_0[0]),.doutb(w_n5651_0[1]),.din(n5651));
	jspl3 jspl3_w_n5652_0(.douta(w_n5652_0[0]),.doutb(w_n5652_0[1]),.doutc(w_n5652_0[2]),.din(n5652));
	jspl jspl_w_n5653_0(.douta(w_n5653_0[0]),.doutb(w_n5653_0[1]),.din(n5653));
	jspl jspl_w_n5657_0(.douta(w_n5657_0[0]),.doutb(w_n5657_0[1]),.din(n5657));
	jspl jspl_w_n5663_0(.douta(w_n5663_0[0]),.doutb(w_n5663_0[1]),.din(n5663));
	jspl jspl_w_n5664_0(.douta(w_n5664_0[0]),.doutb(w_n5664_0[1]),.din(n5664));
	jspl jspl_w_n5666_0(.douta(w_n5666_0[0]),.doutb(w_n5666_0[1]),.din(n5666));
	jspl jspl_w_n5668_0(.douta(w_n5668_0[0]),.doutb(w_n5668_0[1]),.din(n5668));
	jspl jspl_w_n5671_0(.douta(w_n5671_0[0]),.doutb(w_n5671_0[1]),.din(n5671));
	jspl jspl_w_n5677_0(.douta(w_n5677_0[0]),.doutb(w_n5677_0[1]),.din(n5677));
	jspl jspl_w_n5679_0(.douta(w_n5679_0[0]),.doutb(w_n5679_0[1]),.din(n5679));
	jspl3 jspl3_w_n5680_0(.douta(w_n5680_0[0]),.doutb(w_n5680_0[1]),.doutc(w_n5680_0[2]),.din(n5680));
	jspl jspl_w_n5684_0(.douta(w_n5684_0[0]),.doutb(w_n5684_0[1]),.din(n5684));
	jspl jspl_w_n5685_0(.douta(w_n5685_0[0]),.doutb(w_n5685_0[1]),.din(n5685));
	jspl3 jspl3_w_n5686_0(.douta(w_n5686_0[0]),.doutb(w_n5686_0[1]),.doutc(w_n5686_0[2]),.din(n5686));
	jspl jspl_w_n5688_0(.douta(w_n5688_0[0]),.doutb(w_n5688_0[1]),.din(n5688));
	jspl jspl_w_n5693_0(.douta(w_n5693_0[0]),.doutb(w_n5693_0[1]),.din(n5693));
	jspl jspl_w_n5695_0(.douta(w_n5695_0[0]),.doutb(w_n5695_0[1]),.din(n5695));
	jspl jspl_w_n5696_0(.douta(w_n5696_0[0]),.doutb(w_n5696_0[1]),.din(n5696));
	jspl3 jspl3_w_n5697_0(.douta(w_n5697_0[0]),.doutb(w_n5697_0[1]),.doutc(w_n5697_0[2]),.din(n5697));
	jspl jspl_w_n5698_0(.douta(w_n5698_0[0]),.doutb(w_n5698_0[1]),.din(n5698));
	jspl jspl_w_n5702_0(.douta(w_n5702_0[0]),.doutb(w_n5702_0[1]),.din(n5702));
	jspl jspl_w_n5708_0(.douta(w_n5708_0[0]),.doutb(w_n5708_0[1]),.din(n5708));
	jspl jspl_w_n5709_0(.douta(w_n5709_0[0]),.doutb(w_n5709_0[1]),.din(n5709));
	jspl jspl_w_n5711_0(.douta(w_n5711_0[0]),.doutb(w_n5711_0[1]),.din(n5711));
	jspl jspl_w_n5713_0(.douta(w_n5713_0[0]),.doutb(w_n5713_0[1]),.din(n5713));
	jspl jspl_w_n5716_0(.douta(w_n5716_0[0]),.doutb(w_n5716_0[1]),.din(n5716));
	jspl jspl_w_n5722_0(.douta(w_n5722_0[0]),.doutb(w_n5722_0[1]),.din(n5722));
	jspl jspl_w_n5724_0(.douta(w_n5724_0[0]),.doutb(w_n5724_0[1]),.din(n5724));
	jspl3 jspl3_w_n5725_0(.douta(w_n5725_0[0]),.doutb(w_n5725_0[1]),.doutc(w_n5725_0[2]),.din(n5725));
	jspl jspl_w_n5729_0(.douta(w_n5729_0[0]),.doutb(w_n5729_0[1]),.din(n5729));
	jspl jspl_w_n5730_0(.douta(w_n5730_0[0]),.doutb(w_n5730_0[1]),.din(n5730));
	jspl3 jspl3_w_n5731_0(.douta(w_n5731_0[0]),.doutb(w_n5731_0[1]),.doutc(w_n5731_0[2]),.din(n5731));
	jspl jspl_w_n5733_0(.douta(w_n5733_0[0]),.doutb(w_n5733_0[1]),.din(n5733));
	jspl jspl_w_n5738_0(.douta(w_n5738_0[0]),.doutb(w_n5738_0[1]),.din(n5738));
	jspl jspl_w_n5740_0(.douta(w_n5740_0[0]),.doutb(w_n5740_0[1]),.din(n5740));
	jspl jspl_w_n5741_0(.douta(w_n5741_0[0]),.doutb(w_n5741_0[1]),.din(n5741));
	jspl3 jspl3_w_n5742_0(.douta(w_n5742_0[0]),.doutb(w_n5742_0[1]),.doutc(w_n5742_0[2]),.din(n5742));
	jspl jspl_w_n5743_0(.douta(w_n5743_0[0]),.doutb(w_n5743_0[1]),.din(n5743));
	jspl jspl_w_n5747_0(.douta(w_n5747_0[0]),.doutb(w_n5747_0[1]),.din(n5747));
	jspl jspl_w_n5753_0(.douta(w_n5753_0[0]),.doutb(w_n5753_0[1]),.din(n5753));
	jspl jspl_w_n5754_0(.douta(w_n5754_0[0]),.doutb(w_n5754_0[1]),.din(n5754));
	jspl jspl_w_n5756_0(.douta(w_n5756_0[0]),.doutb(w_n5756_0[1]),.din(n5756));
	jspl jspl_w_n5758_0(.douta(w_n5758_0[0]),.doutb(w_n5758_0[1]),.din(n5758));
	jspl jspl_w_n5761_0(.douta(w_n5761_0[0]),.doutb(w_n5761_0[1]),.din(n5761));
	jspl jspl_w_n5767_0(.douta(w_n5767_0[0]),.doutb(w_n5767_0[1]),.din(n5767));
	jspl3 jspl3_w_n5769_0(.douta(w_n5769_0[0]),.doutb(w_n5769_0[1]),.doutc(w_n5769_0[2]),.din(n5769));
	jspl3 jspl3_w_n5769_1(.douta(w_n5769_1[0]),.doutb(w_n5769_1[1]),.doutc(w_n5769_1[2]),.din(w_n5769_0[0]));
	jspl jspl_w_n5772_0(.douta(w_n5772_0[0]),.doutb(w_n5772_0[1]),.din(n5772));
	jspl3 jspl3_w_n5773_0(.douta(w_n5773_0[0]),.doutb(w_n5773_0[1]),.doutc(w_n5773_0[2]),.din(n5773));
	jspl jspl_w_n5774_0(.douta(w_n5774_0[0]),.doutb(w_n5774_0[1]),.din(n5774));
	jspl jspl_w_n5780_0(.douta(w_n5780_0[0]),.doutb(w_n5780_0[1]),.din(n5780));
	jspl3 jspl3_w_n5781_0(.douta(w_n5781_0[0]),.doutb(w_n5781_0[1]),.doutc(w_n5781_0[2]),.din(n5781));
	jspl jspl_w_n5782_0(.douta(w_n5782_0[0]),.doutb(w_n5782_0[1]),.din(n5782));
	jspl jspl_w_n5787_0(.douta(w_n5787_0[0]),.doutb(w_n5787_0[1]),.din(n5787));
	jspl3 jspl3_w_n5788_0(.douta(w_n5788_0[0]),.doutb(w_n5788_0[1]),.doutc(w_n5788_0[2]),.din(n5788));
	jspl3 jspl3_w_n5788_1(.douta(w_n5788_1[0]),.doutb(w_n5788_1[1]),.doutc(w_n5788_1[2]),.din(w_n5788_0[0]));
	jspl3 jspl3_w_n5788_2(.douta(w_n5788_2[0]),.doutb(w_n5788_2[1]),.doutc(w_n5788_2[2]),.din(w_n5788_0[1]));
	jspl3 jspl3_w_n5788_3(.douta(w_n5788_3[0]),.doutb(w_n5788_3[1]),.doutc(w_n5788_3[2]),.din(w_n5788_0[2]));
	jspl3 jspl3_w_n5788_4(.douta(w_n5788_4[0]),.doutb(w_n5788_4[1]),.doutc(w_n5788_4[2]),.din(w_n5788_1[0]));
	jspl3 jspl3_w_n5788_5(.douta(w_n5788_5[0]),.doutb(w_n5788_5[1]),.doutc(w_n5788_5[2]),.din(w_n5788_1[1]));
	jspl3 jspl3_w_n5788_6(.douta(w_n5788_6[0]),.doutb(w_n5788_6[1]),.doutc(w_n5788_6[2]),.din(w_n5788_1[2]));
	jspl3 jspl3_w_n5788_7(.douta(w_n5788_7[0]),.doutb(w_n5788_7[1]),.doutc(w_n5788_7[2]),.din(w_n5788_2[0]));
	jspl3 jspl3_w_n5788_8(.douta(w_n5788_8[0]),.doutb(w_n5788_8[1]),.doutc(w_n5788_8[2]),.din(w_n5788_2[1]));
	jspl3 jspl3_w_n5788_9(.douta(w_n5788_9[0]),.doutb(w_n5788_9[1]),.doutc(w_n5788_9[2]),.din(w_n5788_2[2]));
	jspl3 jspl3_w_n5788_10(.douta(w_n5788_10[0]),.doutb(w_n5788_10[1]),.doutc(w_n5788_10[2]),.din(w_n5788_3[0]));
	jspl3 jspl3_w_n5788_11(.douta(w_n5788_11[0]),.doutb(w_n5788_11[1]),.doutc(w_n5788_11[2]),.din(w_n5788_3[1]));
	jspl3 jspl3_w_n5788_12(.douta(w_n5788_12[0]),.doutb(w_n5788_12[1]),.doutc(w_n5788_12[2]),.din(w_n5788_3[2]));
	jspl3 jspl3_w_n5788_13(.douta(w_n5788_13[0]),.doutb(w_n5788_13[1]),.doutc(w_n5788_13[2]),.din(w_n5788_4[0]));
	jspl3 jspl3_w_n5788_14(.douta(w_n5788_14[0]),.doutb(w_n5788_14[1]),.doutc(w_n5788_14[2]),.din(w_n5788_4[1]));
	jspl3 jspl3_w_n5788_15(.douta(w_n5788_15[0]),.doutb(w_n5788_15[1]),.doutc(w_n5788_15[2]),.din(w_n5788_4[2]));
	jspl3 jspl3_w_n5788_16(.douta(w_n5788_16[0]),.doutb(w_n5788_16[1]),.doutc(w_n5788_16[2]),.din(w_n5788_5[0]));
	jspl3 jspl3_w_n5788_17(.douta(w_n5788_17[0]),.doutb(w_n5788_17[1]),.doutc(w_n5788_17[2]),.din(w_n5788_5[1]));
	jspl3 jspl3_w_n5788_18(.douta(w_n5788_18[0]),.doutb(w_n5788_18[1]),.doutc(w_n5788_18[2]),.din(w_n5788_5[2]));
	jspl3 jspl3_w_n5788_19(.douta(w_n5788_19[0]),.doutb(w_n5788_19[1]),.doutc(w_n5788_19[2]),.din(w_n5788_6[0]));
	jspl3 jspl3_w_n5788_20(.douta(w_n5788_20[0]),.doutb(w_n5788_20[1]),.doutc(w_n5788_20[2]),.din(w_n5788_6[1]));
	jspl3 jspl3_w_n5793_0(.douta(w_n5793_0[0]),.doutb(w_n5793_0[1]),.doutc(w_n5793_0[2]),.din(n5793));
	jspl3 jspl3_w_n5793_1(.douta(w_n5793_1[0]),.doutb(w_n5793_1[1]),.doutc(w_n5793_1[2]),.din(w_n5793_0[0]));
	jspl3 jspl3_w_n5793_2(.douta(w_n5793_2[0]),.doutb(w_n5793_2[1]),.doutc(w_n5793_2[2]),.din(w_n5793_0[1]));
	jspl3 jspl3_w_n5793_3(.douta(w_n5793_3[0]),.doutb(w_n5793_3[1]),.doutc(w_n5793_3[2]),.din(w_n5793_0[2]));
	jspl3 jspl3_w_n5793_4(.douta(w_n5793_4[0]),.doutb(w_n5793_4[1]),.doutc(w_n5793_4[2]),.din(w_n5793_1[0]));
	jspl3 jspl3_w_n5793_5(.douta(w_n5793_5[0]),.doutb(w_n5793_5[1]),.doutc(w_n5793_5[2]),.din(w_n5793_1[1]));
	jspl3 jspl3_w_n5793_6(.douta(w_n5793_6[0]),.doutb(w_n5793_6[1]),.doutc(w_n5793_6[2]),.din(w_n5793_1[2]));
	jspl3 jspl3_w_n5793_7(.douta(w_n5793_7[0]),.doutb(w_n5793_7[1]),.doutc(w_n5793_7[2]),.din(w_n5793_2[0]));
	jspl3 jspl3_w_n5793_8(.douta(w_n5793_8[0]),.doutb(w_n5793_8[1]),.doutc(w_n5793_8[2]),.din(w_n5793_2[1]));
	jspl3 jspl3_w_n5793_9(.douta(w_n5793_9[0]),.doutb(w_n5793_9[1]),.doutc(w_n5793_9[2]),.din(w_n5793_2[2]));
	jspl3 jspl3_w_n5793_10(.douta(w_n5793_10[0]),.doutb(w_n5793_10[1]),.doutc(w_n5793_10[2]),.din(w_n5793_3[0]));
	jspl3 jspl3_w_n5793_11(.douta(w_n5793_11[0]),.doutb(w_n5793_11[1]),.doutc(w_n5793_11[2]),.din(w_n5793_3[1]));
	jspl3 jspl3_w_n5793_12(.douta(w_n5793_12[0]),.doutb(w_n5793_12[1]),.doutc(w_n5793_12[2]),.din(w_n5793_3[2]));
	jspl3 jspl3_w_n5793_13(.douta(w_n5793_13[0]),.doutb(w_n5793_13[1]),.doutc(w_n5793_13[2]),.din(w_n5793_4[0]));
	jspl3 jspl3_w_n5793_14(.douta(w_n5793_14[0]),.doutb(w_n5793_14[1]),.doutc(w_n5793_14[2]),.din(w_n5793_4[1]));
	jspl3 jspl3_w_n5793_15(.douta(w_n5793_15[0]),.doutb(w_n5793_15[1]),.doutc(w_n5793_15[2]),.din(w_n5793_4[2]));
	jspl3 jspl3_w_n5793_16(.douta(w_n5793_16[0]),.doutb(w_n5793_16[1]),.doutc(w_n5793_16[2]),.din(w_n5793_5[0]));
	jspl3 jspl3_w_n5793_17(.douta(w_n5793_17[0]),.doutb(w_n5793_17[1]),.doutc(w_n5793_17[2]),.din(w_n5793_5[1]));
	jspl3 jspl3_w_n5793_18(.douta(w_n5793_18[0]),.doutb(w_n5793_18[1]),.doutc(w_n5793_18[2]),.din(w_n5793_5[2]));
	jspl3 jspl3_w_n5793_19(.douta(w_n5793_19[0]),.doutb(w_n5793_19[1]),.doutc(w_n5793_19[2]),.din(w_n5793_6[0]));
	jspl3 jspl3_w_n5793_20(.douta(w_n5793_20[0]),.doutb(w_n5793_20[1]),.doutc(w_n5793_20[2]),.din(w_n5793_6[1]));
	jspl3 jspl3_w_n5793_21(.douta(w_n5793_21[0]),.doutb(w_n5793_21[1]),.doutc(w_n5793_21[2]),.din(w_n5793_6[2]));
	jspl3 jspl3_w_n5793_22(.douta(w_n5793_22[0]),.doutb(w_n5793_22[1]),.doutc(w_n5793_22[2]),.din(w_n5793_7[0]));
	jspl3 jspl3_w_n5793_23(.douta(w_n5793_23[0]),.doutb(w_n5793_23[1]),.doutc(w_n5793_23[2]),.din(w_n5793_7[1]));
	jspl3 jspl3_w_n5793_24(.douta(w_n5793_24[0]),.doutb(w_n5793_24[1]),.doutc(w_n5793_24[2]),.din(w_n5793_7[2]));
	jspl3 jspl3_w_n5793_25(.douta(w_n5793_25[0]),.doutb(w_n5793_25[1]),.doutc(w_n5793_25[2]),.din(w_n5793_8[0]));
	jspl3 jspl3_w_n5793_26(.douta(w_n5793_26[0]),.doutb(w_n5793_26[1]),.doutc(w_n5793_26[2]),.din(w_n5793_8[1]));
	jspl3 jspl3_w_n5793_27(.douta(w_n5793_27[0]),.doutb(w_n5793_27[1]),.doutc(w_n5793_27[2]),.din(w_n5793_8[2]));
	jspl3 jspl3_w_n5793_28(.douta(w_n5793_28[0]),.doutb(w_n5793_28[1]),.doutc(w_n5793_28[2]),.din(w_n5793_9[0]));
	jspl3 jspl3_w_n5793_29(.douta(w_n5793_29[0]),.doutb(w_n5793_29[1]),.doutc(w_n5793_29[2]),.din(w_n5793_9[1]));
	jspl jspl_w_n5794_0(.douta(w_n5794_0[0]),.doutb(w_n5794_0[1]),.din(n5794));
	jspl jspl_w_n5795_0(.douta(w_n5795_0[0]),.doutb(w_n5795_0[1]),.din(n5795));
	jspl3 jspl3_w_n5797_0(.douta(w_n5797_0[0]),.doutb(w_n5797_0[1]),.doutc(w_n5797_0[2]),.din(n5797));
	jspl jspl_w_n5797_1(.douta(w_n5797_1[0]),.doutb(w_n5797_1[1]),.din(w_n5797_0[0]));
	jspl3 jspl3_w_n5798_0(.douta(w_n5798_0[0]),.doutb(w_n5798_0[1]),.doutc(w_n5798_0[2]),.din(n5798));
	jspl3 jspl3_w_n5802_0(.douta(w_n5802_0[0]),.doutb(w_n5802_0[1]),.doutc(w_n5802_0[2]),.din(n5802));
	jspl jspl_w_n5803_0(.douta(w_n5803_0[0]),.doutb(w_n5803_0[1]),.din(n5803));
	jspl jspl_w_n5805_0(.douta(w_n5805_0[0]),.doutb(w_n5805_0[1]),.din(n5805));
	jspl jspl_w_n5807_0(.douta(w_n5807_0[0]),.doutb(w_n5807_0[1]),.din(n5807));
	jspl jspl_w_n5810_0(.douta(w_n5810_0[0]),.doutb(w_n5810_0[1]),.din(n5810));
	jspl jspl_w_n5815_0(.douta(w_n5815_0[0]),.doutb(w_n5815_0[1]),.din(n5815));
	jspl jspl_w_n5817_0(.douta(w_n5817_0[0]),.doutb(w_n5817_0[1]),.din(n5817));
	jspl jspl_w_n5818_0(.douta(w_n5818_0[0]),.doutb(w_n5818_0[1]),.din(n5818));
	jspl3 jspl3_w_n5819_0(.douta(w_n5819_0[0]),.doutb(w_n5819_0[1]),.doutc(w_n5819_0[2]),.din(n5819));
	jspl jspl_w_n5820_0(.douta(w_n5820_0[0]),.doutb(w_n5820_0[1]),.din(n5820));
	jspl jspl_w_n5824_0(.douta(w_n5824_0[0]),.doutb(w_n5824_0[1]),.din(n5824));
	jspl jspl_w_n5825_0(.douta(w_n5825_0[0]),.doutb(w_n5825_0[1]),.din(n5825));
	jspl jspl_w_n5827_0(.douta(w_n5827_0[0]),.doutb(w_n5827_0[1]),.din(n5827));
	jspl jspl_w_n5831_0(.douta(w_n5831_0[0]),.doutb(w_n5831_0[1]),.din(n5831));
	jspl jspl_w_n5833_0(.douta(w_n5833_0[0]),.doutb(w_n5833_0[1]),.din(n5833));
	jspl jspl_w_n5834_0(.douta(w_n5834_0[0]),.doutb(w_n5834_0[1]),.din(n5834));
	jspl3 jspl3_w_n5835_0(.douta(w_n5835_0[0]),.doutb(w_n5835_0[1]),.doutc(w_n5835_0[2]),.din(n5835));
	jspl jspl_w_n5836_0(.douta(w_n5836_0[0]),.doutb(w_n5836_0[1]),.din(n5836));
	jspl jspl_w_n5840_0(.douta(w_n5840_0[0]),.doutb(w_n5840_0[1]),.din(n5840));
	jspl jspl_w_n5842_0(.douta(w_n5842_0[0]),.doutb(w_n5842_0[1]),.din(n5842));
	jspl jspl_w_n5844_0(.douta(w_n5844_0[0]),.doutb(w_n5844_0[1]),.din(n5844));
	jspl jspl_w_n5846_0(.douta(w_n5846_0[0]),.doutb(w_n5846_0[1]),.din(n5846));
	jspl jspl_w_n5849_0(.douta(w_n5849_0[0]),.doutb(w_n5849_0[1]),.din(n5849));
	jspl jspl_w_n5855_0(.douta(w_n5855_0[0]),.doutb(w_n5855_0[1]),.din(n5855));
	jspl3 jspl3_w_n5857_0(.douta(w_n5857_0[0]),.doutb(w_n5857_0[1]),.doutc(w_n5857_0[2]),.din(n5857));
	jspl jspl_w_n5858_0(.douta(w_n5858_0[0]),.doutb(w_n5858_0[1]),.din(n5858));
	jspl jspl_w_n5863_0(.douta(w_n5863_0[0]),.doutb(w_n5863_0[1]),.din(n5863));
	jspl jspl_w_n5865_0(.douta(w_n5865_0[0]),.doutb(w_n5865_0[1]),.din(n5865));
	jspl jspl_w_n5867_0(.douta(w_n5867_0[0]),.doutb(w_n5867_0[1]),.din(n5867));
	jspl jspl_w_n5871_0(.douta(w_n5871_0[0]),.doutb(w_n5871_0[1]),.din(n5871));
	jspl jspl_w_n5873_0(.douta(w_n5873_0[0]),.doutb(w_n5873_0[1]),.din(n5873));
	jspl jspl_w_n5874_0(.douta(w_n5874_0[0]),.doutb(w_n5874_0[1]),.din(n5874));
	jspl3 jspl3_w_n5875_0(.douta(w_n5875_0[0]),.doutb(w_n5875_0[1]),.doutc(w_n5875_0[2]),.din(n5875));
	jspl jspl_w_n5876_0(.douta(w_n5876_0[0]),.doutb(w_n5876_0[1]),.din(n5876));
	jspl jspl_w_n5882_0(.douta(w_n5882_0[0]),.doutb(w_n5882_0[1]),.din(n5882));
	jspl jspl_w_n5883_0(.douta(w_n5883_0[0]),.doutb(w_n5883_0[1]),.din(n5883));
	jspl jspl_w_n5885_0(.douta(w_n5885_0[0]),.doutb(w_n5885_0[1]),.din(n5885));
	jspl jspl_w_n5887_0(.douta(w_n5887_0[0]),.doutb(w_n5887_0[1]),.din(n5887));
	jspl jspl_w_n5889_0(.douta(w_n5889_0[0]),.doutb(w_n5889_0[1]),.din(n5889));
	jspl jspl_w_n5895_0(.douta(w_n5895_0[0]),.doutb(w_n5895_0[1]),.din(n5895));
	jspl jspl_w_n5897_0(.douta(w_n5897_0[0]),.doutb(w_n5897_0[1]),.din(n5897));
	jspl3 jspl3_w_n5898_0(.douta(w_n5898_0[0]),.doutb(w_n5898_0[1]),.doutc(w_n5898_0[2]),.din(n5898));
	jspl jspl_w_n5901_0(.douta(w_n5901_0[0]),.doutb(w_n5901_0[1]),.din(n5901));
	jspl jspl_w_n5902_0(.douta(w_n5902_0[0]),.doutb(w_n5902_0[1]),.din(n5902));
	jspl3 jspl3_w_n5903_0(.douta(w_n5903_0[0]),.doutb(w_n5903_0[1]),.doutc(w_n5903_0[2]),.din(n5903));
	jspl jspl_w_n5905_0(.douta(w_n5905_0[0]),.doutb(w_n5905_0[1]),.din(n5905));
	jspl jspl_w_n5909_0(.douta(w_n5909_0[0]),.doutb(w_n5909_0[1]),.din(n5909));
	jspl jspl_w_n5911_0(.douta(w_n5911_0[0]),.doutb(w_n5911_0[1]),.din(n5911));
	jspl jspl_w_n5912_0(.douta(w_n5912_0[0]),.doutb(w_n5912_0[1]),.din(n5912));
	jspl3 jspl3_w_n5913_0(.douta(w_n5913_0[0]),.doutb(w_n5913_0[1]),.doutc(w_n5913_0[2]),.din(n5913));
	jspl jspl_w_n5914_0(.douta(w_n5914_0[0]),.doutb(w_n5914_0[1]),.din(n5914));
	jspl jspl_w_n5917_0(.douta(w_n5917_0[0]),.doutb(w_n5917_0[1]),.din(n5917));
	jspl jspl_w_n5923_0(.douta(w_n5923_0[0]),.doutb(w_n5923_0[1]),.din(n5923));
	jspl jspl_w_n5924_0(.douta(w_n5924_0[0]),.doutb(w_n5924_0[1]),.din(n5924));
	jspl jspl_w_n5926_0(.douta(w_n5926_0[0]),.doutb(w_n5926_0[1]),.din(n5926));
	jspl jspl_w_n5928_0(.douta(w_n5928_0[0]),.doutb(w_n5928_0[1]),.din(n5928));
	jspl jspl_w_n5930_0(.douta(w_n5930_0[0]),.doutb(w_n5930_0[1]),.din(n5930));
	jspl jspl_w_n5936_0(.douta(w_n5936_0[0]),.doutb(w_n5936_0[1]),.din(n5936));
	jspl jspl_w_n5938_0(.douta(w_n5938_0[0]),.doutb(w_n5938_0[1]),.din(n5938));
	jspl3 jspl3_w_n5939_0(.douta(w_n5939_0[0]),.doutb(w_n5939_0[1]),.doutc(w_n5939_0[2]),.din(n5939));
	jspl jspl_w_n5942_0(.douta(w_n5942_0[0]),.doutb(w_n5942_0[1]),.din(n5942));
	jspl jspl_w_n5943_0(.douta(w_n5943_0[0]),.doutb(w_n5943_0[1]),.din(n5943));
	jspl3 jspl3_w_n5944_0(.douta(w_n5944_0[0]),.doutb(w_n5944_0[1]),.doutc(w_n5944_0[2]),.din(n5944));
	jspl jspl_w_n5946_0(.douta(w_n5946_0[0]),.doutb(w_n5946_0[1]),.din(n5946));
	jspl jspl_w_n5950_0(.douta(w_n5950_0[0]),.doutb(w_n5950_0[1]),.din(n5950));
	jspl jspl_w_n5952_0(.douta(w_n5952_0[0]),.doutb(w_n5952_0[1]),.din(n5952));
	jspl jspl_w_n5953_0(.douta(w_n5953_0[0]),.doutb(w_n5953_0[1]),.din(n5953));
	jspl3 jspl3_w_n5954_0(.douta(w_n5954_0[0]),.doutb(w_n5954_0[1]),.doutc(w_n5954_0[2]),.din(n5954));
	jspl jspl_w_n5955_0(.douta(w_n5955_0[0]),.doutb(w_n5955_0[1]),.din(n5955));
	jspl jspl_w_n5958_0(.douta(w_n5958_0[0]),.doutb(w_n5958_0[1]),.din(n5958));
	jspl jspl_w_n5964_0(.douta(w_n5964_0[0]),.doutb(w_n5964_0[1]),.din(n5964));
	jspl jspl_w_n5965_0(.douta(w_n5965_0[0]),.doutb(w_n5965_0[1]),.din(n5965));
	jspl jspl_w_n5967_0(.douta(w_n5967_0[0]),.doutb(w_n5967_0[1]),.din(n5967));
	jspl jspl_w_n5969_0(.douta(w_n5969_0[0]),.doutb(w_n5969_0[1]),.din(n5969));
	jspl jspl_w_n5971_0(.douta(w_n5971_0[0]),.doutb(w_n5971_0[1]),.din(n5971));
	jspl jspl_w_n5977_0(.douta(w_n5977_0[0]),.doutb(w_n5977_0[1]),.din(n5977));
	jspl jspl_w_n5979_0(.douta(w_n5979_0[0]),.doutb(w_n5979_0[1]),.din(n5979));
	jspl3 jspl3_w_n5980_0(.douta(w_n5980_0[0]),.doutb(w_n5980_0[1]),.doutc(w_n5980_0[2]),.din(n5980));
	jspl jspl_w_n5983_0(.douta(w_n5983_0[0]),.doutb(w_n5983_0[1]),.din(n5983));
	jspl jspl_w_n5984_0(.douta(w_n5984_0[0]),.doutb(w_n5984_0[1]),.din(n5984));
	jspl3 jspl3_w_n5985_0(.douta(w_n5985_0[0]),.doutb(w_n5985_0[1]),.doutc(w_n5985_0[2]),.din(n5985));
	jspl jspl_w_n5987_0(.douta(w_n5987_0[0]),.doutb(w_n5987_0[1]),.din(n5987));
	jspl jspl_w_n5991_0(.douta(w_n5991_0[0]),.doutb(w_n5991_0[1]),.din(n5991));
	jspl jspl_w_n5993_0(.douta(w_n5993_0[0]),.doutb(w_n5993_0[1]),.din(n5993));
	jspl jspl_w_n5994_0(.douta(w_n5994_0[0]),.doutb(w_n5994_0[1]),.din(n5994));
	jspl3 jspl3_w_n5995_0(.douta(w_n5995_0[0]),.doutb(w_n5995_0[1]),.doutc(w_n5995_0[2]),.din(n5995));
	jspl jspl_w_n5996_0(.douta(w_n5996_0[0]),.doutb(w_n5996_0[1]),.din(n5996));
	jspl jspl_w_n5999_0(.douta(w_n5999_0[0]),.doutb(w_n5999_0[1]),.din(n5999));
	jspl jspl_w_n6005_0(.douta(w_n6005_0[0]),.doutb(w_n6005_0[1]),.din(n6005));
	jspl jspl_w_n6006_0(.douta(w_n6006_0[0]),.doutb(w_n6006_0[1]),.din(n6006));
	jspl jspl_w_n6008_0(.douta(w_n6008_0[0]),.doutb(w_n6008_0[1]),.din(n6008));
	jspl jspl_w_n6010_0(.douta(w_n6010_0[0]),.doutb(w_n6010_0[1]),.din(n6010));
	jspl jspl_w_n6012_0(.douta(w_n6012_0[0]),.doutb(w_n6012_0[1]),.din(n6012));
	jspl jspl_w_n6018_0(.douta(w_n6018_0[0]),.doutb(w_n6018_0[1]),.din(n6018));
	jspl jspl_w_n6020_0(.douta(w_n6020_0[0]),.doutb(w_n6020_0[1]),.din(n6020));
	jspl3 jspl3_w_n6021_0(.douta(w_n6021_0[0]),.doutb(w_n6021_0[1]),.doutc(w_n6021_0[2]),.din(n6021));
	jspl jspl_w_n6024_0(.douta(w_n6024_0[0]),.doutb(w_n6024_0[1]),.din(n6024));
	jspl jspl_w_n6025_0(.douta(w_n6025_0[0]),.doutb(w_n6025_0[1]),.din(n6025));
	jspl3 jspl3_w_n6026_0(.douta(w_n6026_0[0]),.doutb(w_n6026_0[1]),.doutc(w_n6026_0[2]),.din(n6026));
	jspl jspl_w_n6028_0(.douta(w_n6028_0[0]),.doutb(w_n6028_0[1]),.din(n6028));
	jspl jspl_w_n6032_0(.douta(w_n6032_0[0]),.doutb(w_n6032_0[1]),.din(n6032));
	jspl jspl_w_n6034_0(.douta(w_n6034_0[0]),.doutb(w_n6034_0[1]),.din(n6034));
	jspl jspl_w_n6035_0(.douta(w_n6035_0[0]),.doutb(w_n6035_0[1]),.din(n6035));
	jspl3 jspl3_w_n6036_0(.douta(w_n6036_0[0]),.doutb(w_n6036_0[1]),.doutc(w_n6036_0[2]),.din(n6036));
	jspl jspl_w_n6037_0(.douta(w_n6037_0[0]),.doutb(w_n6037_0[1]),.din(n6037));
	jspl jspl_w_n6040_0(.douta(w_n6040_0[0]),.doutb(w_n6040_0[1]),.din(n6040));
	jspl jspl_w_n6046_0(.douta(w_n6046_0[0]),.doutb(w_n6046_0[1]),.din(n6046));
	jspl jspl_w_n6047_0(.douta(w_n6047_0[0]),.doutb(w_n6047_0[1]),.din(n6047));
	jspl jspl_w_n6049_0(.douta(w_n6049_0[0]),.doutb(w_n6049_0[1]),.din(n6049));
	jspl jspl_w_n6051_0(.douta(w_n6051_0[0]),.doutb(w_n6051_0[1]),.din(n6051));
	jspl jspl_w_n6053_0(.douta(w_n6053_0[0]),.doutb(w_n6053_0[1]),.din(n6053));
	jspl jspl_w_n6059_0(.douta(w_n6059_0[0]),.doutb(w_n6059_0[1]),.din(n6059));
	jspl jspl_w_n6061_0(.douta(w_n6061_0[0]),.doutb(w_n6061_0[1]),.din(n6061));
	jspl3 jspl3_w_n6062_0(.douta(w_n6062_0[0]),.doutb(w_n6062_0[1]),.doutc(w_n6062_0[2]),.din(n6062));
	jspl jspl_w_n6065_0(.douta(w_n6065_0[0]),.doutb(w_n6065_0[1]),.din(n6065));
	jspl jspl_w_n6066_0(.douta(w_n6066_0[0]),.doutb(w_n6066_0[1]),.din(n6066));
	jspl3 jspl3_w_n6067_0(.douta(w_n6067_0[0]),.doutb(w_n6067_0[1]),.doutc(w_n6067_0[2]),.din(n6067));
	jspl jspl_w_n6069_0(.douta(w_n6069_0[0]),.doutb(w_n6069_0[1]),.din(n6069));
	jspl jspl_w_n6073_0(.douta(w_n6073_0[0]),.doutb(w_n6073_0[1]),.din(n6073));
	jspl jspl_w_n6075_0(.douta(w_n6075_0[0]),.doutb(w_n6075_0[1]),.din(n6075));
	jspl jspl_w_n6076_0(.douta(w_n6076_0[0]),.doutb(w_n6076_0[1]),.din(n6076));
	jspl3 jspl3_w_n6077_0(.douta(w_n6077_0[0]),.doutb(w_n6077_0[1]),.doutc(w_n6077_0[2]),.din(n6077));
	jspl jspl_w_n6078_0(.douta(w_n6078_0[0]),.doutb(w_n6078_0[1]),.din(n6078));
	jspl jspl_w_n6081_0(.douta(w_n6081_0[0]),.doutb(w_n6081_0[1]),.din(n6081));
	jspl jspl_w_n6087_0(.douta(w_n6087_0[0]),.doutb(w_n6087_0[1]),.din(n6087));
	jspl jspl_w_n6088_0(.douta(w_n6088_0[0]),.doutb(w_n6088_0[1]),.din(n6088));
	jspl jspl_w_n6090_0(.douta(w_n6090_0[0]),.doutb(w_n6090_0[1]),.din(n6090));
	jspl jspl_w_n6092_0(.douta(w_n6092_0[0]),.doutb(w_n6092_0[1]),.din(n6092));
	jspl jspl_w_n6094_0(.douta(w_n6094_0[0]),.doutb(w_n6094_0[1]),.din(n6094));
	jspl jspl_w_n6100_0(.douta(w_n6100_0[0]),.doutb(w_n6100_0[1]),.din(n6100));
	jspl3 jspl3_w_n6102_0(.douta(w_n6102_0[0]),.doutb(w_n6102_0[1]),.doutc(w_n6102_0[2]),.din(n6102));
	jspl jspl_w_n6107_0(.douta(w_n6107_0[0]),.doutb(w_n6107_0[1]),.din(n6107));
	jspl3 jspl3_w_n6109_0(.douta(w_n6109_0[0]),.doutb(w_n6109_0[1]),.doutc(w_n6109_0[2]),.din(n6109));
	jspl3 jspl3_w_n6113_0(.douta(w_n6113_0[0]),.doutb(w_n6113_0[1]),.doutc(w_n6113_0[2]),.din(n6113));
	jspl jspl_w_n6114_0(.douta(w_n6114_0[0]),.doutb(w_n6114_0[1]),.din(n6114));
	jspl jspl_w_n6119_0(.douta(w_n6119_0[0]),.doutb(w_n6119_0[1]),.din(n6119));
	jspl3 jspl3_w_n6120_0(.douta(w_n6120_0[0]),.doutb(w_n6120_0[1]),.doutc(w_n6120_0[2]),.din(n6120));
	jspl jspl_w_n6125_0(.douta(w_n6125_0[0]),.doutb(w_n6125_0[1]),.din(n6125));
	jspl jspl_w_n6132_0(.douta(w_n6132_0[0]),.doutb(w_n6132_0[1]),.din(n6132));
	jspl3 jspl3_w_n6134_0(.douta(w_n6134_0[0]),.doutb(w_n6134_0[1]),.doutc(w_n6134_0[2]),.din(n6134));
	jspl jspl_w_n6134_1(.douta(w_n6134_1[0]),.doutb(w_n6134_1[1]),.din(w_n6134_0[0]));
	jspl jspl_w_n6135_0(.douta(w_n6135_0[0]),.doutb(w_n6135_0[1]),.din(n6135));
	jspl3 jspl3_w_n6138_0(.douta(w_n6138_0[0]),.doutb(w_n6138_0[1]),.doutc(w_n6138_0[2]),.din(n6138));
	jspl jspl_w_n6139_0(.douta(w_n6139_0[0]),.doutb(w_n6139_0[1]),.din(n6139));
	jspl jspl_w_n6140_0(.douta(w_n6140_0[0]),.doutb(w_n6140_0[1]),.din(n6140));
	jspl jspl_w_n6141_0(.douta(w_n6141_0[0]),.doutb(w_n6141_0[1]),.din(n6141));
	jspl jspl_w_n6143_0(.douta(w_n6143_0[0]),.doutb(w_n6143_0[1]),.din(n6143));
	jspl jspl_w_n6145_0(.douta(w_n6145_0[0]),.doutb(w_n6145_0[1]),.din(n6145));
	jspl jspl_w_n6154_0(.douta(w_n6154_0[0]),.doutb(w_n6154_0[1]),.din(n6154));
	jspl jspl_w_n6156_0(.douta(w_n6156_0[0]),.doutb(w_n6156_0[1]),.din(n6156));
	jspl jspl_w_n6157_0(.douta(w_n6157_0[0]),.doutb(w_n6157_0[1]),.din(n6157));
	jspl3 jspl3_w_n6158_0(.douta(w_n6158_0[0]),.doutb(w_n6158_0[1]),.doutc(w_n6158_0[2]),.din(n6158));
	jspl jspl_w_n6159_0(.douta(w_n6159_0[0]),.doutb(w_n6159_0[1]),.din(n6159));
	jspl jspl_w_n6162_0(.douta(w_n6162_0[0]),.doutb(w_n6162_0[1]),.din(n6162));
	jspl jspl_w_n6164_0(.douta(w_n6164_0[0]),.doutb(w_n6164_0[1]),.din(n6164));
	jspl jspl_w_n6166_0(.douta(w_n6166_0[0]),.doutb(w_n6166_0[1]),.din(n6166));
	jspl jspl_w_n6169_0(.douta(w_n6169_0[0]),.doutb(w_n6169_0[1]),.din(n6169));
	jspl jspl_w_n6175_0(.douta(w_n6175_0[0]),.doutb(w_n6175_0[1]),.din(n6175));
	jspl3 jspl3_w_n6177_0(.douta(w_n6177_0[0]),.doutb(w_n6177_0[1]),.doutc(w_n6177_0[2]),.din(n6177));
	jspl jspl_w_n6178_0(.douta(w_n6178_0[0]),.doutb(w_n6178_0[1]),.din(n6178));
	jspl jspl_w_n6183_0(.douta(w_n6183_0[0]),.doutb(w_n6183_0[1]),.din(n6183));
	jspl jspl_w_n6184_0(.douta(w_n6184_0[0]),.doutb(w_n6184_0[1]),.din(n6184));
	jspl jspl_w_n6186_0(.douta(w_n6186_0[0]),.doutb(w_n6186_0[1]),.din(n6186));
	jspl jspl_w_n6188_0(.douta(w_n6188_0[0]),.doutb(w_n6188_0[1]),.din(n6188));
	jspl jspl_w_n6191_0(.douta(w_n6191_0[0]),.doutb(w_n6191_0[1]),.din(n6191));
	jspl jspl_w_n6197_0(.douta(w_n6197_0[0]),.doutb(w_n6197_0[1]),.din(n6197));
	jspl3 jspl3_w_n6199_0(.douta(w_n6199_0[0]),.doutb(w_n6199_0[1]),.doutc(w_n6199_0[2]),.din(n6199));
	jspl jspl_w_n6200_0(.douta(w_n6200_0[0]),.doutb(w_n6200_0[1]),.din(n6200));
	jspl jspl_w_n6204_0(.douta(w_n6204_0[0]),.doutb(w_n6204_0[1]),.din(n6204));
	jspl jspl_w_n6205_0(.douta(w_n6205_0[0]),.doutb(w_n6205_0[1]),.din(n6205));
	jspl jspl_w_n6207_0(.douta(w_n6207_0[0]),.doutb(w_n6207_0[1]),.din(n6207));
	jspl jspl_w_n6212_0(.douta(w_n6212_0[0]),.doutb(w_n6212_0[1]),.din(n6212));
	jspl jspl_w_n6214_0(.douta(w_n6214_0[0]),.doutb(w_n6214_0[1]),.din(n6214));
	jspl jspl_w_n6215_0(.douta(w_n6215_0[0]),.doutb(w_n6215_0[1]),.din(n6215));
	jspl3 jspl3_w_n6216_0(.douta(w_n6216_0[0]),.doutb(w_n6216_0[1]),.doutc(w_n6216_0[2]),.din(n6216));
	jspl jspl_w_n6217_0(.douta(w_n6217_0[0]),.doutb(w_n6217_0[1]),.din(n6217));
	jspl jspl_w_n6221_0(.douta(w_n6221_0[0]),.doutb(w_n6221_0[1]),.din(n6221));
	jspl jspl_w_n6222_0(.douta(w_n6222_0[0]),.doutb(w_n6222_0[1]),.din(n6222));
	jspl jspl_w_n6224_0(.douta(w_n6224_0[0]),.doutb(w_n6224_0[1]),.din(n6224));
	jspl jspl_w_n6226_0(.douta(w_n6226_0[0]),.doutb(w_n6226_0[1]),.din(n6226));
	jspl jspl_w_n6229_0(.douta(w_n6229_0[0]),.doutb(w_n6229_0[1]),.din(n6229));
	jspl jspl_w_n6235_0(.douta(w_n6235_0[0]),.doutb(w_n6235_0[1]),.din(n6235));
	jspl jspl_w_n6237_0(.douta(w_n6237_0[0]),.doutb(w_n6237_0[1]),.din(n6237));
	jspl3 jspl3_w_n6238_0(.douta(w_n6238_0[0]),.doutb(w_n6238_0[1]),.doutc(w_n6238_0[2]),.din(n6238));
	jspl jspl_w_n6242_0(.douta(w_n6242_0[0]),.doutb(w_n6242_0[1]),.din(n6242));
	jspl jspl_w_n6243_0(.douta(w_n6243_0[0]),.doutb(w_n6243_0[1]),.din(n6243));
	jspl3 jspl3_w_n6244_0(.douta(w_n6244_0[0]),.doutb(w_n6244_0[1]),.doutc(w_n6244_0[2]),.din(n6244));
	jspl jspl_w_n6246_0(.douta(w_n6246_0[0]),.doutb(w_n6246_0[1]),.din(n6246));
	jspl jspl_w_n6251_0(.douta(w_n6251_0[0]),.doutb(w_n6251_0[1]),.din(n6251));
	jspl jspl_w_n6253_0(.douta(w_n6253_0[0]),.doutb(w_n6253_0[1]),.din(n6253));
	jspl jspl_w_n6254_0(.douta(w_n6254_0[0]),.doutb(w_n6254_0[1]),.din(n6254));
	jspl3 jspl3_w_n6255_0(.douta(w_n6255_0[0]),.doutb(w_n6255_0[1]),.doutc(w_n6255_0[2]),.din(n6255));
	jspl jspl_w_n6256_0(.douta(w_n6256_0[0]),.doutb(w_n6256_0[1]),.din(n6256));
	jspl jspl_w_n6260_0(.douta(w_n6260_0[0]),.doutb(w_n6260_0[1]),.din(n6260));
	jspl jspl_w_n6266_0(.douta(w_n6266_0[0]),.doutb(w_n6266_0[1]),.din(n6266));
	jspl jspl_w_n6267_0(.douta(w_n6267_0[0]),.doutb(w_n6267_0[1]),.din(n6267));
	jspl jspl_w_n6269_0(.douta(w_n6269_0[0]),.doutb(w_n6269_0[1]),.din(n6269));
	jspl jspl_w_n6271_0(.douta(w_n6271_0[0]),.doutb(w_n6271_0[1]),.din(n6271));
	jspl jspl_w_n6274_0(.douta(w_n6274_0[0]),.doutb(w_n6274_0[1]),.din(n6274));
	jspl jspl_w_n6280_0(.douta(w_n6280_0[0]),.doutb(w_n6280_0[1]),.din(n6280));
	jspl jspl_w_n6282_0(.douta(w_n6282_0[0]),.doutb(w_n6282_0[1]),.din(n6282));
	jspl3 jspl3_w_n6283_0(.douta(w_n6283_0[0]),.doutb(w_n6283_0[1]),.doutc(w_n6283_0[2]),.din(n6283));
	jspl jspl_w_n6287_0(.douta(w_n6287_0[0]),.doutb(w_n6287_0[1]),.din(n6287));
	jspl jspl_w_n6288_0(.douta(w_n6288_0[0]),.doutb(w_n6288_0[1]),.din(n6288));
	jspl3 jspl3_w_n6289_0(.douta(w_n6289_0[0]),.doutb(w_n6289_0[1]),.doutc(w_n6289_0[2]),.din(n6289));
	jspl jspl_w_n6291_0(.douta(w_n6291_0[0]),.doutb(w_n6291_0[1]),.din(n6291));
	jspl jspl_w_n6296_0(.douta(w_n6296_0[0]),.doutb(w_n6296_0[1]),.din(n6296));
	jspl jspl_w_n6298_0(.douta(w_n6298_0[0]),.doutb(w_n6298_0[1]),.din(n6298));
	jspl jspl_w_n6299_0(.douta(w_n6299_0[0]),.doutb(w_n6299_0[1]),.din(n6299));
	jspl3 jspl3_w_n6300_0(.douta(w_n6300_0[0]),.doutb(w_n6300_0[1]),.doutc(w_n6300_0[2]),.din(n6300));
	jspl jspl_w_n6301_0(.douta(w_n6301_0[0]),.doutb(w_n6301_0[1]),.din(n6301));
	jspl jspl_w_n6305_0(.douta(w_n6305_0[0]),.doutb(w_n6305_0[1]),.din(n6305));
	jspl jspl_w_n6311_0(.douta(w_n6311_0[0]),.doutb(w_n6311_0[1]),.din(n6311));
	jspl jspl_w_n6312_0(.douta(w_n6312_0[0]),.doutb(w_n6312_0[1]),.din(n6312));
	jspl jspl_w_n6314_0(.douta(w_n6314_0[0]),.doutb(w_n6314_0[1]),.din(n6314));
	jspl jspl_w_n6316_0(.douta(w_n6316_0[0]),.doutb(w_n6316_0[1]),.din(n6316));
	jspl jspl_w_n6319_0(.douta(w_n6319_0[0]),.doutb(w_n6319_0[1]),.din(n6319));
	jspl jspl_w_n6325_0(.douta(w_n6325_0[0]),.doutb(w_n6325_0[1]),.din(n6325));
	jspl jspl_w_n6327_0(.douta(w_n6327_0[0]),.doutb(w_n6327_0[1]),.din(n6327));
	jspl3 jspl3_w_n6328_0(.douta(w_n6328_0[0]),.doutb(w_n6328_0[1]),.doutc(w_n6328_0[2]),.din(n6328));
	jspl jspl_w_n6332_0(.douta(w_n6332_0[0]),.doutb(w_n6332_0[1]),.din(n6332));
	jspl jspl_w_n6333_0(.douta(w_n6333_0[0]),.doutb(w_n6333_0[1]),.din(n6333));
	jspl3 jspl3_w_n6334_0(.douta(w_n6334_0[0]),.doutb(w_n6334_0[1]),.doutc(w_n6334_0[2]),.din(n6334));
	jspl jspl_w_n6336_0(.douta(w_n6336_0[0]),.doutb(w_n6336_0[1]),.din(n6336));
	jspl jspl_w_n6341_0(.douta(w_n6341_0[0]),.doutb(w_n6341_0[1]),.din(n6341));
	jspl jspl_w_n6343_0(.douta(w_n6343_0[0]),.doutb(w_n6343_0[1]),.din(n6343));
	jspl jspl_w_n6344_0(.douta(w_n6344_0[0]),.doutb(w_n6344_0[1]),.din(n6344));
	jspl3 jspl3_w_n6345_0(.douta(w_n6345_0[0]),.doutb(w_n6345_0[1]),.doutc(w_n6345_0[2]),.din(n6345));
	jspl jspl_w_n6346_0(.douta(w_n6346_0[0]),.doutb(w_n6346_0[1]),.din(n6346));
	jspl jspl_w_n6350_0(.douta(w_n6350_0[0]),.doutb(w_n6350_0[1]),.din(n6350));
	jspl jspl_w_n6356_0(.douta(w_n6356_0[0]),.doutb(w_n6356_0[1]),.din(n6356));
	jspl jspl_w_n6357_0(.douta(w_n6357_0[0]),.doutb(w_n6357_0[1]),.din(n6357));
	jspl jspl_w_n6359_0(.douta(w_n6359_0[0]),.doutb(w_n6359_0[1]),.din(n6359));
	jspl jspl_w_n6361_0(.douta(w_n6361_0[0]),.doutb(w_n6361_0[1]),.din(n6361));
	jspl jspl_w_n6364_0(.douta(w_n6364_0[0]),.doutb(w_n6364_0[1]),.din(n6364));
	jspl jspl_w_n6370_0(.douta(w_n6370_0[0]),.doutb(w_n6370_0[1]),.din(n6370));
	jspl jspl_w_n6372_0(.douta(w_n6372_0[0]),.doutb(w_n6372_0[1]),.din(n6372));
	jspl3 jspl3_w_n6373_0(.douta(w_n6373_0[0]),.doutb(w_n6373_0[1]),.doutc(w_n6373_0[2]),.din(n6373));
	jspl jspl_w_n6377_0(.douta(w_n6377_0[0]),.doutb(w_n6377_0[1]),.din(n6377));
	jspl jspl_w_n6378_0(.douta(w_n6378_0[0]),.doutb(w_n6378_0[1]),.din(n6378));
	jspl3 jspl3_w_n6379_0(.douta(w_n6379_0[0]),.doutb(w_n6379_0[1]),.doutc(w_n6379_0[2]),.din(n6379));
	jspl jspl_w_n6381_0(.douta(w_n6381_0[0]),.doutb(w_n6381_0[1]),.din(n6381));
	jspl jspl_w_n6386_0(.douta(w_n6386_0[0]),.doutb(w_n6386_0[1]),.din(n6386));
	jspl jspl_w_n6388_0(.douta(w_n6388_0[0]),.doutb(w_n6388_0[1]),.din(n6388));
	jspl jspl_w_n6389_0(.douta(w_n6389_0[0]),.doutb(w_n6389_0[1]),.din(n6389));
	jspl3 jspl3_w_n6390_0(.douta(w_n6390_0[0]),.doutb(w_n6390_0[1]),.doutc(w_n6390_0[2]),.din(n6390));
	jspl jspl_w_n6391_0(.douta(w_n6391_0[0]),.doutb(w_n6391_0[1]),.din(n6391));
	jspl jspl_w_n6395_0(.douta(w_n6395_0[0]),.doutb(w_n6395_0[1]),.din(n6395));
	jspl jspl_w_n6401_0(.douta(w_n6401_0[0]),.doutb(w_n6401_0[1]),.din(n6401));
	jspl jspl_w_n6402_0(.douta(w_n6402_0[0]),.doutb(w_n6402_0[1]),.din(n6402));
	jspl jspl_w_n6404_0(.douta(w_n6404_0[0]),.doutb(w_n6404_0[1]),.din(n6404));
	jspl jspl_w_n6406_0(.douta(w_n6406_0[0]),.doutb(w_n6406_0[1]),.din(n6406));
	jspl jspl_w_n6409_0(.douta(w_n6409_0[0]),.doutb(w_n6409_0[1]),.din(n6409));
	jspl jspl_w_n6415_0(.douta(w_n6415_0[0]),.doutb(w_n6415_0[1]),.din(n6415));
	jspl jspl_w_n6417_0(.douta(w_n6417_0[0]),.doutb(w_n6417_0[1]),.din(n6417));
	jspl3 jspl3_w_n6418_0(.douta(w_n6418_0[0]),.doutb(w_n6418_0[1]),.doutc(w_n6418_0[2]),.din(n6418));
	jspl jspl_w_n6422_0(.douta(w_n6422_0[0]),.doutb(w_n6422_0[1]),.din(n6422));
	jspl jspl_w_n6423_0(.douta(w_n6423_0[0]),.doutb(w_n6423_0[1]),.din(n6423));
	jspl3 jspl3_w_n6424_0(.douta(w_n6424_0[0]),.doutb(w_n6424_0[1]),.doutc(w_n6424_0[2]),.din(n6424));
	jspl jspl_w_n6426_0(.douta(w_n6426_0[0]),.doutb(w_n6426_0[1]),.din(n6426));
	jspl jspl_w_n6431_0(.douta(w_n6431_0[0]),.doutb(w_n6431_0[1]),.din(n6431));
	jspl jspl_w_n6433_0(.douta(w_n6433_0[0]),.doutb(w_n6433_0[1]),.din(n6433));
	jspl jspl_w_n6434_0(.douta(w_n6434_0[0]),.doutb(w_n6434_0[1]),.din(n6434));
	jspl3 jspl3_w_n6435_0(.douta(w_n6435_0[0]),.doutb(w_n6435_0[1]),.doutc(w_n6435_0[2]),.din(n6435));
	jspl jspl_w_n6436_0(.douta(w_n6436_0[0]),.doutb(w_n6436_0[1]),.din(n6436));
	jspl jspl_w_n6440_0(.douta(w_n6440_0[0]),.doutb(w_n6440_0[1]),.din(n6440));
	jspl jspl_w_n6446_0(.douta(w_n6446_0[0]),.doutb(w_n6446_0[1]),.din(n6446));
	jspl jspl_w_n6447_0(.douta(w_n6447_0[0]),.doutb(w_n6447_0[1]),.din(n6447));
	jspl jspl_w_n6449_0(.douta(w_n6449_0[0]),.doutb(w_n6449_0[1]),.din(n6449));
	jspl jspl_w_n6451_0(.douta(w_n6451_0[0]),.doutb(w_n6451_0[1]),.din(n6451));
	jspl jspl_w_n6454_0(.douta(w_n6454_0[0]),.doutb(w_n6454_0[1]),.din(n6454));
	jspl jspl_w_n6460_0(.douta(w_n6460_0[0]),.doutb(w_n6460_0[1]),.din(n6460));
	jspl jspl_w_n6462_0(.douta(w_n6462_0[0]),.doutb(w_n6462_0[1]),.din(n6462));
	jspl3 jspl3_w_n6463_0(.douta(w_n6463_0[0]),.doutb(w_n6463_0[1]),.doutc(w_n6463_0[2]),.din(n6463));
	jspl jspl_w_n6467_0(.douta(w_n6467_0[0]),.doutb(w_n6467_0[1]),.din(n6467));
	jspl jspl_w_n6468_0(.douta(w_n6468_0[0]),.doutb(w_n6468_0[1]),.din(n6468));
	jspl3 jspl3_w_n6469_0(.douta(w_n6469_0[0]),.doutb(w_n6469_0[1]),.doutc(w_n6469_0[2]),.din(n6469));
	jspl jspl_w_n6471_0(.douta(w_n6471_0[0]),.doutb(w_n6471_0[1]),.din(n6471));
	jspl jspl_w_n6476_0(.douta(w_n6476_0[0]),.doutb(w_n6476_0[1]),.din(n6476));
	jspl jspl_w_n6478_0(.douta(w_n6478_0[0]),.doutb(w_n6478_0[1]),.din(n6478));
	jspl jspl_w_n6479_0(.douta(w_n6479_0[0]),.doutb(w_n6479_0[1]),.din(n6479));
	jspl3 jspl3_w_n6480_0(.douta(w_n6480_0[0]),.doutb(w_n6480_0[1]),.doutc(w_n6480_0[2]),.din(n6480));
	jspl3 jspl3_w_n6480_1(.douta(w_n6480_1[0]),.doutb(w_n6480_1[1]),.doutc(w_n6480_1[2]),.din(w_n6480_0[0]));
	jspl jspl_w_n6483_0(.douta(w_n6483_0[0]),.doutb(w_n6483_0[1]),.din(n6483));
	jspl3 jspl3_w_n6484_0(.douta(w_n6484_0[0]),.doutb(w_n6484_0[1]),.doutc(w_n6484_0[2]),.din(n6484));
	jspl jspl_w_n6485_0(.douta(w_n6485_0[0]),.doutb(w_n6485_0[1]),.din(n6485));
	jspl jspl_w_n6486_0(.douta(w_n6486_0[0]),.doutb(w_n6486_0[1]),.din(n6486));
	jspl jspl_w_n6492_0(.douta(w_n6492_0[0]),.doutb(w_n6492_0[1]),.din(n6492));
	jspl3 jspl3_w_n6493_0(.douta(w_n6493_0[0]),.doutb(w_n6493_0[1]),.doutc(w_n6493_0[2]),.din(n6493));
	jspl jspl_w_n6494_0(.douta(w_n6494_0[0]),.doutb(w_n6494_0[1]),.din(n6494));
	jspl jspl_w_n6499_0(.douta(w_n6499_0[0]),.doutb(w_n6499_0[1]),.din(n6499));
	jspl3 jspl3_w_n6500_0(.douta(w_n6500_0[0]),.doutb(w_n6500_0[1]),.doutc(w_n6500_0[2]),.din(n6500));
	jspl3 jspl3_w_n6500_1(.douta(w_n6500_1[0]),.doutb(w_n6500_1[1]),.doutc(w_n6500_1[2]),.din(w_n6500_0[0]));
	jspl3 jspl3_w_n6500_2(.douta(w_n6500_2[0]),.doutb(w_n6500_2[1]),.doutc(w_n6500_2[2]),.din(w_n6500_0[1]));
	jspl3 jspl3_w_n6500_3(.douta(w_n6500_3[0]),.doutb(w_n6500_3[1]),.doutc(w_n6500_3[2]),.din(w_n6500_0[2]));
	jspl3 jspl3_w_n6500_4(.douta(w_n6500_4[0]),.doutb(w_n6500_4[1]),.doutc(w_n6500_4[2]),.din(w_n6500_1[0]));
	jspl3 jspl3_w_n6500_5(.douta(w_n6500_5[0]),.doutb(w_n6500_5[1]),.doutc(w_n6500_5[2]),.din(w_n6500_1[1]));
	jspl3 jspl3_w_n6500_6(.douta(w_n6500_6[0]),.doutb(w_n6500_6[1]),.doutc(w_n6500_6[2]),.din(w_n6500_1[2]));
	jspl3 jspl3_w_n6500_7(.douta(w_n6500_7[0]),.doutb(w_n6500_7[1]),.doutc(w_n6500_7[2]),.din(w_n6500_2[0]));
	jspl3 jspl3_w_n6500_8(.douta(w_n6500_8[0]),.doutb(w_n6500_8[1]),.doutc(w_n6500_8[2]),.din(w_n6500_2[1]));
	jspl3 jspl3_w_n6500_9(.douta(w_n6500_9[0]),.doutb(w_n6500_9[1]),.doutc(w_n6500_9[2]),.din(w_n6500_2[2]));
	jspl3 jspl3_w_n6500_10(.douta(w_n6500_10[0]),.doutb(w_n6500_10[1]),.doutc(w_n6500_10[2]),.din(w_n6500_3[0]));
	jspl3 jspl3_w_n6500_11(.douta(w_n6500_11[0]),.doutb(w_n6500_11[1]),.doutc(w_n6500_11[2]),.din(w_n6500_3[1]));
	jspl3 jspl3_w_n6500_12(.douta(w_n6500_12[0]),.doutb(w_n6500_12[1]),.doutc(w_n6500_12[2]),.din(w_n6500_3[2]));
	jspl3 jspl3_w_n6500_13(.douta(w_n6500_13[0]),.doutb(w_n6500_13[1]),.doutc(w_n6500_13[2]),.din(w_n6500_4[0]));
	jspl3 jspl3_w_n6500_14(.douta(w_n6500_14[0]),.doutb(w_n6500_14[1]),.doutc(w_n6500_14[2]),.din(w_n6500_4[1]));
	jspl3 jspl3_w_n6500_15(.douta(w_n6500_15[0]),.doutb(w_n6500_15[1]),.doutc(w_n6500_15[2]),.din(w_n6500_4[2]));
	jspl3 jspl3_w_n6500_16(.douta(w_n6500_16[0]),.doutb(w_n6500_16[1]),.doutc(w_n6500_16[2]),.din(w_n6500_5[0]));
	jspl3 jspl3_w_n6500_17(.douta(w_n6500_17[0]),.doutb(w_n6500_17[1]),.doutc(w_n6500_17[2]),.din(w_n6500_5[1]));
	jspl3 jspl3_w_n6500_18(.douta(w_n6500_18[0]),.doutb(w_n6500_18[1]),.doutc(w_n6500_18[2]),.din(w_n6500_5[2]));
	jspl jspl_w_n6500_19(.douta(w_n6500_19[0]),.doutb(w_n6500_19[1]),.din(w_n6500_6[0]));
	jspl3 jspl3_w_n6505_0(.douta(w_n6505_0[0]),.doutb(w_n6505_0[1]),.doutc(w_n6505_0[2]),.din(n6505));
	jspl3 jspl3_w_n6505_1(.douta(w_n6505_1[0]),.doutb(w_n6505_1[1]),.doutc(w_n6505_1[2]),.din(w_n6505_0[0]));
	jspl3 jspl3_w_n6505_2(.douta(w_n6505_2[0]),.doutb(w_n6505_2[1]),.doutc(w_n6505_2[2]),.din(w_n6505_0[1]));
	jspl3 jspl3_w_n6505_3(.douta(w_n6505_3[0]),.doutb(w_n6505_3[1]),.doutc(w_n6505_3[2]),.din(w_n6505_0[2]));
	jspl3 jspl3_w_n6505_4(.douta(w_n6505_4[0]),.doutb(w_n6505_4[1]),.doutc(w_n6505_4[2]),.din(w_n6505_1[0]));
	jspl3 jspl3_w_n6505_5(.douta(w_n6505_5[0]),.doutb(w_n6505_5[1]),.doutc(w_n6505_5[2]),.din(w_n6505_1[1]));
	jspl3 jspl3_w_n6505_6(.douta(w_n6505_6[0]),.doutb(w_n6505_6[1]),.doutc(w_n6505_6[2]),.din(w_n6505_1[2]));
	jspl3 jspl3_w_n6505_7(.douta(w_n6505_7[0]),.doutb(w_n6505_7[1]),.doutc(w_n6505_7[2]),.din(w_n6505_2[0]));
	jspl3 jspl3_w_n6505_8(.douta(w_n6505_8[0]),.doutb(w_n6505_8[1]),.doutc(w_n6505_8[2]),.din(w_n6505_2[1]));
	jspl3 jspl3_w_n6505_9(.douta(w_n6505_9[0]),.doutb(w_n6505_9[1]),.doutc(w_n6505_9[2]),.din(w_n6505_2[2]));
	jspl3 jspl3_w_n6505_10(.douta(w_n6505_10[0]),.doutb(w_n6505_10[1]),.doutc(w_n6505_10[2]),.din(w_n6505_3[0]));
	jspl3 jspl3_w_n6505_11(.douta(w_n6505_11[0]),.doutb(w_n6505_11[1]),.doutc(w_n6505_11[2]),.din(w_n6505_3[1]));
	jspl3 jspl3_w_n6505_12(.douta(w_n6505_12[0]),.doutb(w_n6505_12[1]),.doutc(w_n6505_12[2]),.din(w_n6505_3[2]));
	jspl3 jspl3_w_n6505_13(.douta(w_n6505_13[0]),.doutb(w_n6505_13[1]),.doutc(w_n6505_13[2]),.din(w_n6505_4[0]));
	jspl3 jspl3_w_n6505_14(.douta(w_n6505_14[0]),.doutb(w_n6505_14[1]),.doutc(w_n6505_14[2]),.din(w_n6505_4[1]));
	jspl3 jspl3_w_n6505_15(.douta(w_n6505_15[0]),.doutb(w_n6505_15[1]),.doutc(w_n6505_15[2]),.din(w_n6505_4[2]));
	jspl3 jspl3_w_n6505_16(.douta(w_n6505_16[0]),.doutb(w_n6505_16[1]),.doutc(w_n6505_16[2]),.din(w_n6505_5[0]));
	jspl3 jspl3_w_n6505_17(.douta(w_n6505_17[0]),.doutb(w_n6505_17[1]),.doutc(w_n6505_17[2]),.din(w_n6505_5[1]));
	jspl3 jspl3_w_n6505_18(.douta(w_n6505_18[0]),.doutb(w_n6505_18[1]),.doutc(w_n6505_18[2]),.din(w_n6505_5[2]));
	jspl3 jspl3_w_n6505_19(.douta(w_n6505_19[0]),.doutb(w_n6505_19[1]),.doutc(w_n6505_19[2]),.din(w_n6505_6[0]));
	jspl3 jspl3_w_n6505_20(.douta(w_n6505_20[0]),.doutb(w_n6505_20[1]),.doutc(w_n6505_20[2]),.din(w_n6505_6[1]));
	jspl3 jspl3_w_n6505_21(.douta(w_n6505_21[0]),.doutb(w_n6505_21[1]),.doutc(w_n6505_21[2]),.din(w_n6505_6[2]));
	jspl3 jspl3_w_n6505_22(.douta(w_n6505_22[0]),.doutb(w_n6505_22[1]),.doutc(w_n6505_22[2]),.din(w_n6505_7[0]));
	jspl3 jspl3_w_n6505_23(.douta(w_n6505_23[0]),.doutb(w_n6505_23[1]),.doutc(w_n6505_23[2]),.din(w_n6505_7[1]));
	jspl3 jspl3_w_n6505_24(.douta(w_n6505_24[0]),.doutb(w_n6505_24[1]),.doutc(w_n6505_24[2]),.din(w_n6505_7[2]));
	jspl3 jspl3_w_n6505_25(.douta(w_n6505_25[0]),.doutb(w_n6505_25[1]),.doutc(w_n6505_25[2]),.din(w_n6505_8[0]));
	jspl3 jspl3_w_n6505_26(.douta(w_n6505_26[0]),.doutb(w_n6505_26[1]),.doutc(w_n6505_26[2]),.din(w_n6505_8[1]));
	jspl3 jspl3_w_n6505_27(.douta(w_n6505_27[0]),.doutb(w_n6505_27[1]),.doutc(w_n6505_27[2]),.din(w_n6505_8[2]));
	jspl jspl_w_n6505_28(.douta(w_n6505_28[0]),.doutb(w_n6505_28[1]),.din(w_n6505_9[0]));
	jspl jspl_w_n6508_0(.douta(w_n6508_0[0]),.doutb(w_n6508_0[1]),.din(n6508));
	jspl3 jspl3_w_n6510_0(.douta(w_n6510_0[0]),.doutb(w_n6510_0[1]),.doutc(w_n6510_0[2]),.din(n6510));
	jspl jspl_w_n6510_1(.douta(w_n6510_1[0]),.doutb(w_n6510_1[1]),.din(w_n6510_0[0]));
	jspl3 jspl3_w_n6511_0(.douta(w_n6511_0[0]),.doutb(w_n6511_0[1]),.doutc(w_n6511_0[2]),.din(n6511));
	jspl3 jspl3_w_n6515_0(.douta(w_n6515_0[0]),.doutb(w_n6515_0[1]),.doutc(w_n6515_0[2]),.din(n6515));
	jspl jspl_w_n6516_0(.douta(w_n6516_0[0]),.doutb(w_n6516_0[1]),.din(n6516));
	jspl jspl_w_n6517_0(.douta(w_n6517_0[0]),.doutb(w_n6517_0[1]),.din(n6517));
	jspl jspl_w_n6518_0(.douta(w_n6518_0[0]),.doutb(w_n6518_0[1]),.din(n6518));
	jspl jspl_w_n6520_0(.douta(w_n6520_0[0]),.doutb(w_n6520_0[1]),.din(n6520));
	jspl jspl_w_n6522_0(.douta(w_n6522_0[0]),.doutb(w_n6522_0[1]),.din(n6522));
	jspl jspl_w_n6524_0(.douta(w_n6524_0[0]),.doutb(w_n6524_0[1]),.din(n6524));
	jspl jspl_w_n6527_0(.douta(w_n6527_0[0]),.doutb(w_n6527_0[1]),.din(n6527));
	jspl jspl_w_n6532_0(.douta(w_n6532_0[0]),.doutb(w_n6532_0[1]),.din(n6532));
	jspl3 jspl3_w_n6534_0(.douta(w_n6534_0[0]),.doutb(w_n6534_0[1]),.doutc(w_n6534_0[2]),.din(n6534));
	jspl jspl_w_n6535_0(.douta(w_n6535_0[0]),.doutb(w_n6535_0[1]),.din(n6535));
	jspl jspl_w_n6539_0(.douta(w_n6539_0[0]),.doutb(w_n6539_0[1]),.din(n6539));
	jspl jspl_w_n6540_0(.douta(w_n6540_0[0]),.doutb(w_n6540_0[1]),.din(n6540));
	jspl jspl_w_n6542_0(.douta(w_n6542_0[0]),.doutb(w_n6542_0[1]),.din(n6542));
	jspl jspl_w_n6544_0(.douta(w_n6544_0[0]),.doutb(w_n6544_0[1]),.din(n6544));
	jspl jspl_w_n6547_0(.douta(w_n6547_0[0]),.doutb(w_n6547_0[1]),.din(n6547));
	jspl jspl_w_n6553_0(.douta(w_n6553_0[0]),.doutb(w_n6553_0[1]),.din(n6553));
	jspl3 jspl3_w_n6555_0(.douta(w_n6555_0[0]),.doutb(w_n6555_0[1]),.doutc(w_n6555_0[2]),.din(n6555));
	jspl jspl_w_n6556_0(.douta(w_n6556_0[0]),.doutb(w_n6556_0[1]),.din(n6556));
	jspl jspl_w_n6559_0(.douta(w_n6559_0[0]),.doutb(w_n6559_0[1]),.din(n6559));
	jspl jspl_w_n6561_0(.douta(w_n6561_0[0]),.doutb(w_n6561_0[1]),.din(n6561));
	jspl jspl_w_n6565_0(.douta(w_n6565_0[0]),.doutb(w_n6565_0[1]),.din(n6565));
	jspl jspl_w_n6567_0(.douta(w_n6567_0[0]),.doutb(w_n6567_0[1]),.din(n6567));
	jspl jspl_w_n6568_0(.douta(w_n6568_0[0]),.doutb(w_n6568_0[1]),.din(n6568));
	jspl3 jspl3_w_n6569_0(.douta(w_n6569_0[0]),.doutb(w_n6569_0[1]),.doutc(w_n6569_0[2]),.din(n6569));
	jspl jspl_w_n6570_0(.douta(w_n6570_0[0]),.doutb(w_n6570_0[1]),.din(n6570));
	jspl jspl_w_n6575_0(.douta(w_n6575_0[0]),.doutb(w_n6575_0[1]),.din(n6575));
	jspl jspl_w_n6577_0(.douta(w_n6577_0[0]),.doutb(w_n6577_0[1]),.din(n6577));
	jspl jspl_w_n6579_0(.douta(w_n6579_0[0]),.doutb(w_n6579_0[1]),.din(n6579));
	jspl jspl_w_n6583_0(.douta(w_n6583_0[0]),.doutb(w_n6583_0[1]),.din(n6583));
	jspl jspl_w_n6585_0(.douta(w_n6585_0[0]),.doutb(w_n6585_0[1]),.din(n6585));
	jspl jspl_w_n6586_0(.douta(w_n6586_0[0]),.doutb(w_n6586_0[1]),.din(n6586));
	jspl3 jspl3_w_n6587_0(.douta(w_n6587_0[0]),.doutb(w_n6587_0[1]),.doutc(w_n6587_0[2]),.din(n6587));
	jspl jspl_w_n6588_0(.douta(w_n6588_0[0]),.doutb(w_n6588_0[1]),.din(n6588));
	jspl jspl_w_n6594_0(.douta(w_n6594_0[0]),.doutb(w_n6594_0[1]),.din(n6594));
	jspl jspl_w_n6595_0(.douta(w_n6595_0[0]),.doutb(w_n6595_0[1]),.din(n6595));
	jspl jspl_w_n6597_0(.douta(w_n6597_0[0]),.doutb(w_n6597_0[1]),.din(n6597));
	jspl jspl_w_n6599_0(.douta(w_n6599_0[0]),.doutb(w_n6599_0[1]),.din(n6599));
	jspl jspl_w_n6601_0(.douta(w_n6601_0[0]),.doutb(w_n6601_0[1]),.din(n6601));
	jspl jspl_w_n6607_0(.douta(w_n6607_0[0]),.doutb(w_n6607_0[1]),.din(n6607));
	jspl jspl_w_n6609_0(.douta(w_n6609_0[0]),.doutb(w_n6609_0[1]),.din(n6609));
	jspl3 jspl3_w_n6610_0(.douta(w_n6610_0[0]),.doutb(w_n6610_0[1]),.doutc(w_n6610_0[2]),.din(n6610));
	jspl jspl_w_n6613_0(.douta(w_n6613_0[0]),.doutb(w_n6613_0[1]),.din(n6613));
	jspl jspl_w_n6614_0(.douta(w_n6614_0[0]),.doutb(w_n6614_0[1]),.din(n6614));
	jspl3 jspl3_w_n6615_0(.douta(w_n6615_0[0]),.doutb(w_n6615_0[1]),.doutc(w_n6615_0[2]),.din(n6615));
	jspl jspl_w_n6617_0(.douta(w_n6617_0[0]),.doutb(w_n6617_0[1]),.din(n6617));
	jspl jspl_w_n6621_0(.douta(w_n6621_0[0]),.doutb(w_n6621_0[1]),.din(n6621));
	jspl jspl_w_n6623_0(.douta(w_n6623_0[0]),.doutb(w_n6623_0[1]),.din(n6623));
	jspl jspl_w_n6624_0(.douta(w_n6624_0[0]),.doutb(w_n6624_0[1]),.din(n6624));
	jspl3 jspl3_w_n6625_0(.douta(w_n6625_0[0]),.doutb(w_n6625_0[1]),.doutc(w_n6625_0[2]),.din(n6625));
	jspl jspl_w_n6626_0(.douta(w_n6626_0[0]),.doutb(w_n6626_0[1]),.din(n6626));
	jspl jspl_w_n6629_0(.douta(w_n6629_0[0]),.doutb(w_n6629_0[1]),.din(n6629));
	jspl jspl_w_n6635_0(.douta(w_n6635_0[0]),.doutb(w_n6635_0[1]),.din(n6635));
	jspl jspl_w_n6636_0(.douta(w_n6636_0[0]),.doutb(w_n6636_0[1]),.din(n6636));
	jspl jspl_w_n6638_0(.douta(w_n6638_0[0]),.doutb(w_n6638_0[1]),.din(n6638));
	jspl jspl_w_n6640_0(.douta(w_n6640_0[0]),.doutb(w_n6640_0[1]),.din(n6640));
	jspl jspl_w_n6642_0(.douta(w_n6642_0[0]),.doutb(w_n6642_0[1]),.din(n6642));
	jspl jspl_w_n6648_0(.douta(w_n6648_0[0]),.doutb(w_n6648_0[1]),.din(n6648));
	jspl jspl_w_n6650_0(.douta(w_n6650_0[0]),.doutb(w_n6650_0[1]),.din(n6650));
	jspl3 jspl3_w_n6651_0(.douta(w_n6651_0[0]),.doutb(w_n6651_0[1]),.doutc(w_n6651_0[2]),.din(n6651));
	jspl jspl_w_n6654_0(.douta(w_n6654_0[0]),.doutb(w_n6654_0[1]),.din(n6654));
	jspl jspl_w_n6655_0(.douta(w_n6655_0[0]),.doutb(w_n6655_0[1]),.din(n6655));
	jspl3 jspl3_w_n6656_0(.douta(w_n6656_0[0]),.doutb(w_n6656_0[1]),.doutc(w_n6656_0[2]),.din(n6656));
	jspl jspl_w_n6658_0(.douta(w_n6658_0[0]),.doutb(w_n6658_0[1]),.din(n6658));
	jspl jspl_w_n6662_0(.douta(w_n6662_0[0]),.doutb(w_n6662_0[1]),.din(n6662));
	jspl jspl_w_n6664_0(.douta(w_n6664_0[0]),.doutb(w_n6664_0[1]),.din(n6664));
	jspl jspl_w_n6665_0(.douta(w_n6665_0[0]),.doutb(w_n6665_0[1]),.din(n6665));
	jspl3 jspl3_w_n6666_0(.douta(w_n6666_0[0]),.doutb(w_n6666_0[1]),.doutc(w_n6666_0[2]),.din(n6666));
	jspl jspl_w_n6667_0(.douta(w_n6667_0[0]),.doutb(w_n6667_0[1]),.din(n6667));
	jspl jspl_w_n6670_0(.douta(w_n6670_0[0]),.doutb(w_n6670_0[1]),.din(n6670));
	jspl jspl_w_n6676_0(.douta(w_n6676_0[0]),.doutb(w_n6676_0[1]),.din(n6676));
	jspl jspl_w_n6677_0(.douta(w_n6677_0[0]),.doutb(w_n6677_0[1]),.din(n6677));
	jspl jspl_w_n6679_0(.douta(w_n6679_0[0]),.doutb(w_n6679_0[1]),.din(n6679));
	jspl jspl_w_n6681_0(.douta(w_n6681_0[0]),.doutb(w_n6681_0[1]),.din(n6681));
	jspl jspl_w_n6683_0(.douta(w_n6683_0[0]),.doutb(w_n6683_0[1]),.din(n6683));
	jspl jspl_w_n6689_0(.douta(w_n6689_0[0]),.doutb(w_n6689_0[1]),.din(n6689));
	jspl jspl_w_n6691_0(.douta(w_n6691_0[0]),.doutb(w_n6691_0[1]),.din(n6691));
	jspl3 jspl3_w_n6692_0(.douta(w_n6692_0[0]),.doutb(w_n6692_0[1]),.doutc(w_n6692_0[2]),.din(n6692));
	jspl jspl_w_n6695_0(.douta(w_n6695_0[0]),.doutb(w_n6695_0[1]),.din(n6695));
	jspl jspl_w_n6696_0(.douta(w_n6696_0[0]),.doutb(w_n6696_0[1]),.din(n6696));
	jspl3 jspl3_w_n6697_0(.douta(w_n6697_0[0]),.doutb(w_n6697_0[1]),.doutc(w_n6697_0[2]),.din(n6697));
	jspl jspl_w_n6699_0(.douta(w_n6699_0[0]),.doutb(w_n6699_0[1]),.din(n6699));
	jspl jspl_w_n6703_0(.douta(w_n6703_0[0]),.doutb(w_n6703_0[1]),.din(n6703));
	jspl jspl_w_n6705_0(.douta(w_n6705_0[0]),.doutb(w_n6705_0[1]),.din(n6705));
	jspl jspl_w_n6706_0(.douta(w_n6706_0[0]),.doutb(w_n6706_0[1]),.din(n6706));
	jspl3 jspl3_w_n6707_0(.douta(w_n6707_0[0]),.doutb(w_n6707_0[1]),.doutc(w_n6707_0[2]),.din(n6707));
	jspl jspl_w_n6708_0(.douta(w_n6708_0[0]),.doutb(w_n6708_0[1]),.din(n6708));
	jspl jspl_w_n6711_0(.douta(w_n6711_0[0]),.doutb(w_n6711_0[1]),.din(n6711));
	jspl jspl_w_n6717_0(.douta(w_n6717_0[0]),.doutb(w_n6717_0[1]),.din(n6717));
	jspl jspl_w_n6718_0(.douta(w_n6718_0[0]),.doutb(w_n6718_0[1]),.din(n6718));
	jspl jspl_w_n6720_0(.douta(w_n6720_0[0]),.doutb(w_n6720_0[1]),.din(n6720));
	jspl jspl_w_n6722_0(.douta(w_n6722_0[0]),.doutb(w_n6722_0[1]),.din(n6722));
	jspl jspl_w_n6724_0(.douta(w_n6724_0[0]),.doutb(w_n6724_0[1]),.din(n6724));
	jspl jspl_w_n6730_0(.douta(w_n6730_0[0]),.doutb(w_n6730_0[1]),.din(n6730));
	jspl jspl_w_n6732_0(.douta(w_n6732_0[0]),.doutb(w_n6732_0[1]),.din(n6732));
	jspl3 jspl3_w_n6733_0(.douta(w_n6733_0[0]),.doutb(w_n6733_0[1]),.doutc(w_n6733_0[2]),.din(n6733));
	jspl jspl_w_n6736_0(.douta(w_n6736_0[0]),.doutb(w_n6736_0[1]),.din(n6736));
	jspl jspl_w_n6737_0(.douta(w_n6737_0[0]),.doutb(w_n6737_0[1]),.din(n6737));
	jspl3 jspl3_w_n6738_0(.douta(w_n6738_0[0]),.doutb(w_n6738_0[1]),.doutc(w_n6738_0[2]),.din(n6738));
	jspl jspl_w_n6740_0(.douta(w_n6740_0[0]),.doutb(w_n6740_0[1]),.din(n6740));
	jspl jspl_w_n6744_0(.douta(w_n6744_0[0]),.doutb(w_n6744_0[1]),.din(n6744));
	jspl jspl_w_n6746_0(.douta(w_n6746_0[0]),.doutb(w_n6746_0[1]),.din(n6746));
	jspl jspl_w_n6747_0(.douta(w_n6747_0[0]),.doutb(w_n6747_0[1]),.din(n6747));
	jspl3 jspl3_w_n6748_0(.douta(w_n6748_0[0]),.doutb(w_n6748_0[1]),.doutc(w_n6748_0[2]),.din(n6748));
	jspl jspl_w_n6749_0(.douta(w_n6749_0[0]),.doutb(w_n6749_0[1]),.din(n6749));
	jspl jspl_w_n6752_0(.douta(w_n6752_0[0]),.doutb(w_n6752_0[1]),.din(n6752));
	jspl jspl_w_n6758_0(.douta(w_n6758_0[0]),.doutb(w_n6758_0[1]),.din(n6758));
	jspl jspl_w_n6759_0(.douta(w_n6759_0[0]),.doutb(w_n6759_0[1]),.din(n6759));
	jspl jspl_w_n6761_0(.douta(w_n6761_0[0]),.doutb(w_n6761_0[1]),.din(n6761));
	jspl jspl_w_n6763_0(.douta(w_n6763_0[0]),.doutb(w_n6763_0[1]),.din(n6763));
	jspl jspl_w_n6765_0(.douta(w_n6765_0[0]),.doutb(w_n6765_0[1]),.din(n6765));
	jspl jspl_w_n6771_0(.douta(w_n6771_0[0]),.doutb(w_n6771_0[1]),.din(n6771));
	jspl jspl_w_n6773_0(.douta(w_n6773_0[0]),.doutb(w_n6773_0[1]),.din(n6773));
	jspl3 jspl3_w_n6774_0(.douta(w_n6774_0[0]),.doutb(w_n6774_0[1]),.doutc(w_n6774_0[2]),.din(n6774));
	jspl jspl_w_n6777_0(.douta(w_n6777_0[0]),.doutb(w_n6777_0[1]),.din(n6777));
	jspl jspl_w_n6778_0(.douta(w_n6778_0[0]),.doutb(w_n6778_0[1]),.din(n6778));
	jspl3 jspl3_w_n6779_0(.douta(w_n6779_0[0]),.doutb(w_n6779_0[1]),.doutc(w_n6779_0[2]),.din(n6779));
	jspl jspl_w_n6781_0(.douta(w_n6781_0[0]),.doutb(w_n6781_0[1]),.din(n6781));
	jspl jspl_w_n6785_0(.douta(w_n6785_0[0]),.doutb(w_n6785_0[1]),.din(n6785));
	jspl jspl_w_n6787_0(.douta(w_n6787_0[0]),.doutb(w_n6787_0[1]),.din(n6787));
	jspl jspl_w_n6788_0(.douta(w_n6788_0[0]),.doutb(w_n6788_0[1]),.din(n6788));
	jspl3 jspl3_w_n6789_0(.douta(w_n6789_0[0]),.doutb(w_n6789_0[1]),.doutc(w_n6789_0[2]),.din(n6789));
	jspl jspl_w_n6790_0(.douta(w_n6790_0[0]),.doutb(w_n6790_0[1]),.din(n6790));
	jspl jspl_w_n6793_0(.douta(w_n6793_0[0]),.doutb(w_n6793_0[1]),.din(n6793));
	jspl jspl_w_n6799_0(.douta(w_n6799_0[0]),.doutb(w_n6799_0[1]),.din(n6799));
	jspl jspl_w_n6800_0(.douta(w_n6800_0[0]),.doutb(w_n6800_0[1]),.din(n6800));
	jspl jspl_w_n6802_0(.douta(w_n6802_0[0]),.doutb(w_n6802_0[1]),.din(n6802));
	jspl jspl_w_n6804_0(.douta(w_n6804_0[0]),.doutb(w_n6804_0[1]),.din(n6804));
	jspl jspl_w_n6806_0(.douta(w_n6806_0[0]),.doutb(w_n6806_0[1]),.din(n6806));
	jspl jspl_w_n6812_0(.douta(w_n6812_0[0]),.doutb(w_n6812_0[1]),.din(n6812));
	jspl jspl_w_n6814_0(.douta(w_n6814_0[0]),.doutb(w_n6814_0[1]),.din(n6814));
	jspl3 jspl3_w_n6815_0(.douta(w_n6815_0[0]),.doutb(w_n6815_0[1]),.doutc(w_n6815_0[2]),.din(n6815));
	jspl jspl_w_n6818_0(.douta(w_n6818_0[0]),.doutb(w_n6818_0[1]),.din(n6818));
	jspl jspl_w_n6819_0(.douta(w_n6819_0[0]),.doutb(w_n6819_0[1]),.din(n6819));
	jspl3 jspl3_w_n6820_0(.douta(w_n6820_0[0]),.doutb(w_n6820_0[1]),.doutc(w_n6820_0[2]),.din(n6820));
	jspl jspl_w_n6822_0(.douta(w_n6822_0[0]),.doutb(w_n6822_0[1]),.din(n6822));
	jspl jspl_w_n6826_0(.douta(w_n6826_0[0]),.doutb(w_n6826_0[1]),.din(n6826));
	jspl jspl_w_n6828_0(.douta(w_n6828_0[0]),.doutb(w_n6828_0[1]),.din(n6828));
	jspl jspl_w_n6829_0(.douta(w_n6829_0[0]),.doutb(w_n6829_0[1]),.din(n6829));
	jspl3 jspl3_w_n6830_0(.douta(w_n6830_0[0]),.doutb(w_n6830_0[1]),.doutc(w_n6830_0[2]),.din(n6830));
	jspl jspl_w_n6834_0(.douta(w_n6834_0[0]),.doutb(w_n6834_0[1]),.din(n6834));
	jspl jspl_w_n6840_0(.douta(w_n6840_0[0]),.doutb(w_n6840_0[1]),.din(n6840));
	jspl3 jspl3_w_n6842_0(.douta(w_n6842_0[0]),.doutb(w_n6842_0[1]),.doutc(w_n6842_0[2]),.din(n6842));
	jspl jspl_w_n6844_0(.douta(w_n6844_0[0]),.doutb(w_n6844_0[1]),.din(n6844));
	jspl3 jspl3_w_n6849_0(.douta(w_n6849_0[0]),.doutb(w_n6849_0[1]),.doutc(w_n6849_0[2]),.din(n6849));
	jspl jspl_w_n6850_0(.douta(w_n6850_0[0]),.doutb(w_n6850_0[1]),.din(n6850));
	jspl jspl_w_n6851_0(.douta(w_n6851_0[0]),.doutb(w_n6851_0[1]),.din(n6851));
	jspl jspl_w_n6856_0(.douta(w_n6856_0[0]),.doutb(w_n6856_0[1]),.din(n6856));
	jspl3 jspl3_w_n6857_0(.douta(w_n6857_0[0]),.doutb(w_n6857_0[1]),.doutc(w_n6857_0[2]),.din(n6857));
	jspl jspl_w_n6862_0(.douta(w_n6862_0[0]),.doutb(w_n6862_0[1]),.din(n6862));
	jspl jspl_w_n6869_0(.douta(w_n6869_0[0]),.doutb(w_n6869_0[1]),.din(n6869));
	jspl3 jspl3_w_n6872_0(.douta(w_n6872_0[0]),.doutb(w_n6872_0[1]),.doutc(w_n6872_0[2]),.din(n6872));
	jspl jspl_w_n6872_1(.douta(w_n6872_1[0]),.doutb(w_n6872_1[1]),.din(w_n6872_0[0]));
	jspl jspl_w_n6873_0(.douta(w_n6873_0[0]),.doutb(w_n6873_0[1]),.din(n6873));
	jspl3 jspl3_w_n6876_0(.douta(w_n6876_0[0]),.doutb(w_n6876_0[1]),.doutc(w_n6876_0[2]),.din(n6876));
	jspl jspl_w_n6877_0(.douta(w_n6877_0[0]),.doutb(w_n6877_0[1]),.din(n6877));
	jspl jspl_w_n6878_0(.douta(w_n6878_0[0]),.doutb(w_n6878_0[1]),.din(n6878));
	jspl jspl_w_n6879_0(.douta(w_n6879_0[0]),.doutb(w_n6879_0[1]),.din(n6879));
	jspl jspl_w_n6881_0(.douta(w_n6881_0[0]),.doutb(w_n6881_0[1]),.din(n6881));
	jspl jspl_w_n6883_0(.douta(w_n6883_0[0]),.doutb(w_n6883_0[1]),.din(n6883));
	jspl jspl_w_n6885_0(.douta(w_n6885_0[0]),.doutb(w_n6885_0[1]),.din(n6885));
	jspl jspl_w_n6894_0(.douta(w_n6894_0[0]),.doutb(w_n6894_0[1]),.din(n6894));
	jspl3 jspl3_w_n6896_0(.douta(w_n6896_0[0]),.doutb(w_n6896_0[1]),.doutc(w_n6896_0[2]),.din(n6896));
	jspl jspl_w_n6897_0(.douta(w_n6897_0[0]),.doutb(w_n6897_0[1]),.din(n6897));
	jspl jspl_w_n6901_0(.douta(w_n6901_0[0]),.doutb(w_n6901_0[1]),.din(n6901));
	jspl jspl_w_n6903_0(.douta(w_n6903_0[0]),.doutb(w_n6903_0[1]),.din(n6903));
	jspl jspl_w_n6905_0(.douta(w_n6905_0[0]),.doutb(w_n6905_0[1]),.din(n6905));
	jspl jspl_w_n6910_0(.douta(w_n6910_0[0]),.doutb(w_n6910_0[1]),.din(n6910));
	jspl jspl_w_n6912_0(.douta(w_n6912_0[0]),.doutb(w_n6912_0[1]),.din(n6912));
	jspl jspl_w_n6913_0(.douta(w_n6913_0[0]),.doutb(w_n6913_0[1]),.din(n6913));
	jspl3 jspl3_w_n6914_0(.douta(w_n6914_0[0]),.doutb(w_n6914_0[1]),.doutc(w_n6914_0[2]),.din(n6914));
	jspl jspl_w_n6915_0(.douta(w_n6915_0[0]),.doutb(w_n6915_0[1]),.din(n6915));
	jspl jspl_w_n6920_0(.douta(w_n6920_0[0]),.doutb(w_n6920_0[1]),.din(n6920));
	jspl jspl_w_n6921_0(.douta(w_n6921_0[0]),.doutb(w_n6921_0[1]),.din(n6921));
	jspl jspl_w_n6923_0(.douta(w_n6923_0[0]),.doutb(w_n6923_0[1]),.din(n6923));
	jspl jspl_w_n6928_0(.douta(w_n6928_0[0]),.doutb(w_n6928_0[1]),.din(n6928));
	jspl jspl_w_n6930_0(.douta(w_n6930_0[0]),.doutb(w_n6930_0[1]),.din(n6930));
	jspl jspl_w_n6931_0(.douta(w_n6931_0[0]),.doutb(w_n6931_0[1]),.din(n6931));
	jspl3 jspl3_w_n6932_0(.douta(w_n6932_0[0]),.doutb(w_n6932_0[1]),.doutc(w_n6932_0[2]),.din(n6932));
	jspl jspl_w_n6933_0(.douta(w_n6933_0[0]),.doutb(w_n6933_0[1]),.din(n6933));
	jspl jspl_w_n6935_0(.douta(w_n6935_0[0]),.doutb(w_n6935_0[1]),.din(n6935));
	jspl jspl_w_n6937_0(.douta(w_n6937_0[0]),.doutb(w_n6937_0[1]),.din(n6937));
	jspl jspl_w_n6939_0(.douta(w_n6939_0[0]),.doutb(w_n6939_0[1]),.din(n6939));
	jspl jspl_w_n6942_0(.douta(w_n6942_0[0]),.doutb(w_n6942_0[1]),.din(n6942));
	jspl jspl_w_n6948_0(.douta(w_n6948_0[0]),.doutb(w_n6948_0[1]),.din(n6948));
	jspl3 jspl3_w_n6950_0(.douta(w_n6950_0[0]),.doutb(w_n6950_0[1]),.doutc(w_n6950_0[2]),.din(n6950));
	jspl jspl_w_n6951_0(.douta(w_n6951_0[0]),.doutb(w_n6951_0[1]),.din(n6951));
	jspl jspl_w_n6955_0(.douta(w_n6955_0[0]),.doutb(w_n6955_0[1]),.din(n6955));
	jspl jspl_w_n6956_0(.douta(w_n6956_0[0]),.doutb(w_n6956_0[1]),.din(n6956));
	jspl jspl_w_n6958_0(.douta(w_n6958_0[0]),.doutb(w_n6958_0[1]),.din(n6958));
	jspl jspl_w_n6960_0(.douta(w_n6960_0[0]),.doutb(w_n6960_0[1]),.din(n6960));
	jspl jspl_w_n6963_0(.douta(w_n6963_0[0]),.doutb(w_n6963_0[1]),.din(n6963));
	jspl jspl_w_n6969_0(.douta(w_n6969_0[0]),.doutb(w_n6969_0[1]),.din(n6969));
	jspl jspl_w_n6971_0(.douta(w_n6971_0[0]),.doutb(w_n6971_0[1]),.din(n6971));
	jspl3 jspl3_w_n6972_0(.douta(w_n6972_0[0]),.doutb(w_n6972_0[1]),.doutc(w_n6972_0[2]),.din(n6972));
	jspl jspl_w_n6976_0(.douta(w_n6976_0[0]),.doutb(w_n6976_0[1]),.din(n6976));
	jspl jspl_w_n6977_0(.douta(w_n6977_0[0]),.doutb(w_n6977_0[1]),.din(n6977));
	jspl3 jspl3_w_n6978_0(.douta(w_n6978_0[0]),.doutb(w_n6978_0[1]),.doutc(w_n6978_0[2]),.din(n6978));
	jspl jspl_w_n6980_0(.douta(w_n6980_0[0]),.doutb(w_n6980_0[1]),.din(n6980));
	jspl jspl_w_n6985_0(.douta(w_n6985_0[0]),.doutb(w_n6985_0[1]),.din(n6985));
	jspl jspl_w_n6987_0(.douta(w_n6987_0[0]),.doutb(w_n6987_0[1]),.din(n6987));
	jspl jspl_w_n6988_0(.douta(w_n6988_0[0]),.doutb(w_n6988_0[1]),.din(n6988));
	jspl3 jspl3_w_n6989_0(.douta(w_n6989_0[0]),.doutb(w_n6989_0[1]),.doutc(w_n6989_0[2]),.din(n6989));
	jspl jspl_w_n6990_0(.douta(w_n6990_0[0]),.doutb(w_n6990_0[1]),.din(n6990));
	jspl jspl_w_n6994_0(.douta(w_n6994_0[0]),.doutb(w_n6994_0[1]),.din(n6994));
	jspl jspl_w_n7000_0(.douta(w_n7000_0[0]),.doutb(w_n7000_0[1]),.din(n7000));
	jspl jspl_w_n7001_0(.douta(w_n7001_0[0]),.doutb(w_n7001_0[1]),.din(n7001));
	jspl jspl_w_n7003_0(.douta(w_n7003_0[0]),.doutb(w_n7003_0[1]),.din(n7003));
	jspl jspl_w_n7005_0(.douta(w_n7005_0[0]),.doutb(w_n7005_0[1]),.din(n7005));
	jspl jspl_w_n7008_0(.douta(w_n7008_0[0]),.doutb(w_n7008_0[1]),.din(n7008));
	jspl jspl_w_n7014_0(.douta(w_n7014_0[0]),.doutb(w_n7014_0[1]),.din(n7014));
	jspl jspl_w_n7016_0(.douta(w_n7016_0[0]),.doutb(w_n7016_0[1]),.din(n7016));
	jspl3 jspl3_w_n7017_0(.douta(w_n7017_0[0]),.doutb(w_n7017_0[1]),.doutc(w_n7017_0[2]),.din(n7017));
	jspl jspl_w_n7021_0(.douta(w_n7021_0[0]),.doutb(w_n7021_0[1]),.din(n7021));
	jspl jspl_w_n7022_0(.douta(w_n7022_0[0]),.doutb(w_n7022_0[1]),.din(n7022));
	jspl3 jspl3_w_n7023_0(.douta(w_n7023_0[0]),.doutb(w_n7023_0[1]),.doutc(w_n7023_0[2]),.din(n7023));
	jspl jspl_w_n7025_0(.douta(w_n7025_0[0]),.doutb(w_n7025_0[1]),.din(n7025));
	jspl jspl_w_n7030_0(.douta(w_n7030_0[0]),.doutb(w_n7030_0[1]),.din(n7030));
	jspl jspl_w_n7032_0(.douta(w_n7032_0[0]),.doutb(w_n7032_0[1]),.din(n7032));
	jspl jspl_w_n7033_0(.douta(w_n7033_0[0]),.doutb(w_n7033_0[1]),.din(n7033));
	jspl3 jspl3_w_n7034_0(.douta(w_n7034_0[0]),.doutb(w_n7034_0[1]),.doutc(w_n7034_0[2]),.din(n7034));
	jspl jspl_w_n7035_0(.douta(w_n7035_0[0]),.doutb(w_n7035_0[1]),.din(n7035));
	jspl jspl_w_n7039_0(.douta(w_n7039_0[0]),.doutb(w_n7039_0[1]),.din(n7039));
	jspl jspl_w_n7045_0(.douta(w_n7045_0[0]),.doutb(w_n7045_0[1]),.din(n7045));
	jspl jspl_w_n7046_0(.douta(w_n7046_0[0]),.doutb(w_n7046_0[1]),.din(n7046));
	jspl jspl_w_n7048_0(.douta(w_n7048_0[0]),.doutb(w_n7048_0[1]),.din(n7048));
	jspl jspl_w_n7050_0(.douta(w_n7050_0[0]),.doutb(w_n7050_0[1]),.din(n7050));
	jspl jspl_w_n7053_0(.douta(w_n7053_0[0]),.doutb(w_n7053_0[1]),.din(n7053));
	jspl jspl_w_n7059_0(.douta(w_n7059_0[0]),.doutb(w_n7059_0[1]),.din(n7059));
	jspl jspl_w_n7061_0(.douta(w_n7061_0[0]),.doutb(w_n7061_0[1]),.din(n7061));
	jspl3 jspl3_w_n7062_0(.douta(w_n7062_0[0]),.doutb(w_n7062_0[1]),.doutc(w_n7062_0[2]),.din(n7062));
	jspl jspl_w_n7066_0(.douta(w_n7066_0[0]),.doutb(w_n7066_0[1]),.din(n7066));
	jspl jspl_w_n7067_0(.douta(w_n7067_0[0]),.doutb(w_n7067_0[1]),.din(n7067));
	jspl3 jspl3_w_n7068_0(.douta(w_n7068_0[0]),.doutb(w_n7068_0[1]),.doutc(w_n7068_0[2]),.din(n7068));
	jspl jspl_w_n7070_0(.douta(w_n7070_0[0]),.doutb(w_n7070_0[1]),.din(n7070));
	jspl jspl_w_n7075_0(.douta(w_n7075_0[0]),.doutb(w_n7075_0[1]),.din(n7075));
	jspl jspl_w_n7077_0(.douta(w_n7077_0[0]),.doutb(w_n7077_0[1]),.din(n7077));
	jspl jspl_w_n7078_0(.douta(w_n7078_0[0]),.doutb(w_n7078_0[1]),.din(n7078));
	jspl3 jspl3_w_n7079_0(.douta(w_n7079_0[0]),.doutb(w_n7079_0[1]),.doutc(w_n7079_0[2]),.din(n7079));
	jspl jspl_w_n7080_0(.douta(w_n7080_0[0]),.doutb(w_n7080_0[1]),.din(n7080));
	jspl jspl_w_n7084_0(.douta(w_n7084_0[0]),.doutb(w_n7084_0[1]),.din(n7084));
	jspl jspl_w_n7090_0(.douta(w_n7090_0[0]),.doutb(w_n7090_0[1]),.din(n7090));
	jspl jspl_w_n7091_0(.douta(w_n7091_0[0]),.doutb(w_n7091_0[1]),.din(n7091));
	jspl jspl_w_n7093_0(.douta(w_n7093_0[0]),.doutb(w_n7093_0[1]),.din(n7093));
	jspl jspl_w_n7095_0(.douta(w_n7095_0[0]),.doutb(w_n7095_0[1]),.din(n7095));
	jspl jspl_w_n7098_0(.douta(w_n7098_0[0]),.doutb(w_n7098_0[1]),.din(n7098));
	jspl jspl_w_n7104_0(.douta(w_n7104_0[0]),.doutb(w_n7104_0[1]),.din(n7104));
	jspl jspl_w_n7106_0(.douta(w_n7106_0[0]),.doutb(w_n7106_0[1]),.din(n7106));
	jspl3 jspl3_w_n7107_0(.douta(w_n7107_0[0]),.doutb(w_n7107_0[1]),.doutc(w_n7107_0[2]),.din(n7107));
	jspl jspl_w_n7111_0(.douta(w_n7111_0[0]),.doutb(w_n7111_0[1]),.din(n7111));
	jspl jspl_w_n7112_0(.douta(w_n7112_0[0]),.doutb(w_n7112_0[1]),.din(n7112));
	jspl3 jspl3_w_n7113_0(.douta(w_n7113_0[0]),.doutb(w_n7113_0[1]),.doutc(w_n7113_0[2]),.din(n7113));
	jspl jspl_w_n7115_0(.douta(w_n7115_0[0]),.doutb(w_n7115_0[1]),.din(n7115));
	jspl jspl_w_n7120_0(.douta(w_n7120_0[0]),.doutb(w_n7120_0[1]),.din(n7120));
	jspl jspl_w_n7122_0(.douta(w_n7122_0[0]),.doutb(w_n7122_0[1]),.din(n7122));
	jspl jspl_w_n7123_0(.douta(w_n7123_0[0]),.doutb(w_n7123_0[1]),.din(n7123));
	jspl3 jspl3_w_n7124_0(.douta(w_n7124_0[0]),.doutb(w_n7124_0[1]),.doutc(w_n7124_0[2]),.din(n7124));
	jspl jspl_w_n7125_0(.douta(w_n7125_0[0]),.doutb(w_n7125_0[1]),.din(n7125));
	jspl jspl_w_n7129_0(.douta(w_n7129_0[0]),.doutb(w_n7129_0[1]),.din(n7129));
	jspl jspl_w_n7135_0(.douta(w_n7135_0[0]),.doutb(w_n7135_0[1]),.din(n7135));
	jspl jspl_w_n7136_0(.douta(w_n7136_0[0]),.doutb(w_n7136_0[1]),.din(n7136));
	jspl jspl_w_n7138_0(.douta(w_n7138_0[0]),.doutb(w_n7138_0[1]),.din(n7138));
	jspl jspl_w_n7140_0(.douta(w_n7140_0[0]),.doutb(w_n7140_0[1]),.din(n7140));
	jspl jspl_w_n7143_0(.douta(w_n7143_0[0]),.doutb(w_n7143_0[1]),.din(n7143));
	jspl jspl_w_n7149_0(.douta(w_n7149_0[0]),.doutb(w_n7149_0[1]),.din(n7149));
	jspl jspl_w_n7151_0(.douta(w_n7151_0[0]),.doutb(w_n7151_0[1]),.din(n7151));
	jspl3 jspl3_w_n7152_0(.douta(w_n7152_0[0]),.doutb(w_n7152_0[1]),.doutc(w_n7152_0[2]),.din(n7152));
	jspl jspl_w_n7156_0(.douta(w_n7156_0[0]),.doutb(w_n7156_0[1]),.din(n7156));
	jspl jspl_w_n7157_0(.douta(w_n7157_0[0]),.doutb(w_n7157_0[1]),.din(n7157));
	jspl3 jspl3_w_n7158_0(.douta(w_n7158_0[0]),.doutb(w_n7158_0[1]),.doutc(w_n7158_0[2]),.din(n7158));
	jspl jspl_w_n7160_0(.douta(w_n7160_0[0]),.doutb(w_n7160_0[1]),.din(n7160));
	jspl jspl_w_n7165_0(.douta(w_n7165_0[0]),.doutb(w_n7165_0[1]),.din(n7165));
	jspl jspl_w_n7167_0(.douta(w_n7167_0[0]),.doutb(w_n7167_0[1]),.din(n7167));
	jspl jspl_w_n7168_0(.douta(w_n7168_0[0]),.doutb(w_n7168_0[1]),.din(n7168));
	jspl3 jspl3_w_n7169_0(.douta(w_n7169_0[0]),.doutb(w_n7169_0[1]),.doutc(w_n7169_0[2]),.din(n7169));
	jspl jspl_w_n7170_0(.douta(w_n7170_0[0]),.doutb(w_n7170_0[1]),.din(n7170));
	jspl jspl_w_n7174_0(.douta(w_n7174_0[0]),.doutb(w_n7174_0[1]),.din(n7174));
	jspl jspl_w_n7180_0(.douta(w_n7180_0[0]),.doutb(w_n7180_0[1]),.din(n7180));
	jspl jspl_w_n7181_0(.douta(w_n7181_0[0]),.doutb(w_n7181_0[1]),.din(n7181));
	jspl jspl_w_n7183_0(.douta(w_n7183_0[0]),.doutb(w_n7183_0[1]),.din(n7183));
	jspl jspl_w_n7185_0(.douta(w_n7185_0[0]),.doutb(w_n7185_0[1]),.din(n7185));
	jspl jspl_w_n7188_0(.douta(w_n7188_0[0]),.doutb(w_n7188_0[1]),.din(n7188));
	jspl jspl_w_n7194_0(.douta(w_n7194_0[0]),.doutb(w_n7194_0[1]),.din(n7194));
	jspl jspl_w_n7196_0(.douta(w_n7196_0[0]),.doutb(w_n7196_0[1]),.din(n7196));
	jspl3 jspl3_w_n7197_0(.douta(w_n7197_0[0]),.doutb(w_n7197_0[1]),.doutc(w_n7197_0[2]),.din(n7197));
	jspl jspl_w_n7201_0(.douta(w_n7201_0[0]),.doutb(w_n7201_0[1]),.din(n7201));
	jspl jspl_w_n7202_0(.douta(w_n7202_0[0]),.doutb(w_n7202_0[1]),.din(n7202));
	jspl3 jspl3_w_n7203_0(.douta(w_n7203_0[0]),.doutb(w_n7203_0[1]),.doutc(w_n7203_0[2]),.din(n7203));
	jspl jspl_w_n7205_0(.douta(w_n7205_0[0]),.doutb(w_n7205_0[1]),.din(n7205));
	jspl jspl_w_n7210_0(.douta(w_n7210_0[0]),.doutb(w_n7210_0[1]),.din(n7210));
	jspl jspl_w_n7212_0(.douta(w_n7212_0[0]),.doutb(w_n7212_0[1]),.din(n7212));
	jspl jspl_w_n7213_0(.douta(w_n7213_0[0]),.doutb(w_n7213_0[1]),.din(n7213));
	jspl3 jspl3_w_n7214_0(.douta(w_n7214_0[0]),.doutb(w_n7214_0[1]),.doutc(w_n7214_0[2]),.din(n7214));
	jspl jspl_w_n7215_0(.douta(w_n7215_0[0]),.doutb(w_n7215_0[1]),.din(n7215));
	jspl jspl_w_n7219_0(.douta(w_n7219_0[0]),.doutb(w_n7219_0[1]),.din(n7219));
	jspl jspl_w_n7225_0(.douta(w_n7225_0[0]),.doutb(w_n7225_0[1]),.din(n7225));
	jspl jspl_w_n7226_0(.douta(w_n7226_0[0]),.doutb(w_n7226_0[1]),.din(n7226));
	jspl jspl_w_n7228_0(.douta(w_n7228_0[0]),.doutb(w_n7228_0[1]),.din(n7228));
	jspl jspl_w_n7230_0(.douta(w_n7230_0[0]),.doutb(w_n7230_0[1]),.din(n7230));
	jspl jspl_w_n7233_0(.douta(w_n7233_0[0]),.doutb(w_n7233_0[1]),.din(n7233));
	jspl jspl_w_n7239_0(.douta(w_n7239_0[0]),.doutb(w_n7239_0[1]),.din(n7239));
	jspl3 jspl3_w_n7241_0(.douta(w_n7241_0[0]),.doutb(w_n7241_0[1]),.doutc(w_n7241_0[2]),.din(n7241));
	jspl3 jspl3_w_n7241_1(.douta(w_n7241_1[0]),.doutb(w_n7241_1[1]),.doutc(w_n7241_1[2]),.din(w_n7241_0[0]));
	jspl jspl_w_n7244_0(.douta(w_n7244_0[0]),.doutb(w_n7244_0[1]),.din(n7244));
	jspl3 jspl3_w_n7245_0(.douta(w_n7245_0[0]),.doutb(w_n7245_0[1]),.doutc(w_n7245_0[2]),.din(n7245));
	jspl jspl_w_n7246_0(.douta(w_n7246_0[0]),.doutb(w_n7246_0[1]),.din(n7246));
	jspl jspl_w_n7252_0(.douta(w_n7252_0[0]),.doutb(w_n7252_0[1]),.din(n7252));
	jspl3 jspl3_w_n7253_0(.douta(w_n7253_0[0]),.doutb(w_n7253_0[1]),.doutc(w_n7253_0[2]),.din(n7253));
	jspl jspl_w_n7254_0(.douta(w_n7254_0[0]),.doutb(w_n7254_0[1]),.din(n7254));
	jspl jspl_w_n7259_0(.douta(w_n7259_0[0]),.doutb(w_n7259_0[1]),.din(n7259));
	jspl3 jspl3_w_n7260_0(.douta(w_n7260_0[0]),.doutb(w_n7260_0[1]),.doutc(w_n7260_0[2]),.din(n7260));
	jspl3 jspl3_w_n7260_1(.douta(w_n7260_1[0]),.doutb(w_n7260_1[1]),.doutc(w_n7260_1[2]),.din(w_n7260_0[0]));
	jspl3 jspl3_w_n7260_2(.douta(w_n7260_2[0]),.doutb(w_n7260_2[1]),.doutc(w_n7260_2[2]),.din(w_n7260_0[1]));
	jspl3 jspl3_w_n7260_3(.douta(w_n7260_3[0]),.doutb(w_n7260_3[1]),.doutc(w_n7260_3[2]),.din(w_n7260_0[2]));
	jspl3 jspl3_w_n7260_4(.douta(w_n7260_4[0]),.doutb(w_n7260_4[1]),.doutc(w_n7260_4[2]),.din(w_n7260_1[0]));
	jspl3 jspl3_w_n7260_5(.douta(w_n7260_5[0]),.doutb(w_n7260_5[1]),.doutc(w_n7260_5[2]),.din(w_n7260_1[1]));
	jspl3 jspl3_w_n7260_6(.douta(w_n7260_6[0]),.doutb(w_n7260_6[1]),.doutc(w_n7260_6[2]),.din(w_n7260_1[2]));
	jspl3 jspl3_w_n7260_7(.douta(w_n7260_7[0]),.doutb(w_n7260_7[1]),.doutc(w_n7260_7[2]),.din(w_n7260_2[0]));
	jspl3 jspl3_w_n7260_8(.douta(w_n7260_8[0]),.doutb(w_n7260_8[1]),.doutc(w_n7260_8[2]),.din(w_n7260_2[1]));
	jspl3 jspl3_w_n7260_9(.douta(w_n7260_9[0]),.doutb(w_n7260_9[1]),.doutc(w_n7260_9[2]),.din(w_n7260_2[2]));
	jspl3 jspl3_w_n7260_10(.douta(w_n7260_10[0]),.doutb(w_n7260_10[1]),.doutc(w_n7260_10[2]),.din(w_n7260_3[0]));
	jspl3 jspl3_w_n7260_11(.douta(w_n7260_11[0]),.doutb(w_n7260_11[1]),.doutc(w_n7260_11[2]),.din(w_n7260_3[1]));
	jspl3 jspl3_w_n7260_12(.douta(w_n7260_12[0]),.doutb(w_n7260_12[1]),.doutc(w_n7260_12[2]),.din(w_n7260_3[2]));
	jspl3 jspl3_w_n7260_13(.douta(w_n7260_13[0]),.doutb(w_n7260_13[1]),.doutc(w_n7260_13[2]),.din(w_n7260_4[0]));
	jspl3 jspl3_w_n7260_14(.douta(w_n7260_14[0]),.doutb(w_n7260_14[1]),.doutc(w_n7260_14[2]),.din(w_n7260_4[1]));
	jspl3 jspl3_w_n7260_15(.douta(w_n7260_15[0]),.doutb(w_n7260_15[1]),.doutc(w_n7260_15[2]),.din(w_n7260_4[2]));
	jspl3 jspl3_w_n7260_16(.douta(w_n7260_16[0]),.doutb(w_n7260_16[1]),.doutc(w_n7260_16[2]),.din(w_n7260_5[0]));
	jspl3 jspl3_w_n7260_17(.douta(w_n7260_17[0]),.doutb(w_n7260_17[1]),.doutc(w_n7260_17[2]),.din(w_n7260_5[1]));
	jspl jspl_w_n7260_18(.douta(w_n7260_18[0]),.doutb(w_n7260_18[1]),.din(w_n7260_5[2]));
	jspl3 jspl3_w_n7265_0(.douta(w_n7265_0[0]),.doutb(w_n7265_0[1]),.doutc(w_n7265_0[2]),.din(n7265));
	jspl3 jspl3_w_n7265_1(.douta(w_n7265_1[0]),.doutb(w_n7265_1[1]),.doutc(w_n7265_1[2]),.din(w_n7265_0[0]));
	jspl3 jspl3_w_n7265_2(.douta(w_n7265_2[0]),.doutb(w_n7265_2[1]),.doutc(w_n7265_2[2]),.din(w_n7265_0[1]));
	jspl3 jspl3_w_n7265_3(.douta(w_n7265_3[0]),.doutb(w_n7265_3[1]),.doutc(w_n7265_3[2]),.din(w_n7265_0[2]));
	jspl3 jspl3_w_n7265_4(.douta(w_n7265_4[0]),.doutb(w_n7265_4[1]),.doutc(w_n7265_4[2]),.din(w_n7265_1[0]));
	jspl3 jspl3_w_n7265_5(.douta(w_n7265_5[0]),.doutb(w_n7265_5[1]),.doutc(w_n7265_5[2]),.din(w_n7265_1[1]));
	jspl3 jspl3_w_n7265_6(.douta(w_n7265_6[0]),.doutb(w_n7265_6[1]),.doutc(w_n7265_6[2]),.din(w_n7265_1[2]));
	jspl3 jspl3_w_n7265_7(.douta(w_n7265_7[0]),.doutb(w_n7265_7[1]),.doutc(w_n7265_7[2]),.din(w_n7265_2[0]));
	jspl3 jspl3_w_n7265_8(.douta(w_n7265_8[0]),.doutb(w_n7265_8[1]),.doutc(w_n7265_8[2]),.din(w_n7265_2[1]));
	jspl3 jspl3_w_n7265_9(.douta(w_n7265_9[0]),.doutb(w_n7265_9[1]),.doutc(w_n7265_9[2]),.din(w_n7265_2[2]));
	jspl3 jspl3_w_n7265_10(.douta(w_n7265_10[0]),.doutb(w_n7265_10[1]),.doutc(w_n7265_10[2]),.din(w_n7265_3[0]));
	jspl3 jspl3_w_n7265_11(.douta(w_n7265_11[0]),.doutb(w_n7265_11[1]),.doutc(w_n7265_11[2]),.din(w_n7265_3[1]));
	jspl3 jspl3_w_n7265_12(.douta(w_n7265_12[0]),.doutb(w_n7265_12[1]),.doutc(w_n7265_12[2]),.din(w_n7265_3[2]));
	jspl3 jspl3_w_n7265_13(.douta(w_n7265_13[0]),.doutb(w_n7265_13[1]),.doutc(w_n7265_13[2]),.din(w_n7265_4[0]));
	jspl3 jspl3_w_n7265_14(.douta(w_n7265_14[0]),.doutb(w_n7265_14[1]),.doutc(w_n7265_14[2]),.din(w_n7265_4[1]));
	jspl3 jspl3_w_n7265_15(.douta(w_n7265_15[0]),.doutb(w_n7265_15[1]),.doutc(w_n7265_15[2]),.din(w_n7265_4[2]));
	jspl3 jspl3_w_n7265_16(.douta(w_n7265_16[0]),.doutb(w_n7265_16[1]),.doutc(w_n7265_16[2]),.din(w_n7265_5[0]));
	jspl3 jspl3_w_n7265_17(.douta(w_n7265_17[0]),.doutb(w_n7265_17[1]),.doutc(w_n7265_17[2]),.din(w_n7265_5[1]));
	jspl3 jspl3_w_n7265_18(.douta(w_n7265_18[0]),.doutb(w_n7265_18[1]),.doutc(w_n7265_18[2]),.din(w_n7265_5[2]));
	jspl3 jspl3_w_n7265_19(.douta(w_n7265_19[0]),.doutb(w_n7265_19[1]),.doutc(w_n7265_19[2]),.din(w_n7265_6[0]));
	jspl3 jspl3_w_n7265_20(.douta(w_n7265_20[0]),.doutb(w_n7265_20[1]),.doutc(w_n7265_20[2]),.din(w_n7265_6[1]));
	jspl3 jspl3_w_n7265_21(.douta(w_n7265_21[0]),.doutb(w_n7265_21[1]),.doutc(w_n7265_21[2]),.din(w_n7265_6[2]));
	jspl3 jspl3_w_n7265_22(.douta(w_n7265_22[0]),.doutb(w_n7265_22[1]),.doutc(w_n7265_22[2]),.din(w_n7265_7[0]));
	jspl3 jspl3_w_n7265_23(.douta(w_n7265_23[0]),.doutb(w_n7265_23[1]),.doutc(w_n7265_23[2]),.din(w_n7265_7[1]));
	jspl3 jspl3_w_n7265_24(.douta(w_n7265_24[0]),.doutb(w_n7265_24[1]),.doutc(w_n7265_24[2]),.din(w_n7265_7[2]));
	jspl3 jspl3_w_n7265_25(.douta(w_n7265_25[0]),.doutb(w_n7265_25[1]),.doutc(w_n7265_25[2]),.din(w_n7265_8[0]));
	jspl3 jspl3_w_n7265_26(.douta(w_n7265_26[0]),.doutb(w_n7265_26[1]),.doutc(w_n7265_26[2]),.din(w_n7265_8[1]));
	jspl3 jspl3_w_n7265_27(.douta(w_n7265_27[0]),.doutb(w_n7265_27[1]),.doutc(w_n7265_27[2]),.din(w_n7265_8[2]));
	jspl jspl_w_n7265_28(.douta(w_n7265_28[0]),.doutb(w_n7265_28[1]),.din(w_n7265_9[0]));
	jspl jspl_w_n7269_0(.douta(w_n7269_0[0]),.doutb(w_n7269_0[1]),.din(n7269));
	jspl3 jspl3_w_n7271_0(.douta(w_n7271_0[0]),.doutb(w_n7271_0[1]),.doutc(w_n7271_0[2]),.din(n7271));
	jspl jspl_w_n7271_1(.douta(w_n7271_1[0]),.doutb(w_n7271_1[1]),.din(w_n7271_0[0]));
	jspl3 jspl3_w_n7272_0(.douta(w_n7272_0[0]),.doutb(w_n7272_0[1]),.doutc(w_n7272_0[2]),.din(n7272));
	jspl3 jspl3_w_n7276_0(.douta(w_n7276_0[0]),.doutb(w_n7276_0[1]),.doutc(w_n7276_0[2]),.din(n7276));
	jspl jspl_w_n7277_0(.douta(w_n7277_0[0]),.doutb(w_n7277_0[1]),.din(n7277));
	jspl jspl_w_n7278_0(.douta(w_n7278_0[0]),.doutb(w_n7278_0[1]),.din(n7278));
	jspl jspl_w_n7279_0(.douta(w_n7279_0[0]),.doutb(w_n7279_0[1]),.din(n7279));
	jspl jspl_w_n7281_0(.douta(w_n7281_0[0]),.doutb(w_n7281_0[1]),.din(n7281));
	jspl jspl_w_n7283_0(.douta(w_n7283_0[0]),.doutb(w_n7283_0[1]),.din(n7283));
	jspl jspl_w_n7285_0(.douta(w_n7285_0[0]),.doutb(w_n7285_0[1]),.din(n7285));
	jspl jspl_w_n7288_0(.douta(w_n7288_0[0]),.doutb(w_n7288_0[1]),.din(n7288));
	jspl jspl_w_n7293_0(.douta(w_n7293_0[0]),.doutb(w_n7293_0[1]),.din(n7293));
	jspl3 jspl3_w_n7295_0(.douta(w_n7295_0[0]),.doutb(w_n7295_0[1]),.doutc(w_n7295_0[2]),.din(n7295));
	jspl jspl_w_n7296_0(.douta(w_n7296_0[0]),.doutb(w_n7296_0[1]),.din(n7296));
	jspl jspl_w_n7300_0(.douta(w_n7300_0[0]),.doutb(w_n7300_0[1]),.din(n7300));
	jspl jspl_w_n7301_0(.douta(w_n7301_0[0]),.doutb(w_n7301_0[1]),.din(n7301));
	jspl jspl_w_n7303_0(.douta(w_n7303_0[0]),.doutb(w_n7303_0[1]),.din(n7303));
	jspl jspl_w_n7307_0(.douta(w_n7307_0[0]),.doutb(w_n7307_0[1]),.din(n7307));
	jspl jspl_w_n7309_0(.douta(w_n7309_0[0]),.doutb(w_n7309_0[1]),.din(n7309));
	jspl jspl_w_n7310_0(.douta(w_n7310_0[0]),.doutb(w_n7310_0[1]),.din(n7310));
	jspl3 jspl3_w_n7311_0(.douta(w_n7311_0[0]),.doutb(w_n7311_0[1]),.doutc(w_n7311_0[2]),.din(n7311));
	jspl jspl_w_n7312_0(.douta(w_n7312_0[0]),.doutb(w_n7312_0[1]),.din(n7312));
	jspl jspl_w_n7316_0(.douta(w_n7316_0[0]),.doutb(w_n7316_0[1]),.din(n7316));
	jspl jspl_w_n7318_0(.douta(w_n7318_0[0]),.doutb(w_n7318_0[1]),.din(n7318));
	jspl jspl_w_n7320_0(.douta(w_n7320_0[0]),.doutb(w_n7320_0[1]),.din(n7320));
	jspl jspl_w_n7322_0(.douta(w_n7322_0[0]),.doutb(w_n7322_0[1]),.din(n7322));
	jspl jspl_w_n7325_0(.douta(w_n7325_0[0]),.doutb(w_n7325_0[1]),.din(n7325));
	jspl jspl_w_n7331_0(.douta(w_n7331_0[0]),.doutb(w_n7331_0[1]),.din(n7331));
	jspl3 jspl3_w_n7333_0(.douta(w_n7333_0[0]),.doutb(w_n7333_0[1]),.doutc(w_n7333_0[2]),.din(n7333));
	jspl jspl_w_n7334_0(.douta(w_n7334_0[0]),.doutb(w_n7334_0[1]),.din(n7334));
	jspl jspl_w_n7339_0(.douta(w_n7339_0[0]),.doutb(w_n7339_0[1]),.din(n7339));
	jspl jspl_w_n7341_0(.douta(w_n7341_0[0]),.doutb(w_n7341_0[1]),.din(n7341));
	jspl jspl_w_n7343_0(.douta(w_n7343_0[0]),.doutb(w_n7343_0[1]),.din(n7343));
	jspl jspl_w_n7345_0(.douta(w_n7345_0[0]),.doutb(w_n7345_0[1]),.din(n7345));
	jspl jspl_w_n7347_0(.douta(w_n7347_0[0]),.doutb(w_n7347_0[1]),.din(n7347));
	jspl jspl_w_n7353_0(.douta(w_n7353_0[0]),.doutb(w_n7353_0[1]),.din(n7353));
	jspl3 jspl3_w_n7355_0(.douta(w_n7355_0[0]),.doutb(w_n7355_0[1]),.doutc(w_n7355_0[2]),.din(n7355));
	jspl jspl_w_n7356_0(.douta(w_n7356_0[0]),.doutb(w_n7356_0[1]),.din(n7356));
	jspl jspl_w_n7358_0(.douta(w_n7358_0[0]),.doutb(w_n7358_0[1]),.din(n7358));
	jspl jspl_w_n7360_0(.douta(w_n7360_0[0]),.doutb(w_n7360_0[1]),.din(n7360));
	jspl jspl_w_n7364_0(.douta(w_n7364_0[0]),.doutb(w_n7364_0[1]),.din(n7364));
	jspl jspl_w_n7366_0(.douta(w_n7366_0[0]),.doutb(w_n7366_0[1]),.din(n7366));
	jspl jspl_w_n7367_0(.douta(w_n7367_0[0]),.doutb(w_n7367_0[1]),.din(n7367));
	jspl jspl_w_n7368_0(.douta(w_n7368_0[0]),.doutb(w_n7368_0[1]),.din(n7368));
	jspl3 jspl3_w_n7369_0(.douta(w_n7369_0[0]),.doutb(w_n7369_0[1]),.doutc(w_n7369_0[2]),.din(n7369));
	jspl jspl_w_n7372_0(.douta(w_n7372_0[0]),.doutb(w_n7372_0[1]),.din(n7372));
	jspl jspl_w_n7373_0(.douta(w_n7373_0[0]),.doutb(w_n7373_0[1]),.din(n7373));
	jspl3 jspl3_w_n7374_0(.douta(w_n7374_0[0]),.doutb(w_n7374_0[1]),.doutc(w_n7374_0[2]),.din(n7374));
	jspl jspl_w_n7376_0(.douta(w_n7376_0[0]),.doutb(w_n7376_0[1]),.din(n7376));
	jspl jspl_w_n7380_0(.douta(w_n7380_0[0]),.doutb(w_n7380_0[1]),.din(n7380));
	jspl jspl_w_n7382_0(.douta(w_n7382_0[0]),.doutb(w_n7382_0[1]),.din(n7382));
	jspl jspl_w_n7383_0(.douta(w_n7383_0[0]),.doutb(w_n7383_0[1]),.din(n7383));
	jspl3 jspl3_w_n7384_0(.douta(w_n7384_0[0]),.doutb(w_n7384_0[1]),.doutc(w_n7384_0[2]),.din(n7384));
	jspl jspl_w_n7385_0(.douta(w_n7385_0[0]),.doutb(w_n7385_0[1]),.din(n7385));
	jspl jspl_w_n7388_0(.douta(w_n7388_0[0]),.doutb(w_n7388_0[1]),.din(n7388));
	jspl jspl_w_n7394_0(.douta(w_n7394_0[0]),.doutb(w_n7394_0[1]),.din(n7394));
	jspl jspl_w_n7395_0(.douta(w_n7395_0[0]),.doutb(w_n7395_0[1]),.din(n7395));
	jspl jspl_w_n7397_0(.douta(w_n7397_0[0]),.doutb(w_n7397_0[1]),.din(n7397));
	jspl jspl_w_n7399_0(.douta(w_n7399_0[0]),.doutb(w_n7399_0[1]),.din(n7399));
	jspl jspl_w_n7401_0(.douta(w_n7401_0[0]),.doutb(w_n7401_0[1]),.din(n7401));
	jspl jspl_w_n7407_0(.douta(w_n7407_0[0]),.doutb(w_n7407_0[1]),.din(n7407));
	jspl jspl_w_n7409_0(.douta(w_n7409_0[0]),.doutb(w_n7409_0[1]),.din(n7409));
	jspl3 jspl3_w_n7410_0(.douta(w_n7410_0[0]),.doutb(w_n7410_0[1]),.doutc(w_n7410_0[2]),.din(n7410));
	jspl jspl_w_n7413_0(.douta(w_n7413_0[0]),.doutb(w_n7413_0[1]),.din(n7413));
	jspl jspl_w_n7414_0(.douta(w_n7414_0[0]),.doutb(w_n7414_0[1]),.din(n7414));
	jspl3 jspl3_w_n7415_0(.douta(w_n7415_0[0]),.doutb(w_n7415_0[1]),.doutc(w_n7415_0[2]),.din(n7415));
	jspl jspl_w_n7417_0(.douta(w_n7417_0[0]),.doutb(w_n7417_0[1]),.din(n7417));
	jspl jspl_w_n7421_0(.douta(w_n7421_0[0]),.doutb(w_n7421_0[1]),.din(n7421));
	jspl jspl_w_n7423_0(.douta(w_n7423_0[0]),.doutb(w_n7423_0[1]),.din(n7423));
	jspl jspl_w_n7424_0(.douta(w_n7424_0[0]),.doutb(w_n7424_0[1]),.din(n7424));
	jspl3 jspl3_w_n7425_0(.douta(w_n7425_0[0]),.doutb(w_n7425_0[1]),.doutc(w_n7425_0[2]),.din(n7425));
	jspl jspl_w_n7426_0(.douta(w_n7426_0[0]),.doutb(w_n7426_0[1]),.din(n7426));
	jspl jspl_w_n7429_0(.douta(w_n7429_0[0]),.doutb(w_n7429_0[1]),.din(n7429));
	jspl jspl_w_n7435_0(.douta(w_n7435_0[0]),.doutb(w_n7435_0[1]),.din(n7435));
	jspl jspl_w_n7436_0(.douta(w_n7436_0[0]),.doutb(w_n7436_0[1]),.din(n7436));
	jspl jspl_w_n7438_0(.douta(w_n7438_0[0]),.doutb(w_n7438_0[1]),.din(n7438));
	jspl jspl_w_n7440_0(.douta(w_n7440_0[0]),.doutb(w_n7440_0[1]),.din(n7440));
	jspl jspl_w_n7442_0(.douta(w_n7442_0[0]),.doutb(w_n7442_0[1]),.din(n7442));
	jspl jspl_w_n7448_0(.douta(w_n7448_0[0]),.doutb(w_n7448_0[1]),.din(n7448));
	jspl jspl_w_n7450_0(.douta(w_n7450_0[0]),.doutb(w_n7450_0[1]),.din(n7450));
	jspl3 jspl3_w_n7451_0(.douta(w_n7451_0[0]),.doutb(w_n7451_0[1]),.doutc(w_n7451_0[2]),.din(n7451));
	jspl jspl_w_n7454_0(.douta(w_n7454_0[0]),.doutb(w_n7454_0[1]),.din(n7454));
	jspl jspl_w_n7455_0(.douta(w_n7455_0[0]),.doutb(w_n7455_0[1]),.din(n7455));
	jspl3 jspl3_w_n7456_0(.douta(w_n7456_0[0]),.doutb(w_n7456_0[1]),.doutc(w_n7456_0[2]),.din(n7456));
	jspl jspl_w_n7458_0(.douta(w_n7458_0[0]),.doutb(w_n7458_0[1]),.din(n7458));
	jspl jspl_w_n7462_0(.douta(w_n7462_0[0]),.doutb(w_n7462_0[1]),.din(n7462));
	jspl jspl_w_n7464_0(.douta(w_n7464_0[0]),.doutb(w_n7464_0[1]),.din(n7464));
	jspl jspl_w_n7465_0(.douta(w_n7465_0[0]),.doutb(w_n7465_0[1]),.din(n7465));
	jspl3 jspl3_w_n7466_0(.douta(w_n7466_0[0]),.doutb(w_n7466_0[1]),.doutc(w_n7466_0[2]),.din(n7466));
	jspl jspl_w_n7467_0(.douta(w_n7467_0[0]),.doutb(w_n7467_0[1]),.din(n7467));
	jspl jspl_w_n7470_0(.douta(w_n7470_0[0]),.doutb(w_n7470_0[1]),.din(n7470));
	jspl jspl_w_n7476_0(.douta(w_n7476_0[0]),.doutb(w_n7476_0[1]),.din(n7476));
	jspl jspl_w_n7477_0(.douta(w_n7477_0[0]),.doutb(w_n7477_0[1]),.din(n7477));
	jspl jspl_w_n7479_0(.douta(w_n7479_0[0]),.doutb(w_n7479_0[1]),.din(n7479));
	jspl jspl_w_n7481_0(.douta(w_n7481_0[0]),.doutb(w_n7481_0[1]),.din(n7481));
	jspl jspl_w_n7483_0(.douta(w_n7483_0[0]),.doutb(w_n7483_0[1]),.din(n7483));
	jspl jspl_w_n7489_0(.douta(w_n7489_0[0]),.doutb(w_n7489_0[1]),.din(n7489));
	jspl jspl_w_n7491_0(.douta(w_n7491_0[0]),.doutb(w_n7491_0[1]),.din(n7491));
	jspl3 jspl3_w_n7492_0(.douta(w_n7492_0[0]),.doutb(w_n7492_0[1]),.doutc(w_n7492_0[2]),.din(n7492));
	jspl jspl_w_n7495_0(.douta(w_n7495_0[0]),.doutb(w_n7495_0[1]),.din(n7495));
	jspl jspl_w_n7496_0(.douta(w_n7496_0[0]),.doutb(w_n7496_0[1]),.din(n7496));
	jspl3 jspl3_w_n7497_0(.douta(w_n7497_0[0]),.doutb(w_n7497_0[1]),.doutc(w_n7497_0[2]),.din(n7497));
	jspl jspl_w_n7499_0(.douta(w_n7499_0[0]),.doutb(w_n7499_0[1]),.din(n7499));
	jspl jspl_w_n7503_0(.douta(w_n7503_0[0]),.doutb(w_n7503_0[1]),.din(n7503));
	jspl jspl_w_n7505_0(.douta(w_n7505_0[0]),.doutb(w_n7505_0[1]),.din(n7505));
	jspl jspl_w_n7506_0(.douta(w_n7506_0[0]),.doutb(w_n7506_0[1]),.din(n7506));
	jspl3 jspl3_w_n7507_0(.douta(w_n7507_0[0]),.doutb(w_n7507_0[1]),.doutc(w_n7507_0[2]),.din(n7507));
	jspl jspl_w_n7508_0(.douta(w_n7508_0[0]),.doutb(w_n7508_0[1]),.din(n7508));
	jspl jspl_w_n7511_0(.douta(w_n7511_0[0]),.doutb(w_n7511_0[1]),.din(n7511));
	jspl jspl_w_n7517_0(.douta(w_n7517_0[0]),.doutb(w_n7517_0[1]),.din(n7517));
	jspl jspl_w_n7518_0(.douta(w_n7518_0[0]),.doutb(w_n7518_0[1]),.din(n7518));
	jspl jspl_w_n7520_0(.douta(w_n7520_0[0]),.doutb(w_n7520_0[1]),.din(n7520));
	jspl jspl_w_n7522_0(.douta(w_n7522_0[0]),.doutb(w_n7522_0[1]),.din(n7522));
	jspl jspl_w_n7524_0(.douta(w_n7524_0[0]),.doutb(w_n7524_0[1]),.din(n7524));
	jspl jspl_w_n7530_0(.douta(w_n7530_0[0]),.doutb(w_n7530_0[1]),.din(n7530));
	jspl jspl_w_n7532_0(.douta(w_n7532_0[0]),.doutb(w_n7532_0[1]),.din(n7532));
	jspl3 jspl3_w_n7533_0(.douta(w_n7533_0[0]),.doutb(w_n7533_0[1]),.doutc(w_n7533_0[2]),.din(n7533));
	jspl jspl_w_n7536_0(.douta(w_n7536_0[0]),.doutb(w_n7536_0[1]),.din(n7536));
	jspl jspl_w_n7537_0(.douta(w_n7537_0[0]),.doutb(w_n7537_0[1]),.din(n7537));
	jspl3 jspl3_w_n7538_0(.douta(w_n7538_0[0]),.doutb(w_n7538_0[1]),.doutc(w_n7538_0[2]),.din(n7538));
	jspl jspl_w_n7540_0(.douta(w_n7540_0[0]),.doutb(w_n7540_0[1]),.din(n7540));
	jspl jspl_w_n7544_0(.douta(w_n7544_0[0]),.doutb(w_n7544_0[1]),.din(n7544));
	jspl jspl_w_n7546_0(.douta(w_n7546_0[0]),.doutb(w_n7546_0[1]),.din(n7546));
	jspl jspl_w_n7547_0(.douta(w_n7547_0[0]),.doutb(w_n7547_0[1]),.din(n7547));
	jspl3 jspl3_w_n7548_0(.douta(w_n7548_0[0]),.doutb(w_n7548_0[1]),.doutc(w_n7548_0[2]),.din(n7548));
	jspl jspl_w_n7549_0(.douta(w_n7549_0[0]),.doutb(w_n7549_0[1]),.din(n7549));
	jspl jspl_w_n7552_0(.douta(w_n7552_0[0]),.doutb(w_n7552_0[1]),.din(n7552));
	jspl jspl_w_n7558_0(.douta(w_n7558_0[0]),.doutb(w_n7558_0[1]),.din(n7558));
	jspl jspl_w_n7559_0(.douta(w_n7559_0[0]),.doutb(w_n7559_0[1]),.din(n7559));
	jspl jspl_w_n7561_0(.douta(w_n7561_0[0]),.doutb(w_n7561_0[1]),.din(n7561));
	jspl jspl_w_n7563_0(.douta(w_n7563_0[0]),.doutb(w_n7563_0[1]),.din(n7563));
	jspl jspl_w_n7565_0(.douta(w_n7565_0[0]),.doutb(w_n7565_0[1]),.din(n7565));
	jspl jspl_w_n7571_0(.douta(w_n7571_0[0]),.doutb(w_n7571_0[1]),.din(n7571));
	jspl jspl_w_n7573_0(.douta(w_n7573_0[0]),.doutb(w_n7573_0[1]),.din(n7573));
	jspl3 jspl3_w_n7574_0(.douta(w_n7574_0[0]),.doutb(w_n7574_0[1]),.doutc(w_n7574_0[2]),.din(n7574));
	jspl jspl_w_n7577_0(.douta(w_n7577_0[0]),.doutb(w_n7577_0[1]),.din(n7577));
	jspl jspl_w_n7578_0(.douta(w_n7578_0[0]),.doutb(w_n7578_0[1]),.din(n7578));
	jspl3 jspl3_w_n7579_0(.douta(w_n7579_0[0]),.doutb(w_n7579_0[1]),.doutc(w_n7579_0[2]),.din(n7579));
	jspl jspl_w_n7581_0(.douta(w_n7581_0[0]),.doutb(w_n7581_0[1]),.din(n7581));
	jspl jspl_w_n7585_0(.douta(w_n7585_0[0]),.doutb(w_n7585_0[1]),.din(n7585));
	jspl jspl_w_n7587_0(.douta(w_n7587_0[0]),.doutb(w_n7587_0[1]),.din(n7587));
	jspl jspl_w_n7588_0(.douta(w_n7588_0[0]),.doutb(w_n7588_0[1]),.din(n7588));
	jspl3 jspl3_w_n7589_0(.douta(w_n7589_0[0]),.doutb(w_n7589_0[1]),.doutc(w_n7589_0[2]),.din(n7589));
	jspl jspl_w_n7590_0(.douta(w_n7590_0[0]),.doutb(w_n7590_0[1]),.din(n7590));
	jspl jspl_w_n7593_0(.douta(w_n7593_0[0]),.doutb(w_n7593_0[1]),.din(n7593));
	jspl jspl_w_n7599_0(.douta(w_n7599_0[0]),.doutb(w_n7599_0[1]),.din(n7599));
	jspl jspl_w_n7600_0(.douta(w_n7600_0[0]),.doutb(w_n7600_0[1]),.din(n7600));
	jspl jspl_w_n7602_0(.douta(w_n7602_0[0]),.doutb(w_n7602_0[1]),.din(n7602));
	jspl jspl_w_n7604_0(.douta(w_n7604_0[0]),.doutb(w_n7604_0[1]),.din(n7604));
	jspl jspl_w_n7606_0(.douta(w_n7606_0[0]),.doutb(w_n7606_0[1]),.din(n7606));
	jspl jspl_w_n7612_0(.douta(w_n7612_0[0]),.doutb(w_n7612_0[1]),.din(n7612));
	jspl3 jspl3_w_n7614_0(.douta(w_n7614_0[0]),.doutb(w_n7614_0[1]),.doutc(w_n7614_0[2]),.din(n7614));
	jspl jspl_w_n7619_0(.douta(w_n7619_0[0]),.doutb(w_n7619_0[1]),.din(n7619));
	jspl3 jspl3_w_n7621_0(.douta(w_n7621_0[0]),.doutb(w_n7621_0[1]),.doutc(w_n7621_0[2]),.din(n7621));
	jspl3 jspl3_w_n7625_0(.douta(w_n7625_0[0]),.doutb(w_n7625_0[1]),.doutc(w_n7625_0[2]),.din(n7625));
	jspl jspl_w_n7626_0(.douta(w_n7626_0[0]),.doutb(w_n7626_0[1]),.din(n7626));
	jspl jspl_w_n7631_0(.douta(w_n7631_0[0]),.doutb(w_n7631_0[1]),.din(n7631));
	jspl3 jspl3_w_n7632_0(.douta(w_n7632_0[0]),.doutb(w_n7632_0[1]),.doutc(w_n7632_0[2]),.din(n7632));
	jspl jspl_w_n7637_0(.douta(w_n7637_0[0]),.doutb(w_n7637_0[1]),.din(n7637));
	jspl jspl_w_n7645_0(.douta(w_n7645_0[0]),.doutb(w_n7645_0[1]),.din(n7645));
	jspl3 jspl3_w_n7647_0(.douta(w_n7647_0[0]),.doutb(w_n7647_0[1]),.doutc(w_n7647_0[2]),.din(n7647));
	jspl jspl_w_n7647_1(.douta(w_n7647_1[0]),.doutb(w_n7647_1[1]),.din(w_n7647_0[0]));
	jspl jspl_w_n7648_0(.douta(w_n7648_0[0]),.doutb(w_n7648_0[1]),.din(n7648));
	jspl3 jspl3_w_n7651_0(.douta(w_n7651_0[0]),.doutb(w_n7651_0[1]),.doutc(w_n7651_0[2]),.din(n7651));
	jspl jspl_w_n7652_0(.douta(w_n7652_0[0]),.doutb(w_n7652_0[1]),.din(n7652));
	jspl jspl_w_n7653_0(.douta(w_n7653_0[0]),.doutb(w_n7653_0[1]),.din(n7653));
	jspl jspl_w_n7654_0(.douta(w_n7654_0[0]),.doutb(w_n7654_0[1]),.din(n7654));
	jspl jspl_w_n7656_0(.douta(w_n7656_0[0]),.doutb(w_n7656_0[1]),.din(n7656));
	jspl jspl_w_n7658_0(.douta(w_n7658_0[0]),.doutb(w_n7658_0[1]),.din(n7658));
	jspl jspl_w_n7660_0(.douta(w_n7660_0[0]),.doutb(w_n7660_0[1]),.din(n7660));
	jspl jspl_w_n7669_0(.douta(w_n7669_0[0]),.doutb(w_n7669_0[1]),.din(n7669));
	jspl3 jspl3_w_n7671_0(.douta(w_n7671_0[0]),.doutb(w_n7671_0[1]),.doutc(w_n7671_0[2]),.din(n7671));
	jspl jspl_w_n7672_0(.douta(w_n7672_0[0]),.doutb(w_n7672_0[1]),.din(n7672));
	jspl jspl_w_n7676_0(.douta(w_n7676_0[0]),.doutb(w_n7676_0[1]),.din(n7676));
	jspl jspl_w_n7678_0(.douta(w_n7678_0[0]),.doutb(w_n7678_0[1]),.din(n7678));
	jspl jspl_w_n7680_0(.douta(w_n7680_0[0]),.doutb(w_n7680_0[1]),.din(n7680));
	jspl jspl_w_n7685_0(.douta(w_n7685_0[0]),.doutb(w_n7685_0[1]),.din(n7685));
	jspl jspl_w_n7687_0(.douta(w_n7687_0[0]),.doutb(w_n7687_0[1]),.din(n7687));
	jspl jspl_w_n7688_0(.douta(w_n7688_0[0]),.doutb(w_n7688_0[1]),.din(n7688));
	jspl3 jspl3_w_n7689_0(.douta(w_n7689_0[0]),.doutb(w_n7689_0[1]),.doutc(w_n7689_0[2]),.din(n7689));
	jspl jspl_w_n7690_0(.douta(w_n7690_0[0]),.doutb(w_n7690_0[1]),.din(n7690));
	jspl jspl_w_n7695_0(.douta(w_n7695_0[0]),.doutb(w_n7695_0[1]),.din(n7695));
	jspl jspl_w_n7696_0(.douta(w_n7696_0[0]),.doutb(w_n7696_0[1]),.din(n7696));
	jspl jspl_w_n7698_0(.douta(w_n7698_0[0]),.doutb(w_n7698_0[1]),.din(n7698));
	jspl jspl_w_n7700_0(.douta(w_n7700_0[0]),.doutb(w_n7700_0[1]),.din(n7700));
	jspl jspl_w_n7703_0(.douta(w_n7703_0[0]),.doutb(w_n7703_0[1]),.din(n7703));
	jspl jspl_w_n7709_0(.douta(w_n7709_0[0]),.doutb(w_n7709_0[1]),.din(n7709));
	jspl3 jspl3_w_n7711_0(.douta(w_n7711_0[0]),.doutb(w_n7711_0[1]),.doutc(w_n7711_0[2]),.din(n7711));
	jspl jspl_w_n7712_0(.douta(w_n7712_0[0]),.doutb(w_n7712_0[1]),.din(n7712));
	jspl jspl_w_n7716_0(.douta(w_n7716_0[0]),.doutb(w_n7716_0[1]),.din(n7716));
	jspl jspl_w_n7717_0(.douta(w_n7717_0[0]),.doutb(w_n7717_0[1]),.din(n7717));
	jspl jspl_w_n7719_0(.douta(w_n7719_0[0]),.doutb(w_n7719_0[1]),.din(n7719));
	jspl jspl_w_n7724_0(.douta(w_n7724_0[0]),.doutb(w_n7724_0[1]),.din(n7724));
	jspl jspl_w_n7726_0(.douta(w_n7726_0[0]),.doutb(w_n7726_0[1]),.din(n7726));
	jspl jspl_w_n7727_0(.douta(w_n7727_0[0]),.doutb(w_n7727_0[1]),.din(n7727));
	jspl3 jspl3_w_n7728_0(.douta(w_n7728_0[0]),.doutb(w_n7728_0[1]),.doutc(w_n7728_0[2]),.din(n7728));
	jspl jspl_w_n7729_0(.douta(w_n7729_0[0]),.doutb(w_n7729_0[1]),.din(n7729));
	jspl jspl_w_n7733_0(.douta(w_n7733_0[0]),.doutb(w_n7733_0[1]),.din(n7733));
	jspl jspl_w_n7734_0(.douta(w_n7734_0[0]),.doutb(w_n7734_0[1]),.din(n7734));
	jspl jspl_w_n7736_0(.douta(w_n7736_0[0]),.doutb(w_n7736_0[1]),.din(n7736));
	jspl jspl_w_n7741_0(.douta(w_n7741_0[0]),.doutb(w_n7741_0[1]),.din(n7741));
	jspl jspl_w_n7743_0(.douta(w_n7743_0[0]),.doutb(w_n7743_0[1]),.din(n7743));
	jspl jspl_w_n7744_0(.douta(w_n7744_0[0]),.doutb(w_n7744_0[1]),.din(n7744));
	jspl3 jspl3_w_n7745_0(.douta(w_n7745_0[0]),.doutb(w_n7745_0[1]),.doutc(w_n7745_0[2]),.din(n7745));
	jspl jspl_w_n7746_0(.douta(w_n7746_0[0]),.doutb(w_n7746_0[1]),.din(n7746));
	jspl jspl_w_n7748_0(.douta(w_n7748_0[0]),.doutb(w_n7748_0[1]),.din(n7748));
	jspl jspl_w_n7750_0(.douta(w_n7750_0[0]),.doutb(w_n7750_0[1]),.din(n7750));
	jspl jspl_w_n7752_0(.douta(w_n7752_0[0]),.doutb(w_n7752_0[1]),.din(n7752));
	jspl jspl_w_n7755_0(.douta(w_n7755_0[0]),.doutb(w_n7755_0[1]),.din(n7755));
	jspl jspl_w_n7761_0(.douta(w_n7761_0[0]),.doutb(w_n7761_0[1]),.din(n7761));
	jspl3 jspl3_w_n7763_0(.douta(w_n7763_0[0]),.doutb(w_n7763_0[1]),.doutc(w_n7763_0[2]),.din(n7763));
	jspl jspl_w_n7764_0(.douta(w_n7764_0[0]),.doutb(w_n7764_0[1]),.din(n7764));
	jspl jspl_w_n7768_0(.douta(w_n7768_0[0]),.doutb(w_n7768_0[1]),.din(n7768));
	jspl jspl_w_n7774_0(.douta(w_n7774_0[0]),.doutb(w_n7774_0[1]),.din(n7774));
	jspl jspl_w_n7775_0(.douta(w_n7775_0[0]),.doutb(w_n7775_0[1]),.din(n7775));
	jspl jspl_w_n7777_0(.douta(w_n7777_0[0]),.doutb(w_n7777_0[1]),.din(n7777));
	jspl jspl_w_n7779_0(.douta(w_n7779_0[0]),.doutb(w_n7779_0[1]),.din(n7779));
	jspl jspl_w_n7782_0(.douta(w_n7782_0[0]),.doutb(w_n7782_0[1]),.din(n7782));
	jspl jspl_w_n7788_0(.douta(w_n7788_0[0]),.doutb(w_n7788_0[1]),.din(n7788));
	jspl jspl_w_n7790_0(.douta(w_n7790_0[0]),.doutb(w_n7790_0[1]),.din(n7790));
	jspl3 jspl3_w_n7791_0(.douta(w_n7791_0[0]),.doutb(w_n7791_0[1]),.doutc(w_n7791_0[2]),.din(n7791));
	jspl jspl_w_n7795_0(.douta(w_n7795_0[0]),.doutb(w_n7795_0[1]),.din(n7795));
	jspl jspl_w_n7796_0(.douta(w_n7796_0[0]),.doutb(w_n7796_0[1]),.din(n7796));
	jspl3 jspl3_w_n7797_0(.douta(w_n7797_0[0]),.doutb(w_n7797_0[1]),.doutc(w_n7797_0[2]),.din(n7797));
	jspl jspl_w_n7799_0(.douta(w_n7799_0[0]),.doutb(w_n7799_0[1]),.din(n7799));
	jspl jspl_w_n7804_0(.douta(w_n7804_0[0]),.doutb(w_n7804_0[1]),.din(n7804));
	jspl jspl_w_n7806_0(.douta(w_n7806_0[0]),.doutb(w_n7806_0[1]),.din(n7806));
	jspl jspl_w_n7807_0(.douta(w_n7807_0[0]),.doutb(w_n7807_0[1]),.din(n7807));
	jspl3 jspl3_w_n7808_0(.douta(w_n7808_0[0]),.doutb(w_n7808_0[1]),.doutc(w_n7808_0[2]),.din(n7808));
	jspl jspl_w_n7809_0(.douta(w_n7809_0[0]),.doutb(w_n7809_0[1]),.din(n7809));
	jspl jspl_w_n7813_0(.douta(w_n7813_0[0]),.doutb(w_n7813_0[1]),.din(n7813));
	jspl jspl_w_n7819_0(.douta(w_n7819_0[0]),.doutb(w_n7819_0[1]),.din(n7819));
	jspl jspl_w_n7820_0(.douta(w_n7820_0[0]),.doutb(w_n7820_0[1]),.din(n7820));
	jspl jspl_w_n7822_0(.douta(w_n7822_0[0]),.doutb(w_n7822_0[1]),.din(n7822));
	jspl jspl_w_n7824_0(.douta(w_n7824_0[0]),.doutb(w_n7824_0[1]),.din(n7824));
	jspl jspl_w_n7827_0(.douta(w_n7827_0[0]),.doutb(w_n7827_0[1]),.din(n7827));
	jspl jspl_w_n7833_0(.douta(w_n7833_0[0]),.doutb(w_n7833_0[1]),.din(n7833));
	jspl jspl_w_n7835_0(.douta(w_n7835_0[0]),.doutb(w_n7835_0[1]),.din(n7835));
	jspl3 jspl3_w_n7836_0(.douta(w_n7836_0[0]),.doutb(w_n7836_0[1]),.doutc(w_n7836_0[2]),.din(n7836));
	jspl jspl_w_n7840_0(.douta(w_n7840_0[0]),.doutb(w_n7840_0[1]),.din(n7840));
	jspl jspl_w_n7841_0(.douta(w_n7841_0[0]),.doutb(w_n7841_0[1]),.din(n7841));
	jspl3 jspl3_w_n7842_0(.douta(w_n7842_0[0]),.doutb(w_n7842_0[1]),.doutc(w_n7842_0[2]),.din(n7842));
	jspl jspl_w_n7844_0(.douta(w_n7844_0[0]),.doutb(w_n7844_0[1]),.din(n7844));
	jspl jspl_w_n7849_0(.douta(w_n7849_0[0]),.doutb(w_n7849_0[1]),.din(n7849));
	jspl jspl_w_n7851_0(.douta(w_n7851_0[0]),.doutb(w_n7851_0[1]),.din(n7851));
	jspl jspl_w_n7852_0(.douta(w_n7852_0[0]),.doutb(w_n7852_0[1]),.din(n7852));
	jspl3 jspl3_w_n7853_0(.douta(w_n7853_0[0]),.doutb(w_n7853_0[1]),.doutc(w_n7853_0[2]),.din(n7853));
	jspl jspl_w_n7854_0(.douta(w_n7854_0[0]),.doutb(w_n7854_0[1]),.din(n7854));
	jspl jspl_w_n7858_0(.douta(w_n7858_0[0]),.doutb(w_n7858_0[1]),.din(n7858));
	jspl jspl_w_n7864_0(.douta(w_n7864_0[0]),.doutb(w_n7864_0[1]),.din(n7864));
	jspl jspl_w_n7865_0(.douta(w_n7865_0[0]),.doutb(w_n7865_0[1]),.din(n7865));
	jspl jspl_w_n7867_0(.douta(w_n7867_0[0]),.doutb(w_n7867_0[1]),.din(n7867));
	jspl jspl_w_n7869_0(.douta(w_n7869_0[0]),.doutb(w_n7869_0[1]),.din(n7869));
	jspl jspl_w_n7872_0(.douta(w_n7872_0[0]),.doutb(w_n7872_0[1]),.din(n7872));
	jspl jspl_w_n7878_0(.douta(w_n7878_0[0]),.doutb(w_n7878_0[1]),.din(n7878));
	jspl jspl_w_n7880_0(.douta(w_n7880_0[0]),.doutb(w_n7880_0[1]),.din(n7880));
	jspl3 jspl3_w_n7881_0(.douta(w_n7881_0[0]),.doutb(w_n7881_0[1]),.doutc(w_n7881_0[2]),.din(n7881));
	jspl jspl_w_n7885_0(.douta(w_n7885_0[0]),.doutb(w_n7885_0[1]),.din(n7885));
	jspl jspl_w_n7886_0(.douta(w_n7886_0[0]),.doutb(w_n7886_0[1]),.din(n7886));
	jspl3 jspl3_w_n7887_0(.douta(w_n7887_0[0]),.doutb(w_n7887_0[1]),.doutc(w_n7887_0[2]),.din(n7887));
	jspl jspl_w_n7889_0(.douta(w_n7889_0[0]),.doutb(w_n7889_0[1]),.din(n7889));
	jspl jspl_w_n7894_0(.douta(w_n7894_0[0]),.doutb(w_n7894_0[1]),.din(n7894));
	jspl jspl_w_n7896_0(.douta(w_n7896_0[0]),.doutb(w_n7896_0[1]),.din(n7896));
	jspl jspl_w_n7897_0(.douta(w_n7897_0[0]),.doutb(w_n7897_0[1]),.din(n7897));
	jspl3 jspl3_w_n7898_0(.douta(w_n7898_0[0]),.doutb(w_n7898_0[1]),.doutc(w_n7898_0[2]),.din(n7898));
	jspl jspl_w_n7899_0(.douta(w_n7899_0[0]),.doutb(w_n7899_0[1]),.din(n7899));
	jspl jspl_w_n7903_0(.douta(w_n7903_0[0]),.doutb(w_n7903_0[1]),.din(n7903));
	jspl jspl_w_n7909_0(.douta(w_n7909_0[0]),.doutb(w_n7909_0[1]),.din(n7909));
	jspl jspl_w_n7910_0(.douta(w_n7910_0[0]),.doutb(w_n7910_0[1]),.din(n7910));
	jspl jspl_w_n7912_0(.douta(w_n7912_0[0]),.doutb(w_n7912_0[1]),.din(n7912));
	jspl jspl_w_n7914_0(.douta(w_n7914_0[0]),.doutb(w_n7914_0[1]),.din(n7914));
	jspl jspl_w_n7917_0(.douta(w_n7917_0[0]),.doutb(w_n7917_0[1]),.din(n7917));
	jspl jspl_w_n7923_0(.douta(w_n7923_0[0]),.doutb(w_n7923_0[1]),.din(n7923));
	jspl jspl_w_n7925_0(.douta(w_n7925_0[0]),.doutb(w_n7925_0[1]),.din(n7925));
	jspl3 jspl3_w_n7926_0(.douta(w_n7926_0[0]),.doutb(w_n7926_0[1]),.doutc(w_n7926_0[2]),.din(n7926));
	jspl jspl_w_n7930_0(.douta(w_n7930_0[0]),.doutb(w_n7930_0[1]),.din(n7930));
	jspl jspl_w_n7931_0(.douta(w_n7931_0[0]),.doutb(w_n7931_0[1]),.din(n7931));
	jspl3 jspl3_w_n7932_0(.douta(w_n7932_0[0]),.doutb(w_n7932_0[1]),.doutc(w_n7932_0[2]),.din(n7932));
	jspl jspl_w_n7934_0(.douta(w_n7934_0[0]),.doutb(w_n7934_0[1]),.din(n7934));
	jspl jspl_w_n7939_0(.douta(w_n7939_0[0]),.doutb(w_n7939_0[1]),.din(n7939));
	jspl jspl_w_n7941_0(.douta(w_n7941_0[0]),.doutb(w_n7941_0[1]),.din(n7941));
	jspl jspl_w_n7942_0(.douta(w_n7942_0[0]),.doutb(w_n7942_0[1]),.din(n7942));
	jspl3 jspl3_w_n7943_0(.douta(w_n7943_0[0]),.doutb(w_n7943_0[1]),.doutc(w_n7943_0[2]),.din(n7943));
	jspl jspl_w_n7944_0(.douta(w_n7944_0[0]),.doutb(w_n7944_0[1]),.din(n7944));
	jspl jspl_w_n7948_0(.douta(w_n7948_0[0]),.doutb(w_n7948_0[1]),.din(n7948));
	jspl jspl_w_n7954_0(.douta(w_n7954_0[0]),.doutb(w_n7954_0[1]),.din(n7954));
	jspl jspl_w_n7955_0(.douta(w_n7955_0[0]),.doutb(w_n7955_0[1]),.din(n7955));
	jspl jspl_w_n7957_0(.douta(w_n7957_0[0]),.doutb(w_n7957_0[1]),.din(n7957));
	jspl jspl_w_n7959_0(.douta(w_n7959_0[0]),.doutb(w_n7959_0[1]),.din(n7959));
	jspl jspl_w_n7962_0(.douta(w_n7962_0[0]),.doutb(w_n7962_0[1]),.din(n7962));
	jspl jspl_w_n7968_0(.douta(w_n7968_0[0]),.doutb(w_n7968_0[1]),.din(n7968));
	jspl jspl_w_n7970_0(.douta(w_n7970_0[0]),.doutb(w_n7970_0[1]),.din(n7970));
	jspl3 jspl3_w_n7971_0(.douta(w_n7971_0[0]),.doutb(w_n7971_0[1]),.doutc(w_n7971_0[2]),.din(n7971));
	jspl jspl_w_n7975_0(.douta(w_n7975_0[0]),.doutb(w_n7975_0[1]),.din(n7975));
	jspl jspl_w_n7976_0(.douta(w_n7976_0[0]),.doutb(w_n7976_0[1]),.din(n7976));
	jspl3 jspl3_w_n7977_0(.douta(w_n7977_0[0]),.doutb(w_n7977_0[1]),.doutc(w_n7977_0[2]),.din(n7977));
	jspl jspl_w_n7979_0(.douta(w_n7979_0[0]),.doutb(w_n7979_0[1]),.din(n7979));
	jspl jspl_w_n7984_0(.douta(w_n7984_0[0]),.doutb(w_n7984_0[1]),.din(n7984));
	jspl jspl_w_n7986_0(.douta(w_n7986_0[0]),.doutb(w_n7986_0[1]),.din(n7986));
	jspl jspl_w_n7987_0(.douta(w_n7987_0[0]),.doutb(w_n7987_0[1]),.din(n7987));
	jspl3 jspl3_w_n7988_0(.douta(w_n7988_0[0]),.doutb(w_n7988_0[1]),.doutc(w_n7988_0[2]),.din(n7988));
	jspl jspl_w_n7989_0(.douta(w_n7989_0[0]),.doutb(w_n7989_0[1]),.din(n7989));
	jspl jspl_w_n7993_0(.douta(w_n7993_0[0]),.doutb(w_n7993_0[1]),.din(n7993));
	jspl jspl_w_n7999_0(.douta(w_n7999_0[0]),.doutb(w_n7999_0[1]),.din(n7999));
	jspl jspl_w_n8000_0(.douta(w_n8000_0[0]),.doutb(w_n8000_0[1]),.din(n8000));
	jspl jspl_w_n8002_0(.douta(w_n8002_0[0]),.doutb(w_n8002_0[1]),.din(n8002));
	jspl jspl_w_n8004_0(.douta(w_n8004_0[0]),.doutb(w_n8004_0[1]),.din(n8004));
	jspl jspl_w_n8007_0(.douta(w_n8007_0[0]),.doutb(w_n8007_0[1]),.din(n8007));
	jspl jspl_w_n8013_0(.douta(w_n8013_0[0]),.doutb(w_n8013_0[1]),.din(n8013));
	jspl jspl_w_n8015_0(.douta(w_n8015_0[0]),.doutb(w_n8015_0[1]),.din(n8015));
	jspl3 jspl3_w_n8016_0(.douta(w_n8016_0[0]),.doutb(w_n8016_0[1]),.doutc(w_n8016_0[2]),.din(n8016));
	jspl jspl_w_n8020_0(.douta(w_n8020_0[0]),.doutb(w_n8020_0[1]),.din(n8020));
	jspl jspl_w_n8021_0(.douta(w_n8021_0[0]),.doutb(w_n8021_0[1]),.din(n8021));
	jspl3 jspl3_w_n8022_0(.douta(w_n8022_0[0]),.doutb(w_n8022_0[1]),.doutc(w_n8022_0[2]),.din(n8022));
	jspl jspl_w_n8024_0(.douta(w_n8024_0[0]),.doutb(w_n8024_0[1]),.din(n8024));
	jspl jspl_w_n8029_0(.douta(w_n8029_0[0]),.doutb(w_n8029_0[1]),.din(n8029));
	jspl jspl_w_n8031_0(.douta(w_n8031_0[0]),.doutb(w_n8031_0[1]),.din(n8031));
	jspl jspl_w_n8032_0(.douta(w_n8032_0[0]),.doutb(w_n8032_0[1]),.din(n8032));
	jspl3 jspl3_w_n8033_0(.douta(w_n8033_0[0]),.doutb(w_n8033_0[1]),.doutc(w_n8033_0[2]),.din(n8033));
	jspl3 jspl3_w_n8033_1(.douta(w_n8033_1[0]),.doutb(w_n8033_1[1]),.doutc(w_n8033_1[2]),.din(w_n8033_0[0]));
	jspl jspl_w_n8036_0(.douta(w_n8036_0[0]),.doutb(w_n8036_0[1]),.din(n8036));
	jspl3 jspl3_w_n8037_0(.douta(w_n8037_0[0]),.doutb(w_n8037_0[1]),.doutc(w_n8037_0[2]),.din(n8037));
	jspl jspl_w_n8038_0(.douta(w_n8038_0[0]),.doutb(w_n8038_0[1]),.din(n8038));
	jspl jspl_w_n8039_0(.douta(w_n8039_0[0]),.doutb(w_n8039_0[1]),.din(n8039));
	jspl jspl_w_n8045_0(.douta(w_n8045_0[0]),.doutb(w_n8045_0[1]),.din(n8045));
	jspl3 jspl3_w_n8046_0(.douta(w_n8046_0[0]),.doutb(w_n8046_0[1]),.doutc(w_n8046_0[2]),.din(n8046));
	jspl jspl_w_n8047_0(.douta(w_n8047_0[0]),.doutb(w_n8047_0[1]),.din(n8047));
	jspl jspl_w_n8052_0(.douta(w_n8052_0[0]),.doutb(w_n8052_0[1]),.din(n8052));
	jspl3 jspl3_w_n8053_0(.douta(w_n8053_0[0]),.doutb(w_n8053_0[1]),.doutc(w_n8053_0[2]),.din(n8053));
	jspl3 jspl3_w_n8053_1(.douta(w_n8053_1[0]),.doutb(w_n8053_1[1]),.doutc(w_n8053_1[2]),.din(w_n8053_0[0]));
	jspl3 jspl3_w_n8053_2(.douta(w_n8053_2[0]),.doutb(w_n8053_2[1]),.doutc(w_n8053_2[2]),.din(w_n8053_0[1]));
	jspl3 jspl3_w_n8053_3(.douta(w_n8053_3[0]),.doutb(w_n8053_3[1]),.doutc(w_n8053_3[2]),.din(w_n8053_0[2]));
	jspl3 jspl3_w_n8053_4(.douta(w_n8053_4[0]),.doutb(w_n8053_4[1]),.doutc(w_n8053_4[2]),.din(w_n8053_1[0]));
	jspl3 jspl3_w_n8053_5(.douta(w_n8053_5[0]),.doutb(w_n8053_5[1]),.doutc(w_n8053_5[2]),.din(w_n8053_1[1]));
	jspl3 jspl3_w_n8053_6(.douta(w_n8053_6[0]),.doutb(w_n8053_6[1]),.doutc(w_n8053_6[2]),.din(w_n8053_1[2]));
	jspl3 jspl3_w_n8053_7(.douta(w_n8053_7[0]),.doutb(w_n8053_7[1]),.doutc(w_n8053_7[2]),.din(w_n8053_2[0]));
	jspl3 jspl3_w_n8053_8(.douta(w_n8053_8[0]),.doutb(w_n8053_8[1]),.doutc(w_n8053_8[2]),.din(w_n8053_2[1]));
	jspl3 jspl3_w_n8053_9(.douta(w_n8053_9[0]),.doutb(w_n8053_9[1]),.doutc(w_n8053_9[2]),.din(w_n8053_2[2]));
	jspl3 jspl3_w_n8053_10(.douta(w_n8053_10[0]),.doutb(w_n8053_10[1]),.doutc(w_n8053_10[2]),.din(w_n8053_3[0]));
	jspl3 jspl3_w_n8053_11(.douta(w_n8053_11[0]),.doutb(w_n8053_11[1]),.doutc(w_n8053_11[2]),.din(w_n8053_3[1]));
	jspl3 jspl3_w_n8053_12(.douta(w_n8053_12[0]),.doutb(w_n8053_12[1]),.doutc(w_n8053_12[2]),.din(w_n8053_3[2]));
	jspl3 jspl3_w_n8053_13(.douta(w_n8053_13[0]),.doutb(w_n8053_13[1]),.doutc(w_n8053_13[2]),.din(w_n8053_4[0]));
	jspl3 jspl3_w_n8053_14(.douta(w_n8053_14[0]),.doutb(w_n8053_14[1]),.doutc(w_n8053_14[2]),.din(w_n8053_4[1]));
	jspl3 jspl3_w_n8053_15(.douta(w_n8053_15[0]),.doutb(w_n8053_15[1]),.doutc(w_n8053_15[2]),.din(w_n8053_4[2]));
	jspl3 jspl3_w_n8053_16(.douta(w_n8053_16[0]),.doutb(w_n8053_16[1]),.doutc(w_n8053_16[2]),.din(w_n8053_5[0]));
	jspl3 jspl3_w_n8058_0(.douta(w_n8058_0[0]),.doutb(w_n8058_0[1]),.doutc(w_n8058_0[2]),.din(n8058));
	jspl3 jspl3_w_n8058_1(.douta(w_n8058_1[0]),.doutb(w_n8058_1[1]),.doutc(w_n8058_1[2]),.din(w_n8058_0[0]));
	jspl3 jspl3_w_n8058_2(.douta(w_n8058_2[0]),.doutb(w_n8058_2[1]),.doutc(w_n8058_2[2]),.din(w_n8058_0[1]));
	jspl3 jspl3_w_n8058_3(.douta(w_n8058_3[0]),.doutb(w_n8058_3[1]),.doutc(w_n8058_3[2]),.din(w_n8058_0[2]));
	jspl3 jspl3_w_n8058_4(.douta(w_n8058_4[0]),.doutb(w_n8058_4[1]),.doutc(w_n8058_4[2]),.din(w_n8058_1[0]));
	jspl3 jspl3_w_n8058_5(.douta(w_n8058_5[0]),.doutb(w_n8058_5[1]),.doutc(w_n8058_5[2]),.din(w_n8058_1[1]));
	jspl3 jspl3_w_n8058_6(.douta(w_n8058_6[0]),.doutb(w_n8058_6[1]),.doutc(w_n8058_6[2]),.din(w_n8058_1[2]));
	jspl3 jspl3_w_n8058_7(.douta(w_n8058_7[0]),.doutb(w_n8058_7[1]),.doutc(w_n8058_7[2]),.din(w_n8058_2[0]));
	jspl3 jspl3_w_n8058_8(.douta(w_n8058_8[0]),.doutb(w_n8058_8[1]),.doutc(w_n8058_8[2]),.din(w_n8058_2[1]));
	jspl3 jspl3_w_n8058_9(.douta(w_n8058_9[0]),.doutb(w_n8058_9[1]),.doutc(w_n8058_9[2]),.din(w_n8058_2[2]));
	jspl3 jspl3_w_n8058_10(.douta(w_n8058_10[0]),.doutb(w_n8058_10[1]),.doutc(w_n8058_10[2]),.din(w_n8058_3[0]));
	jspl3 jspl3_w_n8058_11(.douta(w_n8058_11[0]),.doutb(w_n8058_11[1]),.doutc(w_n8058_11[2]),.din(w_n8058_3[1]));
	jspl3 jspl3_w_n8058_12(.douta(w_n8058_12[0]),.doutb(w_n8058_12[1]),.doutc(w_n8058_12[2]),.din(w_n8058_3[2]));
	jspl3 jspl3_w_n8058_13(.douta(w_n8058_13[0]),.doutb(w_n8058_13[1]),.doutc(w_n8058_13[2]),.din(w_n8058_4[0]));
	jspl3 jspl3_w_n8058_14(.douta(w_n8058_14[0]),.doutb(w_n8058_14[1]),.doutc(w_n8058_14[2]),.din(w_n8058_4[1]));
	jspl3 jspl3_w_n8058_15(.douta(w_n8058_15[0]),.doutb(w_n8058_15[1]),.doutc(w_n8058_15[2]),.din(w_n8058_4[2]));
	jspl3 jspl3_w_n8058_16(.douta(w_n8058_16[0]),.doutb(w_n8058_16[1]),.doutc(w_n8058_16[2]),.din(w_n8058_5[0]));
	jspl3 jspl3_w_n8058_17(.douta(w_n8058_17[0]),.doutb(w_n8058_17[1]),.doutc(w_n8058_17[2]),.din(w_n8058_5[1]));
	jspl3 jspl3_w_n8058_18(.douta(w_n8058_18[0]),.doutb(w_n8058_18[1]),.doutc(w_n8058_18[2]),.din(w_n8058_5[2]));
	jspl3 jspl3_w_n8058_19(.douta(w_n8058_19[0]),.doutb(w_n8058_19[1]),.doutc(w_n8058_19[2]),.din(w_n8058_6[0]));
	jspl3 jspl3_w_n8058_20(.douta(w_n8058_20[0]),.doutb(w_n8058_20[1]),.doutc(w_n8058_20[2]),.din(w_n8058_6[1]));
	jspl3 jspl3_w_n8058_21(.douta(w_n8058_21[0]),.doutb(w_n8058_21[1]),.doutc(w_n8058_21[2]),.din(w_n8058_6[2]));
	jspl3 jspl3_w_n8058_22(.douta(w_n8058_22[0]),.doutb(w_n8058_22[1]),.doutc(w_n8058_22[2]),.din(w_n8058_7[0]));
	jspl3 jspl3_w_n8058_23(.douta(w_n8058_23[0]),.doutb(w_n8058_23[1]),.doutc(w_n8058_23[2]),.din(w_n8058_7[1]));
	jspl3 jspl3_w_n8058_24(.douta(w_n8058_24[0]),.doutb(w_n8058_24[1]),.doutc(w_n8058_24[2]),.din(w_n8058_7[2]));
	jspl3 jspl3_w_n8058_25(.douta(w_n8058_25[0]),.doutb(w_n8058_25[1]),.doutc(w_n8058_25[2]),.din(w_n8058_8[0]));
	jspl3 jspl3_w_n8058_26(.douta(w_n8058_26[0]),.doutb(w_n8058_26[1]),.doutc(w_n8058_26[2]),.din(w_n8058_8[1]));
	jspl jspl_w_n8058_27(.douta(w_n8058_27[0]),.doutb(w_n8058_27[1]),.din(w_n8058_8[2]));
	jspl jspl_w_n8061_0(.douta(w_n8061_0[0]),.doutb(w_n8061_0[1]),.din(n8061));
	jspl3 jspl3_w_n8063_0(.douta(w_n8063_0[0]),.doutb(w_n8063_0[1]),.doutc(w_n8063_0[2]),.din(n8063));
	jspl jspl_w_n8063_1(.douta(w_n8063_1[0]),.doutb(w_n8063_1[1]),.din(w_n8063_0[0]));
	jspl3 jspl3_w_n8064_0(.douta(w_n8064_0[0]),.doutb(w_n8064_0[1]),.doutc(w_n8064_0[2]),.din(n8064));
	jspl3 jspl3_w_n8068_0(.douta(w_n8068_0[0]),.doutb(w_n8068_0[1]),.doutc(w_n8068_0[2]),.din(n8068));
	jspl jspl_w_n8069_0(.douta(w_n8069_0[0]),.doutb(w_n8069_0[1]),.din(n8069));
	jspl jspl_w_n8070_0(.douta(w_n8070_0[0]),.doutb(w_n8070_0[1]),.din(n8070));
	jspl jspl_w_n8071_0(.douta(w_n8071_0[0]),.doutb(w_n8071_0[1]),.din(n8071));
	jspl jspl_w_n8073_0(.douta(w_n8073_0[0]),.doutb(w_n8073_0[1]),.din(n8073));
	jspl jspl_w_n8075_0(.douta(w_n8075_0[0]),.doutb(w_n8075_0[1]),.din(n8075));
	jspl jspl_w_n8077_0(.douta(w_n8077_0[0]),.doutb(w_n8077_0[1]),.din(n8077));
	jspl jspl_w_n8080_0(.douta(w_n8080_0[0]),.doutb(w_n8080_0[1]),.din(n8080));
	jspl jspl_w_n8085_0(.douta(w_n8085_0[0]),.doutb(w_n8085_0[1]),.din(n8085));
	jspl3 jspl3_w_n8087_0(.douta(w_n8087_0[0]),.doutb(w_n8087_0[1]),.doutc(w_n8087_0[2]),.din(n8087));
	jspl jspl_w_n8088_0(.douta(w_n8088_0[0]),.doutb(w_n8088_0[1]),.din(n8088));
	jspl jspl_w_n8092_0(.douta(w_n8092_0[0]),.doutb(w_n8092_0[1]),.din(n8092));
	jspl jspl_w_n8093_0(.douta(w_n8093_0[0]),.doutb(w_n8093_0[1]),.din(n8093));
	jspl jspl_w_n8095_0(.douta(w_n8095_0[0]),.doutb(w_n8095_0[1]),.din(n8095));
	jspl jspl_w_n8099_0(.douta(w_n8099_0[0]),.doutb(w_n8099_0[1]),.din(n8099));
	jspl jspl_w_n8101_0(.douta(w_n8101_0[0]),.doutb(w_n8101_0[1]),.din(n8101));
	jspl jspl_w_n8102_0(.douta(w_n8102_0[0]),.doutb(w_n8102_0[1]),.din(n8102));
	jspl3 jspl3_w_n8103_0(.douta(w_n8103_0[0]),.doutb(w_n8103_0[1]),.doutc(w_n8103_0[2]),.din(n8103));
	jspl jspl_w_n8104_0(.douta(w_n8104_0[0]),.doutb(w_n8104_0[1]),.din(n8104));
	jspl jspl_w_n8108_0(.douta(w_n8108_0[0]),.doutb(w_n8108_0[1]),.din(n8108));
	jspl jspl_w_n8110_0(.douta(w_n8110_0[0]),.doutb(w_n8110_0[1]),.din(n8110));
	jspl jspl_w_n8112_0(.douta(w_n8112_0[0]),.doutb(w_n8112_0[1]),.din(n8112));
	jspl jspl_w_n8114_0(.douta(w_n8114_0[0]),.doutb(w_n8114_0[1]),.din(n8114));
	jspl jspl_w_n8117_0(.douta(w_n8117_0[0]),.doutb(w_n8117_0[1]),.din(n8117));
	jspl jspl_w_n8123_0(.douta(w_n8123_0[0]),.doutb(w_n8123_0[1]),.din(n8123));
	jspl3 jspl3_w_n8125_0(.douta(w_n8125_0[0]),.doutb(w_n8125_0[1]),.doutc(w_n8125_0[2]),.din(n8125));
	jspl jspl_w_n8126_0(.douta(w_n8126_0[0]),.doutb(w_n8126_0[1]),.din(n8126));
	jspl jspl_w_n8131_0(.douta(w_n8131_0[0]),.doutb(w_n8131_0[1]),.din(n8131));
	jspl jspl_w_n8133_0(.douta(w_n8133_0[0]),.doutb(w_n8133_0[1]),.din(n8133));
	jspl jspl_w_n8135_0(.douta(w_n8135_0[0]),.doutb(w_n8135_0[1]),.din(n8135));
	jspl jspl_w_n8139_0(.douta(w_n8139_0[0]),.doutb(w_n8139_0[1]),.din(n8139));
	jspl jspl_w_n8141_0(.douta(w_n8141_0[0]),.doutb(w_n8141_0[1]),.din(n8141));
	jspl jspl_w_n8142_0(.douta(w_n8142_0[0]),.doutb(w_n8142_0[1]),.din(n8142));
	jspl3 jspl3_w_n8143_0(.douta(w_n8143_0[0]),.doutb(w_n8143_0[1]),.doutc(w_n8143_0[2]),.din(n8143));
	jspl jspl_w_n8144_0(.douta(w_n8144_0[0]),.doutb(w_n8144_0[1]),.din(n8144));
	jspl jspl_w_n8150_0(.douta(w_n8150_0[0]),.doutb(w_n8150_0[1]),.din(n8150));
	jspl jspl_w_n8151_0(.douta(w_n8151_0[0]),.doutb(w_n8151_0[1]),.din(n8151));
	jspl jspl_w_n8153_0(.douta(w_n8153_0[0]),.doutb(w_n8153_0[1]),.din(n8153));
	jspl jspl_w_n8155_0(.douta(w_n8155_0[0]),.doutb(w_n8155_0[1]),.din(n8155));
	jspl jspl_w_n8157_0(.douta(w_n8157_0[0]),.doutb(w_n8157_0[1]),.din(n8157));
	jspl jspl_w_n8163_0(.douta(w_n8163_0[0]),.doutb(w_n8163_0[1]),.din(n8163));
	jspl jspl_w_n8165_0(.douta(w_n8165_0[0]),.doutb(w_n8165_0[1]),.din(n8165));
	jspl3 jspl3_w_n8166_0(.douta(w_n8166_0[0]),.doutb(w_n8166_0[1]),.doutc(w_n8166_0[2]),.din(n8166));
	jspl jspl_w_n8169_0(.douta(w_n8169_0[0]),.doutb(w_n8169_0[1]),.din(n8169));
	jspl jspl_w_n8170_0(.douta(w_n8170_0[0]),.doutb(w_n8170_0[1]),.din(n8170));
	jspl3 jspl3_w_n8171_0(.douta(w_n8171_0[0]),.doutb(w_n8171_0[1]),.doutc(w_n8171_0[2]),.din(n8171));
	jspl jspl_w_n8173_0(.douta(w_n8173_0[0]),.doutb(w_n8173_0[1]),.din(n8173));
	jspl jspl_w_n8175_0(.douta(w_n8175_0[0]),.doutb(w_n8175_0[1]),.din(n8175));
	jspl jspl_w_n8177_0(.douta(w_n8177_0[0]),.doutb(w_n8177_0[1]),.din(n8177));
	jspl jspl_w_n8183_0(.douta(w_n8183_0[0]),.doutb(w_n8183_0[1]),.din(n8183));
	jspl3 jspl3_w_n8185_0(.douta(w_n8185_0[0]),.doutb(w_n8185_0[1]),.doutc(w_n8185_0[2]),.din(n8185));
	jspl jspl_w_n8186_0(.douta(w_n8186_0[0]),.doutb(w_n8186_0[1]),.din(n8186));
	jspl jspl_w_n8188_0(.douta(w_n8188_0[0]),.doutb(w_n8188_0[1]),.din(n8188));
	jspl jspl_w_n8190_0(.douta(w_n8190_0[0]),.doutb(w_n8190_0[1]),.din(n8190));
	jspl jspl_w_n8194_0(.douta(w_n8194_0[0]),.doutb(w_n8194_0[1]),.din(n8194));
	jspl jspl_w_n8196_0(.douta(w_n8196_0[0]),.doutb(w_n8196_0[1]),.din(n8196));
	jspl jspl_w_n8197_0(.douta(w_n8197_0[0]),.doutb(w_n8197_0[1]),.din(n8197));
	jspl jspl_w_n8198_0(.douta(w_n8198_0[0]),.doutb(w_n8198_0[1]),.din(n8198));
	jspl3 jspl3_w_n8199_0(.douta(w_n8199_0[0]),.doutb(w_n8199_0[1]),.doutc(w_n8199_0[2]),.din(n8199));
	jspl jspl_w_n8202_0(.douta(w_n8202_0[0]),.doutb(w_n8202_0[1]),.din(n8202));
	jspl jspl_w_n8203_0(.douta(w_n8203_0[0]),.doutb(w_n8203_0[1]),.din(n8203));
	jspl3 jspl3_w_n8204_0(.douta(w_n8204_0[0]),.doutb(w_n8204_0[1]),.doutc(w_n8204_0[2]),.din(n8204));
	jspl jspl_w_n8206_0(.douta(w_n8206_0[0]),.doutb(w_n8206_0[1]),.din(n8206));
	jspl jspl_w_n8210_0(.douta(w_n8210_0[0]),.doutb(w_n8210_0[1]),.din(n8210));
	jspl jspl_w_n8212_0(.douta(w_n8212_0[0]),.doutb(w_n8212_0[1]),.din(n8212));
	jspl jspl_w_n8213_0(.douta(w_n8213_0[0]),.doutb(w_n8213_0[1]),.din(n8213));
	jspl3 jspl3_w_n8214_0(.douta(w_n8214_0[0]),.doutb(w_n8214_0[1]),.doutc(w_n8214_0[2]),.din(n8214));
	jspl jspl_w_n8215_0(.douta(w_n8215_0[0]),.doutb(w_n8215_0[1]),.din(n8215));
	jspl jspl_w_n8218_0(.douta(w_n8218_0[0]),.doutb(w_n8218_0[1]),.din(n8218));
	jspl jspl_w_n8224_0(.douta(w_n8224_0[0]),.doutb(w_n8224_0[1]),.din(n8224));
	jspl jspl_w_n8225_0(.douta(w_n8225_0[0]),.doutb(w_n8225_0[1]),.din(n8225));
	jspl jspl_w_n8227_0(.douta(w_n8227_0[0]),.doutb(w_n8227_0[1]),.din(n8227));
	jspl jspl_w_n8229_0(.douta(w_n8229_0[0]),.doutb(w_n8229_0[1]),.din(n8229));
	jspl jspl_w_n8231_0(.douta(w_n8231_0[0]),.doutb(w_n8231_0[1]),.din(n8231));
	jspl jspl_w_n8237_0(.douta(w_n8237_0[0]),.doutb(w_n8237_0[1]),.din(n8237));
	jspl jspl_w_n8239_0(.douta(w_n8239_0[0]),.doutb(w_n8239_0[1]),.din(n8239));
	jspl3 jspl3_w_n8240_0(.douta(w_n8240_0[0]),.doutb(w_n8240_0[1]),.doutc(w_n8240_0[2]),.din(n8240));
	jspl jspl_w_n8243_0(.douta(w_n8243_0[0]),.doutb(w_n8243_0[1]),.din(n8243));
	jspl jspl_w_n8244_0(.douta(w_n8244_0[0]),.doutb(w_n8244_0[1]),.din(n8244));
	jspl3 jspl3_w_n8245_0(.douta(w_n8245_0[0]),.doutb(w_n8245_0[1]),.doutc(w_n8245_0[2]),.din(n8245));
	jspl jspl_w_n8247_0(.douta(w_n8247_0[0]),.doutb(w_n8247_0[1]),.din(n8247));
	jspl jspl_w_n8251_0(.douta(w_n8251_0[0]),.doutb(w_n8251_0[1]),.din(n8251));
	jspl jspl_w_n8253_0(.douta(w_n8253_0[0]),.doutb(w_n8253_0[1]),.din(n8253));
	jspl jspl_w_n8254_0(.douta(w_n8254_0[0]),.doutb(w_n8254_0[1]),.din(n8254));
	jspl3 jspl3_w_n8255_0(.douta(w_n8255_0[0]),.doutb(w_n8255_0[1]),.doutc(w_n8255_0[2]),.din(n8255));
	jspl jspl_w_n8256_0(.douta(w_n8256_0[0]),.doutb(w_n8256_0[1]),.din(n8256));
	jspl jspl_w_n8259_0(.douta(w_n8259_0[0]),.doutb(w_n8259_0[1]),.din(n8259));
	jspl jspl_w_n8265_0(.douta(w_n8265_0[0]),.doutb(w_n8265_0[1]),.din(n8265));
	jspl jspl_w_n8266_0(.douta(w_n8266_0[0]),.doutb(w_n8266_0[1]),.din(n8266));
	jspl jspl_w_n8268_0(.douta(w_n8268_0[0]),.doutb(w_n8268_0[1]),.din(n8268));
	jspl jspl_w_n8270_0(.douta(w_n8270_0[0]),.doutb(w_n8270_0[1]),.din(n8270));
	jspl jspl_w_n8272_0(.douta(w_n8272_0[0]),.doutb(w_n8272_0[1]),.din(n8272));
	jspl jspl_w_n8278_0(.douta(w_n8278_0[0]),.doutb(w_n8278_0[1]),.din(n8278));
	jspl jspl_w_n8280_0(.douta(w_n8280_0[0]),.doutb(w_n8280_0[1]),.din(n8280));
	jspl3 jspl3_w_n8281_0(.douta(w_n8281_0[0]),.doutb(w_n8281_0[1]),.doutc(w_n8281_0[2]),.din(n8281));
	jspl jspl_w_n8284_0(.douta(w_n8284_0[0]),.doutb(w_n8284_0[1]),.din(n8284));
	jspl jspl_w_n8285_0(.douta(w_n8285_0[0]),.doutb(w_n8285_0[1]),.din(n8285));
	jspl3 jspl3_w_n8286_0(.douta(w_n8286_0[0]),.doutb(w_n8286_0[1]),.doutc(w_n8286_0[2]),.din(n8286));
	jspl jspl_w_n8288_0(.douta(w_n8288_0[0]),.doutb(w_n8288_0[1]),.din(n8288));
	jspl jspl_w_n8292_0(.douta(w_n8292_0[0]),.doutb(w_n8292_0[1]),.din(n8292));
	jspl jspl_w_n8294_0(.douta(w_n8294_0[0]),.doutb(w_n8294_0[1]),.din(n8294));
	jspl jspl_w_n8295_0(.douta(w_n8295_0[0]),.doutb(w_n8295_0[1]),.din(n8295));
	jspl3 jspl3_w_n8296_0(.douta(w_n8296_0[0]),.doutb(w_n8296_0[1]),.doutc(w_n8296_0[2]),.din(n8296));
	jspl jspl_w_n8297_0(.douta(w_n8297_0[0]),.doutb(w_n8297_0[1]),.din(n8297));
	jspl jspl_w_n8300_0(.douta(w_n8300_0[0]),.doutb(w_n8300_0[1]),.din(n8300));
	jspl jspl_w_n8306_0(.douta(w_n8306_0[0]),.doutb(w_n8306_0[1]),.din(n8306));
	jspl jspl_w_n8307_0(.douta(w_n8307_0[0]),.doutb(w_n8307_0[1]),.din(n8307));
	jspl jspl_w_n8309_0(.douta(w_n8309_0[0]),.doutb(w_n8309_0[1]),.din(n8309));
	jspl jspl_w_n8311_0(.douta(w_n8311_0[0]),.doutb(w_n8311_0[1]),.din(n8311));
	jspl jspl_w_n8313_0(.douta(w_n8313_0[0]),.doutb(w_n8313_0[1]),.din(n8313));
	jspl jspl_w_n8319_0(.douta(w_n8319_0[0]),.doutb(w_n8319_0[1]),.din(n8319));
	jspl jspl_w_n8321_0(.douta(w_n8321_0[0]),.doutb(w_n8321_0[1]),.din(n8321));
	jspl3 jspl3_w_n8322_0(.douta(w_n8322_0[0]),.doutb(w_n8322_0[1]),.doutc(w_n8322_0[2]),.din(n8322));
	jspl jspl_w_n8325_0(.douta(w_n8325_0[0]),.doutb(w_n8325_0[1]),.din(n8325));
	jspl jspl_w_n8326_0(.douta(w_n8326_0[0]),.doutb(w_n8326_0[1]),.din(n8326));
	jspl3 jspl3_w_n8327_0(.douta(w_n8327_0[0]),.doutb(w_n8327_0[1]),.doutc(w_n8327_0[2]),.din(n8327));
	jspl jspl_w_n8329_0(.douta(w_n8329_0[0]),.doutb(w_n8329_0[1]),.din(n8329));
	jspl jspl_w_n8333_0(.douta(w_n8333_0[0]),.doutb(w_n8333_0[1]),.din(n8333));
	jspl jspl_w_n8335_0(.douta(w_n8335_0[0]),.doutb(w_n8335_0[1]),.din(n8335));
	jspl jspl_w_n8336_0(.douta(w_n8336_0[0]),.doutb(w_n8336_0[1]),.din(n8336));
	jspl3 jspl3_w_n8337_0(.douta(w_n8337_0[0]),.doutb(w_n8337_0[1]),.doutc(w_n8337_0[2]),.din(n8337));
	jspl jspl_w_n8338_0(.douta(w_n8338_0[0]),.doutb(w_n8338_0[1]),.din(n8338));
	jspl jspl_w_n8341_0(.douta(w_n8341_0[0]),.doutb(w_n8341_0[1]),.din(n8341));
	jspl jspl_w_n8347_0(.douta(w_n8347_0[0]),.doutb(w_n8347_0[1]),.din(n8347));
	jspl jspl_w_n8348_0(.douta(w_n8348_0[0]),.doutb(w_n8348_0[1]),.din(n8348));
	jspl jspl_w_n8350_0(.douta(w_n8350_0[0]),.doutb(w_n8350_0[1]),.din(n8350));
	jspl jspl_w_n8352_0(.douta(w_n8352_0[0]),.doutb(w_n8352_0[1]),.din(n8352));
	jspl jspl_w_n8354_0(.douta(w_n8354_0[0]),.doutb(w_n8354_0[1]),.din(n8354));
	jspl jspl_w_n8360_0(.douta(w_n8360_0[0]),.doutb(w_n8360_0[1]),.din(n8360));
	jspl jspl_w_n8362_0(.douta(w_n8362_0[0]),.doutb(w_n8362_0[1]),.din(n8362));
	jspl3 jspl3_w_n8363_0(.douta(w_n8363_0[0]),.doutb(w_n8363_0[1]),.doutc(w_n8363_0[2]),.din(n8363));
	jspl jspl_w_n8366_0(.douta(w_n8366_0[0]),.doutb(w_n8366_0[1]),.din(n8366));
	jspl jspl_w_n8367_0(.douta(w_n8367_0[0]),.doutb(w_n8367_0[1]),.din(n8367));
	jspl3 jspl3_w_n8368_0(.douta(w_n8368_0[0]),.doutb(w_n8368_0[1]),.doutc(w_n8368_0[2]),.din(n8368));
	jspl jspl_w_n8370_0(.douta(w_n8370_0[0]),.doutb(w_n8370_0[1]),.din(n8370));
	jspl jspl_w_n8374_0(.douta(w_n8374_0[0]),.doutb(w_n8374_0[1]),.din(n8374));
	jspl jspl_w_n8376_0(.douta(w_n8376_0[0]),.doutb(w_n8376_0[1]),.din(n8376));
	jspl jspl_w_n8377_0(.douta(w_n8377_0[0]),.doutb(w_n8377_0[1]),.din(n8377));
	jspl3 jspl3_w_n8378_0(.douta(w_n8378_0[0]),.doutb(w_n8378_0[1]),.doutc(w_n8378_0[2]),.din(n8378));
	jspl jspl_w_n8379_0(.douta(w_n8379_0[0]),.doutb(w_n8379_0[1]),.din(n8379));
	jspl jspl_w_n8382_0(.douta(w_n8382_0[0]),.doutb(w_n8382_0[1]),.din(n8382));
	jspl jspl_w_n8388_0(.douta(w_n8388_0[0]),.doutb(w_n8388_0[1]),.din(n8388));
	jspl jspl_w_n8389_0(.douta(w_n8389_0[0]),.doutb(w_n8389_0[1]),.din(n8389));
	jspl jspl_w_n8391_0(.douta(w_n8391_0[0]),.doutb(w_n8391_0[1]),.din(n8391));
	jspl jspl_w_n8393_0(.douta(w_n8393_0[0]),.doutb(w_n8393_0[1]),.din(n8393));
	jspl jspl_w_n8395_0(.douta(w_n8395_0[0]),.doutb(w_n8395_0[1]),.din(n8395));
	jspl jspl_w_n8401_0(.douta(w_n8401_0[0]),.doutb(w_n8401_0[1]),.din(n8401));
	jspl jspl_w_n8403_0(.douta(w_n8403_0[0]),.doutb(w_n8403_0[1]),.din(n8403));
	jspl3 jspl3_w_n8404_0(.douta(w_n8404_0[0]),.doutb(w_n8404_0[1]),.doutc(w_n8404_0[2]),.din(n8404));
	jspl jspl_w_n8407_0(.douta(w_n8407_0[0]),.doutb(w_n8407_0[1]),.din(n8407));
	jspl jspl_w_n8408_0(.douta(w_n8408_0[0]),.doutb(w_n8408_0[1]),.din(n8408));
	jspl3 jspl3_w_n8409_0(.douta(w_n8409_0[0]),.doutb(w_n8409_0[1]),.doutc(w_n8409_0[2]),.din(n8409));
	jspl jspl_w_n8411_0(.douta(w_n8411_0[0]),.doutb(w_n8411_0[1]),.din(n8411));
	jspl jspl_w_n8415_0(.douta(w_n8415_0[0]),.doutb(w_n8415_0[1]),.din(n8415));
	jspl jspl_w_n8417_0(.douta(w_n8417_0[0]),.doutb(w_n8417_0[1]),.din(n8417));
	jspl jspl_w_n8418_0(.douta(w_n8418_0[0]),.doutb(w_n8418_0[1]),.din(n8418));
	jspl3 jspl3_w_n8419_0(.douta(w_n8419_0[0]),.doutb(w_n8419_0[1]),.doutc(w_n8419_0[2]),.din(n8419));
	jspl jspl_w_n8423_0(.douta(w_n8423_0[0]),.doutb(w_n8423_0[1]),.din(n8423));
	jspl jspl_w_n8429_0(.douta(w_n8429_0[0]),.doutb(w_n8429_0[1]),.din(n8429));
	jspl3 jspl3_w_n8431_0(.douta(w_n8431_0[0]),.doutb(w_n8431_0[1]),.doutc(w_n8431_0[2]),.din(n8431));
	jspl jspl_w_n8433_0(.douta(w_n8433_0[0]),.doutb(w_n8433_0[1]),.din(n8433));
	jspl3 jspl3_w_n8438_0(.douta(w_n8438_0[0]),.doutb(w_n8438_0[1]),.doutc(w_n8438_0[2]),.din(n8438));
	jspl jspl_w_n8439_0(.douta(w_n8439_0[0]),.doutb(w_n8439_0[1]),.din(n8439));
	jspl jspl_w_n8440_0(.douta(w_n8440_0[0]),.doutb(w_n8440_0[1]),.din(n8440));
	jspl jspl_w_n8445_0(.douta(w_n8445_0[0]),.doutb(w_n8445_0[1]),.din(n8445));
	jspl3 jspl3_w_n8446_0(.douta(w_n8446_0[0]),.doutb(w_n8446_0[1]),.doutc(w_n8446_0[2]),.din(n8446));
	jspl jspl_w_n8451_0(.douta(w_n8451_0[0]),.doutb(w_n8451_0[1]),.din(n8451));
	jspl jspl_w_n8458_0(.douta(w_n8458_0[0]),.doutb(w_n8458_0[1]),.din(n8458));
	jspl3 jspl3_w_n8460_0(.douta(w_n8460_0[0]),.doutb(w_n8460_0[1]),.doutc(w_n8460_0[2]),.din(n8460));
	jspl jspl_w_n8460_1(.douta(w_n8460_1[0]),.doutb(w_n8460_1[1]),.din(w_n8460_0[0]));
	jspl jspl_w_n8461_0(.douta(w_n8461_0[0]),.doutb(w_n8461_0[1]),.din(n8461));
	jspl3 jspl3_w_n8464_0(.douta(w_n8464_0[0]),.doutb(w_n8464_0[1]),.doutc(w_n8464_0[2]),.din(n8464));
	jspl jspl_w_n8465_0(.douta(w_n8465_0[0]),.doutb(w_n8465_0[1]),.din(n8465));
	jspl jspl_w_n8466_0(.douta(w_n8466_0[0]),.doutb(w_n8466_0[1]),.din(n8466));
	jspl jspl_w_n8467_0(.douta(w_n8467_0[0]),.doutb(w_n8467_0[1]),.din(n8467));
	jspl jspl_w_n8469_0(.douta(w_n8469_0[0]),.doutb(w_n8469_0[1]),.din(n8469));
	jspl jspl_w_n8471_0(.douta(w_n8471_0[0]),.doutb(w_n8471_0[1]),.din(n8471));
	jspl jspl_w_n8473_0(.douta(w_n8473_0[0]),.doutb(w_n8473_0[1]),.din(n8473));
	jspl jspl_w_n8482_0(.douta(w_n8482_0[0]),.doutb(w_n8482_0[1]),.din(n8482));
	jspl3 jspl3_w_n8484_0(.douta(w_n8484_0[0]),.doutb(w_n8484_0[1]),.doutc(w_n8484_0[2]),.din(n8484));
	jspl jspl_w_n8485_0(.douta(w_n8485_0[0]),.doutb(w_n8485_0[1]),.din(n8485));
	jspl jspl_w_n8489_0(.douta(w_n8489_0[0]),.doutb(w_n8489_0[1]),.din(n8489));
	jspl jspl_w_n8491_0(.douta(w_n8491_0[0]),.doutb(w_n8491_0[1]),.din(n8491));
	jspl jspl_w_n8493_0(.douta(w_n8493_0[0]),.doutb(w_n8493_0[1]),.din(n8493));
	jspl jspl_w_n8498_0(.douta(w_n8498_0[0]),.doutb(w_n8498_0[1]),.din(n8498));
	jspl jspl_w_n8500_0(.douta(w_n8500_0[0]),.doutb(w_n8500_0[1]),.din(n8500));
	jspl jspl_w_n8501_0(.douta(w_n8501_0[0]),.doutb(w_n8501_0[1]),.din(n8501));
	jspl3 jspl3_w_n8502_0(.douta(w_n8502_0[0]),.doutb(w_n8502_0[1]),.doutc(w_n8502_0[2]),.din(n8502));
	jspl jspl_w_n8503_0(.douta(w_n8503_0[0]),.doutb(w_n8503_0[1]),.din(n8503));
	jspl jspl_w_n8508_0(.douta(w_n8508_0[0]),.doutb(w_n8508_0[1]),.din(n8508));
	jspl jspl_w_n8509_0(.douta(w_n8509_0[0]),.doutb(w_n8509_0[1]),.din(n8509));
	jspl jspl_w_n8511_0(.douta(w_n8511_0[0]),.doutb(w_n8511_0[1]),.din(n8511));
	jspl jspl_w_n8513_0(.douta(w_n8513_0[0]),.doutb(w_n8513_0[1]),.din(n8513));
	jspl jspl_w_n8516_0(.douta(w_n8516_0[0]),.doutb(w_n8516_0[1]),.din(n8516));
	jspl jspl_w_n8522_0(.douta(w_n8522_0[0]),.doutb(w_n8522_0[1]),.din(n8522));
	jspl3 jspl3_w_n8524_0(.douta(w_n8524_0[0]),.doutb(w_n8524_0[1]),.doutc(w_n8524_0[2]),.din(n8524));
	jspl jspl_w_n8525_0(.douta(w_n8525_0[0]),.doutb(w_n8525_0[1]),.din(n8525));
	jspl jspl_w_n8529_0(.douta(w_n8529_0[0]),.doutb(w_n8529_0[1]),.din(n8529));
	jspl jspl_w_n8530_0(.douta(w_n8530_0[0]),.doutb(w_n8530_0[1]),.din(n8530));
	jspl jspl_w_n8532_0(.douta(w_n8532_0[0]),.doutb(w_n8532_0[1]),.din(n8532));
	jspl jspl_w_n8537_0(.douta(w_n8537_0[0]),.doutb(w_n8537_0[1]),.din(n8537));
	jspl jspl_w_n8539_0(.douta(w_n8539_0[0]),.doutb(w_n8539_0[1]),.din(n8539));
	jspl jspl_w_n8540_0(.douta(w_n8540_0[0]),.doutb(w_n8540_0[1]),.din(n8540));
	jspl3 jspl3_w_n8541_0(.douta(w_n8541_0[0]),.doutb(w_n8541_0[1]),.doutc(w_n8541_0[2]),.din(n8541));
	jspl jspl_w_n8542_0(.douta(w_n8542_0[0]),.doutb(w_n8542_0[1]),.din(n8542));
	jspl jspl_w_n8546_0(.douta(w_n8546_0[0]),.doutb(w_n8546_0[1]),.din(n8546));
	jspl jspl_w_n8547_0(.douta(w_n8547_0[0]),.doutb(w_n8547_0[1]),.din(n8547));
	jspl jspl_w_n8549_0(.douta(w_n8549_0[0]),.doutb(w_n8549_0[1]),.din(n8549));
	jspl jspl_w_n8551_0(.douta(w_n8551_0[0]),.doutb(w_n8551_0[1]),.din(n8551));
	jspl jspl_w_n8554_0(.douta(w_n8554_0[0]),.doutb(w_n8554_0[1]),.din(n8554));
	jspl jspl_w_n8560_0(.douta(w_n8560_0[0]),.doutb(w_n8560_0[1]),.din(n8560));
	jspl jspl_w_n8562_0(.douta(w_n8562_0[0]),.doutb(w_n8562_0[1]),.din(n8562));
	jspl3 jspl3_w_n8563_0(.douta(w_n8563_0[0]),.doutb(w_n8563_0[1]),.doutc(w_n8563_0[2]),.din(n8563));
	jspl jspl_w_n8567_0(.douta(w_n8567_0[0]),.doutb(w_n8567_0[1]),.din(n8567));
	jspl jspl_w_n8568_0(.douta(w_n8568_0[0]),.doutb(w_n8568_0[1]),.din(n8568));
	jspl3 jspl3_w_n8569_0(.douta(w_n8569_0[0]),.doutb(w_n8569_0[1]),.doutc(w_n8569_0[2]),.din(n8569));
	jspl jspl_w_n8571_0(.douta(w_n8571_0[0]),.doutb(w_n8571_0[1]),.din(n8571));
	jspl jspl_w_n8576_0(.douta(w_n8576_0[0]),.doutb(w_n8576_0[1]),.din(n8576));
	jspl jspl_w_n8578_0(.douta(w_n8578_0[0]),.doutb(w_n8578_0[1]),.din(n8578));
	jspl jspl_w_n8579_0(.douta(w_n8579_0[0]),.doutb(w_n8579_0[1]),.din(n8579));
	jspl3 jspl3_w_n8580_0(.douta(w_n8580_0[0]),.doutb(w_n8580_0[1]),.doutc(w_n8580_0[2]),.din(n8580));
	jspl jspl_w_n8581_0(.douta(w_n8581_0[0]),.doutb(w_n8581_0[1]),.din(n8581));
	jspl jspl_w_n8585_0(.douta(w_n8585_0[0]),.doutb(w_n8585_0[1]),.din(n8585));
	jspl jspl_w_n8591_0(.douta(w_n8591_0[0]),.doutb(w_n8591_0[1]),.din(n8591));
	jspl jspl_w_n8592_0(.douta(w_n8592_0[0]),.doutb(w_n8592_0[1]),.din(n8592));
	jspl jspl_w_n8594_0(.douta(w_n8594_0[0]),.doutb(w_n8594_0[1]),.din(n8594));
	jspl jspl_w_n8599_0(.douta(w_n8599_0[0]),.doutb(w_n8599_0[1]),.din(n8599));
	jspl jspl_w_n8601_0(.douta(w_n8601_0[0]),.doutb(w_n8601_0[1]),.din(n8601));
	jspl jspl_w_n8602_0(.douta(w_n8602_0[0]),.doutb(w_n8602_0[1]),.din(n8602));
	jspl3 jspl3_w_n8603_0(.douta(w_n8603_0[0]),.doutb(w_n8603_0[1]),.doutc(w_n8603_0[2]),.din(n8603));
	jspl jspl_w_n8604_0(.douta(w_n8604_0[0]),.doutb(w_n8604_0[1]),.din(n8604));
	jspl jspl_w_n8607_0(.douta(w_n8607_0[0]),.doutb(w_n8607_0[1]),.din(n8607));
	jspl jspl_w_n8609_0(.douta(w_n8609_0[0]),.doutb(w_n8609_0[1]),.din(n8609));
	jspl jspl_w_n8611_0(.douta(w_n8611_0[0]),.doutb(w_n8611_0[1]),.din(n8611));
	jspl jspl_w_n8614_0(.douta(w_n8614_0[0]),.doutb(w_n8614_0[1]),.din(n8614));
	jspl jspl_w_n8620_0(.douta(w_n8620_0[0]),.doutb(w_n8620_0[1]),.din(n8620));
	jspl3 jspl3_w_n8622_0(.douta(w_n8622_0[0]),.doutb(w_n8622_0[1]),.doutc(w_n8622_0[2]),.din(n8622));
	jspl jspl_w_n8623_0(.douta(w_n8623_0[0]),.doutb(w_n8623_0[1]),.din(n8623));
	jspl jspl_w_n8627_0(.douta(w_n8627_0[0]),.doutb(w_n8627_0[1]),.din(n8627));
	jspl jspl_w_n8633_0(.douta(w_n8633_0[0]),.doutb(w_n8633_0[1]),.din(n8633));
	jspl jspl_w_n8634_0(.douta(w_n8634_0[0]),.doutb(w_n8634_0[1]),.din(n8634));
	jspl jspl_w_n8636_0(.douta(w_n8636_0[0]),.doutb(w_n8636_0[1]),.din(n8636));
	jspl jspl_w_n8638_0(.douta(w_n8638_0[0]),.doutb(w_n8638_0[1]),.din(n8638));
	jspl jspl_w_n8641_0(.douta(w_n8641_0[0]),.doutb(w_n8641_0[1]),.din(n8641));
	jspl jspl_w_n8647_0(.douta(w_n8647_0[0]),.doutb(w_n8647_0[1]),.din(n8647));
	jspl jspl_w_n8649_0(.douta(w_n8649_0[0]),.doutb(w_n8649_0[1]),.din(n8649));
	jspl3 jspl3_w_n8650_0(.douta(w_n8650_0[0]),.doutb(w_n8650_0[1]),.doutc(w_n8650_0[2]),.din(n8650));
	jspl jspl_w_n8654_0(.douta(w_n8654_0[0]),.doutb(w_n8654_0[1]),.din(n8654));
	jspl jspl_w_n8655_0(.douta(w_n8655_0[0]),.doutb(w_n8655_0[1]),.din(n8655));
	jspl3 jspl3_w_n8656_0(.douta(w_n8656_0[0]),.doutb(w_n8656_0[1]),.doutc(w_n8656_0[2]),.din(n8656));
	jspl jspl_w_n8658_0(.douta(w_n8658_0[0]),.doutb(w_n8658_0[1]),.din(n8658));
	jspl jspl_w_n8663_0(.douta(w_n8663_0[0]),.doutb(w_n8663_0[1]),.din(n8663));
	jspl jspl_w_n8665_0(.douta(w_n8665_0[0]),.doutb(w_n8665_0[1]),.din(n8665));
	jspl jspl_w_n8666_0(.douta(w_n8666_0[0]),.doutb(w_n8666_0[1]),.din(n8666));
	jspl3 jspl3_w_n8667_0(.douta(w_n8667_0[0]),.doutb(w_n8667_0[1]),.doutc(w_n8667_0[2]),.din(n8667));
	jspl jspl_w_n8668_0(.douta(w_n8668_0[0]),.doutb(w_n8668_0[1]),.din(n8668));
	jspl jspl_w_n8672_0(.douta(w_n8672_0[0]),.doutb(w_n8672_0[1]),.din(n8672));
	jspl jspl_w_n8678_0(.douta(w_n8678_0[0]),.doutb(w_n8678_0[1]),.din(n8678));
	jspl jspl_w_n8679_0(.douta(w_n8679_0[0]),.doutb(w_n8679_0[1]),.din(n8679));
	jspl jspl_w_n8681_0(.douta(w_n8681_0[0]),.doutb(w_n8681_0[1]),.din(n8681));
	jspl jspl_w_n8683_0(.douta(w_n8683_0[0]),.doutb(w_n8683_0[1]),.din(n8683));
	jspl jspl_w_n8686_0(.douta(w_n8686_0[0]),.doutb(w_n8686_0[1]),.din(n8686));
	jspl jspl_w_n8692_0(.douta(w_n8692_0[0]),.doutb(w_n8692_0[1]),.din(n8692));
	jspl jspl_w_n8694_0(.douta(w_n8694_0[0]),.doutb(w_n8694_0[1]),.din(n8694));
	jspl3 jspl3_w_n8695_0(.douta(w_n8695_0[0]),.doutb(w_n8695_0[1]),.doutc(w_n8695_0[2]),.din(n8695));
	jspl jspl_w_n8699_0(.douta(w_n8699_0[0]),.doutb(w_n8699_0[1]),.din(n8699));
	jspl jspl_w_n8700_0(.douta(w_n8700_0[0]),.doutb(w_n8700_0[1]),.din(n8700));
	jspl3 jspl3_w_n8701_0(.douta(w_n8701_0[0]),.doutb(w_n8701_0[1]),.doutc(w_n8701_0[2]),.din(n8701));
	jspl jspl_w_n8703_0(.douta(w_n8703_0[0]),.doutb(w_n8703_0[1]),.din(n8703));
	jspl jspl_w_n8708_0(.douta(w_n8708_0[0]),.doutb(w_n8708_0[1]),.din(n8708));
	jspl jspl_w_n8710_0(.douta(w_n8710_0[0]),.doutb(w_n8710_0[1]),.din(n8710));
	jspl jspl_w_n8711_0(.douta(w_n8711_0[0]),.doutb(w_n8711_0[1]),.din(n8711));
	jspl3 jspl3_w_n8712_0(.douta(w_n8712_0[0]),.doutb(w_n8712_0[1]),.doutc(w_n8712_0[2]),.din(n8712));
	jspl jspl_w_n8713_0(.douta(w_n8713_0[0]),.doutb(w_n8713_0[1]),.din(n8713));
	jspl jspl_w_n8717_0(.douta(w_n8717_0[0]),.doutb(w_n8717_0[1]),.din(n8717));
	jspl jspl_w_n8723_0(.douta(w_n8723_0[0]),.doutb(w_n8723_0[1]),.din(n8723));
	jspl jspl_w_n8724_0(.douta(w_n8724_0[0]),.doutb(w_n8724_0[1]),.din(n8724));
	jspl jspl_w_n8726_0(.douta(w_n8726_0[0]),.doutb(w_n8726_0[1]),.din(n8726));
	jspl jspl_w_n8728_0(.douta(w_n8728_0[0]),.doutb(w_n8728_0[1]),.din(n8728));
	jspl jspl_w_n8731_0(.douta(w_n8731_0[0]),.doutb(w_n8731_0[1]),.din(n8731));
	jspl jspl_w_n8737_0(.douta(w_n8737_0[0]),.doutb(w_n8737_0[1]),.din(n8737));
	jspl jspl_w_n8739_0(.douta(w_n8739_0[0]),.doutb(w_n8739_0[1]),.din(n8739));
	jspl3 jspl3_w_n8740_0(.douta(w_n8740_0[0]),.doutb(w_n8740_0[1]),.doutc(w_n8740_0[2]),.din(n8740));
	jspl jspl_w_n8744_0(.douta(w_n8744_0[0]),.doutb(w_n8744_0[1]),.din(n8744));
	jspl jspl_w_n8745_0(.douta(w_n8745_0[0]),.doutb(w_n8745_0[1]),.din(n8745));
	jspl3 jspl3_w_n8746_0(.douta(w_n8746_0[0]),.doutb(w_n8746_0[1]),.doutc(w_n8746_0[2]),.din(n8746));
	jspl jspl_w_n8748_0(.douta(w_n8748_0[0]),.doutb(w_n8748_0[1]),.din(n8748));
	jspl jspl_w_n8753_0(.douta(w_n8753_0[0]),.doutb(w_n8753_0[1]),.din(n8753));
	jspl jspl_w_n8755_0(.douta(w_n8755_0[0]),.doutb(w_n8755_0[1]),.din(n8755));
	jspl jspl_w_n8756_0(.douta(w_n8756_0[0]),.doutb(w_n8756_0[1]),.din(n8756));
	jspl3 jspl3_w_n8757_0(.douta(w_n8757_0[0]),.doutb(w_n8757_0[1]),.doutc(w_n8757_0[2]),.din(n8757));
	jspl jspl_w_n8758_0(.douta(w_n8758_0[0]),.doutb(w_n8758_0[1]),.din(n8758));
	jspl jspl_w_n8762_0(.douta(w_n8762_0[0]),.doutb(w_n8762_0[1]),.din(n8762));
	jspl jspl_w_n8768_0(.douta(w_n8768_0[0]),.doutb(w_n8768_0[1]),.din(n8768));
	jspl jspl_w_n8769_0(.douta(w_n8769_0[0]),.doutb(w_n8769_0[1]),.din(n8769));
	jspl jspl_w_n8771_0(.douta(w_n8771_0[0]),.doutb(w_n8771_0[1]),.din(n8771));
	jspl jspl_w_n8773_0(.douta(w_n8773_0[0]),.doutb(w_n8773_0[1]),.din(n8773));
	jspl jspl_w_n8776_0(.douta(w_n8776_0[0]),.doutb(w_n8776_0[1]),.din(n8776));
	jspl jspl_w_n8782_0(.douta(w_n8782_0[0]),.doutb(w_n8782_0[1]),.din(n8782));
	jspl jspl_w_n8784_0(.douta(w_n8784_0[0]),.doutb(w_n8784_0[1]),.din(n8784));
	jspl3 jspl3_w_n8785_0(.douta(w_n8785_0[0]),.doutb(w_n8785_0[1]),.doutc(w_n8785_0[2]),.din(n8785));
	jspl jspl_w_n8789_0(.douta(w_n8789_0[0]),.doutb(w_n8789_0[1]),.din(n8789));
	jspl jspl_w_n8790_0(.douta(w_n8790_0[0]),.doutb(w_n8790_0[1]),.din(n8790));
	jspl3 jspl3_w_n8791_0(.douta(w_n8791_0[0]),.doutb(w_n8791_0[1]),.doutc(w_n8791_0[2]),.din(n8791));
	jspl jspl_w_n8793_0(.douta(w_n8793_0[0]),.doutb(w_n8793_0[1]),.din(n8793));
	jspl jspl_w_n8798_0(.douta(w_n8798_0[0]),.doutb(w_n8798_0[1]),.din(n8798));
	jspl jspl_w_n8800_0(.douta(w_n8800_0[0]),.doutb(w_n8800_0[1]),.din(n8800));
	jspl jspl_w_n8801_0(.douta(w_n8801_0[0]),.doutb(w_n8801_0[1]),.din(n8801));
	jspl3 jspl3_w_n8802_0(.douta(w_n8802_0[0]),.doutb(w_n8802_0[1]),.doutc(w_n8802_0[2]),.din(n8802));
	jspl jspl_w_n8803_0(.douta(w_n8803_0[0]),.doutb(w_n8803_0[1]),.din(n8803));
	jspl jspl_w_n8807_0(.douta(w_n8807_0[0]),.doutb(w_n8807_0[1]),.din(n8807));
	jspl jspl_w_n8813_0(.douta(w_n8813_0[0]),.doutb(w_n8813_0[1]),.din(n8813));
	jspl jspl_w_n8814_0(.douta(w_n8814_0[0]),.doutb(w_n8814_0[1]),.din(n8814));
	jspl jspl_w_n8816_0(.douta(w_n8816_0[0]),.doutb(w_n8816_0[1]),.din(n8816));
	jspl jspl_w_n8818_0(.douta(w_n8818_0[0]),.doutb(w_n8818_0[1]),.din(n8818));
	jspl jspl_w_n8821_0(.douta(w_n8821_0[0]),.doutb(w_n8821_0[1]),.din(n8821));
	jspl jspl_w_n8827_0(.douta(w_n8827_0[0]),.doutb(w_n8827_0[1]),.din(n8827));
	jspl jspl_w_n8829_0(.douta(w_n8829_0[0]),.doutb(w_n8829_0[1]),.din(n8829));
	jspl3 jspl3_w_n8830_0(.douta(w_n8830_0[0]),.doutb(w_n8830_0[1]),.doutc(w_n8830_0[2]),.din(n8830));
	jspl jspl_w_n8834_0(.douta(w_n8834_0[0]),.doutb(w_n8834_0[1]),.din(n8834));
	jspl jspl_w_n8835_0(.douta(w_n8835_0[0]),.doutb(w_n8835_0[1]),.din(n8835));
	jspl3 jspl3_w_n8836_0(.douta(w_n8836_0[0]),.doutb(w_n8836_0[1]),.doutc(w_n8836_0[2]),.din(n8836));
	jspl jspl_w_n8838_0(.douta(w_n8838_0[0]),.doutb(w_n8838_0[1]),.din(n8838));
	jspl jspl_w_n8843_0(.douta(w_n8843_0[0]),.doutb(w_n8843_0[1]),.din(n8843));
	jspl jspl_w_n8845_0(.douta(w_n8845_0[0]),.doutb(w_n8845_0[1]),.din(n8845));
	jspl jspl_w_n8846_0(.douta(w_n8846_0[0]),.doutb(w_n8846_0[1]),.din(n8846));
	jspl3 jspl3_w_n8847_0(.douta(w_n8847_0[0]),.doutb(w_n8847_0[1]),.doutc(w_n8847_0[2]),.din(n8847));
	jspl jspl_w_n8848_0(.douta(w_n8848_0[0]),.doutb(w_n8848_0[1]),.din(n8848));
	jspl jspl_w_n8852_0(.douta(w_n8852_0[0]),.doutb(w_n8852_0[1]),.din(n8852));
	jspl jspl_w_n8858_0(.douta(w_n8858_0[0]),.doutb(w_n8858_0[1]),.din(n8858));
	jspl jspl_w_n8859_0(.douta(w_n8859_0[0]),.doutb(w_n8859_0[1]),.din(n8859));
	jspl jspl_w_n8861_0(.douta(w_n8861_0[0]),.doutb(w_n8861_0[1]),.din(n8861));
	jspl jspl_w_n8863_0(.douta(w_n8863_0[0]),.doutb(w_n8863_0[1]),.din(n8863));
	jspl jspl_w_n8866_0(.douta(w_n8866_0[0]),.doutb(w_n8866_0[1]),.din(n8866));
	jspl jspl_w_n8872_0(.douta(w_n8872_0[0]),.doutb(w_n8872_0[1]),.din(n8872));
	jspl3 jspl3_w_n8874_0(.douta(w_n8874_0[0]),.doutb(w_n8874_0[1]),.doutc(w_n8874_0[2]),.din(n8874));
	jspl3 jspl3_w_n8874_1(.douta(w_n8874_1[0]),.doutb(w_n8874_1[1]),.doutc(w_n8874_1[2]),.din(w_n8874_0[0]));
	jspl jspl_w_n8877_0(.douta(w_n8877_0[0]),.doutb(w_n8877_0[1]),.din(n8877));
	jspl3 jspl3_w_n8878_0(.douta(w_n8878_0[0]),.doutb(w_n8878_0[1]),.doutc(w_n8878_0[2]),.din(n8878));
	jspl jspl_w_n8879_0(.douta(w_n8879_0[0]),.doutb(w_n8879_0[1]),.din(n8879));
	jspl jspl_w_n8885_0(.douta(w_n8885_0[0]),.doutb(w_n8885_0[1]),.din(n8885));
	jspl3 jspl3_w_n8886_0(.douta(w_n8886_0[0]),.doutb(w_n8886_0[1]),.doutc(w_n8886_0[2]),.din(n8886));
	jspl jspl_w_n8887_0(.douta(w_n8887_0[0]),.doutb(w_n8887_0[1]),.din(n8887));
	jspl jspl_w_n8892_0(.douta(w_n8892_0[0]),.doutb(w_n8892_0[1]),.din(n8892));
	jspl3 jspl3_w_n8893_0(.douta(w_n8893_0[0]),.doutb(w_n8893_0[1]),.doutc(w_n8893_0[2]),.din(n8893));
	jspl3 jspl3_w_n8893_1(.douta(w_n8893_1[0]),.doutb(w_n8893_1[1]),.doutc(w_n8893_1[2]),.din(w_n8893_0[0]));
	jspl3 jspl3_w_n8893_2(.douta(w_n8893_2[0]),.doutb(w_n8893_2[1]),.doutc(w_n8893_2[2]),.din(w_n8893_0[1]));
	jspl3 jspl3_w_n8893_3(.douta(w_n8893_3[0]),.doutb(w_n8893_3[1]),.doutc(w_n8893_3[2]),.din(w_n8893_0[2]));
	jspl3 jspl3_w_n8893_4(.douta(w_n8893_4[0]),.doutb(w_n8893_4[1]),.doutc(w_n8893_4[2]),.din(w_n8893_1[0]));
	jspl3 jspl3_w_n8893_5(.douta(w_n8893_5[0]),.doutb(w_n8893_5[1]),.doutc(w_n8893_5[2]),.din(w_n8893_1[1]));
	jspl3 jspl3_w_n8893_6(.douta(w_n8893_6[0]),.doutb(w_n8893_6[1]),.doutc(w_n8893_6[2]),.din(w_n8893_1[2]));
	jspl3 jspl3_w_n8893_7(.douta(w_n8893_7[0]),.doutb(w_n8893_7[1]),.doutc(w_n8893_7[2]),.din(w_n8893_2[0]));
	jspl3 jspl3_w_n8893_8(.douta(w_n8893_8[0]),.doutb(w_n8893_8[1]),.doutc(w_n8893_8[2]),.din(w_n8893_2[1]));
	jspl3 jspl3_w_n8893_9(.douta(w_n8893_9[0]),.doutb(w_n8893_9[1]),.doutc(w_n8893_9[2]),.din(w_n8893_2[2]));
	jspl3 jspl3_w_n8893_10(.douta(w_n8893_10[0]),.doutb(w_n8893_10[1]),.doutc(w_n8893_10[2]),.din(w_n8893_3[0]));
	jspl3 jspl3_w_n8893_11(.douta(w_n8893_11[0]),.doutb(w_n8893_11[1]),.doutc(w_n8893_11[2]),.din(w_n8893_3[1]));
	jspl3 jspl3_w_n8893_12(.douta(w_n8893_12[0]),.doutb(w_n8893_12[1]),.doutc(w_n8893_12[2]),.din(w_n8893_3[2]));
	jspl3 jspl3_w_n8893_13(.douta(w_n8893_13[0]),.doutb(w_n8893_13[1]),.doutc(w_n8893_13[2]),.din(w_n8893_4[0]));
	jspl3 jspl3_w_n8893_14(.douta(w_n8893_14[0]),.doutb(w_n8893_14[1]),.doutc(w_n8893_14[2]),.din(w_n8893_4[1]));
	jspl3 jspl3_w_n8893_15(.douta(w_n8893_15[0]),.doutb(w_n8893_15[1]),.doutc(w_n8893_15[2]),.din(w_n8893_4[2]));
	jspl3 jspl3_w_n8898_0(.douta(w_n8898_0[0]),.doutb(w_n8898_0[1]),.doutc(w_n8898_0[2]),.din(n8898));
	jspl3 jspl3_w_n8898_1(.douta(w_n8898_1[0]),.doutb(w_n8898_1[1]),.doutc(w_n8898_1[2]),.din(w_n8898_0[0]));
	jspl3 jspl3_w_n8898_2(.douta(w_n8898_2[0]),.doutb(w_n8898_2[1]),.doutc(w_n8898_2[2]),.din(w_n8898_0[1]));
	jspl3 jspl3_w_n8898_3(.douta(w_n8898_3[0]),.doutb(w_n8898_3[1]),.doutc(w_n8898_3[2]),.din(w_n8898_0[2]));
	jspl3 jspl3_w_n8898_4(.douta(w_n8898_4[0]),.doutb(w_n8898_4[1]),.doutc(w_n8898_4[2]),.din(w_n8898_1[0]));
	jspl3 jspl3_w_n8898_5(.douta(w_n8898_5[0]),.doutb(w_n8898_5[1]),.doutc(w_n8898_5[2]),.din(w_n8898_1[1]));
	jspl3 jspl3_w_n8898_6(.douta(w_n8898_6[0]),.doutb(w_n8898_6[1]),.doutc(w_n8898_6[2]),.din(w_n8898_1[2]));
	jspl3 jspl3_w_n8898_7(.douta(w_n8898_7[0]),.doutb(w_n8898_7[1]),.doutc(w_n8898_7[2]),.din(w_n8898_2[0]));
	jspl3 jspl3_w_n8898_8(.douta(w_n8898_8[0]),.doutb(w_n8898_8[1]),.doutc(w_n8898_8[2]),.din(w_n8898_2[1]));
	jspl3 jspl3_w_n8898_9(.douta(w_n8898_9[0]),.doutb(w_n8898_9[1]),.doutc(w_n8898_9[2]),.din(w_n8898_2[2]));
	jspl3 jspl3_w_n8898_10(.douta(w_n8898_10[0]),.doutb(w_n8898_10[1]),.doutc(w_n8898_10[2]),.din(w_n8898_3[0]));
	jspl3 jspl3_w_n8898_11(.douta(w_n8898_11[0]),.doutb(w_n8898_11[1]),.doutc(w_n8898_11[2]),.din(w_n8898_3[1]));
	jspl3 jspl3_w_n8898_12(.douta(w_n8898_12[0]),.doutb(w_n8898_12[1]),.doutc(w_n8898_12[2]),.din(w_n8898_3[2]));
	jspl3 jspl3_w_n8898_13(.douta(w_n8898_13[0]),.doutb(w_n8898_13[1]),.doutc(w_n8898_13[2]),.din(w_n8898_4[0]));
	jspl3 jspl3_w_n8898_14(.douta(w_n8898_14[0]),.doutb(w_n8898_14[1]),.doutc(w_n8898_14[2]),.din(w_n8898_4[1]));
	jspl3 jspl3_w_n8898_15(.douta(w_n8898_15[0]),.doutb(w_n8898_15[1]),.doutc(w_n8898_15[2]),.din(w_n8898_4[2]));
	jspl3 jspl3_w_n8898_16(.douta(w_n8898_16[0]),.doutb(w_n8898_16[1]),.doutc(w_n8898_16[2]),.din(w_n8898_5[0]));
	jspl3 jspl3_w_n8898_17(.douta(w_n8898_17[0]),.doutb(w_n8898_17[1]),.doutc(w_n8898_17[2]),.din(w_n8898_5[1]));
	jspl3 jspl3_w_n8898_18(.douta(w_n8898_18[0]),.doutb(w_n8898_18[1]),.doutc(w_n8898_18[2]),.din(w_n8898_5[2]));
	jspl3 jspl3_w_n8898_19(.douta(w_n8898_19[0]),.doutb(w_n8898_19[1]),.doutc(w_n8898_19[2]),.din(w_n8898_6[0]));
	jspl3 jspl3_w_n8898_20(.douta(w_n8898_20[0]),.doutb(w_n8898_20[1]),.doutc(w_n8898_20[2]),.din(w_n8898_6[1]));
	jspl3 jspl3_w_n8898_21(.douta(w_n8898_21[0]),.doutb(w_n8898_21[1]),.doutc(w_n8898_21[2]),.din(w_n8898_6[2]));
	jspl3 jspl3_w_n8898_22(.douta(w_n8898_22[0]),.doutb(w_n8898_22[1]),.doutc(w_n8898_22[2]),.din(w_n8898_7[0]));
	jspl3 jspl3_w_n8898_23(.douta(w_n8898_23[0]),.doutb(w_n8898_23[1]),.doutc(w_n8898_23[2]),.din(w_n8898_7[1]));
	jspl3 jspl3_w_n8898_24(.douta(w_n8898_24[0]),.doutb(w_n8898_24[1]),.doutc(w_n8898_24[2]),.din(w_n8898_7[2]));
	jspl3 jspl3_w_n8898_25(.douta(w_n8898_25[0]),.doutb(w_n8898_25[1]),.doutc(w_n8898_25[2]),.din(w_n8898_8[0]));
	jspl3 jspl3_w_n8898_26(.douta(w_n8898_26[0]),.doutb(w_n8898_26[1]),.doutc(w_n8898_26[2]),.din(w_n8898_8[1]));
	jspl jspl_w_n8898_27(.douta(w_n8898_27[0]),.doutb(w_n8898_27[1]),.din(w_n8898_8[2]));
	jspl jspl_w_n8901_0(.douta(w_n8901_0[0]),.doutb(w_n8901_0[1]),.din(n8901));
	jspl3 jspl3_w_n8903_0(.douta(w_n8903_0[0]),.doutb(w_n8903_0[1]),.doutc(w_n8903_0[2]),.din(n8903));
	jspl jspl_w_n8903_1(.douta(w_n8903_1[0]),.doutb(w_n8903_1[1]),.din(w_n8903_0[0]));
	jspl3 jspl3_w_n8904_0(.douta(w_n8904_0[0]),.doutb(w_n8904_0[1]),.doutc(w_n8904_0[2]),.din(n8904));
	jspl3 jspl3_w_n8908_0(.douta(w_n8908_0[0]),.doutb(w_n8908_0[1]),.doutc(w_n8908_0[2]),.din(n8908));
	jspl jspl_w_n8909_0(.douta(w_n8909_0[0]),.doutb(w_n8909_0[1]),.din(n8909));
	jspl jspl_w_n8910_0(.douta(w_n8910_0[0]),.doutb(w_n8910_0[1]),.din(n8910));
	jspl jspl_w_n8911_0(.douta(w_n8911_0[0]),.doutb(w_n8911_0[1]),.din(n8911));
	jspl jspl_w_n8913_0(.douta(w_n8913_0[0]),.doutb(w_n8913_0[1]),.din(n8913));
	jspl jspl_w_n8915_0(.douta(w_n8915_0[0]),.doutb(w_n8915_0[1]),.din(n8915));
	jspl jspl_w_n8917_0(.douta(w_n8917_0[0]),.doutb(w_n8917_0[1]),.din(n8917));
	jspl jspl_w_n8920_0(.douta(w_n8920_0[0]),.doutb(w_n8920_0[1]),.din(n8920));
	jspl jspl_w_n8925_0(.douta(w_n8925_0[0]),.doutb(w_n8925_0[1]),.din(n8925));
	jspl3 jspl3_w_n8927_0(.douta(w_n8927_0[0]),.doutb(w_n8927_0[1]),.doutc(w_n8927_0[2]),.din(n8927));
	jspl jspl_w_n8928_0(.douta(w_n8928_0[0]),.doutb(w_n8928_0[1]),.din(n8928));
	jspl jspl_w_n8932_0(.douta(w_n8932_0[0]),.doutb(w_n8932_0[1]),.din(n8932));
	jspl jspl_w_n8933_0(.douta(w_n8933_0[0]),.doutb(w_n8933_0[1]),.din(n8933));
	jspl jspl_w_n8935_0(.douta(w_n8935_0[0]),.doutb(w_n8935_0[1]),.din(n8935));
	jspl jspl_w_n8939_0(.douta(w_n8939_0[0]),.doutb(w_n8939_0[1]),.din(n8939));
	jspl jspl_w_n8941_0(.douta(w_n8941_0[0]),.doutb(w_n8941_0[1]),.din(n8941));
	jspl jspl_w_n8942_0(.douta(w_n8942_0[0]),.doutb(w_n8942_0[1]),.din(n8942));
	jspl3 jspl3_w_n8943_0(.douta(w_n8943_0[0]),.doutb(w_n8943_0[1]),.doutc(w_n8943_0[2]),.din(n8943));
	jspl jspl_w_n8944_0(.douta(w_n8944_0[0]),.doutb(w_n8944_0[1]),.din(n8944));
	jspl jspl_w_n8948_0(.douta(w_n8948_0[0]),.doutb(w_n8948_0[1]),.din(n8948));
	jspl jspl_w_n8950_0(.douta(w_n8950_0[0]),.doutb(w_n8950_0[1]),.din(n8950));
	jspl jspl_w_n8952_0(.douta(w_n8952_0[0]),.doutb(w_n8952_0[1]),.din(n8952));
	jspl jspl_w_n8954_0(.douta(w_n8954_0[0]),.doutb(w_n8954_0[1]),.din(n8954));
	jspl jspl_w_n8957_0(.douta(w_n8957_0[0]),.doutb(w_n8957_0[1]),.din(n8957));
	jspl jspl_w_n8963_0(.douta(w_n8963_0[0]),.doutb(w_n8963_0[1]),.din(n8963));
	jspl3 jspl3_w_n8965_0(.douta(w_n8965_0[0]),.doutb(w_n8965_0[1]),.doutc(w_n8965_0[2]),.din(n8965));
	jspl jspl_w_n8966_0(.douta(w_n8966_0[0]),.doutb(w_n8966_0[1]),.din(n8966));
	jspl jspl_w_n8971_0(.douta(w_n8971_0[0]),.doutb(w_n8971_0[1]),.din(n8971));
	jspl jspl_w_n8973_0(.douta(w_n8973_0[0]),.doutb(w_n8973_0[1]),.din(n8973));
	jspl jspl_w_n8975_0(.douta(w_n8975_0[0]),.doutb(w_n8975_0[1]),.din(n8975));
	jspl jspl_w_n8979_0(.douta(w_n8979_0[0]),.doutb(w_n8979_0[1]),.din(n8979));
	jspl jspl_w_n8981_0(.douta(w_n8981_0[0]),.doutb(w_n8981_0[1]),.din(n8981));
	jspl jspl_w_n8982_0(.douta(w_n8982_0[0]),.doutb(w_n8982_0[1]),.din(n8982));
	jspl3 jspl3_w_n8983_0(.douta(w_n8983_0[0]),.doutb(w_n8983_0[1]),.doutc(w_n8983_0[2]),.din(n8983));
	jspl jspl_w_n8984_0(.douta(w_n8984_0[0]),.doutb(w_n8984_0[1]),.din(n8984));
	jspl jspl_w_n8990_0(.douta(w_n8990_0[0]),.doutb(w_n8990_0[1]),.din(n8990));
	jspl jspl_w_n8991_0(.douta(w_n8991_0[0]),.doutb(w_n8991_0[1]),.din(n8991));
	jspl jspl_w_n8993_0(.douta(w_n8993_0[0]),.doutb(w_n8993_0[1]),.din(n8993));
	jspl jspl_w_n8995_0(.douta(w_n8995_0[0]),.doutb(w_n8995_0[1]),.din(n8995));
	jspl jspl_w_n8997_0(.douta(w_n8997_0[0]),.doutb(w_n8997_0[1]),.din(n8997));
	jspl jspl_w_n9003_0(.douta(w_n9003_0[0]),.doutb(w_n9003_0[1]),.din(n9003));
	jspl jspl_w_n9005_0(.douta(w_n9005_0[0]),.doutb(w_n9005_0[1]),.din(n9005));
	jspl3 jspl3_w_n9006_0(.douta(w_n9006_0[0]),.doutb(w_n9006_0[1]),.doutc(w_n9006_0[2]),.din(n9006));
	jspl jspl_w_n9009_0(.douta(w_n9009_0[0]),.doutb(w_n9009_0[1]),.din(n9009));
	jspl jspl_w_n9010_0(.douta(w_n9010_0[0]),.doutb(w_n9010_0[1]),.din(n9010));
	jspl3 jspl3_w_n9011_0(.douta(w_n9011_0[0]),.doutb(w_n9011_0[1]),.doutc(w_n9011_0[2]),.din(n9011));
	jspl jspl_w_n9013_0(.douta(w_n9013_0[0]),.doutb(w_n9013_0[1]),.din(n9013));
	jspl jspl_w_n9017_0(.douta(w_n9017_0[0]),.doutb(w_n9017_0[1]),.din(n9017));
	jspl jspl_w_n9019_0(.douta(w_n9019_0[0]),.doutb(w_n9019_0[1]),.din(n9019));
	jspl jspl_w_n9020_0(.douta(w_n9020_0[0]),.doutb(w_n9020_0[1]),.din(n9020));
	jspl3 jspl3_w_n9021_0(.douta(w_n9021_0[0]),.doutb(w_n9021_0[1]),.doutc(w_n9021_0[2]),.din(n9021));
	jspl jspl_w_n9022_0(.douta(w_n9022_0[0]),.doutb(w_n9022_0[1]),.din(n9022));
	jspl jspl_w_n9025_0(.douta(w_n9025_0[0]),.doutb(w_n9025_0[1]),.din(n9025));
	jspl jspl_w_n9031_0(.douta(w_n9031_0[0]),.doutb(w_n9031_0[1]),.din(n9031));
	jspl jspl_w_n9032_0(.douta(w_n9032_0[0]),.doutb(w_n9032_0[1]),.din(n9032));
	jspl jspl_w_n9034_0(.douta(w_n9034_0[0]),.doutb(w_n9034_0[1]),.din(n9034));
	jspl jspl_w_n9036_0(.douta(w_n9036_0[0]),.doutb(w_n9036_0[1]),.din(n9036));
	jspl jspl_w_n9038_0(.douta(w_n9038_0[0]),.doutb(w_n9038_0[1]),.din(n9038));
	jspl jspl_w_n9044_0(.douta(w_n9044_0[0]),.doutb(w_n9044_0[1]),.din(n9044));
	jspl jspl_w_n9046_0(.douta(w_n9046_0[0]),.doutb(w_n9046_0[1]),.din(n9046));
	jspl3 jspl3_w_n9047_0(.douta(w_n9047_0[0]),.doutb(w_n9047_0[1]),.doutc(w_n9047_0[2]),.din(n9047));
	jspl jspl_w_n9050_0(.douta(w_n9050_0[0]),.doutb(w_n9050_0[1]),.din(n9050));
	jspl jspl_w_n9051_0(.douta(w_n9051_0[0]),.doutb(w_n9051_0[1]),.din(n9051));
	jspl3 jspl3_w_n9052_0(.douta(w_n9052_0[0]),.doutb(w_n9052_0[1]),.doutc(w_n9052_0[2]),.din(n9052));
	jspl jspl_w_n9054_0(.douta(w_n9054_0[0]),.doutb(w_n9054_0[1]),.din(n9054));
	jspl jspl_w_n9056_0(.douta(w_n9056_0[0]),.doutb(w_n9056_0[1]),.din(n9056));
	jspl jspl_w_n9058_0(.douta(w_n9058_0[0]),.doutb(w_n9058_0[1]),.din(n9058));
	jspl jspl_w_n9064_0(.douta(w_n9064_0[0]),.doutb(w_n9064_0[1]),.din(n9064));
	jspl3 jspl3_w_n9066_0(.douta(w_n9066_0[0]),.doutb(w_n9066_0[1]),.doutc(w_n9066_0[2]),.din(n9066));
	jspl jspl_w_n9067_0(.douta(w_n9067_0[0]),.doutb(w_n9067_0[1]),.din(n9067));
	jspl jspl_w_n9070_0(.douta(w_n9070_0[0]),.doutb(w_n9070_0[1]),.din(n9070));
	jspl jspl_w_n9072_0(.douta(w_n9072_0[0]),.doutb(w_n9072_0[1]),.din(n9072));
	jspl jspl_w_n9076_0(.douta(w_n9076_0[0]),.doutb(w_n9076_0[1]),.din(n9076));
	jspl jspl_w_n9078_0(.douta(w_n9078_0[0]),.doutb(w_n9078_0[1]),.din(n9078));
	jspl jspl_w_n9079_0(.douta(w_n9079_0[0]),.doutb(w_n9079_0[1]),.din(n9079));
	jspl jspl_w_n9080_0(.douta(w_n9080_0[0]),.doutb(w_n9080_0[1]),.din(n9080));
	jspl3 jspl3_w_n9081_0(.douta(w_n9081_0[0]),.doutb(w_n9081_0[1]),.doutc(w_n9081_0[2]),.din(n9081));
	jspl jspl_w_n9084_0(.douta(w_n9084_0[0]),.doutb(w_n9084_0[1]),.din(n9084));
	jspl jspl_w_n9085_0(.douta(w_n9085_0[0]),.doutb(w_n9085_0[1]),.din(n9085));
	jspl3 jspl3_w_n9086_0(.douta(w_n9086_0[0]),.doutb(w_n9086_0[1]),.doutc(w_n9086_0[2]),.din(n9086));
	jspl jspl_w_n9088_0(.douta(w_n9088_0[0]),.doutb(w_n9088_0[1]),.din(n9088));
	jspl jspl_w_n9092_0(.douta(w_n9092_0[0]),.doutb(w_n9092_0[1]),.din(n9092));
	jspl jspl_w_n9094_0(.douta(w_n9094_0[0]),.doutb(w_n9094_0[1]),.din(n9094));
	jspl jspl_w_n9095_0(.douta(w_n9095_0[0]),.doutb(w_n9095_0[1]),.din(n9095));
	jspl3 jspl3_w_n9096_0(.douta(w_n9096_0[0]),.doutb(w_n9096_0[1]),.doutc(w_n9096_0[2]),.din(n9096));
	jspl jspl_w_n9097_0(.douta(w_n9097_0[0]),.doutb(w_n9097_0[1]),.din(n9097));
	jspl jspl_w_n9100_0(.douta(w_n9100_0[0]),.doutb(w_n9100_0[1]),.din(n9100));
	jspl jspl_w_n9106_0(.douta(w_n9106_0[0]),.doutb(w_n9106_0[1]),.din(n9106));
	jspl jspl_w_n9107_0(.douta(w_n9107_0[0]),.doutb(w_n9107_0[1]),.din(n9107));
	jspl jspl_w_n9109_0(.douta(w_n9109_0[0]),.doutb(w_n9109_0[1]),.din(n9109));
	jspl jspl_w_n9111_0(.douta(w_n9111_0[0]),.doutb(w_n9111_0[1]),.din(n9111));
	jspl jspl_w_n9113_0(.douta(w_n9113_0[0]),.doutb(w_n9113_0[1]),.din(n9113));
	jspl jspl_w_n9119_0(.douta(w_n9119_0[0]),.doutb(w_n9119_0[1]),.din(n9119));
	jspl jspl_w_n9121_0(.douta(w_n9121_0[0]),.doutb(w_n9121_0[1]),.din(n9121));
	jspl3 jspl3_w_n9122_0(.douta(w_n9122_0[0]),.doutb(w_n9122_0[1]),.doutc(w_n9122_0[2]),.din(n9122));
	jspl jspl_w_n9125_0(.douta(w_n9125_0[0]),.doutb(w_n9125_0[1]),.din(n9125));
	jspl jspl_w_n9126_0(.douta(w_n9126_0[0]),.doutb(w_n9126_0[1]),.din(n9126));
	jspl3 jspl3_w_n9127_0(.douta(w_n9127_0[0]),.doutb(w_n9127_0[1]),.doutc(w_n9127_0[2]),.din(n9127));
	jspl jspl_w_n9129_0(.douta(w_n9129_0[0]),.doutb(w_n9129_0[1]),.din(n9129));
	jspl jspl_w_n9133_0(.douta(w_n9133_0[0]),.doutb(w_n9133_0[1]),.din(n9133));
	jspl jspl_w_n9135_0(.douta(w_n9135_0[0]),.doutb(w_n9135_0[1]),.din(n9135));
	jspl jspl_w_n9136_0(.douta(w_n9136_0[0]),.doutb(w_n9136_0[1]),.din(n9136));
	jspl3 jspl3_w_n9137_0(.douta(w_n9137_0[0]),.doutb(w_n9137_0[1]),.doutc(w_n9137_0[2]),.din(n9137));
	jspl jspl_w_n9138_0(.douta(w_n9138_0[0]),.doutb(w_n9138_0[1]),.din(n9138));
	jspl jspl_w_n9141_0(.douta(w_n9141_0[0]),.doutb(w_n9141_0[1]),.din(n9141));
	jspl jspl_w_n9147_0(.douta(w_n9147_0[0]),.doutb(w_n9147_0[1]),.din(n9147));
	jspl jspl_w_n9148_0(.douta(w_n9148_0[0]),.doutb(w_n9148_0[1]),.din(n9148));
	jspl jspl_w_n9150_0(.douta(w_n9150_0[0]),.doutb(w_n9150_0[1]),.din(n9150));
	jspl jspl_w_n9152_0(.douta(w_n9152_0[0]),.doutb(w_n9152_0[1]),.din(n9152));
	jspl jspl_w_n9154_0(.douta(w_n9154_0[0]),.doutb(w_n9154_0[1]),.din(n9154));
	jspl jspl_w_n9160_0(.douta(w_n9160_0[0]),.doutb(w_n9160_0[1]),.din(n9160));
	jspl jspl_w_n9162_0(.douta(w_n9162_0[0]),.doutb(w_n9162_0[1]),.din(n9162));
	jspl3 jspl3_w_n9163_0(.douta(w_n9163_0[0]),.doutb(w_n9163_0[1]),.doutc(w_n9163_0[2]),.din(n9163));
	jspl jspl_w_n9166_0(.douta(w_n9166_0[0]),.doutb(w_n9166_0[1]),.din(n9166));
	jspl jspl_w_n9167_0(.douta(w_n9167_0[0]),.doutb(w_n9167_0[1]),.din(n9167));
	jspl3 jspl3_w_n9168_0(.douta(w_n9168_0[0]),.doutb(w_n9168_0[1]),.doutc(w_n9168_0[2]),.din(n9168));
	jspl jspl_w_n9170_0(.douta(w_n9170_0[0]),.doutb(w_n9170_0[1]),.din(n9170));
	jspl jspl_w_n9174_0(.douta(w_n9174_0[0]),.doutb(w_n9174_0[1]),.din(n9174));
	jspl jspl_w_n9176_0(.douta(w_n9176_0[0]),.doutb(w_n9176_0[1]),.din(n9176));
	jspl jspl_w_n9177_0(.douta(w_n9177_0[0]),.doutb(w_n9177_0[1]),.din(n9177));
	jspl3 jspl3_w_n9178_0(.douta(w_n9178_0[0]),.doutb(w_n9178_0[1]),.doutc(w_n9178_0[2]),.din(n9178));
	jspl jspl_w_n9179_0(.douta(w_n9179_0[0]),.doutb(w_n9179_0[1]),.din(n9179));
	jspl jspl_w_n9182_0(.douta(w_n9182_0[0]),.doutb(w_n9182_0[1]),.din(n9182));
	jspl jspl_w_n9188_0(.douta(w_n9188_0[0]),.doutb(w_n9188_0[1]),.din(n9188));
	jspl jspl_w_n9189_0(.douta(w_n9189_0[0]),.doutb(w_n9189_0[1]),.din(n9189));
	jspl jspl_w_n9191_0(.douta(w_n9191_0[0]),.doutb(w_n9191_0[1]),.din(n9191));
	jspl jspl_w_n9193_0(.douta(w_n9193_0[0]),.doutb(w_n9193_0[1]),.din(n9193));
	jspl jspl_w_n9195_0(.douta(w_n9195_0[0]),.doutb(w_n9195_0[1]),.din(n9195));
	jspl jspl_w_n9201_0(.douta(w_n9201_0[0]),.doutb(w_n9201_0[1]),.din(n9201));
	jspl jspl_w_n9203_0(.douta(w_n9203_0[0]),.doutb(w_n9203_0[1]),.din(n9203));
	jspl3 jspl3_w_n9204_0(.douta(w_n9204_0[0]),.doutb(w_n9204_0[1]),.doutc(w_n9204_0[2]),.din(n9204));
	jspl jspl_w_n9207_0(.douta(w_n9207_0[0]),.doutb(w_n9207_0[1]),.din(n9207));
	jspl jspl_w_n9208_0(.douta(w_n9208_0[0]),.doutb(w_n9208_0[1]),.din(n9208));
	jspl3 jspl3_w_n9209_0(.douta(w_n9209_0[0]),.doutb(w_n9209_0[1]),.doutc(w_n9209_0[2]),.din(n9209));
	jspl jspl_w_n9211_0(.douta(w_n9211_0[0]),.doutb(w_n9211_0[1]),.din(n9211));
	jspl jspl_w_n9215_0(.douta(w_n9215_0[0]),.doutb(w_n9215_0[1]),.din(n9215));
	jspl jspl_w_n9217_0(.douta(w_n9217_0[0]),.doutb(w_n9217_0[1]),.din(n9217));
	jspl jspl_w_n9218_0(.douta(w_n9218_0[0]),.doutb(w_n9218_0[1]),.din(n9218));
	jspl3 jspl3_w_n9219_0(.douta(w_n9219_0[0]),.doutb(w_n9219_0[1]),.doutc(w_n9219_0[2]),.din(n9219));
	jspl jspl_w_n9220_0(.douta(w_n9220_0[0]),.doutb(w_n9220_0[1]),.din(n9220));
	jspl jspl_w_n9223_0(.douta(w_n9223_0[0]),.doutb(w_n9223_0[1]),.din(n9223));
	jspl jspl_w_n9229_0(.douta(w_n9229_0[0]),.doutb(w_n9229_0[1]),.din(n9229));
	jspl jspl_w_n9230_0(.douta(w_n9230_0[0]),.doutb(w_n9230_0[1]),.din(n9230));
	jspl jspl_w_n9232_0(.douta(w_n9232_0[0]),.doutb(w_n9232_0[1]),.din(n9232));
	jspl jspl_w_n9234_0(.douta(w_n9234_0[0]),.doutb(w_n9234_0[1]),.din(n9234));
	jspl jspl_w_n9236_0(.douta(w_n9236_0[0]),.doutb(w_n9236_0[1]),.din(n9236));
	jspl jspl_w_n9242_0(.douta(w_n9242_0[0]),.doutb(w_n9242_0[1]),.din(n9242));
	jspl jspl_w_n9244_0(.douta(w_n9244_0[0]),.doutb(w_n9244_0[1]),.din(n9244));
	jspl3 jspl3_w_n9245_0(.douta(w_n9245_0[0]),.doutb(w_n9245_0[1]),.doutc(w_n9245_0[2]),.din(n9245));
	jspl jspl_w_n9248_0(.douta(w_n9248_0[0]),.doutb(w_n9248_0[1]),.din(n9248));
	jspl jspl_w_n9249_0(.douta(w_n9249_0[0]),.doutb(w_n9249_0[1]),.din(n9249));
	jspl3 jspl3_w_n9250_0(.douta(w_n9250_0[0]),.doutb(w_n9250_0[1]),.doutc(w_n9250_0[2]),.din(n9250));
	jspl jspl_w_n9252_0(.douta(w_n9252_0[0]),.doutb(w_n9252_0[1]),.din(n9252));
	jspl jspl_w_n9256_0(.douta(w_n9256_0[0]),.doutb(w_n9256_0[1]),.din(n9256));
	jspl jspl_w_n9258_0(.douta(w_n9258_0[0]),.doutb(w_n9258_0[1]),.din(n9258));
	jspl jspl_w_n9259_0(.douta(w_n9259_0[0]),.doutb(w_n9259_0[1]),.din(n9259));
	jspl3 jspl3_w_n9260_0(.douta(w_n9260_0[0]),.doutb(w_n9260_0[1]),.doutc(w_n9260_0[2]),.din(n9260));
	jspl jspl_w_n9261_0(.douta(w_n9261_0[0]),.doutb(w_n9261_0[1]),.din(n9261));
	jspl jspl_w_n9264_0(.douta(w_n9264_0[0]),.doutb(w_n9264_0[1]),.din(n9264));
	jspl jspl_w_n9270_0(.douta(w_n9270_0[0]),.doutb(w_n9270_0[1]),.din(n9270));
	jspl jspl_w_n9271_0(.douta(w_n9271_0[0]),.doutb(w_n9271_0[1]),.din(n9271));
	jspl jspl_w_n9273_0(.douta(w_n9273_0[0]),.doutb(w_n9273_0[1]),.din(n9273));
	jspl jspl_w_n9275_0(.douta(w_n9275_0[0]),.doutb(w_n9275_0[1]),.din(n9275));
	jspl jspl_w_n9277_0(.douta(w_n9277_0[0]),.doutb(w_n9277_0[1]),.din(n9277));
	jspl jspl_w_n9283_0(.douta(w_n9283_0[0]),.doutb(w_n9283_0[1]),.din(n9283));
	jspl3 jspl3_w_n9285_0(.douta(w_n9285_0[0]),.doutb(w_n9285_0[1]),.doutc(w_n9285_0[2]),.din(n9285));
	jspl jspl_w_n9290_0(.douta(w_n9290_0[0]),.doutb(w_n9290_0[1]),.din(n9290));
	jspl3 jspl3_w_n9292_0(.douta(w_n9292_0[0]),.doutb(w_n9292_0[1]),.doutc(w_n9292_0[2]),.din(n9292));
	jspl3 jspl3_w_n9296_0(.douta(w_n9296_0[0]),.doutb(w_n9296_0[1]),.doutc(w_n9296_0[2]),.din(n9296));
	jspl jspl_w_n9297_0(.douta(w_n9297_0[0]),.doutb(w_n9297_0[1]),.din(n9297));
	jspl jspl_w_n9302_0(.douta(w_n9302_0[0]),.doutb(w_n9302_0[1]),.din(n9302));
	jspl3 jspl3_w_n9303_0(.douta(w_n9303_0[0]),.doutb(w_n9303_0[1]),.doutc(w_n9303_0[2]),.din(n9303));
	jspl jspl_w_n9308_0(.douta(w_n9308_0[0]),.doutb(w_n9308_0[1]),.din(n9308));
	jspl jspl_w_n9315_0(.douta(w_n9315_0[0]),.doutb(w_n9315_0[1]),.din(n9315));
	jspl3 jspl3_w_n9318_0(.douta(w_n9318_0[0]),.doutb(w_n9318_0[1]),.doutc(w_n9318_0[2]),.din(n9318));
	jspl jspl_w_n9318_1(.douta(w_n9318_1[0]),.doutb(w_n9318_1[1]),.din(w_n9318_0[0]));
	jspl jspl_w_n9319_0(.douta(w_n9319_0[0]),.doutb(w_n9319_0[1]),.din(n9319));
	jspl3 jspl3_w_n9322_0(.douta(w_n9322_0[0]),.doutb(w_n9322_0[1]),.doutc(w_n9322_0[2]),.din(n9322));
	jspl jspl_w_n9323_0(.douta(w_n9323_0[0]),.doutb(w_n9323_0[1]),.din(n9323));
	jspl jspl_w_n9324_0(.douta(w_n9324_0[0]),.doutb(w_n9324_0[1]),.din(n9324));
	jspl jspl_w_n9325_0(.douta(w_n9325_0[0]),.doutb(w_n9325_0[1]),.din(n9325));
	jspl jspl_w_n9327_0(.douta(w_n9327_0[0]),.doutb(w_n9327_0[1]),.din(n9327));
	jspl jspl_w_n9329_0(.douta(w_n9329_0[0]),.doutb(w_n9329_0[1]),.din(n9329));
	jspl jspl_w_n9331_0(.douta(w_n9331_0[0]),.doutb(w_n9331_0[1]),.din(n9331));
	jspl jspl_w_n9340_0(.douta(w_n9340_0[0]),.doutb(w_n9340_0[1]),.din(n9340));
	jspl3 jspl3_w_n9342_0(.douta(w_n9342_0[0]),.doutb(w_n9342_0[1]),.doutc(w_n9342_0[2]),.din(n9342));
	jspl jspl_w_n9343_0(.douta(w_n9343_0[0]),.doutb(w_n9343_0[1]),.din(n9343));
	jspl jspl_w_n9347_0(.douta(w_n9347_0[0]),.doutb(w_n9347_0[1]),.din(n9347));
	jspl jspl_w_n9349_0(.douta(w_n9349_0[0]),.doutb(w_n9349_0[1]),.din(n9349));
	jspl jspl_w_n9351_0(.douta(w_n9351_0[0]),.doutb(w_n9351_0[1]),.din(n9351));
	jspl jspl_w_n9356_0(.douta(w_n9356_0[0]),.doutb(w_n9356_0[1]),.din(n9356));
	jspl jspl_w_n9358_0(.douta(w_n9358_0[0]),.doutb(w_n9358_0[1]),.din(n9358));
	jspl jspl_w_n9359_0(.douta(w_n9359_0[0]),.doutb(w_n9359_0[1]),.din(n9359));
	jspl3 jspl3_w_n9360_0(.douta(w_n9360_0[0]),.doutb(w_n9360_0[1]),.doutc(w_n9360_0[2]),.din(n9360));
	jspl jspl_w_n9361_0(.douta(w_n9361_0[0]),.doutb(w_n9361_0[1]),.din(n9361));
	jspl jspl_w_n9366_0(.douta(w_n9366_0[0]),.doutb(w_n9366_0[1]),.din(n9366));
	jspl jspl_w_n9367_0(.douta(w_n9367_0[0]),.doutb(w_n9367_0[1]),.din(n9367));
	jspl jspl_w_n9369_0(.douta(w_n9369_0[0]),.doutb(w_n9369_0[1]),.din(n9369));
	jspl jspl_w_n9371_0(.douta(w_n9371_0[0]),.doutb(w_n9371_0[1]),.din(n9371));
	jspl jspl_w_n9374_0(.douta(w_n9374_0[0]),.doutb(w_n9374_0[1]),.din(n9374));
	jspl jspl_w_n9380_0(.douta(w_n9380_0[0]),.doutb(w_n9380_0[1]),.din(n9380));
	jspl3 jspl3_w_n9382_0(.douta(w_n9382_0[0]),.doutb(w_n9382_0[1]),.doutc(w_n9382_0[2]),.din(n9382));
	jspl jspl_w_n9383_0(.douta(w_n9383_0[0]),.doutb(w_n9383_0[1]),.din(n9383));
	jspl jspl_w_n9387_0(.douta(w_n9387_0[0]),.doutb(w_n9387_0[1]),.din(n9387));
	jspl jspl_w_n9388_0(.douta(w_n9388_0[0]),.doutb(w_n9388_0[1]),.din(n9388));
	jspl jspl_w_n9390_0(.douta(w_n9390_0[0]),.doutb(w_n9390_0[1]),.din(n9390));
	jspl jspl_w_n9395_0(.douta(w_n9395_0[0]),.doutb(w_n9395_0[1]),.din(n9395));
	jspl jspl_w_n9397_0(.douta(w_n9397_0[0]),.doutb(w_n9397_0[1]),.din(n9397));
	jspl jspl_w_n9398_0(.douta(w_n9398_0[0]),.doutb(w_n9398_0[1]),.din(n9398));
	jspl3 jspl3_w_n9399_0(.douta(w_n9399_0[0]),.doutb(w_n9399_0[1]),.doutc(w_n9399_0[2]),.din(n9399));
	jspl jspl_w_n9400_0(.douta(w_n9400_0[0]),.doutb(w_n9400_0[1]),.din(n9400));
	jspl jspl_w_n9404_0(.douta(w_n9404_0[0]),.doutb(w_n9404_0[1]),.din(n9404));
	jspl jspl_w_n9405_0(.douta(w_n9405_0[0]),.doutb(w_n9405_0[1]),.din(n9405));
	jspl jspl_w_n9407_0(.douta(w_n9407_0[0]),.doutb(w_n9407_0[1]),.din(n9407));
	jspl jspl_w_n9409_0(.douta(w_n9409_0[0]),.doutb(w_n9409_0[1]),.din(n9409));
	jspl jspl_w_n9412_0(.douta(w_n9412_0[0]),.doutb(w_n9412_0[1]),.din(n9412));
	jspl jspl_w_n9418_0(.douta(w_n9418_0[0]),.doutb(w_n9418_0[1]),.din(n9418));
	jspl jspl_w_n9420_0(.douta(w_n9420_0[0]),.doutb(w_n9420_0[1]),.din(n9420));
	jspl3 jspl3_w_n9421_0(.douta(w_n9421_0[0]),.doutb(w_n9421_0[1]),.doutc(w_n9421_0[2]),.din(n9421));
	jspl jspl_w_n9425_0(.douta(w_n9425_0[0]),.doutb(w_n9425_0[1]),.din(n9425));
	jspl jspl_w_n9426_0(.douta(w_n9426_0[0]),.doutb(w_n9426_0[1]),.din(n9426));
	jspl3 jspl3_w_n9427_0(.douta(w_n9427_0[0]),.doutb(w_n9427_0[1]),.doutc(w_n9427_0[2]),.din(n9427));
	jspl jspl_w_n9429_0(.douta(w_n9429_0[0]),.doutb(w_n9429_0[1]),.din(n9429));
	jspl jspl_w_n9434_0(.douta(w_n9434_0[0]),.doutb(w_n9434_0[1]),.din(n9434));
	jspl jspl_w_n9436_0(.douta(w_n9436_0[0]),.doutb(w_n9436_0[1]),.din(n9436));
	jspl jspl_w_n9437_0(.douta(w_n9437_0[0]),.doutb(w_n9437_0[1]),.din(n9437));
	jspl3 jspl3_w_n9438_0(.douta(w_n9438_0[0]),.doutb(w_n9438_0[1]),.doutc(w_n9438_0[2]),.din(n9438));
	jspl jspl_w_n9439_0(.douta(w_n9439_0[0]),.doutb(w_n9439_0[1]),.din(n9439));
	jspl jspl_w_n9443_0(.douta(w_n9443_0[0]),.doutb(w_n9443_0[1]),.din(n9443));
	jspl jspl_w_n9449_0(.douta(w_n9449_0[0]),.doutb(w_n9449_0[1]),.din(n9449));
	jspl jspl_w_n9450_0(.douta(w_n9450_0[0]),.doutb(w_n9450_0[1]),.din(n9450));
	jspl jspl_w_n9452_0(.douta(w_n9452_0[0]),.doutb(w_n9452_0[1]),.din(n9452));
	jspl jspl_w_n9454_0(.douta(w_n9454_0[0]),.doutb(w_n9454_0[1]),.din(n9454));
	jspl jspl_w_n9457_0(.douta(w_n9457_0[0]),.doutb(w_n9457_0[1]),.din(n9457));
	jspl jspl_w_n9463_0(.douta(w_n9463_0[0]),.doutb(w_n9463_0[1]),.din(n9463));
	jspl jspl_w_n9465_0(.douta(w_n9465_0[0]),.doutb(w_n9465_0[1]),.din(n9465));
	jspl3 jspl3_w_n9466_0(.douta(w_n9466_0[0]),.doutb(w_n9466_0[1]),.doutc(w_n9466_0[2]),.din(n9466));
	jspl jspl_w_n9470_0(.douta(w_n9470_0[0]),.doutb(w_n9470_0[1]),.din(n9470));
	jspl jspl_w_n9471_0(.douta(w_n9471_0[0]),.doutb(w_n9471_0[1]),.din(n9471));
	jspl3 jspl3_w_n9472_0(.douta(w_n9472_0[0]),.doutb(w_n9472_0[1]),.doutc(w_n9472_0[2]),.din(n9472));
	jspl jspl_w_n9474_0(.douta(w_n9474_0[0]),.doutb(w_n9474_0[1]),.din(n9474));
	jspl jspl_w_n9479_0(.douta(w_n9479_0[0]),.doutb(w_n9479_0[1]),.din(n9479));
	jspl jspl_w_n9481_0(.douta(w_n9481_0[0]),.doutb(w_n9481_0[1]),.din(n9481));
	jspl jspl_w_n9482_0(.douta(w_n9482_0[0]),.doutb(w_n9482_0[1]),.din(n9482));
	jspl3 jspl3_w_n9483_0(.douta(w_n9483_0[0]),.doutb(w_n9483_0[1]),.doutc(w_n9483_0[2]),.din(n9483));
	jspl jspl_w_n9484_0(.douta(w_n9484_0[0]),.doutb(w_n9484_0[1]),.din(n9484));
	jspl jspl_w_n9488_0(.douta(w_n9488_0[0]),.doutb(w_n9488_0[1]),.din(n9488));
	jspl jspl_w_n9494_0(.douta(w_n9494_0[0]),.doutb(w_n9494_0[1]),.din(n9494));
	jspl jspl_w_n9495_0(.douta(w_n9495_0[0]),.doutb(w_n9495_0[1]),.din(n9495));
	jspl jspl_w_n9497_0(.douta(w_n9497_0[0]),.doutb(w_n9497_0[1]),.din(n9497));
	jspl jspl_w_n9502_0(.douta(w_n9502_0[0]),.doutb(w_n9502_0[1]),.din(n9502));
	jspl jspl_w_n9504_0(.douta(w_n9504_0[0]),.doutb(w_n9504_0[1]),.din(n9504));
	jspl jspl_w_n9505_0(.douta(w_n9505_0[0]),.doutb(w_n9505_0[1]),.din(n9505));
	jspl3 jspl3_w_n9506_0(.douta(w_n9506_0[0]),.doutb(w_n9506_0[1]),.doutc(w_n9506_0[2]),.din(n9506));
	jspl jspl_w_n9507_0(.douta(w_n9507_0[0]),.doutb(w_n9507_0[1]),.din(n9507));
	jspl jspl_w_n9509_0(.douta(w_n9509_0[0]),.doutb(w_n9509_0[1]),.din(n9509));
	jspl jspl_w_n9511_0(.douta(w_n9511_0[0]),.doutb(w_n9511_0[1]),.din(n9511));
	jspl jspl_w_n9513_0(.douta(w_n9513_0[0]),.doutb(w_n9513_0[1]),.din(n9513));
	jspl jspl_w_n9516_0(.douta(w_n9516_0[0]),.doutb(w_n9516_0[1]),.din(n9516));
	jspl jspl_w_n9522_0(.douta(w_n9522_0[0]),.doutb(w_n9522_0[1]),.din(n9522));
	jspl3 jspl3_w_n9524_0(.douta(w_n9524_0[0]),.doutb(w_n9524_0[1]),.doutc(w_n9524_0[2]),.din(n9524));
	jspl jspl_w_n9525_0(.douta(w_n9525_0[0]),.doutb(w_n9525_0[1]),.din(n9525));
	jspl jspl_w_n9529_0(.douta(w_n9529_0[0]),.doutb(w_n9529_0[1]),.din(n9529));
	jspl jspl_w_n9535_0(.douta(w_n9535_0[0]),.doutb(w_n9535_0[1]),.din(n9535));
	jspl jspl_w_n9536_0(.douta(w_n9536_0[0]),.doutb(w_n9536_0[1]),.din(n9536));
	jspl jspl_w_n9538_0(.douta(w_n9538_0[0]),.doutb(w_n9538_0[1]),.din(n9538));
	jspl jspl_w_n9540_0(.douta(w_n9540_0[0]),.doutb(w_n9540_0[1]),.din(n9540));
	jspl jspl_w_n9543_0(.douta(w_n9543_0[0]),.doutb(w_n9543_0[1]),.din(n9543));
	jspl jspl_w_n9549_0(.douta(w_n9549_0[0]),.doutb(w_n9549_0[1]),.din(n9549));
	jspl jspl_w_n9551_0(.douta(w_n9551_0[0]),.doutb(w_n9551_0[1]),.din(n9551));
	jspl3 jspl3_w_n9552_0(.douta(w_n9552_0[0]),.doutb(w_n9552_0[1]),.doutc(w_n9552_0[2]),.din(n9552));
	jspl jspl_w_n9556_0(.douta(w_n9556_0[0]),.doutb(w_n9556_0[1]),.din(n9556));
	jspl jspl_w_n9557_0(.douta(w_n9557_0[0]),.doutb(w_n9557_0[1]),.din(n9557));
	jspl3 jspl3_w_n9558_0(.douta(w_n9558_0[0]),.doutb(w_n9558_0[1]),.doutc(w_n9558_0[2]),.din(n9558));
	jspl jspl_w_n9560_0(.douta(w_n9560_0[0]),.doutb(w_n9560_0[1]),.din(n9560));
	jspl jspl_w_n9565_0(.douta(w_n9565_0[0]),.doutb(w_n9565_0[1]),.din(n9565));
	jspl jspl_w_n9567_0(.douta(w_n9567_0[0]),.doutb(w_n9567_0[1]),.din(n9567));
	jspl jspl_w_n9568_0(.douta(w_n9568_0[0]),.doutb(w_n9568_0[1]),.din(n9568));
	jspl3 jspl3_w_n9569_0(.douta(w_n9569_0[0]),.doutb(w_n9569_0[1]),.doutc(w_n9569_0[2]),.din(n9569));
	jspl jspl_w_n9570_0(.douta(w_n9570_0[0]),.doutb(w_n9570_0[1]),.din(n9570));
	jspl jspl_w_n9574_0(.douta(w_n9574_0[0]),.doutb(w_n9574_0[1]),.din(n9574));
	jspl jspl_w_n9580_0(.douta(w_n9580_0[0]),.doutb(w_n9580_0[1]),.din(n9580));
	jspl jspl_w_n9581_0(.douta(w_n9581_0[0]),.doutb(w_n9581_0[1]),.din(n9581));
	jspl jspl_w_n9583_0(.douta(w_n9583_0[0]),.doutb(w_n9583_0[1]),.din(n9583));
	jspl jspl_w_n9585_0(.douta(w_n9585_0[0]),.doutb(w_n9585_0[1]),.din(n9585));
	jspl jspl_w_n9588_0(.douta(w_n9588_0[0]),.doutb(w_n9588_0[1]),.din(n9588));
	jspl jspl_w_n9594_0(.douta(w_n9594_0[0]),.doutb(w_n9594_0[1]),.din(n9594));
	jspl jspl_w_n9596_0(.douta(w_n9596_0[0]),.doutb(w_n9596_0[1]),.din(n9596));
	jspl3 jspl3_w_n9597_0(.douta(w_n9597_0[0]),.doutb(w_n9597_0[1]),.doutc(w_n9597_0[2]),.din(n9597));
	jspl jspl_w_n9601_0(.douta(w_n9601_0[0]),.doutb(w_n9601_0[1]),.din(n9601));
	jspl jspl_w_n9602_0(.douta(w_n9602_0[0]),.doutb(w_n9602_0[1]),.din(n9602));
	jspl3 jspl3_w_n9603_0(.douta(w_n9603_0[0]),.doutb(w_n9603_0[1]),.doutc(w_n9603_0[2]),.din(n9603));
	jspl jspl_w_n9605_0(.douta(w_n9605_0[0]),.doutb(w_n9605_0[1]),.din(n9605));
	jspl jspl_w_n9610_0(.douta(w_n9610_0[0]),.doutb(w_n9610_0[1]),.din(n9610));
	jspl jspl_w_n9612_0(.douta(w_n9612_0[0]),.doutb(w_n9612_0[1]),.din(n9612));
	jspl jspl_w_n9613_0(.douta(w_n9613_0[0]),.doutb(w_n9613_0[1]),.din(n9613));
	jspl3 jspl3_w_n9614_0(.douta(w_n9614_0[0]),.doutb(w_n9614_0[1]),.doutc(w_n9614_0[2]),.din(n9614));
	jspl jspl_w_n9615_0(.douta(w_n9615_0[0]),.doutb(w_n9615_0[1]),.din(n9615));
	jspl jspl_w_n9619_0(.douta(w_n9619_0[0]),.doutb(w_n9619_0[1]),.din(n9619));
	jspl jspl_w_n9625_0(.douta(w_n9625_0[0]),.doutb(w_n9625_0[1]),.din(n9625));
	jspl jspl_w_n9626_0(.douta(w_n9626_0[0]),.doutb(w_n9626_0[1]),.din(n9626));
	jspl jspl_w_n9628_0(.douta(w_n9628_0[0]),.doutb(w_n9628_0[1]),.din(n9628));
	jspl jspl_w_n9630_0(.douta(w_n9630_0[0]),.doutb(w_n9630_0[1]),.din(n9630));
	jspl jspl_w_n9633_0(.douta(w_n9633_0[0]),.doutb(w_n9633_0[1]),.din(n9633));
	jspl jspl_w_n9639_0(.douta(w_n9639_0[0]),.doutb(w_n9639_0[1]),.din(n9639));
	jspl jspl_w_n9641_0(.douta(w_n9641_0[0]),.doutb(w_n9641_0[1]),.din(n9641));
	jspl3 jspl3_w_n9642_0(.douta(w_n9642_0[0]),.doutb(w_n9642_0[1]),.doutc(w_n9642_0[2]),.din(n9642));
	jspl jspl_w_n9646_0(.douta(w_n9646_0[0]),.doutb(w_n9646_0[1]),.din(n9646));
	jspl jspl_w_n9647_0(.douta(w_n9647_0[0]),.doutb(w_n9647_0[1]),.din(n9647));
	jspl3 jspl3_w_n9648_0(.douta(w_n9648_0[0]),.doutb(w_n9648_0[1]),.doutc(w_n9648_0[2]),.din(n9648));
	jspl jspl_w_n9650_0(.douta(w_n9650_0[0]),.doutb(w_n9650_0[1]),.din(n9650));
	jspl jspl_w_n9655_0(.douta(w_n9655_0[0]),.doutb(w_n9655_0[1]),.din(n9655));
	jspl jspl_w_n9657_0(.douta(w_n9657_0[0]),.doutb(w_n9657_0[1]),.din(n9657));
	jspl jspl_w_n9658_0(.douta(w_n9658_0[0]),.doutb(w_n9658_0[1]),.din(n9658));
	jspl3 jspl3_w_n9659_0(.douta(w_n9659_0[0]),.doutb(w_n9659_0[1]),.doutc(w_n9659_0[2]),.din(n9659));
	jspl jspl_w_n9660_0(.douta(w_n9660_0[0]),.doutb(w_n9660_0[1]),.din(n9660));
	jspl jspl_w_n9664_0(.douta(w_n9664_0[0]),.doutb(w_n9664_0[1]),.din(n9664));
	jspl jspl_w_n9670_0(.douta(w_n9670_0[0]),.doutb(w_n9670_0[1]),.din(n9670));
	jspl jspl_w_n9671_0(.douta(w_n9671_0[0]),.doutb(w_n9671_0[1]),.din(n9671));
	jspl jspl_w_n9673_0(.douta(w_n9673_0[0]),.doutb(w_n9673_0[1]),.din(n9673));
	jspl jspl_w_n9675_0(.douta(w_n9675_0[0]),.doutb(w_n9675_0[1]),.din(n9675));
	jspl jspl_w_n9678_0(.douta(w_n9678_0[0]),.doutb(w_n9678_0[1]),.din(n9678));
	jspl jspl_w_n9684_0(.douta(w_n9684_0[0]),.doutb(w_n9684_0[1]),.din(n9684));
	jspl jspl_w_n9686_0(.douta(w_n9686_0[0]),.doutb(w_n9686_0[1]),.din(n9686));
	jspl3 jspl3_w_n9687_0(.douta(w_n9687_0[0]),.doutb(w_n9687_0[1]),.doutc(w_n9687_0[2]),.din(n9687));
	jspl jspl_w_n9691_0(.douta(w_n9691_0[0]),.doutb(w_n9691_0[1]),.din(n9691));
	jspl jspl_w_n9692_0(.douta(w_n9692_0[0]),.doutb(w_n9692_0[1]),.din(n9692));
	jspl3 jspl3_w_n9693_0(.douta(w_n9693_0[0]),.doutb(w_n9693_0[1]),.doutc(w_n9693_0[2]),.din(n9693));
	jspl jspl_w_n9695_0(.douta(w_n9695_0[0]),.doutb(w_n9695_0[1]),.din(n9695));
	jspl jspl_w_n9700_0(.douta(w_n9700_0[0]),.doutb(w_n9700_0[1]),.din(n9700));
	jspl jspl_w_n9702_0(.douta(w_n9702_0[0]),.doutb(w_n9702_0[1]),.din(n9702));
	jspl jspl_w_n9703_0(.douta(w_n9703_0[0]),.doutb(w_n9703_0[1]),.din(n9703));
	jspl3 jspl3_w_n9704_0(.douta(w_n9704_0[0]),.doutb(w_n9704_0[1]),.doutc(w_n9704_0[2]),.din(n9704));
	jspl jspl_w_n9705_0(.douta(w_n9705_0[0]),.doutb(w_n9705_0[1]),.din(n9705));
	jspl jspl_w_n9709_0(.douta(w_n9709_0[0]),.doutb(w_n9709_0[1]),.din(n9709));
	jspl jspl_w_n9715_0(.douta(w_n9715_0[0]),.doutb(w_n9715_0[1]),.din(n9715));
	jspl jspl_w_n9716_0(.douta(w_n9716_0[0]),.doutb(w_n9716_0[1]),.din(n9716));
	jspl jspl_w_n9718_0(.douta(w_n9718_0[0]),.doutb(w_n9718_0[1]),.din(n9718));
	jspl jspl_w_n9720_0(.douta(w_n9720_0[0]),.doutb(w_n9720_0[1]),.din(n9720));
	jspl jspl_w_n9723_0(.douta(w_n9723_0[0]),.doutb(w_n9723_0[1]),.din(n9723));
	jspl jspl_w_n9729_0(.douta(w_n9729_0[0]),.doutb(w_n9729_0[1]),.din(n9729));
	jspl jspl_w_n9731_0(.douta(w_n9731_0[0]),.doutb(w_n9731_0[1]),.din(n9731));
	jspl3 jspl3_w_n9732_0(.douta(w_n9732_0[0]),.doutb(w_n9732_0[1]),.doutc(w_n9732_0[2]),.din(n9732));
	jspl jspl_w_n9736_0(.douta(w_n9736_0[0]),.doutb(w_n9736_0[1]),.din(n9736));
	jspl jspl_w_n9737_0(.douta(w_n9737_0[0]),.doutb(w_n9737_0[1]),.din(n9737));
	jspl3 jspl3_w_n9738_0(.douta(w_n9738_0[0]),.doutb(w_n9738_0[1]),.doutc(w_n9738_0[2]),.din(n9738));
	jspl jspl_w_n9740_0(.douta(w_n9740_0[0]),.doutb(w_n9740_0[1]),.din(n9740));
	jspl jspl_w_n9745_0(.douta(w_n9745_0[0]),.doutb(w_n9745_0[1]),.din(n9745));
	jspl jspl_w_n9747_0(.douta(w_n9747_0[0]),.doutb(w_n9747_0[1]),.din(n9747));
	jspl jspl_w_n9748_0(.douta(w_n9748_0[0]),.doutb(w_n9748_0[1]),.din(n9748));
	jspl3 jspl3_w_n9749_0(.douta(w_n9749_0[0]),.doutb(w_n9749_0[1]),.doutc(w_n9749_0[2]),.din(n9749));
	jspl3 jspl3_w_n9749_1(.douta(w_n9749_1[0]),.doutb(w_n9749_1[1]),.doutc(w_n9749_1[2]),.din(w_n9749_0[0]));
	jspl jspl_w_n9752_0(.douta(w_n9752_0[0]),.doutb(w_n9752_0[1]),.din(n9752));
	jspl3 jspl3_w_n9753_0(.douta(w_n9753_0[0]),.doutb(w_n9753_0[1]),.doutc(w_n9753_0[2]),.din(n9753));
	jspl jspl_w_n9754_0(.douta(w_n9754_0[0]),.doutb(w_n9754_0[1]),.din(n9754));
	jspl jspl_w_n9755_0(.douta(w_n9755_0[0]),.doutb(w_n9755_0[1]),.din(n9755));
	jspl jspl_w_n9761_0(.douta(w_n9761_0[0]),.doutb(w_n9761_0[1]),.din(n9761));
	jspl3 jspl3_w_n9762_0(.douta(w_n9762_0[0]),.doutb(w_n9762_0[1]),.doutc(w_n9762_0[2]),.din(n9762));
	jspl jspl_w_n9763_0(.douta(w_n9763_0[0]),.doutb(w_n9763_0[1]),.din(n9763));
	jspl jspl_w_n9768_0(.douta(w_n9768_0[0]),.doutb(w_n9768_0[1]),.din(n9768));
	jspl3 jspl3_w_n9769_0(.douta(w_n9769_0[0]),.doutb(w_n9769_0[1]),.doutc(w_n9769_0[2]),.din(n9769));
	jspl3 jspl3_w_n9769_1(.douta(w_n9769_1[0]),.doutb(w_n9769_1[1]),.doutc(w_n9769_1[2]),.din(w_n9769_0[0]));
	jspl3 jspl3_w_n9769_2(.douta(w_n9769_2[0]),.doutb(w_n9769_2[1]),.doutc(w_n9769_2[2]),.din(w_n9769_0[1]));
	jspl3 jspl3_w_n9769_3(.douta(w_n9769_3[0]),.doutb(w_n9769_3[1]),.doutc(w_n9769_3[2]),.din(w_n9769_0[2]));
	jspl3 jspl3_w_n9769_4(.douta(w_n9769_4[0]),.doutb(w_n9769_4[1]),.doutc(w_n9769_4[2]),.din(w_n9769_1[0]));
	jspl3 jspl3_w_n9769_5(.douta(w_n9769_5[0]),.doutb(w_n9769_5[1]),.doutc(w_n9769_5[2]),.din(w_n9769_1[1]));
	jspl3 jspl3_w_n9769_6(.douta(w_n9769_6[0]),.doutb(w_n9769_6[1]),.doutc(w_n9769_6[2]),.din(w_n9769_1[2]));
	jspl3 jspl3_w_n9769_7(.douta(w_n9769_7[0]),.doutb(w_n9769_7[1]),.doutc(w_n9769_7[2]),.din(w_n9769_2[0]));
	jspl3 jspl3_w_n9769_8(.douta(w_n9769_8[0]),.doutb(w_n9769_8[1]),.doutc(w_n9769_8[2]),.din(w_n9769_2[1]));
	jspl3 jspl3_w_n9769_9(.douta(w_n9769_9[0]),.doutb(w_n9769_9[1]),.doutc(w_n9769_9[2]),.din(w_n9769_2[2]));
	jspl3 jspl3_w_n9769_10(.douta(w_n9769_10[0]),.doutb(w_n9769_10[1]),.doutc(w_n9769_10[2]),.din(w_n9769_3[0]));
	jspl3 jspl3_w_n9769_11(.douta(w_n9769_11[0]),.doutb(w_n9769_11[1]),.doutc(w_n9769_11[2]),.din(w_n9769_3[1]));
	jspl3 jspl3_w_n9769_12(.douta(w_n9769_12[0]),.doutb(w_n9769_12[1]),.doutc(w_n9769_12[2]),.din(w_n9769_3[2]));
	jspl3 jspl3_w_n9769_13(.douta(w_n9769_13[0]),.doutb(w_n9769_13[1]),.doutc(w_n9769_13[2]),.din(w_n9769_4[0]));
	jspl jspl_w_n9769_14(.douta(w_n9769_14[0]),.doutb(w_n9769_14[1]),.din(w_n9769_4[1]));
	jspl3 jspl3_w_n9774_0(.douta(w_n9774_0[0]),.doutb(w_n9774_0[1]),.doutc(w_n9774_0[2]),.din(n9774));
	jspl3 jspl3_w_n9774_1(.douta(w_n9774_1[0]),.doutb(w_n9774_1[1]),.doutc(w_n9774_1[2]),.din(w_n9774_0[0]));
	jspl3 jspl3_w_n9774_2(.douta(w_n9774_2[0]),.doutb(w_n9774_2[1]),.doutc(w_n9774_2[2]),.din(w_n9774_0[1]));
	jspl3 jspl3_w_n9774_3(.douta(w_n9774_3[0]),.doutb(w_n9774_3[1]),.doutc(w_n9774_3[2]),.din(w_n9774_0[2]));
	jspl3 jspl3_w_n9774_4(.douta(w_n9774_4[0]),.doutb(w_n9774_4[1]),.doutc(w_n9774_4[2]),.din(w_n9774_1[0]));
	jspl3 jspl3_w_n9774_5(.douta(w_n9774_5[0]),.doutb(w_n9774_5[1]),.doutc(w_n9774_5[2]),.din(w_n9774_1[1]));
	jspl3 jspl3_w_n9774_6(.douta(w_n9774_6[0]),.doutb(w_n9774_6[1]),.doutc(w_n9774_6[2]),.din(w_n9774_1[2]));
	jspl3 jspl3_w_n9774_7(.douta(w_n9774_7[0]),.doutb(w_n9774_7[1]),.doutc(w_n9774_7[2]),.din(w_n9774_2[0]));
	jspl3 jspl3_w_n9774_8(.douta(w_n9774_8[0]),.doutb(w_n9774_8[1]),.doutc(w_n9774_8[2]),.din(w_n9774_2[1]));
	jspl3 jspl3_w_n9774_9(.douta(w_n9774_9[0]),.doutb(w_n9774_9[1]),.doutc(w_n9774_9[2]),.din(w_n9774_2[2]));
	jspl3 jspl3_w_n9774_10(.douta(w_n9774_10[0]),.doutb(w_n9774_10[1]),.doutc(w_n9774_10[2]),.din(w_n9774_3[0]));
	jspl3 jspl3_w_n9774_11(.douta(w_n9774_11[0]),.doutb(w_n9774_11[1]),.doutc(w_n9774_11[2]),.din(w_n9774_3[1]));
	jspl3 jspl3_w_n9774_12(.douta(w_n9774_12[0]),.doutb(w_n9774_12[1]),.doutc(w_n9774_12[2]),.din(w_n9774_3[2]));
	jspl3 jspl3_w_n9774_13(.douta(w_n9774_13[0]),.doutb(w_n9774_13[1]),.doutc(w_n9774_13[2]),.din(w_n9774_4[0]));
	jspl3 jspl3_w_n9774_14(.douta(w_n9774_14[0]),.doutb(w_n9774_14[1]),.doutc(w_n9774_14[2]),.din(w_n9774_4[1]));
	jspl3 jspl3_w_n9774_15(.douta(w_n9774_15[0]),.doutb(w_n9774_15[1]),.doutc(w_n9774_15[2]),.din(w_n9774_4[2]));
	jspl3 jspl3_w_n9774_16(.douta(w_n9774_16[0]),.doutb(w_n9774_16[1]),.doutc(w_n9774_16[2]),.din(w_n9774_5[0]));
	jspl3 jspl3_w_n9774_17(.douta(w_n9774_17[0]),.doutb(w_n9774_17[1]),.doutc(w_n9774_17[2]),.din(w_n9774_5[1]));
	jspl3 jspl3_w_n9774_18(.douta(w_n9774_18[0]),.doutb(w_n9774_18[1]),.doutc(w_n9774_18[2]),.din(w_n9774_5[2]));
	jspl3 jspl3_w_n9774_19(.douta(w_n9774_19[0]),.doutb(w_n9774_19[1]),.doutc(w_n9774_19[2]),.din(w_n9774_6[0]));
	jspl3 jspl3_w_n9774_20(.douta(w_n9774_20[0]),.doutb(w_n9774_20[1]),.doutc(w_n9774_20[2]),.din(w_n9774_6[1]));
	jspl3 jspl3_w_n9774_21(.douta(w_n9774_21[0]),.doutb(w_n9774_21[1]),.doutc(w_n9774_21[2]),.din(w_n9774_6[2]));
	jspl3 jspl3_w_n9774_22(.douta(w_n9774_22[0]),.doutb(w_n9774_22[1]),.doutc(w_n9774_22[2]),.din(w_n9774_7[0]));
	jspl3 jspl3_w_n9774_23(.douta(w_n9774_23[0]),.doutb(w_n9774_23[1]),.doutc(w_n9774_23[2]),.din(w_n9774_7[1]));
	jspl3 jspl3_w_n9774_24(.douta(w_n9774_24[0]),.doutb(w_n9774_24[1]),.doutc(w_n9774_24[2]),.din(w_n9774_7[2]));
	jspl3 jspl3_w_n9774_25(.douta(w_n9774_25[0]),.doutb(w_n9774_25[1]),.doutc(w_n9774_25[2]),.din(w_n9774_8[0]));
	jspl jspl_w_n9778_0(.douta(w_n9778_0[0]),.doutb(w_n9778_0[1]),.din(n9778));
	jspl3 jspl3_w_n9780_0(.douta(w_n9780_0[0]),.doutb(w_n9780_0[1]),.doutc(w_n9780_0[2]),.din(n9780));
	jspl jspl_w_n9780_1(.douta(w_n9780_1[0]),.doutb(w_n9780_1[1]),.din(w_n9780_0[0]));
	jspl3 jspl3_w_n9781_0(.douta(w_n9781_0[0]),.doutb(w_n9781_0[1]),.doutc(w_n9781_0[2]),.din(n9781));
	jspl3 jspl3_w_n9785_0(.douta(w_n9785_0[0]),.doutb(w_n9785_0[1]),.doutc(w_n9785_0[2]),.din(n9785));
	jspl jspl_w_n9786_0(.douta(w_n9786_0[0]),.doutb(w_n9786_0[1]),.din(n9786));
	jspl jspl_w_n9787_0(.douta(w_n9787_0[0]),.doutb(w_n9787_0[1]),.din(n9787));
	jspl jspl_w_n9788_0(.douta(w_n9788_0[0]),.doutb(w_n9788_0[1]),.din(n9788));
	jspl jspl_w_n9790_0(.douta(w_n9790_0[0]),.doutb(w_n9790_0[1]),.din(n9790));
	jspl jspl_w_n9792_0(.douta(w_n9792_0[0]),.doutb(w_n9792_0[1]),.din(n9792));
	jspl jspl_w_n9794_0(.douta(w_n9794_0[0]),.doutb(w_n9794_0[1]),.din(n9794));
	jspl jspl_w_n9797_0(.douta(w_n9797_0[0]),.doutb(w_n9797_0[1]),.din(n9797));
	jspl jspl_w_n9802_0(.douta(w_n9802_0[0]),.doutb(w_n9802_0[1]),.din(n9802));
	jspl3 jspl3_w_n9804_0(.douta(w_n9804_0[0]),.doutb(w_n9804_0[1]),.doutc(w_n9804_0[2]),.din(n9804));
	jspl jspl_w_n9805_0(.douta(w_n9805_0[0]),.doutb(w_n9805_0[1]),.din(n9805));
	jspl jspl_w_n9809_0(.douta(w_n9809_0[0]),.doutb(w_n9809_0[1]),.din(n9809));
	jspl jspl_w_n9810_0(.douta(w_n9810_0[0]),.doutb(w_n9810_0[1]),.din(n9810));
	jspl jspl_w_n9812_0(.douta(w_n9812_0[0]),.doutb(w_n9812_0[1]),.din(n9812));
	jspl jspl_w_n9816_0(.douta(w_n9816_0[0]),.doutb(w_n9816_0[1]),.din(n9816));
	jspl jspl_w_n9818_0(.douta(w_n9818_0[0]),.doutb(w_n9818_0[1]),.din(n9818));
	jspl jspl_w_n9819_0(.douta(w_n9819_0[0]),.doutb(w_n9819_0[1]),.din(n9819));
	jspl3 jspl3_w_n9820_0(.douta(w_n9820_0[0]),.doutb(w_n9820_0[1]),.doutc(w_n9820_0[2]),.din(n9820));
	jspl jspl_w_n9821_0(.douta(w_n9821_0[0]),.doutb(w_n9821_0[1]),.din(n9821));
	jspl jspl_w_n9825_0(.douta(w_n9825_0[0]),.doutb(w_n9825_0[1]),.din(n9825));
	jspl jspl_w_n9827_0(.douta(w_n9827_0[0]),.doutb(w_n9827_0[1]),.din(n9827));
	jspl jspl_w_n9829_0(.douta(w_n9829_0[0]),.doutb(w_n9829_0[1]),.din(n9829));
	jspl jspl_w_n9831_0(.douta(w_n9831_0[0]),.doutb(w_n9831_0[1]),.din(n9831));
	jspl jspl_w_n9834_0(.douta(w_n9834_0[0]),.doutb(w_n9834_0[1]),.din(n9834));
	jspl jspl_w_n9840_0(.douta(w_n9840_0[0]),.doutb(w_n9840_0[1]),.din(n9840));
	jspl3 jspl3_w_n9842_0(.douta(w_n9842_0[0]),.doutb(w_n9842_0[1]),.doutc(w_n9842_0[2]),.din(n9842));
	jspl jspl_w_n9843_0(.douta(w_n9843_0[0]),.doutb(w_n9843_0[1]),.din(n9843));
	jspl jspl_w_n9848_0(.douta(w_n9848_0[0]),.doutb(w_n9848_0[1]),.din(n9848));
	jspl jspl_w_n9850_0(.douta(w_n9850_0[0]),.doutb(w_n9850_0[1]),.din(n9850));
	jspl jspl_w_n9852_0(.douta(w_n9852_0[0]),.doutb(w_n9852_0[1]),.din(n9852));
	jspl jspl_w_n9856_0(.douta(w_n9856_0[0]),.doutb(w_n9856_0[1]),.din(n9856));
	jspl jspl_w_n9858_0(.douta(w_n9858_0[0]),.doutb(w_n9858_0[1]),.din(n9858));
	jspl jspl_w_n9859_0(.douta(w_n9859_0[0]),.doutb(w_n9859_0[1]),.din(n9859));
	jspl3 jspl3_w_n9860_0(.douta(w_n9860_0[0]),.doutb(w_n9860_0[1]),.doutc(w_n9860_0[2]),.din(n9860));
	jspl jspl_w_n9861_0(.douta(w_n9861_0[0]),.doutb(w_n9861_0[1]),.din(n9861));
	jspl jspl_w_n9867_0(.douta(w_n9867_0[0]),.doutb(w_n9867_0[1]),.din(n9867));
	jspl jspl_w_n9868_0(.douta(w_n9868_0[0]),.doutb(w_n9868_0[1]),.din(n9868));
	jspl jspl_w_n9870_0(.douta(w_n9870_0[0]),.doutb(w_n9870_0[1]),.din(n9870));
	jspl jspl_w_n9872_0(.douta(w_n9872_0[0]),.doutb(w_n9872_0[1]),.din(n9872));
	jspl jspl_w_n9874_0(.douta(w_n9874_0[0]),.doutb(w_n9874_0[1]),.din(n9874));
	jspl jspl_w_n9880_0(.douta(w_n9880_0[0]),.doutb(w_n9880_0[1]),.din(n9880));
	jspl jspl_w_n9882_0(.douta(w_n9882_0[0]),.doutb(w_n9882_0[1]),.din(n9882));
	jspl3 jspl3_w_n9883_0(.douta(w_n9883_0[0]),.doutb(w_n9883_0[1]),.doutc(w_n9883_0[2]),.din(n9883));
	jspl jspl_w_n9886_0(.douta(w_n9886_0[0]),.doutb(w_n9886_0[1]),.din(n9886));
	jspl jspl_w_n9887_0(.douta(w_n9887_0[0]),.doutb(w_n9887_0[1]),.din(n9887));
	jspl3 jspl3_w_n9888_0(.douta(w_n9888_0[0]),.doutb(w_n9888_0[1]),.doutc(w_n9888_0[2]),.din(n9888));
	jspl jspl_w_n9890_0(.douta(w_n9890_0[0]),.doutb(w_n9890_0[1]),.din(n9890));
	jspl jspl_w_n9894_0(.douta(w_n9894_0[0]),.doutb(w_n9894_0[1]),.din(n9894));
	jspl jspl_w_n9896_0(.douta(w_n9896_0[0]),.doutb(w_n9896_0[1]),.din(n9896));
	jspl jspl_w_n9897_0(.douta(w_n9897_0[0]),.doutb(w_n9897_0[1]),.din(n9897));
	jspl3 jspl3_w_n9898_0(.douta(w_n9898_0[0]),.doutb(w_n9898_0[1]),.doutc(w_n9898_0[2]),.din(n9898));
	jspl jspl_w_n9899_0(.douta(w_n9899_0[0]),.doutb(w_n9899_0[1]),.din(n9899));
	jspl jspl_w_n9902_0(.douta(w_n9902_0[0]),.doutb(w_n9902_0[1]),.din(n9902));
	jspl jspl_w_n9908_0(.douta(w_n9908_0[0]),.doutb(w_n9908_0[1]),.din(n9908));
	jspl jspl_w_n9909_0(.douta(w_n9909_0[0]),.doutb(w_n9909_0[1]),.din(n9909));
	jspl jspl_w_n9911_0(.douta(w_n9911_0[0]),.doutb(w_n9911_0[1]),.din(n9911));
	jspl jspl_w_n9913_0(.douta(w_n9913_0[0]),.doutb(w_n9913_0[1]),.din(n9913));
	jspl jspl_w_n9915_0(.douta(w_n9915_0[0]),.doutb(w_n9915_0[1]),.din(n9915));
	jspl jspl_w_n9921_0(.douta(w_n9921_0[0]),.doutb(w_n9921_0[1]),.din(n9921));
	jspl jspl_w_n9923_0(.douta(w_n9923_0[0]),.doutb(w_n9923_0[1]),.din(n9923));
	jspl3 jspl3_w_n9924_0(.douta(w_n9924_0[0]),.doutb(w_n9924_0[1]),.doutc(w_n9924_0[2]),.din(n9924));
	jspl jspl_w_n9927_0(.douta(w_n9927_0[0]),.doutb(w_n9927_0[1]),.din(n9927));
	jspl jspl_w_n9928_0(.douta(w_n9928_0[0]),.doutb(w_n9928_0[1]),.din(n9928));
	jspl3 jspl3_w_n9929_0(.douta(w_n9929_0[0]),.doutb(w_n9929_0[1]),.doutc(w_n9929_0[2]),.din(n9929));
	jspl jspl_w_n9931_0(.douta(w_n9931_0[0]),.doutb(w_n9931_0[1]),.din(n9931));
	jspl jspl_w_n9935_0(.douta(w_n9935_0[0]),.doutb(w_n9935_0[1]),.din(n9935));
	jspl jspl_w_n9937_0(.douta(w_n9937_0[0]),.doutb(w_n9937_0[1]),.din(n9937));
	jspl jspl_w_n9938_0(.douta(w_n9938_0[0]),.doutb(w_n9938_0[1]),.din(n9938));
	jspl3 jspl3_w_n9939_0(.douta(w_n9939_0[0]),.doutb(w_n9939_0[1]),.doutc(w_n9939_0[2]),.din(n9939));
	jspl jspl_w_n9940_0(.douta(w_n9940_0[0]),.doutb(w_n9940_0[1]),.din(n9940));
	jspl jspl_w_n9943_0(.douta(w_n9943_0[0]),.doutb(w_n9943_0[1]),.din(n9943));
	jspl jspl_w_n9949_0(.douta(w_n9949_0[0]),.doutb(w_n9949_0[1]),.din(n9949));
	jspl jspl_w_n9950_0(.douta(w_n9950_0[0]),.doutb(w_n9950_0[1]),.din(n9950));
	jspl jspl_w_n9952_0(.douta(w_n9952_0[0]),.doutb(w_n9952_0[1]),.din(n9952));
	jspl jspl_w_n9954_0(.douta(w_n9954_0[0]),.doutb(w_n9954_0[1]),.din(n9954));
	jspl jspl_w_n9956_0(.douta(w_n9956_0[0]),.doutb(w_n9956_0[1]),.din(n9956));
	jspl jspl_w_n9962_0(.douta(w_n9962_0[0]),.doutb(w_n9962_0[1]),.din(n9962));
	jspl jspl_w_n9964_0(.douta(w_n9964_0[0]),.doutb(w_n9964_0[1]),.din(n9964));
	jspl3 jspl3_w_n9965_0(.douta(w_n9965_0[0]),.doutb(w_n9965_0[1]),.doutc(w_n9965_0[2]),.din(n9965));
	jspl jspl_w_n9968_0(.douta(w_n9968_0[0]),.doutb(w_n9968_0[1]),.din(n9968));
	jspl jspl_w_n9969_0(.douta(w_n9969_0[0]),.doutb(w_n9969_0[1]),.din(n9969));
	jspl3 jspl3_w_n9970_0(.douta(w_n9970_0[0]),.doutb(w_n9970_0[1]),.doutc(w_n9970_0[2]),.din(n9970));
	jspl jspl_w_n9972_0(.douta(w_n9972_0[0]),.doutb(w_n9972_0[1]),.din(n9972));
	jspl jspl_w_n9974_0(.douta(w_n9974_0[0]),.doutb(w_n9974_0[1]),.din(n9974));
	jspl jspl_w_n9976_0(.douta(w_n9976_0[0]),.doutb(w_n9976_0[1]),.din(n9976));
	jspl jspl_w_n9982_0(.douta(w_n9982_0[0]),.doutb(w_n9982_0[1]),.din(n9982));
	jspl3 jspl3_w_n9984_0(.douta(w_n9984_0[0]),.doutb(w_n9984_0[1]),.doutc(w_n9984_0[2]),.din(n9984));
	jspl jspl_w_n9985_0(.douta(w_n9985_0[0]),.doutb(w_n9985_0[1]),.din(n9985));
	jspl jspl_w_n9987_0(.douta(w_n9987_0[0]),.doutb(w_n9987_0[1]),.din(n9987));
	jspl jspl_w_n9989_0(.douta(w_n9989_0[0]),.doutb(w_n9989_0[1]),.din(n9989));
	jspl jspl_w_n9993_0(.douta(w_n9993_0[0]),.doutb(w_n9993_0[1]),.din(n9993));
	jspl jspl_w_n9995_0(.douta(w_n9995_0[0]),.doutb(w_n9995_0[1]),.din(n9995));
	jspl jspl_w_n9996_0(.douta(w_n9996_0[0]),.doutb(w_n9996_0[1]),.din(n9996));
	jspl jspl_w_n9997_0(.douta(w_n9997_0[0]),.doutb(w_n9997_0[1]),.din(n9997));
	jspl3 jspl3_w_n9998_0(.douta(w_n9998_0[0]),.doutb(w_n9998_0[1]),.doutc(w_n9998_0[2]),.din(n9998));
	jspl jspl_w_n10001_0(.douta(w_n10001_0[0]),.doutb(w_n10001_0[1]),.din(n10001));
	jspl jspl_w_n10002_0(.douta(w_n10002_0[0]),.doutb(w_n10002_0[1]),.din(n10002));
	jspl3 jspl3_w_n10003_0(.douta(w_n10003_0[0]),.doutb(w_n10003_0[1]),.doutc(w_n10003_0[2]),.din(n10003));
	jspl jspl_w_n10005_0(.douta(w_n10005_0[0]),.doutb(w_n10005_0[1]),.din(n10005));
	jspl jspl_w_n10009_0(.douta(w_n10009_0[0]),.doutb(w_n10009_0[1]),.din(n10009));
	jspl jspl_w_n10011_0(.douta(w_n10011_0[0]),.doutb(w_n10011_0[1]),.din(n10011));
	jspl jspl_w_n10012_0(.douta(w_n10012_0[0]),.doutb(w_n10012_0[1]),.din(n10012));
	jspl3 jspl3_w_n10013_0(.douta(w_n10013_0[0]),.doutb(w_n10013_0[1]),.doutc(w_n10013_0[2]),.din(n10013));
	jspl jspl_w_n10014_0(.douta(w_n10014_0[0]),.doutb(w_n10014_0[1]),.din(n10014));
	jspl jspl_w_n10017_0(.douta(w_n10017_0[0]),.doutb(w_n10017_0[1]),.din(n10017));
	jspl jspl_w_n10023_0(.douta(w_n10023_0[0]),.doutb(w_n10023_0[1]),.din(n10023));
	jspl jspl_w_n10024_0(.douta(w_n10024_0[0]),.doutb(w_n10024_0[1]),.din(n10024));
	jspl jspl_w_n10026_0(.douta(w_n10026_0[0]),.doutb(w_n10026_0[1]),.din(n10026));
	jspl jspl_w_n10028_0(.douta(w_n10028_0[0]),.doutb(w_n10028_0[1]),.din(n10028));
	jspl jspl_w_n10030_0(.douta(w_n10030_0[0]),.doutb(w_n10030_0[1]),.din(n10030));
	jspl jspl_w_n10036_0(.douta(w_n10036_0[0]),.doutb(w_n10036_0[1]),.din(n10036));
	jspl jspl_w_n10038_0(.douta(w_n10038_0[0]),.doutb(w_n10038_0[1]),.din(n10038));
	jspl3 jspl3_w_n10039_0(.douta(w_n10039_0[0]),.doutb(w_n10039_0[1]),.doutc(w_n10039_0[2]),.din(n10039));
	jspl jspl_w_n10042_0(.douta(w_n10042_0[0]),.doutb(w_n10042_0[1]),.din(n10042));
	jspl jspl_w_n10043_0(.douta(w_n10043_0[0]),.doutb(w_n10043_0[1]),.din(n10043));
	jspl3 jspl3_w_n10044_0(.douta(w_n10044_0[0]),.doutb(w_n10044_0[1]),.doutc(w_n10044_0[2]),.din(n10044));
	jspl jspl_w_n10046_0(.douta(w_n10046_0[0]),.doutb(w_n10046_0[1]),.din(n10046));
	jspl jspl_w_n10050_0(.douta(w_n10050_0[0]),.doutb(w_n10050_0[1]),.din(n10050));
	jspl jspl_w_n10052_0(.douta(w_n10052_0[0]),.doutb(w_n10052_0[1]),.din(n10052));
	jspl jspl_w_n10053_0(.douta(w_n10053_0[0]),.doutb(w_n10053_0[1]),.din(n10053));
	jspl3 jspl3_w_n10054_0(.douta(w_n10054_0[0]),.doutb(w_n10054_0[1]),.doutc(w_n10054_0[2]),.din(n10054));
	jspl jspl_w_n10055_0(.douta(w_n10055_0[0]),.doutb(w_n10055_0[1]),.din(n10055));
	jspl jspl_w_n10058_0(.douta(w_n10058_0[0]),.doutb(w_n10058_0[1]),.din(n10058));
	jspl jspl_w_n10064_0(.douta(w_n10064_0[0]),.doutb(w_n10064_0[1]),.din(n10064));
	jspl jspl_w_n10065_0(.douta(w_n10065_0[0]),.doutb(w_n10065_0[1]),.din(n10065));
	jspl jspl_w_n10067_0(.douta(w_n10067_0[0]),.doutb(w_n10067_0[1]),.din(n10067));
	jspl jspl_w_n10069_0(.douta(w_n10069_0[0]),.doutb(w_n10069_0[1]),.din(n10069));
	jspl jspl_w_n10071_0(.douta(w_n10071_0[0]),.doutb(w_n10071_0[1]),.din(n10071));
	jspl jspl_w_n10077_0(.douta(w_n10077_0[0]),.doutb(w_n10077_0[1]),.din(n10077));
	jspl jspl_w_n10079_0(.douta(w_n10079_0[0]),.doutb(w_n10079_0[1]),.din(n10079));
	jspl3 jspl3_w_n10080_0(.douta(w_n10080_0[0]),.doutb(w_n10080_0[1]),.doutc(w_n10080_0[2]),.din(n10080));
	jspl jspl_w_n10083_0(.douta(w_n10083_0[0]),.doutb(w_n10083_0[1]),.din(n10083));
	jspl jspl_w_n10084_0(.douta(w_n10084_0[0]),.doutb(w_n10084_0[1]),.din(n10084));
	jspl3 jspl3_w_n10085_0(.douta(w_n10085_0[0]),.doutb(w_n10085_0[1]),.doutc(w_n10085_0[2]),.din(n10085));
	jspl jspl_w_n10087_0(.douta(w_n10087_0[0]),.doutb(w_n10087_0[1]),.din(n10087));
	jspl jspl_w_n10091_0(.douta(w_n10091_0[0]),.doutb(w_n10091_0[1]),.din(n10091));
	jspl jspl_w_n10093_0(.douta(w_n10093_0[0]),.doutb(w_n10093_0[1]),.din(n10093));
	jspl jspl_w_n10094_0(.douta(w_n10094_0[0]),.doutb(w_n10094_0[1]),.din(n10094));
	jspl3 jspl3_w_n10095_0(.douta(w_n10095_0[0]),.doutb(w_n10095_0[1]),.doutc(w_n10095_0[2]),.din(n10095));
	jspl jspl_w_n10096_0(.douta(w_n10096_0[0]),.doutb(w_n10096_0[1]),.din(n10096));
	jspl jspl_w_n10099_0(.douta(w_n10099_0[0]),.doutb(w_n10099_0[1]),.din(n10099));
	jspl jspl_w_n10105_0(.douta(w_n10105_0[0]),.doutb(w_n10105_0[1]),.din(n10105));
	jspl jspl_w_n10106_0(.douta(w_n10106_0[0]),.doutb(w_n10106_0[1]),.din(n10106));
	jspl jspl_w_n10108_0(.douta(w_n10108_0[0]),.doutb(w_n10108_0[1]),.din(n10108));
	jspl jspl_w_n10110_0(.douta(w_n10110_0[0]),.doutb(w_n10110_0[1]),.din(n10110));
	jspl jspl_w_n10112_0(.douta(w_n10112_0[0]),.doutb(w_n10112_0[1]),.din(n10112));
	jspl jspl_w_n10118_0(.douta(w_n10118_0[0]),.doutb(w_n10118_0[1]),.din(n10118));
	jspl jspl_w_n10120_0(.douta(w_n10120_0[0]),.doutb(w_n10120_0[1]),.din(n10120));
	jspl3 jspl3_w_n10121_0(.douta(w_n10121_0[0]),.doutb(w_n10121_0[1]),.doutc(w_n10121_0[2]),.din(n10121));
	jspl jspl_w_n10124_0(.douta(w_n10124_0[0]),.doutb(w_n10124_0[1]),.din(n10124));
	jspl jspl_w_n10125_0(.douta(w_n10125_0[0]),.doutb(w_n10125_0[1]),.din(n10125));
	jspl3 jspl3_w_n10126_0(.douta(w_n10126_0[0]),.doutb(w_n10126_0[1]),.doutc(w_n10126_0[2]),.din(n10126));
	jspl jspl_w_n10128_0(.douta(w_n10128_0[0]),.doutb(w_n10128_0[1]),.din(n10128));
	jspl jspl_w_n10132_0(.douta(w_n10132_0[0]),.doutb(w_n10132_0[1]),.din(n10132));
	jspl jspl_w_n10134_0(.douta(w_n10134_0[0]),.doutb(w_n10134_0[1]),.din(n10134));
	jspl jspl_w_n10135_0(.douta(w_n10135_0[0]),.doutb(w_n10135_0[1]),.din(n10135));
	jspl3 jspl3_w_n10136_0(.douta(w_n10136_0[0]),.doutb(w_n10136_0[1]),.doutc(w_n10136_0[2]),.din(n10136));
	jspl jspl_w_n10137_0(.douta(w_n10137_0[0]),.doutb(w_n10137_0[1]),.din(n10137));
	jspl jspl_w_n10140_0(.douta(w_n10140_0[0]),.doutb(w_n10140_0[1]),.din(n10140));
	jspl jspl_w_n10146_0(.douta(w_n10146_0[0]),.doutb(w_n10146_0[1]),.din(n10146));
	jspl jspl_w_n10147_0(.douta(w_n10147_0[0]),.doutb(w_n10147_0[1]),.din(n10147));
	jspl jspl_w_n10149_0(.douta(w_n10149_0[0]),.doutb(w_n10149_0[1]),.din(n10149));
	jspl jspl_w_n10151_0(.douta(w_n10151_0[0]),.doutb(w_n10151_0[1]),.din(n10151));
	jspl jspl_w_n10153_0(.douta(w_n10153_0[0]),.doutb(w_n10153_0[1]),.din(n10153));
	jspl jspl_w_n10159_0(.douta(w_n10159_0[0]),.doutb(w_n10159_0[1]),.din(n10159));
	jspl jspl_w_n10161_0(.douta(w_n10161_0[0]),.doutb(w_n10161_0[1]),.din(n10161));
	jspl3 jspl3_w_n10162_0(.douta(w_n10162_0[0]),.doutb(w_n10162_0[1]),.doutc(w_n10162_0[2]),.din(n10162));
	jspl jspl_w_n10165_0(.douta(w_n10165_0[0]),.doutb(w_n10165_0[1]),.din(n10165));
	jspl jspl_w_n10166_0(.douta(w_n10166_0[0]),.doutb(w_n10166_0[1]),.din(n10166));
	jspl3 jspl3_w_n10167_0(.douta(w_n10167_0[0]),.doutb(w_n10167_0[1]),.doutc(w_n10167_0[2]),.din(n10167));
	jspl jspl_w_n10169_0(.douta(w_n10169_0[0]),.doutb(w_n10169_0[1]),.din(n10169));
	jspl jspl_w_n10173_0(.douta(w_n10173_0[0]),.doutb(w_n10173_0[1]),.din(n10173));
	jspl jspl_w_n10175_0(.douta(w_n10175_0[0]),.doutb(w_n10175_0[1]),.din(n10175));
	jspl jspl_w_n10176_0(.douta(w_n10176_0[0]),.doutb(w_n10176_0[1]),.din(n10176));
	jspl3 jspl3_w_n10177_0(.douta(w_n10177_0[0]),.doutb(w_n10177_0[1]),.doutc(w_n10177_0[2]),.din(n10177));
	jspl jspl_w_n10181_0(.douta(w_n10181_0[0]),.doutb(w_n10181_0[1]),.din(n10181));
	jspl jspl_w_n10187_0(.douta(w_n10187_0[0]),.doutb(w_n10187_0[1]),.din(n10187));
	jspl3 jspl3_w_n10189_0(.douta(w_n10189_0[0]),.doutb(w_n10189_0[1]),.doutc(w_n10189_0[2]),.din(n10189));
	jspl jspl_w_n10191_0(.douta(w_n10191_0[0]),.doutb(w_n10191_0[1]),.din(n10191));
	jspl3 jspl3_w_n10196_0(.douta(w_n10196_0[0]),.doutb(w_n10196_0[1]),.doutc(w_n10196_0[2]),.din(n10196));
	jspl jspl_w_n10197_0(.douta(w_n10197_0[0]),.doutb(w_n10197_0[1]),.din(n10197));
	jspl jspl_w_n10198_0(.douta(w_n10198_0[0]),.doutb(w_n10198_0[1]),.din(n10198));
	jspl jspl_w_n10203_0(.douta(w_n10203_0[0]),.doutb(w_n10203_0[1]),.din(n10203));
	jspl3 jspl3_w_n10204_0(.douta(w_n10204_0[0]),.doutb(w_n10204_0[1]),.doutc(w_n10204_0[2]),.din(n10204));
	jspl jspl_w_n10209_0(.douta(w_n10209_0[0]),.doutb(w_n10209_0[1]),.din(n10209));
	jspl jspl_w_n10217_0(.douta(w_n10217_0[0]),.doutb(w_n10217_0[1]),.din(n10217));
	jspl3 jspl3_w_n10219_0(.douta(w_n10219_0[0]),.doutb(w_n10219_0[1]),.doutc(w_n10219_0[2]),.din(n10219));
	jspl jspl_w_n10219_1(.douta(w_n10219_1[0]),.doutb(w_n10219_1[1]),.din(w_n10219_0[0]));
	jspl jspl_w_n10220_0(.douta(w_n10220_0[0]),.doutb(w_n10220_0[1]),.din(n10220));
	jspl3 jspl3_w_n10223_0(.douta(w_n10223_0[0]),.doutb(w_n10223_0[1]),.doutc(w_n10223_0[2]),.din(n10223));
	jspl jspl_w_n10224_0(.douta(w_n10224_0[0]),.doutb(w_n10224_0[1]),.din(n10224));
	jspl jspl_w_n10225_0(.douta(w_n10225_0[0]),.doutb(w_n10225_0[1]),.din(n10225));
	jspl jspl_w_n10226_0(.douta(w_n10226_0[0]),.doutb(w_n10226_0[1]),.din(n10226));
	jspl jspl_w_n10228_0(.douta(w_n10228_0[0]),.doutb(w_n10228_0[1]),.din(n10228));
	jspl jspl_w_n10230_0(.douta(w_n10230_0[0]),.doutb(w_n10230_0[1]),.din(n10230));
	jspl jspl_w_n10232_0(.douta(w_n10232_0[0]),.doutb(w_n10232_0[1]),.din(n10232));
	jspl jspl_w_n10241_0(.douta(w_n10241_0[0]),.doutb(w_n10241_0[1]),.din(n10241));
	jspl3 jspl3_w_n10243_0(.douta(w_n10243_0[0]),.doutb(w_n10243_0[1]),.doutc(w_n10243_0[2]),.din(n10243));
	jspl jspl_w_n10244_0(.douta(w_n10244_0[0]),.doutb(w_n10244_0[1]),.din(n10244));
	jspl jspl_w_n10248_0(.douta(w_n10248_0[0]),.doutb(w_n10248_0[1]),.din(n10248));
	jspl jspl_w_n10250_0(.douta(w_n10250_0[0]),.doutb(w_n10250_0[1]),.din(n10250));
	jspl jspl_w_n10252_0(.douta(w_n10252_0[0]),.doutb(w_n10252_0[1]),.din(n10252));
	jspl jspl_w_n10257_0(.douta(w_n10257_0[0]),.doutb(w_n10257_0[1]),.din(n10257));
	jspl jspl_w_n10259_0(.douta(w_n10259_0[0]),.doutb(w_n10259_0[1]),.din(n10259));
	jspl jspl_w_n10260_0(.douta(w_n10260_0[0]),.doutb(w_n10260_0[1]),.din(n10260));
	jspl3 jspl3_w_n10261_0(.douta(w_n10261_0[0]),.doutb(w_n10261_0[1]),.doutc(w_n10261_0[2]),.din(n10261));
	jspl jspl_w_n10262_0(.douta(w_n10262_0[0]),.doutb(w_n10262_0[1]),.din(n10262));
	jspl jspl_w_n10267_0(.douta(w_n10267_0[0]),.doutb(w_n10267_0[1]),.din(n10267));
	jspl jspl_w_n10268_0(.douta(w_n10268_0[0]),.doutb(w_n10268_0[1]),.din(n10268));
	jspl jspl_w_n10270_0(.douta(w_n10270_0[0]),.doutb(w_n10270_0[1]),.din(n10270));
	jspl jspl_w_n10272_0(.douta(w_n10272_0[0]),.doutb(w_n10272_0[1]),.din(n10272));
	jspl jspl_w_n10275_0(.douta(w_n10275_0[0]),.doutb(w_n10275_0[1]),.din(n10275));
	jspl jspl_w_n10281_0(.douta(w_n10281_0[0]),.doutb(w_n10281_0[1]),.din(n10281));
	jspl3 jspl3_w_n10283_0(.douta(w_n10283_0[0]),.doutb(w_n10283_0[1]),.doutc(w_n10283_0[2]),.din(n10283));
	jspl jspl_w_n10284_0(.douta(w_n10284_0[0]),.doutb(w_n10284_0[1]),.din(n10284));
	jspl jspl_w_n10288_0(.douta(w_n10288_0[0]),.doutb(w_n10288_0[1]),.din(n10288));
	jspl jspl_w_n10289_0(.douta(w_n10289_0[0]),.doutb(w_n10289_0[1]),.din(n10289));
	jspl jspl_w_n10291_0(.douta(w_n10291_0[0]),.doutb(w_n10291_0[1]),.din(n10291));
	jspl jspl_w_n10296_0(.douta(w_n10296_0[0]),.doutb(w_n10296_0[1]),.din(n10296));
	jspl jspl_w_n10298_0(.douta(w_n10298_0[0]),.doutb(w_n10298_0[1]),.din(n10298));
	jspl jspl_w_n10299_0(.douta(w_n10299_0[0]),.doutb(w_n10299_0[1]),.din(n10299));
	jspl3 jspl3_w_n10300_0(.douta(w_n10300_0[0]),.doutb(w_n10300_0[1]),.doutc(w_n10300_0[2]),.din(n10300));
	jspl jspl_w_n10301_0(.douta(w_n10301_0[0]),.doutb(w_n10301_0[1]),.din(n10301));
	jspl jspl_w_n10305_0(.douta(w_n10305_0[0]),.doutb(w_n10305_0[1]),.din(n10305));
	jspl jspl_w_n10306_0(.douta(w_n10306_0[0]),.doutb(w_n10306_0[1]),.din(n10306));
	jspl jspl_w_n10308_0(.douta(w_n10308_0[0]),.doutb(w_n10308_0[1]),.din(n10308));
	jspl jspl_w_n10310_0(.douta(w_n10310_0[0]),.doutb(w_n10310_0[1]),.din(n10310));
	jspl jspl_w_n10313_0(.douta(w_n10313_0[0]),.doutb(w_n10313_0[1]),.din(n10313));
	jspl jspl_w_n10319_0(.douta(w_n10319_0[0]),.doutb(w_n10319_0[1]),.din(n10319));
	jspl jspl_w_n10321_0(.douta(w_n10321_0[0]),.doutb(w_n10321_0[1]),.din(n10321));
	jspl3 jspl3_w_n10322_0(.douta(w_n10322_0[0]),.doutb(w_n10322_0[1]),.doutc(w_n10322_0[2]),.din(n10322));
	jspl jspl_w_n10326_0(.douta(w_n10326_0[0]),.doutb(w_n10326_0[1]),.din(n10326));
	jspl jspl_w_n10327_0(.douta(w_n10327_0[0]),.doutb(w_n10327_0[1]),.din(n10327));
	jspl3 jspl3_w_n10328_0(.douta(w_n10328_0[0]),.doutb(w_n10328_0[1]),.doutc(w_n10328_0[2]),.din(n10328));
	jspl jspl_w_n10330_0(.douta(w_n10330_0[0]),.doutb(w_n10330_0[1]),.din(n10330));
	jspl jspl_w_n10335_0(.douta(w_n10335_0[0]),.doutb(w_n10335_0[1]),.din(n10335));
	jspl jspl_w_n10337_0(.douta(w_n10337_0[0]),.doutb(w_n10337_0[1]),.din(n10337));
	jspl jspl_w_n10338_0(.douta(w_n10338_0[0]),.doutb(w_n10338_0[1]),.din(n10338));
	jspl3 jspl3_w_n10339_0(.douta(w_n10339_0[0]),.doutb(w_n10339_0[1]),.doutc(w_n10339_0[2]),.din(n10339));
	jspl jspl_w_n10340_0(.douta(w_n10340_0[0]),.doutb(w_n10340_0[1]),.din(n10340));
	jspl jspl_w_n10344_0(.douta(w_n10344_0[0]),.doutb(w_n10344_0[1]),.din(n10344));
	jspl jspl_w_n10350_0(.douta(w_n10350_0[0]),.doutb(w_n10350_0[1]),.din(n10350));
	jspl jspl_w_n10351_0(.douta(w_n10351_0[0]),.doutb(w_n10351_0[1]),.din(n10351));
	jspl jspl_w_n10353_0(.douta(w_n10353_0[0]),.doutb(w_n10353_0[1]),.din(n10353));
	jspl jspl_w_n10355_0(.douta(w_n10355_0[0]),.doutb(w_n10355_0[1]),.din(n10355));
	jspl jspl_w_n10358_0(.douta(w_n10358_0[0]),.doutb(w_n10358_0[1]),.din(n10358));
	jspl jspl_w_n10364_0(.douta(w_n10364_0[0]),.doutb(w_n10364_0[1]),.din(n10364));
	jspl jspl_w_n10366_0(.douta(w_n10366_0[0]),.doutb(w_n10366_0[1]),.din(n10366));
	jspl3 jspl3_w_n10367_0(.douta(w_n10367_0[0]),.doutb(w_n10367_0[1]),.doutc(w_n10367_0[2]),.din(n10367));
	jspl jspl_w_n10371_0(.douta(w_n10371_0[0]),.doutb(w_n10371_0[1]),.din(n10371));
	jspl jspl_w_n10372_0(.douta(w_n10372_0[0]),.doutb(w_n10372_0[1]),.din(n10372));
	jspl3 jspl3_w_n10373_0(.douta(w_n10373_0[0]),.doutb(w_n10373_0[1]),.doutc(w_n10373_0[2]),.din(n10373));
	jspl jspl_w_n10375_0(.douta(w_n10375_0[0]),.doutb(w_n10375_0[1]),.din(n10375));
	jspl jspl_w_n10380_0(.douta(w_n10380_0[0]),.doutb(w_n10380_0[1]),.din(n10380));
	jspl jspl_w_n10382_0(.douta(w_n10382_0[0]),.doutb(w_n10382_0[1]),.din(n10382));
	jspl jspl_w_n10383_0(.douta(w_n10383_0[0]),.doutb(w_n10383_0[1]),.din(n10383));
	jspl3 jspl3_w_n10384_0(.douta(w_n10384_0[0]),.doutb(w_n10384_0[1]),.doutc(w_n10384_0[2]),.din(n10384));
	jspl jspl_w_n10385_0(.douta(w_n10385_0[0]),.doutb(w_n10385_0[1]),.din(n10385));
	jspl jspl_w_n10389_0(.douta(w_n10389_0[0]),.doutb(w_n10389_0[1]),.din(n10389));
	jspl jspl_w_n10395_0(.douta(w_n10395_0[0]),.doutb(w_n10395_0[1]),.din(n10395));
	jspl jspl_w_n10396_0(.douta(w_n10396_0[0]),.doutb(w_n10396_0[1]),.din(n10396));
	jspl jspl_w_n10398_0(.douta(w_n10398_0[0]),.doutb(w_n10398_0[1]),.din(n10398));
	jspl jspl_w_n10400_0(.douta(w_n10400_0[0]),.doutb(w_n10400_0[1]),.din(n10400));
	jspl jspl_w_n10403_0(.douta(w_n10403_0[0]),.doutb(w_n10403_0[1]),.din(n10403));
	jspl jspl_w_n10409_0(.douta(w_n10409_0[0]),.doutb(w_n10409_0[1]),.din(n10409));
	jspl jspl_w_n10411_0(.douta(w_n10411_0[0]),.doutb(w_n10411_0[1]),.din(n10411));
	jspl3 jspl3_w_n10412_0(.douta(w_n10412_0[0]),.doutb(w_n10412_0[1]),.doutc(w_n10412_0[2]),.din(n10412));
	jspl jspl_w_n10416_0(.douta(w_n10416_0[0]),.doutb(w_n10416_0[1]),.din(n10416));
	jspl jspl_w_n10417_0(.douta(w_n10417_0[0]),.doutb(w_n10417_0[1]),.din(n10417));
	jspl3 jspl3_w_n10418_0(.douta(w_n10418_0[0]),.doutb(w_n10418_0[1]),.doutc(w_n10418_0[2]),.din(n10418));
	jspl jspl_w_n10420_0(.douta(w_n10420_0[0]),.doutb(w_n10420_0[1]),.din(n10420));
	jspl jspl_w_n10425_0(.douta(w_n10425_0[0]),.doutb(w_n10425_0[1]),.din(n10425));
	jspl jspl_w_n10427_0(.douta(w_n10427_0[0]),.doutb(w_n10427_0[1]),.din(n10427));
	jspl jspl_w_n10428_0(.douta(w_n10428_0[0]),.doutb(w_n10428_0[1]),.din(n10428));
	jspl3 jspl3_w_n10429_0(.douta(w_n10429_0[0]),.doutb(w_n10429_0[1]),.doutc(w_n10429_0[2]),.din(n10429));
	jspl jspl_w_n10430_0(.douta(w_n10430_0[0]),.doutb(w_n10430_0[1]),.din(n10430));
	jspl jspl_w_n10434_0(.douta(w_n10434_0[0]),.doutb(w_n10434_0[1]),.din(n10434));
	jspl jspl_w_n10440_0(.douta(w_n10440_0[0]),.doutb(w_n10440_0[1]),.din(n10440));
	jspl jspl_w_n10441_0(.douta(w_n10441_0[0]),.doutb(w_n10441_0[1]),.din(n10441));
	jspl jspl_w_n10443_0(.douta(w_n10443_0[0]),.doutb(w_n10443_0[1]),.din(n10443));
	jspl jspl_w_n10448_0(.douta(w_n10448_0[0]),.doutb(w_n10448_0[1]),.din(n10448));
	jspl jspl_w_n10450_0(.douta(w_n10450_0[0]),.doutb(w_n10450_0[1]),.din(n10450));
	jspl jspl_w_n10451_0(.douta(w_n10451_0[0]),.doutb(w_n10451_0[1]),.din(n10451));
	jspl3 jspl3_w_n10452_0(.douta(w_n10452_0[0]),.doutb(w_n10452_0[1]),.doutc(w_n10452_0[2]),.din(n10452));
	jspl jspl_w_n10453_0(.douta(w_n10453_0[0]),.doutb(w_n10453_0[1]),.din(n10453));
	jspl jspl_w_n10455_0(.douta(w_n10455_0[0]),.doutb(w_n10455_0[1]),.din(n10455));
	jspl jspl_w_n10457_0(.douta(w_n10457_0[0]),.doutb(w_n10457_0[1]),.din(n10457));
	jspl jspl_w_n10459_0(.douta(w_n10459_0[0]),.doutb(w_n10459_0[1]),.din(n10459));
	jspl jspl_w_n10462_0(.douta(w_n10462_0[0]),.doutb(w_n10462_0[1]),.din(n10462));
	jspl jspl_w_n10468_0(.douta(w_n10468_0[0]),.doutb(w_n10468_0[1]),.din(n10468));
	jspl3 jspl3_w_n10470_0(.douta(w_n10470_0[0]),.doutb(w_n10470_0[1]),.doutc(w_n10470_0[2]),.din(n10470));
	jspl jspl_w_n10471_0(.douta(w_n10471_0[0]),.doutb(w_n10471_0[1]),.din(n10471));
	jspl jspl_w_n10475_0(.douta(w_n10475_0[0]),.doutb(w_n10475_0[1]),.din(n10475));
	jspl jspl_w_n10481_0(.douta(w_n10481_0[0]),.doutb(w_n10481_0[1]),.din(n10481));
	jspl jspl_w_n10482_0(.douta(w_n10482_0[0]),.doutb(w_n10482_0[1]),.din(n10482));
	jspl jspl_w_n10484_0(.douta(w_n10484_0[0]),.doutb(w_n10484_0[1]),.din(n10484));
	jspl jspl_w_n10486_0(.douta(w_n10486_0[0]),.doutb(w_n10486_0[1]),.din(n10486));
	jspl jspl_w_n10489_0(.douta(w_n10489_0[0]),.doutb(w_n10489_0[1]),.din(n10489));
	jspl jspl_w_n10495_0(.douta(w_n10495_0[0]),.doutb(w_n10495_0[1]),.din(n10495));
	jspl jspl_w_n10497_0(.douta(w_n10497_0[0]),.doutb(w_n10497_0[1]),.din(n10497));
	jspl3 jspl3_w_n10498_0(.douta(w_n10498_0[0]),.doutb(w_n10498_0[1]),.doutc(w_n10498_0[2]),.din(n10498));
	jspl jspl_w_n10502_0(.douta(w_n10502_0[0]),.doutb(w_n10502_0[1]),.din(n10502));
	jspl jspl_w_n10503_0(.douta(w_n10503_0[0]),.doutb(w_n10503_0[1]),.din(n10503));
	jspl3 jspl3_w_n10504_0(.douta(w_n10504_0[0]),.doutb(w_n10504_0[1]),.doutc(w_n10504_0[2]),.din(n10504));
	jspl jspl_w_n10506_0(.douta(w_n10506_0[0]),.doutb(w_n10506_0[1]),.din(n10506));
	jspl jspl_w_n10511_0(.douta(w_n10511_0[0]),.doutb(w_n10511_0[1]),.din(n10511));
	jspl jspl_w_n10513_0(.douta(w_n10513_0[0]),.doutb(w_n10513_0[1]),.din(n10513));
	jspl jspl_w_n10514_0(.douta(w_n10514_0[0]),.doutb(w_n10514_0[1]),.din(n10514));
	jspl3 jspl3_w_n10515_0(.douta(w_n10515_0[0]),.doutb(w_n10515_0[1]),.doutc(w_n10515_0[2]),.din(n10515));
	jspl jspl_w_n10516_0(.douta(w_n10516_0[0]),.doutb(w_n10516_0[1]),.din(n10516));
	jspl jspl_w_n10520_0(.douta(w_n10520_0[0]),.doutb(w_n10520_0[1]),.din(n10520));
	jspl jspl_w_n10526_0(.douta(w_n10526_0[0]),.doutb(w_n10526_0[1]),.din(n10526));
	jspl jspl_w_n10527_0(.douta(w_n10527_0[0]),.doutb(w_n10527_0[1]),.din(n10527));
	jspl jspl_w_n10529_0(.douta(w_n10529_0[0]),.doutb(w_n10529_0[1]),.din(n10529));
	jspl jspl_w_n10531_0(.douta(w_n10531_0[0]),.doutb(w_n10531_0[1]),.din(n10531));
	jspl jspl_w_n10534_0(.douta(w_n10534_0[0]),.doutb(w_n10534_0[1]),.din(n10534));
	jspl jspl_w_n10540_0(.douta(w_n10540_0[0]),.doutb(w_n10540_0[1]),.din(n10540));
	jspl jspl_w_n10542_0(.douta(w_n10542_0[0]),.doutb(w_n10542_0[1]),.din(n10542));
	jspl3 jspl3_w_n10543_0(.douta(w_n10543_0[0]),.doutb(w_n10543_0[1]),.doutc(w_n10543_0[2]),.din(n10543));
	jspl jspl_w_n10547_0(.douta(w_n10547_0[0]),.doutb(w_n10547_0[1]),.din(n10547));
	jspl jspl_w_n10548_0(.douta(w_n10548_0[0]),.doutb(w_n10548_0[1]),.din(n10548));
	jspl3 jspl3_w_n10549_0(.douta(w_n10549_0[0]),.doutb(w_n10549_0[1]),.doutc(w_n10549_0[2]),.din(n10549));
	jspl jspl_w_n10551_0(.douta(w_n10551_0[0]),.doutb(w_n10551_0[1]),.din(n10551));
	jspl jspl_w_n10556_0(.douta(w_n10556_0[0]),.doutb(w_n10556_0[1]),.din(n10556));
	jspl jspl_w_n10558_0(.douta(w_n10558_0[0]),.doutb(w_n10558_0[1]),.din(n10558));
	jspl jspl_w_n10559_0(.douta(w_n10559_0[0]),.doutb(w_n10559_0[1]),.din(n10559));
	jspl3 jspl3_w_n10560_0(.douta(w_n10560_0[0]),.doutb(w_n10560_0[1]),.doutc(w_n10560_0[2]),.din(n10560));
	jspl jspl_w_n10561_0(.douta(w_n10561_0[0]),.doutb(w_n10561_0[1]),.din(n10561));
	jspl jspl_w_n10565_0(.douta(w_n10565_0[0]),.doutb(w_n10565_0[1]),.din(n10565));
	jspl jspl_w_n10571_0(.douta(w_n10571_0[0]),.doutb(w_n10571_0[1]),.din(n10571));
	jspl jspl_w_n10572_0(.douta(w_n10572_0[0]),.doutb(w_n10572_0[1]),.din(n10572));
	jspl jspl_w_n10574_0(.douta(w_n10574_0[0]),.doutb(w_n10574_0[1]),.din(n10574));
	jspl jspl_w_n10576_0(.douta(w_n10576_0[0]),.doutb(w_n10576_0[1]),.din(n10576));
	jspl jspl_w_n10579_0(.douta(w_n10579_0[0]),.doutb(w_n10579_0[1]),.din(n10579));
	jspl jspl_w_n10585_0(.douta(w_n10585_0[0]),.doutb(w_n10585_0[1]),.din(n10585));
	jspl jspl_w_n10587_0(.douta(w_n10587_0[0]),.doutb(w_n10587_0[1]),.din(n10587));
	jspl3 jspl3_w_n10588_0(.douta(w_n10588_0[0]),.doutb(w_n10588_0[1]),.doutc(w_n10588_0[2]),.din(n10588));
	jspl jspl_w_n10592_0(.douta(w_n10592_0[0]),.doutb(w_n10592_0[1]),.din(n10592));
	jspl jspl_w_n10593_0(.douta(w_n10593_0[0]),.doutb(w_n10593_0[1]),.din(n10593));
	jspl3 jspl3_w_n10594_0(.douta(w_n10594_0[0]),.doutb(w_n10594_0[1]),.doutc(w_n10594_0[2]),.din(n10594));
	jspl jspl_w_n10596_0(.douta(w_n10596_0[0]),.doutb(w_n10596_0[1]),.din(n10596));
	jspl jspl_w_n10601_0(.douta(w_n10601_0[0]),.doutb(w_n10601_0[1]),.din(n10601));
	jspl jspl_w_n10603_0(.douta(w_n10603_0[0]),.doutb(w_n10603_0[1]),.din(n10603));
	jspl jspl_w_n10604_0(.douta(w_n10604_0[0]),.doutb(w_n10604_0[1]),.din(n10604));
	jspl3 jspl3_w_n10605_0(.douta(w_n10605_0[0]),.doutb(w_n10605_0[1]),.doutc(w_n10605_0[2]),.din(n10605));
	jspl jspl_w_n10606_0(.douta(w_n10606_0[0]),.doutb(w_n10606_0[1]),.din(n10606));
	jspl jspl_w_n10610_0(.douta(w_n10610_0[0]),.doutb(w_n10610_0[1]),.din(n10610));
	jspl jspl_w_n10616_0(.douta(w_n10616_0[0]),.doutb(w_n10616_0[1]),.din(n10616));
	jspl jspl_w_n10617_0(.douta(w_n10617_0[0]),.doutb(w_n10617_0[1]),.din(n10617));
	jspl jspl_w_n10619_0(.douta(w_n10619_0[0]),.doutb(w_n10619_0[1]),.din(n10619));
	jspl jspl_w_n10621_0(.douta(w_n10621_0[0]),.doutb(w_n10621_0[1]),.din(n10621));
	jspl jspl_w_n10624_0(.douta(w_n10624_0[0]),.doutb(w_n10624_0[1]),.din(n10624));
	jspl jspl_w_n10630_0(.douta(w_n10630_0[0]),.doutb(w_n10630_0[1]),.din(n10630));
	jspl jspl_w_n10632_0(.douta(w_n10632_0[0]),.doutb(w_n10632_0[1]),.din(n10632));
	jspl3 jspl3_w_n10633_0(.douta(w_n10633_0[0]),.doutb(w_n10633_0[1]),.doutc(w_n10633_0[2]),.din(n10633));
	jspl jspl_w_n10637_0(.douta(w_n10637_0[0]),.doutb(w_n10637_0[1]),.din(n10637));
	jspl jspl_w_n10638_0(.douta(w_n10638_0[0]),.doutb(w_n10638_0[1]),.din(n10638));
	jspl3 jspl3_w_n10639_0(.douta(w_n10639_0[0]),.doutb(w_n10639_0[1]),.doutc(w_n10639_0[2]),.din(n10639));
	jspl jspl_w_n10641_0(.douta(w_n10641_0[0]),.doutb(w_n10641_0[1]),.din(n10641));
	jspl jspl_w_n10646_0(.douta(w_n10646_0[0]),.doutb(w_n10646_0[1]),.din(n10646));
	jspl jspl_w_n10648_0(.douta(w_n10648_0[0]),.doutb(w_n10648_0[1]),.din(n10648));
	jspl jspl_w_n10649_0(.douta(w_n10649_0[0]),.doutb(w_n10649_0[1]),.din(n10649));
	jspl3 jspl3_w_n10650_0(.douta(w_n10650_0[0]),.doutb(w_n10650_0[1]),.doutc(w_n10650_0[2]),.din(n10650));
	jspl jspl_w_n10651_0(.douta(w_n10651_0[0]),.doutb(w_n10651_0[1]),.din(n10651));
	jspl jspl_w_n10655_0(.douta(w_n10655_0[0]),.doutb(w_n10655_0[1]),.din(n10655));
	jspl jspl_w_n10661_0(.douta(w_n10661_0[0]),.doutb(w_n10661_0[1]),.din(n10661));
	jspl jspl_w_n10662_0(.douta(w_n10662_0[0]),.doutb(w_n10662_0[1]),.din(n10662));
	jspl jspl_w_n10664_0(.douta(w_n10664_0[0]),.doutb(w_n10664_0[1]),.din(n10664));
	jspl jspl_w_n10666_0(.douta(w_n10666_0[0]),.doutb(w_n10666_0[1]),.din(n10666));
	jspl jspl_w_n10669_0(.douta(w_n10669_0[0]),.doutb(w_n10669_0[1]),.din(n10669));
	jspl jspl_w_n10675_0(.douta(w_n10675_0[0]),.doutb(w_n10675_0[1]),.din(n10675));
	jspl3 jspl3_w_n10677_0(.douta(w_n10677_0[0]),.doutb(w_n10677_0[1]),.doutc(w_n10677_0[2]),.din(n10677));
	jspl3 jspl3_w_n10677_1(.douta(w_n10677_1[0]),.doutb(w_n10677_1[1]),.doutc(w_n10677_1[2]),.din(w_n10677_0[0]));
	jspl jspl_w_n10680_0(.douta(w_n10680_0[0]),.doutb(w_n10680_0[1]),.din(n10680));
	jspl3 jspl3_w_n10681_0(.douta(w_n10681_0[0]),.doutb(w_n10681_0[1]),.doutc(w_n10681_0[2]),.din(n10681));
	jspl jspl_w_n10682_0(.douta(w_n10682_0[0]),.doutb(w_n10682_0[1]),.din(n10682));
	jspl jspl_w_n10688_0(.douta(w_n10688_0[0]),.doutb(w_n10688_0[1]),.din(n10688));
	jspl3 jspl3_w_n10689_0(.douta(w_n10689_0[0]),.doutb(w_n10689_0[1]),.doutc(w_n10689_0[2]),.din(n10689));
	jspl jspl_w_n10690_0(.douta(w_n10690_0[0]),.doutb(w_n10690_0[1]),.din(n10690));
	jspl jspl_w_n10695_0(.douta(w_n10695_0[0]),.doutb(w_n10695_0[1]),.din(n10695));
	jspl3 jspl3_w_n10696_0(.douta(w_n10696_0[0]),.doutb(w_n10696_0[1]),.doutc(w_n10696_0[2]),.din(n10696));
	jspl3 jspl3_w_n10696_1(.douta(w_n10696_1[0]),.doutb(w_n10696_1[1]),.doutc(w_n10696_1[2]),.din(w_n10696_0[0]));
	jspl3 jspl3_w_n10696_2(.douta(w_n10696_2[0]),.doutb(w_n10696_2[1]),.doutc(w_n10696_2[2]),.din(w_n10696_0[1]));
	jspl3 jspl3_w_n10696_3(.douta(w_n10696_3[0]),.doutb(w_n10696_3[1]),.doutc(w_n10696_3[2]),.din(w_n10696_0[2]));
	jspl3 jspl3_w_n10696_4(.douta(w_n10696_4[0]),.doutb(w_n10696_4[1]),.doutc(w_n10696_4[2]),.din(w_n10696_1[0]));
	jspl3 jspl3_w_n10696_5(.douta(w_n10696_5[0]),.doutb(w_n10696_5[1]),.doutc(w_n10696_5[2]),.din(w_n10696_1[1]));
	jspl3 jspl3_w_n10696_6(.douta(w_n10696_6[0]),.doutb(w_n10696_6[1]),.doutc(w_n10696_6[2]),.din(w_n10696_1[2]));
	jspl3 jspl3_w_n10696_7(.douta(w_n10696_7[0]),.doutb(w_n10696_7[1]),.doutc(w_n10696_7[2]),.din(w_n10696_2[0]));
	jspl3 jspl3_w_n10696_8(.douta(w_n10696_8[0]),.doutb(w_n10696_8[1]),.doutc(w_n10696_8[2]),.din(w_n10696_2[1]));
	jspl3 jspl3_w_n10696_9(.douta(w_n10696_9[0]),.doutb(w_n10696_9[1]),.doutc(w_n10696_9[2]),.din(w_n10696_2[2]));
	jspl3 jspl3_w_n10696_10(.douta(w_n10696_10[0]),.doutb(w_n10696_10[1]),.doutc(w_n10696_10[2]),.din(w_n10696_3[0]));
	jspl3 jspl3_w_n10696_11(.douta(w_n10696_11[0]),.doutb(w_n10696_11[1]),.doutc(w_n10696_11[2]),.din(w_n10696_3[1]));
	jspl3 jspl3_w_n10696_12(.douta(w_n10696_12[0]),.doutb(w_n10696_12[1]),.doutc(w_n10696_12[2]),.din(w_n10696_3[2]));
	jspl jspl_w_n10696_13(.douta(w_n10696_13[0]),.doutb(w_n10696_13[1]),.din(w_n10696_4[0]));
	jspl3 jspl3_w_n10701_0(.douta(w_n10701_0[0]),.doutb(w_n10701_0[1]),.doutc(w_n10701_0[2]),.din(n10701));
	jspl3 jspl3_w_n10701_1(.douta(w_n10701_1[0]),.doutb(w_n10701_1[1]),.doutc(w_n10701_1[2]),.din(w_n10701_0[0]));
	jspl3 jspl3_w_n10701_2(.douta(w_n10701_2[0]),.doutb(w_n10701_2[1]),.doutc(w_n10701_2[2]),.din(w_n10701_0[1]));
	jspl3 jspl3_w_n10701_3(.douta(w_n10701_3[0]),.doutb(w_n10701_3[1]),.doutc(w_n10701_3[2]),.din(w_n10701_0[2]));
	jspl3 jspl3_w_n10701_4(.douta(w_n10701_4[0]),.doutb(w_n10701_4[1]),.doutc(w_n10701_4[2]),.din(w_n10701_1[0]));
	jspl3 jspl3_w_n10701_5(.douta(w_n10701_5[0]),.doutb(w_n10701_5[1]),.doutc(w_n10701_5[2]),.din(w_n10701_1[1]));
	jspl3 jspl3_w_n10701_6(.douta(w_n10701_6[0]),.doutb(w_n10701_6[1]),.doutc(w_n10701_6[2]),.din(w_n10701_1[2]));
	jspl3 jspl3_w_n10701_7(.douta(w_n10701_7[0]),.doutb(w_n10701_7[1]),.doutc(w_n10701_7[2]),.din(w_n10701_2[0]));
	jspl3 jspl3_w_n10701_8(.douta(w_n10701_8[0]),.doutb(w_n10701_8[1]),.doutc(w_n10701_8[2]),.din(w_n10701_2[1]));
	jspl3 jspl3_w_n10701_9(.douta(w_n10701_9[0]),.doutb(w_n10701_9[1]),.doutc(w_n10701_9[2]),.din(w_n10701_2[2]));
	jspl3 jspl3_w_n10701_10(.douta(w_n10701_10[0]),.doutb(w_n10701_10[1]),.doutc(w_n10701_10[2]),.din(w_n10701_3[0]));
	jspl3 jspl3_w_n10701_11(.douta(w_n10701_11[0]),.doutb(w_n10701_11[1]),.doutc(w_n10701_11[2]),.din(w_n10701_3[1]));
	jspl3 jspl3_w_n10701_12(.douta(w_n10701_12[0]),.doutb(w_n10701_12[1]),.doutc(w_n10701_12[2]),.din(w_n10701_3[2]));
	jspl3 jspl3_w_n10701_13(.douta(w_n10701_13[0]),.doutb(w_n10701_13[1]),.doutc(w_n10701_13[2]),.din(w_n10701_4[0]));
	jspl3 jspl3_w_n10701_14(.douta(w_n10701_14[0]),.doutb(w_n10701_14[1]),.doutc(w_n10701_14[2]),.din(w_n10701_4[1]));
	jspl3 jspl3_w_n10701_15(.douta(w_n10701_15[0]),.doutb(w_n10701_15[1]),.doutc(w_n10701_15[2]),.din(w_n10701_4[2]));
	jspl3 jspl3_w_n10701_16(.douta(w_n10701_16[0]),.doutb(w_n10701_16[1]),.doutc(w_n10701_16[2]),.din(w_n10701_5[0]));
	jspl3 jspl3_w_n10701_17(.douta(w_n10701_17[0]),.doutb(w_n10701_17[1]),.doutc(w_n10701_17[2]),.din(w_n10701_5[1]));
	jspl3 jspl3_w_n10701_18(.douta(w_n10701_18[0]),.doutb(w_n10701_18[1]),.doutc(w_n10701_18[2]),.din(w_n10701_5[2]));
	jspl3 jspl3_w_n10701_19(.douta(w_n10701_19[0]),.doutb(w_n10701_19[1]),.doutc(w_n10701_19[2]),.din(w_n10701_6[0]));
	jspl3 jspl3_w_n10701_20(.douta(w_n10701_20[0]),.doutb(w_n10701_20[1]),.doutc(w_n10701_20[2]),.din(w_n10701_6[1]));
	jspl3 jspl3_w_n10701_21(.douta(w_n10701_21[0]),.doutb(w_n10701_21[1]),.doutc(w_n10701_21[2]),.din(w_n10701_6[2]));
	jspl3 jspl3_w_n10701_22(.douta(w_n10701_22[0]),.doutb(w_n10701_22[1]),.doutc(w_n10701_22[2]),.din(w_n10701_7[0]));
	jspl3 jspl3_w_n10701_23(.douta(w_n10701_23[0]),.doutb(w_n10701_23[1]),.doutc(w_n10701_23[2]),.din(w_n10701_7[1]));
	jspl3 jspl3_w_n10701_24(.douta(w_n10701_24[0]),.doutb(w_n10701_24[1]),.doutc(w_n10701_24[2]),.din(w_n10701_7[2]));
	jspl3 jspl3_w_n10701_25(.douta(w_n10701_25[0]),.doutb(w_n10701_25[1]),.doutc(w_n10701_25[2]),.din(w_n10701_8[0]));
	jspl jspl_w_n10704_0(.douta(w_n10704_0[0]),.doutb(w_n10704_0[1]),.din(n10704));
	jspl3 jspl3_w_n10706_0(.douta(w_n10706_0[0]),.doutb(w_n10706_0[1]),.doutc(w_n10706_0[2]),.din(n10706));
	jspl jspl_w_n10706_1(.douta(w_n10706_1[0]),.doutb(w_n10706_1[1]),.din(w_n10706_0[0]));
	jspl3 jspl3_w_n10707_0(.douta(w_n10707_0[0]),.doutb(w_n10707_0[1]),.doutc(w_n10707_0[2]),.din(n10707));
	jspl3 jspl3_w_n10711_0(.douta(w_n10711_0[0]),.doutb(w_n10711_0[1]),.doutc(w_n10711_0[2]),.din(n10711));
	jspl jspl_w_n10712_0(.douta(w_n10712_0[0]),.doutb(w_n10712_0[1]),.din(n10712));
	jspl jspl_w_n10713_0(.douta(w_n10713_0[0]),.doutb(w_n10713_0[1]),.din(n10713));
	jspl jspl_w_n10714_0(.douta(w_n10714_0[0]),.doutb(w_n10714_0[1]),.din(n10714));
	jspl jspl_w_n10716_0(.douta(w_n10716_0[0]),.doutb(w_n10716_0[1]),.din(n10716));
	jspl jspl_w_n10718_0(.douta(w_n10718_0[0]),.doutb(w_n10718_0[1]),.din(n10718));
	jspl jspl_w_n10720_0(.douta(w_n10720_0[0]),.doutb(w_n10720_0[1]),.din(n10720));
	jspl jspl_w_n10723_0(.douta(w_n10723_0[0]),.doutb(w_n10723_0[1]),.din(n10723));
	jspl jspl_w_n10728_0(.douta(w_n10728_0[0]),.doutb(w_n10728_0[1]),.din(n10728));
	jspl3 jspl3_w_n10730_0(.douta(w_n10730_0[0]),.doutb(w_n10730_0[1]),.doutc(w_n10730_0[2]),.din(n10730));
	jspl jspl_w_n10731_0(.douta(w_n10731_0[0]),.doutb(w_n10731_0[1]),.din(n10731));
	jspl jspl_w_n10735_0(.douta(w_n10735_0[0]),.doutb(w_n10735_0[1]),.din(n10735));
	jspl jspl_w_n10736_0(.douta(w_n10736_0[0]),.doutb(w_n10736_0[1]),.din(n10736));
	jspl jspl_w_n10738_0(.douta(w_n10738_0[0]),.doutb(w_n10738_0[1]),.din(n10738));
	jspl jspl_w_n10742_0(.douta(w_n10742_0[0]),.doutb(w_n10742_0[1]),.din(n10742));
	jspl jspl_w_n10744_0(.douta(w_n10744_0[0]),.doutb(w_n10744_0[1]),.din(n10744));
	jspl jspl_w_n10745_0(.douta(w_n10745_0[0]),.doutb(w_n10745_0[1]),.din(n10745));
	jspl3 jspl3_w_n10746_0(.douta(w_n10746_0[0]),.doutb(w_n10746_0[1]),.doutc(w_n10746_0[2]),.din(n10746));
	jspl jspl_w_n10747_0(.douta(w_n10747_0[0]),.doutb(w_n10747_0[1]),.din(n10747));
	jspl jspl_w_n10751_0(.douta(w_n10751_0[0]),.doutb(w_n10751_0[1]),.din(n10751));
	jspl jspl_w_n10753_0(.douta(w_n10753_0[0]),.doutb(w_n10753_0[1]),.din(n10753));
	jspl jspl_w_n10755_0(.douta(w_n10755_0[0]),.doutb(w_n10755_0[1]),.din(n10755));
	jspl jspl_w_n10757_0(.douta(w_n10757_0[0]),.doutb(w_n10757_0[1]),.din(n10757));
	jspl jspl_w_n10760_0(.douta(w_n10760_0[0]),.doutb(w_n10760_0[1]),.din(n10760));
	jspl jspl_w_n10766_0(.douta(w_n10766_0[0]),.doutb(w_n10766_0[1]),.din(n10766));
	jspl3 jspl3_w_n10768_0(.douta(w_n10768_0[0]),.doutb(w_n10768_0[1]),.doutc(w_n10768_0[2]),.din(n10768));
	jspl jspl_w_n10769_0(.douta(w_n10769_0[0]),.doutb(w_n10769_0[1]),.din(n10769));
	jspl jspl_w_n10774_0(.douta(w_n10774_0[0]),.doutb(w_n10774_0[1]),.din(n10774));
	jspl jspl_w_n10776_0(.douta(w_n10776_0[0]),.doutb(w_n10776_0[1]),.din(n10776));
	jspl jspl_w_n10778_0(.douta(w_n10778_0[0]),.doutb(w_n10778_0[1]),.din(n10778));
	jspl jspl_w_n10782_0(.douta(w_n10782_0[0]),.doutb(w_n10782_0[1]),.din(n10782));
	jspl jspl_w_n10784_0(.douta(w_n10784_0[0]),.doutb(w_n10784_0[1]),.din(n10784));
	jspl jspl_w_n10785_0(.douta(w_n10785_0[0]),.doutb(w_n10785_0[1]),.din(n10785));
	jspl3 jspl3_w_n10786_0(.douta(w_n10786_0[0]),.doutb(w_n10786_0[1]),.doutc(w_n10786_0[2]),.din(n10786));
	jspl jspl_w_n10787_0(.douta(w_n10787_0[0]),.doutb(w_n10787_0[1]),.din(n10787));
	jspl jspl_w_n10793_0(.douta(w_n10793_0[0]),.doutb(w_n10793_0[1]),.din(n10793));
	jspl jspl_w_n10794_0(.douta(w_n10794_0[0]),.doutb(w_n10794_0[1]),.din(n10794));
	jspl jspl_w_n10796_0(.douta(w_n10796_0[0]),.doutb(w_n10796_0[1]),.din(n10796));
	jspl jspl_w_n10798_0(.douta(w_n10798_0[0]),.doutb(w_n10798_0[1]),.din(n10798));
	jspl jspl_w_n10800_0(.douta(w_n10800_0[0]),.doutb(w_n10800_0[1]),.din(n10800));
	jspl jspl_w_n10806_0(.douta(w_n10806_0[0]),.doutb(w_n10806_0[1]),.din(n10806));
	jspl jspl_w_n10808_0(.douta(w_n10808_0[0]),.doutb(w_n10808_0[1]),.din(n10808));
	jspl3 jspl3_w_n10809_0(.douta(w_n10809_0[0]),.doutb(w_n10809_0[1]),.doutc(w_n10809_0[2]),.din(n10809));
	jspl jspl_w_n10812_0(.douta(w_n10812_0[0]),.doutb(w_n10812_0[1]),.din(n10812));
	jspl jspl_w_n10813_0(.douta(w_n10813_0[0]),.doutb(w_n10813_0[1]),.din(n10813));
	jspl3 jspl3_w_n10814_0(.douta(w_n10814_0[0]),.doutb(w_n10814_0[1]),.doutc(w_n10814_0[2]),.din(n10814));
	jspl jspl_w_n10816_0(.douta(w_n10816_0[0]),.doutb(w_n10816_0[1]),.din(n10816));
	jspl jspl_w_n10820_0(.douta(w_n10820_0[0]),.doutb(w_n10820_0[1]),.din(n10820));
	jspl jspl_w_n10822_0(.douta(w_n10822_0[0]),.doutb(w_n10822_0[1]),.din(n10822));
	jspl jspl_w_n10823_0(.douta(w_n10823_0[0]),.doutb(w_n10823_0[1]),.din(n10823));
	jspl3 jspl3_w_n10824_0(.douta(w_n10824_0[0]),.doutb(w_n10824_0[1]),.doutc(w_n10824_0[2]),.din(n10824));
	jspl jspl_w_n10825_0(.douta(w_n10825_0[0]),.doutb(w_n10825_0[1]),.din(n10825));
	jspl jspl_w_n10828_0(.douta(w_n10828_0[0]),.doutb(w_n10828_0[1]),.din(n10828));
	jspl jspl_w_n10834_0(.douta(w_n10834_0[0]),.doutb(w_n10834_0[1]),.din(n10834));
	jspl jspl_w_n10835_0(.douta(w_n10835_0[0]),.doutb(w_n10835_0[1]),.din(n10835));
	jspl jspl_w_n10837_0(.douta(w_n10837_0[0]),.doutb(w_n10837_0[1]),.din(n10837));
	jspl jspl_w_n10839_0(.douta(w_n10839_0[0]),.doutb(w_n10839_0[1]),.din(n10839));
	jspl jspl_w_n10841_0(.douta(w_n10841_0[0]),.doutb(w_n10841_0[1]),.din(n10841));
	jspl jspl_w_n10847_0(.douta(w_n10847_0[0]),.doutb(w_n10847_0[1]),.din(n10847));
	jspl jspl_w_n10849_0(.douta(w_n10849_0[0]),.doutb(w_n10849_0[1]),.din(n10849));
	jspl3 jspl3_w_n10850_0(.douta(w_n10850_0[0]),.doutb(w_n10850_0[1]),.doutc(w_n10850_0[2]),.din(n10850));
	jspl jspl_w_n10853_0(.douta(w_n10853_0[0]),.doutb(w_n10853_0[1]),.din(n10853));
	jspl jspl_w_n10854_0(.douta(w_n10854_0[0]),.doutb(w_n10854_0[1]),.din(n10854));
	jspl3 jspl3_w_n10855_0(.douta(w_n10855_0[0]),.doutb(w_n10855_0[1]),.doutc(w_n10855_0[2]),.din(n10855));
	jspl jspl_w_n10857_0(.douta(w_n10857_0[0]),.doutb(w_n10857_0[1]),.din(n10857));
	jspl jspl_w_n10861_0(.douta(w_n10861_0[0]),.doutb(w_n10861_0[1]),.din(n10861));
	jspl jspl_w_n10863_0(.douta(w_n10863_0[0]),.doutb(w_n10863_0[1]),.din(n10863));
	jspl jspl_w_n10864_0(.douta(w_n10864_0[0]),.doutb(w_n10864_0[1]),.din(n10864));
	jspl3 jspl3_w_n10865_0(.douta(w_n10865_0[0]),.doutb(w_n10865_0[1]),.doutc(w_n10865_0[2]),.din(n10865));
	jspl jspl_w_n10866_0(.douta(w_n10866_0[0]),.doutb(w_n10866_0[1]),.din(n10866));
	jspl jspl_w_n10869_0(.douta(w_n10869_0[0]),.doutb(w_n10869_0[1]),.din(n10869));
	jspl jspl_w_n10875_0(.douta(w_n10875_0[0]),.doutb(w_n10875_0[1]),.din(n10875));
	jspl jspl_w_n10876_0(.douta(w_n10876_0[0]),.doutb(w_n10876_0[1]),.din(n10876));
	jspl jspl_w_n10878_0(.douta(w_n10878_0[0]),.doutb(w_n10878_0[1]),.din(n10878));
	jspl jspl_w_n10880_0(.douta(w_n10880_0[0]),.doutb(w_n10880_0[1]),.din(n10880));
	jspl jspl_w_n10882_0(.douta(w_n10882_0[0]),.doutb(w_n10882_0[1]),.din(n10882));
	jspl jspl_w_n10888_0(.douta(w_n10888_0[0]),.doutb(w_n10888_0[1]),.din(n10888));
	jspl jspl_w_n10890_0(.douta(w_n10890_0[0]),.doutb(w_n10890_0[1]),.din(n10890));
	jspl3 jspl3_w_n10891_0(.douta(w_n10891_0[0]),.doutb(w_n10891_0[1]),.doutc(w_n10891_0[2]),.din(n10891));
	jspl jspl_w_n10894_0(.douta(w_n10894_0[0]),.doutb(w_n10894_0[1]),.din(n10894));
	jspl jspl_w_n10895_0(.douta(w_n10895_0[0]),.doutb(w_n10895_0[1]),.din(n10895));
	jspl3 jspl3_w_n10896_0(.douta(w_n10896_0[0]),.doutb(w_n10896_0[1]),.doutc(w_n10896_0[2]),.din(n10896));
	jspl jspl_w_n10898_0(.douta(w_n10898_0[0]),.doutb(w_n10898_0[1]),.din(n10898));
	jspl jspl_w_n10902_0(.douta(w_n10902_0[0]),.doutb(w_n10902_0[1]),.din(n10902));
	jspl jspl_w_n10904_0(.douta(w_n10904_0[0]),.doutb(w_n10904_0[1]),.din(n10904));
	jspl jspl_w_n10905_0(.douta(w_n10905_0[0]),.doutb(w_n10905_0[1]),.din(n10905));
	jspl3 jspl3_w_n10906_0(.douta(w_n10906_0[0]),.doutb(w_n10906_0[1]),.doutc(w_n10906_0[2]),.din(n10906));
	jspl jspl_w_n10907_0(.douta(w_n10907_0[0]),.doutb(w_n10907_0[1]),.din(n10907));
	jspl jspl_w_n10910_0(.douta(w_n10910_0[0]),.doutb(w_n10910_0[1]),.din(n10910));
	jspl jspl_w_n10916_0(.douta(w_n10916_0[0]),.doutb(w_n10916_0[1]),.din(n10916));
	jspl jspl_w_n10917_0(.douta(w_n10917_0[0]),.doutb(w_n10917_0[1]),.din(n10917));
	jspl jspl_w_n10919_0(.douta(w_n10919_0[0]),.doutb(w_n10919_0[1]),.din(n10919));
	jspl jspl_w_n10921_0(.douta(w_n10921_0[0]),.doutb(w_n10921_0[1]),.din(n10921));
	jspl jspl_w_n10923_0(.douta(w_n10923_0[0]),.doutb(w_n10923_0[1]),.din(n10923));
	jspl jspl_w_n10929_0(.douta(w_n10929_0[0]),.doutb(w_n10929_0[1]),.din(n10929));
	jspl jspl_w_n10931_0(.douta(w_n10931_0[0]),.doutb(w_n10931_0[1]),.din(n10931));
	jspl3 jspl3_w_n10932_0(.douta(w_n10932_0[0]),.doutb(w_n10932_0[1]),.doutc(w_n10932_0[2]),.din(n10932));
	jspl jspl_w_n10935_0(.douta(w_n10935_0[0]),.doutb(w_n10935_0[1]),.din(n10935));
	jspl jspl_w_n10936_0(.douta(w_n10936_0[0]),.doutb(w_n10936_0[1]),.din(n10936));
	jspl3 jspl3_w_n10937_0(.douta(w_n10937_0[0]),.doutb(w_n10937_0[1]),.doutc(w_n10937_0[2]),.din(n10937));
	jspl jspl_w_n10939_0(.douta(w_n10939_0[0]),.doutb(w_n10939_0[1]),.din(n10939));
	jspl jspl_w_n10941_0(.douta(w_n10941_0[0]),.doutb(w_n10941_0[1]),.din(n10941));
	jspl jspl_w_n10943_0(.douta(w_n10943_0[0]),.doutb(w_n10943_0[1]),.din(n10943));
	jspl jspl_w_n10949_0(.douta(w_n10949_0[0]),.doutb(w_n10949_0[1]),.din(n10949));
	jspl3 jspl3_w_n10951_0(.douta(w_n10951_0[0]),.doutb(w_n10951_0[1]),.doutc(w_n10951_0[2]),.din(n10951));
	jspl jspl_w_n10952_0(.douta(w_n10952_0[0]),.doutb(w_n10952_0[1]),.din(n10952));
	jspl jspl_w_n10954_0(.douta(w_n10954_0[0]),.doutb(w_n10954_0[1]),.din(n10954));
	jspl jspl_w_n10956_0(.douta(w_n10956_0[0]),.doutb(w_n10956_0[1]),.din(n10956));
	jspl jspl_w_n10960_0(.douta(w_n10960_0[0]),.doutb(w_n10960_0[1]),.din(n10960));
	jspl jspl_w_n10962_0(.douta(w_n10962_0[0]),.doutb(w_n10962_0[1]),.din(n10962));
	jspl jspl_w_n10963_0(.douta(w_n10963_0[0]),.doutb(w_n10963_0[1]),.din(n10963));
	jspl jspl_w_n10964_0(.douta(w_n10964_0[0]),.doutb(w_n10964_0[1]),.din(n10964));
	jspl3 jspl3_w_n10965_0(.douta(w_n10965_0[0]),.doutb(w_n10965_0[1]),.doutc(w_n10965_0[2]),.din(n10965));
	jspl jspl_w_n10968_0(.douta(w_n10968_0[0]),.doutb(w_n10968_0[1]),.din(n10968));
	jspl jspl_w_n10969_0(.douta(w_n10969_0[0]),.doutb(w_n10969_0[1]),.din(n10969));
	jspl3 jspl3_w_n10970_0(.douta(w_n10970_0[0]),.doutb(w_n10970_0[1]),.doutc(w_n10970_0[2]),.din(n10970));
	jspl jspl_w_n10972_0(.douta(w_n10972_0[0]),.doutb(w_n10972_0[1]),.din(n10972));
	jspl jspl_w_n10976_0(.douta(w_n10976_0[0]),.doutb(w_n10976_0[1]),.din(n10976));
	jspl jspl_w_n10978_0(.douta(w_n10978_0[0]),.doutb(w_n10978_0[1]),.din(n10978));
	jspl jspl_w_n10979_0(.douta(w_n10979_0[0]),.doutb(w_n10979_0[1]),.din(n10979));
	jspl3 jspl3_w_n10980_0(.douta(w_n10980_0[0]),.doutb(w_n10980_0[1]),.doutc(w_n10980_0[2]),.din(n10980));
	jspl jspl_w_n10981_0(.douta(w_n10981_0[0]),.doutb(w_n10981_0[1]),.din(n10981));
	jspl jspl_w_n10984_0(.douta(w_n10984_0[0]),.doutb(w_n10984_0[1]),.din(n10984));
	jspl jspl_w_n10990_0(.douta(w_n10990_0[0]),.doutb(w_n10990_0[1]),.din(n10990));
	jspl jspl_w_n10991_0(.douta(w_n10991_0[0]),.doutb(w_n10991_0[1]),.din(n10991));
	jspl jspl_w_n10993_0(.douta(w_n10993_0[0]),.doutb(w_n10993_0[1]),.din(n10993));
	jspl jspl_w_n10995_0(.douta(w_n10995_0[0]),.doutb(w_n10995_0[1]),.din(n10995));
	jspl jspl_w_n10997_0(.douta(w_n10997_0[0]),.doutb(w_n10997_0[1]),.din(n10997));
	jspl jspl_w_n11003_0(.douta(w_n11003_0[0]),.doutb(w_n11003_0[1]),.din(n11003));
	jspl jspl_w_n11005_0(.douta(w_n11005_0[0]),.doutb(w_n11005_0[1]),.din(n11005));
	jspl3 jspl3_w_n11006_0(.douta(w_n11006_0[0]),.doutb(w_n11006_0[1]),.doutc(w_n11006_0[2]),.din(n11006));
	jspl jspl_w_n11009_0(.douta(w_n11009_0[0]),.doutb(w_n11009_0[1]),.din(n11009));
	jspl jspl_w_n11010_0(.douta(w_n11010_0[0]),.doutb(w_n11010_0[1]),.din(n11010));
	jspl3 jspl3_w_n11011_0(.douta(w_n11011_0[0]),.doutb(w_n11011_0[1]),.doutc(w_n11011_0[2]),.din(n11011));
	jspl jspl_w_n11013_0(.douta(w_n11013_0[0]),.doutb(w_n11013_0[1]),.din(n11013));
	jspl jspl_w_n11017_0(.douta(w_n11017_0[0]),.doutb(w_n11017_0[1]),.din(n11017));
	jspl jspl_w_n11019_0(.douta(w_n11019_0[0]),.doutb(w_n11019_0[1]),.din(n11019));
	jspl jspl_w_n11020_0(.douta(w_n11020_0[0]),.doutb(w_n11020_0[1]),.din(n11020));
	jspl3 jspl3_w_n11021_0(.douta(w_n11021_0[0]),.doutb(w_n11021_0[1]),.doutc(w_n11021_0[2]),.din(n11021));
	jspl jspl_w_n11022_0(.douta(w_n11022_0[0]),.doutb(w_n11022_0[1]),.din(n11022));
	jspl jspl_w_n11025_0(.douta(w_n11025_0[0]),.doutb(w_n11025_0[1]),.din(n11025));
	jspl jspl_w_n11031_0(.douta(w_n11031_0[0]),.doutb(w_n11031_0[1]),.din(n11031));
	jspl jspl_w_n11032_0(.douta(w_n11032_0[0]),.doutb(w_n11032_0[1]),.din(n11032));
	jspl jspl_w_n11034_0(.douta(w_n11034_0[0]),.doutb(w_n11034_0[1]),.din(n11034));
	jspl jspl_w_n11036_0(.douta(w_n11036_0[0]),.doutb(w_n11036_0[1]),.din(n11036));
	jspl jspl_w_n11038_0(.douta(w_n11038_0[0]),.doutb(w_n11038_0[1]),.din(n11038));
	jspl jspl_w_n11044_0(.douta(w_n11044_0[0]),.doutb(w_n11044_0[1]),.din(n11044));
	jspl jspl_w_n11046_0(.douta(w_n11046_0[0]),.doutb(w_n11046_0[1]),.din(n11046));
	jspl3 jspl3_w_n11047_0(.douta(w_n11047_0[0]),.doutb(w_n11047_0[1]),.doutc(w_n11047_0[2]),.din(n11047));
	jspl jspl_w_n11050_0(.douta(w_n11050_0[0]),.doutb(w_n11050_0[1]),.din(n11050));
	jspl jspl_w_n11051_0(.douta(w_n11051_0[0]),.doutb(w_n11051_0[1]),.din(n11051));
	jspl3 jspl3_w_n11052_0(.douta(w_n11052_0[0]),.doutb(w_n11052_0[1]),.doutc(w_n11052_0[2]),.din(n11052));
	jspl jspl_w_n11054_0(.douta(w_n11054_0[0]),.doutb(w_n11054_0[1]),.din(n11054));
	jspl jspl_w_n11058_0(.douta(w_n11058_0[0]),.doutb(w_n11058_0[1]),.din(n11058));
	jspl jspl_w_n11060_0(.douta(w_n11060_0[0]),.doutb(w_n11060_0[1]),.din(n11060));
	jspl jspl_w_n11061_0(.douta(w_n11061_0[0]),.doutb(w_n11061_0[1]),.din(n11061));
	jspl3 jspl3_w_n11062_0(.douta(w_n11062_0[0]),.doutb(w_n11062_0[1]),.doutc(w_n11062_0[2]),.din(n11062));
	jspl jspl_w_n11063_0(.douta(w_n11063_0[0]),.doutb(w_n11063_0[1]),.din(n11063));
	jspl jspl_w_n11066_0(.douta(w_n11066_0[0]),.doutb(w_n11066_0[1]),.din(n11066));
	jspl jspl_w_n11072_0(.douta(w_n11072_0[0]),.doutb(w_n11072_0[1]),.din(n11072));
	jspl jspl_w_n11073_0(.douta(w_n11073_0[0]),.doutb(w_n11073_0[1]),.din(n11073));
	jspl jspl_w_n11075_0(.douta(w_n11075_0[0]),.doutb(w_n11075_0[1]),.din(n11075));
	jspl jspl_w_n11077_0(.douta(w_n11077_0[0]),.doutb(w_n11077_0[1]),.din(n11077));
	jspl jspl_w_n11079_0(.douta(w_n11079_0[0]),.doutb(w_n11079_0[1]),.din(n11079));
	jspl jspl_w_n11085_0(.douta(w_n11085_0[0]),.doutb(w_n11085_0[1]),.din(n11085));
	jspl jspl_w_n11087_0(.douta(w_n11087_0[0]),.doutb(w_n11087_0[1]),.din(n11087));
	jspl3 jspl3_w_n11088_0(.douta(w_n11088_0[0]),.doutb(w_n11088_0[1]),.doutc(w_n11088_0[2]),.din(n11088));
	jspl jspl_w_n11091_0(.douta(w_n11091_0[0]),.doutb(w_n11091_0[1]),.din(n11091));
	jspl jspl_w_n11092_0(.douta(w_n11092_0[0]),.doutb(w_n11092_0[1]),.din(n11092));
	jspl3 jspl3_w_n11093_0(.douta(w_n11093_0[0]),.doutb(w_n11093_0[1]),.doutc(w_n11093_0[2]),.din(n11093));
	jspl jspl_w_n11095_0(.douta(w_n11095_0[0]),.doutb(w_n11095_0[1]),.din(n11095));
	jspl jspl_w_n11099_0(.douta(w_n11099_0[0]),.doutb(w_n11099_0[1]),.din(n11099));
	jspl jspl_w_n11101_0(.douta(w_n11101_0[0]),.doutb(w_n11101_0[1]),.din(n11101));
	jspl jspl_w_n11102_0(.douta(w_n11102_0[0]),.doutb(w_n11102_0[1]),.din(n11102));
	jspl3 jspl3_w_n11103_0(.douta(w_n11103_0[0]),.doutb(w_n11103_0[1]),.doutc(w_n11103_0[2]),.din(n11103));
	jspl jspl_w_n11104_0(.douta(w_n11104_0[0]),.doutb(w_n11104_0[1]),.din(n11104));
	jspl jspl_w_n11107_0(.douta(w_n11107_0[0]),.doutb(w_n11107_0[1]),.din(n11107));
	jspl jspl_w_n11113_0(.douta(w_n11113_0[0]),.doutb(w_n11113_0[1]),.din(n11113));
	jspl jspl_w_n11114_0(.douta(w_n11114_0[0]),.doutb(w_n11114_0[1]),.din(n11114));
	jspl jspl_w_n11116_0(.douta(w_n11116_0[0]),.doutb(w_n11116_0[1]),.din(n11116));
	jspl jspl_w_n11118_0(.douta(w_n11118_0[0]),.doutb(w_n11118_0[1]),.din(n11118));
	jspl jspl_w_n11120_0(.douta(w_n11120_0[0]),.doutb(w_n11120_0[1]),.din(n11120));
	jspl jspl_w_n11126_0(.douta(w_n11126_0[0]),.doutb(w_n11126_0[1]),.din(n11126));
	jspl3 jspl3_w_n11128_0(.douta(w_n11128_0[0]),.doutb(w_n11128_0[1]),.doutc(w_n11128_0[2]),.din(n11128));
	jspl jspl_w_n11133_0(.douta(w_n11133_0[0]),.doutb(w_n11133_0[1]),.din(n11133));
	jspl3 jspl3_w_n11135_0(.douta(w_n11135_0[0]),.doutb(w_n11135_0[1]),.doutc(w_n11135_0[2]),.din(n11135));
	jspl3 jspl3_w_n11139_0(.douta(w_n11139_0[0]),.doutb(w_n11139_0[1]),.doutc(w_n11139_0[2]),.din(n11139));
	jspl jspl_w_n11140_0(.douta(w_n11140_0[0]),.doutb(w_n11140_0[1]),.din(n11140));
	jspl jspl_w_n11145_0(.douta(w_n11145_0[0]),.doutb(w_n11145_0[1]),.din(n11145));
	jspl3 jspl3_w_n11146_0(.douta(w_n11146_0[0]),.doutb(w_n11146_0[1]),.doutc(w_n11146_0[2]),.din(n11146));
	jspl jspl_w_n11151_0(.douta(w_n11151_0[0]),.doutb(w_n11151_0[1]),.din(n11151));
	jspl jspl_w_n11158_0(.douta(w_n11158_0[0]),.doutb(w_n11158_0[1]),.din(n11158));
	jspl3 jspl3_w_n11160_0(.douta(w_n11160_0[0]),.doutb(w_n11160_0[1]),.doutc(w_n11160_0[2]),.din(n11160));
	jspl jspl_w_n11160_1(.douta(w_n11160_1[0]),.doutb(w_n11160_1[1]),.din(w_n11160_0[0]));
	jspl jspl_w_n11161_0(.douta(w_n11161_0[0]),.doutb(w_n11161_0[1]),.din(n11161));
	jspl3 jspl3_w_n11164_0(.douta(w_n11164_0[0]),.doutb(w_n11164_0[1]),.doutc(w_n11164_0[2]),.din(n11164));
	jspl jspl_w_n11165_0(.douta(w_n11165_0[0]),.doutb(w_n11165_0[1]),.din(n11165));
	jspl jspl_w_n11166_0(.douta(w_n11166_0[0]),.doutb(w_n11166_0[1]),.din(n11166));
	jspl jspl_w_n11167_0(.douta(w_n11167_0[0]),.doutb(w_n11167_0[1]),.din(n11167));
	jspl jspl_w_n11169_0(.douta(w_n11169_0[0]),.doutb(w_n11169_0[1]),.din(n11169));
	jspl jspl_w_n11171_0(.douta(w_n11171_0[0]),.doutb(w_n11171_0[1]),.din(n11171));
	jspl jspl_w_n11173_0(.douta(w_n11173_0[0]),.doutb(w_n11173_0[1]),.din(n11173));
	jspl jspl_w_n11182_0(.douta(w_n11182_0[0]),.doutb(w_n11182_0[1]),.din(n11182));
	jspl3 jspl3_w_n11184_0(.douta(w_n11184_0[0]),.doutb(w_n11184_0[1]),.doutc(w_n11184_0[2]),.din(n11184));
	jspl jspl_w_n11185_0(.douta(w_n11185_0[0]),.doutb(w_n11185_0[1]),.din(n11185));
	jspl jspl_w_n11189_0(.douta(w_n11189_0[0]),.doutb(w_n11189_0[1]),.din(n11189));
	jspl jspl_w_n11191_0(.douta(w_n11191_0[0]),.doutb(w_n11191_0[1]),.din(n11191));
	jspl jspl_w_n11193_0(.douta(w_n11193_0[0]),.doutb(w_n11193_0[1]),.din(n11193));
	jspl jspl_w_n11198_0(.douta(w_n11198_0[0]),.doutb(w_n11198_0[1]),.din(n11198));
	jspl jspl_w_n11200_0(.douta(w_n11200_0[0]),.doutb(w_n11200_0[1]),.din(n11200));
	jspl jspl_w_n11201_0(.douta(w_n11201_0[0]),.doutb(w_n11201_0[1]),.din(n11201));
	jspl3 jspl3_w_n11202_0(.douta(w_n11202_0[0]),.doutb(w_n11202_0[1]),.doutc(w_n11202_0[2]),.din(n11202));
	jspl jspl_w_n11203_0(.douta(w_n11203_0[0]),.doutb(w_n11203_0[1]),.din(n11203));
	jspl jspl_w_n11208_0(.douta(w_n11208_0[0]),.doutb(w_n11208_0[1]),.din(n11208));
	jspl jspl_w_n11209_0(.douta(w_n11209_0[0]),.doutb(w_n11209_0[1]),.din(n11209));
	jspl jspl_w_n11211_0(.douta(w_n11211_0[0]),.doutb(w_n11211_0[1]),.din(n11211));
	jspl jspl_w_n11213_0(.douta(w_n11213_0[0]),.doutb(w_n11213_0[1]),.din(n11213));
	jspl jspl_w_n11216_0(.douta(w_n11216_0[0]),.doutb(w_n11216_0[1]),.din(n11216));
	jspl jspl_w_n11222_0(.douta(w_n11222_0[0]),.doutb(w_n11222_0[1]),.din(n11222));
	jspl3 jspl3_w_n11224_0(.douta(w_n11224_0[0]),.doutb(w_n11224_0[1]),.doutc(w_n11224_0[2]),.din(n11224));
	jspl jspl_w_n11225_0(.douta(w_n11225_0[0]),.doutb(w_n11225_0[1]),.din(n11225));
	jspl jspl_w_n11229_0(.douta(w_n11229_0[0]),.doutb(w_n11229_0[1]),.din(n11229));
	jspl jspl_w_n11230_0(.douta(w_n11230_0[0]),.doutb(w_n11230_0[1]),.din(n11230));
	jspl jspl_w_n11232_0(.douta(w_n11232_0[0]),.doutb(w_n11232_0[1]),.din(n11232));
	jspl jspl_w_n11237_0(.douta(w_n11237_0[0]),.doutb(w_n11237_0[1]),.din(n11237));
	jspl jspl_w_n11239_0(.douta(w_n11239_0[0]),.doutb(w_n11239_0[1]),.din(n11239));
	jspl jspl_w_n11240_0(.douta(w_n11240_0[0]),.doutb(w_n11240_0[1]),.din(n11240));
	jspl3 jspl3_w_n11241_0(.douta(w_n11241_0[0]),.doutb(w_n11241_0[1]),.doutc(w_n11241_0[2]),.din(n11241));
	jspl jspl_w_n11242_0(.douta(w_n11242_0[0]),.doutb(w_n11242_0[1]),.din(n11242));
	jspl jspl_w_n11246_0(.douta(w_n11246_0[0]),.doutb(w_n11246_0[1]),.din(n11246));
	jspl jspl_w_n11247_0(.douta(w_n11247_0[0]),.doutb(w_n11247_0[1]),.din(n11247));
	jspl jspl_w_n11249_0(.douta(w_n11249_0[0]),.doutb(w_n11249_0[1]),.din(n11249));
	jspl jspl_w_n11251_0(.douta(w_n11251_0[0]),.doutb(w_n11251_0[1]),.din(n11251));
	jspl jspl_w_n11254_0(.douta(w_n11254_0[0]),.doutb(w_n11254_0[1]),.din(n11254));
	jspl jspl_w_n11260_0(.douta(w_n11260_0[0]),.doutb(w_n11260_0[1]),.din(n11260));
	jspl jspl_w_n11262_0(.douta(w_n11262_0[0]),.doutb(w_n11262_0[1]),.din(n11262));
	jspl3 jspl3_w_n11263_0(.douta(w_n11263_0[0]),.doutb(w_n11263_0[1]),.doutc(w_n11263_0[2]),.din(n11263));
	jspl jspl_w_n11267_0(.douta(w_n11267_0[0]),.doutb(w_n11267_0[1]),.din(n11267));
	jspl jspl_w_n11268_0(.douta(w_n11268_0[0]),.doutb(w_n11268_0[1]),.din(n11268));
	jspl3 jspl3_w_n11269_0(.douta(w_n11269_0[0]),.doutb(w_n11269_0[1]),.doutc(w_n11269_0[2]),.din(n11269));
	jspl jspl_w_n11271_0(.douta(w_n11271_0[0]),.doutb(w_n11271_0[1]),.din(n11271));
	jspl jspl_w_n11276_0(.douta(w_n11276_0[0]),.doutb(w_n11276_0[1]),.din(n11276));
	jspl jspl_w_n11278_0(.douta(w_n11278_0[0]),.doutb(w_n11278_0[1]),.din(n11278));
	jspl jspl_w_n11279_0(.douta(w_n11279_0[0]),.doutb(w_n11279_0[1]),.din(n11279));
	jspl3 jspl3_w_n11280_0(.douta(w_n11280_0[0]),.doutb(w_n11280_0[1]),.doutc(w_n11280_0[2]),.din(n11280));
	jspl jspl_w_n11281_0(.douta(w_n11281_0[0]),.doutb(w_n11281_0[1]),.din(n11281));
	jspl jspl_w_n11285_0(.douta(w_n11285_0[0]),.doutb(w_n11285_0[1]),.din(n11285));
	jspl jspl_w_n11291_0(.douta(w_n11291_0[0]),.doutb(w_n11291_0[1]),.din(n11291));
	jspl jspl_w_n11292_0(.douta(w_n11292_0[0]),.doutb(w_n11292_0[1]),.din(n11292));
	jspl jspl_w_n11294_0(.douta(w_n11294_0[0]),.doutb(w_n11294_0[1]),.din(n11294));
	jspl jspl_w_n11296_0(.douta(w_n11296_0[0]),.doutb(w_n11296_0[1]),.din(n11296));
	jspl jspl_w_n11299_0(.douta(w_n11299_0[0]),.doutb(w_n11299_0[1]),.din(n11299));
	jspl jspl_w_n11305_0(.douta(w_n11305_0[0]),.doutb(w_n11305_0[1]),.din(n11305));
	jspl jspl_w_n11307_0(.douta(w_n11307_0[0]),.doutb(w_n11307_0[1]),.din(n11307));
	jspl3 jspl3_w_n11308_0(.douta(w_n11308_0[0]),.doutb(w_n11308_0[1]),.doutc(w_n11308_0[2]),.din(n11308));
	jspl jspl_w_n11312_0(.douta(w_n11312_0[0]),.doutb(w_n11312_0[1]),.din(n11312));
	jspl jspl_w_n11313_0(.douta(w_n11313_0[0]),.doutb(w_n11313_0[1]),.din(n11313));
	jspl3 jspl3_w_n11314_0(.douta(w_n11314_0[0]),.doutb(w_n11314_0[1]),.doutc(w_n11314_0[2]),.din(n11314));
	jspl jspl_w_n11316_0(.douta(w_n11316_0[0]),.doutb(w_n11316_0[1]),.din(n11316));
	jspl jspl_w_n11321_0(.douta(w_n11321_0[0]),.doutb(w_n11321_0[1]),.din(n11321));
	jspl jspl_w_n11323_0(.douta(w_n11323_0[0]),.doutb(w_n11323_0[1]),.din(n11323));
	jspl jspl_w_n11324_0(.douta(w_n11324_0[0]),.doutb(w_n11324_0[1]),.din(n11324));
	jspl3 jspl3_w_n11325_0(.douta(w_n11325_0[0]),.doutb(w_n11325_0[1]),.doutc(w_n11325_0[2]),.din(n11325));
	jspl jspl_w_n11326_0(.douta(w_n11326_0[0]),.doutb(w_n11326_0[1]),.din(n11326));
	jspl jspl_w_n11330_0(.douta(w_n11330_0[0]),.doutb(w_n11330_0[1]),.din(n11330));
	jspl jspl_w_n11336_0(.douta(w_n11336_0[0]),.doutb(w_n11336_0[1]),.din(n11336));
	jspl jspl_w_n11337_0(.douta(w_n11337_0[0]),.doutb(w_n11337_0[1]),.din(n11337));
	jspl jspl_w_n11339_0(.douta(w_n11339_0[0]),.doutb(w_n11339_0[1]),.din(n11339));
	jspl jspl_w_n11341_0(.douta(w_n11341_0[0]),.doutb(w_n11341_0[1]),.din(n11341));
	jspl jspl_w_n11344_0(.douta(w_n11344_0[0]),.doutb(w_n11344_0[1]),.din(n11344));
	jspl jspl_w_n11350_0(.douta(w_n11350_0[0]),.doutb(w_n11350_0[1]),.din(n11350));
	jspl jspl_w_n11352_0(.douta(w_n11352_0[0]),.doutb(w_n11352_0[1]),.din(n11352));
	jspl3 jspl3_w_n11353_0(.douta(w_n11353_0[0]),.doutb(w_n11353_0[1]),.doutc(w_n11353_0[2]),.din(n11353));
	jspl jspl_w_n11357_0(.douta(w_n11357_0[0]),.doutb(w_n11357_0[1]),.din(n11357));
	jspl jspl_w_n11358_0(.douta(w_n11358_0[0]),.doutb(w_n11358_0[1]),.din(n11358));
	jspl3 jspl3_w_n11359_0(.douta(w_n11359_0[0]),.doutb(w_n11359_0[1]),.doutc(w_n11359_0[2]),.din(n11359));
	jspl jspl_w_n11361_0(.douta(w_n11361_0[0]),.doutb(w_n11361_0[1]),.din(n11361));
	jspl jspl_w_n11366_0(.douta(w_n11366_0[0]),.doutb(w_n11366_0[1]),.din(n11366));
	jspl jspl_w_n11368_0(.douta(w_n11368_0[0]),.doutb(w_n11368_0[1]),.din(n11368));
	jspl jspl_w_n11369_0(.douta(w_n11369_0[0]),.doutb(w_n11369_0[1]),.din(n11369));
	jspl3 jspl3_w_n11370_0(.douta(w_n11370_0[0]),.doutb(w_n11370_0[1]),.doutc(w_n11370_0[2]),.din(n11370));
	jspl jspl_w_n11371_0(.douta(w_n11371_0[0]),.doutb(w_n11371_0[1]),.din(n11371));
	jspl jspl_w_n11375_0(.douta(w_n11375_0[0]),.doutb(w_n11375_0[1]),.din(n11375));
	jspl jspl_w_n11381_0(.douta(w_n11381_0[0]),.doutb(w_n11381_0[1]),.din(n11381));
	jspl jspl_w_n11382_0(.douta(w_n11382_0[0]),.doutb(w_n11382_0[1]),.din(n11382));
	jspl jspl_w_n11384_0(.douta(w_n11384_0[0]),.doutb(w_n11384_0[1]),.din(n11384));
	jspl jspl_w_n11386_0(.douta(w_n11386_0[0]),.doutb(w_n11386_0[1]),.din(n11386));
	jspl jspl_w_n11389_0(.douta(w_n11389_0[0]),.doutb(w_n11389_0[1]),.din(n11389));
	jspl jspl_w_n11395_0(.douta(w_n11395_0[0]),.doutb(w_n11395_0[1]),.din(n11395));
	jspl jspl_w_n11397_0(.douta(w_n11397_0[0]),.doutb(w_n11397_0[1]),.din(n11397));
	jspl3 jspl3_w_n11398_0(.douta(w_n11398_0[0]),.doutb(w_n11398_0[1]),.doutc(w_n11398_0[2]),.din(n11398));
	jspl jspl_w_n11402_0(.douta(w_n11402_0[0]),.doutb(w_n11402_0[1]),.din(n11402));
	jspl jspl_w_n11403_0(.douta(w_n11403_0[0]),.doutb(w_n11403_0[1]),.din(n11403));
	jspl3 jspl3_w_n11404_0(.douta(w_n11404_0[0]),.doutb(w_n11404_0[1]),.doutc(w_n11404_0[2]),.din(n11404));
	jspl jspl_w_n11406_0(.douta(w_n11406_0[0]),.doutb(w_n11406_0[1]),.din(n11406));
	jspl jspl_w_n11411_0(.douta(w_n11411_0[0]),.doutb(w_n11411_0[1]),.din(n11411));
	jspl jspl_w_n11413_0(.douta(w_n11413_0[0]),.doutb(w_n11413_0[1]),.din(n11413));
	jspl jspl_w_n11414_0(.douta(w_n11414_0[0]),.doutb(w_n11414_0[1]),.din(n11414));
	jspl3 jspl3_w_n11415_0(.douta(w_n11415_0[0]),.doutb(w_n11415_0[1]),.doutc(w_n11415_0[2]),.din(n11415));
	jspl jspl_w_n11416_0(.douta(w_n11416_0[0]),.doutb(w_n11416_0[1]),.din(n11416));
	jspl jspl_w_n11420_0(.douta(w_n11420_0[0]),.doutb(w_n11420_0[1]),.din(n11420));
	jspl jspl_w_n11426_0(.douta(w_n11426_0[0]),.doutb(w_n11426_0[1]),.din(n11426));
	jspl jspl_w_n11427_0(.douta(w_n11427_0[0]),.doutb(w_n11427_0[1]),.din(n11427));
	jspl jspl_w_n11429_0(.douta(w_n11429_0[0]),.doutb(w_n11429_0[1]),.din(n11429));
	jspl jspl_w_n11434_0(.douta(w_n11434_0[0]),.doutb(w_n11434_0[1]),.din(n11434));
	jspl jspl_w_n11436_0(.douta(w_n11436_0[0]),.doutb(w_n11436_0[1]),.din(n11436));
	jspl jspl_w_n11437_0(.douta(w_n11437_0[0]),.doutb(w_n11437_0[1]),.din(n11437));
	jspl3 jspl3_w_n11438_0(.douta(w_n11438_0[0]),.doutb(w_n11438_0[1]),.doutc(w_n11438_0[2]),.din(n11438));
	jspl jspl_w_n11439_0(.douta(w_n11439_0[0]),.doutb(w_n11439_0[1]),.din(n11439));
	jspl jspl_w_n11442_0(.douta(w_n11442_0[0]),.doutb(w_n11442_0[1]),.din(n11442));
	jspl jspl_w_n11444_0(.douta(w_n11444_0[0]),.doutb(w_n11444_0[1]),.din(n11444));
	jspl jspl_w_n11446_0(.douta(w_n11446_0[0]),.doutb(w_n11446_0[1]),.din(n11446));
	jspl jspl_w_n11449_0(.douta(w_n11449_0[0]),.doutb(w_n11449_0[1]),.din(n11449));
	jspl jspl_w_n11455_0(.douta(w_n11455_0[0]),.doutb(w_n11455_0[1]),.din(n11455));
	jspl3 jspl3_w_n11457_0(.douta(w_n11457_0[0]),.doutb(w_n11457_0[1]),.doutc(w_n11457_0[2]),.din(n11457));
	jspl jspl_w_n11458_0(.douta(w_n11458_0[0]),.doutb(w_n11458_0[1]),.din(n11458));
	jspl jspl_w_n11462_0(.douta(w_n11462_0[0]),.doutb(w_n11462_0[1]),.din(n11462));
	jspl jspl_w_n11468_0(.douta(w_n11468_0[0]),.doutb(w_n11468_0[1]),.din(n11468));
	jspl jspl_w_n11469_0(.douta(w_n11469_0[0]),.doutb(w_n11469_0[1]),.din(n11469));
	jspl jspl_w_n11471_0(.douta(w_n11471_0[0]),.doutb(w_n11471_0[1]),.din(n11471));
	jspl jspl_w_n11473_0(.douta(w_n11473_0[0]),.doutb(w_n11473_0[1]),.din(n11473));
	jspl jspl_w_n11476_0(.douta(w_n11476_0[0]),.doutb(w_n11476_0[1]),.din(n11476));
	jspl jspl_w_n11482_0(.douta(w_n11482_0[0]),.doutb(w_n11482_0[1]),.din(n11482));
	jspl jspl_w_n11484_0(.douta(w_n11484_0[0]),.doutb(w_n11484_0[1]),.din(n11484));
	jspl3 jspl3_w_n11485_0(.douta(w_n11485_0[0]),.doutb(w_n11485_0[1]),.doutc(w_n11485_0[2]),.din(n11485));
	jspl jspl_w_n11489_0(.douta(w_n11489_0[0]),.doutb(w_n11489_0[1]),.din(n11489));
	jspl jspl_w_n11490_0(.douta(w_n11490_0[0]),.doutb(w_n11490_0[1]),.din(n11490));
	jspl3 jspl3_w_n11491_0(.douta(w_n11491_0[0]),.doutb(w_n11491_0[1]),.doutc(w_n11491_0[2]),.din(n11491));
	jspl jspl_w_n11493_0(.douta(w_n11493_0[0]),.doutb(w_n11493_0[1]),.din(n11493));
	jspl jspl_w_n11498_0(.douta(w_n11498_0[0]),.doutb(w_n11498_0[1]),.din(n11498));
	jspl jspl_w_n11500_0(.douta(w_n11500_0[0]),.doutb(w_n11500_0[1]),.din(n11500));
	jspl jspl_w_n11501_0(.douta(w_n11501_0[0]),.doutb(w_n11501_0[1]),.din(n11501));
	jspl3 jspl3_w_n11502_0(.douta(w_n11502_0[0]),.doutb(w_n11502_0[1]),.doutc(w_n11502_0[2]),.din(n11502));
	jspl jspl_w_n11503_0(.douta(w_n11503_0[0]),.doutb(w_n11503_0[1]),.din(n11503));
	jspl jspl_w_n11507_0(.douta(w_n11507_0[0]),.doutb(w_n11507_0[1]),.din(n11507));
	jspl jspl_w_n11513_0(.douta(w_n11513_0[0]),.doutb(w_n11513_0[1]),.din(n11513));
	jspl jspl_w_n11514_0(.douta(w_n11514_0[0]),.doutb(w_n11514_0[1]),.din(n11514));
	jspl jspl_w_n11516_0(.douta(w_n11516_0[0]),.doutb(w_n11516_0[1]),.din(n11516));
	jspl jspl_w_n11518_0(.douta(w_n11518_0[0]),.doutb(w_n11518_0[1]),.din(n11518));
	jspl jspl_w_n11521_0(.douta(w_n11521_0[0]),.doutb(w_n11521_0[1]),.din(n11521));
	jspl jspl_w_n11527_0(.douta(w_n11527_0[0]),.doutb(w_n11527_0[1]),.din(n11527));
	jspl jspl_w_n11529_0(.douta(w_n11529_0[0]),.doutb(w_n11529_0[1]),.din(n11529));
	jspl3 jspl3_w_n11530_0(.douta(w_n11530_0[0]),.doutb(w_n11530_0[1]),.doutc(w_n11530_0[2]),.din(n11530));
	jspl jspl_w_n11534_0(.douta(w_n11534_0[0]),.doutb(w_n11534_0[1]),.din(n11534));
	jspl jspl_w_n11535_0(.douta(w_n11535_0[0]),.doutb(w_n11535_0[1]),.din(n11535));
	jspl3 jspl3_w_n11536_0(.douta(w_n11536_0[0]),.doutb(w_n11536_0[1]),.doutc(w_n11536_0[2]),.din(n11536));
	jspl jspl_w_n11538_0(.douta(w_n11538_0[0]),.doutb(w_n11538_0[1]),.din(n11538));
	jspl jspl_w_n11543_0(.douta(w_n11543_0[0]),.doutb(w_n11543_0[1]),.din(n11543));
	jspl jspl_w_n11545_0(.douta(w_n11545_0[0]),.doutb(w_n11545_0[1]),.din(n11545));
	jspl jspl_w_n11546_0(.douta(w_n11546_0[0]),.doutb(w_n11546_0[1]),.din(n11546));
	jspl3 jspl3_w_n11547_0(.douta(w_n11547_0[0]),.doutb(w_n11547_0[1]),.doutc(w_n11547_0[2]),.din(n11547));
	jspl jspl_w_n11548_0(.douta(w_n11548_0[0]),.doutb(w_n11548_0[1]),.din(n11548));
	jspl jspl_w_n11552_0(.douta(w_n11552_0[0]),.doutb(w_n11552_0[1]),.din(n11552));
	jspl jspl_w_n11558_0(.douta(w_n11558_0[0]),.doutb(w_n11558_0[1]),.din(n11558));
	jspl jspl_w_n11559_0(.douta(w_n11559_0[0]),.doutb(w_n11559_0[1]),.din(n11559));
	jspl jspl_w_n11561_0(.douta(w_n11561_0[0]),.doutb(w_n11561_0[1]),.din(n11561));
	jspl jspl_w_n11563_0(.douta(w_n11563_0[0]),.doutb(w_n11563_0[1]),.din(n11563));
	jspl jspl_w_n11566_0(.douta(w_n11566_0[0]),.doutb(w_n11566_0[1]),.din(n11566));
	jspl jspl_w_n11572_0(.douta(w_n11572_0[0]),.doutb(w_n11572_0[1]),.din(n11572));
	jspl jspl_w_n11574_0(.douta(w_n11574_0[0]),.doutb(w_n11574_0[1]),.din(n11574));
	jspl3 jspl3_w_n11575_0(.douta(w_n11575_0[0]),.doutb(w_n11575_0[1]),.doutc(w_n11575_0[2]),.din(n11575));
	jspl jspl_w_n11579_0(.douta(w_n11579_0[0]),.doutb(w_n11579_0[1]),.din(n11579));
	jspl jspl_w_n11580_0(.douta(w_n11580_0[0]),.doutb(w_n11580_0[1]),.din(n11580));
	jspl3 jspl3_w_n11581_0(.douta(w_n11581_0[0]),.doutb(w_n11581_0[1]),.doutc(w_n11581_0[2]),.din(n11581));
	jspl jspl_w_n11583_0(.douta(w_n11583_0[0]),.doutb(w_n11583_0[1]),.din(n11583));
	jspl jspl_w_n11588_0(.douta(w_n11588_0[0]),.doutb(w_n11588_0[1]),.din(n11588));
	jspl jspl_w_n11590_0(.douta(w_n11590_0[0]),.doutb(w_n11590_0[1]),.din(n11590));
	jspl jspl_w_n11591_0(.douta(w_n11591_0[0]),.doutb(w_n11591_0[1]),.din(n11591));
	jspl3 jspl3_w_n11592_0(.douta(w_n11592_0[0]),.doutb(w_n11592_0[1]),.doutc(w_n11592_0[2]),.din(n11592));
	jspl jspl_w_n11593_0(.douta(w_n11593_0[0]),.doutb(w_n11593_0[1]),.din(n11593));
	jspl jspl_w_n11597_0(.douta(w_n11597_0[0]),.doutb(w_n11597_0[1]),.din(n11597));
	jspl jspl_w_n11603_0(.douta(w_n11603_0[0]),.doutb(w_n11603_0[1]),.din(n11603));
	jspl jspl_w_n11604_0(.douta(w_n11604_0[0]),.doutb(w_n11604_0[1]),.din(n11604));
	jspl jspl_w_n11606_0(.douta(w_n11606_0[0]),.doutb(w_n11606_0[1]),.din(n11606));
	jspl jspl_w_n11608_0(.douta(w_n11608_0[0]),.doutb(w_n11608_0[1]),.din(n11608));
	jspl jspl_w_n11611_0(.douta(w_n11611_0[0]),.doutb(w_n11611_0[1]),.din(n11611));
	jspl jspl_w_n11617_0(.douta(w_n11617_0[0]),.doutb(w_n11617_0[1]),.din(n11617));
	jspl jspl_w_n11619_0(.douta(w_n11619_0[0]),.doutb(w_n11619_0[1]),.din(n11619));
	jspl3 jspl3_w_n11620_0(.douta(w_n11620_0[0]),.doutb(w_n11620_0[1]),.doutc(w_n11620_0[2]),.din(n11620));
	jspl jspl_w_n11624_0(.douta(w_n11624_0[0]),.doutb(w_n11624_0[1]),.din(n11624));
	jspl jspl_w_n11625_0(.douta(w_n11625_0[0]),.doutb(w_n11625_0[1]),.din(n11625));
	jspl3 jspl3_w_n11626_0(.douta(w_n11626_0[0]),.doutb(w_n11626_0[1]),.doutc(w_n11626_0[2]),.din(n11626));
	jspl jspl_w_n11628_0(.douta(w_n11628_0[0]),.doutb(w_n11628_0[1]),.din(n11628));
	jspl jspl_w_n11633_0(.douta(w_n11633_0[0]),.doutb(w_n11633_0[1]),.din(n11633));
	jspl jspl_w_n11635_0(.douta(w_n11635_0[0]),.doutb(w_n11635_0[1]),.din(n11635));
	jspl jspl_w_n11636_0(.douta(w_n11636_0[0]),.doutb(w_n11636_0[1]),.din(n11636));
	jspl3 jspl3_w_n11637_0(.douta(w_n11637_0[0]),.doutb(w_n11637_0[1]),.doutc(w_n11637_0[2]),.din(n11637));
	jspl3 jspl3_w_n11637_1(.douta(w_n11637_1[0]),.doutb(w_n11637_1[1]),.doutc(w_n11637_1[2]),.din(w_n11637_0[0]));
	jspl jspl_w_n11640_0(.douta(w_n11640_0[0]),.doutb(w_n11640_0[1]),.din(n11640));
	jspl3 jspl3_w_n11641_0(.douta(w_n11641_0[0]),.doutb(w_n11641_0[1]),.doutc(w_n11641_0[2]),.din(n11641));
	jspl jspl_w_n11642_0(.douta(w_n11642_0[0]),.doutb(w_n11642_0[1]),.din(n11642));
	jspl jspl_w_n11643_0(.douta(w_n11643_0[0]),.doutb(w_n11643_0[1]),.din(n11643));
	jspl jspl_w_n11649_0(.douta(w_n11649_0[0]),.doutb(w_n11649_0[1]),.din(n11649));
	jspl3 jspl3_w_n11650_0(.douta(w_n11650_0[0]),.doutb(w_n11650_0[1]),.doutc(w_n11650_0[2]),.din(n11650));
	jspl jspl_w_n11651_0(.douta(w_n11651_0[0]),.doutb(w_n11651_0[1]),.din(n11651));
	jspl jspl_w_n11656_0(.douta(w_n11656_0[0]),.doutb(w_n11656_0[1]),.din(n11656));
	jspl3 jspl3_w_n11657_0(.douta(w_n11657_0[0]),.doutb(w_n11657_0[1]),.doutc(w_n11657_0[2]),.din(n11657));
	jspl3 jspl3_w_n11657_1(.douta(w_n11657_1[0]),.doutb(w_n11657_1[1]),.doutc(w_n11657_1[2]),.din(w_n11657_0[0]));
	jspl3 jspl3_w_n11657_2(.douta(w_n11657_2[0]),.doutb(w_n11657_2[1]),.doutc(w_n11657_2[2]),.din(w_n11657_0[1]));
	jspl3 jspl3_w_n11657_3(.douta(w_n11657_3[0]),.doutb(w_n11657_3[1]),.doutc(w_n11657_3[2]),.din(w_n11657_0[2]));
	jspl3 jspl3_w_n11657_4(.douta(w_n11657_4[0]),.doutb(w_n11657_4[1]),.doutc(w_n11657_4[2]),.din(w_n11657_1[0]));
	jspl3 jspl3_w_n11657_5(.douta(w_n11657_5[0]),.doutb(w_n11657_5[1]),.doutc(w_n11657_5[2]),.din(w_n11657_1[1]));
	jspl3 jspl3_w_n11657_6(.douta(w_n11657_6[0]),.doutb(w_n11657_6[1]),.doutc(w_n11657_6[2]),.din(w_n11657_1[2]));
	jspl3 jspl3_w_n11657_7(.douta(w_n11657_7[0]),.doutb(w_n11657_7[1]),.doutc(w_n11657_7[2]),.din(w_n11657_2[0]));
	jspl3 jspl3_w_n11657_8(.douta(w_n11657_8[0]),.doutb(w_n11657_8[1]),.doutc(w_n11657_8[2]),.din(w_n11657_2[1]));
	jspl3 jspl3_w_n11657_9(.douta(w_n11657_9[0]),.doutb(w_n11657_9[1]),.doutc(w_n11657_9[2]),.din(w_n11657_2[2]));
	jspl3 jspl3_w_n11657_10(.douta(w_n11657_10[0]),.doutb(w_n11657_10[1]),.doutc(w_n11657_10[2]),.din(w_n11657_3[0]));
	jspl3 jspl3_w_n11657_11(.douta(w_n11657_11[0]),.doutb(w_n11657_11[1]),.doutc(w_n11657_11[2]),.din(w_n11657_3[1]));
	jspl3 jspl3_w_n11662_0(.douta(w_n11662_0[0]),.doutb(w_n11662_0[1]),.doutc(w_n11662_0[2]),.din(n11662));
	jspl3 jspl3_w_n11662_1(.douta(w_n11662_1[0]),.doutb(w_n11662_1[1]),.doutc(w_n11662_1[2]),.din(w_n11662_0[0]));
	jspl3 jspl3_w_n11662_2(.douta(w_n11662_2[0]),.doutb(w_n11662_2[1]),.doutc(w_n11662_2[2]),.din(w_n11662_0[1]));
	jspl3 jspl3_w_n11662_3(.douta(w_n11662_3[0]),.doutb(w_n11662_3[1]),.doutc(w_n11662_3[2]),.din(w_n11662_0[2]));
	jspl3 jspl3_w_n11662_4(.douta(w_n11662_4[0]),.doutb(w_n11662_4[1]),.doutc(w_n11662_4[2]),.din(w_n11662_1[0]));
	jspl3 jspl3_w_n11662_5(.douta(w_n11662_5[0]),.doutb(w_n11662_5[1]),.doutc(w_n11662_5[2]),.din(w_n11662_1[1]));
	jspl3 jspl3_w_n11662_6(.douta(w_n11662_6[0]),.doutb(w_n11662_6[1]),.doutc(w_n11662_6[2]),.din(w_n11662_1[2]));
	jspl3 jspl3_w_n11662_7(.douta(w_n11662_7[0]),.doutb(w_n11662_7[1]),.doutc(w_n11662_7[2]),.din(w_n11662_2[0]));
	jspl3 jspl3_w_n11662_8(.douta(w_n11662_8[0]),.doutb(w_n11662_8[1]),.doutc(w_n11662_8[2]),.din(w_n11662_2[1]));
	jspl3 jspl3_w_n11662_9(.douta(w_n11662_9[0]),.doutb(w_n11662_9[1]),.doutc(w_n11662_9[2]),.din(w_n11662_2[2]));
	jspl3 jspl3_w_n11662_10(.douta(w_n11662_10[0]),.doutb(w_n11662_10[1]),.doutc(w_n11662_10[2]),.din(w_n11662_3[0]));
	jspl3 jspl3_w_n11662_11(.douta(w_n11662_11[0]),.doutb(w_n11662_11[1]),.doutc(w_n11662_11[2]),.din(w_n11662_3[1]));
	jspl3 jspl3_w_n11662_12(.douta(w_n11662_12[0]),.doutb(w_n11662_12[1]),.doutc(w_n11662_12[2]),.din(w_n11662_3[2]));
	jspl3 jspl3_w_n11662_13(.douta(w_n11662_13[0]),.doutb(w_n11662_13[1]),.doutc(w_n11662_13[2]),.din(w_n11662_4[0]));
	jspl3 jspl3_w_n11662_14(.douta(w_n11662_14[0]),.doutb(w_n11662_14[1]),.doutc(w_n11662_14[2]),.din(w_n11662_4[1]));
	jspl3 jspl3_w_n11662_15(.douta(w_n11662_15[0]),.doutb(w_n11662_15[1]),.doutc(w_n11662_15[2]),.din(w_n11662_4[2]));
	jspl3 jspl3_w_n11662_16(.douta(w_n11662_16[0]),.doutb(w_n11662_16[1]),.doutc(w_n11662_16[2]),.din(w_n11662_5[0]));
	jspl3 jspl3_w_n11662_17(.douta(w_n11662_17[0]),.doutb(w_n11662_17[1]),.doutc(w_n11662_17[2]),.din(w_n11662_5[1]));
	jspl3 jspl3_w_n11662_18(.douta(w_n11662_18[0]),.doutb(w_n11662_18[1]),.doutc(w_n11662_18[2]),.din(w_n11662_5[2]));
	jspl3 jspl3_w_n11662_19(.douta(w_n11662_19[0]),.doutb(w_n11662_19[1]),.doutc(w_n11662_19[2]),.din(w_n11662_6[0]));
	jspl3 jspl3_w_n11662_20(.douta(w_n11662_20[0]),.doutb(w_n11662_20[1]),.doutc(w_n11662_20[2]),.din(w_n11662_6[1]));
	jspl3 jspl3_w_n11662_21(.douta(w_n11662_21[0]),.doutb(w_n11662_21[1]),.doutc(w_n11662_21[2]),.din(w_n11662_6[2]));
	jspl3 jspl3_w_n11662_22(.douta(w_n11662_22[0]),.doutb(w_n11662_22[1]),.doutc(w_n11662_22[2]),.din(w_n11662_7[0]));
	jspl3 jspl3_w_n11662_23(.douta(w_n11662_23[0]),.doutb(w_n11662_23[1]),.doutc(w_n11662_23[2]),.din(w_n11662_7[1]));
	jspl jspl_w_n11662_24(.douta(w_n11662_24[0]),.doutb(w_n11662_24[1]),.din(w_n11662_7[2]));
	jspl jspl_w_n11665_0(.douta(w_n11665_0[0]),.doutb(w_n11665_0[1]),.din(n11665));
	jspl3 jspl3_w_n11667_0(.douta(w_n11667_0[0]),.doutb(w_n11667_0[1]),.doutc(w_n11667_0[2]),.din(n11667));
	jspl jspl_w_n11667_1(.douta(w_n11667_1[0]),.doutb(w_n11667_1[1]),.din(w_n11667_0[0]));
	jspl3 jspl3_w_n11668_0(.douta(w_n11668_0[0]),.doutb(w_n11668_0[1]),.doutc(w_n11668_0[2]),.din(n11668));
	jspl3 jspl3_w_n11672_0(.douta(w_n11672_0[0]),.doutb(w_n11672_0[1]),.doutc(w_n11672_0[2]),.din(n11672));
	jspl jspl_w_n11673_0(.douta(w_n11673_0[0]),.doutb(w_n11673_0[1]),.din(n11673));
	jspl jspl_w_n11674_0(.douta(w_n11674_0[0]),.doutb(w_n11674_0[1]),.din(n11674));
	jspl jspl_w_n11675_0(.douta(w_n11675_0[0]),.doutb(w_n11675_0[1]),.din(n11675));
	jspl jspl_w_n11677_0(.douta(w_n11677_0[0]),.doutb(w_n11677_0[1]),.din(n11677));
	jspl jspl_w_n11679_0(.douta(w_n11679_0[0]),.doutb(w_n11679_0[1]),.din(n11679));
	jspl jspl_w_n11681_0(.douta(w_n11681_0[0]),.doutb(w_n11681_0[1]),.din(n11681));
	jspl jspl_w_n11684_0(.douta(w_n11684_0[0]),.doutb(w_n11684_0[1]),.din(n11684));
	jspl jspl_w_n11689_0(.douta(w_n11689_0[0]),.doutb(w_n11689_0[1]),.din(n11689));
	jspl3 jspl3_w_n11691_0(.douta(w_n11691_0[0]),.doutb(w_n11691_0[1]),.doutc(w_n11691_0[2]),.din(n11691));
	jspl jspl_w_n11692_0(.douta(w_n11692_0[0]),.doutb(w_n11692_0[1]),.din(n11692));
	jspl jspl_w_n11696_0(.douta(w_n11696_0[0]),.doutb(w_n11696_0[1]),.din(n11696));
	jspl jspl_w_n11697_0(.douta(w_n11697_0[0]),.doutb(w_n11697_0[1]),.din(n11697));
	jspl jspl_w_n11699_0(.douta(w_n11699_0[0]),.doutb(w_n11699_0[1]),.din(n11699));
	jspl jspl_w_n11703_0(.douta(w_n11703_0[0]),.doutb(w_n11703_0[1]),.din(n11703));
	jspl jspl_w_n11705_0(.douta(w_n11705_0[0]),.doutb(w_n11705_0[1]),.din(n11705));
	jspl jspl_w_n11706_0(.douta(w_n11706_0[0]),.doutb(w_n11706_0[1]),.din(n11706));
	jspl3 jspl3_w_n11707_0(.douta(w_n11707_0[0]),.doutb(w_n11707_0[1]),.doutc(w_n11707_0[2]),.din(n11707));
	jspl jspl_w_n11708_0(.douta(w_n11708_0[0]),.doutb(w_n11708_0[1]),.din(n11708));
	jspl jspl_w_n11712_0(.douta(w_n11712_0[0]),.doutb(w_n11712_0[1]),.din(n11712));
	jspl jspl_w_n11714_0(.douta(w_n11714_0[0]),.doutb(w_n11714_0[1]),.din(n11714));
	jspl jspl_w_n11716_0(.douta(w_n11716_0[0]),.doutb(w_n11716_0[1]),.din(n11716));
	jspl jspl_w_n11718_0(.douta(w_n11718_0[0]),.doutb(w_n11718_0[1]),.din(n11718));
	jspl jspl_w_n11721_0(.douta(w_n11721_0[0]),.doutb(w_n11721_0[1]),.din(n11721));
	jspl jspl_w_n11727_0(.douta(w_n11727_0[0]),.doutb(w_n11727_0[1]),.din(n11727));
	jspl3 jspl3_w_n11729_0(.douta(w_n11729_0[0]),.doutb(w_n11729_0[1]),.doutc(w_n11729_0[2]),.din(n11729));
	jspl jspl_w_n11730_0(.douta(w_n11730_0[0]),.doutb(w_n11730_0[1]),.din(n11730));
	jspl jspl_w_n11735_0(.douta(w_n11735_0[0]),.doutb(w_n11735_0[1]),.din(n11735));
	jspl jspl_w_n11737_0(.douta(w_n11737_0[0]),.doutb(w_n11737_0[1]),.din(n11737));
	jspl jspl_w_n11739_0(.douta(w_n11739_0[0]),.doutb(w_n11739_0[1]),.din(n11739));
	jspl jspl_w_n11743_0(.douta(w_n11743_0[0]),.doutb(w_n11743_0[1]),.din(n11743));
	jspl jspl_w_n11745_0(.douta(w_n11745_0[0]),.doutb(w_n11745_0[1]),.din(n11745));
	jspl jspl_w_n11746_0(.douta(w_n11746_0[0]),.doutb(w_n11746_0[1]),.din(n11746));
	jspl3 jspl3_w_n11747_0(.douta(w_n11747_0[0]),.doutb(w_n11747_0[1]),.doutc(w_n11747_0[2]),.din(n11747));
	jspl jspl_w_n11748_0(.douta(w_n11748_0[0]),.doutb(w_n11748_0[1]),.din(n11748));
	jspl jspl_w_n11754_0(.douta(w_n11754_0[0]),.doutb(w_n11754_0[1]),.din(n11754));
	jspl jspl_w_n11755_0(.douta(w_n11755_0[0]),.doutb(w_n11755_0[1]),.din(n11755));
	jspl jspl_w_n11757_0(.douta(w_n11757_0[0]),.doutb(w_n11757_0[1]),.din(n11757));
	jspl jspl_w_n11759_0(.douta(w_n11759_0[0]),.doutb(w_n11759_0[1]),.din(n11759));
	jspl jspl_w_n11761_0(.douta(w_n11761_0[0]),.doutb(w_n11761_0[1]),.din(n11761));
	jspl jspl_w_n11767_0(.douta(w_n11767_0[0]),.doutb(w_n11767_0[1]),.din(n11767));
	jspl jspl_w_n11769_0(.douta(w_n11769_0[0]),.doutb(w_n11769_0[1]),.din(n11769));
	jspl3 jspl3_w_n11770_0(.douta(w_n11770_0[0]),.doutb(w_n11770_0[1]),.doutc(w_n11770_0[2]),.din(n11770));
	jspl jspl_w_n11773_0(.douta(w_n11773_0[0]),.doutb(w_n11773_0[1]),.din(n11773));
	jspl jspl_w_n11774_0(.douta(w_n11774_0[0]),.doutb(w_n11774_0[1]),.din(n11774));
	jspl3 jspl3_w_n11775_0(.douta(w_n11775_0[0]),.doutb(w_n11775_0[1]),.doutc(w_n11775_0[2]),.din(n11775));
	jspl jspl_w_n11777_0(.douta(w_n11777_0[0]),.doutb(w_n11777_0[1]),.din(n11777));
	jspl jspl_w_n11781_0(.douta(w_n11781_0[0]),.doutb(w_n11781_0[1]),.din(n11781));
	jspl jspl_w_n11783_0(.douta(w_n11783_0[0]),.doutb(w_n11783_0[1]),.din(n11783));
	jspl jspl_w_n11784_0(.douta(w_n11784_0[0]),.doutb(w_n11784_0[1]),.din(n11784));
	jspl3 jspl3_w_n11785_0(.douta(w_n11785_0[0]),.doutb(w_n11785_0[1]),.doutc(w_n11785_0[2]),.din(n11785));
	jspl jspl_w_n11786_0(.douta(w_n11786_0[0]),.doutb(w_n11786_0[1]),.din(n11786));
	jspl jspl_w_n11789_0(.douta(w_n11789_0[0]),.doutb(w_n11789_0[1]),.din(n11789));
	jspl jspl_w_n11795_0(.douta(w_n11795_0[0]),.doutb(w_n11795_0[1]),.din(n11795));
	jspl jspl_w_n11796_0(.douta(w_n11796_0[0]),.doutb(w_n11796_0[1]),.din(n11796));
	jspl jspl_w_n11798_0(.douta(w_n11798_0[0]),.doutb(w_n11798_0[1]),.din(n11798));
	jspl jspl_w_n11800_0(.douta(w_n11800_0[0]),.doutb(w_n11800_0[1]),.din(n11800));
	jspl jspl_w_n11802_0(.douta(w_n11802_0[0]),.doutb(w_n11802_0[1]),.din(n11802));
	jspl jspl_w_n11808_0(.douta(w_n11808_0[0]),.doutb(w_n11808_0[1]),.din(n11808));
	jspl jspl_w_n11810_0(.douta(w_n11810_0[0]),.doutb(w_n11810_0[1]),.din(n11810));
	jspl3 jspl3_w_n11811_0(.douta(w_n11811_0[0]),.doutb(w_n11811_0[1]),.doutc(w_n11811_0[2]),.din(n11811));
	jspl jspl_w_n11814_0(.douta(w_n11814_0[0]),.doutb(w_n11814_0[1]),.din(n11814));
	jspl jspl_w_n11815_0(.douta(w_n11815_0[0]),.doutb(w_n11815_0[1]),.din(n11815));
	jspl3 jspl3_w_n11816_0(.douta(w_n11816_0[0]),.doutb(w_n11816_0[1]),.doutc(w_n11816_0[2]),.din(n11816));
	jspl jspl_w_n11818_0(.douta(w_n11818_0[0]),.doutb(w_n11818_0[1]),.din(n11818));
	jspl jspl_w_n11822_0(.douta(w_n11822_0[0]),.doutb(w_n11822_0[1]),.din(n11822));
	jspl jspl_w_n11824_0(.douta(w_n11824_0[0]),.doutb(w_n11824_0[1]),.din(n11824));
	jspl jspl_w_n11825_0(.douta(w_n11825_0[0]),.doutb(w_n11825_0[1]),.din(n11825));
	jspl3 jspl3_w_n11826_0(.douta(w_n11826_0[0]),.doutb(w_n11826_0[1]),.doutc(w_n11826_0[2]),.din(n11826));
	jspl jspl_w_n11827_0(.douta(w_n11827_0[0]),.doutb(w_n11827_0[1]),.din(n11827));
	jspl jspl_w_n11830_0(.douta(w_n11830_0[0]),.doutb(w_n11830_0[1]),.din(n11830));
	jspl jspl_w_n11836_0(.douta(w_n11836_0[0]),.doutb(w_n11836_0[1]),.din(n11836));
	jspl jspl_w_n11837_0(.douta(w_n11837_0[0]),.doutb(w_n11837_0[1]),.din(n11837));
	jspl jspl_w_n11839_0(.douta(w_n11839_0[0]),.doutb(w_n11839_0[1]),.din(n11839));
	jspl jspl_w_n11841_0(.douta(w_n11841_0[0]),.doutb(w_n11841_0[1]),.din(n11841));
	jspl jspl_w_n11843_0(.douta(w_n11843_0[0]),.doutb(w_n11843_0[1]),.din(n11843));
	jspl jspl_w_n11849_0(.douta(w_n11849_0[0]),.doutb(w_n11849_0[1]),.din(n11849));
	jspl jspl_w_n11851_0(.douta(w_n11851_0[0]),.doutb(w_n11851_0[1]),.din(n11851));
	jspl3 jspl3_w_n11852_0(.douta(w_n11852_0[0]),.doutb(w_n11852_0[1]),.doutc(w_n11852_0[2]),.din(n11852));
	jspl jspl_w_n11855_0(.douta(w_n11855_0[0]),.doutb(w_n11855_0[1]),.din(n11855));
	jspl jspl_w_n11856_0(.douta(w_n11856_0[0]),.doutb(w_n11856_0[1]),.din(n11856));
	jspl3 jspl3_w_n11857_0(.douta(w_n11857_0[0]),.doutb(w_n11857_0[1]),.doutc(w_n11857_0[2]),.din(n11857));
	jspl jspl_w_n11859_0(.douta(w_n11859_0[0]),.doutb(w_n11859_0[1]),.din(n11859));
	jspl jspl_w_n11863_0(.douta(w_n11863_0[0]),.doutb(w_n11863_0[1]),.din(n11863));
	jspl jspl_w_n11865_0(.douta(w_n11865_0[0]),.doutb(w_n11865_0[1]),.din(n11865));
	jspl jspl_w_n11866_0(.douta(w_n11866_0[0]),.doutb(w_n11866_0[1]),.din(n11866));
	jspl3 jspl3_w_n11867_0(.douta(w_n11867_0[0]),.doutb(w_n11867_0[1]),.doutc(w_n11867_0[2]),.din(n11867));
	jspl jspl_w_n11868_0(.douta(w_n11868_0[0]),.doutb(w_n11868_0[1]),.din(n11868));
	jspl jspl_w_n11871_0(.douta(w_n11871_0[0]),.doutb(w_n11871_0[1]),.din(n11871));
	jspl jspl_w_n11877_0(.douta(w_n11877_0[0]),.doutb(w_n11877_0[1]),.din(n11877));
	jspl jspl_w_n11878_0(.douta(w_n11878_0[0]),.doutb(w_n11878_0[1]),.din(n11878));
	jspl jspl_w_n11880_0(.douta(w_n11880_0[0]),.doutb(w_n11880_0[1]),.din(n11880));
	jspl jspl_w_n11882_0(.douta(w_n11882_0[0]),.doutb(w_n11882_0[1]),.din(n11882));
	jspl jspl_w_n11884_0(.douta(w_n11884_0[0]),.doutb(w_n11884_0[1]),.din(n11884));
	jspl jspl_w_n11890_0(.douta(w_n11890_0[0]),.doutb(w_n11890_0[1]),.din(n11890));
	jspl jspl_w_n11892_0(.douta(w_n11892_0[0]),.doutb(w_n11892_0[1]),.din(n11892));
	jspl3 jspl3_w_n11893_0(.douta(w_n11893_0[0]),.doutb(w_n11893_0[1]),.doutc(w_n11893_0[2]),.din(n11893));
	jspl jspl_w_n11896_0(.douta(w_n11896_0[0]),.doutb(w_n11896_0[1]),.din(n11896));
	jspl jspl_w_n11897_0(.douta(w_n11897_0[0]),.doutb(w_n11897_0[1]),.din(n11897));
	jspl3 jspl3_w_n11898_0(.douta(w_n11898_0[0]),.doutb(w_n11898_0[1]),.doutc(w_n11898_0[2]),.din(n11898));
	jspl jspl_w_n11900_0(.douta(w_n11900_0[0]),.doutb(w_n11900_0[1]),.din(n11900));
	jspl jspl_w_n11904_0(.douta(w_n11904_0[0]),.doutb(w_n11904_0[1]),.din(n11904));
	jspl jspl_w_n11906_0(.douta(w_n11906_0[0]),.doutb(w_n11906_0[1]),.din(n11906));
	jspl jspl_w_n11907_0(.douta(w_n11907_0[0]),.doutb(w_n11907_0[1]),.din(n11907));
	jspl3 jspl3_w_n11908_0(.douta(w_n11908_0[0]),.doutb(w_n11908_0[1]),.doutc(w_n11908_0[2]),.din(n11908));
	jspl jspl_w_n11909_0(.douta(w_n11909_0[0]),.doutb(w_n11909_0[1]),.din(n11909));
	jspl jspl_w_n11912_0(.douta(w_n11912_0[0]),.doutb(w_n11912_0[1]),.din(n11912));
	jspl jspl_w_n11918_0(.douta(w_n11918_0[0]),.doutb(w_n11918_0[1]),.din(n11918));
	jspl jspl_w_n11919_0(.douta(w_n11919_0[0]),.doutb(w_n11919_0[1]),.din(n11919));
	jspl jspl_w_n11921_0(.douta(w_n11921_0[0]),.doutb(w_n11921_0[1]),.din(n11921));
	jspl jspl_w_n11923_0(.douta(w_n11923_0[0]),.doutb(w_n11923_0[1]),.din(n11923));
	jspl jspl_w_n11925_0(.douta(w_n11925_0[0]),.doutb(w_n11925_0[1]),.din(n11925));
	jspl jspl_w_n11931_0(.douta(w_n11931_0[0]),.doutb(w_n11931_0[1]),.din(n11931));
	jspl jspl_w_n11933_0(.douta(w_n11933_0[0]),.doutb(w_n11933_0[1]),.din(n11933));
	jspl3 jspl3_w_n11934_0(.douta(w_n11934_0[0]),.doutb(w_n11934_0[1]),.doutc(w_n11934_0[2]),.din(n11934));
	jspl jspl_w_n11937_0(.douta(w_n11937_0[0]),.doutb(w_n11937_0[1]),.din(n11937));
	jspl jspl_w_n11938_0(.douta(w_n11938_0[0]),.doutb(w_n11938_0[1]),.din(n11938));
	jspl3 jspl3_w_n11939_0(.douta(w_n11939_0[0]),.doutb(w_n11939_0[1]),.doutc(w_n11939_0[2]),.din(n11939));
	jspl jspl_w_n11941_0(.douta(w_n11941_0[0]),.doutb(w_n11941_0[1]),.din(n11941));
	jspl jspl_w_n11943_0(.douta(w_n11943_0[0]),.doutb(w_n11943_0[1]),.din(n11943));
	jspl jspl_w_n11945_0(.douta(w_n11945_0[0]),.doutb(w_n11945_0[1]),.din(n11945));
	jspl jspl_w_n11951_0(.douta(w_n11951_0[0]),.doutb(w_n11951_0[1]),.din(n11951));
	jspl3 jspl3_w_n11953_0(.douta(w_n11953_0[0]),.doutb(w_n11953_0[1]),.doutc(w_n11953_0[2]),.din(n11953));
	jspl jspl_w_n11954_0(.douta(w_n11954_0[0]),.doutb(w_n11954_0[1]),.din(n11954));
	jspl jspl_w_n11957_0(.douta(w_n11957_0[0]),.doutb(w_n11957_0[1]),.din(n11957));
	jspl jspl_w_n11959_0(.douta(w_n11959_0[0]),.doutb(w_n11959_0[1]),.din(n11959));
	jspl jspl_w_n11963_0(.douta(w_n11963_0[0]),.doutb(w_n11963_0[1]),.din(n11963));
	jspl jspl_w_n11965_0(.douta(w_n11965_0[0]),.doutb(w_n11965_0[1]),.din(n11965));
	jspl jspl_w_n11966_0(.douta(w_n11966_0[0]),.doutb(w_n11966_0[1]),.din(n11966));
	jspl jspl_w_n11967_0(.douta(w_n11967_0[0]),.doutb(w_n11967_0[1]),.din(n11967));
	jspl3 jspl3_w_n11968_0(.douta(w_n11968_0[0]),.doutb(w_n11968_0[1]),.doutc(w_n11968_0[2]),.din(n11968));
	jspl jspl_w_n11971_0(.douta(w_n11971_0[0]),.doutb(w_n11971_0[1]),.din(n11971));
	jspl jspl_w_n11972_0(.douta(w_n11972_0[0]),.doutb(w_n11972_0[1]),.din(n11972));
	jspl3 jspl3_w_n11973_0(.douta(w_n11973_0[0]),.doutb(w_n11973_0[1]),.doutc(w_n11973_0[2]),.din(n11973));
	jspl jspl_w_n11975_0(.douta(w_n11975_0[0]),.doutb(w_n11975_0[1]),.din(n11975));
	jspl jspl_w_n11979_0(.douta(w_n11979_0[0]),.doutb(w_n11979_0[1]),.din(n11979));
	jspl jspl_w_n11981_0(.douta(w_n11981_0[0]),.doutb(w_n11981_0[1]),.din(n11981));
	jspl jspl_w_n11982_0(.douta(w_n11982_0[0]),.doutb(w_n11982_0[1]),.din(n11982));
	jspl3 jspl3_w_n11983_0(.douta(w_n11983_0[0]),.doutb(w_n11983_0[1]),.doutc(w_n11983_0[2]),.din(n11983));
	jspl jspl_w_n11984_0(.douta(w_n11984_0[0]),.doutb(w_n11984_0[1]),.din(n11984));
	jspl jspl_w_n11987_0(.douta(w_n11987_0[0]),.doutb(w_n11987_0[1]),.din(n11987));
	jspl jspl_w_n11993_0(.douta(w_n11993_0[0]),.doutb(w_n11993_0[1]),.din(n11993));
	jspl jspl_w_n11994_0(.douta(w_n11994_0[0]),.doutb(w_n11994_0[1]),.din(n11994));
	jspl jspl_w_n11996_0(.douta(w_n11996_0[0]),.doutb(w_n11996_0[1]),.din(n11996));
	jspl jspl_w_n11998_0(.douta(w_n11998_0[0]),.doutb(w_n11998_0[1]),.din(n11998));
	jspl jspl_w_n12000_0(.douta(w_n12000_0[0]),.doutb(w_n12000_0[1]),.din(n12000));
	jspl jspl_w_n12006_0(.douta(w_n12006_0[0]),.doutb(w_n12006_0[1]),.din(n12006));
	jspl jspl_w_n12008_0(.douta(w_n12008_0[0]),.doutb(w_n12008_0[1]),.din(n12008));
	jspl3 jspl3_w_n12009_0(.douta(w_n12009_0[0]),.doutb(w_n12009_0[1]),.doutc(w_n12009_0[2]),.din(n12009));
	jspl jspl_w_n12012_0(.douta(w_n12012_0[0]),.doutb(w_n12012_0[1]),.din(n12012));
	jspl jspl_w_n12013_0(.douta(w_n12013_0[0]),.doutb(w_n12013_0[1]),.din(n12013));
	jspl3 jspl3_w_n12014_0(.douta(w_n12014_0[0]),.doutb(w_n12014_0[1]),.doutc(w_n12014_0[2]),.din(n12014));
	jspl jspl_w_n12016_0(.douta(w_n12016_0[0]),.doutb(w_n12016_0[1]),.din(n12016));
	jspl jspl_w_n12020_0(.douta(w_n12020_0[0]),.doutb(w_n12020_0[1]),.din(n12020));
	jspl jspl_w_n12022_0(.douta(w_n12022_0[0]),.doutb(w_n12022_0[1]),.din(n12022));
	jspl jspl_w_n12023_0(.douta(w_n12023_0[0]),.doutb(w_n12023_0[1]),.din(n12023));
	jspl3 jspl3_w_n12024_0(.douta(w_n12024_0[0]),.doutb(w_n12024_0[1]),.doutc(w_n12024_0[2]),.din(n12024));
	jspl jspl_w_n12025_0(.douta(w_n12025_0[0]),.doutb(w_n12025_0[1]),.din(n12025));
	jspl jspl_w_n12028_0(.douta(w_n12028_0[0]),.doutb(w_n12028_0[1]),.din(n12028));
	jspl jspl_w_n12034_0(.douta(w_n12034_0[0]),.doutb(w_n12034_0[1]),.din(n12034));
	jspl jspl_w_n12035_0(.douta(w_n12035_0[0]),.doutb(w_n12035_0[1]),.din(n12035));
	jspl jspl_w_n12037_0(.douta(w_n12037_0[0]),.doutb(w_n12037_0[1]),.din(n12037));
	jspl jspl_w_n12039_0(.douta(w_n12039_0[0]),.doutb(w_n12039_0[1]),.din(n12039));
	jspl jspl_w_n12041_0(.douta(w_n12041_0[0]),.doutb(w_n12041_0[1]),.din(n12041));
	jspl jspl_w_n12047_0(.douta(w_n12047_0[0]),.doutb(w_n12047_0[1]),.din(n12047));
	jspl jspl_w_n12049_0(.douta(w_n12049_0[0]),.doutb(w_n12049_0[1]),.din(n12049));
	jspl3 jspl3_w_n12050_0(.douta(w_n12050_0[0]),.doutb(w_n12050_0[1]),.doutc(w_n12050_0[2]),.din(n12050));
	jspl jspl_w_n12053_0(.douta(w_n12053_0[0]),.doutb(w_n12053_0[1]),.din(n12053));
	jspl jspl_w_n12054_0(.douta(w_n12054_0[0]),.doutb(w_n12054_0[1]),.din(n12054));
	jspl3 jspl3_w_n12055_0(.douta(w_n12055_0[0]),.doutb(w_n12055_0[1]),.doutc(w_n12055_0[2]),.din(n12055));
	jspl jspl_w_n12057_0(.douta(w_n12057_0[0]),.doutb(w_n12057_0[1]),.din(n12057));
	jspl jspl_w_n12061_0(.douta(w_n12061_0[0]),.doutb(w_n12061_0[1]),.din(n12061));
	jspl jspl_w_n12063_0(.douta(w_n12063_0[0]),.doutb(w_n12063_0[1]),.din(n12063));
	jspl jspl_w_n12064_0(.douta(w_n12064_0[0]),.doutb(w_n12064_0[1]),.din(n12064));
	jspl3 jspl3_w_n12065_0(.douta(w_n12065_0[0]),.doutb(w_n12065_0[1]),.doutc(w_n12065_0[2]),.din(n12065));
	jspl jspl_w_n12066_0(.douta(w_n12066_0[0]),.doutb(w_n12066_0[1]),.din(n12066));
	jspl jspl_w_n12069_0(.douta(w_n12069_0[0]),.doutb(w_n12069_0[1]),.din(n12069));
	jspl jspl_w_n12075_0(.douta(w_n12075_0[0]),.doutb(w_n12075_0[1]),.din(n12075));
	jspl jspl_w_n12076_0(.douta(w_n12076_0[0]),.doutb(w_n12076_0[1]),.din(n12076));
	jspl jspl_w_n12078_0(.douta(w_n12078_0[0]),.doutb(w_n12078_0[1]),.din(n12078));
	jspl jspl_w_n12080_0(.douta(w_n12080_0[0]),.doutb(w_n12080_0[1]),.din(n12080));
	jspl jspl_w_n12082_0(.douta(w_n12082_0[0]),.doutb(w_n12082_0[1]),.din(n12082));
	jspl jspl_w_n12088_0(.douta(w_n12088_0[0]),.doutb(w_n12088_0[1]),.din(n12088));
	jspl jspl_w_n12090_0(.douta(w_n12090_0[0]),.doutb(w_n12090_0[1]),.din(n12090));
	jspl3 jspl3_w_n12091_0(.douta(w_n12091_0[0]),.doutb(w_n12091_0[1]),.doutc(w_n12091_0[2]),.din(n12091));
	jspl jspl_w_n12094_0(.douta(w_n12094_0[0]),.doutb(w_n12094_0[1]),.din(n12094));
	jspl jspl_w_n12095_0(.douta(w_n12095_0[0]),.doutb(w_n12095_0[1]),.din(n12095));
	jspl3 jspl3_w_n12096_0(.douta(w_n12096_0[0]),.doutb(w_n12096_0[1]),.doutc(w_n12096_0[2]),.din(n12096));
	jspl jspl_w_n12098_0(.douta(w_n12098_0[0]),.doutb(w_n12098_0[1]),.din(n12098));
	jspl jspl_w_n12102_0(.douta(w_n12102_0[0]),.doutb(w_n12102_0[1]),.din(n12102));
	jspl jspl_w_n12104_0(.douta(w_n12104_0[0]),.doutb(w_n12104_0[1]),.din(n12104));
	jspl jspl_w_n12105_0(.douta(w_n12105_0[0]),.doutb(w_n12105_0[1]),.din(n12105));
	jspl3 jspl3_w_n12106_0(.douta(w_n12106_0[0]),.doutb(w_n12106_0[1]),.doutc(w_n12106_0[2]),.din(n12106));
	jspl jspl_w_n12110_0(.douta(w_n12110_0[0]),.doutb(w_n12110_0[1]),.din(n12110));
	jspl jspl_w_n12116_0(.douta(w_n12116_0[0]),.doutb(w_n12116_0[1]),.din(n12116));
	jspl3 jspl3_w_n12118_0(.douta(w_n12118_0[0]),.doutb(w_n12118_0[1]),.doutc(w_n12118_0[2]),.din(n12118));
	jspl jspl_w_n12120_0(.douta(w_n12120_0[0]),.doutb(w_n12120_0[1]),.din(n12120));
	jspl3 jspl3_w_n12125_0(.douta(w_n12125_0[0]),.doutb(w_n12125_0[1]),.doutc(w_n12125_0[2]),.din(n12125));
	jspl jspl_w_n12126_0(.douta(w_n12126_0[0]),.doutb(w_n12126_0[1]),.din(n12126));
	jspl jspl_w_n12127_0(.douta(w_n12127_0[0]),.doutb(w_n12127_0[1]),.din(n12127));
	jspl jspl_w_n12132_0(.douta(w_n12132_0[0]),.doutb(w_n12132_0[1]),.din(n12132));
	jspl3 jspl3_w_n12133_0(.douta(w_n12133_0[0]),.doutb(w_n12133_0[1]),.doutc(w_n12133_0[2]),.din(n12133));
	jspl jspl_w_n12138_0(.douta(w_n12138_0[0]),.doutb(w_n12138_0[1]),.din(n12138));
	jspl jspl_w_n12145_0(.douta(w_n12145_0[0]),.doutb(w_n12145_0[1]),.din(n12145));
	jspl3 jspl3_w_n12148_0(.douta(w_n12148_0[0]),.doutb(w_n12148_0[1]),.doutc(w_n12148_0[2]),.din(n12148));
	jspl jspl_w_n12148_1(.douta(w_n12148_1[0]),.doutb(w_n12148_1[1]),.din(w_n12148_0[0]));
	jspl jspl_w_n12149_0(.douta(w_n12149_0[0]),.doutb(w_n12149_0[1]),.din(n12149));
	jspl3 jspl3_w_n12152_0(.douta(w_n12152_0[0]),.doutb(w_n12152_0[1]),.doutc(w_n12152_0[2]),.din(n12152));
	jspl jspl_w_n12153_0(.douta(w_n12153_0[0]),.doutb(w_n12153_0[1]),.din(n12153));
	jspl jspl_w_n12154_0(.douta(w_n12154_0[0]),.doutb(w_n12154_0[1]),.din(n12154));
	jspl jspl_w_n12155_0(.douta(w_n12155_0[0]),.doutb(w_n12155_0[1]),.din(n12155));
	jspl jspl_w_n12157_0(.douta(w_n12157_0[0]),.doutb(w_n12157_0[1]),.din(n12157));
	jspl jspl_w_n12159_0(.douta(w_n12159_0[0]),.doutb(w_n12159_0[1]),.din(n12159));
	jspl jspl_w_n12161_0(.douta(w_n12161_0[0]),.doutb(w_n12161_0[1]),.din(n12161));
	jspl jspl_w_n12170_0(.douta(w_n12170_0[0]),.doutb(w_n12170_0[1]),.din(n12170));
	jspl3 jspl3_w_n12172_0(.douta(w_n12172_0[0]),.doutb(w_n12172_0[1]),.doutc(w_n12172_0[2]),.din(n12172));
	jspl jspl_w_n12173_0(.douta(w_n12173_0[0]),.doutb(w_n12173_0[1]),.din(n12173));
	jspl jspl_w_n12177_0(.douta(w_n12177_0[0]),.doutb(w_n12177_0[1]),.din(n12177));
	jspl jspl_w_n12179_0(.douta(w_n12179_0[0]),.doutb(w_n12179_0[1]),.din(n12179));
	jspl jspl_w_n12181_0(.douta(w_n12181_0[0]),.doutb(w_n12181_0[1]),.din(n12181));
	jspl jspl_w_n12186_0(.douta(w_n12186_0[0]),.doutb(w_n12186_0[1]),.din(n12186));
	jspl jspl_w_n12188_0(.douta(w_n12188_0[0]),.doutb(w_n12188_0[1]),.din(n12188));
	jspl jspl_w_n12189_0(.douta(w_n12189_0[0]),.doutb(w_n12189_0[1]),.din(n12189));
	jspl3 jspl3_w_n12190_0(.douta(w_n12190_0[0]),.doutb(w_n12190_0[1]),.doutc(w_n12190_0[2]),.din(n12190));
	jspl jspl_w_n12191_0(.douta(w_n12191_0[0]),.doutb(w_n12191_0[1]),.din(n12191));
	jspl jspl_w_n12196_0(.douta(w_n12196_0[0]),.doutb(w_n12196_0[1]),.din(n12196));
	jspl jspl_w_n12197_0(.douta(w_n12197_0[0]),.doutb(w_n12197_0[1]),.din(n12197));
	jspl jspl_w_n12199_0(.douta(w_n12199_0[0]),.doutb(w_n12199_0[1]),.din(n12199));
	jspl jspl_w_n12201_0(.douta(w_n12201_0[0]),.doutb(w_n12201_0[1]),.din(n12201));
	jspl jspl_w_n12204_0(.douta(w_n12204_0[0]),.doutb(w_n12204_0[1]),.din(n12204));
	jspl jspl_w_n12210_0(.douta(w_n12210_0[0]),.doutb(w_n12210_0[1]),.din(n12210));
	jspl3 jspl3_w_n12212_0(.douta(w_n12212_0[0]),.doutb(w_n12212_0[1]),.doutc(w_n12212_0[2]),.din(n12212));
	jspl jspl_w_n12213_0(.douta(w_n12213_0[0]),.doutb(w_n12213_0[1]),.din(n12213));
	jspl jspl_w_n12217_0(.douta(w_n12217_0[0]),.doutb(w_n12217_0[1]),.din(n12217));
	jspl jspl_w_n12218_0(.douta(w_n12218_0[0]),.doutb(w_n12218_0[1]),.din(n12218));
	jspl jspl_w_n12220_0(.douta(w_n12220_0[0]),.doutb(w_n12220_0[1]),.din(n12220));
	jspl jspl_w_n12225_0(.douta(w_n12225_0[0]),.doutb(w_n12225_0[1]),.din(n12225));
	jspl jspl_w_n12227_0(.douta(w_n12227_0[0]),.doutb(w_n12227_0[1]),.din(n12227));
	jspl jspl_w_n12228_0(.douta(w_n12228_0[0]),.doutb(w_n12228_0[1]),.din(n12228));
	jspl3 jspl3_w_n12229_0(.douta(w_n12229_0[0]),.doutb(w_n12229_0[1]),.doutc(w_n12229_0[2]),.din(n12229));
	jspl jspl_w_n12230_0(.douta(w_n12230_0[0]),.doutb(w_n12230_0[1]),.din(n12230));
	jspl jspl_w_n12234_0(.douta(w_n12234_0[0]),.doutb(w_n12234_0[1]),.din(n12234));
	jspl jspl_w_n12235_0(.douta(w_n12235_0[0]),.doutb(w_n12235_0[1]),.din(n12235));
	jspl jspl_w_n12237_0(.douta(w_n12237_0[0]),.doutb(w_n12237_0[1]),.din(n12237));
	jspl jspl_w_n12239_0(.douta(w_n12239_0[0]),.doutb(w_n12239_0[1]),.din(n12239));
	jspl jspl_w_n12242_0(.douta(w_n12242_0[0]),.doutb(w_n12242_0[1]),.din(n12242));
	jspl jspl_w_n12248_0(.douta(w_n12248_0[0]),.doutb(w_n12248_0[1]),.din(n12248));
	jspl jspl_w_n12250_0(.douta(w_n12250_0[0]),.doutb(w_n12250_0[1]),.din(n12250));
	jspl3 jspl3_w_n12251_0(.douta(w_n12251_0[0]),.doutb(w_n12251_0[1]),.doutc(w_n12251_0[2]),.din(n12251));
	jspl jspl_w_n12255_0(.douta(w_n12255_0[0]),.doutb(w_n12255_0[1]),.din(n12255));
	jspl jspl_w_n12256_0(.douta(w_n12256_0[0]),.doutb(w_n12256_0[1]),.din(n12256));
	jspl3 jspl3_w_n12257_0(.douta(w_n12257_0[0]),.doutb(w_n12257_0[1]),.doutc(w_n12257_0[2]),.din(n12257));
	jspl jspl_w_n12259_0(.douta(w_n12259_0[0]),.doutb(w_n12259_0[1]),.din(n12259));
	jspl jspl_w_n12264_0(.douta(w_n12264_0[0]),.doutb(w_n12264_0[1]),.din(n12264));
	jspl jspl_w_n12266_0(.douta(w_n12266_0[0]),.doutb(w_n12266_0[1]),.din(n12266));
	jspl jspl_w_n12267_0(.douta(w_n12267_0[0]),.doutb(w_n12267_0[1]),.din(n12267));
	jspl3 jspl3_w_n12268_0(.douta(w_n12268_0[0]),.doutb(w_n12268_0[1]),.doutc(w_n12268_0[2]),.din(n12268));
	jspl jspl_w_n12269_0(.douta(w_n12269_0[0]),.doutb(w_n12269_0[1]),.din(n12269));
	jspl jspl_w_n12273_0(.douta(w_n12273_0[0]),.doutb(w_n12273_0[1]),.din(n12273));
	jspl jspl_w_n12279_0(.douta(w_n12279_0[0]),.doutb(w_n12279_0[1]),.din(n12279));
	jspl jspl_w_n12280_0(.douta(w_n12280_0[0]),.doutb(w_n12280_0[1]),.din(n12280));
	jspl jspl_w_n12282_0(.douta(w_n12282_0[0]),.doutb(w_n12282_0[1]),.din(n12282));
	jspl jspl_w_n12284_0(.douta(w_n12284_0[0]),.doutb(w_n12284_0[1]),.din(n12284));
	jspl jspl_w_n12287_0(.douta(w_n12287_0[0]),.doutb(w_n12287_0[1]),.din(n12287));
	jspl jspl_w_n12293_0(.douta(w_n12293_0[0]),.doutb(w_n12293_0[1]),.din(n12293));
	jspl jspl_w_n12295_0(.douta(w_n12295_0[0]),.doutb(w_n12295_0[1]),.din(n12295));
	jspl3 jspl3_w_n12296_0(.douta(w_n12296_0[0]),.doutb(w_n12296_0[1]),.doutc(w_n12296_0[2]),.din(n12296));
	jspl jspl_w_n12300_0(.douta(w_n12300_0[0]),.doutb(w_n12300_0[1]),.din(n12300));
	jspl jspl_w_n12301_0(.douta(w_n12301_0[0]),.doutb(w_n12301_0[1]),.din(n12301));
	jspl3 jspl3_w_n12302_0(.douta(w_n12302_0[0]),.doutb(w_n12302_0[1]),.doutc(w_n12302_0[2]),.din(n12302));
	jspl jspl_w_n12304_0(.douta(w_n12304_0[0]),.doutb(w_n12304_0[1]),.din(n12304));
	jspl jspl_w_n12309_0(.douta(w_n12309_0[0]),.doutb(w_n12309_0[1]),.din(n12309));
	jspl jspl_w_n12311_0(.douta(w_n12311_0[0]),.doutb(w_n12311_0[1]),.din(n12311));
	jspl jspl_w_n12312_0(.douta(w_n12312_0[0]),.doutb(w_n12312_0[1]),.din(n12312));
	jspl3 jspl3_w_n12313_0(.douta(w_n12313_0[0]),.doutb(w_n12313_0[1]),.doutc(w_n12313_0[2]),.din(n12313));
	jspl jspl_w_n12314_0(.douta(w_n12314_0[0]),.doutb(w_n12314_0[1]),.din(n12314));
	jspl jspl_w_n12318_0(.douta(w_n12318_0[0]),.doutb(w_n12318_0[1]),.din(n12318));
	jspl jspl_w_n12324_0(.douta(w_n12324_0[0]),.doutb(w_n12324_0[1]),.din(n12324));
	jspl jspl_w_n12325_0(.douta(w_n12325_0[0]),.doutb(w_n12325_0[1]),.din(n12325));
	jspl jspl_w_n12327_0(.douta(w_n12327_0[0]),.doutb(w_n12327_0[1]),.din(n12327));
	jspl jspl_w_n12329_0(.douta(w_n12329_0[0]),.doutb(w_n12329_0[1]),.din(n12329));
	jspl jspl_w_n12332_0(.douta(w_n12332_0[0]),.doutb(w_n12332_0[1]),.din(n12332));
	jspl jspl_w_n12338_0(.douta(w_n12338_0[0]),.doutb(w_n12338_0[1]),.din(n12338));
	jspl jspl_w_n12340_0(.douta(w_n12340_0[0]),.doutb(w_n12340_0[1]),.din(n12340));
	jspl3 jspl3_w_n12341_0(.douta(w_n12341_0[0]),.doutb(w_n12341_0[1]),.doutc(w_n12341_0[2]),.din(n12341));
	jspl jspl_w_n12345_0(.douta(w_n12345_0[0]),.doutb(w_n12345_0[1]),.din(n12345));
	jspl jspl_w_n12346_0(.douta(w_n12346_0[0]),.doutb(w_n12346_0[1]),.din(n12346));
	jspl3 jspl3_w_n12347_0(.douta(w_n12347_0[0]),.doutb(w_n12347_0[1]),.doutc(w_n12347_0[2]),.din(n12347));
	jspl jspl_w_n12349_0(.douta(w_n12349_0[0]),.doutb(w_n12349_0[1]),.din(n12349));
	jspl jspl_w_n12354_0(.douta(w_n12354_0[0]),.doutb(w_n12354_0[1]),.din(n12354));
	jspl jspl_w_n12356_0(.douta(w_n12356_0[0]),.doutb(w_n12356_0[1]),.din(n12356));
	jspl jspl_w_n12357_0(.douta(w_n12357_0[0]),.doutb(w_n12357_0[1]),.din(n12357));
	jspl3 jspl3_w_n12358_0(.douta(w_n12358_0[0]),.doutb(w_n12358_0[1]),.doutc(w_n12358_0[2]),.din(n12358));
	jspl jspl_w_n12359_0(.douta(w_n12359_0[0]),.doutb(w_n12359_0[1]),.din(n12359));
	jspl jspl_w_n12363_0(.douta(w_n12363_0[0]),.doutb(w_n12363_0[1]),.din(n12363));
	jspl jspl_w_n12369_0(.douta(w_n12369_0[0]),.doutb(w_n12369_0[1]),.din(n12369));
	jspl jspl_w_n12370_0(.douta(w_n12370_0[0]),.doutb(w_n12370_0[1]),.din(n12370));
	jspl jspl_w_n12372_0(.douta(w_n12372_0[0]),.doutb(w_n12372_0[1]),.din(n12372));
	jspl jspl_w_n12374_0(.douta(w_n12374_0[0]),.doutb(w_n12374_0[1]),.din(n12374));
	jspl jspl_w_n12377_0(.douta(w_n12377_0[0]),.doutb(w_n12377_0[1]),.din(n12377));
	jspl jspl_w_n12383_0(.douta(w_n12383_0[0]),.doutb(w_n12383_0[1]),.din(n12383));
	jspl jspl_w_n12385_0(.douta(w_n12385_0[0]),.doutb(w_n12385_0[1]),.din(n12385));
	jspl3 jspl3_w_n12386_0(.douta(w_n12386_0[0]),.doutb(w_n12386_0[1]),.doutc(w_n12386_0[2]),.din(n12386));
	jspl jspl_w_n12390_0(.douta(w_n12390_0[0]),.doutb(w_n12390_0[1]),.din(n12390));
	jspl jspl_w_n12391_0(.douta(w_n12391_0[0]),.doutb(w_n12391_0[1]),.din(n12391));
	jspl3 jspl3_w_n12392_0(.douta(w_n12392_0[0]),.doutb(w_n12392_0[1]),.doutc(w_n12392_0[2]),.din(n12392));
	jspl jspl_w_n12394_0(.douta(w_n12394_0[0]),.doutb(w_n12394_0[1]),.din(n12394));
	jspl jspl_w_n12399_0(.douta(w_n12399_0[0]),.doutb(w_n12399_0[1]),.din(n12399));
	jspl jspl_w_n12401_0(.douta(w_n12401_0[0]),.doutb(w_n12401_0[1]),.din(n12401));
	jspl jspl_w_n12402_0(.douta(w_n12402_0[0]),.doutb(w_n12402_0[1]),.din(n12402));
	jspl3 jspl3_w_n12403_0(.douta(w_n12403_0[0]),.doutb(w_n12403_0[1]),.doutc(w_n12403_0[2]),.din(n12403));
	jspl jspl_w_n12404_0(.douta(w_n12404_0[0]),.doutb(w_n12404_0[1]),.din(n12404));
	jspl jspl_w_n12408_0(.douta(w_n12408_0[0]),.doutb(w_n12408_0[1]),.din(n12408));
	jspl jspl_w_n12414_0(.douta(w_n12414_0[0]),.doutb(w_n12414_0[1]),.din(n12414));
	jspl jspl_w_n12415_0(.douta(w_n12415_0[0]),.doutb(w_n12415_0[1]),.din(n12415));
	jspl jspl_w_n12417_0(.douta(w_n12417_0[0]),.doutb(w_n12417_0[1]),.din(n12417));
	jspl jspl_w_n12419_0(.douta(w_n12419_0[0]),.doutb(w_n12419_0[1]),.din(n12419));
	jspl jspl_w_n12422_0(.douta(w_n12422_0[0]),.doutb(w_n12422_0[1]),.din(n12422));
	jspl jspl_w_n12428_0(.douta(w_n12428_0[0]),.doutb(w_n12428_0[1]),.din(n12428));
	jspl jspl_w_n12430_0(.douta(w_n12430_0[0]),.doutb(w_n12430_0[1]),.din(n12430));
	jspl3 jspl3_w_n12431_0(.douta(w_n12431_0[0]),.doutb(w_n12431_0[1]),.doutc(w_n12431_0[2]),.din(n12431));
	jspl jspl_w_n12435_0(.douta(w_n12435_0[0]),.doutb(w_n12435_0[1]),.din(n12435));
	jspl jspl_w_n12436_0(.douta(w_n12436_0[0]),.doutb(w_n12436_0[1]),.din(n12436));
	jspl3 jspl3_w_n12437_0(.douta(w_n12437_0[0]),.doutb(w_n12437_0[1]),.doutc(w_n12437_0[2]),.din(n12437));
	jspl jspl_w_n12439_0(.douta(w_n12439_0[0]),.doutb(w_n12439_0[1]),.din(n12439));
	jspl jspl_w_n12444_0(.douta(w_n12444_0[0]),.doutb(w_n12444_0[1]),.din(n12444));
	jspl jspl_w_n12446_0(.douta(w_n12446_0[0]),.doutb(w_n12446_0[1]),.din(n12446));
	jspl jspl_w_n12447_0(.douta(w_n12447_0[0]),.doutb(w_n12447_0[1]),.din(n12447));
	jspl3 jspl3_w_n12448_0(.douta(w_n12448_0[0]),.doutb(w_n12448_0[1]),.doutc(w_n12448_0[2]),.din(n12448));
	jspl jspl_w_n12449_0(.douta(w_n12449_0[0]),.doutb(w_n12449_0[1]),.din(n12449));
	jspl jspl_w_n12453_0(.douta(w_n12453_0[0]),.doutb(w_n12453_0[1]),.din(n12453));
	jspl jspl_w_n12459_0(.douta(w_n12459_0[0]),.doutb(w_n12459_0[1]),.din(n12459));
	jspl jspl_w_n12460_0(.douta(w_n12460_0[0]),.doutb(w_n12460_0[1]),.din(n12460));
	jspl jspl_w_n12462_0(.douta(w_n12462_0[0]),.doutb(w_n12462_0[1]),.din(n12462));
	jspl jspl_w_n12467_0(.douta(w_n12467_0[0]),.doutb(w_n12467_0[1]),.din(n12467));
	jspl jspl_w_n12469_0(.douta(w_n12469_0[0]),.doutb(w_n12469_0[1]),.din(n12469));
	jspl jspl_w_n12470_0(.douta(w_n12470_0[0]),.doutb(w_n12470_0[1]),.din(n12470));
	jspl3 jspl3_w_n12471_0(.douta(w_n12471_0[0]),.doutb(w_n12471_0[1]),.doutc(w_n12471_0[2]),.din(n12471));
	jspl jspl_w_n12472_0(.douta(w_n12472_0[0]),.doutb(w_n12472_0[1]),.din(n12472));
	jspl jspl_w_n12474_0(.douta(w_n12474_0[0]),.doutb(w_n12474_0[1]),.din(n12474));
	jspl jspl_w_n12476_0(.douta(w_n12476_0[0]),.doutb(w_n12476_0[1]),.din(n12476));
	jspl jspl_w_n12478_0(.douta(w_n12478_0[0]),.doutb(w_n12478_0[1]),.din(n12478));
	jspl jspl_w_n12481_0(.douta(w_n12481_0[0]),.doutb(w_n12481_0[1]),.din(n12481));
	jspl jspl_w_n12487_0(.douta(w_n12487_0[0]),.doutb(w_n12487_0[1]),.din(n12487));
	jspl3 jspl3_w_n12489_0(.douta(w_n12489_0[0]),.doutb(w_n12489_0[1]),.doutc(w_n12489_0[2]),.din(n12489));
	jspl jspl_w_n12490_0(.douta(w_n12490_0[0]),.doutb(w_n12490_0[1]),.din(n12490));
	jspl jspl_w_n12494_0(.douta(w_n12494_0[0]),.doutb(w_n12494_0[1]),.din(n12494));
	jspl jspl_w_n12500_0(.douta(w_n12500_0[0]),.doutb(w_n12500_0[1]),.din(n12500));
	jspl jspl_w_n12501_0(.douta(w_n12501_0[0]),.doutb(w_n12501_0[1]),.din(n12501));
	jspl jspl_w_n12503_0(.douta(w_n12503_0[0]),.doutb(w_n12503_0[1]),.din(n12503));
	jspl jspl_w_n12505_0(.douta(w_n12505_0[0]),.doutb(w_n12505_0[1]),.din(n12505));
	jspl jspl_w_n12508_0(.douta(w_n12508_0[0]),.doutb(w_n12508_0[1]),.din(n12508));
	jspl jspl_w_n12514_0(.douta(w_n12514_0[0]),.doutb(w_n12514_0[1]),.din(n12514));
	jspl jspl_w_n12516_0(.douta(w_n12516_0[0]),.doutb(w_n12516_0[1]),.din(n12516));
	jspl3 jspl3_w_n12517_0(.douta(w_n12517_0[0]),.doutb(w_n12517_0[1]),.doutc(w_n12517_0[2]),.din(n12517));
	jspl jspl_w_n12521_0(.douta(w_n12521_0[0]),.doutb(w_n12521_0[1]),.din(n12521));
	jspl jspl_w_n12522_0(.douta(w_n12522_0[0]),.doutb(w_n12522_0[1]),.din(n12522));
	jspl3 jspl3_w_n12523_0(.douta(w_n12523_0[0]),.doutb(w_n12523_0[1]),.doutc(w_n12523_0[2]),.din(n12523));
	jspl jspl_w_n12525_0(.douta(w_n12525_0[0]),.doutb(w_n12525_0[1]),.din(n12525));
	jspl jspl_w_n12530_0(.douta(w_n12530_0[0]),.doutb(w_n12530_0[1]),.din(n12530));
	jspl jspl_w_n12532_0(.douta(w_n12532_0[0]),.doutb(w_n12532_0[1]),.din(n12532));
	jspl jspl_w_n12533_0(.douta(w_n12533_0[0]),.doutb(w_n12533_0[1]),.din(n12533));
	jspl3 jspl3_w_n12534_0(.douta(w_n12534_0[0]),.doutb(w_n12534_0[1]),.doutc(w_n12534_0[2]),.din(n12534));
	jspl jspl_w_n12535_0(.douta(w_n12535_0[0]),.doutb(w_n12535_0[1]),.din(n12535));
	jspl jspl_w_n12539_0(.douta(w_n12539_0[0]),.doutb(w_n12539_0[1]),.din(n12539));
	jspl jspl_w_n12545_0(.douta(w_n12545_0[0]),.doutb(w_n12545_0[1]),.din(n12545));
	jspl jspl_w_n12546_0(.douta(w_n12546_0[0]),.doutb(w_n12546_0[1]),.din(n12546));
	jspl jspl_w_n12548_0(.douta(w_n12548_0[0]),.doutb(w_n12548_0[1]),.din(n12548));
	jspl jspl_w_n12550_0(.douta(w_n12550_0[0]),.doutb(w_n12550_0[1]),.din(n12550));
	jspl jspl_w_n12553_0(.douta(w_n12553_0[0]),.doutb(w_n12553_0[1]),.din(n12553));
	jspl jspl_w_n12559_0(.douta(w_n12559_0[0]),.doutb(w_n12559_0[1]),.din(n12559));
	jspl jspl_w_n12561_0(.douta(w_n12561_0[0]),.doutb(w_n12561_0[1]),.din(n12561));
	jspl3 jspl3_w_n12562_0(.douta(w_n12562_0[0]),.doutb(w_n12562_0[1]),.doutc(w_n12562_0[2]),.din(n12562));
	jspl jspl_w_n12566_0(.douta(w_n12566_0[0]),.doutb(w_n12566_0[1]),.din(n12566));
	jspl jspl_w_n12567_0(.douta(w_n12567_0[0]),.doutb(w_n12567_0[1]),.din(n12567));
	jspl3 jspl3_w_n12568_0(.douta(w_n12568_0[0]),.doutb(w_n12568_0[1]),.doutc(w_n12568_0[2]),.din(n12568));
	jspl jspl_w_n12570_0(.douta(w_n12570_0[0]),.doutb(w_n12570_0[1]),.din(n12570));
	jspl jspl_w_n12575_0(.douta(w_n12575_0[0]),.doutb(w_n12575_0[1]),.din(n12575));
	jspl jspl_w_n12577_0(.douta(w_n12577_0[0]),.doutb(w_n12577_0[1]),.din(n12577));
	jspl jspl_w_n12578_0(.douta(w_n12578_0[0]),.doutb(w_n12578_0[1]),.din(n12578));
	jspl3 jspl3_w_n12579_0(.douta(w_n12579_0[0]),.doutb(w_n12579_0[1]),.doutc(w_n12579_0[2]),.din(n12579));
	jspl jspl_w_n12580_0(.douta(w_n12580_0[0]),.doutb(w_n12580_0[1]),.din(n12580));
	jspl jspl_w_n12584_0(.douta(w_n12584_0[0]),.doutb(w_n12584_0[1]),.din(n12584));
	jspl jspl_w_n12590_0(.douta(w_n12590_0[0]),.doutb(w_n12590_0[1]),.din(n12590));
	jspl jspl_w_n12591_0(.douta(w_n12591_0[0]),.doutb(w_n12591_0[1]),.din(n12591));
	jspl jspl_w_n12593_0(.douta(w_n12593_0[0]),.doutb(w_n12593_0[1]),.din(n12593));
	jspl jspl_w_n12595_0(.douta(w_n12595_0[0]),.doutb(w_n12595_0[1]),.din(n12595));
	jspl jspl_w_n12598_0(.douta(w_n12598_0[0]),.doutb(w_n12598_0[1]),.din(n12598));
	jspl jspl_w_n12604_0(.douta(w_n12604_0[0]),.doutb(w_n12604_0[1]),.din(n12604));
	jspl jspl_w_n12606_0(.douta(w_n12606_0[0]),.doutb(w_n12606_0[1]),.din(n12606));
	jspl3 jspl3_w_n12607_0(.douta(w_n12607_0[0]),.doutb(w_n12607_0[1]),.doutc(w_n12607_0[2]),.din(n12607));
	jspl jspl_w_n12611_0(.douta(w_n12611_0[0]),.doutb(w_n12611_0[1]),.din(n12611));
	jspl jspl_w_n12612_0(.douta(w_n12612_0[0]),.doutb(w_n12612_0[1]),.din(n12612));
	jspl3 jspl3_w_n12613_0(.douta(w_n12613_0[0]),.doutb(w_n12613_0[1]),.doutc(w_n12613_0[2]),.din(n12613));
	jspl jspl_w_n12615_0(.douta(w_n12615_0[0]),.doutb(w_n12615_0[1]),.din(n12615));
	jspl jspl_w_n12620_0(.douta(w_n12620_0[0]),.doutb(w_n12620_0[1]),.din(n12620));
	jspl jspl_w_n12622_0(.douta(w_n12622_0[0]),.doutb(w_n12622_0[1]),.din(n12622));
	jspl jspl_w_n12623_0(.douta(w_n12623_0[0]),.doutb(w_n12623_0[1]),.din(n12623));
	jspl3 jspl3_w_n12624_0(.douta(w_n12624_0[0]),.doutb(w_n12624_0[1]),.doutc(w_n12624_0[2]),.din(n12624));
	jspl jspl_w_n12625_0(.douta(w_n12625_0[0]),.doutb(w_n12625_0[1]),.din(n12625));
	jspl jspl_w_n12629_0(.douta(w_n12629_0[0]),.doutb(w_n12629_0[1]),.din(n12629));
	jspl jspl_w_n12635_0(.douta(w_n12635_0[0]),.doutb(w_n12635_0[1]),.din(n12635));
	jspl jspl_w_n12636_0(.douta(w_n12636_0[0]),.doutb(w_n12636_0[1]),.din(n12636));
	jspl jspl_w_n12638_0(.douta(w_n12638_0[0]),.doutb(w_n12638_0[1]),.din(n12638));
	jspl jspl_w_n12640_0(.douta(w_n12640_0[0]),.doutb(w_n12640_0[1]),.din(n12640));
	jspl jspl_w_n12643_0(.douta(w_n12643_0[0]),.doutb(w_n12643_0[1]),.din(n12643));
	jspl jspl_w_n12649_0(.douta(w_n12649_0[0]),.doutb(w_n12649_0[1]),.din(n12649));
	jspl3 jspl3_w_n12651_0(.douta(w_n12651_0[0]),.doutb(w_n12651_0[1]),.doutc(w_n12651_0[2]),.din(n12651));
	jspl3 jspl3_w_n12651_1(.douta(w_n12651_1[0]),.doutb(w_n12651_1[1]),.doutc(w_n12651_1[2]),.din(w_n12651_0[0]));
	jspl jspl_w_n12654_0(.douta(w_n12654_0[0]),.doutb(w_n12654_0[1]),.din(n12654));
	jspl3 jspl3_w_n12655_0(.douta(w_n12655_0[0]),.doutb(w_n12655_0[1]),.doutc(w_n12655_0[2]),.din(n12655));
	jspl jspl_w_n12656_0(.douta(w_n12656_0[0]),.doutb(w_n12656_0[1]),.din(n12656));
	jspl jspl_w_n12662_0(.douta(w_n12662_0[0]),.doutb(w_n12662_0[1]),.din(n12662));
	jspl3 jspl3_w_n12663_0(.douta(w_n12663_0[0]),.doutb(w_n12663_0[1]),.doutc(w_n12663_0[2]),.din(n12663));
	jspl jspl_w_n12664_0(.douta(w_n12664_0[0]),.doutb(w_n12664_0[1]),.din(n12664));
	jspl jspl_w_n12669_0(.douta(w_n12669_0[0]),.doutb(w_n12669_0[1]),.din(n12669));
	jspl3 jspl3_w_n12670_0(.douta(w_n12670_0[0]),.doutb(w_n12670_0[1]),.doutc(w_n12670_0[2]),.din(n12670));
	jspl3 jspl3_w_n12670_1(.douta(w_n12670_1[0]),.doutb(w_n12670_1[1]),.doutc(w_n12670_1[2]),.din(w_n12670_0[0]));
	jspl3 jspl3_w_n12670_2(.douta(w_n12670_2[0]),.doutb(w_n12670_2[1]),.doutc(w_n12670_2[2]),.din(w_n12670_0[1]));
	jspl3 jspl3_w_n12670_3(.douta(w_n12670_3[0]),.doutb(w_n12670_3[1]),.doutc(w_n12670_3[2]),.din(w_n12670_0[2]));
	jspl3 jspl3_w_n12670_4(.douta(w_n12670_4[0]),.doutb(w_n12670_4[1]),.doutc(w_n12670_4[2]),.din(w_n12670_1[0]));
	jspl3 jspl3_w_n12670_5(.douta(w_n12670_5[0]),.doutb(w_n12670_5[1]),.doutc(w_n12670_5[2]),.din(w_n12670_1[1]));
	jspl3 jspl3_w_n12670_6(.douta(w_n12670_6[0]),.doutb(w_n12670_6[1]),.doutc(w_n12670_6[2]),.din(w_n12670_1[2]));
	jspl3 jspl3_w_n12670_7(.douta(w_n12670_7[0]),.doutb(w_n12670_7[1]),.doutc(w_n12670_7[2]),.din(w_n12670_2[0]));
	jspl3 jspl3_w_n12670_8(.douta(w_n12670_8[0]),.doutb(w_n12670_8[1]),.doutc(w_n12670_8[2]),.din(w_n12670_2[1]));
	jspl3 jspl3_w_n12670_9(.douta(w_n12670_9[0]),.doutb(w_n12670_9[1]),.doutc(w_n12670_9[2]),.din(w_n12670_2[2]));
	jspl3 jspl3_w_n12670_10(.douta(w_n12670_10[0]),.doutb(w_n12670_10[1]),.doutc(w_n12670_10[2]),.din(w_n12670_3[0]));
	jspl3 jspl3_w_n12675_0(.douta(w_n12675_0[0]),.doutb(w_n12675_0[1]),.doutc(w_n12675_0[2]),.din(n12675));
	jspl3 jspl3_w_n12675_1(.douta(w_n12675_1[0]),.doutb(w_n12675_1[1]),.doutc(w_n12675_1[2]),.din(w_n12675_0[0]));
	jspl3 jspl3_w_n12675_2(.douta(w_n12675_2[0]),.doutb(w_n12675_2[1]),.doutc(w_n12675_2[2]),.din(w_n12675_0[1]));
	jspl3 jspl3_w_n12675_3(.douta(w_n12675_3[0]),.doutb(w_n12675_3[1]),.doutc(w_n12675_3[2]),.din(w_n12675_0[2]));
	jspl3 jspl3_w_n12675_4(.douta(w_n12675_4[0]),.doutb(w_n12675_4[1]),.doutc(w_n12675_4[2]),.din(w_n12675_1[0]));
	jspl3 jspl3_w_n12675_5(.douta(w_n12675_5[0]),.doutb(w_n12675_5[1]),.doutc(w_n12675_5[2]),.din(w_n12675_1[1]));
	jspl3 jspl3_w_n12675_6(.douta(w_n12675_6[0]),.doutb(w_n12675_6[1]),.doutc(w_n12675_6[2]),.din(w_n12675_1[2]));
	jspl3 jspl3_w_n12675_7(.douta(w_n12675_7[0]),.doutb(w_n12675_7[1]),.doutc(w_n12675_7[2]),.din(w_n12675_2[0]));
	jspl3 jspl3_w_n12675_8(.douta(w_n12675_8[0]),.doutb(w_n12675_8[1]),.doutc(w_n12675_8[2]),.din(w_n12675_2[1]));
	jspl3 jspl3_w_n12675_9(.douta(w_n12675_9[0]),.doutb(w_n12675_9[1]),.doutc(w_n12675_9[2]),.din(w_n12675_2[2]));
	jspl3 jspl3_w_n12675_10(.douta(w_n12675_10[0]),.doutb(w_n12675_10[1]),.doutc(w_n12675_10[2]),.din(w_n12675_3[0]));
	jspl3 jspl3_w_n12675_11(.douta(w_n12675_11[0]),.doutb(w_n12675_11[1]),.doutc(w_n12675_11[2]),.din(w_n12675_3[1]));
	jspl3 jspl3_w_n12675_12(.douta(w_n12675_12[0]),.doutb(w_n12675_12[1]),.doutc(w_n12675_12[2]),.din(w_n12675_3[2]));
	jspl3 jspl3_w_n12675_13(.douta(w_n12675_13[0]),.doutb(w_n12675_13[1]),.doutc(w_n12675_13[2]),.din(w_n12675_4[0]));
	jspl3 jspl3_w_n12675_14(.douta(w_n12675_14[0]),.doutb(w_n12675_14[1]),.doutc(w_n12675_14[2]),.din(w_n12675_4[1]));
	jspl3 jspl3_w_n12675_15(.douta(w_n12675_15[0]),.doutb(w_n12675_15[1]),.doutc(w_n12675_15[2]),.din(w_n12675_4[2]));
	jspl3 jspl3_w_n12675_16(.douta(w_n12675_16[0]),.doutb(w_n12675_16[1]),.doutc(w_n12675_16[2]),.din(w_n12675_5[0]));
	jspl3 jspl3_w_n12675_17(.douta(w_n12675_17[0]),.doutb(w_n12675_17[1]),.doutc(w_n12675_17[2]),.din(w_n12675_5[1]));
	jspl3 jspl3_w_n12675_18(.douta(w_n12675_18[0]),.doutb(w_n12675_18[1]),.doutc(w_n12675_18[2]),.din(w_n12675_5[2]));
	jspl3 jspl3_w_n12675_19(.douta(w_n12675_19[0]),.doutb(w_n12675_19[1]),.doutc(w_n12675_19[2]),.din(w_n12675_6[0]));
	jspl3 jspl3_w_n12675_20(.douta(w_n12675_20[0]),.doutb(w_n12675_20[1]),.doutc(w_n12675_20[2]),.din(w_n12675_6[1]));
	jspl3 jspl3_w_n12675_21(.douta(w_n12675_21[0]),.doutb(w_n12675_21[1]),.doutc(w_n12675_21[2]),.din(w_n12675_6[2]));
	jspl3 jspl3_w_n12675_22(.douta(w_n12675_22[0]),.doutb(w_n12675_22[1]),.doutc(w_n12675_22[2]),.din(w_n12675_7[0]));
	jspl3 jspl3_w_n12675_23(.douta(w_n12675_23[0]),.doutb(w_n12675_23[1]),.doutc(w_n12675_23[2]),.din(w_n12675_7[1]));
	jspl jspl_w_n12675_24(.douta(w_n12675_24[0]),.doutb(w_n12675_24[1]),.din(w_n12675_7[2]));
	jspl jspl_w_n12679_0(.douta(w_n12679_0[0]),.doutb(w_n12679_0[1]),.din(n12679));
	jspl3 jspl3_w_n12681_0(.douta(w_n12681_0[0]),.doutb(w_n12681_0[1]),.doutc(w_n12681_0[2]),.din(n12681));
	jspl jspl_w_n12681_1(.douta(w_n12681_1[0]),.doutb(w_n12681_1[1]),.din(w_n12681_0[0]));
	jspl3 jspl3_w_n12682_0(.douta(w_n12682_0[0]),.doutb(w_n12682_0[1]),.doutc(w_n12682_0[2]),.din(n12682));
	jspl3 jspl3_w_n12686_0(.douta(w_n12686_0[0]),.doutb(w_n12686_0[1]),.doutc(w_n12686_0[2]),.din(n12686));
	jspl jspl_w_n12687_0(.douta(w_n12687_0[0]),.doutb(w_n12687_0[1]),.din(n12687));
	jspl jspl_w_n12688_0(.douta(w_n12688_0[0]),.doutb(w_n12688_0[1]),.din(n12688));
	jspl jspl_w_n12689_0(.douta(w_n12689_0[0]),.doutb(w_n12689_0[1]),.din(n12689));
	jspl jspl_w_n12691_0(.douta(w_n12691_0[0]),.doutb(w_n12691_0[1]),.din(n12691));
	jspl jspl_w_n12693_0(.douta(w_n12693_0[0]),.doutb(w_n12693_0[1]),.din(n12693));
	jspl jspl_w_n12695_0(.douta(w_n12695_0[0]),.doutb(w_n12695_0[1]),.din(n12695));
	jspl jspl_w_n12698_0(.douta(w_n12698_0[0]),.doutb(w_n12698_0[1]),.din(n12698));
	jspl jspl_w_n12703_0(.douta(w_n12703_0[0]),.doutb(w_n12703_0[1]),.din(n12703));
	jspl3 jspl3_w_n12705_0(.douta(w_n12705_0[0]),.doutb(w_n12705_0[1]),.doutc(w_n12705_0[2]),.din(n12705));
	jspl jspl_w_n12706_0(.douta(w_n12706_0[0]),.doutb(w_n12706_0[1]),.din(n12706));
	jspl jspl_w_n12710_0(.douta(w_n12710_0[0]),.doutb(w_n12710_0[1]),.din(n12710));
	jspl jspl_w_n12711_0(.douta(w_n12711_0[0]),.doutb(w_n12711_0[1]),.din(n12711));
	jspl jspl_w_n12713_0(.douta(w_n12713_0[0]),.doutb(w_n12713_0[1]),.din(n12713));
	jspl jspl_w_n12717_0(.douta(w_n12717_0[0]),.doutb(w_n12717_0[1]),.din(n12717));
	jspl jspl_w_n12719_0(.douta(w_n12719_0[0]),.doutb(w_n12719_0[1]),.din(n12719));
	jspl jspl_w_n12720_0(.douta(w_n12720_0[0]),.doutb(w_n12720_0[1]),.din(n12720));
	jspl3 jspl3_w_n12721_0(.douta(w_n12721_0[0]),.doutb(w_n12721_0[1]),.doutc(w_n12721_0[2]),.din(n12721));
	jspl jspl_w_n12722_0(.douta(w_n12722_0[0]),.doutb(w_n12722_0[1]),.din(n12722));
	jspl jspl_w_n12726_0(.douta(w_n12726_0[0]),.doutb(w_n12726_0[1]),.din(n12726));
	jspl jspl_w_n12728_0(.douta(w_n12728_0[0]),.doutb(w_n12728_0[1]),.din(n12728));
	jspl jspl_w_n12730_0(.douta(w_n12730_0[0]),.doutb(w_n12730_0[1]),.din(n12730));
	jspl jspl_w_n12732_0(.douta(w_n12732_0[0]),.doutb(w_n12732_0[1]),.din(n12732));
	jspl jspl_w_n12735_0(.douta(w_n12735_0[0]),.doutb(w_n12735_0[1]),.din(n12735));
	jspl jspl_w_n12741_0(.douta(w_n12741_0[0]),.doutb(w_n12741_0[1]),.din(n12741));
	jspl3 jspl3_w_n12743_0(.douta(w_n12743_0[0]),.doutb(w_n12743_0[1]),.doutc(w_n12743_0[2]),.din(n12743));
	jspl jspl_w_n12744_0(.douta(w_n12744_0[0]),.doutb(w_n12744_0[1]),.din(n12744));
	jspl jspl_w_n12749_0(.douta(w_n12749_0[0]),.doutb(w_n12749_0[1]),.din(n12749));
	jspl jspl_w_n12751_0(.douta(w_n12751_0[0]),.doutb(w_n12751_0[1]),.din(n12751));
	jspl jspl_w_n12753_0(.douta(w_n12753_0[0]),.doutb(w_n12753_0[1]),.din(n12753));
	jspl jspl_w_n12757_0(.douta(w_n12757_0[0]),.doutb(w_n12757_0[1]),.din(n12757));
	jspl jspl_w_n12759_0(.douta(w_n12759_0[0]),.doutb(w_n12759_0[1]),.din(n12759));
	jspl jspl_w_n12760_0(.douta(w_n12760_0[0]),.doutb(w_n12760_0[1]),.din(n12760));
	jspl3 jspl3_w_n12761_0(.douta(w_n12761_0[0]),.doutb(w_n12761_0[1]),.doutc(w_n12761_0[2]),.din(n12761));
	jspl jspl_w_n12762_0(.douta(w_n12762_0[0]),.doutb(w_n12762_0[1]),.din(n12762));
	jspl jspl_w_n12768_0(.douta(w_n12768_0[0]),.doutb(w_n12768_0[1]),.din(n12768));
	jspl jspl_w_n12769_0(.douta(w_n12769_0[0]),.doutb(w_n12769_0[1]),.din(n12769));
	jspl jspl_w_n12771_0(.douta(w_n12771_0[0]),.doutb(w_n12771_0[1]),.din(n12771));
	jspl jspl_w_n12773_0(.douta(w_n12773_0[0]),.doutb(w_n12773_0[1]),.din(n12773));
	jspl jspl_w_n12775_0(.douta(w_n12775_0[0]),.doutb(w_n12775_0[1]),.din(n12775));
	jspl jspl_w_n12781_0(.douta(w_n12781_0[0]),.doutb(w_n12781_0[1]),.din(n12781));
	jspl jspl_w_n12783_0(.douta(w_n12783_0[0]),.doutb(w_n12783_0[1]),.din(n12783));
	jspl3 jspl3_w_n12784_0(.douta(w_n12784_0[0]),.doutb(w_n12784_0[1]),.doutc(w_n12784_0[2]),.din(n12784));
	jspl jspl_w_n12787_0(.douta(w_n12787_0[0]),.doutb(w_n12787_0[1]),.din(n12787));
	jspl jspl_w_n12788_0(.douta(w_n12788_0[0]),.doutb(w_n12788_0[1]),.din(n12788));
	jspl3 jspl3_w_n12789_0(.douta(w_n12789_0[0]),.doutb(w_n12789_0[1]),.doutc(w_n12789_0[2]),.din(n12789));
	jspl jspl_w_n12791_0(.douta(w_n12791_0[0]),.doutb(w_n12791_0[1]),.din(n12791));
	jspl jspl_w_n12795_0(.douta(w_n12795_0[0]),.doutb(w_n12795_0[1]),.din(n12795));
	jspl jspl_w_n12797_0(.douta(w_n12797_0[0]),.doutb(w_n12797_0[1]),.din(n12797));
	jspl jspl_w_n12798_0(.douta(w_n12798_0[0]),.doutb(w_n12798_0[1]),.din(n12798));
	jspl3 jspl3_w_n12799_0(.douta(w_n12799_0[0]),.doutb(w_n12799_0[1]),.doutc(w_n12799_0[2]),.din(n12799));
	jspl jspl_w_n12800_0(.douta(w_n12800_0[0]),.doutb(w_n12800_0[1]),.din(n12800));
	jspl jspl_w_n12803_0(.douta(w_n12803_0[0]),.doutb(w_n12803_0[1]),.din(n12803));
	jspl jspl_w_n12809_0(.douta(w_n12809_0[0]),.doutb(w_n12809_0[1]),.din(n12809));
	jspl jspl_w_n12810_0(.douta(w_n12810_0[0]),.doutb(w_n12810_0[1]),.din(n12810));
	jspl jspl_w_n12812_0(.douta(w_n12812_0[0]),.doutb(w_n12812_0[1]),.din(n12812));
	jspl jspl_w_n12814_0(.douta(w_n12814_0[0]),.doutb(w_n12814_0[1]),.din(n12814));
	jspl jspl_w_n12816_0(.douta(w_n12816_0[0]),.doutb(w_n12816_0[1]),.din(n12816));
	jspl jspl_w_n12822_0(.douta(w_n12822_0[0]),.doutb(w_n12822_0[1]),.din(n12822));
	jspl jspl_w_n12824_0(.douta(w_n12824_0[0]),.doutb(w_n12824_0[1]),.din(n12824));
	jspl3 jspl3_w_n12825_0(.douta(w_n12825_0[0]),.doutb(w_n12825_0[1]),.doutc(w_n12825_0[2]),.din(n12825));
	jspl jspl_w_n12828_0(.douta(w_n12828_0[0]),.doutb(w_n12828_0[1]),.din(n12828));
	jspl jspl_w_n12829_0(.douta(w_n12829_0[0]),.doutb(w_n12829_0[1]),.din(n12829));
	jspl3 jspl3_w_n12830_0(.douta(w_n12830_0[0]),.doutb(w_n12830_0[1]),.doutc(w_n12830_0[2]),.din(n12830));
	jspl jspl_w_n12832_0(.douta(w_n12832_0[0]),.doutb(w_n12832_0[1]),.din(n12832));
	jspl jspl_w_n12836_0(.douta(w_n12836_0[0]),.doutb(w_n12836_0[1]),.din(n12836));
	jspl jspl_w_n12838_0(.douta(w_n12838_0[0]),.doutb(w_n12838_0[1]),.din(n12838));
	jspl jspl_w_n12839_0(.douta(w_n12839_0[0]),.doutb(w_n12839_0[1]),.din(n12839));
	jspl3 jspl3_w_n12840_0(.douta(w_n12840_0[0]),.doutb(w_n12840_0[1]),.doutc(w_n12840_0[2]),.din(n12840));
	jspl jspl_w_n12841_0(.douta(w_n12841_0[0]),.doutb(w_n12841_0[1]),.din(n12841));
	jspl jspl_w_n12844_0(.douta(w_n12844_0[0]),.doutb(w_n12844_0[1]),.din(n12844));
	jspl jspl_w_n12850_0(.douta(w_n12850_0[0]),.doutb(w_n12850_0[1]),.din(n12850));
	jspl jspl_w_n12851_0(.douta(w_n12851_0[0]),.doutb(w_n12851_0[1]),.din(n12851));
	jspl jspl_w_n12853_0(.douta(w_n12853_0[0]),.doutb(w_n12853_0[1]),.din(n12853));
	jspl jspl_w_n12855_0(.douta(w_n12855_0[0]),.doutb(w_n12855_0[1]),.din(n12855));
	jspl jspl_w_n12857_0(.douta(w_n12857_0[0]),.doutb(w_n12857_0[1]),.din(n12857));
	jspl jspl_w_n12863_0(.douta(w_n12863_0[0]),.doutb(w_n12863_0[1]),.din(n12863));
	jspl jspl_w_n12865_0(.douta(w_n12865_0[0]),.doutb(w_n12865_0[1]),.din(n12865));
	jspl3 jspl3_w_n12866_0(.douta(w_n12866_0[0]),.doutb(w_n12866_0[1]),.doutc(w_n12866_0[2]),.din(n12866));
	jspl jspl_w_n12869_0(.douta(w_n12869_0[0]),.doutb(w_n12869_0[1]),.din(n12869));
	jspl jspl_w_n12870_0(.douta(w_n12870_0[0]),.doutb(w_n12870_0[1]),.din(n12870));
	jspl3 jspl3_w_n12871_0(.douta(w_n12871_0[0]),.doutb(w_n12871_0[1]),.doutc(w_n12871_0[2]),.din(n12871));
	jspl jspl_w_n12873_0(.douta(w_n12873_0[0]),.doutb(w_n12873_0[1]),.din(n12873));
	jspl jspl_w_n12877_0(.douta(w_n12877_0[0]),.doutb(w_n12877_0[1]),.din(n12877));
	jspl jspl_w_n12879_0(.douta(w_n12879_0[0]),.doutb(w_n12879_0[1]),.din(n12879));
	jspl jspl_w_n12880_0(.douta(w_n12880_0[0]),.doutb(w_n12880_0[1]),.din(n12880));
	jspl3 jspl3_w_n12881_0(.douta(w_n12881_0[0]),.doutb(w_n12881_0[1]),.doutc(w_n12881_0[2]),.din(n12881));
	jspl jspl_w_n12882_0(.douta(w_n12882_0[0]),.doutb(w_n12882_0[1]),.din(n12882));
	jspl jspl_w_n12885_0(.douta(w_n12885_0[0]),.doutb(w_n12885_0[1]),.din(n12885));
	jspl jspl_w_n12891_0(.douta(w_n12891_0[0]),.doutb(w_n12891_0[1]),.din(n12891));
	jspl jspl_w_n12892_0(.douta(w_n12892_0[0]),.doutb(w_n12892_0[1]),.din(n12892));
	jspl jspl_w_n12894_0(.douta(w_n12894_0[0]),.doutb(w_n12894_0[1]),.din(n12894));
	jspl jspl_w_n12896_0(.douta(w_n12896_0[0]),.doutb(w_n12896_0[1]),.din(n12896));
	jspl jspl_w_n12898_0(.douta(w_n12898_0[0]),.doutb(w_n12898_0[1]),.din(n12898));
	jspl jspl_w_n12904_0(.douta(w_n12904_0[0]),.doutb(w_n12904_0[1]),.din(n12904));
	jspl jspl_w_n12906_0(.douta(w_n12906_0[0]),.doutb(w_n12906_0[1]),.din(n12906));
	jspl3 jspl3_w_n12907_0(.douta(w_n12907_0[0]),.doutb(w_n12907_0[1]),.doutc(w_n12907_0[2]),.din(n12907));
	jspl jspl_w_n12910_0(.douta(w_n12910_0[0]),.doutb(w_n12910_0[1]),.din(n12910));
	jspl jspl_w_n12911_0(.douta(w_n12911_0[0]),.doutb(w_n12911_0[1]),.din(n12911));
	jspl3 jspl3_w_n12912_0(.douta(w_n12912_0[0]),.doutb(w_n12912_0[1]),.doutc(w_n12912_0[2]),.din(n12912));
	jspl jspl_w_n12914_0(.douta(w_n12914_0[0]),.doutb(w_n12914_0[1]),.din(n12914));
	jspl jspl_w_n12918_0(.douta(w_n12918_0[0]),.doutb(w_n12918_0[1]),.din(n12918));
	jspl jspl_w_n12920_0(.douta(w_n12920_0[0]),.doutb(w_n12920_0[1]),.din(n12920));
	jspl jspl_w_n12921_0(.douta(w_n12921_0[0]),.doutb(w_n12921_0[1]),.din(n12921));
	jspl3 jspl3_w_n12922_0(.douta(w_n12922_0[0]),.doutb(w_n12922_0[1]),.doutc(w_n12922_0[2]),.din(n12922));
	jspl jspl_w_n12923_0(.douta(w_n12923_0[0]),.doutb(w_n12923_0[1]),.din(n12923));
	jspl jspl_w_n12926_0(.douta(w_n12926_0[0]),.doutb(w_n12926_0[1]),.din(n12926));
	jspl jspl_w_n12932_0(.douta(w_n12932_0[0]),.doutb(w_n12932_0[1]),.din(n12932));
	jspl jspl_w_n12933_0(.douta(w_n12933_0[0]),.doutb(w_n12933_0[1]),.din(n12933));
	jspl jspl_w_n12935_0(.douta(w_n12935_0[0]),.doutb(w_n12935_0[1]),.din(n12935));
	jspl jspl_w_n12937_0(.douta(w_n12937_0[0]),.doutb(w_n12937_0[1]),.din(n12937));
	jspl jspl_w_n12939_0(.douta(w_n12939_0[0]),.doutb(w_n12939_0[1]),.din(n12939));
	jspl jspl_w_n12945_0(.douta(w_n12945_0[0]),.doutb(w_n12945_0[1]),.din(n12945));
	jspl jspl_w_n12947_0(.douta(w_n12947_0[0]),.doutb(w_n12947_0[1]),.din(n12947));
	jspl3 jspl3_w_n12948_0(.douta(w_n12948_0[0]),.doutb(w_n12948_0[1]),.doutc(w_n12948_0[2]),.din(n12948));
	jspl jspl_w_n12951_0(.douta(w_n12951_0[0]),.doutb(w_n12951_0[1]),.din(n12951));
	jspl jspl_w_n12952_0(.douta(w_n12952_0[0]),.doutb(w_n12952_0[1]),.din(n12952));
	jspl3 jspl3_w_n12953_0(.douta(w_n12953_0[0]),.doutb(w_n12953_0[1]),.doutc(w_n12953_0[2]),.din(n12953));
	jspl jspl_w_n12955_0(.douta(w_n12955_0[0]),.doutb(w_n12955_0[1]),.din(n12955));
	jspl jspl_w_n12959_0(.douta(w_n12959_0[0]),.doutb(w_n12959_0[1]),.din(n12959));
	jspl jspl_w_n12961_0(.douta(w_n12961_0[0]),.doutb(w_n12961_0[1]),.din(n12961));
	jspl jspl_w_n12962_0(.douta(w_n12962_0[0]),.doutb(w_n12962_0[1]),.din(n12962));
	jspl3 jspl3_w_n12963_0(.douta(w_n12963_0[0]),.doutb(w_n12963_0[1]),.doutc(w_n12963_0[2]),.din(n12963));
	jspl jspl_w_n12964_0(.douta(w_n12964_0[0]),.doutb(w_n12964_0[1]),.din(n12964));
	jspl jspl_w_n12967_0(.douta(w_n12967_0[0]),.doutb(w_n12967_0[1]),.din(n12967));
	jspl jspl_w_n12973_0(.douta(w_n12973_0[0]),.doutb(w_n12973_0[1]),.din(n12973));
	jspl jspl_w_n12974_0(.douta(w_n12974_0[0]),.doutb(w_n12974_0[1]),.din(n12974));
	jspl jspl_w_n12976_0(.douta(w_n12976_0[0]),.doutb(w_n12976_0[1]),.din(n12976));
	jspl jspl_w_n12978_0(.douta(w_n12978_0[0]),.doutb(w_n12978_0[1]),.din(n12978));
	jspl jspl_w_n12980_0(.douta(w_n12980_0[0]),.doutb(w_n12980_0[1]),.din(n12980));
	jspl jspl_w_n12986_0(.douta(w_n12986_0[0]),.doutb(w_n12986_0[1]),.din(n12986));
	jspl jspl_w_n12988_0(.douta(w_n12988_0[0]),.doutb(w_n12988_0[1]),.din(n12988));
	jspl3 jspl3_w_n12989_0(.douta(w_n12989_0[0]),.doutb(w_n12989_0[1]),.doutc(w_n12989_0[2]),.din(n12989));
	jspl jspl_w_n12992_0(.douta(w_n12992_0[0]),.doutb(w_n12992_0[1]),.din(n12992));
	jspl jspl_w_n12993_0(.douta(w_n12993_0[0]),.doutb(w_n12993_0[1]),.din(n12993));
	jspl3 jspl3_w_n12994_0(.douta(w_n12994_0[0]),.doutb(w_n12994_0[1]),.doutc(w_n12994_0[2]),.din(n12994));
	jspl jspl_w_n12996_0(.douta(w_n12996_0[0]),.doutb(w_n12996_0[1]),.din(n12996));
	jspl jspl_w_n12998_0(.douta(w_n12998_0[0]),.doutb(w_n12998_0[1]),.din(n12998));
	jspl jspl_w_n13000_0(.douta(w_n13000_0[0]),.doutb(w_n13000_0[1]),.din(n13000));
	jspl jspl_w_n13006_0(.douta(w_n13006_0[0]),.doutb(w_n13006_0[1]),.din(n13006));
	jspl3 jspl3_w_n13008_0(.douta(w_n13008_0[0]),.doutb(w_n13008_0[1]),.doutc(w_n13008_0[2]),.din(n13008));
	jspl jspl_w_n13009_0(.douta(w_n13009_0[0]),.doutb(w_n13009_0[1]),.din(n13009));
	jspl jspl_w_n13011_0(.douta(w_n13011_0[0]),.doutb(w_n13011_0[1]),.din(n13011));
	jspl jspl_w_n13013_0(.douta(w_n13013_0[0]),.doutb(w_n13013_0[1]),.din(n13013));
	jspl jspl_w_n13017_0(.douta(w_n13017_0[0]),.doutb(w_n13017_0[1]),.din(n13017));
	jspl jspl_w_n13019_0(.douta(w_n13019_0[0]),.doutb(w_n13019_0[1]),.din(n13019));
	jspl jspl_w_n13020_0(.douta(w_n13020_0[0]),.doutb(w_n13020_0[1]),.din(n13020));
	jspl jspl_w_n13021_0(.douta(w_n13021_0[0]),.doutb(w_n13021_0[1]),.din(n13021));
	jspl3 jspl3_w_n13022_0(.douta(w_n13022_0[0]),.doutb(w_n13022_0[1]),.doutc(w_n13022_0[2]),.din(n13022));
	jspl jspl_w_n13025_0(.douta(w_n13025_0[0]),.doutb(w_n13025_0[1]),.din(n13025));
	jspl jspl_w_n13026_0(.douta(w_n13026_0[0]),.doutb(w_n13026_0[1]),.din(n13026));
	jspl3 jspl3_w_n13027_0(.douta(w_n13027_0[0]),.doutb(w_n13027_0[1]),.doutc(w_n13027_0[2]),.din(n13027));
	jspl jspl_w_n13029_0(.douta(w_n13029_0[0]),.doutb(w_n13029_0[1]),.din(n13029));
	jspl jspl_w_n13033_0(.douta(w_n13033_0[0]),.doutb(w_n13033_0[1]),.din(n13033));
	jspl jspl_w_n13035_0(.douta(w_n13035_0[0]),.doutb(w_n13035_0[1]),.din(n13035));
	jspl jspl_w_n13036_0(.douta(w_n13036_0[0]),.doutb(w_n13036_0[1]),.din(n13036));
	jspl3 jspl3_w_n13037_0(.douta(w_n13037_0[0]),.doutb(w_n13037_0[1]),.doutc(w_n13037_0[2]),.din(n13037));
	jspl jspl_w_n13038_0(.douta(w_n13038_0[0]),.doutb(w_n13038_0[1]),.din(n13038));
	jspl jspl_w_n13041_0(.douta(w_n13041_0[0]),.doutb(w_n13041_0[1]),.din(n13041));
	jspl jspl_w_n13047_0(.douta(w_n13047_0[0]),.doutb(w_n13047_0[1]),.din(n13047));
	jspl jspl_w_n13048_0(.douta(w_n13048_0[0]),.doutb(w_n13048_0[1]),.din(n13048));
	jspl jspl_w_n13050_0(.douta(w_n13050_0[0]),.doutb(w_n13050_0[1]),.din(n13050));
	jspl jspl_w_n13052_0(.douta(w_n13052_0[0]),.doutb(w_n13052_0[1]),.din(n13052));
	jspl jspl_w_n13054_0(.douta(w_n13054_0[0]),.doutb(w_n13054_0[1]),.din(n13054));
	jspl jspl_w_n13060_0(.douta(w_n13060_0[0]),.doutb(w_n13060_0[1]),.din(n13060));
	jspl jspl_w_n13062_0(.douta(w_n13062_0[0]),.doutb(w_n13062_0[1]),.din(n13062));
	jspl3 jspl3_w_n13063_0(.douta(w_n13063_0[0]),.doutb(w_n13063_0[1]),.doutc(w_n13063_0[2]),.din(n13063));
	jspl jspl_w_n13066_0(.douta(w_n13066_0[0]),.doutb(w_n13066_0[1]),.din(n13066));
	jspl jspl_w_n13067_0(.douta(w_n13067_0[0]),.doutb(w_n13067_0[1]),.din(n13067));
	jspl3 jspl3_w_n13068_0(.douta(w_n13068_0[0]),.doutb(w_n13068_0[1]),.doutc(w_n13068_0[2]),.din(n13068));
	jspl jspl_w_n13070_0(.douta(w_n13070_0[0]),.doutb(w_n13070_0[1]),.din(n13070));
	jspl jspl_w_n13074_0(.douta(w_n13074_0[0]),.doutb(w_n13074_0[1]),.din(n13074));
	jspl jspl_w_n13076_0(.douta(w_n13076_0[0]),.doutb(w_n13076_0[1]),.din(n13076));
	jspl jspl_w_n13077_0(.douta(w_n13077_0[0]),.doutb(w_n13077_0[1]),.din(n13077));
	jspl3 jspl3_w_n13078_0(.douta(w_n13078_0[0]),.doutb(w_n13078_0[1]),.doutc(w_n13078_0[2]),.din(n13078));
	jspl jspl_w_n13079_0(.douta(w_n13079_0[0]),.doutb(w_n13079_0[1]),.din(n13079));
	jspl jspl_w_n13082_0(.douta(w_n13082_0[0]),.doutb(w_n13082_0[1]),.din(n13082));
	jspl jspl_w_n13088_0(.douta(w_n13088_0[0]),.doutb(w_n13088_0[1]),.din(n13088));
	jspl jspl_w_n13089_0(.douta(w_n13089_0[0]),.doutb(w_n13089_0[1]),.din(n13089));
	jspl jspl_w_n13091_0(.douta(w_n13091_0[0]),.doutb(w_n13091_0[1]),.din(n13091));
	jspl jspl_w_n13093_0(.douta(w_n13093_0[0]),.doutb(w_n13093_0[1]),.din(n13093));
	jspl jspl_w_n13095_0(.douta(w_n13095_0[0]),.doutb(w_n13095_0[1]),.din(n13095));
	jspl jspl_w_n13101_0(.douta(w_n13101_0[0]),.doutb(w_n13101_0[1]),.din(n13101));
	jspl jspl_w_n13103_0(.douta(w_n13103_0[0]),.doutb(w_n13103_0[1]),.din(n13103));
	jspl3 jspl3_w_n13104_0(.douta(w_n13104_0[0]),.doutb(w_n13104_0[1]),.doutc(w_n13104_0[2]),.din(n13104));
	jspl jspl_w_n13107_0(.douta(w_n13107_0[0]),.doutb(w_n13107_0[1]),.din(n13107));
	jspl jspl_w_n13108_0(.douta(w_n13108_0[0]),.doutb(w_n13108_0[1]),.din(n13108));
	jspl3 jspl3_w_n13109_0(.douta(w_n13109_0[0]),.doutb(w_n13109_0[1]),.doutc(w_n13109_0[2]),.din(n13109));
	jspl jspl_w_n13111_0(.douta(w_n13111_0[0]),.doutb(w_n13111_0[1]),.din(n13111));
	jspl jspl_w_n13115_0(.douta(w_n13115_0[0]),.doutb(w_n13115_0[1]),.din(n13115));
	jspl jspl_w_n13117_0(.douta(w_n13117_0[0]),.doutb(w_n13117_0[1]),.din(n13117));
	jspl jspl_w_n13118_0(.douta(w_n13118_0[0]),.doutb(w_n13118_0[1]),.din(n13118));
	jspl3 jspl3_w_n13119_0(.douta(w_n13119_0[0]),.doutb(w_n13119_0[1]),.doutc(w_n13119_0[2]),.din(n13119));
	jspl jspl_w_n13120_0(.douta(w_n13120_0[0]),.doutb(w_n13120_0[1]),.din(n13120));
	jspl jspl_w_n13123_0(.douta(w_n13123_0[0]),.doutb(w_n13123_0[1]),.din(n13123));
	jspl jspl_w_n13129_0(.douta(w_n13129_0[0]),.doutb(w_n13129_0[1]),.din(n13129));
	jspl jspl_w_n13130_0(.douta(w_n13130_0[0]),.doutb(w_n13130_0[1]),.din(n13130));
	jspl jspl_w_n13132_0(.douta(w_n13132_0[0]),.doutb(w_n13132_0[1]),.din(n13132));
	jspl jspl_w_n13134_0(.douta(w_n13134_0[0]),.doutb(w_n13134_0[1]),.din(n13134));
	jspl jspl_w_n13136_0(.douta(w_n13136_0[0]),.doutb(w_n13136_0[1]),.din(n13136));
	jspl jspl_w_n13142_0(.douta(w_n13142_0[0]),.doutb(w_n13142_0[1]),.din(n13142));
	jspl3 jspl3_w_n13144_0(.douta(w_n13144_0[0]),.doutb(w_n13144_0[1]),.doutc(w_n13144_0[2]),.din(n13144));
	jspl jspl_w_n13149_0(.douta(w_n13149_0[0]),.doutb(w_n13149_0[1]),.din(n13149));
	jspl3 jspl3_w_n13151_0(.douta(w_n13151_0[0]),.doutb(w_n13151_0[1]),.doutc(w_n13151_0[2]),.din(n13151));
	jspl3 jspl3_w_n13155_0(.douta(w_n13155_0[0]),.doutb(w_n13155_0[1]),.doutc(w_n13155_0[2]),.din(n13155));
	jspl jspl_w_n13156_0(.douta(w_n13156_0[0]),.doutb(w_n13156_0[1]),.din(n13156));
	jspl jspl_w_n13161_0(.douta(w_n13161_0[0]),.doutb(w_n13161_0[1]),.din(n13161));
	jspl3 jspl3_w_n13162_0(.douta(w_n13162_0[0]),.doutb(w_n13162_0[1]),.doutc(w_n13162_0[2]),.din(n13162));
	jspl jspl_w_n13167_0(.douta(w_n13167_0[0]),.doutb(w_n13167_0[1]),.din(n13167));
	jspl jspl_w_n13175_0(.douta(w_n13175_0[0]),.doutb(w_n13175_0[1]),.din(n13175));
	jspl3 jspl3_w_n13177_0(.douta(w_n13177_0[0]),.doutb(w_n13177_0[1]),.doutc(w_n13177_0[2]),.din(n13177));
	jspl jspl_w_n13177_1(.douta(w_n13177_1[0]),.doutb(w_n13177_1[1]),.din(w_n13177_0[0]));
	jspl jspl_w_n13178_0(.douta(w_n13178_0[0]),.doutb(w_n13178_0[1]),.din(n13178));
	jspl3 jspl3_w_n13181_0(.douta(w_n13181_0[0]),.doutb(w_n13181_0[1]),.doutc(w_n13181_0[2]),.din(n13181));
	jspl jspl_w_n13182_0(.douta(w_n13182_0[0]),.doutb(w_n13182_0[1]),.din(n13182));
	jspl jspl_w_n13183_0(.douta(w_n13183_0[0]),.doutb(w_n13183_0[1]),.din(n13183));
	jspl jspl_w_n13184_0(.douta(w_n13184_0[0]),.doutb(w_n13184_0[1]),.din(n13184));
	jspl jspl_w_n13186_0(.douta(w_n13186_0[0]),.doutb(w_n13186_0[1]),.din(n13186));
	jspl jspl_w_n13188_0(.douta(w_n13188_0[0]),.doutb(w_n13188_0[1]),.din(n13188));
	jspl jspl_w_n13190_0(.douta(w_n13190_0[0]),.doutb(w_n13190_0[1]),.din(n13190));
	jspl jspl_w_n13199_0(.douta(w_n13199_0[0]),.doutb(w_n13199_0[1]),.din(n13199));
	jspl3 jspl3_w_n13201_0(.douta(w_n13201_0[0]),.doutb(w_n13201_0[1]),.doutc(w_n13201_0[2]),.din(n13201));
	jspl jspl_w_n13202_0(.douta(w_n13202_0[0]),.doutb(w_n13202_0[1]),.din(n13202));
	jspl jspl_w_n13206_0(.douta(w_n13206_0[0]),.doutb(w_n13206_0[1]),.din(n13206));
	jspl jspl_w_n13208_0(.douta(w_n13208_0[0]),.doutb(w_n13208_0[1]),.din(n13208));
	jspl jspl_w_n13210_0(.douta(w_n13210_0[0]),.doutb(w_n13210_0[1]),.din(n13210));
	jspl jspl_w_n13215_0(.douta(w_n13215_0[0]),.doutb(w_n13215_0[1]),.din(n13215));
	jspl jspl_w_n13217_0(.douta(w_n13217_0[0]),.doutb(w_n13217_0[1]),.din(n13217));
	jspl jspl_w_n13218_0(.douta(w_n13218_0[0]),.doutb(w_n13218_0[1]),.din(n13218));
	jspl3 jspl3_w_n13219_0(.douta(w_n13219_0[0]),.doutb(w_n13219_0[1]),.doutc(w_n13219_0[2]),.din(n13219));
	jspl jspl_w_n13220_0(.douta(w_n13220_0[0]),.doutb(w_n13220_0[1]),.din(n13220));
	jspl jspl_w_n13225_0(.douta(w_n13225_0[0]),.doutb(w_n13225_0[1]),.din(n13225));
	jspl jspl_w_n13226_0(.douta(w_n13226_0[0]),.doutb(w_n13226_0[1]),.din(n13226));
	jspl jspl_w_n13228_0(.douta(w_n13228_0[0]),.doutb(w_n13228_0[1]),.din(n13228));
	jspl jspl_w_n13230_0(.douta(w_n13230_0[0]),.doutb(w_n13230_0[1]),.din(n13230));
	jspl jspl_w_n13233_0(.douta(w_n13233_0[0]),.doutb(w_n13233_0[1]),.din(n13233));
	jspl jspl_w_n13239_0(.douta(w_n13239_0[0]),.doutb(w_n13239_0[1]),.din(n13239));
	jspl3 jspl3_w_n13241_0(.douta(w_n13241_0[0]),.doutb(w_n13241_0[1]),.doutc(w_n13241_0[2]),.din(n13241));
	jspl jspl_w_n13242_0(.douta(w_n13242_0[0]),.doutb(w_n13242_0[1]),.din(n13242));
	jspl jspl_w_n13246_0(.douta(w_n13246_0[0]),.doutb(w_n13246_0[1]),.din(n13246));
	jspl jspl_w_n13247_0(.douta(w_n13247_0[0]),.doutb(w_n13247_0[1]),.din(n13247));
	jspl jspl_w_n13249_0(.douta(w_n13249_0[0]),.doutb(w_n13249_0[1]),.din(n13249));
	jspl jspl_w_n13254_0(.douta(w_n13254_0[0]),.doutb(w_n13254_0[1]),.din(n13254));
	jspl jspl_w_n13256_0(.douta(w_n13256_0[0]),.doutb(w_n13256_0[1]),.din(n13256));
	jspl jspl_w_n13257_0(.douta(w_n13257_0[0]),.doutb(w_n13257_0[1]),.din(n13257));
	jspl3 jspl3_w_n13258_0(.douta(w_n13258_0[0]),.doutb(w_n13258_0[1]),.doutc(w_n13258_0[2]),.din(n13258));
	jspl jspl_w_n13259_0(.douta(w_n13259_0[0]),.doutb(w_n13259_0[1]),.din(n13259));
	jspl jspl_w_n13263_0(.douta(w_n13263_0[0]),.doutb(w_n13263_0[1]),.din(n13263));
	jspl jspl_w_n13264_0(.douta(w_n13264_0[0]),.doutb(w_n13264_0[1]),.din(n13264));
	jspl jspl_w_n13266_0(.douta(w_n13266_0[0]),.doutb(w_n13266_0[1]),.din(n13266));
	jspl jspl_w_n13268_0(.douta(w_n13268_0[0]),.doutb(w_n13268_0[1]),.din(n13268));
	jspl jspl_w_n13271_0(.douta(w_n13271_0[0]),.doutb(w_n13271_0[1]),.din(n13271));
	jspl jspl_w_n13277_0(.douta(w_n13277_0[0]),.doutb(w_n13277_0[1]),.din(n13277));
	jspl jspl_w_n13279_0(.douta(w_n13279_0[0]),.doutb(w_n13279_0[1]),.din(n13279));
	jspl3 jspl3_w_n13280_0(.douta(w_n13280_0[0]),.doutb(w_n13280_0[1]),.doutc(w_n13280_0[2]),.din(n13280));
	jspl jspl_w_n13284_0(.douta(w_n13284_0[0]),.doutb(w_n13284_0[1]),.din(n13284));
	jspl jspl_w_n13285_0(.douta(w_n13285_0[0]),.doutb(w_n13285_0[1]),.din(n13285));
	jspl3 jspl3_w_n13286_0(.douta(w_n13286_0[0]),.doutb(w_n13286_0[1]),.doutc(w_n13286_0[2]),.din(n13286));
	jspl jspl_w_n13288_0(.douta(w_n13288_0[0]),.doutb(w_n13288_0[1]),.din(n13288));
	jspl jspl_w_n13293_0(.douta(w_n13293_0[0]),.doutb(w_n13293_0[1]),.din(n13293));
	jspl jspl_w_n13295_0(.douta(w_n13295_0[0]),.doutb(w_n13295_0[1]),.din(n13295));
	jspl jspl_w_n13296_0(.douta(w_n13296_0[0]),.doutb(w_n13296_0[1]),.din(n13296));
	jspl3 jspl3_w_n13297_0(.douta(w_n13297_0[0]),.doutb(w_n13297_0[1]),.doutc(w_n13297_0[2]),.din(n13297));
	jspl jspl_w_n13298_0(.douta(w_n13298_0[0]),.doutb(w_n13298_0[1]),.din(n13298));
	jspl jspl_w_n13302_0(.douta(w_n13302_0[0]),.doutb(w_n13302_0[1]),.din(n13302));
	jspl jspl_w_n13308_0(.douta(w_n13308_0[0]),.doutb(w_n13308_0[1]),.din(n13308));
	jspl jspl_w_n13309_0(.douta(w_n13309_0[0]),.doutb(w_n13309_0[1]),.din(n13309));
	jspl jspl_w_n13311_0(.douta(w_n13311_0[0]),.doutb(w_n13311_0[1]),.din(n13311));
	jspl jspl_w_n13313_0(.douta(w_n13313_0[0]),.doutb(w_n13313_0[1]),.din(n13313));
	jspl jspl_w_n13316_0(.douta(w_n13316_0[0]),.doutb(w_n13316_0[1]),.din(n13316));
	jspl jspl_w_n13322_0(.douta(w_n13322_0[0]),.doutb(w_n13322_0[1]),.din(n13322));
	jspl jspl_w_n13324_0(.douta(w_n13324_0[0]),.doutb(w_n13324_0[1]),.din(n13324));
	jspl3 jspl3_w_n13325_0(.douta(w_n13325_0[0]),.doutb(w_n13325_0[1]),.doutc(w_n13325_0[2]),.din(n13325));
	jspl jspl_w_n13329_0(.douta(w_n13329_0[0]),.doutb(w_n13329_0[1]),.din(n13329));
	jspl jspl_w_n13330_0(.douta(w_n13330_0[0]),.doutb(w_n13330_0[1]),.din(n13330));
	jspl3 jspl3_w_n13331_0(.douta(w_n13331_0[0]),.doutb(w_n13331_0[1]),.doutc(w_n13331_0[2]),.din(n13331));
	jspl jspl_w_n13333_0(.douta(w_n13333_0[0]),.doutb(w_n13333_0[1]),.din(n13333));
	jspl jspl_w_n13338_0(.douta(w_n13338_0[0]),.doutb(w_n13338_0[1]),.din(n13338));
	jspl jspl_w_n13340_0(.douta(w_n13340_0[0]),.doutb(w_n13340_0[1]),.din(n13340));
	jspl jspl_w_n13341_0(.douta(w_n13341_0[0]),.doutb(w_n13341_0[1]),.din(n13341));
	jspl3 jspl3_w_n13342_0(.douta(w_n13342_0[0]),.doutb(w_n13342_0[1]),.doutc(w_n13342_0[2]),.din(n13342));
	jspl jspl_w_n13343_0(.douta(w_n13343_0[0]),.doutb(w_n13343_0[1]),.din(n13343));
	jspl jspl_w_n13347_0(.douta(w_n13347_0[0]),.doutb(w_n13347_0[1]),.din(n13347));
	jspl jspl_w_n13353_0(.douta(w_n13353_0[0]),.doutb(w_n13353_0[1]),.din(n13353));
	jspl jspl_w_n13354_0(.douta(w_n13354_0[0]),.doutb(w_n13354_0[1]),.din(n13354));
	jspl jspl_w_n13356_0(.douta(w_n13356_0[0]),.doutb(w_n13356_0[1]),.din(n13356));
	jspl jspl_w_n13358_0(.douta(w_n13358_0[0]),.doutb(w_n13358_0[1]),.din(n13358));
	jspl jspl_w_n13361_0(.douta(w_n13361_0[0]),.doutb(w_n13361_0[1]),.din(n13361));
	jspl jspl_w_n13367_0(.douta(w_n13367_0[0]),.doutb(w_n13367_0[1]),.din(n13367));
	jspl jspl_w_n13369_0(.douta(w_n13369_0[0]),.doutb(w_n13369_0[1]),.din(n13369));
	jspl3 jspl3_w_n13370_0(.douta(w_n13370_0[0]),.doutb(w_n13370_0[1]),.doutc(w_n13370_0[2]),.din(n13370));
	jspl jspl_w_n13374_0(.douta(w_n13374_0[0]),.doutb(w_n13374_0[1]),.din(n13374));
	jspl jspl_w_n13375_0(.douta(w_n13375_0[0]),.doutb(w_n13375_0[1]),.din(n13375));
	jspl3 jspl3_w_n13376_0(.douta(w_n13376_0[0]),.doutb(w_n13376_0[1]),.doutc(w_n13376_0[2]),.din(n13376));
	jspl jspl_w_n13378_0(.douta(w_n13378_0[0]),.doutb(w_n13378_0[1]),.din(n13378));
	jspl jspl_w_n13383_0(.douta(w_n13383_0[0]),.doutb(w_n13383_0[1]),.din(n13383));
	jspl jspl_w_n13385_0(.douta(w_n13385_0[0]),.doutb(w_n13385_0[1]),.din(n13385));
	jspl jspl_w_n13386_0(.douta(w_n13386_0[0]),.doutb(w_n13386_0[1]),.din(n13386));
	jspl3 jspl3_w_n13387_0(.douta(w_n13387_0[0]),.doutb(w_n13387_0[1]),.doutc(w_n13387_0[2]),.din(n13387));
	jspl jspl_w_n13388_0(.douta(w_n13388_0[0]),.doutb(w_n13388_0[1]),.din(n13388));
	jspl jspl_w_n13392_0(.douta(w_n13392_0[0]),.doutb(w_n13392_0[1]),.din(n13392));
	jspl jspl_w_n13398_0(.douta(w_n13398_0[0]),.doutb(w_n13398_0[1]),.din(n13398));
	jspl jspl_w_n13399_0(.douta(w_n13399_0[0]),.doutb(w_n13399_0[1]),.din(n13399));
	jspl jspl_w_n13401_0(.douta(w_n13401_0[0]),.doutb(w_n13401_0[1]),.din(n13401));
	jspl jspl_w_n13403_0(.douta(w_n13403_0[0]),.doutb(w_n13403_0[1]),.din(n13403));
	jspl jspl_w_n13406_0(.douta(w_n13406_0[0]),.doutb(w_n13406_0[1]),.din(n13406));
	jspl jspl_w_n13412_0(.douta(w_n13412_0[0]),.doutb(w_n13412_0[1]),.din(n13412));
	jspl jspl_w_n13414_0(.douta(w_n13414_0[0]),.doutb(w_n13414_0[1]),.din(n13414));
	jspl3 jspl3_w_n13415_0(.douta(w_n13415_0[0]),.doutb(w_n13415_0[1]),.doutc(w_n13415_0[2]),.din(n13415));
	jspl jspl_w_n13419_0(.douta(w_n13419_0[0]),.doutb(w_n13419_0[1]),.din(n13419));
	jspl jspl_w_n13420_0(.douta(w_n13420_0[0]),.doutb(w_n13420_0[1]),.din(n13420));
	jspl3 jspl3_w_n13421_0(.douta(w_n13421_0[0]),.doutb(w_n13421_0[1]),.doutc(w_n13421_0[2]),.din(n13421));
	jspl jspl_w_n13423_0(.douta(w_n13423_0[0]),.doutb(w_n13423_0[1]),.din(n13423));
	jspl jspl_w_n13428_0(.douta(w_n13428_0[0]),.doutb(w_n13428_0[1]),.din(n13428));
	jspl jspl_w_n13430_0(.douta(w_n13430_0[0]),.doutb(w_n13430_0[1]),.din(n13430));
	jspl jspl_w_n13431_0(.douta(w_n13431_0[0]),.doutb(w_n13431_0[1]),.din(n13431));
	jspl3 jspl3_w_n13432_0(.douta(w_n13432_0[0]),.doutb(w_n13432_0[1]),.doutc(w_n13432_0[2]),.din(n13432));
	jspl jspl_w_n13433_0(.douta(w_n13433_0[0]),.doutb(w_n13433_0[1]),.din(n13433));
	jspl jspl_w_n13437_0(.douta(w_n13437_0[0]),.doutb(w_n13437_0[1]),.din(n13437));
	jspl jspl_w_n13443_0(.douta(w_n13443_0[0]),.doutb(w_n13443_0[1]),.din(n13443));
	jspl jspl_w_n13444_0(.douta(w_n13444_0[0]),.doutb(w_n13444_0[1]),.din(n13444));
	jspl jspl_w_n13446_0(.douta(w_n13446_0[0]),.doutb(w_n13446_0[1]),.din(n13446));
	jspl jspl_w_n13448_0(.douta(w_n13448_0[0]),.doutb(w_n13448_0[1]),.din(n13448));
	jspl jspl_w_n13451_0(.douta(w_n13451_0[0]),.doutb(w_n13451_0[1]),.din(n13451));
	jspl jspl_w_n13457_0(.douta(w_n13457_0[0]),.doutb(w_n13457_0[1]),.din(n13457));
	jspl jspl_w_n13459_0(.douta(w_n13459_0[0]),.doutb(w_n13459_0[1]),.din(n13459));
	jspl3 jspl3_w_n13460_0(.douta(w_n13460_0[0]),.doutb(w_n13460_0[1]),.doutc(w_n13460_0[2]),.din(n13460));
	jspl jspl_w_n13464_0(.douta(w_n13464_0[0]),.doutb(w_n13464_0[1]),.din(n13464));
	jspl jspl_w_n13465_0(.douta(w_n13465_0[0]),.doutb(w_n13465_0[1]),.din(n13465));
	jspl3 jspl3_w_n13466_0(.douta(w_n13466_0[0]),.doutb(w_n13466_0[1]),.doutc(w_n13466_0[2]),.din(n13466));
	jspl jspl_w_n13468_0(.douta(w_n13468_0[0]),.doutb(w_n13468_0[1]),.din(n13468));
	jspl jspl_w_n13473_0(.douta(w_n13473_0[0]),.doutb(w_n13473_0[1]),.din(n13473));
	jspl jspl_w_n13475_0(.douta(w_n13475_0[0]),.doutb(w_n13475_0[1]),.din(n13475));
	jspl jspl_w_n13476_0(.douta(w_n13476_0[0]),.doutb(w_n13476_0[1]),.din(n13476));
	jspl3 jspl3_w_n13477_0(.douta(w_n13477_0[0]),.doutb(w_n13477_0[1]),.doutc(w_n13477_0[2]),.din(n13477));
	jspl jspl_w_n13478_0(.douta(w_n13478_0[0]),.doutb(w_n13478_0[1]),.din(n13478));
	jspl jspl_w_n13482_0(.douta(w_n13482_0[0]),.doutb(w_n13482_0[1]),.din(n13482));
	jspl jspl_w_n13488_0(.douta(w_n13488_0[0]),.doutb(w_n13488_0[1]),.din(n13488));
	jspl jspl_w_n13489_0(.douta(w_n13489_0[0]),.doutb(w_n13489_0[1]),.din(n13489));
	jspl jspl_w_n13491_0(.douta(w_n13491_0[0]),.doutb(w_n13491_0[1]),.din(n13491));
	jspl jspl_w_n13493_0(.douta(w_n13493_0[0]),.doutb(w_n13493_0[1]),.din(n13493));
	jspl jspl_w_n13496_0(.douta(w_n13496_0[0]),.doutb(w_n13496_0[1]),.din(n13496));
	jspl jspl_w_n13502_0(.douta(w_n13502_0[0]),.doutb(w_n13502_0[1]),.din(n13502));
	jspl jspl_w_n13504_0(.douta(w_n13504_0[0]),.doutb(w_n13504_0[1]),.din(n13504));
	jspl3 jspl3_w_n13505_0(.douta(w_n13505_0[0]),.doutb(w_n13505_0[1]),.doutc(w_n13505_0[2]),.din(n13505));
	jspl jspl_w_n13509_0(.douta(w_n13509_0[0]),.doutb(w_n13509_0[1]),.din(n13509));
	jspl jspl_w_n13510_0(.douta(w_n13510_0[0]),.doutb(w_n13510_0[1]),.din(n13510));
	jspl3 jspl3_w_n13511_0(.douta(w_n13511_0[0]),.doutb(w_n13511_0[1]),.doutc(w_n13511_0[2]),.din(n13511));
	jspl jspl_w_n13513_0(.douta(w_n13513_0[0]),.doutb(w_n13513_0[1]),.din(n13513));
	jspl jspl_w_n13518_0(.douta(w_n13518_0[0]),.doutb(w_n13518_0[1]),.din(n13518));
	jspl jspl_w_n13520_0(.douta(w_n13520_0[0]),.doutb(w_n13520_0[1]),.din(n13520));
	jspl jspl_w_n13521_0(.douta(w_n13521_0[0]),.doutb(w_n13521_0[1]),.din(n13521));
	jspl3 jspl3_w_n13522_0(.douta(w_n13522_0[0]),.doutb(w_n13522_0[1]),.doutc(w_n13522_0[2]),.din(n13522));
	jspl jspl_w_n13523_0(.douta(w_n13523_0[0]),.doutb(w_n13523_0[1]),.din(n13523));
	jspl jspl_w_n13527_0(.douta(w_n13527_0[0]),.doutb(w_n13527_0[1]),.din(n13527));
	jspl jspl_w_n13533_0(.douta(w_n13533_0[0]),.doutb(w_n13533_0[1]),.din(n13533));
	jspl jspl_w_n13534_0(.douta(w_n13534_0[0]),.doutb(w_n13534_0[1]),.din(n13534));
	jspl jspl_w_n13536_0(.douta(w_n13536_0[0]),.doutb(w_n13536_0[1]),.din(n13536));
	jspl jspl_w_n13541_0(.douta(w_n13541_0[0]),.doutb(w_n13541_0[1]),.din(n13541));
	jspl jspl_w_n13543_0(.douta(w_n13543_0[0]),.doutb(w_n13543_0[1]),.din(n13543));
	jspl jspl_w_n13544_0(.douta(w_n13544_0[0]),.doutb(w_n13544_0[1]),.din(n13544));
	jspl3 jspl3_w_n13545_0(.douta(w_n13545_0[0]),.doutb(w_n13545_0[1]),.doutc(w_n13545_0[2]),.din(n13545));
	jspl jspl_w_n13546_0(.douta(w_n13546_0[0]),.doutb(w_n13546_0[1]),.din(n13546));
	jspl jspl_w_n13548_0(.douta(w_n13548_0[0]),.doutb(w_n13548_0[1]),.din(n13548));
	jspl jspl_w_n13550_0(.douta(w_n13550_0[0]),.doutb(w_n13550_0[1]),.din(n13550));
	jspl jspl_w_n13552_0(.douta(w_n13552_0[0]),.doutb(w_n13552_0[1]),.din(n13552));
	jspl jspl_w_n13555_0(.douta(w_n13555_0[0]),.doutb(w_n13555_0[1]),.din(n13555));
	jspl jspl_w_n13561_0(.douta(w_n13561_0[0]),.doutb(w_n13561_0[1]),.din(n13561));
	jspl3 jspl3_w_n13563_0(.douta(w_n13563_0[0]),.doutb(w_n13563_0[1]),.doutc(w_n13563_0[2]),.din(n13563));
	jspl jspl_w_n13564_0(.douta(w_n13564_0[0]),.doutb(w_n13564_0[1]),.din(n13564));
	jspl jspl_w_n13568_0(.douta(w_n13568_0[0]),.doutb(w_n13568_0[1]),.din(n13568));
	jspl jspl_w_n13574_0(.douta(w_n13574_0[0]),.doutb(w_n13574_0[1]),.din(n13574));
	jspl jspl_w_n13575_0(.douta(w_n13575_0[0]),.doutb(w_n13575_0[1]),.din(n13575));
	jspl jspl_w_n13577_0(.douta(w_n13577_0[0]),.doutb(w_n13577_0[1]),.din(n13577));
	jspl jspl_w_n13579_0(.douta(w_n13579_0[0]),.doutb(w_n13579_0[1]),.din(n13579));
	jspl jspl_w_n13582_0(.douta(w_n13582_0[0]),.doutb(w_n13582_0[1]),.din(n13582));
	jspl jspl_w_n13588_0(.douta(w_n13588_0[0]),.doutb(w_n13588_0[1]),.din(n13588));
	jspl jspl_w_n13590_0(.douta(w_n13590_0[0]),.doutb(w_n13590_0[1]),.din(n13590));
	jspl3 jspl3_w_n13591_0(.douta(w_n13591_0[0]),.doutb(w_n13591_0[1]),.doutc(w_n13591_0[2]),.din(n13591));
	jspl jspl_w_n13595_0(.douta(w_n13595_0[0]),.doutb(w_n13595_0[1]),.din(n13595));
	jspl jspl_w_n13596_0(.douta(w_n13596_0[0]),.doutb(w_n13596_0[1]),.din(n13596));
	jspl3 jspl3_w_n13597_0(.douta(w_n13597_0[0]),.doutb(w_n13597_0[1]),.doutc(w_n13597_0[2]),.din(n13597));
	jspl jspl_w_n13599_0(.douta(w_n13599_0[0]),.doutb(w_n13599_0[1]),.din(n13599));
	jspl jspl_w_n13604_0(.douta(w_n13604_0[0]),.doutb(w_n13604_0[1]),.din(n13604));
	jspl jspl_w_n13606_0(.douta(w_n13606_0[0]),.doutb(w_n13606_0[1]),.din(n13606));
	jspl jspl_w_n13607_0(.douta(w_n13607_0[0]),.doutb(w_n13607_0[1]),.din(n13607));
	jspl3 jspl3_w_n13608_0(.douta(w_n13608_0[0]),.doutb(w_n13608_0[1]),.doutc(w_n13608_0[2]),.din(n13608));
	jspl jspl_w_n13609_0(.douta(w_n13609_0[0]),.doutb(w_n13609_0[1]),.din(n13609));
	jspl jspl_w_n13613_0(.douta(w_n13613_0[0]),.doutb(w_n13613_0[1]),.din(n13613));
	jspl jspl_w_n13619_0(.douta(w_n13619_0[0]),.doutb(w_n13619_0[1]),.din(n13619));
	jspl jspl_w_n13620_0(.douta(w_n13620_0[0]),.doutb(w_n13620_0[1]),.din(n13620));
	jspl jspl_w_n13622_0(.douta(w_n13622_0[0]),.doutb(w_n13622_0[1]),.din(n13622));
	jspl jspl_w_n13624_0(.douta(w_n13624_0[0]),.doutb(w_n13624_0[1]),.din(n13624));
	jspl jspl_w_n13627_0(.douta(w_n13627_0[0]),.doutb(w_n13627_0[1]),.din(n13627));
	jspl jspl_w_n13633_0(.douta(w_n13633_0[0]),.doutb(w_n13633_0[1]),.din(n13633));
	jspl jspl_w_n13635_0(.douta(w_n13635_0[0]),.doutb(w_n13635_0[1]),.din(n13635));
	jspl3 jspl3_w_n13636_0(.douta(w_n13636_0[0]),.doutb(w_n13636_0[1]),.doutc(w_n13636_0[2]),.din(n13636));
	jspl jspl_w_n13640_0(.douta(w_n13640_0[0]),.doutb(w_n13640_0[1]),.din(n13640));
	jspl jspl_w_n13641_0(.douta(w_n13641_0[0]),.doutb(w_n13641_0[1]),.din(n13641));
	jspl3 jspl3_w_n13642_0(.douta(w_n13642_0[0]),.doutb(w_n13642_0[1]),.doutc(w_n13642_0[2]),.din(n13642));
	jspl jspl_w_n13644_0(.douta(w_n13644_0[0]),.doutb(w_n13644_0[1]),.din(n13644));
	jspl jspl_w_n13649_0(.douta(w_n13649_0[0]),.doutb(w_n13649_0[1]),.din(n13649));
	jspl jspl_w_n13651_0(.douta(w_n13651_0[0]),.doutb(w_n13651_0[1]),.din(n13651));
	jspl jspl_w_n13652_0(.douta(w_n13652_0[0]),.doutb(w_n13652_0[1]),.din(n13652));
	jspl3 jspl3_w_n13653_0(.douta(w_n13653_0[0]),.doutb(w_n13653_0[1]),.doutc(w_n13653_0[2]),.din(n13653));
	jspl jspl_w_n13654_0(.douta(w_n13654_0[0]),.doutb(w_n13654_0[1]),.din(n13654));
	jspl jspl_w_n13658_0(.douta(w_n13658_0[0]),.doutb(w_n13658_0[1]),.din(n13658));
	jspl jspl_w_n13664_0(.douta(w_n13664_0[0]),.doutb(w_n13664_0[1]),.din(n13664));
	jspl jspl_w_n13665_0(.douta(w_n13665_0[0]),.doutb(w_n13665_0[1]),.din(n13665));
	jspl jspl_w_n13667_0(.douta(w_n13667_0[0]),.doutb(w_n13667_0[1]),.din(n13667));
	jspl jspl_w_n13669_0(.douta(w_n13669_0[0]),.doutb(w_n13669_0[1]),.din(n13669));
	jspl jspl_w_n13672_0(.douta(w_n13672_0[0]),.doutb(w_n13672_0[1]),.din(n13672));
	jspl jspl_w_n13678_0(.douta(w_n13678_0[0]),.doutb(w_n13678_0[1]),.din(n13678));
	jspl jspl_w_n13680_0(.douta(w_n13680_0[0]),.doutb(w_n13680_0[1]),.din(n13680));
	jspl3 jspl3_w_n13681_0(.douta(w_n13681_0[0]),.doutb(w_n13681_0[1]),.doutc(w_n13681_0[2]),.din(n13681));
	jspl jspl_w_n13685_0(.douta(w_n13685_0[0]),.doutb(w_n13685_0[1]),.din(n13685));
	jspl jspl_w_n13686_0(.douta(w_n13686_0[0]),.doutb(w_n13686_0[1]),.din(n13686));
	jspl3 jspl3_w_n13687_0(.douta(w_n13687_0[0]),.doutb(w_n13687_0[1]),.doutc(w_n13687_0[2]),.din(n13687));
	jspl jspl_w_n13689_0(.douta(w_n13689_0[0]),.doutb(w_n13689_0[1]),.din(n13689));
	jspl jspl_w_n13694_0(.douta(w_n13694_0[0]),.doutb(w_n13694_0[1]),.din(n13694));
	jspl jspl_w_n13696_0(.douta(w_n13696_0[0]),.doutb(w_n13696_0[1]),.din(n13696));
	jspl jspl_w_n13697_0(.douta(w_n13697_0[0]),.doutb(w_n13697_0[1]),.din(n13697));
	jspl3 jspl3_w_n13698_0(.douta(w_n13698_0[0]),.doutb(w_n13698_0[1]),.doutc(w_n13698_0[2]),.din(n13698));
	jspl3 jspl3_w_n13698_1(.douta(w_n13698_1[0]),.doutb(w_n13698_1[1]),.doutc(w_n13698_1[2]),.din(w_n13698_0[0]));
	jspl jspl_w_n13701_0(.douta(w_n13701_0[0]),.doutb(w_n13701_0[1]),.din(n13701));
	jspl3 jspl3_w_n13702_0(.douta(w_n13702_0[0]),.doutb(w_n13702_0[1]),.doutc(w_n13702_0[2]),.din(n13702));
	jspl jspl_w_n13703_0(.douta(w_n13703_0[0]),.doutb(w_n13703_0[1]),.din(n13703));
	jspl jspl_w_n13704_0(.douta(w_n13704_0[0]),.doutb(w_n13704_0[1]),.din(n13704));
	jspl jspl_w_n13710_0(.douta(w_n13710_0[0]),.doutb(w_n13710_0[1]),.din(n13710));
	jspl3 jspl3_w_n13711_0(.douta(w_n13711_0[0]),.doutb(w_n13711_0[1]),.doutc(w_n13711_0[2]),.din(n13711));
	jspl jspl_w_n13712_0(.douta(w_n13712_0[0]),.doutb(w_n13712_0[1]),.din(n13712));
	jspl jspl_w_n13717_0(.douta(w_n13717_0[0]),.doutb(w_n13717_0[1]),.din(n13717));
	jspl3 jspl3_w_n13718_0(.douta(w_n13718_0[0]),.doutb(w_n13718_0[1]),.doutc(w_n13718_0[2]),.din(n13718));
	jspl3 jspl3_w_n13718_1(.douta(w_n13718_1[0]),.doutb(w_n13718_1[1]),.doutc(w_n13718_1[2]),.din(w_n13718_0[0]));
	jspl3 jspl3_w_n13718_2(.douta(w_n13718_2[0]),.doutb(w_n13718_2[1]),.doutc(w_n13718_2[2]),.din(w_n13718_0[1]));
	jspl3 jspl3_w_n13718_3(.douta(w_n13718_3[0]),.doutb(w_n13718_3[1]),.doutc(w_n13718_3[2]),.din(w_n13718_0[2]));
	jspl3 jspl3_w_n13718_4(.douta(w_n13718_4[0]),.doutb(w_n13718_4[1]),.doutc(w_n13718_4[2]),.din(w_n13718_1[0]));
	jspl3 jspl3_w_n13718_5(.douta(w_n13718_5[0]),.doutb(w_n13718_5[1]),.doutc(w_n13718_5[2]),.din(w_n13718_1[1]));
	jspl3 jspl3_w_n13718_6(.douta(w_n13718_6[0]),.doutb(w_n13718_6[1]),.doutc(w_n13718_6[2]),.din(w_n13718_1[2]));
	jspl3 jspl3_w_n13718_7(.douta(w_n13718_7[0]),.doutb(w_n13718_7[1]),.doutc(w_n13718_7[2]),.din(w_n13718_2[0]));
	jspl3 jspl3_w_n13718_8(.douta(w_n13718_8[0]),.doutb(w_n13718_8[1]),.doutc(w_n13718_8[2]),.din(w_n13718_2[1]));
	jspl jspl_w_n13718_9(.douta(w_n13718_9[0]),.doutb(w_n13718_9[1]),.din(w_n13718_2[2]));
	jspl3 jspl3_w_n13723_0(.douta(w_n13723_0[0]),.doutb(w_n13723_0[1]),.doutc(w_n13723_0[2]),.din(n13723));
	jspl3 jspl3_w_n13723_1(.douta(w_n13723_1[0]),.doutb(w_n13723_1[1]),.doutc(w_n13723_1[2]),.din(w_n13723_0[0]));
	jspl3 jspl3_w_n13723_2(.douta(w_n13723_2[0]),.doutb(w_n13723_2[1]),.doutc(w_n13723_2[2]),.din(w_n13723_0[1]));
	jspl3 jspl3_w_n13723_3(.douta(w_n13723_3[0]),.doutb(w_n13723_3[1]),.doutc(w_n13723_3[2]),.din(w_n13723_0[2]));
	jspl3 jspl3_w_n13723_4(.douta(w_n13723_4[0]),.doutb(w_n13723_4[1]),.doutc(w_n13723_4[2]),.din(w_n13723_1[0]));
	jspl3 jspl3_w_n13723_5(.douta(w_n13723_5[0]),.doutb(w_n13723_5[1]),.doutc(w_n13723_5[2]),.din(w_n13723_1[1]));
	jspl3 jspl3_w_n13723_6(.douta(w_n13723_6[0]),.doutb(w_n13723_6[1]),.doutc(w_n13723_6[2]),.din(w_n13723_1[2]));
	jspl3 jspl3_w_n13723_7(.douta(w_n13723_7[0]),.doutb(w_n13723_7[1]),.doutc(w_n13723_7[2]),.din(w_n13723_2[0]));
	jspl3 jspl3_w_n13723_8(.douta(w_n13723_8[0]),.doutb(w_n13723_8[1]),.doutc(w_n13723_8[2]),.din(w_n13723_2[1]));
	jspl3 jspl3_w_n13723_9(.douta(w_n13723_9[0]),.doutb(w_n13723_9[1]),.doutc(w_n13723_9[2]),.din(w_n13723_2[2]));
	jspl3 jspl3_w_n13723_10(.douta(w_n13723_10[0]),.doutb(w_n13723_10[1]),.doutc(w_n13723_10[2]),.din(w_n13723_3[0]));
	jspl3 jspl3_w_n13723_11(.douta(w_n13723_11[0]),.doutb(w_n13723_11[1]),.doutc(w_n13723_11[2]),.din(w_n13723_3[1]));
	jspl3 jspl3_w_n13723_12(.douta(w_n13723_12[0]),.doutb(w_n13723_12[1]),.doutc(w_n13723_12[2]),.din(w_n13723_3[2]));
	jspl3 jspl3_w_n13723_13(.douta(w_n13723_13[0]),.doutb(w_n13723_13[1]),.doutc(w_n13723_13[2]),.din(w_n13723_4[0]));
	jspl3 jspl3_w_n13723_14(.douta(w_n13723_14[0]),.doutb(w_n13723_14[1]),.doutc(w_n13723_14[2]),.din(w_n13723_4[1]));
	jspl3 jspl3_w_n13723_15(.douta(w_n13723_15[0]),.doutb(w_n13723_15[1]),.doutc(w_n13723_15[2]),.din(w_n13723_4[2]));
	jspl3 jspl3_w_n13723_16(.douta(w_n13723_16[0]),.doutb(w_n13723_16[1]),.doutc(w_n13723_16[2]),.din(w_n13723_5[0]));
	jspl3 jspl3_w_n13723_17(.douta(w_n13723_17[0]),.doutb(w_n13723_17[1]),.doutc(w_n13723_17[2]),.din(w_n13723_5[1]));
	jspl3 jspl3_w_n13723_18(.douta(w_n13723_18[0]),.doutb(w_n13723_18[1]),.doutc(w_n13723_18[2]),.din(w_n13723_5[2]));
	jspl3 jspl3_w_n13723_19(.douta(w_n13723_19[0]),.doutb(w_n13723_19[1]),.doutc(w_n13723_19[2]),.din(w_n13723_6[0]));
	jspl3 jspl3_w_n13723_20(.douta(w_n13723_20[0]),.doutb(w_n13723_20[1]),.doutc(w_n13723_20[2]),.din(w_n13723_6[1]));
	jspl3 jspl3_w_n13723_21(.douta(w_n13723_21[0]),.doutb(w_n13723_21[1]),.doutc(w_n13723_21[2]),.din(w_n13723_6[2]));
	jspl3 jspl3_w_n13723_22(.douta(w_n13723_22[0]),.doutb(w_n13723_22[1]),.doutc(w_n13723_22[2]),.din(w_n13723_7[0]));
	jspl jspl_w_n13726_0(.douta(w_n13726_0[0]),.doutb(w_n13726_0[1]),.din(n13726));
	jspl3 jspl3_w_n13728_0(.douta(w_n13728_0[0]),.doutb(w_n13728_0[1]),.doutc(w_n13728_0[2]),.din(n13728));
	jspl jspl_w_n13728_1(.douta(w_n13728_1[0]),.doutb(w_n13728_1[1]),.din(w_n13728_0[0]));
	jspl3 jspl3_w_n13729_0(.douta(w_n13729_0[0]),.doutb(w_n13729_0[1]),.doutc(w_n13729_0[2]),.din(n13729));
	jspl3 jspl3_w_n13733_0(.douta(w_n13733_0[0]),.doutb(w_n13733_0[1]),.doutc(w_n13733_0[2]),.din(n13733));
	jspl jspl_w_n13734_0(.douta(w_n13734_0[0]),.doutb(w_n13734_0[1]),.din(n13734));
	jspl jspl_w_n13735_0(.douta(w_n13735_0[0]),.doutb(w_n13735_0[1]),.din(n13735));
	jspl jspl_w_n13736_0(.douta(w_n13736_0[0]),.doutb(w_n13736_0[1]),.din(n13736));
	jspl jspl_w_n13738_0(.douta(w_n13738_0[0]),.doutb(w_n13738_0[1]),.din(n13738));
	jspl jspl_w_n13740_0(.douta(w_n13740_0[0]),.doutb(w_n13740_0[1]),.din(n13740));
	jspl jspl_w_n13742_0(.douta(w_n13742_0[0]),.doutb(w_n13742_0[1]),.din(n13742));
	jspl jspl_w_n13745_0(.douta(w_n13745_0[0]),.doutb(w_n13745_0[1]),.din(n13745));
	jspl jspl_w_n13750_0(.douta(w_n13750_0[0]),.doutb(w_n13750_0[1]),.din(n13750));
	jspl3 jspl3_w_n13752_0(.douta(w_n13752_0[0]),.doutb(w_n13752_0[1]),.doutc(w_n13752_0[2]),.din(n13752));
	jspl jspl_w_n13753_0(.douta(w_n13753_0[0]),.doutb(w_n13753_0[1]),.din(n13753));
	jspl jspl_w_n13757_0(.douta(w_n13757_0[0]),.doutb(w_n13757_0[1]),.din(n13757));
	jspl jspl_w_n13758_0(.douta(w_n13758_0[0]),.doutb(w_n13758_0[1]),.din(n13758));
	jspl jspl_w_n13760_0(.douta(w_n13760_0[0]),.doutb(w_n13760_0[1]),.din(n13760));
	jspl jspl_w_n13764_0(.douta(w_n13764_0[0]),.doutb(w_n13764_0[1]),.din(n13764));
	jspl jspl_w_n13766_0(.douta(w_n13766_0[0]),.doutb(w_n13766_0[1]),.din(n13766));
	jspl jspl_w_n13767_0(.douta(w_n13767_0[0]),.doutb(w_n13767_0[1]),.din(n13767));
	jspl3 jspl3_w_n13768_0(.douta(w_n13768_0[0]),.doutb(w_n13768_0[1]),.doutc(w_n13768_0[2]),.din(n13768));
	jspl jspl_w_n13769_0(.douta(w_n13769_0[0]),.doutb(w_n13769_0[1]),.din(n13769));
	jspl jspl_w_n13773_0(.douta(w_n13773_0[0]),.doutb(w_n13773_0[1]),.din(n13773));
	jspl jspl_w_n13775_0(.douta(w_n13775_0[0]),.doutb(w_n13775_0[1]),.din(n13775));
	jspl jspl_w_n13777_0(.douta(w_n13777_0[0]),.doutb(w_n13777_0[1]),.din(n13777));
	jspl jspl_w_n13779_0(.douta(w_n13779_0[0]),.doutb(w_n13779_0[1]),.din(n13779));
	jspl jspl_w_n13782_0(.douta(w_n13782_0[0]),.doutb(w_n13782_0[1]),.din(n13782));
	jspl jspl_w_n13788_0(.douta(w_n13788_0[0]),.doutb(w_n13788_0[1]),.din(n13788));
	jspl3 jspl3_w_n13790_0(.douta(w_n13790_0[0]),.doutb(w_n13790_0[1]),.doutc(w_n13790_0[2]),.din(n13790));
	jspl jspl_w_n13791_0(.douta(w_n13791_0[0]),.doutb(w_n13791_0[1]),.din(n13791));
	jspl jspl_w_n13796_0(.douta(w_n13796_0[0]),.doutb(w_n13796_0[1]),.din(n13796));
	jspl jspl_w_n13798_0(.douta(w_n13798_0[0]),.doutb(w_n13798_0[1]),.din(n13798));
	jspl jspl_w_n13800_0(.douta(w_n13800_0[0]),.doutb(w_n13800_0[1]),.din(n13800));
	jspl jspl_w_n13804_0(.douta(w_n13804_0[0]),.doutb(w_n13804_0[1]),.din(n13804));
	jspl jspl_w_n13806_0(.douta(w_n13806_0[0]),.doutb(w_n13806_0[1]),.din(n13806));
	jspl jspl_w_n13807_0(.douta(w_n13807_0[0]),.doutb(w_n13807_0[1]),.din(n13807));
	jspl3 jspl3_w_n13808_0(.douta(w_n13808_0[0]),.doutb(w_n13808_0[1]),.doutc(w_n13808_0[2]),.din(n13808));
	jspl jspl_w_n13809_0(.douta(w_n13809_0[0]),.doutb(w_n13809_0[1]),.din(n13809));
	jspl jspl_w_n13815_0(.douta(w_n13815_0[0]),.doutb(w_n13815_0[1]),.din(n13815));
	jspl jspl_w_n13816_0(.douta(w_n13816_0[0]),.doutb(w_n13816_0[1]),.din(n13816));
	jspl jspl_w_n13818_0(.douta(w_n13818_0[0]),.doutb(w_n13818_0[1]),.din(n13818));
	jspl jspl_w_n13820_0(.douta(w_n13820_0[0]),.doutb(w_n13820_0[1]),.din(n13820));
	jspl jspl_w_n13822_0(.douta(w_n13822_0[0]),.doutb(w_n13822_0[1]),.din(n13822));
	jspl jspl_w_n13828_0(.douta(w_n13828_0[0]),.doutb(w_n13828_0[1]),.din(n13828));
	jspl jspl_w_n13830_0(.douta(w_n13830_0[0]),.doutb(w_n13830_0[1]),.din(n13830));
	jspl3 jspl3_w_n13831_0(.douta(w_n13831_0[0]),.doutb(w_n13831_0[1]),.doutc(w_n13831_0[2]),.din(n13831));
	jspl jspl_w_n13834_0(.douta(w_n13834_0[0]),.doutb(w_n13834_0[1]),.din(n13834));
	jspl jspl_w_n13835_0(.douta(w_n13835_0[0]),.doutb(w_n13835_0[1]),.din(n13835));
	jspl3 jspl3_w_n13836_0(.douta(w_n13836_0[0]),.doutb(w_n13836_0[1]),.doutc(w_n13836_0[2]),.din(n13836));
	jspl jspl_w_n13838_0(.douta(w_n13838_0[0]),.doutb(w_n13838_0[1]),.din(n13838));
	jspl jspl_w_n13842_0(.douta(w_n13842_0[0]),.doutb(w_n13842_0[1]),.din(n13842));
	jspl jspl_w_n13844_0(.douta(w_n13844_0[0]),.doutb(w_n13844_0[1]),.din(n13844));
	jspl jspl_w_n13845_0(.douta(w_n13845_0[0]),.doutb(w_n13845_0[1]),.din(n13845));
	jspl3 jspl3_w_n13846_0(.douta(w_n13846_0[0]),.doutb(w_n13846_0[1]),.doutc(w_n13846_0[2]),.din(n13846));
	jspl jspl_w_n13847_0(.douta(w_n13847_0[0]),.doutb(w_n13847_0[1]),.din(n13847));
	jspl jspl_w_n13850_0(.douta(w_n13850_0[0]),.doutb(w_n13850_0[1]),.din(n13850));
	jspl jspl_w_n13856_0(.douta(w_n13856_0[0]),.doutb(w_n13856_0[1]),.din(n13856));
	jspl jspl_w_n13857_0(.douta(w_n13857_0[0]),.doutb(w_n13857_0[1]),.din(n13857));
	jspl jspl_w_n13859_0(.douta(w_n13859_0[0]),.doutb(w_n13859_0[1]),.din(n13859));
	jspl jspl_w_n13861_0(.douta(w_n13861_0[0]),.doutb(w_n13861_0[1]),.din(n13861));
	jspl jspl_w_n13863_0(.douta(w_n13863_0[0]),.doutb(w_n13863_0[1]),.din(n13863));
	jspl jspl_w_n13869_0(.douta(w_n13869_0[0]),.doutb(w_n13869_0[1]),.din(n13869));
	jspl jspl_w_n13871_0(.douta(w_n13871_0[0]),.doutb(w_n13871_0[1]),.din(n13871));
	jspl3 jspl3_w_n13872_0(.douta(w_n13872_0[0]),.doutb(w_n13872_0[1]),.doutc(w_n13872_0[2]),.din(n13872));
	jspl jspl_w_n13875_0(.douta(w_n13875_0[0]),.doutb(w_n13875_0[1]),.din(n13875));
	jspl jspl_w_n13876_0(.douta(w_n13876_0[0]),.doutb(w_n13876_0[1]),.din(n13876));
	jspl3 jspl3_w_n13877_0(.douta(w_n13877_0[0]),.doutb(w_n13877_0[1]),.doutc(w_n13877_0[2]),.din(n13877));
	jspl jspl_w_n13879_0(.douta(w_n13879_0[0]),.doutb(w_n13879_0[1]),.din(n13879));
	jspl jspl_w_n13883_0(.douta(w_n13883_0[0]),.doutb(w_n13883_0[1]),.din(n13883));
	jspl jspl_w_n13885_0(.douta(w_n13885_0[0]),.doutb(w_n13885_0[1]),.din(n13885));
	jspl jspl_w_n13886_0(.douta(w_n13886_0[0]),.doutb(w_n13886_0[1]),.din(n13886));
	jspl3 jspl3_w_n13887_0(.douta(w_n13887_0[0]),.doutb(w_n13887_0[1]),.doutc(w_n13887_0[2]),.din(n13887));
	jspl jspl_w_n13888_0(.douta(w_n13888_0[0]),.doutb(w_n13888_0[1]),.din(n13888));
	jspl jspl_w_n13891_0(.douta(w_n13891_0[0]),.doutb(w_n13891_0[1]),.din(n13891));
	jspl jspl_w_n13897_0(.douta(w_n13897_0[0]),.doutb(w_n13897_0[1]),.din(n13897));
	jspl jspl_w_n13898_0(.douta(w_n13898_0[0]),.doutb(w_n13898_0[1]),.din(n13898));
	jspl jspl_w_n13900_0(.douta(w_n13900_0[0]),.doutb(w_n13900_0[1]),.din(n13900));
	jspl jspl_w_n13902_0(.douta(w_n13902_0[0]),.doutb(w_n13902_0[1]),.din(n13902));
	jspl jspl_w_n13904_0(.douta(w_n13904_0[0]),.doutb(w_n13904_0[1]),.din(n13904));
	jspl jspl_w_n13910_0(.douta(w_n13910_0[0]),.doutb(w_n13910_0[1]),.din(n13910));
	jspl jspl_w_n13912_0(.douta(w_n13912_0[0]),.doutb(w_n13912_0[1]),.din(n13912));
	jspl3 jspl3_w_n13913_0(.douta(w_n13913_0[0]),.doutb(w_n13913_0[1]),.doutc(w_n13913_0[2]),.din(n13913));
	jspl jspl_w_n13916_0(.douta(w_n13916_0[0]),.doutb(w_n13916_0[1]),.din(n13916));
	jspl jspl_w_n13917_0(.douta(w_n13917_0[0]),.doutb(w_n13917_0[1]),.din(n13917));
	jspl3 jspl3_w_n13918_0(.douta(w_n13918_0[0]),.doutb(w_n13918_0[1]),.doutc(w_n13918_0[2]),.din(n13918));
	jspl jspl_w_n13920_0(.douta(w_n13920_0[0]),.doutb(w_n13920_0[1]),.din(n13920));
	jspl jspl_w_n13924_0(.douta(w_n13924_0[0]),.doutb(w_n13924_0[1]),.din(n13924));
	jspl jspl_w_n13926_0(.douta(w_n13926_0[0]),.doutb(w_n13926_0[1]),.din(n13926));
	jspl jspl_w_n13927_0(.douta(w_n13927_0[0]),.doutb(w_n13927_0[1]),.din(n13927));
	jspl3 jspl3_w_n13928_0(.douta(w_n13928_0[0]),.doutb(w_n13928_0[1]),.doutc(w_n13928_0[2]),.din(n13928));
	jspl jspl_w_n13929_0(.douta(w_n13929_0[0]),.doutb(w_n13929_0[1]),.din(n13929));
	jspl jspl_w_n13932_0(.douta(w_n13932_0[0]),.doutb(w_n13932_0[1]),.din(n13932));
	jspl jspl_w_n13938_0(.douta(w_n13938_0[0]),.doutb(w_n13938_0[1]),.din(n13938));
	jspl jspl_w_n13939_0(.douta(w_n13939_0[0]),.doutb(w_n13939_0[1]),.din(n13939));
	jspl jspl_w_n13941_0(.douta(w_n13941_0[0]),.doutb(w_n13941_0[1]),.din(n13941));
	jspl jspl_w_n13943_0(.douta(w_n13943_0[0]),.doutb(w_n13943_0[1]),.din(n13943));
	jspl jspl_w_n13945_0(.douta(w_n13945_0[0]),.doutb(w_n13945_0[1]),.din(n13945));
	jspl jspl_w_n13951_0(.douta(w_n13951_0[0]),.doutb(w_n13951_0[1]),.din(n13951));
	jspl jspl_w_n13953_0(.douta(w_n13953_0[0]),.doutb(w_n13953_0[1]),.din(n13953));
	jspl3 jspl3_w_n13954_0(.douta(w_n13954_0[0]),.doutb(w_n13954_0[1]),.doutc(w_n13954_0[2]),.din(n13954));
	jspl jspl_w_n13957_0(.douta(w_n13957_0[0]),.doutb(w_n13957_0[1]),.din(n13957));
	jspl jspl_w_n13958_0(.douta(w_n13958_0[0]),.doutb(w_n13958_0[1]),.din(n13958));
	jspl3 jspl3_w_n13959_0(.douta(w_n13959_0[0]),.doutb(w_n13959_0[1]),.doutc(w_n13959_0[2]),.din(n13959));
	jspl jspl_w_n13961_0(.douta(w_n13961_0[0]),.doutb(w_n13961_0[1]),.din(n13961));
	jspl jspl_w_n13965_0(.douta(w_n13965_0[0]),.doutb(w_n13965_0[1]),.din(n13965));
	jspl jspl_w_n13967_0(.douta(w_n13967_0[0]),.doutb(w_n13967_0[1]),.din(n13967));
	jspl jspl_w_n13968_0(.douta(w_n13968_0[0]),.doutb(w_n13968_0[1]),.din(n13968));
	jspl3 jspl3_w_n13969_0(.douta(w_n13969_0[0]),.doutb(w_n13969_0[1]),.doutc(w_n13969_0[2]),.din(n13969));
	jspl jspl_w_n13970_0(.douta(w_n13970_0[0]),.doutb(w_n13970_0[1]),.din(n13970));
	jspl jspl_w_n13973_0(.douta(w_n13973_0[0]),.doutb(w_n13973_0[1]),.din(n13973));
	jspl jspl_w_n13979_0(.douta(w_n13979_0[0]),.doutb(w_n13979_0[1]),.din(n13979));
	jspl jspl_w_n13980_0(.douta(w_n13980_0[0]),.doutb(w_n13980_0[1]),.din(n13980));
	jspl jspl_w_n13982_0(.douta(w_n13982_0[0]),.doutb(w_n13982_0[1]),.din(n13982));
	jspl jspl_w_n13984_0(.douta(w_n13984_0[0]),.doutb(w_n13984_0[1]),.din(n13984));
	jspl jspl_w_n13986_0(.douta(w_n13986_0[0]),.doutb(w_n13986_0[1]),.din(n13986));
	jspl jspl_w_n13992_0(.douta(w_n13992_0[0]),.doutb(w_n13992_0[1]),.din(n13992));
	jspl jspl_w_n13994_0(.douta(w_n13994_0[0]),.doutb(w_n13994_0[1]),.din(n13994));
	jspl3 jspl3_w_n13995_0(.douta(w_n13995_0[0]),.doutb(w_n13995_0[1]),.doutc(w_n13995_0[2]),.din(n13995));
	jspl jspl_w_n13998_0(.douta(w_n13998_0[0]),.doutb(w_n13998_0[1]),.din(n13998));
	jspl jspl_w_n13999_0(.douta(w_n13999_0[0]),.doutb(w_n13999_0[1]),.din(n13999));
	jspl3 jspl3_w_n14000_0(.douta(w_n14000_0[0]),.doutb(w_n14000_0[1]),.doutc(w_n14000_0[2]),.din(n14000));
	jspl jspl_w_n14002_0(.douta(w_n14002_0[0]),.doutb(w_n14002_0[1]),.din(n14002));
	jspl jspl_w_n14006_0(.douta(w_n14006_0[0]),.doutb(w_n14006_0[1]),.din(n14006));
	jspl jspl_w_n14008_0(.douta(w_n14008_0[0]),.doutb(w_n14008_0[1]),.din(n14008));
	jspl jspl_w_n14009_0(.douta(w_n14009_0[0]),.doutb(w_n14009_0[1]),.din(n14009));
	jspl3 jspl3_w_n14010_0(.douta(w_n14010_0[0]),.doutb(w_n14010_0[1]),.doutc(w_n14010_0[2]),.din(n14010));
	jspl jspl_w_n14011_0(.douta(w_n14011_0[0]),.doutb(w_n14011_0[1]),.din(n14011));
	jspl jspl_w_n14014_0(.douta(w_n14014_0[0]),.doutb(w_n14014_0[1]),.din(n14014));
	jspl jspl_w_n14020_0(.douta(w_n14020_0[0]),.doutb(w_n14020_0[1]),.din(n14020));
	jspl jspl_w_n14021_0(.douta(w_n14021_0[0]),.doutb(w_n14021_0[1]),.din(n14021));
	jspl jspl_w_n14023_0(.douta(w_n14023_0[0]),.doutb(w_n14023_0[1]),.din(n14023));
	jspl jspl_w_n14025_0(.douta(w_n14025_0[0]),.doutb(w_n14025_0[1]),.din(n14025));
	jspl jspl_w_n14027_0(.douta(w_n14027_0[0]),.doutb(w_n14027_0[1]),.din(n14027));
	jspl jspl_w_n14033_0(.douta(w_n14033_0[0]),.doutb(w_n14033_0[1]),.din(n14033));
	jspl jspl_w_n14035_0(.douta(w_n14035_0[0]),.doutb(w_n14035_0[1]),.din(n14035));
	jspl3 jspl3_w_n14036_0(.douta(w_n14036_0[0]),.doutb(w_n14036_0[1]),.doutc(w_n14036_0[2]),.din(n14036));
	jspl jspl_w_n14039_0(.douta(w_n14039_0[0]),.doutb(w_n14039_0[1]),.din(n14039));
	jspl jspl_w_n14040_0(.douta(w_n14040_0[0]),.doutb(w_n14040_0[1]),.din(n14040));
	jspl3 jspl3_w_n14041_0(.douta(w_n14041_0[0]),.doutb(w_n14041_0[1]),.doutc(w_n14041_0[2]),.din(n14041));
	jspl jspl_w_n14043_0(.douta(w_n14043_0[0]),.doutb(w_n14043_0[1]),.din(n14043));
	jspl jspl_w_n14047_0(.douta(w_n14047_0[0]),.doutb(w_n14047_0[1]),.din(n14047));
	jspl jspl_w_n14049_0(.douta(w_n14049_0[0]),.doutb(w_n14049_0[1]),.din(n14049));
	jspl jspl_w_n14050_0(.douta(w_n14050_0[0]),.doutb(w_n14050_0[1]),.din(n14050));
	jspl3 jspl3_w_n14051_0(.douta(w_n14051_0[0]),.doutb(w_n14051_0[1]),.doutc(w_n14051_0[2]),.din(n14051));
	jspl jspl_w_n14052_0(.douta(w_n14052_0[0]),.doutb(w_n14052_0[1]),.din(n14052));
	jspl jspl_w_n14055_0(.douta(w_n14055_0[0]),.doutb(w_n14055_0[1]),.din(n14055));
	jspl jspl_w_n14061_0(.douta(w_n14061_0[0]),.doutb(w_n14061_0[1]),.din(n14061));
	jspl jspl_w_n14062_0(.douta(w_n14062_0[0]),.doutb(w_n14062_0[1]),.din(n14062));
	jspl jspl_w_n14064_0(.douta(w_n14064_0[0]),.doutb(w_n14064_0[1]),.din(n14064));
	jspl jspl_w_n14066_0(.douta(w_n14066_0[0]),.doutb(w_n14066_0[1]),.din(n14066));
	jspl jspl_w_n14068_0(.douta(w_n14068_0[0]),.doutb(w_n14068_0[1]),.din(n14068));
	jspl jspl_w_n14074_0(.douta(w_n14074_0[0]),.doutb(w_n14074_0[1]),.din(n14074));
	jspl jspl_w_n14076_0(.douta(w_n14076_0[0]),.doutb(w_n14076_0[1]),.din(n14076));
	jspl3 jspl3_w_n14077_0(.douta(w_n14077_0[0]),.doutb(w_n14077_0[1]),.doutc(w_n14077_0[2]),.din(n14077));
	jspl jspl_w_n14080_0(.douta(w_n14080_0[0]),.doutb(w_n14080_0[1]),.din(n14080));
	jspl jspl_w_n14081_0(.douta(w_n14081_0[0]),.doutb(w_n14081_0[1]),.din(n14081));
	jspl3 jspl3_w_n14082_0(.douta(w_n14082_0[0]),.doutb(w_n14082_0[1]),.doutc(w_n14082_0[2]),.din(n14082));
	jspl jspl_w_n14084_0(.douta(w_n14084_0[0]),.doutb(w_n14084_0[1]),.din(n14084));
	jspl jspl_w_n14086_0(.douta(w_n14086_0[0]),.doutb(w_n14086_0[1]),.din(n14086));
	jspl jspl_w_n14088_0(.douta(w_n14088_0[0]),.doutb(w_n14088_0[1]),.din(n14088));
	jspl jspl_w_n14094_0(.douta(w_n14094_0[0]),.doutb(w_n14094_0[1]),.din(n14094));
	jspl3 jspl3_w_n14096_0(.douta(w_n14096_0[0]),.doutb(w_n14096_0[1]),.doutc(w_n14096_0[2]),.din(n14096));
	jspl jspl_w_n14097_0(.douta(w_n14097_0[0]),.doutb(w_n14097_0[1]),.din(n14097));
	jspl jspl_w_n14099_0(.douta(w_n14099_0[0]),.doutb(w_n14099_0[1]),.din(n14099));
	jspl jspl_w_n14101_0(.douta(w_n14101_0[0]),.doutb(w_n14101_0[1]),.din(n14101));
	jspl jspl_w_n14105_0(.douta(w_n14105_0[0]),.doutb(w_n14105_0[1]),.din(n14105));
	jspl jspl_w_n14107_0(.douta(w_n14107_0[0]),.doutb(w_n14107_0[1]),.din(n14107));
	jspl jspl_w_n14108_0(.douta(w_n14108_0[0]),.doutb(w_n14108_0[1]),.din(n14108));
	jspl jspl_w_n14109_0(.douta(w_n14109_0[0]),.doutb(w_n14109_0[1]),.din(n14109));
	jspl3 jspl3_w_n14110_0(.douta(w_n14110_0[0]),.doutb(w_n14110_0[1]),.doutc(w_n14110_0[2]),.din(n14110));
	jspl jspl_w_n14113_0(.douta(w_n14113_0[0]),.doutb(w_n14113_0[1]),.din(n14113));
	jspl jspl_w_n14114_0(.douta(w_n14114_0[0]),.doutb(w_n14114_0[1]),.din(n14114));
	jspl3 jspl3_w_n14115_0(.douta(w_n14115_0[0]),.doutb(w_n14115_0[1]),.doutc(w_n14115_0[2]),.din(n14115));
	jspl jspl_w_n14117_0(.douta(w_n14117_0[0]),.doutb(w_n14117_0[1]),.din(n14117));
	jspl jspl_w_n14121_0(.douta(w_n14121_0[0]),.doutb(w_n14121_0[1]),.din(n14121));
	jspl jspl_w_n14123_0(.douta(w_n14123_0[0]),.doutb(w_n14123_0[1]),.din(n14123));
	jspl jspl_w_n14124_0(.douta(w_n14124_0[0]),.doutb(w_n14124_0[1]),.din(n14124));
	jspl3 jspl3_w_n14125_0(.douta(w_n14125_0[0]),.doutb(w_n14125_0[1]),.doutc(w_n14125_0[2]),.din(n14125));
	jspl jspl_w_n14126_0(.douta(w_n14126_0[0]),.doutb(w_n14126_0[1]),.din(n14126));
	jspl jspl_w_n14129_0(.douta(w_n14129_0[0]),.doutb(w_n14129_0[1]),.din(n14129));
	jspl jspl_w_n14135_0(.douta(w_n14135_0[0]),.doutb(w_n14135_0[1]),.din(n14135));
	jspl jspl_w_n14136_0(.douta(w_n14136_0[0]),.doutb(w_n14136_0[1]),.din(n14136));
	jspl jspl_w_n14138_0(.douta(w_n14138_0[0]),.doutb(w_n14138_0[1]),.din(n14138));
	jspl jspl_w_n14140_0(.douta(w_n14140_0[0]),.doutb(w_n14140_0[1]),.din(n14140));
	jspl jspl_w_n14142_0(.douta(w_n14142_0[0]),.doutb(w_n14142_0[1]),.din(n14142));
	jspl jspl_w_n14148_0(.douta(w_n14148_0[0]),.doutb(w_n14148_0[1]),.din(n14148));
	jspl jspl_w_n14150_0(.douta(w_n14150_0[0]),.doutb(w_n14150_0[1]),.din(n14150));
	jspl3 jspl3_w_n14151_0(.douta(w_n14151_0[0]),.doutb(w_n14151_0[1]),.doutc(w_n14151_0[2]),.din(n14151));
	jspl jspl_w_n14154_0(.douta(w_n14154_0[0]),.doutb(w_n14154_0[1]),.din(n14154));
	jspl jspl_w_n14155_0(.douta(w_n14155_0[0]),.doutb(w_n14155_0[1]),.din(n14155));
	jspl3 jspl3_w_n14156_0(.douta(w_n14156_0[0]),.doutb(w_n14156_0[1]),.doutc(w_n14156_0[2]),.din(n14156));
	jspl jspl_w_n14158_0(.douta(w_n14158_0[0]),.doutb(w_n14158_0[1]),.din(n14158));
	jspl jspl_w_n14162_0(.douta(w_n14162_0[0]),.doutb(w_n14162_0[1]),.din(n14162));
	jspl jspl_w_n14164_0(.douta(w_n14164_0[0]),.doutb(w_n14164_0[1]),.din(n14164));
	jspl jspl_w_n14165_0(.douta(w_n14165_0[0]),.doutb(w_n14165_0[1]),.din(n14165));
	jspl3 jspl3_w_n14166_0(.douta(w_n14166_0[0]),.doutb(w_n14166_0[1]),.doutc(w_n14166_0[2]),.din(n14166));
	jspl jspl_w_n14167_0(.douta(w_n14167_0[0]),.doutb(w_n14167_0[1]),.din(n14167));
	jspl jspl_w_n14170_0(.douta(w_n14170_0[0]),.doutb(w_n14170_0[1]),.din(n14170));
	jspl jspl_w_n14176_0(.douta(w_n14176_0[0]),.doutb(w_n14176_0[1]),.din(n14176));
	jspl jspl_w_n14177_0(.douta(w_n14177_0[0]),.doutb(w_n14177_0[1]),.din(n14177));
	jspl jspl_w_n14179_0(.douta(w_n14179_0[0]),.doutb(w_n14179_0[1]),.din(n14179));
	jspl jspl_w_n14181_0(.douta(w_n14181_0[0]),.doutb(w_n14181_0[1]),.din(n14181));
	jspl jspl_w_n14183_0(.douta(w_n14183_0[0]),.doutb(w_n14183_0[1]),.din(n14183));
	jspl jspl_w_n14189_0(.douta(w_n14189_0[0]),.doutb(w_n14189_0[1]),.din(n14189));
	jspl jspl_w_n14191_0(.douta(w_n14191_0[0]),.doutb(w_n14191_0[1]),.din(n14191));
	jspl3 jspl3_w_n14192_0(.douta(w_n14192_0[0]),.doutb(w_n14192_0[1]),.doutc(w_n14192_0[2]),.din(n14192));
	jspl jspl_w_n14195_0(.douta(w_n14195_0[0]),.doutb(w_n14195_0[1]),.din(n14195));
	jspl jspl_w_n14196_0(.douta(w_n14196_0[0]),.doutb(w_n14196_0[1]),.din(n14196));
	jspl3 jspl3_w_n14197_0(.douta(w_n14197_0[0]),.doutb(w_n14197_0[1]),.doutc(w_n14197_0[2]),.din(n14197));
	jspl jspl_w_n14199_0(.douta(w_n14199_0[0]),.doutb(w_n14199_0[1]),.din(n14199));
	jspl jspl_w_n14203_0(.douta(w_n14203_0[0]),.doutb(w_n14203_0[1]),.din(n14203));
	jspl jspl_w_n14205_0(.douta(w_n14205_0[0]),.doutb(w_n14205_0[1]),.din(n14205));
	jspl jspl_w_n14206_0(.douta(w_n14206_0[0]),.doutb(w_n14206_0[1]),.din(n14206));
	jspl3 jspl3_w_n14207_0(.douta(w_n14207_0[0]),.doutb(w_n14207_0[1]),.doutc(w_n14207_0[2]),.din(n14207));
	jspl jspl_w_n14211_0(.douta(w_n14211_0[0]),.doutb(w_n14211_0[1]),.din(n14211));
	jspl jspl_w_n14217_0(.douta(w_n14217_0[0]),.doutb(w_n14217_0[1]),.din(n14217));
	jspl3 jspl3_w_n14219_0(.douta(w_n14219_0[0]),.doutb(w_n14219_0[1]),.doutc(w_n14219_0[2]),.din(n14219));
	jspl jspl_w_n14221_0(.douta(w_n14221_0[0]),.doutb(w_n14221_0[1]),.din(n14221));
	jspl3 jspl3_w_n14226_0(.douta(w_n14226_0[0]),.doutb(w_n14226_0[1]),.doutc(w_n14226_0[2]),.din(n14226));
	jspl jspl_w_n14227_0(.douta(w_n14227_0[0]),.doutb(w_n14227_0[1]),.din(n14227));
	jspl jspl_w_n14228_0(.douta(w_n14228_0[0]),.doutb(w_n14228_0[1]),.din(n14228));
	jspl jspl_w_n14233_0(.douta(w_n14233_0[0]),.doutb(w_n14233_0[1]),.din(n14233));
	jspl3 jspl3_w_n14234_0(.douta(w_n14234_0[0]),.doutb(w_n14234_0[1]),.doutc(w_n14234_0[2]),.din(n14234));
	jspl jspl_w_n14239_0(.douta(w_n14239_0[0]),.doutb(w_n14239_0[1]),.din(n14239));
	jspl jspl_w_n14246_0(.douta(w_n14246_0[0]),.doutb(w_n14246_0[1]),.din(n14246));
	jspl3 jspl3_w_n14248_0(.douta(w_n14248_0[0]),.doutb(w_n14248_0[1]),.doutc(w_n14248_0[2]),.din(n14248));
	jspl jspl_w_n14248_1(.douta(w_n14248_1[0]),.doutb(w_n14248_1[1]),.din(w_n14248_0[0]));
	jspl jspl_w_n14249_0(.douta(w_n14249_0[0]),.doutb(w_n14249_0[1]),.din(n14249));
	jspl3 jspl3_w_n14252_0(.douta(w_n14252_0[0]),.doutb(w_n14252_0[1]),.doutc(w_n14252_0[2]),.din(n14252));
	jspl jspl_w_n14253_0(.douta(w_n14253_0[0]),.doutb(w_n14253_0[1]),.din(n14253));
	jspl jspl_w_n14254_0(.douta(w_n14254_0[0]),.doutb(w_n14254_0[1]),.din(n14254));
	jspl jspl_w_n14255_0(.douta(w_n14255_0[0]),.doutb(w_n14255_0[1]),.din(n14255));
	jspl jspl_w_n14257_0(.douta(w_n14257_0[0]),.doutb(w_n14257_0[1]),.din(n14257));
	jspl jspl_w_n14259_0(.douta(w_n14259_0[0]),.doutb(w_n14259_0[1]),.din(n14259));
	jspl jspl_w_n14261_0(.douta(w_n14261_0[0]),.doutb(w_n14261_0[1]),.din(n14261));
	jspl jspl_w_n14270_0(.douta(w_n14270_0[0]),.doutb(w_n14270_0[1]),.din(n14270));
	jspl3 jspl3_w_n14272_0(.douta(w_n14272_0[0]),.doutb(w_n14272_0[1]),.doutc(w_n14272_0[2]),.din(n14272));
	jspl jspl_w_n14273_0(.douta(w_n14273_0[0]),.doutb(w_n14273_0[1]),.din(n14273));
	jspl jspl_w_n14277_0(.douta(w_n14277_0[0]),.doutb(w_n14277_0[1]),.din(n14277));
	jspl jspl_w_n14279_0(.douta(w_n14279_0[0]),.doutb(w_n14279_0[1]),.din(n14279));
	jspl jspl_w_n14281_0(.douta(w_n14281_0[0]),.doutb(w_n14281_0[1]),.din(n14281));
	jspl jspl_w_n14286_0(.douta(w_n14286_0[0]),.doutb(w_n14286_0[1]),.din(n14286));
	jspl jspl_w_n14288_0(.douta(w_n14288_0[0]),.doutb(w_n14288_0[1]),.din(n14288));
	jspl jspl_w_n14289_0(.douta(w_n14289_0[0]),.doutb(w_n14289_0[1]),.din(n14289));
	jspl3 jspl3_w_n14290_0(.douta(w_n14290_0[0]),.doutb(w_n14290_0[1]),.doutc(w_n14290_0[2]),.din(n14290));
	jspl jspl_w_n14291_0(.douta(w_n14291_0[0]),.doutb(w_n14291_0[1]),.din(n14291));
	jspl jspl_w_n14296_0(.douta(w_n14296_0[0]),.doutb(w_n14296_0[1]),.din(n14296));
	jspl jspl_w_n14297_0(.douta(w_n14297_0[0]),.doutb(w_n14297_0[1]),.din(n14297));
	jspl jspl_w_n14299_0(.douta(w_n14299_0[0]),.doutb(w_n14299_0[1]),.din(n14299));
	jspl jspl_w_n14301_0(.douta(w_n14301_0[0]),.doutb(w_n14301_0[1]),.din(n14301));
	jspl jspl_w_n14304_0(.douta(w_n14304_0[0]),.doutb(w_n14304_0[1]),.din(n14304));
	jspl jspl_w_n14310_0(.douta(w_n14310_0[0]),.doutb(w_n14310_0[1]),.din(n14310));
	jspl3 jspl3_w_n14312_0(.douta(w_n14312_0[0]),.doutb(w_n14312_0[1]),.doutc(w_n14312_0[2]),.din(n14312));
	jspl jspl_w_n14313_0(.douta(w_n14313_0[0]),.doutb(w_n14313_0[1]),.din(n14313));
	jspl jspl_w_n14317_0(.douta(w_n14317_0[0]),.doutb(w_n14317_0[1]),.din(n14317));
	jspl jspl_w_n14318_0(.douta(w_n14318_0[0]),.doutb(w_n14318_0[1]),.din(n14318));
	jspl jspl_w_n14320_0(.douta(w_n14320_0[0]),.doutb(w_n14320_0[1]),.din(n14320));
	jspl jspl_w_n14325_0(.douta(w_n14325_0[0]),.doutb(w_n14325_0[1]),.din(n14325));
	jspl jspl_w_n14327_0(.douta(w_n14327_0[0]),.doutb(w_n14327_0[1]),.din(n14327));
	jspl jspl_w_n14328_0(.douta(w_n14328_0[0]),.doutb(w_n14328_0[1]),.din(n14328));
	jspl3 jspl3_w_n14329_0(.douta(w_n14329_0[0]),.doutb(w_n14329_0[1]),.doutc(w_n14329_0[2]),.din(n14329));
	jspl jspl_w_n14330_0(.douta(w_n14330_0[0]),.doutb(w_n14330_0[1]),.din(n14330));
	jspl jspl_w_n14334_0(.douta(w_n14334_0[0]),.doutb(w_n14334_0[1]),.din(n14334));
	jspl jspl_w_n14335_0(.douta(w_n14335_0[0]),.doutb(w_n14335_0[1]),.din(n14335));
	jspl jspl_w_n14337_0(.douta(w_n14337_0[0]),.doutb(w_n14337_0[1]),.din(n14337));
	jspl jspl_w_n14339_0(.douta(w_n14339_0[0]),.doutb(w_n14339_0[1]),.din(n14339));
	jspl jspl_w_n14342_0(.douta(w_n14342_0[0]),.doutb(w_n14342_0[1]),.din(n14342));
	jspl jspl_w_n14348_0(.douta(w_n14348_0[0]),.doutb(w_n14348_0[1]),.din(n14348));
	jspl jspl_w_n14350_0(.douta(w_n14350_0[0]),.doutb(w_n14350_0[1]),.din(n14350));
	jspl3 jspl3_w_n14351_0(.douta(w_n14351_0[0]),.doutb(w_n14351_0[1]),.doutc(w_n14351_0[2]),.din(n14351));
	jspl jspl_w_n14355_0(.douta(w_n14355_0[0]),.doutb(w_n14355_0[1]),.din(n14355));
	jspl jspl_w_n14356_0(.douta(w_n14356_0[0]),.doutb(w_n14356_0[1]),.din(n14356));
	jspl3 jspl3_w_n14357_0(.douta(w_n14357_0[0]),.doutb(w_n14357_0[1]),.doutc(w_n14357_0[2]),.din(n14357));
	jspl jspl_w_n14359_0(.douta(w_n14359_0[0]),.doutb(w_n14359_0[1]),.din(n14359));
	jspl jspl_w_n14364_0(.douta(w_n14364_0[0]),.doutb(w_n14364_0[1]),.din(n14364));
	jspl jspl_w_n14366_0(.douta(w_n14366_0[0]),.doutb(w_n14366_0[1]),.din(n14366));
	jspl jspl_w_n14367_0(.douta(w_n14367_0[0]),.doutb(w_n14367_0[1]),.din(n14367));
	jspl3 jspl3_w_n14368_0(.douta(w_n14368_0[0]),.doutb(w_n14368_0[1]),.doutc(w_n14368_0[2]),.din(n14368));
	jspl jspl_w_n14369_0(.douta(w_n14369_0[0]),.doutb(w_n14369_0[1]),.din(n14369));
	jspl jspl_w_n14373_0(.douta(w_n14373_0[0]),.doutb(w_n14373_0[1]),.din(n14373));
	jspl jspl_w_n14379_0(.douta(w_n14379_0[0]),.doutb(w_n14379_0[1]),.din(n14379));
	jspl jspl_w_n14380_0(.douta(w_n14380_0[0]),.doutb(w_n14380_0[1]),.din(n14380));
	jspl jspl_w_n14382_0(.douta(w_n14382_0[0]),.doutb(w_n14382_0[1]),.din(n14382));
	jspl jspl_w_n14384_0(.douta(w_n14384_0[0]),.doutb(w_n14384_0[1]),.din(n14384));
	jspl jspl_w_n14387_0(.douta(w_n14387_0[0]),.doutb(w_n14387_0[1]),.din(n14387));
	jspl jspl_w_n14393_0(.douta(w_n14393_0[0]),.doutb(w_n14393_0[1]),.din(n14393));
	jspl jspl_w_n14395_0(.douta(w_n14395_0[0]),.doutb(w_n14395_0[1]),.din(n14395));
	jspl3 jspl3_w_n14396_0(.douta(w_n14396_0[0]),.doutb(w_n14396_0[1]),.doutc(w_n14396_0[2]),.din(n14396));
	jspl jspl_w_n14400_0(.douta(w_n14400_0[0]),.doutb(w_n14400_0[1]),.din(n14400));
	jspl jspl_w_n14401_0(.douta(w_n14401_0[0]),.doutb(w_n14401_0[1]),.din(n14401));
	jspl3 jspl3_w_n14402_0(.douta(w_n14402_0[0]),.doutb(w_n14402_0[1]),.doutc(w_n14402_0[2]),.din(n14402));
	jspl jspl_w_n14404_0(.douta(w_n14404_0[0]),.doutb(w_n14404_0[1]),.din(n14404));
	jspl jspl_w_n14409_0(.douta(w_n14409_0[0]),.doutb(w_n14409_0[1]),.din(n14409));
	jspl jspl_w_n14411_0(.douta(w_n14411_0[0]),.doutb(w_n14411_0[1]),.din(n14411));
	jspl jspl_w_n14412_0(.douta(w_n14412_0[0]),.doutb(w_n14412_0[1]),.din(n14412));
	jspl3 jspl3_w_n14413_0(.douta(w_n14413_0[0]),.doutb(w_n14413_0[1]),.doutc(w_n14413_0[2]),.din(n14413));
	jspl jspl_w_n14414_0(.douta(w_n14414_0[0]),.doutb(w_n14414_0[1]),.din(n14414));
	jspl jspl_w_n14418_0(.douta(w_n14418_0[0]),.doutb(w_n14418_0[1]),.din(n14418));
	jspl jspl_w_n14424_0(.douta(w_n14424_0[0]),.doutb(w_n14424_0[1]),.din(n14424));
	jspl jspl_w_n14425_0(.douta(w_n14425_0[0]),.doutb(w_n14425_0[1]),.din(n14425));
	jspl jspl_w_n14427_0(.douta(w_n14427_0[0]),.doutb(w_n14427_0[1]),.din(n14427));
	jspl jspl_w_n14429_0(.douta(w_n14429_0[0]),.doutb(w_n14429_0[1]),.din(n14429));
	jspl jspl_w_n14432_0(.douta(w_n14432_0[0]),.doutb(w_n14432_0[1]),.din(n14432));
	jspl jspl_w_n14438_0(.douta(w_n14438_0[0]),.doutb(w_n14438_0[1]),.din(n14438));
	jspl jspl_w_n14440_0(.douta(w_n14440_0[0]),.doutb(w_n14440_0[1]),.din(n14440));
	jspl3 jspl3_w_n14441_0(.douta(w_n14441_0[0]),.doutb(w_n14441_0[1]),.doutc(w_n14441_0[2]),.din(n14441));
	jspl jspl_w_n14445_0(.douta(w_n14445_0[0]),.doutb(w_n14445_0[1]),.din(n14445));
	jspl jspl_w_n14446_0(.douta(w_n14446_0[0]),.doutb(w_n14446_0[1]),.din(n14446));
	jspl3 jspl3_w_n14447_0(.douta(w_n14447_0[0]),.doutb(w_n14447_0[1]),.doutc(w_n14447_0[2]),.din(n14447));
	jspl jspl_w_n14449_0(.douta(w_n14449_0[0]),.doutb(w_n14449_0[1]),.din(n14449));
	jspl jspl_w_n14454_0(.douta(w_n14454_0[0]),.doutb(w_n14454_0[1]),.din(n14454));
	jspl jspl_w_n14456_0(.douta(w_n14456_0[0]),.doutb(w_n14456_0[1]),.din(n14456));
	jspl jspl_w_n14457_0(.douta(w_n14457_0[0]),.doutb(w_n14457_0[1]),.din(n14457));
	jspl3 jspl3_w_n14458_0(.douta(w_n14458_0[0]),.doutb(w_n14458_0[1]),.doutc(w_n14458_0[2]),.din(n14458));
	jspl jspl_w_n14459_0(.douta(w_n14459_0[0]),.doutb(w_n14459_0[1]),.din(n14459));
	jspl jspl_w_n14463_0(.douta(w_n14463_0[0]),.doutb(w_n14463_0[1]),.din(n14463));
	jspl jspl_w_n14469_0(.douta(w_n14469_0[0]),.doutb(w_n14469_0[1]),.din(n14469));
	jspl jspl_w_n14470_0(.douta(w_n14470_0[0]),.doutb(w_n14470_0[1]),.din(n14470));
	jspl jspl_w_n14472_0(.douta(w_n14472_0[0]),.doutb(w_n14472_0[1]),.din(n14472));
	jspl jspl_w_n14474_0(.douta(w_n14474_0[0]),.doutb(w_n14474_0[1]),.din(n14474));
	jspl jspl_w_n14477_0(.douta(w_n14477_0[0]),.doutb(w_n14477_0[1]),.din(n14477));
	jspl jspl_w_n14483_0(.douta(w_n14483_0[0]),.doutb(w_n14483_0[1]),.din(n14483));
	jspl jspl_w_n14485_0(.douta(w_n14485_0[0]),.doutb(w_n14485_0[1]),.din(n14485));
	jspl3 jspl3_w_n14486_0(.douta(w_n14486_0[0]),.doutb(w_n14486_0[1]),.doutc(w_n14486_0[2]),.din(n14486));
	jspl jspl_w_n14490_0(.douta(w_n14490_0[0]),.doutb(w_n14490_0[1]),.din(n14490));
	jspl jspl_w_n14491_0(.douta(w_n14491_0[0]),.doutb(w_n14491_0[1]),.din(n14491));
	jspl3 jspl3_w_n14492_0(.douta(w_n14492_0[0]),.doutb(w_n14492_0[1]),.doutc(w_n14492_0[2]),.din(n14492));
	jspl jspl_w_n14494_0(.douta(w_n14494_0[0]),.doutb(w_n14494_0[1]),.din(n14494));
	jspl jspl_w_n14499_0(.douta(w_n14499_0[0]),.doutb(w_n14499_0[1]),.din(n14499));
	jspl jspl_w_n14501_0(.douta(w_n14501_0[0]),.doutb(w_n14501_0[1]),.din(n14501));
	jspl jspl_w_n14502_0(.douta(w_n14502_0[0]),.doutb(w_n14502_0[1]),.din(n14502));
	jspl3 jspl3_w_n14503_0(.douta(w_n14503_0[0]),.doutb(w_n14503_0[1]),.doutc(w_n14503_0[2]),.din(n14503));
	jspl jspl_w_n14504_0(.douta(w_n14504_0[0]),.doutb(w_n14504_0[1]),.din(n14504));
	jspl jspl_w_n14508_0(.douta(w_n14508_0[0]),.doutb(w_n14508_0[1]),.din(n14508));
	jspl jspl_w_n14514_0(.douta(w_n14514_0[0]),.doutb(w_n14514_0[1]),.din(n14514));
	jspl jspl_w_n14515_0(.douta(w_n14515_0[0]),.doutb(w_n14515_0[1]),.din(n14515));
	jspl jspl_w_n14517_0(.douta(w_n14517_0[0]),.doutb(w_n14517_0[1]),.din(n14517));
	jspl jspl_w_n14519_0(.douta(w_n14519_0[0]),.doutb(w_n14519_0[1]),.din(n14519));
	jspl jspl_w_n14522_0(.douta(w_n14522_0[0]),.doutb(w_n14522_0[1]),.din(n14522));
	jspl jspl_w_n14528_0(.douta(w_n14528_0[0]),.doutb(w_n14528_0[1]),.din(n14528));
	jspl jspl_w_n14530_0(.douta(w_n14530_0[0]),.doutb(w_n14530_0[1]),.din(n14530));
	jspl3 jspl3_w_n14531_0(.douta(w_n14531_0[0]),.doutb(w_n14531_0[1]),.doutc(w_n14531_0[2]),.din(n14531));
	jspl jspl_w_n14535_0(.douta(w_n14535_0[0]),.doutb(w_n14535_0[1]),.din(n14535));
	jspl jspl_w_n14536_0(.douta(w_n14536_0[0]),.doutb(w_n14536_0[1]),.din(n14536));
	jspl3 jspl3_w_n14537_0(.douta(w_n14537_0[0]),.doutb(w_n14537_0[1]),.doutc(w_n14537_0[2]),.din(n14537));
	jspl jspl_w_n14539_0(.douta(w_n14539_0[0]),.doutb(w_n14539_0[1]),.din(n14539));
	jspl jspl_w_n14544_0(.douta(w_n14544_0[0]),.doutb(w_n14544_0[1]),.din(n14544));
	jspl jspl_w_n14546_0(.douta(w_n14546_0[0]),.doutb(w_n14546_0[1]),.din(n14546));
	jspl jspl_w_n14547_0(.douta(w_n14547_0[0]),.doutb(w_n14547_0[1]),.din(n14547));
	jspl3 jspl3_w_n14548_0(.douta(w_n14548_0[0]),.doutb(w_n14548_0[1]),.doutc(w_n14548_0[2]),.din(n14548));
	jspl jspl_w_n14549_0(.douta(w_n14549_0[0]),.doutb(w_n14549_0[1]),.din(n14549));
	jspl jspl_w_n14553_0(.douta(w_n14553_0[0]),.doutb(w_n14553_0[1]),.din(n14553));
	jspl jspl_w_n14559_0(.douta(w_n14559_0[0]),.doutb(w_n14559_0[1]),.din(n14559));
	jspl jspl_w_n14560_0(.douta(w_n14560_0[0]),.doutb(w_n14560_0[1]),.din(n14560));
	jspl jspl_w_n14562_0(.douta(w_n14562_0[0]),.doutb(w_n14562_0[1]),.din(n14562));
	jspl jspl_w_n14564_0(.douta(w_n14564_0[0]),.doutb(w_n14564_0[1]),.din(n14564));
	jspl jspl_w_n14567_0(.douta(w_n14567_0[0]),.doutb(w_n14567_0[1]),.din(n14567));
	jspl jspl_w_n14573_0(.douta(w_n14573_0[0]),.doutb(w_n14573_0[1]),.din(n14573));
	jspl jspl_w_n14575_0(.douta(w_n14575_0[0]),.doutb(w_n14575_0[1]),.din(n14575));
	jspl3 jspl3_w_n14576_0(.douta(w_n14576_0[0]),.doutb(w_n14576_0[1]),.doutc(w_n14576_0[2]),.din(n14576));
	jspl jspl_w_n14580_0(.douta(w_n14580_0[0]),.doutb(w_n14580_0[1]),.din(n14580));
	jspl jspl_w_n14581_0(.douta(w_n14581_0[0]),.doutb(w_n14581_0[1]),.din(n14581));
	jspl3 jspl3_w_n14582_0(.douta(w_n14582_0[0]),.doutb(w_n14582_0[1]),.doutc(w_n14582_0[2]),.din(n14582));
	jspl jspl_w_n14584_0(.douta(w_n14584_0[0]),.doutb(w_n14584_0[1]),.din(n14584));
	jspl jspl_w_n14589_0(.douta(w_n14589_0[0]),.doutb(w_n14589_0[1]),.din(n14589));
	jspl jspl_w_n14591_0(.douta(w_n14591_0[0]),.doutb(w_n14591_0[1]),.din(n14591));
	jspl jspl_w_n14592_0(.douta(w_n14592_0[0]),.doutb(w_n14592_0[1]),.din(n14592));
	jspl3 jspl3_w_n14593_0(.douta(w_n14593_0[0]),.doutb(w_n14593_0[1]),.doutc(w_n14593_0[2]),.din(n14593));
	jspl jspl_w_n14594_0(.douta(w_n14594_0[0]),.doutb(w_n14594_0[1]),.din(n14594));
	jspl jspl_w_n14598_0(.douta(w_n14598_0[0]),.doutb(w_n14598_0[1]),.din(n14598));
	jspl jspl_w_n14604_0(.douta(w_n14604_0[0]),.doutb(w_n14604_0[1]),.din(n14604));
	jspl jspl_w_n14605_0(.douta(w_n14605_0[0]),.doutb(w_n14605_0[1]),.din(n14605));
	jspl jspl_w_n14607_0(.douta(w_n14607_0[0]),.doutb(w_n14607_0[1]),.din(n14607));
	jspl jspl_w_n14609_0(.douta(w_n14609_0[0]),.doutb(w_n14609_0[1]),.din(n14609));
	jspl jspl_w_n14612_0(.douta(w_n14612_0[0]),.doutb(w_n14612_0[1]),.din(n14612));
	jspl jspl_w_n14618_0(.douta(w_n14618_0[0]),.doutb(w_n14618_0[1]),.din(n14618));
	jspl jspl_w_n14620_0(.douta(w_n14620_0[0]),.doutb(w_n14620_0[1]),.din(n14620));
	jspl3 jspl3_w_n14621_0(.douta(w_n14621_0[0]),.doutb(w_n14621_0[1]),.doutc(w_n14621_0[2]),.din(n14621));
	jspl jspl_w_n14625_0(.douta(w_n14625_0[0]),.doutb(w_n14625_0[1]),.din(n14625));
	jspl jspl_w_n14626_0(.douta(w_n14626_0[0]),.doutb(w_n14626_0[1]),.din(n14626));
	jspl3 jspl3_w_n14627_0(.douta(w_n14627_0[0]),.doutb(w_n14627_0[1]),.doutc(w_n14627_0[2]),.din(n14627));
	jspl jspl_w_n14629_0(.douta(w_n14629_0[0]),.doutb(w_n14629_0[1]),.din(n14629));
	jspl jspl_w_n14634_0(.douta(w_n14634_0[0]),.doutb(w_n14634_0[1]),.din(n14634));
	jspl jspl_w_n14636_0(.douta(w_n14636_0[0]),.doutb(w_n14636_0[1]),.din(n14636));
	jspl jspl_w_n14637_0(.douta(w_n14637_0[0]),.doutb(w_n14637_0[1]),.din(n14637));
	jspl3 jspl3_w_n14638_0(.douta(w_n14638_0[0]),.doutb(w_n14638_0[1]),.doutc(w_n14638_0[2]),.din(n14638));
	jspl jspl_w_n14639_0(.douta(w_n14639_0[0]),.doutb(w_n14639_0[1]),.din(n14639));
	jspl jspl_w_n14643_0(.douta(w_n14643_0[0]),.doutb(w_n14643_0[1]),.din(n14643));
	jspl jspl_w_n14649_0(.douta(w_n14649_0[0]),.doutb(w_n14649_0[1]),.din(n14649));
	jspl jspl_w_n14650_0(.douta(w_n14650_0[0]),.doutb(w_n14650_0[1]),.din(n14650));
	jspl jspl_w_n14652_0(.douta(w_n14652_0[0]),.doutb(w_n14652_0[1]),.din(n14652));
	jspl jspl_w_n14657_0(.douta(w_n14657_0[0]),.doutb(w_n14657_0[1]),.din(n14657));
	jspl jspl_w_n14659_0(.douta(w_n14659_0[0]),.doutb(w_n14659_0[1]),.din(n14659));
	jspl jspl_w_n14660_0(.douta(w_n14660_0[0]),.doutb(w_n14660_0[1]),.din(n14660));
	jspl3 jspl3_w_n14661_0(.douta(w_n14661_0[0]),.doutb(w_n14661_0[1]),.doutc(w_n14661_0[2]),.din(n14661));
	jspl jspl_w_n14662_0(.douta(w_n14662_0[0]),.doutb(w_n14662_0[1]),.din(n14662));
	jspl jspl_w_n14665_0(.douta(w_n14665_0[0]),.doutb(w_n14665_0[1]),.din(n14665));
	jspl jspl_w_n14667_0(.douta(w_n14667_0[0]),.doutb(w_n14667_0[1]),.din(n14667));
	jspl jspl_w_n14669_0(.douta(w_n14669_0[0]),.doutb(w_n14669_0[1]),.din(n14669));
	jspl jspl_w_n14672_0(.douta(w_n14672_0[0]),.doutb(w_n14672_0[1]),.din(n14672));
	jspl jspl_w_n14678_0(.douta(w_n14678_0[0]),.doutb(w_n14678_0[1]),.din(n14678));
	jspl3 jspl3_w_n14680_0(.douta(w_n14680_0[0]),.doutb(w_n14680_0[1]),.doutc(w_n14680_0[2]),.din(n14680));
	jspl jspl_w_n14681_0(.douta(w_n14681_0[0]),.doutb(w_n14681_0[1]),.din(n14681));
	jspl jspl_w_n14685_0(.douta(w_n14685_0[0]),.doutb(w_n14685_0[1]),.din(n14685));
	jspl jspl_w_n14691_0(.douta(w_n14691_0[0]),.doutb(w_n14691_0[1]),.din(n14691));
	jspl jspl_w_n14692_0(.douta(w_n14692_0[0]),.doutb(w_n14692_0[1]),.din(n14692));
	jspl jspl_w_n14694_0(.douta(w_n14694_0[0]),.doutb(w_n14694_0[1]),.din(n14694));
	jspl jspl_w_n14696_0(.douta(w_n14696_0[0]),.doutb(w_n14696_0[1]),.din(n14696));
	jspl jspl_w_n14699_0(.douta(w_n14699_0[0]),.doutb(w_n14699_0[1]),.din(n14699));
	jspl jspl_w_n14705_0(.douta(w_n14705_0[0]),.doutb(w_n14705_0[1]),.din(n14705));
	jspl jspl_w_n14707_0(.douta(w_n14707_0[0]),.doutb(w_n14707_0[1]),.din(n14707));
	jspl3 jspl3_w_n14708_0(.douta(w_n14708_0[0]),.doutb(w_n14708_0[1]),.doutc(w_n14708_0[2]),.din(n14708));
	jspl jspl_w_n14712_0(.douta(w_n14712_0[0]),.doutb(w_n14712_0[1]),.din(n14712));
	jspl jspl_w_n14713_0(.douta(w_n14713_0[0]),.doutb(w_n14713_0[1]),.din(n14713));
	jspl3 jspl3_w_n14714_0(.douta(w_n14714_0[0]),.doutb(w_n14714_0[1]),.doutc(w_n14714_0[2]),.din(n14714));
	jspl jspl_w_n14716_0(.douta(w_n14716_0[0]),.doutb(w_n14716_0[1]),.din(n14716));
	jspl jspl_w_n14721_0(.douta(w_n14721_0[0]),.doutb(w_n14721_0[1]),.din(n14721));
	jspl jspl_w_n14723_0(.douta(w_n14723_0[0]),.doutb(w_n14723_0[1]),.din(n14723));
	jspl jspl_w_n14724_0(.douta(w_n14724_0[0]),.doutb(w_n14724_0[1]),.din(n14724));
	jspl3 jspl3_w_n14725_0(.douta(w_n14725_0[0]),.doutb(w_n14725_0[1]),.doutc(w_n14725_0[2]),.din(n14725));
	jspl jspl_w_n14726_0(.douta(w_n14726_0[0]),.doutb(w_n14726_0[1]),.din(n14726));
	jspl jspl_w_n14730_0(.douta(w_n14730_0[0]),.doutb(w_n14730_0[1]),.din(n14730));
	jspl jspl_w_n14736_0(.douta(w_n14736_0[0]),.doutb(w_n14736_0[1]),.din(n14736));
	jspl jspl_w_n14737_0(.douta(w_n14737_0[0]),.doutb(w_n14737_0[1]),.din(n14737));
	jspl jspl_w_n14739_0(.douta(w_n14739_0[0]),.doutb(w_n14739_0[1]),.din(n14739));
	jspl jspl_w_n14741_0(.douta(w_n14741_0[0]),.doutb(w_n14741_0[1]),.din(n14741));
	jspl jspl_w_n14744_0(.douta(w_n14744_0[0]),.doutb(w_n14744_0[1]),.din(n14744));
	jspl jspl_w_n14750_0(.douta(w_n14750_0[0]),.doutb(w_n14750_0[1]),.din(n14750));
	jspl jspl_w_n14752_0(.douta(w_n14752_0[0]),.doutb(w_n14752_0[1]),.din(n14752));
	jspl3 jspl3_w_n14753_0(.douta(w_n14753_0[0]),.doutb(w_n14753_0[1]),.doutc(w_n14753_0[2]),.din(n14753));
	jspl jspl_w_n14757_0(.douta(w_n14757_0[0]),.doutb(w_n14757_0[1]),.din(n14757));
	jspl jspl_w_n14758_0(.douta(w_n14758_0[0]),.doutb(w_n14758_0[1]),.din(n14758));
	jspl3 jspl3_w_n14759_0(.douta(w_n14759_0[0]),.doutb(w_n14759_0[1]),.doutc(w_n14759_0[2]),.din(n14759));
	jspl jspl_w_n14761_0(.douta(w_n14761_0[0]),.doutb(w_n14761_0[1]),.din(n14761));
	jspl jspl_w_n14766_0(.douta(w_n14766_0[0]),.doutb(w_n14766_0[1]),.din(n14766));
	jspl jspl_w_n14768_0(.douta(w_n14768_0[0]),.doutb(w_n14768_0[1]),.din(n14768));
	jspl jspl_w_n14769_0(.douta(w_n14769_0[0]),.doutb(w_n14769_0[1]),.din(n14769));
	jspl3 jspl3_w_n14770_0(.douta(w_n14770_0[0]),.doutb(w_n14770_0[1]),.doutc(w_n14770_0[2]),.din(n14770));
	jspl jspl_w_n14771_0(.douta(w_n14771_0[0]),.doutb(w_n14771_0[1]),.din(n14771));
	jspl jspl_w_n14775_0(.douta(w_n14775_0[0]),.doutb(w_n14775_0[1]),.din(n14775));
	jspl jspl_w_n14781_0(.douta(w_n14781_0[0]),.doutb(w_n14781_0[1]),.din(n14781));
	jspl jspl_w_n14782_0(.douta(w_n14782_0[0]),.doutb(w_n14782_0[1]),.din(n14782));
	jspl jspl_w_n14784_0(.douta(w_n14784_0[0]),.doutb(w_n14784_0[1]),.din(n14784));
	jspl jspl_w_n14786_0(.douta(w_n14786_0[0]),.doutb(w_n14786_0[1]),.din(n14786));
	jspl jspl_w_n14789_0(.douta(w_n14789_0[0]),.doutb(w_n14789_0[1]),.din(n14789));
	jspl jspl_w_n14795_0(.douta(w_n14795_0[0]),.doutb(w_n14795_0[1]),.din(n14795));
	jspl3 jspl3_w_n14797_0(.douta(w_n14797_0[0]),.doutb(w_n14797_0[1]),.doutc(w_n14797_0[2]),.din(n14797));
	jspl3 jspl3_w_n14797_1(.douta(w_n14797_1[0]),.doutb(w_n14797_1[1]),.doutc(w_n14797_1[2]),.din(w_n14797_0[0]));
	jspl jspl_w_n14800_0(.douta(w_n14800_0[0]),.doutb(w_n14800_0[1]),.din(n14800));
	jspl3 jspl3_w_n14801_0(.douta(w_n14801_0[0]),.doutb(w_n14801_0[1]),.doutc(w_n14801_0[2]),.din(n14801));
	jspl jspl_w_n14802_0(.douta(w_n14802_0[0]),.doutb(w_n14802_0[1]),.din(n14802));
	jspl jspl_w_n14808_0(.douta(w_n14808_0[0]),.doutb(w_n14808_0[1]),.din(n14808));
	jspl3 jspl3_w_n14809_0(.douta(w_n14809_0[0]),.doutb(w_n14809_0[1]),.doutc(w_n14809_0[2]),.din(n14809));
	jspl jspl_w_n14810_0(.douta(w_n14810_0[0]),.doutb(w_n14810_0[1]),.din(n14810));
	jspl jspl_w_n14815_0(.douta(w_n14815_0[0]),.doutb(w_n14815_0[1]),.din(n14815));
	jspl3 jspl3_w_n14816_0(.douta(w_n14816_0[0]),.doutb(w_n14816_0[1]),.doutc(w_n14816_0[2]),.din(n14816));
	jspl3 jspl3_w_n14816_1(.douta(w_n14816_1[0]),.doutb(w_n14816_1[1]),.doutc(w_n14816_1[2]),.din(w_n14816_0[0]));
	jspl3 jspl3_w_n14816_2(.douta(w_n14816_2[0]),.doutb(w_n14816_2[1]),.doutc(w_n14816_2[2]),.din(w_n14816_0[1]));
	jspl3 jspl3_w_n14816_3(.douta(w_n14816_3[0]),.doutb(w_n14816_3[1]),.doutc(w_n14816_3[2]),.din(w_n14816_0[2]));
	jspl3 jspl3_w_n14816_4(.douta(w_n14816_4[0]),.doutb(w_n14816_4[1]),.doutc(w_n14816_4[2]),.din(w_n14816_1[0]));
	jspl3 jspl3_w_n14816_5(.douta(w_n14816_5[0]),.doutb(w_n14816_5[1]),.doutc(w_n14816_5[2]),.din(w_n14816_1[1]));
	jspl3 jspl3_w_n14816_6(.douta(w_n14816_6[0]),.doutb(w_n14816_6[1]),.doutc(w_n14816_6[2]),.din(w_n14816_1[2]));
	jspl3 jspl3_w_n14816_7(.douta(w_n14816_7[0]),.doutb(w_n14816_7[1]),.doutc(w_n14816_7[2]),.din(w_n14816_2[0]));
	jspl jspl_w_n14816_8(.douta(w_n14816_8[0]),.doutb(w_n14816_8[1]),.din(w_n14816_2[1]));
	jspl3 jspl3_w_n14821_0(.douta(w_n14821_0[0]),.doutb(w_n14821_0[1]),.doutc(w_n14821_0[2]),.din(n14821));
	jspl3 jspl3_w_n14821_1(.douta(w_n14821_1[0]),.doutb(w_n14821_1[1]),.doutc(w_n14821_1[2]),.din(w_n14821_0[0]));
	jspl3 jspl3_w_n14821_2(.douta(w_n14821_2[0]),.doutb(w_n14821_2[1]),.doutc(w_n14821_2[2]),.din(w_n14821_0[1]));
	jspl3 jspl3_w_n14821_3(.douta(w_n14821_3[0]),.doutb(w_n14821_3[1]),.doutc(w_n14821_3[2]),.din(w_n14821_0[2]));
	jspl3 jspl3_w_n14821_4(.douta(w_n14821_4[0]),.doutb(w_n14821_4[1]),.doutc(w_n14821_4[2]),.din(w_n14821_1[0]));
	jspl3 jspl3_w_n14821_5(.douta(w_n14821_5[0]),.doutb(w_n14821_5[1]),.doutc(w_n14821_5[2]),.din(w_n14821_1[1]));
	jspl3 jspl3_w_n14821_6(.douta(w_n14821_6[0]),.doutb(w_n14821_6[1]),.doutc(w_n14821_6[2]),.din(w_n14821_1[2]));
	jspl3 jspl3_w_n14821_7(.douta(w_n14821_7[0]),.doutb(w_n14821_7[1]),.doutc(w_n14821_7[2]),.din(w_n14821_2[0]));
	jspl3 jspl3_w_n14821_8(.douta(w_n14821_8[0]),.doutb(w_n14821_8[1]),.doutc(w_n14821_8[2]),.din(w_n14821_2[1]));
	jspl3 jspl3_w_n14821_9(.douta(w_n14821_9[0]),.doutb(w_n14821_9[1]),.doutc(w_n14821_9[2]),.din(w_n14821_2[2]));
	jspl3 jspl3_w_n14821_10(.douta(w_n14821_10[0]),.doutb(w_n14821_10[1]),.doutc(w_n14821_10[2]),.din(w_n14821_3[0]));
	jspl3 jspl3_w_n14821_11(.douta(w_n14821_11[0]),.doutb(w_n14821_11[1]),.doutc(w_n14821_11[2]),.din(w_n14821_3[1]));
	jspl3 jspl3_w_n14821_12(.douta(w_n14821_12[0]),.doutb(w_n14821_12[1]),.doutc(w_n14821_12[2]),.din(w_n14821_3[2]));
	jspl3 jspl3_w_n14821_13(.douta(w_n14821_13[0]),.doutb(w_n14821_13[1]),.doutc(w_n14821_13[2]),.din(w_n14821_4[0]));
	jspl3 jspl3_w_n14821_14(.douta(w_n14821_14[0]),.doutb(w_n14821_14[1]),.doutc(w_n14821_14[2]),.din(w_n14821_4[1]));
	jspl3 jspl3_w_n14821_15(.douta(w_n14821_15[0]),.doutb(w_n14821_15[1]),.doutc(w_n14821_15[2]),.din(w_n14821_4[2]));
	jspl3 jspl3_w_n14821_16(.douta(w_n14821_16[0]),.doutb(w_n14821_16[1]),.doutc(w_n14821_16[2]),.din(w_n14821_5[0]));
	jspl3 jspl3_w_n14821_17(.douta(w_n14821_17[0]),.doutb(w_n14821_17[1]),.doutc(w_n14821_17[2]),.din(w_n14821_5[1]));
	jspl3 jspl3_w_n14821_18(.douta(w_n14821_18[0]),.doutb(w_n14821_18[1]),.doutc(w_n14821_18[2]),.din(w_n14821_5[2]));
	jspl3 jspl3_w_n14821_19(.douta(w_n14821_19[0]),.doutb(w_n14821_19[1]),.doutc(w_n14821_19[2]),.din(w_n14821_6[0]));
	jspl3 jspl3_w_n14821_20(.douta(w_n14821_20[0]),.doutb(w_n14821_20[1]),.doutc(w_n14821_20[2]),.din(w_n14821_6[1]));
	jspl3 jspl3_w_n14821_21(.douta(w_n14821_21[0]),.doutb(w_n14821_21[1]),.doutc(w_n14821_21[2]),.din(w_n14821_6[2]));
	jspl3 jspl3_w_n14821_22(.douta(w_n14821_22[0]),.doutb(w_n14821_22[1]),.doutc(w_n14821_22[2]),.din(w_n14821_7[0]));
	jspl jspl_w_n14824_0(.douta(w_n14824_0[0]),.doutb(w_n14824_0[1]),.din(n14824));
	jspl3 jspl3_w_n14826_0(.douta(w_n14826_0[0]),.doutb(w_n14826_0[1]),.doutc(w_n14826_0[2]),.din(n14826));
	jspl jspl_w_n14826_1(.douta(w_n14826_1[0]),.doutb(w_n14826_1[1]),.din(w_n14826_0[0]));
	jspl3 jspl3_w_n14827_0(.douta(w_n14827_0[0]),.doutb(w_n14827_0[1]),.doutc(w_n14827_0[2]),.din(n14827));
	jspl3 jspl3_w_n14831_0(.douta(w_n14831_0[0]),.doutb(w_n14831_0[1]),.doutc(w_n14831_0[2]),.din(n14831));
	jspl jspl_w_n14832_0(.douta(w_n14832_0[0]),.doutb(w_n14832_0[1]),.din(n14832));
	jspl jspl_w_n14833_0(.douta(w_n14833_0[0]),.doutb(w_n14833_0[1]),.din(n14833));
	jspl jspl_w_n14834_0(.douta(w_n14834_0[0]),.doutb(w_n14834_0[1]),.din(n14834));
	jspl jspl_w_n14836_0(.douta(w_n14836_0[0]),.doutb(w_n14836_0[1]),.din(n14836));
	jspl jspl_w_n14838_0(.douta(w_n14838_0[0]),.doutb(w_n14838_0[1]),.din(n14838));
	jspl jspl_w_n14840_0(.douta(w_n14840_0[0]),.doutb(w_n14840_0[1]),.din(n14840));
	jspl jspl_w_n14843_0(.douta(w_n14843_0[0]),.doutb(w_n14843_0[1]),.din(n14843));
	jspl jspl_w_n14848_0(.douta(w_n14848_0[0]),.doutb(w_n14848_0[1]),.din(n14848));
	jspl3 jspl3_w_n14850_0(.douta(w_n14850_0[0]),.doutb(w_n14850_0[1]),.doutc(w_n14850_0[2]),.din(n14850));
	jspl jspl_w_n14851_0(.douta(w_n14851_0[0]),.doutb(w_n14851_0[1]),.din(n14851));
	jspl jspl_w_n14855_0(.douta(w_n14855_0[0]),.doutb(w_n14855_0[1]),.din(n14855));
	jspl jspl_w_n14856_0(.douta(w_n14856_0[0]),.doutb(w_n14856_0[1]),.din(n14856));
	jspl jspl_w_n14858_0(.douta(w_n14858_0[0]),.doutb(w_n14858_0[1]),.din(n14858));
	jspl jspl_w_n14862_0(.douta(w_n14862_0[0]),.doutb(w_n14862_0[1]),.din(n14862));
	jspl jspl_w_n14864_0(.douta(w_n14864_0[0]),.doutb(w_n14864_0[1]),.din(n14864));
	jspl jspl_w_n14865_0(.douta(w_n14865_0[0]),.doutb(w_n14865_0[1]),.din(n14865));
	jspl3 jspl3_w_n14866_0(.douta(w_n14866_0[0]),.doutb(w_n14866_0[1]),.doutc(w_n14866_0[2]),.din(n14866));
	jspl jspl_w_n14867_0(.douta(w_n14867_0[0]),.doutb(w_n14867_0[1]),.din(n14867));
	jspl jspl_w_n14871_0(.douta(w_n14871_0[0]),.doutb(w_n14871_0[1]),.din(n14871));
	jspl jspl_w_n14873_0(.douta(w_n14873_0[0]),.doutb(w_n14873_0[1]),.din(n14873));
	jspl jspl_w_n14875_0(.douta(w_n14875_0[0]),.doutb(w_n14875_0[1]),.din(n14875));
	jspl jspl_w_n14877_0(.douta(w_n14877_0[0]),.doutb(w_n14877_0[1]),.din(n14877));
	jspl jspl_w_n14880_0(.douta(w_n14880_0[0]),.doutb(w_n14880_0[1]),.din(n14880));
	jspl jspl_w_n14886_0(.douta(w_n14886_0[0]),.doutb(w_n14886_0[1]),.din(n14886));
	jspl3 jspl3_w_n14888_0(.douta(w_n14888_0[0]),.doutb(w_n14888_0[1]),.doutc(w_n14888_0[2]),.din(n14888));
	jspl jspl_w_n14889_0(.douta(w_n14889_0[0]),.doutb(w_n14889_0[1]),.din(n14889));
	jspl jspl_w_n14894_0(.douta(w_n14894_0[0]),.doutb(w_n14894_0[1]),.din(n14894));
	jspl jspl_w_n14896_0(.douta(w_n14896_0[0]),.doutb(w_n14896_0[1]),.din(n14896));
	jspl jspl_w_n14898_0(.douta(w_n14898_0[0]),.doutb(w_n14898_0[1]),.din(n14898));
	jspl jspl_w_n14902_0(.douta(w_n14902_0[0]),.doutb(w_n14902_0[1]),.din(n14902));
	jspl jspl_w_n14904_0(.douta(w_n14904_0[0]),.doutb(w_n14904_0[1]),.din(n14904));
	jspl jspl_w_n14905_0(.douta(w_n14905_0[0]),.doutb(w_n14905_0[1]),.din(n14905));
	jspl3 jspl3_w_n14906_0(.douta(w_n14906_0[0]),.doutb(w_n14906_0[1]),.doutc(w_n14906_0[2]),.din(n14906));
	jspl jspl_w_n14907_0(.douta(w_n14907_0[0]),.doutb(w_n14907_0[1]),.din(n14907));
	jspl jspl_w_n14913_0(.douta(w_n14913_0[0]),.doutb(w_n14913_0[1]),.din(n14913));
	jspl jspl_w_n14914_0(.douta(w_n14914_0[0]),.doutb(w_n14914_0[1]),.din(n14914));
	jspl jspl_w_n14916_0(.douta(w_n14916_0[0]),.doutb(w_n14916_0[1]),.din(n14916));
	jspl jspl_w_n14918_0(.douta(w_n14918_0[0]),.doutb(w_n14918_0[1]),.din(n14918));
	jspl jspl_w_n14920_0(.douta(w_n14920_0[0]),.doutb(w_n14920_0[1]),.din(n14920));
	jspl jspl_w_n14926_0(.douta(w_n14926_0[0]),.doutb(w_n14926_0[1]),.din(n14926));
	jspl jspl_w_n14928_0(.douta(w_n14928_0[0]),.doutb(w_n14928_0[1]),.din(n14928));
	jspl3 jspl3_w_n14929_0(.douta(w_n14929_0[0]),.doutb(w_n14929_0[1]),.doutc(w_n14929_0[2]),.din(n14929));
	jspl jspl_w_n14932_0(.douta(w_n14932_0[0]),.doutb(w_n14932_0[1]),.din(n14932));
	jspl jspl_w_n14933_0(.douta(w_n14933_0[0]),.doutb(w_n14933_0[1]),.din(n14933));
	jspl3 jspl3_w_n14934_0(.douta(w_n14934_0[0]),.doutb(w_n14934_0[1]),.doutc(w_n14934_0[2]),.din(n14934));
	jspl jspl_w_n14936_0(.douta(w_n14936_0[0]),.doutb(w_n14936_0[1]),.din(n14936));
	jspl jspl_w_n14940_0(.douta(w_n14940_0[0]),.doutb(w_n14940_0[1]),.din(n14940));
	jspl jspl_w_n14942_0(.douta(w_n14942_0[0]),.doutb(w_n14942_0[1]),.din(n14942));
	jspl jspl_w_n14943_0(.douta(w_n14943_0[0]),.doutb(w_n14943_0[1]),.din(n14943));
	jspl3 jspl3_w_n14944_0(.douta(w_n14944_0[0]),.doutb(w_n14944_0[1]),.doutc(w_n14944_0[2]),.din(n14944));
	jspl jspl_w_n14945_0(.douta(w_n14945_0[0]),.doutb(w_n14945_0[1]),.din(n14945));
	jspl jspl_w_n14948_0(.douta(w_n14948_0[0]),.doutb(w_n14948_0[1]),.din(n14948));
	jspl jspl_w_n14954_0(.douta(w_n14954_0[0]),.doutb(w_n14954_0[1]),.din(n14954));
	jspl jspl_w_n14955_0(.douta(w_n14955_0[0]),.doutb(w_n14955_0[1]),.din(n14955));
	jspl jspl_w_n14957_0(.douta(w_n14957_0[0]),.doutb(w_n14957_0[1]),.din(n14957));
	jspl jspl_w_n14959_0(.douta(w_n14959_0[0]),.doutb(w_n14959_0[1]),.din(n14959));
	jspl jspl_w_n14961_0(.douta(w_n14961_0[0]),.doutb(w_n14961_0[1]),.din(n14961));
	jspl jspl_w_n14967_0(.douta(w_n14967_0[0]),.doutb(w_n14967_0[1]),.din(n14967));
	jspl jspl_w_n14969_0(.douta(w_n14969_0[0]),.doutb(w_n14969_0[1]),.din(n14969));
	jspl3 jspl3_w_n14970_0(.douta(w_n14970_0[0]),.doutb(w_n14970_0[1]),.doutc(w_n14970_0[2]),.din(n14970));
	jspl jspl_w_n14973_0(.douta(w_n14973_0[0]),.doutb(w_n14973_0[1]),.din(n14973));
	jspl jspl_w_n14974_0(.douta(w_n14974_0[0]),.doutb(w_n14974_0[1]),.din(n14974));
	jspl3 jspl3_w_n14975_0(.douta(w_n14975_0[0]),.doutb(w_n14975_0[1]),.doutc(w_n14975_0[2]),.din(n14975));
	jspl jspl_w_n14977_0(.douta(w_n14977_0[0]),.doutb(w_n14977_0[1]),.din(n14977));
	jspl jspl_w_n14981_0(.douta(w_n14981_0[0]),.doutb(w_n14981_0[1]),.din(n14981));
	jspl jspl_w_n14983_0(.douta(w_n14983_0[0]),.doutb(w_n14983_0[1]),.din(n14983));
	jspl jspl_w_n14984_0(.douta(w_n14984_0[0]),.doutb(w_n14984_0[1]),.din(n14984));
	jspl3 jspl3_w_n14985_0(.douta(w_n14985_0[0]),.doutb(w_n14985_0[1]),.doutc(w_n14985_0[2]),.din(n14985));
	jspl jspl_w_n14986_0(.douta(w_n14986_0[0]),.doutb(w_n14986_0[1]),.din(n14986));
	jspl jspl_w_n14989_0(.douta(w_n14989_0[0]),.doutb(w_n14989_0[1]),.din(n14989));
	jspl jspl_w_n14995_0(.douta(w_n14995_0[0]),.doutb(w_n14995_0[1]),.din(n14995));
	jspl jspl_w_n14996_0(.douta(w_n14996_0[0]),.doutb(w_n14996_0[1]),.din(n14996));
	jspl jspl_w_n14998_0(.douta(w_n14998_0[0]),.doutb(w_n14998_0[1]),.din(n14998));
	jspl jspl_w_n15000_0(.douta(w_n15000_0[0]),.doutb(w_n15000_0[1]),.din(n15000));
	jspl jspl_w_n15002_0(.douta(w_n15002_0[0]),.doutb(w_n15002_0[1]),.din(n15002));
	jspl jspl_w_n15008_0(.douta(w_n15008_0[0]),.doutb(w_n15008_0[1]),.din(n15008));
	jspl jspl_w_n15010_0(.douta(w_n15010_0[0]),.doutb(w_n15010_0[1]),.din(n15010));
	jspl3 jspl3_w_n15011_0(.douta(w_n15011_0[0]),.doutb(w_n15011_0[1]),.doutc(w_n15011_0[2]),.din(n15011));
	jspl jspl_w_n15014_0(.douta(w_n15014_0[0]),.doutb(w_n15014_0[1]),.din(n15014));
	jspl jspl_w_n15015_0(.douta(w_n15015_0[0]),.doutb(w_n15015_0[1]),.din(n15015));
	jspl3 jspl3_w_n15016_0(.douta(w_n15016_0[0]),.doutb(w_n15016_0[1]),.doutc(w_n15016_0[2]),.din(n15016));
	jspl jspl_w_n15018_0(.douta(w_n15018_0[0]),.doutb(w_n15018_0[1]),.din(n15018));
	jspl jspl_w_n15022_0(.douta(w_n15022_0[0]),.doutb(w_n15022_0[1]),.din(n15022));
	jspl jspl_w_n15024_0(.douta(w_n15024_0[0]),.doutb(w_n15024_0[1]),.din(n15024));
	jspl jspl_w_n15025_0(.douta(w_n15025_0[0]),.doutb(w_n15025_0[1]),.din(n15025));
	jspl3 jspl3_w_n15026_0(.douta(w_n15026_0[0]),.doutb(w_n15026_0[1]),.doutc(w_n15026_0[2]),.din(n15026));
	jspl jspl_w_n15027_0(.douta(w_n15027_0[0]),.doutb(w_n15027_0[1]),.din(n15027));
	jspl jspl_w_n15030_0(.douta(w_n15030_0[0]),.doutb(w_n15030_0[1]),.din(n15030));
	jspl jspl_w_n15036_0(.douta(w_n15036_0[0]),.doutb(w_n15036_0[1]),.din(n15036));
	jspl jspl_w_n15037_0(.douta(w_n15037_0[0]),.doutb(w_n15037_0[1]),.din(n15037));
	jspl jspl_w_n15039_0(.douta(w_n15039_0[0]),.doutb(w_n15039_0[1]),.din(n15039));
	jspl jspl_w_n15041_0(.douta(w_n15041_0[0]),.doutb(w_n15041_0[1]),.din(n15041));
	jspl jspl_w_n15043_0(.douta(w_n15043_0[0]),.doutb(w_n15043_0[1]),.din(n15043));
	jspl jspl_w_n15049_0(.douta(w_n15049_0[0]),.doutb(w_n15049_0[1]),.din(n15049));
	jspl jspl_w_n15051_0(.douta(w_n15051_0[0]),.doutb(w_n15051_0[1]),.din(n15051));
	jspl3 jspl3_w_n15052_0(.douta(w_n15052_0[0]),.doutb(w_n15052_0[1]),.doutc(w_n15052_0[2]),.din(n15052));
	jspl jspl_w_n15055_0(.douta(w_n15055_0[0]),.doutb(w_n15055_0[1]),.din(n15055));
	jspl jspl_w_n15056_0(.douta(w_n15056_0[0]),.doutb(w_n15056_0[1]),.din(n15056));
	jspl3 jspl3_w_n15057_0(.douta(w_n15057_0[0]),.doutb(w_n15057_0[1]),.doutc(w_n15057_0[2]),.din(n15057));
	jspl jspl_w_n15059_0(.douta(w_n15059_0[0]),.doutb(w_n15059_0[1]),.din(n15059));
	jspl jspl_w_n15063_0(.douta(w_n15063_0[0]),.doutb(w_n15063_0[1]),.din(n15063));
	jspl jspl_w_n15065_0(.douta(w_n15065_0[0]),.doutb(w_n15065_0[1]),.din(n15065));
	jspl jspl_w_n15066_0(.douta(w_n15066_0[0]),.doutb(w_n15066_0[1]),.din(n15066));
	jspl3 jspl3_w_n15067_0(.douta(w_n15067_0[0]),.doutb(w_n15067_0[1]),.doutc(w_n15067_0[2]),.din(n15067));
	jspl jspl_w_n15068_0(.douta(w_n15068_0[0]),.doutb(w_n15068_0[1]),.din(n15068));
	jspl jspl_w_n15071_0(.douta(w_n15071_0[0]),.doutb(w_n15071_0[1]),.din(n15071));
	jspl jspl_w_n15077_0(.douta(w_n15077_0[0]),.doutb(w_n15077_0[1]),.din(n15077));
	jspl jspl_w_n15078_0(.douta(w_n15078_0[0]),.doutb(w_n15078_0[1]),.din(n15078));
	jspl jspl_w_n15080_0(.douta(w_n15080_0[0]),.doutb(w_n15080_0[1]),.din(n15080));
	jspl jspl_w_n15082_0(.douta(w_n15082_0[0]),.doutb(w_n15082_0[1]),.din(n15082));
	jspl jspl_w_n15084_0(.douta(w_n15084_0[0]),.doutb(w_n15084_0[1]),.din(n15084));
	jspl jspl_w_n15090_0(.douta(w_n15090_0[0]),.doutb(w_n15090_0[1]),.din(n15090));
	jspl jspl_w_n15092_0(.douta(w_n15092_0[0]),.doutb(w_n15092_0[1]),.din(n15092));
	jspl3 jspl3_w_n15093_0(.douta(w_n15093_0[0]),.doutb(w_n15093_0[1]),.doutc(w_n15093_0[2]),.din(n15093));
	jspl jspl_w_n15096_0(.douta(w_n15096_0[0]),.doutb(w_n15096_0[1]),.din(n15096));
	jspl jspl_w_n15097_0(.douta(w_n15097_0[0]),.doutb(w_n15097_0[1]),.din(n15097));
	jspl3 jspl3_w_n15098_0(.douta(w_n15098_0[0]),.doutb(w_n15098_0[1]),.doutc(w_n15098_0[2]),.din(n15098));
	jspl jspl_w_n15100_0(.douta(w_n15100_0[0]),.doutb(w_n15100_0[1]),.din(n15100));
	jspl jspl_w_n15104_0(.douta(w_n15104_0[0]),.doutb(w_n15104_0[1]),.din(n15104));
	jspl jspl_w_n15106_0(.douta(w_n15106_0[0]),.doutb(w_n15106_0[1]),.din(n15106));
	jspl jspl_w_n15107_0(.douta(w_n15107_0[0]),.doutb(w_n15107_0[1]),.din(n15107));
	jspl3 jspl3_w_n15108_0(.douta(w_n15108_0[0]),.doutb(w_n15108_0[1]),.doutc(w_n15108_0[2]),.din(n15108));
	jspl jspl_w_n15109_0(.douta(w_n15109_0[0]),.doutb(w_n15109_0[1]),.din(n15109));
	jspl jspl_w_n15112_0(.douta(w_n15112_0[0]),.doutb(w_n15112_0[1]),.din(n15112));
	jspl jspl_w_n15118_0(.douta(w_n15118_0[0]),.doutb(w_n15118_0[1]),.din(n15118));
	jspl jspl_w_n15119_0(.douta(w_n15119_0[0]),.doutb(w_n15119_0[1]),.din(n15119));
	jspl jspl_w_n15121_0(.douta(w_n15121_0[0]),.doutb(w_n15121_0[1]),.din(n15121));
	jspl jspl_w_n15123_0(.douta(w_n15123_0[0]),.doutb(w_n15123_0[1]),.din(n15123));
	jspl jspl_w_n15125_0(.douta(w_n15125_0[0]),.doutb(w_n15125_0[1]),.din(n15125));
	jspl jspl_w_n15131_0(.douta(w_n15131_0[0]),.doutb(w_n15131_0[1]),.din(n15131));
	jspl jspl_w_n15133_0(.douta(w_n15133_0[0]),.doutb(w_n15133_0[1]),.din(n15133));
	jspl3 jspl3_w_n15134_0(.douta(w_n15134_0[0]),.doutb(w_n15134_0[1]),.doutc(w_n15134_0[2]),.din(n15134));
	jspl jspl_w_n15137_0(.douta(w_n15137_0[0]),.doutb(w_n15137_0[1]),.din(n15137));
	jspl jspl_w_n15138_0(.douta(w_n15138_0[0]),.doutb(w_n15138_0[1]),.din(n15138));
	jspl3 jspl3_w_n15139_0(.douta(w_n15139_0[0]),.doutb(w_n15139_0[1]),.doutc(w_n15139_0[2]),.din(n15139));
	jspl jspl_w_n15141_0(.douta(w_n15141_0[0]),.doutb(w_n15141_0[1]),.din(n15141));
	jspl jspl_w_n15145_0(.douta(w_n15145_0[0]),.doutb(w_n15145_0[1]),.din(n15145));
	jspl jspl_w_n15147_0(.douta(w_n15147_0[0]),.doutb(w_n15147_0[1]),.din(n15147));
	jspl jspl_w_n15148_0(.douta(w_n15148_0[0]),.doutb(w_n15148_0[1]),.din(n15148));
	jspl3 jspl3_w_n15149_0(.douta(w_n15149_0[0]),.doutb(w_n15149_0[1]),.doutc(w_n15149_0[2]),.din(n15149));
	jspl jspl_w_n15150_0(.douta(w_n15150_0[0]),.doutb(w_n15150_0[1]),.din(n15150));
	jspl jspl_w_n15153_0(.douta(w_n15153_0[0]),.doutb(w_n15153_0[1]),.din(n15153));
	jspl jspl_w_n15159_0(.douta(w_n15159_0[0]),.doutb(w_n15159_0[1]),.din(n15159));
	jspl jspl_w_n15160_0(.douta(w_n15160_0[0]),.doutb(w_n15160_0[1]),.din(n15160));
	jspl jspl_w_n15162_0(.douta(w_n15162_0[0]),.doutb(w_n15162_0[1]),.din(n15162));
	jspl jspl_w_n15164_0(.douta(w_n15164_0[0]),.doutb(w_n15164_0[1]),.din(n15164));
	jspl jspl_w_n15166_0(.douta(w_n15166_0[0]),.doutb(w_n15166_0[1]),.din(n15166));
	jspl jspl_w_n15172_0(.douta(w_n15172_0[0]),.doutb(w_n15172_0[1]),.din(n15172));
	jspl jspl_w_n15174_0(.douta(w_n15174_0[0]),.doutb(w_n15174_0[1]),.din(n15174));
	jspl3 jspl3_w_n15175_0(.douta(w_n15175_0[0]),.doutb(w_n15175_0[1]),.doutc(w_n15175_0[2]),.din(n15175));
	jspl jspl_w_n15178_0(.douta(w_n15178_0[0]),.doutb(w_n15178_0[1]),.din(n15178));
	jspl jspl_w_n15179_0(.douta(w_n15179_0[0]),.doutb(w_n15179_0[1]),.din(n15179));
	jspl3 jspl3_w_n15180_0(.douta(w_n15180_0[0]),.doutb(w_n15180_0[1]),.doutc(w_n15180_0[2]),.din(n15180));
	jspl jspl_w_n15182_0(.douta(w_n15182_0[0]),.doutb(w_n15182_0[1]),.din(n15182));
	jspl jspl_w_n15186_0(.douta(w_n15186_0[0]),.doutb(w_n15186_0[1]),.din(n15186));
	jspl jspl_w_n15188_0(.douta(w_n15188_0[0]),.doutb(w_n15188_0[1]),.din(n15188));
	jspl jspl_w_n15189_0(.douta(w_n15189_0[0]),.doutb(w_n15189_0[1]),.din(n15189));
	jspl3 jspl3_w_n15190_0(.douta(w_n15190_0[0]),.doutb(w_n15190_0[1]),.doutc(w_n15190_0[2]),.din(n15190));
	jspl jspl_w_n15191_0(.douta(w_n15191_0[0]),.doutb(w_n15191_0[1]),.din(n15191));
	jspl jspl_w_n15194_0(.douta(w_n15194_0[0]),.doutb(w_n15194_0[1]),.din(n15194));
	jspl jspl_w_n15200_0(.douta(w_n15200_0[0]),.doutb(w_n15200_0[1]),.din(n15200));
	jspl jspl_w_n15201_0(.douta(w_n15201_0[0]),.doutb(w_n15201_0[1]),.din(n15201));
	jspl jspl_w_n15203_0(.douta(w_n15203_0[0]),.doutb(w_n15203_0[1]),.din(n15203));
	jspl jspl_w_n15205_0(.douta(w_n15205_0[0]),.doutb(w_n15205_0[1]),.din(n15205));
	jspl jspl_w_n15207_0(.douta(w_n15207_0[0]),.doutb(w_n15207_0[1]),.din(n15207));
	jspl jspl_w_n15213_0(.douta(w_n15213_0[0]),.doutb(w_n15213_0[1]),.din(n15213));
	jspl jspl_w_n15215_0(.douta(w_n15215_0[0]),.doutb(w_n15215_0[1]),.din(n15215));
	jspl3 jspl3_w_n15216_0(.douta(w_n15216_0[0]),.doutb(w_n15216_0[1]),.doutc(w_n15216_0[2]),.din(n15216));
	jspl jspl_w_n15219_0(.douta(w_n15219_0[0]),.doutb(w_n15219_0[1]),.din(n15219));
	jspl jspl_w_n15220_0(.douta(w_n15220_0[0]),.doutb(w_n15220_0[1]),.din(n15220));
	jspl3 jspl3_w_n15221_0(.douta(w_n15221_0[0]),.doutb(w_n15221_0[1]),.doutc(w_n15221_0[2]),.din(n15221));
	jspl jspl_w_n15223_0(.douta(w_n15223_0[0]),.doutb(w_n15223_0[1]),.din(n15223));
	jspl jspl_w_n15225_0(.douta(w_n15225_0[0]),.doutb(w_n15225_0[1]),.din(n15225));
	jspl jspl_w_n15227_0(.douta(w_n15227_0[0]),.doutb(w_n15227_0[1]),.din(n15227));
	jspl jspl_w_n15233_0(.douta(w_n15233_0[0]),.doutb(w_n15233_0[1]),.din(n15233));
	jspl3 jspl3_w_n15235_0(.douta(w_n15235_0[0]),.doutb(w_n15235_0[1]),.doutc(w_n15235_0[2]),.din(n15235));
	jspl jspl_w_n15236_0(.douta(w_n15236_0[0]),.doutb(w_n15236_0[1]),.din(n15236));
	jspl jspl_w_n15239_0(.douta(w_n15239_0[0]),.doutb(w_n15239_0[1]),.din(n15239));
	jspl jspl_w_n15241_0(.douta(w_n15241_0[0]),.doutb(w_n15241_0[1]),.din(n15241));
	jspl jspl_w_n15245_0(.douta(w_n15245_0[0]),.doutb(w_n15245_0[1]),.din(n15245));
	jspl jspl_w_n15247_0(.douta(w_n15247_0[0]),.doutb(w_n15247_0[1]),.din(n15247));
	jspl jspl_w_n15248_0(.douta(w_n15248_0[0]),.doutb(w_n15248_0[1]),.din(n15248));
	jspl jspl_w_n15249_0(.douta(w_n15249_0[0]),.doutb(w_n15249_0[1]),.din(n15249));
	jspl3 jspl3_w_n15250_0(.douta(w_n15250_0[0]),.doutb(w_n15250_0[1]),.doutc(w_n15250_0[2]),.din(n15250));
	jspl jspl_w_n15253_0(.douta(w_n15253_0[0]),.doutb(w_n15253_0[1]),.din(n15253));
	jspl jspl_w_n15254_0(.douta(w_n15254_0[0]),.doutb(w_n15254_0[1]),.din(n15254));
	jspl3 jspl3_w_n15255_0(.douta(w_n15255_0[0]),.doutb(w_n15255_0[1]),.doutc(w_n15255_0[2]),.din(n15255));
	jspl jspl_w_n15257_0(.douta(w_n15257_0[0]),.doutb(w_n15257_0[1]),.din(n15257));
	jspl jspl_w_n15261_0(.douta(w_n15261_0[0]),.doutb(w_n15261_0[1]),.din(n15261));
	jspl jspl_w_n15263_0(.douta(w_n15263_0[0]),.doutb(w_n15263_0[1]),.din(n15263));
	jspl jspl_w_n15264_0(.douta(w_n15264_0[0]),.doutb(w_n15264_0[1]),.din(n15264));
	jspl3 jspl3_w_n15265_0(.douta(w_n15265_0[0]),.doutb(w_n15265_0[1]),.doutc(w_n15265_0[2]),.din(n15265));
	jspl jspl_w_n15266_0(.douta(w_n15266_0[0]),.doutb(w_n15266_0[1]),.din(n15266));
	jspl jspl_w_n15269_0(.douta(w_n15269_0[0]),.doutb(w_n15269_0[1]),.din(n15269));
	jspl jspl_w_n15275_0(.douta(w_n15275_0[0]),.doutb(w_n15275_0[1]),.din(n15275));
	jspl jspl_w_n15276_0(.douta(w_n15276_0[0]),.doutb(w_n15276_0[1]),.din(n15276));
	jspl jspl_w_n15278_0(.douta(w_n15278_0[0]),.doutb(w_n15278_0[1]),.din(n15278));
	jspl jspl_w_n15280_0(.douta(w_n15280_0[0]),.doutb(w_n15280_0[1]),.din(n15280));
	jspl jspl_w_n15282_0(.douta(w_n15282_0[0]),.doutb(w_n15282_0[1]),.din(n15282));
	jspl jspl_w_n15288_0(.douta(w_n15288_0[0]),.doutb(w_n15288_0[1]),.din(n15288));
	jspl jspl_w_n15290_0(.douta(w_n15290_0[0]),.doutb(w_n15290_0[1]),.din(n15290));
	jspl3 jspl3_w_n15291_0(.douta(w_n15291_0[0]),.doutb(w_n15291_0[1]),.doutc(w_n15291_0[2]),.din(n15291));
	jspl jspl_w_n15294_0(.douta(w_n15294_0[0]),.doutb(w_n15294_0[1]),.din(n15294));
	jspl jspl_w_n15295_0(.douta(w_n15295_0[0]),.doutb(w_n15295_0[1]),.din(n15295));
	jspl3 jspl3_w_n15296_0(.douta(w_n15296_0[0]),.doutb(w_n15296_0[1]),.doutc(w_n15296_0[2]),.din(n15296));
	jspl jspl_w_n15298_0(.douta(w_n15298_0[0]),.doutb(w_n15298_0[1]),.din(n15298));
	jspl jspl_w_n15302_0(.douta(w_n15302_0[0]),.doutb(w_n15302_0[1]),.din(n15302));
	jspl jspl_w_n15304_0(.douta(w_n15304_0[0]),.doutb(w_n15304_0[1]),.din(n15304));
	jspl jspl_w_n15305_0(.douta(w_n15305_0[0]),.doutb(w_n15305_0[1]),.din(n15305));
	jspl3 jspl3_w_n15306_0(.douta(w_n15306_0[0]),.doutb(w_n15306_0[1]),.doutc(w_n15306_0[2]),.din(n15306));
	jspl jspl_w_n15307_0(.douta(w_n15307_0[0]),.doutb(w_n15307_0[1]),.din(n15307));
	jspl jspl_w_n15310_0(.douta(w_n15310_0[0]),.doutb(w_n15310_0[1]),.din(n15310));
	jspl jspl_w_n15316_0(.douta(w_n15316_0[0]),.doutb(w_n15316_0[1]),.din(n15316));
	jspl jspl_w_n15317_0(.douta(w_n15317_0[0]),.doutb(w_n15317_0[1]),.din(n15317));
	jspl jspl_w_n15319_0(.douta(w_n15319_0[0]),.doutb(w_n15319_0[1]),.din(n15319));
	jspl jspl_w_n15321_0(.douta(w_n15321_0[0]),.doutb(w_n15321_0[1]),.din(n15321));
	jspl jspl_w_n15323_0(.douta(w_n15323_0[0]),.doutb(w_n15323_0[1]),.din(n15323));
	jspl jspl_w_n15329_0(.douta(w_n15329_0[0]),.doutb(w_n15329_0[1]),.din(n15329));
	jspl3 jspl3_w_n15331_0(.douta(w_n15331_0[0]),.doutb(w_n15331_0[1]),.doutc(w_n15331_0[2]),.din(n15331));
	jspl jspl_w_n15336_0(.douta(w_n15336_0[0]),.doutb(w_n15336_0[1]),.din(n15336));
	jspl3 jspl3_w_n15338_0(.douta(w_n15338_0[0]),.doutb(w_n15338_0[1]),.doutc(w_n15338_0[2]),.din(n15338));
	jspl3 jspl3_w_n15342_0(.douta(w_n15342_0[0]),.doutb(w_n15342_0[1]),.doutc(w_n15342_0[2]),.din(n15342));
	jspl jspl_w_n15343_0(.douta(w_n15343_0[0]),.doutb(w_n15343_0[1]),.din(n15343));
	jspl jspl_w_n15348_0(.douta(w_n15348_0[0]),.doutb(w_n15348_0[1]),.din(n15348));
	jspl3 jspl3_w_n15349_0(.douta(w_n15349_0[0]),.doutb(w_n15349_0[1]),.doutc(w_n15349_0[2]),.din(n15349));
	jspl jspl_w_n15354_0(.douta(w_n15354_0[0]),.doutb(w_n15354_0[1]),.din(n15354));
	jspl jspl_w_n15361_0(.douta(w_n15361_0[0]),.doutb(w_n15361_0[1]),.din(n15361));
	jspl3 jspl3_w_n15364_0(.douta(w_n15364_0[0]),.doutb(w_n15364_0[1]),.doutc(w_n15364_0[2]),.din(n15364));
	jspl jspl_w_n15364_1(.douta(w_n15364_1[0]),.doutb(w_n15364_1[1]),.din(w_n15364_0[0]));
	jspl jspl_w_n15365_0(.douta(w_n15365_0[0]),.doutb(w_n15365_0[1]),.din(n15365));
	jspl3 jspl3_w_n15368_0(.douta(w_n15368_0[0]),.doutb(w_n15368_0[1]),.doutc(w_n15368_0[2]),.din(n15368));
	jspl jspl_w_n15369_0(.douta(w_n15369_0[0]),.doutb(w_n15369_0[1]),.din(n15369));
	jspl jspl_w_n15370_0(.douta(w_n15370_0[0]),.doutb(w_n15370_0[1]),.din(n15370));
	jspl jspl_w_n15371_0(.douta(w_n15371_0[0]),.doutb(w_n15371_0[1]),.din(n15371));
	jspl jspl_w_n15373_0(.douta(w_n15373_0[0]),.doutb(w_n15373_0[1]),.din(n15373));
	jspl jspl_w_n15375_0(.douta(w_n15375_0[0]),.doutb(w_n15375_0[1]),.din(n15375));
	jspl jspl_w_n15377_0(.douta(w_n15377_0[0]),.doutb(w_n15377_0[1]),.din(n15377));
	jspl jspl_w_n15386_0(.douta(w_n15386_0[0]),.doutb(w_n15386_0[1]),.din(n15386));
	jspl3 jspl3_w_n15388_0(.douta(w_n15388_0[0]),.doutb(w_n15388_0[1]),.doutc(w_n15388_0[2]),.din(n15388));
	jspl jspl_w_n15389_0(.douta(w_n15389_0[0]),.doutb(w_n15389_0[1]),.din(n15389));
	jspl jspl_w_n15393_0(.douta(w_n15393_0[0]),.doutb(w_n15393_0[1]),.din(n15393));
	jspl jspl_w_n15395_0(.douta(w_n15395_0[0]),.doutb(w_n15395_0[1]),.din(n15395));
	jspl jspl_w_n15397_0(.douta(w_n15397_0[0]),.doutb(w_n15397_0[1]),.din(n15397));
	jspl jspl_w_n15402_0(.douta(w_n15402_0[0]),.doutb(w_n15402_0[1]),.din(n15402));
	jspl jspl_w_n15404_0(.douta(w_n15404_0[0]),.doutb(w_n15404_0[1]),.din(n15404));
	jspl jspl_w_n15405_0(.douta(w_n15405_0[0]),.doutb(w_n15405_0[1]),.din(n15405));
	jspl3 jspl3_w_n15406_0(.douta(w_n15406_0[0]),.doutb(w_n15406_0[1]),.doutc(w_n15406_0[2]),.din(n15406));
	jspl jspl_w_n15407_0(.douta(w_n15407_0[0]),.doutb(w_n15407_0[1]),.din(n15407));
	jspl jspl_w_n15412_0(.douta(w_n15412_0[0]),.doutb(w_n15412_0[1]),.din(n15412));
	jspl jspl_w_n15413_0(.douta(w_n15413_0[0]),.doutb(w_n15413_0[1]),.din(n15413));
	jspl jspl_w_n15415_0(.douta(w_n15415_0[0]),.doutb(w_n15415_0[1]),.din(n15415));
	jspl jspl_w_n15417_0(.douta(w_n15417_0[0]),.doutb(w_n15417_0[1]),.din(n15417));
	jspl jspl_w_n15420_0(.douta(w_n15420_0[0]),.doutb(w_n15420_0[1]),.din(n15420));
	jspl jspl_w_n15426_0(.douta(w_n15426_0[0]),.doutb(w_n15426_0[1]),.din(n15426));
	jspl3 jspl3_w_n15428_0(.douta(w_n15428_0[0]),.doutb(w_n15428_0[1]),.doutc(w_n15428_0[2]),.din(n15428));
	jspl jspl_w_n15429_0(.douta(w_n15429_0[0]),.doutb(w_n15429_0[1]),.din(n15429));
	jspl jspl_w_n15433_0(.douta(w_n15433_0[0]),.doutb(w_n15433_0[1]),.din(n15433));
	jspl jspl_w_n15434_0(.douta(w_n15434_0[0]),.doutb(w_n15434_0[1]),.din(n15434));
	jspl jspl_w_n15436_0(.douta(w_n15436_0[0]),.doutb(w_n15436_0[1]),.din(n15436));
	jspl jspl_w_n15441_0(.douta(w_n15441_0[0]),.doutb(w_n15441_0[1]),.din(n15441));
	jspl jspl_w_n15443_0(.douta(w_n15443_0[0]),.doutb(w_n15443_0[1]),.din(n15443));
	jspl jspl_w_n15444_0(.douta(w_n15444_0[0]),.doutb(w_n15444_0[1]),.din(n15444));
	jspl3 jspl3_w_n15445_0(.douta(w_n15445_0[0]),.doutb(w_n15445_0[1]),.doutc(w_n15445_0[2]),.din(n15445));
	jspl jspl_w_n15446_0(.douta(w_n15446_0[0]),.doutb(w_n15446_0[1]),.din(n15446));
	jspl jspl_w_n15450_0(.douta(w_n15450_0[0]),.doutb(w_n15450_0[1]),.din(n15450));
	jspl jspl_w_n15451_0(.douta(w_n15451_0[0]),.doutb(w_n15451_0[1]),.din(n15451));
	jspl jspl_w_n15453_0(.douta(w_n15453_0[0]),.doutb(w_n15453_0[1]),.din(n15453));
	jspl jspl_w_n15455_0(.douta(w_n15455_0[0]),.doutb(w_n15455_0[1]),.din(n15455));
	jspl jspl_w_n15458_0(.douta(w_n15458_0[0]),.doutb(w_n15458_0[1]),.din(n15458));
	jspl jspl_w_n15464_0(.douta(w_n15464_0[0]),.doutb(w_n15464_0[1]),.din(n15464));
	jspl jspl_w_n15466_0(.douta(w_n15466_0[0]),.doutb(w_n15466_0[1]),.din(n15466));
	jspl3 jspl3_w_n15467_0(.douta(w_n15467_0[0]),.doutb(w_n15467_0[1]),.doutc(w_n15467_0[2]),.din(n15467));
	jspl jspl_w_n15471_0(.douta(w_n15471_0[0]),.doutb(w_n15471_0[1]),.din(n15471));
	jspl jspl_w_n15472_0(.douta(w_n15472_0[0]),.doutb(w_n15472_0[1]),.din(n15472));
	jspl3 jspl3_w_n15473_0(.douta(w_n15473_0[0]),.doutb(w_n15473_0[1]),.doutc(w_n15473_0[2]),.din(n15473));
	jspl jspl_w_n15475_0(.douta(w_n15475_0[0]),.doutb(w_n15475_0[1]),.din(n15475));
	jspl jspl_w_n15480_0(.douta(w_n15480_0[0]),.doutb(w_n15480_0[1]),.din(n15480));
	jspl jspl_w_n15482_0(.douta(w_n15482_0[0]),.doutb(w_n15482_0[1]),.din(n15482));
	jspl jspl_w_n15483_0(.douta(w_n15483_0[0]),.doutb(w_n15483_0[1]),.din(n15483));
	jspl3 jspl3_w_n15484_0(.douta(w_n15484_0[0]),.doutb(w_n15484_0[1]),.doutc(w_n15484_0[2]),.din(n15484));
	jspl jspl_w_n15485_0(.douta(w_n15485_0[0]),.doutb(w_n15485_0[1]),.din(n15485));
	jspl jspl_w_n15489_0(.douta(w_n15489_0[0]),.doutb(w_n15489_0[1]),.din(n15489));
	jspl jspl_w_n15495_0(.douta(w_n15495_0[0]),.doutb(w_n15495_0[1]),.din(n15495));
	jspl jspl_w_n15496_0(.douta(w_n15496_0[0]),.doutb(w_n15496_0[1]),.din(n15496));
	jspl jspl_w_n15498_0(.douta(w_n15498_0[0]),.doutb(w_n15498_0[1]),.din(n15498));
	jspl jspl_w_n15500_0(.douta(w_n15500_0[0]),.doutb(w_n15500_0[1]),.din(n15500));
	jspl jspl_w_n15503_0(.douta(w_n15503_0[0]),.doutb(w_n15503_0[1]),.din(n15503));
	jspl jspl_w_n15509_0(.douta(w_n15509_0[0]),.doutb(w_n15509_0[1]),.din(n15509));
	jspl jspl_w_n15511_0(.douta(w_n15511_0[0]),.doutb(w_n15511_0[1]),.din(n15511));
	jspl3 jspl3_w_n15512_0(.douta(w_n15512_0[0]),.doutb(w_n15512_0[1]),.doutc(w_n15512_0[2]),.din(n15512));
	jspl jspl_w_n15516_0(.douta(w_n15516_0[0]),.doutb(w_n15516_0[1]),.din(n15516));
	jspl jspl_w_n15517_0(.douta(w_n15517_0[0]),.doutb(w_n15517_0[1]),.din(n15517));
	jspl3 jspl3_w_n15518_0(.douta(w_n15518_0[0]),.doutb(w_n15518_0[1]),.doutc(w_n15518_0[2]),.din(n15518));
	jspl jspl_w_n15520_0(.douta(w_n15520_0[0]),.doutb(w_n15520_0[1]),.din(n15520));
	jspl jspl_w_n15525_0(.douta(w_n15525_0[0]),.doutb(w_n15525_0[1]),.din(n15525));
	jspl jspl_w_n15527_0(.douta(w_n15527_0[0]),.doutb(w_n15527_0[1]),.din(n15527));
	jspl jspl_w_n15528_0(.douta(w_n15528_0[0]),.doutb(w_n15528_0[1]),.din(n15528));
	jspl3 jspl3_w_n15529_0(.douta(w_n15529_0[0]),.doutb(w_n15529_0[1]),.doutc(w_n15529_0[2]),.din(n15529));
	jspl jspl_w_n15530_0(.douta(w_n15530_0[0]),.doutb(w_n15530_0[1]),.din(n15530));
	jspl jspl_w_n15534_0(.douta(w_n15534_0[0]),.doutb(w_n15534_0[1]),.din(n15534));
	jspl jspl_w_n15540_0(.douta(w_n15540_0[0]),.doutb(w_n15540_0[1]),.din(n15540));
	jspl jspl_w_n15541_0(.douta(w_n15541_0[0]),.doutb(w_n15541_0[1]),.din(n15541));
	jspl jspl_w_n15543_0(.douta(w_n15543_0[0]),.doutb(w_n15543_0[1]),.din(n15543));
	jspl jspl_w_n15545_0(.douta(w_n15545_0[0]),.doutb(w_n15545_0[1]),.din(n15545));
	jspl jspl_w_n15548_0(.douta(w_n15548_0[0]),.doutb(w_n15548_0[1]),.din(n15548));
	jspl jspl_w_n15554_0(.douta(w_n15554_0[0]),.doutb(w_n15554_0[1]),.din(n15554));
	jspl jspl_w_n15556_0(.douta(w_n15556_0[0]),.doutb(w_n15556_0[1]),.din(n15556));
	jspl3 jspl3_w_n15557_0(.douta(w_n15557_0[0]),.doutb(w_n15557_0[1]),.doutc(w_n15557_0[2]),.din(n15557));
	jspl jspl_w_n15561_0(.douta(w_n15561_0[0]),.doutb(w_n15561_0[1]),.din(n15561));
	jspl jspl_w_n15562_0(.douta(w_n15562_0[0]),.doutb(w_n15562_0[1]),.din(n15562));
	jspl3 jspl3_w_n15563_0(.douta(w_n15563_0[0]),.doutb(w_n15563_0[1]),.doutc(w_n15563_0[2]),.din(n15563));
	jspl jspl_w_n15565_0(.douta(w_n15565_0[0]),.doutb(w_n15565_0[1]),.din(n15565));
	jspl jspl_w_n15570_0(.douta(w_n15570_0[0]),.doutb(w_n15570_0[1]),.din(n15570));
	jspl jspl_w_n15572_0(.douta(w_n15572_0[0]),.doutb(w_n15572_0[1]),.din(n15572));
	jspl jspl_w_n15573_0(.douta(w_n15573_0[0]),.doutb(w_n15573_0[1]),.din(n15573));
	jspl3 jspl3_w_n15574_0(.douta(w_n15574_0[0]),.doutb(w_n15574_0[1]),.doutc(w_n15574_0[2]),.din(n15574));
	jspl jspl_w_n15575_0(.douta(w_n15575_0[0]),.doutb(w_n15575_0[1]),.din(n15575));
	jspl jspl_w_n15579_0(.douta(w_n15579_0[0]),.doutb(w_n15579_0[1]),.din(n15579));
	jspl jspl_w_n15585_0(.douta(w_n15585_0[0]),.doutb(w_n15585_0[1]),.din(n15585));
	jspl jspl_w_n15586_0(.douta(w_n15586_0[0]),.doutb(w_n15586_0[1]),.din(n15586));
	jspl jspl_w_n15588_0(.douta(w_n15588_0[0]),.doutb(w_n15588_0[1]),.din(n15588));
	jspl jspl_w_n15590_0(.douta(w_n15590_0[0]),.doutb(w_n15590_0[1]),.din(n15590));
	jspl jspl_w_n15593_0(.douta(w_n15593_0[0]),.doutb(w_n15593_0[1]),.din(n15593));
	jspl jspl_w_n15599_0(.douta(w_n15599_0[0]),.doutb(w_n15599_0[1]),.din(n15599));
	jspl jspl_w_n15601_0(.douta(w_n15601_0[0]),.doutb(w_n15601_0[1]),.din(n15601));
	jspl3 jspl3_w_n15602_0(.douta(w_n15602_0[0]),.doutb(w_n15602_0[1]),.doutc(w_n15602_0[2]),.din(n15602));
	jspl jspl_w_n15606_0(.douta(w_n15606_0[0]),.doutb(w_n15606_0[1]),.din(n15606));
	jspl jspl_w_n15607_0(.douta(w_n15607_0[0]),.doutb(w_n15607_0[1]),.din(n15607));
	jspl3 jspl3_w_n15608_0(.douta(w_n15608_0[0]),.doutb(w_n15608_0[1]),.doutc(w_n15608_0[2]),.din(n15608));
	jspl jspl_w_n15610_0(.douta(w_n15610_0[0]),.doutb(w_n15610_0[1]),.din(n15610));
	jspl jspl_w_n15615_0(.douta(w_n15615_0[0]),.doutb(w_n15615_0[1]),.din(n15615));
	jspl jspl_w_n15617_0(.douta(w_n15617_0[0]),.doutb(w_n15617_0[1]),.din(n15617));
	jspl jspl_w_n15618_0(.douta(w_n15618_0[0]),.doutb(w_n15618_0[1]),.din(n15618));
	jspl3 jspl3_w_n15619_0(.douta(w_n15619_0[0]),.doutb(w_n15619_0[1]),.doutc(w_n15619_0[2]),.din(n15619));
	jspl jspl_w_n15620_0(.douta(w_n15620_0[0]),.doutb(w_n15620_0[1]),.din(n15620));
	jspl jspl_w_n15624_0(.douta(w_n15624_0[0]),.doutb(w_n15624_0[1]),.din(n15624));
	jspl jspl_w_n15630_0(.douta(w_n15630_0[0]),.doutb(w_n15630_0[1]),.din(n15630));
	jspl jspl_w_n15631_0(.douta(w_n15631_0[0]),.doutb(w_n15631_0[1]),.din(n15631));
	jspl jspl_w_n15633_0(.douta(w_n15633_0[0]),.doutb(w_n15633_0[1]),.din(n15633));
	jspl jspl_w_n15635_0(.douta(w_n15635_0[0]),.doutb(w_n15635_0[1]),.din(n15635));
	jspl jspl_w_n15638_0(.douta(w_n15638_0[0]),.doutb(w_n15638_0[1]),.din(n15638));
	jspl jspl_w_n15644_0(.douta(w_n15644_0[0]),.doutb(w_n15644_0[1]),.din(n15644));
	jspl jspl_w_n15646_0(.douta(w_n15646_0[0]),.doutb(w_n15646_0[1]),.din(n15646));
	jspl3 jspl3_w_n15647_0(.douta(w_n15647_0[0]),.doutb(w_n15647_0[1]),.doutc(w_n15647_0[2]),.din(n15647));
	jspl jspl_w_n15651_0(.douta(w_n15651_0[0]),.doutb(w_n15651_0[1]),.din(n15651));
	jspl jspl_w_n15652_0(.douta(w_n15652_0[0]),.doutb(w_n15652_0[1]),.din(n15652));
	jspl3 jspl3_w_n15653_0(.douta(w_n15653_0[0]),.doutb(w_n15653_0[1]),.doutc(w_n15653_0[2]),.din(n15653));
	jspl jspl_w_n15655_0(.douta(w_n15655_0[0]),.doutb(w_n15655_0[1]),.din(n15655));
	jspl jspl_w_n15660_0(.douta(w_n15660_0[0]),.doutb(w_n15660_0[1]),.din(n15660));
	jspl jspl_w_n15662_0(.douta(w_n15662_0[0]),.doutb(w_n15662_0[1]),.din(n15662));
	jspl jspl_w_n15663_0(.douta(w_n15663_0[0]),.doutb(w_n15663_0[1]),.din(n15663));
	jspl3 jspl3_w_n15664_0(.douta(w_n15664_0[0]),.doutb(w_n15664_0[1]),.doutc(w_n15664_0[2]),.din(n15664));
	jspl jspl_w_n15665_0(.douta(w_n15665_0[0]),.doutb(w_n15665_0[1]),.din(n15665));
	jspl jspl_w_n15669_0(.douta(w_n15669_0[0]),.doutb(w_n15669_0[1]),.din(n15669));
	jspl jspl_w_n15675_0(.douta(w_n15675_0[0]),.doutb(w_n15675_0[1]),.din(n15675));
	jspl jspl_w_n15676_0(.douta(w_n15676_0[0]),.doutb(w_n15676_0[1]),.din(n15676));
	jspl jspl_w_n15678_0(.douta(w_n15678_0[0]),.doutb(w_n15678_0[1]),.din(n15678));
	jspl jspl_w_n15680_0(.douta(w_n15680_0[0]),.doutb(w_n15680_0[1]),.din(n15680));
	jspl jspl_w_n15683_0(.douta(w_n15683_0[0]),.doutb(w_n15683_0[1]),.din(n15683));
	jspl jspl_w_n15689_0(.douta(w_n15689_0[0]),.doutb(w_n15689_0[1]),.din(n15689));
	jspl jspl_w_n15691_0(.douta(w_n15691_0[0]),.doutb(w_n15691_0[1]),.din(n15691));
	jspl3 jspl3_w_n15692_0(.douta(w_n15692_0[0]),.doutb(w_n15692_0[1]),.doutc(w_n15692_0[2]),.din(n15692));
	jspl jspl_w_n15696_0(.douta(w_n15696_0[0]),.doutb(w_n15696_0[1]),.din(n15696));
	jspl jspl_w_n15697_0(.douta(w_n15697_0[0]),.doutb(w_n15697_0[1]),.din(n15697));
	jspl3 jspl3_w_n15698_0(.douta(w_n15698_0[0]),.doutb(w_n15698_0[1]),.doutc(w_n15698_0[2]),.din(n15698));
	jspl jspl_w_n15700_0(.douta(w_n15700_0[0]),.doutb(w_n15700_0[1]),.din(n15700));
	jspl jspl_w_n15705_0(.douta(w_n15705_0[0]),.doutb(w_n15705_0[1]),.din(n15705));
	jspl jspl_w_n15707_0(.douta(w_n15707_0[0]),.doutb(w_n15707_0[1]),.din(n15707));
	jspl jspl_w_n15708_0(.douta(w_n15708_0[0]),.doutb(w_n15708_0[1]),.din(n15708));
	jspl3 jspl3_w_n15709_0(.douta(w_n15709_0[0]),.doutb(w_n15709_0[1]),.doutc(w_n15709_0[2]),.din(n15709));
	jspl jspl_w_n15710_0(.douta(w_n15710_0[0]),.doutb(w_n15710_0[1]),.din(n15710));
	jspl jspl_w_n15714_0(.douta(w_n15714_0[0]),.doutb(w_n15714_0[1]),.din(n15714));
	jspl jspl_w_n15720_0(.douta(w_n15720_0[0]),.doutb(w_n15720_0[1]),.din(n15720));
	jspl jspl_w_n15721_0(.douta(w_n15721_0[0]),.doutb(w_n15721_0[1]),.din(n15721));
	jspl jspl_w_n15723_0(.douta(w_n15723_0[0]),.doutb(w_n15723_0[1]),.din(n15723));
	jspl jspl_w_n15725_0(.douta(w_n15725_0[0]),.doutb(w_n15725_0[1]),.din(n15725));
	jspl jspl_w_n15728_0(.douta(w_n15728_0[0]),.doutb(w_n15728_0[1]),.din(n15728));
	jspl jspl_w_n15734_0(.douta(w_n15734_0[0]),.doutb(w_n15734_0[1]),.din(n15734));
	jspl jspl_w_n15736_0(.douta(w_n15736_0[0]),.doutb(w_n15736_0[1]),.din(n15736));
	jspl3 jspl3_w_n15737_0(.douta(w_n15737_0[0]),.doutb(w_n15737_0[1]),.doutc(w_n15737_0[2]),.din(n15737));
	jspl jspl_w_n15741_0(.douta(w_n15741_0[0]),.doutb(w_n15741_0[1]),.din(n15741));
	jspl jspl_w_n15742_0(.douta(w_n15742_0[0]),.doutb(w_n15742_0[1]),.din(n15742));
	jspl3 jspl3_w_n15743_0(.douta(w_n15743_0[0]),.doutb(w_n15743_0[1]),.doutc(w_n15743_0[2]),.din(n15743));
	jspl jspl_w_n15745_0(.douta(w_n15745_0[0]),.doutb(w_n15745_0[1]),.din(n15745));
	jspl jspl_w_n15750_0(.douta(w_n15750_0[0]),.doutb(w_n15750_0[1]),.din(n15750));
	jspl jspl_w_n15752_0(.douta(w_n15752_0[0]),.doutb(w_n15752_0[1]),.din(n15752));
	jspl jspl_w_n15753_0(.douta(w_n15753_0[0]),.doutb(w_n15753_0[1]),.din(n15753));
	jspl3 jspl3_w_n15754_0(.douta(w_n15754_0[0]),.doutb(w_n15754_0[1]),.doutc(w_n15754_0[2]),.din(n15754));
	jspl jspl_w_n15755_0(.douta(w_n15755_0[0]),.doutb(w_n15755_0[1]),.din(n15755));
	jspl jspl_w_n15759_0(.douta(w_n15759_0[0]),.doutb(w_n15759_0[1]),.din(n15759));
	jspl jspl_w_n15765_0(.douta(w_n15765_0[0]),.doutb(w_n15765_0[1]),.din(n15765));
	jspl jspl_w_n15766_0(.douta(w_n15766_0[0]),.doutb(w_n15766_0[1]),.din(n15766));
	jspl jspl_w_n15768_0(.douta(w_n15768_0[0]),.doutb(w_n15768_0[1]),.din(n15768));
	jspl jspl_w_n15770_0(.douta(w_n15770_0[0]),.doutb(w_n15770_0[1]),.din(n15770));
	jspl jspl_w_n15773_0(.douta(w_n15773_0[0]),.doutb(w_n15773_0[1]),.din(n15773));
	jspl jspl_w_n15779_0(.douta(w_n15779_0[0]),.doutb(w_n15779_0[1]),.din(n15779));
	jspl jspl_w_n15781_0(.douta(w_n15781_0[0]),.doutb(w_n15781_0[1]),.din(n15781));
	jspl3 jspl3_w_n15782_0(.douta(w_n15782_0[0]),.doutb(w_n15782_0[1]),.doutc(w_n15782_0[2]),.din(n15782));
	jspl jspl_w_n15786_0(.douta(w_n15786_0[0]),.doutb(w_n15786_0[1]),.din(n15786));
	jspl jspl_w_n15787_0(.douta(w_n15787_0[0]),.doutb(w_n15787_0[1]),.din(n15787));
	jspl3 jspl3_w_n15788_0(.douta(w_n15788_0[0]),.doutb(w_n15788_0[1]),.doutc(w_n15788_0[2]),.din(n15788));
	jspl jspl_w_n15790_0(.douta(w_n15790_0[0]),.doutb(w_n15790_0[1]),.din(n15790));
	jspl jspl_w_n15795_0(.douta(w_n15795_0[0]),.doutb(w_n15795_0[1]),.din(n15795));
	jspl jspl_w_n15797_0(.douta(w_n15797_0[0]),.doutb(w_n15797_0[1]),.din(n15797));
	jspl jspl_w_n15798_0(.douta(w_n15798_0[0]),.doutb(w_n15798_0[1]),.din(n15798));
	jspl3 jspl3_w_n15799_0(.douta(w_n15799_0[0]),.doutb(w_n15799_0[1]),.doutc(w_n15799_0[2]),.din(n15799));
	jspl jspl_w_n15800_0(.douta(w_n15800_0[0]),.doutb(w_n15800_0[1]),.din(n15800));
	jspl jspl_w_n15804_0(.douta(w_n15804_0[0]),.doutb(w_n15804_0[1]),.din(n15804));
	jspl jspl_w_n15810_0(.douta(w_n15810_0[0]),.doutb(w_n15810_0[1]),.din(n15810));
	jspl jspl_w_n15811_0(.douta(w_n15811_0[0]),.doutb(w_n15811_0[1]),.din(n15811));
	jspl jspl_w_n15813_0(.douta(w_n15813_0[0]),.doutb(w_n15813_0[1]),.din(n15813));
	jspl jspl_w_n15818_0(.douta(w_n15818_0[0]),.doutb(w_n15818_0[1]),.din(n15818));
	jspl jspl_w_n15820_0(.douta(w_n15820_0[0]),.doutb(w_n15820_0[1]),.din(n15820));
	jspl jspl_w_n15821_0(.douta(w_n15821_0[0]),.doutb(w_n15821_0[1]),.din(n15821));
	jspl3 jspl3_w_n15822_0(.douta(w_n15822_0[0]),.doutb(w_n15822_0[1]),.doutc(w_n15822_0[2]),.din(n15822));
	jspl jspl_w_n15823_0(.douta(w_n15823_0[0]),.doutb(w_n15823_0[1]),.din(n15823));
	jspl jspl_w_n15825_0(.douta(w_n15825_0[0]),.doutb(w_n15825_0[1]),.din(n15825));
	jspl jspl_w_n15827_0(.douta(w_n15827_0[0]),.doutb(w_n15827_0[1]),.din(n15827));
	jspl jspl_w_n15829_0(.douta(w_n15829_0[0]),.doutb(w_n15829_0[1]),.din(n15829));
	jspl jspl_w_n15832_0(.douta(w_n15832_0[0]),.doutb(w_n15832_0[1]),.din(n15832));
	jspl jspl_w_n15838_0(.douta(w_n15838_0[0]),.doutb(w_n15838_0[1]),.din(n15838));
	jspl3 jspl3_w_n15840_0(.douta(w_n15840_0[0]),.doutb(w_n15840_0[1]),.doutc(w_n15840_0[2]),.din(n15840));
	jspl jspl_w_n15841_0(.douta(w_n15841_0[0]),.doutb(w_n15841_0[1]),.din(n15841));
	jspl jspl_w_n15845_0(.douta(w_n15845_0[0]),.doutb(w_n15845_0[1]),.din(n15845));
	jspl jspl_w_n15851_0(.douta(w_n15851_0[0]),.doutb(w_n15851_0[1]),.din(n15851));
	jspl jspl_w_n15852_0(.douta(w_n15852_0[0]),.doutb(w_n15852_0[1]),.din(n15852));
	jspl jspl_w_n15854_0(.douta(w_n15854_0[0]),.doutb(w_n15854_0[1]),.din(n15854));
	jspl jspl_w_n15856_0(.douta(w_n15856_0[0]),.doutb(w_n15856_0[1]),.din(n15856));
	jspl jspl_w_n15859_0(.douta(w_n15859_0[0]),.doutb(w_n15859_0[1]),.din(n15859));
	jspl jspl_w_n15865_0(.douta(w_n15865_0[0]),.doutb(w_n15865_0[1]),.din(n15865));
	jspl jspl_w_n15867_0(.douta(w_n15867_0[0]),.doutb(w_n15867_0[1]),.din(n15867));
	jspl3 jspl3_w_n15868_0(.douta(w_n15868_0[0]),.doutb(w_n15868_0[1]),.doutc(w_n15868_0[2]),.din(n15868));
	jspl jspl_w_n15872_0(.douta(w_n15872_0[0]),.doutb(w_n15872_0[1]),.din(n15872));
	jspl jspl_w_n15873_0(.douta(w_n15873_0[0]),.doutb(w_n15873_0[1]),.din(n15873));
	jspl3 jspl3_w_n15874_0(.douta(w_n15874_0[0]),.doutb(w_n15874_0[1]),.doutc(w_n15874_0[2]),.din(n15874));
	jspl jspl_w_n15876_0(.douta(w_n15876_0[0]),.doutb(w_n15876_0[1]),.din(n15876));
	jspl jspl_w_n15881_0(.douta(w_n15881_0[0]),.doutb(w_n15881_0[1]),.din(n15881));
	jspl jspl_w_n15883_0(.douta(w_n15883_0[0]),.doutb(w_n15883_0[1]),.din(n15883));
	jspl jspl_w_n15884_0(.douta(w_n15884_0[0]),.doutb(w_n15884_0[1]),.din(n15884));
	jspl3 jspl3_w_n15885_0(.douta(w_n15885_0[0]),.doutb(w_n15885_0[1]),.doutc(w_n15885_0[2]),.din(n15885));
	jspl jspl_w_n15886_0(.douta(w_n15886_0[0]),.doutb(w_n15886_0[1]),.din(n15886));
	jspl jspl_w_n15890_0(.douta(w_n15890_0[0]),.doutb(w_n15890_0[1]),.din(n15890));
	jspl jspl_w_n15896_0(.douta(w_n15896_0[0]),.doutb(w_n15896_0[1]),.din(n15896));
	jspl jspl_w_n15897_0(.douta(w_n15897_0[0]),.doutb(w_n15897_0[1]),.din(n15897));
	jspl jspl_w_n15899_0(.douta(w_n15899_0[0]),.doutb(w_n15899_0[1]),.din(n15899));
	jspl jspl_w_n15901_0(.douta(w_n15901_0[0]),.doutb(w_n15901_0[1]),.din(n15901));
	jspl jspl_w_n15904_0(.douta(w_n15904_0[0]),.doutb(w_n15904_0[1]),.din(n15904));
	jspl jspl_w_n15910_0(.douta(w_n15910_0[0]),.doutb(w_n15910_0[1]),.din(n15910));
	jspl jspl_w_n15912_0(.douta(w_n15912_0[0]),.doutb(w_n15912_0[1]),.din(n15912));
	jspl3 jspl3_w_n15913_0(.douta(w_n15913_0[0]),.doutb(w_n15913_0[1]),.doutc(w_n15913_0[2]),.din(n15913));
	jspl jspl_w_n15917_0(.douta(w_n15917_0[0]),.doutb(w_n15917_0[1]),.din(n15917));
	jspl jspl_w_n15918_0(.douta(w_n15918_0[0]),.doutb(w_n15918_0[1]),.din(n15918));
	jspl3 jspl3_w_n15919_0(.douta(w_n15919_0[0]),.doutb(w_n15919_0[1]),.doutc(w_n15919_0[2]),.din(n15919));
	jspl jspl_w_n15921_0(.douta(w_n15921_0[0]),.doutb(w_n15921_0[1]),.din(n15921));
	jspl jspl_w_n15926_0(.douta(w_n15926_0[0]),.doutb(w_n15926_0[1]),.din(n15926));
	jspl jspl_w_n15928_0(.douta(w_n15928_0[0]),.doutb(w_n15928_0[1]),.din(n15928));
	jspl jspl_w_n15929_0(.douta(w_n15929_0[0]),.doutb(w_n15929_0[1]),.din(n15929));
	jspl3 jspl3_w_n15930_0(.douta(w_n15930_0[0]),.doutb(w_n15930_0[1]),.doutc(w_n15930_0[2]),.din(n15930));
	jspl3 jspl3_w_n15930_1(.douta(w_n15930_1[0]),.doutb(w_n15930_1[1]),.doutc(w_n15930_1[2]),.din(w_n15930_0[0]));
	jspl jspl_w_n15933_0(.douta(w_n15933_0[0]),.doutb(w_n15933_0[1]),.din(n15933));
	jspl3 jspl3_w_n15934_0(.douta(w_n15934_0[0]),.doutb(w_n15934_0[1]),.doutc(w_n15934_0[2]),.din(n15934));
	jspl jspl_w_n15935_0(.douta(w_n15935_0[0]),.doutb(w_n15935_0[1]),.din(n15935));
	jspl jspl_w_n15936_0(.douta(w_n15936_0[0]),.doutb(w_n15936_0[1]),.din(n15936));
	jspl jspl_w_n15942_0(.douta(w_n15942_0[0]),.doutb(w_n15942_0[1]),.din(n15942));
	jspl3 jspl3_w_n15943_0(.douta(w_n15943_0[0]),.doutb(w_n15943_0[1]),.doutc(w_n15943_0[2]),.din(n15943));
	jspl jspl_w_n15944_0(.douta(w_n15944_0[0]),.doutb(w_n15944_0[1]),.din(n15944));
	jspl jspl_w_n15949_0(.douta(w_n15949_0[0]),.doutb(w_n15949_0[1]),.din(n15949));
	jspl3 jspl3_w_n15950_0(.douta(w_n15950_0[0]),.doutb(w_n15950_0[1]),.doutc(w_n15950_0[2]),.din(n15950));
	jspl3 jspl3_w_n15950_1(.douta(w_n15950_1[0]),.doutb(w_n15950_1[1]),.doutc(w_n15950_1[2]),.din(w_n15950_0[0]));
	jspl3 jspl3_w_n15950_2(.douta(w_n15950_2[0]),.doutb(w_n15950_2[1]),.doutc(w_n15950_2[2]),.din(w_n15950_0[1]));
	jspl3 jspl3_w_n15950_3(.douta(w_n15950_3[0]),.doutb(w_n15950_3[1]),.doutc(w_n15950_3[2]),.din(w_n15950_0[2]));
	jspl3 jspl3_w_n15950_4(.douta(w_n15950_4[0]),.doutb(w_n15950_4[1]),.doutc(w_n15950_4[2]),.din(w_n15950_1[0]));
	jspl3 jspl3_w_n15950_5(.douta(w_n15950_5[0]),.doutb(w_n15950_5[1]),.doutc(w_n15950_5[2]),.din(w_n15950_1[1]));
	jspl3 jspl3_w_n15950_6(.douta(w_n15950_6[0]),.doutb(w_n15950_6[1]),.doutc(w_n15950_6[2]),.din(w_n15950_1[2]));
	jspl3 jspl3_w_n15955_0(.douta(w_n15955_0[0]),.doutb(w_n15955_0[1]),.doutc(w_n15955_0[2]),.din(n15955));
	jspl3 jspl3_w_n15955_1(.douta(w_n15955_1[0]),.doutb(w_n15955_1[1]),.doutc(w_n15955_1[2]),.din(w_n15955_0[0]));
	jspl3 jspl3_w_n15955_2(.douta(w_n15955_2[0]),.doutb(w_n15955_2[1]),.doutc(w_n15955_2[2]),.din(w_n15955_0[1]));
	jspl3 jspl3_w_n15955_3(.douta(w_n15955_3[0]),.doutb(w_n15955_3[1]),.doutc(w_n15955_3[2]),.din(w_n15955_0[2]));
	jspl3 jspl3_w_n15955_4(.douta(w_n15955_4[0]),.doutb(w_n15955_4[1]),.doutc(w_n15955_4[2]),.din(w_n15955_1[0]));
	jspl3 jspl3_w_n15955_5(.douta(w_n15955_5[0]),.doutb(w_n15955_5[1]),.doutc(w_n15955_5[2]),.din(w_n15955_1[1]));
	jspl3 jspl3_w_n15955_6(.douta(w_n15955_6[0]),.doutb(w_n15955_6[1]),.doutc(w_n15955_6[2]),.din(w_n15955_1[2]));
	jspl3 jspl3_w_n15955_7(.douta(w_n15955_7[0]),.doutb(w_n15955_7[1]),.doutc(w_n15955_7[2]),.din(w_n15955_2[0]));
	jspl3 jspl3_w_n15955_8(.douta(w_n15955_8[0]),.doutb(w_n15955_8[1]),.doutc(w_n15955_8[2]),.din(w_n15955_2[1]));
	jspl3 jspl3_w_n15955_9(.douta(w_n15955_9[0]),.doutb(w_n15955_9[1]),.doutc(w_n15955_9[2]),.din(w_n15955_2[2]));
	jspl3 jspl3_w_n15955_10(.douta(w_n15955_10[0]),.doutb(w_n15955_10[1]),.doutc(w_n15955_10[2]),.din(w_n15955_3[0]));
	jspl3 jspl3_w_n15955_11(.douta(w_n15955_11[0]),.doutb(w_n15955_11[1]),.doutc(w_n15955_11[2]),.din(w_n15955_3[1]));
	jspl3 jspl3_w_n15955_12(.douta(w_n15955_12[0]),.doutb(w_n15955_12[1]),.doutc(w_n15955_12[2]),.din(w_n15955_3[2]));
	jspl3 jspl3_w_n15955_13(.douta(w_n15955_13[0]),.doutb(w_n15955_13[1]),.doutc(w_n15955_13[2]),.din(w_n15955_4[0]));
	jspl3 jspl3_w_n15955_14(.douta(w_n15955_14[0]),.doutb(w_n15955_14[1]),.doutc(w_n15955_14[2]),.din(w_n15955_4[1]));
	jspl3 jspl3_w_n15955_15(.douta(w_n15955_15[0]),.doutb(w_n15955_15[1]),.doutc(w_n15955_15[2]),.din(w_n15955_4[2]));
	jspl3 jspl3_w_n15955_16(.douta(w_n15955_16[0]),.doutb(w_n15955_16[1]),.doutc(w_n15955_16[2]),.din(w_n15955_5[0]));
	jspl3 jspl3_w_n15955_17(.douta(w_n15955_17[0]),.doutb(w_n15955_17[1]),.doutc(w_n15955_17[2]),.din(w_n15955_5[1]));
	jspl3 jspl3_w_n15955_18(.douta(w_n15955_18[0]),.doutb(w_n15955_18[1]),.doutc(w_n15955_18[2]),.din(w_n15955_5[2]));
	jspl3 jspl3_w_n15955_19(.douta(w_n15955_19[0]),.doutb(w_n15955_19[1]),.doutc(w_n15955_19[2]),.din(w_n15955_6[0]));
	jspl3 jspl3_w_n15955_20(.douta(w_n15955_20[0]),.doutb(w_n15955_20[1]),.doutc(w_n15955_20[2]),.din(w_n15955_6[1]));
	jspl jspl_w_n15955_21(.douta(w_n15955_21[0]),.doutb(w_n15955_21[1]),.din(w_n15955_6[2]));
	jspl jspl_w_n15959_0(.douta(w_n15959_0[0]),.doutb(w_n15959_0[1]),.din(n15959));
	jspl3 jspl3_w_n15961_0(.douta(w_n15961_0[0]),.doutb(w_n15961_0[1]),.doutc(w_n15961_0[2]),.din(n15961));
	jspl jspl_w_n15961_1(.douta(w_n15961_1[0]),.doutb(w_n15961_1[1]),.din(w_n15961_0[0]));
	jspl3 jspl3_w_n15962_0(.douta(w_n15962_0[0]),.doutb(w_n15962_0[1]),.doutc(w_n15962_0[2]),.din(n15962));
	jspl3 jspl3_w_n15966_0(.douta(w_n15966_0[0]),.doutb(w_n15966_0[1]),.doutc(w_n15966_0[2]),.din(n15966));
	jspl jspl_w_n15967_0(.douta(w_n15967_0[0]),.doutb(w_n15967_0[1]),.din(n15967));
	jspl jspl_w_n15968_0(.douta(w_n15968_0[0]),.doutb(w_n15968_0[1]),.din(n15968));
	jspl jspl_w_n15969_0(.douta(w_n15969_0[0]),.doutb(w_n15969_0[1]),.din(n15969));
	jspl jspl_w_n15971_0(.douta(w_n15971_0[0]),.doutb(w_n15971_0[1]),.din(n15971));
	jspl jspl_w_n15973_0(.douta(w_n15973_0[0]),.doutb(w_n15973_0[1]),.din(n15973));
	jspl jspl_w_n15975_0(.douta(w_n15975_0[0]),.doutb(w_n15975_0[1]),.din(n15975));
	jspl jspl_w_n15978_0(.douta(w_n15978_0[0]),.doutb(w_n15978_0[1]),.din(n15978));
	jspl jspl_w_n15983_0(.douta(w_n15983_0[0]),.doutb(w_n15983_0[1]),.din(n15983));
	jspl3 jspl3_w_n15985_0(.douta(w_n15985_0[0]),.doutb(w_n15985_0[1]),.doutc(w_n15985_0[2]),.din(n15985));
	jspl jspl_w_n15986_0(.douta(w_n15986_0[0]),.doutb(w_n15986_0[1]),.din(n15986));
	jspl jspl_w_n15990_0(.douta(w_n15990_0[0]),.doutb(w_n15990_0[1]),.din(n15990));
	jspl jspl_w_n15991_0(.douta(w_n15991_0[0]),.doutb(w_n15991_0[1]),.din(n15991));
	jspl jspl_w_n15993_0(.douta(w_n15993_0[0]),.doutb(w_n15993_0[1]),.din(n15993));
	jspl jspl_w_n15997_0(.douta(w_n15997_0[0]),.doutb(w_n15997_0[1]),.din(n15997));
	jspl jspl_w_n15999_0(.douta(w_n15999_0[0]),.doutb(w_n15999_0[1]),.din(n15999));
	jspl jspl_w_n16000_0(.douta(w_n16000_0[0]),.doutb(w_n16000_0[1]),.din(n16000));
	jspl3 jspl3_w_n16001_0(.douta(w_n16001_0[0]),.doutb(w_n16001_0[1]),.doutc(w_n16001_0[2]),.din(n16001));
	jspl jspl_w_n16002_0(.douta(w_n16002_0[0]),.doutb(w_n16002_0[1]),.din(n16002));
	jspl jspl_w_n16006_0(.douta(w_n16006_0[0]),.doutb(w_n16006_0[1]),.din(n16006));
	jspl jspl_w_n16008_0(.douta(w_n16008_0[0]),.doutb(w_n16008_0[1]),.din(n16008));
	jspl jspl_w_n16010_0(.douta(w_n16010_0[0]),.doutb(w_n16010_0[1]),.din(n16010));
	jspl jspl_w_n16012_0(.douta(w_n16012_0[0]),.doutb(w_n16012_0[1]),.din(n16012));
	jspl jspl_w_n16015_0(.douta(w_n16015_0[0]),.doutb(w_n16015_0[1]),.din(n16015));
	jspl jspl_w_n16021_0(.douta(w_n16021_0[0]),.doutb(w_n16021_0[1]),.din(n16021));
	jspl3 jspl3_w_n16023_0(.douta(w_n16023_0[0]),.doutb(w_n16023_0[1]),.doutc(w_n16023_0[2]),.din(n16023));
	jspl jspl_w_n16024_0(.douta(w_n16024_0[0]),.doutb(w_n16024_0[1]),.din(n16024));
	jspl jspl_w_n16029_0(.douta(w_n16029_0[0]),.doutb(w_n16029_0[1]),.din(n16029));
	jspl jspl_w_n16031_0(.douta(w_n16031_0[0]),.doutb(w_n16031_0[1]),.din(n16031));
	jspl jspl_w_n16033_0(.douta(w_n16033_0[0]),.doutb(w_n16033_0[1]),.din(n16033));
	jspl jspl_w_n16037_0(.douta(w_n16037_0[0]),.doutb(w_n16037_0[1]),.din(n16037));
	jspl jspl_w_n16039_0(.douta(w_n16039_0[0]),.doutb(w_n16039_0[1]),.din(n16039));
	jspl jspl_w_n16040_0(.douta(w_n16040_0[0]),.doutb(w_n16040_0[1]),.din(n16040));
	jspl3 jspl3_w_n16041_0(.douta(w_n16041_0[0]),.doutb(w_n16041_0[1]),.doutc(w_n16041_0[2]),.din(n16041));
	jspl jspl_w_n16042_0(.douta(w_n16042_0[0]),.doutb(w_n16042_0[1]),.din(n16042));
	jspl jspl_w_n16048_0(.douta(w_n16048_0[0]),.doutb(w_n16048_0[1]),.din(n16048));
	jspl jspl_w_n16049_0(.douta(w_n16049_0[0]),.doutb(w_n16049_0[1]),.din(n16049));
	jspl jspl_w_n16051_0(.douta(w_n16051_0[0]),.doutb(w_n16051_0[1]),.din(n16051));
	jspl jspl_w_n16053_0(.douta(w_n16053_0[0]),.doutb(w_n16053_0[1]),.din(n16053));
	jspl jspl_w_n16055_0(.douta(w_n16055_0[0]),.doutb(w_n16055_0[1]),.din(n16055));
	jspl jspl_w_n16061_0(.douta(w_n16061_0[0]),.doutb(w_n16061_0[1]),.din(n16061));
	jspl jspl_w_n16063_0(.douta(w_n16063_0[0]),.doutb(w_n16063_0[1]),.din(n16063));
	jspl3 jspl3_w_n16064_0(.douta(w_n16064_0[0]),.doutb(w_n16064_0[1]),.doutc(w_n16064_0[2]),.din(n16064));
	jspl jspl_w_n16067_0(.douta(w_n16067_0[0]),.doutb(w_n16067_0[1]),.din(n16067));
	jspl jspl_w_n16068_0(.douta(w_n16068_0[0]),.doutb(w_n16068_0[1]),.din(n16068));
	jspl3 jspl3_w_n16069_0(.douta(w_n16069_0[0]),.doutb(w_n16069_0[1]),.doutc(w_n16069_0[2]),.din(n16069));
	jspl jspl_w_n16071_0(.douta(w_n16071_0[0]),.doutb(w_n16071_0[1]),.din(n16071));
	jspl jspl_w_n16075_0(.douta(w_n16075_0[0]),.doutb(w_n16075_0[1]),.din(n16075));
	jspl jspl_w_n16077_0(.douta(w_n16077_0[0]),.doutb(w_n16077_0[1]),.din(n16077));
	jspl jspl_w_n16078_0(.douta(w_n16078_0[0]),.doutb(w_n16078_0[1]),.din(n16078));
	jspl3 jspl3_w_n16079_0(.douta(w_n16079_0[0]),.doutb(w_n16079_0[1]),.doutc(w_n16079_0[2]),.din(n16079));
	jspl jspl_w_n16080_0(.douta(w_n16080_0[0]),.doutb(w_n16080_0[1]),.din(n16080));
	jspl jspl_w_n16083_0(.douta(w_n16083_0[0]),.doutb(w_n16083_0[1]),.din(n16083));
	jspl jspl_w_n16089_0(.douta(w_n16089_0[0]),.doutb(w_n16089_0[1]),.din(n16089));
	jspl jspl_w_n16090_0(.douta(w_n16090_0[0]),.doutb(w_n16090_0[1]),.din(n16090));
	jspl jspl_w_n16092_0(.douta(w_n16092_0[0]),.doutb(w_n16092_0[1]),.din(n16092));
	jspl jspl_w_n16094_0(.douta(w_n16094_0[0]),.doutb(w_n16094_0[1]),.din(n16094));
	jspl jspl_w_n16096_0(.douta(w_n16096_0[0]),.doutb(w_n16096_0[1]),.din(n16096));
	jspl jspl_w_n16102_0(.douta(w_n16102_0[0]),.doutb(w_n16102_0[1]),.din(n16102));
	jspl jspl_w_n16104_0(.douta(w_n16104_0[0]),.doutb(w_n16104_0[1]),.din(n16104));
	jspl3 jspl3_w_n16105_0(.douta(w_n16105_0[0]),.doutb(w_n16105_0[1]),.doutc(w_n16105_0[2]),.din(n16105));
	jspl jspl_w_n16108_0(.douta(w_n16108_0[0]),.doutb(w_n16108_0[1]),.din(n16108));
	jspl jspl_w_n16109_0(.douta(w_n16109_0[0]),.doutb(w_n16109_0[1]),.din(n16109));
	jspl3 jspl3_w_n16110_0(.douta(w_n16110_0[0]),.doutb(w_n16110_0[1]),.doutc(w_n16110_0[2]),.din(n16110));
	jspl jspl_w_n16112_0(.douta(w_n16112_0[0]),.doutb(w_n16112_0[1]),.din(n16112));
	jspl jspl_w_n16116_0(.douta(w_n16116_0[0]),.doutb(w_n16116_0[1]),.din(n16116));
	jspl jspl_w_n16118_0(.douta(w_n16118_0[0]),.doutb(w_n16118_0[1]),.din(n16118));
	jspl jspl_w_n16119_0(.douta(w_n16119_0[0]),.doutb(w_n16119_0[1]),.din(n16119));
	jspl3 jspl3_w_n16120_0(.douta(w_n16120_0[0]),.doutb(w_n16120_0[1]),.doutc(w_n16120_0[2]),.din(n16120));
	jspl jspl_w_n16121_0(.douta(w_n16121_0[0]),.doutb(w_n16121_0[1]),.din(n16121));
	jspl jspl_w_n16124_0(.douta(w_n16124_0[0]),.doutb(w_n16124_0[1]),.din(n16124));
	jspl jspl_w_n16130_0(.douta(w_n16130_0[0]),.doutb(w_n16130_0[1]),.din(n16130));
	jspl jspl_w_n16131_0(.douta(w_n16131_0[0]),.doutb(w_n16131_0[1]),.din(n16131));
	jspl jspl_w_n16133_0(.douta(w_n16133_0[0]),.doutb(w_n16133_0[1]),.din(n16133));
	jspl jspl_w_n16135_0(.douta(w_n16135_0[0]),.doutb(w_n16135_0[1]),.din(n16135));
	jspl jspl_w_n16137_0(.douta(w_n16137_0[0]),.doutb(w_n16137_0[1]),.din(n16137));
	jspl jspl_w_n16143_0(.douta(w_n16143_0[0]),.doutb(w_n16143_0[1]),.din(n16143));
	jspl jspl_w_n16145_0(.douta(w_n16145_0[0]),.doutb(w_n16145_0[1]),.din(n16145));
	jspl3 jspl3_w_n16146_0(.douta(w_n16146_0[0]),.doutb(w_n16146_0[1]),.doutc(w_n16146_0[2]),.din(n16146));
	jspl jspl_w_n16149_0(.douta(w_n16149_0[0]),.doutb(w_n16149_0[1]),.din(n16149));
	jspl jspl_w_n16150_0(.douta(w_n16150_0[0]),.doutb(w_n16150_0[1]),.din(n16150));
	jspl3 jspl3_w_n16151_0(.douta(w_n16151_0[0]),.doutb(w_n16151_0[1]),.doutc(w_n16151_0[2]),.din(n16151));
	jspl jspl_w_n16153_0(.douta(w_n16153_0[0]),.doutb(w_n16153_0[1]),.din(n16153));
	jspl jspl_w_n16157_0(.douta(w_n16157_0[0]),.doutb(w_n16157_0[1]),.din(n16157));
	jspl jspl_w_n16159_0(.douta(w_n16159_0[0]),.doutb(w_n16159_0[1]),.din(n16159));
	jspl jspl_w_n16160_0(.douta(w_n16160_0[0]),.doutb(w_n16160_0[1]),.din(n16160));
	jspl3 jspl3_w_n16161_0(.douta(w_n16161_0[0]),.doutb(w_n16161_0[1]),.doutc(w_n16161_0[2]),.din(n16161));
	jspl jspl_w_n16162_0(.douta(w_n16162_0[0]),.doutb(w_n16162_0[1]),.din(n16162));
	jspl jspl_w_n16165_0(.douta(w_n16165_0[0]),.doutb(w_n16165_0[1]),.din(n16165));
	jspl jspl_w_n16171_0(.douta(w_n16171_0[0]),.doutb(w_n16171_0[1]),.din(n16171));
	jspl jspl_w_n16172_0(.douta(w_n16172_0[0]),.doutb(w_n16172_0[1]),.din(n16172));
	jspl jspl_w_n16174_0(.douta(w_n16174_0[0]),.doutb(w_n16174_0[1]),.din(n16174));
	jspl jspl_w_n16176_0(.douta(w_n16176_0[0]),.doutb(w_n16176_0[1]),.din(n16176));
	jspl jspl_w_n16178_0(.douta(w_n16178_0[0]),.doutb(w_n16178_0[1]),.din(n16178));
	jspl jspl_w_n16184_0(.douta(w_n16184_0[0]),.doutb(w_n16184_0[1]),.din(n16184));
	jspl jspl_w_n16186_0(.douta(w_n16186_0[0]),.doutb(w_n16186_0[1]),.din(n16186));
	jspl3 jspl3_w_n16187_0(.douta(w_n16187_0[0]),.doutb(w_n16187_0[1]),.doutc(w_n16187_0[2]),.din(n16187));
	jspl jspl_w_n16190_0(.douta(w_n16190_0[0]),.doutb(w_n16190_0[1]),.din(n16190));
	jspl jspl_w_n16191_0(.douta(w_n16191_0[0]),.doutb(w_n16191_0[1]),.din(n16191));
	jspl3 jspl3_w_n16192_0(.douta(w_n16192_0[0]),.doutb(w_n16192_0[1]),.doutc(w_n16192_0[2]),.din(n16192));
	jspl jspl_w_n16194_0(.douta(w_n16194_0[0]),.doutb(w_n16194_0[1]),.din(n16194));
	jspl jspl_w_n16198_0(.douta(w_n16198_0[0]),.doutb(w_n16198_0[1]),.din(n16198));
	jspl jspl_w_n16200_0(.douta(w_n16200_0[0]),.doutb(w_n16200_0[1]),.din(n16200));
	jspl jspl_w_n16201_0(.douta(w_n16201_0[0]),.doutb(w_n16201_0[1]),.din(n16201));
	jspl3 jspl3_w_n16202_0(.douta(w_n16202_0[0]),.doutb(w_n16202_0[1]),.doutc(w_n16202_0[2]),.din(n16202));
	jspl jspl_w_n16203_0(.douta(w_n16203_0[0]),.doutb(w_n16203_0[1]),.din(n16203));
	jspl jspl_w_n16206_0(.douta(w_n16206_0[0]),.doutb(w_n16206_0[1]),.din(n16206));
	jspl jspl_w_n16212_0(.douta(w_n16212_0[0]),.doutb(w_n16212_0[1]),.din(n16212));
	jspl jspl_w_n16213_0(.douta(w_n16213_0[0]),.doutb(w_n16213_0[1]),.din(n16213));
	jspl jspl_w_n16215_0(.douta(w_n16215_0[0]),.doutb(w_n16215_0[1]),.din(n16215));
	jspl jspl_w_n16217_0(.douta(w_n16217_0[0]),.doutb(w_n16217_0[1]),.din(n16217));
	jspl jspl_w_n16219_0(.douta(w_n16219_0[0]),.doutb(w_n16219_0[1]),.din(n16219));
	jspl jspl_w_n16225_0(.douta(w_n16225_0[0]),.doutb(w_n16225_0[1]),.din(n16225));
	jspl jspl_w_n16227_0(.douta(w_n16227_0[0]),.doutb(w_n16227_0[1]),.din(n16227));
	jspl3 jspl3_w_n16228_0(.douta(w_n16228_0[0]),.doutb(w_n16228_0[1]),.doutc(w_n16228_0[2]),.din(n16228));
	jspl jspl_w_n16231_0(.douta(w_n16231_0[0]),.doutb(w_n16231_0[1]),.din(n16231));
	jspl jspl_w_n16232_0(.douta(w_n16232_0[0]),.doutb(w_n16232_0[1]),.din(n16232));
	jspl3 jspl3_w_n16233_0(.douta(w_n16233_0[0]),.doutb(w_n16233_0[1]),.doutc(w_n16233_0[2]),.din(n16233));
	jspl jspl_w_n16235_0(.douta(w_n16235_0[0]),.doutb(w_n16235_0[1]),.din(n16235));
	jspl jspl_w_n16239_0(.douta(w_n16239_0[0]),.doutb(w_n16239_0[1]),.din(n16239));
	jspl jspl_w_n16241_0(.douta(w_n16241_0[0]),.doutb(w_n16241_0[1]),.din(n16241));
	jspl jspl_w_n16242_0(.douta(w_n16242_0[0]),.doutb(w_n16242_0[1]),.din(n16242));
	jspl3 jspl3_w_n16243_0(.douta(w_n16243_0[0]),.doutb(w_n16243_0[1]),.doutc(w_n16243_0[2]),.din(n16243));
	jspl jspl_w_n16244_0(.douta(w_n16244_0[0]),.doutb(w_n16244_0[1]),.din(n16244));
	jspl jspl_w_n16247_0(.douta(w_n16247_0[0]),.doutb(w_n16247_0[1]),.din(n16247));
	jspl jspl_w_n16253_0(.douta(w_n16253_0[0]),.doutb(w_n16253_0[1]),.din(n16253));
	jspl jspl_w_n16254_0(.douta(w_n16254_0[0]),.doutb(w_n16254_0[1]),.din(n16254));
	jspl jspl_w_n16256_0(.douta(w_n16256_0[0]),.doutb(w_n16256_0[1]),.din(n16256));
	jspl jspl_w_n16258_0(.douta(w_n16258_0[0]),.doutb(w_n16258_0[1]),.din(n16258));
	jspl jspl_w_n16260_0(.douta(w_n16260_0[0]),.doutb(w_n16260_0[1]),.din(n16260));
	jspl jspl_w_n16266_0(.douta(w_n16266_0[0]),.doutb(w_n16266_0[1]),.din(n16266));
	jspl jspl_w_n16268_0(.douta(w_n16268_0[0]),.doutb(w_n16268_0[1]),.din(n16268));
	jspl3 jspl3_w_n16269_0(.douta(w_n16269_0[0]),.doutb(w_n16269_0[1]),.doutc(w_n16269_0[2]),.din(n16269));
	jspl jspl_w_n16272_0(.douta(w_n16272_0[0]),.doutb(w_n16272_0[1]),.din(n16272));
	jspl jspl_w_n16273_0(.douta(w_n16273_0[0]),.doutb(w_n16273_0[1]),.din(n16273));
	jspl3 jspl3_w_n16274_0(.douta(w_n16274_0[0]),.doutb(w_n16274_0[1]),.doutc(w_n16274_0[2]),.din(n16274));
	jspl jspl_w_n16276_0(.douta(w_n16276_0[0]),.doutb(w_n16276_0[1]),.din(n16276));
	jspl jspl_w_n16280_0(.douta(w_n16280_0[0]),.doutb(w_n16280_0[1]),.din(n16280));
	jspl jspl_w_n16282_0(.douta(w_n16282_0[0]),.doutb(w_n16282_0[1]),.din(n16282));
	jspl jspl_w_n16283_0(.douta(w_n16283_0[0]),.doutb(w_n16283_0[1]),.din(n16283));
	jspl3 jspl3_w_n16284_0(.douta(w_n16284_0[0]),.doutb(w_n16284_0[1]),.doutc(w_n16284_0[2]),.din(n16284));
	jspl jspl_w_n16285_0(.douta(w_n16285_0[0]),.doutb(w_n16285_0[1]),.din(n16285));
	jspl jspl_w_n16288_0(.douta(w_n16288_0[0]),.doutb(w_n16288_0[1]),.din(n16288));
	jspl jspl_w_n16294_0(.douta(w_n16294_0[0]),.doutb(w_n16294_0[1]),.din(n16294));
	jspl jspl_w_n16295_0(.douta(w_n16295_0[0]),.doutb(w_n16295_0[1]),.din(n16295));
	jspl jspl_w_n16297_0(.douta(w_n16297_0[0]),.doutb(w_n16297_0[1]),.din(n16297));
	jspl jspl_w_n16299_0(.douta(w_n16299_0[0]),.doutb(w_n16299_0[1]),.din(n16299));
	jspl jspl_w_n16301_0(.douta(w_n16301_0[0]),.doutb(w_n16301_0[1]),.din(n16301));
	jspl jspl_w_n16307_0(.douta(w_n16307_0[0]),.doutb(w_n16307_0[1]),.din(n16307));
	jspl jspl_w_n16309_0(.douta(w_n16309_0[0]),.doutb(w_n16309_0[1]),.din(n16309));
	jspl3 jspl3_w_n16310_0(.douta(w_n16310_0[0]),.doutb(w_n16310_0[1]),.doutc(w_n16310_0[2]),.din(n16310));
	jspl jspl_w_n16313_0(.douta(w_n16313_0[0]),.doutb(w_n16313_0[1]),.din(n16313));
	jspl jspl_w_n16314_0(.douta(w_n16314_0[0]),.doutb(w_n16314_0[1]),.din(n16314));
	jspl3 jspl3_w_n16315_0(.douta(w_n16315_0[0]),.doutb(w_n16315_0[1]),.doutc(w_n16315_0[2]),.din(n16315));
	jspl jspl_w_n16317_0(.douta(w_n16317_0[0]),.doutb(w_n16317_0[1]),.din(n16317));
	jspl jspl_w_n16321_0(.douta(w_n16321_0[0]),.doutb(w_n16321_0[1]),.din(n16321));
	jspl jspl_w_n16323_0(.douta(w_n16323_0[0]),.doutb(w_n16323_0[1]),.din(n16323));
	jspl jspl_w_n16324_0(.douta(w_n16324_0[0]),.doutb(w_n16324_0[1]),.din(n16324));
	jspl3 jspl3_w_n16325_0(.douta(w_n16325_0[0]),.doutb(w_n16325_0[1]),.doutc(w_n16325_0[2]),.din(n16325));
	jspl jspl_w_n16326_0(.douta(w_n16326_0[0]),.doutb(w_n16326_0[1]),.din(n16326));
	jspl jspl_w_n16329_0(.douta(w_n16329_0[0]),.doutb(w_n16329_0[1]),.din(n16329));
	jspl jspl_w_n16335_0(.douta(w_n16335_0[0]),.doutb(w_n16335_0[1]),.din(n16335));
	jspl jspl_w_n16336_0(.douta(w_n16336_0[0]),.doutb(w_n16336_0[1]),.din(n16336));
	jspl jspl_w_n16338_0(.douta(w_n16338_0[0]),.doutb(w_n16338_0[1]),.din(n16338));
	jspl jspl_w_n16340_0(.douta(w_n16340_0[0]),.doutb(w_n16340_0[1]),.din(n16340));
	jspl jspl_w_n16342_0(.douta(w_n16342_0[0]),.doutb(w_n16342_0[1]),.din(n16342));
	jspl jspl_w_n16348_0(.douta(w_n16348_0[0]),.doutb(w_n16348_0[1]),.din(n16348));
	jspl jspl_w_n16350_0(.douta(w_n16350_0[0]),.doutb(w_n16350_0[1]),.din(n16350));
	jspl3 jspl3_w_n16351_0(.douta(w_n16351_0[0]),.doutb(w_n16351_0[1]),.doutc(w_n16351_0[2]),.din(n16351));
	jspl jspl_w_n16354_0(.douta(w_n16354_0[0]),.doutb(w_n16354_0[1]),.din(n16354));
	jspl jspl_w_n16355_0(.douta(w_n16355_0[0]),.doutb(w_n16355_0[1]),.din(n16355));
	jspl3 jspl3_w_n16356_0(.douta(w_n16356_0[0]),.doutb(w_n16356_0[1]),.doutc(w_n16356_0[2]),.din(n16356));
	jspl jspl_w_n16358_0(.douta(w_n16358_0[0]),.doutb(w_n16358_0[1]),.din(n16358));
	jspl jspl_w_n16362_0(.douta(w_n16362_0[0]),.doutb(w_n16362_0[1]),.din(n16362));
	jspl jspl_w_n16364_0(.douta(w_n16364_0[0]),.doutb(w_n16364_0[1]),.din(n16364));
	jspl jspl_w_n16365_0(.douta(w_n16365_0[0]),.doutb(w_n16365_0[1]),.din(n16365));
	jspl3 jspl3_w_n16366_0(.douta(w_n16366_0[0]),.doutb(w_n16366_0[1]),.doutc(w_n16366_0[2]),.din(n16366));
	jspl jspl_w_n16367_0(.douta(w_n16367_0[0]),.doutb(w_n16367_0[1]),.din(n16367));
	jspl jspl_w_n16370_0(.douta(w_n16370_0[0]),.doutb(w_n16370_0[1]),.din(n16370));
	jspl jspl_w_n16376_0(.douta(w_n16376_0[0]),.doutb(w_n16376_0[1]),.din(n16376));
	jspl jspl_w_n16377_0(.douta(w_n16377_0[0]),.doutb(w_n16377_0[1]),.din(n16377));
	jspl jspl_w_n16379_0(.douta(w_n16379_0[0]),.doutb(w_n16379_0[1]),.din(n16379));
	jspl jspl_w_n16381_0(.douta(w_n16381_0[0]),.doutb(w_n16381_0[1]),.din(n16381));
	jspl jspl_w_n16383_0(.douta(w_n16383_0[0]),.doutb(w_n16383_0[1]),.din(n16383));
	jspl jspl_w_n16389_0(.douta(w_n16389_0[0]),.doutb(w_n16389_0[1]),.din(n16389));
	jspl jspl_w_n16391_0(.douta(w_n16391_0[0]),.doutb(w_n16391_0[1]),.din(n16391));
	jspl3 jspl3_w_n16392_0(.douta(w_n16392_0[0]),.doutb(w_n16392_0[1]),.doutc(w_n16392_0[2]),.din(n16392));
	jspl jspl_w_n16395_0(.douta(w_n16395_0[0]),.doutb(w_n16395_0[1]),.din(n16395));
	jspl jspl_w_n16396_0(.douta(w_n16396_0[0]),.doutb(w_n16396_0[1]),.din(n16396));
	jspl3 jspl3_w_n16397_0(.douta(w_n16397_0[0]),.doutb(w_n16397_0[1]),.doutc(w_n16397_0[2]),.din(n16397));
	jspl jspl_w_n16399_0(.douta(w_n16399_0[0]),.doutb(w_n16399_0[1]),.din(n16399));
	jspl jspl_w_n16401_0(.douta(w_n16401_0[0]),.doutb(w_n16401_0[1]),.din(n16401));
	jspl jspl_w_n16403_0(.douta(w_n16403_0[0]),.doutb(w_n16403_0[1]),.din(n16403));
	jspl jspl_w_n16409_0(.douta(w_n16409_0[0]),.doutb(w_n16409_0[1]),.din(n16409));
	jspl3 jspl3_w_n16411_0(.douta(w_n16411_0[0]),.doutb(w_n16411_0[1]),.doutc(w_n16411_0[2]),.din(n16411));
	jspl jspl_w_n16412_0(.douta(w_n16412_0[0]),.doutb(w_n16412_0[1]),.din(n16412));
	jspl jspl_w_n16414_0(.douta(w_n16414_0[0]),.doutb(w_n16414_0[1]),.din(n16414));
	jspl jspl_w_n16416_0(.douta(w_n16416_0[0]),.doutb(w_n16416_0[1]),.din(n16416));
	jspl jspl_w_n16420_0(.douta(w_n16420_0[0]),.doutb(w_n16420_0[1]),.din(n16420));
	jspl jspl_w_n16422_0(.douta(w_n16422_0[0]),.doutb(w_n16422_0[1]),.din(n16422));
	jspl jspl_w_n16423_0(.douta(w_n16423_0[0]),.doutb(w_n16423_0[1]),.din(n16423));
	jspl jspl_w_n16424_0(.douta(w_n16424_0[0]),.doutb(w_n16424_0[1]),.din(n16424));
	jspl3 jspl3_w_n16425_0(.douta(w_n16425_0[0]),.doutb(w_n16425_0[1]),.doutc(w_n16425_0[2]),.din(n16425));
	jspl jspl_w_n16428_0(.douta(w_n16428_0[0]),.doutb(w_n16428_0[1]),.din(n16428));
	jspl jspl_w_n16429_0(.douta(w_n16429_0[0]),.doutb(w_n16429_0[1]),.din(n16429));
	jspl3 jspl3_w_n16430_0(.douta(w_n16430_0[0]),.doutb(w_n16430_0[1]),.doutc(w_n16430_0[2]),.din(n16430));
	jspl jspl_w_n16432_0(.douta(w_n16432_0[0]),.doutb(w_n16432_0[1]),.din(n16432));
	jspl jspl_w_n16436_0(.douta(w_n16436_0[0]),.doutb(w_n16436_0[1]),.din(n16436));
	jspl jspl_w_n16438_0(.douta(w_n16438_0[0]),.doutb(w_n16438_0[1]),.din(n16438));
	jspl jspl_w_n16439_0(.douta(w_n16439_0[0]),.doutb(w_n16439_0[1]),.din(n16439));
	jspl3 jspl3_w_n16440_0(.douta(w_n16440_0[0]),.doutb(w_n16440_0[1]),.doutc(w_n16440_0[2]),.din(n16440));
	jspl jspl_w_n16441_0(.douta(w_n16441_0[0]),.doutb(w_n16441_0[1]),.din(n16441));
	jspl jspl_w_n16444_0(.douta(w_n16444_0[0]),.doutb(w_n16444_0[1]),.din(n16444));
	jspl jspl_w_n16450_0(.douta(w_n16450_0[0]),.doutb(w_n16450_0[1]),.din(n16450));
	jspl jspl_w_n16451_0(.douta(w_n16451_0[0]),.doutb(w_n16451_0[1]),.din(n16451));
	jspl jspl_w_n16453_0(.douta(w_n16453_0[0]),.doutb(w_n16453_0[1]),.din(n16453));
	jspl jspl_w_n16455_0(.douta(w_n16455_0[0]),.doutb(w_n16455_0[1]),.din(n16455));
	jspl jspl_w_n16457_0(.douta(w_n16457_0[0]),.doutb(w_n16457_0[1]),.din(n16457));
	jspl jspl_w_n16463_0(.douta(w_n16463_0[0]),.doutb(w_n16463_0[1]),.din(n16463));
	jspl jspl_w_n16465_0(.douta(w_n16465_0[0]),.doutb(w_n16465_0[1]),.din(n16465));
	jspl3 jspl3_w_n16466_0(.douta(w_n16466_0[0]),.doutb(w_n16466_0[1]),.doutc(w_n16466_0[2]),.din(n16466));
	jspl jspl_w_n16469_0(.douta(w_n16469_0[0]),.doutb(w_n16469_0[1]),.din(n16469));
	jspl jspl_w_n16470_0(.douta(w_n16470_0[0]),.doutb(w_n16470_0[1]),.din(n16470));
	jspl3 jspl3_w_n16471_0(.douta(w_n16471_0[0]),.doutb(w_n16471_0[1]),.doutc(w_n16471_0[2]),.din(n16471));
	jspl jspl_w_n16473_0(.douta(w_n16473_0[0]),.doutb(w_n16473_0[1]),.din(n16473));
	jspl jspl_w_n16477_0(.douta(w_n16477_0[0]),.doutb(w_n16477_0[1]),.din(n16477));
	jspl jspl_w_n16479_0(.douta(w_n16479_0[0]),.doutb(w_n16479_0[1]),.din(n16479));
	jspl jspl_w_n16480_0(.douta(w_n16480_0[0]),.doutb(w_n16480_0[1]),.din(n16480));
	jspl3 jspl3_w_n16481_0(.douta(w_n16481_0[0]),.doutb(w_n16481_0[1]),.doutc(w_n16481_0[2]),.din(n16481));
	jspl jspl_w_n16485_0(.douta(w_n16485_0[0]),.doutb(w_n16485_0[1]),.din(n16485));
	jspl jspl_w_n16491_0(.douta(w_n16491_0[0]),.doutb(w_n16491_0[1]),.din(n16491));
	jspl3 jspl3_w_n16493_0(.douta(w_n16493_0[0]),.doutb(w_n16493_0[1]),.doutc(w_n16493_0[2]),.din(n16493));
	jspl jspl_w_n16495_0(.douta(w_n16495_0[0]),.doutb(w_n16495_0[1]),.din(n16495));
	jspl3 jspl3_w_n16500_0(.douta(w_n16500_0[0]),.doutb(w_n16500_0[1]),.doutc(w_n16500_0[2]),.din(n16500));
	jspl jspl_w_n16501_0(.douta(w_n16501_0[0]),.doutb(w_n16501_0[1]),.din(n16501));
	jspl jspl_w_n16502_0(.douta(w_n16502_0[0]),.doutb(w_n16502_0[1]),.din(n16502));
	jspl jspl_w_n16507_0(.douta(w_n16507_0[0]),.doutb(w_n16507_0[1]),.din(n16507));
	jspl3 jspl3_w_n16508_0(.douta(w_n16508_0[0]),.doutb(w_n16508_0[1]),.doutc(w_n16508_0[2]),.din(n16508));
	jspl jspl_w_n16513_0(.douta(w_n16513_0[0]),.doutb(w_n16513_0[1]),.din(n16513));
	jspl jspl_w_n16521_0(.douta(w_n16521_0[0]),.doutb(w_n16521_0[1]),.din(n16521));
	jspl3 jspl3_w_n16523_0(.douta(w_n16523_0[0]),.doutb(w_n16523_0[1]),.doutc(w_n16523_0[2]),.din(n16523));
	jspl jspl_w_n16523_1(.douta(w_n16523_1[0]),.doutb(w_n16523_1[1]),.din(w_n16523_0[0]));
	jspl jspl_w_n16524_0(.douta(w_n16524_0[0]),.doutb(w_n16524_0[1]),.din(n16524));
	jspl3 jspl3_w_n16527_0(.douta(w_n16527_0[0]),.doutb(w_n16527_0[1]),.doutc(w_n16527_0[2]),.din(n16527));
	jspl jspl_w_n16528_0(.douta(w_n16528_0[0]),.doutb(w_n16528_0[1]),.din(n16528));
	jspl jspl_w_n16529_0(.douta(w_n16529_0[0]),.doutb(w_n16529_0[1]),.din(n16529));
	jspl jspl_w_n16530_0(.douta(w_n16530_0[0]),.doutb(w_n16530_0[1]),.din(n16530));
	jspl jspl_w_n16532_0(.douta(w_n16532_0[0]),.doutb(w_n16532_0[1]),.din(n16532));
	jspl jspl_w_n16534_0(.douta(w_n16534_0[0]),.doutb(w_n16534_0[1]),.din(n16534));
	jspl jspl_w_n16536_0(.douta(w_n16536_0[0]),.doutb(w_n16536_0[1]),.din(n16536));
	jspl jspl_w_n16545_0(.douta(w_n16545_0[0]),.doutb(w_n16545_0[1]),.din(n16545));
	jspl3 jspl3_w_n16547_0(.douta(w_n16547_0[0]),.doutb(w_n16547_0[1]),.doutc(w_n16547_0[2]),.din(n16547));
	jspl jspl_w_n16548_0(.douta(w_n16548_0[0]),.doutb(w_n16548_0[1]),.din(n16548));
	jspl jspl_w_n16552_0(.douta(w_n16552_0[0]),.doutb(w_n16552_0[1]),.din(n16552));
	jspl jspl_w_n16554_0(.douta(w_n16554_0[0]),.doutb(w_n16554_0[1]),.din(n16554));
	jspl jspl_w_n16556_0(.douta(w_n16556_0[0]),.doutb(w_n16556_0[1]),.din(n16556));
	jspl jspl_w_n16561_0(.douta(w_n16561_0[0]),.doutb(w_n16561_0[1]),.din(n16561));
	jspl jspl_w_n16563_0(.douta(w_n16563_0[0]),.doutb(w_n16563_0[1]),.din(n16563));
	jspl jspl_w_n16564_0(.douta(w_n16564_0[0]),.doutb(w_n16564_0[1]),.din(n16564));
	jspl3 jspl3_w_n16565_0(.douta(w_n16565_0[0]),.doutb(w_n16565_0[1]),.doutc(w_n16565_0[2]),.din(n16565));
	jspl jspl_w_n16566_0(.douta(w_n16566_0[0]),.doutb(w_n16566_0[1]),.din(n16566));
	jspl jspl_w_n16571_0(.douta(w_n16571_0[0]),.doutb(w_n16571_0[1]),.din(n16571));
	jspl jspl_w_n16572_0(.douta(w_n16572_0[0]),.doutb(w_n16572_0[1]),.din(n16572));
	jspl jspl_w_n16574_0(.douta(w_n16574_0[0]),.doutb(w_n16574_0[1]),.din(n16574));
	jspl jspl_w_n16576_0(.douta(w_n16576_0[0]),.doutb(w_n16576_0[1]),.din(n16576));
	jspl jspl_w_n16579_0(.douta(w_n16579_0[0]),.doutb(w_n16579_0[1]),.din(n16579));
	jspl jspl_w_n16585_0(.douta(w_n16585_0[0]),.doutb(w_n16585_0[1]),.din(n16585));
	jspl3 jspl3_w_n16587_0(.douta(w_n16587_0[0]),.doutb(w_n16587_0[1]),.doutc(w_n16587_0[2]),.din(n16587));
	jspl jspl_w_n16588_0(.douta(w_n16588_0[0]),.doutb(w_n16588_0[1]),.din(n16588));
	jspl jspl_w_n16592_0(.douta(w_n16592_0[0]),.doutb(w_n16592_0[1]),.din(n16592));
	jspl jspl_w_n16593_0(.douta(w_n16593_0[0]),.doutb(w_n16593_0[1]),.din(n16593));
	jspl jspl_w_n16595_0(.douta(w_n16595_0[0]),.doutb(w_n16595_0[1]),.din(n16595));
	jspl jspl_w_n16600_0(.douta(w_n16600_0[0]),.doutb(w_n16600_0[1]),.din(n16600));
	jspl jspl_w_n16602_0(.douta(w_n16602_0[0]),.doutb(w_n16602_0[1]),.din(n16602));
	jspl jspl_w_n16603_0(.douta(w_n16603_0[0]),.doutb(w_n16603_0[1]),.din(n16603));
	jspl3 jspl3_w_n16604_0(.douta(w_n16604_0[0]),.doutb(w_n16604_0[1]),.doutc(w_n16604_0[2]),.din(n16604));
	jspl jspl_w_n16605_0(.douta(w_n16605_0[0]),.doutb(w_n16605_0[1]),.din(n16605));
	jspl jspl_w_n16609_0(.douta(w_n16609_0[0]),.doutb(w_n16609_0[1]),.din(n16609));
	jspl jspl_w_n16610_0(.douta(w_n16610_0[0]),.doutb(w_n16610_0[1]),.din(n16610));
	jspl jspl_w_n16612_0(.douta(w_n16612_0[0]),.doutb(w_n16612_0[1]),.din(n16612));
	jspl jspl_w_n16614_0(.douta(w_n16614_0[0]),.doutb(w_n16614_0[1]),.din(n16614));
	jspl jspl_w_n16617_0(.douta(w_n16617_0[0]),.doutb(w_n16617_0[1]),.din(n16617));
	jspl jspl_w_n16623_0(.douta(w_n16623_0[0]),.doutb(w_n16623_0[1]),.din(n16623));
	jspl jspl_w_n16625_0(.douta(w_n16625_0[0]),.doutb(w_n16625_0[1]),.din(n16625));
	jspl3 jspl3_w_n16626_0(.douta(w_n16626_0[0]),.doutb(w_n16626_0[1]),.doutc(w_n16626_0[2]),.din(n16626));
	jspl jspl_w_n16630_0(.douta(w_n16630_0[0]),.doutb(w_n16630_0[1]),.din(n16630));
	jspl jspl_w_n16631_0(.douta(w_n16631_0[0]),.doutb(w_n16631_0[1]),.din(n16631));
	jspl3 jspl3_w_n16632_0(.douta(w_n16632_0[0]),.doutb(w_n16632_0[1]),.doutc(w_n16632_0[2]),.din(n16632));
	jspl jspl_w_n16634_0(.douta(w_n16634_0[0]),.doutb(w_n16634_0[1]),.din(n16634));
	jspl jspl_w_n16639_0(.douta(w_n16639_0[0]),.doutb(w_n16639_0[1]),.din(n16639));
	jspl jspl_w_n16641_0(.douta(w_n16641_0[0]),.doutb(w_n16641_0[1]),.din(n16641));
	jspl jspl_w_n16642_0(.douta(w_n16642_0[0]),.doutb(w_n16642_0[1]),.din(n16642));
	jspl3 jspl3_w_n16643_0(.douta(w_n16643_0[0]),.doutb(w_n16643_0[1]),.doutc(w_n16643_0[2]),.din(n16643));
	jspl jspl_w_n16644_0(.douta(w_n16644_0[0]),.doutb(w_n16644_0[1]),.din(n16644));
	jspl jspl_w_n16648_0(.douta(w_n16648_0[0]),.doutb(w_n16648_0[1]),.din(n16648));
	jspl jspl_w_n16654_0(.douta(w_n16654_0[0]),.doutb(w_n16654_0[1]),.din(n16654));
	jspl jspl_w_n16655_0(.douta(w_n16655_0[0]),.doutb(w_n16655_0[1]),.din(n16655));
	jspl jspl_w_n16657_0(.douta(w_n16657_0[0]),.doutb(w_n16657_0[1]),.din(n16657));
	jspl jspl_w_n16659_0(.douta(w_n16659_0[0]),.doutb(w_n16659_0[1]),.din(n16659));
	jspl jspl_w_n16662_0(.douta(w_n16662_0[0]),.doutb(w_n16662_0[1]),.din(n16662));
	jspl jspl_w_n16668_0(.douta(w_n16668_0[0]),.doutb(w_n16668_0[1]),.din(n16668));
	jspl jspl_w_n16670_0(.douta(w_n16670_0[0]),.doutb(w_n16670_0[1]),.din(n16670));
	jspl3 jspl3_w_n16671_0(.douta(w_n16671_0[0]),.doutb(w_n16671_0[1]),.doutc(w_n16671_0[2]),.din(n16671));
	jspl jspl_w_n16675_0(.douta(w_n16675_0[0]),.doutb(w_n16675_0[1]),.din(n16675));
	jspl jspl_w_n16676_0(.douta(w_n16676_0[0]),.doutb(w_n16676_0[1]),.din(n16676));
	jspl3 jspl3_w_n16677_0(.douta(w_n16677_0[0]),.doutb(w_n16677_0[1]),.doutc(w_n16677_0[2]),.din(n16677));
	jspl jspl_w_n16679_0(.douta(w_n16679_0[0]),.doutb(w_n16679_0[1]),.din(n16679));
	jspl jspl_w_n16684_0(.douta(w_n16684_0[0]),.doutb(w_n16684_0[1]),.din(n16684));
	jspl jspl_w_n16686_0(.douta(w_n16686_0[0]),.doutb(w_n16686_0[1]),.din(n16686));
	jspl jspl_w_n16687_0(.douta(w_n16687_0[0]),.doutb(w_n16687_0[1]),.din(n16687));
	jspl3 jspl3_w_n16688_0(.douta(w_n16688_0[0]),.doutb(w_n16688_0[1]),.doutc(w_n16688_0[2]),.din(n16688));
	jspl jspl_w_n16689_0(.douta(w_n16689_0[0]),.doutb(w_n16689_0[1]),.din(n16689));
	jspl jspl_w_n16693_0(.douta(w_n16693_0[0]),.doutb(w_n16693_0[1]),.din(n16693));
	jspl jspl_w_n16699_0(.douta(w_n16699_0[0]),.doutb(w_n16699_0[1]),.din(n16699));
	jspl jspl_w_n16700_0(.douta(w_n16700_0[0]),.doutb(w_n16700_0[1]),.din(n16700));
	jspl jspl_w_n16702_0(.douta(w_n16702_0[0]),.doutb(w_n16702_0[1]),.din(n16702));
	jspl jspl_w_n16704_0(.douta(w_n16704_0[0]),.doutb(w_n16704_0[1]),.din(n16704));
	jspl jspl_w_n16707_0(.douta(w_n16707_0[0]),.doutb(w_n16707_0[1]),.din(n16707));
	jspl jspl_w_n16713_0(.douta(w_n16713_0[0]),.doutb(w_n16713_0[1]),.din(n16713));
	jspl jspl_w_n16715_0(.douta(w_n16715_0[0]),.doutb(w_n16715_0[1]),.din(n16715));
	jspl3 jspl3_w_n16716_0(.douta(w_n16716_0[0]),.doutb(w_n16716_0[1]),.doutc(w_n16716_0[2]),.din(n16716));
	jspl jspl_w_n16720_0(.douta(w_n16720_0[0]),.doutb(w_n16720_0[1]),.din(n16720));
	jspl jspl_w_n16721_0(.douta(w_n16721_0[0]),.doutb(w_n16721_0[1]),.din(n16721));
	jspl3 jspl3_w_n16722_0(.douta(w_n16722_0[0]),.doutb(w_n16722_0[1]),.doutc(w_n16722_0[2]),.din(n16722));
	jspl jspl_w_n16724_0(.douta(w_n16724_0[0]),.doutb(w_n16724_0[1]),.din(n16724));
	jspl jspl_w_n16729_0(.douta(w_n16729_0[0]),.doutb(w_n16729_0[1]),.din(n16729));
	jspl jspl_w_n16731_0(.douta(w_n16731_0[0]),.doutb(w_n16731_0[1]),.din(n16731));
	jspl jspl_w_n16732_0(.douta(w_n16732_0[0]),.doutb(w_n16732_0[1]),.din(n16732));
	jspl3 jspl3_w_n16733_0(.douta(w_n16733_0[0]),.doutb(w_n16733_0[1]),.doutc(w_n16733_0[2]),.din(n16733));
	jspl jspl_w_n16734_0(.douta(w_n16734_0[0]),.doutb(w_n16734_0[1]),.din(n16734));
	jspl jspl_w_n16738_0(.douta(w_n16738_0[0]),.doutb(w_n16738_0[1]),.din(n16738));
	jspl jspl_w_n16744_0(.douta(w_n16744_0[0]),.doutb(w_n16744_0[1]),.din(n16744));
	jspl jspl_w_n16745_0(.douta(w_n16745_0[0]),.doutb(w_n16745_0[1]),.din(n16745));
	jspl jspl_w_n16747_0(.douta(w_n16747_0[0]),.doutb(w_n16747_0[1]),.din(n16747));
	jspl jspl_w_n16749_0(.douta(w_n16749_0[0]),.doutb(w_n16749_0[1]),.din(n16749));
	jspl jspl_w_n16752_0(.douta(w_n16752_0[0]),.doutb(w_n16752_0[1]),.din(n16752));
	jspl jspl_w_n16758_0(.douta(w_n16758_0[0]),.doutb(w_n16758_0[1]),.din(n16758));
	jspl jspl_w_n16760_0(.douta(w_n16760_0[0]),.doutb(w_n16760_0[1]),.din(n16760));
	jspl3 jspl3_w_n16761_0(.douta(w_n16761_0[0]),.doutb(w_n16761_0[1]),.doutc(w_n16761_0[2]),.din(n16761));
	jspl jspl_w_n16765_0(.douta(w_n16765_0[0]),.doutb(w_n16765_0[1]),.din(n16765));
	jspl jspl_w_n16766_0(.douta(w_n16766_0[0]),.doutb(w_n16766_0[1]),.din(n16766));
	jspl3 jspl3_w_n16767_0(.douta(w_n16767_0[0]),.doutb(w_n16767_0[1]),.doutc(w_n16767_0[2]),.din(n16767));
	jspl jspl_w_n16769_0(.douta(w_n16769_0[0]),.doutb(w_n16769_0[1]),.din(n16769));
	jspl jspl_w_n16774_0(.douta(w_n16774_0[0]),.doutb(w_n16774_0[1]),.din(n16774));
	jspl jspl_w_n16776_0(.douta(w_n16776_0[0]),.doutb(w_n16776_0[1]),.din(n16776));
	jspl jspl_w_n16777_0(.douta(w_n16777_0[0]),.doutb(w_n16777_0[1]),.din(n16777));
	jspl3 jspl3_w_n16778_0(.douta(w_n16778_0[0]),.doutb(w_n16778_0[1]),.doutc(w_n16778_0[2]),.din(n16778));
	jspl jspl_w_n16779_0(.douta(w_n16779_0[0]),.doutb(w_n16779_0[1]),.din(n16779));
	jspl jspl_w_n16783_0(.douta(w_n16783_0[0]),.doutb(w_n16783_0[1]),.din(n16783));
	jspl jspl_w_n16789_0(.douta(w_n16789_0[0]),.doutb(w_n16789_0[1]),.din(n16789));
	jspl jspl_w_n16790_0(.douta(w_n16790_0[0]),.doutb(w_n16790_0[1]),.din(n16790));
	jspl jspl_w_n16792_0(.douta(w_n16792_0[0]),.doutb(w_n16792_0[1]),.din(n16792));
	jspl jspl_w_n16794_0(.douta(w_n16794_0[0]),.doutb(w_n16794_0[1]),.din(n16794));
	jspl jspl_w_n16797_0(.douta(w_n16797_0[0]),.doutb(w_n16797_0[1]),.din(n16797));
	jspl jspl_w_n16803_0(.douta(w_n16803_0[0]),.doutb(w_n16803_0[1]),.din(n16803));
	jspl jspl_w_n16805_0(.douta(w_n16805_0[0]),.doutb(w_n16805_0[1]),.din(n16805));
	jspl3 jspl3_w_n16806_0(.douta(w_n16806_0[0]),.doutb(w_n16806_0[1]),.doutc(w_n16806_0[2]),.din(n16806));
	jspl jspl_w_n16810_0(.douta(w_n16810_0[0]),.doutb(w_n16810_0[1]),.din(n16810));
	jspl jspl_w_n16811_0(.douta(w_n16811_0[0]),.doutb(w_n16811_0[1]),.din(n16811));
	jspl3 jspl3_w_n16812_0(.douta(w_n16812_0[0]),.doutb(w_n16812_0[1]),.doutc(w_n16812_0[2]),.din(n16812));
	jspl jspl_w_n16814_0(.douta(w_n16814_0[0]),.doutb(w_n16814_0[1]),.din(n16814));
	jspl jspl_w_n16819_0(.douta(w_n16819_0[0]),.doutb(w_n16819_0[1]),.din(n16819));
	jspl jspl_w_n16821_0(.douta(w_n16821_0[0]),.doutb(w_n16821_0[1]),.din(n16821));
	jspl jspl_w_n16822_0(.douta(w_n16822_0[0]),.doutb(w_n16822_0[1]),.din(n16822));
	jspl3 jspl3_w_n16823_0(.douta(w_n16823_0[0]),.doutb(w_n16823_0[1]),.doutc(w_n16823_0[2]),.din(n16823));
	jspl jspl_w_n16824_0(.douta(w_n16824_0[0]),.doutb(w_n16824_0[1]),.din(n16824));
	jspl jspl_w_n16828_0(.douta(w_n16828_0[0]),.doutb(w_n16828_0[1]),.din(n16828));
	jspl jspl_w_n16834_0(.douta(w_n16834_0[0]),.doutb(w_n16834_0[1]),.din(n16834));
	jspl jspl_w_n16835_0(.douta(w_n16835_0[0]),.doutb(w_n16835_0[1]),.din(n16835));
	jspl jspl_w_n16837_0(.douta(w_n16837_0[0]),.doutb(w_n16837_0[1]),.din(n16837));
	jspl jspl_w_n16839_0(.douta(w_n16839_0[0]),.doutb(w_n16839_0[1]),.din(n16839));
	jspl jspl_w_n16842_0(.douta(w_n16842_0[0]),.doutb(w_n16842_0[1]),.din(n16842));
	jspl jspl_w_n16848_0(.douta(w_n16848_0[0]),.doutb(w_n16848_0[1]),.din(n16848));
	jspl jspl_w_n16850_0(.douta(w_n16850_0[0]),.doutb(w_n16850_0[1]),.din(n16850));
	jspl3 jspl3_w_n16851_0(.douta(w_n16851_0[0]),.doutb(w_n16851_0[1]),.doutc(w_n16851_0[2]),.din(n16851));
	jspl jspl_w_n16855_0(.douta(w_n16855_0[0]),.doutb(w_n16855_0[1]),.din(n16855));
	jspl jspl_w_n16856_0(.douta(w_n16856_0[0]),.doutb(w_n16856_0[1]),.din(n16856));
	jspl3 jspl3_w_n16857_0(.douta(w_n16857_0[0]),.doutb(w_n16857_0[1]),.doutc(w_n16857_0[2]),.din(n16857));
	jspl jspl_w_n16859_0(.douta(w_n16859_0[0]),.doutb(w_n16859_0[1]),.din(n16859));
	jspl jspl_w_n16864_0(.douta(w_n16864_0[0]),.doutb(w_n16864_0[1]),.din(n16864));
	jspl jspl_w_n16866_0(.douta(w_n16866_0[0]),.doutb(w_n16866_0[1]),.din(n16866));
	jspl jspl_w_n16867_0(.douta(w_n16867_0[0]),.doutb(w_n16867_0[1]),.din(n16867));
	jspl3 jspl3_w_n16868_0(.douta(w_n16868_0[0]),.doutb(w_n16868_0[1]),.doutc(w_n16868_0[2]),.din(n16868));
	jspl jspl_w_n16869_0(.douta(w_n16869_0[0]),.doutb(w_n16869_0[1]),.din(n16869));
	jspl jspl_w_n16873_0(.douta(w_n16873_0[0]),.doutb(w_n16873_0[1]),.din(n16873));
	jspl jspl_w_n16879_0(.douta(w_n16879_0[0]),.doutb(w_n16879_0[1]),.din(n16879));
	jspl jspl_w_n16880_0(.douta(w_n16880_0[0]),.doutb(w_n16880_0[1]),.din(n16880));
	jspl jspl_w_n16882_0(.douta(w_n16882_0[0]),.doutb(w_n16882_0[1]),.din(n16882));
	jspl jspl_w_n16884_0(.douta(w_n16884_0[0]),.doutb(w_n16884_0[1]),.din(n16884));
	jspl jspl_w_n16887_0(.douta(w_n16887_0[0]),.doutb(w_n16887_0[1]),.din(n16887));
	jspl jspl_w_n16893_0(.douta(w_n16893_0[0]),.doutb(w_n16893_0[1]),.din(n16893));
	jspl jspl_w_n16895_0(.douta(w_n16895_0[0]),.doutb(w_n16895_0[1]),.din(n16895));
	jspl3 jspl3_w_n16896_0(.douta(w_n16896_0[0]),.doutb(w_n16896_0[1]),.doutc(w_n16896_0[2]),.din(n16896));
	jspl jspl_w_n16900_0(.douta(w_n16900_0[0]),.doutb(w_n16900_0[1]),.din(n16900));
	jspl jspl_w_n16901_0(.douta(w_n16901_0[0]),.doutb(w_n16901_0[1]),.din(n16901));
	jspl3 jspl3_w_n16902_0(.douta(w_n16902_0[0]),.doutb(w_n16902_0[1]),.doutc(w_n16902_0[2]),.din(n16902));
	jspl jspl_w_n16904_0(.douta(w_n16904_0[0]),.doutb(w_n16904_0[1]),.din(n16904));
	jspl jspl_w_n16909_0(.douta(w_n16909_0[0]),.doutb(w_n16909_0[1]),.din(n16909));
	jspl jspl_w_n16911_0(.douta(w_n16911_0[0]),.doutb(w_n16911_0[1]),.din(n16911));
	jspl jspl_w_n16912_0(.douta(w_n16912_0[0]),.doutb(w_n16912_0[1]),.din(n16912));
	jspl3 jspl3_w_n16913_0(.douta(w_n16913_0[0]),.doutb(w_n16913_0[1]),.doutc(w_n16913_0[2]),.din(n16913));
	jspl jspl_w_n16914_0(.douta(w_n16914_0[0]),.doutb(w_n16914_0[1]),.din(n16914));
	jspl jspl_w_n16918_0(.douta(w_n16918_0[0]),.doutb(w_n16918_0[1]),.din(n16918));
	jspl jspl_w_n16924_0(.douta(w_n16924_0[0]),.doutb(w_n16924_0[1]),.din(n16924));
	jspl jspl_w_n16925_0(.douta(w_n16925_0[0]),.doutb(w_n16925_0[1]),.din(n16925));
	jspl jspl_w_n16927_0(.douta(w_n16927_0[0]),.doutb(w_n16927_0[1]),.din(n16927));
	jspl jspl_w_n16929_0(.douta(w_n16929_0[0]),.doutb(w_n16929_0[1]),.din(n16929));
	jspl jspl_w_n16932_0(.douta(w_n16932_0[0]),.doutb(w_n16932_0[1]),.din(n16932));
	jspl jspl_w_n16938_0(.douta(w_n16938_0[0]),.doutb(w_n16938_0[1]),.din(n16938));
	jspl jspl_w_n16940_0(.douta(w_n16940_0[0]),.doutb(w_n16940_0[1]),.din(n16940));
	jspl3 jspl3_w_n16941_0(.douta(w_n16941_0[0]),.doutb(w_n16941_0[1]),.doutc(w_n16941_0[2]),.din(n16941));
	jspl jspl_w_n16945_0(.douta(w_n16945_0[0]),.doutb(w_n16945_0[1]),.din(n16945));
	jspl jspl_w_n16946_0(.douta(w_n16946_0[0]),.doutb(w_n16946_0[1]),.din(n16946));
	jspl3 jspl3_w_n16947_0(.douta(w_n16947_0[0]),.doutb(w_n16947_0[1]),.doutc(w_n16947_0[2]),.din(n16947));
	jspl jspl_w_n16949_0(.douta(w_n16949_0[0]),.doutb(w_n16949_0[1]),.din(n16949));
	jspl jspl_w_n16954_0(.douta(w_n16954_0[0]),.doutb(w_n16954_0[1]),.din(n16954));
	jspl jspl_w_n16956_0(.douta(w_n16956_0[0]),.doutb(w_n16956_0[1]),.din(n16956));
	jspl jspl_w_n16957_0(.douta(w_n16957_0[0]),.doutb(w_n16957_0[1]),.din(n16957));
	jspl3 jspl3_w_n16958_0(.douta(w_n16958_0[0]),.doutb(w_n16958_0[1]),.doutc(w_n16958_0[2]),.din(n16958));
	jspl jspl_w_n16959_0(.douta(w_n16959_0[0]),.doutb(w_n16959_0[1]),.din(n16959));
	jspl jspl_w_n16963_0(.douta(w_n16963_0[0]),.doutb(w_n16963_0[1]),.din(n16963));
	jspl jspl_w_n16969_0(.douta(w_n16969_0[0]),.doutb(w_n16969_0[1]),.din(n16969));
	jspl jspl_w_n16970_0(.douta(w_n16970_0[0]),.doutb(w_n16970_0[1]),.din(n16970));
	jspl jspl_w_n16972_0(.douta(w_n16972_0[0]),.doutb(w_n16972_0[1]),.din(n16972));
	jspl jspl_w_n16974_0(.douta(w_n16974_0[0]),.doutb(w_n16974_0[1]),.din(n16974));
	jspl jspl_w_n16977_0(.douta(w_n16977_0[0]),.doutb(w_n16977_0[1]),.din(n16977));
	jspl jspl_w_n16983_0(.douta(w_n16983_0[0]),.doutb(w_n16983_0[1]),.din(n16983));
	jspl jspl_w_n16985_0(.douta(w_n16985_0[0]),.doutb(w_n16985_0[1]),.din(n16985));
	jspl3 jspl3_w_n16986_0(.douta(w_n16986_0[0]),.doutb(w_n16986_0[1]),.doutc(w_n16986_0[2]),.din(n16986));
	jspl jspl_w_n16990_0(.douta(w_n16990_0[0]),.doutb(w_n16990_0[1]),.din(n16990));
	jspl jspl_w_n16991_0(.douta(w_n16991_0[0]),.doutb(w_n16991_0[1]),.din(n16991));
	jspl3 jspl3_w_n16992_0(.douta(w_n16992_0[0]),.doutb(w_n16992_0[1]),.doutc(w_n16992_0[2]),.din(n16992));
	jspl jspl_w_n16994_0(.douta(w_n16994_0[0]),.doutb(w_n16994_0[1]),.din(n16994));
	jspl jspl_w_n16999_0(.douta(w_n16999_0[0]),.doutb(w_n16999_0[1]),.din(n16999));
	jspl jspl_w_n17001_0(.douta(w_n17001_0[0]),.doutb(w_n17001_0[1]),.din(n17001));
	jspl jspl_w_n17002_0(.douta(w_n17002_0[0]),.doutb(w_n17002_0[1]),.din(n17002));
	jspl3 jspl3_w_n17003_0(.douta(w_n17003_0[0]),.doutb(w_n17003_0[1]),.doutc(w_n17003_0[2]),.din(n17003));
	jspl jspl_w_n17004_0(.douta(w_n17004_0[0]),.doutb(w_n17004_0[1]),.din(n17004));
	jspl jspl_w_n17008_0(.douta(w_n17008_0[0]),.doutb(w_n17008_0[1]),.din(n17008));
	jspl jspl_w_n17014_0(.douta(w_n17014_0[0]),.doutb(w_n17014_0[1]),.din(n17014));
	jspl jspl_w_n17015_0(.douta(w_n17015_0[0]),.doutb(w_n17015_0[1]),.din(n17015));
	jspl jspl_w_n17017_0(.douta(w_n17017_0[0]),.doutb(w_n17017_0[1]),.din(n17017));
	jspl jspl_w_n17022_0(.douta(w_n17022_0[0]),.doutb(w_n17022_0[1]),.din(n17022));
	jspl jspl_w_n17024_0(.douta(w_n17024_0[0]),.doutb(w_n17024_0[1]),.din(n17024));
	jspl jspl_w_n17025_0(.douta(w_n17025_0[0]),.doutb(w_n17025_0[1]),.din(n17025));
	jspl3 jspl3_w_n17026_0(.douta(w_n17026_0[0]),.doutb(w_n17026_0[1]),.doutc(w_n17026_0[2]),.din(n17026));
	jspl jspl_w_n17027_0(.douta(w_n17027_0[0]),.doutb(w_n17027_0[1]),.din(n17027));
	jspl jspl_w_n17029_0(.douta(w_n17029_0[0]),.doutb(w_n17029_0[1]),.din(n17029));
	jspl jspl_w_n17031_0(.douta(w_n17031_0[0]),.doutb(w_n17031_0[1]),.din(n17031));
	jspl jspl_w_n17033_0(.douta(w_n17033_0[0]),.doutb(w_n17033_0[1]),.din(n17033));
	jspl jspl_w_n17036_0(.douta(w_n17036_0[0]),.doutb(w_n17036_0[1]),.din(n17036));
	jspl jspl_w_n17042_0(.douta(w_n17042_0[0]),.doutb(w_n17042_0[1]),.din(n17042));
	jspl3 jspl3_w_n17044_0(.douta(w_n17044_0[0]),.doutb(w_n17044_0[1]),.doutc(w_n17044_0[2]),.din(n17044));
	jspl jspl_w_n17045_0(.douta(w_n17045_0[0]),.doutb(w_n17045_0[1]),.din(n17045));
	jspl jspl_w_n17049_0(.douta(w_n17049_0[0]),.doutb(w_n17049_0[1]),.din(n17049));
	jspl jspl_w_n17055_0(.douta(w_n17055_0[0]),.doutb(w_n17055_0[1]),.din(n17055));
	jspl jspl_w_n17056_0(.douta(w_n17056_0[0]),.doutb(w_n17056_0[1]),.din(n17056));
	jspl jspl_w_n17058_0(.douta(w_n17058_0[0]),.doutb(w_n17058_0[1]),.din(n17058));
	jspl jspl_w_n17060_0(.douta(w_n17060_0[0]),.doutb(w_n17060_0[1]),.din(n17060));
	jspl jspl_w_n17063_0(.douta(w_n17063_0[0]),.doutb(w_n17063_0[1]),.din(n17063));
	jspl jspl_w_n17069_0(.douta(w_n17069_0[0]),.doutb(w_n17069_0[1]),.din(n17069));
	jspl jspl_w_n17071_0(.douta(w_n17071_0[0]),.doutb(w_n17071_0[1]),.din(n17071));
	jspl3 jspl3_w_n17072_0(.douta(w_n17072_0[0]),.doutb(w_n17072_0[1]),.doutc(w_n17072_0[2]),.din(n17072));
	jspl jspl_w_n17076_0(.douta(w_n17076_0[0]),.doutb(w_n17076_0[1]),.din(n17076));
	jspl jspl_w_n17077_0(.douta(w_n17077_0[0]),.doutb(w_n17077_0[1]),.din(n17077));
	jspl3 jspl3_w_n17078_0(.douta(w_n17078_0[0]),.doutb(w_n17078_0[1]),.doutc(w_n17078_0[2]),.din(n17078));
	jspl jspl_w_n17080_0(.douta(w_n17080_0[0]),.doutb(w_n17080_0[1]),.din(n17080));
	jspl jspl_w_n17085_0(.douta(w_n17085_0[0]),.doutb(w_n17085_0[1]),.din(n17085));
	jspl jspl_w_n17087_0(.douta(w_n17087_0[0]),.doutb(w_n17087_0[1]),.din(n17087));
	jspl jspl_w_n17088_0(.douta(w_n17088_0[0]),.doutb(w_n17088_0[1]),.din(n17088));
	jspl3 jspl3_w_n17089_0(.douta(w_n17089_0[0]),.doutb(w_n17089_0[1]),.doutc(w_n17089_0[2]),.din(n17089));
	jspl jspl_w_n17090_0(.douta(w_n17090_0[0]),.doutb(w_n17090_0[1]),.din(n17090));
	jspl jspl_w_n17094_0(.douta(w_n17094_0[0]),.doutb(w_n17094_0[1]),.din(n17094));
	jspl jspl_w_n17100_0(.douta(w_n17100_0[0]),.doutb(w_n17100_0[1]),.din(n17100));
	jspl jspl_w_n17101_0(.douta(w_n17101_0[0]),.doutb(w_n17101_0[1]),.din(n17101));
	jspl jspl_w_n17103_0(.douta(w_n17103_0[0]),.doutb(w_n17103_0[1]),.din(n17103));
	jspl jspl_w_n17105_0(.douta(w_n17105_0[0]),.doutb(w_n17105_0[1]),.din(n17105));
	jspl jspl_w_n17108_0(.douta(w_n17108_0[0]),.doutb(w_n17108_0[1]),.din(n17108));
	jspl jspl_w_n17114_0(.douta(w_n17114_0[0]),.doutb(w_n17114_0[1]),.din(n17114));
	jspl3 jspl3_w_n17116_0(.douta(w_n17116_0[0]),.doutb(w_n17116_0[1]),.doutc(w_n17116_0[2]),.din(n17116));
	jspl3 jspl3_w_n17116_1(.douta(w_n17116_1[0]),.doutb(w_n17116_1[1]),.doutc(w_n17116_1[2]),.din(w_n17116_0[0]));
	jspl jspl_w_n17119_0(.douta(w_n17119_0[0]),.doutb(w_n17119_0[1]),.din(n17119));
	jspl3 jspl3_w_n17120_0(.douta(w_n17120_0[0]),.doutb(w_n17120_0[1]),.doutc(w_n17120_0[2]),.din(n17120));
	jspl jspl_w_n17121_0(.douta(w_n17121_0[0]),.doutb(w_n17121_0[1]),.din(n17121));
	jspl jspl_w_n17127_0(.douta(w_n17127_0[0]),.doutb(w_n17127_0[1]),.din(n17127));
	jspl3 jspl3_w_n17128_0(.douta(w_n17128_0[0]),.doutb(w_n17128_0[1]),.doutc(w_n17128_0[2]),.din(n17128));
	jspl jspl_w_n17129_0(.douta(w_n17129_0[0]),.doutb(w_n17129_0[1]),.din(n17129));
	jspl jspl_w_n17134_0(.douta(w_n17134_0[0]),.doutb(w_n17134_0[1]),.din(n17134));
	jspl3 jspl3_w_n17135_0(.douta(w_n17135_0[0]),.doutb(w_n17135_0[1]),.doutc(w_n17135_0[2]),.din(n17135));
	jspl3 jspl3_w_n17135_1(.douta(w_n17135_1[0]),.doutb(w_n17135_1[1]),.doutc(w_n17135_1[2]),.din(w_n17135_0[0]));
	jspl3 jspl3_w_n17135_2(.douta(w_n17135_2[0]),.doutb(w_n17135_2[1]),.doutc(w_n17135_2[2]),.din(w_n17135_0[1]));
	jspl3 jspl3_w_n17135_3(.douta(w_n17135_3[0]),.doutb(w_n17135_3[1]),.doutc(w_n17135_3[2]),.din(w_n17135_0[2]));
	jspl3 jspl3_w_n17135_4(.douta(w_n17135_4[0]),.doutb(w_n17135_4[1]),.doutc(w_n17135_4[2]),.din(w_n17135_1[0]));
	jspl jspl_w_n17135_5(.douta(w_n17135_5[0]),.doutb(w_n17135_5[1]),.din(w_n17135_1[1]));
	jspl3 jspl3_w_n17140_0(.douta(w_n17140_0[0]),.doutb(w_n17140_0[1]),.doutc(w_n17140_0[2]),.din(n17140));
	jspl3 jspl3_w_n17140_1(.douta(w_n17140_1[0]),.doutb(w_n17140_1[1]),.doutc(w_n17140_1[2]),.din(w_n17140_0[0]));
	jspl3 jspl3_w_n17140_2(.douta(w_n17140_2[0]),.doutb(w_n17140_2[1]),.doutc(w_n17140_2[2]),.din(w_n17140_0[1]));
	jspl3 jspl3_w_n17140_3(.douta(w_n17140_3[0]),.doutb(w_n17140_3[1]),.doutc(w_n17140_3[2]),.din(w_n17140_0[2]));
	jspl3 jspl3_w_n17140_4(.douta(w_n17140_4[0]),.doutb(w_n17140_4[1]),.doutc(w_n17140_4[2]),.din(w_n17140_1[0]));
	jspl3 jspl3_w_n17140_5(.douta(w_n17140_5[0]),.doutb(w_n17140_5[1]),.doutc(w_n17140_5[2]),.din(w_n17140_1[1]));
	jspl3 jspl3_w_n17140_6(.douta(w_n17140_6[0]),.doutb(w_n17140_6[1]),.doutc(w_n17140_6[2]),.din(w_n17140_1[2]));
	jspl3 jspl3_w_n17140_7(.douta(w_n17140_7[0]),.doutb(w_n17140_7[1]),.doutc(w_n17140_7[2]),.din(w_n17140_2[0]));
	jspl3 jspl3_w_n17140_8(.douta(w_n17140_8[0]),.doutb(w_n17140_8[1]),.doutc(w_n17140_8[2]),.din(w_n17140_2[1]));
	jspl3 jspl3_w_n17140_9(.douta(w_n17140_9[0]),.doutb(w_n17140_9[1]),.doutc(w_n17140_9[2]),.din(w_n17140_2[2]));
	jspl3 jspl3_w_n17140_10(.douta(w_n17140_10[0]),.doutb(w_n17140_10[1]),.doutc(w_n17140_10[2]),.din(w_n17140_3[0]));
	jspl3 jspl3_w_n17140_11(.douta(w_n17140_11[0]),.doutb(w_n17140_11[1]),.doutc(w_n17140_11[2]),.din(w_n17140_3[1]));
	jspl3 jspl3_w_n17140_12(.douta(w_n17140_12[0]),.doutb(w_n17140_12[1]),.doutc(w_n17140_12[2]),.din(w_n17140_3[2]));
	jspl3 jspl3_w_n17140_13(.douta(w_n17140_13[0]),.doutb(w_n17140_13[1]),.doutc(w_n17140_13[2]),.din(w_n17140_4[0]));
	jspl3 jspl3_w_n17140_14(.douta(w_n17140_14[0]),.doutb(w_n17140_14[1]),.doutc(w_n17140_14[2]),.din(w_n17140_4[1]));
	jspl3 jspl3_w_n17140_15(.douta(w_n17140_15[0]),.doutb(w_n17140_15[1]),.doutc(w_n17140_15[2]),.din(w_n17140_4[2]));
	jspl3 jspl3_w_n17140_16(.douta(w_n17140_16[0]),.doutb(w_n17140_16[1]),.doutc(w_n17140_16[2]),.din(w_n17140_5[0]));
	jspl3 jspl3_w_n17140_17(.douta(w_n17140_17[0]),.doutb(w_n17140_17[1]),.doutc(w_n17140_17[2]),.din(w_n17140_5[1]));
	jspl3 jspl3_w_n17140_18(.douta(w_n17140_18[0]),.doutb(w_n17140_18[1]),.doutc(w_n17140_18[2]),.din(w_n17140_5[2]));
	jspl3 jspl3_w_n17140_19(.douta(w_n17140_19[0]),.doutb(w_n17140_19[1]),.doutc(w_n17140_19[2]),.din(w_n17140_6[0]));
	jspl3 jspl3_w_n17140_20(.douta(w_n17140_20[0]),.doutb(w_n17140_20[1]),.doutc(w_n17140_20[2]),.din(w_n17140_6[1]));
	jspl jspl_w_n17143_0(.douta(w_n17143_0[0]),.doutb(w_n17143_0[1]),.din(n17143));
	jspl3 jspl3_w_n17145_0(.douta(w_n17145_0[0]),.doutb(w_n17145_0[1]),.doutc(w_n17145_0[2]),.din(n17145));
	jspl jspl_w_n17145_1(.douta(w_n17145_1[0]),.doutb(w_n17145_1[1]),.din(w_n17145_0[0]));
	jspl3 jspl3_w_n17146_0(.douta(w_n17146_0[0]),.doutb(w_n17146_0[1]),.doutc(w_n17146_0[2]),.din(n17146));
	jspl3 jspl3_w_n17150_0(.douta(w_n17150_0[0]),.doutb(w_n17150_0[1]),.doutc(w_n17150_0[2]),.din(n17150));
	jspl jspl_w_n17151_0(.douta(w_n17151_0[0]),.doutb(w_n17151_0[1]),.din(n17151));
	jspl jspl_w_n17152_0(.douta(w_n17152_0[0]),.doutb(w_n17152_0[1]),.din(n17152));
	jspl jspl_w_n17153_0(.douta(w_n17153_0[0]),.doutb(w_n17153_0[1]),.din(n17153));
	jspl jspl_w_n17155_0(.douta(w_n17155_0[0]),.doutb(w_n17155_0[1]),.din(n17155));
	jspl jspl_w_n17157_0(.douta(w_n17157_0[0]),.doutb(w_n17157_0[1]),.din(n17157));
	jspl jspl_w_n17159_0(.douta(w_n17159_0[0]),.doutb(w_n17159_0[1]),.din(n17159));
	jspl jspl_w_n17162_0(.douta(w_n17162_0[0]),.doutb(w_n17162_0[1]),.din(n17162));
	jspl jspl_w_n17167_0(.douta(w_n17167_0[0]),.doutb(w_n17167_0[1]),.din(n17167));
	jspl3 jspl3_w_n17169_0(.douta(w_n17169_0[0]),.doutb(w_n17169_0[1]),.doutc(w_n17169_0[2]),.din(n17169));
	jspl jspl_w_n17170_0(.douta(w_n17170_0[0]),.doutb(w_n17170_0[1]),.din(n17170));
	jspl jspl_w_n17174_0(.douta(w_n17174_0[0]),.doutb(w_n17174_0[1]),.din(n17174));
	jspl jspl_w_n17175_0(.douta(w_n17175_0[0]),.doutb(w_n17175_0[1]),.din(n17175));
	jspl jspl_w_n17177_0(.douta(w_n17177_0[0]),.doutb(w_n17177_0[1]),.din(n17177));
	jspl jspl_w_n17181_0(.douta(w_n17181_0[0]),.doutb(w_n17181_0[1]),.din(n17181));
	jspl jspl_w_n17183_0(.douta(w_n17183_0[0]),.doutb(w_n17183_0[1]),.din(n17183));
	jspl jspl_w_n17184_0(.douta(w_n17184_0[0]),.doutb(w_n17184_0[1]),.din(n17184));
	jspl3 jspl3_w_n17185_0(.douta(w_n17185_0[0]),.doutb(w_n17185_0[1]),.doutc(w_n17185_0[2]),.din(n17185));
	jspl jspl_w_n17186_0(.douta(w_n17186_0[0]),.doutb(w_n17186_0[1]),.din(n17186));
	jspl jspl_w_n17190_0(.douta(w_n17190_0[0]),.doutb(w_n17190_0[1]),.din(n17190));
	jspl jspl_w_n17192_0(.douta(w_n17192_0[0]),.doutb(w_n17192_0[1]),.din(n17192));
	jspl jspl_w_n17194_0(.douta(w_n17194_0[0]),.doutb(w_n17194_0[1]),.din(n17194));
	jspl jspl_w_n17196_0(.douta(w_n17196_0[0]),.doutb(w_n17196_0[1]),.din(n17196));
	jspl jspl_w_n17199_0(.douta(w_n17199_0[0]),.doutb(w_n17199_0[1]),.din(n17199));
	jspl jspl_w_n17205_0(.douta(w_n17205_0[0]),.doutb(w_n17205_0[1]),.din(n17205));
	jspl3 jspl3_w_n17207_0(.douta(w_n17207_0[0]),.doutb(w_n17207_0[1]),.doutc(w_n17207_0[2]),.din(n17207));
	jspl jspl_w_n17208_0(.douta(w_n17208_0[0]),.doutb(w_n17208_0[1]),.din(n17208));
	jspl jspl_w_n17213_0(.douta(w_n17213_0[0]),.doutb(w_n17213_0[1]),.din(n17213));
	jspl jspl_w_n17215_0(.douta(w_n17215_0[0]),.doutb(w_n17215_0[1]),.din(n17215));
	jspl jspl_w_n17217_0(.douta(w_n17217_0[0]),.doutb(w_n17217_0[1]),.din(n17217));
	jspl jspl_w_n17221_0(.douta(w_n17221_0[0]),.doutb(w_n17221_0[1]),.din(n17221));
	jspl jspl_w_n17223_0(.douta(w_n17223_0[0]),.doutb(w_n17223_0[1]),.din(n17223));
	jspl jspl_w_n17224_0(.douta(w_n17224_0[0]),.doutb(w_n17224_0[1]),.din(n17224));
	jspl3 jspl3_w_n17225_0(.douta(w_n17225_0[0]),.doutb(w_n17225_0[1]),.doutc(w_n17225_0[2]),.din(n17225));
	jspl jspl_w_n17226_0(.douta(w_n17226_0[0]),.doutb(w_n17226_0[1]),.din(n17226));
	jspl jspl_w_n17232_0(.douta(w_n17232_0[0]),.doutb(w_n17232_0[1]),.din(n17232));
	jspl jspl_w_n17233_0(.douta(w_n17233_0[0]),.doutb(w_n17233_0[1]),.din(n17233));
	jspl jspl_w_n17235_0(.douta(w_n17235_0[0]),.doutb(w_n17235_0[1]),.din(n17235));
	jspl jspl_w_n17237_0(.douta(w_n17237_0[0]),.doutb(w_n17237_0[1]),.din(n17237));
	jspl jspl_w_n17239_0(.douta(w_n17239_0[0]),.doutb(w_n17239_0[1]),.din(n17239));
	jspl jspl_w_n17245_0(.douta(w_n17245_0[0]),.doutb(w_n17245_0[1]),.din(n17245));
	jspl jspl_w_n17247_0(.douta(w_n17247_0[0]),.doutb(w_n17247_0[1]),.din(n17247));
	jspl3 jspl3_w_n17248_0(.douta(w_n17248_0[0]),.doutb(w_n17248_0[1]),.doutc(w_n17248_0[2]),.din(n17248));
	jspl jspl_w_n17251_0(.douta(w_n17251_0[0]),.doutb(w_n17251_0[1]),.din(n17251));
	jspl jspl_w_n17252_0(.douta(w_n17252_0[0]),.doutb(w_n17252_0[1]),.din(n17252));
	jspl3 jspl3_w_n17253_0(.douta(w_n17253_0[0]),.doutb(w_n17253_0[1]),.doutc(w_n17253_0[2]),.din(n17253));
	jspl jspl_w_n17255_0(.douta(w_n17255_0[0]),.doutb(w_n17255_0[1]),.din(n17255));
	jspl jspl_w_n17259_0(.douta(w_n17259_0[0]),.doutb(w_n17259_0[1]),.din(n17259));
	jspl jspl_w_n17261_0(.douta(w_n17261_0[0]),.doutb(w_n17261_0[1]),.din(n17261));
	jspl jspl_w_n17262_0(.douta(w_n17262_0[0]),.doutb(w_n17262_0[1]),.din(n17262));
	jspl3 jspl3_w_n17263_0(.douta(w_n17263_0[0]),.doutb(w_n17263_0[1]),.doutc(w_n17263_0[2]),.din(n17263));
	jspl jspl_w_n17264_0(.douta(w_n17264_0[0]),.doutb(w_n17264_0[1]),.din(n17264));
	jspl jspl_w_n17267_0(.douta(w_n17267_0[0]),.doutb(w_n17267_0[1]),.din(n17267));
	jspl jspl_w_n17273_0(.douta(w_n17273_0[0]),.doutb(w_n17273_0[1]),.din(n17273));
	jspl jspl_w_n17274_0(.douta(w_n17274_0[0]),.doutb(w_n17274_0[1]),.din(n17274));
	jspl jspl_w_n17276_0(.douta(w_n17276_0[0]),.doutb(w_n17276_0[1]),.din(n17276));
	jspl jspl_w_n17278_0(.douta(w_n17278_0[0]),.doutb(w_n17278_0[1]),.din(n17278));
	jspl jspl_w_n17280_0(.douta(w_n17280_0[0]),.doutb(w_n17280_0[1]),.din(n17280));
	jspl jspl_w_n17286_0(.douta(w_n17286_0[0]),.doutb(w_n17286_0[1]),.din(n17286));
	jspl jspl_w_n17288_0(.douta(w_n17288_0[0]),.doutb(w_n17288_0[1]),.din(n17288));
	jspl3 jspl3_w_n17289_0(.douta(w_n17289_0[0]),.doutb(w_n17289_0[1]),.doutc(w_n17289_0[2]),.din(n17289));
	jspl jspl_w_n17292_0(.douta(w_n17292_0[0]),.doutb(w_n17292_0[1]),.din(n17292));
	jspl jspl_w_n17293_0(.douta(w_n17293_0[0]),.doutb(w_n17293_0[1]),.din(n17293));
	jspl3 jspl3_w_n17294_0(.douta(w_n17294_0[0]),.doutb(w_n17294_0[1]),.doutc(w_n17294_0[2]),.din(n17294));
	jspl jspl_w_n17296_0(.douta(w_n17296_0[0]),.doutb(w_n17296_0[1]),.din(n17296));
	jspl jspl_w_n17300_0(.douta(w_n17300_0[0]),.doutb(w_n17300_0[1]),.din(n17300));
	jspl jspl_w_n17302_0(.douta(w_n17302_0[0]),.doutb(w_n17302_0[1]),.din(n17302));
	jspl jspl_w_n17303_0(.douta(w_n17303_0[0]),.doutb(w_n17303_0[1]),.din(n17303));
	jspl3 jspl3_w_n17304_0(.douta(w_n17304_0[0]),.doutb(w_n17304_0[1]),.doutc(w_n17304_0[2]),.din(n17304));
	jspl jspl_w_n17305_0(.douta(w_n17305_0[0]),.doutb(w_n17305_0[1]),.din(n17305));
	jspl jspl_w_n17308_0(.douta(w_n17308_0[0]),.doutb(w_n17308_0[1]),.din(n17308));
	jspl jspl_w_n17314_0(.douta(w_n17314_0[0]),.doutb(w_n17314_0[1]),.din(n17314));
	jspl jspl_w_n17315_0(.douta(w_n17315_0[0]),.doutb(w_n17315_0[1]),.din(n17315));
	jspl jspl_w_n17317_0(.douta(w_n17317_0[0]),.doutb(w_n17317_0[1]),.din(n17317));
	jspl jspl_w_n17319_0(.douta(w_n17319_0[0]),.doutb(w_n17319_0[1]),.din(n17319));
	jspl jspl_w_n17321_0(.douta(w_n17321_0[0]),.doutb(w_n17321_0[1]),.din(n17321));
	jspl jspl_w_n17327_0(.douta(w_n17327_0[0]),.doutb(w_n17327_0[1]),.din(n17327));
	jspl jspl_w_n17329_0(.douta(w_n17329_0[0]),.doutb(w_n17329_0[1]),.din(n17329));
	jspl3 jspl3_w_n17330_0(.douta(w_n17330_0[0]),.doutb(w_n17330_0[1]),.doutc(w_n17330_0[2]),.din(n17330));
	jspl jspl_w_n17333_0(.douta(w_n17333_0[0]),.doutb(w_n17333_0[1]),.din(n17333));
	jspl jspl_w_n17334_0(.douta(w_n17334_0[0]),.doutb(w_n17334_0[1]),.din(n17334));
	jspl3 jspl3_w_n17335_0(.douta(w_n17335_0[0]),.doutb(w_n17335_0[1]),.doutc(w_n17335_0[2]),.din(n17335));
	jspl jspl_w_n17337_0(.douta(w_n17337_0[0]),.doutb(w_n17337_0[1]),.din(n17337));
	jspl jspl_w_n17341_0(.douta(w_n17341_0[0]),.doutb(w_n17341_0[1]),.din(n17341));
	jspl jspl_w_n17343_0(.douta(w_n17343_0[0]),.doutb(w_n17343_0[1]),.din(n17343));
	jspl jspl_w_n17344_0(.douta(w_n17344_0[0]),.doutb(w_n17344_0[1]),.din(n17344));
	jspl3 jspl3_w_n17345_0(.douta(w_n17345_0[0]),.doutb(w_n17345_0[1]),.doutc(w_n17345_0[2]),.din(n17345));
	jspl jspl_w_n17346_0(.douta(w_n17346_0[0]),.doutb(w_n17346_0[1]),.din(n17346));
	jspl jspl_w_n17349_0(.douta(w_n17349_0[0]),.doutb(w_n17349_0[1]),.din(n17349));
	jspl jspl_w_n17355_0(.douta(w_n17355_0[0]),.doutb(w_n17355_0[1]),.din(n17355));
	jspl jspl_w_n17356_0(.douta(w_n17356_0[0]),.doutb(w_n17356_0[1]),.din(n17356));
	jspl jspl_w_n17358_0(.douta(w_n17358_0[0]),.doutb(w_n17358_0[1]),.din(n17358));
	jspl jspl_w_n17360_0(.douta(w_n17360_0[0]),.doutb(w_n17360_0[1]),.din(n17360));
	jspl jspl_w_n17362_0(.douta(w_n17362_0[0]),.doutb(w_n17362_0[1]),.din(n17362));
	jspl jspl_w_n17368_0(.douta(w_n17368_0[0]),.doutb(w_n17368_0[1]),.din(n17368));
	jspl jspl_w_n17370_0(.douta(w_n17370_0[0]),.doutb(w_n17370_0[1]),.din(n17370));
	jspl3 jspl3_w_n17371_0(.douta(w_n17371_0[0]),.doutb(w_n17371_0[1]),.doutc(w_n17371_0[2]),.din(n17371));
	jspl jspl_w_n17374_0(.douta(w_n17374_0[0]),.doutb(w_n17374_0[1]),.din(n17374));
	jspl jspl_w_n17375_0(.douta(w_n17375_0[0]),.doutb(w_n17375_0[1]),.din(n17375));
	jspl3 jspl3_w_n17376_0(.douta(w_n17376_0[0]),.doutb(w_n17376_0[1]),.doutc(w_n17376_0[2]),.din(n17376));
	jspl jspl_w_n17378_0(.douta(w_n17378_0[0]),.doutb(w_n17378_0[1]),.din(n17378));
	jspl jspl_w_n17382_0(.douta(w_n17382_0[0]),.doutb(w_n17382_0[1]),.din(n17382));
	jspl jspl_w_n17384_0(.douta(w_n17384_0[0]),.doutb(w_n17384_0[1]),.din(n17384));
	jspl jspl_w_n17385_0(.douta(w_n17385_0[0]),.doutb(w_n17385_0[1]),.din(n17385));
	jspl3 jspl3_w_n17386_0(.douta(w_n17386_0[0]),.doutb(w_n17386_0[1]),.doutc(w_n17386_0[2]),.din(n17386));
	jspl jspl_w_n17387_0(.douta(w_n17387_0[0]),.doutb(w_n17387_0[1]),.din(n17387));
	jspl jspl_w_n17390_0(.douta(w_n17390_0[0]),.doutb(w_n17390_0[1]),.din(n17390));
	jspl jspl_w_n17396_0(.douta(w_n17396_0[0]),.doutb(w_n17396_0[1]),.din(n17396));
	jspl jspl_w_n17397_0(.douta(w_n17397_0[0]),.doutb(w_n17397_0[1]),.din(n17397));
	jspl jspl_w_n17399_0(.douta(w_n17399_0[0]),.doutb(w_n17399_0[1]),.din(n17399));
	jspl jspl_w_n17401_0(.douta(w_n17401_0[0]),.doutb(w_n17401_0[1]),.din(n17401));
	jspl jspl_w_n17403_0(.douta(w_n17403_0[0]),.doutb(w_n17403_0[1]),.din(n17403));
	jspl jspl_w_n17409_0(.douta(w_n17409_0[0]),.doutb(w_n17409_0[1]),.din(n17409));
	jspl jspl_w_n17411_0(.douta(w_n17411_0[0]),.doutb(w_n17411_0[1]),.din(n17411));
	jspl3 jspl3_w_n17412_0(.douta(w_n17412_0[0]),.doutb(w_n17412_0[1]),.doutc(w_n17412_0[2]),.din(n17412));
	jspl jspl_w_n17415_0(.douta(w_n17415_0[0]),.doutb(w_n17415_0[1]),.din(n17415));
	jspl jspl_w_n17416_0(.douta(w_n17416_0[0]),.doutb(w_n17416_0[1]),.din(n17416));
	jspl3 jspl3_w_n17417_0(.douta(w_n17417_0[0]),.doutb(w_n17417_0[1]),.doutc(w_n17417_0[2]),.din(n17417));
	jspl jspl_w_n17419_0(.douta(w_n17419_0[0]),.doutb(w_n17419_0[1]),.din(n17419));
	jspl jspl_w_n17423_0(.douta(w_n17423_0[0]),.doutb(w_n17423_0[1]),.din(n17423));
	jspl jspl_w_n17425_0(.douta(w_n17425_0[0]),.doutb(w_n17425_0[1]),.din(n17425));
	jspl jspl_w_n17426_0(.douta(w_n17426_0[0]),.doutb(w_n17426_0[1]),.din(n17426));
	jspl3 jspl3_w_n17427_0(.douta(w_n17427_0[0]),.doutb(w_n17427_0[1]),.doutc(w_n17427_0[2]),.din(n17427));
	jspl jspl_w_n17428_0(.douta(w_n17428_0[0]),.doutb(w_n17428_0[1]),.din(n17428));
	jspl jspl_w_n17431_0(.douta(w_n17431_0[0]),.doutb(w_n17431_0[1]),.din(n17431));
	jspl jspl_w_n17437_0(.douta(w_n17437_0[0]),.doutb(w_n17437_0[1]),.din(n17437));
	jspl jspl_w_n17438_0(.douta(w_n17438_0[0]),.doutb(w_n17438_0[1]),.din(n17438));
	jspl jspl_w_n17440_0(.douta(w_n17440_0[0]),.doutb(w_n17440_0[1]),.din(n17440));
	jspl jspl_w_n17442_0(.douta(w_n17442_0[0]),.doutb(w_n17442_0[1]),.din(n17442));
	jspl jspl_w_n17444_0(.douta(w_n17444_0[0]),.doutb(w_n17444_0[1]),.din(n17444));
	jspl jspl_w_n17450_0(.douta(w_n17450_0[0]),.doutb(w_n17450_0[1]),.din(n17450));
	jspl jspl_w_n17452_0(.douta(w_n17452_0[0]),.doutb(w_n17452_0[1]),.din(n17452));
	jspl3 jspl3_w_n17453_0(.douta(w_n17453_0[0]),.doutb(w_n17453_0[1]),.doutc(w_n17453_0[2]),.din(n17453));
	jspl jspl_w_n17456_0(.douta(w_n17456_0[0]),.doutb(w_n17456_0[1]),.din(n17456));
	jspl jspl_w_n17457_0(.douta(w_n17457_0[0]),.doutb(w_n17457_0[1]),.din(n17457));
	jspl3 jspl3_w_n17458_0(.douta(w_n17458_0[0]),.doutb(w_n17458_0[1]),.doutc(w_n17458_0[2]),.din(n17458));
	jspl jspl_w_n17460_0(.douta(w_n17460_0[0]),.doutb(w_n17460_0[1]),.din(n17460));
	jspl jspl_w_n17464_0(.douta(w_n17464_0[0]),.doutb(w_n17464_0[1]),.din(n17464));
	jspl jspl_w_n17466_0(.douta(w_n17466_0[0]),.doutb(w_n17466_0[1]),.din(n17466));
	jspl jspl_w_n17467_0(.douta(w_n17467_0[0]),.doutb(w_n17467_0[1]),.din(n17467));
	jspl3 jspl3_w_n17468_0(.douta(w_n17468_0[0]),.doutb(w_n17468_0[1]),.doutc(w_n17468_0[2]),.din(n17468));
	jspl jspl_w_n17469_0(.douta(w_n17469_0[0]),.doutb(w_n17469_0[1]),.din(n17469));
	jspl jspl_w_n17472_0(.douta(w_n17472_0[0]),.doutb(w_n17472_0[1]),.din(n17472));
	jspl jspl_w_n17478_0(.douta(w_n17478_0[0]),.doutb(w_n17478_0[1]),.din(n17478));
	jspl jspl_w_n17479_0(.douta(w_n17479_0[0]),.doutb(w_n17479_0[1]),.din(n17479));
	jspl jspl_w_n17481_0(.douta(w_n17481_0[0]),.doutb(w_n17481_0[1]),.din(n17481));
	jspl jspl_w_n17483_0(.douta(w_n17483_0[0]),.doutb(w_n17483_0[1]),.din(n17483));
	jspl jspl_w_n17485_0(.douta(w_n17485_0[0]),.doutb(w_n17485_0[1]),.din(n17485));
	jspl jspl_w_n17491_0(.douta(w_n17491_0[0]),.doutb(w_n17491_0[1]),.din(n17491));
	jspl jspl_w_n17493_0(.douta(w_n17493_0[0]),.doutb(w_n17493_0[1]),.din(n17493));
	jspl3 jspl3_w_n17494_0(.douta(w_n17494_0[0]),.doutb(w_n17494_0[1]),.doutc(w_n17494_0[2]),.din(n17494));
	jspl jspl_w_n17497_0(.douta(w_n17497_0[0]),.doutb(w_n17497_0[1]),.din(n17497));
	jspl jspl_w_n17498_0(.douta(w_n17498_0[0]),.doutb(w_n17498_0[1]),.din(n17498));
	jspl3 jspl3_w_n17499_0(.douta(w_n17499_0[0]),.doutb(w_n17499_0[1]),.doutc(w_n17499_0[2]),.din(n17499));
	jspl jspl_w_n17501_0(.douta(w_n17501_0[0]),.doutb(w_n17501_0[1]),.din(n17501));
	jspl jspl_w_n17505_0(.douta(w_n17505_0[0]),.doutb(w_n17505_0[1]),.din(n17505));
	jspl jspl_w_n17507_0(.douta(w_n17507_0[0]),.doutb(w_n17507_0[1]),.din(n17507));
	jspl jspl_w_n17508_0(.douta(w_n17508_0[0]),.doutb(w_n17508_0[1]),.din(n17508));
	jspl3 jspl3_w_n17509_0(.douta(w_n17509_0[0]),.doutb(w_n17509_0[1]),.doutc(w_n17509_0[2]),.din(n17509));
	jspl jspl_w_n17510_0(.douta(w_n17510_0[0]),.doutb(w_n17510_0[1]),.din(n17510));
	jspl jspl_w_n17513_0(.douta(w_n17513_0[0]),.doutb(w_n17513_0[1]),.din(n17513));
	jspl jspl_w_n17519_0(.douta(w_n17519_0[0]),.doutb(w_n17519_0[1]),.din(n17519));
	jspl jspl_w_n17520_0(.douta(w_n17520_0[0]),.doutb(w_n17520_0[1]),.din(n17520));
	jspl jspl_w_n17522_0(.douta(w_n17522_0[0]),.doutb(w_n17522_0[1]),.din(n17522));
	jspl jspl_w_n17524_0(.douta(w_n17524_0[0]),.doutb(w_n17524_0[1]),.din(n17524));
	jspl jspl_w_n17526_0(.douta(w_n17526_0[0]),.doutb(w_n17526_0[1]),.din(n17526));
	jspl jspl_w_n17532_0(.douta(w_n17532_0[0]),.doutb(w_n17532_0[1]),.din(n17532));
	jspl jspl_w_n17534_0(.douta(w_n17534_0[0]),.doutb(w_n17534_0[1]),.din(n17534));
	jspl3 jspl3_w_n17535_0(.douta(w_n17535_0[0]),.doutb(w_n17535_0[1]),.doutc(w_n17535_0[2]),.din(n17535));
	jspl jspl_w_n17538_0(.douta(w_n17538_0[0]),.doutb(w_n17538_0[1]),.din(n17538));
	jspl jspl_w_n17539_0(.douta(w_n17539_0[0]),.doutb(w_n17539_0[1]),.din(n17539));
	jspl3 jspl3_w_n17540_0(.douta(w_n17540_0[0]),.doutb(w_n17540_0[1]),.doutc(w_n17540_0[2]),.din(n17540));
	jspl jspl_w_n17542_0(.douta(w_n17542_0[0]),.doutb(w_n17542_0[1]),.din(n17542));
	jspl jspl_w_n17546_0(.douta(w_n17546_0[0]),.doutb(w_n17546_0[1]),.din(n17546));
	jspl jspl_w_n17548_0(.douta(w_n17548_0[0]),.doutb(w_n17548_0[1]),.din(n17548));
	jspl jspl_w_n17549_0(.douta(w_n17549_0[0]),.doutb(w_n17549_0[1]),.din(n17549));
	jspl3 jspl3_w_n17550_0(.douta(w_n17550_0[0]),.doutb(w_n17550_0[1]),.doutc(w_n17550_0[2]),.din(n17550));
	jspl jspl_w_n17551_0(.douta(w_n17551_0[0]),.doutb(w_n17551_0[1]),.din(n17551));
	jspl jspl_w_n17554_0(.douta(w_n17554_0[0]),.doutb(w_n17554_0[1]),.din(n17554));
	jspl jspl_w_n17560_0(.douta(w_n17560_0[0]),.doutb(w_n17560_0[1]),.din(n17560));
	jspl jspl_w_n17561_0(.douta(w_n17561_0[0]),.doutb(w_n17561_0[1]),.din(n17561));
	jspl jspl_w_n17563_0(.douta(w_n17563_0[0]),.doutb(w_n17563_0[1]),.din(n17563));
	jspl jspl_w_n17565_0(.douta(w_n17565_0[0]),.doutb(w_n17565_0[1]),.din(n17565));
	jspl jspl_w_n17567_0(.douta(w_n17567_0[0]),.doutb(w_n17567_0[1]),.din(n17567));
	jspl jspl_w_n17573_0(.douta(w_n17573_0[0]),.doutb(w_n17573_0[1]),.din(n17573));
	jspl jspl_w_n17575_0(.douta(w_n17575_0[0]),.doutb(w_n17575_0[1]),.din(n17575));
	jspl3 jspl3_w_n17576_0(.douta(w_n17576_0[0]),.doutb(w_n17576_0[1]),.doutc(w_n17576_0[2]),.din(n17576));
	jspl jspl_w_n17579_0(.douta(w_n17579_0[0]),.doutb(w_n17579_0[1]),.din(n17579));
	jspl jspl_w_n17580_0(.douta(w_n17580_0[0]),.doutb(w_n17580_0[1]),.din(n17580));
	jspl3 jspl3_w_n17581_0(.douta(w_n17581_0[0]),.doutb(w_n17581_0[1]),.doutc(w_n17581_0[2]),.din(n17581));
	jspl jspl_w_n17583_0(.douta(w_n17583_0[0]),.doutb(w_n17583_0[1]),.din(n17583));
	jspl jspl_w_n17587_0(.douta(w_n17587_0[0]),.doutb(w_n17587_0[1]),.din(n17587));
	jspl jspl_w_n17589_0(.douta(w_n17589_0[0]),.doutb(w_n17589_0[1]),.din(n17589));
	jspl jspl_w_n17590_0(.douta(w_n17590_0[0]),.doutb(w_n17590_0[1]),.din(n17590));
	jspl3 jspl3_w_n17591_0(.douta(w_n17591_0[0]),.doutb(w_n17591_0[1]),.doutc(w_n17591_0[2]),.din(n17591));
	jspl jspl_w_n17592_0(.douta(w_n17592_0[0]),.doutb(w_n17592_0[1]),.din(n17592));
	jspl jspl_w_n17595_0(.douta(w_n17595_0[0]),.doutb(w_n17595_0[1]),.din(n17595));
	jspl jspl_w_n17601_0(.douta(w_n17601_0[0]),.doutb(w_n17601_0[1]),.din(n17601));
	jspl jspl_w_n17602_0(.douta(w_n17602_0[0]),.doutb(w_n17602_0[1]),.din(n17602));
	jspl jspl_w_n17604_0(.douta(w_n17604_0[0]),.doutb(w_n17604_0[1]),.din(n17604));
	jspl jspl_w_n17606_0(.douta(w_n17606_0[0]),.doutb(w_n17606_0[1]),.din(n17606));
	jspl jspl_w_n17608_0(.douta(w_n17608_0[0]),.doutb(w_n17608_0[1]),.din(n17608));
	jspl jspl_w_n17614_0(.douta(w_n17614_0[0]),.doutb(w_n17614_0[1]),.din(n17614));
	jspl jspl_w_n17616_0(.douta(w_n17616_0[0]),.doutb(w_n17616_0[1]),.din(n17616));
	jspl3 jspl3_w_n17617_0(.douta(w_n17617_0[0]),.doutb(w_n17617_0[1]),.doutc(w_n17617_0[2]),.din(n17617));
	jspl jspl_w_n17620_0(.douta(w_n17620_0[0]),.doutb(w_n17620_0[1]),.din(n17620));
	jspl jspl_w_n17621_0(.douta(w_n17621_0[0]),.doutb(w_n17621_0[1]),.din(n17621));
	jspl3 jspl3_w_n17622_0(.douta(w_n17622_0[0]),.doutb(w_n17622_0[1]),.doutc(w_n17622_0[2]),.din(n17622));
	jspl jspl_w_n17624_0(.douta(w_n17624_0[0]),.doutb(w_n17624_0[1]),.din(n17624));
	jspl jspl_w_n17626_0(.douta(w_n17626_0[0]),.doutb(w_n17626_0[1]),.din(n17626));
	jspl jspl_w_n17628_0(.douta(w_n17628_0[0]),.doutb(w_n17628_0[1]),.din(n17628));
	jspl jspl_w_n17634_0(.douta(w_n17634_0[0]),.doutb(w_n17634_0[1]),.din(n17634));
	jspl3 jspl3_w_n17636_0(.douta(w_n17636_0[0]),.doutb(w_n17636_0[1]),.doutc(w_n17636_0[2]),.din(n17636));
	jspl jspl_w_n17637_0(.douta(w_n17637_0[0]),.doutb(w_n17637_0[1]),.din(n17637));
	jspl jspl_w_n17639_0(.douta(w_n17639_0[0]),.doutb(w_n17639_0[1]),.din(n17639));
	jspl jspl_w_n17641_0(.douta(w_n17641_0[0]),.doutb(w_n17641_0[1]),.din(n17641));
	jspl jspl_w_n17645_0(.douta(w_n17645_0[0]),.doutb(w_n17645_0[1]),.din(n17645));
	jspl jspl_w_n17647_0(.douta(w_n17647_0[0]),.doutb(w_n17647_0[1]),.din(n17647));
	jspl jspl_w_n17648_0(.douta(w_n17648_0[0]),.doutb(w_n17648_0[1]),.din(n17648));
	jspl jspl_w_n17649_0(.douta(w_n17649_0[0]),.doutb(w_n17649_0[1]),.din(n17649));
	jspl3 jspl3_w_n17650_0(.douta(w_n17650_0[0]),.doutb(w_n17650_0[1]),.doutc(w_n17650_0[2]),.din(n17650));
	jspl jspl_w_n17653_0(.douta(w_n17653_0[0]),.doutb(w_n17653_0[1]),.din(n17653));
	jspl jspl_w_n17654_0(.douta(w_n17654_0[0]),.doutb(w_n17654_0[1]),.din(n17654));
	jspl3 jspl3_w_n17655_0(.douta(w_n17655_0[0]),.doutb(w_n17655_0[1]),.doutc(w_n17655_0[2]),.din(n17655));
	jspl jspl_w_n17657_0(.douta(w_n17657_0[0]),.doutb(w_n17657_0[1]),.din(n17657));
	jspl jspl_w_n17661_0(.douta(w_n17661_0[0]),.doutb(w_n17661_0[1]),.din(n17661));
	jspl jspl_w_n17663_0(.douta(w_n17663_0[0]),.doutb(w_n17663_0[1]),.din(n17663));
	jspl jspl_w_n17664_0(.douta(w_n17664_0[0]),.doutb(w_n17664_0[1]),.din(n17664));
	jspl3 jspl3_w_n17665_0(.douta(w_n17665_0[0]),.doutb(w_n17665_0[1]),.doutc(w_n17665_0[2]),.din(n17665));
	jspl jspl_w_n17666_0(.douta(w_n17666_0[0]),.doutb(w_n17666_0[1]),.din(n17666));
	jspl jspl_w_n17669_0(.douta(w_n17669_0[0]),.doutb(w_n17669_0[1]),.din(n17669));
	jspl jspl_w_n17675_0(.douta(w_n17675_0[0]),.doutb(w_n17675_0[1]),.din(n17675));
	jspl jspl_w_n17676_0(.douta(w_n17676_0[0]),.doutb(w_n17676_0[1]),.din(n17676));
	jspl jspl_w_n17678_0(.douta(w_n17678_0[0]),.doutb(w_n17678_0[1]),.din(n17678));
	jspl jspl_w_n17680_0(.douta(w_n17680_0[0]),.doutb(w_n17680_0[1]),.din(n17680));
	jspl jspl_w_n17682_0(.douta(w_n17682_0[0]),.doutb(w_n17682_0[1]),.din(n17682));
	jspl jspl_w_n17688_0(.douta(w_n17688_0[0]),.doutb(w_n17688_0[1]),.din(n17688));
	jspl3 jspl3_w_n17690_0(.douta(w_n17690_0[0]),.doutb(w_n17690_0[1]),.doutc(w_n17690_0[2]),.din(n17690));
	jspl jspl_w_n17695_0(.douta(w_n17695_0[0]),.doutb(w_n17695_0[1]),.din(n17695));
	jspl3 jspl3_w_n17697_0(.douta(w_n17697_0[0]),.doutb(w_n17697_0[1]),.doutc(w_n17697_0[2]),.din(n17697));
	jspl3 jspl3_w_n17701_0(.douta(w_n17701_0[0]),.doutb(w_n17701_0[1]),.doutc(w_n17701_0[2]),.din(n17701));
	jspl jspl_w_n17702_0(.douta(w_n17702_0[0]),.doutb(w_n17702_0[1]),.din(n17702));
	jspl jspl_w_n17707_0(.douta(w_n17707_0[0]),.doutb(w_n17707_0[1]),.din(n17707));
	jspl3 jspl3_w_n17708_0(.douta(w_n17708_0[0]),.doutb(w_n17708_0[1]),.doutc(w_n17708_0[2]),.din(n17708));
	jspl jspl_w_n17713_0(.douta(w_n17713_0[0]),.doutb(w_n17713_0[1]),.din(n17713));
	jspl jspl_w_n17720_0(.douta(w_n17720_0[0]),.doutb(w_n17720_0[1]),.din(n17720));
	jspl3 jspl3_w_n17722_0(.douta(w_n17722_0[0]),.doutb(w_n17722_0[1]),.doutc(w_n17722_0[2]),.din(n17722));
	jspl jspl_w_n17722_1(.douta(w_n17722_1[0]),.doutb(w_n17722_1[1]),.din(w_n17722_0[0]));
	jspl jspl_w_n17723_0(.douta(w_n17723_0[0]),.doutb(w_n17723_0[1]),.din(n17723));
	jspl3 jspl3_w_n17726_0(.douta(w_n17726_0[0]),.doutb(w_n17726_0[1]),.doutc(w_n17726_0[2]),.din(n17726));
	jspl jspl_w_n17727_0(.douta(w_n17727_0[0]),.doutb(w_n17727_0[1]),.din(n17727));
	jspl jspl_w_n17728_0(.douta(w_n17728_0[0]),.doutb(w_n17728_0[1]),.din(n17728));
	jspl jspl_w_n17729_0(.douta(w_n17729_0[0]),.doutb(w_n17729_0[1]),.din(n17729));
	jspl jspl_w_n17731_0(.douta(w_n17731_0[0]),.doutb(w_n17731_0[1]),.din(n17731));
	jspl jspl_w_n17733_0(.douta(w_n17733_0[0]),.doutb(w_n17733_0[1]),.din(n17733));
	jspl jspl_w_n17735_0(.douta(w_n17735_0[0]),.doutb(w_n17735_0[1]),.din(n17735));
	jspl jspl_w_n17744_0(.douta(w_n17744_0[0]),.doutb(w_n17744_0[1]),.din(n17744));
	jspl3 jspl3_w_n17746_0(.douta(w_n17746_0[0]),.doutb(w_n17746_0[1]),.doutc(w_n17746_0[2]),.din(n17746));
	jspl jspl_w_n17747_0(.douta(w_n17747_0[0]),.doutb(w_n17747_0[1]),.din(n17747));
	jspl jspl_w_n17751_0(.douta(w_n17751_0[0]),.doutb(w_n17751_0[1]),.din(n17751));
	jspl jspl_w_n17753_0(.douta(w_n17753_0[0]),.doutb(w_n17753_0[1]),.din(n17753));
	jspl jspl_w_n17755_0(.douta(w_n17755_0[0]),.doutb(w_n17755_0[1]),.din(n17755));
	jspl jspl_w_n17760_0(.douta(w_n17760_0[0]),.doutb(w_n17760_0[1]),.din(n17760));
	jspl jspl_w_n17762_0(.douta(w_n17762_0[0]),.doutb(w_n17762_0[1]),.din(n17762));
	jspl jspl_w_n17763_0(.douta(w_n17763_0[0]),.doutb(w_n17763_0[1]),.din(n17763));
	jspl3 jspl3_w_n17764_0(.douta(w_n17764_0[0]),.doutb(w_n17764_0[1]),.doutc(w_n17764_0[2]),.din(n17764));
	jspl jspl_w_n17765_0(.douta(w_n17765_0[0]),.doutb(w_n17765_0[1]),.din(n17765));
	jspl jspl_w_n17770_0(.douta(w_n17770_0[0]),.doutb(w_n17770_0[1]),.din(n17770));
	jspl jspl_w_n17771_0(.douta(w_n17771_0[0]),.doutb(w_n17771_0[1]),.din(n17771));
	jspl jspl_w_n17773_0(.douta(w_n17773_0[0]),.doutb(w_n17773_0[1]),.din(n17773));
	jspl jspl_w_n17775_0(.douta(w_n17775_0[0]),.doutb(w_n17775_0[1]),.din(n17775));
	jspl jspl_w_n17778_0(.douta(w_n17778_0[0]),.doutb(w_n17778_0[1]),.din(n17778));
	jspl jspl_w_n17784_0(.douta(w_n17784_0[0]),.doutb(w_n17784_0[1]),.din(n17784));
	jspl3 jspl3_w_n17786_0(.douta(w_n17786_0[0]),.doutb(w_n17786_0[1]),.doutc(w_n17786_0[2]),.din(n17786));
	jspl jspl_w_n17787_0(.douta(w_n17787_0[0]),.doutb(w_n17787_0[1]),.din(n17787));
	jspl jspl_w_n17791_0(.douta(w_n17791_0[0]),.doutb(w_n17791_0[1]),.din(n17791));
	jspl jspl_w_n17792_0(.douta(w_n17792_0[0]),.doutb(w_n17792_0[1]),.din(n17792));
	jspl jspl_w_n17794_0(.douta(w_n17794_0[0]),.doutb(w_n17794_0[1]),.din(n17794));
	jspl jspl_w_n17799_0(.douta(w_n17799_0[0]),.doutb(w_n17799_0[1]),.din(n17799));
	jspl jspl_w_n17801_0(.douta(w_n17801_0[0]),.doutb(w_n17801_0[1]),.din(n17801));
	jspl jspl_w_n17802_0(.douta(w_n17802_0[0]),.doutb(w_n17802_0[1]),.din(n17802));
	jspl3 jspl3_w_n17803_0(.douta(w_n17803_0[0]),.doutb(w_n17803_0[1]),.doutc(w_n17803_0[2]),.din(n17803));
	jspl jspl_w_n17804_0(.douta(w_n17804_0[0]),.doutb(w_n17804_0[1]),.din(n17804));
	jspl jspl_w_n17808_0(.douta(w_n17808_0[0]),.doutb(w_n17808_0[1]),.din(n17808));
	jspl jspl_w_n17809_0(.douta(w_n17809_0[0]),.doutb(w_n17809_0[1]),.din(n17809));
	jspl jspl_w_n17811_0(.douta(w_n17811_0[0]),.doutb(w_n17811_0[1]),.din(n17811));
	jspl jspl_w_n17813_0(.douta(w_n17813_0[0]),.doutb(w_n17813_0[1]),.din(n17813));
	jspl jspl_w_n17816_0(.douta(w_n17816_0[0]),.doutb(w_n17816_0[1]),.din(n17816));
	jspl jspl_w_n17822_0(.douta(w_n17822_0[0]),.doutb(w_n17822_0[1]),.din(n17822));
	jspl jspl_w_n17824_0(.douta(w_n17824_0[0]),.doutb(w_n17824_0[1]),.din(n17824));
	jspl3 jspl3_w_n17825_0(.douta(w_n17825_0[0]),.doutb(w_n17825_0[1]),.doutc(w_n17825_0[2]),.din(n17825));
	jspl jspl_w_n17829_0(.douta(w_n17829_0[0]),.doutb(w_n17829_0[1]),.din(n17829));
	jspl jspl_w_n17830_0(.douta(w_n17830_0[0]),.doutb(w_n17830_0[1]),.din(n17830));
	jspl3 jspl3_w_n17831_0(.douta(w_n17831_0[0]),.doutb(w_n17831_0[1]),.doutc(w_n17831_0[2]),.din(n17831));
	jspl jspl_w_n17833_0(.douta(w_n17833_0[0]),.doutb(w_n17833_0[1]),.din(n17833));
	jspl jspl_w_n17838_0(.douta(w_n17838_0[0]),.doutb(w_n17838_0[1]),.din(n17838));
	jspl jspl_w_n17840_0(.douta(w_n17840_0[0]),.doutb(w_n17840_0[1]),.din(n17840));
	jspl jspl_w_n17841_0(.douta(w_n17841_0[0]),.doutb(w_n17841_0[1]),.din(n17841));
	jspl3 jspl3_w_n17842_0(.douta(w_n17842_0[0]),.doutb(w_n17842_0[1]),.doutc(w_n17842_0[2]),.din(n17842));
	jspl jspl_w_n17843_0(.douta(w_n17843_0[0]),.doutb(w_n17843_0[1]),.din(n17843));
	jspl jspl_w_n17847_0(.douta(w_n17847_0[0]),.doutb(w_n17847_0[1]),.din(n17847));
	jspl jspl_w_n17853_0(.douta(w_n17853_0[0]),.doutb(w_n17853_0[1]),.din(n17853));
	jspl jspl_w_n17854_0(.douta(w_n17854_0[0]),.doutb(w_n17854_0[1]),.din(n17854));
	jspl jspl_w_n17856_0(.douta(w_n17856_0[0]),.doutb(w_n17856_0[1]),.din(n17856));
	jspl jspl_w_n17858_0(.douta(w_n17858_0[0]),.doutb(w_n17858_0[1]),.din(n17858));
	jspl jspl_w_n17861_0(.douta(w_n17861_0[0]),.doutb(w_n17861_0[1]),.din(n17861));
	jspl jspl_w_n17867_0(.douta(w_n17867_0[0]),.doutb(w_n17867_0[1]),.din(n17867));
	jspl jspl_w_n17869_0(.douta(w_n17869_0[0]),.doutb(w_n17869_0[1]),.din(n17869));
	jspl3 jspl3_w_n17870_0(.douta(w_n17870_0[0]),.doutb(w_n17870_0[1]),.doutc(w_n17870_0[2]),.din(n17870));
	jspl jspl_w_n17874_0(.douta(w_n17874_0[0]),.doutb(w_n17874_0[1]),.din(n17874));
	jspl jspl_w_n17875_0(.douta(w_n17875_0[0]),.doutb(w_n17875_0[1]),.din(n17875));
	jspl3 jspl3_w_n17876_0(.douta(w_n17876_0[0]),.doutb(w_n17876_0[1]),.doutc(w_n17876_0[2]),.din(n17876));
	jspl jspl_w_n17878_0(.douta(w_n17878_0[0]),.doutb(w_n17878_0[1]),.din(n17878));
	jspl jspl_w_n17883_0(.douta(w_n17883_0[0]),.doutb(w_n17883_0[1]),.din(n17883));
	jspl jspl_w_n17885_0(.douta(w_n17885_0[0]),.doutb(w_n17885_0[1]),.din(n17885));
	jspl jspl_w_n17886_0(.douta(w_n17886_0[0]),.doutb(w_n17886_0[1]),.din(n17886));
	jspl3 jspl3_w_n17887_0(.douta(w_n17887_0[0]),.doutb(w_n17887_0[1]),.doutc(w_n17887_0[2]),.din(n17887));
	jspl jspl_w_n17888_0(.douta(w_n17888_0[0]),.doutb(w_n17888_0[1]),.din(n17888));
	jspl jspl_w_n17892_0(.douta(w_n17892_0[0]),.doutb(w_n17892_0[1]),.din(n17892));
	jspl jspl_w_n17898_0(.douta(w_n17898_0[0]),.doutb(w_n17898_0[1]),.din(n17898));
	jspl jspl_w_n17899_0(.douta(w_n17899_0[0]),.doutb(w_n17899_0[1]),.din(n17899));
	jspl jspl_w_n17901_0(.douta(w_n17901_0[0]),.doutb(w_n17901_0[1]),.din(n17901));
	jspl jspl_w_n17903_0(.douta(w_n17903_0[0]),.doutb(w_n17903_0[1]),.din(n17903));
	jspl jspl_w_n17906_0(.douta(w_n17906_0[0]),.doutb(w_n17906_0[1]),.din(n17906));
	jspl jspl_w_n17912_0(.douta(w_n17912_0[0]),.doutb(w_n17912_0[1]),.din(n17912));
	jspl jspl_w_n17914_0(.douta(w_n17914_0[0]),.doutb(w_n17914_0[1]),.din(n17914));
	jspl3 jspl3_w_n17915_0(.douta(w_n17915_0[0]),.doutb(w_n17915_0[1]),.doutc(w_n17915_0[2]),.din(n17915));
	jspl jspl_w_n17919_0(.douta(w_n17919_0[0]),.doutb(w_n17919_0[1]),.din(n17919));
	jspl jspl_w_n17920_0(.douta(w_n17920_0[0]),.doutb(w_n17920_0[1]),.din(n17920));
	jspl3 jspl3_w_n17921_0(.douta(w_n17921_0[0]),.doutb(w_n17921_0[1]),.doutc(w_n17921_0[2]),.din(n17921));
	jspl jspl_w_n17923_0(.douta(w_n17923_0[0]),.doutb(w_n17923_0[1]),.din(n17923));
	jspl jspl_w_n17928_0(.douta(w_n17928_0[0]),.doutb(w_n17928_0[1]),.din(n17928));
	jspl jspl_w_n17930_0(.douta(w_n17930_0[0]),.doutb(w_n17930_0[1]),.din(n17930));
	jspl jspl_w_n17931_0(.douta(w_n17931_0[0]),.doutb(w_n17931_0[1]),.din(n17931));
	jspl3 jspl3_w_n17932_0(.douta(w_n17932_0[0]),.doutb(w_n17932_0[1]),.doutc(w_n17932_0[2]),.din(n17932));
	jspl jspl_w_n17933_0(.douta(w_n17933_0[0]),.doutb(w_n17933_0[1]),.din(n17933));
	jspl jspl_w_n17937_0(.douta(w_n17937_0[0]),.doutb(w_n17937_0[1]),.din(n17937));
	jspl jspl_w_n17943_0(.douta(w_n17943_0[0]),.doutb(w_n17943_0[1]),.din(n17943));
	jspl jspl_w_n17944_0(.douta(w_n17944_0[0]),.doutb(w_n17944_0[1]),.din(n17944));
	jspl jspl_w_n17946_0(.douta(w_n17946_0[0]),.doutb(w_n17946_0[1]),.din(n17946));
	jspl jspl_w_n17948_0(.douta(w_n17948_0[0]),.doutb(w_n17948_0[1]),.din(n17948));
	jspl jspl_w_n17951_0(.douta(w_n17951_0[0]),.doutb(w_n17951_0[1]),.din(n17951));
	jspl jspl_w_n17957_0(.douta(w_n17957_0[0]),.doutb(w_n17957_0[1]),.din(n17957));
	jspl jspl_w_n17959_0(.douta(w_n17959_0[0]),.doutb(w_n17959_0[1]),.din(n17959));
	jspl3 jspl3_w_n17960_0(.douta(w_n17960_0[0]),.doutb(w_n17960_0[1]),.doutc(w_n17960_0[2]),.din(n17960));
	jspl jspl_w_n17964_0(.douta(w_n17964_0[0]),.doutb(w_n17964_0[1]),.din(n17964));
	jspl jspl_w_n17965_0(.douta(w_n17965_0[0]),.doutb(w_n17965_0[1]),.din(n17965));
	jspl3 jspl3_w_n17966_0(.douta(w_n17966_0[0]),.doutb(w_n17966_0[1]),.doutc(w_n17966_0[2]),.din(n17966));
	jspl jspl_w_n17968_0(.douta(w_n17968_0[0]),.doutb(w_n17968_0[1]),.din(n17968));
	jspl jspl_w_n17973_0(.douta(w_n17973_0[0]),.doutb(w_n17973_0[1]),.din(n17973));
	jspl jspl_w_n17975_0(.douta(w_n17975_0[0]),.doutb(w_n17975_0[1]),.din(n17975));
	jspl jspl_w_n17976_0(.douta(w_n17976_0[0]),.doutb(w_n17976_0[1]),.din(n17976));
	jspl3 jspl3_w_n17977_0(.douta(w_n17977_0[0]),.doutb(w_n17977_0[1]),.doutc(w_n17977_0[2]),.din(n17977));
	jspl jspl_w_n17978_0(.douta(w_n17978_0[0]),.doutb(w_n17978_0[1]),.din(n17978));
	jspl jspl_w_n17982_0(.douta(w_n17982_0[0]),.doutb(w_n17982_0[1]),.din(n17982));
	jspl jspl_w_n17988_0(.douta(w_n17988_0[0]),.doutb(w_n17988_0[1]),.din(n17988));
	jspl jspl_w_n17989_0(.douta(w_n17989_0[0]),.doutb(w_n17989_0[1]),.din(n17989));
	jspl jspl_w_n17991_0(.douta(w_n17991_0[0]),.doutb(w_n17991_0[1]),.din(n17991));
	jspl jspl_w_n17993_0(.douta(w_n17993_0[0]),.doutb(w_n17993_0[1]),.din(n17993));
	jspl jspl_w_n17996_0(.douta(w_n17996_0[0]),.doutb(w_n17996_0[1]),.din(n17996));
	jspl jspl_w_n18002_0(.douta(w_n18002_0[0]),.doutb(w_n18002_0[1]),.din(n18002));
	jspl jspl_w_n18004_0(.douta(w_n18004_0[0]),.doutb(w_n18004_0[1]),.din(n18004));
	jspl3 jspl3_w_n18005_0(.douta(w_n18005_0[0]),.doutb(w_n18005_0[1]),.doutc(w_n18005_0[2]),.din(n18005));
	jspl jspl_w_n18009_0(.douta(w_n18009_0[0]),.doutb(w_n18009_0[1]),.din(n18009));
	jspl jspl_w_n18010_0(.douta(w_n18010_0[0]),.doutb(w_n18010_0[1]),.din(n18010));
	jspl3 jspl3_w_n18011_0(.douta(w_n18011_0[0]),.doutb(w_n18011_0[1]),.doutc(w_n18011_0[2]),.din(n18011));
	jspl jspl_w_n18013_0(.douta(w_n18013_0[0]),.doutb(w_n18013_0[1]),.din(n18013));
	jspl jspl_w_n18018_0(.douta(w_n18018_0[0]),.doutb(w_n18018_0[1]),.din(n18018));
	jspl jspl_w_n18020_0(.douta(w_n18020_0[0]),.doutb(w_n18020_0[1]),.din(n18020));
	jspl jspl_w_n18021_0(.douta(w_n18021_0[0]),.doutb(w_n18021_0[1]),.din(n18021));
	jspl3 jspl3_w_n18022_0(.douta(w_n18022_0[0]),.doutb(w_n18022_0[1]),.doutc(w_n18022_0[2]),.din(n18022));
	jspl jspl_w_n18023_0(.douta(w_n18023_0[0]),.doutb(w_n18023_0[1]),.din(n18023));
	jspl jspl_w_n18027_0(.douta(w_n18027_0[0]),.doutb(w_n18027_0[1]),.din(n18027));
	jspl jspl_w_n18033_0(.douta(w_n18033_0[0]),.doutb(w_n18033_0[1]),.din(n18033));
	jspl jspl_w_n18034_0(.douta(w_n18034_0[0]),.doutb(w_n18034_0[1]),.din(n18034));
	jspl jspl_w_n18036_0(.douta(w_n18036_0[0]),.doutb(w_n18036_0[1]),.din(n18036));
	jspl jspl_w_n18038_0(.douta(w_n18038_0[0]),.doutb(w_n18038_0[1]),.din(n18038));
	jspl jspl_w_n18041_0(.douta(w_n18041_0[0]),.doutb(w_n18041_0[1]),.din(n18041));
	jspl jspl_w_n18047_0(.douta(w_n18047_0[0]),.doutb(w_n18047_0[1]),.din(n18047));
	jspl jspl_w_n18049_0(.douta(w_n18049_0[0]),.doutb(w_n18049_0[1]),.din(n18049));
	jspl3 jspl3_w_n18050_0(.douta(w_n18050_0[0]),.doutb(w_n18050_0[1]),.doutc(w_n18050_0[2]),.din(n18050));
	jspl jspl_w_n18054_0(.douta(w_n18054_0[0]),.doutb(w_n18054_0[1]),.din(n18054));
	jspl jspl_w_n18055_0(.douta(w_n18055_0[0]),.doutb(w_n18055_0[1]),.din(n18055));
	jspl3 jspl3_w_n18056_0(.douta(w_n18056_0[0]),.doutb(w_n18056_0[1]),.doutc(w_n18056_0[2]),.din(n18056));
	jspl jspl_w_n18058_0(.douta(w_n18058_0[0]),.doutb(w_n18058_0[1]),.din(n18058));
	jspl jspl_w_n18063_0(.douta(w_n18063_0[0]),.doutb(w_n18063_0[1]),.din(n18063));
	jspl jspl_w_n18065_0(.douta(w_n18065_0[0]),.doutb(w_n18065_0[1]),.din(n18065));
	jspl jspl_w_n18066_0(.douta(w_n18066_0[0]),.doutb(w_n18066_0[1]),.din(n18066));
	jspl3 jspl3_w_n18067_0(.douta(w_n18067_0[0]),.doutb(w_n18067_0[1]),.doutc(w_n18067_0[2]),.din(n18067));
	jspl jspl_w_n18068_0(.douta(w_n18068_0[0]),.doutb(w_n18068_0[1]),.din(n18068));
	jspl jspl_w_n18072_0(.douta(w_n18072_0[0]),.doutb(w_n18072_0[1]),.din(n18072));
	jspl jspl_w_n18078_0(.douta(w_n18078_0[0]),.doutb(w_n18078_0[1]),.din(n18078));
	jspl jspl_w_n18079_0(.douta(w_n18079_0[0]),.doutb(w_n18079_0[1]),.din(n18079));
	jspl jspl_w_n18081_0(.douta(w_n18081_0[0]),.doutb(w_n18081_0[1]),.din(n18081));
	jspl jspl_w_n18083_0(.douta(w_n18083_0[0]),.doutb(w_n18083_0[1]),.din(n18083));
	jspl jspl_w_n18086_0(.douta(w_n18086_0[0]),.doutb(w_n18086_0[1]),.din(n18086));
	jspl jspl_w_n18092_0(.douta(w_n18092_0[0]),.doutb(w_n18092_0[1]),.din(n18092));
	jspl jspl_w_n18094_0(.douta(w_n18094_0[0]),.doutb(w_n18094_0[1]),.din(n18094));
	jspl3 jspl3_w_n18095_0(.douta(w_n18095_0[0]),.doutb(w_n18095_0[1]),.doutc(w_n18095_0[2]),.din(n18095));
	jspl jspl_w_n18099_0(.douta(w_n18099_0[0]),.doutb(w_n18099_0[1]),.din(n18099));
	jspl jspl_w_n18100_0(.douta(w_n18100_0[0]),.doutb(w_n18100_0[1]),.din(n18100));
	jspl3 jspl3_w_n18101_0(.douta(w_n18101_0[0]),.doutb(w_n18101_0[1]),.doutc(w_n18101_0[2]),.din(n18101));
	jspl jspl_w_n18103_0(.douta(w_n18103_0[0]),.doutb(w_n18103_0[1]),.din(n18103));
	jspl jspl_w_n18108_0(.douta(w_n18108_0[0]),.doutb(w_n18108_0[1]),.din(n18108));
	jspl jspl_w_n18110_0(.douta(w_n18110_0[0]),.doutb(w_n18110_0[1]),.din(n18110));
	jspl jspl_w_n18111_0(.douta(w_n18111_0[0]),.doutb(w_n18111_0[1]),.din(n18111));
	jspl3 jspl3_w_n18112_0(.douta(w_n18112_0[0]),.doutb(w_n18112_0[1]),.doutc(w_n18112_0[2]),.din(n18112));
	jspl jspl_w_n18113_0(.douta(w_n18113_0[0]),.doutb(w_n18113_0[1]),.din(n18113));
	jspl jspl_w_n18117_0(.douta(w_n18117_0[0]),.doutb(w_n18117_0[1]),.din(n18117));
	jspl jspl_w_n18123_0(.douta(w_n18123_0[0]),.doutb(w_n18123_0[1]),.din(n18123));
	jspl jspl_w_n18124_0(.douta(w_n18124_0[0]),.doutb(w_n18124_0[1]),.din(n18124));
	jspl jspl_w_n18126_0(.douta(w_n18126_0[0]),.doutb(w_n18126_0[1]),.din(n18126));
	jspl jspl_w_n18128_0(.douta(w_n18128_0[0]),.doutb(w_n18128_0[1]),.din(n18128));
	jspl jspl_w_n18131_0(.douta(w_n18131_0[0]),.doutb(w_n18131_0[1]),.din(n18131));
	jspl jspl_w_n18137_0(.douta(w_n18137_0[0]),.doutb(w_n18137_0[1]),.din(n18137));
	jspl jspl_w_n18139_0(.douta(w_n18139_0[0]),.doutb(w_n18139_0[1]),.din(n18139));
	jspl3 jspl3_w_n18140_0(.douta(w_n18140_0[0]),.doutb(w_n18140_0[1]),.doutc(w_n18140_0[2]),.din(n18140));
	jspl jspl_w_n18144_0(.douta(w_n18144_0[0]),.doutb(w_n18144_0[1]),.din(n18144));
	jspl jspl_w_n18145_0(.douta(w_n18145_0[0]),.doutb(w_n18145_0[1]),.din(n18145));
	jspl3 jspl3_w_n18146_0(.douta(w_n18146_0[0]),.doutb(w_n18146_0[1]),.doutc(w_n18146_0[2]),.din(n18146));
	jspl jspl_w_n18148_0(.douta(w_n18148_0[0]),.doutb(w_n18148_0[1]),.din(n18148));
	jspl jspl_w_n18153_0(.douta(w_n18153_0[0]),.doutb(w_n18153_0[1]),.din(n18153));
	jspl jspl_w_n18155_0(.douta(w_n18155_0[0]),.doutb(w_n18155_0[1]),.din(n18155));
	jspl jspl_w_n18156_0(.douta(w_n18156_0[0]),.doutb(w_n18156_0[1]),.din(n18156));
	jspl3 jspl3_w_n18157_0(.douta(w_n18157_0[0]),.doutb(w_n18157_0[1]),.doutc(w_n18157_0[2]),.din(n18157));
	jspl jspl_w_n18158_0(.douta(w_n18158_0[0]),.doutb(w_n18158_0[1]),.din(n18158));
	jspl jspl_w_n18162_0(.douta(w_n18162_0[0]),.doutb(w_n18162_0[1]),.din(n18162));
	jspl jspl_w_n18168_0(.douta(w_n18168_0[0]),.doutb(w_n18168_0[1]),.din(n18168));
	jspl jspl_w_n18169_0(.douta(w_n18169_0[0]),.doutb(w_n18169_0[1]),.din(n18169));
	jspl jspl_w_n18171_0(.douta(w_n18171_0[0]),.doutb(w_n18171_0[1]),.din(n18171));
	jspl jspl_w_n18173_0(.douta(w_n18173_0[0]),.doutb(w_n18173_0[1]),.din(n18173));
	jspl jspl_w_n18176_0(.douta(w_n18176_0[0]),.doutb(w_n18176_0[1]),.din(n18176));
	jspl jspl_w_n18182_0(.douta(w_n18182_0[0]),.doutb(w_n18182_0[1]),.din(n18182));
	jspl jspl_w_n18184_0(.douta(w_n18184_0[0]),.doutb(w_n18184_0[1]),.din(n18184));
	jspl3 jspl3_w_n18185_0(.douta(w_n18185_0[0]),.doutb(w_n18185_0[1]),.doutc(w_n18185_0[2]),.din(n18185));
	jspl jspl_w_n18189_0(.douta(w_n18189_0[0]),.doutb(w_n18189_0[1]),.din(n18189));
	jspl jspl_w_n18190_0(.douta(w_n18190_0[0]),.doutb(w_n18190_0[1]),.din(n18190));
	jspl3 jspl3_w_n18191_0(.douta(w_n18191_0[0]),.doutb(w_n18191_0[1]),.doutc(w_n18191_0[2]),.din(n18191));
	jspl jspl_w_n18193_0(.douta(w_n18193_0[0]),.doutb(w_n18193_0[1]),.din(n18193));
	jspl jspl_w_n18198_0(.douta(w_n18198_0[0]),.doutb(w_n18198_0[1]),.din(n18198));
	jspl jspl_w_n18200_0(.douta(w_n18200_0[0]),.doutb(w_n18200_0[1]),.din(n18200));
	jspl jspl_w_n18201_0(.douta(w_n18201_0[0]),.doutb(w_n18201_0[1]),.din(n18201));
	jspl3 jspl3_w_n18202_0(.douta(w_n18202_0[0]),.doutb(w_n18202_0[1]),.doutc(w_n18202_0[2]),.din(n18202));
	jspl jspl_w_n18203_0(.douta(w_n18203_0[0]),.doutb(w_n18203_0[1]),.din(n18203));
	jspl jspl_w_n18207_0(.douta(w_n18207_0[0]),.doutb(w_n18207_0[1]),.din(n18207));
	jspl jspl_w_n18213_0(.douta(w_n18213_0[0]),.doutb(w_n18213_0[1]),.din(n18213));
	jspl jspl_w_n18214_0(.douta(w_n18214_0[0]),.doutb(w_n18214_0[1]),.din(n18214));
	jspl jspl_w_n18216_0(.douta(w_n18216_0[0]),.doutb(w_n18216_0[1]),.din(n18216));
	jspl jspl_w_n18218_0(.douta(w_n18218_0[0]),.doutb(w_n18218_0[1]),.din(n18218));
	jspl jspl_w_n18221_0(.douta(w_n18221_0[0]),.doutb(w_n18221_0[1]),.din(n18221));
	jspl jspl_w_n18227_0(.douta(w_n18227_0[0]),.doutb(w_n18227_0[1]),.din(n18227));
	jspl jspl_w_n18229_0(.douta(w_n18229_0[0]),.doutb(w_n18229_0[1]),.din(n18229));
	jspl3 jspl3_w_n18230_0(.douta(w_n18230_0[0]),.doutb(w_n18230_0[1]),.doutc(w_n18230_0[2]),.din(n18230));
	jspl jspl_w_n18234_0(.douta(w_n18234_0[0]),.doutb(w_n18234_0[1]),.din(n18234));
	jspl jspl_w_n18235_0(.douta(w_n18235_0[0]),.doutb(w_n18235_0[1]),.din(n18235));
	jspl3 jspl3_w_n18236_0(.douta(w_n18236_0[0]),.doutb(w_n18236_0[1]),.doutc(w_n18236_0[2]),.din(n18236));
	jspl jspl_w_n18238_0(.douta(w_n18238_0[0]),.doutb(w_n18238_0[1]),.din(n18238));
	jspl jspl_w_n18243_0(.douta(w_n18243_0[0]),.doutb(w_n18243_0[1]),.din(n18243));
	jspl jspl_w_n18245_0(.douta(w_n18245_0[0]),.doutb(w_n18245_0[1]),.din(n18245));
	jspl jspl_w_n18246_0(.douta(w_n18246_0[0]),.doutb(w_n18246_0[1]),.din(n18246));
	jspl3 jspl3_w_n18247_0(.douta(w_n18247_0[0]),.doutb(w_n18247_0[1]),.doutc(w_n18247_0[2]),.din(n18247));
	jspl jspl_w_n18248_0(.douta(w_n18248_0[0]),.doutb(w_n18248_0[1]),.din(n18248));
	jspl jspl_w_n18252_0(.douta(w_n18252_0[0]),.doutb(w_n18252_0[1]),.din(n18252));
	jspl jspl_w_n18258_0(.douta(w_n18258_0[0]),.doutb(w_n18258_0[1]),.din(n18258));
	jspl jspl_w_n18259_0(.douta(w_n18259_0[0]),.doutb(w_n18259_0[1]),.din(n18259));
	jspl jspl_w_n18261_0(.douta(w_n18261_0[0]),.doutb(w_n18261_0[1]),.din(n18261));
	jspl jspl_w_n18266_0(.douta(w_n18266_0[0]),.doutb(w_n18266_0[1]),.din(n18266));
	jspl jspl_w_n18268_0(.douta(w_n18268_0[0]),.doutb(w_n18268_0[1]),.din(n18268));
	jspl jspl_w_n18269_0(.douta(w_n18269_0[0]),.doutb(w_n18269_0[1]),.din(n18269));
	jspl3 jspl3_w_n18270_0(.douta(w_n18270_0[0]),.doutb(w_n18270_0[1]),.doutc(w_n18270_0[2]),.din(n18270));
	jspl jspl_w_n18271_0(.douta(w_n18271_0[0]),.doutb(w_n18271_0[1]),.din(n18271));
	jspl jspl_w_n18274_0(.douta(w_n18274_0[0]),.doutb(w_n18274_0[1]),.din(n18274));
	jspl jspl_w_n18276_0(.douta(w_n18276_0[0]),.doutb(w_n18276_0[1]),.din(n18276));
	jspl jspl_w_n18278_0(.douta(w_n18278_0[0]),.doutb(w_n18278_0[1]),.din(n18278));
	jspl jspl_w_n18281_0(.douta(w_n18281_0[0]),.doutb(w_n18281_0[1]),.din(n18281));
	jspl jspl_w_n18287_0(.douta(w_n18287_0[0]),.doutb(w_n18287_0[1]),.din(n18287));
	jspl3 jspl3_w_n18289_0(.douta(w_n18289_0[0]),.doutb(w_n18289_0[1]),.doutc(w_n18289_0[2]),.din(n18289));
	jspl jspl_w_n18290_0(.douta(w_n18290_0[0]),.doutb(w_n18290_0[1]),.din(n18290));
	jspl jspl_w_n18294_0(.douta(w_n18294_0[0]),.doutb(w_n18294_0[1]),.din(n18294));
	jspl jspl_w_n18300_0(.douta(w_n18300_0[0]),.doutb(w_n18300_0[1]),.din(n18300));
	jspl jspl_w_n18301_0(.douta(w_n18301_0[0]),.doutb(w_n18301_0[1]),.din(n18301));
	jspl jspl_w_n18303_0(.douta(w_n18303_0[0]),.doutb(w_n18303_0[1]),.din(n18303));
	jspl jspl_w_n18305_0(.douta(w_n18305_0[0]),.doutb(w_n18305_0[1]),.din(n18305));
	jspl jspl_w_n18308_0(.douta(w_n18308_0[0]),.doutb(w_n18308_0[1]),.din(n18308));
	jspl jspl_w_n18314_0(.douta(w_n18314_0[0]),.doutb(w_n18314_0[1]),.din(n18314));
	jspl jspl_w_n18316_0(.douta(w_n18316_0[0]),.doutb(w_n18316_0[1]),.din(n18316));
	jspl3 jspl3_w_n18317_0(.douta(w_n18317_0[0]),.doutb(w_n18317_0[1]),.doutc(w_n18317_0[2]),.din(n18317));
	jspl jspl_w_n18321_0(.douta(w_n18321_0[0]),.doutb(w_n18321_0[1]),.din(n18321));
	jspl jspl_w_n18322_0(.douta(w_n18322_0[0]),.doutb(w_n18322_0[1]),.din(n18322));
	jspl3 jspl3_w_n18323_0(.douta(w_n18323_0[0]),.doutb(w_n18323_0[1]),.doutc(w_n18323_0[2]),.din(n18323));
	jspl jspl_w_n18325_0(.douta(w_n18325_0[0]),.doutb(w_n18325_0[1]),.din(n18325));
	jspl jspl_w_n18330_0(.douta(w_n18330_0[0]),.doutb(w_n18330_0[1]),.din(n18330));
	jspl jspl_w_n18332_0(.douta(w_n18332_0[0]),.doutb(w_n18332_0[1]),.din(n18332));
	jspl jspl_w_n18333_0(.douta(w_n18333_0[0]),.doutb(w_n18333_0[1]),.din(n18333));
	jspl3 jspl3_w_n18334_0(.douta(w_n18334_0[0]),.doutb(w_n18334_0[1]),.doutc(w_n18334_0[2]),.din(n18334));
	jspl3 jspl3_w_n18334_1(.douta(w_n18334_1[0]),.doutb(w_n18334_1[1]),.doutc(w_n18334_1[2]),.din(w_n18334_0[0]));
	jspl jspl_w_n18337_0(.douta(w_n18337_0[0]),.doutb(w_n18337_0[1]),.din(n18337));
	jspl3 jspl3_w_n18338_0(.douta(w_n18338_0[0]),.doutb(w_n18338_0[1]),.doutc(w_n18338_0[2]),.din(n18338));
	jspl jspl_w_n18339_0(.douta(w_n18339_0[0]),.doutb(w_n18339_0[1]),.din(n18339));
	jspl jspl_w_n18340_0(.douta(w_n18340_0[0]),.doutb(w_n18340_0[1]),.din(n18340));
	jspl3 jspl3_w_n18347_0(.douta(w_n18347_0[0]),.doutb(w_n18347_0[1]),.doutc(w_n18347_0[2]),.din(n18347));
	jspl jspl_w_n18348_0(.douta(w_n18348_0[0]),.doutb(w_n18348_0[1]),.din(n18348));
	jspl3 jspl3_w_n18356_0(.douta(w_n18356_0[0]),.doutb(w_n18356_0[1]),.doutc(w_n18356_0[2]),.din(n18356));
	jspl3 jspl3_w_n18356_1(.douta(w_n18356_1[0]),.doutb(w_n18356_1[1]),.doutc(w_n18356_1[2]),.din(w_n18356_0[0]));
	jspl3 jspl3_w_n18356_2(.douta(w_n18356_2[0]),.doutb(w_n18356_2[1]),.doutc(w_n18356_2[2]),.din(w_n18356_0[1]));
	jspl3 jspl3_w_n18356_3(.douta(w_n18356_3[0]),.doutb(w_n18356_3[1]),.doutc(w_n18356_3[2]),.din(w_n18356_0[2]));
	jspl3 jspl3_w_n18356_4(.douta(w_n18356_4[0]),.doutb(w_n18356_4[1]),.doutc(w_n18356_4[2]),.din(w_n18356_1[0]));
	jspl3 jspl3_w_n18356_5(.douta(w_n18356_5[0]),.doutb(w_n18356_5[1]),.doutc(w_n18356_5[2]),.din(w_n18356_1[1]));
	jspl3 jspl3_w_n18356_6(.douta(w_n18356_6[0]),.doutb(w_n18356_6[1]),.doutc(w_n18356_6[2]),.din(w_n18356_1[2]));
	jspl3 jspl3_w_n18356_7(.douta(w_n18356_7[0]),.doutb(w_n18356_7[1]),.doutc(w_n18356_7[2]),.din(w_n18356_2[0]));
	jspl3 jspl3_w_n18356_8(.douta(w_n18356_8[0]),.doutb(w_n18356_8[1]),.doutc(w_n18356_8[2]),.din(w_n18356_2[1]));
	jspl3 jspl3_w_n18356_9(.douta(w_n18356_9[0]),.doutb(w_n18356_9[1]),.doutc(w_n18356_9[2]),.din(w_n18356_2[2]));
	jspl3 jspl3_w_n18356_10(.douta(w_n18356_10[0]),.doutb(w_n18356_10[1]),.doutc(w_n18356_10[2]),.din(w_n18356_3[0]));
	jspl3 jspl3_w_n18356_11(.douta(w_n18356_11[0]),.doutb(w_n18356_11[1]),.doutc(w_n18356_11[2]),.din(w_n18356_3[1]));
	jspl3 jspl3_w_n18356_12(.douta(w_n18356_12[0]),.doutb(w_n18356_12[1]),.doutc(w_n18356_12[2]),.din(w_n18356_3[2]));
	jspl3 jspl3_w_n18356_13(.douta(w_n18356_13[0]),.doutb(w_n18356_13[1]),.doutc(w_n18356_13[2]),.din(w_n18356_4[0]));
	jspl3 jspl3_w_n18356_14(.douta(w_n18356_14[0]),.doutb(w_n18356_14[1]),.doutc(w_n18356_14[2]),.din(w_n18356_4[1]));
	jspl3 jspl3_w_n18356_15(.douta(w_n18356_15[0]),.doutb(w_n18356_15[1]),.doutc(w_n18356_15[2]),.din(w_n18356_4[2]));
	jspl3 jspl3_w_n18356_16(.douta(w_n18356_16[0]),.doutb(w_n18356_16[1]),.doutc(w_n18356_16[2]),.din(w_n18356_5[0]));
	jspl3 jspl3_w_n18356_17(.douta(w_n18356_17[0]),.doutb(w_n18356_17[1]),.doutc(w_n18356_17[2]),.din(w_n18356_5[1]));
	jspl3 jspl3_w_n18356_18(.douta(w_n18356_18[0]),.doutb(w_n18356_18[1]),.doutc(w_n18356_18[2]),.din(w_n18356_5[2]));
	jspl jspl_w_n18356_19(.douta(w_n18356_19[0]),.doutb(w_n18356_19[1]),.din(w_n18356_6[0]));
	jspl jspl_w_n18359_0(.douta(w_n18359_0[0]),.doutb(w_n18359_0[1]),.din(n18359));
	jspl3 jspl3_w_n18360_0(.douta(w_n18360_0[0]),.doutb(w_n18360_0[1]),.doutc(w_n18360_0[2]),.din(n18360));
	jspl3 jspl3_w_n18360_1(.douta(w_n18360_1[0]),.doutb(w_n18360_1[1]),.doutc(w_n18360_1[2]),.din(w_n18360_0[0]));
	jspl3 jspl3_w_n18360_2(.douta(w_n18360_2[0]),.doutb(w_n18360_2[1]),.doutc(w_n18360_2[2]),.din(w_n18360_0[1]));
	jspl3 jspl3_w_n18360_3(.douta(w_n18360_3[0]),.doutb(w_n18360_3[1]),.doutc(w_n18360_3[2]),.din(w_n18360_0[2]));
	jspl3 jspl3_w_n18362_0(.douta(w_n18362_0[0]),.doutb(w_n18362_0[1]),.doutc(w_n18362_0[2]),.din(n18362));
	jspl jspl_w_n18362_1(.douta(w_n18362_1[0]),.doutb(w_n18362_1[1]),.din(w_n18362_0[0]));
	jspl3 jspl3_w_n18363_0(.douta(w_n18363_0[0]),.doutb(w_n18363_0[1]),.doutc(w_n18363_0[2]),.din(n18363));
	jspl3 jspl3_w_n18367_0(.douta(w_n18367_0[0]),.doutb(w_n18367_0[1]),.doutc(w_n18367_0[2]),.din(n18367));
	jspl jspl_w_n18368_0(.douta(w_n18368_0[0]),.doutb(w_n18368_0[1]),.din(n18368));
	jspl jspl_w_n18369_0(.douta(w_n18369_0[0]),.doutb(w_n18369_0[1]),.din(n18369));
	jspl jspl_w_n18370_0(.douta(w_n18370_0[0]),.doutb(w_n18370_0[1]),.din(n18370));
	jspl jspl_w_n18372_0(.douta(w_n18372_0[0]),.doutb(w_n18372_0[1]),.din(n18372));
	jspl jspl_w_n18374_0(.douta(w_n18374_0[0]),.doutb(w_n18374_0[1]),.din(n18374));
	jspl jspl_w_n18376_0(.douta(w_n18376_0[0]),.doutb(w_n18376_0[1]),.din(n18376));
	jspl jspl_w_n18381_0(.douta(w_n18381_0[0]),.doutb(w_n18381_0[1]),.din(n18381));
	jspl3 jspl3_w_n18383_0(.douta(w_n18383_0[0]),.doutb(w_n18383_0[1]),.doutc(w_n18383_0[2]),.din(n18383));
	jspl jspl_w_n18384_0(.douta(w_n18384_0[0]),.doutb(w_n18384_0[1]),.din(n18384));
	jspl jspl_w_n18388_0(.douta(w_n18388_0[0]),.doutb(w_n18388_0[1]),.din(n18388));
	jspl jspl_w_n18389_0(.douta(w_n18389_0[0]),.doutb(w_n18389_0[1]),.din(n18389));
	jspl jspl_w_n18391_0(.douta(w_n18391_0[0]),.doutb(w_n18391_0[1]),.din(n18391));
	jspl jspl_w_n18395_0(.douta(w_n18395_0[0]),.doutb(w_n18395_0[1]),.din(n18395));
	jspl jspl_w_n18397_0(.douta(w_n18397_0[0]),.doutb(w_n18397_0[1]),.din(n18397));
	jspl jspl_w_n18398_0(.douta(w_n18398_0[0]),.doutb(w_n18398_0[1]),.din(n18398));
	jspl3 jspl3_w_n18399_0(.douta(w_n18399_0[0]),.doutb(w_n18399_0[1]),.doutc(w_n18399_0[2]),.din(n18399));
	jspl jspl_w_n18400_0(.douta(w_n18400_0[0]),.doutb(w_n18400_0[1]),.din(n18400));
	jspl jspl_w_n18404_0(.douta(w_n18404_0[0]),.doutb(w_n18404_0[1]),.din(n18404));
	jspl jspl_w_n18406_0(.douta(w_n18406_0[0]),.doutb(w_n18406_0[1]),.din(n18406));
	jspl jspl_w_n18408_0(.douta(w_n18408_0[0]),.doutb(w_n18408_0[1]),.din(n18408));
	jspl jspl_w_n18410_0(.douta(w_n18410_0[0]),.doutb(w_n18410_0[1]),.din(n18410));
	jspl jspl_w_n18412_0(.douta(w_n18412_0[0]),.doutb(w_n18412_0[1]),.din(n18412));
	jspl jspl_w_n18418_0(.douta(w_n18418_0[0]),.doutb(w_n18418_0[1]),.din(n18418));
	jspl3 jspl3_w_n18420_0(.douta(w_n18420_0[0]),.doutb(w_n18420_0[1]),.doutc(w_n18420_0[2]),.din(n18420));
	jspl jspl_w_n18421_0(.douta(w_n18421_0[0]),.doutb(w_n18421_0[1]),.din(n18421));
	jspl jspl_w_n18426_0(.douta(w_n18426_0[0]),.doutb(w_n18426_0[1]),.din(n18426));
	jspl jspl_w_n18428_0(.douta(w_n18428_0[0]),.doutb(w_n18428_0[1]),.din(n18428));
	jspl jspl_w_n18430_0(.douta(w_n18430_0[0]),.doutb(w_n18430_0[1]),.din(n18430));
	jspl jspl_w_n18434_0(.douta(w_n18434_0[0]),.doutb(w_n18434_0[1]),.din(n18434));
	jspl jspl_w_n18436_0(.douta(w_n18436_0[0]),.doutb(w_n18436_0[1]),.din(n18436));
	jspl jspl_w_n18437_0(.douta(w_n18437_0[0]),.doutb(w_n18437_0[1]),.din(n18437));
	jspl3 jspl3_w_n18438_0(.douta(w_n18438_0[0]),.doutb(w_n18438_0[1]),.doutc(w_n18438_0[2]),.din(n18438));
	jspl jspl_w_n18439_0(.douta(w_n18439_0[0]),.doutb(w_n18439_0[1]),.din(n18439));
	jspl jspl_w_n18445_0(.douta(w_n18445_0[0]),.doutb(w_n18445_0[1]),.din(n18445));
	jspl jspl_w_n18446_0(.douta(w_n18446_0[0]),.doutb(w_n18446_0[1]),.din(n18446));
	jspl jspl_w_n18448_0(.douta(w_n18448_0[0]),.doutb(w_n18448_0[1]),.din(n18448));
	jspl jspl_w_n18450_0(.douta(w_n18450_0[0]),.doutb(w_n18450_0[1]),.din(n18450));
	jspl jspl_w_n18452_0(.douta(w_n18452_0[0]),.doutb(w_n18452_0[1]),.din(n18452));
	jspl jspl_w_n18458_0(.douta(w_n18458_0[0]),.doutb(w_n18458_0[1]),.din(n18458));
	jspl jspl_w_n18460_0(.douta(w_n18460_0[0]),.doutb(w_n18460_0[1]),.din(n18460));
	jspl3 jspl3_w_n18461_0(.douta(w_n18461_0[0]),.doutb(w_n18461_0[1]),.doutc(w_n18461_0[2]),.din(n18461));
	jspl jspl_w_n18464_0(.douta(w_n18464_0[0]),.doutb(w_n18464_0[1]),.din(n18464));
	jspl jspl_w_n18465_0(.douta(w_n18465_0[0]),.doutb(w_n18465_0[1]),.din(n18465));
	jspl3 jspl3_w_n18466_0(.douta(w_n18466_0[0]),.doutb(w_n18466_0[1]),.doutc(w_n18466_0[2]),.din(n18466));
	jspl jspl_w_n18468_0(.douta(w_n18468_0[0]),.doutb(w_n18468_0[1]),.din(n18468));
	jspl jspl_w_n18472_0(.douta(w_n18472_0[0]),.doutb(w_n18472_0[1]),.din(n18472));
	jspl jspl_w_n18474_0(.douta(w_n18474_0[0]),.doutb(w_n18474_0[1]),.din(n18474));
	jspl jspl_w_n18475_0(.douta(w_n18475_0[0]),.doutb(w_n18475_0[1]),.din(n18475));
	jspl3 jspl3_w_n18476_0(.douta(w_n18476_0[0]),.doutb(w_n18476_0[1]),.doutc(w_n18476_0[2]),.din(n18476));
	jspl jspl_w_n18477_0(.douta(w_n18477_0[0]),.doutb(w_n18477_0[1]),.din(n18477));
	jspl jspl_w_n18480_0(.douta(w_n18480_0[0]),.doutb(w_n18480_0[1]),.din(n18480));
	jspl jspl_w_n18486_0(.douta(w_n18486_0[0]),.doutb(w_n18486_0[1]),.din(n18486));
	jspl jspl_w_n18487_0(.douta(w_n18487_0[0]),.doutb(w_n18487_0[1]),.din(n18487));
	jspl jspl_w_n18489_0(.douta(w_n18489_0[0]),.doutb(w_n18489_0[1]),.din(n18489));
	jspl jspl_w_n18491_0(.douta(w_n18491_0[0]),.doutb(w_n18491_0[1]),.din(n18491));
	jspl jspl_w_n18493_0(.douta(w_n18493_0[0]),.doutb(w_n18493_0[1]),.din(n18493));
	jspl jspl_w_n18499_0(.douta(w_n18499_0[0]),.doutb(w_n18499_0[1]),.din(n18499));
	jspl jspl_w_n18501_0(.douta(w_n18501_0[0]),.doutb(w_n18501_0[1]),.din(n18501));
	jspl3 jspl3_w_n18502_0(.douta(w_n18502_0[0]),.doutb(w_n18502_0[1]),.doutc(w_n18502_0[2]),.din(n18502));
	jspl jspl_w_n18505_0(.douta(w_n18505_0[0]),.doutb(w_n18505_0[1]),.din(n18505));
	jspl jspl_w_n18506_0(.douta(w_n18506_0[0]),.doutb(w_n18506_0[1]),.din(n18506));
	jspl3 jspl3_w_n18507_0(.douta(w_n18507_0[0]),.doutb(w_n18507_0[1]),.doutc(w_n18507_0[2]),.din(n18507));
	jspl jspl_w_n18509_0(.douta(w_n18509_0[0]),.doutb(w_n18509_0[1]),.din(n18509));
	jspl jspl_w_n18513_0(.douta(w_n18513_0[0]),.doutb(w_n18513_0[1]),.din(n18513));
	jspl jspl_w_n18515_0(.douta(w_n18515_0[0]),.doutb(w_n18515_0[1]),.din(n18515));
	jspl jspl_w_n18516_0(.douta(w_n18516_0[0]),.doutb(w_n18516_0[1]),.din(n18516));
	jspl3 jspl3_w_n18517_0(.douta(w_n18517_0[0]),.doutb(w_n18517_0[1]),.doutc(w_n18517_0[2]),.din(n18517));
	jspl jspl_w_n18518_0(.douta(w_n18518_0[0]),.doutb(w_n18518_0[1]),.din(n18518));
	jspl jspl_w_n18521_0(.douta(w_n18521_0[0]),.doutb(w_n18521_0[1]),.din(n18521));
	jspl jspl_w_n18527_0(.douta(w_n18527_0[0]),.doutb(w_n18527_0[1]),.din(n18527));
	jspl jspl_w_n18528_0(.douta(w_n18528_0[0]),.doutb(w_n18528_0[1]),.din(n18528));
	jspl jspl_w_n18530_0(.douta(w_n18530_0[0]),.doutb(w_n18530_0[1]),.din(n18530));
	jspl jspl_w_n18532_0(.douta(w_n18532_0[0]),.doutb(w_n18532_0[1]),.din(n18532));
	jspl jspl_w_n18534_0(.douta(w_n18534_0[0]),.doutb(w_n18534_0[1]),.din(n18534));
	jspl jspl_w_n18540_0(.douta(w_n18540_0[0]),.doutb(w_n18540_0[1]),.din(n18540));
	jspl jspl_w_n18542_0(.douta(w_n18542_0[0]),.doutb(w_n18542_0[1]),.din(n18542));
	jspl3 jspl3_w_n18543_0(.douta(w_n18543_0[0]),.doutb(w_n18543_0[1]),.doutc(w_n18543_0[2]),.din(n18543));
	jspl jspl_w_n18546_0(.douta(w_n18546_0[0]),.doutb(w_n18546_0[1]),.din(n18546));
	jspl jspl_w_n18547_0(.douta(w_n18547_0[0]),.doutb(w_n18547_0[1]),.din(n18547));
	jspl3 jspl3_w_n18548_0(.douta(w_n18548_0[0]),.doutb(w_n18548_0[1]),.doutc(w_n18548_0[2]),.din(n18548));
	jspl jspl_w_n18550_0(.douta(w_n18550_0[0]),.doutb(w_n18550_0[1]),.din(n18550));
	jspl jspl_w_n18554_0(.douta(w_n18554_0[0]),.doutb(w_n18554_0[1]),.din(n18554));
	jspl jspl_w_n18556_0(.douta(w_n18556_0[0]),.doutb(w_n18556_0[1]),.din(n18556));
	jspl jspl_w_n18557_0(.douta(w_n18557_0[0]),.doutb(w_n18557_0[1]),.din(n18557));
	jspl3 jspl3_w_n18558_0(.douta(w_n18558_0[0]),.doutb(w_n18558_0[1]),.doutc(w_n18558_0[2]),.din(n18558));
	jspl jspl_w_n18559_0(.douta(w_n18559_0[0]),.doutb(w_n18559_0[1]),.din(n18559));
	jspl jspl_w_n18562_0(.douta(w_n18562_0[0]),.doutb(w_n18562_0[1]),.din(n18562));
	jspl jspl_w_n18568_0(.douta(w_n18568_0[0]),.doutb(w_n18568_0[1]),.din(n18568));
	jspl jspl_w_n18569_0(.douta(w_n18569_0[0]),.doutb(w_n18569_0[1]),.din(n18569));
	jspl jspl_w_n18571_0(.douta(w_n18571_0[0]),.doutb(w_n18571_0[1]),.din(n18571));
	jspl jspl_w_n18573_0(.douta(w_n18573_0[0]),.doutb(w_n18573_0[1]),.din(n18573));
	jspl jspl_w_n18575_0(.douta(w_n18575_0[0]),.doutb(w_n18575_0[1]),.din(n18575));
	jspl jspl_w_n18581_0(.douta(w_n18581_0[0]),.doutb(w_n18581_0[1]),.din(n18581));
	jspl jspl_w_n18583_0(.douta(w_n18583_0[0]),.doutb(w_n18583_0[1]),.din(n18583));
	jspl3 jspl3_w_n18584_0(.douta(w_n18584_0[0]),.doutb(w_n18584_0[1]),.doutc(w_n18584_0[2]),.din(n18584));
	jspl jspl_w_n18587_0(.douta(w_n18587_0[0]),.doutb(w_n18587_0[1]),.din(n18587));
	jspl jspl_w_n18588_0(.douta(w_n18588_0[0]),.doutb(w_n18588_0[1]),.din(n18588));
	jspl3 jspl3_w_n18589_0(.douta(w_n18589_0[0]),.doutb(w_n18589_0[1]),.doutc(w_n18589_0[2]),.din(n18589));
	jspl jspl_w_n18591_0(.douta(w_n18591_0[0]),.doutb(w_n18591_0[1]),.din(n18591));
	jspl jspl_w_n18595_0(.douta(w_n18595_0[0]),.doutb(w_n18595_0[1]),.din(n18595));
	jspl jspl_w_n18597_0(.douta(w_n18597_0[0]),.doutb(w_n18597_0[1]),.din(n18597));
	jspl jspl_w_n18598_0(.douta(w_n18598_0[0]),.doutb(w_n18598_0[1]),.din(n18598));
	jspl3 jspl3_w_n18599_0(.douta(w_n18599_0[0]),.doutb(w_n18599_0[1]),.doutc(w_n18599_0[2]),.din(n18599));
	jspl jspl_w_n18600_0(.douta(w_n18600_0[0]),.doutb(w_n18600_0[1]),.din(n18600));
	jspl jspl_w_n18603_0(.douta(w_n18603_0[0]),.doutb(w_n18603_0[1]),.din(n18603));
	jspl jspl_w_n18609_0(.douta(w_n18609_0[0]),.doutb(w_n18609_0[1]),.din(n18609));
	jspl jspl_w_n18610_0(.douta(w_n18610_0[0]),.doutb(w_n18610_0[1]),.din(n18610));
	jspl jspl_w_n18612_0(.douta(w_n18612_0[0]),.doutb(w_n18612_0[1]),.din(n18612));
	jspl jspl_w_n18614_0(.douta(w_n18614_0[0]),.doutb(w_n18614_0[1]),.din(n18614));
	jspl jspl_w_n18616_0(.douta(w_n18616_0[0]),.doutb(w_n18616_0[1]),.din(n18616));
	jspl jspl_w_n18622_0(.douta(w_n18622_0[0]),.doutb(w_n18622_0[1]),.din(n18622));
	jspl jspl_w_n18624_0(.douta(w_n18624_0[0]),.doutb(w_n18624_0[1]),.din(n18624));
	jspl3 jspl3_w_n18625_0(.douta(w_n18625_0[0]),.doutb(w_n18625_0[1]),.doutc(w_n18625_0[2]),.din(n18625));
	jspl jspl_w_n18628_0(.douta(w_n18628_0[0]),.doutb(w_n18628_0[1]),.din(n18628));
	jspl jspl_w_n18629_0(.douta(w_n18629_0[0]),.doutb(w_n18629_0[1]),.din(n18629));
	jspl3 jspl3_w_n18630_0(.douta(w_n18630_0[0]),.doutb(w_n18630_0[1]),.doutc(w_n18630_0[2]),.din(n18630));
	jspl jspl_w_n18632_0(.douta(w_n18632_0[0]),.doutb(w_n18632_0[1]),.din(n18632));
	jspl jspl_w_n18636_0(.douta(w_n18636_0[0]),.doutb(w_n18636_0[1]),.din(n18636));
	jspl jspl_w_n18638_0(.douta(w_n18638_0[0]),.doutb(w_n18638_0[1]),.din(n18638));
	jspl jspl_w_n18639_0(.douta(w_n18639_0[0]),.doutb(w_n18639_0[1]),.din(n18639));
	jspl3 jspl3_w_n18640_0(.douta(w_n18640_0[0]),.doutb(w_n18640_0[1]),.doutc(w_n18640_0[2]),.din(n18640));
	jspl jspl_w_n18641_0(.douta(w_n18641_0[0]),.doutb(w_n18641_0[1]),.din(n18641));
	jspl jspl_w_n18644_0(.douta(w_n18644_0[0]),.doutb(w_n18644_0[1]),.din(n18644));
	jspl jspl_w_n18650_0(.douta(w_n18650_0[0]),.doutb(w_n18650_0[1]),.din(n18650));
	jspl jspl_w_n18651_0(.douta(w_n18651_0[0]),.doutb(w_n18651_0[1]),.din(n18651));
	jspl jspl_w_n18653_0(.douta(w_n18653_0[0]),.doutb(w_n18653_0[1]),.din(n18653));
	jspl jspl_w_n18655_0(.douta(w_n18655_0[0]),.doutb(w_n18655_0[1]),.din(n18655));
	jspl jspl_w_n18657_0(.douta(w_n18657_0[0]),.doutb(w_n18657_0[1]),.din(n18657));
	jspl jspl_w_n18663_0(.douta(w_n18663_0[0]),.doutb(w_n18663_0[1]),.din(n18663));
	jspl jspl_w_n18665_0(.douta(w_n18665_0[0]),.doutb(w_n18665_0[1]),.din(n18665));
	jspl3 jspl3_w_n18666_0(.douta(w_n18666_0[0]),.doutb(w_n18666_0[1]),.doutc(w_n18666_0[2]),.din(n18666));
	jspl jspl_w_n18669_0(.douta(w_n18669_0[0]),.doutb(w_n18669_0[1]),.din(n18669));
	jspl jspl_w_n18670_0(.douta(w_n18670_0[0]),.doutb(w_n18670_0[1]),.din(n18670));
	jspl3 jspl3_w_n18671_0(.douta(w_n18671_0[0]),.doutb(w_n18671_0[1]),.doutc(w_n18671_0[2]),.din(n18671));
	jspl jspl_w_n18673_0(.douta(w_n18673_0[0]),.doutb(w_n18673_0[1]),.din(n18673));
	jspl jspl_w_n18677_0(.douta(w_n18677_0[0]),.doutb(w_n18677_0[1]),.din(n18677));
	jspl jspl_w_n18679_0(.douta(w_n18679_0[0]),.doutb(w_n18679_0[1]),.din(n18679));
	jspl jspl_w_n18680_0(.douta(w_n18680_0[0]),.doutb(w_n18680_0[1]),.din(n18680));
	jspl3 jspl3_w_n18681_0(.douta(w_n18681_0[0]),.doutb(w_n18681_0[1]),.doutc(w_n18681_0[2]),.din(n18681));
	jspl jspl_w_n18682_0(.douta(w_n18682_0[0]),.doutb(w_n18682_0[1]),.din(n18682));
	jspl jspl_w_n18685_0(.douta(w_n18685_0[0]),.doutb(w_n18685_0[1]),.din(n18685));
	jspl jspl_w_n18691_0(.douta(w_n18691_0[0]),.doutb(w_n18691_0[1]),.din(n18691));
	jspl jspl_w_n18692_0(.douta(w_n18692_0[0]),.doutb(w_n18692_0[1]),.din(n18692));
	jspl jspl_w_n18694_0(.douta(w_n18694_0[0]),.doutb(w_n18694_0[1]),.din(n18694));
	jspl jspl_w_n18696_0(.douta(w_n18696_0[0]),.doutb(w_n18696_0[1]),.din(n18696));
	jspl jspl_w_n18698_0(.douta(w_n18698_0[0]),.doutb(w_n18698_0[1]),.din(n18698));
	jspl jspl_w_n18704_0(.douta(w_n18704_0[0]),.doutb(w_n18704_0[1]),.din(n18704));
	jspl jspl_w_n18706_0(.douta(w_n18706_0[0]),.doutb(w_n18706_0[1]),.din(n18706));
	jspl3 jspl3_w_n18707_0(.douta(w_n18707_0[0]),.doutb(w_n18707_0[1]),.doutc(w_n18707_0[2]),.din(n18707));
	jspl jspl_w_n18710_0(.douta(w_n18710_0[0]),.doutb(w_n18710_0[1]),.din(n18710));
	jspl jspl_w_n18711_0(.douta(w_n18711_0[0]),.doutb(w_n18711_0[1]),.din(n18711));
	jspl3 jspl3_w_n18712_0(.douta(w_n18712_0[0]),.doutb(w_n18712_0[1]),.doutc(w_n18712_0[2]),.din(n18712));
	jspl jspl_w_n18714_0(.douta(w_n18714_0[0]),.doutb(w_n18714_0[1]),.din(n18714));
	jspl jspl_w_n18718_0(.douta(w_n18718_0[0]),.doutb(w_n18718_0[1]),.din(n18718));
	jspl jspl_w_n18720_0(.douta(w_n18720_0[0]),.doutb(w_n18720_0[1]),.din(n18720));
	jspl jspl_w_n18721_0(.douta(w_n18721_0[0]),.doutb(w_n18721_0[1]),.din(n18721));
	jspl3 jspl3_w_n18722_0(.douta(w_n18722_0[0]),.doutb(w_n18722_0[1]),.doutc(w_n18722_0[2]),.din(n18722));
	jspl jspl_w_n18723_0(.douta(w_n18723_0[0]),.doutb(w_n18723_0[1]),.din(n18723));
	jspl jspl_w_n18726_0(.douta(w_n18726_0[0]),.doutb(w_n18726_0[1]),.din(n18726));
	jspl jspl_w_n18732_0(.douta(w_n18732_0[0]),.doutb(w_n18732_0[1]),.din(n18732));
	jspl jspl_w_n18733_0(.douta(w_n18733_0[0]),.doutb(w_n18733_0[1]),.din(n18733));
	jspl jspl_w_n18735_0(.douta(w_n18735_0[0]),.doutb(w_n18735_0[1]),.din(n18735));
	jspl jspl_w_n18737_0(.douta(w_n18737_0[0]),.doutb(w_n18737_0[1]),.din(n18737));
	jspl jspl_w_n18739_0(.douta(w_n18739_0[0]),.doutb(w_n18739_0[1]),.din(n18739));
	jspl jspl_w_n18745_0(.douta(w_n18745_0[0]),.doutb(w_n18745_0[1]),.din(n18745));
	jspl jspl_w_n18747_0(.douta(w_n18747_0[0]),.doutb(w_n18747_0[1]),.din(n18747));
	jspl3 jspl3_w_n18748_0(.douta(w_n18748_0[0]),.doutb(w_n18748_0[1]),.doutc(w_n18748_0[2]),.din(n18748));
	jspl jspl_w_n18751_0(.douta(w_n18751_0[0]),.doutb(w_n18751_0[1]),.din(n18751));
	jspl jspl_w_n18752_0(.douta(w_n18752_0[0]),.doutb(w_n18752_0[1]),.din(n18752));
	jspl3 jspl3_w_n18753_0(.douta(w_n18753_0[0]),.doutb(w_n18753_0[1]),.doutc(w_n18753_0[2]),.din(n18753));
	jspl jspl_w_n18755_0(.douta(w_n18755_0[0]),.doutb(w_n18755_0[1]),.din(n18755));
	jspl jspl_w_n18759_0(.douta(w_n18759_0[0]),.doutb(w_n18759_0[1]),.din(n18759));
	jspl jspl_w_n18761_0(.douta(w_n18761_0[0]),.doutb(w_n18761_0[1]),.din(n18761));
	jspl jspl_w_n18762_0(.douta(w_n18762_0[0]),.doutb(w_n18762_0[1]),.din(n18762));
	jspl3 jspl3_w_n18763_0(.douta(w_n18763_0[0]),.doutb(w_n18763_0[1]),.doutc(w_n18763_0[2]),.din(n18763));
	jspl jspl_w_n18764_0(.douta(w_n18764_0[0]),.doutb(w_n18764_0[1]),.din(n18764));
	jspl jspl_w_n18767_0(.douta(w_n18767_0[0]),.doutb(w_n18767_0[1]),.din(n18767));
	jspl jspl_w_n18773_0(.douta(w_n18773_0[0]),.doutb(w_n18773_0[1]),.din(n18773));
	jspl jspl_w_n18774_0(.douta(w_n18774_0[0]),.doutb(w_n18774_0[1]),.din(n18774));
	jspl jspl_w_n18776_0(.douta(w_n18776_0[0]),.doutb(w_n18776_0[1]),.din(n18776));
	jspl jspl_w_n18778_0(.douta(w_n18778_0[0]),.doutb(w_n18778_0[1]),.din(n18778));
	jspl jspl_w_n18780_0(.douta(w_n18780_0[0]),.doutb(w_n18780_0[1]),.din(n18780));
	jspl jspl_w_n18786_0(.douta(w_n18786_0[0]),.doutb(w_n18786_0[1]),.din(n18786));
	jspl jspl_w_n18788_0(.douta(w_n18788_0[0]),.doutb(w_n18788_0[1]),.din(n18788));
	jspl3 jspl3_w_n18789_0(.douta(w_n18789_0[0]),.doutb(w_n18789_0[1]),.doutc(w_n18789_0[2]),.din(n18789));
	jspl jspl_w_n18792_0(.douta(w_n18792_0[0]),.doutb(w_n18792_0[1]),.din(n18792));
	jspl jspl_w_n18793_0(.douta(w_n18793_0[0]),.doutb(w_n18793_0[1]),.din(n18793));
	jspl3 jspl3_w_n18794_0(.douta(w_n18794_0[0]),.doutb(w_n18794_0[1]),.doutc(w_n18794_0[2]),.din(n18794));
	jspl jspl_w_n18796_0(.douta(w_n18796_0[0]),.doutb(w_n18796_0[1]),.din(n18796));
	jspl jspl_w_n18800_0(.douta(w_n18800_0[0]),.doutb(w_n18800_0[1]),.din(n18800));
	jspl jspl_w_n18802_0(.douta(w_n18802_0[0]),.doutb(w_n18802_0[1]),.din(n18802));
	jspl jspl_w_n18803_0(.douta(w_n18803_0[0]),.doutb(w_n18803_0[1]),.din(n18803));
	jspl3 jspl3_w_n18804_0(.douta(w_n18804_0[0]),.doutb(w_n18804_0[1]),.doutc(w_n18804_0[2]),.din(n18804));
	jspl jspl_w_n18805_0(.douta(w_n18805_0[0]),.doutb(w_n18805_0[1]),.din(n18805));
	jspl jspl_w_n18808_0(.douta(w_n18808_0[0]),.doutb(w_n18808_0[1]),.din(n18808));
	jspl jspl_w_n18814_0(.douta(w_n18814_0[0]),.doutb(w_n18814_0[1]),.din(n18814));
	jspl jspl_w_n18815_0(.douta(w_n18815_0[0]),.doutb(w_n18815_0[1]),.din(n18815));
	jspl jspl_w_n18817_0(.douta(w_n18817_0[0]),.doutb(w_n18817_0[1]),.din(n18817));
	jspl jspl_w_n18819_0(.douta(w_n18819_0[0]),.doutb(w_n18819_0[1]),.din(n18819));
	jspl jspl_w_n18821_0(.douta(w_n18821_0[0]),.doutb(w_n18821_0[1]),.din(n18821));
	jspl jspl_w_n18827_0(.douta(w_n18827_0[0]),.doutb(w_n18827_0[1]),.din(n18827));
	jspl jspl_w_n18829_0(.douta(w_n18829_0[0]),.doutb(w_n18829_0[1]),.din(n18829));
	jspl3 jspl3_w_n18830_0(.douta(w_n18830_0[0]),.doutb(w_n18830_0[1]),.doutc(w_n18830_0[2]),.din(n18830));
	jspl jspl_w_n18833_0(.douta(w_n18833_0[0]),.doutb(w_n18833_0[1]),.din(n18833));
	jspl jspl_w_n18834_0(.douta(w_n18834_0[0]),.doutb(w_n18834_0[1]),.din(n18834));
	jspl3 jspl3_w_n18835_0(.douta(w_n18835_0[0]),.doutb(w_n18835_0[1]),.doutc(w_n18835_0[2]),.din(n18835));
	jspl jspl_w_n18837_0(.douta(w_n18837_0[0]),.doutb(w_n18837_0[1]),.din(n18837));
	jspl jspl_w_n18841_0(.douta(w_n18841_0[0]),.doutb(w_n18841_0[1]),.din(n18841));
	jspl jspl_w_n18843_0(.douta(w_n18843_0[0]),.doutb(w_n18843_0[1]),.din(n18843));
	jspl jspl_w_n18844_0(.douta(w_n18844_0[0]),.doutb(w_n18844_0[1]),.din(n18844));
	jspl3 jspl3_w_n18845_0(.douta(w_n18845_0[0]),.doutb(w_n18845_0[1]),.doutc(w_n18845_0[2]),.din(n18845));
	jspl jspl_w_n18846_0(.douta(w_n18846_0[0]),.doutb(w_n18846_0[1]),.din(n18846));
	jspl jspl_w_n18849_0(.douta(w_n18849_0[0]),.doutb(w_n18849_0[1]),.din(n18849));
	jspl jspl_w_n18855_0(.douta(w_n18855_0[0]),.doutb(w_n18855_0[1]),.din(n18855));
	jspl jspl_w_n18856_0(.douta(w_n18856_0[0]),.doutb(w_n18856_0[1]),.din(n18856));
	jspl jspl_w_n18858_0(.douta(w_n18858_0[0]),.doutb(w_n18858_0[1]),.din(n18858));
	jspl jspl_w_n18860_0(.douta(w_n18860_0[0]),.doutb(w_n18860_0[1]),.din(n18860));
	jspl jspl_w_n18862_0(.douta(w_n18862_0[0]),.doutb(w_n18862_0[1]),.din(n18862));
	jspl jspl_w_n18868_0(.douta(w_n18868_0[0]),.doutb(w_n18868_0[1]),.din(n18868));
	jspl jspl_w_n18870_0(.douta(w_n18870_0[0]),.doutb(w_n18870_0[1]),.din(n18870));
	jspl3 jspl3_w_n18871_0(.douta(w_n18871_0[0]),.doutb(w_n18871_0[1]),.doutc(w_n18871_0[2]),.din(n18871));
	jspl jspl_w_n18874_0(.douta(w_n18874_0[0]),.doutb(w_n18874_0[1]),.din(n18874));
	jspl jspl_w_n18875_0(.douta(w_n18875_0[0]),.doutb(w_n18875_0[1]),.din(n18875));
	jspl3 jspl3_w_n18876_0(.douta(w_n18876_0[0]),.doutb(w_n18876_0[1]),.doutc(w_n18876_0[2]),.din(n18876));
	jspl jspl_w_n18878_0(.douta(w_n18878_0[0]),.doutb(w_n18878_0[1]),.din(n18878));
	jspl jspl_w_n18880_0(.douta(w_n18880_0[0]),.doutb(w_n18880_0[1]),.din(n18880));
	jspl jspl_w_n18882_0(.douta(w_n18882_0[0]),.doutb(w_n18882_0[1]),.din(n18882));
	jspl jspl_w_n18888_0(.douta(w_n18888_0[0]),.doutb(w_n18888_0[1]),.din(n18888));
	jspl3 jspl3_w_n18890_0(.douta(w_n18890_0[0]),.doutb(w_n18890_0[1]),.doutc(w_n18890_0[2]),.din(n18890));
	jspl jspl_w_n18891_0(.douta(w_n18891_0[0]),.doutb(w_n18891_0[1]),.din(n18891));
	jspl jspl_w_n18894_0(.douta(w_n18894_0[0]),.doutb(w_n18894_0[1]),.din(n18894));
	jspl jspl_w_n18896_0(.douta(w_n18896_0[0]),.doutb(w_n18896_0[1]),.din(n18896));
	jspl jspl_w_n18900_0(.douta(w_n18900_0[0]),.doutb(w_n18900_0[1]),.din(n18900));
	jspl jspl_w_n18902_0(.douta(w_n18902_0[0]),.doutb(w_n18902_0[1]),.din(n18902));
	jspl jspl_w_n18903_0(.douta(w_n18903_0[0]),.doutb(w_n18903_0[1]),.din(n18903));
	jspl jspl_w_n18904_0(.douta(w_n18904_0[0]),.doutb(w_n18904_0[1]),.din(n18904));
	jspl3 jspl3_w_n18905_0(.douta(w_n18905_0[0]),.doutb(w_n18905_0[1]),.doutc(w_n18905_0[2]),.din(n18905));
	jspl jspl_w_n18908_0(.douta(w_n18908_0[0]),.doutb(w_n18908_0[1]),.din(n18908));
	jspl jspl_w_n18909_0(.douta(w_n18909_0[0]),.doutb(w_n18909_0[1]),.din(n18909));
	jspl3 jspl3_w_n18910_0(.douta(w_n18910_0[0]),.doutb(w_n18910_0[1]),.doutc(w_n18910_0[2]),.din(n18910));
	jspl jspl_w_n18912_0(.douta(w_n18912_0[0]),.doutb(w_n18912_0[1]),.din(n18912));
	jspl jspl_w_n18916_0(.douta(w_n18916_0[0]),.doutb(w_n18916_0[1]),.din(n18916));
	jspl jspl_w_n18918_0(.douta(w_n18918_0[0]),.doutb(w_n18918_0[1]),.din(n18918));
	jspl jspl_w_n18919_0(.douta(w_n18919_0[0]),.doutb(w_n18919_0[1]),.din(n18919));
	jspl3 jspl3_w_n18920_0(.douta(w_n18920_0[0]),.doutb(w_n18920_0[1]),.doutc(w_n18920_0[2]),.din(n18920));
	jspl jspl_w_n18924_0(.douta(w_n18924_0[0]),.doutb(w_n18924_0[1]),.din(n18924));
	jspl jspl_w_n18930_0(.douta(w_n18930_0[0]),.doutb(w_n18930_0[1]),.din(n18930));
	jspl3 jspl3_w_n18932_0(.douta(w_n18932_0[0]),.doutb(w_n18932_0[1]),.doutc(w_n18932_0[2]),.din(n18932));
	jspl jspl_w_n18934_0(.douta(w_n18934_0[0]),.doutb(w_n18934_0[1]),.din(n18934));
	jspl3 jspl3_w_n18939_0(.douta(w_n18939_0[0]),.doutb(w_n18939_0[1]),.doutc(w_n18939_0[2]),.din(n18939));
	jspl jspl_w_n18940_0(.douta(w_n18940_0[0]),.doutb(w_n18940_0[1]),.din(n18940));
	jspl jspl_w_n18942_0(.douta(w_n18942_0[0]),.doutb(w_n18942_0[1]),.din(n18942));
	jspl jspl_w_n18948_0(.douta(w_n18948_0[0]),.doutb(w_n18948_0[1]),.din(n18948));
	jspl jspl_w_n18958_0(.douta(w_n18958_0[0]),.doutb(w_n18958_0[1]),.din(n18958));
	jspl3 jspl3_w_n18961_0(.douta(w_n18961_0[0]),.doutb(w_n18961_0[1]),.doutc(w_n18961_0[2]),.din(n18961));
	jspl jspl_w_n18961_1(.douta(w_n18961_1[0]),.doutb(w_n18961_1[1]),.din(w_n18961_0[0]));
	jspl jspl_w_n18962_0(.douta(w_n18962_0[0]),.doutb(w_n18962_0[1]),.din(n18962));
	jspl3 jspl3_w_n18965_0(.douta(w_n18965_0[0]),.doutb(w_n18965_0[1]),.doutc(w_n18965_0[2]),.din(n18965));
	jspl jspl_w_n18966_0(.douta(w_n18966_0[0]),.doutb(w_n18966_0[1]),.din(n18966));
	jspl jspl_w_n18967_0(.douta(w_n18967_0[0]),.doutb(w_n18967_0[1]),.din(n18967));
	jspl jspl_w_n18968_0(.douta(w_n18968_0[0]),.doutb(w_n18968_0[1]),.din(n18968));
	jspl jspl_w_n18970_0(.douta(w_n18970_0[0]),.doutb(w_n18970_0[1]),.din(n18970));
	jspl jspl_w_n18972_0(.douta(w_n18972_0[0]),.doutb(w_n18972_0[1]),.din(n18972));
	jspl jspl_w_n18974_0(.douta(w_n18974_0[0]),.doutb(w_n18974_0[1]),.din(n18974));
	jspl3 jspl3_w_n18976_0(.douta(w_n18976_0[0]),.doutb(w_n18976_0[1]),.doutc(w_n18976_0[2]),.din(n18976));
	jspl3 jspl3_w_n18976_1(.douta(w_n18976_1[0]),.doutb(w_n18976_1[1]),.doutc(w_n18976_1[2]),.din(w_n18976_0[0]));
	jspl3 jspl3_w_n18976_2(.douta(w_n18976_2[0]),.doutb(w_n18976_2[1]),.doutc(w_n18976_2[2]),.din(w_n18976_0[1]));
	jspl jspl_w_n18979_0(.douta(w_n18979_0[0]),.doutb(w_n18979_0[1]),.din(n18979));
	jspl3 jspl3_w_n18981_0(.douta(w_n18981_0[0]),.doutb(w_n18981_0[1]),.doutc(w_n18981_0[2]),.din(n18981));
	jspl jspl_w_n18982_0(.douta(w_n18982_0[0]),.doutb(w_n18982_0[1]),.din(n18982));
	jspl jspl_w_n18986_0(.douta(w_n18986_0[0]),.doutb(w_n18986_0[1]),.din(n18986));
	jspl jspl_w_n18988_0(.douta(w_n18988_0[0]),.doutb(w_n18988_0[1]),.din(n18988));
	jspl jspl_w_n18990_0(.douta(w_n18990_0[0]),.doutb(w_n18990_0[1]),.din(n18990));
	jspl jspl_w_n18995_0(.douta(w_n18995_0[0]),.doutb(w_n18995_0[1]),.din(n18995));
	jspl jspl_w_n18997_0(.douta(w_n18997_0[0]),.doutb(w_n18997_0[1]),.din(n18997));
	jspl jspl_w_n18998_0(.douta(w_n18998_0[0]),.doutb(w_n18998_0[1]),.din(n18998));
	jspl3 jspl3_w_n18999_0(.douta(w_n18999_0[0]),.doutb(w_n18999_0[1]),.doutc(w_n18999_0[2]),.din(n18999));
	jspl jspl_w_n19000_0(.douta(w_n19000_0[0]),.doutb(w_n19000_0[1]),.din(n19000));
	jspl jspl_w_n19005_0(.douta(w_n19005_0[0]),.doutb(w_n19005_0[1]),.din(n19005));
	jspl jspl_w_n19006_0(.douta(w_n19006_0[0]),.doutb(w_n19006_0[1]),.din(n19006));
	jspl jspl_w_n19008_0(.douta(w_n19008_0[0]),.doutb(w_n19008_0[1]),.din(n19008));
	jspl jspl_w_n19010_0(.douta(w_n19010_0[0]),.doutb(w_n19010_0[1]),.din(n19010));
	jspl jspl_w_n19013_0(.douta(w_n19013_0[0]),.doutb(w_n19013_0[1]),.din(n19013));
	jspl jspl_w_n19019_0(.douta(w_n19019_0[0]),.doutb(w_n19019_0[1]),.din(n19019));
	jspl3 jspl3_w_n19021_0(.douta(w_n19021_0[0]),.doutb(w_n19021_0[1]),.doutc(w_n19021_0[2]),.din(n19021));
	jspl jspl_w_n19022_0(.douta(w_n19022_0[0]),.doutb(w_n19022_0[1]),.din(n19022));
	jspl jspl_w_n19026_0(.douta(w_n19026_0[0]),.doutb(w_n19026_0[1]),.din(n19026));
	jspl jspl_w_n19027_0(.douta(w_n19027_0[0]),.doutb(w_n19027_0[1]),.din(n19027));
	jspl jspl_w_n19029_0(.douta(w_n19029_0[0]),.doutb(w_n19029_0[1]),.din(n19029));
	jspl jspl_w_n19034_0(.douta(w_n19034_0[0]),.doutb(w_n19034_0[1]),.din(n19034));
	jspl jspl_w_n19036_0(.douta(w_n19036_0[0]),.doutb(w_n19036_0[1]),.din(n19036));
	jspl jspl_w_n19037_0(.douta(w_n19037_0[0]),.doutb(w_n19037_0[1]),.din(n19037));
	jspl3 jspl3_w_n19038_0(.douta(w_n19038_0[0]),.doutb(w_n19038_0[1]),.doutc(w_n19038_0[2]),.din(n19038));
	jspl jspl_w_n19039_0(.douta(w_n19039_0[0]),.doutb(w_n19039_0[1]),.din(n19039));
	jspl jspl_w_n19043_0(.douta(w_n19043_0[0]),.doutb(w_n19043_0[1]),.din(n19043));
	jspl jspl_w_n19044_0(.douta(w_n19044_0[0]),.doutb(w_n19044_0[1]),.din(n19044));
	jspl jspl_w_n19046_0(.douta(w_n19046_0[0]),.doutb(w_n19046_0[1]),.din(n19046));
	jspl jspl_w_n19048_0(.douta(w_n19048_0[0]),.doutb(w_n19048_0[1]),.din(n19048));
	jspl jspl_w_n19051_0(.douta(w_n19051_0[0]),.doutb(w_n19051_0[1]),.din(n19051));
	jspl jspl_w_n19057_0(.douta(w_n19057_0[0]),.doutb(w_n19057_0[1]),.din(n19057));
	jspl jspl_w_n19059_0(.douta(w_n19059_0[0]),.doutb(w_n19059_0[1]),.din(n19059));
	jspl3 jspl3_w_n19060_0(.douta(w_n19060_0[0]),.doutb(w_n19060_0[1]),.doutc(w_n19060_0[2]),.din(n19060));
	jspl jspl_w_n19064_0(.douta(w_n19064_0[0]),.doutb(w_n19064_0[1]),.din(n19064));
	jspl jspl_w_n19065_0(.douta(w_n19065_0[0]),.doutb(w_n19065_0[1]),.din(n19065));
	jspl3 jspl3_w_n19066_0(.douta(w_n19066_0[0]),.doutb(w_n19066_0[1]),.doutc(w_n19066_0[2]),.din(n19066));
	jspl jspl_w_n19068_0(.douta(w_n19068_0[0]),.doutb(w_n19068_0[1]),.din(n19068));
	jspl jspl_w_n19073_0(.douta(w_n19073_0[0]),.doutb(w_n19073_0[1]),.din(n19073));
	jspl jspl_w_n19075_0(.douta(w_n19075_0[0]),.doutb(w_n19075_0[1]),.din(n19075));
	jspl jspl_w_n19076_0(.douta(w_n19076_0[0]),.doutb(w_n19076_0[1]),.din(n19076));
	jspl3 jspl3_w_n19077_0(.douta(w_n19077_0[0]),.doutb(w_n19077_0[1]),.doutc(w_n19077_0[2]),.din(n19077));
	jspl jspl_w_n19078_0(.douta(w_n19078_0[0]),.doutb(w_n19078_0[1]),.din(n19078));
	jspl jspl_w_n19082_0(.douta(w_n19082_0[0]),.doutb(w_n19082_0[1]),.din(n19082));
	jspl jspl_w_n19088_0(.douta(w_n19088_0[0]),.doutb(w_n19088_0[1]),.din(n19088));
	jspl jspl_w_n19089_0(.douta(w_n19089_0[0]),.doutb(w_n19089_0[1]),.din(n19089));
	jspl jspl_w_n19091_0(.douta(w_n19091_0[0]),.doutb(w_n19091_0[1]),.din(n19091));
	jspl jspl_w_n19093_0(.douta(w_n19093_0[0]),.doutb(w_n19093_0[1]),.din(n19093));
	jspl jspl_w_n19096_0(.douta(w_n19096_0[0]),.doutb(w_n19096_0[1]),.din(n19096));
	jspl jspl_w_n19102_0(.douta(w_n19102_0[0]),.doutb(w_n19102_0[1]),.din(n19102));
	jspl jspl_w_n19104_0(.douta(w_n19104_0[0]),.doutb(w_n19104_0[1]),.din(n19104));
	jspl3 jspl3_w_n19105_0(.douta(w_n19105_0[0]),.doutb(w_n19105_0[1]),.doutc(w_n19105_0[2]),.din(n19105));
	jspl jspl_w_n19109_0(.douta(w_n19109_0[0]),.doutb(w_n19109_0[1]),.din(n19109));
	jspl jspl_w_n19110_0(.douta(w_n19110_0[0]),.doutb(w_n19110_0[1]),.din(n19110));
	jspl3 jspl3_w_n19111_0(.douta(w_n19111_0[0]),.doutb(w_n19111_0[1]),.doutc(w_n19111_0[2]),.din(n19111));
	jspl jspl_w_n19113_0(.douta(w_n19113_0[0]),.doutb(w_n19113_0[1]),.din(n19113));
	jspl jspl_w_n19118_0(.douta(w_n19118_0[0]),.doutb(w_n19118_0[1]),.din(n19118));
	jspl jspl_w_n19120_0(.douta(w_n19120_0[0]),.doutb(w_n19120_0[1]),.din(n19120));
	jspl jspl_w_n19121_0(.douta(w_n19121_0[0]),.doutb(w_n19121_0[1]),.din(n19121));
	jspl3 jspl3_w_n19122_0(.douta(w_n19122_0[0]),.doutb(w_n19122_0[1]),.doutc(w_n19122_0[2]),.din(n19122));
	jspl jspl_w_n19123_0(.douta(w_n19123_0[0]),.doutb(w_n19123_0[1]),.din(n19123));
	jspl jspl_w_n19127_0(.douta(w_n19127_0[0]),.doutb(w_n19127_0[1]),.din(n19127));
	jspl jspl_w_n19133_0(.douta(w_n19133_0[0]),.doutb(w_n19133_0[1]),.din(n19133));
	jspl jspl_w_n19134_0(.douta(w_n19134_0[0]),.doutb(w_n19134_0[1]),.din(n19134));
	jspl jspl_w_n19136_0(.douta(w_n19136_0[0]),.doutb(w_n19136_0[1]),.din(n19136));
	jspl jspl_w_n19138_0(.douta(w_n19138_0[0]),.doutb(w_n19138_0[1]),.din(n19138));
	jspl jspl_w_n19141_0(.douta(w_n19141_0[0]),.doutb(w_n19141_0[1]),.din(n19141));
	jspl jspl_w_n19147_0(.douta(w_n19147_0[0]),.doutb(w_n19147_0[1]),.din(n19147));
	jspl jspl_w_n19149_0(.douta(w_n19149_0[0]),.doutb(w_n19149_0[1]),.din(n19149));
	jspl3 jspl3_w_n19150_0(.douta(w_n19150_0[0]),.doutb(w_n19150_0[1]),.doutc(w_n19150_0[2]),.din(n19150));
	jspl jspl_w_n19154_0(.douta(w_n19154_0[0]),.doutb(w_n19154_0[1]),.din(n19154));
	jspl jspl_w_n19155_0(.douta(w_n19155_0[0]),.doutb(w_n19155_0[1]),.din(n19155));
	jspl3 jspl3_w_n19156_0(.douta(w_n19156_0[0]),.doutb(w_n19156_0[1]),.doutc(w_n19156_0[2]),.din(n19156));
	jspl jspl_w_n19158_0(.douta(w_n19158_0[0]),.doutb(w_n19158_0[1]),.din(n19158));
	jspl jspl_w_n19163_0(.douta(w_n19163_0[0]),.doutb(w_n19163_0[1]),.din(n19163));
	jspl jspl_w_n19165_0(.douta(w_n19165_0[0]),.doutb(w_n19165_0[1]),.din(n19165));
	jspl jspl_w_n19166_0(.douta(w_n19166_0[0]),.doutb(w_n19166_0[1]),.din(n19166));
	jspl3 jspl3_w_n19167_0(.douta(w_n19167_0[0]),.doutb(w_n19167_0[1]),.doutc(w_n19167_0[2]),.din(n19167));
	jspl jspl_w_n19168_0(.douta(w_n19168_0[0]),.doutb(w_n19168_0[1]),.din(n19168));
	jspl jspl_w_n19172_0(.douta(w_n19172_0[0]),.doutb(w_n19172_0[1]),.din(n19172));
	jspl jspl_w_n19178_0(.douta(w_n19178_0[0]),.doutb(w_n19178_0[1]),.din(n19178));
	jspl jspl_w_n19179_0(.douta(w_n19179_0[0]),.doutb(w_n19179_0[1]),.din(n19179));
	jspl jspl_w_n19181_0(.douta(w_n19181_0[0]),.doutb(w_n19181_0[1]),.din(n19181));
	jspl jspl_w_n19183_0(.douta(w_n19183_0[0]),.doutb(w_n19183_0[1]),.din(n19183));
	jspl jspl_w_n19186_0(.douta(w_n19186_0[0]),.doutb(w_n19186_0[1]),.din(n19186));
	jspl jspl_w_n19192_0(.douta(w_n19192_0[0]),.doutb(w_n19192_0[1]),.din(n19192));
	jspl jspl_w_n19194_0(.douta(w_n19194_0[0]),.doutb(w_n19194_0[1]),.din(n19194));
	jspl3 jspl3_w_n19195_0(.douta(w_n19195_0[0]),.doutb(w_n19195_0[1]),.doutc(w_n19195_0[2]),.din(n19195));
	jspl jspl_w_n19199_0(.douta(w_n19199_0[0]),.doutb(w_n19199_0[1]),.din(n19199));
	jspl jspl_w_n19200_0(.douta(w_n19200_0[0]),.doutb(w_n19200_0[1]),.din(n19200));
	jspl3 jspl3_w_n19201_0(.douta(w_n19201_0[0]),.doutb(w_n19201_0[1]),.doutc(w_n19201_0[2]),.din(n19201));
	jspl jspl_w_n19203_0(.douta(w_n19203_0[0]),.doutb(w_n19203_0[1]),.din(n19203));
	jspl jspl_w_n19208_0(.douta(w_n19208_0[0]),.doutb(w_n19208_0[1]),.din(n19208));
	jspl jspl_w_n19210_0(.douta(w_n19210_0[0]),.doutb(w_n19210_0[1]),.din(n19210));
	jspl jspl_w_n19211_0(.douta(w_n19211_0[0]),.doutb(w_n19211_0[1]),.din(n19211));
	jspl3 jspl3_w_n19212_0(.douta(w_n19212_0[0]),.doutb(w_n19212_0[1]),.doutc(w_n19212_0[2]),.din(n19212));
	jspl jspl_w_n19213_0(.douta(w_n19213_0[0]),.doutb(w_n19213_0[1]),.din(n19213));
	jspl jspl_w_n19217_0(.douta(w_n19217_0[0]),.doutb(w_n19217_0[1]),.din(n19217));
	jspl jspl_w_n19223_0(.douta(w_n19223_0[0]),.doutb(w_n19223_0[1]),.din(n19223));
	jspl jspl_w_n19224_0(.douta(w_n19224_0[0]),.doutb(w_n19224_0[1]),.din(n19224));
	jspl jspl_w_n19226_0(.douta(w_n19226_0[0]),.doutb(w_n19226_0[1]),.din(n19226));
	jspl jspl_w_n19228_0(.douta(w_n19228_0[0]),.doutb(w_n19228_0[1]),.din(n19228));
	jspl jspl_w_n19231_0(.douta(w_n19231_0[0]),.doutb(w_n19231_0[1]),.din(n19231));
	jspl jspl_w_n19237_0(.douta(w_n19237_0[0]),.doutb(w_n19237_0[1]),.din(n19237));
	jspl jspl_w_n19239_0(.douta(w_n19239_0[0]),.doutb(w_n19239_0[1]),.din(n19239));
	jspl3 jspl3_w_n19240_0(.douta(w_n19240_0[0]),.doutb(w_n19240_0[1]),.doutc(w_n19240_0[2]),.din(n19240));
	jspl jspl_w_n19244_0(.douta(w_n19244_0[0]),.doutb(w_n19244_0[1]),.din(n19244));
	jspl jspl_w_n19245_0(.douta(w_n19245_0[0]),.doutb(w_n19245_0[1]),.din(n19245));
	jspl3 jspl3_w_n19246_0(.douta(w_n19246_0[0]),.doutb(w_n19246_0[1]),.doutc(w_n19246_0[2]),.din(n19246));
	jspl jspl_w_n19248_0(.douta(w_n19248_0[0]),.doutb(w_n19248_0[1]),.din(n19248));
	jspl jspl_w_n19253_0(.douta(w_n19253_0[0]),.doutb(w_n19253_0[1]),.din(n19253));
	jspl jspl_w_n19255_0(.douta(w_n19255_0[0]),.doutb(w_n19255_0[1]),.din(n19255));
	jspl jspl_w_n19256_0(.douta(w_n19256_0[0]),.doutb(w_n19256_0[1]),.din(n19256));
	jspl3 jspl3_w_n19257_0(.douta(w_n19257_0[0]),.doutb(w_n19257_0[1]),.doutc(w_n19257_0[2]),.din(n19257));
	jspl jspl_w_n19258_0(.douta(w_n19258_0[0]),.doutb(w_n19258_0[1]),.din(n19258));
	jspl jspl_w_n19262_0(.douta(w_n19262_0[0]),.doutb(w_n19262_0[1]),.din(n19262));
	jspl jspl_w_n19268_0(.douta(w_n19268_0[0]),.doutb(w_n19268_0[1]),.din(n19268));
	jspl jspl_w_n19269_0(.douta(w_n19269_0[0]),.doutb(w_n19269_0[1]),.din(n19269));
	jspl jspl_w_n19271_0(.douta(w_n19271_0[0]),.doutb(w_n19271_0[1]),.din(n19271));
	jspl jspl_w_n19273_0(.douta(w_n19273_0[0]),.doutb(w_n19273_0[1]),.din(n19273));
	jspl jspl_w_n19276_0(.douta(w_n19276_0[0]),.doutb(w_n19276_0[1]),.din(n19276));
	jspl jspl_w_n19282_0(.douta(w_n19282_0[0]),.doutb(w_n19282_0[1]),.din(n19282));
	jspl jspl_w_n19284_0(.douta(w_n19284_0[0]),.doutb(w_n19284_0[1]),.din(n19284));
	jspl3 jspl3_w_n19285_0(.douta(w_n19285_0[0]),.doutb(w_n19285_0[1]),.doutc(w_n19285_0[2]),.din(n19285));
	jspl jspl_w_n19289_0(.douta(w_n19289_0[0]),.doutb(w_n19289_0[1]),.din(n19289));
	jspl jspl_w_n19290_0(.douta(w_n19290_0[0]),.doutb(w_n19290_0[1]),.din(n19290));
	jspl3 jspl3_w_n19291_0(.douta(w_n19291_0[0]),.doutb(w_n19291_0[1]),.doutc(w_n19291_0[2]),.din(n19291));
	jspl jspl_w_n19293_0(.douta(w_n19293_0[0]),.doutb(w_n19293_0[1]),.din(n19293));
	jspl jspl_w_n19298_0(.douta(w_n19298_0[0]),.doutb(w_n19298_0[1]),.din(n19298));
	jspl jspl_w_n19300_0(.douta(w_n19300_0[0]),.doutb(w_n19300_0[1]),.din(n19300));
	jspl jspl_w_n19301_0(.douta(w_n19301_0[0]),.doutb(w_n19301_0[1]),.din(n19301));
	jspl3 jspl3_w_n19302_0(.douta(w_n19302_0[0]),.doutb(w_n19302_0[1]),.doutc(w_n19302_0[2]),.din(n19302));
	jspl jspl_w_n19303_0(.douta(w_n19303_0[0]),.doutb(w_n19303_0[1]),.din(n19303));
	jspl jspl_w_n19307_0(.douta(w_n19307_0[0]),.doutb(w_n19307_0[1]),.din(n19307));
	jspl jspl_w_n19313_0(.douta(w_n19313_0[0]),.doutb(w_n19313_0[1]),.din(n19313));
	jspl jspl_w_n19314_0(.douta(w_n19314_0[0]),.doutb(w_n19314_0[1]),.din(n19314));
	jspl jspl_w_n19316_0(.douta(w_n19316_0[0]),.doutb(w_n19316_0[1]),.din(n19316));
	jspl jspl_w_n19318_0(.douta(w_n19318_0[0]),.doutb(w_n19318_0[1]),.din(n19318));
	jspl jspl_w_n19321_0(.douta(w_n19321_0[0]),.doutb(w_n19321_0[1]),.din(n19321));
	jspl jspl_w_n19327_0(.douta(w_n19327_0[0]),.doutb(w_n19327_0[1]),.din(n19327));
	jspl jspl_w_n19329_0(.douta(w_n19329_0[0]),.doutb(w_n19329_0[1]),.din(n19329));
	jspl3 jspl3_w_n19330_0(.douta(w_n19330_0[0]),.doutb(w_n19330_0[1]),.doutc(w_n19330_0[2]),.din(n19330));
	jspl jspl_w_n19334_0(.douta(w_n19334_0[0]),.doutb(w_n19334_0[1]),.din(n19334));
	jspl jspl_w_n19335_0(.douta(w_n19335_0[0]),.doutb(w_n19335_0[1]),.din(n19335));
	jspl3 jspl3_w_n19336_0(.douta(w_n19336_0[0]),.doutb(w_n19336_0[1]),.doutc(w_n19336_0[2]),.din(n19336));
	jspl jspl_w_n19338_0(.douta(w_n19338_0[0]),.doutb(w_n19338_0[1]),.din(n19338));
	jspl jspl_w_n19343_0(.douta(w_n19343_0[0]),.doutb(w_n19343_0[1]),.din(n19343));
	jspl jspl_w_n19345_0(.douta(w_n19345_0[0]),.doutb(w_n19345_0[1]),.din(n19345));
	jspl jspl_w_n19346_0(.douta(w_n19346_0[0]),.doutb(w_n19346_0[1]),.din(n19346));
	jspl3 jspl3_w_n19347_0(.douta(w_n19347_0[0]),.doutb(w_n19347_0[1]),.doutc(w_n19347_0[2]),.din(n19347));
	jspl jspl_w_n19348_0(.douta(w_n19348_0[0]),.doutb(w_n19348_0[1]),.din(n19348));
	jspl jspl_w_n19352_0(.douta(w_n19352_0[0]),.doutb(w_n19352_0[1]),.din(n19352));
	jspl jspl_w_n19358_0(.douta(w_n19358_0[0]),.doutb(w_n19358_0[1]),.din(n19358));
	jspl jspl_w_n19359_0(.douta(w_n19359_0[0]),.doutb(w_n19359_0[1]),.din(n19359));
	jspl jspl_w_n19361_0(.douta(w_n19361_0[0]),.doutb(w_n19361_0[1]),.din(n19361));
	jspl jspl_w_n19363_0(.douta(w_n19363_0[0]),.doutb(w_n19363_0[1]),.din(n19363));
	jspl jspl_w_n19366_0(.douta(w_n19366_0[0]),.doutb(w_n19366_0[1]),.din(n19366));
	jspl jspl_w_n19372_0(.douta(w_n19372_0[0]),.doutb(w_n19372_0[1]),.din(n19372));
	jspl jspl_w_n19374_0(.douta(w_n19374_0[0]),.doutb(w_n19374_0[1]),.din(n19374));
	jspl3 jspl3_w_n19375_0(.douta(w_n19375_0[0]),.doutb(w_n19375_0[1]),.doutc(w_n19375_0[2]),.din(n19375));
	jspl jspl_w_n19379_0(.douta(w_n19379_0[0]),.doutb(w_n19379_0[1]),.din(n19379));
	jspl jspl_w_n19380_0(.douta(w_n19380_0[0]),.doutb(w_n19380_0[1]),.din(n19380));
	jspl3 jspl3_w_n19381_0(.douta(w_n19381_0[0]),.doutb(w_n19381_0[1]),.doutc(w_n19381_0[2]),.din(n19381));
	jspl jspl_w_n19383_0(.douta(w_n19383_0[0]),.doutb(w_n19383_0[1]),.din(n19383));
	jspl jspl_w_n19388_0(.douta(w_n19388_0[0]),.doutb(w_n19388_0[1]),.din(n19388));
	jspl jspl_w_n19390_0(.douta(w_n19390_0[0]),.doutb(w_n19390_0[1]),.din(n19390));
	jspl jspl_w_n19391_0(.douta(w_n19391_0[0]),.doutb(w_n19391_0[1]),.din(n19391));
	jspl3 jspl3_w_n19392_0(.douta(w_n19392_0[0]),.doutb(w_n19392_0[1]),.doutc(w_n19392_0[2]),.din(n19392));
	jspl jspl_w_n19393_0(.douta(w_n19393_0[0]),.doutb(w_n19393_0[1]),.din(n19393));
	jspl jspl_w_n19397_0(.douta(w_n19397_0[0]),.doutb(w_n19397_0[1]),.din(n19397));
	jspl jspl_w_n19403_0(.douta(w_n19403_0[0]),.doutb(w_n19403_0[1]),.din(n19403));
	jspl jspl_w_n19404_0(.douta(w_n19404_0[0]),.doutb(w_n19404_0[1]),.din(n19404));
	jspl jspl_w_n19406_0(.douta(w_n19406_0[0]),.doutb(w_n19406_0[1]),.din(n19406));
	jspl jspl_w_n19408_0(.douta(w_n19408_0[0]),.doutb(w_n19408_0[1]),.din(n19408));
	jspl jspl_w_n19411_0(.douta(w_n19411_0[0]),.doutb(w_n19411_0[1]),.din(n19411));
	jspl jspl_w_n19417_0(.douta(w_n19417_0[0]),.doutb(w_n19417_0[1]),.din(n19417));
	jspl jspl_w_n19419_0(.douta(w_n19419_0[0]),.doutb(w_n19419_0[1]),.din(n19419));
	jspl3 jspl3_w_n19420_0(.douta(w_n19420_0[0]),.doutb(w_n19420_0[1]),.doutc(w_n19420_0[2]),.din(n19420));
	jspl jspl_w_n19424_0(.douta(w_n19424_0[0]),.doutb(w_n19424_0[1]),.din(n19424));
	jspl jspl_w_n19425_0(.douta(w_n19425_0[0]),.doutb(w_n19425_0[1]),.din(n19425));
	jspl3 jspl3_w_n19426_0(.douta(w_n19426_0[0]),.doutb(w_n19426_0[1]),.doutc(w_n19426_0[2]),.din(n19426));
	jspl jspl_w_n19428_0(.douta(w_n19428_0[0]),.doutb(w_n19428_0[1]),.din(n19428));
	jspl jspl_w_n19433_0(.douta(w_n19433_0[0]),.doutb(w_n19433_0[1]),.din(n19433));
	jspl jspl_w_n19435_0(.douta(w_n19435_0[0]),.doutb(w_n19435_0[1]),.din(n19435));
	jspl jspl_w_n19436_0(.douta(w_n19436_0[0]),.doutb(w_n19436_0[1]),.din(n19436));
	jspl3 jspl3_w_n19437_0(.douta(w_n19437_0[0]),.doutb(w_n19437_0[1]),.doutc(w_n19437_0[2]),.din(n19437));
	jspl jspl_w_n19438_0(.douta(w_n19438_0[0]),.doutb(w_n19438_0[1]),.din(n19438));
	jspl jspl_w_n19442_0(.douta(w_n19442_0[0]),.doutb(w_n19442_0[1]),.din(n19442));
	jspl jspl_w_n19448_0(.douta(w_n19448_0[0]),.doutb(w_n19448_0[1]),.din(n19448));
	jspl jspl_w_n19449_0(.douta(w_n19449_0[0]),.doutb(w_n19449_0[1]),.din(n19449));
	jspl jspl_w_n19451_0(.douta(w_n19451_0[0]),.doutb(w_n19451_0[1]),.din(n19451));
	jspl jspl_w_n19453_0(.douta(w_n19453_0[0]),.doutb(w_n19453_0[1]),.din(n19453));
	jspl jspl_w_n19456_0(.douta(w_n19456_0[0]),.doutb(w_n19456_0[1]),.din(n19456));
	jspl jspl_w_n19462_0(.douta(w_n19462_0[0]),.doutb(w_n19462_0[1]),.din(n19462));
	jspl jspl_w_n19464_0(.douta(w_n19464_0[0]),.doutb(w_n19464_0[1]),.din(n19464));
	jspl3 jspl3_w_n19465_0(.douta(w_n19465_0[0]),.doutb(w_n19465_0[1]),.doutc(w_n19465_0[2]),.din(n19465));
	jspl jspl_w_n19469_0(.douta(w_n19469_0[0]),.doutb(w_n19469_0[1]),.din(n19469));
	jspl jspl_w_n19470_0(.douta(w_n19470_0[0]),.doutb(w_n19470_0[1]),.din(n19470));
	jspl3 jspl3_w_n19471_0(.douta(w_n19471_0[0]),.doutb(w_n19471_0[1]),.doutc(w_n19471_0[2]),.din(n19471));
	jspl jspl_w_n19473_0(.douta(w_n19473_0[0]),.doutb(w_n19473_0[1]),.din(n19473));
	jspl jspl_w_n19478_0(.douta(w_n19478_0[0]),.doutb(w_n19478_0[1]),.din(n19478));
	jspl jspl_w_n19480_0(.douta(w_n19480_0[0]),.doutb(w_n19480_0[1]),.din(n19480));
	jspl jspl_w_n19481_0(.douta(w_n19481_0[0]),.doutb(w_n19481_0[1]),.din(n19481));
	jspl3 jspl3_w_n19482_0(.douta(w_n19482_0[0]),.doutb(w_n19482_0[1]),.doutc(w_n19482_0[2]),.din(n19482));
	jspl jspl_w_n19483_0(.douta(w_n19483_0[0]),.doutb(w_n19483_0[1]),.din(n19483));
	jspl jspl_w_n19487_0(.douta(w_n19487_0[0]),.doutb(w_n19487_0[1]),.din(n19487));
	jspl jspl_w_n19493_0(.douta(w_n19493_0[0]),.doutb(w_n19493_0[1]),.din(n19493));
	jspl jspl_w_n19494_0(.douta(w_n19494_0[0]),.doutb(w_n19494_0[1]),.din(n19494));
	jspl jspl_w_n19496_0(.douta(w_n19496_0[0]),.doutb(w_n19496_0[1]),.din(n19496));
	jspl jspl_w_n19498_0(.douta(w_n19498_0[0]),.doutb(w_n19498_0[1]),.din(n19498));
	jspl jspl_w_n19501_0(.douta(w_n19501_0[0]),.doutb(w_n19501_0[1]),.din(n19501));
	jspl jspl_w_n19507_0(.douta(w_n19507_0[0]),.doutb(w_n19507_0[1]),.din(n19507));
	jspl jspl_w_n19509_0(.douta(w_n19509_0[0]),.doutb(w_n19509_0[1]),.din(n19509));
	jspl3 jspl3_w_n19510_0(.douta(w_n19510_0[0]),.doutb(w_n19510_0[1]),.doutc(w_n19510_0[2]),.din(n19510));
	jspl jspl_w_n19514_0(.douta(w_n19514_0[0]),.doutb(w_n19514_0[1]),.din(n19514));
	jspl jspl_w_n19515_0(.douta(w_n19515_0[0]),.doutb(w_n19515_0[1]),.din(n19515));
	jspl3 jspl3_w_n19516_0(.douta(w_n19516_0[0]),.doutb(w_n19516_0[1]),.doutc(w_n19516_0[2]),.din(n19516));
	jspl jspl_w_n19518_0(.douta(w_n19518_0[0]),.doutb(w_n19518_0[1]),.din(n19518));
	jspl jspl_w_n19523_0(.douta(w_n19523_0[0]),.doutb(w_n19523_0[1]),.din(n19523));
	jspl jspl_w_n19525_0(.douta(w_n19525_0[0]),.doutb(w_n19525_0[1]),.din(n19525));
	jspl jspl_w_n19526_0(.douta(w_n19526_0[0]),.doutb(w_n19526_0[1]),.din(n19526));
	jspl3 jspl3_w_n19527_0(.douta(w_n19527_0[0]),.doutb(w_n19527_0[1]),.doutc(w_n19527_0[2]),.din(n19527));
	jspl jspl_w_n19528_0(.douta(w_n19528_0[0]),.doutb(w_n19528_0[1]),.din(n19528));
	jspl jspl_w_n19532_0(.douta(w_n19532_0[0]),.doutb(w_n19532_0[1]),.din(n19532));
	jspl jspl_w_n19538_0(.douta(w_n19538_0[0]),.doutb(w_n19538_0[1]),.din(n19538));
	jspl jspl_w_n19539_0(.douta(w_n19539_0[0]),.doutb(w_n19539_0[1]),.din(n19539));
	jspl jspl_w_n19541_0(.douta(w_n19541_0[0]),.doutb(w_n19541_0[1]),.din(n19541));
	jspl jspl_w_n19546_0(.douta(w_n19546_0[0]),.doutb(w_n19546_0[1]),.din(n19546));
	jspl jspl_w_n19548_0(.douta(w_n19548_0[0]),.doutb(w_n19548_0[1]),.din(n19548));
	jspl jspl_w_n19549_0(.douta(w_n19549_0[0]),.doutb(w_n19549_0[1]),.din(n19549));
	jspl3 jspl3_w_n19550_0(.douta(w_n19550_0[0]),.doutb(w_n19550_0[1]),.doutc(w_n19550_0[2]),.din(n19550));
	jspl jspl_w_n19551_0(.douta(w_n19551_0[0]),.doutb(w_n19551_0[1]),.din(n19551));
	jspl jspl_w_n19553_0(.douta(w_n19553_0[0]),.doutb(w_n19553_0[1]),.din(n19553));
	jspl jspl_w_n19555_0(.douta(w_n19555_0[0]),.doutb(w_n19555_0[1]),.din(n19555));
	jspl jspl_w_n19557_0(.douta(w_n19557_0[0]),.doutb(w_n19557_0[1]),.din(n19557));
	jspl jspl_w_n19560_0(.douta(w_n19560_0[0]),.doutb(w_n19560_0[1]),.din(n19560));
	jspl jspl_w_n19566_0(.douta(w_n19566_0[0]),.doutb(w_n19566_0[1]),.din(n19566));
	jspl3 jspl3_w_n19568_0(.douta(w_n19568_0[0]),.doutb(w_n19568_0[1]),.doutc(w_n19568_0[2]),.din(n19568));
	jspl jspl_w_n19569_0(.douta(w_n19569_0[0]),.doutb(w_n19569_0[1]),.din(n19569));
	jspl jspl_w_n19573_0(.douta(w_n19573_0[0]),.doutb(w_n19573_0[1]),.din(n19573));
	jspl jspl_w_n19579_0(.douta(w_n19579_0[0]),.doutb(w_n19579_0[1]),.din(n19579));
	jspl jspl_w_n19580_0(.douta(w_n19580_0[0]),.doutb(w_n19580_0[1]),.din(n19580));
	jspl jspl_w_n19582_0(.douta(w_n19582_0[0]),.doutb(w_n19582_0[1]),.din(n19582));
	jspl jspl_w_n19584_0(.douta(w_n19584_0[0]),.doutb(w_n19584_0[1]),.din(n19584));
	jspl jspl_w_n19587_0(.douta(w_n19587_0[0]),.doutb(w_n19587_0[1]),.din(n19587));
	jspl jspl_w_n19593_0(.douta(w_n19593_0[0]),.doutb(w_n19593_0[1]),.din(n19593));
	jspl3 jspl3_w_n19595_0(.douta(w_n19595_0[0]),.doutb(w_n19595_0[1]),.doutc(w_n19595_0[2]),.din(n19595));
	jspl3 jspl3_w_n19595_1(.douta(w_n19595_1[0]),.doutb(w_n19595_1[1]),.doutc(w_n19595_1[2]),.din(w_n19595_0[0]));
	jspl jspl_w_n19598_0(.douta(w_n19598_0[0]),.doutb(w_n19598_0[1]),.din(n19598));
	jspl3 jspl3_w_n19599_0(.douta(w_n19599_0[0]),.doutb(w_n19599_0[1]),.doutc(w_n19599_0[2]),.din(n19599));
	jspl jspl_w_n19600_0(.douta(w_n19600_0[0]),.doutb(w_n19600_0[1]),.din(n19600));
	jspl3 jspl3_w_n19607_0(.douta(w_n19607_0[0]),.doutb(w_n19607_0[1]),.doutc(w_n19607_0[2]),.din(n19607));
	jspl jspl_w_n19608_0(.douta(w_n19608_0[0]),.doutb(w_n19608_0[1]),.din(n19608));
	jspl3 jspl3_w_n19616_0(.douta(w_n19616_0[0]),.doutb(w_n19616_0[1]),.doutc(w_n19616_0[2]),.din(n19616));
	jspl3 jspl3_w_n19616_1(.douta(w_n19616_1[0]),.doutb(w_n19616_1[1]),.doutc(w_n19616_1[2]),.din(w_n19616_0[0]));
	jspl3 jspl3_w_n19616_2(.douta(w_n19616_2[0]),.doutb(w_n19616_2[1]),.doutc(w_n19616_2[2]),.din(w_n19616_0[1]));
	jspl3 jspl3_w_n19616_3(.douta(w_n19616_3[0]),.doutb(w_n19616_3[1]),.doutc(w_n19616_3[2]),.din(w_n19616_0[2]));
	jspl3 jspl3_w_n19616_4(.douta(w_n19616_4[0]),.doutb(w_n19616_4[1]),.doutc(w_n19616_4[2]),.din(w_n19616_1[0]));
	jspl3 jspl3_w_n19616_5(.douta(w_n19616_5[0]),.doutb(w_n19616_5[1]),.doutc(w_n19616_5[2]),.din(w_n19616_1[1]));
	jspl3 jspl3_w_n19616_6(.douta(w_n19616_6[0]),.doutb(w_n19616_6[1]),.doutc(w_n19616_6[2]),.din(w_n19616_1[2]));
	jspl3 jspl3_w_n19616_7(.douta(w_n19616_7[0]),.doutb(w_n19616_7[1]),.doutc(w_n19616_7[2]),.din(w_n19616_2[0]));
	jspl3 jspl3_w_n19616_8(.douta(w_n19616_8[0]),.doutb(w_n19616_8[1]),.doutc(w_n19616_8[2]),.din(w_n19616_2[1]));
	jspl3 jspl3_w_n19616_9(.douta(w_n19616_9[0]),.doutb(w_n19616_9[1]),.doutc(w_n19616_9[2]),.din(w_n19616_2[2]));
	jspl3 jspl3_w_n19616_10(.douta(w_n19616_10[0]),.doutb(w_n19616_10[1]),.doutc(w_n19616_10[2]),.din(w_n19616_3[0]));
	jspl3 jspl3_w_n19616_11(.douta(w_n19616_11[0]),.doutb(w_n19616_11[1]),.doutc(w_n19616_11[2]),.din(w_n19616_3[1]));
	jspl3 jspl3_w_n19616_12(.douta(w_n19616_12[0]),.doutb(w_n19616_12[1]),.doutc(w_n19616_12[2]),.din(w_n19616_3[2]));
	jspl3 jspl3_w_n19616_13(.douta(w_n19616_13[0]),.doutb(w_n19616_13[1]),.doutc(w_n19616_13[2]),.din(w_n19616_4[0]));
	jspl3 jspl3_w_n19616_14(.douta(w_n19616_14[0]),.doutb(w_n19616_14[1]),.doutc(w_n19616_14[2]),.din(w_n19616_4[1]));
	jspl3 jspl3_w_n19616_15(.douta(w_n19616_15[0]),.doutb(w_n19616_15[1]),.doutc(w_n19616_15[2]),.din(w_n19616_4[2]));
	jspl3 jspl3_w_n19616_16(.douta(w_n19616_16[0]),.doutb(w_n19616_16[1]),.doutc(w_n19616_16[2]),.din(w_n19616_5[0]));
	jspl3 jspl3_w_n19616_17(.douta(w_n19616_17[0]),.doutb(w_n19616_17[1]),.doutc(w_n19616_17[2]),.din(w_n19616_5[1]));
	jspl3 jspl3_w_n19616_18(.douta(w_n19616_18[0]),.doutb(w_n19616_18[1]),.doutc(w_n19616_18[2]),.din(w_n19616_5[2]));
	jspl jspl_w_n19620_0(.douta(w_n19620_0[0]),.doutb(w_n19620_0[1]),.din(n19620));
	jspl3 jspl3_w_n19622_0(.douta(w_n19622_0[0]),.doutb(w_n19622_0[1]),.doutc(w_n19622_0[2]),.din(n19622));
	jspl jspl_w_n19622_1(.douta(w_n19622_1[0]),.doutb(w_n19622_1[1]),.din(w_n19622_0[0]));
	jspl3 jspl3_w_n19623_0(.douta(w_n19623_0[0]),.doutb(w_n19623_0[1]),.doutc(w_n19623_0[2]),.din(n19623));
	jspl3 jspl3_w_n19627_0(.douta(w_n19627_0[0]),.doutb(w_n19627_0[1]),.doutc(w_n19627_0[2]),.din(n19627));
	jspl jspl_w_n19628_0(.douta(w_n19628_0[0]),.doutb(w_n19628_0[1]),.din(n19628));
	jspl jspl_w_n19629_0(.douta(w_n19629_0[0]),.doutb(w_n19629_0[1]),.din(n19629));
	jspl jspl_w_n19630_0(.douta(w_n19630_0[0]),.doutb(w_n19630_0[1]),.din(n19630));
	jspl jspl_w_n19632_0(.douta(w_n19632_0[0]),.doutb(w_n19632_0[1]),.din(n19632));
	jspl jspl_w_n19634_0(.douta(w_n19634_0[0]),.doutb(w_n19634_0[1]),.din(n19634));
	jspl jspl_w_n19636_0(.douta(w_n19636_0[0]),.doutb(w_n19636_0[1]),.din(n19636));
	jspl jspl_w_n19641_0(.douta(w_n19641_0[0]),.doutb(w_n19641_0[1]),.din(n19641));
	jspl3 jspl3_w_n19643_0(.douta(w_n19643_0[0]),.doutb(w_n19643_0[1]),.doutc(w_n19643_0[2]),.din(n19643));
	jspl jspl_w_n19644_0(.douta(w_n19644_0[0]),.doutb(w_n19644_0[1]),.din(n19644));
	jspl jspl_w_n19648_0(.douta(w_n19648_0[0]),.doutb(w_n19648_0[1]),.din(n19648));
	jspl jspl_w_n19649_0(.douta(w_n19649_0[0]),.doutb(w_n19649_0[1]),.din(n19649));
	jspl jspl_w_n19651_0(.douta(w_n19651_0[0]),.doutb(w_n19651_0[1]),.din(n19651));
	jspl jspl_w_n19655_0(.douta(w_n19655_0[0]),.doutb(w_n19655_0[1]),.din(n19655));
	jspl jspl_w_n19657_0(.douta(w_n19657_0[0]),.doutb(w_n19657_0[1]),.din(n19657));
	jspl jspl_w_n19658_0(.douta(w_n19658_0[0]),.doutb(w_n19658_0[1]),.din(n19658));
	jspl3 jspl3_w_n19659_0(.douta(w_n19659_0[0]),.doutb(w_n19659_0[1]),.doutc(w_n19659_0[2]),.din(n19659));
	jspl jspl_w_n19660_0(.douta(w_n19660_0[0]),.doutb(w_n19660_0[1]),.din(n19660));
	jspl jspl_w_n19664_0(.douta(w_n19664_0[0]),.doutb(w_n19664_0[1]),.din(n19664));
	jspl jspl_w_n19666_0(.douta(w_n19666_0[0]),.doutb(w_n19666_0[1]),.din(n19666));
	jspl jspl_w_n19668_0(.douta(w_n19668_0[0]),.doutb(w_n19668_0[1]),.din(n19668));
	jspl jspl_w_n19670_0(.douta(w_n19670_0[0]),.doutb(w_n19670_0[1]),.din(n19670));
	jspl jspl_w_n19672_0(.douta(w_n19672_0[0]),.doutb(w_n19672_0[1]),.din(n19672));
	jspl jspl_w_n19678_0(.douta(w_n19678_0[0]),.doutb(w_n19678_0[1]),.din(n19678));
	jspl3 jspl3_w_n19680_0(.douta(w_n19680_0[0]),.doutb(w_n19680_0[1]),.doutc(w_n19680_0[2]),.din(n19680));
	jspl jspl_w_n19681_0(.douta(w_n19681_0[0]),.doutb(w_n19681_0[1]),.din(n19681));
	jspl jspl_w_n19686_0(.douta(w_n19686_0[0]),.doutb(w_n19686_0[1]),.din(n19686));
	jspl jspl_w_n19688_0(.douta(w_n19688_0[0]),.doutb(w_n19688_0[1]),.din(n19688));
	jspl jspl_w_n19690_0(.douta(w_n19690_0[0]),.doutb(w_n19690_0[1]),.din(n19690));
	jspl jspl_w_n19694_0(.douta(w_n19694_0[0]),.doutb(w_n19694_0[1]),.din(n19694));
	jspl jspl_w_n19696_0(.douta(w_n19696_0[0]),.doutb(w_n19696_0[1]),.din(n19696));
	jspl jspl_w_n19697_0(.douta(w_n19697_0[0]),.doutb(w_n19697_0[1]),.din(n19697));
	jspl3 jspl3_w_n19698_0(.douta(w_n19698_0[0]),.doutb(w_n19698_0[1]),.doutc(w_n19698_0[2]),.din(n19698));
	jspl jspl_w_n19699_0(.douta(w_n19699_0[0]),.doutb(w_n19699_0[1]),.din(n19699));
	jspl jspl_w_n19705_0(.douta(w_n19705_0[0]),.doutb(w_n19705_0[1]),.din(n19705));
	jspl jspl_w_n19706_0(.douta(w_n19706_0[0]),.doutb(w_n19706_0[1]),.din(n19706));
	jspl jspl_w_n19708_0(.douta(w_n19708_0[0]),.doutb(w_n19708_0[1]),.din(n19708));
	jspl jspl_w_n19710_0(.douta(w_n19710_0[0]),.doutb(w_n19710_0[1]),.din(n19710));
	jspl jspl_w_n19712_0(.douta(w_n19712_0[0]),.doutb(w_n19712_0[1]),.din(n19712));
	jspl jspl_w_n19718_0(.douta(w_n19718_0[0]),.doutb(w_n19718_0[1]),.din(n19718));
	jspl jspl_w_n19720_0(.douta(w_n19720_0[0]),.doutb(w_n19720_0[1]),.din(n19720));
	jspl3 jspl3_w_n19721_0(.douta(w_n19721_0[0]),.doutb(w_n19721_0[1]),.doutc(w_n19721_0[2]),.din(n19721));
	jspl jspl_w_n19724_0(.douta(w_n19724_0[0]),.doutb(w_n19724_0[1]),.din(n19724));
	jspl jspl_w_n19725_0(.douta(w_n19725_0[0]),.doutb(w_n19725_0[1]),.din(n19725));
	jspl3 jspl3_w_n19726_0(.douta(w_n19726_0[0]),.doutb(w_n19726_0[1]),.doutc(w_n19726_0[2]),.din(n19726));
	jspl jspl_w_n19728_0(.douta(w_n19728_0[0]),.doutb(w_n19728_0[1]),.din(n19728));
	jspl jspl_w_n19732_0(.douta(w_n19732_0[0]),.doutb(w_n19732_0[1]),.din(n19732));
	jspl jspl_w_n19734_0(.douta(w_n19734_0[0]),.doutb(w_n19734_0[1]),.din(n19734));
	jspl jspl_w_n19735_0(.douta(w_n19735_0[0]),.doutb(w_n19735_0[1]),.din(n19735));
	jspl3 jspl3_w_n19736_0(.douta(w_n19736_0[0]),.doutb(w_n19736_0[1]),.doutc(w_n19736_0[2]),.din(n19736));
	jspl jspl_w_n19737_0(.douta(w_n19737_0[0]),.doutb(w_n19737_0[1]),.din(n19737));
	jspl jspl_w_n19740_0(.douta(w_n19740_0[0]),.doutb(w_n19740_0[1]),.din(n19740));
	jspl jspl_w_n19746_0(.douta(w_n19746_0[0]),.doutb(w_n19746_0[1]),.din(n19746));
	jspl jspl_w_n19747_0(.douta(w_n19747_0[0]),.doutb(w_n19747_0[1]),.din(n19747));
	jspl jspl_w_n19749_0(.douta(w_n19749_0[0]),.doutb(w_n19749_0[1]),.din(n19749));
	jspl jspl_w_n19751_0(.douta(w_n19751_0[0]),.doutb(w_n19751_0[1]),.din(n19751));
	jspl jspl_w_n19753_0(.douta(w_n19753_0[0]),.doutb(w_n19753_0[1]),.din(n19753));
	jspl jspl_w_n19759_0(.douta(w_n19759_0[0]),.doutb(w_n19759_0[1]),.din(n19759));
	jspl jspl_w_n19761_0(.douta(w_n19761_0[0]),.doutb(w_n19761_0[1]),.din(n19761));
	jspl3 jspl3_w_n19762_0(.douta(w_n19762_0[0]),.doutb(w_n19762_0[1]),.doutc(w_n19762_0[2]),.din(n19762));
	jspl jspl_w_n19765_0(.douta(w_n19765_0[0]),.doutb(w_n19765_0[1]),.din(n19765));
	jspl jspl_w_n19766_0(.douta(w_n19766_0[0]),.doutb(w_n19766_0[1]),.din(n19766));
	jspl3 jspl3_w_n19767_0(.douta(w_n19767_0[0]),.doutb(w_n19767_0[1]),.doutc(w_n19767_0[2]),.din(n19767));
	jspl jspl_w_n19769_0(.douta(w_n19769_0[0]),.doutb(w_n19769_0[1]),.din(n19769));
	jspl jspl_w_n19773_0(.douta(w_n19773_0[0]),.doutb(w_n19773_0[1]),.din(n19773));
	jspl jspl_w_n19775_0(.douta(w_n19775_0[0]),.doutb(w_n19775_0[1]),.din(n19775));
	jspl jspl_w_n19776_0(.douta(w_n19776_0[0]),.doutb(w_n19776_0[1]),.din(n19776));
	jspl3 jspl3_w_n19777_0(.douta(w_n19777_0[0]),.doutb(w_n19777_0[1]),.doutc(w_n19777_0[2]),.din(n19777));
	jspl jspl_w_n19778_0(.douta(w_n19778_0[0]),.doutb(w_n19778_0[1]),.din(n19778));
	jspl jspl_w_n19781_0(.douta(w_n19781_0[0]),.doutb(w_n19781_0[1]),.din(n19781));
	jspl jspl_w_n19787_0(.douta(w_n19787_0[0]),.doutb(w_n19787_0[1]),.din(n19787));
	jspl jspl_w_n19788_0(.douta(w_n19788_0[0]),.doutb(w_n19788_0[1]),.din(n19788));
	jspl jspl_w_n19790_0(.douta(w_n19790_0[0]),.doutb(w_n19790_0[1]),.din(n19790));
	jspl jspl_w_n19792_0(.douta(w_n19792_0[0]),.doutb(w_n19792_0[1]),.din(n19792));
	jspl jspl_w_n19794_0(.douta(w_n19794_0[0]),.doutb(w_n19794_0[1]),.din(n19794));
	jspl jspl_w_n19800_0(.douta(w_n19800_0[0]),.doutb(w_n19800_0[1]),.din(n19800));
	jspl jspl_w_n19802_0(.douta(w_n19802_0[0]),.doutb(w_n19802_0[1]),.din(n19802));
	jspl3 jspl3_w_n19803_0(.douta(w_n19803_0[0]),.doutb(w_n19803_0[1]),.doutc(w_n19803_0[2]),.din(n19803));
	jspl jspl_w_n19806_0(.douta(w_n19806_0[0]),.doutb(w_n19806_0[1]),.din(n19806));
	jspl jspl_w_n19807_0(.douta(w_n19807_0[0]),.doutb(w_n19807_0[1]),.din(n19807));
	jspl3 jspl3_w_n19808_0(.douta(w_n19808_0[0]),.doutb(w_n19808_0[1]),.doutc(w_n19808_0[2]),.din(n19808));
	jspl jspl_w_n19810_0(.douta(w_n19810_0[0]),.doutb(w_n19810_0[1]),.din(n19810));
	jspl jspl_w_n19814_0(.douta(w_n19814_0[0]),.doutb(w_n19814_0[1]),.din(n19814));
	jspl jspl_w_n19816_0(.douta(w_n19816_0[0]),.doutb(w_n19816_0[1]),.din(n19816));
	jspl jspl_w_n19817_0(.douta(w_n19817_0[0]),.doutb(w_n19817_0[1]),.din(n19817));
	jspl3 jspl3_w_n19818_0(.douta(w_n19818_0[0]),.doutb(w_n19818_0[1]),.doutc(w_n19818_0[2]),.din(n19818));
	jspl jspl_w_n19819_0(.douta(w_n19819_0[0]),.doutb(w_n19819_0[1]),.din(n19819));
	jspl jspl_w_n19822_0(.douta(w_n19822_0[0]),.doutb(w_n19822_0[1]),.din(n19822));
	jspl jspl_w_n19828_0(.douta(w_n19828_0[0]),.doutb(w_n19828_0[1]),.din(n19828));
	jspl jspl_w_n19829_0(.douta(w_n19829_0[0]),.doutb(w_n19829_0[1]),.din(n19829));
	jspl jspl_w_n19831_0(.douta(w_n19831_0[0]),.doutb(w_n19831_0[1]),.din(n19831));
	jspl jspl_w_n19833_0(.douta(w_n19833_0[0]),.doutb(w_n19833_0[1]),.din(n19833));
	jspl jspl_w_n19835_0(.douta(w_n19835_0[0]),.doutb(w_n19835_0[1]),.din(n19835));
	jspl jspl_w_n19841_0(.douta(w_n19841_0[0]),.doutb(w_n19841_0[1]),.din(n19841));
	jspl jspl_w_n19843_0(.douta(w_n19843_0[0]),.doutb(w_n19843_0[1]),.din(n19843));
	jspl3 jspl3_w_n19844_0(.douta(w_n19844_0[0]),.doutb(w_n19844_0[1]),.doutc(w_n19844_0[2]),.din(n19844));
	jspl jspl_w_n19847_0(.douta(w_n19847_0[0]),.doutb(w_n19847_0[1]),.din(n19847));
	jspl jspl_w_n19848_0(.douta(w_n19848_0[0]),.doutb(w_n19848_0[1]),.din(n19848));
	jspl3 jspl3_w_n19849_0(.douta(w_n19849_0[0]),.doutb(w_n19849_0[1]),.doutc(w_n19849_0[2]),.din(n19849));
	jspl jspl_w_n19851_0(.douta(w_n19851_0[0]),.doutb(w_n19851_0[1]),.din(n19851));
	jspl jspl_w_n19855_0(.douta(w_n19855_0[0]),.doutb(w_n19855_0[1]),.din(n19855));
	jspl jspl_w_n19857_0(.douta(w_n19857_0[0]),.doutb(w_n19857_0[1]),.din(n19857));
	jspl jspl_w_n19858_0(.douta(w_n19858_0[0]),.doutb(w_n19858_0[1]),.din(n19858));
	jspl3 jspl3_w_n19859_0(.douta(w_n19859_0[0]),.doutb(w_n19859_0[1]),.doutc(w_n19859_0[2]),.din(n19859));
	jspl jspl_w_n19860_0(.douta(w_n19860_0[0]),.doutb(w_n19860_0[1]),.din(n19860));
	jspl jspl_w_n19863_0(.douta(w_n19863_0[0]),.doutb(w_n19863_0[1]),.din(n19863));
	jspl jspl_w_n19869_0(.douta(w_n19869_0[0]),.doutb(w_n19869_0[1]),.din(n19869));
	jspl jspl_w_n19870_0(.douta(w_n19870_0[0]),.doutb(w_n19870_0[1]),.din(n19870));
	jspl jspl_w_n19872_0(.douta(w_n19872_0[0]),.doutb(w_n19872_0[1]),.din(n19872));
	jspl jspl_w_n19874_0(.douta(w_n19874_0[0]),.doutb(w_n19874_0[1]),.din(n19874));
	jspl jspl_w_n19876_0(.douta(w_n19876_0[0]),.doutb(w_n19876_0[1]),.din(n19876));
	jspl jspl_w_n19882_0(.douta(w_n19882_0[0]),.doutb(w_n19882_0[1]),.din(n19882));
	jspl jspl_w_n19884_0(.douta(w_n19884_0[0]),.doutb(w_n19884_0[1]),.din(n19884));
	jspl3 jspl3_w_n19885_0(.douta(w_n19885_0[0]),.doutb(w_n19885_0[1]),.doutc(w_n19885_0[2]),.din(n19885));
	jspl jspl_w_n19888_0(.douta(w_n19888_0[0]),.doutb(w_n19888_0[1]),.din(n19888));
	jspl jspl_w_n19889_0(.douta(w_n19889_0[0]),.doutb(w_n19889_0[1]),.din(n19889));
	jspl3 jspl3_w_n19890_0(.douta(w_n19890_0[0]),.doutb(w_n19890_0[1]),.doutc(w_n19890_0[2]),.din(n19890));
	jspl jspl_w_n19892_0(.douta(w_n19892_0[0]),.doutb(w_n19892_0[1]),.din(n19892));
	jspl jspl_w_n19896_0(.douta(w_n19896_0[0]),.doutb(w_n19896_0[1]),.din(n19896));
	jspl jspl_w_n19898_0(.douta(w_n19898_0[0]),.doutb(w_n19898_0[1]),.din(n19898));
	jspl jspl_w_n19899_0(.douta(w_n19899_0[0]),.doutb(w_n19899_0[1]),.din(n19899));
	jspl3 jspl3_w_n19900_0(.douta(w_n19900_0[0]),.doutb(w_n19900_0[1]),.doutc(w_n19900_0[2]),.din(n19900));
	jspl jspl_w_n19901_0(.douta(w_n19901_0[0]),.doutb(w_n19901_0[1]),.din(n19901));
	jspl jspl_w_n19904_0(.douta(w_n19904_0[0]),.doutb(w_n19904_0[1]),.din(n19904));
	jspl jspl_w_n19910_0(.douta(w_n19910_0[0]),.doutb(w_n19910_0[1]),.din(n19910));
	jspl jspl_w_n19911_0(.douta(w_n19911_0[0]),.doutb(w_n19911_0[1]),.din(n19911));
	jspl jspl_w_n19913_0(.douta(w_n19913_0[0]),.doutb(w_n19913_0[1]),.din(n19913));
	jspl jspl_w_n19915_0(.douta(w_n19915_0[0]),.doutb(w_n19915_0[1]),.din(n19915));
	jspl jspl_w_n19917_0(.douta(w_n19917_0[0]),.doutb(w_n19917_0[1]),.din(n19917));
	jspl jspl_w_n19923_0(.douta(w_n19923_0[0]),.doutb(w_n19923_0[1]),.din(n19923));
	jspl jspl_w_n19925_0(.douta(w_n19925_0[0]),.doutb(w_n19925_0[1]),.din(n19925));
	jspl3 jspl3_w_n19926_0(.douta(w_n19926_0[0]),.doutb(w_n19926_0[1]),.doutc(w_n19926_0[2]),.din(n19926));
	jspl jspl_w_n19929_0(.douta(w_n19929_0[0]),.doutb(w_n19929_0[1]),.din(n19929));
	jspl jspl_w_n19930_0(.douta(w_n19930_0[0]),.doutb(w_n19930_0[1]),.din(n19930));
	jspl3 jspl3_w_n19931_0(.douta(w_n19931_0[0]),.doutb(w_n19931_0[1]),.doutc(w_n19931_0[2]),.din(n19931));
	jspl jspl_w_n19933_0(.douta(w_n19933_0[0]),.doutb(w_n19933_0[1]),.din(n19933));
	jspl jspl_w_n19937_0(.douta(w_n19937_0[0]),.doutb(w_n19937_0[1]),.din(n19937));
	jspl jspl_w_n19939_0(.douta(w_n19939_0[0]),.doutb(w_n19939_0[1]),.din(n19939));
	jspl jspl_w_n19940_0(.douta(w_n19940_0[0]),.doutb(w_n19940_0[1]),.din(n19940));
	jspl3 jspl3_w_n19941_0(.douta(w_n19941_0[0]),.doutb(w_n19941_0[1]),.doutc(w_n19941_0[2]),.din(n19941));
	jspl jspl_w_n19942_0(.douta(w_n19942_0[0]),.doutb(w_n19942_0[1]),.din(n19942));
	jspl jspl_w_n19945_0(.douta(w_n19945_0[0]),.doutb(w_n19945_0[1]),.din(n19945));
	jspl jspl_w_n19951_0(.douta(w_n19951_0[0]),.doutb(w_n19951_0[1]),.din(n19951));
	jspl jspl_w_n19952_0(.douta(w_n19952_0[0]),.doutb(w_n19952_0[1]),.din(n19952));
	jspl jspl_w_n19954_0(.douta(w_n19954_0[0]),.doutb(w_n19954_0[1]),.din(n19954));
	jspl jspl_w_n19956_0(.douta(w_n19956_0[0]),.doutb(w_n19956_0[1]),.din(n19956));
	jspl jspl_w_n19958_0(.douta(w_n19958_0[0]),.doutb(w_n19958_0[1]),.din(n19958));
	jspl jspl_w_n19964_0(.douta(w_n19964_0[0]),.doutb(w_n19964_0[1]),.din(n19964));
	jspl jspl_w_n19966_0(.douta(w_n19966_0[0]),.doutb(w_n19966_0[1]),.din(n19966));
	jspl3 jspl3_w_n19967_0(.douta(w_n19967_0[0]),.doutb(w_n19967_0[1]),.doutc(w_n19967_0[2]),.din(n19967));
	jspl jspl_w_n19970_0(.douta(w_n19970_0[0]),.doutb(w_n19970_0[1]),.din(n19970));
	jspl jspl_w_n19971_0(.douta(w_n19971_0[0]),.doutb(w_n19971_0[1]),.din(n19971));
	jspl3 jspl3_w_n19972_0(.douta(w_n19972_0[0]),.doutb(w_n19972_0[1]),.doutc(w_n19972_0[2]),.din(n19972));
	jspl jspl_w_n19974_0(.douta(w_n19974_0[0]),.doutb(w_n19974_0[1]),.din(n19974));
	jspl jspl_w_n19978_0(.douta(w_n19978_0[0]),.doutb(w_n19978_0[1]),.din(n19978));
	jspl jspl_w_n19980_0(.douta(w_n19980_0[0]),.doutb(w_n19980_0[1]),.din(n19980));
	jspl jspl_w_n19981_0(.douta(w_n19981_0[0]),.doutb(w_n19981_0[1]),.din(n19981));
	jspl3 jspl3_w_n19982_0(.douta(w_n19982_0[0]),.doutb(w_n19982_0[1]),.doutc(w_n19982_0[2]),.din(n19982));
	jspl jspl_w_n19983_0(.douta(w_n19983_0[0]),.doutb(w_n19983_0[1]),.din(n19983));
	jspl jspl_w_n19986_0(.douta(w_n19986_0[0]),.doutb(w_n19986_0[1]),.din(n19986));
	jspl jspl_w_n19992_0(.douta(w_n19992_0[0]),.doutb(w_n19992_0[1]),.din(n19992));
	jspl jspl_w_n19993_0(.douta(w_n19993_0[0]),.doutb(w_n19993_0[1]),.din(n19993));
	jspl jspl_w_n19995_0(.douta(w_n19995_0[0]),.doutb(w_n19995_0[1]),.din(n19995));
	jspl jspl_w_n19997_0(.douta(w_n19997_0[0]),.doutb(w_n19997_0[1]),.din(n19997));
	jspl jspl_w_n19999_0(.douta(w_n19999_0[0]),.doutb(w_n19999_0[1]),.din(n19999));
	jspl jspl_w_n20005_0(.douta(w_n20005_0[0]),.doutb(w_n20005_0[1]),.din(n20005));
	jspl jspl_w_n20007_0(.douta(w_n20007_0[0]),.doutb(w_n20007_0[1]),.din(n20007));
	jspl3 jspl3_w_n20008_0(.douta(w_n20008_0[0]),.doutb(w_n20008_0[1]),.doutc(w_n20008_0[2]),.din(n20008));
	jspl jspl_w_n20011_0(.douta(w_n20011_0[0]),.doutb(w_n20011_0[1]),.din(n20011));
	jspl jspl_w_n20012_0(.douta(w_n20012_0[0]),.doutb(w_n20012_0[1]),.din(n20012));
	jspl3 jspl3_w_n20013_0(.douta(w_n20013_0[0]),.doutb(w_n20013_0[1]),.doutc(w_n20013_0[2]),.din(n20013));
	jspl jspl_w_n20015_0(.douta(w_n20015_0[0]),.doutb(w_n20015_0[1]),.din(n20015));
	jspl jspl_w_n20019_0(.douta(w_n20019_0[0]),.doutb(w_n20019_0[1]),.din(n20019));
	jspl jspl_w_n20021_0(.douta(w_n20021_0[0]),.doutb(w_n20021_0[1]),.din(n20021));
	jspl jspl_w_n20022_0(.douta(w_n20022_0[0]),.doutb(w_n20022_0[1]),.din(n20022));
	jspl3 jspl3_w_n20023_0(.douta(w_n20023_0[0]),.doutb(w_n20023_0[1]),.doutc(w_n20023_0[2]),.din(n20023));
	jspl jspl_w_n20024_0(.douta(w_n20024_0[0]),.doutb(w_n20024_0[1]),.din(n20024));
	jspl jspl_w_n20027_0(.douta(w_n20027_0[0]),.doutb(w_n20027_0[1]),.din(n20027));
	jspl jspl_w_n20033_0(.douta(w_n20033_0[0]),.doutb(w_n20033_0[1]),.din(n20033));
	jspl jspl_w_n20034_0(.douta(w_n20034_0[0]),.doutb(w_n20034_0[1]),.din(n20034));
	jspl jspl_w_n20036_0(.douta(w_n20036_0[0]),.doutb(w_n20036_0[1]),.din(n20036));
	jspl jspl_w_n20038_0(.douta(w_n20038_0[0]),.doutb(w_n20038_0[1]),.din(n20038));
	jspl jspl_w_n20040_0(.douta(w_n20040_0[0]),.doutb(w_n20040_0[1]),.din(n20040));
	jspl jspl_w_n20046_0(.douta(w_n20046_0[0]),.doutb(w_n20046_0[1]),.din(n20046));
	jspl jspl_w_n20048_0(.douta(w_n20048_0[0]),.doutb(w_n20048_0[1]),.din(n20048));
	jspl3 jspl3_w_n20049_0(.douta(w_n20049_0[0]),.doutb(w_n20049_0[1]),.doutc(w_n20049_0[2]),.din(n20049));
	jspl jspl_w_n20052_0(.douta(w_n20052_0[0]),.doutb(w_n20052_0[1]),.din(n20052));
	jspl jspl_w_n20053_0(.douta(w_n20053_0[0]),.doutb(w_n20053_0[1]),.din(n20053));
	jspl3 jspl3_w_n20054_0(.douta(w_n20054_0[0]),.doutb(w_n20054_0[1]),.doutc(w_n20054_0[2]),.din(n20054));
	jspl jspl_w_n20056_0(.douta(w_n20056_0[0]),.doutb(w_n20056_0[1]),.din(n20056));
	jspl jspl_w_n20060_0(.douta(w_n20060_0[0]),.doutb(w_n20060_0[1]),.din(n20060));
	jspl jspl_w_n20062_0(.douta(w_n20062_0[0]),.doutb(w_n20062_0[1]),.din(n20062));
	jspl jspl_w_n20063_0(.douta(w_n20063_0[0]),.doutb(w_n20063_0[1]),.din(n20063));
	jspl3 jspl3_w_n20064_0(.douta(w_n20064_0[0]),.doutb(w_n20064_0[1]),.doutc(w_n20064_0[2]),.din(n20064));
	jspl jspl_w_n20065_0(.douta(w_n20065_0[0]),.doutb(w_n20065_0[1]),.din(n20065));
	jspl jspl_w_n20068_0(.douta(w_n20068_0[0]),.doutb(w_n20068_0[1]),.din(n20068));
	jspl jspl_w_n20074_0(.douta(w_n20074_0[0]),.doutb(w_n20074_0[1]),.din(n20074));
	jspl jspl_w_n20075_0(.douta(w_n20075_0[0]),.doutb(w_n20075_0[1]),.din(n20075));
	jspl jspl_w_n20077_0(.douta(w_n20077_0[0]),.doutb(w_n20077_0[1]),.din(n20077));
	jspl jspl_w_n20079_0(.douta(w_n20079_0[0]),.doutb(w_n20079_0[1]),.din(n20079));
	jspl jspl_w_n20081_0(.douta(w_n20081_0[0]),.doutb(w_n20081_0[1]),.din(n20081));
	jspl jspl_w_n20087_0(.douta(w_n20087_0[0]),.doutb(w_n20087_0[1]),.din(n20087));
	jspl jspl_w_n20089_0(.douta(w_n20089_0[0]),.doutb(w_n20089_0[1]),.din(n20089));
	jspl3 jspl3_w_n20090_0(.douta(w_n20090_0[0]),.doutb(w_n20090_0[1]),.doutc(w_n20090_0[2]),.din(n20090));
	jspl jspl_w_n20093_0(.douta(w_n20093_0[0]),.doutb(w_n20093_0[1]),.din(n20093));
	jspl jspl_w_n20094_0(.douta(w_n20094_0[0]),.doutb(w_n20094_0[1]),.din(n20094));
	jspl3 jspl3_w_n20095_0(.douta(w_n20095_0[0]),.doutb(w_n20095_0[1]),.doutc(w_n20095_0[2]),.din(n20095));
	jspl jspl_w_n20097_0(.douta(w_n20097_0[0]),.doutb(w_n20097_0[1]),.din(n20097));
	jspl jspl_w_n20101_0(.douta(w_n20101_0[0]),.doutb(w_n20101_0[1]),.din(n20101));
	jspl jspl_w_n20103_0(.douta(w_n20103_0[0]),.doutb(w_n20103_0[1]),.din(n20103));
	jspl jspl_w_n20104_0(.douta(w_n20104_0[0]),.doutb(w_n20104_0[1]),.din(n20104));
	jspl3 jspl3_w_n20105_0(.douta(w_n20105_0[0]),.doutb(w_n20105_0[1]),.doutc(w_n20105_0[2]),.din(n20105));
	jspl jspl_w_n20106_0(.douta(w_n20106_0[0]),.doutb(w_n20106_0[1]),.din(n20106));
	jspl jspl_w_n20109_0(.douta(w_n20109_0[0]),.doutb(w_n20109_0[1]),.din(n20109));
	jspl jspl_w_n20115_0(.douta(w_n20115_0[0]),.doutb(w_n20115_0[1]),.din(n20115));
	jspl jspl_w_n20116_0(.douta(w_n20116_0[0]),.doutb(w_n20116_0[1]),.din(n20116));
	jspl jspl_w_n20118_0(.douta(w_n20118_0[0]),.doutb(w_n20118_0[1]),.din(n20118));
	jspl jspl_w_n20120_0(.douta(w_n20120_0[0]),.doutb(w_n20120_0[1]),.din(n20120));
	jspl jspl_w_n20122_0(.douta(w_n20122_0[0]),.doutb(w_n20122_0[1]),.din(n20122));
	jspl jspl_w_n20128_0(.douta(w_n20128_0[0]),.doutb(w_n20128_0[1]),.din(n20128));
	jspl jspl_w_n20130_0(.douta(w_n20130_0[0]),.doutb(w_n20130_0[1]),.din(n20130));
	jspl3 jspl3_w_n20131_0(.douta(w_n20131_0[0]),.doutb(w_n20131_0[1]),.doutc(w_n20131_0[2]),.din(n20131));
	jspl jspl_w_n20134_0(.douta(w_n20134_0[0]),.doutb(w_n20134_0[1]),.din(n20134));
	jspl jspl_w_n20135_0(.douta(w_n20135_0[0]),.doutb(w_n20135_0[1]),.din(n20135));
	jspl3 jspl3_w_n20136_0(.douta(w_n20136_0[0]),.doutb(w_n20136_0[1]),.doutc(w_n20136_0[2]),.din(n20136));
	jspl jspl_w_n20138_0(.douta(w_n20138_0[0]),.doutb(w_n20138_0[1]),.din(n20138));
	jspl jspl_w_n20142_0(.douta(w_n20142_0[0]),.doutb(w_n20142_0[1]),.din(n20142));
	jspl jspl_w_n20144_0(.douta(w_n20144_0[0]),.doutb(w_n20144_0[1]),.din(n20144));
	jspl jspl_w_n20145_0(.douta(w_n20145_0[0]),.doutb(w_n20145_0[1]),.din(n20145));
	jspl3 jspl3_w_n20146_0(.douta(w_n20146_0[0]),.doutb(w_n20146_0[1]),.doutc(w_n20146_0[2]),.din(n20146));
	jspl jspl_w_n20147_0(.douta(w_n20147_0[0]),.doutb(w_n20147_0[1]),.din(n20147));
	jspl jspl_w_n20150_0(.douta(w_n20150_0[0]),.doutb(w_n20150_0[1]),.din(n20150));
	jspl jspl_w_n20156_0(.douta(w_n20156_0[0]),.doutb(w_n20156_0[1]),.din(n20156));
	jspl jspl_w_n20157_0(.douta(w_n20157_0[0]),.doutb(w_n20157_0[1]),.din(n20157));
	jspl jspl_w_n20159_0(.douta(w_n20159_0[0]),.doutb(w_n20159_0[1]),.din(n20159));
	jspl jspl_w_n20161_0(.douta(w_n20161_0[0]),.doutb(w_n20161_0[1]),.din(n20161));
	jspl jspl_w_n20163_0(.douta(w_n20163_0[0]),.doutb(w_n20163_0[1]),.din(n20163));
	jspl jspl_w_n20169_0(.douta(w_n20169_0[0]),.doutb(w_n20169_0[1]),.din(n20169));
	jspl jspl_w_n20171_0(.douta(w_n20171_0[0]),.doutb(w_n20171_0[1]),.din(n20171));
	jspl3 jspl3_w_n20172_0(.douta(w_n20172_0[0]),.doutb(w_n20172_0[1]),.doutc(w_n20172_0[2]),.din(n20172));
	jspl jspl_w_n20175_0(.douta(w_n20175_0[0]),.doutb(w_n20175_0[1]),.din(n20175));
	jspl jspl_w_n20176_0(.douta(w_n20176_0[0]),.doutb(w_n20176_0[1]),.din(n20176));
	jspl3 jspl3_w_n20177_0(.douta(w_n20177_0[0]),.doutb(w_n20177_0[1]),.doutc(w_n20177_0[2]),.din(n20177));
	jspl jspl_w_n20179_0(.douta(w_n20179_0[0]),.doutb(w_n20179_0[1]),.din(n20179));
	jspl jspl_w_n20181_0(.douta(w_n20181_0[0]),.doutb(w_n20181_0[1]),.din(n20181));
	jspl jspl_w_n20183_0(.douta(w_n20183_0[0]),.doutb(w_n20183_0[1]),.din(n20183));
	jspl jspl_w_n20189_0(.douta(w_n20189_0[0]),.doutb(w_n20189_0[1]),.din(n20189));
	jspl3 jspl3_w_n20191_0(.douta(w_n20191_0[0]),.doutb(w_n20191_0[1]),.doutc(w_n20191_0[2]),.din(n20191));
	jspl jspl_w_n20192_0(.douta(w_n20192_0[0]),.doutb(w_n20192_0[1]),.din(n20192));
	jspl jspl_w_n20194_0(.douta(w_n20194_0[0]),.doutb(w_n20194_0[1]),.din(n20194));
	jspl jspl_w_n20196_0(.douta(w_n20196_0[0]),.doutb(w_n20196_0[1]),.din(n20196));
	jspl jspl_w_n20200_0(.douta(w_n20200_0[0]),.doutb(w_n20200_0[1]),.din(n20200));
	jspl jspl_w_n20202_0(.douta(w_n20202_0[0]),.doutb(w_n20202_0[1]),.din(n20202));
	jspl jspl_w_n20203_0(.douta(w_n20203_0[0]),.doutb(w_n20203_0[1]),.din(n20203));
	jspl3 jspl3_w_n20204_0(.douta(w_n20204_0[0]),.doutb(w_n20204_0[1]),.doutc(w_n20204_0[2]),.din(n20204));
	jspl jspl_w_n20209_0(.douta(w_n20209_0[0]),.doutb(w_n20209_0[1]),.din(n20209));
	jspl3 jspl3_w_n20211_0(.douta(w_n20211_0[0]),.doutb(w_n20211_0[1]),.doutc(w_n20211_0[2]),.din(n20211));
	jspl3 jspl3_w_n20215_0(.douta(w_n20215_0[0]),.doutb(w_n20215_0[1]),.doutc(w_n20215_0[2]),.din(n20215));
	jspl jspl_w_n20217_0(.douta(w_n20217_0[0]),.doutb(w_n20217_0[1]),.din(n20217));
	jspl jspl_w_n20223_0(.douta(w_n20223_0[0]),.doutb(w_n20223_0[1]),.din(n20223));
	jspl jspl_w_n20234_0(.douta(w_n20234_0[0]),.doutb(w_n20234_0[1]),.din(n20234));
	jspl jspl_w_n20236_0(.douta(w_n20236_0[0]),.doutb(w_n20236_0[1]),.din(n20236));
	jspl jspl_w_n20237_0(.douta(w_n20237_0[0]),.doutb(w_n20237_0[1]),.din(n20237));
	jspl3 jspl3_w_n20240_0(.douta(w_n20240_0[0]),.doutb(w_n20240_0[1]),.doutc(w_n20240_0[2]),.din(n20240));
	jspl jspl_w_n20241_0(.douta(w_n20241_0[0]),.doutb(w_n20241_0[1]),.din(n20241));
	jspl jspl_w_n20242_0(.douta(w_n20242_0[0]),.doutb(w_n20242_0[1]),.din(n20242));
	jspl jspl_w_n20243_0(.douta(w_n20243_0[0]),.doutb(w_n20243_0[1]),.din(n20243));
	jspl jspl_w_n20245_0(.douta(w_n20245_0[0]),.doutb(w_n20245_0[1]),.din(n20245));
	jspl jspl_w_n20247_0(.douta(w_n20247_0[0]),.doutb(w_n20247_0[1]),.din(n20247));
	jspl jspl_w_n20249_0(.douta(w_n20249_0[0]),.doutb(w_n20249_0[1]),.din(n20249));
	jspl3 jspl3_w_n20251_0(.douta(w_n20251_0[0]),.doutb(w_n20251_0[1]),.doutc(w_n20251_0[2]),.din(n20251));
	jspl jspl_w_n20251_1(.douta(w_n20251_1[0]),.doutb(w_n20251_1[1]),.din(w_n20251_0[0]));
	jspl jspl_w_n20254_0(.douta(w_n20254_0[0]),.doutb(w_n20254_0[1]),.din(n20254));
	jspl3 jspl3_w_n20256_0(.douta(w_n20256_0[0]),.doutb(w_n20256_0[1]),.doutc(w_n20256_0[2]),.din(n20256));
	jspl jspl_w_n20257_0(.douta(w_n20257_0[0]),.doutb(w_n20257_0[1]),.din(n20257));
	jspl jspl_w_n20262_0(.douta(w_n20262_0[0]),.doutb(w_n20262_0[1]),.din(n20262));
	jspl jspl_w_n20263_0(.douta(w_n20263_0[0]),.doutb(w_n20263_0[1]),.din(n20263));
	jspl jspl_w_n20265_0(.douta(w_n20265_0[0]),.doutb(w_n20265_0[1]),.din(n20265));
	jspl jspl_w_n20269_0(.douta(w_n20269_0[0]),.doutb(w_n20269_0[1]),.din(n20269));
	jspl jspl_w_n20272_0(.douta(w_n20272_0[0]),.doutb(w_n20272_0[1]),.din(n20272));
	jspl jspl_w_n20273_0(.douta(w_n20273_0[0]),.doutb(w_n20273_0[1]),.din(n20273));
	jspl3 jspl3_w_n20274_0(.douta(w_n20274_0[0]),.doutb(w_n20274_0[1]),.doutc(w_n20274_0[2]),.din(n20274));
	jspl jspl_w_n20275_0(.douta(w_n20275_0[0]),.doutb(w_n20275_0[1]),.din(n20275));
	jspl jspl_w_n20280_0(.douta(w_n20280_0[0]),.doutb(w_n20280_0[1]),.din(n20280));
	jspl jspl_w_n20281_0(.douta(w_n20281_0[0]),.doutb(w_n20281_0[1]),.din(n20281));
	jspl jspl_w_n20283_0(.douta(w_n20283_0[0]),.doutb(w_n20283_0[1]),.din(n20283));
	jspl jspl_w_n20285_0(.douta(w_n20285_0[0]),.doutb(w_n20285_0[1]),.din(n20285));
	jspl jspl_w_n20288_0(.douta(w_n20288_0[0]),.doutb(w_n20288_0[1]),.din(n20288));
	jspl jspl_w_n20294_0(.douta(w_n20294_0[0]),.doutb(w_n20294_0[1]),.din(n20294));
	jspl3 jspl3_w_n20296_0(.douta(w_n20296_0[0]),.doutb(w_n20296_0[1]),.doutc(w_n20296_0[2]),.din(n20296));
	jspl jspl_w_n20297_0(.douta(w_n20297_0[0]),.doutb(w_n20297_0[1]),.din(n20297));
	jspl jspl_w_n20301_0(.douta(w_n20301_0[0]),.doutb(w_n20301_0[1]),.din(n20301));
	jspl jspl_w_n20302_0(.douta(w_n20302_0[0]),.doutb(w_n20302_0[1]),.din(n20302));
	jspl jspl_w_n20304_0(.douta(w_n20304_0[0]),.doutb(w_n20304_0[1]),.din(n20304));
	jspl jspl_w_n20308_0(.douta(w_n20308_0[0]),.doutb(w_n20308_0[1]),.din(n20308));
	jspl jspl_w_n20311_0(.douta(w_n20311_0[0]),.doutb(w_n20311_0[1]),.din(n20311));
	jspl jspl_w_n20312_0(.douta(w_n20312_0[0]),.doutb(w_n20312_0[1]),.din(n20312));
	jspl3 jspl3_w_n20313_0(.douta(w_n20313_0[0]),.doutb(w_n20313_0[1]),.doutc(w_n20313_0[2]),.din(n20313));
	jspl jspl_w_n20314_0(.douta(w_n20314_0[0]),.doutb(w_n20314_0[1]),.din(n20314));
	jspl jspl_w_n20318_0(.douta(w_n20318_0[0]),.doutb(w_n20318_0[1]),.din(n20318));
	jspl jspl_w_n20319_0(.douta(w_n20319_0[0]),.doutb(w_n20319_0[1]),.din(n20319));
	jspl jspl_w_n20321_0(.douta(w_n20321_0[0]),.doutb(w_n20321_0[1]),.din(n20321));
	jspl jspl_w_n20323_0(.douta(w_n20323_0[0]),.doutb(w_n20323_0[1]),.din(n20323));
	jspl jspl_w_n20326_0(.douta(w_n20326_0[0]),.doutb(w_n20326_0[1]),.din(n20326));
	jspl jspl_w_n20332_0(.douta(w_n20332_0[0]),.doutb(w_n20332_0[1]),.din(n20332));
	jspl jspl_w_n20334_0(.douta(w_n20334_0[0]),.doutb(w_n20334_0[1]),.din(n20334));
	jspl3 jspl3_w_n20335_0(.douta(w_n20335_0[0]),.doutb(w_n20335_0[1]),.doutc(w_n20335_0[2]),.din(n20335));
	jspl jspl_w_n20338_0(.douta(w_n20338_0[0]),.doutb(w_n20338_0[1]),.din(n20338));
	jspl jspl_w_n20340_0(.douta(w_n20340_0[0]),.doutb(w_n20340_0[1]),.din(n20340));
	jspl3 jspl3_w_n20341_0(.douta(w_n20341_0[0]),.doutb(w_n20341_0[1]),.doutc(w_n20341_0[2]),.din(n20341));
	jspl jspl_w_n20343_0(.douta(w_n20343_0[0]),.doutb(w_n20343_0[1]),.din(n20343));
	jspl jspl_w_n20347_0(.douta(w_n20347_0[0]),.doutb(w_n20347_0[1]),.din(n20347));
	jspl jspl_w_n20350_0(.douta(w_n20350_0[0]),.doutb(w_n20350_0[1]),.din(n20350));
	jspl jspl_w_n20351_0(.douta(w_n20351_0[0]),.doutb(w_n20351_0[1]),.din(n20351));
	jspl3 jspl3_w_n20352_0(.douta(w_n20352_0[0]),.doutb(w_n20352_0[1]),.doutc(w_n20352_0[2]),.din(n20352));
	jspl jspl_w_n20353_0(.douta(w_n20353_0[0]),.doutb(w_n20353_0[1]),.din(n20353));
	jspl jspl_w_n20357_0(.douta(w_n20357_0[0]),.doutb(w_n20357_0[1]),.din(n20357));
	jspl jspl_w_n20363_0(.douta(w_n20363_0[0]),.doutb(w_n20363_0[1]),.din(n20363));
	jspl jspl_w_n20364_0(.douta(w_n20364_0[0]),.doutb(w_n20364_0[1]),.din(n20364));
	jspl jspl_w_n20366_0(.douta(w_n20366_0[0]),.doutb(w_n20366_0[1]),.din(n20366));
	jspl jspl_w_n20368_0(.douta(w_n20368_0[0]),.doutb(w_n20368_0[1]),.din(n20368));
	jspl jspl_w_n20371_0(.douta(w_n20371_0[0]),.doutb(w_n20371_0[1]),.din(n20371));
	jspl jspl_w_n20377_0(.douta(w_n20377_0[0]),.doutb(w_n20377_0[1]),.din(n20377));
	jspl jspl_w_n20379_0(.douta(w_n20379_0[0]),.doutb(w_n20379_0[1]),.din(n20379));
	jspl3 jspl3_w_n20380_0(.douta(w_n20380_0[0]),.doutb(w_n20380_0[1]),.doutc(w_n20380_0[2]),.din(n20380));
	jspl jspl_w_n20383_0(.douta(w_n20383_0[0]),.doutb(w_n20383_0[1]),.din(n20383));
	jspl jspl_w_n20385_0(.douta(w_n20385_0[0]),.doutb(w_n20385_0[1]),.din(n20385));
	jspl3 jspl3_w_n20386_0(.douta(w_n20386_0[0]),.doutb(w_n20386_0[1]),.doutc(w_n20386_0[2]),.din(n20386));
	jspl jspl_w_n20388_0(.douta(w_n20388_0[0]),.doutb(w_n20388_0[1]),.din(n20388));
	jspl jspl_w_n20392_0(.douta(w_n20392_0[0]),.doutb(w_n20392_0[1]),.din(n20392));
	jspl jspl_w_n20395_0(.douta(w_n20395_0[0]),.doutb(w_n20395_0[1]),.din(n20395));
	jspl jspl_w_n20396_0(.douta(w_n20396_0[0]),.doutb(w_n20396_0[1]),.din(n20396));
	jspl3 jspl3_w_n20397_0(.douta(w_n20397_0[0]),.doutb(w_n20397_0[1]),.doutc(w_n20397_0[2]),.din(n20397));
	jspl jspl_w_n20398_0(.douta(w_n20398_0[0]),.doutb(w_n20398_0[1]),.din(n20398));
	jspl jspl_w_n20402_0(.douta(w_n20402_0[0]),.doutb(w_n20402_0[1]),.din(n20402));
	jspl jspl_w_n20408_0(.douta(w_n20408_0[0]),.doutb(w_n20408_0[1]),.din(n20408));
	jspl jspl_w_n20409_0(.douta(w_n20409_0[0]),.doutb(w_n20409_0[1]),.din(n20409));
	jspl jspl_w_n20411_0(.douta(w_n20411_0[0]),.doutb(w_n20411_0[1]),.din(n20411));
	jspl jspl_w_n20413_0(.douta(w_n20413_0[0]),.doutb(w_n20413_0[1]),.din(n20413));
	jspl jspl_w_n20416_0(.douta(w_n20416_0[0]),.doutb(w_n20416_0[1]),.din(n20416));
	jspl jspl_w_n20422_0(.douta(w_n20422_0[0]),.doutb(w_n20422_0[1]),.din(n20422));
	jspl jspl_w_n20424_0(.douta(w_n20424_0[0]),.doutb(w_n20424_0[1]),.din(n20424));
	jspl3 jspl3_w_n20425_0(.douta(w_n20425_0[0]),.doutb(w_n20425_0[1]),.doutc(w_n20425_0[2]),.din(n20425));
	jspl jspl_w_n20428_0(.douta(w_n20428_0[0]),.doutb(w_n20428_0[1]),.din(n20428));
	jspl jspl_w_n20430_0(.douta(w_n20430_0[0]),.doutb(w_n20430_0[1]),.din(n20430));
	jspl3 jspl3_w_n20431_0(.douta(w_n20431_0[0]),.doutb(w_n20431_0[1]),.doutc(w_n20431_0[2]),.din(n20431));
	jspl jspl_w_n20433_0(.douta(w_n20433_0[0]),.doutb(w_n20433_0[1]),.din(n20433));
	jspl jspl_w_n20437_0(.douta(w_n20437_0[0]),.doutb(w_n20437_0[1]),.din(n20437));
	jspl jspl_w_n20440_0(.douta(w_n20440_0[0]),.doutb(w_n20440_0[1]),.din(n20440));
	jspl jspl_w_n20441_0(.douta(w_n20441_0[0]),.doutb(w_n20441_0[1]),.din(n20441));
	jspl3 jspl3_w_n20442_0(.douta(w_n20442_0[0]),.doutb(w_n20442_0[1]),.doutc(w_n20442_0[2]),.din(n20442));
	jspl jspl_w_n20443_0(.douta(w_n20443_0[0]),.doutb(w_n20443_0[1]),.din(n20443));
	jspl jspl_w_n20447_0(.douta(w_n20447_0[0]),.doutb(w_n20447_0[1]),.din(n20447));
	jspl jspl_w_n20453_0(.douta(w_n20453_0[0]),.doutb(w_n20453_0[1]),.din(n20453));
	jspl jspl_w_n20454_0(.douta(w_n20454_0[0]),.doutb(w_n20454_0[1]),.din(n20454));
	jspl jspl_w_n20456_0(.douta(w_n20456_0[0]),.doutb(w_n20456_0[1]),.din(n20456));
	jspl jspl_w_n20458_0(.douta(w_n20458_0[0]),.doutb(w_n20458_0[1]),.din(n20458));
	jspl jspl_w_n20461_0(.douta(w_n20461_0[0]),.doutb(w_n20461_0[1]),.din(n20461));
	jspl jspl_w_n20467_0(.douta(w_n20467_0[0]),.doutb(w_n20467_0[1]),.din(n20467));
	jspl jspl_w_n20469_0(.douta(w_n20469_0[0]),.doutb(w_n20469_0[1]),.din(n20469));
	jspl3 jspl3_w_n20470_0(.douta(w_n20470_0[0]),.doutb(w_n20470_0[1]),.doutc(w_n20470_0[2]),.din(n20470));
	jspl jspl_w_n20473_0(.douta(w_n20473_0[0]),.doutb(w_n20473_0[1]),.din(n20473));
	jspl jspl_w_n20475_0(.douta(w_n20475_0[0]),.doutb(w_n20475_0[1]),.din(n20475));
	jspl3 jspl3_w_n20476_0(.douta(w_n20476_0[0]),.doutb(w_n20476_0[1]),.doutc(w_n20476_0[2]),.din(n20476));
	jspl jspl_w_n20478_0(.douta(w_n20478_0[0]),.doutb(w_n20478_0[1]),.din(n20478));
	jspl jspl_w_n20482_0(.douta(w_n20482_0[0]),.doutb(w_n20482_0[1]),.din(n20482));
	jspl jspl_w_n20485_0(.douta(w_n20485_0[0]),.doutb(w_n20485_0[1]),.din(n20485));
	jspl jspl_w_n20486_0(.douta(w_n20486_0[0]),.doutb(w_n20486_0[1]),.din(n20486));
	jspl3 jspl3_w_n20487_0(.douta(w_n20487_0[0]),.doutb(w_n20487_0[1]),.doutc(w_n20487_0[2]),.din(n20487));
	jspl jspl_w_n20488_0(.douta(w_n20488_0[0]),.doutb(w_n20488_0[1]),.din(n20488));
	jspl jspl_w_n20492_0(.douta(w_n20492_0[0]),.doutb(w_n20492_0[1]),.din(n20492));
	jspl jspl_w_n20498_0(.douta(w_n20498_0[0]),.doutb(w_n20498_0[1]),.din(n20498));
	jspl jspl_w_n20499_0(.douta(w_n20499_0[0]),.doutb(w_n20499_0[1]),.din(n20499));
	jspl jspl_w_n20501_0(.douta(w_n20501_0[0]),.doutb(w_n20501_0[1]),.din(n20501));
	jspl jspl_w_n20503_0(.douta(w_n20503_0[0]),.doutb(w_n20503_0[1]),.din(n20503));
	jspl jspl_w_n20506_0(.douta(w_n20506_0[0]),.doutb(w_n20506_0[1]),.din(n20506));
	jspl jspl_w_n20512_0(.douta(w_n20512_0[0]),.doutb(w_n20512_0[1]),.din(n20512));
	jspl jspl_w_n20514_0(.douta(w_n20514_0[0]),.doutb(w_n20514_0[1]),.din(n20514));
	jspl3 jspl3_w_n20515_0(.douta(w_n20515_0[0]),.doutb(w_n20515_0[1]),.doutc(w_n20515_0[2]),.din(n20515));
	jspl jspl_w_n20518_0(.douta(w_n20518_0[0]),.doutb(w_n20518_0[1]),.din(n20518));
	jspl jspl_w_n20520_0(.douta(w_n20520_0[0]),.doutb(w_n20520_0[1]),.din(n20520));
	jspl3 jspl3_w_n20521_0(.douta(w_n20521_0[0]),.doutb(w_n20521_0[1]),.doutc(w_n20521_0[2]),.din(n20521));
	jspl jspl_w_n20523_0(.douta(w_n20523_0[0]),.doutb(w_n20523_0[1]),.din(n20523));
	jspl jspl_w_n20527_0(.douta(w_n20527_0[0]),.doutb(w_n20527_0[1]),.din(n20527));
	jspl jspl_w_n20530_0(.douta(w_n20530_0[0]),.doutb(w_n20530_0[1]),.din(n20530));
	jspl jspl_w_n20531_0(.douta(w_n20531_0[0]),.doutb(w_n20531_0[1]),.din(n20531));
	jspl3 jspl3_w_n20532_0(.douta(w_n20532_0[0]),.doutb(w_n20532_0[1]),.doutc(w_n20532_0[2]),.din(n20532));
	jspl jspl_w_n20533_0(.douta(w_n20533_0[0]),.doutb(w_n20533_0[1]),.din(n20533));
	jspl jspl_w_n20537_0(.douta(w_n20537_0[0]),.doutb(w_n20537_0[1]),.din(n20537));
	jspl jspl_w_n20543_0(.douta(w_n20543_0[0]),.doutb(w_n20543_0[1]),.din(n20543));
	jspl jspl_w_n20544_0(.douta(w_n20544_0[0]),.doutb(w_n20544_0[1]),.din(n20544));
	jspl jspl_w_n20546_0(.douta(w_n20546_0[0]),.doutb(w_n20546_0[1]),.din(n20546));
	jspl jspl_w_n20548_0(.douta(w_n20548_0[0]),.doutb(w_n20548_0[1]),.din(n20548));
	jspl jspl_w_n20551_0(.douta(w_n20551_0[0]),.doutb(w_n20551_0[1]),.din(n20551));
	jspl jspl_w_n20557_0(.douta(w_n20557_0[0]),.doutb(w_n20557_0[1]),.din(n20557));
	jspl jspl_w_n20559_0(.douta(w_n20559_0[0]),.doutb(w_n20559_0[1]),.din(n20559));
	jspl3 jspl3_w_n20560_0(.douta(w_n20560_0[0]),.doutb(w_n20560_0[1]),.doutc(w_n20560_0[2]),.din(n20560));
	jspl jspl_w_n20563_0(.douta(w_n20563_0[0]),.doutb(w_n20563_0[1]),.din(n20563));
	jspl jspl_w_n20565_0(.douta(w_n20565_0[0]),.doutb(w_n20565_0[1]),.din(n20565));
	jspl3 jspl3_w_n20566_0(.douta(w_n20566_0[0]),.doutb(w_n20566_0[1]),.doutc(w_n20566_0[2]),.din(n20566));
	jspl jspl_w_n20568_0(.douta(w_n20568_0[0]),.doutb(w_n20568_0[1]),.din(n20568));
	jspl jspl_w_n20572_0(.douta(w_n20572_0[0]),.doutb(w_n20572_0[1]),.din(n20572));
	jspl jspl_w_n20575_0(.douta(w_n20575_0[0]),.doutb(w_n20575_0[1]),.din(n20575));
	jspl jspl_w_n20576_0(.douta(w_n20576_0[0]),.doutb(w_n20576_0[1]),.din(n20576));
	jspl3 jspl3_w_n20577_0(.douta(w_n20577_0[0]),.doutb(w_n20577_0[1]),.doutc(w_n20577_0[2]),.din(n20577));
	jspl jspl_w_n20578_0(.douta(w_n20578_0[0]),.doutb(w_n20578_0[1]),.din(n20578));
	jspl jspl_w_n20582_0(.douta(w_n20582_0[0]),.doutb(w_n20582_0[1]),.din(n20582));
	jspl jspl_w_n20588_0(.douta(w_n20588_0[0]),.doutb(w_n20588_0[1]),.din(n20588));
	jspl jspl_w_n20589_0(.douta(w_n20589_0[0]),.doutb(w_n20589_0[1]),.din(n20589));
	jspl jspl_w_n20591_0(.douta(w_n20591_0[0]),.doutb(w_n20591_0[1]),.din(n20591));
	jspl jspl_w_n20593_0(.douta(w_n20593_0[0]),.doutb(w_n20593_0[1]),.din(n20593));
	jspl jspl_w_n20596_0(.douta(w_n20596_0[0]),.doutb(w_n20596_0[1]),.din(n20596));
	jspl jspl_w_n20602_0(.douta(w_n20602_0[0]),.doutb(w_n20602_0[1]),.din(n20602));
	jspl jspl_w_n20604_0(.douta(w_n20604_0[0]),.doutb(w_n20604_0[1]),.din(n20604));
	jspl3 jspl3_w_n20605_0(.douta(w_n20605_0[0]),.doutb(w_n20605_0[1]),.doutc(w_n20605_0[2]),.din(n20605));
	jspl jspl_w_n20608_0(.douta(w_n20608_0[0]),.doutb(w_n20608_0[1]),.din(n20608));
	jspl jspl_w_n20610_0(.douta(w_n20610_0[0]),.doutb(w_n20610_0[1]),.din(n20610));
	jspl3 jspl3_w_n20611_0(.douta(w_n20611_0[0]),.doutb(w_n20611_0[1]),.doutc(w_n20611_0[2]),.din(n20611));
	jspl jspl_w_n20613_0(.douta(w_n20613_0[0]),.doutb(w_n20613_0[1]),.din(n20613));
	jspl jspl_w_n20617_0(.douta(w_n20617_0[0]),.doutb(w_n20617_0[1]),.din(n20617));
	jspl jspl_w_n20620_0(.douta(w_n20620_0[0]),.doutb(w_n20620_0[1]),.din(n20620));
	jspl jspl_w_n20621_0(.douta(w_n20621_0[0]),.doutb(w_n20621_0[1]),.din(n20621));
	jspl3 jspl3_w_n20622_0(.douta(w_n20622_0[0]),.doutb(w_n20622_0[1]),.doutc(w_n20622_0[2]),.din(n20622));
	jspl jspl_w_n20623_0(.douta(w_n20623_0[0]),.doutb(w_n20623_0[1]),.din(n20623));
	jspl jspl_w_n20627_0(.douta(w_n20627_0[0]),.doutb(w_n20627_0[1]),.din(n20627));
	jspl jspl_w_n20633_0(.douta(w_n20633_0[0]),.doutb(w_n20633_0[1]),.din(n20633));
	jspl jspl_w_n20634_0(.douta(w_n20634_0[0]),.doutb(w_n20634_0[1]),.din(n20634));
	jspl jspl_w_n20636_0(.douta(w_n20636_0[0]),.doutb(w_n20636_0[1]),.din(n20636));
	jspl jspl_w_n20638_0(.douta(w_n20638_0[0]),.doutb(w_n20638_0[1]),.din(n20638));
	jspl jspl_w_n20641_0(.douta(w_n20641_0[0]),.doutb(w_n20641_0[1]),.din(n20641));
	jspl jspl_w_n20647_0(.douta(w_n20647_0[0]),.doutb(w_n20647_0[1]),.din(n20647));
	jspl jspl_w_n20649_0(.douta(w_n20649_0[0]),.doutb(w_n20649_0[1]),.din(n20649));
	jspl3 jspl3_w_n20650_0(.douta(w_n20650_0[0]),.doutb(w_n20650_0[1]),.doutc(w_n20650_0[2]),.din(n20650));
	jspl jspl_w_n20653_0(.douta(w_n20653_0[0]),.doutb(w_n20653_0[1]),.din(n20653));
	jspl jspl_w_n20655_0(.douta(w_n20655_0[0]),.doutb(w_n20655_0[1]),.din(n20655));
	jspl3 jspl3_w_n20656_0(.douta(w_n20656_0[0]),.doutb(w_n20656_0[1]),.doutc(w_n20656_0[2]),.din(n20656));
	jspl jspl_w_n20658_0(.douta(w_n20658_0[0]),.doutb(w_n20658_0[1]),.din(n20658));
	jspl jspl_w_n20662_0(.douta(w_n20662_0[0]),.doutb(w_n20662_0[1]),.din(n20662));
	jspl jspl_w_n20665_0(.douta(w_n20665_0[0]),.doutb(w_n20665_0[1]),.din(n20665));
	jspl jspl_w_n20666_0(.douta(w_n20666_0[0]),.doutb(w_n20666_0[1]),.din(n20666));
	jspl3 jspl3_w_n20667_0(.douta(w_n20667_0[0]),.doutb(w_n20667_0[1]),.doutc(w_n20667_0[2]),.din(n20667));
	jspl jspl_w_n20668_0(.douta(w_n20668_0[0]),.doutb(w_n20668_0[1]),.din(n20668));
	jspl jspl_w_n20672_0(.douta(w_n20672_0[0]),.doutb(w_n20672_0[1]),.din(n20672));
	jspl jspl_w_n20678_0(.douta(w_n20678_0[0]),.doutb(w_n20678_0[1]),.din(n20678));
	jspl jspl_w_n20679_0(.douta(w_n20679_0[0]),.doutb(w_n20679_0[1]),.din(n20679));
	jspl jspl_w_n20681_0(.douta(w_n20681_0[0]),.doutb(w_n20681_0[1]),.din(n20681));
	jspl jspl_w_n20683_0(.douta(w_n20683_0[0]),.doutb(w_n20683_0[1]),.din(n20683));
	jspl jspl_w_n20686_0(.douta(w_n20686_0[0]),.doutb(w_n20686_0[1]),.din(n20686));
	jspl jspl_w_n20692_0(.douta(w_n20692_0[0]),.doutb(w_n20692_0[1]),.din(n20692));
	jspl jspl_w_n20694_0(.douta(w_n20694_0[0]),.doutb(w_n20694_0[1]),.din(n20694));
	jspl3 jspl3_w_n20695_0(.douta(w_n20695_0[0]),.doutb(w_n20695_0[1]),.doutc(w_n20695_0[2]),.din(n20695));
	jspl jspl_w_n20698_0(.douta(w_n20698_0[0]),.doutb(w_n20698_0[1]),.din(n20698));
	jspl jspl_w_n20700_0(.douta(w_n20700_0[0]),.doutb(w_n20700_0[1]),.din(n20700));
	jspl3 jspl3_w_n20701_0(.douta(w_n20701_0[0]),.doutb(w_n20701_0[1]),.doutc(w_n20701_0[2]),.din(n20701));
	jspl jspl_w_n20703_0(.douta(w_n20703_0[0]),.doutb(w_n20703_0[1]),.din(n20703));
	jspl jspl_w_n20707_0(.douta(w_n20707_0[0]),.doutb(w_n20707_0[1]),.din(n20707));
	jspl jspl_w_n20710_0(.douta(w_n20710_0[0]),.doutb(w_n20710_0[1]),.din(n20710));
	jspl jspl_w_n20711_0(.douta(w_n20711_0[0]),.doutb(w_n20711_0[1]),.din(n20711));
	jspl3 jspl3_w_n20712_0(.douta(w_n20712_0[0]),.doutb(w_n20712_0[1]),.doutc(w_n20712_0[2]),.din(n20712));
	jspl jspl_w_n20713_0(.douta(w_n20713_0[0]),.doutb(w_n20713_0[1]),.din(n20713));
	jspl jspl_w_n20717_0(.douta(w_n20717_0[0]),.doutb(w_n20717_0[1]),.din(n20717));
	jspl jspl_w_n20723_0(.douta(w_n20723_0[0]),.doutb(w_n20723_0[1]),.din(n20723));
	jspl jspl_w_n20724_0(.douta(w_n20724_0[0]),.doutb(w_n20724_0[1]),.din(n20724));
	jspl jspl_w_n20726_0(.douta(w_n20726_0[0]),.doutb(w_n20726_0[1]),.din(n20726));
	jspl jspl_w_n20728_0(.douta(w_n20728_0[0]),.doutb(w_n20728_0[1]),.din(n20728));
	jspl jspl_w_n20731_0(.douta(w_n20731_0[0]),.doutb(w_n20731_0[1]),.din(n20731));
	jspl jspl_w_n20737_0(.douta(w_n20737_0[0]),.doutb(w_n20737_0[1]),.din(n20737));
	jspl jspl_w_n20739_0(.douta(w_n20739_0[0]),.doutb(w_n20739_0[1]),.din(n20739));
	jspl3 jspl3_w_n20740_0(.douta(w_n20740_0[0]),.doutb(w_n20740_0[1]),.doutc(w_n20740_0[2]),.din(n20740));
	jspl jspl_w_n20743_0(.douta(w_n20743_0[0]),.doutb(w_n20743_0[1]),.din(n20743));
	jspl jspl_w_n20745_0(.douta(w_n20745_0[0]),.doutb(w_n20745_0[1]),.din(n20745));
	jspl3 jspl3_w_n20746_0(.douta(w_n20746_0[0]),.doutb(w_n20746_0[1]),.doutc(w_n20746_0[2]),.din(n20746));
	jspl jspl_w_n20748_0(.douta(w_n20748_0[0]),.doutb(w_n20748_0[1]),.din(n20748));
	jspl jspl_w_n20752_0(.douta(w_n20752_0[0]),.doutb(w_n20752_0[1]),.din(n20752));
	jspl jspl_w_n20755_0(.douta(w_n20755_0[0]),.doutb(w_n20755_0[1]),.din(n20755));
	jspl jspl_w_n20756_0(.douta(w_n20756_0[0]),.doutb(w_n20756_0[1]),.din(n20756));
	jspl3 jspl3_w_n20757_0(.douta(w_n20757_0[0]),.doutb(w_n20757_0[1]),.doutc(w_n20757_0[2]),.din(n20757));
	jspl jspl_w_n20758_0(.douta(w_n20758_0[0]),.doutb(w_n20758_0[1]),.din(n20758));
	jspl jspl_w_n20762_0(.douta(w_n20762_0[0]),.doutb(w_n20762_0[1]),.din(n20762));
	jspl jspl_w_n20768_0(.douta(w_n20768_0[0]),.doutb(w_n20768_0[1]),.din(n20768));
	jspl jspl_w_n20769_0(.douta(w_n20769_0[0]),.doutb(w_n20769_0[1]),.din(n20769));
	jspl jspl_w_n20771_0(.douta(w_n20771_0[0]),.doutb(w_n20771_0[1]),.din(n20771));
	jspl jspl_w_n20773_0(.douta(w_n20773_0[0]),.doutb(w_n20773_0[1]),.din(n20773));
	jspl jspl_w_n20776_0(.douta(w_n20776_0[0]),.doutb(w_n20776_0[1]),.din(n20776));
	jspl jspl_w_n20782_0(.douta(w_n20782_0[0]),.doutb(w_n20782_0[1]),.din(n20782));
	jspl jspl_w_n20784_0(.douta(w_n20784_0[0]),.doutb(w_n20784_0[1]),.din(n20784));
	jspl3 jspl3_w_n20785_0(.douta(w_n20785_0[0]),.doutb(w_n20785_0[1]),.doutc(w_n20785_0[2]),.din(n20785));
	jspl jspl_w_n20788_0(.douta(w_n20788_0[0]),.doutb(w_n20788_0[1]),.din(n20788));
	jspl jspl_w_n20790_0(.douta(w_n20790_0[0]),.doutb(w_n20790_0[1]),.din(n20790));
	jspl3 jspl3_w_n20791_0(.douta(w_n20791_0[0]),.doutb(w_n20791_0[1]),.doutc(w_n20791_0[2]),.din(n20791));
	jspl jspl_w_n20793_0(.douta(w_n20793_0[0]),.doutb(w_n20793_0[1]),.din(n20793));
	jspl jspl_w_n20797_0(.douta(w_n20797_0[0]),.doutb(w_n20797_0[1]),.din(n20797));
	jspl jspl_w_n20800_0(.douta(w_n20800_0[0]),.doutb(w_n20800_0[1]),.din(n20800));
	jspl jspl_w_n20801_0(.douta(w_n20801_0[0]),.doutb(w_n20801_0[1]),.din(n20801));
	jspl3 jspl3_w_n20802_0(.douta(w_n20802_0[0]),.doutb(w_n20802_0[1]),.doutc(w_n20802_0[2]),.din(n20802));
	jspl jspl_w_n20803_0(.douta(w_n20803_0[0]),.doutb(w_n20803_0[1]),.din(n20803));
	jspl jspl_w_n20807_0(.douta(w_n20807_0[0]),.doutb(w_n20807_0[1]),.din(n20807));
	jspl jspl_w_n20813_0(.douta(w_n20813_0[0]),.doutb(w_n20813_0[1]),.din(n20813));
	jspl jspl_w_n20814_0(.douta(w_n20814_0[0]),.doutb(w_n20814_0[1]),.din(n20814));
	jspl jspl_w_n20816_0(.douta(w_n20816_0[0]),.doutb(w_n20816_0[1]),.din(n20816));
	jspl jspl_w_n20818_0(.douta(w_n20818_0[0]),.doutb(w_n20818_0[1]),.din(n20818));
	jspl jspl_w_n20821_0(.douta(w_n20821_0[0]),.doutb(w_n20821_0[1]),.din(n20821));
	jspl jspl_w_n20827_0(.douta(w_n20827_0[0]),.doutb(w_n20827_0[1]),.din(n20827));
	jspl jspl_w_n20829_0(.douta(w_n20829_0[0]),.doutb(w_n20829_0[1]),.din(n20829));
	jspl3 jspl3_w_n20830_0(.douta(w_n20830_0[0]),.doutb(w_n20830_0[1]),.doutc(w_n20830_0[2]),.din(n20830));
	jspl jspl_w_n20833_0(.douta(w_n20833_0[0]),.doutb(w_n20833_0[1]),.din(n20833));
	jspl jspl_w_n20835_0(.douta(w_n20835_0[0]),.doutb(w_n20835_0[1]),.din(n20835));
	jspl3 jspl3_w_n20836_0(.douta(w_n20836_0[0]),.doutb(w_n20836_0[1]),.doutc(w_n20836_0[2]),.din(n20836));
	jspl jspl_w_n20838_0(.douta(w_n20838_0[0]),.doutb(w_n20838_0[1]),.din(n20838));
	jspl jspl_w_n20842_0(.douta(w_n20842_0[0]),.doutb(w_n20842_0[1]),.din(n20842));
	jspl jspl_w_n20845_0(.douta(w_n20845_0[0]),.doutb(w_n20845_0[1]),.din(n20845));
	jspl jspl_w_n20846_0(.douta(w_n20846_0[0]),.doutb(w_n20846_0[1]),.din(n20846));
	jspl3 jspl3_w_n20847_0(.douta(w_n20847_0[0]),.doutb(w_n20847_0[1]),.doutc(w_n20847_0[2]),.din(n20847));
	jspl jspl_w_n20848_0(.douta(w_n20848_0[0]),.doutb(w_n20848_0[1]),.din(n20848));
	jspl jspl_w_n20852_0(.douta(w_n20852_0[0]),.doutb(w_n20852_0[1]),.din(n20852));
	jspl jspl_w_n20858_0(.douta(w_n20858_0[0]),.doutb(w_n20858_0[1]),.din(n20858));
	jspl jspl_w_n20859_0(.douta(w_n20859_0[0]),.doutb(w_n20859_0[1]),.din(n20859));
	jspl jspl_w_n20861_0(.douta(w_n20861_0[0]),.doutb(w_n20861_0[1]),.din(n20861));
	jspl jspl_w_n20865_0(.douta(w_n20865_0[0]),.doutb(w_n20865_0[1]),.din(n20865));
	jspl jspl_w_n20868_0(.douta(w_n20868_0[0]),.doutb(w_n20868_0[1]),.din(n20868));
	jspl jspl_w_n20869_0(.douta(w_n20869_0[0]),.doutb(w_n20869_0[1]),.din(n20869));
	jspl3 jspl3_w_n20870_0(.douta(w_n20870_0[0]),.doutb(w_n20870_0[1]),.doutc(w_n20870_0[2]),.din(n20870));
	jspl jspl_w_n20871_0(.douta(w_n20871_0[0]),.doutb(w_n20871_0[1]),.din(n20871));
	jspl jspl_w_n20873_0(.douta(w_n20873_0[0]),.doutb(w_n20873_0[1]),.din(n20873));
	jspl jspl_w_n20875_0(.douta(w_n20875_0[0]),.doutb(w_n20875_0[1]),.din(n20875));
	jspl jspl_w_n20877_0(.douta(w_n20877_0[0]),.doutb(w_n20877_0[1]),.din(n20877));
	jspl jspl_w_n20880_0(.douta(w_n20880_0[0]),.doutb(w_n20880_0[1]),.din(n20880));
	jspl jspl_w_n20886_0(.douta(w_n20886_0[0]),.doutb(w_n20886_0[1]),.din(n20886));
	jspl3 jspl3_w_n20888_0(.douta(w_n20888_0[0]),.doutb(w_n20888_0[1]),.doutc(w_n20888_0[2]),.din(n20888));
	jspl3 jspl3_w_n20888_1(.douta(w_n20888_1[0]),.doutb(w_n20888_1[1]),.doutc(w_n20888_1[2]),.din(w_n20888_0[0]));
	jspl3 jspl3_w_n20891_0(.douta(w_n20891_0[0]),.doutb(w_n20891_0[1]),.doutc(w_n20891_0[2]),.din(n20891));
	jspl3 jspl3_w_n20892_0(.douta(w_n20892_0[0]),.doutb(w_n20892_0[1]),.doutc(w_n20892_0[2]),.din(n20892));
	jspl jspl_w_n20893_0(.douta(w_n20893_0[0]),.doutb(w_n20893_0[1]),.din(n20893));
	jspl jspl_w_n20894_0(.douta(w_n20894_0[0]),.doutb(w_n20894_0[1]),.din(n20894));
	jspl jspl_w_n20901_0(.douta(w_n20901_0[0]),.doutb(w_n20901_0[1]),.din(n20901));
	jspl jspl_w_n20902_0(.douta(w_n20902_0[0]),.doutb(w_n20902_0[1]),.din(n20902));
	jspl3 jspl3_w_n20910_0(.douta(w_n20910_0[0]),.doutb(w_n20910_0[1]),.doutc(w_n20910_0[2]),.din(n20910));
	jspl3 jspl3_w_n20910_1(.douta(w_n20910_1[0]),.doutb(w_n20910_1[1]),.doutc(w_n20910_1[2]),.din(w_n20910_0[0]));
	jspl3 jspl3_w_n20910_2(.douta(w_n20910_2[0]),.doutb(w_n20910_2[1]),.doutc(w_n20910_2[2]),.din(w_n20910_0[1]));
	jspl3 jspl3_w_n20910_3(.douta(w_n20910_3[0]),.doutb(w_n20910_3[1]),.doutc(w_n20910_3[2]),.din(w_n20910_0[2]));
	jspl3 jspl3_w_n20910_4(.douta(w_n20910_4[0]),.doutb(w_n20910_4[1]),.doutc(w_n20910_4[2]),.din(w_n20910_1[0]));
	jspl3 jspl3_w_n20910_5(.douta(w_n20910_5[0]),.doutb(w_n20910_5[1]),.doutc(w_n20910_5[2]),.din(w_n20910_1[1]));
	jspl3 jspl3_w_n20910_6(.douta(w_n20910_6[0]),.doutb(w_n20910_6[1]),.doutc(w_n20910_6[2]),.din(w_n20910_1[2]));
	jspl3 jspl3_w_n20910_7(.douta(w_n20910_7[0]),.doutb(w_n20910_7[1]),.doutc(w_n20910_7[2]),.din(w_n20910_2[0]));
	jspl3 jspl3_w_n20910_8(.douta(w_n20910_8[0]),.doutb(w_n20910_8[1]),.doutc(w_n20910_8[2]),.din(w_n20910_2[1]));
	jspl3 jspl3_w_n20910_9(.douta(w_n20910_9[0]),.doutb(w_n20910_9[1]),.doutc(w_n20910_9[2]),.din(w_n20910_2[2]));
	jspl3 jspl3_w_n20910_10(.douta(w_n20910_10[0]),.doutb(w_n20910_10[1]),.doutc(w_n20910_10[2]),.din(w_n20910_3[0]));
	jspl3 jspl3_w_n20910_11(.douta(w_n20910_11[0]),.doutb(w_n20910_11[1]),.doutc(w_n20910_11[2]),.din(w_n20910_3[1]));
	jspl3 jspl3_w_n20910_12(.douta(w_n20910_12[0]),.doutb(w_n20910_12[1]),.doutc(w_n20910_12[2]),.din(w_n20910_3[2]));
	jspl3 jspl3_w_n20910_13(.douta(w_n20910_13[0]),.doutb(w_n20910_13[1]),.doutc(w_n20910_13[2]),.din(w_n20910_4[0]));
	jspl3 jspl3_w_n20910_14(.douta(w_n20910_14[0]),.doutb(w_n20910_14[1]),.doutc(w_n20910_14[2]),.din(w_n20910_4[1]));
	jspl3 jspl3_w_n20910_15(.douta(w_n20910_15[0]),.doutb(w_n20910_15[1]),.doutc(w_n20910_15[2]),.din(w_n20910_4[2]));
	jspl3 jspl3_w_n20910_16(.douta(w_n20910_16[0]),.doutb(w_n20910_16[1]),.doutc(w_n20910_16[2]),.din(w_n20910_5[0]));
	jspl3 jspl3_w_n20910_17(.douta(w_n20910_17[0]),.doutb(w_n20910_17[1]),.doutc(w_n20910_17[2]),.din(w_n20910_5[1]));
	jspl jspl_w_n20913_0(.douta(w_n20913_0[0]),.doutb(w_n20913_0[1]),.din(n20913));
	jspl jspl_w_n20918_0(.douta(w_n20918_0[0]),.doutb(w_n20918_0[1]),.din(n20918));
	jspl jspl_w_n20921_0(.douta(w_n20921_0[0]),.doutb(w_n20921_0[1]),.din(n20921));
	jspl jspl_w_n20924_0(.douta(w_n20924_0[0]),.doutb(w_n20924_0[1]),.din(n20924));
	jspl jspl_w_n20934_0(.douta(w_n20934_0[0]),.doutb(w_n20934_0[1]),.din(n20934));
	jspl jspl_w_n20942_0(.douta(w_n20942_0[0]),.doutb(w_n20942_0[1]),.din(n20942));
	jspl jspl_w_n20950_0(.douta(w_n20950_0[0]),.doutb(w_n20950_0[1]),.din(n20950));
	jspl jspl_w_n20955_0(.douta(w_n20955_0[0]),.doutb(w_n20955_0[1]),.din(n20955));
	jspl jspl_w_n20960_0(.douta(w_n20960_0[0]),.doutb(w_n20960_0[1]),.din(n20960));
	jspl jspl_w_n20967_0(.douta(w_n20967_0[0]),.doutb(w_n20967_0[1]),.din(n20967));
	jspl jspl_w_n20975_0(.douta(w_n20975_0[0]),.doutb(w_n20975_0[1]),.din(n20975));
	jspl jspl_w_n20982_0(.douta(w_n20982_0[0]),.doutb(w_n20982_0[1]),.din(n20982));
	jspl jspl_w_n20989_0(.douta(w_n20989_0[0]),.doutb(w_n20989_0[1]),.din(n20989));
	jspl jspl_w_n20994_0(.douta(w_n20994_0[0]),.doutb(w_n20994_0[1]),.din(n20994));
	jspl jspl_w_n21001_0(.douta(w_n21001_0[0]),.doutb(w_n21001_0[1]),.din(n21001));
	jspl jspl_w_n21009_0(.douta(w_n21009_0[0]),.doutb(w_n21009_0[1]),.din(n21009));
	jspl jspl_w_n21016_0(.douta(w_n21016_0[0]),.doutb(w_n21016_0[1]),.din(n21016));
	jspl jspl_w_n21021_0(.douta(w_n21021_0[0]),.doutb(w_n21021_0[1]),.din(n21021));
	jspl jspl_w_n21028_0(.douta(w_n21028_0[0]),.doutb(w_n21028_0[1]),.din(n21028));
	jspl jspl_w_n21033_0(.douta(w_n21033_0[0]),.doutb(w_n21033_0[1]),.din(n21033));
	jspl jspl_w_n21040_0(.douta(w_n21040_0[0]),.doutb(w_n21040_0[1]),.din(n21040));
	jspl jspl_w_n21048_0(.douta(w_n21048_0[0]),.doutb(w_n21048_0[1]),.din(n21048));
	jspl jspl_w_n21055_0(.douta(w_n21055_0[0]),.doutb(w_n21055_0[1]),.din(n21055));
	jspl jspl_w_n21060_0(.douta(w_n21060_0[0]),.doutb(w_n21060_0[1]),.din(n21060));
	jspl jspl_w_n21067_0(.douta(w_n21067_0[0]),.doutb(w_n21067_0[1]),.din(n21067));
	jspl jspl_w_n21072_0(.douta(w_n21072_0[0]),.doutb(w_n21072_0[1]),.din(n21072));
	jspl jspl_w_n21079_0(.douta(w_n21079_0[0]),.doutb(w_n21079_0[1]),.din(n21079));
	jspl jspl_w_n21087_0(.douta(w_n21087_0[0]),.doutb(w_n21087_0[1]),.din(n21087));
	jspl jspl_w_n21094_0(.douta(w_n21094_0[0]),.doutb(w_n21094_0[1]),.din(n21094));
	jspl jspl_w_n21099_0(.douta(w_n21099_0[0]),.doutb(w_n21099_0[1]),.din(n21099));
	jspl jspl_w_n21106_0(.douta(w_n21106_0[0]),.doutb(w_n21106_0[1]),.din(n21106));
	jspl jspl_w_n21111_0(.douta(w_n21111_0[0]),.doutb(w_n21111_0[1]),.din(n21111));
	jspl jspl_w_n21118_0(.douta(w_n21118_0[0]),.doutb(w_n21118_0[1]),.din(n21118));
	jspl jspl_w_n21126_0(.douta(w_n21126_0[0]),.doutb(w_n21126_0[1]),.din(n21126));
	jspl jspl_w_n21133_0(.douta(w_n21133_0[0]),.doutb(w_n21133_0[1]),.din(n21133));
	jspl jspl_w_n21138_0(.douta(w_n21138_0[0]),.doutb(w_n21138_0[1]),.din(n21138));
	jspl jspl_w_n21145_0(.douta(w_n21145_0[0]),.doutb(w_n21145_0[1]),.din(n21145));
	jspl jspl_w_n21150_0(.douta(w_n21150_0[0]),.doutb(w_n21150_0[1]),.din(n21150));
	jspl jspl_w_n21157_0(.douta(w_n21157_0[0]),.doutb(w_n21157_0[1]),.din(n21157));
	jspl jspl_w_n21165_0(.douta(w_n21165_0[0]),.doutb(w_n21165_0[1]),.din(n21165));
	jspl jspl_w_n21172_0(.douta(w_n21172_0[0]),.doutb(w_n21172_0[1]),.din(n21172));
	jspl jspl_w_n21177_0(.douta(w_n21177_0[0]),.doutb(w_n21177_0[1]),.din(n21177));
	jspl jspl_w_n21184_0(.douta(w_n21184_0[0]),.doutb(w_n21184_0[1]),.din(n21184));
	jspl jspl_w_n21189_0(.douta(w_n21189_0[0]),.doutb(w_n21189_0[1]),.din(n21189));
	jspl jspl_w_n21196_0(.douta(w_n21196_0[0]),.doutb(w_n21196_0[1]),.din(n21196));
	jspl jspl_w_n21204_0(.douta(w_n21204_0[0]),.doutb(w_n21204_0[1]),.din(n21204));
	jspl jspl_w_n21211_0(.douta(w_n21211_0[0]),.doutb(w_n21211_0[1]),.din(n21211));
	jspl jspl_w_n21216_0(.douta(w_n21216_0[0]),.doutb(w_n21216_0[1]),.din(n21216));
	jspl jspl_w_n21223_0(.douta(w_n21223_0[0]),.doutb(w_n21223_0[1]),.din(n21223));
	jspl jspl_w_n21228_0(.douta(w_n21228_0[0]),.doutb(w_n21228_0[1]),.din(n21228));
	jspl jspl_w_n21235_0(.douta(w_n21235_0[0]),.doutb(w_n21235_0[1]),.din(n21235));
	jspl jspl_w_n21243_0(.douta(w_n21243_0[0]),.doutb(w_n21243_0[1]),.din(n21243));
	jspl jspl_w_n21250_0(.douta(w_n21250_0[0]),.doutb(w_n21250_0[1]),.din(n21250));
	jspl jspl_w_n21255_0(.douta(w_n21255_0[0]),.doutb(w_n21255_0[1]),.din(n21255));
	jspl jspl_w_n21262_0(.douta(w_n21262_0[0]),.doutb(w_n21262_0[1]),.din(n21262));
	jspl jspl_w_n21267_0(.douta(w_n21267_0[0]),.doutb(w_n21267_0[1]),.din(n21267));
	jspl jspl_w_n21274_0(.douta(w_n21274_0[0]),.doutb(w_n21274_0[1]),.din(n21274));
	jspl jspl_w_n21282_0(.douta(w_n21282_0[0]),.doutb(w_n21282_0[1]),.din(n21282));
	jspl jspl_w_n21289_0(.douta(w_n21289_0[0]),.doutb(w_n21289_0[1]),.din(n21289));
	jspl jspl_w_n21294_0(.douta(w_n21294_0[0]),.doutb(w_n21294_0[1]),.din(n21294));
	jspl jspl_w_n21301_0(.douta(w_n21301_0[0]),.doutb(w_n21301_0[1]),.din(n21301));
	jspl jspl_w_n21306_0(.douta(w_n21306_0[0]),.doutb(w_n21306_0[1]),.din(n21306));
	jspl jspl_w_n21313_0(.douta(w_n21313_0[0]),.doutb(w_n21313_0[1]),.din(n21313));
	jspl jspl_w_n21321_0(.douta(w_n21321_0[0]),.doutb(w_n21321_0[1]),.din(n21321));
	jspl jspl_w_n21328_0(.douta(w_n21328_0[0]),.doutb(w_n21328_0[1]),.din(n21328));
	jspl jspl_w_n21333_0(.douta(w_n21333_0[0]),.doutb(w_n21333_0[1]),.din(n21333));
	jspl jspl_w_n21340_0(.douta(w_n21340_0[0]),.doutb(w_n21340_0[1]),.din(n21340));
	jspl jspl_w_n21345_0(.douta(w_n21345_0[0]),.doutb(w_n21345_0[1]),.din(n21345));
	jspl jspl_w_n21352_0(.douta(w_n21352_0[0]),.doutb(w_n21352_0[1]),.din(n21352));
	jspl jspl_w_n21360_0(.douta(w_n21360_0[0]),.doutb(w_n21360_0[1]),.din(n21360));
	jspl jspl_w_n21367_0(.douta(w_n21367_0[0]),.doutb(w_n21367_0[1]),.din(n21367));
	jspl jspl_w_n21372_0(.douta(w_n21372_0[0]),.doutb(w_n21372_0[1]),.din(n21372));
	jspl jspl_w_n21379_0(.douta(w_n21379_0[0]),.doutb(w_n21379_0[1]),.din(n21379));
	jspl jspl_w_n21384_0(.douta(w_n21384_0[0]),.doutb(w_n21384_0[1]),.din(n21384));
	jspl jspl_w_n21391_0(.douta(w_n21391_0[0]),.doutb(w_n21391_0[1]),.din(n21391));
	jspl jspl_w_n21399_0(.douta(w_n21399_0[0]),.doutb(w_n21399_0[1]),.din(n21399));
	jspl jspl_w_n21406_0(.douta(w_n21406_0[0]),.doutb(w_n21406_0[1]),.din(n21406));
	jspl jspl_w_n21411_0(.douta(w_n21411_0[0]),.doutb(w_n21411_0[1]),.din(n21411));
	jspl jspl_w_n21418_0(.douta(w_n21418_0[0]),.doutb(w_n21418_0[1]),.din(n21418));
	jspl jspl_w_n21423_0(.douta(w_n21423_0[0]),.doutb(w_n21423_0[1]),.din(n21423));
	jspl jspl_w_n21430_0(.douta(w_n21430_0[0]),.doutb(w_n21430_0[1]),.din(n21430));
	jspl jspl_w_n21438_0(.douta(w_n21438_0[0]),.doutb(w_n21438_0[1]),.din(n21438));
	jspl jspl_w_n21445_0(.douta(w_n21445_0[0]),.doutb(w_n21445_0[1]),.din(n21445));
	jspl jspl_w_n21450_0(.douta(w_n21450_0[0]),.doutb(w_n21450_0[1]),.din(n21450));
	jspl jspl_w_n21457_0(.douta(w_n21457_0[0]),.doutb(w_n21457_0[1]),.din(n21457));
	jspl jspl_w_n21462_0(.douta(w_n21462_0[0]),.doutb(w_n21462_0[1]),.din(n21462));
	jspl jspl_w_n21469_0(.douta(w_n21469_0[0]),.doutb(w_n21469_0[1]),.din(n21469));
	jspl jspl_w_n21476_0(.douta(w_n21476_0[0]),.doutb(w_n21476_0[1]),.din(n21476));
	jspl jspl_w_n21481_0(.douta(w_n21481_0[0]),.doutb(w_n21481_0[1]),.din(n21481));
	jspl jspl_w_n21490_0(.douta(w_n21490_0[0]),.doutb(w_n21490_0[1]),.din(n21490));
	jspl jspl_w_n21494_0(.douta(w_n21494_0[0]),.doutb(w_n21494_0[1]),.din(n21494));
	jspl jspl_w_n21496_0(.douta(w_n21496_0[0]),.doutb(w_n21496_0[1]),.din(n21496));
endmodule

