// Benchmark "top" written by ABC on Wed May 27 23:36:55 2020

module gf_decoder ( 
    count0 , count1 , count2 , count3 , count4 , count5 ,
    count6 , count7 ,
    selectp10 , selectp11 , selectp12 , selectp13 ,
    selectp14 , selectp15 , selectp16 , selectp17 ,
    selectp18 , selectp19 , selectp110 , selectp111 ,
    selectp112 , selectp113 , selectp114 , selectp115 ,
    selectp116 , selectp117 , selectp118 , selectp119 ,
    selectp120 , selectp121 , selectp122 , selectp123 ,
    selectp124 , selectp125 , selectp126 , selectp127 ,
    selectp128 , selectp129 , selectp130 , selectp131 ,
    selectp132 , selectp133 , selectp134 , selectp135 ,
    selectp136 , selectp137 , selectp138 , selectp139 ,
    selectp140 , selectp141 , selectp142 , selectp143 ,
    selectp144 , selectp145 , selectp146 , selectp147 ,
    selectp148 , selectp149 , selectp150 , selectp151 ,
    selectp152 , selectp153 , selectp154 , selectp155 ,
    selectp156 , selectp157 , selectp158 , selectp159 ,
    selectp160 , selectp161 , selectp162 , selectp163 ,
    selectp164 , selectp165 , selectp166 , selectp167 ,
    selectp168 , selectp169 , selectp170 , selectp171 ,
    selectp172 , selectp173 , selectp174 , selectp175 ,
    selectp176 , selectp177 , selectp178 , selectp179 ,
    selectp180 , selectp181 , selectp182 , selectp183 ,
    selectp184 , selectp185 , selectp186 , selectp187 ,
    selectp188 , selectp189 , selectp190 , selectp191 ,
    selectp192 , selectp193 , selectp194 , selectp195 ,
    selectp196 , selectp197 , selectp198 , selectp199 ,
    selectp1100 , selectp1101 , selectp1102 , selectp1103 ,
    selectp1104 , selectp1105 , selectp1106 , selectp1107 ,
    selectp1108 , selectp1109 , selectp1110 , selectp1111 ,
    selectp1112 , selectp1113 , selectp1114 , selectp1115 ,
    selectp1116 , selectp1117 , selectp1118 , selectp1119 ,
    selectp1120 , selectp1121 , selectp1122 , selectp1123 ,
    selectp1124 , selectp1125 , selectp1126 , selectp1127 ,
    selectp20 , selectp21 , selectp22 , selectp23 ,
    selectp24 , selectp25 , selectp26 , selectp27 ,
    selectp28 , selectp29 , selectp210 , selectp211 ,
    selectp212 , selectp213 , selectp214 , selectp215 ,
    selectp216 , selectp217 , selectp218 , selectp219 ,
    selectp220 , selectp221 , selectp222 , selectp223 ,
    selectp224 , selectp225 , selectp226 , selectp227 ,
    selectp228 , selectp229 , selectp230 , selectp231 ,
    selectp232 , selectp233 , selectp234 , selectp235 ,
    selectp236 , selectp237 , selectp238 , selectp239 ,
    selectp240 , selectp241 , selectp242 , selectp243 ,
    selectp244 , selectp245 , selectp246 , selectp247 ,
    selectp248 , selectp249 , selectp250 , selectp251 ,
    selectp252 , selectp253 , selectp254 , selectp255 ,
    selectp256 , selectp257 , selectp258 , selectp259 ,
    selectp260 , selectp261 , selectp262 , selectp263 ,
    selectp264 , selectp265 , selectp266 , selectp267 ,
    selectp268 , selectp269 , selectp270 , selectp271 ,
    selectp272 , selectp273 , selectp274 , selectp275 ,
    selectp276 , selectp277 , selectp278 , selectp279 ,
    selectp280 , selectp281 , selectp282 , selectp283 ,
    selectp284 , selectp285 , selectp286 , selectp287 ,
    selectp288 , selectp289 , selectp290 , selectp291 ,
    selectp292 , selectp293 , selectp294 , selectp295 ,
    selectp296 , selectp297 , selectp298 , selectp299 ,
    selectp2100 , selectp2101 , selectp2102 , selectp2103 ,
    selectp2104 , selectp2105 , selectp2106 , selectp2107 ,
    selectp2108 , selectp2109 , selectp2110 , selectp2111 ,
    selectp2112 , selectp2113 , selectp2114 , selectp2115 ,
    selectp2116 , selectp2117 , selectp2118 , selectp2119 ,
    selectp2120 , selectp2121 , selectp2122 , selectp2123 ,
    selectp2124 , selectp2125 , selectp2126 , selectp2127   );
  input  count0 , count1 , count2 , count3 , count4 ,
    count5 , count6 , count7 ;
  output selectp10 , selectp11 , selectp12 , selectp13 ,
    selectp14 , selectp15 , selectp16 , selectp17 ,
    selectp18 , selectp19 , selectp110 , selectp111 ,
    selectp112 , selectp113 , selectp114 , selectp115 ,
    selectp116 , selectp117 , selectp118 , selectp119 ,
    selectp120 , selectp121 , selectp122 , selectp123 ,
    selectp124 , selectp125 , selectp126 , selectp127 ,
    selectp128 , selectp129 , selectp130 , selectp131 ,
    selectp132 , selectp133 , selectp134 , selectp135 ,
    selectp136 , selectp137 , selectp138 , selectp139 ,
    selectp140 , selectp141 , selectp142 , selectp143 ,
    selectp144 , selectp145 , selectp146 , selectp147 ,
    selectp148 , selectp149 , selectp150 , selectp151 ,
    selectp152 , selectp153 , selectp154 , selectp155 ,
    selectp156 , selectp157 , selectp158 , selectp159 ,
    selectp160 , selectp161 , selectp162 , selectp163 ,
    selectp164 , selectp165 , selectp166 , selectp167 ,
    selectp168 , selectp169 , selectp170 , selectp171 ,
    selectp172 , selectp173 , selectp174 , selectp175 ,
    selectp176 , selectp177 , selectp178 , selectp179 ,
    selectp180 , selectp181 , selectp182 , selectp183 ,
    selectp184 , selectp185 , selectp186 , selectp187 ,
    selectp188 , selectp189 , selectp190 , selectp191 ,
    selectp192 , selectp193 , selectp194 , selectp195 ,
    selectp196 , selectp197 , selectp198 , selectp199 ,
    selectp1100 , selectp1101 , selectp1102 , selectp1103 ,
    selectp1104 , selectp1105 , selectp1106 , selectp1107 ,
    selectp1108 , selectp1109 , selectp1110 , selectp1111 ,
    selectp1112 , selectp1113 , selectp1114 , selectp1115 ,
    selectp1116 , selectp1117 , selectp1118 , selectp1119 ,
    selectp1120 , selectp1121 , selectp1122 , selectp1123 ,
    selectp1124 , selectp1125 , selectp1126 , selectp1127 ,
    selectp20 , selectp21 , selectp22 , selectp23 ,
    selectp24 , selectp25 , selectp26 , selectp27 ,
    selectp28 , selectp29 , selectp210 , selectp211 ,
    selectp212 , selectp213 , selectp214 , selectp215 ,
    selectp216 , selectp217 , selectp218 , selectp219 ,
    selectp220 , selectp221 , selectp222 , selectp223 ,
    selectp224 , selectp225 , selectp226 , selectp227 ,
    selectp228 , selectp229 , selectp230 , selectp231 ,
    selectp232 , selectp233 , selectp234 , selectp235 ,
    selectp236 , selectp237 , selectp238 , selectp239 ,
    selectp240 , selectp241 , selectp242 , selectp243 ,
    selectp244 , selectp245 , selectp246 , selectp247 ,
    selectp248 , selectp249 , selectp250 , selectp251 ,
    selectp252 , selectp253 , selectp254 , selectp255 ,
    selectp256 , selectp257 , selectp258 , selectp259 ,
    selectp260 , selectp261 , selectp262 , selectp263 ,
    selectp264 , selectp265 , selectp266 , selectp267 ,
    selectp268 , selectp269 , selectp270 , selectp271 ,
    selectp272 , selectp273 , selectp274 , selectp275 ,
    selectp276 , selectp277 , selectp278 , selectp279 ,
    selectp280 , selectp281 , selectp282 , selectp283 ,
    selectp284 , selectp285 , selectp286 , selectp287 ,
    selectp288 , selectp289 , selectp290 , selectp291 ,
    selectp292 , selectp293 , selectp294 , selectp295 ,
    selectp296 , selectp297 , selectp298 , selectp299 ,
    selectp2100 , selectp2101 , selectp2102 , selectp2103 ,
    selectp2104 , selectp2105 , selectp2106 , selectp2107 ,
    selectp2108 , selectp2109 , selectp2110 , selectp2111 ,
    selectp2112 , selectp2113 , selectp2114 , selectp2115 ,
    selectp2116 , selectp2117 , selectp2118 , selectp2119 ,
    selectp2120 , selectp2121 , selectp2122 , selectp2123 ,
    selectp2124 , selectp2125 , selectp2126 , selectp2127 ;
  wire n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
    n275, n276, n278, n279, n281, n282, n284, n286, n287, n289, n290, n292,
    n294, n296, n297, n299, n301, n302, n304, n306, n308, n310, n312, n314,
    n315, n332, n333, n350, n351, n368, n369, n386, n403, n420, n437, n438,
    n439, n456, n473, n490, n507, n508, n525, n542, n559;
  jnot g000(.din(count4 ), .dout(n264));
  jnot g001(.din(count5 ), .dout(n265));
  jand g002(.dina(n265), .dinb(n264), .dout(n266));
  jnot g003(.din(count6 ), .dout(n267));
  jand g004(.dina(count7 ), .dinb(n267), .dout(n268));
  jand g005(.dina(n268), .dinb(n266), .dout(n269));
  jnot g006(.din(count0 ), .dout(n270));
  jnot g007(.din(count2 ), .dout(n271));
  jand g008(.dina(n271), .dinb(n270), .dout(n272));
  jnot g009(.din(count1 ), .dout(n273));
  jnot g010(.din(count3 ), .dout(n274));
  jand g011(.dina(n274), .dinb(n273), .dout(n275));
  jand g012(.dina(n275), .dinb(n272), .dout(n276));
  jand g013(.dina(n276), .dinb(n269), .dout(selectp10 ));
  jand g014(.dina(n271), .dinb(count0 ), .dout(n278));
  jand g015(.dina(n278), .dinb(n275), .dout(n279));
  jand g016(.dina(n279), .dinb(n269), .dout(selectp11 ));
  jand g017(.dina(n274), .dinb(count1 ), .dout(n281));
  jand g018(.dina(n281), .dinb(n272), .dout(n282));
  jand g019(.dina(n282), .dinb(n269), .dout(selectp12 ));
  jand g020(.dina(n281), .dinb(n278), .dout(n284));
  jand g021(.dina(n284), .dinb(n269), .dout(selectp13 ));
  jand g022(.dina(count2 ), .dinb(n270), .dout(n286));
  jand g023(.dina(n286), .dinb(n275), .dout(n287));
  jand g024(.dina(n287), .dinb(n269), .dout(selectp14 ));
  jand g025(.dina(count2 ), .dinb(count0 ), .dout(n289));
  jand g026(.dina(n289), .dinb(n275), .dout(n290));
  jand g027(.dina(n290), .dinb(n269), .dout(selectp15 ));
  jand g028(.dina(n286), .dinb(n281), .dout(n292));
  jand g029(.dina(n292), .dinb(n269), .dout(selectp16 ));
  jand g030(.dina(n289), .dinb(n281), .dout(n294));
  jand g031(.dina(n294), .dinb(n269), .dout(selectp17 ));
  jand g032(.dina(count3 ), .dinb(n273), .dout(n296));
  jand g033(.dina(n296), .dinb(n272), .dout(n297));
  jand g034(.dina(n297), .dinb(n269), .dout(selectp18 ));
  jand g035(.dina(n296), .dinb(n278), .dout(n299));
  jand g036(.dina(n299), .dinb(n269), .dout(selectp19 ));
  jand g037(.dina(count3 ), .dinb(count1 ), .dout(n301));
  jand g038(.dina(n301), .dinb(n272), .dout(n302));
  jand g039(.dina(n302), .dinb(n269), .dout(selectp110 ));
  jand g040(.dina(n301), .dinb(n278), .dout(n304));
  jand g041(.dina(n304), .dinb(n269), .dout(selectp111 ));
  jand g042(.dina(n296), .dinb(n286), .dout(n306));
  jand g043(.dina(n306), .dinb(n269), .dout(selectp112 ));
  jand g044(.dina(n296), .dinb(n289), .dout(n308));
  jand g045(.dina(n308), .dinb(n269), .dout(selectp113 ));
  jand g046(.dina(n301), .dinb(n286), .dout(n310));
  jand g047(.dina(n310), .dinb(n269), .dout(selectp114 ));
  jand g048(.dina(n301), .dinb(n289), .dout(n312));
  jand g049(.dina(n312), .dinb(n269), .dout(selectp115 ));
  jand g050(.dina(n265), .dinb(count4 ), .dout(n314));
  jand g051(.dina(n314), .dinb(n268), .dout(n315));
  jand g052(.dina(n315), .dinb(n276), .dout(selectp116 ));
  jand g053(.dina(n315), .dinb(n279), .dout(selectp117 ));
  jand g054(.dina(n315), .dinb(n282), .dout(selectp118 ));
  jand g055(.dina(n315), .dinb(n284), .dout(selectp119 ));
  jand g056(.dina(n315), .dinb(n287), .dout(selectp120 ));
  jand g057(.dina(n315), .dinb(n290), .dout(selectp121 ));
  jand g058(.dina(n315), .dinb(n292), .dout(selectp122 ));
  jand g059(.dina(n315), .dinb(n294), .dout(selectp123 ));
  jand g060(.dina(n315), .dinb(n297), .dout(selectp124 ));
  jand g061(.dina(n315), .dinb(n299), .dout(selectp125 ));
  jand g062(.dina(n315), .dinb(n302), .dout(selectp126 ));
  jand g063(.dina(n315), .dinb(n304), .dout(selectp127 ));
  jand g064(.dina(n315), .dinb(n306), .dout(selectp128 ));
  jand g065(.dina(n315), .dinb(n308), .dout(selectp129 ));
  jand g066(.dina(n315), .dinb(n310), .dout(selectp130 ));
  jand g067(.dina(n315), .dinb(n312), .dout(selectp131 ));
  jand g068(.dina(count5 ), .dinb(n264), .dout(n332));
  jand g069(.dina(n332), .dinb(n268), .dout(n333));
  jand g070(.dina(n333), .dinb(n276), .dout(selectp132 ));
  jand g071(.dina(n333), .dinb(n279), .dout(selectp133 ));
  jand g072(.dina(n333), .dinb(n282), .dout(selectp134 ));
  jand g073(.dina(n333), .dinb(n284), .dout(selectp135 ));
  jand g074(.dina(n333), .dinb(n287), .dout(selectp136 ));
  jand g075(.dina(n333), .dinb(n290), .dout(selectp137 ));
  jand g076(.dina(n333), .dinb(n292), .dout(selectp138 ));
  jand g077(.dina(n333), .dinb(n294), .dout(selectp139 ));
  jand g078(.dina(n333), .dinb(n297), .dout(selectp140 ));
  jand g079(.dina(n333), .dinb(n299), .dout(selectp141 ));
  jand g080(.dina(n333), .dinb(n302), .dout(selectp142 ));
  jand g081(.dina(n333), .dinb(n304), .dout(selectp143 ));
  jand g082(.dina(n333), .dinb(n306), .dout(selectp144 ));
  jand g083(.dina(n333), .dinb(n308), .dout(selectp145 ));
  jand g084(.dina(n333), .dinb(n310), .dout(selectp146 ));
  jand g085(.dina(n333), .dinb(n312), .dout(selectp147 ));
  jand g086(.dina(count5 ), .dinb(count4 ), .dout(n350));
  jand g087(.dina(n350), .dinb(n268), .dout(n351));
  jand g088(.dina(n351), .dinb(n276), .dout(selectp148 ));
  jand g089(.dina(n351), .dinb(n279), .dout(selectp149 ));
  jand g090(.dina(n351), .dinb(n282), .dout(selectp150 ));
  jand g091(.dina(n351), .dinb(n284), .dout(selectp151 ));
  jand g092(.dina(n351), .dinb(n287), .dout(selectp152 ));
  jand g093(.dina(n351), .dinb(n290), .dout(selectp153 ));
  jand g094(.dina(n351), .dinb(n292), .dout(selectp154 ));
  jand g095(.dina(n351), .dinb(n294), .dout(selectp155 ));
  jand g096(.dina(n351), .dinb(n297), .dout(selectp156 ));
  jand g097(.dina(n351), .dinb(n299), .dout(selectp157 ));
  jand g098(.dina(n351), .dinb(n302), .dout(selectp158 ));
  jand g099(.dina(n351), .dinb(n304), .dout(selectp159 ));
  jand g100(.dina(n351), .dinb(n306), .dout(selectp160 ));
  jand g101(.dina(n351), .dinb(n308), .dout(selectp161 ));
  jand g102(.dina(n351), .dinb(n310), .dout(selectp162 ));
  jand g103(.dina(n351), .dinb(n312), .dout(selectp163 ));
  jand g104(.dina(count7 ), .dinb(count6 ), .dout(n368));
  jand g105(.dina(n368), .dinb(n266), .dout(n369));
  jand g106(.dina(n369), .dinb(n276), .dout(selectp164 ));
  jand g107(.dina(n369), .dinb(n279), .dout(selectp165 ));
  jand g108(.dina(n369), .dinb(n282), .dout(selectp166 ));
  jand g109(.dina(n369), .dinb(n284), .dout(selectp167 ));
  jand g110(.dina(n369), .dinb(n287), .dout(selectp168 ));
  jand g111(.dina(n369), .dinb(n290), .dout(selectp169 ));
  jand g112(.dina(n369), .dinb(n292), .dout(selectp170 ));
  jand g113(.dina(n369), .dinb(n294), .dout(selectp171 ));
  jand g114(.dina(n369), .dinb(n297), .dout(selectp172 ));
  jand g115(.dina(n369), .dinb(n299), .dout(selectp173 ));
  jand g116(.dina(n369), .dinb(n302), .dout(selectp174 ));
  jand g117(.dina(n369), .dinb(n304), .dout(selectp175 ));
  jand g118(.dina(n369), .dinb(n306), .dout(selectp176 ));
  jand g119(.dina(n369), .dinb(n308), .dout(selectp177 ));
  jand g120(.dina(n369), .dinb(n310), .dout(selectp178 ));
  jand g121(.dina(n369), .dinb(n312), .dout(selectp179 ));
  jand g122(.dina(n368), .dinb(n314), .dout(n386));
  jand g123(.dina(n386), .dinb(n276), .dout(selectp180 ));
  jand g124(.dina(n386), .dinb(n279), .dout(selectp181 ));
  jand g125(.dina(n386), .dinb(n282), .dout(selectp182 ));
  jand g126(.dina(n386), .dinb(n284), .dout(selectp183 ));
  jand g127(.dina(n386), .dinb(n287), .dout(selectp184 ));
  jand g128(.dina(n386), .dinb(n290), .dout(selectp185 ));
  jand g129(.dina(n386), .dinb(n292), .dout(selectp186 ));
  jand g130(.dina(n386), .dinb(n294), .dout(selectp187 ));
  jand g131(.dina(n386), .dinb(n297), .dout(selectp188 ));
  jand g132(.dina(n386), .dinb(n299), .dout(selectp189 ));
  jand g133(.dina(n386), .dinb(n302), .dout(selectp190 ));
  jand g134(.dina(n386), .dinb(n304), .dout(selectp191 ));
  jand g135(.dina(n386), .dinb(n306), .dout(selectp192 ));
  jand g136(.dina(n386), .dinb(n308), .dout(selectp193 ));
  jand g137(.dina(n386), .dinb(n310), .dout(selectp194 ));
  jand g138(.dina(n386), .dinb(n312), .dout(selectp195 ));
  jand g139(.dina(n368), .dinb(n332), .dout(n403));
  jand g140(.dina(n403), .dinb(n276), .dout(selectp196 ));
  jand g141(.dina(n403), .dinb(n279), .dout(selectp197 ));
  jand g142(.dina(n403), .dinb(n282), .dout(selectp198 ));
  jand g143(.dina(n403), .dinb(n284), .dout(selectp199 ));
  jand g144(.dina(n403), .dinb(n287), .dout(selectp1100 ));
  jand g145(.dina(n403), .dinb(n290), .dout(selectp1101 ));
  jand g146(.dina(n403), .dinb(n292), .dout(selectp1102 ));
  jand g147(.dina(n403), .dinb(n294), .dout(selectp1103 ));
  jand g148(.dina(n403), .dinb(n297), .dout(selectp1104 ));
  jand g149(.dina(n403), .dinb(n299), .dout(selectp1105 ));
  jand g150(.dina(n403), .dinb(n302), .dout(selectp1106 ));
  jand g151(.dina(n403), .dinb(n304), .dout(selectp1107 ));
  jand g152(.dina(n403), .dinb(n306), .dout(selectp1108 ));
  jand g153(.dina(n403), .dinb(n308), .dout(selectp1109 ));
  jand g154(.dina(n403), .dinb(n310), .dout(selectp1110 ));
  jand g155(.dina(n403), .dinb(n312), .dout(selectp1111 ));
  jand g156(.dina(n368), .dinb(n350), .dout(n420));
  jand g157(.dina(n420), .dinb(n276), .dout(selectp1112 ));
  jand g158(.dina(n420), .dinb(n279), .dout(selectp1113 ));
  jand g159(.dina(n420), .dinb(n282), .dout(selectp1114 ));
  jand g160(.dina(n420), .dinb(n284), .dout(selectp1115 ));
  jand g161(.dina(n420), .dinb(n287), .dout(selectp1116 ));
  jand g162(.dina(n420), .dinb(n290), .dout(selectp1117 ));
  jand g163(.dina(n420), .dinb(n292), .dout(selectp1118 ));
  jand g164(.dina(n420), .dinb(n294), .dout(selectp1119 ));
  jand g165(.dina(n420), .dinb(n297), .dout(selectp1120 ));
  jand g166(.dina(n420), .dinb(n299), .dout(selectp1121 ));
  jand g167(.dina(n420), .dinb(n302), .dout(selectp1122 ));
  jand g168(.dina(n420), .dinb(n304), .dout(selectp1123 ));
  jand g169(.dina(n420), .dinb(n306), .dout(selectp1124 ));
  jand g170(.dina(n420), .dinb(n308), .dout(selectp1125 ));
  jand g171(.dina(n420), .dinb(n310), .dout(selectp1126 ));
  jand g172(.dina(n420), .dinb(n312), .dout(selectp1127 ));
  jnot g173(.din(count7 ), .dout(n437));
  jand g174(.dina(n437), .dinb(n267), .dout(n438));
  jand g175(.dina(n438), .dinb(n266), .dout(n439));
  jand g176(.dina(n439), .dinb(n276), .dout(selectp20 ));
  jand g177(.dina(n439), .dinb(n279), .dout(selectp21 ));
  jand g178(.dina(n439), .dinb(n282), .dout(selectp22 ));
  jand g179(.dina(n439), .dinb(n284), .dout(selectp23 ));
  jand g180(.dina(n439), .dinb(n287), .dout(selectp24 ));
  jand g181(.dina(n439), .dinb(n290), .dout(selectp25 ));
  jand g182(.dina(n439), .dinb(n292), .dout(selectp26 ));
  jand g183(.dina(n439), .dinb(n294), .dout(selectp27 ));
  jand g184(.dina(n439), .dinb(n297), .dout(selectp28 ));
  jand g185(.dina(n439), .dinb(n299), .dout(selectp29 ));
  jand g186(.dina(n439), .dinb(n302), .dout(selectp210 ));
  jand g187(.dina(n439), .dinb(n304), .dout(selectp211 ));
  jand g188(.dina(n439), .dinb(n306), .dout(selectp212 ));
  jand g189(.dina(n439), .dinb(n308), .dout(selectp213 ));
  jand g190(.dina(n439), .dinb(n310), .dout(selectp214 ));
  jand g191(.dina(n439), .dinb(n312), .dout(selectp215 ));
  jand g192(.dina(n438), .dinb(n314), .dout(n456));
  jand g193(.dina(n456), .dinb(n276), .dout(selectp216 ));
  jand g194(.dina(n456), .dinb(n279), .dout(selectp217 ));
  jand g195(.dina(n456), .dinb(n282), .dout(selectp218 ));
  jand g196(.dina(n456), .dinb(n284), .dout(selectp219 ));
  jand g197(.dina(n456), .dinb(n287), .dout(selectp220 ));
  jand g198(.dina(n456), .dinb(n290), .dout(selectp221 ));
  jand g199(.dina(n456), .dinb(n292), .dout(selectp222 ));
  jand g200(.dina(n456), .dinb(n294), .dout(selectp223 ));
  jand g201(.dina(n456), .dinb(n297), .dout(selectp224 ));
  jand g202(.dina(n456), .dinb(n299), .dout(selectp225 ));
  jand g203(.dina(n456), .dinb(n302), .dout(selectp226 ));
  jand g204(.dina(n456), .dinb(n304), .dout(selectp227 ));
  jand g205(.dina(n456), .dinb(n306), .dout(selectp228 ));
  jand g206(.dina(n456), .dinb(n308), .dout(selectp229 ));
  jand g207(.dina(n456), .dinb(n310), .dout(selectp230 ));
  jand g208(.dina(n456), .dinb(n312), .dout(selectp231 ));
  jand g209(.dina(n438), .dinb(n332), .dout(n473));
  jand g210(.dina(n473), .dinb(n276), .dout(selectp232 ));
  jand g211(.dina(n473), .dinb(n279), .dout(selectp233 ));
  jand g212(.dina(n473), .dinb(n282), .dout(selectp234 ));
  jand g213(.dina(n473), .dinb(n284), .dout(selectp235 ));
  jand g214(.dina(n473), .dinb(n287), .dout(selectp236 ));
  jand g215(.dina(n473), .dinb(n290), .dout(selectp237 ));
  jand g216(.dina(n473), .dinb(n292), .dout(selectp238 ));
  jand g217(.dina(n473), .dinb(n294), .dout(selectp239 ));
  jand g218(.dina(n473), .dinb(n297), .dout(selectp240 ));
  jand g219(.dina(n473), .dinb(n299), .dout(selectp241 ));
  jand g220(.dina(n473), .dinb(n302), .dout(selectp242 ));
  jand g221(.dina(n473), .dinb(n304), .dout(selectp243 ));
  jand g222(.dina(n473), .dinb(n306), .dout(selectp244 ));
  jand g223(.dina(n473), .dinb(n308), .dout(selectp245 ));
  jand g224(.dina(n473), .dinb(n310), .dout(selectp246 ));
  jand g225(.dina(n473), .dinb(n312), .dout(selectp247 ));
  jand g226(.dina(n438), .dinb(n350), .dout(n490));
  jand g227(.dina(n490), .dinb(n276), .dout(selectp248 ));
  jand g228(.dina(n490), .dinb(n279), .dout(selectp249 ));
  jand g229(.dina(n490), .dinb(n282), .dout(selectp250 ));
  jand g230(.dina(n490), .dinb(n284), .dout(selectp251 ));
  jand g231(.dina(n490), .dinb(n287), .dout(selectp252 ));
  jand g232(.dina(n490), .dinb(n290), .dout(selectp253 ));
  jand g233(.dina(n490), .dinb(n292), .dout(selectp254 ));
  jand g234(.dina(n490), .dinb(n294), .dout(selectp255 ));
  jand g235(.dina(n490), .dinb(n297), .dout(selectp256 ));
  jand g236(.dina(n490), .dinb(n299), .dout(selectp257 ));
  jand g237(.dina(n490), .dinb(n302), .dout(selectp258 ));
  jand g238(.dina(n490), .dinb(n304), .dout(selectp259 ));
  jand g239(.dina(n490), .dinb(n306), .dout(selectp260 ));
  jand g240(.dina(n490), .dinb(n308), .dout(selectp261 ));
  jand g241(.dina(n490), .dinb(n310), .dout(selectp262 ));
  jand g242(.dina(n490), .dinb(n312), .dout(selectp263 ));
  jand g243(.dina(n437), .dinb(count6 ), .dout(n507));
  jand g244(.dina(n507), .dinb(n266), .dout(n508));
  jand g245(.dina(n508), .dinb(n276), .dout(selectp264 ));
  jand g246(.dina(n508), .dinb(n279), .dout(selectp265 ));
  jand g247(.dina(n508), .dinb(n282), .dout(selectp266 ));
  jand g248(.dina(n508), .dinb(n284), .dout(selectp267 ));
  jand g249(.dina(n508), .dinb(n287), .dout(selectp268 ));
  jand g250(.dina(n508), .dinb(n290), .dout(selectp269 ));
  jand g251(.dina(n508), .dinb(n292), .dout(selectp270 ));
  jand g252(.dina(n508), .dinb(n294), .dout(selectp271 ));
  jand g253(.dina(n508), .dinb(n297), .dout(selectp272 ));
  jand g254(.dina(n508), .dinb(n299), .dout(selectp273 ));
  jand g255(.dina(n508), .dinb(n302), .dout(selectp274 ));
  jand g256(.dina(n508), .dinb(n304), .dout(selectp275 ));
  jand g257(.dina(n508), .dinb(n306), .dout(selectp276 ));
  jand g258(.dina(n508), .dinb(n308), .dout(selectp277 ));
  jand g259(.dina(n508), .dinb(n310), .dout(selectp278 ));
  jand g260(.dina(n508), .dinb(n312), .dout(selectp279 ));
  jand g261(.dina(n507), .dinb(n314), .dout(n525));
  jand g262(.dina(n525), .dinb(n276), .dout(selectp280 ));
  jand g263(.dina(n525), .dinb(n279), .dout(selectp281 ));
  jand g264(.dina(n525), .dinb(n282), .dout(selectp282 ));
  jand g265(.dina(n525), .dinb(n284), .dout(selectp283 ));
  jand g266(.dina(n525), .dinb(n287), .dout(selectp284 ));
  jand g267(.dina(n525), .dinb(n290), .dout(selectp285 ));
  jand g268(.dina(n525), .dinb(n292), .dout(selectp286 ));
  jand g269(.dina(n525), .dinb(n294), .dout(selectp287 ));
  jand g270(.dina(n525), .dinb(n297), .dout(selectp288 ));
  jand g271(.dina(n525), .dinb(n299), .dout(selectp289 ));
  jand g272(.dina(n525), .dinb(n302), .dout(selectp290 ));
  jand g273(.dina(n525), .dinb(n304), .dout(selectp291 ));
  jand g274(.dina(n525), .dinb(n306), .dout(selectp292 ));
  jand g275(.dina(n525), .dinb(n308), .dout(selectp293 ));
  jand g276(.dina(n525), .dinb(n310), .dout(selectp294 ));
  jand g277(.dina(n525), .dinb(n312), .dout(selectp295 ));
  jand g278(.dina(n507), .dinb(n332), .dout(n542));
  jand g279(.dina(n542), .dinb(n276), .dout(selectp296 ));
  jand g280(.dina(n542), .dinb(n279), .dout(selectp297 ));
  jand g281(.dina(n542), .dinb(n282), .dout(selectp298 ));
  jand g282(.dina(n542), .dinb(n284), .dout(selectp299 ));
  jand g283(.dina(n542), .dinb(n287), .dout(selectp2100 ));
  jand g284(.dina(n542), .dinb(n290), .dout(selectp2101 ));
  jand g285(.dina(n542), .dinb(n292), .dout(selectp2102 ));
  jand g286(.dina(n542), .dinb(n294), .dout(selectp2103 ));
  jand g287(.dina(n542), .dinb(n297), .dout(selectp2104 ));
  jand g288(.dina(n542), .dinb(n299), .dout(selectp2105 ));
  jand g289(.dina(n542), .dinb(n302), .dout(selectp2106 ));
  jand g290(.dina(n542), .dinb(n304), .dout(selectp2107 ));
  jand g291(.dina(n542), .dinb(n306), .dout(selectp2108 ));
  jand g292(.dina(n542), .dinb(n308), .dout(selectp2109 ));
  jand g293(.dina(n542), .dinb(n310), .dout(selectp2110 ));
  jand g294(.dina(n542), .dinb(n312), .dout(selectp2111 ));
  jand g295(.dina(n507), .dinb(n350), .dout(n559));
  jand g296(.dina(n559), .dinb(n276), .dout(selectp2112 ));
  jand g297(.dina(n559), .dinb(n279), .dout(selectp2113 ));
  jand g298(.dina(n559), .dinb(n282), .dout(selectp2114 ));
  jand g299(.dina(n559), .dinb(n284), .dout(selectp2115 ));
  jand g300(.dina(n559), .dinb(n287), .dout(selectp2116 ));
  jand g301(.dina(n559), .dinb(n290), .dout(selectp2117 ));
  jand g302(.dina(n559), .dinb(n292), .dout(selectp2118 ));
  jand g303(.dina(n559), .dinb(n294), .dout(selectp2119 ));
  jand g304(.dina(n559), .dinb(n297), .dout(selectp2120 ));
  jand g305(.dina(n559), .dinb(n299), .dout(selectp2121 ));
  jand g306(.dina(n559), .dinb(n302), .dout(selectp2122 ));
  jand g307(.dina(n559), .dinb(n304), .dout(selectp2123 ));
  jand g308(.dina(n559), .dinb(n306), .dout(selectp2124 ));
  jand g309(.dina(n559), .dinb(n308), .dout(selectp2125 ));
  jand g310(.dina(n559), .dinb(n310), .dout(selectp2126 ));
  jand g311(.dina(n559), .dinb(n312), .dout(selectp2127 ));
endmodule


