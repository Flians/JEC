// Benchmark "c3540" written by ABC on Sun May 24 21:36:35 2020

module c3540 ( 
    G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116,
    G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200,
    G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274,
    G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698,
    G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107,
    G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190,
    G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270,
    G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire n72, n73, n74, n75, n76, n77, n79, n80, n81, n82, n83, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n129, n130, n131, n132, n133, n134, n135, n137, n138, n139,
    n140, n141, n142, n143, n144, n146, n147, n148, n149, n150, n151, n152,
    n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
    n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
    n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
    n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
    n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
    n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
    n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519, n521, n522, n523, n524, n525,
    n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n550,
    n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
    n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
    n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n599, n600,
    n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
    n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
    n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n690, n691, n692, n693, n694, n695, n696, n697,
    n698, n699, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
    n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
    n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
    n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
    n747, n748, n749, n750, n752, n753, n754, n755, n756, n757, n758, n759,
    n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
    n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
    n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
    n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
    n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
    n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
    n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
    n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
    n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
    n869, n870, n871, n872, n873, n874, n875, n876, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
    n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
    n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936, n937, n939, n940, n941, n942,
    n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
    n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
    n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n990, n991,
    n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
    n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
    n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
    n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
    n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
    n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
    n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
    n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
    n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
    n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
    n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1164, n1165,
    n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1174, n1175, n1176,
    n1177, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
    n1188, n1189;
  jnot g0000(.din(G77), .dout(n72));
  jnot g0001(.din(G50), .dout(n73));
  jnot g0002(.din(G58), .dout(n74));
  jnot g0003(.din(G68), .dout(n75));
  jand g0004(.dina(n75), .dinb(n74), .dout(n76));
  jand g0005(.dina(n76), .dinb(n73), .dout(n77));
  jand g0006(.dina(n77), .dinb(n72), .dout(G353));
  jnot g0007(.din(G97), .dout(n79));
  jnot g0008(.din(G107), .dout(n80));
  jand g0009(.dina(n80), .dinb(n79), .dout(n81));
  jnot g0010(.din(n81), .dout(n82));
  jand g0011(.dina(n82), .dinb(G87), .dout(n83));
  jnot g0012(.din(n83), .dout(G355));
  jand g0013(.dina(G20), .dinb(G1), .dout(n85));
  jnot g0014(.din(G226), .dout(n86));
  jor  g0015(.dina(n86), .dinb(n73), .dout(n87));
  jnot g0016(.din(G264), .dout(n88));
  jor  g0017(.dina(n88), .dinb(n80), .dout(n89));
  jand g0018(.dina(n89), .dinb(n87), .dout(n90));
  jnot g0019(.din(G257), .dout(n91));
  jor  g0020(.dina(n91), .dinb(n79), .dout(n92));
  jnot g0021(.din(G238), .dout(n93));
  jor  g0022(.dina(n93), .dinb(n75), .dout(n94));
  jand g0023(.dina(n94), .dinb(n92), .dout(n95));
  jand g0024(.dina(n95), .dinb(n90), .dout(n96));
  jnot g0025(.din(G87), .dout(n97));
  jnot g0026(.din(G250), .dout(n98));
  jor  g0027(.dina(n98), .dinb(n97), .dout(n99));
  jnot g0028(.din(G232), .dout(n100));
  jor  g0029(.dina(n100), .dinb(n74), .dout(n101));
  jand g0030(.dina(n101), .dinb(n99), .dout(n102));
  jnot g0031(.din(G244), .dout(n103));
  jor  g0032(.dina(n103), .dinb(n72), .dout(n104));
  jnot g0033(.din(G116), .dout(n105));
  jnot g0034(.din(G270), .dout(n106));
  jor  g0035(.dina(n106), .dinb(n105), .dout(n107));
  jand g0036(.dina(n107), .dinb(n104), .dout(n108));
  jand g0037(.dina(n108), .dinb(n102), .dout(n109));
  jand g0038(.dina(n109), .dinb(n96), .dout(n110));
  jor  g0039(.dina(n110), .dinb(n85), .dout(n111));
  jnot g0040(.din(G20), .dout(n112));
  jnot g0041(.din(G1), .dout(n113));
  jnot g0042(.din(G13), .dout(n114));
  jor  g0043(.dina(n114), .dinb(n113), .dout(n115));
  jor  g0044(.dina(n115), .dinb(n112), .dout(n116));
  jnot g0045(.din(n76), .dout(n117));
  jand g0046(.dina(n117), .dinb(G50), .dout(n118));
  jnot g0047(.din(n118), .dout(n119));
  jor  g0048(.dina(n119), .dinb(n116), .dout(n120));
  jand g0049(.dina(n114), .dinb(G1), .dout(n121));
  jand g0050(.dina(n121), .dinb(G20), .dout(n122));
  jnot g0051(.din(n122), .dout(n123));
  jand g0052(.dina(n88), .dinb(n91), .dout(n124));
  jor  g0053(.dina(n124), .dinb(n98), .dout(n125));
  jor  g0054(.dina(n125), .dinb(n123), .dout(n126));
  jand g0055(.dina(n126), .dinb(n120), .dout(n127));
  jand g0056(.dina(n127), .dinb(n111), .dout(G361));
  jxor g0057(.dina(G270), .dinb(G264), .dout(n129));
  jxor g0058(.dina(G257), .dinb(n98), .dout(n130));
  jxor g0059(.dina(n130), .dinb(n129), .dout(n131));
  jnot g0060(.din(n131), .dout(n132));
  jxor g0061(.dina(G244), .dinb(G238), .dout(n133));
  jxor g0062(.dina(G232), .dinb(n86), .dout(n134));
  jxor g0063(.dina(n134), .dinb(n133), .dout(n135));
  jxor g0064(.dina(n135), .dinb(n132), .dout(G358));
  jxor g0065(.dina(G68), .dinb(G58), .dout(n137));
  jnot g0066(.din(n137), .dout(n138));
  jxor g0067(.dina(G77), .dinb(G50), .dout(n139));
  jxor g0068(.dina(n139), .dinb(n138), .dout(n140));
  jnot g0069(.din(n140), .dout(n141));
  jxor g0070(.dina(G116), .dinb(G107), .dout(n142));
  jxor g0071(.dina(G97), .dinb(n97), .dout(n143));
  jxor g0072(.dina(n143), .dinb(n142), .dout(n144));
  jxor g0073(.dina(n144), .dinb(n141), .dout(G351));
  jnot g0074(.din(G169), .dout(n146));
  jand g0075(.dina(G13), .dinb(G1), .dout(n147));
  jnot g0076(.din(G33), .dout(n148));
  jnot g0077(.din(G41), .dout(n149));
  jor  g0078(.dina(n149), .dinb(n148), .dout(n150));
  jand g0079(.dina(n150), .dinb(n147), .dout(n151));
  jand g0080(.dina(G1698), .dinb(n148), .dout(n152));
  jand g0081(.dina(n152), .dinb(G244), .dout(n153));
  jnot g0082(.din(G1698), .dout(n154));
  jand g0083(.dina(n154), .dinb(n148), .dout(n155));
  jand g0084(.dina(n155), .dinb(G238), .dout(n156));
  jand g0085(.dina(G116), .dinb(G33), .dout(n157));
  jor  g0086(.dina(n157), .dinb(n156), .dout(n158));
  jor  g0087(.dina(n158), .dinb(n153), .dout(n159));
  jand g0088(.dina(n159), .dinb(n151), .dout(n160));
  jnot g0089(.din(G45), .dout(n161));
  jor  g0090(.dina(n161), .dinb(G1), .dout(n162));
  jand g0091(.dina(n162), .dinb(n98), .dout(n163));
  jnot g0092(.din(n163), .dout(n164));
  jand g0093(.dina(G41), .dinb(G33), .dout(n165));
  jor  g0094(.dina(n165), .dinb(n115), .dout(n166));
  jor  g0095(.dina(n162), .dinb(G274), .dout(n167));
  jand g0096(.dina(n167), .dinb(n166), .dout(n168));
  jand g0097(.dina(n168), .dinb(n164), .dout(n169));
  jor  g0098(.dina(n169), .dinb(n160), .dout(n170));
  jand g0099(.dina(n170), .dinb(n146), .dout(n171));
  jand g0100(.dina(G97), .dinb(G33), .dout(n172));
  jand g0101(.dina(G68), .dinb(n148), .dout(n173));
  jor  g0102(.dina(n173), .dinb(G20), .dout(n174));
  jor  g0103(.dina(n174), .dinb(n172), .dout(n175));
  jnot g0104(.din(n175), .dout(n176));
  jor  g0105(.dina(n112), .dinb(n113), .dout(n177));
  jor  g0106(.dina(n177), .dinb(n148), .dout(n178));
  jand g0107(.dina(n178), .dinb(n115), .dout(n179));
  jand g0108(.dina(n81), .dinb(n97), .dout(n180));
  jand g0109(.dina(n180), .dinb(G20), .dout(n181));
  jor  g0110(.dina(n181), .dinb(n179), .dout(n182));
  jor  g0111(.dina(n182), .dinb(n176), .dout(n183));
  jand g0112(.dina(G20), .dinb(n113), .dout(n184));
  jand g0113(.dina(n184), .dinb(G13), .dout(n185));
  jand g0114(.dina(n185), .dinb(n97), .dout(n186));
  jnot g0115(.din(n186), .dout(n187));
  jand g0116(.dina(n85), .dinb(G33), .dout(n188));
  jor  g0117(.dina(n188), .dinb(n147), .dout(n189));
  jor  g0118(.dina(n185), .dinb(n189), .dout(n190));
  jand g0119(.dina(G33), .dinb(n113), .dout(n191));
  jor  g0120(.dina(n191), .dinb(n97), .dout(n192));
  jor  g0121(.dina(n192), .dinb(n190), .dout(n193));
  jand g0122(.dina(n193), .dinb(n187), .dout(n194));
  jand g0123(.dina(n194), .dinb(n183), .dout(n195));
  jnot g0124(.din(G179), .dout(n196));
  jor  g0125(.dina(n154), .dinb(G33), .dout(n197));
  jor  g0126(.dina(n197), .dinb(n103), .dout(n198));
  jor  g0127(.dina(G1698), .dinb(G33), .dout(n199));
  jor  g0128(.dina(n199), .dinb(n93), .dout(n200));
  jnot g0129(.din(n157), .dout(n201));
  jand g0130(.dina(n201), .dinb(n200), .dout(n202));
  jand g0131(.dina(n202), .dinb(n198), .dout(n203));
  jor  g0132(.dina(n203), .dinb(n166), .dout(n204));
  jnot g0133(.din(G274), .dout(n205));
  jand g0134(.dina(G45), .dinb(n113), .dout(n206));
  jand g0135(.dina(n206), .dinb(n205), .dout(n207));
  jor  g0136(.dina(n207), .dinb(n151), .dout(n208));
  jor  g0137(.dina(n208), .dinb(n163), .dout(n209));
  jand g0138(.dina(n209), .dinb(n204), .dout(n210));
  jand g0139(.dina(n210), .dinb(n196), .dout(n211));
  jor  g0140(.dina(n211), .dinb(n195), .dout(n212));
  jor  g0141(.dina(n212), .dinb(n171), .dout(n213));
  jnot g0142(.din(n195), .dout(n214));
  jand g0143(.dina(n210), .dinb(G190), .dout(n215));
  jand g0144(.dina(n170), .dinb(G200), .dout(n216));
  jor  g0145(.dina(n216), .dinb(n215), .dout(n217));
  jor  g0146(.dina(n217), .dinb(n214), .dout(n218));
  jand g0147(.dina(n218), .dinb(n213), .dout(n219));
  jor  g0148(.dina(n197), .dinb(n98), .dout(n220));
  jand g0149(.dina(G283), .dinb(G33), .dout(n221));
  jnot g0150(.din(n221), .dout(n222));
  jor  g0151(.dina(n199), .dinb(n103), .dout(n223));
  jand g0152(.dina(n223), .dinb(n222), .dout(n224));
  jand g0153(.dina(n224), .dinb(n220), .dout(n225));
  jor  g0154(.dina(n225), .dinb(n166), .dout(n226));
  jor  g0155(.dina(n151), .dinb(n205), .dout(n227));
  jor  g0156(.dina(n162), .dinb(G41), .dout(n228));
  jor  g0157(.dina(n228), .dinb(n227), .dout(n229));
  jand g0158(.dina(n206), .dinb(n149), .dout(n230));
  jor  g0159(.dina(n230), .dinb(n151), .dout(n231));
  jor  g0160(.dina(n231), .dinb(n91), .dout(n232));
  jand g0161(.dina(n232), .dinb(n229), .dout(n233));
  jand g0162(.dina(n233), .dinb(n226), .dout(n234));
  jor  g0163(.dina(n234), .dinb(n146), .dout(n235));
  jand g0164(.dina(n152), .dinb(G250), .dout(n236));
  jand g0165(.dina(n155), .dinb(G244), .dout(n237));
  jor  g0166(.dina(n237), .dinb(n221), .dout(n238));
  jor  g0167(.dina(n238), .dinb(n236), .dout(n239));
  jand g0168(.dina(n239), .dinb(n151), .dout(n240));
  jand g0169(.dina(n166), .dinb(G274), .dout(n241));
  jand g0170(.dina(n230), .dinb(n241), .dout(n242));
  jand g0171(.dina(n228), .dinb(n166), .dout(n243));
  jand g0172(.dina(n243), .dinb(G257), .dout(n244));
  jor  g0173(.dina(n244), .dinb(n242), .dout(n245));
  jor  g0174(.dina(n245), .dinb(n240), .dout(n246));
  jor  g0175(.dina(n246), .dinb(n196), .dout(n247));
  jand g0176(.dina(n247), .dinb(n235), .dout(n248));
  jand g0177(.dina(G107), .dinb(G33), .dout(n249));
  jand g0178(.dina(G77), .dinb(n148), .dout(n250));
  jor  g0179(.dina(n250), .dinb(G20), .dout(n251));
  jor  g0180(.dina(n251), .dinb(n249), .dout(n252));
  jand g0181(.dina(G107), .dinb(G97), .dout(n253));
  jor  g0182(.dina(n253), .dinb(n112), .dout(n254));
  jor  g0183(.dina(n254), .dinb(n81), .dout(n255));
  jand g0184(.dina(n255), .dinb(n252), .dout(n256));
  jand g0185(.dina(n256), .dinb(n189), .dout(n257));
  jnot g0186(.din(n257), .dout(n258));
  jand g0187(.dina(n185), .dinb(n79), .dout(n259));
  jnot g0188(.din(n259), .dout(n260));
  jnot g0189(.din(n191), .dout(n261));
  jand g0190(.dina(n261), .dinb(G97), .dout(n262));
  jnot g0191(.din(n262), .dout(n263));
  jor  g0192(.dina(n263), .dinb(n190), .dout(n264));
  jand g0193(.dina(n264), .dinb(n260), .dout(n265));
  jand g0194(.dina(n265), .dinb(n258), .dout(n266));
  jor  g0195(.dina(n266), .dinb(n248), .dout(n267));
  jand g0196(.dina(n246), .dinb(G200), .dout(n268));
  jor  g0197(.dina(n112), .dinb(G1), .dout(n269));
  jor  g0198(.dina(n269), .dinb(n114), .dout(n270));
  jand g0199(.dina(n270), .dinb(n179), .dout(n271));
  jand g0200(.dina(n262), .dinb(n271), .dout(n272));
  jor  g0201(.dina(n272), .dinb(n259), .dout(n273));
  jor  g0202(.dina(n273), .dinb(n257), .dout(n274));
  jand g0203(.dina(n234), .dinb(G190), .dout(n275));
  jor  g0204(.dina(n275), .dinb(n274), .dout(n276));
  jor  g0205(.dina(n276), .dinb(n268), .dout(n277));
  jand g0206(.dina(n277), .dinb(n267), .dout(n278));
  jand g0207(.dina(n278), .dinb(n219), .dout(n279));
  jand g0208(.dina(n152), .dinb(G264), .dout(n280));
  jand g0209(.dina(G303), .dinb(G33), .dout(n281));
  jand g0210(.dina(n155), .dinb(G257), .dout(n282));
  jor  g0211(.dina(n282), .dinb(n281), .dout(n283));
  jor  g0212(.dina(n283), .dinb(n280), .dout(n284));
  jand g0213(.dina(n284), .dinb(n151), .dout(n285));
  jand g0214(.dina(n243), .dinb(G270), .dout(n286));
  jor  g0215(.dina(n286), .dinb(n242), .dout(n287));
  jor  g0216(.dina(n287), .dinb(n285), .dout(n288));
  jand g0217(.dina(n288), .dinb(n146), .dout(n289));
  jand g0218(.dina(G97), .dinb(n148), .dout(n290));
  jor  g0219(.dina(n290), .dinb(G20), .dout(n291));
  jor  g0220(.dina(n291), .dinb(n221), .dout(n292));
  jand g0221(.dina(n105), .dinb(G20), .dout(n293));
  jnot g0222(.din(n293), .dout(n294));
  jand g0223(.dina(n294), .dinb(n189), .dout(n295));
  jand g0224(.dina(n295), .dinb(n292), .dout(n296));
  jnot g0225(.din(n296), .dout(n297));
  jand g0226(.dina(n185), .dinb(n105), .dout(n298));
  jnot g0227(.din(n298), .dout(n299));
  jor  g0228(.dina(n191), .dinb(n105), .dout(n300));
  jor  g0229(.dina(n300), .dinb(n190), .dout(n301));
  jand g0230(.dina(n301), .dinb(n299), .dout(n302));
  jand g0231(.dina(n302), .dinb(n297), .dout(n303));
  jor  g0232(.dina(n197), .dinb(n88), .dout(n304));
  jnot g0233(.din(n281), .dout(n305));
  jor  g0234(.dina(n199), .dinb(n91), .dout(n306));
  jand g0235(.dina(n306), .dinb(n305), .dout(n307));
  jand g0236(.dina(n307), .dinb(n304), .dout(n308));
  jor  g0237(.dina(n308), .dinb(n166), .dout(n309));
  jor  g0238(.dina(n231), .dinb(n106), .dout(n310));
  jand g0239(.dina(n310), .dinb(n229), .dout(n311));
  jand g0240(.dina(n311), .dinb(n309), .dout(n312));
  jand g0241(.dina(n312), .dinb(n196), .dout(n313));
  jor  g0242(.dina(n313), .dinb(n303), .dout(n314));
  jor  g0243(.dina(n314), .dinb(n289), .dout(n315));
  jand g0244(.dina(n288), .dinb(G200), .dout(n316));
  jnot g0245(.din(n300), .dout(n317));
  jand g0246(.dina(n317), .dinb(n271), .dout(n318));
  jor  g0247(.dina(n318), .dinb(n298), .dout(n319));
  jor  g0248(.dina(n319), .dinb(n296), .dout(n320));
  jand g0249(.dina(n312), .dinb(G190), .dout(n321));
  jor  g0250(.dina(n321), .dinb(n320), .dout(n322));
  jor  g0251(.dina(n322), .dinb(n316), .dout(n323));
  jand g0252(.dina(n323), .dinb(n315), .dout(n324));
  jor  g0253(.dina(n97), .dinb(G33), .dout(n325));
  jand g0254(.dina(n325), .dinb(n112), .dout(n326));
  jand g0255(.dina(n326), .dinb(n201), .dout(n327));
  jor  g0256(.dina(n327), .dinb(n179), .dout(n328));
  jor  g0257(.dina(n328), .dinb(G20), .dout(n329));
  jand g0258(.dina(n329), .dinb(G107), .dout(n330));
  jand g0259(.dina(n328), .dinb(n270), .dout(n331));
  jor  g0260(.dina(n331), .dinb(n330), .dout(n332));
  jand g0261(.dina(n261), .dinb(G107), .dout(n333));
  jand g0262(.dina(n333), .dinb(n271), .dout(n334));
  jnot g0263(.din(n334), .dout(n335));
  jand g0264(.dina(n335), .dinb(n332), .dout(n336));
  jor  g0265(.dina(n197), .dinb(n91), .dout(n337));
  jor  g0266(.dina(n199), .dinb(n98), .dout(n338));
  jand g0267(.dina(G294), .dinb(G33), .dout(n339));
  jnot g0268(.din(n339), .dout(n340));
  jand g0269(.dina(n340), .dinb(n338), .dout(n341));
  jand g0270(.dina(n341), .dinb(n337), .dout(n342));
  jor  g0271(.dina(n342), .dinb(n166), .dout(n343));
  jor  g0272(.dina(n231), .dinb(n88), .dout(n344));
  jand g0273(.dina(n344), .dinb(n229), .dout(n345));
  jand g0274(.dina(n345), .dinb(n343), .dout(n346));
  jand g0275(.dina(n346), .dinb(n196), .dout(n347));
  jand g0276(.dina(n152), .dinb(G257), .dout(n348));
  jand g0277(.dina(n155), .dinb(G250), .dout(n349));
  jor  g0278(.dina(n339), .dinb(n349), .dout(n350));
  jor  g0279(.dina(n350), .dinb(n348), .dout(n351));
  jand g0280(.dina(n351), .dinb(n151), .dout(n352));
  jand g0281(.dina(n243), .dinb(G264), .dout(n353));
  jor  g0282(.dina(n353), .dinb(n242), .dout(n354));
  jor  g0283(.dina(n354), .dinb(n352), .dout(n355));
  jand g0284(.dina(n355), .dinb(n146), .dout(n356));
  jor  g0285(.dina(n356), .dinb(n347), .dout(n357));
  jor  g0286(.dina(n357), .dinb(n336), .dout(n358));
  jand g0287(.dina(G87), .dinb(n148), .dout(n359));
  jor  g0288(.dina(n359), .dinb(G20), .dout(n360));
  jor  g0289(.dina(n360), .dinb(n157), .dout(n361));
  jand g0290(.dina(n361), .dinb(n189), .dout(n362));
  jand g0291(.dina(n362), .dinb(n112), .dout(n363));
  jor  g0292(.dina(n363), .dinb(n80), .dout(n364));
  jor  g0293(.dina(n362), .dinb(n185), .dout(n365));
  jand g0294(.dina(n365), .dinb(n364), .dout(n366));
  jor  g0295(.dina(n334), .dinb(n366), .dout(n367));
  jor  g0296(.dina(n355), .dinb(G190), .dout(n368));
  jor  g0297(.dina(n346), .dinb(G200), .dout(n369));
  jand g0298(.dina(n369), .dinb(n368), .dout(n370));
  jor  g0299(.dina(n370), .dinb(n367), .dout(n371));
  jand g0300(.dina(n371), .dinb(n358), .dout(n372));
  jand g0301(.dina(n372), .dinb(n324), .dout(n373));
  jand g0302(.dina(n373), .dinb(n279), .dout(n374));
  jand g0303(.dina(n155), .dinb(G232), .dout(n375));
  jand g0304(.dina(n152), .dinb(G238), .dout(n376));
  jor  g0305(.dina(n376), .dinb(n249), .dout(n377));
  jor  g0306(.dina(n377), .dinb(n375), .dout(n378));
  jand g0307(.dina(n378), .dinb(n151), .dout(n379));
  jand g0308(.dina(n161), .dinb(n149), .dout(n380));
  jor  g0309(.dina(n380), .dinb(G1), .dout(n381));
  jand g0310(.dina(n381), .dinb(n166), .dout(n382));
  jand g0311(.dina(n382), .dinb(G244), .dout(n383));
  jnot g0312(.din(n381), .dout(n384));
  jand g0313(.dina(n384), .dinb(n241), .dout(n385));
  jor  g0314(.dina(n385), .dinb(n383), .dout(n386));
  jor  g0315(.dina(n386), .dinb(n379), .dout(n387));
  jand g0316(.dina(n387), .dinb(n146), .dout(n388));
  jnot g0317(.din(n388), .dout(n389));
  jand g0318(.dina(G87), .dinb(G33), .dout(n390));
  jand g0319(.dina(G58), .dinb(n148), .dout(n391));
  jor  g0320(.dina(n391), .dinb(G20), .dout(n392));
  jor  g0321(.dina(n392), .dinb(n390), .dout(n393));
  jor  g0322(.dina(G77), .dinb(n112), .dout(n394));
  jand g0323(.dina(n394), .dinb(n189), .dout(n395));
  jand g0324(.dina(n395), .dinb(n393), .dout(n396));
  jand g0325(.dina(n185), .dinb(n72), .dout(n397));
  jand g0326(.dina(n269), .dinb(G77), .dout(n398));
  jand g0327(.dina(n398), .dinb(n271), .dout(n399));
  jor  g0328(.dina(n399), .dinb(n397), .dout(n400));
  jor  g0329(.dina(n400), .dinb(n396), .dout(n401));
  jor  g0330(.dina(n387), .dinb(G179), .dout(n402));
  jand g0331(.dina(n402), .dinb(n401), .dout(n403));
  jand g0332(.dina(n403), .dinb(n389), .dout(n404));
  jnot g0333(.din(n404), .dout(n405));
  jand g0334(.dina(n387), .dinb(G200), .dout(n406));
  jnot g0335(.din(G190), .dout(n407));
  jor  g0336(.dina(n387), .dinb(n407), .dout(n408));
  jnot g0337(.din(n408), .dout(n409));
  jor  g0338(.dina(n409), .dinb(n401), .dout(n410));
  jor  g0339(.dina(n410), .dinb(n406), .dout(n411));
  jand g0340(.dina(n411), .dinb(n405), .dout(n412));
  jand g0341(.dina(n155), .dinb(G226), .dout(n413));
  jand g0342(.dina(n152), .dinb(G232), .dout(n414));
  jor  g0343(.dina(n414), .dinb(n172), .dout(n415));
  jor  g0344(.dina(n415), .dinb(n413), .dout(n416));
  jand g0345(.dina(n416), .dinb(n151), .dout(n417));
  jand g0346(.dina(n382), .dinb(G238), .dout(n418));
  jor  g0347(.dina(n418), .dinb(n385), .dout(n419));
  jor  g0348(.dina(n419), .dinb(n417), .dout(n420));
  jand g0349(.dina(n420), .dinb(n146), .dout(n421));
  jnot g0350(.din(n421), .dout(n422));
  jand g0351(.dina(n269), .dinb(G68), .dout(n423));
  jand g0352(.dina(n423), .dinb(n271), .dout(n424));
  jand g0353(.dina(n148), .dinb(n114), .dout(n425));
  jnot g0354(.din(n425), .dout(n426));
  jand g0355(.dina(n426), .dinb(n85), .dout(n427));
  jor  g0356(.dina(n427), .dinb(n185), .dout(n428));
  jand g0357(.dina(n428), .dinb(n75), .dout(n429));
  jand g0358(.dina(G77), .dinb(G33), .dout(n430));
  jand g0359(.dina(G50), .dinb(n148), .dout(n431));
  jor  g0360(.dina(n431), .dinb(n430), .dout(n432));
  jand g0361(.dina(n432), .dinb(n112), .dout(n433));
  jand g0362(.dina(n433), .dinb(n189), .dout(n434));
  jor  g0363(.dina(n434), .dinb(n429), .dout(n435));
  jor  g0364(.dina(n435), .dinb(n424), .dout(n436));
  jor  g0365(.dina(n420), .dinb(G179), .dout(n437));
  jand g0366(.dina(n437), .dinb(n436), .dout(n438));
  jand g0367(.dina(n438), .dinb(n422), .dout(n439));
  jnot g0368(.din(n439), .dout(n440));
  jand g0369(.dina(n420), .dinb(G200), .dout(n441));
  jor  g0370(.dina(n420), .dinb(n407), .dout(n442));
  jnot g0371(.din(n442), .dout(n443));
  jor  g0372(.dina(n443), .dinb(n436), .dout(n444));
  jor  g0373(.dina(n444), .dinb(n441), .dout(n445));
  jand g0374(.dina(n445), .dinb(n440), .dout(n446));
  jand g0375(.dina(n446), .dinb(n412), .dout(n447));
  jand g0376(.dina(n152), .dinb(G223), .dout(n448));
  jand g0377(.dina(n155), .dinb(G222), .dout(n449));
  jor  g0378(.dina(n449), .dinb(n430), .dout(n450));
  jor  g0379(.dina(n450), .dinb(n448), .dout(n451));
  jand g0380(.dina(n451), .dinb(n151), .dout(n452));
  jand g0381(.dina(n382), .dinb(G226), .dout(n453));
  jor  g0382(.dina(n453), .dinb(n385), .dout(n454));
  jor  g0383(.dina(n454), .dinb(n452), .dout(n455));
  jand g0384(.dina(n455), .dinb(n146), .dout(n456));
  jand g0385(.dina(n269), .dinb(G50), .dout(n457));
  jnot g0386(.din(n457), .dout(n458));
  jor  g0387(.dina(n458), .dinb(n190), .dout(n459));
  jor  g0388(.dina(n77), .dinb(n112), .dout(n460));
  jnot g0389(.din(G150), .dout(n461));
  jand g0390(.dina(n148), .dinb(n112), .dout(n462));
  jnot g0391(.din(n462), .dout(n463));
  jor  g0392(.dina(n463), .dinb(n461), .dout(n464));
  jand g0393(.dina(G33), .dinb(n112), .dout(n465));
  jand g0394(.dina(n465), .dinb(G58), .dout(n466));
  jnot g0395(.din(n466), .dout(n467));
  jand g0396(.dina(n467), .dinb(n464), .dout(n468));
  jand g0397(.dina(n468), .dinb(n460), .dout(n469));
  jor  g0398(.dina(n469), .dinb(n179), .dout(n470));
  jand g0399(.dina(n185), .dinb(n73), .dout(n471));
  jnot g0400(.din(n471), .dout(n472));
  jand g0401(.dina(n472), .dinb(n470), .dout(n473));
  jand g0402(.dina(n473), .dinb(n459), .dout(n474));
  jnot g0403(.din(n455), .dout(n475));
  jand g0404(.dina(n475), .dinb(n196), .dout(n476));
  jor  g0405(.dina(n476), .dinb(n474), .dout(n477));
  jor  g0406(.dina(n477), .dinb(n456), .dout(n478));
  jnot g0407(.din(n474), .dout(n479));
  jand g0408(.dina(n475), .dinb(G190), .dout(n480));
  jand g0409(.dina(n455), .dinb(G200), .dout(n481));
  jor  g0410(.dina(n481), .dinb(n480), .dout(n482));
  jor  g0411(.dina(n482), .dinb(n479), .dout(n483));
  jand g0412(.dina(n483), .dinb(n478), .dout(n484));
  jand g0413(.dina(n152), .dinb(G226), .dout(n485));
  jand g0414(.dina(n155), .dinb(G223), .dout(n486));
  jor  g0415(.dina(n486), .dinb(n390), .dout(n487));
  jor  g0416(.dina(n487), .dinb(n485), .dout(n488));
  jand g0417(.dina(n488), .dinb(n151), .dout(n489));
  jand g0418(.dina(n382), .dinb(G232), .dout(n490));
  jor  g0419(.dina(n490), .dinb(n385), .dout(n491));
  jor  g0420(.dina(n491), .dinb(n489), .dout(n492));
  jand g0421(.dina(n492), .dinb(n146), .dout(n493));
  jand g0422(.dina(n269), .dinb(G58), .dout(n494));
  jnot g0423(.din(n494), .dout(n495));
  jor  g0424(.dina(n495), .dinb(n190), .dout(n496));
  jor  g0425(.dina(n137), .dinb(n112), .dout(n497));
  jand g0426(.dina(n462), .dinb(G159), .dout(n498));
  jand g0427(.dina(n465), .dinb(G68), .dout(n499));
  jor  g0428(.dina(n499), .dinb(n498), .dout(n500));
  jnot g0429(.din(n500), .dout(n501));
  jand g0430(.dina(n501), .dinb(n497), .dout(n502));
  jor  g0431(.dina(n502), .dinb(n179), .dout(n503));
  jand g0432(.dina(n185), .dinb(n74), .dout(n504));
  jnot g0433(.din(n504), .dout(n505));
  jand g0434(.dina(n505), .dinb(n503), .dout(n506));
  jand g0435(.dina(n506), .dinb(n496), .dout(n507));
  jnot g0436(.din(n492), .dout(n508));
  jand g0437(.dina(n508), .dinb(n196), .dout(n509));
  jor  g0438(.dina(n509), .dinb(n507), .dout(n510));
  jor  g0439(.dina(n510), .dinb(n493), .dout(n511));
  jnot g0440(.din(n507), .dout(n512));
  jand g0441(.dina(n508), .dinb(G190), .dout(n513));
  jand g0442(.dina(n492), .dinb(G200), .dout(n514));
  jor  g0443(.dina(n514), .dinb(n513), .dout(n515));
  jor  g0444(.dina(n515), .dinb(n512), .dout(n516));
  jand g0445(.dina(n516), .dinb(n511), .dout(n517));
  jand g0446(.dina(n517), .dinb(n484), .dout(n518));
  jand g0447(.dina(n518), .dinb(n447), .dout(n519));
  jand g0448(.dina(n519), .dinb(n374), .dout(G372));
  jor  g0449(.dina(n355), .dinb(G179), .dout(n521));
  jor  g0450(.dina(n346), .dinb(G169), .dout(n522));
  jand g0451(.dina(n522), .dinb(n521), .dout(n523));
  jand g0452(.dina(n523), .dinb(n367), .dout(n524));
  jor  g0453(.dina(n312), .dinb(G169), .dout(n525));
  jor  g0454(.dina(n288), .dinb(G179), .dout(n526));
  jand g0455(.dina(n526), .dinb(n320), .dout(n527));
  jand g0456(.dina(n527), .dinb(n525), .dout(n528));
  jand g0457(.dina(n371), .dinb(n528), .dout(n529));
  jor  g0458(.dina(n529), .dinb(n524), .dout(n530));
  jand g0459(.dina(n530), .dinb(n279), .dout(n531));
  jnot g0460(.din(n213), .dout(n532));
  jand g0461(.dina(n246), .dinb(G169), .dout(n533));
  jand g0462(.dina(n234), .dinb(G179), .dout(n534));
  jor  g0463(.dina(n534), .dinb(n533), .dout(n535));
  jand g0464(.dina(n274), .dinb(n535), .dout(n536));
  jand g0465(.dina(n536), .dinb(n218), .dout(n537));
  jor  g0466(.dina(n537), .dinb(n532), .dout(n538));
  jor  g0467(.dina(n538), .dinb(n531), .dout(n539));
  jand g0468(.dina(n539), .dinb(n519), .dout(n540));
  jnot g0469(.din(n478), .dout(n541));
  jnot g0470(.din(n511), .dout(n542));
  jor  g0471(.dina(n439), .dinb(n404), .dout(n543));
  jand g0472(.dina(n543), .dinb(n445), .dout(n544));
  jor  g0473(.dina(n544), .dinb(n542), .dout(n545));
  jand g0474(.dina(n545), .dinb(n516), .dout(n546));
  jor  g0475(.dina(n546), .dinb(n541), .dout(n547));
  jand g0476(.dina(n547), .dinb(n483), .dout(n548));
  jor  g0477(.dina(n548), .dinb(n540), .dout(G369));
  jand g0478(.dina(n112), .dinb(G13), .dout(n550));
  jand g0479(.dina(G213), .dinb(n113), .dout(n551));
  jand g0480(.dina(n551), .dinb(n550), .dout(n552));
  jand g0481(.dina(n552), .dinb(G343), .dout(n553));
  jnot g0482(.din(n553), .dout(n554));
  jand g0483(.dina(n554), .dinb(n524), .dout(n555));
  jand g0484(.dina(n554), .dinb(n528), .dout(n556));
  jand g0485(.dina(n553), .dinb(n367), .dout(n557));
  jnot g0486(.din(n557), .dout(n558));
  jand g0487(.dina(n558), .dinb(n372), .dout(n559));
  jand g0488(.dina(n557), .dinb(n523), .dout(n560));
  jor  g0489(.dina(n560), .dinb(n559), .dout(n561));
  jand g0490(.dina(n561), .dinb(n556), .dout(n562));
  jor  g0491(.dina(n562), .dinb(n555), .dout(n563));
  jnot g0492(.din(n561), .dout(n564));
  jnot g0493(.din(G330), .dout(n565));
  jnot g0494(.din(n324), .dout(n566));
  jor  g0495(.dina(n554), .dinb(n303), .dout(n567));
  jnot g0496(.din(n567), .dout(n568));
  jor  g0497(.dina(n568), .dinb(n566), .dout(n569));
  jor  g0498(.dina(n567), .dinb(n315), .dout(n570));
  jand g0499(.dina(n570), .dinb(n569), .dout(n571));
  jor  g0500(.dina(n571), .dinb(n565), .dout(n572));
  jor  g0501(.dina(n572), .dinb(n564), .dout(n573));
  jnot g0502(.din(n573), .dout(n574));
  jor  g0503(.dina(n574), .dinb(n563), .dout(G399));
  jand g0504(.dina(n554), .dinb(n539), .dout(n576));
  jor  g0505(.dina(n553), .dinb(n374), .dout(n577));
  jand g0506(.dina(n346), .dinb(n210), .dout(n578));
  jand g0507(.dina(n578), .dinb(n312), .dout(n579));
  jand g0508(.dina(n579), .dinb(n534), .dout(n580));
  jand g0509(.dina(n288), .dinb(n196), .dout(n581));
  jand g0510(.dina(n355), .dinb(n246), .dout(n582));
  jand g0511(.dina(n582), .dinb(n170), .dout(n583));
  jand g0512(.dina(n583), .dinb(n581), .dout(n584));
  jor  g0513(.dina(n584), .dinb(n554), .dout(n585));
  jor  g0514(.dina(n585), .dinb(n580), .dout(n586));
  jand g0515(.dina(n586), .dinb(G330), .dout(n587));
  jand g0516(.dina(n587), .dinb(n577), .dout(n588));
  jor  g0517(.dina(n588), .dinb(n576), .dout(n589));
  jand g0518(.dina(n589), .dinb(n113), .dout(n590));
  jand g0519(.dina(n122), .dinb(n149), .dout(n591));
  jnot g0520(.din(n591), .dout(n592));
  jand g0521(.dina(n180), .dinb(n105), .dout(n593));
  jand g0522(.dina(n593), .dinb(G1), .dout(n594));
  jand g0523(.dina(n594), .dinb(n592), .dout(n595));
  jand g0524(.dina(n591), .dinb(n118), .dout(n596));
  jor  g0525(.dina(n596), .dinb(n595), .dout(n597));
  jor  g0526(.dina(n597), .dinb(n590), .dout(G364));
  jand g0527(.dina(n571), .dinb(n565), .dout(n599));
  jnot g0528(.din(n599), .dout(n600));
  jand g0529(.dina(n550), .dinb(G45), .dout(n601));
  jor  g0530(.dina(n601), .dinb(n113), .dout(n602));
  jnot g0531(.din(n602), .dout(n603));
  jand g0532(.dina(n603), .dinb(n592), .dout(n604));
  jnot g0533(.din(n604), .dout(n605));
  jand g0534(.dina(n605), .dinb(n572), .dout(n606));
  jand g0535(.dina(n606), .dinb(n600), .dout(n607));
  jand g0536(.dina(n462), .dinb(n114), .dout(n608));
  jand g0537(.dina(n608), .dinb(n571), .dout(n609));
  jnot g0538(.din(n609), .dout(n610));
  jand g0539(.dina(n146), .dinb(G20), .dout(n611));
  jor  g0540(.dina(n611), .dinb(n115), .dout(n612));
  jand g0541(.dina(G179), .dinb(G20), .dout(n613));
  jnot g0542(.din(n613), .dout(n614));
  jand g0543(.dina(G200), .dinb(G20), .dout(n615));
  jand g0544(.dina(n615), .dinb(n614), .dout(n616));
  jand g0545(.dina(n616), .dinb(G190), .dout(n617));
  jand g0546(.dina(n617), .dinb(G303), .dout(n618));
  jand g0547(.dina(n407), .dinb(G20), .dout(n619));
  jnot g0548(.din(n619), .dout(n620));
  jor  g0549(.dina(n615), .dinb(n613), .dout(n621));
  jnot g0550(.din(n621), .dout(n622));
  jand g0551(.dina(n622), .dinb(n620), .dout(n623));
  jand g0552(.dina(n623), .dinb(G294), .dout(n624));
  jnot g0553(.din(G200), .dout(n625));
  jand g0554(.dina(n613), .dinb(n625), .dout(n626));
  jand g0555(.dina(n626), .dinb(G190), .dout(n627));
  jand g0556(.dina(n627), .dinb(G322), .dout(n628));
  jor  g0557(.dina(n628), .dinb(n624), .dout(n629));
  jor  g0558(.dina(n629), .dinb(n618), .dout(n630));
  jand g0559(.dina(n622), .dinb(n619), .dout(n631));
  jand g0560(.dina(n631), .dinb(G329), .dout(n632));
  jor  g0561(.dina(n632), .dinb(n148), .dout(n633));
  jand g0562(.dina(n616), .dinb(n407), .dout(n634));
  jand g0563(.dina(n634), .dinb(G283), .dout(n635));
  jand g0564(.dina(n626), .dinb(n407), .dout(n636));
  jand g0565(.dina(n636), .dinb(G311), .dout(n637));
  jor  g0566(.dina(n637), .dinb(n635), .dout(n638));
  jand g0567(.dina(n613), .dinb(G200), .dout(n639));
  jand g0568(.dina(n639), .dinb(G190), .dout(n640));
  jand g0569(.dina(n640), .dinb(G326), .dout(n641));
  jand g0570(.dina(n639), .dinb(n407), .dout(n642));
  jand g0571(.dina(n642), .dinb(G317), .dout(n643));
  jor  g0572(.dina(n643), .dinb(n641), .dout(n644));
  jor  g0573(.dina(n644), .dinb(n638), .dout(n645));
  jor  g0574(.dina(n645), .dinb(n633), .dout(n646));
  jor  g0575(.dina(n646), .dinb(n630), .dout(n647));
  jand g0576(.dina(n631), .dinb(G159), .dout(n648));
  jand g0577(.dina(n640), .dinb(G50), .dout(n649));
  jand g0578(.dina(n642), .dinb(G68), .dout(n650));
  jor  g0579(.dina(n650), .dinb(n649), .dout(n651));
  jor  g0580(.dina(n651), .dinb(n648), .dout(n652));
  jnot g0581(.din(n652), .dout(n653));
  jand g0582(.dina(n617), .dinb(G87), .dout(n654));
  jnot g0583(.din(n654), .dout(n655));
  jand g0584(.dina(n655), .dinb(n148), .dout(n656));
  jand g0585(.dina(n634), .dinb(G107), .dout(n657));
  jand g0586(.dina(n636), .dinb(G77), .dout(n658));
  jor  g0587(.dina(n658), .dinb(n657), .dout(n659));
  jand g0588(.dina(n627), .dinb(G58), .dout(n660));
  jand g0589(.dina(n623), .dinb(G97), .dout(n661));
  jor  g0590(.dina(n661), .dinb(n660), .dout(n662));
  jor  g0591(.dina(n662), .dinb(n659), .dout(n663));
  jnot g0592(.din(n663), .dout(n664));
  jand g0593(.dina(n664), .dinb(n656), .dout(n665));
  jand g0594(.dina(n665), .dinb(n653), .dout(n666));
  jnot g0595(.din(n666), .dout(n667));
  jand g0596(.dina(n667), .dinb(n647), .dout(n668));
  jor  g0597(.dina(n668), .dinb(n612), .dout(n669));
  jnot g0598(.din(n608), .dout(n670));
  jand g0599(.dina(n612), .dinb(n670), .dout(n671));
  jnot g0600(.din(n671), .dout(n672));
  jand g0601(.dina(n140), .dinb(G45), .dout(n673));
  jand g0602(.dina(n118), .dinb(n161), .dout(n674));
  jand g0603(.dina(n122), .dinb(G33), .dout(n675));
  jnot g0604(.din(n675), .dout(n676));
  jor  g0605(.dina(n676), .dinb(n674), .dout(n677));
  jor  g0606(.dina(n677), .dinb(n673), .dout(n678));
  jand g0607(.dina(n123), .dinb(n105), .dout(n679));
  jand g0608(.dina(n122), .dinb(n148), .dout(n680));
  jand g0609(.dina(n680), .dinb(G355), .dout(n681));
  jor  g0610(.dina(n681), .dinb(n679), .dout(n682));
  jnot g0611(.din(n682), .dout(n683));
  jand g0612(.dina(n683), .dinb(n678), .dout(n684));
  jor  g0613(.dina(n684), .dinb(n672), .dout(n685));
  jand g0614(.dina(n685), .dinb(n604), .dout(n686));
  jand g0615(.dina(n686), .dinb(n669), .dout(n687));
  jand g0616(.dina(n687), .dinb(n610), .dout(n688));
  jor  g0617(.dina(n688), .dinb(n607), .dout(G396));
  jnot g0618(.din(n588), .dout(n690));
  jnot g0619(.din(n401), .dout(n691));
  jor  g0620(.dina(n554), .dinb(n691), .dout(n692));
  jand g0621(.dina(n692), .dinb(n412), .dout(n693));
  jor  g0622(.dina(n692), .dinb(n405), .dout(n694));
  jnot g0623(.din(n694), .dout(n695));
  jor  g0624(.dina(n695), .dinb(n693), .dout(n696));
  jxor g0625(.dina(n696), .dinb(n576), .dout(n697));
  jnot g0626(.din(n697), .dout(n698));
  jand g0627(.dina(n698), .dinb(n690), .dout(n699));
  jor  g0628(.dina(n991), .dinb(n604), .dout(n701));
  jor  g0629(.dina(n701), .dinb(n699), .dout(n702));
  jnot g0630(.din(n696), .dout(n703));
  jand g0631(.dina(n703), .dinb(n425), .dout(n704));
  jnot g0632(.din(n704), .dout(n705));
  jand g0633(.dina(n631), .dinb(G132), .dout(n706));
  jand g0634(.dina(n623), .dinb(G58), .dout(n707));
  jand g0635(.dina(n642), .dinb(G150), .dout(n708));
  jor  g0636(.dina(n708), .dinb(n707), .dout(n709));
  jor  g0637(.dina(n709), .dinb(n706), .dout(n710));
  jand g0638(.dina(n617), .dinb(G50), .dout(n711));
  jor  g0639(.dina(n711), .dinb(G33), .dout(n712));
  jand g0640(.dina(n636), .dinb(G159), .dout(n713));
  jand g0641(.dina(n627), .dinb(G143), .dout(n714));
  jor  g0642(.dina(n714), .dinb(n713), .dout(n715));
  jand g0643(.dina(n640), .dinb(G137), .dout(n716));
  jand g0644(.dina(n634), .dinb(G68), .dout(n717));
  jor  g0645(.dina(n717), .dinb(n716), .dout(n718));
  jor  g0646(.dina(n718), .dinb(n715), .dout(n719));
  jor  g0647(.dina(n719), .dinb(n712), .dout(n720));
  jor  g0648(.dina(n720), .dinb(n710), .dout(n721));
  jand g0649(.dina(n631), .dinb(G311), .dout(n722));
  jand g0650(.dina(n617), .dinb(G107), .dout(n723));
  jand g0651(.dina(n642), .dinb(G283), .dout(n724));
  jor  g0652(.dina(n724), .dinb(n723), .dout(n725));
  jor  g0653(.dina(n725), .dinb(n722), .dout(n726));
  jnot g0654(.din(n726), .dout(n727));
  jand g0655(.dina(n634), .dinb(G87), .dout(n728));
  jnot g0656(.din(n728), .dout(n729));
  jand g0657(.dina(n729), .dinb(G33), .dout(n730));
  jand g0658(.dina(n636), .dinb(G116), .dout(n731));
  jand g0659(.dina(n627), .dinb(G294), .dout(n732));
  jor  g0660(.dina(n732), .dinb(n731), .dout(n733));
  jand g0661(.dina(n640), .dinb(G303), .dout(n734));
  jor  g0662(.dina(n734), .dinb(n661), .dout(n735));
  jor  g0663(.dina(n735), .dinb(n733), .dout(n736));
  jnot g0664(.din(n736), .dout(n737));
  jand g0665(.dina(n737), .dinb(n730), .dout(n738));
  jand g0666(.dina(n738), .dinb(n727), .dout(n739));
  jnot g0667(.din(n739), .dout(n740));
  jand g0668(.dina(n740), .dinb(n721), .dout(n741));
  jor  g0669(.dina(n741), .dinb(n612), .dout(n742));
  jand g0670(.dina(n612), .dinb(n426), .dout(n743));
  jand g0671(.dina(n743), .dinb(n72), .dout(n744));
  jor  g0672(.dina(n744), .dinb(n605), .dout(n745));
  jnot g0673(.din(n745), .dout(n746));
  jand g0674(.dina(n746), .dinb(n742), .dout(n747));
  jand g0675(.dina(n747), .dinb(n705), .dout(n748));
  jnot g0676(.din(n748), .dout(n749));
  jand g0677(.dina(n749), .dinb(n702), .dout(n750));
  jnot g0678(.din(n750), .dout(G384));
  jnot g0679(.din(n552), .dout(n752));
  jand g0680(.dina(n752), .dinb(n542), .dout(n753));
  jand g0681(.dina(n552), .dinb(n512), .dout(n754));
  jnot g0682(.din(n754), .dout(n755));
  jand g0683(.dina(n755), .dinb(n517), .dout(n756));
  jand g0684(.dina(n754), .dinb(n542), .dout(n757));
  jor  g0685(.dina(n757), .dinb(n756), .dout(n758));
  jand g0686(.dina(n696), .dinb(n576), .dout(n759));
  jand g0687(.dina(n553), .dinb(n436), .dout(n760));
  jnot g0688(.din(n760), .dout(n761));
  jand g0689(.dina(n761), .dinb(n446), .dout(n762));
  jand g0690(.dina(n760), .dinb(n439), .dout(n763));
  jor  g0691(.dina(n763), .dinb(n762), .dout(n764));
  jand g0692(.dina(n764), .dinb(n759), .dout(n765));
  jor  g0693(.dina(n764), .dinb(n439), .dout(n766));
  jand g0694(.dina(n554), .dinb(n543), .dout(n767));
  jand g0695(.dina(n767), .dinb(n766), .dout(n768));
  jor  g0696(.dina(n768), .dinb(n765), .dout(n769));
  jand g0697(.dina(n769), .dinb(n758), .dout(n770));
  jor  g0698(.dina(n770), .dinb(n753), .dout(n771));
  jnot g0699(.din(n771), .dout(n772));
  jand g0700(.dina(n576), .dinb(n519), .dout(n773));
  jor  g0701(.dina(n773), .dinb(n548), .dout(n774));
  jand g0702(.dina(n764), .dinb(n696), .dout(n775));
  jand g0703(.dina(n775), .dinb(n758), .dout(n776));
  jxor g0704(.dina(n776), .dinb(n519), .dout(n777));
  jand g0705(.dina(n777), .dinb(n588), .dout(n778));
  jxor g0706(.dina(n778), .dinb(n774), .dout(n779));
  jnot g0707(.din(n779), .dout(n780));
  jor  g0708(.dina(n780), .dinb(n772), .dout(n781));
  jor  g0709(.dina(n779), .dinb(n771), .dout(n782));
  jnot g0710(.din(n121), .dout(n783));
  jand g0711(.dina(n783), .dinb(n116), .dout(n784));
  jand g0712(.dina(n784), .dinb(n782), .dout(n785));
  jand g0713(.dina(n785), .dinb(n781), .dout(n786));
  jand g0714(.dina(G77), .dinb(G50), .dout(n787));
  jand g0715(.dina(n787), .dinb(n137), .dout(n788));
  jand g0716(.dina(G68), .dinb(n73), .dout(n789));
  jor  g0717(.dina(n789), .dinb(n788), .dout(n790));
  jand g0718(.dina(n790), .dinb(n121), .dout(n791));
  jnot g0719(.din(n255), .dout(n792));
  jand g0720(.dina(n147), .dinb(G116), .dout(n793));
  jand g0721(.dina(n793), .dinb(n792), .dout(n794));
  jor  g0722(.dina(n794), .dinb(n791), .dout(n795));
  jor  g0723(.dina(n795), .dinb(n786), .dout(G367));
  jand g0724(.dina(n553), .dinb(n214), .dout(n797));
  jnot g0725(.din(n797), .dout(n798));
  jand g0726(.dina(n798), .dinb(n219), .dout(n799));
  jand g0727(.dina(n797), .dinb(n532), .dout(n800));
  jor  g0728(.dina(n800), .dinb(n799), .dout(n801));
  jnot g0729(.din(n801), .dout(n802));
  jand g0730(.dina(n802), .dinb(n608), .dout(n803));
  jnot g0731(.din(n803), .dout(n804));
  jand g0732(.dina(n631), .dinb(G317), .dout(n805));
  jand g0733(.dina(n623), .dinb(G107), .dout(n806));
  jand g0734(.dina(n642), .dinb(G294), .dout(n807));
  jor  g0735(.dina(n807), .dinb(n806), .dout(n808));
  jor  g0736(.dina(n808), .dinb(n805), .dout(n809));
  jand g0737(.dina(n617), .dinb(G116), .dout(n810));
  jor  g0738(.dina(n810), .dinb(n148), .dout(n811));
  jand g0739(.dina(n636), .dinb(G283), .dout(n812));
  jand g0740(.dina(n627), .dinb(G303), .dout(n813));
  jor  g0741(.dina(n813), .dinb(n812), .dout(n814));
  jand g0742(.dina(n640), .dinb(G311), .dout(n815));
  jand g0743(.dina(n634), .dinb(G97), .dout(n816));
  jor  g0744(.dina(n816), .dinb(n815), .dout(n817));
  jor  g0745(.dina(n817), .dinb(n814), .dout(n818));
  jor  g0746(.dina(n818), .dinb(n811), .dout(n819));
  jor  g0747(.dina(n819), .dinb(n809), .dout(n820));
  jand g0748(.dina(n631), .dinb(G137), .dout(n821));
  jnot g0749(.din(n821), .dout(n822));
  jand g0750(.dina(n623), .dinb(G68), .dout(n823));
  jnot g0751(.din(n823), .dout(n824));
  jand g0752(.dina(n634), .dinb(G77), .dout(n825));
  jnot g0753(.din(n825), .dout(n826));
  jand g0754(.dina(n826), .dinb(n824), .dout(n827));
  jand g0755(.dina(n827), .dinb(n822), .dout(n828));
  jand g0756(.dina(n642), .dinb(G159), .dout(n829));
  jor  g0757(.dina(n829), .dinb(G33), .dout(n830));
  jand g0758(.dina(n640), .dinb(G143), .dout(n831));
  jand g0759(.dina(n627), .dinb(G150), .dout(n832));
  jor  g0760(.dina(n832), .dinb(n831), .dout(n833));
  jand g0761(.dina(n636), .dinb(G50), .dout(n834));
  jand g0762(.dina(n617), .dinb(G58), .dout(n835));
  jor  g0763(.dina(n835), .dinb(n834), .dout(n836));
  jor  g0764(.dina(n836), .dinb(n833), .dout(n837));
  jor  g0765(.dina(n837), .dinb(n830), .dout(n838));
  jnot g0766(.din(n838), .dout(n839));
  jand g0767(.dina(n839), .dinb(n828), .dout(n840));
  jnot g0768(.din(n840), .dout(n841));
  jand g0769(.dina(n841), .dinb(n820), .dout(n842));
  jor  g0770(.dina(n842), .dinb(n612), .dout(n843));
  jand g0771(.dina(n675), .dinb(n131), .dout(n844));
  jand g0772(.dina(n123), .dinb(G87), .dout(n845));
  jor  g0773(.dina(n845), .dinb(n672), .dout(n846));
  jor  g0774(.dina(n846), .dinb(n844), .dout(n847));
  jand g0775(.dina(n847), .dinb(n604), .dout(n848));
  jand g0776(.dina(n848), .dinb(n843), .dout(n849));
  jand g0777(.dina(n849), .dinb(n804), .dout(n850));
  jnot g0778(.din(n589), .dout(n851));
  jxor g0779(.dina(n561), .dinb(n556), .dout(n852));
  jxor g0780(.dina(n852), .dinb(n572), .dout(n853));
  jnot g0781(.din(n853), .dout(n854));
  jand g0782(.dina(n854), .dinb(n851), .dout(n855));
  jnot g0783(.din(n278), .dout(n856));
  jand g0784(.dina(n553), .dinb(n274), .dout(n857));
  jor  g0785(.dina(n857), .dinb(n856), .dout(n858));
  jand g0786(.dina(n553), .dinb(n536), .dout(n859));
  jnot g0787(.din(n859), .dout(n860));
  jand g0788(.dina(n860), .dinb(n858), .dout(n861));
  jxor g0789(.dina(n861), .dinb(n573), .dout(n862));
  jxor g0790(.dina(n862), .dinb(n563), .dout(n863));
  jand g0791(.dina(n863), .dinb(n855), .dout(n864));
  jor  g0792(.dina(n864), .dinb(n589), .dout(n865));
  jand g0793(.dina(n865), .dinb(n591), .dout(n866));
  jor  g0794(.dina(n866), .dinb(n602), .dout(n867));
  jand g0795(.dina(n554), .dinb(n536), .dout(n868));
  jnot g0796(.din(n861), .dout(n869));
  jand g0797(.dina(n869), .dinb(n563), .dout(n870));
  jor  g0798(.dina(n870), .dinb(n868), .dout(n871));
  jor  g0799(.dina(n861), .dinb(n573), .dout(n872));
  jxor g0800(.dina(n872), .dinb(n801), .dout(n873));
  jxor g0801(.dina(n873), .dinb(n871), .dout(n874));
  jnot g0802(.din(n874), .dout(n875));
  jand g0803(.dina(n875), .dinb(n867), .dout(n876));
  jor  g0804(.dina(n876), .dinb(n850), .dout(G387));
  jand g0805(.dina(n853), .dinb(n589), .dout(n878));
  jor  g0806(.dina(n855), .dinb(n592), .dout(n879));
  jor  g0807(.dina(n879), .dinb(n878), .dout(n880));
  jor  g0808(.dina(n853), .dinb(n603), .dout(n881));
  jand g0809(.dina(n608), .dinb(n564), .dout(n882));
  jand g0810(.dina(n631), .dinb(G326), .dout(n883));
  jand g0811(.dina(n623), .dinb(G283), .dout(n884));
  jand g0812(.dina(n627), .dinb(G317), .dout(n885));
  jor  g0813(.dina(n885), .dinb(n884), .dout(n886));
  jor  g0814(.dina(n886), .dinb(n883), .dout(n887));
  jand g0815(.dina(n617), .dinb(G294), .dout(n888));
  jor  g0816(.dina(n888), .dinb(n148), .dout(n889));
  jand g0817(.dina(n634), .dinb(G116), .dout(n890));
  jand g0818(.dina(n636), .dinb(G303), .dout(n891));
  jor  g0819(.dina(n891), .dinb(n890), .dout(n892));
  jand g0820(.dina(n640), .dinb(G322), .dout(n893));
  jand g0821(.dina(n642), .dinb(G311), .dout(n894));
  jor  g0822(.dina(n894), .dinb(n893), .dout(n895));
  jor  g0823(.dina(n895), .dinb(n892), .dout(n896));
  jor  g0824(.dina(n896), .dinb(n889), .dout(n897));
  jor  g0825(.dina(n897), .dinb(n887), .dout(n898));
  jand g0826(.dina(n623), .dinb(G87), .dout(n899));
  jand g0827(.dina(n642), .dinb(G58), .dout(n900));
  jor  g0828(.dina(n900), .dinb(n816), .dout(n901));
  jor  g0829(.dina(n901), .dinb(n899), .dout(n902));
  jand g0830(.dina(n631), .dinb(G150), .dout(n903));
  jor  g0831(.dina(n903), .dinb(G33), .dout(n904));
  jand g0832(.dina(n640), .dinb(G159), .dout(n905));
  jand g0833(.dina(n636), .dinb(G68), .dout(n906));
  jor  g0834(.dina(n906), .dinb(n905), .dout(n907));
  jand g0835(.dina(n627), .dinb(G50), .dout(n908));
  jand g0836(.dina(n617), .dinb(G77), .dout(n909));
  jor  g0837(.dina(n909), .dinb(n908), .dout(n910));
  jor  g0838(.dina(n910), .dinb(n907), .dout(n911));
  jor  g0839(.dina(n911), .dinb(n904), .dout(n912));
  jor  g0840(.dina(n912), .dinb(n902), .dout(n913));
  jand g0841(.dina(n913), .dinb(n898), .dout(n914));
  jor  g0842(.dina(n914), .dinb(n612), .dout(n915));
  jand g0843(.dina(n135), .dinb(G45), .dout(n916));
  jand g0844(.dina(G77), .dinb(G68), .dout(n917));
  jnot g0845(.din(n917), .dout(n918));
  jand g0846(.dina(G58), .dinb(n161), .dout(n919));
  jand g0847(.dina(n919), .dinb(n73), .dout(n920));
  jand g0848(.dina(n920), .dinb(n918), .dout(n921));
  jand g0849(.dina(n921), .dinb(n593), .dout(n922));
  jor  g0850(.dina(n922), .dinb(n676), .dout(n923));
  jor  g0851(.dina(n923), .dinb(n916), .dout(n924));
  jand g0852(.dina(n123), .dinb(n80), .dout(n925));
  jnot g0853(.din(n593), .dout(n926));
  jand g0854(.dina(n680), .dinb(n926), .dout(n927));
  jor  g0855(.dina(n927), .dinb(n925), .dout(n928));
  jnot g0856(.din(n928), .dout(n929));
  jand g0857(.dina(n929), .dinb(n924), .dout(n930));
  jor  g0858(.dina(n930), .dinb(n672), .dout(n931));
  jand g0859(.dina(n931), .dinb(n604), .dout(n932));
  jand g0860(.dina(n932), .dinb(n915), .dout(n933));
  jnot g0861(.din(n933), .dout(n934));
  jor  g0862(.dina(n934), .dinb(n882), .dout(n935));
  jand g0863(.dina(n935), .dinb(n881), .dout(n936));
  jand g0864(.dina(n936), .dinb(n880), .dout(n937));
  jnot g0865(.din(n937), .dout(G393));
  jnot g0866(.din(n855), .dout(n939));
  jnot g0867(.din(n863), .dout(n940));
  jand g0868(.dina(n940), .dinb(n939), .dout(n941));
  jor  g0869(.dina(n864), .dinb(n592), .dout(n942));
  jor  g0870(.dina(n942), .dinb(n941), .dout(n943));
  jor  g0871(.dina(n940), .dinb(n603), .dout(n944));
  jand g0872(.dina(n861), .dinb(n608), .dout(n945));
  jnot g0873(.din(n945), .dout(n946));
  jand g0874(.dina(n623), .dinb(G116), .dout(n947));
  jand g0875(.dina(n617), .dinb(G283), .dout(n948));
  jand g0876(.dina(n642), .dinb(G303), .dout(n949));
  jor  g0877(.dina(n949), .dinb(n948), .dout(n950));
  jor  g0878(.dina(n950), .dinb(n947), .dout(n951));
  jand g0879(.dina(n631), .dinb(G322), .dout(n952));
  jor  g0880(.dina(n952), .dinb(n148), .dout(n953));
  jand g0881(.dina(n636), .dinb(G294), .dout(n954));
  jand g0882(.dina(n627), .dinb(G311), .dout(n955));
  jor  g0883(.dina(n955), .dinb(n954), .dout(n956));
  jand g0884(.dina(n640), .dinb(G317), .dout(n957));
  jor  g0885(.dina(n957), .dinb(n657), .dout(n958));
  jor  g0886(.dina(n958), .dinb(n956), .dout(n959));
  jor  g0887(.dina(n959), .dinb(n953), .dout(n960));
  jor  g0888(.dina(n960), .dinb(n951), .dout(n961));
  jand g0889(.dina(n623), .dinb(G77), .dout(n962));
  jand g0890(.dina(n617), .dinb(G68), .dout(n963));
  jand g0891(.dina(n642), .dinb(G50), .dout(n964));
  jor  g0892(.dina(n964), .dinb(n963), .dout(n965));
  jor  g0893(.dina(n965), .dinb(n962), .dout(n966));
  jand g0894(.dina(n631), .dinb(G143), .dout(n967));
  jor  g0895(.dina(n967), .dinb(G33), .dout(n968));
  jand g0896(.dina(n636), .dinb(G58), .dout(n969));
  jand g0897(.dina(n627), .dinb(G159), .dout(n970));
  jor  g0898(.dina(n970), .dinb(n969), .dout(n971));
  jand g0899(.dina(n640), .dinb(G150), .dout(n972));
  jor  g0900(.dina(n972), .dinb(n728), .dout(n973));
  jor  g0901(.dina(n973), .dinb(n971), .dout(n974));
  jor  g0902(.dina(n974), .dinb(n968), .dout(n975));
  jor  g0903(.dina(n975), .dinb(n966), .dout(n976));
  jand g0904(.dina(n976), .dinb(n961), .dout(n977));
  jor  g0905(.dina(n977), .dinb(n612), .dout(n978));
  jand g0906(.dina(n675), .dinb(n144), .dout(n979));
  jand g0907(.dina(n123), .dinb(G97), .dout(n980));
  jor  g0908(.dina(n980), .dinb(n672), .dout(n981));
  jor  g0909(.dina(n981), .dinb(n979), .dout(n982));
  jand g0910(.dina(n982), .dinb(n604), .dout(n983));
  jand g0911(.dina(n983), .dinb(n978), .dout(n984));
  jand g0912(.dina(n984), .dinb(n946), .dout(n985));
  jnot g0913(.din(n985), .dout(n986));
  jand g0914(.dina(n986), .dinb(n944), .dout(n987));
  jand g0915(.dina(n987), .dinb(n943), .dout(n988));
  jnot g0916(.din(n988), .dout(G390));
  jnot g0917(.din(n758), .dout(n990));
  jand g0918(.dina(n696), .dinb(n588), .dout(n991));
  jand g0919(.dina(n991), .dinb(n764), .dout(n992));
  jxor g0920(.dina(n992), .dinb(n990), .dout(n993));
  jxor g0921(.dina(n993), .dinb(n769), .dout(n994));
  jand g0922(.dina(n589), .dinb(n519), .dout(n995));
  jor  g0923(.dina(n995), .dinb(n548), .dout(n996));
  jand g0924(.dina(n554), .dinb(n404), .dout(n997));
  jor  g0925(.dina(n997), .dinb(n759), .dout(n998));
  jnot g0926(.din(n764), .dout(n999));
  jxor g0927(.dina(n991), .dinb(n999), .dout(n1000));
  jxor g0928(.dina(n1000), .dinb(n998), .dout(n1001));
  jor  g0929(.dina(n1001), .dinb(n996), .dout(n1002));
  jor  g0930(.dina(n1002), .dinb(n994), .dout(n1003));
  jnot g0931(.din(n1003), .dout(n1004));
  jand g0932(.dina(n1002), .dinb(n994), .dout(n1005));
  jor  g0933(.dina(n1005), .dinb(n592), .dout(n1006));
  jor  g0934(.dina(n1006), .dinb(n1004), .dout(n1007));
  jor  g0935(.dina(n994), .dinb(n603), .dout(n1008));
  jand g0936(.dina(n990), .dinb(n425), .dout(n1009));
  jnot g0937(.din(n1009), .dout(n1010));
  jand g0938(.dina(n631), .dinb(G125), .dout(n1011));
  jand g0939(.dina(n623), .dinb(G159), .dout(n1012));
  jand g0940(.dina(n642), .dinb(G137), .dout(n1013));
  jor  g0941(.dina(n1013), .dinb(n1012), .dout(n1014));
  jor  g0942(.dina(n1014), .dinb(n1011), .dout(n1015));
  jand g0943(.dina(n617), .dinb(G150), .dout(n1016));
  jor  g0944(.dina(n1016), .dinb(G33), .dout(n1017));
  jand g0945(.dina(n636), .dinb(G143), .dout(n1018));
  jand g0946(.dina(n627), .dinb(G132), .dout(n1019));
  jor  g0947(.dina(n1019), .dinb(n1018), .dout(n1020));
  jand g0948(.dina(n640), .dinb(G128), .dout(n1021));
  jand g0949(.dina(n634), .dinb(G50), .dout(n1022));
  jor  g0950(.dina(n1022), .dinb(n1021), .dout(n1023));
  jor  g0951(.dina(n1023), .dinb(n1020), .dout(n1024));
  jor  g0952(.dina(n1024), .dinb(n1017), .dout(n1025));
  jor  g0953(.dina(n1025), .dinb(n1015), .dout(n1026));
  jand g0954(.dina(n631), .dinb(G294), .dout(n1027));
  jand g0955(.dina(n642), .dinb(G107), .dout(n1028));
  jor  g0956(.dina(n1028), .dinb(n962), .dout(n1029));
  jor  g0957(.dina(n1029), .dinb(n1027), .dout(n1030));
  jand g0958(.dina(n640), .dinb(G283), .dout(n1031));
  jor  g0959(.dina(n1031), .dinb(n148), .dout(n1032));
  jand g0960(.dina(n636), .dinb(G97), .dout(n1033));
  jand g0961(.dina(n627), .dinb(G116), .dout(n1034));
  jor  g0962(.dina(n1034), .dinb(n1033), .dout(n1035));
  jor  g0963(.dina(n717), .dinb(n654), .dout(n1036));
  jor  g0964(.dina(n1036), .dinb(n1035), .dout(n1037));
  jor  g0965(.dina(n1037), .dinb(n1032), .dout(n1038));
  jor  g0966(.dina(n1038), .dinb(n1030), .dout(n1039));
  jand g0967(.dina(n1039), .dinb(n1026), .dout(n1040));
  jor  g0968(.dina(n1040), .dinb(n612), .dout(n1041));
  jand g0969(.dina(n743), .dinb(n74), .dout(n1042));
  jor  g0970(.dina(n1042), .dinb(n605), .dout(n1043));
  jnot g0971(.din(n1043), .dout(n1044));
  jand g0972(.dina(n1044), .dinb(n1041), .dout(n1045));
  jand g0973(.dina(n1045), .dinb(n1010), .dout(n1046));
  jnot g0974(.din(n1046), .dout(n1047));
  jand g0975(.dina(n1047), .dinb(n1008), .dout(n1048));
  jand g0976(.dina(n1048), .dinb(n1007), .dout(n1049));
  jnot g0977(.din(n1049), .dout(G378));
  jand g0978(.dina(n992), .dinb(n758), .dout(n1051));
  jand g0979(.dina(n552), .dinb(n479), .dout(n1052));
  jnot g0980(.din(n1052), .dout(n1053));
  jand g0981(.dina(n1053), .dinb(n484), .dout(n1054));
  jand g0982(.dina(n1052), .dinb(n541), .dout(n1055));
  jor  g0983(.dina(n1055), .dinb(n1054), .dout(n1056));
  jnot g0984(.din(n1056), .dout(n1057));
  jxor g0985(.dina(n1057), .dinb(n771), .dout(n1058));
  jxor g0986(.dina(n1058), .dinb(n1051), .dout(n1059));
  jor  g0987(.dina(n1059), .dinb(n603), .dout(n1060));
  jnot g0988(.din(n996), .dout(n1061));
  jand g0989(.dina(n1003), .dinb(n1061), .dout(n1062));
  jor  g0990(.dina(n1062), .dinb(n592), .dout(n1063));
  jor  g0991(.dina(n1063), .dinb(n1059), .dout(n1064));
  jand g0992(.dina(n1057), .dinb(n425), .dout(n1065));
  jnot g0993(.din(n612), .dout(n1066));
  jand g0994(.dina(n642), .dinb(G132), .dout(n1067));
  jand g0995(.dina(n627), .dinb(G128), .dout(n1068));
  jand g0996(.dina(n636), .dinb(G137), .dout(n1069));
  jor  g0997(.dina(n1069), .dinb(n1068), .dout(n1070));
  jor  g0998(.dina(n1070), .dinb(n1067), .dout(n1071));
  jnot g0999(.din(n1071), .dout(n1072));
  jand g1000(.dina(n623), .dinb(G150), .dout(n1073));
  jnot g1001(.din(n1073), .dout(n1074));
  jand g1002(.dina(n149), .dinb(n148), .dout(n1075));
  jand g1003(.dina(n1075), .dinb(n1074), .dout(n1076));
  jand g1004(.dina(n640), .dinb(G125), .dout(n1077));
  jand g1005(.dina(n617), .dinb(G143), .dout(n1078));
  jor  g1006(.dina(n1078), .dinb(n1077), .dout(n1079));
  jand g1007(.dina(n631), .dinb(G124), .dout(n1080));
  jand g1008(.dina(n634), .dinb(G159), .dout(n1081));
  jor  g1009(.dina(n1081), .dinb(n1080), .dout(n1082));
  jor  g1010(.dina(n1082), .dinb(n1079), .dout(n1083));
  jnot g1011(.din(n1083), .dout(n1084));
  jand g1012(.dina(n1084), .dinb(n1076), .dout(n1085));
  jand g1013(.dina(n1085), .dinb(n1072), .dout(n1086));
  jand g1014(.dina(n627), .dinb(G107), .dout(n1087));
  jand g1015(.dina(n634), .dinb(G58), .dout(n1088));
  jand g1016(.dina(n636), .dinb(G87), .dout(n1089));
  jor  g1017(.dina(n1089), .dinb(n1088), .dout(n1090));
  jor  g1018(.dina(n1090), .dinb(n1087), .dout(n1091));
  jnot g1019(.din(n1091), .dout(n1092));
  jand g1020(.dina(n642), .dinb(G97), .dout(n1093));
  jnot g1021(.din(n1093), .dout(n1094));
  jand g1022(.dina(n149), .dinb(G33), .dout(n1095));
  jand g1023(.dina(n1095), .dinb(n1094), .dout(n1096));
  jand g1024(.dina(n631), .dinb(G283), .dout(n1097));
  jor  g1025(.dina(n1097), .dinb(n823), .dout(n1098));
  jand g1026(.dina(n640), .dinb(G116), .dout(n1099));
  jor  g1027(.dina(n1099), .dinb(n909), .dout(n1100));
  jor  g1028(.dina(n1100), .dinb(n1098), .dout(n1101));
  jnot g1029(.din(n1101), .dout(n1102));
  jand g1030(.dina(n1102), .dinb(n1096), .dout(n1103));
  jand g1031(.dina(n1103), .dinb(n1092), .dout(n1104));
  jand g1032(.dina(n73), .dinb(G41), .dout(n1105));
  jor  g1033(.dina(n1105), .dinb(n1104), .dout(n1106));
  jor  g1034(.dina(n1106), .dinb(n1086), .dout(n1107));
  jand g1035(.dina(n1107), .dinb(n1066), .dout(n1108));
  jand g1036(.dina(n743), .dinb(n73), .dout(n1109));
  jor  g1037(.dina(n1109), .dinb(n605), .dout(n1110));
  jor  g1038(.dina(n1110), .dinb(n1108), .dout(n1111));
  jor  g1039(.dina(n1111), .dinb(n1065), .dout(n1112));
  jand g1040(.dina(n1112), .dinb(n1064), .dout(n1113));
  jand g1041(.dina(n1113), .dinb(n1060), .dout(n1114));
  jnot g1042(.din(n1114), .dout(G375));
  jand g1043(.dina(n1001), .dinb(n996), .dout(n1116));
  jnot g1044(.din(n1116), .dout(n1117));
  jand g1045(.dina(n1002), .dinb(n591), .dout(n1118));
  jand g1046(.dina(n1118), .dinb(n1117), .dout(n1119));
  jnot g1047(.din(n1119), .dout(n1120));
  jor  g1048(.dina(n1001), .dinb(n603), .dout(n1121));
  jand g1049(.dina(n999), .dinb(n425), .dout(n1122));
  jnot g1050(.din(n1122), .dout(n1123));
  jand g1051(.dina(n623), .dinb(G50), .dout(n1124));
  jand g1052(.dina(n617), .dinb(G159), .dout(n1125));
  jand g1053(.dina(n642), .dinb(G143), .dout(n1126));
  jor  g1054(.dina(n1126), .dinb(n1125), .dout(n1127));
  jor  g1055(.dina(n1127), .dinb(n1124), .dout(n1128));
  jand g1056(.dina(n631), .dinb(G128), .dout(n1129));
  jor  g1057(.dina(n1129), .dinb(G33), .dout(n1130));
  jand g1058(.dina(n636), .dinb(G150), .dout(n1131));
  jand g1059(.dina(n627), .dinb(G137), .dout(n1132));
  jor  g1060(.dina(n1132), .dinb(n1131), .dout(n1133));
  jand g1061(.dina(n640), .dinb(G132), .dout(n1134));
  jor  g1062(.dina(n1134), .dinb(n1088), .dout(n1135));
  jor  g1063(.dina(n1135), .dinb(n1133), .dout(n1136));
  jor  g1064(.dina(n1136), .dinb(n1130), .dout(n1137));
  jor  g1065(.dina(n1137), .dinb(n1128), .dout(n1138));
  jand g1066(.dina(n617), .dinb(G97), .dout(n1139));
  jand g1067(.dina(n640), .dinb(G294), .dout(n1140));
  jand g1068(.dina(n642), .dinb(G116), .dout(n1141));
  jor  g1069(.dina(n1141), .dinb(n1140), .dout(n1142));
  jor  g1070(.dina(n1142), .dinb(n1139), .dout(n1143));
  jand g1071(.dina(n631), .dinb(G303), .dout(n1144));
  jor  g1072(.dina(n1144), .dinb(n148), .dout(n1145));
  jand g1073(.dina(n636), .dinb(G107), .dout(n1146));
  jand g1074(.dina(n627), .dinb(G283), .dout(n1147));
  jor  g1075(.dina(n1147), .dinb(n1146), .dout(n1148));
  jor  g1076(.dina(n899), .dinb(n825), .dout(n1149));
  jor  g1077(.dina(n1149), .dinb(n1148), .dout(n1150));
  jor  g1078(.dina(n1150), .dinb(n1145), .dout(n1151));
  jor  g1079(.dina(n1151), .dinb(n1143), .dout(n1152));
  jand g1080(.dina(n1152), .dinb(n1138), .dout(n1153));
  jor  g1081(.dina(n1153), .dinb(n612), .dout(n1154));
  jand g1082(.dina(n743), .dinb(n75), .dout(n1155));
  jor  g1083(.dina(n1155), .dinb(n605), .dout(n1156));
  jnot g1084(.din(n1156), .dout(n1157));
  jand g1085(.dina(n1157), .dinb(n1154), .dout(n1158));
  jand g1086(.dina(n1158), .dinb(n1123), .dout(n1159));
  jnot g1087(.din(n1159), .dout(n1160));
  jand g1088(.dina(n1160), .dinb(n1121), .dout(n1161));
  jand g1089(.dina(n1161), .dinb(n1120), .dout(n1162));
  jnot g1090(.din(n1162), .dout(G381));
  jand g1091(.dina(n1114), .dinb(n1049), .dout(n1164));
  jnot g1092(.din(G387), .dout(n1165));
  jnot g1093(.din(G396), .dout(n1166));
  jand g1094(.dina(n937), .dinb(n1166), .dout(n1167));
  jand g1095(.dina(n1167), .dinb(n750), .dout(n1168));
  jand g1096(.dina(n1168), .dinb(n988), .dout(n1169));
  jand g1097(.dina(n1169), .dinb(n1162), .dout(n1170));
  jand g1098(.dina(n1170), .dinb(n1165), .dout(n1171));
  jand g1099(.dina(n1171), .dinb(n1164), .dout(n1172));
  jnot g1100(.din(n1172), .dout(G407));
  jnot g1101(.din(G213), .dout(n1174));
  jnot g1102(.din(G343), .dout(n1175));
  jand g1103(.dina(n1164), .dinb(n1175), .dout(n1176));
  jor  g1104(.dina(n1176), .dinb(n1174), .dout(n1177));
  jor  g1105(.dina(n1177), .dinb(n1172), .dout(G409));
  jxor g1106(.dina(n1162), .dinb(G384), .dout(n1179));
  jxor g1107(.dina(n937), .dinb(G396), .dout(n1180));
  jxor g1108(.dina(n988), .dinb(G387), .dout(n1181));
  jxor g1109(.dina(n1181), .dinb(n1180), .dout(n1182));
  jxor g1110(.dina(n1182), .dinb(n1179), .dout(n1183));
  jand g1111(.dina(n1175), .dinb(G213), .dout(n1184));
  jnot g1112(.din(n1184), .dout(n1185));
  jor  g1113(.dina(n1185), .dinb(G2897), .dout(n1186));
  jxor g1114(.dina(n1114), .dinb(n1049), .dout(n1187));
  jor  g1115(.dina(n1187), .dinb(n1184), .dout(n1188));
  jand g1116(.dina(n1188), .dinb(n1186), .dout(n1189));
  jxor g1117(.dina(n1189), .dinb(n1183), .dout(G405));
  jxor g1118(.dina(n1187), .dinb(n1183), .dout(G402));
endmodule


