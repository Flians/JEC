/*

c1908:
	jxor: 78
	jspl: 105
	jspl3: 86
	jnot: 30
	jdff: 163
	jor: 87
	jand: 120

Summary:
	jxor: 78
	jspl: 105
	jspl3: 86
	jnot: 30
	jdff: 163
	jor: 87
	jand: 120

The maximum logic level gap of any gate:
	c1908: 17
*/

module gf_c1908(gclk, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57);
	input gclk;
	input G101;
	input G104;
	input G107;
	input G110;
	input G113;
	input G116;
	input G119;
	input G122;
	input G125;
	input G128;
	input G131;
	input G134;
	input G137;
	input G140;
	input G143;
	input G146;
	input G210;
	input G214;
	input G217;
	input G221;
	input G224;
	input G227;
	input G234;
	input G237;
	input G469;
	input G472;
	input G475;
	input G478;
	input G898;
	input G900;
	input G902;
	input G952;
	input G953;
	output G3;
	output G6;
	output G9;
	output G12;
	output G30;
	output G45;
	output G48;
	output G15;
	output G18;
	output G21;
	output G24;
	output G27;
	output G33;
	output G36;
	output G39;
	output G42;
	output G75;
	output G51;
	output G54;
	output G60;
	output G63;
	output G66;
	output G69;
	output G72;
	output G57;
	wire n58;
	wire n59;
	wire n60;
	wire n61;
	wire n62;
	wire n63;
	wire n64;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n69;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n173;
	wire n174;
	wire n175;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n191;
	wire n192;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n201;
	wire n203;
	wire n204;
	wire n206;
	wire n207;
	wire n208;
	wire n210;
	wire n211;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n220;
	wire n222;
	wire n223;
	wire n224;
	wire n226;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n270;
	wire n271;
	wire n272;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n348;
	wire n349;
	wire n350;
	wire n352;
	wire n353;
	wire n354;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n369;
	wire n370;
	wire n371;
	wire[2:0] w_G101_0;
	wire[2:0] w_G104_0;
	wire[2:0] w_G107_0;
	wire[2:0] w_G110_0;
	wire[2:0] w_G113_0;
	wire[2:0] w_G116_0;
	wire[2:0] w_G119_0;
	wire[2:0] w_G122_0;
	wire[1:0] w_G122_1;
	wire[2:0] w_G125_0;
	wire[2:0] w_G128_0;
	wire[2:0] w_G131_0;
	wire[2:0] w_G134_0;
	wire[2:0] w_G137_0;
	wire[2:0] w_G140_0;
	wire[2:0] w_G143_0;
	wire[2:0] w_G146_0;
	wire[2:0] w_G210_0;
	wire[1:0] w_G214_0;
	wire[2:0] w_G217_0;
	wire[1:0] w_G221_0;
	wire[1:0] w_G224_0;
	wire[1:0] w_G227_0;
	wire[2:0] w_G234_0;
	wire[1:0] w_G234_1;
	wire[2:0] w_G237_0;
	wire[2:0] w_G469_0;
	wire[2:0] w_G472_0;
	wire[2:0] w_G475_0;
	wire[2:0] w_G478_0;
	wire[1:0] w_G898_0;
	wire[1:0] w_G900_0;
	wire[2:0] w_G902_0;
	wire[2:0] w_G902_1;
	wire[2:0] w_G902_2;
	wire[2:0] w_G902_3;
	wire[2:0] w_G952_0;
	wire[2:0] w_G953_0;
	wire[2:0] w_G953_1;
	wire[1:0] w_G953_2;
	wire[2:0] w_n58_0;
	wire[2:0] w_n58_1;
	wire[2:0] w_n58_2;
	wire[1:0] w_n63_0;
	wire[1:0] w_n66_0;
	wire[1:0] w_n67_0;
	wire[1:0] w_n70_0;
	wire[1:0] w_n71_0;
	wire[1:0] w_n73_0;
	wire[1:0] w_n74_0;
	wire[2:0] w_n76_0;
	wire[2:0] w_n76_1;
	wire[1:0] w_n77_0;
	wire[1:0] w_n78_0;
	wire[2:0] w_n81_0;
	wire[1:0] w_n84_0;
	wire[1:0] w_n86_0;
	wire[1:0] w_n90_0;
	wire[1:0] w_n91_0;
	wire[2:0] w_n92_0;
	wire[1:0] w_n92_1;
	wire[2:0] w_n93_0;
	wire[1:0] w_n93_1;
	wire[1:0] w_n94_0;
	wire[2:0] w_n95_0;
	wire[1:0] w_n95_1;
	wire[2:0] w_n96_0;
	wire[1:0] w_n99_0;
	wire[1:0] w_n102_0;
	wire[2:0] w_n103_0;
	wire[2:0] w_n103_1;
	wire[2:0] w_n103_2;
	wire[2:0] w_n103_3;
	wire[1:0] w_n107_0;
	wire[1:0] w_n108_0;
	wire[1:0] w_n109_0;
	wire[1:0] w_n110_0;
	wire[1:0] w_n111_0;
	wire[2:0] w_n112_0;
	wire[1:0] w_n112_1;
	wire[2:0] w_n113_0;
	wire[1:0] w_n118_0;
	wire[1:0] w_n119_0;
	wire[1:0] w_n120_0;
	wire[1:0] w_n121_0;
	wire[2:0] w_n122_0;
	wire[1:0] w_n122_1;
	wire[1:0] w_n124_0;
	wire[1:0] w_n126_0;
	wire[1:0] w_n127_0;
	wire[2:0] w_n130_0;
	wire[1:0] w_n130_1;
	wire[2:0] w_n131_0;
	wire[2:0] w_n131_1;
	wire[1:0] w_n139_0;
	wire[1:0] w_n140_0;
	wire[2:0] w_n141_0;
	wire[1:0] w_n141_1;
	wire[2:0] w_n151_0;
	wire[1:0] w_n152_0;
	wire[2:0] w_n153_0;
	wire[1:0] w_n153_1;
	wire[2:0] w_n154_0;
	wire[1:0] w_n154_1;
	wire[1:0] w_n155_0;
	wire[1:0] w_n156_0;
	wire[1:0] w_n157_0;
	wire[2:0] w_n160_0;
	wire[2:0] w_n160_1;
	wire[2:0] w_n161_0;
	wire[1:0] w_n161_1;
	wire[1:0] w_n162_0;
	wire[2:0] w_n163_0;
	wire[1:0] w_n163_1;
	wire[1:0] w_n164_0;
	wire[2:0] w_n165_0;
	wire[1:0] w_n166_0;
	wire[2:0] w_n168_0;
	wire[1:0] w_n168_1;
	wire[1:0] w_n169_0;
	wire[1:0] w_n170_0;
	wire[1:0] w_n171_0;
	wire[2:0] w_n173_0;
	wire[1:0] w_n173_1;
	wire[1:0] w_n174_0;
	wire[1:0] w_n175_0;
	wire[2:0] w_n177_0;
	wire[1:0] w_n178_0;
	wire[1:0] w_n180_0;
	wire[2:0] w_n182_0;
	wire[2:0] w_n182_1;
	wire[2:0] w_n183_0;
	wire[1:0] w_n184_0;
	wire[1:0] w_n186_0;
	wire[1:0] w_n189_0;
	wire[2:0] w_n191_0;
	wire[2:0] w_n192_0;
	wire[2:0] w_n195_0;
	wire[2:0] w_n197_0;
	wire[1:0] w_n197_1;
	wire[1:0] w_n198_0;
	wire[2:0] w_n199_0;
	wire[1:0] w_n201_0;
	wire[1:0] w_n204_0;
	wire[1:0] w_n206_0;
	wire[1:0] w_n208_0;
	wire[1:0] w_n210_0;
	wire[1:0] w_n211_0;
	wire[2:0] w_n214_0;
	wire[2:0] w_n216_0;
	wire[1:0] w_n216_1;
	wire[1:0] w_n217_0;
	wire[1:0] w_n218_0;
	wire[1:0] w_n220_0;
	wire[1:0] w_n224_0;
	wire[1:0] w_n226_0;
	wire[2:0] w_n242_0;
	wire[2:0] w_n242_1;
	wire[2:0] w_n242_2;
	wire[1:0] w_n243_0;
	wire[1:0] w_n249_0;
	wire[2:0] w_n258_0;
	wire[2:0] w_n265_0;
	wire[2:0] w_n265_1;
	wire[1:0] w_n265_2;
	wire[1:0] w_n274_0;
	wire[2:0] w_n278_0;
	wire[1:0] w_n279_0;
	wire[1:0] w_n280_0;
	wire[2:0] w_n282_0;
	wire[1:0] w_n282_1;
	wire[1:0] w_n286_0;
	wire[2:0] w_n287_0;
	wire[1:0] w_n287_1;
	wire[1:0] w_n288_0;
	wire[2:0] w_n291_0;
	wire[1:0] w_n291_1;
	wire[1:0] w_n292_0;
	wire[1:0] w_n293_0;
	wire[1:0] w_n294_0;
	wire[1:0] w_n297_0;
	wire[1:0] w_n303_0;
	wire[2:0] w_n307_0;
	wire[1:0] w_n313_0;
	wire[2:0] w_n316_0;
	wire[2:0] w_n317_0;
	wire[1:0] w_n322_0;
	wire[1:0] w_n323_0;
	wire[1:0] w_n327_0;
	wire[1:0] w_n329_0;
	wire[1:0] w_n341_0;
	wire w_dff_B_mcx8HXjZ1_0;
	wire w_dff_B_bFOZa4sH6_0;
	wire w_dff_B_grBeq9j94_0;
	wire w_dff_B_9UFfzvlu2_0;
	wire w_dff_B_MLTY3rqi9_0;
	wire w_dff_B_aWYS1ZOy1_1;
	wire w_dff_B_52GnKZf39_1;
	wire w_dff_B_PpmdxMA92_1;
	wire w_dff_B_U0PxIqWc0_1;
	wire w_dff_B_XWZSrCpu1_1;
	wire w_dff_B_AVuulWGR7_1;
	wire w_dff_B_qe0ME2T25_1;
	wire w_dff_B_QKks3Nyo9_1;
	wire w_dff_B_6UoEHvV06_1;
	wire w_dff_B_T0nU5WW41_1;
	wire w_dff_B_4Wvdo2MD6_1;
	wire w_dff_B_r8lSCO022_1;
	wire w_dff_B_k0Z0wKK09_1;
	wire w_dff_B_7VXxI4l23_0;
	wire w_dff_B_i7PbQM5S0_0;
	wire w_dff_B_juNbU65h3_0;
	wire w_dff_B_ZqgcQENp8_0;
	wire w_dff_B_sNEiNVkP9_0;
	wire w_dff_B_uaPcn3RO5_0;
	wire w_dff_B_OQjizde24_0;
	wire w_dff_B_tV1wbGDu1_0;
	wire w_dff_B_ObDKHwKj7_0;
	wire w_dff_B_HoaeaW9F5_0;
	wire w_dff_B_VZ1fJwtq4_0;
	wire w_dff_B_wHVSvMI70_0;
	wire w_dff_A_oVsTq72R1_2;
	wire w_dff_A_0C9ObIdz0_0;
	wire w_dff_A_VTtHXf1F2_0;
	wire w_dff_A_pXh7WgNI4_0;
	wire w_dff_A_v4hP8LCg6_0;
	wire w_dff_A_KvxqVpnN9_0;
	wire w_dff_A_Th9AYmzj6_0;
	wire w_dff_A_aUtnlEKl1_0;
	wire w_dff_A_l0poYgO75_2;
	wire w_dff_A_Ijlgz3FN8_0;
	wire w_dff_A_HS7wqKna6_0;
	wire w_dff_A_cOyKGyYO3_0;
	wire w_dff_A_HYXdyIgm0_0;
	wire w_dff_A_1u6WuHLL3_0;
	wire w_dff_A_J8vR6Aft9_0;
	wire w_dff_A_LMEzXytF4_0;
	wire w_dff_A_YW8W7tRx6_2;
	wire w_dff_A_7jFk8CV00_0;
	wire w_dff_A_yqAu8yh37_0;
	wire w_dff_A_2obB2PTB9_0;
	wire w_dff_A_CcPjPksI8_0;
	wire w_dff_A_YVQrcD270_0;
	wire w_dff_A_dH36MvzL2_0;
	wire w_dff_A_LhoicajQ8_0;
	wire w_dff_A_gGm2HDNQ2_2;
	wire w_dff_A_b5T9GjKi0_0;
	wire w_dff_A_Sk7t9mV98_0;
	wire w_dff_A_lDUlwOQB3_0;
	wire w_dff_A_JuJnZyNl5_0;
	wire w_dff_A_b46OLkIx0_0;
	wire w_dff_A_TRlfbQ617_0;
	wire w_dff_A_TctbjcZR3_0;
	wire w_dff_A_Vp6nTiae6_2;
	wire w_dff_A_24bQa3Bi5_0;
	wire w_dff_A_xrJX33Sg2_0;
	wire w_dff_A_sEvO2muf3_0;
	wire w_dff_A_6J0mkjEY9_0;
	wire w_dff_A_JJVwsxEo3_0;
	wire w_dff_A_WFsMxitT1_0;
	wire w_dff_A_yeCunKXX4_0;
	wire w_dff_A_jKXqwK7t1_2;
	wire w_dff_A_sYAVy6pF3_0;
	wire w_dff_A_KFl9pbzH7_0;
	wire w_dff_A_IFb2x9iA9_0;
	wire w_dff_A_PjYxAS1v3_0;
	wire w_dff_A_tN3SXOc79_0;
	wire w_dff_A_MAPOkg9G3_0;
	wire w_dff_A_GuQUmgZ43_0;
	wire w_dff_A_xLZeIvHB1_2;
	wire w_dff_A_n7FfThNw2_0;
	wire w_dff_A_rv8UR1Ui2_0;
	wire w_dff_A_cTpxm0Z59_0;
	wire w_dff_A_4lzkzswJ4_0;
	wire w_dff_A_g8wPsrTs2_0;
	wire w_dff_A_DKz2k2r71_0;
	wire w_dff_A_UInU27ge7_0;
	wire w_dff_A_iwFOWnuB4_2;
	wire w_dff_A_barZ3sRj6_0;
	wire w_dff_A_CqSBO5hc0_0;
	wire w_dff_A_LUHHYikK1_0;
	wire w_dff_A_PwPyty8z0_0;
	wire w_dff_A_P54LFzTU8_0;
	wire w_dff_A_qdV3DD4Y6_0;
	wire w_dff_A_uAX3FQTh3_0;
	wire w_dff_A_E73ITE3P9_2;
	wire w_dff_A_ySGCkCjc0_0;
	wire w_dff_A_xyA1laYS8_0;
	wire w_dff_A_FS7zwQeQ4_0;
	wire w_dff_A_qtDWqYxR9_0;
	wire w_dff_A_PqOrVhch4_0;
	wire w_dff_A_x8C7AKdU5_0;
	wire w_dff_A_JSgVYWW44_0;
	wire w_dff_A_XOYZZE3e4_2;
	wire w_dff_A_63W526Nc5_0;
	wire w_dff_A_XTsxj5Mo1_0;
	wire w_dff_A_fYeEoUwM2_0;
	wire w_dff_A_SBzPjrmn4_0;
	wire w_dff_A_tgCO6byC4_0;
	wire w_dff_A_ptAm8GdO5_0;
	wire w_dff_A_Eu3Pq5975_0;
	wire w_dff_A_5zLbCwG53_2;
	wire w_dff_A_LweQl56s5_0;
	wire w_dff_A_cgCOdFSo7_0;
	wire w_dff_A_s08SeP1K0_0;
	wire w_dff_A_sUGmBRsO0_0;
	wire w_dff_A_pnuinHEP4_0;
	wire w_dff_A_sUOKxKkw6_0;
	wire w_dff_A_PMMyqFGP2_2;
	wire w_dff_A_e7VnHSKm1_0;
	wire w_dff_A_7OuwsZWL3_0;
	wire w_dff_A_MHfphiOd2_0;
	wire w_dff_A_SBe3M3F32_0;
	wire w_dff_A_FkrH5WKV0_0;
	wire w_dff_A_Cmj6XXNM7_0;
	wire w_dff_A_7SDL1qwd8_0;
	wire w_dff_A_8Vc8w38d7_2;
	wire w_dff_A_gHFDlBjI5_0;
	wire w_dff_A_prqr8yZ23_0;
	wire w_dff_A_BvpQ5XvI6_0;
	wire w_dff_A_XFaziCNF0_0;
	wire w_dff_A_sDqZu0UT6_0;
	wire w_dff_A_pkaiTCoc0_0;
	wire w_dff_A_rBEg7uQw7_0;
	wire w_dff_A_KqOJDCII5_2;
	wire w_dff_A_BJtD2o3t5_0;
	wire w_dff_A_fsUBMFRg8_0;
	wire w_dff_A_U81QikaM4_0;
	wire w_dff_A_enSP1Mit9_0;
	wire w_dff_A_8ZAhcqkK2_0;
	wire w_dff_A_b2nk0cNJ0_0;
	wire w_dff_A_v5lJGdRk4_0;
	wire w_dff_A_K41iITcE1_2;
	wire w_dff_A_V0GzjCRJ0_0;
	wire w_dff_A_nNodPbMX1_0;
	wire w_dff_A_JlUFRsSp1_0;
	wire w_dff_A_5zrBvXGJ2_0;
	wire w_dff_A_ldIo83AH2_0;
	wire w_dff_A_qya9AF8Z2_0;
	wire w_dff_A_6eyP3IdB3_0;
	wire w_dff_A_RLsCUGFu5_2;
	wire w_dff_A_zXDiMy8I2_0;
	wire w_dff_A_TlwsZlB46_0;
	wire w_dff_A_yzDMr6002_0;
	wire w_dff_A_bhmUH3KQ9_0;
	wire w_dff_A_kXM7QATo9_0;
	wire w_dff_A_zVpqac9g1_0;
	wire w_dff_A_d36VfAlB3_0;
	wire w_dff_A_OZrJidH88_2;
	wire w_dff_A_rJpE2Sql2_2;
	wire w_dff_A_6qmy4NLb6_0;
	wire w_dff_A_4zosqtN80_2;
	wire w_dff_A_Etogts5K7_0;
	wire w_dff_A_H21VoaHU2_2;
	jnot g000(.din(w_G902_3[2]),.dout(n58),.clk(gclk));
	jnot g001(.din(w_G221_0[1]),.dout(n59),.clk(gclk));
	jnot g002(.din(w_G234_1[1]),.dout(n60),.clk(gclk));
	jor g003(.dina(w_G953_2[1]),.dinb(n60),.dout(n61),.clk(gclk));
	jor g004(.dina(n61),.dinb(n59),.dout(n62),.clk(gclk));
	jnot g005(.din(w_G110_0[2]),.dout(n63),.clk(gclk));
	jxor g006(.dina(w_G119_0[2]),.dinb(w_n63_0[1]),.dout(n64),.clk(gclk));
	jxor g007(.dina(n64),.dinb(n62),.dout(n65),.clk(gclk));
	jxor g008(.dina(w_G140_0[2]),.dinb(w_G125_0[2]),.dout(n66),.clk(gclk));
	jxor g009(.dina(w_n66_0[1]),.dinb(w_G146_0[2]),.dout(n67),.clk(gclk));
	jxor g010(.dina(w_G137_0[2]),.dinb(w_G128_0[2]),.dout(n68),.clk(gclk));
	jxor g011(.dina(n68),.dinb(w_n67_0[1]),.dout(n69),.clk(gclk));
	jxor g012(.dina(n69),.dinb(n65),.dout(n70),.clk(gclk));
	jand g013(.dina(w_n70_0[1]),.dinb(w_n58_2[2]),.dout(n71),.clk(gclk));
	jand g014(.dina(w_n58_2[1]),.dinb(w_G234_1[0]),.dout(n72),.clk(gclk));
	jnot g015(.din(n72),.dout(n73),.clk(gclk));
	jand g016(.dina(w_n73_0[1]),.dinb(w_G217_0[2]),.dout(n74),.clk(gclk));
	jnot g017(.din(w_n74_0[1]),.dout(n75),.clk(gclk));
	jxor g018(.dina(n75),.dinb(w_n71_0[1]),.dout(n76),.clk(gclk));
	jxor g019(.dina(w_G143_0[2]),.dinb(w_G128_0[1]),.dout(n77),.clk(gclk));
	jxor g020(.dina(w_n77_0[1]),.dinb(w_G146_0[1]),.dout(n78),.clk(gclk));
	jxor g021(.dina(w_G137_0[1]),.dinb(w_G134_0[2]),.dout(n79),.clk(gclk));
	jxor g022(.dina(n79),.dinb(w_G131_0[2]),.dout(n80),.clk(gclk));
	jxor g023(.dina(n80),.dinb(w_n78_0[1]),.dout(n81),.clk(gclk));
	jnot g024(.din(w_G113_0[2]),.dout(n82),.clk(gclk));
	jxor g025(.dina(w_G119_0[1]),.dinb(w_G116_0[2]),.dout(n83),.clk(gclk));
	jxor g026(.dina(n83),.dinb(n82),.dout(n84),.clk(gclk));
	jnot g027(.din(w_G210_0[2]),.dout(n85),.clk(gclk));
	jor g028(.dina(w_G953_2[0]),.dinb(w_G237_0[2]),.dout(n86),.clk(gclk));
	jor g029(.dina(w_n86_0[1]),.dinb(n85),.dout(n87),.clk(gclk));
	jxor g030(.dina(n87),.dinb(w_G101_0[2]),.dout(n88),.clk(gclk));
	jxor g031(.dina(n88),.dinb(w_n84_0[1]),.dout(n89),.clk(gclk));
	jxor g032(.dina(n89),.dinb(w_n81_0[2]),.dout(n90),.clk(gclk));
	jand g033(.dina(w_n90_0[1]),.dinb(w_n58_2[0]),.dout(n91),.clk(gclk));
	jxor g034(.dina(w_n91_0[1]),.dinb(w_G472_0[2]),.dout(n92),.clk(gclk));
	jand g035(.dina(w_n92_1[1]),.dinb(w_n76_1[2]),.dout(n93),.clk(gclk));
	jor g036(.dina(w_G902_3[1]),.dinb(w_G237_0[1]),.dout(n94),.clk(gclk));
	jand g037(.dina(w_n94_0[1]),.dinb(w_G214_0[1]),.dout(n95),.clk(gclk));
	jnot g038(.din(w_n95_1[1]),.dout(n96),.clk(gclk));
	jnot g039(.din(w_G101_0[1]),.dout(n97),.clk(gclk));
	jxor g040(.dina(w_G107_0[2]),.dinb(w_G104_0[2]),.dout(n98),.clk(gclk));
	jxor g041(.dina(n98),.dinb(n97),.dout(n99),.clk(gclk));
	jxor g042(.dina(w_n99_0[1]),.dinb(w_n84_0[0]),.dout(n100),.clk(gclk));
	jxor g043(.dina(w_G122_1[1]),.dinb(w_G110_0[1]),.dout(n101),.clk(gclk));
	jxor g044(.dina(n101),.dinb(n100),.dout(n102),.clk(gclk));
	jnot g045(.din(w_G953_1[2]),.dout(n103),.clk(gclk));
	jand g046(.dina(w_n103_3[2]),.dinb(w_G224_0[1]),.dout(n104),.clk(gclk));
	jxor g047(.dina(w_n78_0[0]),.dinb(w_G125_0[1]),.dout(n105),.clk(gclk));
	jxor g048(.dina(n105),.dinb(n104),.dout(n106),.clk(gclk));
	jxor g049(.dina(n106),.dinb(w_n102_0[1]),.dout(n107),.clk(gclk));
	jand g050(.dina(w_n107_0[1]),.dinb(w_n58_1[2]),.dout(n108),.clk(gclk));
	jand g051(.dina(w_n94_0[0]),.dinb(w_G210_0[1]),.dout(n109),.clk(gclk));
	jxor g052(.dina(w_n109_0[1]),.dinb(w_n108_0[1]),.dout(n110),.clk(gclk));
	jand g053(.dina(w_n110_0[1]),.dinb(w_n96_0[2]),.dout(n111),.clk(gclk));
	jand g054(.dina(w_n73_0[0]),.dinb(w_G221_0[0]),.dout(n112),.clk(gclk));
	jnot g055(.din(w_n112_1[1]),.dout(n113),.clk(gclk));
	jand g056(.dina(w_n103_3[1]),.dinb(w_G227_0[1]),.dout(n114),.clk(gclk));
	jxor g057(.dina(w_G140_0[1]),.dinb(w_n63_0[0]),.dout(n115),.clk(gclk));
	jxor g058(.dina(n115),.dinb(n114),.dout(n116),.clk(gclk));
	jxor g059(.dina(n116),.dinb(w_n99_0[0]),.dout(n117),.clk(gclk));
	jxor g060(.dina(n117),.dinb(w_n81_0[1]),.dout(n118),.clk(gclk));
	jand g061(.dina(w_n118_0[1]),.dinb(w_n58_1[1]),.dout(n119),.clk(gclk));
	jxor g062(.dina(w_n119_0[1]),.dinb(w_G469_0[2]),.dout(n120),.clk(gclk));
	jand g063(.dina(w_n120_0[1]),.dinb(w_n113_0[2]),.dout(n121),.clk(gclk));
	jand g064(.dina(w_n121_0[1]),.dinb(w_n111_0[1]),.dout(n122),.clk(gclk));
	jor g065(.dina(w_n103_3[0]),.dinb(w_G898_0[1]),.dout(n123),.clk(gclk));
	jnot g066(.din(n123),.dout(n124),.clk(gclk));
	jand g067(.dina(w_G237_0[0]),.dinb(w_G234_0[2]),.dout(n125),.clk(gclk));
	jnot g068(.din(n125),.dout(n126),.clk(gclk));
	jand g069(.dina(w_n126_0[1]),.dinb(w_G902_3[0]),.dout(n127),.clk(gclk));
	jand g070(.dina(w_n127_0[1]),.dinb(w_n124_0[1]),.dout(n128),.clk(gclk));
	jand g071(.dina(w_n126_0[0]),.dinb(w_G952_0[2]),.dout(n129),.clk(gclk));
	jand g072(.dina(n129),.dinb(w_n103_2[2]),.dout(n130),.clk(gclk));
	jor g073(.dina(w_n130_1[1]),.dinb(n128),.dout(n131),.clk(gclk));
	jnot g074(.din(w_G478_0[2]),.dout(n132),.clk(gclk));
	jxor g075(.dina(w_n77_0[0]),.dinb(w_G134_0[1]),.dout(n133),.clk(gclk));
	jand g076(.dina(w_n103_2[1]),.dinb(w_G234_0[1]),.dout(n134),.clk(gclk));
	jand g077(.dina(n134),.dinb(w_G217_0[1]),.dout(n135),.clk(gclk));
	jxor g078(.dina(w_G122_1[0]),.dinb(w_G116_0[1]),.dout(n136),.clk(gclk));
	jxor g079(.dina(n136),.dinb(w_G107_0[1]),.dout(n137),.clk(gclk));
	jxor g080(.dina(n137),.dinb(n135),.dout(n138),.clk(gclk));
	jxor g081(.dina(n138),.dinb(n133),.dout(n139),.clk(gclk));
	jand g082(.dina(w_n139_0[1]),.dinb(w_n58_1[0]),.dout(n140),.clk(gclk));
	jxor g083(.dina(w_n140_0[1]),.dinb(n132),.dout(n141),.clk(gclk));
	jnot g084(.din(w_G475_0[2]),.dout(n142),.clk(gclk));
	jxor g085(.dina(w_G122_0[2]),.dinb(w_G113_0[1]),.dout(n143),.clk(gclk));
	jxor g086(.dina(n143),.dinb(w_G104_0[1]),.dout(n144),.clk(gclk));
	jnot g087(.din(w_G214_0[0]),.dout(n145),.clk(gclk));
	jor g088(.dina(w_n86_0[0]),.dinb(n145),.dout(n146),.clk(gclk));
	jnot g089(.din(w_G131_0[1]),.dout(n147),.clk(gclk));
	jxor g090(.dina(w_G143_0[1]),.dinb(n147),.dout(n148),.clk(gclk));
	jxor g091(.dina(n148),.dinb(n146),.dout(n149),.clk(gclk));
	jxor g092(.dina(n149),.dinb(w_n67_0[0]),.dout(n150),.clk(gclk));
	jxor g093(.dina(n150),.dinb(n144),.dout(n151),.clk(gclk));
	jand g094(.dina(w_n151_0[2]),.dinb(w_n58_0[2]),.dout(n152),.clk(gclk));
	jxor g095(.dina(w_n152_0[1]),.dinb(n142),.dout(n153),.clk(gclk));
	jand g096(.dina(w_n153_1[1]),.dinb(w_n141_1[1]),.dout(n154),.clk(gclk));
	jand g097(.dina(w_n154_1[1]),.dinb(w_n131_1[2]),.dout(n155),.clk(gclk));
	jand g098(.dina(w_n155_0[1]),.dinb(w_n122_1[1]),.dout(n156),.clk(gclk));
	jand g099(.dina(w_n156_0[1]),.dinb(w_n93_1[1]),.dout(n157),.clk(gclk));
	jxor g100(.dina(w_n157_0[1]),.dinb(w_G101_0[0]),.dout(w_dff_A_oVsTq72R1_2),.clk(gclk));
	jnot g101(.din(w_G472_0[1]),.dout(n159),.clk(gclk));
	jxor g102(.dina(w_n91_0[0]),.dinb(n159),.dout(n160),.clk(gclk));
	jand g103(.dina(w_n160_1[2]),.dinb(w_n76_1[1]),.dout(n161),.clk(gclk));
	jand g104(.dina(w_n161_1[1]),.dinb(w_n122_1[0]),.dout(n162),.clk(gclk));
	jxor g105(.dina(w_n152_0[0]),.dinb(w_G475_0[1]),.dout(n163),.clk(gclk));
	jand g106(.dina(w_n163_1[1]),.dinb(w_n141_1[0]),.dout(n164),.clk(gclk));
	jand g107(.dina(w_n164_0[1]),.dinb(w_n131_1[1]),.dout(n165),.clk(gclk));
	jand g108(.dina(w_n165_0[2]),.dinb(w_n162_0[1]),.dout(n166),.clk(gclk));
	jxor g109(.dina(w_n166_0[1]),.dinb(w_G104_0[0]),.dout(w_dff_A_l0poYgO75_2),.clk(gclk));
	jxor g110(.dina(w_n140_0[0]),.dinb(w_G478_0[1]),.dout(n168),.clk(gclk));
	jand g111(.dina(w_n153_1[0]),.dinb(w_n168_1[1]),.dout(n169),.clk(gclk));
	jand g112(.dina(w_n169_0[1]),.dinb(w_n131_1[0]),.dout(n170),.clk(gclk));
	jand g113(.dina(w_n170_0[1]),.dinb(w_n162_0[0]),.dout(n171),.clk(gclk));
	jxor g114(.dina(w_n171_0[1]),.dinb(w_G107_0[0]),.dout(w_dff_A_YW8W7tRx6_2),.clk(gclk));
	jxor g115(.dina(w_n74_0[0]),.dinb(w_n71_0[0]),.dout(n173),.clk(gclk));
	jand g116(.dina(w_n160_1[1]),.dinb(w_n173_1[1]),.dout(n174),.clk(gclk));
	jand g117(.dina(w_n174_0[1]),.dinb(w_n156_0[0]),.dout(n175),.clk(gclk));
	jxor g118(.dina(w_n175_0[1]),.dinb(w_G110_0[0]),.dout(w_dff_A_gGm2HDNQ2_2),.clk(gclk));
	jand g119(.dina(w_n92_1[0]),.dinb(w_n173_1[0]),.dout(n177),.clk(gclk));
	jand g120(.dina(w_n177_0[2]),.dinb(w_n122_0[2]),.dout(n178),.clk(gclk));
	jor g121(.dina(w_n103_2[0]),.dinb(w_G900_0[1]),.dout(n179),.clk(gclk));
	jnot g122(.din(n179),.dout(n180),.clk(gclk));
	jand g123(.dina(w_n180_0[1]),.dinb(w_n127_0[0]),.dout(n181),.clk(gclk));
	jor g124(.dina(n181),.dinb(w_n130_1[0]),.dout(n182),.clk(gclk));
	jand g125(.dina(w_n182_1[2]),.dinb(w_n169_0[0]),.dout(n183),.clk(gclk));
	jand g126(.dina(w_n183_0[2]),.dinb(w_n178_0[1]),.dout(n184),.clk(gclk));
	jxor g127(.dina(w_n184_0[1]),.dinb(w_G128_0[0]),.dout(w_dff_A_Vp6nTiae6_2),.clk(gclk));
	jand g128(.dina(w_n163_1[0]),.dinb(w_n168_1[0]),.dout(n186),.clk(gclk));
	jand g129(.dina(w_n186_0[1]),.dinb(w_n93_1[0]),.dout(n187),.clk(gclk));
	jand g130(.dina(n187),.dinb(w_n182_1[1]),.dout(n188),.clk(gclk));
	jand g131(.dina(n188),.dinb(w_n122_0[1]),.dout(n189),.clk(gclk));
	jxor g132(.dina(w_n189_0[1]),.dinb(w_G143_0[0]),.dout(w_dff_A_jKXqwK7t1_2),.clk(gclk));
	jand g133(.dina(w_n182_1[0]),.dinb(w_n164_0[0]),.dout(n191),.clk(gclk));
	jand g134(.dina(w_n191_0[2]),.dinb(w_n178_0[0]),.dout(n192),.clk(gclk));
	jxor g135(.dina(w_n192_0[2]),.dinb(w_G146_0[0]),.dout(w_dff_A_xLZeIvHB1_2),.clk(gclk));
	jnot g136(.din(w_G469_0[1]),.dout(n194),.clk(gclk));
	jxor g137(.dina(w_n119_0[0]),.dinb(n194),.dout(n195),.clk(gclk));
	jand g138(.dina(w_n195_0[2]),.dinb(w_n113_0[1]),.dout(n196),.clk(gclk));
	jand g139(.dina(n196),.dinb(w_n111_0[0]),.dout(n197),.clk(gclk));
	jand g140(.dina(w_n197_1[1]),.dinb(w_n93_0[2]),.dout(n198),.clk(gclk));
	jand g141(.dina(w_n198_0[1]),.dinb(w_n165_0[1]),.dout(n199),.clk(gclk));
	jxor g142(.dina(w_n199_0[2]),.dinb(w_G113_0[0]),.dout(w_dff_A_iwFOWnuB4_2),.clk(gclk));
	jand g143(.dina(w_n198_0[0]),.dinb(w_n170_0[0]),.dout(n201),.clk(gclk));
	jxor g144(.dina(w_n201_0[1]),.dinb(w_G116_0[0]),.dout(w_dff_A_E73ITE3P9_2),.clk(gclk));
	jand g145(.dina(w_n177_0[1]),.dinb(w_n155_0[0]),.dout(n203),.clk(gclk));
	jand g146(.dina(n203),.dinb(w_n197_1[0]),.dout(n204),.clk(gclk));
	jxor g147(.dina(w_n204_0[1]),.dinb(w_G119_0[0]),.dout(w_dff_A_XOYZZE3e4_2),.clk(gclk));
	jand g148(.dina(w_n197_0[2]),.dinb(w_n161_1[0]),.dout(n206),.clk(gclk));
	jand g149(.dina(w_n206_0[1]),.dinb(w_n131_0[2]),.dout(n207),.clk(gclk));
	jand g150(.dina(n207),.dinb(w_n186_0[0]),.dout(n208),.clk(gclk));
	jxor g151(.dina(w_n208_0[1]),.dinb(w_G122_0[1]),.dout(w_dff_A_5zLbCwG53_2),.clk(gclk));
	jand g152(.dina(w_n191_0[1]),.dinb(w_n174_0[0]),.dout(n210),.clk(gclk));
	jand g153(.dina(w_n210_0[1]),.dinb(w_n197_0[1]),.dout(n211),.clk(gclk));
	jxor g154(.dina(w_n211_0[1]),.dinb(w_G125_0[0]),.dout(w_dff_A_PMMyqFGP2_2),.clk(gclk));
	jnot g155(.din(w_n109_0[0]),.dout(n213),.clk(gclk));
	jxor g156(.dina(n213),.dinb(w_n108_0[0]),.dout(n214),.clk(gclk));
	jand g157(.dina(w_n214_0[2]),.dinb(w_n96_0[1]),.dout(n215),.clk(gclk));
	jand g158(.dina(n215),.dinb(w_n121_0[0]),.dout(n216),.clk(gclk));
	jand g159(.dina(w_n216_1[1]),.dinb(w_n93_0[1]),.dout(n217),.clk(gclk));
	jand g160(.dina(w_n217_0[1]),.dinb(w_n191_0[0]),.dout(n218),.clk(gclk));
	jxor g161(.dina(w_n218_0[1]),.dinb(w_G131_0[0]),.dout(w_dff_A_8Vc8w38d7_2),.clk(gclk));
	jand g162(.dina(w_n217_0[0]),.dinb(w_n183_0[1]),.dout(n220),.clk(gclk));
	jxor g163(.dina(w_n220_0[1]),.dinb(w_G134_0[0]),.dout(w_dff_A_KqOJDCII5_2),.clk(gclk));
	jand g164(.dina(w_n177_0[0]),.dinb(w_n154_1[0]),.dout(n222),.clk(gclk));
	jand g165(.dina(n222),.dinb(w_n182_0[2]),.dout(n223),.clk(gclk));
	jand g166(.dina(n223),.dinb(w_n216_1[0]),.dout(n224),.clk(gclk));
	jxor g167(.dina(w_n224_0[1]),.dinb(w_G137_0[0]),.dout(w_dff_A_K41iITcE1_2),.clk(gclk));
	jand g168(.dina(w_n216_0[2]),.dinb(w_n210_0[0]),.dout(n226),.clk(gclk));
	jxor g169(.dina(w_n226_0[1]),.dinb(w_G140_0[0]),.dout(w_dff_A_RLsCUGFu5_2),.clk(gclk));
	jor g170(.dina(w_n171_0[0]),.dinb(w_n157_0[0]),.dout(n228),.clk(gclk));
	jor g171(.dina(n228),.dinb(w_n166_0[0]),.dout(n229),.clk(gclk));
	jor g172(.dina(n229),.dinb(w_n208_0[0]),.dout(n230),.clk(gclk));
	jor g173(.dina(w_n204_0[0]),.dinb(w_n201_0[0]),.dout(n231),.clk(gclk));
	jor g174(.dina(n231),.dinb(w_n175_0[0]),.dout(n232),.clk(gclk));
	jor g175(.dina(n232),.dinb(w_n199_0[1]),.dout(n233),.clk(gclk));
	jor g176(.dina(n233),.dinb(n230),.dout(n234),.clk(gclk));
	jor g177(.dina(w_n226_0[0]),.dinb(w_n224_0[0]),.dout(n235),.clk(gclk));
	jor g178(.dina(n235),.dinb(w_n192_0[1]),.dout(n236),.clk(gclk));
	jor g179(.dina(w_n220_0[0]),.dinb(w_n218_0[0]),.dout(n237),.clk(gclk));
	jor g180(.dina(w_n211_0[0]),.dinb(w_n189_0[0]),.dout(n238),.clk(gclk));
	jor g181(.dina(n238),.dinb(w_n184_0[0]),.dout(n239),.clk(gclk));
	jor g182(.dina(n239),.dinb(n237),.dout(n240),.clk(gclk));
	jor g183(.dina(n240),.dinb(n236),.dout(n241),.clk(gclk));
	jor g184(.dina(n241),.dinb(n234),.dout(n242),.clk(gclk));
	jand g185(.dina(w_n195_0[1]),.dinb(w_n214_0[1]),.dout(n243),.clk(gclk));
	jxor g186(.dina(w_n112_1[0]),.dinb(w_n95_1[0]),.dout(n244),.clk(gclk));
	jand g187(.dina(n244),.dinb(w_n243_0[1]),.dout(n245),.clk(gclk));
	jor g188(.dina(n245),.dinb(w_n216_0[1]),.dout(n246),.clk(gclk));
	jand g189(.dina(n246),.dinb(w_n161_0[2]),.dout(n247),.clk(gclk));
	jand g190(.dina(w_n113_0[0]),.dinb(w_n96_0[0]),.dout(n248),.clk(gclk));
	jand g191(.dina(n248),.dinb(w_n243_0[0]),.dout(n249),.clk(gclk));
	jxor g192(.dina(w_n160_1[0]),.dinb(w_n76_1[0]),.dout(n250),.clk(gclk));
	jand g193(.dina(n250),.dinb(w_n249_0[1]),.dout(n251),.clk(gclk));
	jor g194(.dina(n251),.dinb(w_n206_0[0]),.dout(n252),.clk(gclk));
	jor g195(.dina(n252),.dinb(n247),.dout(n253),.clk(gclk));
	jand g196(.dina(n253),.dinb(w_n154_0[2]),.dout(n254),.clk(gclk));
	jand g197(.dina(n254),.dinb(w_n130_0[2]),.dout(n255),.clk(gclk));
	jor g198(.dina(n255),.dinb(w_n242_2[2]),.dout(n256),.clk(gclk));
	jand g199(.dina(n256),.dinb(w_G952_0[1]),.dout(n257),.clk(gclk));
	jor g200(.dina(w_n153_0[2]),.dinb(w_n141_0[2]),.dout(n258),.clk(gclk));
	jor g201(.dina(w_n154_0[1]),.dinb(w_n130_0[1]),.dout(n259),.clk(gclk));
	jand g202(.dina(n259),.dinb(w_n258_0[2]),.dout(n260),.clk(gclk));
	jand g203(.dina(n260),.dinb(w_n161_0[1]),.dout(n261),.clk(gclk));
	jand g204(.dina(n261),.dinb(w_n249_0[0]),.dout(n262),.clk(gclk));
	jor g205(.dina(n262),.dinb(w_G953_1[1]),.dout(n263),.clk(gclk));
	jor g206(.dina(w_dff_B_MLTY3rqi9_0),.dinb(n257),.dout(w_dff_A_OZrJidH88_2),.clk(gclk));
	jor g207(.dina(w_n103_1[2]),.dinb(w_G952_0[0]),.dout(n265),.clk(gclk));
	jand g208(.dina(w_n242_2[1]),.dinb(w_G210_0[0]),.dout(n266),.clk(gclk));
	jand g209(.dina(n266),.dinb(w_G902_2[2]),.dout(n267),.clk(gclk));
	jxor g210(.dina(n267),.dinb(w_n107_0[0]),.dout(n268),.clk(gclk));
	jand g211(.dina(n268),.dinb(w_n265_2[1]),.dout(G51),.clk(gclk));
	jand g212(.dina(w_n242_2[0]),.dinb(w_G469_0[0]),.dout(n270),.clk(gclk));
	jand g213(.dina(n270),.dinb(w_G902_2[1]),.dout(n271),.clk(gclk));
	jxor g214(.dina(n271),.dinb(w_n118_0[0]),.dout(n272),.clk(gclk));
	jand g215(.dina(n272),.dinb(w_n265_2[0]),.dout(G54),.clk(gclk));
	jand g216(.dina(w_G902_2[0]),.dinb(w_G475_0[0]),.dout(n274),.clk(gclk));
	jand g217(.dina(w_n274_0[1]),.dinb(w_n242_1[2]),.dout(n275),.clk(gclk));
	jor g218(.dina(n275),.dinb(w_n151_0[1]),.dout(n276),.clk(gclk));
	jnot g219(.din(w_n151_0[0]),.dout(n277),.clk(gclk));
	jnot g220(.din(w_n131_0[1]),.dout(n278),.clk(gclk));
	jor g221(.dina(w_n92_0[2]),.dinb(w_n173_0[2]),.dout(n279),.clk(gclk));
	jor g222(.dina(w_n214_0[0]),.dinb(w_n95_0[2]),.dout(n280),.clk(gclk));
	jor g223(.dina(w_n120_0[0]),.dinb(w_n112_0[2]),.dout(n281),.clk(gclk));
	jor g224(.dina(n281),.dinb(w_n280_0[1]),.dout(n282),.clk(gclk));
	jor g225(.dina(w_n282_1[1]),.dinb(w_n279_0[1]),.dout(n283),.clk(gclk));
	jor g226(.dina(n283),.dinb(w_n278_0[2]),.dout(n284),.clk(gclk));
	jor g227(.dina(n284),.dinb(w_n258_0[1]),.dout(n285),.clk(gclk));
	jor g228(.dina(w_n195_0[0]),.dinb(w_n112_0[1]),.dout(n286),.clk(gclk));
	jor g229(.dina(w_n286_0[1]),.dinb(w_n280_0[0]),.dout(n287),.clk(gclk));
	jor g230(.dina(w_n279_0[0]),.dinb(w_n287_1[1]),.dout(n288),.clk(gclk));
	jnot g231(.din(w_n165_0[0]),.dout(n289),.clk(gclk));
	jor g232(.dina(n289),.dinb(w_n288_0[1]),.dout(n290),.clk(gclk));
	jor g233(.dina(w_n160_0[2]),.dinb(w_n173_0[1]),.dout(n291),.clk(gclk));
	jor g234(.dina(w_n163_0[2]),.dinb(w_n168_0[2]),.dout(n292),.clk(gclk));
	jor g235(.dina(w_n292_0[1]),.dinb(w_n278_0[1]),.dout(n293),.clk(gclk));
	jor g236(.dina(w_n293_0[1]),.dinb(w_n287_1[0]),.dout(n294),.clk(gclk));
	jor g237(.dina(w_n294_0[1]),.dinb(w_n291_1[1]),.dout(n295),.clk(gclk));
	jor g238(.dina(w_n163_0[1]),.dinb(w_n141_0[1]),.dout(n296),.clk(gclk));
	jor g239(.dina(n296),.dinb(w_n278_0[0]),.dout(n297),.clk(gclk));
	jor g240(.dina(w_n297_0[1]),.dinb(w_n288_0[0]),.dout(n298),.clk(gclk));
	jand g241(.dina(n298),.dinb(n295),.dout(n299),.clk(gclk));
	jand g242(.dina(n299),.dinb(n290),.dout(n300),.clk(gclk));
	jand g243(.dina(n300),.dinb(n285),.dout(n301),.clk(gclk));
	jnot g244(.din(w_n199_0[0]),.dout(n302),.clk(gclk));
	jor g245(.dina(w_n92_0[1]),.dinb(w_n76_0[2]),.dout(n303),.clk(gclk));
	jor g246(.dina(w_n303_0[1]),.dinb(w_n294_0[0]),.dout(n304),.clk(gclk));
	jor g247(.dina(w_n282_1[0]),.dinb(w_n291_1[0]),.dout(n305),.clk(gclk));
	jor g248(.dina(n305),.dinb(w_n297_0[0]),.dout(n306),.clk(gclk));
	jor g249(.dina(w_n160_0[1]),.dinb(w_n76_0[1]),.dout(n307),.clk(gclk));
	jor g250(.dina(w_n307_0[2]),.dinb(w_n293_0[0]),.dout(n308),.clk(gclk));
	jor g251(.dina(n308),.dinb(w_n282_0[2]),.dout(n309),.clk(gclk));
	jand g252(.dina(n309),.dinb(n306),.dout(n310),.clk(gclk));
	jand g253(.dina(n310),.dinb(n304),.dout(n311),.clk(gclk));
	jand g254(.dina(n311),.dinb(n302),.dout(n312),.clk(gclk));
	jand g255(.dina(n312),.dinb(n301),.dout(n313),.clk(gclk));
	jnot g256(.din(w_n192_0[0]),.dout(n314),.clk(gclk));
	jor g257(.dina(w_n110_0[0]),.dinb(w_n95_0[1]),.dout(n315),.clk(gclk));
	jor g258(.dina(n315),.dinb(w_n286_0[0]),.dout(n316),.clk(gclk));
	jnot g259(.din(w_n182_0[1]),.dout(n317),.clk(gclk));
	jor g260(.dina(w_n307_0[1]),.dinb(w_n292_0[0]),.dout(n318),.clk(gclk));
	jor g261(.dina(n318),.dinb(w_n317_0[2]),.dout(n319),.clk(gclk));
	jor g262(.dina(n319),.dinb(w_n316_0[2]),.dout(n320),.clk(gclk));
	jor g263(.dina(w_n153_0[1]),.dinb(w_n168_0[1]),.dout(n321),.clk(gclk));
	jor g264(.dina(w_n317_0[1]),.dinb(n321),.dout(n322),.clk(gclk));
	jor g265(.dina(w_n322_0[1]),.dinb(w_n303_0[0]),.dout(n323),.clk(gclk));
	jor g266(.dina(w_n316_0[1]),.dinb(w_n323_0[1]),.dout(n324),.clk(gclk));
	jand g267(.dina(n324),.dinb(n320),.dout(n325),.clk(gclk));
	jand g268(.dina(n325),.dinb(n314),.dout(n326),.clk(gclk));
	jor g269(.dina(w_n316_0[0]),.dinb(w_n291_0[2]),.dout(n327),.clk(gclk));
	jor g270(.dina(w_n327_0[1]),.dinb(w_n322_0[0]),.dout(n328),.clk(gclk));
	jnot g271(.din(w_n183_0[0]),.dout(n329),.clk(gclk));
	jor g272(.dina(w_n327_0[0]),.dinb(w_n329_0[1]),.dout(n330),.clk(gclk));
	jand g273(.dina(n330),.dinb(n328),.dout(n331),.clk(gclk));
	jor g274(.dina(w_n307_0[0]),.dinb(w_n287_0[2]),.dout(n332),.clk(gclk));
	jor g275(.dina(w_n329_0[0]),.dinb(n332),.dout(n333),.clk(gclk));
	jor g276(.dina(w_n258_0[0]),.dinb(w_n291_0[1]),.dout(n334),.clk(gclk));
	jor g277(.dina(n334),.dinb(w_n317_0[0]),.dout(n335),.clk(gclk));
	jor g278(.dina(n335),.dinb(w_n287_0[1]),.dout(n336),.clk(gclk));
	jor g279(.dina(w_n323_0[0]),.dinb(w_n282_0[1]),.dout(n337),.clk(gclk));
	jand g280(.dina(n337),.dinb(n336),.dout(n338),.clk(gclk));
	jand g281(.dina(n338),.dinb(n333),.dout(n339),.clk(gclk));
	jand g282(.dina(n339),.dinb(n331),.dout(n340),.clk(gclk));
	jand g283(.dina(n340),.dinb(n326),.dout(n341),.clk(gclk));
	jand g284(.dina(w_n341_0[1]),.dinb(w_n313_0[1]),.dout(n342),.clk(gclk));
	jnot g285(.din(w_n274_0[0]),.dout(n343),.clk(gclk));
	jor g286(.dina(n343),.dinb(n342),.dout(n344),.clk(gclk));
	jor g287(.dina(n344),.dinb(n277),.dout(n345),.clk(gclk));
	jand g288(.dina(n345),.dinb(w_n265_1[2]),.dout(n346),.clk(gclk));
	jand g289(.dina(n346),.dinb(w_dff_B_aWYS1ZOy1_1),.dout(G60),.clk(gclk));
	jand g290(.dina(w_n242_1[1]),.dinb(w_G478_0[0]),.dout(n348),.clk(gclk));
	jand g291(.dina(n348),.dinb(w_G902_1[2]),.dout(n349),.clk(gclk));
	jxor g292(.dina(n349),.dinb(w_n139_0[0]),.dout(n350),.clk(gclk));
	jand g293(.dina(n350),.dinb(w_n265_1[1]),.dout(G63),.clk(gclk));
	jand g294(.dina(w_n242_1[0]),.dinb(w_G217_0[0]),.dout(n352),.clk(gclk));
	jand g295(.dina(n352),.dinb(w_G902_1[1]),.dout(n353),.clk(gclk));
	jxor g296(.dina(n353),.dinb(w_n70_0[0]),.dout(n354),.clk(gclk));
	jand g297(.dina(n354),.dinb(w_n265_1[0]),.dout(G66),.clk(gclk));
	jor g298(.dina(w_n124_0[0]),.dinb(w_n102_0[0]),.dout(n356),.clk(gclk));
	jor g299(.dina(w_n313_0[0]),.dinb(w_G953_1[0]),.dout(n357),.clk(gclk));
	jand g300(.dina(w_G898_0[0]),.dinb(w_G224_0[0]),.dout(n358),.clk(gclk));
	jor g301(.dina(n358),.dinb(w_n103_1[1]),.dout(n359),.clk(gclk));
	jand g302(.dina(n359),.dinb(n357),.dout(n360),.clk(gclk));
	jxor g303(.dina(n360),.dinb(w_dff_B_k0Z0wKK09_1),.dout(w_dff_A_rJpE2Sql2_2),.clk(gclk));
	jor g304(.dina(w_n341_0[0]),.dinb(w_G953_0[2]),.dout(n362),.clk(gclk));
	jand g305(.dina(w_G900_0[0]),.dinb(w_G227_0[0]),.dout(n363),.clk(gclk));
	jor g306(.dina(n363),.dinb(w_n103_1[0]),.dout(n364),.clk(gclk));
	jand g307(.dina(n364),.dinb(n362),.dout(n365),.clk(gclk));
	jxor g308(.dina(w_n81_0[0]),.dinb(w_n66_0[0]),.dout(n366),.clk(gclk));
	jor g309(.dina(n366),.dinb(w_n180_0[0]),.dout(n367),.clk(gclk));
	jxor g310(.dina(w_dff_B_wHVSvMI70_0),.dinb(n365),.dout(w_dff_A_4zosqtN80_2),.clk(gclk));
	jand g311(.dina(w_G902_1[0]),.dinb(w_G472_0[0]),.dout(n369),.clk(gclk));
	jand g312(.dina(n369),.dinb(w_n242_0[2]),.dout(n370),.clk(gclk));
	jxor g313(.dina(n370),.dinb(w_n90_0[0]),.dout(n371),.clk(gclk));
	jand g314(.dina(n371),.dinb(w_n265_0[2]),.dout(w_dff_A_H21VoaHU2_2),.clk(gclk));
	jspl3 jspl3_w_G101_0(.douta(w_G101_0[0]),.doutb(w_G101_0[1]),.doutc(w_G101_0[2]),.din(G101));
	jspl3 jspl3_w_G104_0(.douta(w_G104_0[0]),.doutb(w_G104_0[1]),.doutc(w_G104_0[2]),.din(G104));
	jspl3 jspl3_w_G107_0(.douta(w_G107_0[0]),.doutb(w_G107_0[1]),.doutc(w_G107_0[2]),.din(G107));
	jspl3 jspl3_w_G110_0(.douta(w_G110_0[0]),.doutb(w_G110_0[1]),.doutc(w_G110_0[2]),.din(G110));
	jspl3 jspl3_w_G113_0(.douta(w_G113_0[0]),.doutb(w_G113_0[1]),.doutc(w_G113_0[2]),.din(G113));
	jspl3 jspl3_w_G116_0(.douta(w_G116_0[0]),.doutb(w_G116_0[1]),.doutc(w_G116_0[2]),.din(G116));
	jspl3 jspl3_w_G119_0(.douta(w_G119_0[0]),.doutb(w_G119_0[1]),.doutc(w_G119_0[2]),.din(G119));
	jspl3 jspl3_w_G122_0(.douta(w_G122_0[0]),.doutb(w_G122_0[1]),.doutc(w_G122_0[2]),.din(G122));
	jspl jspl_w_G122_1(.douta(w_G122_1[0]),.doutb(w_G122_1[1]),.din(w_G122_0[0]));
	jspl3 jspl3_w_G125_0(.douta(w_G125_0[0]),.doutb(w_G125_0[1]),.doutc(w_G125_0[2]),.din(G125));
	jspl3 jspl3_w_G128_0(.douta(w_G128_0[0]),.doutb(w_G128_0[1]),.doutc(w_G128_0[2]),.din(G128));
	jspl3 jspl3_w_G131_0(.douta(w_G131_0[0]),.doutb(w_G131_0[1]),.doutc(w_G131_0[2]),.din(G131));
	jspl3 jspl3_w_G134_0(.douta(w_G134_0[0]),.doutb(w_G134_0[1]),.doutc(w_G134_0[2]),.din(G134));
	jspl3 jspl3_w_G137_0(.douta(w_G137_0[0]),.doutb(w_G137_0[1]),.doutc(w_G137_0[2]),.din(G137));
	jspl3 jspl3_w_G140_0(.douta(w_G140_0[0]),.doutb(w_G140_0[1]),.doutc(w_G140_0[2]),.din(G140));
	jspl3 jspl3_w_G143_0(.douta(w_G143_0[0]),.doutb(w_G143_0[1]),.doutc(w_G143_0[2]),.din(G143));
	jspl3 jspl3_w_G146_0(.douta(w_G146_0[0]),.doutb(w_G146_0[1]),.doutc(w_G146_0[2]),.din(G146));
	jspl3 jspl3_w_G210_0(.douta(w_G210_0[0]),.doutb(w_G210_0[1]),.doutc(w_G210_0[2]),.din(G210));
	jspl jspl_w_G214_0(.douta(w_G214_0[0]),.doutb(w_G214_0[1]),.din(G214));
	jspl3 jspl3_w_G217_0(.douta(w_G217_0[0]),.doutb(w_G217_0[1]),.doutc(w_G217_0[2]),.din(G217));
	jspl jspl_w_G221_0(.douta(w_G221_0[0]),.doutb(w_G221_0[1]),.din(G221));
	jspl jspl_w_G224_0(.douta(w_G224_0[0]),.doutb(w_G224_0[1]),.din(G224));
	jspl jspl_w_G227_0(.douta(w_G227_0[0]),.doutb(w_G227_0[1]),.din(G227));
	jspl3 jspl3_w_G234_0(.douta(w_G234_0[0]),.doutb(w_G234_0[1]),.doutc(w_G234_0[2]),.din(G234));
	jspl jspl_w_G234_1(.douta(w_G234_1[0]),.doutb(w_G234_1[1]),.din(w_G234_0[0]));
	jspl3 jspl3_w_G237_0(.douta(w_G237_0[0]),.doutb(w_G237_0[1]),.doutc(w_G237_0[2]),.din(G237));
	jspl3 jspl3_w_G469_0(.douta(w_G469_0[0]),.doutb(w_G469_0[1]),.doutc(w_G469_0[2]),.din(G469));
	jspl3 jspl3_w_G472_0(.douta(w_G472_0[0]),.doutb(w_G472_0[1]),.doutc(w_G472_0[2]),.din(G472));
	jspl3 jspl3_w_G475_0(.douta(w_G475_0[0]),.doutb(w_G475_0[1]),.doutc(w_G475_0[2]),.din(G475));
	jspl3 jspl3_w_G478_0(.douta(w_G478_0[0]),.doutb(w_G478_0[1]),.doutc(w_G478_0[2]),.din(G478));
	jspl jspl_w_G898_0(.douta(w_G898_0[0]),.doutb(w_G898_0[1]),.din(G898));
	jspl jspl_w_G900_0(.douta(w_G900_0[0]),.doutb(w_G900_0[1]),.din(G900));
	jspl3 jspl3_w_G902_0(.douta(w_G902_0[0]),.doutb(w_G902_0[1]),.doutc(w_G902_0[2]),.din(G902));
	jspl3 jspl3_w_G902_1(.douta(w_G902_1[0]),.doutb(w_G902_1[1]),.doutc(w_G902_1[2]),.din(w_G902_0[0]));
	jspl3 jspl3_w_G902_2(.douta(w_G902_2[0]),.doutb(w_G902_2[1]),.doutc(w_G902_2[2]),.din(w_G902_0[1]));
	jspl3 jspl3_w_G902_3(.douta(w_G902_3[0]),.doutb(w_G902_3[1]),.doutc(w_G902_3[2]),.din(w_G902_0[2]));
	jspl3 jspl3_w_G952_0(.douta(w_G952_0[0]),.doutb(w_G952_0[1]),.doutc(w_G952_0[2]),.din(G952));
	jspl3 jspl3_w_G953_0(.douta(w_G953_0[0]),.doutb(w_G953_0[1]),.doutc(w_G953_0[2]),.din(G953));
	jspl3 jspl3_w_G953_1(.douta(w_G953_1[0]),.doutb(w_G953_1[1]),.doutc(w_G953_1[2]),.din(w_G953_0[0]));
	jspl jspl_w_G953_2(.douta(w_G953_2[0]),.doutb(w_G953_2[1]),.din(w_G953_0[1]));
	jspl3 jspl3_w_n58_0(.douta(w_n58_0[0]),.doutb(w_n58_0[1]),.doutc(w_n58_0[2]),.din(n58));
	jspl3 jspl3_w_n58_1(.douta(w_n58_1[0]),.doutb(w_n58_1[1]),.doutc(w_n58_1[2]),.din(w_n58_0[0]));
	jspl3 jspl3_w_n58_2(.douta(w_n58_2[0]),.doutb(w_n58_2[1]),.doutc(w_n58_2[2]),.din(w_n58_0[1]));
	jspl jspl_w_n63_0(.douta(w_n63_0[0]),.doutb(w_n63_0[1]),.din(n63));
	jspl jspl_w_n66_0(.douta(w_n66_0[0]),.doutb(w_n66_0[1]),.din(n66));
	jspl jspl_w_n67_0(.douta(w_n67_0[0]),.doutb(w_n67_0[1]),.din(n67));
	jspl jspl_w_n70_0(.douta(w_n70_0[0]),.doutb(w_n70_0[1]),.din(n70));
	jspl jspl_w_n71_0(.douta(w_n71_0[0]),.doutb(w_n71_0[1]),.din(n71));
	jspl jspl_w_n73_0(.douta(w_n73_0[0]),.doutb(w_n73_0[1]),.din(n73));
	jspl jspl_w_n74_0(.douta(w_n74_0[0]),.doutb(w_n74_0[1]),.din(n74));
	jspl3 jspl3_w_n76_0(.douta(w_n76_0[0]),.doutb(w_n76_0[1]),.doutc(w_n76_0[2]),.din(n76));
	jspl3 jspl3_w_n76_1(.douta(w_n76_1[0]),.doutb(w_n76_1[1]),.doutc(w_n76_1[2]),.din(w_n76_0[0]));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl jspl_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.din(n78));
	jspl3 jspl3_w_n81_0(.douta(w_n81_0[0]),.doutb(w_n81_0[1]),.doutc(w_n81_0[2]),.din(n81));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n90_0(.douta(w_n90_0[0]),.doutb(w_n90_0[1]),.din(n90));
	jspl jspl_w_n91_0(.douta(w_n91_0[0]),.doutb(w_n91_0[1]),.din(n91));
	jspl3 jspl3_w_n92_0(.douta(w_n92_0[0]),.doutb(w_n92_0[1]),.doutc(w_n92_0[2]),.din(n92));
	jspl jspl_w_n92_1(.douta(w_n92_1[0]),.doutb(w_n92_1[1]),.din(w_n92_0[0]));
	jspl3 jspl3_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.doutc(w_n93_0[2]),.din(n93));
	jspl jspl_w_n93_1(.douta(w_n93_1[0]),.doutb(w_n93_1[1]),.din(w_n93_0[0]));
	jspl jspl_w_n94_0(.douta(w_n94_0[0]),.doutb(w_n94_0[1]),.din(n94));
	jspl3 jspl3_w_n95_0(.douta(w_n95_0[0]),.doutb(w_n95_0[1]),.doutc(w_n95_0[2]),.din(n95));
	jspl jspl_w_n95_1(.douta(w_n95_1[0]),.doutb(w_n95_1[1]),.din(w_n95_0[0]));
	jspl3 jspl3_w_n96_0(.douta(w_n96_0[0]),.doutb(w_n96_0[1]),.doutc(w_n96_0[2]),.din(n96));
	jspl jspl_w_n99_0(.douta(w_n99_0[0]),.doutb(w_n99_0[1]),.din(n99));
	jspl jspl_w_n102_0(.douta(w_n102_0[0]),.doutb(w_n102_0[1]),.din(n102));
	jspl3 jspl3_w_n103_0(.douta(w_n103_0[0]),.doutb(w_n103_0[1]),.doutc(w_n103_0[2]),.din(n103));
	jspl3 jspl3_w_n103_1(.douta(w_n103_1[0]),.doutb(w_n103_1[1]),.doutc(w_n103_1[2]),.din(w_n103_0[0]));
	jspl3 jspl3_w_n103_2(.douta(w_n103_2[0]),.doutb(w_n103_2[1]),.doutc(w_n103_2[2]),.din(w_n103_0[1]));
	jspl3 jspl3_w_n103_3(.douta(w_n103_3[0]),.doutb(w_n103_3[1]),.doutc(w_n103_3[2]),.din(w_n103_0[2]));
	jspl jspl_w_n107_0(.douta(w_n107_0[0]),.doutb(w_n107_0[1]),.din(n107));
	jspl jspl_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n109_0(.douta(w_n109_0[0]),.doutb(w_n109_0[1]),.din(n109));
	jspl jspl_w_n110_0(.douta(w_n110_0[0]),.doutb(w_n110_0[1]),.din(n110));
	jspl jspl_w_n111_0(.douta(w_n111_0[0]),.doutb(w_n111_0[1]),.din(n111));
	jspl3 jspl3_w_n112_0(.douta(w_n112_0[0]),.doutb(w_n112_0[1]),.doutc(w_n112_0[2]),.din(n112));
	jspl jspl_w_n112_1(.douta(w_n112_1[0]),.doutb(w_n112_1[1]),.din(w_n112_0[0]));
	jspl3 jspl3_w_n113_0(.douta(w_n113_0[0]),.doutb(w_n113_0[1]),.doutc(w_n113_0[2]),.din(n113));
	jspl jspl_w_n118_0(.douta(w_n118_0[0]),.doutb(w_n118_0[1]),.din(n118));
	jspl jspl_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.din(n119));
	jspl jspl_w_n120_0(.douta(w_n120_0[0]),.doutb(w_n120_0[1]),.din(n120));
	jspl jspl_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.din(n121));
	jspl3 jspl3_w_n122_0(.douta(w_n122_0[0]),.doutb(w_n122_0[1]),.doutc(w_n122_0[2]),.din(n122));
	jspl jspl_w_n122_1(.douta(w_n122_1[0]),.doutb(w_n122_1[1]),.din(w_n122_0[0]));
	jspl jspl_w_n124_0(.douta(w_n124_0[0]),.doutb(w_n124_0[1]),.din(n124));
	jspl jspl_w_n126_0(.douta(w_n126_0[0]),.doutb(w_n126_0[1]),.din(n126));
	jspl jspl_w_n127_0(.douta(w_n127_0[0]),.doutb(w_n127_0[1]),.din(n127));
	jspl3 jspl3_w_n130_0(.douta(w_n130_0[0]),.doutb(w_n130_0[1]),.doutc(w_n130_0[2]),.din(n130));
	jspl jspl_w_n130_1(.douta(w_n130_1[0]),.doutb(w_n130_1[1]),.din(w_n130_0[0]));
	jspl3 jspl3_w_n131_0(.douta(w_n131_0[0]),.doutb(w_n131_0[1]),.doutc(w_n131_0[2]),.din(n131));
	jspl3 jspl3_w_n131_1(.douta(w_n131_1[0]),.doutb(w_n131_1[1]),.doutc(w_n131_1[2]),.din(w_n131_0[0]));
	jspl jspl_w_n139_0(.douta(w_n139_0[0]),.doutb(w_n139_0[1]),.din(n139));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl3 jspl3_w_n141_0(.douta(w_n141_0[0]),.doutb(w_n141_0[1]),.doutc(w_n141_0[2]),.din(n141));
	jspl jspl_w_n141_1(.douta(w_n141_1[0]),.doutb(w_n141_1[1]),.din(w_n141_0[0]));
	jspl3 jspl3_w_n151_0(.douta(w_n151_0[0]),.doutb(w_n151_0[1]),.doutc(w_n151_0[2]),.din(n151));
	jspl jspl_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.din(n152));
	jspl3 jspl3_w_n153_0(.douta(w_n153_0[0]),.doutb(w_n153_0[1]),.doutc(w_n153_0[2]),.din(n153));
	jspl jspl_w_n153_1(.douta(w_n153_1[0]),.doutb(w_n153_1[1]),.din(w_n153_0[0]));
	jspl3 jspl3_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.doutc(w_n154_0[2]),.din(n154));
	jspl jspl_w_n154_1(.douta(w_n154_1[0]),.doutb(w_n154_1[1]),.din(w_n154_0[0]));
	jspl jspl_w_n155_0(.douta(w_n155_0[0]),.doutb(w_n155_0[1]),.din(n155));
	jspl jspl_w_n156_0(.douta(w_n156_0[0]),.doutb(w_n156_0[1]),.din(n156));
	jspl jspl_w_n157_0(.douta(w_n157_0[0]),.doutb(w_n157_0[1]),.din(n157));
	jspl3 jspl3_w_n160_0(.douta(w_n160_0[0]),.doutb(w_n160_0[1]),.doutc(w_n160_0[2]),.din(n160));
	jspl3 jspl3_w_n160_1(.douta(w_n160_1[0]),.doutb(w_n160_1[1]),.doutc(w_n160_1[2]),.din(w_n160_0[0]));
	jspl3 jspl3_w_n161_0(.douta(w_n161_0[0]),.doutb(w_n161_0[1]),.doutc(w_n161_0[2]),.din(n161));
	jspl jspl_w_n161_1(.douta(w_n161_1[0]),.doutb(w_n161_1[1]),.din(w_n161_0[0]));
	jspl jspl_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.din(n162));
	jspl3 jspl3_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.doutc(w_n163_0[2]),.din(n163));
	jspl jspl_w_n163_1(.douta(w_n163_1[0]),.doutb(w_n163_1[1]),.din(w_n163_0[0]));
	jspl jspl_w_n164_0(.douta(w_n164_0[0]),.doutb(w_n164_0[1]),.din(n164));
	jspl3 jspl3_w_n165_0(.douta(w_n165_0[0]),.doutb(w_n165_0[1]),.doutc(w_n165_0[2]),.din(n165));
	jspl jspl_w_n166_0(.douta(w_n166_0[0]),.doutb(w_n166_0[1]),.din(n166));
	jspl3 jspl3_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.doutc(w_n168_0[2]),.din(n168));
	jspl jspl_w_n168_1(.douta(w_n168_1[0]),.doutb(w_n168_1[1]),.din(w_n168_0[0]));
	jspl jspl_w_n169_0(.douta(w_n169_0[0]),.doutb(w_n169_0[1]),.din(n169));
	jspl jspl_w_n170_0(.douta(w_n170_0[0]),.doutb(w_n170_0[1]),.din(n170));
	jspl jspl_w_n171_0(.douta(w_n171_0[0]),.doutb(w_n171_0[1]),.din(n171));
	jspl3 jspl3_w_n173_0(.douta(w_n173_0[0]),.doutb(w_n173_0[1]),.doutc(w_n173_0[2]),.din(n173));
	jspl jspl_w_n173_1(.douta(w_n173_1[0]),.doutb(w_n173_1[1]),.din(w_n173_0[0]));
	jspl jspl_w_n174_0(.douta(w_n174_0[0]),.doutb(w_n174_0[1]),.din(n174));
	jspl jspl_w_n175_0(.douta(w_n175_0[0]),.doutb(w_n175_0[1]),.din(n175));
	jspl3 jspl3_w_n177_0(.douta(w_n177_0[0]),.doutb(w_n177_0[1]),.doutc(w_n177_0[2]),.din(n177));
	jspl jspl_w_n178_0(.douta(w_n178_0[0]),.doutb(w_n178_0[1]),.din(n178));
	jspl jspl_w_n180_0(.douta(w_n180_0[0]),.doutb(w_n180_0[1]),.din(n180));
	jspl3 jspl3_w_n182_0(.douta(w_n182_0[0]),.doutb(w_n182_0[1]),.doutc(w_n182_0[2]),.din(n182));
	jspl3 jspl3_w_n182_1(.douta(w_n182_1[0]),.doutb(w_n182_1[1]),.doutc(w_n182_1[2]),.din(w_n182_0[0]));
	jspl3 jspl3_w_n183_0(.douta(w_n183_0[0]),.doutb(w_n183_0[1]),.doutc(w_n183_0[2]),.din(n183));
	jspl jspl_w_n184_0(.douta(w_n184_0[0]),.doutb(w_n184_0[1]),.din(n184));
	jspl jspl_w_n186_0(.douta(w_n186_0[0]),.doutb(w_n186_0[1]),.din(n186));
	jspl jspl_w_n189_0(.douta(w_n189_0[0]),.doutb(w_n189_0[1]),.din(n189));
	jspl3 jspl3_w_n191_0(.douta(w_n191_0[0]),.doutb(w_n191_0[1]),.doutc(w_n191_0[2]),.din(n191));
	jspl3 jspl3_w_n192_0(.douta(w_n192_0[0]),.doutb(w_n192_0[1]),.doutc(w_n192_0[2]),.din(n192));
	jspl3 jspl3_w_n195_0(.douta(w_n195_0[0]),.doutb(w_n195_0[1]),.doutc(w_n195_0[2]),.din(n195));
	jspl3 jspl3_w_n197_0(.douta(w_n197_0[0]),.doutb(w_n197_0[1]),.doutc(w_n197_0[2]),.din(n197));
	jspl jspl_w_n197_1(.douta(w_n197_1[0]),.doutb(w_n197_1[1]),.din(w_n197_0[0]));
	jspl jspl_w_n198_0(.douta(w_n198_0[0]),.doutb(w_n198_0[1]),.din(n198));
	jspl3 jspl3_w_n199_0(.douta(w_n199_0[0]),.doutb(w_n199_0[1]),.doutc(w_n199_0[2]),.din(n199));
	jspl jspl_w_n201_0(.douta(w_n201_0[0]),.doutb(w_n201_0[1]),.din(n201));
	jspl jspl_w_n204_0(.douta(w_n204_0[0]),.doutb(w_n204_0[1]),.din(n204));
	jspl jspl_w_n206_0(.douta(w_n206_0[0]),.doutb(w_n206_0[1]),.din(n206));
	jspl jspl_w_n208_0(.douta(w_n208_0[0]),.doutb(w_n208_0[1]),.din(n208));
	jspl jspl_w_n210_0(.douta(w_n210_0[0]),.doutb(w_n210_0[1]),.din(n210));
	jspl jspl_w_n211_0(.douta(w_n211_0[0]),.doutb(w_n211_0[1]),.din(n211));
	jspl3 jspl3_w_n214_0(.douta(w_n214_0[0]),.doutb(w_n214_0[1]),.doutc(w_n214_0[2]),.din(n214));
	jspl3 jspl3_w_n216_0(.douta(w_n216_0[0]),.doutb(w_n216_0[1]),.doutc(w_n216_0[2]),.din(n216));
	jspl jspl_w_n216_1(.douta(w_n216_1[0]),.doutb(w_n216_1[1]),.din(w_n216_0[0]));
	jspl jspl_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.din(n217));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.din(n218));
	jspl jspl_w_n220_0(.douta(w_n220_0[0]),.doutb(w_n220_0[1]),.din(n220));
	jspl jspl_w_n224_0(.douta(w_n224_0[0]),.doutb(w_n224_0[1]),.din(n224));
	jspl jspl_w_n226_0(.douta(w_n226_0[0]),.doutb(w_n226_0[1]),.din(n226));
	jspl3 jspl3_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.doutc(w_n242_0[2]),.din(n242));
	jspl3 jspl3_w_n242_1(.douta(w_n242_1[0]),.doutb(w_n242_1[1]),.doutc(w_n242_1[2]),.din(w_n242_0[0]));
	jspl3 jspl3_w_n242_2(.douta(w_n242_2[0]),.doutb(w_n242_2[1]),.doutc(w_n242_2[2]),.din(w_n242_0[1]));
	jspl jspl_w_n243_0(.douta(w_n243_0[0]),.doutb(w_n243_0[1]),.din(n243));
	jspl jspl_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.din(n249));
	jspl3 jspl3_w_n258_0(.douta(w_n258_0[0]),.doutb(w_n258_0[1]),.doutc(w_n258_0[2]),.din(n258));
	jspl3 jspl3_w_n265_0(.douta(w_n265_0[0]),.doutb(w_n265_0[1]),.doutc(w_n265_0[2]),.din(n265));
	jspl3 jspl3_w_n265_1(.douta(w_n265_1[0]),.doutb(w_n265_1[1]),.doutc(w_n265_1[2]),.din(w_n265_0[0]));
	jspl jspl_w_n265_2(.douta(w_n265_2[0]),.doutb(w_n265_2[1]),.din(w_n265_0[1]));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_n274_0[1]),.din(n274));
	jspl3 jspl3_w_n278_0(.douta(w_n278_0[0]),.doutb(w_n278_0[1]),.doutc(w_n278_0[2]),.din(n278));
	jspl jspl_w_n279_0(.douta(w_n279_0[0]),.doutb(w_n279_0[1]),.din(n279));
	jspl jspl_w_n280_0(.douta(w_n280_0[0]),.doutb(w_n280_0[1]),.din(n280));
	jspl3 jspl3_w_n282_0(.douta(w_n282_0[0]),.doutb(w_n282_0[1]),.doutc(w_n282_0[2]),.din(n282));
	jspl jspl_w_n282_1(.douta(w_n282_1[0]),.doutb(w_n282_1[1]),.din(w_n282_0[0]));
	jspl jspl_w_n286_0(.douta(w_n286_0[0]),.doutb(w_n286_0[1]),.din(n286));
	jspl3 jspl3_w_n287_0(.douta(w_n287_0[0]),.doutb(w_n287_0[1]),.doutc(w_n287_0[2]),.din(n287));
	jspl jspl_w_n287_1(.douta(w_n287_1[0]),.doutb(w_n287_1[1]),.din(w_n287_0[0]));
	jspl jspl_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.din(n288));
	jspl3 jspl3_w_n291_0(.douta(w_n291_0[0]),.doutb(w_n291_0[1]),.doutc(w_n291_0[2]),.din(n291));
	jspl jspl_w_n291_1(.douta(w_n291_1[0]),.doutb(w_n291_1[1]),.din(w_n291_0[0]));
	jspl jspl_w_n292_0(.douta(w_n292_0[0]),.doutb(w_n292_0[1]),.din(n292));
	jspl jspl_w_n293_0(.douta(w_n293_0[0]),.doutb(w_n293_0[1]),.din(n293));
	jspl jspl_w_n294_0(.douta(w_n294_0[0]),.doutb(w_n294_0[1]),.din(n294));
	jspl jspl_w_n297_0(.douta(w_n297_0[0]),.doutb(w_n297_0[1]),.din(n297));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.din(n303));
	jspl3 jspl3_w_n307_0(.douta(w_n307_0[0]),.doutb(w_n307_0[1]),.doutc(w_n307_0[2]),.din(n307));
	jspl jspl_w_n313_0(.douta(w_n313_0[0]),.doutb(w_n313_0[1]),.din(n313));
	jspl3 jspl3_w_n316_0(.douta(w_n316_0[0]),.doutb(w_n316_0[1]),.doutc(w_n316_0[2]),.din(n316));
	jspl3 jspl3_w_n317_0(.douta(w_n317_0[0]),.doutb(w_n317_0[1]),.doutc(w_n317_0[2]),.din(n317));
	jspl jspl_w_n322_0(.douta(w_n322_0[0]),.doutb(w_n322_0[1]),.din(n322));
	jspl jspl_w_n323_0(.douta(w_n323_0[0]),.doutb(w_n323_0[1]),.din(n323));
	jspl jspl_w_n327_0(.douta(w_n327_0[0]),.doutb(w_n327_0[1]),.din(n327));
	jspl jspl_w_n329_0(.douta(w_n329_0[0]),.doutb(w_n329_0[1]),.din(n329));
	jspl jspl_w_n341_0(.douta(w_n341_0[0]),.doutb(w_n341_0[1]),.din(n341));
	jdff dff_B_mcx8HXjZ1_0(.din(n263),.dout(w_dff_B_mcx8HXjZ1_0),.clk(gclk));
	jdff dff_B_bFOZa4sH6_0(.din(w_dff_B_mcx8HXjZ1_0),.dout(w_dff_B_bFOZa4sH6_0),.clk(gclk));
	jdff dff_B_grBeq9j94_0(.din(w_dff_B_bFOZa4sH6_0),.dout(w_dff_B_grBeq9j94_0),.clk(gclk));
	jdff dff_B_9UFfzvlu2_0(.din(w_dff_B_grBeq9j94_0),.dout(w_dff_B_9UFfzvlu2_0),.clk(gclk));
	jdff dff_B_MLTY3rqi9_0(.din(w_dff_B_9UFfzvlu2_0),.dout(w_dff_B_MLTY3rqi9_0),.clk(gclk));
	jdff dff_B_aWYS1ZOy1_1(.din(n276),.dout(w_dff_B_aWYS1ZOy1_1),.clk(gclk));
	jdff dff_B_52GnKZf39_1(.din(n356),.dout(w_dff_B_52GnKZf39_1),.clk(gclk));
	jdff dff_B_PpmdxMA92_1(.din(w_dff_B_52GnKZf39_1),.dout(w_dff_B_PpmdxMA92_1),.clk(gclk));
	jdff dff_B_U0PxIqWc0_1(.din(w_dff_B_PpmdxMA92_1),.dout(w_dff_B_U0PxIqWc0_1),.clk(gclk));
	jdff dff_B_XWZSrCpu1_1(.din(w_dff_B_U0PxIqWc0_1),.dout(w_dff_B_XWZSrCpu1_1),.clk(gclk));
	jdff dff_B_AVuulWGR7_1(.din(w_dff_B_XWZSrCpu1_1),.dout(w_dff_B_AVuulWGR7_1),.clk(gclk));
	jdff dff_B_qe0ME2T25_1(.din(w_dff_B_AVuulWGR7_1),.dout(w_dff_B_qe0ME2T25_1),.clk(gclk));
	jdff dff_B_QKks3Nyo9_1(.din(w_dff_B_qe0ME2T25_1),.dout(w_dff_B_QKks3Nyo9_1),.clk(gclk));
	jdff dff_B_6UoEHvV06_1(.din(w_dff_B_QKks3Nyo9_1),.dout(w_dff_B_6UoEHvV06_1),.clk(gclk));
	jdff dff_B_T0nU5WW41_1(.din(w_dff_B_6UoEHvV06_1),.dout(w_dff_B_T0nU5WW41_1),.clk(gclk));
	jdff dff_B_4Wvdo2MD6_1(.din(w_dff_B_T0nU5WW41_1),.dout(w_dff_B_4Wvdo2MD6_1),.clk(gclk));
	jdff dff_B_r8lSCO022_1(.din(w_dff_B_4Wvdo2MD6_1),.dout(w_dff_B_r8lSCO022_1),.clk(gclk));
	jdff dff_B_k0Z0wKK09_1(.din(w_dff_B_r8lSCO022_1),.dout(w_dff_B_k0Z0wKK09_1),.clk(gclk));
	jdff dff_B_7VXxI4l23_0(.din(n367),.dout(w_dff_B_7VXxI4l23_0),.clk(gclk));
	jdff dff_B_i7PbQM5S0_0(.din(w_dff_B_7VXxI4l23_0),.dout(w_dff_B_i7PbQM5S0_0),.clk(gclk));
	jdff dff_B_juNbU65h3_0(.din(w_dff_B_i7PbQM5S0_0),.dout(w_dff_B_juNbU65h3_0),.clk(gclk));
	jdff dff_B_ZqgcQENp8_0(.din(w_dff_B_juNbU65h3_0),.dout(w_dff_B_ZqgcQENp8_0),.clk(gclk));
	jdff dff_B_sNEiNVkP9_0(.din(w_dff_B_ZqgcQENp8_0),.dout(w_dff_B_sNEiNVkP9_0),.clk(gclk));
	jdff dff_B_uaPcn3RO5_0(.din(w_dff_B_sNEiNVkP9_0),.dout(w_dff_B_uaPcn3RO5_0),.clk(gclk));
	jdff dff_B_OQjizde24_0(.din(w_dff_B_uaPcn3RO5_0),.dout(w_dff_B_OQjizde24_0),.clk(gclk));
	jdff dff_B_tV1wbGDu1_0(.din(w_dff_B_OQjizde24_0),.dout(w_dff_B_tV1wbGDu1_0),.clk(gclk));
	jdff dff_B_ObDKHwKj7_0(.din(w_dff_B_tV1wbGDu1_0),.dout(w_dff_B_ObDKHwKj7_0),.clk(gclk));
	jdff dff_B_HoaeaW9F5_0(.din(w_dff_B_ObDKHwKj7_0),.dout(w_dff_B_HoaeaW9F5_0),.clk(gclk));
	jdff dff_B_VZ1fJwtq4_0(.din(w_dff_B_HoaeaW9F5_0),.dout(w_dff_B_VZ1fJwtq4_0),.clk(gclk));
	jdff dff_B_wHVSvMI70_0(.din(w_dff_B_VZ1fJwtq4_0),.dout(w_dff_B_wHVSvMI70_0),.clk(gclk));
	jdff dff_A_oVsTq72R1_2(.dout(w_dff_A_0C9ObIdz0_0),.din(w_dff_A_oVsTq72R1_2),.clk(gclk));
	jdff dff_A_0C9ObIdz0_0(.dout(w_dff_A_VTtHXf1F2_0),.din(w_dff_A_0C9ObIdz0_0),.clk(gclk));
	jdff dff_A_VTtHXf1F2_0(.dout(w_dff_A_pXh7WgNI4_0),.din(w_dff_A_VTtHXf1F2_0),.clk(gclk));
	jdff dff_A_pXh7WgNI4_0(.dout(w_dff_A_v4hP8LCg6_0),.din(w_dff_A_pXh7WgNI4_0),.clk(gclk));
	jdff dff_A_v4hP8LCg6_0(.dout(w_dff_A_KvxqVpnN9_0),.din(w_dff_A_v4hP8LCg6_0),.clk(gclk));
	jdff dff_A_KvxqVpnN9_0(.dout(w_dff_A_Th9AYmzj6_0),.din(w_dff_A_KvxqVpnN9_0),.clk(gclk));
	jdff dff_A_Th9AYmzj6_0(.dout(w_dff_A_aUtnlEKl1_0),.din(w_dff_A_Th9AYmzj6_0),.clk(gclk));
	jdff dff_A_aUtnlEKl1_0(.dout(G3),.din(w_dff_A_aUtnlEKl1_0),.clk(gclk));
	jdff dff_A_l0poYgO75_2(.dout(w_dff_A_Ijlgz3FN8_0),.din(w_dff_A_l0poYgO75_2),.clk(gclk));
	jdff dff_A_Ijlgz3FN8_0(.dout(w_dff_A_HS7wqKna6_0),.din(w_dff_A_Ijlgz3FN8_0),.clk(gclk));
	jdff dff_A_HS7wqKna6_0(.dout(w_dff_A_cOyKGyYO3_0),.din(w_dff_A_HS7wqKna6_0),.clk(gclk));
	jdff dff_A_cOyKGyYO3_0(.dout(w_dff_A_HYXdyIgm0_0),.din(w_dff_A_cOyKGyYO3_0),.clk(gclk));
	jdff dff_A_HYXdyIgm0_0(.dout(w_dff_A_1u6WuHLL3_0),.din(w_dff_A_HYXdyIgm0_0),.clk(gclk));
	jdff dff_A_1u6WuHLL3_0(.dout(w_dff_A_J8vR6Aft9_0),.din(w_dff_A_1u6WuHLL3_0),.clk(gclk));
	jdff dff_A_J8vR6Aft9_0(.dout(w_dff_A_LMEzXytF4_0),.din(w_dff_A_J8vR6Aft9_0),.clk(gclk));
	jdff dff_A_LMEzXytF4_0(.dout(G6),.din(w_dff_A_LMEzXytF4_0),.clk(gclk));
	jdff dff_A_YW8W7tRx6_2(.dout(w_dff_A_7jFk8CV00_0),.din(w_dff_A_YW8W7tRx6_2),.clk(gclk));
	jdff dff_A_7jFk8CV00_0(.dout(w_dff_A_yqAu8yh37_0),.din(w_dff_A_7jFk8CV00_0),.clk(gclk));
	jdff dff_A_yqAu8yh37_0(.dout(w_dff_A_2obB2PTB9_0),.din(w_dff_A_yqAu8yh37_0),.clk(gclk));
	jdff dff_A_2obB2PTB9_0(.dout(w_dff_A_CcPjPksI8_0),.din(w_dff_A_2obB2PTB9_0),.clk(gclk));
	jdff dff_A_CcPjPksI8_0(.dout(w_dff_A_YVQrcD270_0),.din(w_dff_A_CcPjPksI8_0),.clk(gclk));
	jdff dff_A_YVQrcD270_0(.dout(w_dff_A_dH36MvzL2_0),.din(w_dff_A_YVQrcD270_0),.clk(gclk));
	jdff dff_A_dH36MvzL2_0(.dout(w_dff_A_LhoicajQ8_0),.din(w_dff_A_dH36MvzL2_0),.clk(gclk));
	jdff dff_A_LhoicajQ8_0(.dout(G9),.din(w_dff_A_LhoicajQ8_0),.clk(gclk));
	jdff dff_A_gGm2HDNQ2_2(.dout(w_dff_A_b5T9GjKi0_0),.din(w_dff_A_gGm2HDNQ2_2),.clk(gclk));
	jdff dff_A_b5T9GjKi0_0(.dout(w_dff_A_Sk7t9mV98_0),.din(w_dff_A_b5T9GjKi0_0),.clk(gclk));
	jdff dff_A_Sk7t9mV98_0(.dout(w_dff_A_lDUlwOQB3_0),.din(w_dff_A_Sk7t9mV98_0),.clk(gclk));
	jdff dff_A_lDUlwOQB3_0(.dout(w_dff_A_JuJnZyNl5_0),.din(w_dff_A_lDUlwOQB3_0),.clk(gclk));
	jdff dff_A_JuJnZyNl5_0(.dout(w_dff_A_b46OLkIx0_0),.din(w_dff_A_JuJnZyNl5_0),.clk(gclk));
	jdff dff_A_b46OLkIx0_0(.dout(w_dff_A_TRlfbQ617_0),.din(w_dff_A_b46OLkIx0_0),.clk(gclk));
	jdff dff_A_TRlfbQ617_0(.dout(w_dff_A_TctbjcZR3_0),.din(w_dff_A_TRlfbQ617_0),.clk(gclk));
	jdff dff_A_TctbjcZR3_0(.dout(G12),.din(w_dff_A_TctbjcZR3_0),.clk(gclk));
	jdff dff_A_Vp6nTiae6_2(.dout(w_dff_A_24bQa3Bi5_0),.din(w_dff_A_Vp6nTiae6_2),.clk(gclk));
	jdff dff_A_24bQa3Bi5_0(.dout(w_dff_A_xrJX33Sg2_0),.din(w_dff_A_24bQa3Bi5_0),.clk(gclk));
	jdff dff_A_xrJX33Sg2_0(.dout(w_dff_A_sEvO2muf3_0),.din(w_dff_A_xrJX33Sg2_0),.clk(gclk));
	jdff dff_A_sEvO2muf3_0(.dout(w_dff_A_6J0mkjEY9_0),.din(w_dff_A_sEvO2muf3_0),.clk(gclk));
	jdff dff_A_6J0mkjEY9_0(.dout(w_dff_A_JJVwsxEo3_0),.din(w_dff_A_6J0mkjEY9_0),.clk(gclk));
	jdff dff_A_JJVwsxEo3_0(.dout(w_dff_A_WFsMxitT1_0),.din(w_dff_A_JJVwsxEo3_0),.clk(gclk));
	jdff dff_A_WFsMxitT1_0(.dout(w_dff_A_yeCunKXX4_0),.din(w_dff_A_WFsMxitT1_0),.clk(gclk));
	jdff dff_A_yeCunKXX4_0(.dout(G30),.din(w_dff_A_yeCunKXX4_0),.clk(gclk));
	jdff dff_A_jKXqwK7t1_2(.dout(w_dff_A_sYAVy6pF3_0),.din(w_dff_A_jKXqwK7t1_2),.clk(gclk));
	jdff dff_A_sYAVy6pF3_0(.dout(w_dff_A_KFl9pbzH7_0),.din(w_dff_A_sYAVy6pF3_0),.clk(gclk));
	jdff dff_A_KFl9pbzH7_0(.dout(w_dff_A_IFb2x9iA9_0),.din(w_dff_A_KFl9pbzH7_0),.clk(gclk));
	jdff dff_A_IFb2x9iA9_0(.dout(w_dff_A_PjYxAS1v3_0),.din(w_dff_A_IFb2x9iA9_0),.clk(gclk));
	jdff dff_A_PjYxAS1v3_0(.dout(w_dff_A_tN3SXOc79_0),.din(w_dff_A_PjYxAS1v3_0),.clk(gclk));
	jdff dff_A_tN3SXOc79_0(.dout(w_dff_A_MAPOkg9G3_0),.din(w_dff_A_tN3SXOc79_0),.clk(gclk));
	jdff dff_A_MAPOkg9G3_0(.dout(w_dff_A_GuQUmgZ43_0),.din(w_dff_A_MAPOkg9G3_0),.clk(gclk));
	jdff dff_A_GuQUmgZ43_0(.dout(G45),.din(w_dff_A_GuQUmgZ43_0),.clk(gclk));
	jdff dff_A_xLZeIvHB1_2(.dout(w_dff_A_n7FfThNw2_0),.din(w_dff_A_xLZeIvHB1_2),.clk(gclk));
	jdff dff_A_n7FfThNw2_0(.dout(w_dff_A_rv8UR1Ui2_0),.din(w_dff_A_n7FfThNw2_0),.clk(gclk));
	jdff dff_A_rv8UR1Ui2_0(.dout(w_dff_A_cTpxm0Z59_0),.din(w_dff_A_rv8UR1Ui2_0),.clk(gclk));
	jdff dff_A_cTpxm0Z59_0(.dout(w_dff_A_4lzkzswJ4_0),.din(w_dff_A_cTpxm0Z59_0),.clk(gclk));
	jdff dff_A_4lzkzswJ4_0(.dout(w_dff_A_g8wPsrTs2_0),.din(w_dff_A_4lzkzswJ4_0),.clk(gclk));
	jdff dff_A_g8wPsrTs2_0(.dout(w_dff_A_DKz2k2r71_0),.din(w_dff_A_g8wPsrTs2_0),.clk(gclk));
	jdff dff_A_DKz2k2r71_0(.dout(w_dff_A_UInU27ge7_0),.din(w_dff_A_DKz2k2r71_0),.clk(gclk));
	jdff dff_A_UInU27ge7_0(.dout(G48),.din(w_dff_A_UInU27ge7_0),.clk(gclk));
	jdff dff_A_iwFOWnuB4_2(.dout(w_dff_A_barZ3sRj6_0),.din(w_dff_A_iwFOWnuB4_2),.clk(gclk));
	jdff dff_A_barZ3sRj6_0(.dout(w_dff_A_CqSBO5hc0_0),.din(w_dff_A_barZ3sRj6_0),.clk(gclk));
	jdff dff_A_CqSBO5hc0_0(.dout(w_dff_A_LUHHYikK1_0),.din(w_dff_A_CqSBO5hc0_0),.clk(gclk));
	jdff dff_A_LUHHYikK1_0(.dout(w_dff_A_PwPyty8z0_0),.din(w_dff_A_LUHHYikK1_0),.clk(gclk));
	jdff dff_A_PwPyty8z0_0(.dout(w_dff_A_P54LFzTU8_0),.din(w_dff_A_PwPyty8z0_0),.clk(gclk));
	jdff dff_A_P54LFzTU8_0(.dout(w_dff_A_qdV3DD4Y6_0),.din(w_dff_A_P54LFzTU8_0),.clk(gclk));
	jdff dff_A_qdV3DD4Y6_0(.dout(w_dff_A_uAX3FQTh3_0),.din(w_dff_A_qdV3DD4Y6_0),.clk(gclk));
	jdff dff_A_uAX3FQTh3_0(.dout(G15),.din(w_dff_A_uAX3FQTh3_0),.clk(gclk));
	jdff dff_A_E73ITE3P9_2(.dout(w_dff_A_ySGCkCjc0_0),.din(w_dff_A_E73ITE3P9_2),.clk(gclk));
	jdff dff_A_ySGCkCjc0_0(.dout(w_dff_A_xyA1laYS8_0),.din(w_dff_A_ySGCkCjc0_0),.clk(gclk));
	jdff dff_A_xyA1laYS8_0(.dout(w_dff_A_FS7zwQeQ4_0),.din(w_dff_A_xyA1laYS8_0),.clk(gclk));
	jdff dff_A_FS7zwQeQ4_0(.dout(w_dff_A_qtDWqYxR9_0),.din(w_dff_A_FS7zwQeQ4_0),.clk(gclk));
	jdff dff_A_qtDWqYxR9_0(.dout(w_dff_A_PqOrVhch4_0),.din(w_dff_A_qtDWqYxR9_0),.clk(gclk));
	jdff dff_A_PqOrVhch4_0(.dout(w_dff_A_x8C7AKdU5_0),.din(w_dff_A_PqOrVhch4_0),.clk(gclk));
	jdff dff_A_x8C7AKdU5_0(.dout(w_dff_A_JSgVYWW44_0),.din(w_dff_A_x8C7AKdU5_0),.clk(gclk));
	jdff dff_A_JSgVYWW44_0(.dout(G18),.din(w_dff_A_JSgVYWW44_0),.clk(gclk));
	jdff dff_A_XOYZZE3e4_2(.dout(w_dff_A_63W526Nc5_0),.din(w_dff_A_XOYZZE3e4_2),.clk(gclk));
	jdff dff_A_63W526Nc5_0(.dout(w_dff_A_XTsxj5Mo1_0),.din(w_dff_A_63W526Nc5_0),.clk(gclk));
	jdff dff_A_XTsxj5Mo1_0(.dout(w_dff_A_fYeEoUwM2_0),.din(w_dff_A_XTsxj5Mo1_0),.clk(gclk));
	jdff dff_A_fYeEoUwM2_0(.dout(w_dff_A_SBzPjrmn4_0),.din(w_dff_A_fYeEoUwM2_0),.clk(gclk));
	jdff dff_A_SBzPjrmn4_0(.dout(w_dff_A_tgCO6byC4_0),.din(w_dff_A_SBzPjrmn4_0),.clk(gclk));
	jdff dff_A_tgCO6byC4_0(.dout(w_dff_A_ptAm8GdO5_0),.din(w_dff_A_tgCO6byC4_0),.clk(gclk));
	jdff dff_A_ptAm8GdO5_0(.dout(w_dff_A_Eu3Pq5975_0),.din(w_dff_A_ptAm8GdO5_0),.clk(gclk));
	jdff dff_A_Eu3Pq5975_0(.dout(G21),.din(w_dff_A_Eu3Pq5975_0),.clk(gclk));
	jdff dff_A_5zLbCwG53_2(.dout(w_dff_A_LweQl56s5_0),.din(w_dff_A_5zLbCwG53_2),.clk(gclk));
	jdff dff_A_LweQl56s5_0(.dout(w_dff_A_cgCOdFSo7_0),.din(w_dff_A_LweQl56s5_0),.clk(gclk));
	jdff dff_A_cgCOdFSo7_0(.dout(w_dff_A_s08SeP1K0_0),.din(w_dff_A_cgCOdFSo7_0),.clk(gclk));
	jdff dff_A_s08SeP1K0_0(.dout(w_dff_A_sUGmBRsO0_0),.din(w_dff_A_s08SeP1K0_0),.clk(gclk));
	jdff dff_A_sUGmBRsO0_0(.dout(w_dff_A_pnuinHEP4_0),.din(w_dff_A_sUGmBRsO0_0),.clk(gclk));
	jdff dff_A_pnuinHEP4_0(.dout(w_dff_A_sUOKxKkw6_0),.din(w_dff_A_pnuinHEP4_0),.clk(gclk));
	jdff dff_A_sUOKxKkw6_0(.dout(G24),.din(w_dff_A_sUOKxKkw6_0),.clk(gclk));
	jdff dff_A_PMMyqFGP2_2(.dout(w_dff_A_e7VnHSKm1_0),.din(w_dff_A_PMMyqFGP2_2),.clk(gclk));
	jdff dff_A_e7VnHSKm1_0(.dout(w_dff_A_7OuwsZWL3_0),.din(w_dff_A_e7VnHSKm1_0),.clk(gclk));
	jdff dff_A_7OuwsZWL3_0(.dout(w_dff_A_MHfphiOd2_0),.din(w_dff_A_7OuwsZWL3_0),.clk(gclk));
	jdff dff_A_MHfphiOd2_0(.dout(w_dff_A_SBe3M3F32_0),.din(w_dff_A_MHfphiOd2_0),.clk(gclk));
	jdff dff_A_SBe3M3F32_0(.dout(w_dff_A_FkrH5WKV0_0),.din(w_dff_A_SBe3M3F32_0),.clk(gclk));
	jdff dff_A_FkrH5WKV0_0(.dout(w_dff_A_Cmj6XXNM7_0),.din(w_dff_A_FkrH5WKV0_0),.clk(gclk));
	jdff dff_A_Cmj6XXNM7_0(.dout(w_dff_A_7SDL1qwd8_0),.din(w_dff_A_Cmj6XXNM7_0),.clk(gclk));
	jdff dff_A_7SDL1qwd8_0(.dout(G27),.din(w_dff_A_7SDL1qwd8_0),.clk(gclk));
	jdff dff_A_8Vc8w38d7_2(.dout(w_dff_A_gHFDlBjI5_0),.din(w_dff_A_8Vc8w38d7_2),.clk(gclk));
	jdff dff_A_gHFDlBjI5_0(.dout(w_dff_A_prqr8yZ23_0),.din(w_dff_A_gHFDlBjI5_0),.clk(gclk));
	jdff dff_A_prqr8yZ23_0(.dout(w_dff_A_BvpQ5XvI6_0),.din(w_dff_A_prqr8yZ23_0),.clk(gclk));
	jdff dff_A_BvpQ5XvI6_0(.dout(w_dff_A_XFaziCNF0_0),.din(w_dff_A_BvpQ5XvI6_0),.clk(gclk));
	jdff dff_A_XFaziCNF0_0(.dout(w_dff_A_sDqZu0UT6_0),.din(w_dff_A_XFaziCNF0_0),.clk(gclk));
	jdff dff_A_sDqZu0UT6_0(.dout(w_dff_A_pkaiTCoc0_0),.din(w_dff_A_sDqZu0UT6_0),.clk(gclk));
	jdff dff_A_pkaiTCoc0_0(.dout(w_dff_A_rBEg7uQw7_0),.din(w_dff_A_pkaiTCoc0_0),.clk(gclk));
	jdff dff_A_rBEg7uQw7_0(.dout(G33),.din(w_dff_A_rBEg7uQw7_0),.clk(gclk));
	jdff dff_A_KqOJDCII5_2(.dout(w_dff_A_BJtD2o3t5_0),.din(w_dff_A_KqOJDCII5_2),.clk(gclk));
	jdff dff_A_BJtD2o3t5_0(.dout(w_dff_A_fsUBMFRg8_0),.din(w_dff_A_BJtD2o3t5_0),.clk(gclk));
	jdff dff_A_fsUBMFRg8_0(.dout(w_dff_A_U81QikaM4_0),.din(w_dff_A_fsUBMFRg8_0),.clk(gclk));
	jdff dff_A_U81QikaM4_0(.dout(w_dff_A_enSP1Mit9_0),.din(w_dff_A_U81QikaM4_0),.clk(gclk));
	jdff dff_A_enSP1Mit9_0(.dout(w_dff_A_8ZAhcqkK2_0),.din(w_dff_A_enSP1Mit9_0),.clk(gclk));
	jdff dff_A_8ZAhcqkK2_0(.dout(w_dff_A_b2nk0cNJ0_0),.din(w_dff_A_8ZAhcqkK2_0),.clk(gclk));
	jdff dff_A_b2nk0cNJ0_0(.dout(w_dff_A_v5lJGdRk4_0),.din(w_dff_A_b2nk0cNJ0_0),.clk(gclk));
	jdff dff_A_v5lJGdRk4_0(.dout(G36),.din(w_dff_A_v5lJGdRk4_0),.clk(gclk));
	jdff dff_A_K41iITcE1_2(.dout(w_dff_A_V0GzjCRJ0_0),.din(w_dff_A_K41iITcE1_2),.clk(gclk));
	jdff dff_A_V0GzjCRJ0_0(.dout(w_dff_A_nNodPbMX1_0),.din(w_dff_A_V0GzjCRJ0_0),.clk(gclk));
	jdff dff_A_nNodPbMX1_0(.dout(w_dff_A_JlUFRsSp1_0),.din(w_dff_A_nNodPbMX1_0),.clk(gclk));
	jdff dff_A_JlUFRsSp1_0(.dout(w_dff_A_5zrBvXGJ2_0),.din(w_dff_A_JlUFRsSp1_0),.clk(gclk));
	jdff dff_A_5zrBvXGJ2_0(.dout(w_dff_A_ldIo83AH2_0),.din(w_dff_A_5zrBvXGJ2_0),.clk(gclk));
	jdff dff_A_ldIo83AH2_0(.dout(w_dff_A_qya9AF8Z2_0),.din(w_dff_A_ldIo83AH2_0),.clk(gclk));
	jdff dff_A_qya9AF8Z2_0(.dout(w_dff_A_6eyP3IdB3_0),.din(w_dff_A_qya9AF8Z2_0),.clk(gclk));
	jdff dff_A_6eyP3IdB3_0(.dout(G39),.din(w_dff_A_6eyP3IdB3_0),.clk(gclk));
	jdff dff_A_RLsCUGFu5_2(.dout(w_dff_A_zXDiMy8I2_0),.din(w_dff_A_RLsCUGFu5_2),.clk(gclk));
	jdff dff_A_zXDiMy8I2_0(.dout(w_dff_A_TlwsZlB46_0),.din(w_dff_A_zXDiMy8I2_0),.clk(gclk));
	jdff dff_A_TlwsZlB46_0(.dout(w_dff_A_yzDMr6002_0),.din(w_dff_A_TlwsZlB46_0),.clk(gclk));
	jdff dff_A_yzDMr6002_0(.dout(w_dff_A_bhmUH3KQ9_0),.din(w_dff_A_yzDMr6002_0),.clk(gclk));
	jdff dff_A_bhmUH3KQ9_0(.dout(w_dff_A_kXM7QATo9_0),.din(w_dff_A_bhmUH3KQ9_0),.clk(gclk));
	jdff dff_A_kXM7QATo9_0(.dout(w_dff_A_zVpqac9g1_0),.din(w_dff_A_kXM7QATo9_0),.clk(gclk));
	jdff dff_A_zVpqac9g1_0(.dout(w_dff_A_d36VfAlB3_0),.din(w_dff_A_zVpqac9g1_0),.clk(gclk));
	jdff dff_A_d36VfAlB3_0(.dout(G42),.din(w_dff_A_d36VfAlB3_0),.clk(gclk));
	jdff dff_A_OZrJidH88_2(.dout(G75),.din(w_dff_A_OZrJidH88_2),.clk(gclk));
	jdff dff_A_rJpE2Sql2_2(.dout(w_dff_A_6qmy4NLb6_0),.din(w_dff_A_rJpE2Sql2_2),.clk(gclk));
	jdff dff_A_6qmy4NLb6_0(.dout(G69),.din(w_dff_A_6qmy4NLb6_0),.clk(gclk));
	jdff dff_A_4zosqtN80_2(.dout(w_dff_A_Etogts5K7_0),.din(w_dff_A_4zosqtN80_2),.clk(gclk));
	jdff dff_A_Etogts5K7_0(.dout(G72),.din(w_dff_A_Etogts5K7_0),.clk(gclk));
	jdff dff_A_H21VoaHU2_2(.dout(G57),.din(w_dff_A_H21VoaHU2_2),.clk(gclk));
endmodule

