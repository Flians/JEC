/*

c499:
	jxor: 120
	jspl: 54
	jspl3: 64
	jnot: 8
	jdff: 477
	jand: 69
	jor: 2

Summary:
	jxor: 120
	jspl: 54
	jspl3: 64
	jnot: 8
	jdff: 477
	jand: 69
	jor: 2
*/

module c499(gclk, Gid0, Gid1, Gid2, Gid3, Gid4, Gid5, Gid6, Gid7, Gid8, Gid9, Gid10, Gid11, Gid12, Gid13, Gid14, Gid15, Gid16, Gid17, Gid18, Gid19, Gid20, Gid21, Gid22, Gid23, Gid24, Gid25, Gid26, Gid27, Gid28, Gid29, Gid30, Gid31, Gic0, Gic1, Gic2, Gic3, Gic4, Gic5, Gic6, Gic7, Gr, God0, God1, God2, God3, God4, God5, God6, God7, God8, God9, God10, God11, God12, God13, God14, God15, God16, God17, God18, God19, God20, God21, God22, God23, God24, God25, God26, God27, God28, God29, God30, God31);
	input gclk;
	input Gid0;
	input Gid1;
	input Gid2;
	input Gid3;
	input Gid4;
	input Gid5;
	input Gid6;
	input Gid7;
	input Gid8;
	input Gid9;
	input Gid10;
	input Gid11;
	input Gid12;
	input Gid13;
	input Gid14;
	input Gid15;
	input Gid16;
	input Gid17;
	input Gid18;
	input Gid19;
	input Gid20;
	input Gid21;
	input Gid22;
	input Gid23;
	input Gid24;
	input Gid25;
	input Gid26;
	input Gid27;
	input Gid28;
	input Gid29;
	input Gid30;
	input Gid31;
	input Gic0;
	input Gic1;
	input Gic2;
	input Gic3;
	input Gic4;
	input Gic5;
	input Gic6;
	input Gic7;
	input Gr;
	output God0;
	output God1;
	output God2;
	output God3;
	output God4;
	output God5;
	output God6;
	output God7;
	output God8;
	output God9;
	output God10;
	output God11;
	output God12;
	output God13;
	output God14;
	output God15;
	output God16;
	output God17;
	output God18;
	output God19;
	output God20;
	output God21;
	output God22;
	output God23;
	output God24;
	output God25;
	output God26;
	output God27;
	output God28;
	output God29;
	output God30;
	output God31;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n180;
	wire n182;
	wire n184;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n194;
	wire n196;
	wire n198;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n208;
	wire n210;
	wire n212;
	wire n214;
	wire n215;
	wire n217;
	wire n219;
	wire n221;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n236;
	wire n238;
	wire n240;
	wire n242;
	wire n243;
	wire n244;
	wire n246;
	wire n248;
	wire n250;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n257;
	wire n259;
	wire n261;
	wire n263;
	wire n264;
	wire n266;
	wire n268;
	wire n270;
	wire [2:0] w_Gid0_0;
	wire [2:0] w_Gid1_0;
	wire [2:0] w_Gid2_0;
	wire [2:0] w_Gid3_0;
	wire [2:0] w_Gid4_0;
	wire [2:0] w_Gid5_0;
	wire [2:0] w_Gid6_0;
	wire [2:0] w_Gid7_0;
	wire [2:0] w_Gid8_0;
	wire [2:0] w_Gid9_0;
	wire [2:0] w_Gid10_0;
	wire [2:0] w_Gid11_0;
	wire [2:0] w_Gid12_0;
	wire [2:0] w_Gid13_0;
	wire [2:0] w_Gid14_0;
	wire [2:0] w_Gid15_0;
	wire [2:0] w_Gid16_0;
	wire [2:0] w_Gid17_0;
	wire [2:0] w_Gid18_0;
	wire [2:0] w_Gid19_0;
	wire [2:0] w_Gid20_0;
	wire [2:0] w_Gid21_0;
	wire [2:0] w_Gid22_0;
	wire [2:0] w_Gid23_0;
	wire [2:0] w_Gid24_0;
	wire [2:0] w_Gid25_0;
	wire [2:0] w_Gid26_0;
	wire [2:0] w_Gid27_0;
	wire [2:0] w_Gid28_0;
	wire [2:0] w_Gid29_0;
	wire [2:0] w_Gid30_0;
	wire [2:0] w_Gid31_0;
	wire [2:0] w_Gr_0;
	wire [2:0] w_Gr_1;
	wire [2:0] w_Gr_2;
	wire [1:0] w_Gr_3;
	wire [1:0] w_n75_0;
	wire [1:0] w_n76_0;
	wire [1:0] w_n80_0;
	wire [1:0] w_n83_0;
	wire [1:0] w_n84_0;
	wire [2:0] w_n85_0;
	wire [2:0] w_n85_1;
	wire [1:0] w_n85_2;
	wire [1:0] w_n88_0;
	wire [1:0] w_n89_0;
	wire [1:0] w_n94_0;
	wire [1:0] w_n97_0;
	wire [1:0] w_n98_0;
	wire [1:0] w_n99_0;
	wire [1:0] w_n107_0;
	wire [1:0] w_n110_0;
	wire [2:0] w_n112_0;
	wire [2:0] w_n112_1;
	wire [2:0] w_n112_2;
	wire [1:0] w_n113_0;
	wire [1:0] w_n116_0;
	wire [1:0] w_n117_0;
	wire [2:0] w_n121_0;
	wire [2:0] w_n124_0;
	wire [1:0] w_n125_0;
	wire [2:0] w_n126_0;
	wire [2:0] w_n126_1;
	wire [1:0] w_n126_2;
	wire [1:0] w_n128_0;
	wire [1:0] w_n134_0;
	wire [1:0] w_n135_0;
	wire [1:0] w_n136_0;
	wire [1:0] w_n142_0;
	wire [1:0] w_n143_0;
	wire [2:0] w_n147_0;
	wire [2:0] w_n147_1;
	wire [1:0] w_n147_2;
	wire [2:0] w_n149_0;
	wire [2:0] w_n149_1;
	wire [1:0] w_n149_2;
	wire [1:0] w_n153_0;
	wire [1:0] w_n156_0;
	wire [2:0] w_n159_0;
	wire [2:0] w_n166_0;
	wire [2:0] w_n166_1;
	wire [2:0] w_n166_2;
	wire [1:0] w_n169_0;
	wire [1:0] w_n170_0;
	wire [1:0] w_n173_0;
	wire [1:0] w_n174_0;
	wire [1:0] w_n175_0;
	wire [2:0] w_n177_0;
	wire [1:0] w_n177_1;
	wire [2:0] w_n187_0;
	wire [2:0] w_n187_1;
	wire [1:0] w_n187_2;
	wire [1:0] w_n188_0;
	wire [1:0] w_n190_0;
	wire [2:0] w_n191_0;
	wire [1:0] w_n191_1;
	wire [1:0] w_n200_0;
	wire [2:0] w_n202_0;
	wire [2:0] w_n202_1;
	wire [1:0] w_n202_2;
	wire [1:0] w_n203_0;
	wire [2:0] w_n205_0;
	wire [1:0] w_n205_1;
	wire [2:0] w_n214_0;
	wire [1:0] w_n214_1;
	wire [1:0] w_n223_0;
	wire [1:0] w_n231_0;
	wire [1:0] w_n232_0;
	wire [2:0] w_n233_0;
	wire [1:0] w_n233_1;
	wire [1:0] w_n242_0;
	wire [2:0] w_n243_0;
	wire [1:0] w_n243_1;
	wire [1:0] w_n253_0;
	wire [2:0] w_n254_0;
	wire [1:0] w_n254_1;
	wire [2:0] w_n263_0;
	wire [1:0] w_n263_1;
	wire w_dff_A_NMBiPfA08_0;
	wire w_dff_B_i5RHafzQ4_2;
	wire w_dff_B_BlATRo9z6_2;
	wire w_dff_A_XJJO2q9r6_1;
	wire w_dff_B_ovUR52QR4_2;
	wire w_dff_B_9popjFMI6_2;
	wire w_dff_B_VB8GMIr55_2;
	wire w_dff_B_4WY4MvOC7_2;
	wire w_dff_B_zHKyPrEP1_0;
	wire w_dff_A_SWz2spEd1_0;
	wire w_dff_A_rJGPT1mb0_0;
	wire w_dff_A_fXuAndlD2_0;
	wire w_dff_A_P0ku1e5Z3_0;
	wire w_dff_A_oIJUwFqg1_0;
	wire w_dff_A_mkT8y3ij7_0;
	wire w_dff_A_bG008g873_0;
	wire w_dff_A_lQ2q4qAY8_0;
	wire w_dff_A_OJQf32ar2_0;
	wire w_dff_A_vHS6vKCS8_0;
	wire w_dff_A_JeCenFCG2_0;
	wire w_dff_A_0rJHf0kh2_0;
	wire w_dff_A_glL36dua6_0;
	wire w_dff_A_kPJ7yxd81_0;
	wire w_dff_A_fbABUCyq5_0;
	wire w_dff_A_HqOMbToB3_0;
	wire w_dff_A_0pZYsjtK0_0;
	wire w_dff_A_8cGMO4gZ7_0;
	wire w_dff_A_1eqpj8yC3_0;
	wire w_dff_A_ruSJ223S5_0;
	wire w_dff_B_x3t1SBEh7_1;
	wire w_dff_B_0hFeU7G62_1;
	wire w_dff_B_UP2iUJHH5_1;
	wire w_dff_A_SeGZvjhO2_0;
	wire w_dff_A_ioAbq98N2_0;
	wire w_dff_A_w6CKBAb81_0;
	wire w_dff_A_bBbp3GfD5_0;
	wire w_dff_A_KyGKnG4J0_0;
	wire w_dff_B_KaBJ0nU53_2;
	wire w_dff_B_QyfcK6VF0_2;
	wire w_dff_B_dm0QMdOB0_2;
	wire w_dff_B_ZWbj9Uoc7_2;
	wire w_dff_A_OhuAyLz43_0;
	wire w_dff_A_1B1ZXF3c1_0;
	wire w_dff_A_UvrBQeLx0_0;
	wire w_dff_A_F23V6yfT8_0;
	wire w_dff_A_ABa81DUA2_0;
	wire w_dff_B_vwVK4pL53_1;
	wire w_dff_B_cYETG44L4_1;
	wire w_dff_B_SiJKSn8T2_1;
	wire w_dff_A_YVygMPnc2_1;
	wire w_dff_A_tf9Ujzwn5_0;
	wire w_dff_A_VpaXB0Rf4_0;
	wire w_dff_A_DghHOQ6g0_0;
	wire w_dff_A_AKcise4m2_0;
	wire w_dff_A_2B6XvYHh7_0;
	wire w_dff_A_JPw379yx3_0;
	wire w_dff_A_eKtt4Lqq4_2;
	wire w_dff_A_3NFEPZyu6_2;
	wire w_dff_A_cMNxwI0D2_2;
	wire w_dff_A_R0kSpJKS2_2;
	wire w_dff_A_o2C4NKxh7_2;
	wire w_dff_A_PGQM1ifd1_2;
	wire w_dff_A_qTQMxoJR3_0;
	wire w_dff_A_ouv0uQWH6_0;
	wire w_dff_A_IikaIfS06_0;
	wire w_dff_A_nBvOlsvz2_0;
	wire w_dff_A_pbXl2sc08_0;
	wire w_dff_A_ZLfkpWer1_0;
	wire w_dff_A_9JwpWNHu3_0;
	wire w_dff_A_72r887Db9_0;
	wire w_dff_A_f9xfAcPB4_2;
	wire w_dff_A_YTWGeupH2_2;
	wire w_dff_A_Z7YB01u19_2;
	wire w_dff_A_I18bsbrJ5_2;
	wire w_dff_A_YHhTEY4p9_2;
	wire w_dff_A_Dqwi5yCP5_2;
	wire w_dff_B_ywuGzupy7_0;
	wire w_dff_A_gUpsNhdc7_1;
	wire w_dff_A_val0AqY39_0;
	wire w_dff_A_UqUR8uJH8_0;
	wire w_dff_A_na1l1pxG7_0;
	wire w_dff_A_y05OQNLB5_0;
	wire w_dff_A_R84Nkzu12_0;
	wire w_dff_A_PAHZ1fb39_0;
	wire w_dff_A_DvnNR7Gr8_2;
	wire w_dff_A_PaJcP9C26_2;
	wire w_dff_A_BCLd1tN77_2;
	wire w_dff_A_apl5VkCD0_2;
	wire w_dff_A_2CqtsBqC1_2;
	wire w_dff_A_LnCvSuYw3_2;
	wire w_dff_A_EjtYTGZI6_0;
	wire w_dff_A_c6Ggwwcr9_0;
	wire w_dff_A_ubP4lckB7_0;
	wire w_dff_A_OkNIja8V9_0;
	wire w_dff_A_zwdJ1dsv9_0;
	wire w_dff_A_BQgqP7PY5_0;
	wire w_dff_A_nW1BTbHm3_0;
	wire w_dff_A_qzBcH4iu1_0;
	wire w_dff_A_oEJq5Y129_0;
	wire w_dff_A_cP9xoJ6c9_0;
	wire w_dff_A_CZtdIhDC9_2;
	wire w_dff_A_aZRWhOKy2_2;
	wire w_dff_A_ojXkaW671_2;
	wire w_dff_A_AOFrt0zn7_2;
	wire w_dff_A_jsnuzbgw6_2;
	wire w_dff_A_qrpZZJsb1_2;
	wire w_dff_B_aEag40On6_0;
	wire w_dff_A_JFe41pC52_0;
	wire w_dff_A_TpGTez5Y7_0;
	wire w_dff_A_LzW34qYD2_0;
	wire w_dff_A_kjw3uN572_0;
	wire w_dff_A_8d4fuzZb7_0;
	wire w_dff_A_KKZrZLki5_1;
	wire w_dff_A_DwFv3ibl3_0;
	wire w_dff_A_y9kXhS3C8_0;
	wire w_dff_A_lFhZsWmk6_0;
	wire w_dff_A_9qWbDexY4_0;
	wire w_dff_A_MB0ROdsr3_0;
	wire w_dff_A_IqMyPzKM5_0;
	wire w_dff_A_vMPiKgwa6_0;
	wire w_dff_A_AJ1bS1Tf2_0;
	wire w_dff_A_gmCKC0tQ3_0;
	wire w_dff_A_e6qHfjer3_0;
	wire w_dff_A_hCwiAIeo8_0;
	wire w_dff_A_OSZBgw5c7_0;
	wire w_dff_A_MBBxGDym4_0;
	wire w_dff_A_4Vp2CxC63_0;
	wire w_dff_A_sFeDdliz6_0;
	wire w_dff_A_aIeU2GuI8_0;
	wire w_dff_A_VmK0hjed0_0;
	wire w_dff_A_2yHW8bBP8_0;
	wire w_dff_A_Rx7o7aBk2_0;
	wire w_dff_A_xyrjiOJf7_0;
	wire w_dff_A_iR1kW9WG3_0;
	wire w_dff_A_15ngu5GP5_0;
	wire w_dff_A_C9FZG8Ob2_0;
	wire w_dff_A_zapEGAJP3_0;
	wire w_dff_A_zYTxt18W7_0;
	wire w_dff_A_Rav4cdvG2_0;
	wire w_dff_A_EDNiREqN0_0;
	wire w_dff_A_T80GeMZf3_0;
	wire w_dff_A_jVCDhH9e1_0;
	wire w_dff_A_e19BsMgq7_0;
	wire w_dff_A_d9kmoeXH9_0;
	wire w_dff_A_DEuaYAYn5_0;
	wire w_dff_A_otYRCJkc9_0;
	wire w_dff_A_ISGge4cv8_0;
	wire w_dff_A_Izc7Bs5L3_0;
	wire w_dff_A_M5JbCvzC7_0;
	wire w_dff_A_lIWeYeRn9_0;
	wire w_dff_A_9mQzmulA3_0;
	wire w_dff_A_Nw1WuOBJ4_0;
	wire w_dff_A_BbKjK4CH4_0;
	wire w_dff_A_fwCw01320_1;
	wire w_dff_A_WawC5gE02_0;
	wire w_dff_A_XBA1D4Hs8_0;
	wire w_dff_A_abPV91rE8_0;
	wire w_dff_A_uddMyPP02_0;
	wire w_dff_A_2E2xC8s41_0;
	wire w_dff_A_dEpawunY5_0;
	wire w_dff_A_jZY79jdm1_0;
	wire w_dff_A_DqkO5rdd9_0;
	wire w_dff_A_vQT2H2Bo2_0;
	wire w_dff_A_yvg1r0oY8_0;
	wire w_dff_A_M9JpT3z83_0;
	wire w_dff_A_iA9wfDyN9_0;
	wire w_dff_A_PUnlEag12_0;
	wire w_dff_A_nZLuvCrW7_0;
	wire w_dff_A_nawXBPD00_0;
	wire w_dff_A_FNnHyjCW0_0;
	wire w_dff_A_2MM5LQ538_0;
	wire w_dff_A_TG2AqP2S5_0;
	wire w_dff_A_lHCVdao89_0;
	wire w_dff_A_sa4OWoUW2_0;
	wire w_dff_A_At90bml85_0;
	wire w_dff_A_g99eVEKr9_0;
	wire w_dff_A_detPl1vj2_0;
	wire w_dff_A_BrP1Za891_0;
	wire w_dff_A_L1S432cR1_0;
	wire w_dff_A_FYeeoov96_0;
	wire w_dff_A_rJWz5WVA5_0;
	wire w_dff_A_YaCx97Sw6_0;
	wire w_dff_A_HqSsxoLx5_0;
	wire w_dff_A_VnYVtnKV4_0;
	wire w_dff_A_ekJUKZR78_0;
	wire w_dff_A_JFzEI21U0_0;
	wire w_dff_A_K00kppmn0_0;
	wire w_dff_A_T7piVlkW3_0;
	wire w_dff_A_mzTopdh82_0;
	wire w_dff_A_ZdGf52bd0_0;
	wire w_dff_A_TGwAMCYX6_0;
	wire w_dff_A_vIRHxb962_0;
	wire w_dff_A_uAKChElf5_0;
	wire w_dff_A_tDxgDZ2d5_0;
	wire w_dff_B_T5XMTz9U6_2;
	wire w_dff_B_oWdEUL8r0_2;
	wire w_dff_B_PlkuSVZL3_2;
	wire w_dff_B_ieGEsqOi6_2;
	wire w_dff_A_tsBNwBtG2_0;
	wire w_dff_A_Puxh7rF57_0;
	wire w_dff_A_oBVWHtSO2_0;
	wire w_dff_A_nMoVTGIG1_0;
	wire w_dff_A_dORseiiV9_0;
	wire w_dff_A_eZQeiVmw7_0;
	wire w_dff_A_tnkVno0X6_0;
	wire w_dff_A_GHRCWbpx7_0;
	wire w_dff_A_XZ6qsNRu5_0;
	wire w_dff_A_EMPIVIqJ8_0;
	wire w_dff_A_f20EweG96_0;
	wire w_dff_A_w2R96mvP2_0;
	wire w_dff_A_DbO3wBK08_0;
	wire w_dff_A_oAVtPxxh4_0;
	wire w_dff_A_XTq4DLOc6_0;
	wire w_dff_A_fV5EdQbm6_0;
	wire w_dff_A_rMMEiVBk4_0;
	wire w_dff_A_AyDRLz6W7_0;
	wire w_dff_A_el3y4pEh1_0;
	wire w_dff_A_gj6iAReM1_0;
	wire w_dff_A_gSpRsrLF3_0;
	wire w_dff_A_QZC074961_0;
	wire w_dff_A_dKyqDLTN5_0;
	wire w_dff_A_Lvzh2QxO8_0;
	wire w_dff_A_bPr8US7I1_0;
	wire w_dff_A_JSfKqfWp1_0;
	wire w_dff_A_oSOxZfVn1_0;
	wire w_dff_A_9K6Bi0Ku2_0;
	wire w_dff_A_6nhii6ug1_0;
	wire w_dff_A_NUSHHJdk6_0;
	wire w_dff_A_BODOr6t57_0;
	wire w_dff_A_QWwRfLJ86_0;
	wire w_dff_A_J3oXYHUn0_0;
	wire w_dff_A_UXGuyqaF2_0;
	wire w_dff_A_vNMhoonh0_0;
	wire w_dff_A_6VrUZnzh8_0;
	wire w_dff_A_M72686594_0;
	wire w_dff_A_7TGCgdXv9_0;
	wire w_dff_A_qASn3qVF8_0;
	wire w_dff_A_IqBfVVeA8_0;
	wire w_dff_A_y8TAGmVZ6_0;
	wire w_dff_A_Gdi3fesB0_0;
	wire w_dff_A_PT0aD6DI8_0;
	wire w_dff_A_5FgW6ieE7_0;
	wire w_dff_A_lSrRblMA3_0;
	wire w_dff_A_lOTExVOr3_0;
	wire w_dff_A_LN9IRyV51_0;
	wire w_dff_A_OrXtFU6a7_0;
	wire w_dff_A_tz2LsV2S1_0;
	wire w_dff_A_a8r5XbTc3_0;
	wire w_dff_A_le8cFb526_0;
	wire w_dff_A_QLpOZsYA9_0;
	wire w_dff_A_ieqTNxBs4_0;
	wire w_dff_A_qQDJj8Dw7_0;
	wire w_dff_A_3YDIIdKx5_0;
	wire w_dff_A_zp4KvbtE6_0;
	wire w_dff_A_moDb1xJL7_0;
	wire w_dff_A_BfHPJgp10_0;
	wire w_dff_A_H0idetRW4_0;
	wire w_dff_A_1Hq53zEO5_0;
	wire w_dff_A_GkSIZpXT0_0;
	wire w_dff_A_MjREwZlV9_0;
	wire w_dff_A_Ltv5IHHs5_0;
	wire w_dff_A_0LWr4iEd8_0;
	wire w_dff_A_BvQkiO895_0;
	wire w_dff_A_K26Bpe4a1_0;
	wire w_dff_A_gTdOFDtA9_0;
	wire w_dff_A_Ty2NVLIk0_0;
	wire w_dff_A_3a69GPrT9_0;
	wire w_dff_A_sQcirZQE4_0;
	wire w_dff_A_9D5pu5wK5_0;
	wire w_dff_A_YhsIfzh68_0;
	wire w_dff_A_mt8WhnID8_0;
	wire w_dff_A_vKR8mQzE2_0;
	wire w_dff_A_ADdHF0cn6_0;
	wire w_dff_A_yxAveYNq4_0;
	wire w_dff_A_b3bpUASY0_0;
	wire w_dff_A_NIWtCpyz7_0;
	wire w_dff_A_5VKUJ0p35_0;
	wire w_dff_A_AGcqx0bD6_0;
	wire w_dff_A_Wjs34HUv3_0;
	wire w_dff_A_LGdOoEMi9_0;
	wire w_dff_A_JlPhArOH3_0;
	wire w_dff_A_KfyVvEv86_0;
	wire w_dff_A_ZJuoWG3b4_0;
	wire w_dff_A_wATpigAW5_0;
	wire w_dff_A_vzi6ZsXL0_0;
	wire w_dff_A_kEeY6YA29_0;
	wire w_dff_A_itw6IJbQ0_0;
	wire w_dff_A_QpW6nWUx4_0;
	wire w_dff_A_acs7cH5E5_0;
	wire w_dff_A_WpLjAqVQ7_0;
	wire w_dff_A_ZVjywUw11_0;
	wire w_dff_A_wDcYrBrj9_0;
	wire w_dff_A_8JOkLVhU6_0;
	wire w_dff_A_fqtUejUg2_0;
	wire w_dff_A_cTlgOsAY7_0;
	wire w_dff_A_5NKyHsij6_0;
	wire w_dff_A_8B6oZxSU6_0;
	wire w_dff_A_dWpCOdiJ9_0;
	wire w_dff_A_eSunXmXI9_0;
	wire w_dff_A_Re4YqTwz5_0;
	wire w_dff_A_37wqzGLc4_0;
	wire w_dff_A_O4HIr8ym7_0;
	wire w_dff_A_0W2MZB119_0;
	wire w_dff_A_mgt7igOC7_0;
	wire w_dff_A_jGuG0zO77_0;
	wire w_dff_A_XxKcmYcI6_0;
	wire w_dff_A_LAgFhPTz4_0;
	wire w_dff_A_UHOrkYer2_0;
	wire w_dff_A_xoOpm9Gi2_0;
	wire w_dff_A_Y1Mkm3kC6_0;
	wire w_dff_A_AqLVnBYc6_0;
	wire w_dff_A_qRvL5tm91_0;
	wire w_dff_A_FScwOEWx9_0;
	wire w_dff_A_3bTLZVW48_0;
	wire w_dff_A_PErTobiK3_0;
	wire w_dff_A_2hZ8NGte0_0;
	wire w_dff_A_HabnOg7g4_0;
	wire w_dff_A_VLgpElNv1_0;
	wire w_dff_A_krFr8OT08_0;
	wire w_dff_A_kAvTY9CC9_0;
	wire w_dff_A_Zkqq8mmR9_0;
	wire w_dff_A_cR7zXUpb8_0;
	wire w_dff_A_65adcIcR0_0;
	wire w_dff_A_GHemA6K55_0;
	wire w_dff_A_1vLGFCsA4_0;
	wire w_dff_A_E4eC3xkc8_0;
	wire w_dff_A_4WZtkrDt4_0;
	wire w_dff_A_ShH3IoYz8_0;
	wire w_dff_A_0txnnUVh5_0;
	wire w_dff_A_iHsKkUgZ6_0;
	wire w_dff_A_uKUG5bvG9_0;
	wire w_dff_A_Cr5cLS2T5_0;
	wire w_dff_A_SzdnntIp3_0;
	wire w_dff_A_nEVbT2oS9_0;
	wire w_dff_A_xMGmcRnX7_0;
	wire w_dff_A_WgSCMoXA9_0;
	wire w_dff_A_s4xXG9OR1_0;
	wire w_dff_A_G2xG24jo3_0;
	wire w_dff_A_BmtKDlhN1_0;
	wire w_dff_A_gVRjlR0a8_0;
	wire w_dff_A_n1TWzyVW1_0;
	wire w_dff_A_7TIpTwFc4_0;
	wire w_dff_A_YuU7x8F87_0;
	wire w_dff_A_6R0zsxVF9_0;
	wire w_dff_A_xw6AtxjP1_0;
	wire w_dff_A_MnPrF0Qk5_0;
	wire w_dff_A_yqqtw33N2_0;
	wire w_dff_A_GjgBXbrJ4_0;
	wire w_dff_A_Mmr638io0_0;
	wire w_dff_A_KYF4qxz23_0;
	wire w_dff_A_cq6iLv8R3_0;
	wire w_dff_A_0eqBGbxx8_0;
	wire w_dff_A_OqiMJQrW8_0;
	wire w_dff_A_Iv6qHPNr2_0;
	wire w_dff_A_3wcrrLaR8_0;
	wire w_dff_A_9yL4V7Y29_0;
	wire w_dff_A_cq0hTvsx5_0;
	wire w_dff_A_9Iv8Nqpw7_0;
	wire w_dff_A_qnkLrDhc8_0;
	wire w_dff_A_6S0Lt0No0_0;
	wire w_dff_A_e5VntDoQ3_0;
	wire w_dff_A_XTa2fve04_0;
	wire w_dff_A_GVpxtwUU3_0;
	wire w_dff_A_8oVzv6NI7_0;
	wire w_dff_A_pJvjy3wE5_0;
	wire w_dff_A_NUjeNaXw5_0;
	wire w_dff_A_90dF8Ipt2_0;
	wire w_dff_A_cD2QuQWK5_0;
	wire w_dff_A_XESSd1qZ4_0;
	wire w_dff_A_hsz9WMop4_0;
	wire w_dff_A_hQjAgRvx7_0;
	wire w_dff_A_gYxrWJE52_0;
	wire w_dff_A_jTdwQiEG0_0;
	wire w_dff_A_0X6kJbZX4_0;
	wire w_dff_A_EdUY70hO3_0;
	wire w_dff_A_CVbxJ1O45_0;
	wire w_dff_A_gcui7y3n5_0;
	wire w_dff_A_GVlw776V6_0;
	wire w_dff_A_m6f3wyN56_0;
	wire w_dff_A_lVQAAwvx6_0;
	wire w_dff_A_dYihbfry2_0;
	wire w_dff_A_M36QszLj1_0;
	wire w_dff_A_UB4x6zde0_0;
	wire w_dff_A_Z2Gbt3hQ2_0;
	wire w_dff_A_seRokvUL9_0;
	wire w_dff_A_wxPMQh1i0_0;
	wire w_dff_A_HadomRkn7_0;
	wire w_dff_A_758EfMk28_0;
	wire w_dff_A_Ptn8KJ041_0;
	wire w_dff_A_DUyp6x3e6_0;
	wire w_dff_A_NyB8ZLBp1_0;
	wire w_dff_A_QJ25Jemb0_0;
	wire w_dff_A_tTZ8JJQe0_0;
	wire w_dff_A_TKmonJqm9_0;
	wire w_dff_A_FJRfv6Cy4_0;
	wire w_dff_A_ngjVyaGw8_0;
	wire w_dff_A_gWh5xNxq1_0;
	wire w_dff_A_dlcrq6ji8_0;
	wire w_dff_A_QoZwEJHg3_0;
	wire w_dff_A_vjFxjNQc9_0;
	wire w_dff_A_ZXFIpy399_0;
	wire w_dff_A_QNYVDP5p6_0;
	wire w_dff_A_TGHBsxi64_0;
	wire w_dff_A_D1mDlDEh8_0;
	wire w_dff_A_SKytCwvL1_0;
	wire w_dff_A_BVTWiVJ57_0;
	wire w_dff_A_A7INm0il2_0;
	wire w_dff_A_vLmltr8C2_0;
	wire w_dff_A_nhO2seAI0_0;
	wire w_dff_A_NcCUgJXk9_0;
	wire w_dff_A_WVY78wq29_0;
	wire w_dff_A_aVpyQfGI2_0;
	wire w_dff_A_SOQSC0H94_0;
	wire w_dff_A_1YqQOX3r9_0;
	wire w_dff_A_ji6kDrI13_0;
	wire w_dff_A_I5NWxeFm7_0;
	wire w_dff_A_lUT0JhVq9_0;
	wire w_dff_A_ulkHrN5l1_0;
	wire w_dff_A_g8ZbEgGx9_0;
	wire w_dff_A_xnVp2jXP2_0;
	wire w_dff_A_i3LucuSc6_0;
	wire w_dff_A_eweSZZoX1_0;
	wire w_dff_A_Q5ReHvpy0_0;
	wire w_dff_A_7ce1bHCc2_0;
	wire w_dff_A_98gQezI82_0;
	wire w_dff_A_MSB5zrTF4_0;
	wire w_dff_A_bk9yXZWk1_0;
	wire w_dff_A_vSOl8sw32_0;
	wire w_dff_A_LAgxRxxT2_0;
	wire w_dff_A_ye7CMO7g0_0;
	wire w_dff_A_klgElF638_0;
	wire w_dff_A_EZtCkkGH1_0;
	wire w_dff_A_GfpiOfhm2_0;
	wire w_dff_A_qDVnjXPD7_0;
	wire w_dff_A_E2ITO4JA5_0;
	wire w_dff_A_0EfcMfr58_0;
	wire w_dff_A_AhopihAe9_0;
	wire w_dff_A_DtEhTuRv8_0;
	wire w_dff_A_wWcCxshH2_0;
	wire w_dff_A_qPO4PSNX3_0;
	wire w_dff_A_RDLDta620_0;
	wire w_dff_A_6xjoCarB1_0;
	wire w_dff_A_F9k0fKYS0_0;
	wire w_dff_A_pNrvSiDE7_0;
	wire w_dff_A_k7AQR2zg6_0;
	wire w_dff_A_07GujSiq6_0;
	wire w_dff_A_d9tJ19oG6_0;
	wire w_dff_A_4bZsYWwC2_0;
	wire w_dff_A_yrXkfJfI7_0;
	wire w_dff_A_OGfsIYmQ9_0;
	wire w_dff_A_UHLZRS6C6_0;
	wire w_dff_A_A7NXdz0I0_0;
	wire w_dff_A_Vc6VUhUq5_0;
	wire w_dff_A_5YsDD7R00_0;
	wire w_dff_A_zsHJsY5r5_0;
	wire w_dff_A_6axai51y6_0;
	wire w_dff_A_GYMBMKg37_0;
	wire w_dff_A_C9Qh45ec5_0;
	wire w_dff_A_ezaJ1M593_0;
	wire w_dff_A_Hm4zJxb31_0;
	wire w_dff_A_zjSHKnUH1_0;
	wire w_dff_A_hRf3olsM3_2;
	wire w_dff_A_t7J0DVId7_2;
	wire w_dff_A_ploDOSLu9_2;
	wire w_dff_A_2pCzVqwn2_2;
	wire w_dff_A_OfomH9JU3_2;
	wire w_dff_A_Sijv3I9R3_2;
	wire w_dff_A_Hq6WEn2f5_2;
	wire w_dff_A_ZlcuYPlk0_2;
	wire w_dff_A_v119lWYX2_2;
	wire w_dff_A_2zDjjN1h9_2;
	wire w_dff_A_1PIQUTmW3_2;
	wire w_dff_A_hpEz6GPV6_2;
	wire w_dff_A_dHt9uu4k3_2;
	wire w_dff_A_zjQaDcGc0_2;
	wire w_dff_A_DqBCJwMz4_2;
	wire w_dff_A_8mvuxWeY8_2;
	jxor g000(.dina(w_Gid12_0[2]),.dinb(w_Gid8_0[2]),.dout(n73),.clk(gclk));
	jxor g001(.dina(w_Gid4_0[2]),.dinb(w_Gid0_0[2]),.dout(n74),.clk(gclk));
	jxor g002(.dina(n74),.dinb(n73),.dout(n75),.clk(gclk));
	jand g003(.dina(w_Gr_3[1]),.dinb(Gic0),.dout(n76),.clk(gclk));
	jxor g004(.dina(w_n76_0[1]),.dinb(w_n75_0[1]),.dout(n77),.clk(gclk));
	jxor g005(.dina(w_Gid19_0[2]),.dinb(w_Gid18_0[2]),.dout(n78),.clk(gclk));
	jxor g006(.dina(w_Gid17_0[2]),.dinb(w_Gid16_0[2]),.dout(n79),.clk(gclk));
	jxor g007(.dina(n79),.dinb(n78),.dout(n80),.clk(gclk));
	jxor g008(.dina(w_Gid23_0[2]),.dinb(w_Gid22_0[2]),.dout(n81),.clk(gclk));
	jxor g009(.dina(w_Gid21_0[2]),.dinb(w_Gid20_0[2]),.dout(n82),.clk(gclk));
	jxor g010(.dina(n82),.dinb(n81),.dout(n83),.clk(gclk));
	jxor g011(.dina(w_n83_0[1]),.dinb(w_n80_0[1]),.dout(n84),.clk(gclk));
	jxor g012(.dina(w_n84_0[1]),.dinb(n77),.dout(n85),.clk(gclk));
	jxor g013(.dina(w_Gid31_0[2]),.dinb(w_Gid27_0[2]),.dout(n86),.clk(gclk));
	jxor g014(.dina(w_Gid23_0[1]),.dinb(w_Gid19_0[1]),.dout(n87),.clk(gclk));
	jxor g015(.dina(n87),.dinb(n86),.dout(n88),.clk(gclk));
	jand g016(.dina(w_Gr_3[0]),.dinb(Gic7),.dout(n89),.clk(gclk));
	jnot g017(.din(w_n89_0[1]),.dout(n90),.clk(gclk));
	jxor g018(.dina(n90),.dinb(w_n88_0[1]),.dout(n91),.clk(gclk));
	jxor g019(.dina(w_Gid7_0[2]),.dinb(w_Gid6_0[2]),.dout(n92),.clk(gclk));
	jxor g020(.dina(w_Gid5_0[2]),.dinb(w_Gid4_0[1]),.dout(n93),.clk(gclk));
	jxor g021(.dina(n93),.dinb(n92),.dout(n94),.clk(gclk));
	jxor g022(.dina(w_Gid15_0[2]),.dinb(w_Gid14_0[2]),.dout(n95),.clk(gclk));
	jxor g023(.dina(w_Gid13_0[2]),.dinb(w_Gid12_0[1]),.dout(n96),.clk(gclk));
	jxor g024(.dina(n96),.dinb(n95),.dout(n97),.clk(gclk));
	jxor g025(.dina(w_n97_0[1]),.dinb(w_n94_0[1]),.dout(n98),.clk(gclk));
	jxor g026(.dina(w_n98_0[1]),.dinb(n91),.dout(n99),.clk(gclk));
	jxor g027(.dina(w_Gid30_0[2]),.dinb(w_Gid26_0[2]),.dout(n100),.clk(gclk));
	jxor g028(.dina(w_Gid22_0[1]),.dinb(w_Gid18_0[1]),.dout(n101),.clk(gclk));
	jxor g029(.dina(n101),.dinb(n100),.dout(n102),.clk(gclk));
	jand g030(.dina(w_Gr_2[2]),.dinb(Gic6),.dout(n103),.clk(gclk));
	jxor g031(.dina(w_dff_B_ywuGzupy7_0),.dinb(n102),.dout(n104),.clk(gclk));
	jxor g032(.dina(w_Gid3_0[2]),.dinb(w_Gid2_0[2]),.dout(n105),.clk(gclk));
	jxor g033(.dina(w_Gid1_0[2]),.dinb(w_Gid0_0[1]),.dout(n106),.clk(gclk));
	jxor g034(.dina(n106),.dinb(n105),.dout(n107),.clk(gclk));
	jxor g035(.dina(w_Gid11_0[2]),.dinb(w_Gid10_0[2]),.dout(n108),.clk(gclk));
	jxor g036(.dina(w_Gid9_0[2]),.dinb(w_Gid8_0[1]),.dout(n109),.clk(gclk));
	jxor g037(.dina(n109),.dinb(n108),.dout(n110),.clk(gclk));
	jxor g038(.dina(w_n110_0[1]),.dinb(w_n107_0[1]),.dout(n111),.clk(gclk));
	jxor g039(.dina(n111),.dinb(n104),.dout(n112),.clk(gclk));
	jand g040(.dina(w_n112_2[2]),.dinb(w_n99_0[1]),.dout(n113),.clk(gclk));
	jxor g041(.dina(w_Gid13_0[1]),.dinb(w_Gid9_0[1]),.dout(n114),.clk(gclk));
	jxor g042(.dina(w_Gid5_0[1]),.dinb(w_Gid1_0[1]),.dout(n115),.clk(gclk));
	jxor g043(.dina(n115),.dinb(n114),.dout(n116),.clk(gclk));
	jand g044(.dina(w_Gr_2[1]),.dinb(Gic1),.dout(n117),.clk(gclk));
	jxor g045(.dina(w_n117_0[1]),.dinb(w_n116_0[1]),.dout(n118),.clk(gclk));
	jxor g046(.dina(w_Gid31_0[1]),.dinb(w_Gid30_0[1]),.dout(n119),.clk(gclk));
	jxor g047(.dina(w_Gid29_0[2]),.dinb(w_Gid28_0[2]),.dout(n120),.clk(gclk));
	jxor g048(.dina(n120),.dinb(n119),.dout(n121),.clk(gclk));
	jxor g049(.dina(w_Gid27_0[1]),.dinb(w_Gid26_0[1]),.dout(n122),.clk(gclk));
	jxor g050(.dina(w_Gid25_0[2]),.dinb(w_Gid24_0[2]),.dout(n123),.clk(gclk));
	jxor g051(.dina(n123),.dinb(n122),.dout(n124),.clk(gclk));
	jxor g052(.dina(w_n124_0[2]),.dinb(w_n121_0[2]),.dout(n125),.clk(gclk));
	jxor g053(.dina(w_n125_0[1]),.dinb(n118),.dout(n126),.clk(gclk));
	jxor g054(.dina(w_n126_2[1]),.dinb(w_n85_2[1]),.dout(n127),.clk(gclk));
	jand g055(.dina(w_Gr_2[0]),.dinb(Gic3),.dout(n128),.clk(gclk));
	jnot g056(.din(w_n128_0[1]),.dout(n129),.clk(gclk));
	jxor g057(.dina(n129),.dinb(w_n121_0[1]),.dout(n130),.clk(gclk));
	jxor g058(.dina(w_Gid15_0[1]),.dinb(w_Gid11_0[1]),.dout(n131),.clk(gclk));
	jxor g059(.dina(w_Gid7_0[1]),.dinb(w_Gid3_0[1]),.dout(n132),.clk(gclk));
	jxor g060(.dina(n132),.dinb(n131),.dout(n133),.clk(gclk));
	jxor g061(.dina(n133),.dinb(w_n83_0[0]),.dout(n134),.clk(gclk));
	jxor g062(.dina(w_n134_0[1]),.dinb(n130),.dout(n135),.clk(gclk));
	jand g063(.dina(w_Gr_1[2]),.dinb(Gic2),.dout(n136),.clk(gclk));
	jnot g064(.din(w_n136_0[1]),.dout(n137),.clk(gclk));
	jxor g065(.dina(n137),.dinb(w_n124_0[1]),.dout(n138),.clk(gclk));
	jxor g066(.dina(w_Gid14_0[1]),.dinb(w_Gid10_0[1]),.dout(n139),.clk(gclk));
	jxor g067(.dina(w_Gid6_0[1]),.dinb(w_Gid2_0[1]),.dout(n140),.clk(gclk));
	jxor g068(.dina(n140),.dinb(n139),.dout(n141),.clk(gclk));
	jxor g069(.dina(n141),.dinb(w_n80_0[0]),.dout(n142),.clk(gclk));
	jxor g070(.dina(w_n142_0[1]),.dinb(n138),.dout(n143),.clk(gclk));
	jand g071(.dina(w_n143_0[1]),.dinb(w_n135_0[1]),.dout(n144),.clk(gclk));
	jand g072(.dina(n144),.dinb(n127),.dout(n145),.clk(gclk));
	jxor g073(.dina(w_n128_0[0]),.dinb(w_n121_0[0]),.dout(n146),.clk(gclk));
	jxor g074(.dina(w_n134_0[0]),.dinb(n146),.dout(n147),.clk(gclk));
	jxor g075(.dina(w_n136_0[0]),.dinb(w_n124_0[0]),.dout(n148),.clk(gclk));
	jxor g076(.dina(w_n142_0[0]),.dinb(n148),.dout(n149),.clk(gclk));
	jxor g077(.dina(w_n149_2[1]),.dinb(w_n147_2[1]),.dout(n150),.clk(gclk));
	jnot g078(.din(w_n76_0[0]),.dout(n151),.clk(gclk));
	jxor g079(.dina(n151),.dinb(w_n75_0[0]),.dout(n152),.clk(gclk));
	jxor g080(.dina(w_n84_0[0]),.dinb(n152),.dout(n153),.clk(gclk));
	jnot g081(.din(w_n117_0[0]),.dout(n154),.clk(gclk));
	jxor g082(.dina(n154),.dinb(w_n116_0[0]),.dout(n155),.clk(gclk));
	jxor g083(.dina(w_n125_0[0]),.dinb(n155),.dout(n156),.clk(gclk));
	jand g084(.dina(w_n156_0[1]),.dinb(w_n153_0[1]),.dout(n157),.clk(gclk));
	jand g085(.dina(n157),.dinb(n150),.dout(n158),.clk(gclk));
	jor g086(.dina(n158),.dinb(n145),.dout(n159),.clk(gclk));
	jxor g087(.dina(w_Gid28_0[1]),.dinb(w_Gid24_0[1]),.dout(n160),.clk(gclk));
	jxor g088(.dina(w_Gid20_0[1]),.dinb(w_Gid16_0[1]),.dout(n161),.clk(gclk));
	jxor g089(.dina(n161),.dinb(n160),.dout(n162),.clk(gclk));
	jand g090(.dina(w_Gr_1[1]),.dinb(Gic4),.dout(n163),.clk(gclk));
	jxor g091(.dina(w_dff_B_aEag40On6_0),.dinb(n162),.dout(n164),.clk(gclk));
	jxor g092(.dina(w_n107_0[0]),.dinb(w_n94_0[0]),.dout(n165),.clk(gclk));
	jxor g093(.dina(n165),.dinb(n164),.dout(n166),.clk(gclk));
	jxor g094(.dina(w_Gid29_0[1]),.dinb(w_Gid25_0[1]),.dout(n167),.clk(gclk));
	jxor g095(.dina(w_Gid21_0[1]),.dinb(w_Gid17_0[1]),.dout(n168),.clk(gclk));
	jxor g096(.dina(n168),.dinb(n167),.dout(n169),.clk(gclk));
	jand g097(.dina(w_Gr_1[0]),.dinb(Gic5),.dout(n170),.clk(gclk));
	jnot g098(.din(w_n170_0[1]),.dout(n171),.clk(gclk));
	jxor g099(.dina(n171),.dinb(w_n169_0[1]),.dout(n172),.clk(gclk));
	jxor g100(.dina(w_n110_0[0]),.dinb(w_n97_0[0]),.dout(n173),.clk(gclk));
	jxor g101(.dina(w_n173_0[1]),.dinb(n172),.dout(n174),.clk(gclk));
	jand g102(.dina(w_n174_0[1]),.dinb(w_n166_2[2]),.dout(n175),.clk(gclk));
	jand g103(.dina(w_n175_0[1]),.dinb(w_n159_0[2]),.dout(n176),.clk(gclk));
	jand g104(.dina(n176),.dinb(w_n113_0[1]),.dout(n177),.clk(gclk));
	jand g105(.dina(w_n177_1[1]),.dinb(w_n85_2[0]),.dout(n178),.clk(gclk));
	jxor g106(.dina(n178),.dinb(w_Gid0_0[0]),.dout(w_dff_A_hRf3olsM3_2),.clk(gclk));
	jand g107(.dina(w_n177_1[0]),.dinb(w_n126_2[0]),.dout(n180),.clk(gclk));
	jxor g108(.dina(n180),.dinb(w_Gid1_0[0]),.dout(w_dff_A_t7J0DVId7_2),.clk(gclk));
	jand g109(.dina(w_n177_0[2]),.dinb(w_n149_2[0]),.dout(n182),.clk(gclk));
	jxor g110(.dina(n182),.dinb(w_Gid2_0[0]),.dout(w_dff_A_ploDOSLu9_2),.clk(gclk));
	jand g111(.dina(w_n177_0[1]),.dinb(w_n147_2[0]),.dout(n184),.clk(gclk));
	jxor g112(.dina(n184),.dinb(w_Gid3_0[0]),.dout(w_dff_A_2pCzVqwn2_2),.clk(gclk));
	jxor g113(.dina(w_n89_0[0]),.dinb(w_n88_0[0]),.dout(n186),.clk(gclk));
	jxor g114(.dina(w_n98_0[0]),.dinb(n186),.dout(n187),.clk(gclk));
	jnot g115(.din(w_n112_2[1]),.dout(n188),.clk(gclk));
	jand g116(.dina(w_n188_0[1]),.dinb(w_n187_2[1]),.dout(n189),.clk(gclk));
	jand g117(.dina(w_dff_B_zHKyPrEP1_0),.dinb(w_n159_0[1]),.dout(n190),.clk(gclk));
	jand g118(.dina(w_n190_0[1]),.dinb(w_n175_0[0]),.dout(n191),.clk(gclk));
	jand g119(.dina(w_n191_1[1]),.dinb(w_n85_1[2]),.dout(n192),.clk(gclk));
	jxor g120(.dina(n192),.dinb(w_Gid4_0[0]),.dout(w_dff_A_OfomH9JU3_2),.clk(gclk));
	jand g121(.dina(w_n191_1[0]),.dinb(w_n126_1[2]),.dout(n194),.clk(gclk));
	jxor g122(.dina(n194),.dinb(w_Gid5_0[0]),.dout(w_dff_A_Sijv3I9R3_2),.clk(gclk));
	jand g123(.dina(w_n191_0[2]),.dinb(w_n149_1[2]),.dout(n196),.clk(gclk));
	jxor g124(.dina(n196),.dinb(w_Gid6_0[0]),.dout(w_dff_A_Hq6WEn2f5_2),.clk(gclk));
	jand g125(.dina(w_n191_0[1]),.dinb(w_n147_1[2]),.dout(n198),.clk(gclk));
	jxor g126(.dina(n198),.dinb(w_Gid7_0[0]),.dout(w_dff_A_ZlcuYPlk0_2),.clk(gclk));
	jnot g127(.din(w_n166_2[1]),.dout(n200),.clk(gclk));
	jxor g128(.dina(w_n170_0[0]),.dinb(w_n169_0[0]),.dout(n201),.clk(gclk));
	jxor g129(.dina(w_n173_0[0]),.dinb(n201),.dout(n202),.clk(gclk));
	jand g130(.dina(w_n202_2[1]),.dinb(w_n200_0[1]),.dout(n203),.clk(gclk));
	jand g131(.dina(w_n159_0[0]),.dinb(w_n113_0[0]),.dout(n204),.clk(gclk));
	jand g132(.dina(n204),.dinb(w_n203_0[1]),.dout(n205),.clk(gclk));
	jand g133(.dina(w_n205_1[1]),.dinb(w_n85_1[1]),.dout(n206),.clk(gclk));
	jxor g134(.dina(n206),.dinb(w_Gid8_0[0]),.dout(w_dff_A_v119lWYX2_2),.clk(gclk));
	jand g135(.dina(w_n205_1[0]),.dinb(w_n126_1[1]),.dout(n208),.clk(gclk));
	jxor g136(.dina(n208),.dinb(w_Gid9_0[0]),.dout(w_dff_A_2zDjjN1h9_2),.clk(gclk));
	jand g137(.dina(w_n205_0[2]),.dinb(w_n149_1[1]),.dout(n210),.clk(gclk));
	jxor g138(.dina(n210),.dinb(w_Gid10_0[0]),.dout(w_dff_A_1PIQUTmW3_2),.clk(gclk));
	jand g139(.dina(w_n205_0[1]),.dinb(w_n147_1[1]),.dout(n212),.clk(gclk));
	jxor g140(.dina(n212),.dinb(w_Gid11_0[0]),.dout(w_dff_A_hpEz6GPV6_2),.clk(gclk));
	jand g141(.dina(w_n203_0[0]),.dinb(w_n190_0[0]),.dout(n214),.clk(gclk));
	jand g142(.dina(w_n214_1[1]),.dinb(w_n85_1[0]),.dout(n215),.clk(gclk));
	jxor g143(.dina(n215),.dinb(w_Gid12_0[0]),.dout(w_dff_A_dHt9uu4k3_2),.clk(gclk));
	jand g144(.dina(w_n214_1[0]),.dinb(w_n126_1[0]),.dout(n217),.clk(gclk));
	jxor g145(.dina(n217),.dinb(w_Gid13_0[0]),.dout(w_dff_A_zjQaDcGc0_2),.clk(gclk));
	jand g146(.dina(w_n214_0[2]),.dinb(w_n149_1[0]),.dout(n219),.clk(gclk));
	jxor g147(.dina(n219),.dinb(w_Gid14_0[0]),.dout(w_dff_A_DqBCJwMz4_2),.clk(gclk));
	jand g148(.dina(w_n214_0[1]),.dinb(w_n147_1[0]),.dout(n221),.clk(gclk));
	jxor g149(.dina(n221),.dinb(w_Gid15_0[0]),.dout(w_dff_A_8mvuxWeY8_2),.clk(gclk));
	jand g150(.dina(w_n149_0[2]),.dinb(w_n135_0[0]),.dout(n223),.clk(gclk));
	jand g151(.dina(w_n156_0[0]),.dinb(w_n85_0[2]),.dout(n224),.clk(gclk));
	jxor g152(.dina(w_n112_2[0]),.dinb(w_n187_2[0]),.dout(n225),.clk(gclk));
	jand g153(.dina(n225),.dinb(w_n174_0[0]),.dout(n226),.clk(gclk));
	jand g154(.dina(n226),.dinb(w_n200_0[0]),.dout(n227),.clk(gclk));
	jxor g155(.dina(w_n202_2[0]),.dinb(w_n166_2[0]),.dout(n228),.clk(gclk));
	jand g156(.dina(n228),.dinb(w_n99_0[0]),.dout(n229),.clk(gclk));
	jand g157(.dina(n229),.dinb(w_n188_0[0]),.dout(n230),.clk(gclk));
	jor g158(.dina(n230),.dinb(n227),.dout(n231),.clk(gclk));
	jand g159(.dina(w_n231_0[1]),.dinb(w_dff_B_UP2iUJHH5_1),.dout(n232),.clk(gclk));
	jand g160(.dina(w_n232_0[1]),.dinb(w_n223_0[1]),.dout(n233),.clk(gclk));
	jand g161(.dina(w_n233_1[1]),.dinb(w_n166_1[2]),.dout(n234),.clk(gclk));
	jxor g162(.dina(n234),.dinb(w_Gid16_0[0]),.dout(God16),.clk(gclk));
	jand g163(.dina(w_n233_1[0]),.dinb(w_n202_1[2]),.dout(n236),.clk(gclk));
	jxor g164(.dina(n236),.dinb(w_Gid17_0[0]),.dout(God17),.clk(gclk));
	jand g165(.dina(w_n233_0[2]),.dinb(w_n112_1[2]),.dout(n238),.clk(gclk));
	jxor g166(.dina(n238),.dinb(w_Gid18_0[0]),.dout(God18),.clk(gclk));
	jand g167(.dina(w_n233_0[1]),.dinb(w_n187_1[2]),.dout(n240),.clk(gclk));
	jxor g168(.dina(n240),.dinb(w_Gid19_0[0]),.dout(God19),.clk(gclk));
	jand g169(.dina(w_n143_0[0]),.dinb(w_n147_0[2]),.dout(n242),.clk(gclk));
	jand g170(.dina(w_n232_0[0]),.dinb(w_n242_0[1]),.dout(n243),.clk(gclk));
	jand g171(.dina(w_n243_1[1]),.dinb(w_n166_1[1]),.dout(n244),.clk(gclk));
	jxor g172(.dina(n244),.dinb(w_Gid20_0[0]),.dout(God20),.clk(gclk));
	jand g173(.dina(w_n243_1[0]),.dinb(w_n202_1[1]),.dout(n246),.clk(gclk));
	jxor g174(.dina(n246),.dinb(w_Gid21_0[0]),.dout(God21),.clk(gclk));
	jand g175(.dina(w_n243_0[2]),.dinb(w_n112_1[1]),.dout(n248),.clk(gclk));
	jxor g176(.dina(n248),.dinb(w_Gid22_0[0]),.dout(God22),.clk(gclk));
	jand g177(.dina(w_n243_0[1]),.dinb(w_n187_1[1]),.dout(n250),.clk(gclk));
	jxor g178(.dina(n250),.dinb(w_Gid23_0[0]),.dout(God23),.clk(gclk));
	jand g179(.dina(w_n126_0[2]),.dinb(w_n153_0[0]),.dout(n252),.clk(gclk));
	jand g180(.dina(w_n231_0[0]),.dinb(w_dff_B_SiJKSn8T2_1),.dout(n253),.clk(gclk));
	jand g181(.dina(w_n253_0[1]),.dinb(w_n223_0[0]),.dout(n254),.clk(gclk));
	jand g182(.dina(w_n254_1[1]),.dinb(w_n166_1[0]),.dout(n255),.clk(gclk));
	jxor g183(.dina(n255),.dinb(w_Gid24_0[0]),.dout(God24),.clk(gclk));
	jand g184(.dina(w_n254_1[0]),.dinb(w_n202_1[0]),.dout(n257),.clk(gclk));
	jxor g185(.dina(n257),.dinb(w_Gid25_0[0]),.dout(God25),.clk(gclk));
	jand g186(.dina(w_n254_0[2]),.dinb(w_n112_1[0]),.dout(n259),.clk(gclk));
	jxor g187(.dina(n259),.dinb(w_Gid26_0[0]),.dout(God26),.clk(gclk));
	jand g188(.dina(w_n254_0[1]),.dinb(w_n187_1[0]),.dout(n261),.clk(gclk));
	jxor g189(.dina(n261),.dinb(w_Gid27_0[0]),.dout(God27),.clk(gclk));
	jand g190(.dina(w_n253_0[0]),.dinb(w_n242_0[0]),.dout(n263),.clk(gclk));
	jand g191(.dina(w_n263_1[1]),.dinb(w_n166_0[2]),.dout(n264),.clk(gclk));
	jxor g192(.dina(n264),.dinb(w_Gid28_0[0]),.dout(God28),.clk(gclk));
	jand g193(.dina(w_n263_1[0]),.dinb(w_n202_0[2]),.dout(n266),.clk(gclk));
	jxor g194(.dina(n266),.dinb(w_Gid29_0[0]),.dout(God29),.clk(gclk));
	jand g195(.dina(w_n263_0[2]),.dinb(w_n112_0[2]),.dout(n268),.clk(gclk));
	jxor g196(.dina(n268),.dinb(w_Gid30_0[0]),.dout(God30),.clk(gclk));
	jand g197(.dina(w_n263_0[1]),.dinb(w_n187_0[2]),.dout(n270),.clk(gclk));
	jxor g198(.dina(n270),.dinb(w_Gid31_0[0]),.dout(God31),.clk(gclk));
	jspl3 jspl3_w_Gid0_0(.douta(w_dff_A_sa4OWoUW2_0),.doutb(w_Gid0_0[1]),.doutc(w_Gid0_0[2]),.din(Gid0));
	jspl3 jspl3_w_Gid1_0(.douta(w_dff_A_xyrjiOJf7_0),.doutb(w_Gid1_0[1]),.doutc(w_Gid1_0[2]),.din(Gid1));
	jspl3 jspl3_w_Gid2_0(.douta(w_dff_A_gj6iAReM1_0),.doutb(w_Gid2_0[1]),.doutc(w_Gid2_0[2]),.din(Gid2));
	jspl3 jspl3_w_Gid3_0(.douta(w_dff_A_0eqBGbxx8_0),.doutb(w_Gid3_0[1]),.doutc(w_Gid3_0[2]),.din(Gid3));
	jspl3 jspl3_w_Gid4_0(.douta(w_dff_A_yvg1r0oY8_0),.doutb(w_Gid4_0[1]),.doutc(w_Gid4_0[2]),.din(Gid4));
	jspl3 jspl3_w_Gid5_0(.douta(w_dff_A_e6qHfjer3_0),.doutb(w_Gid5_0[1]),.doutc(w_Gid5_0[2]),.din(Gid5));
	jspl3 jspl3_w_Gid6_0(.douta(w_dff_A_EMPIVIqJ8_0),.doutb(w_Gid6_0[1]),.doutc(w_Gid6_0[2]),.din(Gid6));
	jspl3 jspl3_w_Gid7_0(.douta(w_dff_A_7TIpTwFc4_0),.doutb(w_Gid7_0[1]),.doutc(w_Gid7_0[2]),.din(Gid7));
	jspl3 jspl3_w_Gid8_0(.douta(w_dff_A_tDxgDZ2d5_0),.doutb(w_Gid8_0[1]),.doutc(w_Gid8_0[2]),.din(Gid8));
	jspl3 jspl3_w_Gid9_0(.douta(w_dff_A_BbKjK4CH4_0),.doutb(w_Gid9_0[1]),.doutc(w_Gid9_0[2]),.din(Gid9));
	jspl3 jspl3_w_Gid10_0(.douta(w_dff_A_IqBfVVeA8_0),.doutb(w_Gid10_0[1]),.doutc(w_Gid10_0[2]),.din(Gid10));
	jspl3 jspl3_w_Gid11_0(.douta(w_dff_A_gYxrWJE52_0),.doutb(w_Gid11_0[1]),.doutc(w_Gid11_0[2]),.din(Gid11));
	jspl3 jspl3_w_Gid12_0(.douta(w_dff_A_VnYVtnKV4_0),.doutb(w_Gid12_0[1]),.doutc(w_Gid12_0[2]),.din(Gid12));
	jspl3 jspl3_w_Gid13_0(.douta(w_dff_A_e19BsMgq7_0),.doutb(w_Gid13_0[1]),.doutc(w_Gid13_0[2]),.din(Gid13));
	jspl3 jspl3_w_Gid14_0(.douta(w_dff_A_NUSHHJdk6_0),.doutb(w_Gid14_0[1]),.doutc(w_Gid14_0[2]),.din(Gid14));
	jspl3 jspl3_w_Gid15_0(.douta(w_dff_A_XTa2fve04_0),.doutb(w_Gid15_0[1]),.doutc(w_Gid15_0[2]),.din(Gid15));
	jspl3 jspl3_w_Gid16_0(.douta(w_dff_A_MjREwZlV9_0),.doutb(w_Gid16_0[1]),.doutc(w_Gid16_0[2]),.din(Gid16));
	jspl3 jspl3_w_Gid17_0(.douta(w_dff_A_le8cFb526_0),.doutb(w_Gid17_0[1]),.doutc(w_Gid17_0[2]),.din(Gid17));
	jspl3 jspl3_w_Gid18_0(.douta(w_dff_A_KfyVvEv86_0),.doutb(w_Gid18_0[1]),.doutc(w_Gid18_0[2]),.din(Gid18));
	jspl3 jspl3_w_Gid19_0(.douta(w_dff_A_mt8WhnID8_0),.doutb(w_Gid19_0[1]),.doutc(w_Gid19_0[2]),.din(Gid19));
	jspl3 jspl3_w_Gid20_0(.douta(w_dff_A_TKmonJqm9_0),.doutb(w_Gid20_0[1]),.doutc(w_Gid20_0[2]),.din(Gid20));
	jspl3 jspl3_w_Gid21_0(.douta(w_dff_A_UB4x6zde0_0),.doutb(w_Gid21_0[1]),.doutc(w_Gid21_0[2]),.din(Gid21));
	jspl3 jspl3_w_Gid22_0(.douta(w_dff_A_I5NWxeFm7_0),.doutb(w_Gid22_0[1]),.doutc(w_Gid22_0[2]),.din(Gid22));
	jspl3 jspl3_w_Gid23_0(.douta(w_dff_A_SKytCwvL1_0),.doutb(w_Gid23_0[1]),.doutc(w_Gid23_0[2]),.din(Gid23));
	jspl3 jspl3_w_Gid24_0(.douta(w_dff_A_jGuG0zO77_0),.doutb(w_Gid24_0[1]),.doutc(w_Gid24_0[2]),.din(Gid24));
	jspl3 jspl3_w_Gid25_0(.douta(w_dff_A_fqtUejUg2_0),.doutb(w_Gid25_0[1]),.doutc(w_Gid25_0[2]),.din(Gid25));
	jspl3 jspl3_w_Gid26_0(.douta(w_dff_A_4WZtkrDt4_0),.doutb(w_Gid26_0[1]),.doutc(w_Gid26_0[2]),.din(Gid26));
	jspl3 jspl3_w_Gid27_0(.douta(w_dff_A_2hZ8NGte0_0),.doutb(w_Gid27_0[1]),.doutc(w_Gid27_0[2]),.din(Gid27));
	jspl3 jspl3_w_Gid28_0(.douta(w_dff_A_wWcCxshH2_0),.doutb(w_Gid28_0[1]),.doutc(w_Gid28_0[2]),.din(Gid28));
	jspl3 jspl3_w_Gid29_0(.douta(w_dff_A_vSOl8sw32_0),.doutb(w_Gid29_0[1]),.doutc(w_Gid29_0[2]),.din(Gid29));
	jspl3 jspl3_w_Gid30_0(.douta(w_dff_A_zjSHKnUH1_0),.doutb(w_Gid30_0[1]),.doutc(w_Gid30_0[2]),.din(Gid30));
	jspl3 jspl3_w_Gid31_0(.douta(w_dff_A_OGfsIYmQ9_0),.doutb(w_Gid31_0[1]),.doutc(w_Gid31_0[2]),.din(Gid31));
	jspl3 jspl3_w_Gr_0(.douta(w_Gr_0[0]),.doutb(w_Gr_0[1]),.doutc(w_Gr_0[2]),.din(Gr));
	jspl3 jspl3_w_Gr_1(.douta(w_Gr_1[0]),.doutb(w_Gr_1[1]),.doutc(w_Gr_1[2]),.din(w_Gr_0[0]));
	jspl3 jspl3_w_Gr_2(.douta(w_Gr_2[0]),.doutb(w_Gr_2[1]),.doutc(w_Gr_2[2]),.din(w_Gr_0[1]));
	jspl jspl_w_Gr_3(.douta(w_Gr_3[0]),.doutb(w_Gr_3[1]),.din(w_Gr_0[2]));
	jspl jspl_w_n75_0(.douta(w_n75_0[0]),.doutb(w_n75_0[1]),.din(n75));
	jspl jspl_w_n76_0(.douta(w_n76_0[0]),.doutb(w_dff_A_fwCw01320_1),.din(n76));
	jspl jspl_w_n80_0(.douta(w_n80_0[0]),.doutb(w_n80_0[1]),.din(n80));
	jspl jspl_w_n83_0(.douta(w_n83_0[0]),.doutb(w_n83_0[1]),.din(n83));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.din(n84));
	jspl3 jspl3_w_n85_0(.douta(w_dff_A_KyGKnG4J0_0),.doutb(w_n85_0[1]),.doutc(w_n85_0[2]),.din(n85));
	jspl3 jspl3_w_n85_1(.douta(w_n85_1[0]),.doutb(w_n85_1[1]),.doutc(w_n85_1[2]),.din(w_n85_0[0]));
	jspl jspl_w_n85_2(.douta(w_dff_A_ruSJ223S5_0),.doutb(w_n85_2[1]),.din(w_n85_0[1]));
	jspl jspl_w_n88_0(.douta(w_n88_0[0]),.doutb(w_n88_0[1]),.din(n88));
	jspl jspl_w_n89_0(.douta(w_dff_A_EjtYTGZI6_0),.doutb(w_n89_0[1]),.din(n89));
	jspl jspl_w_n94_0(.douta(w_n94_0[0]),.doutb(w_n94_0[1]),.din(n94));
	jspl jspl_w_n97_0(.douta(w_n97_0[0]),.doutb(w_n97_0[1]),.din(n97));
	jspl jspl_w_n98_0(.douta(w_n98_0[0]),.doutb(w_n98_0[1]),.din(n98));
	jspl jspl_w_n99_0(.douta(w_dff_A_qTQMxoJR3_0),.doutb(w_n99_0[1]),.din(n99));
	jspl jspl_w_n107_0(.douta(w_n107_0[0]),.doutb(w_n107_0[1]),.din(n107));
	jspl jspl_w_n110_0(.douta(w_n110_0[0]),.doutb(w_n110_0[1]),.din(n110));
	jspl3 jspl3_w_n112_0(.douta(w_dff_A_72r887Db9_0),.doutb(w_n112_0[1]),.doutc(w_dff_A_Dqwi5yCP5_2),.din(n112));
	jspl3 jspl3_w_n112_1(.douta(w_n112_1[0]),.doutb(w_n112_1[1]),.doutc(w_n112_1[2]),.din(w_n112_0[0]));
	jspl3 jspl3_w_n112_2(.douta(w_n112_2[0]),.doutb(w_n112_2[1]),.doutc(w_n112_2[2]),.din(w_n112_0[1]));
	jspl jspl_w_n113_0(.douta(w_n113_0[0]),.doutb(w_dff_A_XJJO2q9r6_1),.din(w_dff_B_9popjFMI6_2));
	jspl jspl_w_n116_0(.douta(w_n116_0[0]),.doutb(w_n116_0[1]),.din(n116));
	jspl jspl_w_n117_0(.douta(w_n117_0[0]),.doutb(w_dff_A_KKZrZLki5_1),.din(n117));
	jspl3 jspl3_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.doutc(w_n121_0[2]),.din(n121));
	jspl3 jspl3_w_n124_0(.douta(w_n124_0[0]),.doutb(w_n124_0[1]),.doutc(w_n124_0[2]),.din(n124));
	jspl jspl_w_n125_0(.douta(w_n125_0[0]),.doutb(w_n125_0[1]),.din(n125));
	jspl3 jspl3_w_n126_0(.douta(w_dff_A_8d4fuzZb7_0),.doutb(w_n126_0[1]),.doutc(w_n126_0[2]),.din(n126));
	jspl3 jspl3_w_n126_1(.douta(w_n126_1[0]),.doutb(w_n126_1[1]),.doutc(w_n126_1[2]),.din(w_n126_0[0]));
	jspl jspl_w_n126_2(.douta(w_dff_A_fbABUCyq5_0),.doutb(w_n126_2[1]),.din(w_n126_0[1]));
	jspl jspl_w_n128_0(.douta(w_dff_A_lUT0JhVq9_0),.doutb(w_n128_0[1]),.din(n128));
	jspl jspl_w_n134_0(.douta(w_n134_0[0]),.doutb(w_n134_0[1]),.din(n134));
	jspl jspl_w_n135_0(.douta(w_n135_0[0]),.doutb(w_n135_0[1]),.din(n135));
	jspl jspl_w_n136_0(.douta(w_dff_A_ZJuoWG3b4_0),.doutb(w_n136_0[1]),.din(n136));
	jspl jspl_w_n142_0(.douta(w_n142_0[0]),.doutb(w_n142_0[1]),.din(n142));
	jspl jspl_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.din(n143));
	jspl3 jspl3_w_n147_0(.douta(w_dff_A_Cr5cLS2T5_0),.doutb(w_n147_0[1]),.doutc(w_n147_0[2]),.din(n147));
	jspl3 jspl3_w_n147_1(.douta(w_n147_1[0]),.doutb(w_n147_1[1]),.doutc(w_n147_1[2]),.din(w_n147_0[0]));
	jspl jspl_w_n147_2(.douta(w_dff_A_vHS6vKCS8_0),.doutb(w_n147_2[1]),.din(w_n147_0[1]));
	jspl3 jspl3_w_n149_0(.douta(w_dff_A_ABa81DUA2_0),.doutb(w_n149_0[1]),.doutc(w_n149_0[2]),.din(n149));
	jspl3 jspl3_w_n149_1(.douta(w_n149_1[0]),.doutb(w_n149_1[1]),.doutc(w_n149_1[2]),.din(w_n149_0[0]));
	jspl jspl_w_n149_2(.douta(w_dff_A_oIJUwFqg1_0),.doutb(w_n149_2[1]),.din(w_n149_0[1]));
	jspl jspl_w_n153_0(.douta(w_n153_0[0]),.doutb(w_n153_0[1]),.din(n153));
	jspl jspl_w_n156_0(.douta(w_n156_0[0]),.doutb(w_n156_0[1]),.din(n156));
	jspl3 jspl3_w_n159_0(.douta(w_n159_0[0]),.doutb(w_n159_0[1]),.doutc(w_n159_0[2]),.din(n159));
	jspl3 jspl3_w_n166_0(.douta(w_dff_A_cP9xoJ6c9_0),.doutb(w_n166_0[1]),.doutc(w_dff_A_qrpZZJsb1_2),.din(n166));
	jspl3 jspl3_w_n166_1(.douta(w_n166_1[0]),.doutb(w_n166_1[1]),.doutc(w_n166_1[2]),.din(w_n166_0[0]));
	jspl3 jspl3_w_n166_2(.douta(w_n166_2[0]),.doutb(w_n166_2[1]),.doutc(w_n166_2[2]),.din(w_n166_0[1]));
	jspl jspl_w_n169_0(.douta(w_n169_0[0]),.doutb(w_n169_0[1]),.din(n169));
	jspl jspl_w_n170_0(.douta(w_dff_A_ubP4lckB7_0),.doutb(w_n170_0[1]),.din(n170));
	jspl jspl_w_n173_0(.douta(w_n173_0[0]),.doutb(w_n173_0[1]),.din(n173));
	jspl jspl_w_n174_0(.douta(w_dff_A_c6Ggwwcr9_0),.doutb(w_n174_0[1]),.din(n174));
	jspl jspl_w_n175_0(.douta(w_dff_A_NMBiPfA08_0),.doutb(w_n175_0[1]),.din(w_dff_B_BlATRo9z6_2));
	jspl3 jspl3_w_n177_0(.douta(w_n177_0[0]),.doutb(w_n177_0[1]),.doutc(w_n177_0[2]),.din(n177));
	jspl jspl_w_n177_1(.douta(w_n177_1[0]),.doutb(w_n177_1[1]),.din(w_n177_0[0]));
	jspl3 jspl3_w_n187_0(.douta(w_dff_A_PAHZ1fb39_0),.doutb(w_n187_0[1]),.doutc(w_dff_A_LnCvSuYw3_2),.din(n187));
	jspl3 jspl3_w_n187_1(.douta(w_n187_1[0]),.doutb(w_n187_1[1]),.doutc(w_n187_1[2]),.din(w_n187_0[0]));
	jspl jspl_w_n187_2(.douta(w_n187_2[0]),.doutb(w_dff_A_gUpsNhdc7_1),.din(w_n187_0[1]));
	jspl jspl_w_n188_0(.douta(w_dff_A_ouv0uQWH6_0),.doutb(w_n188_0[1]),.din(n188));
	jspl jspl_w_n190_0(.douta(w_n190_0[0]),.doutb(w_n190_0[1]),.din(n190));
	jspl3 jspl3_w_n191_0(.douta(w_n191_0[0]),.doutb(w_n191_0[1]),.doutc(w_n191_0[2]),.din(n191));
	jspl jspl_w_n191_1(.douta(w_n191_1[0]),.doutb(w_n191_1[1]),.din(w_n191_0[0]));
	jspl jspl_w_n200_0(.douta(w_dff_A_OkNIja8V9_0),.doutb(w_n200_0[1]),.din(n200));
	jspl3 jspl3_w_n202_0(.douta(w_dff_A_JPw379yx3_0),.doutb(w_n202_0[1]),.doutc(w_dff_A_PGQM1ifd1_2),.din(n202));
	jspl3 jspl3_w_n202_1(.douta(w_n202_1[0]),.doutb(w_n202_1[1]),.doutc(w_n202_1[2]),.din(w_n202_0[0]));
	jspl jspl_w_n202_2(.douta(w_n202_2[0]),.doutb(w_dff_A_YVygMPnc2_1),.din(w_n202_0[1]));
	jspl jspl_w_n203_0(.douta(w_n203_0[0]),.doutb(w_n203_0[1]),.din(w_dff_B_4WY4MvOC7_2));
	jspl3 jspl3_w_n205_0(.douta(w_n205_0[0]),.doutb(w_n205_0[1]),.doutc(w_n205_0[2]),.din(n205));
	jspl jspl_w_n205_1(.douta(w_n205_1[0]),.doutb(w_n205_1[1]),.din(w_n205_0[0]));
	jspl3 jspl3_w_n214_0(.douta(w_n214_0[0]),.doutb(w_n214_0[1]),.doutc(w_n214_0[2]),.din(n214));
	jspl jspl_w_n214_1(.douta(w_n214_1[0]),.doutb(w_n214_1[1]),.din(w_n214_0[0]));
	jspl jspl_w_n223_0(.douta(w_n223_0[0]),.doutb(w_n223_0[1]),.din(w_dff_B_ZWbj9Uoc7_2));
	jspl jspl_w_n231_0(.douta(w_n231_0[0]),.doutb(w_n231_0[1]),.din(n231));
	jspl jspl_w_n232_0(.douta(w_n232_0[0]),.doutb(w_n232_0[1]),.din(n232));
	jspl3 jspl3_w_n233_0(.douta(w_n233_0[0]),.doutb(w_n233_0[1]),.doutc(w_n233_0[2]),.din(n233));
	jspl jspl_w_n233_1(.douta(w_n233_1[0]),.doutb(w_n233_1[1]),.din(w_n233_0[0]));
	jspl jspl_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.din(w_dff_B_ieGEsqOi6_2));
	jspl3 jspl3_w_n243_0(.douta(w_n243_0[0]),.doutb(w_n243_0[1]),.doutc(w_n243_0[2]),.din(n243));
	jspl jspl_w_n243_1(.douta(w_n243_1[0]),.doutb(w_n243_1[1]),.din(w_n243_0[0]));
	jspl jspl_w_n253_0(.douta(w_n253_0[0]),.doutb(w_n253_0[1]),.din(n253));
	jspl3 jspl3_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.doutc(w_n254_0[2]),.din(n254));
	jspl jspl_w_n254_1(.douta(w_n254_1[0]),.doutb(w_n254_1[1]),.din(w_n254_0[0]));
	jspl3 jspl3_w_n263_0(.douta(w_n263_0[0]),.doutb(w_n263_0[1]),.doutc(w_n263_0[2]),.din(n263));
	jspl jspl_w_n263_1(.douta(w_n263_1[0]),.doutb(w_n263_1[1]),.din(w_n263_0[0]));
	jdff dff_A_NMBiPfA08_0(.dout(w_n175_0[0]),.din(w_dff_A_NMBiPfA08_0),.clk(gclk));
	jdff dff_B_i5RHafzQ4_2(.din(n175),.dout(w_dff_B_i5RHafzQ4_2),.clk(gclk));
	jdff dff_B_BlATRo9z6_2(.din(w_dff_B_i5RHafzQ4_2),.dout(w_dff_B_BlATRo9z6_2),.clk(gclk));
	jdff dff_A_XJJO2q9r6_1(.dout(w_n113_0[1]),.din(w_dff_A_XJJO2q9r6_1),.clk(gclk));
	jdff dff_B_ovUR52QR4_2(.din(n113),.dout(w_dff_B_ovUR52QR4_2),.clk(gclk));
	jdff dff_B_9popjFMI6_2(.din(w_dff_B_ovUR52QR4_2),.dout(w_dff_B_9popjFMI6_2),.clk(gclk));
	jdff dff_B_VB8GMIr55_2(.din(n203),.dout(w_dff_B_VB8GMIr55_2),.clk(gclk));
	jdff dff_B_4WY4MvOC7_2(.din(w_dff_B_VB8GMIr55_2),.dout(w_dff_B_4WY4MvOC7_2),.clk(gclk));
	jdff dff_B_zHKyPrEP1_0(.din(n189),.dout(w_dff_B_zHKyPrEP1_0),.clk(gclk));
	jdff dff_A_SWz2spEd1_0(.dout(w_n149_2[0]),.din(w_dff_A_SWz2spEd1_0),.clk(gclk));
	jdff dff_A_rJGPT1mb0_0(.dout(w_dff_A_SWz2spEd1_0),.din(w_dff_A_rJGPT1mb0_0),.clk(gclk));
	jdff dff_A_fXuAndlD2_0(.dout(w_dff_A_rJGPT1mb0_0),.din(w_dff_A_fXuAndlD2_0),.clk(gclk));
	jdff dff_A_P0ku1e5Z3_0(.dout(w_dff_A_fXuAndlD2_0),.din(w_dff_A_P0ku1e5Z3_0),.clk(gclk));
	jdff dff_A_oIJUwFqg1_0(.dout(w_dff_A_P0ku1e5Z3_0),.din(w_dff_A_oIJUwFqg1_0),.clk(gclk));
	jdff dff_A_mkT8y3ij7_0(.dout(w_n147_2[0]),.din(w_dff_A_mkT8y3ij7_0),.clk(gclk));
	jdff dff_A_bG008g873_0(.dout(w_dff_A_mkT8y3ij7_0),.din(w_dff_A_bG008g873_0),.clk(gclk));
	jdff dff_A_lQ2q4qAY8_0(.dout(w_dff_A_bG008g873_0),.din(w_dff_A_lQ2q4qAY8_0),.clk(gclk));
	jdff dff_A_OJQf32ar2_0(.dout(w_dff_A_lQ2q4qAY8_0),.din(w_dff_A_OJQf32ar2_0),.clk(gclk));
	jdff dff_A_vHS6vKCS8_0(.dout(w_dff_A_OJQf32ar2_0),.din(w_dff_A_vHS6vKCS8_0),.clk(gclk));
	jdff dff_A_JeCenFCG2_0(.dout(w_n126_2[0]),.din(w_dff_A_JeCenFCG2_0),.clk(gclk));
	jdff dff_A_0rJHf0kh2_0(.dout(w_dff_A_JeCenFCG2_0),.din(w_dff_A_0rJHf0kh2_0),.clk(gclk));
	jdff dff_A_glL36dua6_0(.dout(w_dff_A_0rJHf0kh2_0),.din(w_dff_A_glL36dua6_0),.clk(gclk));
	jdff dff_A_kPJ7yxd81_0(.dout(w_dff_A_glL36dua6_0),.din(w_dff_A_kPJ7yxd81_0),.clk(gclk));
	jdff dff_A_fbABUCyq5_0(.dout(w_dff_A_kPJ7yxd81_0),.din(w_dff_A_fbABUCyq5_0),.clk(gclk));
	jdff dff_A_HqOMbToB3_0(.dout(w_n85_2[0]),.din(w_dff_A_HqOMbToB3_0),.clk(gclk));
	jdff dff_A_0pZYsjtK0_0(.dout(w_dff_A_HqOMbToB3_0),.din(w_dff_A_0pZYsjtK0_0),.clk(gclk));
	jdff dff_A_8cGMO4gZ7_0(.dout(w_dff_A_0pZYsjtK0_0),.din(w_dff_A_8cGMO4gZ7_0),.clk(gclk));
	jdff dff_A_1eqpj8yC3_0(.dout(w_dff_A_8cGMO4gZ7_0),.din(w_dff_A_1eqpj8yC3_0),.clk(gclk));
	jdff dff_A_ruSJ223S5_0(.dout(w_dff_A_1eqpj8yC3_0),.din(w_dff_A_ruSJ223S5_0),.clk(gclk));
	jdff dff_B_x3t1SBEh7_1(.din(n224),.dout(w_dff_B_x3t1SBEh7_1),.clk(gclk));
	jdff dff_B_0hFeU7G62_1(.din(w_dff_B_x3t1SBEh7_1),.dout(w_dff_B_0hFeU7G62_1),.clk(gclk));
	jdff dff_B_UP2iUJHH5_1(.din(w_dff_B_0hFeU7G62_1),.dout(w_dff_B_UP2iUJHH5_1),.clk(gclk));
	jdff dff_A_SeGZvjhO2_0(.dout(w_n85_0[0]),.din(w_dff_A_SeGZvjhO2_0),.clk(gclk));
	jdff dff_A_ioAbq98N2_0(.dout(w_dff_A_SeGZvjhO2_0),.din(w_dff_A_ioAbq98N2_0),.clk(gclk));
	jdff dff_A_w6CKBAb81_0(.dout(w_dff_A_ioAbq98N2_0),.din(w_dff_A_w6CKBAb81_0),.clk(gclk));
	jdff dff_A_bBbp3GfD5_0(.dout(w_dff_A_w6CKBAb81_0),.din(w_dff_A_bBbp3GfD5_0),.clk(gclk));
	jdff dff_A_KyGKnG4J0_0(.dout(w_dff_A_bBbp3GfD5_0),.din(w_dff_A_KyGKnG4J0_0),.clk(gclk));
	jdff dff_B_KaBJ0nU53_2(.din(n223),.dout(w_dff_B_KaBJ0nU53_2),.clk(gclk));
	jdff dff_B_QyfcK6VF0_2(.din(w_dff_B_KaBJ0nU53_2),.dout(w_dff_B_QyfcK6VF0_2),.clk(gclk));
	jdff dff_B_dm0QMdOB0_2(.din(w_dff_B_QyfcK6VF0_2),.dout(w_dff_B_dm0QMdOB0_2),.clk(gclk));
	jdff dff_B_ZWbj9Uoc7_2(.din(w_dff_B_dm0QMdOB0_2),.dout(w_dff_B_ZWbj9Uoc7_2),.clk(gclk));
	jdff dff_A_OhuAyLz43_0(.dout(w_n149_0[0]),.din(w_dff_A_OhuAyLz43_0),.clk(gclk));
	jdff dff_A_1B1ZXF3c1_0(.dout(w_dff_A_OhuAyLz43_0),.din(w_dff_A_1B1ZXF3c1_0),.clk(gclk));
	jdff dff_A_UvrBQeLx0_0(.dout(w_dff_A_1B1ZXF3c1_0),.din(w_dff_A_UvrBQeLx0_0),.clk(gclk));
	jdff dff_A_F23V6yfT8_0(.dout(w_dff_A_UvrBQeLx0_0),.din(w_dff_A_F23V6yfT8_0),.clk(gclk));
	jdff dff_A_ABa81DUA2_0(.dout(w_dff_A_F23V6yfT8_0),.din(w_dff_A_ABa81DUA2_0),.clk(gclk));
	jdff dff_B_vwVK4pL53_1(.din(n252),.dout(w_dff_B_vwVK4pL53_1),.clk(gclk));
	jdff dff_B_cYETG44L4_1(.din(w_dff_B_vwVK4pL53_1),.dout(w_dff_B_cYETG44L4_1),.clk(gclk));
	jdff dff_B_SiJKSn8T2_1(.din(w_dff_B_cYETG44L4_1),.dout(w_dff_B_SiJKSn8T2_1),.clk(gclk));
	jdff dff_A_YVygMPnc2_1(.dout(w_n202_2[1]),.din(w_dff_A_YVygMPnc2_1),.clk(gclk));
	jdff dff_A_tf9Ujzwn5_0(.dout(w_n202_0[0]),.din(w_dff_A_tf9Ujzwn5_0),.clk(gclk));
	jdff dff_A_VpaXB0Rf4_0(.dout(w_dff_A_tf9Ujzwn5_0),.din(w_dff_A_VpaXB0Rf4_0),.clk(gclk));
	jdff dff_A_DghHOQ6g0_0(.dout(w_dff_A_VpaXB0Rf4_0),.din(w_dff_A_DghHOQ6g0_0),.clk(gclk));
	jdff dff_A_AKcise4m2_0(.dout(w_dff_A_DghHOQ6g0_0),.din(w_dff_A_AKcise4m2_0),.clk(gclk));
	jdff dff_A_2B6XvYHh7_0(.dout(w_dff_A_AKcise4m2_0),.din(w_dff_A_2B6XvYHh7_0),.clk(gclk));
	jdff dff_A_JPw379yx3_0(.dout(w_dff_A_2B6XvYHh7_0),.din(w_dff_A_JPw379yx3_0),.clk(gclk));
	jdff dff_A_eKtt4Lqq4_2(.dout(w_n202_0[2]),.din(w_dff_A_eKtt4Lqq4_2),.clk(gclk));
	jdff dff_A_3NFEPZyu6_2(.dout(w_dff_A_eKtt4Lqq4_2),.din(w_dff_A_3NFEPZyu6_2),.clk(gclk));
	jdff dff_A_cMNxwI0D2_2(.dout(w_dff_A_3NFEPZyu6_2),.din(w_dff_A_cMNxwI0D2_2),.clk(gclk));
	jdff dff_A_R0kSpJKS2_2(.dout(w_dff_A_cMNxwI0D2_2),.din(w_dff_A_R0kSpJKS2_2),.clk(gclk));
	jdff dff_A_o2C4NKxh7_2(.dout(w_dff_A_R0kSpJKS2_2),.din(w_dff_A_o2C4NKxh7_2),.clk(gclk));
	jdff dff_A_PGQM1ifd1_2(.dout(w_dff_A_o2C4NKxh7_2),.din(w_dff_A_PGQM1ifd1_2),.clk(gclk));
	jdff dff_A_qTQMxoJR3_0(.dout(w_n99_0[0]),.din(w_dff_A_qTQMxoJR3_0),.clk(gclk));
	jdff dff_A_ouv0uQWH6_0(.dout(w_n188_0[0]),.din(w_dff_A_ouv0uQWH6_0),.clk(gclk));
	jdff dff_A_IikaIfS06_0(.dout(w_n112_0[0]),.din(w_dff_A_IikaIfS06_0),.clk(gclk));
	jdff dff_A_nBvOlsvz2_0(.dout(w_dff_A_IikaIfS06_0),.din(w_dff_A_nBvOlsvz2_0),.clk(gclk));
	jdff dff_A_pbXl2sc08_0(.dout(w_dff_A_nBvOlsvz2_0),.din(w_dff_A_pbXl2sc08_0),.clk(gclk));
	jdff dff_A_ZLfkpWer1_0(.dout(w_dff_A_pbXl2sc08_0),.din(w_dff_A_ZLfkpWer1_0),.clk(gclk));
	jdff dff_A_9JwpWNHu3_0(.dout(w_dff_A_ZLfkpWer1_0),.din(w_dff_A_9JwpWNHu3_0),.clk(gclk));
	jdff dff_A_72r887Db9_0(.dout(w_dff_A_9JwpWNHu3_0),.din(w_dff_A_72r887Db9_0),.clk(gclk));
	jdff dff_A_f9xfAcPB4_2(.dout(w_n112_0[2]),.din(w_dff_A_f9xfAcPB4_2),.clk(gclk));
	jdff dff_A_YTWGeupH2_2(.dout(w_dff_A_f9xfAcPB4_2),.din(w_dff_A_YTWGeupH2_2),.clk(gclk));
	jdff dff_A_Z7YB01u19_2(.dout(w_dff_A_YTWGeupH2_2),.din(w_dff_A_Z7YB01u19_2),.clk(gclk));
	jdff dff_A_I18bsbrJ5_2(.dout(w_dff_A_Z7YB01u19_2),.din(w_dff_A_I18bsbrJ5_2),.clk(gclk));
	jdff dff_A_YHhTEY4p9_2(.dout(w_dff_A_I18bsbrJ5_2),.din(w_dff_A_YHhTEY4p9_2),.clk(gclk));
	jdff dff_A_Dqwi5yCP5_2(.dout(w_dff_A_YHhTEY4p9_2),.din(w_dff_A_Dqwi5yCP5_2),.clk(gclk));
	jdff dff_B_ywuGzupy7_0(.din(n103),.dout(w_dff_B_ywuGzupy7_0),.clk(gclk));
	jdff dff_A_gUpsNhdc7_1(.dout(w_n187_2[1]),.din(w_dff_A_gUpsNhdc7_1),.clk(gclk));
	jdff dff_A_val0AqY39_0(.dout(w_n187_0[0]),.din(w_dff_A_val0AqY39_0),.clk(gclk));
	jdff dff_A_UqUR8uJH8_0(.dout(w_dff_A_val0AqY39_0),.din(w_dff_A_UqUR8uJH8_0),.clk(gclk));
	jdff dff_A_na1l1pxG7_0(.dout(w_dff_A_UqUR8uJH8_0),.din(w_dff_A_na1l1pxG7_0),.clk(gclk));
	jdff dff_A_y05OQNLB5_0(.dout(w_dff_A_na1l1pxG7_0),.din(w_dff_A_y05OQNLB5_0),.clk(gclk));
	jdff dff_A_R84Nkzu12_0(.dout(w_dff_A_y05OQNLB5_0),.din(w_dff_A_R84Nkzu12_0),.clk(gclk));
	jdff dff_A_PAHZ1fb39_0(.dout(w_dff_A_R84Nkzu12_0),.din(w_dff_A_PAHZ1fb39_0),.clk(gclk));
	jdff dff_A_DvnNR7Gr8_2(.dout(w_n187_0[2]),.din(w_dff_A_DvnNR7Gr8_2),.clk(gclk));
	jdff dff_A_PaJcP9C26_2(.dout(w_dff_A_DvnNR7Gr8_2),.din(w_dff_A_PaJcP9C26_2),.clk(gclk));
	jdff dff_A_BCLd1tN77_2(.dout(w_dff_A_PaJcP9C26_2),.din(w_dff_A_BCLd1tN77_2),.clk(gclk));
	jdff dff_A_apl5VkCD0_2(.dout(w_dff_A_BCLd1tN77_2),.din(w_dff_A_apl5VkCD0_2),.clk(gclk));
	jdff dff_A_2CqtsBqC1_2(.dout(w_dff_A_apl5VkCD0_2),.din(w_dff_A_2CqtsBqC1_2),.clk(gclk));
	jdff dff_A_LnCvSuYw3_2(.dout(w_dff_A_2CqtsBqC1_2),.din(w_dff_A_LnCvSuYw3_2),.clk(gclk));
	jdff dff_A_EjtYTGZI6_0(.dout(w_n89_0[0]),.din(w_dff_A_EjtYTGZI6_0),.clk(gclk));
	jdff dff_A_c6Ggwwcr9_0(.dout(w_n174_0[0]),.din(w_dff_A_c6Ggwwcr9_0),.clk(gclk));
	jdff dff_A_ubP4lckB7_0(.dout(w_n170_0[0]),.din(w_dff_A_ubP4lckB7_0),.clk(gclk));
	jdff dff_A_OkNIja8V9_0(.dout(w_n200_0[0]),.din(w_dff_A_OkNIja8V9_0),.clk(gclk));
	jdff dff_A_zwdJ1dsv9_0(.dout(w_n166_0[0]),.din(w_dff_A_zwdJ1dsv9_0),.clk(gclk));
	jdff dff_A_BQgqP7PY5_0(.dout(w_dff_A_zwdJ1dsv9_0),.din(w_dff_A_BQgqP7PY5_0),.clk(gclk));
	jdff dff_A_nW1BTbHm3_0(.dout(w_dff_A_BQgqP7PY5_0),.din(w_dff_A_nW1BTbHm3_0),.clk(gclk));
	jdff dff_A_qzBcH4iu1_0(.dout(w_dff_A_nW1BTbHm3_0),.din(w_dff_A_qzBcH4iu1_0),.clk(gclk));
	jdff dff_A_oEJq5Y129_0(.dout(w_dff_A_qzBcH4iu1_0),.din(w_dff_A_oEJq5Y129_0),.clk(gclk));
	jdff dff_A_cP9xoJ6c9_0(.dout(w_dff_A_oEJq5Y129_0),.din(w_dff_A_cP9xoJ6c9_0),.clk(gclk));
	jdff dff_A_CZtdIhDC9_2(.dout(w_n166_0[2]),.din(w_dff_A_CZtdIhDC9_2),.clk(gclk));
	jdff dff_A_aZRWhOKy2_2(.dout(w_dff_A_CZtdIhDC9_2),.din(w_dff_A_aZRWhOKy2_2),.clk(gclk));
	jdff dff_A_ojXkaW671_2(.dout(w_dff_A_aZRWhOKy2_2),.din(w_dff_A_ojXkaW671_2),.clk(gclk));
	jdff dff_A_AOFrt0zn7_2(.dout(w_dff_A_ojXkaW671_2),.din(w_dff_A_AOFrt0zn7_2),.clk(gclk));
	jdff dff_A_jsnuzbgw6_2(.dout(w_dff_A_AOFrt0zn7_2),.din(w_dff_A_jsnuzbgw6_2),.clk(gclk));
	jdff dff_A_qrpZZJsb1_2(.dout(w_dff_A_jsnuzbgw6_2),.din(w_dff_A_qrpZZJsb1_2),.clk(gclk));
	jdff dff_B_aEag40On6_0(.din(n163),.dout(w_dff_B_aEag40On6_0),.clk(gclk));
	jdff dff_A_JFe41pC52_0(.dout(w_n126_0[0]),.din(w_dff_A_JFe41pC52_0),.clk(gclk));
	jdff dff_A_TpGTez5Y7_0(.dout(w_dff_A_JFe41pC52_0),.din(w_dff_A_TpGTez5Y7_0),.clk(gclk));
	jdff dff_A_LzW34qYD2_0(.dout(w_dff_A_TpGTez5Y7_0),.din(w_dff_A_LzW34qYD2_0),.clk(gclk));
	jdff dff_A_kjw3uN572_0(.dout(w_dff_A_LzW34qYD2_0),.din(w_dff_A_kjw3uN572_0),.clk(gclk));
	jdff dff_A_8d4fuzZb7_0(.dout(w_dff_A_kjw3uN572_0),.din(w_dff_A_8d4fuzZb7_0),.clk(gclk));
	jdff dff_A_KKZrZLki5_1(.dout(w_n117_0[1]),.din(w_dff_A_KKZrZLki5_1),.clk(gclk));
	jdff dff_A_DwFv3ibl3_0(.dout(w_Gid5_0[0]),.din(w_dff_A_DwFv3ibl3_0),.clk(gclk));
	jdff dff_A_y9kXhS3C8_0(.dout(w_dff_A_DwFv3ibl3_0),.din(w_dff_A_y9kXhS3C8_0),.clk(gclk));
	jdff dff_A_lFhZsWmk6_0(.dout(w_dff_A_y9kXhS3C8_0),.din(w_dff_A_lFhZsWmk6_0),.clk(gclk));
	jdff dff_A_9qWbDexY4_0(.dout(w_dff_A_lFhZsWmk6_0),.din(w_dff_A_9qWbDexY4_0),.clk(gclk));
	jdff dff_A_MB0ROdsr3_0(.dout(w_dff_A_9qWbDexY4_0),.din(w_dff_A_MB0ROdsr3_0),.clk(gclk));
	jdff dff_A_IqMyPzKM5_0(.dout(w_dff_A_MB0ROdsr3_0),.din(w_dff_A_IqMyPzKM5_0),.clk(gclk));
	jdff dff_A_vMPiKgwa6_0(.dout(w_dff_A_IqMyPzKM5_0),.din(w_dff_A_vMPiKgwa6_0),.clk(gclk));
	jdff dff_A_AJ1bS1Tf2_0(.dout(w_dff_A_vMPiKgwa6_0),.din(w_dff_A_AJ1bS1Tf2_0),.clk(gclk));
	jdff dff_A_gmCKC0tQ3_0(.dout(w_dff_A_AJ1bS1Tf2_0),.din(w_dff_A_gmCKC0tQ3_0),.clk(gclk));
	jdff dff_A_e6qHfjer3_0(.dout(w_dff_A_gmCKC0tQ3_0),.din(w_dff_A_e6qHfjer3_0),.clk(gclk));
	jdff dff_A_hCwiAIeo8_0(.dout(w_Gid1_0[0]),.din(w_dff_A_hCwiAIeo8_0),.clk(gclk));
	jdff dff_A_OSZBgw5c7_0(.dout(w_dff_A_hCwiAIeo8_0),.din(w_dff_A_OSZBgw5c7_0),.clk(gclk));
	jdff dff_A_MBBxGDym4_0(.dout(w_dff_A_OSZBgw5c7_0),.din(w_dff_A_MBBxGDym4_0),.clk(gclk));
	jdff dff_A_4Vp2CxC63_0(.dout(w_dff_A_MBBxGDym4_0),.din(w_dff_A_4Vp2CxC63_0),.clk(gclk));
	jdff dff_A_sFeDdliz6_0(.dout(w_dff_A_4Vp2CxC63_0),.din(w_dff_A_sFeDdliz6_0),.clk(gclk));
	jdff dff_A_aIeU2GuI8_0(.dout(w_dff_A_sFeDdliz6_0),.din(w_dff_A_aIeU2GuI8_0),.clk(gclk));
	jdff dff_A_VmK0hjed0_0(.dout(w_dff_A_aIeU2GuI8_0),.din(w_dff_A_VmK0hjed0_0),.clk(gclk));
	jdff dff_A_2yHW8bBP8_0(.dout(w_dff_A_VmK0hjed0_0),.din(w_dff_A_2yHW8bBP8_0),.clk(gclk));
	jdff dff_A_Rx7o7aBk2_0(.dout(w_dff_A_2yHW8bBP8_0),.din(w_dff_A_Rx7o7aBk2_0),.clk(gclk));
	jdff dff_A_xyrjiOJf7_0(.dout(w_dff_A_Rx7o7aBk2_0),.din(w_dff_A_xyrjiOJf7_0),.clk(gclk));
	jdff dff_A_iR1kW9WG3_0(.dout(w_Gid13_0[0]),.din(w_dff_A_iR1kW9WG3_0),.clk(gclk));
	jdff dff_A_15ngu5GP5_0(.dout(w_dff_A_iR1kW9WG3_0),.din(w_dff_A_15ngu5GP5_0),.clk(gclk));
	jdff dff_A_C9FZG8Ob2_0(.dout(w_dff_A_15ngu5GP5_0),.din(w_dff_A_C9FZG8Ob2_0),.clk(gclk));
	jdff dff_A_zapEGAJP3_0(.dout(w_dff_A_C9FZG8Ob2_0),.din(w_dff_A_zapEGAJP3_0),.clk(gclk));
	jdff dff_A_zYTxt18W7_0(.dout(w_dff_A_zapEGAJP3_0),.din(w_dff_A_zYTxt18W7_0),.clk(gclk));
	jdff dff_A_Rav4cdvG2_0(.dout(w_dff_A_zYTxt18W7_0),.din(w_dff_A_Rav4cdvG2_0),.clk(gclk));
	jdff dff_A_EDNiREqN0_0(.dout(w_dff_A_Rav4cdvG2_0),.din(w_dff_A_EDNiREqN0_0),.clk(gclk));
	jdff dff_A_T80GeMZf3_0(.dout(w_dff_A_EDNiREqN0_0),.din(w_dff_A_T80GeMZf3_0),.clk(gclk));
	jdff dff_A_jVCDhH9e1_0(.dout(w_dff_A_T80GeMZf3_0),.din(w_dff_A_jVCDhH9e1_0),.clk(gclk));
	jdff dff_A_e19BsMgq7_0(.dout(w_dff_A_jVCDhH9e1_0),.din(w_dff_A_e19BsMgq7_0),.clk(gclk));
	jdff dff_A_d9kmoeXH9_0(.dout(w_Gid9_0[0]),.din(w_dff_A_d9kmoeXH9_0),.clk(gclk));
	jdff dff_A_DEuaYAYn5_0(.dout(w_dff_A_d9kmoeXH9_0),.din(w_dff_A_DEuaYAYn5_0),.clk(gclk));
	jdff dff_A_otYRCJkc9_0(.dout(w_dff_A_DEuaYAYn5_0),.din(w_dff_A_otYRCJkc9_0),.clk(gclk));
	jdff dff_A_ISGge4cv8_0(.dout(w_dff_A_otYRCJkc9_0),.din(w_dff_A_ISGge4cv8_0),.clk(gclk));
	jdff dff_A_Izc7Bs5L3_0(.dout(w_dff_A_ISGge4cv8_0),.din(w_dff_A_Izc7Bs5L3_0),.clk(gclk));
	jdff dff_A_M5JbCvzC7_0(.dout(w_dff_A_Izc7Bs5L3_0),.din(w_dff_A_M5JbCvzC7_0),.clk(gclk));
	jdff dff_A_lIWeYeRn9_0(.dout(w_dff_A_M5JbCvzC7_0),.din(w_dff_A_lIWeYeRn9_0),.clk(gclk));
	jdff dff_A_9mQzmulA3_0(.dout(w_dff_A_lIWeYeRn9_0),.din(w_dff_A_9mQzmulA3_0),.clk(gclk));
	jdff dff_A_Nw1WuOBJ4_0(.dout(w_dff_A_9mQzmulA3_0),.din(w_dff_A_Nw1WuOBJ4_0),.clk(gclk));
	jdff dff_A_BbKjK4CH4_0(.dout(w_dff_A_Nw1WuOBJ4_0),.din(w_dff_A_BbKjK4CH4_0),.clk(gclk));
	jdff dff_A_fwCw01320_1(.dout(w_n76_0[1]),.din(w_dff_A_fwCw01320_1),.clk(gclk));
	jdff dff_A_WawC5gE02_0(.dout(w_Gid4_0[0]),.din(w_dff_A_WawC5gE02_0),.clk(gclk));
	jdff dff_A_XBA1D4Hs8_0(.dout(w_dff_A_WawC5gE02_0),.din(w_dff_A_XBA1D4Hs8_0),.clk(gclk));
	jdff dff_A_abPV91rE8_0(.dout(w_dff_A_XBA1D4Hs8_0),.din(w_dff_A_abPV91rE8_0),.clk(gclk));
	jdff dff_A_uddMyPP02_0(.dout(w_dff_A_abPV91rE8_0),.din(w_dff_A_uddMyPP02_0),.clk(gclk));
	jdff dff_A_2E2xC8s41_0(.dout(w_dff_A_uddMyPP02_0),.din(w_dff_A_2E2xC8s41_0),.clk(gclk));
	jdff dff_A_dEpawunY5_0(.dout(w_dff_A_2E2xC8s41_0),.din(w_dff_A_dEpawunY5_0),.clk(gclk));
	jdff dff_A_jZY79jdm1_0(.dout(w_dff_A_dEpawunY5_0),.din(w_dff_A_jZY79jdm1_0),.clk(gclk));
	jdff dff_A_DqkO5rdd9_0(.dout(w_dff_A_jZY79jdm1_0),.din(w_dff_A_DqkO5rdd9_0),.clk(gclk));
	jdff dff_A_vQT2H2Bo2_0(.dout(w_dff_A_DqkO5rdd9_0),.din(w_dff_A_vQT2H2Bo2_0),.clk(gclk));
	jdff dff_A_yvg1r0oY8_0(.dout(w_dff_A_vQT2H2Bo2_0),.din(w_dff_A_yvg1r0oY8_0),.clk(gclk));
	jdff dff_A_M9JpT3z83_0(.dout(w_Gid0_0[0]),.din(w_dff_A_M9JpT3z83_0),.clk(gclk));
	jdff dff_A_iA9wfDyN9_0(.dout(w_dff_A_M9JpT3z83_0),.din(w_dff_A_iA9wfDyN9_0),.clk(gclk));
	jdff dff_A_PUnlEag12_0(.dout(w_dff_A_iA9wfDyN9_0),.din(w_dff_A_PUnlEag12_0),.clk(gclk));
	jdff dff_A_nZLuvCrW7_0(.dout(w_dff_A_PUnlEag12_0),.din(w_dff_A_nZLuvCrW7_0),.clk(gclk));
	jdff dff_A_nawXBPD00_0(.dout(w_dff_A_nZLuvCrW7_0),.din(w_dff_A_nawXBPD00_0),.clk(gclk));
	jdff dff_A_FNnHyjCW0_0(.dout(w_dff_A_nawXBPD00_0),.din(w_dff_A_FNnHyjCW0_0),.clk(gclk));
	jdff dff_A_2MM5LQ538_0(.dout(w_dff_A_FNnHyjCW0_0),.din(w_dff_A_2MM5LQ538_0),.clk(gclk));
	jdff dff_A_TG2AqP2S5_0(.dout(w_dff_A_2MM5LQ538_0),.din(w_dff_A_TG2AqP2S5_0),.clk(gclk));
	jdff dff_A_lHCVdao89_0(.dout(w_dff_A_TG2AqP2S5_0),.din(w_dff_A_lHCVdao89_0),.clk(gclk));
	jdff dff_A_sa4OWoUW2_0(.dout(w_dff_A_lHCVdao89_0),.din(w_dff_A_sa4OWoUW2_0),.clk(gclk));
	jdff dff_A_At90bml85_0(.dout(w_Gid12_0[0]),.din(w_dff_A_At90bml85_0),.clk(gclk));
	jdff dff_A_g99eVEKr9_0(.dout(w_dff_A_At90bml85_0),.din(w_dff_A_g99eVEKr9_0),.clk(gclk));
	jdff dff_A_detPl1vj2_0(.dout(w_dff_A_g99eVEKr9_0),.din(w_dff_A_detPl1vj2_0),.clk(gclk));
	jdff dff_A_BrP1Za891_0(.dout(w_dff_A_detPl1vj2_0),.din(w_dff_A_BrP1Za891_0),.clk(gclk));
	jdff dff_A_L1S432cR1_0(.dout(w_dff_A_BrP1Za891_0),.din(w_dff_A_L1S432cR1_0),.clk(gclk));
	jdff dff_A_FYeeoov96_0(.dout(w_dff_A_L1S432cR1_0),.din(w_dff_A_FYeeoov96_0),.clk(gclk));
	jdff dff_A_rJWz5WVA5_0(.dout(w_dff_A_FYeeoov96_0),.din(w_dff_A_rJWz5WVA5_0),.clk(gclk));
	jdff dff_A_YaCx97Sw6_0(.dout(w_dff_A_rJWz5WVA5_0),.din(w_dff_A_YaCx97Sw6_0),.clk(gclk));
	jdff dff_A_HqSsxoLx5_0(.dout(w_dff_A_YaCx97Sw6_0),.din(w_dff_A_HqSsxoLx5_0),.clk(gclk));
	jdff dff_A_VnYVtnKV4_0(.dout(w_dff_A_HqSsxoLx5_0),.din(w_dff_A_VnYVtnKV4_0),.clk(gclk));
	jdff dff_A_ekJUKZR78_0(.dout(w_Gid8_0[0]),.din(w_dff_A_ekJUKZR78_0),.clk(gclk));
	jdff dff_A_JFzEI21U0_0(.dout(w_dff_A_ekJUKZR78_0),.din(w_dff_A_JFzEI21U0_0),.clk(gclk));
	jdff dff_A_K00kppmn0_0(.dout(w_dff_A_JFzEI21U0_0),.din(w_dff_A_K00kppmn0_0),.clk(gclk));
	jdff dff_A_T7piVlkW3_0(.dout(w_dff_A_K00kppmn0_0),.din(w_dff_A_T7piVlkW3_0),.clk(gclk));
	jdff dff_A_mzTopdh82_0(.dout(w_dff_A_T7piVlkW3_0),.din(w_dff_A_mzTopdh82_0),.clk(gclk));
	jdff dff_A_ZdGf52bd0_0(.dout(w_dff_A_mzTopdh82_0),.din(w_dff_A_ZdGf52bd0_0),.clk(gclk));
	jdff dff_A_TGwAMCYX6_0(.dout(w_dff_A_ZdGf52bd0_0),.din(w_dff_A_TGwAMCYX6_0),.clk(gclk));
	jdff dff_A_vIRHxb962_0(.dout(w_dff_A_TGwAMCYX6_0),.din(w_dff_A_vIRHxb962_0),.clk(gclk));
	jdff dff_A_uAKChElf5_0(.dout(w_dff_A_vIRHxb962_0),.din(w_dff_A_uAKChElf5_0),.clk(gclk));
	jdff dff_A_tDxgDZ2d5_0(.dout(w_dff_A_uAKChElf5_0),.din(w_dff_A_tDxgDZ2d5_0),.clk(gclk));
	jdff dff_B_T5XMTz9U6_2(.din(n242),.dout(w_dff_B_T5XMTz9U6_2),.clk(gclk));
	jdff dff_B_oWdEUL8r0_2(.din(w_dff_B_T5XMTz9U6_2),.dout(w_dff_B_oWdEUL8r0_2),.clk(gclk));
	jdff dff_B_PlkuSVZL3_2(.din(w_dff_B_oWdEUL8r0_2),.dout(w_dff_B_PlkuSVZL3_2),.clk(gclk));
	jdff dff_B_ieGEsqOi6_2(.din(w_dff_B_PlkuSVZL3_2),.dout(w_dff_B_ieGEsqOi6_2),.clk(gclk));
	jdff dff_A_tsBNwBtG2_0(.dout(w_Gid6_0[0]),.din(w_dff_A_tsBNwBtG2_0),.clk(gclk));
	jdff dff_A_Puxh7rF57_0(.dout(w_dff_A_tsBNwBtG2_0),.din(w_dff_A_Puxh7rF57_0),.clk(gclk));
	jdff dff_A_oBVWHtSO2_0(.dout(w_dff_A_Puxh7rF57_0),.din(w_dff_A_oBVWHtSO2_0),.clk(gclk));
	jdff dff_A_nMoVTGIG1_0(.dout(w_dff_A_oBVWHtSO2_0),.din(w_dff_A_nMoVTGIG1_0),.clk(gclk));
	jdff dff_A_dORseiiV9_0(.dout(w_dff_A_nMoVTGIG1_0),.din(w_dff_A_dORseiiV9_0),.clk(gclk));
	jdff dff_A_eZQeiVmw7_0(.dout(w_dff_A_dORseiiV9_0),.din(w_dff_A_eZQeiVmw7_0),.clk(gclk));
	jdff dff_A_tnkVno0X6_0(.dout(w_dff_A_eZQeiVmw7_0),.din(w_dff_A_tnkVno0X6_0),.clk(gclk));
	jdff dff_A_GHRCWbpx7_0(.dout(w_dff_A_tnkVno0X6_0),.din(w_dff_A_GHRCWbpx7_0),.clk(gclk));
	jdff dff_A_XZ6qsNRu5_0(.dout(w_dff_A_GHRCWbpx7_0),.din(w_dff_A_XZ6qsNRu5_0),.clk(gclk));
	jdff dff_A_EMPIVIqJ8_0(.dout(w_dff_A_XZ6qsNRu5_0),.din(w_dff_A_EMPIVIqJ8_0),.clk(gclk));
	jdff dff_A_f20EweG96_0(.dout(w_Gid2_0[0]),.din(w_dff_A_f20EweG96_0),.clk(gclk));
	jdff dff_A_w2R96mvP2_0(.dout(w_dff_A_f20EweG96_0),.din(w_dff_A_w2R96mvP2_0),.clk(gclk));
	jdff dff_A_DbO3wBK08_0(.dout(w_dff_A_w2R96mvP2_0),.din(w_dff_A_DbO3wBK08_0),.clk(gclk));
	jdff dff_A_oAVtPxxh4_0(.dout(w_dff_A_DbO3wBK08_0),.din(w_dff_A_oAVtPxxh4_0),.clk(gclk));
	jdff dff_A_XTq4DLOc6_0(.dout(w_dff_A_oAVtPxxh4_0),.din(w_dff_A_XTq4DLOc6_0),.clk(gclk));
	jdff dff_A_fV5EdQbm6_0(.dout(w_dff_A_XTq4DLOc6_0),.din(w_dff_A_fV5EdQbm6_0),.clk(gclk));
	jdff dff_A_rMMEiVBk4_0(.dout(w_dff_A_fV5EdQbm6_0),.din(w_dff_A_rMMEiVBk4_0),.clk(gclk));
	jdff dff_A_AyDRLz6W7_0(.dout(w_dff_A_rMMEiVBk4_0),.din(w_dff_A_AyDRLz6W7_0),.clk(gclk));
	jdff dff_A_el3y4pEh1_0(.dout(w_dff_A_AyDRLz6W7_0),.din(w_dff_A_el3y4pEh1_0),.clk(gclk));
	jdff dff_A_gj6iAReM1_0(.dout(w_dff_A_el3y4pEh1_0),.din(w_dff_A_gj6iAReM1_0),.clk(gclk));
	jdff dff_A_gSpRsrLF3_0(.dout(w_Gid14_0[0]),.din(w_dff_A_gSpRsrLF3_0),.clk(gclk));
	jdff dff_A_QZC074961_0(.dout(w_dff_A_gSpRsrLF3_0),.din(w_dff_A_QZC074961_0),.clk(gclk));
	jdff dff_A_dKyqDLTN5_0(.dout(w_dff_A_QZC074961_0),.din(w_dff_A_dKyqDLTN5_0),.clk(gclk));
	jdff dff_A_Lvzh2QxO8_0(.dout(w_dff_A_dKyqDLTN5_0),.din(w_dff_A_Lvzh2QxO8_0),.clk(gclk));
	jdff dff_A_bPr8US7I1_0(.dout(w_dff_A_Lvzh2QxO8_0),.din(w_dff_A_bPr8US7I1_0),.clk(gclk));
	jdff dff_A_JSfKqfWp1_0(.dout(w_dff_A_bPr8US7I1_0),.din(w_dff_A_JSfKqfWp1_0),.clk(gclk));
	jdff dff_A_oSOxZfVn1_0(.dout(w_dff_A_JSfKqfWp1_0),.din(w_dff_A_oSOxZfVn1_0),.clk(gclk));
	jdff dff_A_9K6Bi0Ku2_0(.dout(w_dff_A_oSOxZfVn1_0),.din(w_dff_A_9K6Bi0Ku2_0),.clk(gclk));
	jdff dff_A_6nhii6ug1_0(.dout(w_dff_A_9K6Bi0Ku2_0),.din(w_dff_A_6nhii6ug1_0),.clk(gclk));
	jdff dff_A_NUSHHJdk6_0(.dout(w_dff_A_6nhii6ug1_0),.din(w_dff_A_NUSHHJdk6_0),.clk(gclk));
	jdff dff_A_BODOr6t57_0(.dout(w_Gid10_0[0]),.din(w_dff_A_BODOr6t57_0),.clk(gclk));
	jdff dff_A_QWwRfLJ86_0(.dout(w_dff_A_BODOr6t57_0),.din(w_dff_A_QWwRfLJ86_0),.clk(gclk));
	jdff dff_A_J3oXYHUn0_0(.dout(w_dff_A_QWwRfLJ86_0),.din(w_dff_A_J3oXYHUn0_0),.clk(gclk));
	jdff dff_A_UXGuyqaF2_0(.dout(w_dff_A_J3oXYHUn0_0),.din(w_dff_A_UXGuyqaF2_0),.clk(gclk));
	jdff dff_A_vNMhoonh0_0(.dout(w_dff_A_UXGuyqaF2_0),.din(w_dff_A_vNMhoonh0_0),.clk(gclk));
	jdff dff_A_6VrUZnzh8_0(.dout(w_dff_A_vNMhoonh0_0),.din(w_dff_A_6VrUZnzh8_0),.clk(gclk));
	jdff dff_A_M72686594_0(.dout(w_dff_A_6VrUZnzh8_0),.din(w_dff_A_M72686594_0),.clk(gclk));
	jdff dff_A_7TGCgdXv9_0(.dout(w_dff_A_M72686594_0),.din(w_dff_A_7TGCgdXv9_0),.clk(gclk));
	jdff dff_A_qASn3qVF8_0(.dout(w_dff_A_7TGCgdXv9_0),.din(w_dff_A_qASn3qVF8_0),.clk(gclk));
	jdff dff_A_IqBfVVeA8_0(.dout(w_dff_A_qASn3qVF8_0),.din(w_dff_A_IqBfVVeA8_0),.clk(gclk));
	jdff dff_A_y8TAGmVZ6_0(.dout(w_Gid17_0[0]),.din(w_dff_A_y8TAGmVZ6_0),.clk(gclk));
	jdff dff_A_Gdi3fesB0_0(.dout(w_dff_A_y8TAGmVZ6_0),.din(w_dff_A_Gdi3fesB0_0),.clk(gclk));
	jdff dff_A_PT0aD6DI8_0(.dout(w_dff_A_Gdi3fesB0_0),.din(w_dff_A_PT0aD6DI8_0),.clk(gclk));
	jdff dff_A_5FgW6ieE7_0(.dout(w_dff_A_PT0aD6DI8_0),.din(w_dff_A_5FgW6ieE7_0),.clk(gclk));
	jdff dff_A_lSrRblMA3_0(.dout(w_dff_A_5FgW6ieE7_0),.din(w_dff_A_lSrRblMA3_0),.clk(gclk));
	jdff dff_A_lOTExVOr3_0(.dout(w_dff_A_lSrRblMA3_0),.din(w_dff_A_lOTExVOr3_0),.clk(gclk));
	jdff dff_A_LN9IRyV51_0(.dout(w_dff_A_lOTExVOr3_0),.din(w_dff_A_LN9IRyV51_0),.clk(gclk));
	jdff dff_A_OrXtFU6a7_0(.dout(w_dff_A_LN9IRyV51_0),.din(w_dff_A_OrXtFU6a7_0),.clk(gclk));
	jdff dff_A_tz2LsV2S1_0(.dout(w_dff_A_OrXtFU6a7_0),.din(w_dff_A_tz2LsV2S1_0),.clk(gclk));
	jdff dff_A_a8r5XbTc3_0(.dout(w_dff_A_tz2LsV2S1_0),.din(w_dff_A_a8r5XbTc3_0),.clk(gclk));
	jdff dff_A_le8cFb526_0(.dout(w_dff_A_a8r5XbTc3_0),.din(w_dff_A_le8cFb526_0),.clk(gclk));
	jdff dff_A_QLpOZsYA9_0(.dout(w_Gid16_0[0]),.din(w_dff_A_QLpOZsYA9_0),.clk(gclk));
	jdff dff_A_ieqTNxBs4_0(.dout(w_dff_A_QLpOZsYA9_0),.din(w_dff_A_ieqTNxBs4_0),.clk(gclk));
	jdff dff_A_qQDJj8Dw7_0(.dout(w_dff_A_ieqTNxBs4_0),.din(w_dff_A_qQDJj8Dw7_0),.clk(gclk));
	jdff dff_A_3YDIIdKx5_0(.dout(w_dff_A_qQDJj8Dw7_0),.din(w_dff_A_3YDIIdKx5_0),.clk(gclk));
	jdff dff_A_zp4KvbtE6_0(.dout(w_dff_A_3YDIIdKx5_0),.din(w_dff_A_zp4KvbtE6_0),.clk(gclk));
	jdff dff_A_moDb1xJL7_0(.dout(w_dff_A_zp4KvbtE6_0),.din(w_dff_A_moDb1xJL7_0),.clk(gclk));
	jdff dff_A_BfHPJgp10_0(.dout(w_dff_A_moDb1xJL7_0),.din(w_dff_A_BfHPJgp10_0),.clk(gclk));
	jdff dff_A_H0idetRW4_0(.dout(w_dff_A_BfHPJgp10_0),.din(w_dff_A_H0idetRW4_0),.clk(gclk));
	jdff dff_A_1Hq53zEO5_0(.dout(w_dff_A_H0idetRW4_0),.din(w_dff_A_1Hq53zEO5_0),.clk(gclk));
	jdff dff_A_GkSIZpXT0_0(.dout(w_dff_A_1Hq53zEO5_0),.din(w_dff_A_GkSIZpXT0_0),.clk(gclk));
	jdff dff_A_MjREwZlV9_0(.dout(w_dff_A_GkSIZpXT0_0),.din(w_dff_A_MjREwZlV9_0),.clk(gclk));
	jdff dff_A_Ltv5IHHs5_0(.dout(w_Gid19_0[0]),.din(w_dff_A_Ltv5IHHs5_0),.clk(gclk));
	jdff dff_A_0LWr4iEd8_0(.dout(w_dff_A_Ltv5IHHs5_0),.din(w_dff_A_0LWr4iEd8_0),.clk(gclk));
	jdff dff_A_BvQkiO895_0(.dout(w_dff_A_0LWr4iEd8_0),.din(w_dff_A_BvQkiO895_0),.clk(gclk));
	jdff dff_A_K26Bpe4a1_0(.dout(w_dff_A_BvQkiO895_0),.din(w_dff_A_K26Bpe4a1_0),.clk(gclk));
	jdff dff_A_gTdOFDtA9_0(.dout(w_dff_A_K26Bpe4a1_0),.din(w_dff_A_gTdOFDtA9_0),.clk(gclk));
	jdff dff_A_Ty2NVLIk0_0(.dout(w_dff_A_gTdOFDtA9_0),.din(w_dff_A_Ty2NVLIk0_0),.clk(gclk));
	jdff dff_A_3a69GPrT9_0(.dout(w_dff_A_Ty2NVLIk0_0),.din(w_dff_A_3a69GPrT9_0),.clk(gclk));
	jdff dff_A_sQcirZQE4_0(.dout(w_dff_A_3a69GPrT9_0),.din(w_dff_A_sQcirZQE4_0),.clk(gclk));
	jdff dff_A_9D5pu5wK5_0(.dout(w_dff_A_sQcirZQE4_0),.din(w_dff_A_9D5pu5wK5_0),.clk(gclk));
	jdff dff_A_YhsIfzh68_0(.dout(w_dff_A_9D5pu5wK5_0),.din(w_dff_A_YhsIfzh68_0),.clk(gclk));
	jdff dff_A_mt8WhnID8_0(.dout(w_dff_A_YhsIfzh68_0),.din(w_dff_A_mt8WhnID8_0),.clk(gclk));
	jdff dff_A_vKR8mQzE2_0(.dout(w_Gid18_0[0]),.din(w_dff_A_vKR8mQzE2_0),.clk(gclk));
	jdff dff_A_ADdHF0cn6_0(.dout(w_dff_A_vKR8mQzE2_0),.din(w_dff_A_ADdHF0cn6_0),.clk(gclk));
	jdff dff_A_yxAveYNq4_0(.dout(w_dff_A_ADdHF0cn6_0),.din(w_dff_A_yxAveYNq4_0),.clk(gclk));
	jdff dff_A_b3bpUASY0_0(.dout(w_dff_A_yxAveYNq4_0),.din(w_dff_A_b3bpUASY0_0),.clk(gclk));
	jdff dff_A_NIWtCpyz7_0(.dout(w_dff_A_b3bpUASY0_0),.din(w_dff_A_NIWtCpyz7_0),.clk(gclk));
	jdff dff_A_5VKUJ0p35_0(.dout(w_dff_A_NIWtCpyz7_0),.din(w_dff_A_5VKUJ0p35_0),.clk(gclk));
	jdff dff_A_AGcqx0bD6_0(.dout(w_dff_A_5VKUJ0p35_0),.din(w_dff_A_AGcqx0bD6_0),.clk(gclk));
	jdff dff_A_Wjs34HUv3_0(.dout(w_dff_A_AGcqx0bD6_0),.din(w_dff_A_Wjs34HUv3_0),.clk(gclk));
	jdff dff_A_LGdOoEMi9_0(.dout(w_dff_A_Wjs34HUv3_0),.din(w_dff_A_LGdOoEMi9_0),.clk(gclk));
	jdff dff_A_JlPhArOH3_0(.dout(w_dff_A_LGdOoEMi9_0),.din(w_dff_A_JlPhArOH3_0),.clk(gclk));
	jdff dff_A_KfyVvEv86_0(.dout(w_dff_A_JlPhArOH3_0),.din(w_dff_A_KfyVvEv86_0),.clk(gclk));
	jdff dff_A_ZJuoWG3b4_0(.dout(w_n136_0[0]),.din(w_dff_A_ZJuoWG3b4_0),.clk(gclk));
	jdff dff_A_wATpigAW5_0(.dout(w_Gid25_0[0]),.din(w_dff_A_wATpigAW5_0),.clk(gclk));
	jdff dff_A_vzi6ZsXL0_0(.dout(w_dff_A_wATpigAW5_0),.din(w_dff_A_vzi6ZsXL0_0),.clk(gclk));
	jdff dff_A_kEeY6YA29_0(.dout(w_dff_A_vzi6ZsXL0_0),.din(w_dff_A_kEeY6YA29_0),.clk(gclk));
	jdff dff_A_itw6IJbQ0_0(.dout(w_dff_A_kEeY6YA29_0),.din(w_dff_A_itw6IJbQ0_0),.clk(gclk));
	jdff dff_A_QpW6nWUx4_0(.dout(w_dff_A_itw6IJbQ0_0),.din(w_dff_A_QpW6nWUx4_0),.clk(gclk));
	jdff dff_A_acs7cH5E5_0(.dout(w_dff_A_QpW6nWUx4_0),.din(w_dff_A_acs7cH5E5_0),.clk(gclk));
	jdff dff_A_WpLjAqVQ7_0(.dout(w_dff_A_acs7cH5E5_0),.din(w_dff_A_WpLjAqVQ7_0),.clk(gclk));
	jdff dff_A_ZVjywUw11_0(.dout(w_dff_A_WpLjAqVQ7_0),.din(w_dff_A_ZVjywUw11_0),.clk(gclk));
	jdff dff_A_wDcYrBrj9_0(.dout(w_dff_A_ZVjywUw11_0),.din(w_dff_A_wDcYrBrj9_0),.clk(gclk));
	jdff dff_A_8JOkLVhU6_0(.dout(w_dff_A_wDcYrBrj9_0),.din(w_dff_A_8JOkLVhU6_0),.clk(gclk));
	jdff dff_A_fqtUejUg2_0(.dout(w_dff_A_8JOkLVhU6_0),.din(w_dff_A_fqtUejUg2_0),.clk(gclk));
	jdff dff_A_cTlgOsAY7_0(.dout(w_Gid24_0[0]),.din(w_dff_A_cTlgOsAY7_0),.clk(gclk));
	jdff dff_A_5NKyHsij6_0(.dout(w_dff_A_cTlgOsAY7_0),.din(w_dff_A_5NKyHsij6_0),.clk(gclk));
	jdff dff_A_8B6oZxSU6_0(.dout(w_dff_A_5NKyHsij6_0),.din(w_dff_A_8B6oZxSU6_0),.clk(gclk));
	jdff dff_A_dWpCOdiJ9_0(.dout(w_dff_A_8B6oZxSU6_0),.din(w_dff_A_dWpCOdiJ9_0),.clk(gclk));
	jdff dff_A_eSunXmXI9_0(.dout(w_dff_A_dWpCOdiJ9_0),.din(w_dff_A_eSunXmXI9_0),.clk(gclk));
	jdff dff_A_Re4YqTwz5_0(.dout(w_dff_A_eSunXmXI9_0),.din(w_dff_A_Re4YqTwz5_0),.clk(gclk));
	jdff dff_A_37wqzGLc4_0(.dout(w_dff_A_Re4YqTwz5_0),.din(w_dff_A_37wqzGLc4_0),.clk(gclk));
	jdff dff_A_O4HIr8ym7_0(.dout(w_dff_A_37wqzGLc4_0),.din(w_dff_A_O4HIr8ym7_0),.clk(gclk));
	jdff dff_A_0W2MZB119_0(.dout(w_dff_A_O4HIr8ym7_0),.din(w_dff_A_0W2MZB119_0),.clk(gclk));
	jdff dff_A_mgt7igOC7_0(.dout(w_dff_A_0W2MZB119_0),.din(w_dff_A_mgt7igOC7_0),.clk(gclk));
	jdff dff_A_jGuG0zO77_0(.dout(w_dff_A_mgt7igOC7_0),.din(w_dff_A_jGuG0zO77_0),.clk(gclk));
	jdff dff_A_XxKcmYcI6_0(.dout(w_Gid27_0[0]),.din(w_dff_A_XxKcmYcI6_0),.clk(gclk));
	jdff dff_A_LAgFhPTz4_0(.dout(w_dff_A_XxKcmYcI6_0),.din(w_dff_A_LAgFhPTz4_0),.clk(gclk));
	jdff dff_A_UHOrkYer2_0(.dout(w_dff_A_LAgFhPTz4_0),.din(w_dff_A_UHOrkYer2_0),.clk(gclk));
	jdff dff_A_xoOpm9Gi2_0(.dout(w_dff_A_UHOrkYer2_0),.din(w_dff_A_xoOpm9Gi2_0),.clk(gclk));
	jdff dff_A_Y1Mkm3kC6_0(.dout(w_dff_A_xoOpm9Gi2_0),.din(w_dff_A_Y1Mkm3kC6_0),.clk(gclk));
	jdff dff_A_AqLVnBYc6_0(.dout(w_dff_A_Y1Mkm3kC6_0),.din(w_dff_A_AqLVnBYc6_0),.clk(gclk));
	jdff dff_A_qRvL5tm91_0(.dout(w_dff_A_AqLVnBYc6_0),.din(w_dff_A_qRvL5tm91_0),.clk(gclk));
	jdff dff_A_FScwOEWx9_0(.dout(w_dff_A_qRvL5tm91_0),.din(w_dff_A_FScwOEWx9_0),.clk(gclk));
	jdff dff_A_3bTLZVW48_0(.dout(w_dff_A_FScwOEWx9_0),.din(w_dff_A_3bTLZVW48_0),.clk(gclk));
	jdff dff_A_PErTobiK3_0(.dout(w_dff_A_3bTLZVW48_0),.din(w_dff_A_PErTobiK3_0),.clk(gclk));
	jdff dff_A_2hZ8NGte0_0(.dout(w_dff_A_PErTobiK3_0),.din(w_dff_A_2hZ8NGte0_0),.clk(gclk));
	jdff dff_A_HabnOg7g4_0(.dout(w_Gid26_0[0]),.din(w_dff_A_HabnOg7g4_0),.clk(gclk));
	jdff dff_A_VLgpElNv1_0(.dout(w_dff_A_HabnOg7g4_0),.din(w_dff_A_VLgpElNv1_0),.clk(gclk));
	jdff dff_A_krFr8OT08_0(.dout(w_dff_A_VLgpElNv1_0),.din(w_dff_A_krFr8OT08_0),.clk(gclk));
	jdff dff_A_kAvTY9CC9_0(.dout(w_dff_A_krFr8OT08_0),.din(w_dff_A_kAvTY9CC9_0),.clk(gclk));
	jdff dff_A_Zkqq8mmR9_0(.dout(w_dff_A_kAvTY9CC9_0),.din(w_dff_A_Zkqq8mmR9_0),.clk(gclk));
	jdff dff_A_cR7zXUpb8_0(.dout(w_dff_A_Zkqq8mmR9_0),.din(w_dff_A_cR7zXUpb8_0),.clk(gclk));
	jdff dff_A_65adcIcR0_0(.dout(w_dff_A_cR7zXUpb8_0),.din(w_dff_A_65adcIcR0_0),.clk(gclk));
	jdff dff_A_GHemA6K55_0(.dout(w_dff_A_65adcIcR0_0),.din(w_dff_A_GHemA6K55_0),.clk(gclk));
	jdff dff_A_1vLGFCsA4_0(.dout(w_dff_A_GHemA6K55_0),.din(w_dff_A_1vLGFCsA4_0),.clk(gclk));
	jdff dff_A_E4eC3xkc8_0(.dout(w_dff_A_1vLGFCsA4_0),.din(w_dff_A_E4eC3xkc8_0),.clk(gclk));
	jdff dff_A_4WZtkrDt4_0(.dout(w_dff_A_E4eC3xkc8_0),.din(w_dff_A_4WZtkrDt4_0),.clk(gclk));
	jdff dff_A_ShH3IoYz8_0(.dout(w_n147_0[0]),.din(w_dff_A_ShH3IoYz8_0),.clk(gclk));
	jdff dff_A_0txnnUVh5_0(.dout(w_dff_A_ShH3IoYz8_0),.din(w_dff_A_0txnnUVh5_0),.clk(gclk));
	jdff dff_A_iHsKkUgZ6_0(.dout(w_dff_A_0txnnUVh5_0),.din(w_dff_A_iHsKkUgZ6_0),.clk(gclk));
	jdff dff_A_uKUG5bvG9_0(.dout(w_dff_A_iHsKkUgZ6_0),.din(w_dff_A_uKUG5bvG9_0),.clk(gclk));
	jdff dff_A_Cr5cLS2T5_0(.dout(w_dff_A_uKUG5bvG9_0),.din(w_dff_A_Cr5cLS2T5_0),.clk(gclk));
	jdff dff_A_SzdnntIp3_0(.dout(w_Gid7_0[0]),.din(w_dff_A_SzdnntIp3_0),.clk(gclk));
	jdff dff_A_nEVbT2oS9_0(.dout(w_dff_A_SzdnntIp3_0),.din(w_dff_A_nEVbT2oS9_0),.clk(gclk));
	jdff dff_A_xMGmcRnX7_0(.dout(w_dff_A_nEVbT2oS9_0),.din(w_dff_A_xMGmcRnX7_0),.clk(gclk));
	jdff dff_A_WgSCMoXA9_0(.dout(w_dff_A_xMGmcRnX7_0),.din(w_dff_A_WgSCMoXA9_0),.clk(gclk));
	jdff dff_A_s4xXG9OR1_0(.dout(w_dff_A_WgSCMoXA9_0),.din(w_dff_A_s4xXG9OR1_0),.clk(gclk));
	jdff dff_A_G2xG24jo3_0(.dout(w_dff_A_s4xXG9OR1_0),.din(w_dff_A_G2xG24jo3_0),.clk(gclk));
	jdff dff_A_BmtKDlhN1_0(.dout(w_dff_A_G2xG24jo3_0),.din(w_dff_A_BmtKDlhN1_0),.clk(gclk));
	jdff dff_A_gVRjlR0a8_0(.dout(w_dff_A_BmtKDlhN1_0),.din(w_dff_A_gVRjlR0a8_0),.clk(gclk));
	jdff dff_A_n1TWzyVW1_0(.dout(w_dff_A_gVRjlR0a8_0),.din(w_dff_A_n1TWzyVW1_0),.clk(gclk));
	jdff dff_A_7TIpTwFc4_0(.dout(w_dff_A_n1TWzyVW1_0),.din(w_dff_A_7TIpTwFc4_0),.clk(gclk));
	jdff dff_A_YuU7x8F87_0(.dout(w_Gid3_0[0]),.din(w_dff_A_YuU7x8F87_0),.clk(gclk));
	jdff dff_A_6R0zsxVF9_0(.dout(w_dff_A_YuU7x8F87_0),.din(w_dff_A_6R0zsxVF9_0),.clk(gclk));
	jdff dff_A_xw6AtxjP1_0(.dout(w_dff_A_6R0zsxVF9_0),.din(w_dff_A_xw6AtxjP1_0),.clk(gclk));
	jdff dff_A_MnPrF0Qk5_0(.dout(w_dff_A_xw6AtxjP1_0),.din(w_dff_A_MnPrF0Qk5_0),.clk(gclk));
	jdff dff_A_yqqtw33N2_0(.dout(w_dff_A_MnPrF0Qk5_0),.din(w_dff_A_yqqtw33N2_0),.clk(gclk));
	jdff dff_A_GjgBXbrJ4_0(.dout(w_dff_A_yqqtw33N2_0),.din(w_dff_A_GjgBXbrJ4_0),.clk(gclk));
	jdff dff_A_Mmr638io0_0(.dout(w_dff_A_GjgBXbrJ4_0),.din(w_dff_A_Mmr638io0_0),.clk(gclk));
	jdff dff_A_KYF4qxz23_0(.dout(w_dff_A_Mmr638io0_0),.din(w_dff_A_KYF4qxz23_0),.clk(gclk));
	jdff dff_A_cq6iLv8R3_0(.dout(w_dff_A_KYF4qxz23_0),.din(w_dff_A_cq6iLv8R3_0),.clk(gclk));
	jdff dff_A_0eqBGbxx8_0(.dout(w_dff_A_cq6iLv8R3_0),.din(w_dff_A_0eqBGbxx8_0),.clk(gclk));
	jdff dff_A_OqiMJQrW8_0(.dout(w_Gid15_0[0]),.din(w_dff_A_OqiMJQrW8_0),.clk(gclk));
	jdff dff_A_Iv6qHPNr2_0(.dout(w_dff_A_OqiMJQrW8_0),.din(w_dff_A_Iv6qHPNr2_0),.clk(gclk));
	jdff dff_A_3wcrrLaR8_0(.dout(w_dff_A_Iv6qHPNr2_0),.din(w_dff_A_3wcrrLaR8_0),.clk(gclk));
	jdff dff_A_9yL4V7Y29_0(.dout(w_dff_A_3wcrrLaR8_0),.din(w_dff_A_9yL4V7Y29_0),.clk(gclk));
	jdff dff_A_cq0hTvsx5_0(.dout(w_dff_A_9yL4V7Y29_0),.din(w_dff_A_cq0hTvsx5_0),.clk(gclk));
	jdff dff_A_9Iv8Nqpw7_0(.dout(w_dff_A_cq0hTvsx5_0),.din(w_dff_A_9Iv8Nqpw7_0),.clk(gclk));
	jdff dff_A_qnkLrDhc8_0(.dout(w_dff_A_9Iv8Nqpw7_0),.din(w_dff_A_qnkLrDhc8_0),.clk(gclk));
	jdff dff_A_6S0Lt0No0_0(.dout(w_dff_A_qnkLrDhc8_0),.din(w_dff_A_6S0Lt0No0_0),.clk(gclk));
	jdff dff_A_e5VntDoQ3_0(.dout(w_dff_A_6S0Lt0No0_0),.din(w_dff_A_e5VntDoQ3_0),.clk(gclk));
	jdff dff_A_XTa2fve04_0(.dout(w_dff_A_e5VntDoQ3_0),.din(w_dff_A_XTa2fve04_0),.clk(gclk));
	jdff dff_A_GVpxtwUU3_0(.dout(w_Gid11_0[0]),.din(w_dff_A_GVpxtwUU3_0),.clk(gclk));
	jdff dff_A_8oVzv6NI7_0(.dout(w_dff_A_GVpxtwUU3_0),.din(w_dff_A_8oVzv6NI7_0),.clk(gclk));
	jdff dff_A_pJvjy3wE5_0(.dout(w_dff_A_8oVzv6NI7_0),.din(w_dff_A_pJvjy3wE5_0),.clk(gclk));
	jdff dff_A_NUjeNaXw5_0(.dout(w_dff_A_pJvjy3wE5_0),.din(w_dff_A_NUjeNaXw5_0),.clk(gclk));
	jdff dff_A_90dF8Ipt2_0(.dout(w_dff_A_NUjeNaXw5_0),.din(w_dff_A_90dF8Ipt2_0),.clk(gclk));
	jdff dff_A_cD2QuQWK5_0(.dout(w_dff_A_90dF8Ipt2_0),.din(w_dff_A_cD2QuQWK5_0),.clk(gclk));
	jdff dff_A_XESSd1qZ4_0(.dout(w_dff_A_cD2QuQWK5_0),.din(w_dff_A_XESSd1qZ4_0),.clk(gclk));
	jdff dff_A_hsz9WMop4_0(.dout(w_dff_A_XESSd1qZ4_0),.din(w_dff_A_hsz9WMop4_0),.clk(gclk));
	jdff dff_A_hQjAgRvx7_0(.dout(w_dff_A_hsz9WMop4_0),.din(w_dff_A_hQjAgRvx7_0),.clk(gclk));
	jdff dff_A_gYxrWJE52_0(.dout(w_dff_A_hQjAgRvx7_0),.din(w_dff_A_gYxrWJE52_0),.clk(gclk));
	jdff dff_A_jTdwQiEG0_0(.dout(w_Gid21_0[0]),.din(w_dff_A_jTdwQiEG0_0),.clk(gclk));
	jdff dff_A_0X6kJbZX4_0(.dout(w_dff_A_jTdwQiEG0_0),.din(w_dff_A_0X6kJbZX4_0),.clk(gclk));
	jdff dff_A_EdUY70hO3_0(.dout(w_dff_A_0X6kJbZX4_0),.din(w_dff_A_EdUY70hO3_0),.clk(gclk));
	jdff dff_A_CVbxJ1O45_0(.dout(w_dff_A_EdUY70hO3_0),.din(w_dff_A_CVbxJ1O45_0),.clk(gclk));
	jdff dff_A_gcui7y3n5_0(.dout(w_dff_A_CVbxJ1O45_0),.din(w_dff_A_gcui7y3n5_0),.clk(gclk));
	jdff dff_A_GVlw776V6_0(.dout(w_dff_A_gcui7y3n5_0),.din(w_dff_A_GVlw776V6_0),.clk(gclk));
	jdff dff_A_m6f3wyN56_0(.dout(w_dff_A_GVlw776V6_0),.din(w_dff_A_m6f3wyN56_0),.clk(gclk));
	jdff dff_A_lVQAAwvx6_0(.dout(w_dff_A_m6f3wyN56_0),.din(w_dff_A_lVQAAwvx6_0),.clk(gclk));
	jdff dff_A_dYihbfry2_0(.dout(w_dff_A_lVQAAwvx6_0),.din(w_dff_A_dYihbfry2_0),.clk(gclk));
	jdff dff_A_M36QszLj1_0(.dout(w_dff_A_dYihbfry2_0),.din(w_dff_A_M36QszLj1_0),.clk(gclk));
	jdff dff_A_UB4x6zde0_0(.dout(w_dff_A_M36QszLj1_0),.din(w_dff_A_UB4x6zde0_0),.clk(gclk));
	jdff dff_A_Z2Gbt3hQ2_0(.dout(w_Gid20_0[0]),.din(w_dff_A_Z2Gbt3hQ2_0),.clk(gclk));
	jdff dff_A_seRokvUL9_0(.dout(w_dff_A_Z2Gbt3hQ2_0),.din(w_dff_A_seRokvUL9_0),.clk(gclk));
	jdff dff_A_wxPMQh1i0_0(.dout(w_dff_A_seRokvUL9_0),.din(w_dff_A_wxPMQh1i0_0),.clk(gclk));
	jdff dff_A_HadomRkn7_0(.dout(w_dff_A_wxPMQh1i0_0),.din(w_dff_A_HadomRkn7_0),.clk(gclk));
	jdff dff_A_758EfMk28_0(.dout(w_dff_A_HadomRkn7_0),.din(w_dff_A_758EfMk28_0),.clk(gclk));
	jdff dff_A_Ptn8KJ041_0(.dout(w_dff_A_758EfMk28_0),.din(w_dff_A_Ptn8KJ041_0),.clk(gclk));
	jdff dff_A_DUyp6x3e6_0(.dout(w_dff_A_Ptn8KJ041_0),.din(w_dff_A_DUyp6x3e6_0),.clk(gclk));
	jdff dff_A_NyB8ZLBp1_0(.dout(w_dff_A_DUyp6x3e6_0),.din(w_dff_A_NyB8ZLBp1_0),.clk(gclk));
	jdff dff_A_QJ25Jemb0_0(.dout(w_dff_A_NyB8ZLBp1_0),.din(w_dff_A_QJ25Jemb0_0),.clk(gclk));
	jdff dff_A_tTZ8JJQe0_0(.dout(w_dff_A_QJ25Jemb0_0),.din(w_dff_A_tTZ8JJQe0_0),.clk(gclk));
	jdff dff_A_TKmonJqm9_0(.dout(w_dff_A_tTZ8JJQe0_0),.din(w_dff_A_TKmonJqm9_0),.clk(gclk));
	jdff dff_A_FJRfv6Cy4_0(.dout(w_Gid23_0[0]),.din(w_dff_A_FJRfv6Cy4_0),.clk(gclk));
	jdff dff_A_ngjVyaGw8_0(.dout(w_dff_A_FJRfv6Cy4_0),.din(w_dff_A_ngjVyaGw8_0),.clk(gclk));
	jdff dff_A_gWh5xNxq1_0(.dout(w_dff_A_ngjVyaGw8_0),.din(w_dff_A_gWh5xNxq1_0),.clk(gclk));
	jdff dff_A_dlcrq6ji8_0(.dout(w_dff_A_gWh5xNxq1_0),.din(w_dff_A_dlcrq6ji8_0),.clk(gclk));
	jdff dff_A_QoZwEJHg3_0(.dout(w_dff_A_dlcrq6ji8_0),.din(w_dff_A_QoZwEJHg3_0),.clk(gclk));
	jdff dff_A_vjFxjNQc9_0(.dout(w_dff_A_QoZwEJHg3_0),.din(w_dff_A_vjFxjNQc9_0),.clk(gclk));
	jdff dff_A_ZXFIpy399_0(.dout(w_dff_A_vjFxjNQc9_0),.din(w_dff_A_ZXFIpy399_0),.clk(gclk));
	jdff dff_A_QNYVDP5p6_0(.dout(w_dff_A_ZXFIpy399_0),.din(w_dff_A_QNYVDP5p6_0),.clk(gclk));
	jdff dff_A_TGHBsxi64_0(.dout(w_dff_A_QNYVDP5p6_0),.din(w_dff_A_TGHBsxi64_0),.clk(gclk));
	jdff dff_A_D1mDlDEh8_0(.dout(w_dff_A_TGHBsxi64_0),.din(w_dff_A_D1mDlDEh8_0),.clk(gclk));
	jdff dff_A_SKytCwvL1_0(.dout(w_dff_A_D1mDlDEh8_0),.din(w_dff_A_SKytCwvL1_0),.clk(gclk));
	jdff dff_A_BVTWiVJ57_0(.dout(w_Gid22_0[0]),.din(w_dff_A_BVTWiVJ57_0),.clk(gclk));
	jdff dff_A_A7INm0il2_0(.dout(w_dff_A_BVTWiVJ57_0),.din(w_dff_A_A7INm0il2_0),.clk(gclk));
	jdff dff_A_vLmltr8C2_0(.dout(w_dff_A_A7INm0il2_0),.din(w_dff_A_vLmltr8C2_0),.clk(gclk));
	jdff dff_A_nhO2seAI0_0(.dout(w_dff_A_vLmltr8C2_0),.din(w_dff_A_nhO2seAI0_0),.clk(gclk));
	jdff dff_A_NcCUgJXk9_0(.dout(w_dff_A_nhO2seAI0_0),.din(w_dff_A_NcCUgJXk9_0),.clk(gclk));
	jdff dff_A_WVY78wq29_0(.dout(w_dff_A_NcCUgJXk9_0),.din(w_dff_A_WVY78wq29_0),.clk(gclk));
	jdff dff_A_aVpyQfGI2_0(.dout(w_dff_A_WVY78wq29_0),.din(w_dff_A_aVpyQfGI2_0),.clk(gclk));
	jdff dff_A_SOQSC0H94_0(.dout(w_dff_A_aVpyQfGI2_0),.din(w_dff_A_SOQSC0H94_0),.clk(gclk));
	jdff dff_A_1YqQOX3r9_0(.dout(w_dff_A_SOQSC0H94_0),.din(w_dff_A_1YqQOX3r9_0),.clk(gclk));
	jdff dff_A_ji6kDrI13_0(.dout(w_dff_A_1YqQOX3r9_0),.din(w_dff_A_ji6kDrI13_0),.clk(gclk));
	jdff dff_A_I5NWxeFm7_0(.dout(w_dff_A_ji6kDrI13_0),.din(w_dff_A_I5NWxeFm7_0),.clk(gclk));
	jdff dff_A_lUT0JhVq9_0(.dout(w_n128_0[0]),.din(w_dff_A_lUT0JhVq9_0),.clk(gclk));
	jdff dff_A_ulkHrN5l1_0(.dout(w_Gid29_0[0]),.din(w_dff_A_ulkHrN5l1_0),.clk(gclk));
	jdff dff_A_g8ZbEgGx9_0(.dout(w_dff_A_ulkHrN5l1_0),.din(w_dff_A_g8ZbEgGx9_0),.clk(gclk));
	jdff dff_A_xnVp2jXP2_0(.dout(w_dff_A_g8ZbEgGx9_0),.din(w_dff_A_xnVp2jXP2_0),.clk(gclk));
	jdff dff_A_i3LucuSc6_0(.dout(w_dff_A_xnVp2jXP2_0),.din(w_dff_A_i3LucuSc6_0),.clk(gclk));
	jdff dff_A_eweSZZoX1_0(.dout(w_dff_A_i3LucuSc6_0),.din(w_dff_A_eweSZZoX1_0),.clk(gclk));
	jdff dff_A_Q5ReHvpy0_0(.dout(w_dff_A_eweSZZoX1_0),.din(w_dff_A_Q5ReHvpy0_0),.clk(gclk));
	jdff dff_A_7ce1bHCc2_0(.dout(w_dff_A_Q5ReHvpy0_0),.din(w_dff_A_7ce1bHCc2_0),.clk(gclk));
	jdff dff_A_98gQezI82_0(.dout(w_dff_A_7ce1bHCc2_0),.din(w_dff_A_98gQezI82_0),.clk(gclk));
	jdff dff_A_MSB5zrTF4_0(.dout(w_dff_A_98gQezI82_0),.din(w_dff_A_MSB5zrTF4_0),.clk(gclk));
	jdff dff_A_bk9yXZWk1_0(.dout(w_dff_A_MSB5zrTF4_0),.din(w_dff_A_bk9yXZWk1_0),.clk(gclk));
	jdff dff_A_vSOl8sw32_0(.dout(w_dff_A_bk9yXZWk1_0),.din(w_dff_A_vSOl8sw32_0),.clk(gclk));
	jdff dff_A_LAgxRxxT2_0(.dout(w_Gid28_0[0]),.din(w_dff_A_LAgxRxxT2_0),.clk(gclk));
	jdff dff_A_ye7CMO7g0_0(.dout(w_dff_A_LAgxRxxT2_0),.din(w_dff_A_ye7CMO7g0_0),.clk(gclk));
	jdff dff_A_klgElF638_0(.dout(w_dff_A_ye7CMO7g0_0),.din(w_dff_A_klgElF638_0),.clk(gclk));
	jdff dff_A_EZtCkkGH1_0(.dout(w_dff_A_klgElF638_0),.din(w_dff_A_EZtCkkGH1_0),.clk(gclk));
	jdff dff_A_GfpiOfhm2_0(.dout(w_dff_A_EZtCkkGH1_0),.din(w_dff_A_GfpiOfhm2_0),.clk(gclk));
	jdff dff_A_qDVnjXPD7_0(.dout(w_dff_A_GfpiOfhm2_0),.din(w_dff_A_qDVnjXPD7_0),.clk(gclk));
	jdff dff_A_E2ITO4JA5_0(.dout(w_dff_A_qDVnjXPD7_0),.din(w_dff_A_E2ITO4JA5_0),.clk(gclk));
	jdff dff_A_0EfcMfr58_0(.dout(w_dff_A_E2ITO4JA5_0),.din(w_dff_A_0EfcMfr58_0),.clk(gclk));
	jdff dff_A_AhopihAe9_0(.dout(w_dff_A_0EfcMfr58_0),.din(w_dff_A_AhopihAe9_0),.clk(gclk));
	jdff dff_A_DtEhTuRv8_0(.dout(w_dff_A_AhopihAe9_0),.din(w_dff_A_DtEhTuRv8_0),.clk(gclk));
	jdff dff_A_wWcCxshH2_0(.dout(w_dff_A_DtEhTuRv8_0),.din(w_dff_A_wWcCxshH2_0),.clk(gclk));
	jdff dff_A_qPO4PSNX3_0(.dout(w_Gid31_0[0]),.din(w_dff_A_qPO4PSNX3_0),.clk(gclk));
	jdff dff_A_RDLDta620_0(.dout(w_dff_A_qPO4PSNX3_0),.din(w_dff_A_RDLDta620_0),.clk(gclk));
	jdff dff_A_6xjoCarB1_0(.dout(w_dff_A_RDLDta620_0),.din(w_dff_A_6xjoCarB1_0),.clk(gclk));
	jdff dff_A_F9k0fKYS0_0(.dout(w_dff_A_6xjoCarB1_0),.din(w_dff_A_F9k0fKYS0_0),.clk(gclk));
	jdff dff_A_pNrvSiDE7_0(.dout(w_dff_A_F9k0fKYS0_0),.din(w_dff_A_pNrvSiDE7_0),.clk(gclk));
	jdff dff_A_k7AQR2zg6_0(.dout(w_dff_A_pNrvSiDE7_0),.din(w_dff_A_k7AQR2zg6_0),.clk(gclk));
	jdff dff_A_07GujSiq6_0(.dout(w_dff_A_k7AQR2zg6_0),.din(w_dff_A_07GujSiq6_0),.clk(gclk));
	jdff dff_A_d9tJ19oG6_0(.dout(w_dff_A_07GujSiq6_0),.din(w_dff_A_d9tJ19oG6_0),.clk(gclk));
	jdff dff_A_4bZsYWwC2_0(.dout(w_dff_A_d9tJ19oG6_0),.din(w_dff_A_4bZsYWwC2_0),.clk(gclk));
	jdff dff_A_yrXkfJfI7_0(.dout(w_dff_A_4bZsYWwC2_0),.din(w_dff_A_yrXkfJfI7_0),.clk(gclk));
	jdff dff_A_OGfsIYmQ9_0(.dout(w_dff_A_yrXkfJfI7_0),.din(w_dff_A_OGfsIYmQ9_0),.clk(gclk));
	jdff dff_A_UHLZRS6C6_0(.dout(w_Gid30_0[0]),.din(w_dff_A_UHLZRS6C6_0),.clk(gclk));
	jdff dff_A_A7NXdz0I0_0(.dout(w_dff_A_UHLZRS6C6_0),.din(w_dff_A_A7NXdz0I0_0),.clk(gclk));
	jdff dff_A_Vc6VUhUq5_0(.dout(w_dff_A_A7NXdz0I0_0),.din(w_dff_A_Vc6VUhUq5_0),.clk(gclk));
	jdff dff_A_5YsDD7R00_0(.dout(w_dff_A_Vc6VUhUq5_0),.din(w_dff_A_5YsDD7R00_0),.clk(gclk));
	jdff dff_A_zsHJsY5r5_0(.dout(w_dff_A_5YsDD7R00_0),.din(w_dff_A_zsHJsY5r5_0),.clk(gclk));
	jdff dff_A_6axai51y6_0(.dout(w_dff_A_zsHJsY5r5_0),.din(w_dff_A_6axai51y6_0),.clk(gclk));
	jdff dff_A_GYMBMKg37_0(.dout(w_dff_A_6axai51y6_0),.din(w_dff_A_GYMBMKg37_0),.clk(gclk));
	jdff dff_A_C9Qh45ec5_0(.dout(w_dff_A_GYMBMKg37_0),.din(w_dff_A_C9Qh45ec5_0),.clk(gclk));
	jdff dff_A_ezaJ1M593_0(.dout(w_dff_A_C9Qh45ec5_0),.din(w_dff_A_ezaJ1M593_0),.clk(gclk));
	jdff dff_A_Hm4zJxb31_0(.dout(w_dff_A_ezaJ1M593_0),.din(w_dff_A_Hm4zJxb31_0),.clk(gclk));
	jdff dff_A_zjSHKnUH1_0(.dout(w_dff_A_Hm4zJxb31_0),.din(w_dff_A_zjSHKnUH1_0),.clk(gclk));
	jdff dff_A_hRf3olsM3_2(.dout(God0),.din(w_dff_A_hRf3olsM3_2),.clk(gclk));
	jdff dff_A_t7J0DVId7_2(.dout(God1),.din(w_dff_A_t7J0DVId7_2),.clk(gclk));
	jdff dff_A_ploDOSLu9_2(.dout(God2),.din(w_dff_A_ploDOSLu9_2),.clk(gclk));
	jdff dff_A_2pCzVqwn2_2(.dout(God3),.din(w_dff_A_2pCzVqwn2_2),.clk(gclk));
	jdff dff_A_OfomH9JU3_2(.dout(God4),.din(w_dff_A_OfomH9JU3_2),.clk(gclk));
	jdff dff_A_Sijv3I9R3_2(.dout(God5),.din(w_dff_A_Sijv3I9R3_2),.clk(gclk));
	jdff dff_A_Hq6WEn2f5_2(.dout(God6),.din(w_dff_A_Hq6WEn2f5_2),.clk(gclk));
	jdff dff_A_ZlcuYPlk0_2(.dout(God7),.din(w_dff_A_ZlcuYPlk0_2),.clk(gclk));
	jdff dff_A_v119lWYX2_2(.dout(God8),.din(w_dff_A_v119lWYX2_2),.clk(gclk));
	jdff dff_A_2zDjjN1h9_2(.dout(God9),.din(w_dff_A_2zDjjN1h9_2),.clk(gclk));
	jdff dff_A_1PIQUTmW3_2(.dout(God10),.din(w_dff_A_1PIQUTmW3_2),.clk(gclk));
	jdff dff_A_hpEz6GPV6_2(.dout(God11),.din(w_dff_A_hpEz6GPV6_2),.clk(gclk));
	jdff dff_A_dHt9uu4k3_2(.dout(God12),.din(w_dff_A_dHt9uu4k3_2),.clk(gclk));
	jdff dff_A_zjQaDcGc0_2(.dout(God13),.din(w_dff_A_zjQaDcGc0_2),.clk(gclk));
	jdff dff_A_DqBCJwMz4_2(.dout(God14),.din(w_dff_A_DqBCJwMz4_2),.clk(gclk));
	jdff dff_A_8mvuxWeY8_2(.dout(God15),.din(w_dff_A_8mvuxWeY8_2),.clk(gclk));
endmodule

