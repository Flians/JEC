// Benchmark "top" written by ABC on Thu May 28 22:01:08 2020

module gf_sqrt (a, asqrt);
  input [127:0] a;
  output [63:0] asqrt;
  wire n192, n193, n194, n195, n197, n198, n199, n200, n201, n202, n203,
    n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
    n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
    n228, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n259, n260, n261, n262, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
    n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n333, n335, n336, n337, n338, n339, n340,
    n342, n343, n345, n346, n347, n349, n350, n351, n352, n353, n354, n355,
    n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
    n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
    n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
    n393, n394, n395, n396, n397, n399, n400, n401, n402, n403, n404, n405,
    n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
    n430, n431, n432, n433, n434, n435, n436, n437, n438, n440, n441, n442,
    n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
    n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
    n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
    n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
    n503, n504, n505, n506, n507, n508, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
    n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n582, n583, n584, n586, n587, n588,
    n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
    n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
    n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727, n728, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
    n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
    n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
    n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
    n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
    n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
    n806, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
    n819, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
    n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
    n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
    n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
    n869, n870, n871, n872, n873, n874, n875, n876, n878, n879, n880, n881,
    n882, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
    n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
    n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
    n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
    n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
    n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
    n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
    n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
    n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
    n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
    n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
    n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
    n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
    n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
    n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
    n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
    n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
    n1103, n1104, n1105, n1106, n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
    n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
    n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
    n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
    n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
    n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
    n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
    n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
    n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
    n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
    n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
    n1254, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
    n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
    n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
    n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
    n1315, n1316, n1319, n1320, n1321, n1322, n1323, n1325, n1326, n1327,
    n1328, n1329, n1330, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
    n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
    n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
    n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
    n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
    n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
    n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
    n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
    n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
    n1419, n1420, n1421, n1422, n1423, n1424, n1426, n1427, n1428, n1429,
    n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1440, n1441,
    n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
    n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
    n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
    n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
    n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
    n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
    n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
    n1513, n1514, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
    n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
    n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
    n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
    n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
    n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
    n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
    n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
    n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
    n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
    n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
    n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
    n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
    n1674, n1675, n1676, n1677, n1678, n1679, n1681, n1682, n1683, n1684,
    n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
    n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
    n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
    n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
    n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
    n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
    n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
    n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
    n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
    n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
    n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
    n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
    n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
    n1815, n1816, n1817, n1818, n1819, n1821, n1822, n1823, n1824, n1825,
    n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
    n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
    n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
    n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
    n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
    n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
    n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
    n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
    n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
    n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
    n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
    n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
    n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
    n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
    n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
    n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
    n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
    n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
    n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
    n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
    n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
    n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
    n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
    n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
    n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
    n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
    n2096, n2097, n2098, n2099, n2100, n2101, n2103, n2104, n2105, n2106,
    n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
    n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
    n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
    n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
    n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
    n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
    n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
    n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
    n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
    n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
    n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
    n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
    n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
    n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
    n2248, n2249, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
    n2260, n2261, n2262, n2263, n2265, n2266, n2267, n2268, n2269, n2270,
    n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
    n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
    n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
    n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
    n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
    n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
    n2341, n2342, n2343, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
    n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
    n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
    n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
    n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
    n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
    n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
    n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
    n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
    n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
    n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
    n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
    n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
    n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
    n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
    n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
    n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
    n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
    n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
    n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
    n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
    n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
    n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
    n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
    n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
    n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
    n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
    n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
    n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
    n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
    n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
    n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
    n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
    n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
    n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
    n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
    n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
    n2713, n2714, n2715, n2716, n2717, n2719, n2720, n2721, n2722, n2723,
    n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2733, n2734, n2735,
    n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2746,
    n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
    n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
    n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
    n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
    n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
    n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
    n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
    n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
    n2827, n2828, n2829, n2830, n2831, n2833, n2834, n2835, n2836, n2837,
    n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
    n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
    n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
    n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
    n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
    n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
    n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
    n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
    n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
    n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
    n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
    n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
    n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
    n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
    n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
    n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
    n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
    n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
    n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
    n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
    n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
    n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
    n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
    n3068, n3069, n3070, n3071, n3072, n3073, n3075, n3076, n3077, n3078,
    n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
    n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
    n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
    n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
    n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
    n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
    n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
    n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
    n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
    n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
    n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
    n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
    n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
    n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
    n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
    n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
    n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3257, n3258, n3259,
    n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
    n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
    n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
    n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
    n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
    n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
    n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
    n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
    n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
    n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
    n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
    n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
    n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
    n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
    n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
    n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
    n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
    n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
    n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
    n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
    n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
    n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
    n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
    n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
    n3520, n3521, n3522, n3523, n3524, n3526, n3527, n3528, n3529, n3530,
    n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
    n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
    n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
    n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
    n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
    n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
    n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
    n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
    n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
    n3631, n3635, n3636, n3637, n3638, n3639, n3640, n3642, n3643, n3644,
    n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
    n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
    n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
    n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
    n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
    n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
    n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
    n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
    n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
    n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
    n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
    n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
    n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
    n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
    n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
    n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
    n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
    n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
    n3825, n3826, n3827, n3828, n3829, n3830, n3832, n3833, n3834, n3835,
    n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
    n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
    n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
    n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
    n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
    n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
    n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
    n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
    n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
    n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
    n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
    n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
    n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
    n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
    n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
    n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
    n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
    n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
    n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
    n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
    n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
    n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
    n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
    n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
    n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
    n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
    n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
    n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
    n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
    n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
    n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
    n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
    n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
    n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
    n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
    n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
    n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
    n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
    n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
    n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
    n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
    n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
    n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
    n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
    n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
    n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
    n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
    n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
    n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
    n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
    n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
    n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
    n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
    n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
    n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
    n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
    n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
    n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
    n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
    n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
    n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
    n4447, n4448, n4449, n4450, n4452, n4453, n4454, n4455, n4456, n4457,
    n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
    n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
    n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
    n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
    n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
    n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
    n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
    n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
    n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
    n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
    n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
    n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
    n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
    n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
    n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
    n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
    n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
    n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
    n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
    n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
    n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
    n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
    n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
    n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
    n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
    n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
    n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
    n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
    n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
    n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
    n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
    n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
    n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
    n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
    n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
    n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
    n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
    n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
    n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
    n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
    n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
    n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
    n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
    n4888, n4889, n4890, n4891, n4892, n4894, n4895, n4896, n4897, n4898,
    n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
    n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
    n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
    n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
    n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
    n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
    n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
    n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
    n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
    n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
    n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
    n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
    n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
    n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
    n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
    n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
    n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
    n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
    n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
    n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
    n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5107, n5108, n5109,
    n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5121,
    n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
    n5132, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
    n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
    n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
    n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
    n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
    n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
    n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
    n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
    n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
    n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
    n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
    n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
    n5253, n5254, n5255, n5256, n5257, n5259, n5260, n5261, n5262, n5263,
    n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
    n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
    n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
    n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
    n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
    n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
    n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
    n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
    n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
    n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
    n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
    n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
    n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
    n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
    n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
    n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
    n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
    n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
    n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
    n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
    n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
    n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
    n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
    n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
    n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
    n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
    n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
    n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
    n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
    n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
    n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
    n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
    n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
    n5594, n5595, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
    n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
    n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
    n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
    n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
    n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
    n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
    n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
    n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
    n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
    n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
    n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
    n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
    n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
    n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
    n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
    n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
    n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
    n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
    n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
    n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
    n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
    n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
    n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
    n5836, n5837, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
    n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5856, n5857, n5858,
    n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
    n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
    n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
    n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
    n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
    n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
    n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
    n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
    n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
    n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
    n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
    n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
    n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5989,
    n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
    n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
    n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
    n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
    n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
    n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
    n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
    n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
    n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
    n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
    n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
    n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
    n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
    n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
    n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
    n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
    n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
    n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
    n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
    n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
    n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
    n6200, n6201, n6202, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
    n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
    n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
    n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
    n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
    n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
    n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
    n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
    n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
    n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
    n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
    n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
    n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
    n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
    n6341, n6342, n6343, n6344, n6345, n6348, n6349, n6351, n6352, n6353,
    n6354, n6355, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
    n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
    n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
    n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
    n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
    n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
    n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
    n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
    n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
    n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
    n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
    n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
    n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
    n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
    n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
    n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
    n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
    n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
    n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
    n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
    n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
    n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
    n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
    n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
    n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
    n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
    n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
    n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
    n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
    n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
    n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
    n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
    n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
    n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
    n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
    n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
    n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
    n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
    n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
    n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
    n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
    n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
    n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
    n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
    n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
    n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
    n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
    n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
    n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
    n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
    n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
    n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
    n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
    n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
    n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
    n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
    n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
    n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
    n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
    n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
    n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
    n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
    n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
    n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
    n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
    n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
    n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
    n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
    n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
    n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
    n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
    n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
    n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
    n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
    n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
    n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
    n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
    n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
    n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7145, n7146,
    n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
    n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
    n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
    n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
    n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
    n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
    n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
    n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
    n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
    n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
    n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
    n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
    n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
    n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
    n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
    n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
    n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
    n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
    n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
    n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
    n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
    n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
    n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
    n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
    n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
    n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
    n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7417,
    n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
    n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
    n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
    n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
    n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
    n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
    n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
    n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
    n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
    n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
    n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
    n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
    n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
    n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
    n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
    n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
    n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
    n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
    n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
    n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
    n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
    n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
    n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
    n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
    n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
    n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
    n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
    n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
    n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
    n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
    n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
    n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
    n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
    n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
    n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
    n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
    n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
    n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
    n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
    n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
    n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
    n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
    n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
    n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
    n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
    n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
    n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
    n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
    n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
    n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
    n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
    n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
    n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
    n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
    n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
    n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
    n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
    n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
    n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
    n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
    n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
    n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
    n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
    n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
    n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
    n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
    n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
    n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
    n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
    n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
    n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
    n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
    n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
    n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
    n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
    n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
    n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
    n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
    n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
    n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
    n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
    n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
    n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
    n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
    n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
    n8269, n8270, n8271, n8272, n8274, n8275, n8276, n8277, n8278, n8279,
    n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
    n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
    n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
    n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
    n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
    n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
    n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
    n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
    n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
    n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
    n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
    n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
    n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
    n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
    n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
    n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
    n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
    n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
    n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
    n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
    n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
    n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
    n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
    n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
    n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
    n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
    n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
    n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
    n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
    n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
    n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
    n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
    n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
    n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
    n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
    n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
    n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
    n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
    n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
    n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
    n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
    n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
    n8700, n8701, n8702, n8703, n8704, n8705, n8707, n8708, n8709, n8710,
    n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
    n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
    n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
    n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
    n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
    n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
    n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
    n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
    n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
    n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
    n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
    n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
    n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
    n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
    n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
    n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
    n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8882, n8883,
    n8884, n8885, n8886, n8887, n8888, n8890, n8891, n8892, n8893, n8894,
    n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
    n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
    n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
    n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
    n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
    n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
    n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
    n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
    n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
    n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
    n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
    n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
    n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
    n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
    n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
    n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
    n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
    n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
    n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
    n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
    n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
    n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
    n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
    n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
    n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
    n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
    n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
    n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
    n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9184, n9185,
    n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
    n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
    n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
    n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
    n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
    n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
    n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
    n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
    n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
    n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
    n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
    n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
    n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
    n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
    n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
    n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
    n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
    n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
    n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
    n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
    n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
    n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
    n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
    n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
    n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
    n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
    n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
    n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
    n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
    n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
    n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
    n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
    n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
    n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
    n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
    n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
    n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
    n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
    n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
    n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
    n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
    n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
    n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
    n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
    n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
    n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
    n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
    n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
    n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
    n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
    n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
    n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
    n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
    n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
    n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
    n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
    n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
    n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
    n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
    n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
    n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
    n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
    n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
    n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9824, n9825, n9826,
    n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
    n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
    n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
    n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
    n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
    n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
    n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
    n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
    n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
    n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
    n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
    n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
    n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
    n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
    n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
    n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
    n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
    n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
    n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
    n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
    n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
    n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
    n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
    n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
    n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
    n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
    n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
    n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
    n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
    n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
    n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
    n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
    n10132, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
    n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
    n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
    n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
    n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
    n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
    n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
    n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
    n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
    n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
    n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
    n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
    n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
    n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
    n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
    n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
    n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
    n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
    n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
    n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
    n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
    n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
    n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
    n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
    n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
    n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
    n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
    n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
    n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
    n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
    n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
    n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
    n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
    n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
    n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
    n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
    n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
    n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
    n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
    n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
    n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
    n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
    n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
    n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
    n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
    n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
    n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
    n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
    n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
    n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
    n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
    n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
    n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
    n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
    n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
    n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
    n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
    n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
    n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
    n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
    n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
    n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
    n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
    n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
    n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
    n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
    n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
    n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
    n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
    n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
    n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
    n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
    n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
    n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
    n10799, n10800, n10801, n10802, n10803, n10805, n10806, n10807, n10808,
    n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
    n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
    n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
    n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
    n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
    n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
    n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
    n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
    n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
    n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
    n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
    n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
    n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
    n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
    n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
    n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
    n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
    n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
    n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
    n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
    n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
    n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
    n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
    n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
    n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
    n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
    n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
    n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
    n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
    n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
    n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
    n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
    n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
    n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
    n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
    n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
    n11133, n11134, n11135, n11137, n11138, n11139, n11140, n11141, n11142,
    n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
    n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
    n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
    n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
    n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
    n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
    n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
    n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
    n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
    n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
    n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
    n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
    n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
    n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
    n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
    n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
    n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
    n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
    n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
    n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
    n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
    n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
    n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
    n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
    n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
    n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
    n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
    n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
    n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
    n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
    n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
    n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
    n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
    n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
    n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
    n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
    n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
    n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
    n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
    n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
    n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
    n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
    n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
    n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
    n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
    n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
    n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
    n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
    n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
    n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
    n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
    n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
    n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
    n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
    n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
    n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
    n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11656,
    n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
    n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
    n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
    n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
    n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
    n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
    n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
    n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
    n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
    n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
    n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
    n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
    n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
    n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
    n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
    n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
    n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
    n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
    n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
    n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
    n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
    n11846, n11847, n11851, n11852, n11853, n11854, n11855, n11856, n11858,
    n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
    n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
    n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
    n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
    n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
    n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
    n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
    n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
    n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
    n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
    n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
    n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
    n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
    n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
    n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
    n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
    n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
    n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
    n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
    n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
    n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
    n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
    n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
    n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
    n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
    n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
    n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
    n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
    n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
    n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
    n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
    n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
    n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
    n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
    n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
    n12174, n12175, n12176, n12177, n12179, n12180, n12181, n12182, n12183,
    n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12193, n12194,
    n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
    n12204, n12205, n12206, n12207, n12209, n12210, n12211, n12212, n12213,
    n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
    n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
    n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
    n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
    n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
    n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
    n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
    n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
    n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
    n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
    n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
    n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
    n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
    n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
    n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
    n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
    n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
    n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
    n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
    n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
    n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
    n12403, n12404, n12405, n12406, n12407, n12408, n12410, n12411, n12412,
    n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
    n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
    n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
    n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
    n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
    n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
    n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
    n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
    n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
    n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
    n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
    n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
    n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
    n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
    n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
    n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
    n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
    n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
    n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
    n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
    n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
    n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
    n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
    n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
    n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
    n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
    n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
    n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
    n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
    n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
    n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
    n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
    n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
    n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
    n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
    n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
    n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
    n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
    n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
    n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
    n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
    n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
    n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
    n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
    n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
    n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
    n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
    n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
    n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
    n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
    n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
    n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
    n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
    n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
    n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
    n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
    n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
    n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
    n12935, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
    n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
    n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
    n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
    n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
    n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
    n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
    n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
    n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
    n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
    n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
    n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
    n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
    n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
    n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
    n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
    n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
    n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
    n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
    n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
    n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
    n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
    n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
    n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
    n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
    n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
    n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
    n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
    n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
    n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
    n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
    n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
    n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
    n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
    n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
    n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
    n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
    n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
    n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
    n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13296,
    n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
    n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
    n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
    n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
    n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
    n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
    n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
    n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
    n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
    n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
    n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
    n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
    n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
    n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
    n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
    n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
    n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
    n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
    n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
    n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
    n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
    n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
    n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
    n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
    n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
    n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
    n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
    n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
    n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
    n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
    n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
    n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
    n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
    n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
    n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
    n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
    n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
    n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
    n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
    n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
    n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
    n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
    n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
    n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
    n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
    n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
    n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
    n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
    n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
    n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
    n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
    n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
    n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
    n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
    n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
    n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
    n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
    n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
    n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
    n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
    n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
    n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
    n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
    n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
    n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
    n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
    n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
    n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
    n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
    n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
    n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
    n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
    n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
    n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
    n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
    n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
    n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
    n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
    n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
    n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
    n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
    n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
    n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
    n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
    n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
    n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14070, n14071,
    n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
    n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
    n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
    n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
    n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
    n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
    n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
    n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
    n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
    n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
    n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
    n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
    n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
    n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
    n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
    n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
    n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
    n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
    n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
    n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
    n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
    n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
    n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
    n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
    n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
    n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
    n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
    n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
    n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
    n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
    n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
    n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
    n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
    n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
    n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
    n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
    n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
    n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
    n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
    n14423, n14424, n14425, n14426, n14427, n14429, n14430, n14431, n14432,
    n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14443,
    n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
    n14453, n14454, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
    n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
    n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
    n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
    n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
    n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
    n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
    n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
    n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
    n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
    n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
    n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
    n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
    n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
    n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
    n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
    n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
    n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
    n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
    n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
    n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
    n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
    n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
    n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
    n14670, n14671, n14672, n14674, n14675, n14676, n14677, n14678, n14679,
    n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
    n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
    n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
    n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
    n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
    n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
    n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
    n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
    n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
    n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
    n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
    n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
    n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
    n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
    n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
    n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
    n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
    n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
    n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
    n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
    n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
    n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
    n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
    n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
    n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
    n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
    n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
    n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
    n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
    n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
    n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
    n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
    n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
    n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
    n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
    n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
    n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
    n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
    n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
    n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
    n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
    n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
    n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
    n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
    n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
    n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
    n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
    n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
    n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
    n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
    n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
    n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
    n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
    n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
    n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
    n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
    n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
    n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
    n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
    n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
    n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
    n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
    n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15247,
    n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
    n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
    n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
    n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
    n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
    n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
    n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
    n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
    n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
    n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
    n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
    n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
    n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
    n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
    n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
    n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
    n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
    n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
    n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
    n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
    n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
    n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
    n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
    n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
    n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
    n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
    n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
    n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
    n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
    n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
    n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
    n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
    n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
    n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
    n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
    n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
    n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
    n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
    n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
    n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
    n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
    n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
    n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
    n15635, n15636, n15637, n15638, n15639, n15641, n15642, n15643, n15644,
    n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
    n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662,
    n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
    n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
    n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
    n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
    n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
    n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
    n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
    n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734,
    n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
    n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
    n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
    n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
    n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
    n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
    n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
    n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806,
    n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
    n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
    n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
    n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
    n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
    n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
    n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
    n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
    n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
    n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
    n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
    n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
    n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
    n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
    n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
    n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
    n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
    n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
    n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
    n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
    n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
    n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
    n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
    n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
    n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
    n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
    n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
    n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
    n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
    n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
    n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
    n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094,
    n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
    n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
    n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
    n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
    n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
    n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
    n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
    n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
    n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
    n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
    n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
    n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
    n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
    n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
    n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
    n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238,
    n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
    n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
    n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
    n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
    n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
    n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
    n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
    n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
    n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
    n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
    n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
    n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
    n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
    n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
    n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
    n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
    n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
    n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
    n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
    n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
    n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
    n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
    n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
    n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
    n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
    n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
    n16473, n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
    n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
    n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
    n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
    n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518,
    n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
    n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
    n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
    n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
    n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
    n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
    n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581,
    n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
    n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
    n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
    n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
    n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
    n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
    n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
    n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653,
    n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662,
    n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
    n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
    n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
    n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
    n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
    n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
    n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725,
    n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734,
    n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
    n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
    n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
    n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
    n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
    n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
    n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797,
    n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806,
    n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
    n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
    n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
    n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
    n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
    n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
    n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869,
    n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
    n16880, n16881, n16882, n16885, n16886, n16887, n16888, n16889, n16890,
    n16891, n16892, n16893, n16894, n16895, n16896, n16898, n16899, n16900,
    n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909,
    n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918,
    n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
    n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
    n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
    n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
    n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
    n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
    n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
    n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990,
    n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
    n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
    n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
    n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
    n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
    n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
    n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
    n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062,
    n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
    n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
    n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
    n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
    n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
    n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116,
    n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
    n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17134, n17135,
    n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
    n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
    n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
    n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
    n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180,
    n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
    n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198,
    n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
    n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
    n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
    n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
    n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
    n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
    n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
    n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
    n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
    n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
    n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
    n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
    n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
    n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
    n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
    n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
    n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
    n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
    n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
    n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
    n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
    n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
    n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
    n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
    n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
    n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
    n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
    n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
    n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
    n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
    n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
    n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
    n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
    n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
    n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
    n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
    n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
    n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
    n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
    n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
    n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
    n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
    n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
    n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
    n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
    n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612,
    n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
    n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
    n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
    n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
    n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
    n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
    n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
    n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
    n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
    n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
    n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
    n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
    n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
    n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
    n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
    n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756,
    n17757, n17758, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
    n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
    n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
    n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
    n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
    n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
    n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820,
    n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
    n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
    n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
    n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
    n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
    n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
    n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
    n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892,
    n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
    n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
    n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
    n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
    n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
    n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
    n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
    n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964,
    n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
    n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
    n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
    n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
    n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
    n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
    n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
    n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036,
    n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
    n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
    n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063,
    n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
    n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
    n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
    n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
    n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108,
    n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
    n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
    n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
    n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
    n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
    n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
    n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
    n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18180, n18181,
    n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
    n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
    n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
    n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
    n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
    n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
    n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
    n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
    n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
    n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
    n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
    n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
    n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
    n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
    n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
    n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
    n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
    n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
    n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
    n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
    n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
    n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
    n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
    n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
    n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
    n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
    n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
    n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
    n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
    n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
    n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
    n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
    n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
    n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
    n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
    n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
    n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
    n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
    n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
    n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
    n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
    n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
    n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
    n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
    n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
    n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
    n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
    n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
    n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
    n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
    n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
    n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
    n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
    n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
    n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
    n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
    n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694,
    n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
    n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
    n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
    n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
    n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
    n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
    n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
    n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766,
    n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
    n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
    n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
    n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
    n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
    n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
    n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
    n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838,
    n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
    n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
    n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
    n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
    n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
    n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
    n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
    n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
    n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
    n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
    n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
    n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946,
    n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
    n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
    n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
    n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
    n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
    n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
    n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
    n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018,
    n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
    n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
    n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
    n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
    n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
    n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
    n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
    n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
    n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
    n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109,
    n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118,
    n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127,
    n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,
    n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
    n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154,
    n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
    n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
    n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181,
    n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190,
    n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199,
    n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208,
    n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
    n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226,
    n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
    n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
    n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
    n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262,
    n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271,
    n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280,
    n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
    n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298,
    n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
    n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316,
    n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
    n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334,
    n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
    n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352,
    n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
    n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370,
    n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
    n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388,
    n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
    n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406,
    n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
    n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424,
    n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
    n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442,
    n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
    n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
    n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
    n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478,
    n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
    n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
    n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
    n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
    n19515, n19516, n19520, n19521, n19522, n19523, n19524, n19525, n19526,
    n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
    n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
    n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
    n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562,
    n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
    n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580,
    n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
    n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598,
    n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607,
    n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
    n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
    n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
    n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
    n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
    n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
    n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
    n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
    n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
    n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
    n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
    n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
    n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724,
    n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
    n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
    n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
    n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
    n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
    n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
    n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
    n19788, n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
    n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807,
    n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
    n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
    n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834,
    n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
    n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852,
    n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861,
    n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870,
    n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879,
    n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
    n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
    n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906,
    n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
    n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924,
    n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933,
    n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
    n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951,
    n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
    n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
    n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978,
    n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
    n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996,
    n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005,
    n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014,
    n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023,
    n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032,
    n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
    n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
    n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
    n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068,
    n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077,
    n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
    n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095,
    n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104,
    n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
    n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
    n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
    n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140,
    n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149,
    n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158,
    n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167,
    n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176,
    n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
    n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
    n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
    n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212,
    n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221,
    n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
    n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239,
    n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,
    n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
    n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
    n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
    n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
    n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293,
    n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
    n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311,
    n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320,
    n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
    n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338,
    n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
    n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356,
    n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365,
    n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
    n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383,
    n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,
    n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
    n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
    n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
    n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428,
    n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437,
    n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
    n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20455, n20456,
    n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
    n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
    n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
    n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
    n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
    n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
    n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519,
    n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,
    n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
    n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
    n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
    n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
    n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573,
    n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
    n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591,
    n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,
    n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
    n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
    n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
    n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
    n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645,
    n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
    n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663,
    n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672,
    n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
    n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
    n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
    n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
    n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717,
    n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
    n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735,
    n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
    n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
    n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
    n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
    n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
    n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789,
    n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
    n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807,
    n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
    n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
    n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
    n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
    n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
    n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861,
    n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
    n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879,
    n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888,
    n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
    n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20907,
    n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916,
    n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925,
    n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934,
    n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943,
    n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952,
    n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
    n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970,
    n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
    n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988,
    n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997,
    n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006,
    n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015,
    n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024,
    n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
    n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
    n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
    n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060,
    n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069,
    n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078,
    n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087,
    n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096,
    n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
    n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114,
    n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
    n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132,
    n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141,
    n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150,
    n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159,
    n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168,
    n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
    n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186,
    n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195,
    n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204,
    n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213,
    n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222,
    n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231,
    n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240,
    n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
    n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258,
    n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267,
    n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276,
    n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285,
    n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294,
    n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303,
    n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312,
    n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
    n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330,
    n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339,
    n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348,
    n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357,
    n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366,
    n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375,
    n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384,
    n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
    n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402,
    n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411,
    n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420,
    n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429,
    n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438,
    n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447,
    n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456,
    n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
    n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474,
    n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483,
    n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492,
    n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501,
    n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510,
    n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519,
    n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528,
    n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
    n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546,
    n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555,
    n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564,
    n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573,
    n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582,
    n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591,
    n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600,
    n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
    n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618,
    n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627,
    n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636,
    n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645,
    n21646, n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21654,
    n21655, n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663,
    n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672,
    n21673, n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
    n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690,
    n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699,
    n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708,
    n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717,
    n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726,
    n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735,
    n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744,
    n21745, n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
    n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762,
    n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771,
    n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780,
    n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788, n21789,
    n21790, n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21798,
    n21799, n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807,
    n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816,
    n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
    n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834,
    n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843,
    n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852,
    n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860, n21861,
    n21862, n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870,
    n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21880,
    n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
    n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898,
    n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907,
    n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916,
    n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925,
    n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934,
    n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943,
    n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952,
    n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
    n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970,
    n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979,
    n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988,
    n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997,
    n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006,
    n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015,
    n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024,
    n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
    n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042,
    n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051,
    n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060,
    n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069,
    n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078,
    n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087,
    n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096,
    n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
    n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114,
    n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123,
    n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132,
    n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141,
    n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150,
    n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159,
    n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168,
    n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
    n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186,
    n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195,
    n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204,
    n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213,
    n22214, n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222,
    n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231,
    n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240,
    n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
    n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258,
    n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267,
    n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276,
    n22277, n22278, n22279, n22280, n22281, n22282, n22283, n22284, n22285,
    n22286, n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294,
    n22295, n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303,
    n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312,
    n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
    n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330,
    n22331, n22332, n22334, n22335, n22336, n22337, n22338, n22339, n22340,
    n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348, n22349,
    n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357, n22358,
    n22359, n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367,
    n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376,
    n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
    n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394,
    n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403,
    n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411, n22412,
    n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22420, n22421,
    n22422, n22423, n22424, n22425, n22426, n22427, n22428, n22429, n22430,
    n22431, n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439,
    n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448,
    n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
    n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466,
    n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475,
    n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483, n22484,
    n22485, n22486, n22487, n22488, n22489, n22490, n22491, n22492, n22493,
    n22494, n22495, n22496, n22497, n22498, n22499, n22500, n22501, n22502,
    n22503, n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511,
    n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520,
    n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
    n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538,
    n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547,
    n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556,
    n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564, n22565,
    n22566, n22567, n22568, n22569, n22570, n22571, n22572, n22573, n22574,
    n22575, n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583,
    n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592,
    n22593, n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
    n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610,
    n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619,
    n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628,
    n22629, n22630, n22631, n22632, n22633, n22634, n22635, n22636, n22637,
    n22638, n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646,
    n22647, n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655,
    n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664,
    n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
    n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682,
    n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691,
    n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699, n22700,
    n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708, n22709,
    n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717, n22718,
    n22719, n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727,
    n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736,
    n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
    n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754,
    n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763,
    n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771, n22772,
    n22773, n22774, n22775, n22776, n22777, n22778, n22779, n22780, n22781,
    n22782, n22783, n22784, n22785, n22786, n22787, n22788, n22789, n22790,
    n22791, n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799,
    n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808,
    n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
    n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825, n22826,
    n22827, n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835,
    n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843, n22844,
    n22845, n22846, n22847, n22848, n22849, n22850, n22851, n22852, n22853,
    n22854, n22855, n22856, n22857, n22858, n22859, n22860, n22861, n22862,
    n22863, n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871,
    n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22879, n22880,
    n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
    n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898,
    n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907,
    n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915, n22916,
    n22917, n22918, n22919, n22920, n22921, n22922, n22923, n22924, n22925,
    n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933, n22934,
    n22935, n22936, n22937, n22938, n22939, n22940, n22941, n22942, n22943,
    n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952,
    n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
    n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970,
    n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979,
    n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987, n22988,
    n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997,
    n22998, n22999, n23000, n23001, n23002, n23003, n23004, n23005, n23006,
    n23007, n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015,
    n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023, n23024,
    n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
    n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041, n23042,
    n23043, n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051,
    n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059, n23060,
    n23061, n23062, n23063, n23064, n23065, n23066, n23067, n23068, n23069,
    n23070, n23071, n23072, n23073, n23074, n23075, n23076, n23077, n23078,
    n23079, n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087,
    n23088, n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096,
    n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
    n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114,
    n23115, n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123,
    n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131, n23132,
    n23133, n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141,
    n23142, n23143, n23144, n23145, n23146, n23147, n23148, n23149, n23150,
    n23151, n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159,
    n23160, n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168,
    n23169, n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
    n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185, n23186,
    n23187, n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195,
    n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203, n23204,
    n23205, n23206, n23207, n23208, n23209, n23210, n23211, n23212, n23213,
    n23214, n23215, n23216, n23217, n23218, n23219, n23220, n23221, n23222,
    n23223, n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231,
    n23232, n23233, n23234, n23235, n23236, n23237, n23238, n23239, n23240,
    n23241, n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
    n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257, n23258,
    n23259, n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267,
    n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275, n23276,
    n23277, n23278, n23279, n23280, n23281, n23282, n23283, n23284, n23285,
    n23286, n23287, n23288, n23289, n23290, n23291, n23292, n23293, n23294,
    n23295, n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303,
    n23304, n23305, n23306, n23307, n23308, n23309, n23310, n23311, n23312,
    n23313, n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
    n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329, n23330,
    n23331, n23332, n23333, n23334, n23335, n23336, n23338, n23339, n23340,
    n23341, n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349,
    n23350, n23351, n23352, n23353, n23354, n23355, n23356, n23357, n23358,
    n23359, n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367,
    n23368, n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376,
    n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
    n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394,
    n23395, n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403,
    n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411, n23412,
    n23413, n23414, n23415, n23416, n23417, n23418, n23419, n23420, n23421,
    n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23429, n23430,
    n23431, n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439,
    n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448,
    n23449, n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
    n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465, n23466,
    n23467, n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475,
    n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483, n23484,
    n23485, n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23493,
    n23494, n23495, n23496, n23497, n23498, n23499, n23500, n23501, n23502,
    n23503, n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511,
    n23512, n23513, n23514, n23515, n23516, n23517, n23518, n23519, n23520,
    n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
    n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538,
    n23539, n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547,
    n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555, n23556,
    n23557, n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565,
    n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573, n23574,
    n23575, n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583,
    n23584, n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23592,
    n23593, n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
    n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609, n23610,
    n23611, n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619,
    n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627, n23628,
    n23629, n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637,
    n23638, n23639, n23640, n23641, n23642, n23643, n23644, n23645, n23646,
    n23647, n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655,
    n23656, n23657, n23658, n23659, n23660, n23661, n23662, n23663, n23664,
    n23665, n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
    n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681, n23682,
    n23683, n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691,
    n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699, n23700,
    n23701, n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709,
    n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717, n23718,
    n23719, n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727,
    n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735, n23736,
    n23737, n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
    n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753, n23754,
    n23755, n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763,
    n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771, n23772,
    n23773, n23774, n23775, n23776, n23777, n23778, n23779, n23780, n23781,
    n23782, n23783, n23784, n23785, n23786, n23787, n23788, n23789, n23790,
    n23791, n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799,
    n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23808, n23809,
    n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817, n23818,
    n23819, n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827,
    n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835, n23836,
    n23837, n23838, n23839, n23840, n23841, n23842, n23843, n23844, n23845,
    n23846, n23847, n23848, n23849, n23850, n23851, n23852, n23853, n23854,
    n23855, n23856, n23857, n23858, n23859, n23860, n23861, n23862, n23863,
    n23864, n23865, n23866, n23867, n23868, n23869, n23870, n23871, n23872,
    n23873, n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
    n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889, n23890,
    n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899,
    n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907, n23908,
    n23909, n23910, n23911, n23912, n23913, n23914, n23915, n23916, n23917,
    n23918, n23919, n23920, n23921, n23922, n23923, n23924, n23925, n23926,
    n23927, n23928, n23929, n23930, n23931, n23932, n23933, n23934, n23935,
    n23936, n23937, n23938, n23939, n23940, n23941, n23942, n23943, n23944,
    n23945, n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
    n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961, n23962,
    n23963, n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971,
    n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979, n23980,
    n23981, n23982, n23983, n23984, n23985, n23986, n23987, n23988, n23989,
    n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997, n23998,
    n23999, n24000, n24001, n24002, n24003, n24004, n24005, n24006, n24007,
    n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015, n24016,
    n24017, n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
    n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033, n24034,
    n24035, n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043,
    n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051, n24052,
    n24053, n24054, n24055, n24056, n24057, n24058, n24059, n24060, n24061,
    n24062, n24063, n24064, n24065, n24066, n24067, n24068, n24069, n24070,
    n24071, n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079,
    n24080, n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088,
    n24089, n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
    n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105, n24106,
    n24107, n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115,
    n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123, n24124,
    n24125, n24126, n24127, n24128, n24129, n24130, n24131, n24132, n24133,
    n24134, n24135, n24136, n24137, n24138, n24139, n24140, n24141, n24142,
    n24143, n24144, n24145, n24146, n24147, n24148, n24149, n24150, n24151,
    n24152, n24153, n24154, n24155, n24156, n24157, n24158, n24159, n24160,
    n24161, n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
    n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177, n24178,
    n24179, n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187,
    n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195, n24196,
    n24197, n24198, n24199, n24200, n24201, n24202, n24203, n24204, n24205,
    n24206, n24207, n24208, n24209, n24210, n24211, n24212, n24213, n24214,
    n24215, n24216, n24217, n24218, n24219, n24220, n24221, n24222, n24223,
    n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231, n24232,
    n24233, n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
    n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249, n24250,
    n24251, n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259,
    n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267, n24268,
    n24269, n24270, n24271, n24272, n24273, n24274, n24275, n24276, n24277,
    n24278, n24279, n24280, n24281, n24282, n24283, n24284, n24285, n24286,
    n24287, n24288, n24289, n24290, n24291, n24292, n24293, n24294, n24295,
    n24296, n24297, n24298, n24299, n24300, n24301, n24302, n24303, n24304,
    n24305, n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
    n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322,
    n24323, n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331,
    n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339, n24340,
    n24341, n24342, n24343, n24344, n24345, n24346, n24347, n24348, n24349,
    n24350, n24351, n24352, n24353, n24354, n24355, n24356, n24357, n24358,
    n24359, n24360, n24361, n24362, n24363, n24364, n24365, n24366, n24367,
    n24368, n24369, n24370, n24371, n24372, n24373, n24374, n24375, n24376,
    n24377, n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
    n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393, n24394,
    n24395, n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403,
    n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411, n24412,
    n24413, n24414, n24415, n24416, n24417, n24418, n24419, n24420, n24421,
    n24422, n24423, n24424, n24425, n24426, n24427, n24428, n24429, n24430,
    n24431, n24432, n24433, n24434, n24435, n24436, n24437, n24438, n24439,
    n24440, n24441, n24442, n24443, n24444, n24445, n24446, n24447, n24448,
    n24449, n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
    n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24466,
    n24467, n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475,
    n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483, n24484,
    n24485, n24486, n24487, n24488, n24489, n24490, n24491, n24492, n24493,
    n24494, n24495, n24496, n24497, n24498, n24499, n24500, n24501, n24502,
    n24503, n24504, n24505, n24506, n24507, n24508, n24509, n24510, n24511,
    n24512, n24513, n24514, n24515, n24516, n24517, n24518, n24519, n24520,
    n24521, n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
    n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537, n24538,
    n24539, n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547,
    n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555, n24556,
    n24557, n24558, n24559, n24560, n24561, n24562, n24563, n24564, n24565,
    n24566, n24567, n24568, n24569, n24570, n24571, n24572, n24573, n24574,
    n24575, n24576, n24577, n24578, n24579, n24580, n24581, n24582, n24583,
    n24584, n24585, n24586, n24587, n24588, n24589, n24590, n24591, n24592,
    n24593, n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
    n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609, n24610,
    n24611, n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619,
    n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627, n24628,
    n24629, n24630, n24631, n24632, n24633, n24634, n24635, n24636, n24637,
    n24638, n24639, n24640, n24641, n24642, n24643, n24644, n24645, n24646,
    n24647, n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655,
    n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24663, n24664,
    n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
    n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682,
    n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691,
    n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699, n24700,
    n24701, n24702, n24703, n24704, n24705, n24706, n24707, n24708, n24709,
    n24710, n24711, n24712, n24713, n24714, n24715, n24716, n24717, n24718,
    n24719, n24720, n24721, n24722, n24723, n24724, n24725, n24726, n24727,
    n24728, n24729, n24730, n24731, n24732, n24733, n24734, n24735, n24736,
    n24737, n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
    n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753, n24754,
    n24755, n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763,
    n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771, n24772,
    n24773, n24774, n24775, n24776, n24777, n24778, n24779, n24780, n24781,
    n24782, n24783, n24784, n24785, n24786, n24787, n24788, n24789, n24790,
    n24791, n24792, n24793, n24794, n24795, n24796, n24797, n24798, n24799,
    n24800, n24801, n24802, n24803, n24804, n24805, n24806, n24807, n24808,
    n24809, n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
    n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24826,
    n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835,
    n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843, n24844,
    n24845, n24846, n24848, n24849, n24850, n24851, n24852, n24853, n24854,
    n24855, n24856, n24857, n24858, n24859, n24860, n24861, n24862, n24863,
    n24864, n24865, n24866, n24867, n24868, n24869, n24870, n24871, n24872,
    n24873, n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
    n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889, n24890,
    n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899,
    n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907, n24908,
    n24909, n24910, n24911, n24912, n24913, n24914, n24915, n24916, n24917,
    n24918, n24919, n24920, n24921, n24922, n24923, n24924, n24925, n24926,
    n24927, n24928, n24929, n24930, n24931, n24932, n24933, n24934, n24935,
    n24936, n24937, n24938, n24939, n24940, n24941, n24942, n24943, n24944,
    n24945, n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
    n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962,
    n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971,
    n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979, n24980,
    n24981, n24982, n24983, n24984, n24985, n24986, n24987, n24988, n24989,
    n24990, n24991, n24992, n24993, n24994, n24995, n24996, n24997, n24998,
    n24999, n25000, n25001, n25002, n25003, n25004, n25005, n25006, n25007,
    n25008, n25009, n25010, n25011, n25012, n25013, n25014, n25015, n25016,
    n25017, n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
    n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033, n25034,
    n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042, n25043,
    n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051, n25052,
    n25053, n25054, n25055, n25056, n25057, n25058, n25059, n25060, n25061,
    n25062, n25063, n25064, n25065, n25066, n25067, n25068, n25069, n25070,
    n25071, n25072, n25073, n25074, n25075, n25076, n25077, n25078, n25079,
    n25080, n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25088,
    n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
    n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106,
    n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115,
    n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123, n25124,
    n25125, n25126, n25127, n25128, n25129, n25130, n25131, n25132, n25133,
    n25134, n25135, n25136, n25137, n25138, n25139, n25140, n25141, n25142,
    n25143, n25144, n25145, n25146, n25147, n25148, n25149, n25150, n25151,
    n25152, n25153, n25154, n25155, n25156, n25157, n25158, n25159, n25160,
    n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
    n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178,
    n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187,
    n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195, n25196,
    n25197, n25198, n25199, n25200, n25201, n25202, n25203, n25204, n25205,
    n25206, n25207, n25208, n25209, n25210, n25211, n25212, n25213, n25214,
    n25215, n25216, n25217, n25218, n25219, n25220, n25221, n25222, n25223,
    n25224, n25225, n25226, n25227, n25228, n25229, n25230, n25231, n25232,
    n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
    n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250,
    n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259,
    n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267, n25268,
    n25269, n25270, n25271, n25272, n25273, n25274, n25275, n25276, n25277,
    n25278, n25279, n25280, n25281, n25282, n25283, n25284, n25285, n25286,
    n25287, n25288, n25289, n25290, n25291, n25292, n25293, n25294, n25295,
    n25296, n25297, n25298, n25299, n25300;
  jand g00000(.dina(a[127] ), .dinb(a[126] ), .dout(n192));
  jnot g00001(.din(a[126] ), .dout(n193));
  jor  g00002(.dina(a[125] ), .dinb(a[124] ), .dout(n194));
  jand g00003(.dina(n194), .dinb(n193), .dout(n195));
  jor  g00004(.dina(n195), .dinb(n192), .dout(asqrt[62] ));
  jnot g00005(.din(a[127] ), .dout(n197));
  jnot g00006(.din(a[124] ), .dout(n198));
  jnot g00007(.din(a[125] ), .dout(n199));
  jand g00008(.dina(n199), .dinb(n198), .dout(n200));
  jand g00009(.dina(n200), .dinb(a[126] ), .dout(n201));
  jor  g00010(.dina(n201), .dinb(n197), .dout(n202));
  jor  g00011(.dina(n202), .dinb(n195), .dout(n203));
  jnot g00012(.din(n203), .dout(n204));
  jand g00013(.dina(asqrt[62] ), .dinb(n198), .dout(n205));
  jor  g00014(.dina(n205), .dinb(n199), .dout(n206));
  jand g00015(.dina(n200), .dinb(n192), .dout(n207));
  jnot g00016(.din(n207), .dout(n208));
  jand g00017(.dina(n208), .dinb(n206), .dout(n209));
  jand g00018(.dina(asqrt[62] ), .dinb(a[124] ), .dout(n210));
  jnot g00019(.din(a[122] ), .dout(n211));
  jnot g00020(.din(a[123] ), .dout(n212));
  jand g00021(.dina(n198), .dinb(n212), .dout(n213));
  jand g00022(.dina(n213), .dinb(n211), .dout(n214));
  jor  g00023(.dina(n214), .dinb(n210), .dout(n215));
  jor  g00024(.dina(n215), .dinb(n209), .dout(n216));
  jnot g00025(.din(n216), .dout(n217));
  jand g00026(.dina(n197), .dinb(n193), .dout(n218));
  jnot g00027(.din(n192), .dout(n219));
  jor  g00028(.dina(n200), .dinb(a[126] ), .dout(n220));
  jand g00029(.dina(n220), .dinb(n219), .dout(n221));
  jor  g00030(.dina(n221), .dinb(a[124] ), .dout(n222));
  jand g00031(.dina(n222), .dinb(a[125] ), .dout(n223));
  jor  g00032(.dina(n207), .dinb(n223), .dout(n224));
  jnot g00033(.din(n215), .dout(n225));
  jor  g00034(.dina(n225), .dinb(n224), .dout(n226));
  jand g00035(.dina(n226), .dinb(n218), .dout(n227));
  jor  g00036(.dina(n227), .dinb(n217), .dout(n228));
  jor  g00037(.dina(n228), .dinb(n204), .dout(asqrt[61] ));
  jnot g00038(.din(n218), .dout(asqrt[63] ));
  jand g00039(.dina(n225), .dinb(n204), .dout(n231));
  jor  g00040(.dina(n231), .dinb(n224), .dout(n232));
  jand g00041(.dina(n232), .dinb(asqrt[63] ), .dout(n233));
  jand g00042(.dina(n233), .dinb(n216), .dout(n234));
  jand g00043(.dina(n215), .dinb(n209), .dout(n235));
  jand g00044(.dina(n235), .dinb(n204), .dout(n236));
  jor  g00045(.dina(n235), .dinb(asqrt[63] ), .dout(n237));
  jand g00046(.dina(n237), .dinb(n216), .dout(n238));
  jand g00047(.dina(n238), .dinb(n203), .dout(n239));
  jor  g00048(.dina(n239), .dinb(n211), .dout(n240));
  jnot g00049(.din(a[120] ), .dout(n241));
  jnot g00050(.din(a[121] ), .dout(n242));
  jand g00051(.dina(n242), .dinb(n241), .dout(n243));
  jand g00052(.dina(n243), .dinb(n211), .dout(n244));
  jnot g00053(.din(n244), .dout(n245));
  jand g00054(.dina(n245), .dinb(n240), .dout(n246));
  jor  g00055(.dina(n246), .dinb(n221), .dout(n247));
  jand g00056(.dina(n246), .dinb(n221), .dout(n248));
  jor  g00057(.dina(n239), .dinb(a[122] ), .dout(n249));
  jxor g00058(.dina(n249), .dinb(n212), .dout(n250));
  jor  g00059(.dina(n250), .dinb(n248), .dout(n251));
  jand g00060(.dina(n251), .dinb(n247), .dout(n252));
  jor  g00061(.dina(n249), .dinb(a[123] ), .dout(n253));
  jor  g00062(.dina(asqrt[61] ), .dinb(n221), .dout(n254));
  jand g00063(.dina(n254), .dinb(n253), .dout(n255));
  jxor g00064(.dina(n255), .dinb(n198), .dout(n256));
  jor  g00065(.dina(n256), .dinb(n252), .dout(n257));
  jor  g00066(.dina(n257), .dinb(n217), .dout(n258));
  jor  g00067(.dina(n258), .dinb(n236), .dout(n259));
  jand g00068(.dina(n259), .dinb(n218), .dout(n260));
  jand g00069(.dina(n256), .dinb(n252), .dout(n261));
  jor  g00070(.dina(n261), .dinb(n260), .dout(n262));
  jor  g00071(.dina(n262), .dinb(n234), .dout(asqrt[60] ));
  jnot g00072(.din(n250), .dout(n264));
  jxor g00073(.dina(n246), .dinb(n221), .dout(n265));
  jand g00074(.dina(n265), .dinb(asqrt[60] ), .dout(n266));
  jxor g00075(.dina(n266), .dinb(n264), .dout(n267));
  jnot g00076(.din(a[118] ), .dout(n268));
  jnot g00077(.din(a[119] ), .dout(n269));
  jand g00078(.dina(n269), .dinb(n268), .dout(n270));
  jand g00079(.dina(n270), .dinb(n241), .dout(n271));
  jand g00080(.dina(asqrt[60] ), .dinb(a[120] ), .dout(n272));
  jor  g00081(.dina(n272), .dinb(n271), .dout(n273));
  jand g00082(.dina(n273), .dinb(asqrt[61] ), .dout(n274));
  jor  g00083(.dina(n273), .dinb(asqrt[61] ), .dout(n275));
  jand g00084(.dina(asqrt[60] ), .dinb(n241), .dout(n276));
  jor  g00085(.dina(n276), .dinb(n242), .dout(n277));
  jnot g00086(.din(n243), .dout(n278));
  jnot g00087(.din(n234), .dout(n279));
  jnot g00088(.din(n236), .dout(n280));
  jnot g00089(.din(n247), .dout(n281));
  jand g00090(.dina(asqrt[61] ), .dinb(a[122] ), .dout(n282));
  jor  g00091(.dina(n244), .dinb(n282), .dout(n283));
  jor  g00092(.dina(n283), .dinb(asqrt[62] ), .dout(n284));
  jand g00093(.dina(n264), .dinb(n284), .dout(n285));
  jor  g00094(.dina(n285), .dinb(n281), .dout(n286));
  jnot g00095(.din(n256), .dout(n287));
  jand g00096(.dina(n287), .dinb(n286), .dout(n288));
  jand g00097(.dina(n288), .dinb(n216), .dout(n289));
  jand g00098(.dina(n289), .dinb(n280), .dout(n290));
  jor  g00099(.dina(n290), .dinb(asqrt[63] ), .dout(n291));
  jnot g00100(.din(n261), .dout(n292));
  jand g00101(.dina(n292), .dinb(n291), .dout(n293));
  jand g00102(.dina(n293), .dinb(n279), .dout(n294));
  jor  g00103(.dina(n294), .dinb(n278), .dout(n295));
  jand g00104(.dina(n295), .dinb(n277), .dout(n296));
  jand g00105(.dina(n296), .dinb(n275), .dout(n297));
  jor  g00106(.dina(n297), .dinb(n274), .dout(n298));
  jand g00107(.dina(n298), .dinb(asqrt[62] ), .dout(n299));
  jor  g00108(.dina(n298), .dinb(asqrt[62] ), .dout(n300));
  jor  g00109(.dina(asqrt[60] ), .dinb(n239), .dout(n301));
  jand g00110(.dina(n301), .dinb(n295), .dout(n302));
  jxor g00111(.dina(n302), .dinb(n211), .dout(n303));
  jnot g00112(.din(n303), .dout(n304));
  jand g00113(.dina(n304), .dinb(n300), .dout(n305));
  jor  g00114(.dina(n305), .dinb(n299), .dout(n306));
  jor  g00115(.dina(n306), .dinb(n267), .dout(n307));
  jand g00116(.dina(n307), .dinb(asqrt[63] ), .dout(n308));
  jnot g00117(.din(n308), .dout(n309));
  jnot g00118(.din(n307), .dout(n310));
  jnot g00119(.din(n267), .dout(n311));
  jnot g00120(.din(n299), .dout(n312));
  jnot g00121(.din(n274), .dout(n313));
  jnot g00122(.din(n271), .dout(n314));
  jor  g00123(.dina(n294), .dinb(n241), .dout(n315));
  jand g00124(.dina(n315), .dinb(n314), .dout(n316));
  jand g00125(.dina(n316), .dinb(n239), .dout(n317));
  jor  g00126(.dina(n294), .dinb(a[120] ), .dout(n318));
  jand g00127(.dina(n318), .dinb(a[121] ), .dout(n319));
  jand g00128(.dina(asqrt[60] ), .dinb(n243), .dout(n320));
  jor  g00129(.dina(n320), .dinb(n319), .dout(n321));
  jor  g00130(.dina(n321), .dinb(n317), .dout(n322));
  jand g00131(.dina(n322), .dinb(n313), .dout(n323));
  jand g00132(.dina(n323), .dinb(n221), .dout(n324));
  jor  g00133(.dina(n303), .dinb(n324), .dout(n325));
  jand g00134(.dina(n325), .dinb(n312), .dout(n326));
  jor  g00135(.dina(n326), .dinb(n311), .dout(n327));
  jxor g00136(.dina(n256), .dinb(n252), .dout(n328));
  jor  g00137(.dina(n328), .dinb(n294), .dout(n329));
  jnot g00138(.din(n329), .dout(n330));
  jor  g00139(.dina(n330), .dinb(n327), .dout(n331));
  jand g00140(.dina(n331), .dinb(n309), .dout(n333));
  jor  g00141(.dina(n260), .dinb(n330), .dout(n335));
  jnot g00142(.din(n335), .dout(n336));
  jor  g00143(.dina(n336), .dinb(n333), .dout(n337));
  jand g00144(.dina(n294), .dinb(n287), .dout(n338));
  jnot g00145(.din(n338), .dout(n339));
  jor  g00146(.dina(n339), .dinb(n333), .dout(n340));
  jand g00147(.dina(n340), .dinb(n337), .dout(asqrt[59] ));
  jand g00148(.dina(n306), .dinb(n267), .dout(n342));
  jand g00149(.dina(asqrt[59] ), .dinb(n342), .dout(n343));
  jor  g00150(.dina(n333), .dinb(n343), .dout(n345));
  jnot g00151(.din(n345), .dout(n346));
  jand g00152(.dina(n329), .dinb(n342), .dout(n347));
  jor  g00153(.dina(n347), .dinb(n308), .dout(n349));
  jand g00154(.dina(n335), .dinb(n349), .dout(n350));
  jand g00155(.dina(n338), .dinb(n349), .dout(n351));
  jor  g00156(.dina(n351), .dinb(n350), .dout(n352));
  jor  g00157(.dina(n352), .dinb(n268), .dout(n353));
  jnot g00158(.din(a[116] ), .dout(n354));
  jnot g00159(.din(a[117] ), .dout(n355));
  jand g00160(.dina(n355), .dinb(n354), .dout(n356));
  jand g00161(.dina(n356), .dinb(n268), .dout(n357));
  jnot g00162(.din(n357), .dout(n358));
  jand g00163(.dina(n358), .dinb(n353), .dout(n359));
  jor  g00164(.dina(n359), .dinb(n294), .dout(n360));
  jand g00165(.dina(n359), .dinb(n294), .dout(n361));
  jor  g00166(.dina(n352), .dinb(a[118] ), .dout(n362));
  jand g00167(.dina(n362), .dinb(a[119] ), .dout(n363));
  jand g00168(.dina(asqrt[59] ), .dinb(n270), .dout(n364));
  jor  g00169(.dina(n364), .dinb(n363), .dout(n365));
  jor  g00170(.dina(n365), .dinb(n361), .dout(n366));
  jand g00171(.dina(n366), .dinb(n360), .dout(n367));
  jor  g00172(.dina(n367), .dinb(n239), .dout(n368));
  jand g00173(.dina(n367), .dinb(n239), .dout(n369));
  jnot g00174(.din(n270), .dout(n370));
  jor  g00175(.dina(n352), .dinb(n370), .dout(n371));
  jand g00176(.dina(n371), .dinb(n337), .dout(n372));
  jxor g00177(.dina(n372), .dinb(n241), .dout(n373));
  jor  g00178(.dina(n373), .dinb(n369), .dout(n374));
  jand g00179(.dina(n374), .dinb(n368), .dout(n375));
  jor  g00180(.dina(n375), .dinb(n221), .dout(n376));
  jand g00181(.dina(n375), .dinb(n221), .dout(n377));
  jxor g00182(.dina(n273), .dinb(n239), .dout(n378));
  jor  g00183(.dina(n378), .dinb(n352), .dout(n379));
  jxor g00184(.dina(n379), .dinb(n321), .dout(n380));
  jnot g00185(.din(n380), .dout(n381));
  jor  g00186(.dina(n381), .dinb(n377), .dout(n382));
  jand g00187(.dina(n382), .dinb(n376), .dout(n383));
  jxor g00188(.dina(n298), .dinb(n221), .dout(n384));
  jor  g00189(.dina(n384), .dinb(n352), .dout(n385));
  jxor g00190(.dina(n385), .dinb(n304), .dout(n386));
  jand g00191(.dina(n386), .dinb(n383), .dout(n387));
  jor  g00192(.dina(n387), .dinb(n218), .dout(n388));
  jor  g00193(.dina(n386), .dinb(n383), .dout(n389));
  jor  g00194(.dina(n343), .dinb(n310), .dout(n390));
  jor  g00195(.dina(n390), .dinb(n389), .dout(n391));
  jand g00196(.dina(n391), .dinb(n388), .dout(n393));
  jor  g00197(.dina(n393), .dinb(n346), .dout(n394));
  jand g00198(.dina(n352), .dinb(n267), .dout(n395));
  jnot g00199(.din(n395), .dout(n396));
  jor  g00200(.dina(n396), .dinb(n393), .dout(n397));
  jand g00201(.dina(n397), .dinb(n394), .dout(asqrt[58] ));
  jnot g00202(.din(n376), .dout(n399));
  jnot g00203(.din(n368), .dout(n400));
  jnot g00204(.din(n360), .dout(n401));
  jand g00205(.dina(asqrt[59] ), .dinb(a[118] ), .dout(n402));
  jor  g00206(.dina(n357), .dinb(n402), .dout(n403));
  jor  g00207(.dina(n403), .dinb(asqrt[60] ), .dout(n404));
  jand g00208(.dina(asqrt[59] ), .dinb(n268), .dout(n405));
  jor  g00209(.dina(n405), .dinb(n269), .dout(n406));
  jand g00210(.dina(n371), .dinb(n406), .dout(n407));
  jand g00211(.dina(n407), .dinb(n404), .dout(n408));
  jor  g00212(.dina(n408), .dinb(n401), .dout(n409));
  jor  g00213(.dina(n409), .dinb(asqrt[61] ), .dout(n410));
  jnot g00214(.din(n373), .dout(n411));
  jand g00215(.dina(n411), .dinb(n410), .dout(n412));
  jor  g00216(.dina(n412), .dinb(n400), .dout(n413));
  jor  g00217(.dina(n413), .dinb(asqrt[62] ), .dout(n414));
  jand g00218(.dina(n380), .dinb(n414), .dout(n415));
  jor  g00219(.dina(n415), .dinb(n399), .dout(n416));
  jnot g00220(.din(n386), .dout(n417));
  jand g00221(.dina(n417), .dinb(n416), .dout(n418));
  jand g00222(.dina(asqrt[58] ), .dinb(n418), .dout(n419));
  jxor g00223(.dina(n375), .dinb(n221), .dout(n420));
  jand g00224(.dina(n420), .dinb(asqrt[58] ), .dout(n421));
  jxor g00225(.dina(n421), .dinb(n380), .dout(n422));
  jnot g00226(.din(n422), .dout(n423));
  jand g00227(.dina(asqrt[58] ), .dinb(a[116] ), .dout(n424));
  jnot g00228(.din(a[114] ), .dout(n425));
  jnot g00229(.din(a[115] ), .dout(n426));
  jand g00230(.dina(n426), .dinb(n425), .dout(n427));
  jand g00231(.dina(n427), .dinb(n354), .dout(n428));
  jor  g00232(.dina(n428), .dinb(n424), .dout(n429));
  jand g00233(.dina(n429), .dinb(asqrt[59] ), .dout(n430));
  jor  g00234(.dina(n429), .dinb(asqrt[59] ), .dout(n431));
  jand g00235(.dina(asqrt[58] ), .dinb(n354), .dout(n432));
  jor  g00236(.dina(n432), .dinb(n355), .dout(n433));
  jnot g00237(.din(n356), .dout(n434));
  jnot g00238(.din(n388), .dout(n435));
  jnot g00239(.din(n387), .dout(n436));
  jnot g00240(.din(n390), .dout(n437));
  jand g00241(.dina(n437), .dinb(n418), .dout(n438));
  jor  g00242(.dina(n438), .dinb(n435), .dout(n440));
  jand g00243(.dina(n440), .dinb(n345), .dout(n441));
  jand g00244(.dina(n395), .dinb(n440), .dout(n442));
  jor  g00245(.dina(n442), .dinb(n441), .dout(n443));
  jor  g00246(.dina(n443), .dinb(n434), .dout(n444));
  jand g00247(.dina(n444), .dinb(n433), .dout(n445));
  jand g00248(.dina(n445), .dinb(n431), .dout(n446));
  jor  g00249(.dina(n446), .dinb(n430), .dout(n447));
  jand g00250(.dina(n447), .dinb(asqrt[60] ), .dout(n448));
  jor  g00251(.dina(n447), .dinb(asqrt[60] ), .dout(n449));
  jand g00252(.dina(asqrt[58] ), .dinb(n356), .dout(n450));
  jor  g00253(.dina(n450), .dinb(n441), .dout(n451));
  jxor g00254(.dina(n451), .dinb(a[118] ), .dout(n452));
  jnot g00255(.din(n452), .dout(n453));
  jand g00256(.dina(n453), .dinb(n449), .dout(n454));
  jor  g00257(.dina(n454), .dinb(n448), .dout(n455));
  jand g00258(.dina(n455), .dinb(asqrt[61] ), .dout(n456));
  jor  g00259(.dina(n455), .dinb(asqrt[61] ), .dout(n457));
  jxor g00260(.dina(n359), .dinb(n294), .dout(n458));
  jand g00261(.dina(n458), .dinb(asqrt[58] ), .dout(n459));
  jxor g00262(.dina(n459), .dinb(n407), .dout(n460));
  jand g00263(.dina(n460), .dinb(n457), .dout(n461));
  jor  g00264(.dina(n461), .dinb(n456), .dout(n462));
  jand g00265(.dina(n462), .dinb(asqrt[62] ), .dout(n463));
  jnot g00266(.din(n463), .dout(n464));
  jnot g00267(.din(n456), .dout(n465));
  jnot g00268(.din(n448), .dout(n466));
  jnot g00269(.din(n430), .dout(n467));
  jor  g00270(.dina(n443), .dinb(n354), .dout(n468));
  jnot g00271(.din(n428), .dout(n469));
  jand g00272(.dina(n469), .dinb(n468), .dout(n470));
  jand g00273(.dina(n470), .dinb(n352), .dout(n471));
  jor  g00274(.dina(n443), .dinb(a[116] ), .dout(n472));
  jand g00275(.dina(n472), .dinb(a[117] ), .dout(n473));
  jor  g00276(.dina(n450), .dinb(n473), .dout(n474));
  jor  g00277(.dina(n474), .dinb(n471), .dout(n475));
  jand g00278(.dina(n475), .dinb(n467), .dout(n476));
  jand g00279(.dina(n476), .dinb(n294), .dout(n477));
  jor  g00280(.dina(n452), .dinb(n477), .dout(n478));
  jand g00281(.dina(n478), .dinb(n466), .dout(n479));
  jand g00282(.dina(n479), .dinb(n239), .dout(n480));
  jnot g00283(.din(n460), .dout(n481));
  jor  g00284(.dina(n481), .dinb(n480), .dout(n482));
  jand g00285(.dina(n482), .dinb(n465), .dout(n483));
  jand g00286(.dina(n483), .dinb(n221), .dout(n484));
  jxor g00287(.dina(n367), .dinb(n239), .dout(n485));
  jand g00288(.dina(n485), .dinb(asqrt[58] ), .dout(n486));
  jxor g00289(.dina(n486), .dinb(n373), .dout(n487));
  jor  g00290(.dina(n487), .dinb(n484), .dout(n488));
  jand g00291(.dina(n488), .dinb(n464), .dout(n489));
  jor  g00292(.dina(n489), .dinb(n423), .dout(n490));
  jor  g00293(.dina(n490), .dinb(n387), .dout(n491));
  jor  g00294(.dina(n491), .dinb(n419), .dout(n492));
  jand g00295(.dina(n492), .dinb(n218), .dout(n493));
  jand g00296(.dina(n443), .dinb(n386), .dout(n494));
  jnot g00297(.din(n494), .dout(n495));
  jor  g00298(.dina(n462), .dinb(asqrt[62] ), .dout(n496));
  jnot g00299(.din(n487), .dout(n497));
  jand g00300(.dina(n497), .dinb(n496), .dout(n498));
  jor  g00301(.dina(n498), .dinb(n463), .dout(n499));
  jor  g00302(.dina(n499), .dinb(n422), .dout(n500));
  jand g00303(.dina(n500), .dinb(n495), .dout(n501));
  jand g00304(.dina(n443), .dinb(n383), .dout(n502));
  jnot g00305(.din(n502), .dout(n503));
  jand g00306(.dina(n389), .dinb(n435), .dout(n504));
  jand g00307(.dina(n504), .dinb(n503), .dout(n505));
  jnot g00308(.din(n505), .dout(n506));
  jand g00309(.dina(n506), .dinb(n501), .dout(n507));
  jnot g00310(.din(n507), .dout(n508));
  jor  g00311(.dina(n508), .dinb(n493), .dout(asqrt[57] ));
  jnot g00312(.din(n419), .dout(n510));
  jand g00313(.dina(n499), .dinb(n422), .dout(n511));
  jand g00314(.dina(n511), .dinb(n436), .dout(n512));
  jand g00315(.dina(n512), .dinb(n510), .dout(n513));
  jor  g00316(.dina(n513), .dinb(asqrt[63] ), .dout(n514));
  jand g00317(.dina(n507), .dinb(n514), .dout(n515));
  jxor g00318(.dina(n462), .dinb(n221), .dout(n516));
  jor  g00319(.dina(n516), .dinb(n515), .dout(n517));
  jxor g00320(.dina(n517), .dinb(n487), .dout(n518));
  jnot g00321(.din(n518), .dout(n519));
  jor  g00322(.dina(n515), .dinb(n425), .dout(n520));
  jnot g00323(.din(a[112] ), .dout(n521));
  jnot g00324(.din(a[113] ), .dout(n522));
  jand g00325(.dina(n522), .dinb(n521), .dout(n523));
  jand g00326(.dina(n523), .dinb(n425), .dout(n524));
  jnot g00327(.din(n524), .dout(n525));
  jand g00328(.dina(n525), .dinb(n520), .dout(n526));
  jor  g00329(.dina(n526), .dinb(n443), .dout(n527));
  jand g00330(.dina(n526), .dinb(n443), .dout(n528));
  jor  g00331(.dina(n515), .dinb(a[114] ), .dout(n529));
  jand g00332(.dina(n529), .dinb(a[115] ), .dout(n530));
  jand g00333(.dina(asqrt[57] ), .dinb(n427), .dout(n531));
  jor  g00334(.dina(n531), .dinb(n530), .dout(n532));
  jor  g00335(.dina(n532), .dinb(n528), .dout(n533));
  jand g00336(.dina(n533), .dinb(n527), .dout(n534));
  jor  g00337(.dina(n534), .dinb(n352), .dout(n535));
  jand g00338(.dina(n534), .dinb(n352), .dout(n536));
  jnot g00339(.din(n427), .dout(n537));
  jor  g00340(.dina(n515), .dinb(n537), .dout(n538));
  jnot g00341(.din(n500), .dout(n539));
  jor  g00342(.dina(n504), .dinb(n443), .dout(n540));
  jor  g00343(.dina(n540), .dinb(n539), .dout(n541));
  jor  g00344(.dina(n541), .dinb(n493), .dout(n542));
  jand g00345(.dina(n542), .dinb(n538), .dout(n543));
  jxor g00346(.dina(n543), .dinb(n354), .dout(n544));
  jor  g00347(.dina(n544), .dinb(n536), .dout(n545));
  jand g00348(.dina(n545), .dinb(n535), .dout(n546));
  jor  g00349(.dina(n546), .dinb(n294), .dout(n547));
  jand g00350(.dina(n546), .dinb(n294), .dout(n548));
  jxor g00351(.dina(n429), .dinb(n352), .dout(n549));
  jor  g00352(.dina(n549), .dinb(n515), .dout(n550));
  jxor g00353(.dina(n550), .dinb(n474), .dout(n551));
  jnot g00354(.din(n551), .dout(n552));
  jor  g00355(.dina(n552), .dinb(n548), .dout(n553));
  jand g00356(.dina(n553), .dinb(n547), .dout(n554));
  jor  g00357(.dina(n554), .dinb(n239), .dout(n555));
  jand g00358(.dina(n554), .dinb(n239), .dout(n556));
  jxor g00359(.dina(n447), .dinb(n294), .dout(n557));
  jor  g00360(.dina(n557), .dinb(n515), .dout(n558));
  jxor g00361(.dina(n558), .dinb(n453), .dout(n559));
  jor  g00362(.dina(n559), .dinb(n556), .dout(n560));
  jand g00363(.dina(n560), .dinb(n555), .dout(n561));
  jor  g00364(.dina(n561), .dinb(n221), .dout(n562));
  jand g00365(.dina(n561), .dinb(n221), .dout(n563));
  jxor g00366(.dina(n455), .dinb(n239), .dout(n564));
  jor  g00367(.dina(n564), .dinb(n515), .dout(n565));
  jxor g00368(.dina(n565), .dinb(n481), .dout(n566));
  jnot g00369(.din(n566), .dout(n567));
  jor  g00370(.dina(n567), .dinb(n563), .dout(n568));
  jand g00371(.dina(n568), .dinb(n562), .dout(n569));
  jor  g00372(.dina(n569), .dinb(n519), .dout(n570));
  jand g00373(.dina(asqrt[57] ), .dinb(n511), .dout(n571));
  jor  g00374(.dina(n571), .dinb(n539), .dout(n572));
  jor  g00375(.dina(n572), .dinb(n570), .dout(n573));
  jand g00376(.dina(n573), .dinb(n218), .dout(n574));
  jand g00377(.dina(n515), .dinb(n423), .dout(n575));
  jand g00378(.dina(n569), .dinb(n519), .dout(n576));
  jor  g00379(.dina(n576), .dinb(n575), .dout(n577));
  jand g00380(.dina(n515), .dinb(n489), .dout(n578));
  jand g00381(.dina(n490), .dinb(asqrt[63] ), .dout(n579));
  jand g00382(.dina(n579), .dinb(n500), .dout(n580));
  jnot g00383(.din(n580), .dout(n581));
  jor  g00384(.dina(n581), .dinb(n578), .dout(n582));
  jnot g00385(.din(n582), .dout(n583));
  jor  g00386(.dina(n583), .dinb(n577), .dout(n584));
  jor  g00387(.dina(n584), .dinb(n574), .dout(asqrt[56] ));
  jxor g00388(.dina(n561), .dinb(n221), .dout(n586));
  jand g00389(.dina(n586), .dinb(asqrt[56] ), .dout(n587));
  jxor g00390(.dina(n587), .dinb(n566), .dout(n588));
  jnot g00391(.din(a[110] ), .dout(n589));
  jnot g00392(.din(a[111] ), .dout(n590));
  jand g00393(.dina(n590), .dinb(n589), .dout(n591));
  jand g00394(.dina(n591), .dinb(n521), .dout(n592));
  jand g00395(.dina(asqrt[56] ), .dinb(a[112] ), .dout(n593));
  jor  g00396(.dina(n593), .dinb(n592), .dout(n594));
  jand g00397(.dina(n594), .dinb(asqrt[57] ), .dout(n595));
  jor  g00398(.dina(n594), .dinb(asqrt[57] ), .dout(n596));
  jand g00399(.dina(asqrt[56] ), .dinb(n521), .dout(n597));
  jor  g00400(.dina(n597), .dinb(n522), .dout(n598));
  jnot g00401(.din(n523), .dout(n599));
  jnot g00402(.din(n562), .dout(n600));
  jnot g00403(.din(n555), .dout(n601));
  jnot g00404(.din(n547), .dout(n602));
  jnot g00405(.din(n535), .dout(n603));
  jnot g00406(.din(n527), .dout(n604));
  jand g00407(.dina(asqrt[57] ), .dinb(a[114] ), .dout(n605));
  jor  g00408(.dina(n524), .dinb(n605), .dout(n606));
  jor  g00409(.dina(n606), .dinb(asqrt[58] ), .dout(n607));
  jand g00410(.dina(asqrt[57] ), .dinb(n425), .dout(n608));
  jor  g00411(.dina(n608), .dinb(n426), .dout(n609));
  jand g00412(.dina(n538), .dinb(n609), .dout(n610));
  jand g00413(.dina(n610), .dinb(n607), .dout(n611));
  jor  g00414(.dina(n611), .dinb(n604), .dout(n612));
  jor  g00415(.dina(n612), .dinb(asqrt[59] ), .dout(n613));
  jnot g00416(.din(n544), .dout(n614));
  jand g00417(.dina(n614), .dinb(n613), .dout(n615));
  jor  g00418(.dina(n615), .dinb(n603), .dout(n616));
  jor  g00419(.dina(n616), .dinb(asqrt[60] ), .dout(n617));
  jand g00420(.dina(n551), .dinb(n617), .dout(n618));
  jor  g00421(.dina(n618), .dinb(n602), .dout(n619));
  jor  g00422(.dina(n619), .dinb(asqrt[61] ), .dout(n620));
  jnot g00423(.din(n559), .dout(n621));
  jand g00424(.dina(n621), .dinb(n620), .dout(n622));
  jor  g00425(.dina(n622), .dinb(n601), .dout(n623));
  jor  g00426(.dina(n623), .dinb(asqrt[62] ), .dout(n624));
  jand g00427(.dina(n566), .dinb(n624), .dout(n625));
  jor  g00428(.dina(n625), .dinb(n600), .dout(n626));
  jand g00429(.dina(n626), .dinb(n518), .dout(n627));
  jnot g00430(.din(n572), .dout(n628));
  jand g00431(.dina(n628), .dinb(n627), .dout(n629));
  jor  g00432(.dina(n629), .dinb(asqrt[63] ), .dout(n630));
  jnot g00433(.din(n575), .dout(n631));
  jor  g00434(.dina(n626), .dinb(n518), .dout(n632));
  jand g00435(.dina(n632), .dinb(n631), .dout(n633));
  jand g00436(.dina(n582), .dinb(n633), .dout(n634));
  jand g00437(.dina(n634), .dinb(n630), .dout(n635));
  jor  g00438(.dina(n635), .dinb(n599), .dout(n636));
  jand g00439(.dina(n636), .dinb(n598), .dout(n637));
  jand g00440(.dina(n637), .dinb(n596), .dout(n638));
  jor  g00441(.dina(n638), .dinb(n595), .dout(n639));
  jand g00442(.dina(n639), .dinb(asqrt[58] ), .dout(n640));
  jor  g00443(.dina(n639), .dinb(asqrt[58] ), .dout(n641));
  jand g00444(.dina(asqrt[56] ), .dinb(n523), .dout(n642));
  jand g00445(.dina(n581), .dinb(asqrt[57] ), .dout(n643));
  jand g00446(.dina(n643), .dinb(n632), .dout(n644));
  jand g00447(.dina(n644), .dinb(n630), .dout(n645));
  jor  g00448(.dina(n645), .dinb(n642), .dout(n646));
  jxor g00449(.dina(n646), .dinb(a[114] ), .dout(n647));
  jnot g00450(.din(n647), .dout(n648));
  jand g00451(.dina(n648), .dinb(n641), .dout(n649));
  jor  g00452(.dina(n649), .dinb(n640), .dout(n650));
  jand g00453(.dina(n650), .dinb(asqrt[59] ), .dout(n651));
  jor  g00454(.dina(n650), .dinb(asqrt[59] ), .dout(n652));
  jxor g00455(.dina(n526), .dinb(n443), .dout(n653));
  jand g00456(.dina(n653), .dinb(asqrt[56] ), .dout(n654));
  jxor g00457(.dina(n654), .dinb(n610), .dout(n655));
  jand g00458(.dina(n655), .dinb(n652), .dout(n656));
  jor  g00459(.dina(n656), .dinb(n651), .dout(n657));
  jand g00460(.dina(n657), .dinb(asqrt[60] ), .dout(n658));
  jor  g00461(.dina(n657), .dinb(asqrt[60] ), .dout(n659));
  jxor g00462(.dina(n534), .dinb(n352), .dout(n660));
  jand g00463(.dina(n660), .dinb(asqrt[56] ), .dout(n661));
  jxor g00464(.dina(n661), .dinb(n544), .dout(n662));
  jnot g00465(.din(n662), .dout(n663));
  jand g00466(.dina(n663), .dinb(n659), .dout(n664));
  jor  g00467(.dina(n664), .dinb(n658), .dout(n665));
  jand g00468(.dina(n665), .dinb(asqrt[61] ), .dout(n666));
  jor  g00469(.dina(n665), .dinb(asqrt[61] ), .dout(n667));
  jxor g00470(.dina(n546), .dinb(n294), .dout(n668));
  jand g00471(.dina(n668), .dinb(asqrt[56] ), .dout(n669));
  jxor g00472(.dina(n669), .dinb(n551), .dout(n670));
  jand g00473(.dina(n670), .dinb(n667), .dout(n671));
  jor  g00474(.dina(n671), .dinb(n666), .dout(n672));
  jand g00475(.dina(n672), .dinb(asqrt[62] ), .dout(n673));
  jor  g00476(.dina(n672), .dinb(asqrt[62] ), .dout(n674));
  jxor g00477(.dina(n554), .dinb(n239), .dout(n675));
  jand g00478(.dina(n675), .dinb(asqrt[56] ), .dout(n676));
  jxor g00479(.dina(n676), .dinb(n559), .dout(n677));
  jnot g00480(.din(n677), .dout(n678));
  jand g00481(.dina(n678), .dinb(n674), .dout(n679));
  jor  g00482(.dina(n679), .dinb(n673), .dout(n680));
  jor  g00483(.dina(n680), .dinb(n588), .dout(n681));
  jnot g00484(.din(n681), .dout(n682));
  jand g00485(.dina(n635), .dinb(n569), .dout(n683));
  jnot g00486(.din(n683), .dout(n684));
  jand g00487(.dina(n570), .dinb(asqrt[63] ), .dout(n685));
  jand g00488(.dina(n685), .dinb(n632), .dout(n686));
  jand g00489(.dina(n686), .dinb(n684), .dout(n687));
  jnot g00490(.din(n588), .dout(n688));
  jnot g00491(.din(n673), .dout(n689));
  jnot g00492(.din(n666), .dout(n690));
  jnot g00493(.din(n658), .dout(n691));
  jnot g00494(.din(n651), .dout(n692));
  jnot g00495(.din(n640), .dout(n693));
  jnot g00496(.din(n595), .dout(n694));
  jnot g00497(.din(n592), .dout(n695));
  jor  g00498(.dina(n635), .dinb(n521), .dout(n696));
  jand g00499(.dina(n696), .dinb(n695), .dout(n697));
  jand g00500(.dina(n697), .dinb(n515), .dout(n698));
  jor  g00501(.dina(n635), .dinb(a[112] ), .dout(n699));
  jand g00502(.dina(n699), .dinb(a[113] ), .dout(n700));
  jor  g00503(.dina(n642), .dinb(n700), .dout(n701));
  jor  g00504(.dina(n701), .dinb(n698), .dout(n702));
  jand g00505(.dina(n702), .dinb(n694), .dout(n703));
  jand g00506(.dina(n703), .dinb(n443), .dout(n704));
  jor  g00507(.dina(n647), .dinb(n704), .dout(n705));
  jand g00508(.dina(n705), .dinb(n693), .dout(n706));
  jand g00509(.dina(n706), .dinb(n352), .dout(n707));
  jnot g00510(.din(n655), .dout(n708));
  jor  g00511(.dina(n708), .dinb(n707), .dout(n709));
  jand g00512(.dina(n709), .dinb(n692), .dout(n710));
  jand g00513(.dina(n710), .dinb(n294), .dout(n711));
  jor  g00514(.dina(n662), .dinb(n711), .dout(n712));
  jand g00515(.dina(n712), .dinb(n691), .dout(n713));
  jand g00516(.dina(n713), .dinb(n239), .dout(n714));
  jnot g00517(.din(n670), .dout(n715));
  jor  g00518(.dina(n715), .dinb(n714), .dout(n716));
  jand g00519(.dina(n716), .dinb(n690), .dout(n717));
  jand g00520(.dina(n717), .dinb(n221), .dout(n718));
  jor  g00521(.dina(n677), .dinb(n718), .dout(n719));
  jand g00522(.dina(n719), .dinb(n689), .dout(n720));
  jor  g00523(.dina(n720), .dinb(n688), .dout(n721));
  jand g00524(.dina(asqrt[56] ), .dinb(n627), .dout(n722));
  jor  g00525(.dina(n722), .dinb(n576), .dout(n723));
  jor  g00526(.dina(n723), .dinb(n721), .dout(n724));
  jand g00527(.dina(n724), .dinb(n218), .dout(n725));
  jand g00528(.dina(n635), .dinb(n519), .dout(n726));
  jor  g00529(.dina(n726), .dinb(n725), .dout(n727));
  jor  g00530(.dina(n727), .dinb(n687), .dout(n728));
  jor  g00531(.dina(n728), .dinb(n682), .dout(asqrt[55] ));
  jnot g00532(.din(a[108] ), .dout(n730));
  jnot g00533(.din(a[109] ), .dout(n731));
  jand g00534(.dina(n731), .dinb(n730), .dout(n732));
  jand g00535(.dina(n732), .dinb(n589), .dout(n733));
  jnot g00536(.din(n733), .dout(n734));
  jnot g00537(.din(n687), .dout(n735));
  jand g00538(.dina(n680), .dinb(n588), .dout(n736));
  jnot g00539(.din(n723), .dout(n737));
  jand g00540(.dina(n737), .dinb(n736), .dout(n738));
  jor  g00541(.dina(n738), .dinb(asqrt[63] ), .dout(n739));
  jnot g00542(.din(n726), .dout(n740));
  jand g00543(.dina(n740), .dinb(n739), .dout(n741));
  jand g00544(.dina(n741), .dinb(n735), .dout(n742));
  jand g00545(.dina(n742), .dinb(n681), .dout(n743));
  jor  g00546(.dina(n743), .dinb(n589), .dout(n744));
  jand g00547(.dina(n744), .dinb(n734), .dout(n745));
  jor  g00548(.dina(n745), .dinb(n635), .dout(n746));
  jand g00549(.dina(n745), .dinb(n635), .dout(n747));
  jor  g00550(.dina(n743), .dinb(a[110] ), .dout(n748));
  jand g00551(.dina(n748), .dinb(a[111] ), .dout(n749));
  jand g00552(.dina(asqrt[55] ), .dinb(n591), .dout(n750));
  jor  g00553(.dina(n750), .dinb(n749), .dout(n751));
  jor  g00554(.dina(n751), .dinb(n747), .dout(n752));
  jand g00555(.dina(n752), .dinb(n746), .dout(n753));
  jor  g00556(.dina(n753), .dinb(n515), .dout(n754));
  jand g00557(.dina(n753), .dinb(n515), .dout(n755));
  jnot g00558(.din(n591), .dout(n756));
  jor  g00559(.dina(n743), .dinb(n756), .dout(n757));
  jor  g00560(.dina(n682), .dinb(n635), .dout(n758));
  jor  g00561(.dina(n758), .dinb(n686), .dout(n759));
  jor  g00562(.dina(n759), .dinb(n725), .dout(n760));
  jand g00563(.dina(n760), .dinb(n757), .dout(n761));
  jxor g00564(.dina(n761), .dinb(n521), .dout(n762));
  jor  g00565(.dina(n762), .dinb(n755), .dout(n763));
  jand g00566(.dina(n763), .dinb(n754), .dout(n764));
  jor  g00567(.dina(n764), .dinb(n443), .dout(n765));
  jand g00568(.dina(n764), .dinb(n443), .dout(n766));
  jxor g00569(.dina(n594), .dinb(n515), .dout(n767));
  jor  g00570(.dina(n767), .dinb(n743), .dout(n768));
  jxor g00571(.dina(n768), .dinb(n701), .dout(n769));
  jnot g00572(.din(n769), .dout(n770));
  jor  g00573(.dina(n770), .dinb(n766), .dout(n771));
  jand g00574(.dina(n771), .dinb(n765), .dout(n772));
  jor  g00575(.dina(n772), .dinb(n352), .dout(n773));
  jand g00576(.dina(n772), .dinb(n352), .dout(n774));
  jxor g00577(.dina(n639), .dinb(n443), .dout(n775));
  jor  g00578(.dina(n775), .dinb(n743), .dout(n776));
  jxor g00579(.dina(n776), .dinb(n648), .dout(n777));
  jor  g00580(.dina(n777), .dinb(n774), .dout(n778));
  jand g00581(.dina(n778), .dinb(n773), .dout(n779));
  jor  g00582(.dina(n779), .dinb(n294), .dout(n780));
  jand g00583(.dina(n779), .dinb(n294), .dout(n781));
  jxor g00584(.dina(n650), .dinb(n352), .dout(n782));
  jor  g00585(.dina(n782), .dinb(n743), .dout(n783));
  jxor g00586(.dina(n783), .dinb(n708), .dout(n784));
  jnot g00587(.din(n784), .dout(n785));
  jor  g00588(.dina(n785), .dinb(n781), .dout(n786));
  jand g00589(.dina(n786), .dinb(n780), .dout(n787));
  jor  g00590(.dina(n787), .dinb(n239), .dout(n788));
  jand g00591(.dina(n787), .dinb(n239), .dout(n789));
  jxor g00592(.dina(n657), .dinb(n294), .dout(n790));
  jor  g00593(.dina(n790), .dinb(n743), .dout(n791));
  jxor g00594(.dina(n791), .dinb(n663), .dout(n792));
  jor  g00595(.dina(n792), .dinb(n789), .dout(n793));
  jand g00596(.dina(n793), .dinb(n788), .dout(n794));
  jor  g00597(.dina(n794), .dinb(n221), .dout(n795));
  jand g00598(.dina(n794), .dinb(n221), .dout(n796));
  jxor g00599(.dina(n665), .dinb(n239), .dout(n797));
  jor  g00600(.dina(n797), .dinb(n743), .dout(n798));
  jxor g00601(.dina(n798), .dinb(n715), .dout(n799));
  jnot g00602(.din(n799), .dout(n800));
  jor  g00603(.dina(n800), .dinb(n796), .dout(n801));
  jand g00604(.dina(n801), .dinb(n795), .dout(n802));
  jxor g00605(.dina(n672), .dinb(n221), .dout(n803));
  jor  g00606(.dina(n803), .dinb(n743), .dout(n804));
  jxor g00607(.dina(n804), .dinb(n678), .dout(n805));
  jand g00608(.dina(n805), .dinb(n802), .dout(n806));
  jand g00609(.dina(n728), .dinb(n736), .dout(n808));
  jor  g00610(.dina(n805), .dinb(n802), .dout(n809));
  jor  g00611(.dina(n809), .dinb(n682), .dout(n810));
  jor  g00612(.dina(n810), .dinb(n808), .dout(n811));
  jand g00613(.dina(n811), .dinb(n218), .dout(n812));
  jand g00614(.dina(n742), .dinb(n720), .dout(n813));
  jand g00615(.dina(n721), .dinb(asqrt[63] ), .dout(n814));
  jand g00616(.dina(n814), .dinb(n681), .dout(n815));
  jnot g00617(.din(n815), .dout(n816));
  jor  g00618(.dina(n816), .dinb(n813), .dout(n817));
  jnot g00619(.din(n817), .dout(n818));
  jor  g00620(.dina(n818), .dinb(n812), .dout(n819));
  jor  g00621(.dina(n819), .dinb(n806), .dout(asqrt[54] ));
  jnot g00622(.din(n795), .dout(n822));
  jnot g00623(.din(n788), .dout(n823));
  jnot g00624(.din(n780), .dout(n824));
  jnot g00625(.din(n773), .dout(n825));
  jnot g00626(.din(n765), .dout(n826));
  jnot g00627(.din(n754), .dout(n827));
  jnot g00628(.din(n746), .dout(n828));
  jand g00629(.dina(asqrt[55] ), .dinb(a[110] ), .dout(n829));
  jor  g00630(.dina(n829), .dinb(n733), .dout(n830));
  jor  g00631(.dina(n830), .dinb(asqrt[56] ), .dout(n831));
  jand g00632(.dina(asqrt[55] ), .dinb(n589), .dout(n832));
  jor  g00633(.dina(n832), .dinb(n590), .dout(n833));
  jand g00634(.dina(n757), .dinb(n833), .dout(n834));
  jand g00635(.dina(n834), .dinb(n831), .dout(n835));
  jor  g00636(.dina(n835), .dinb(n828), .dout(n836));
  jor  g00637(.dina(n836), .dinb(asqrt[57] ), .dout(n837));
  jnot g00638(.din(n762), .dout(n838));
  jand g00639(.dina(n838), .dinb(n837), .dout(n839));
  jor  g00640(.dina(n839), .dinb(n827), .dout(n840));
  jor  g00641(.dina(n840), .dinb(asqrt[58] ), .dout(n841));
  jand g00642(.dina(n769), .dinb(n841), .dout(n842));
  jor  g00643(.dina(n842), .dinb(n826), .dout(n843));
  jor  g00644(.dina(n843), .dinb(asqrt[59] ), .dout(n844));
  jnot g00645(.din(n777), .dout(n845));
  jand g00646(.dina(n845), .dinb(n844), .dout(n846));
  jor  g00647(.dina(n846), .dinb(n825), .dout(n847));
  jor  g00648(.dina(n847), .dinb(asqrt[60] ), .dout(n848));
  jand g00649(.dina(n784), .dinb(n848), .dout(n849));
  jor  g00650(.dina(n849), .dinb(n824), .dout(n850));
  jor  g00651(.dina(n850), .dinb(asqrt[61] ), .dout(n851));
  jnot g00652(.din(n792), .dout(n852));
  jand g00653(.dina(n852), .dinb(n851), .dout(n853));
  jor  g00654(.dina(n853), .dinb(n823), .dout(n854));
  jor  g00655(.dina(n854), .dinb(asqrt[62] ), .dout(n855));
  jand g00656(.dina(n799), .dinb(n855), .dout(n856));
  jor  g00657(.dina(n856), .dinb(n822), .dout(n857));
  jnot g00658(.din(n805), .dout(n858));
  jand g00659(.dina(n858), .dinb(n857), .dout(n859));
  jand g00660(.dina(n819), .dinb(n859), .dout(n860));
  jxor g00661(.dina(n794), .dinb(n221), .dout(n861));
  jand g00662(.dina(n861), .dinb(asqrt[54] ), .dout(n862));
  jxor g00663(.dina(n862), .dinb(n799), .dout(n863));
  jnot g00664(.din(n863), .dout(n864));
  jnot g00665(.din(a[106] ), .dout(n865));
  jnot g00666(.din(a[107] ), .dout(n866));
  jand g00667(.dina(n866), .dinb(n865), .dout(n867));
  jand g00668(.dina(n867), .dinb(n730), .dout(n868));
  jand g00669(.dina(asqrt[54] ), .dinb(a[108] ), .dout(n869));
  jor  g00670(.dina(n869), .dinb(n868), .dout(n870));
  jand g00671(.dina(n870), .dinb(asqrt[55] ), .dout(n871));
  jor  g00672(.dina(n870), .dinb(asqrt[55] ), .dout(n872));
  jand g00673(.dina(asqrt[54] ), .dinb(n730), .dout(n873));
  jor  g00674(.dina(n873), .dinb(n731), .dout(n874));
  jnot g00675(.din(n732), .dout(n875));
  jnot g00676(.din(n806), .dout(n876));
  jnot g00677(.din(n808), .dout(n878));
  jand g00678(.dina(n859), .dinb(n681), .dout(n879));
  jand g00679(.dina(n879), .dinb(n878), .dout(n880));
  jor  g00680(.dina(n880), .dinb(asqrt[63] ), .dout(n881));
  jand g00681(.dina(n817), .dinb(n881), .dout(n882));
  jand g00682(.dina(n882), .dinb(n876), .dout(n884));
  jor  g00683(.dina(n884), .dinb(n875), .dout(n885));
  jand g00684(.dina(n885), .dinb(n874), .dout(n886));
  jand g00685(.dina(n886), .dinb(n872), .dout(n887));
  jor  g00686(.dina(n887), .dinb(n871), .dout(n888));
  jand g00687(.dina(n888), .dinb(asqrt[56] ), .dout(n889));
  jor  g00688(.dina(n888), .dinb(asqrt[56] ), .dout(n890));
  jand g00689(.dina(asqrt[54] ), .dinb(n732), .dout(n891));
  jand g00690(.dina(n816), .dinb(n876), .dout(n892));
  jand g00691(.dina(n892), .dinb(n881), .dout(n893));
  jand g00692(.dina(n893), .dinb(asqrt[55] ), .dout(n894));
  jor  g00693(.dina(n894), .dinb(n891), .dout(n895));
  jxor g00694(.dina(n895), .dinb(a[110] ), .dout(n896));
  jnot g00695(.din(n896), .dout(n897));
  jand g00696(.dina(n897), .dinb(n890), .dout(n898));
  jor  g00697(.dina(n898), .dinb(n889), .dout(n899));
  jand g00698(.dina(n899), .dinb(asqrt[57] ), .dout(n900));
  jor  g00699(.dina(n899), .dinb(asqrt[57] ), .dout(n901));
  jxor g00700(.dina(n745), .dinb(n635), .dout(n902));
  jand g00701(.dina(n902), .dinb(asqrt[54] ), .dout(n903));
  jxor g00702(.dina(n903), .dinb(n834), .dout(n904));
  jand g00703(.dina(n904), .dinb(n901), .dout(n905));
  jor  g00704(.dina(n905), .dinb(n900), .dout(n906));
  jand g00705(.dina(n906), .dinb(asqrt[58] ), .dout(n907));
  jor  g00706(.dina(n906), .dinb(asqrt[58] ), .dout(n908));
  jxor g00707(.dina(n753), .dinb(n515), .dout(n909));
  jand g00708(.dina(n909), .dinb(asqrt[54] ), .dout(n910));
  jxor g00709(.dina(n910), .dinb(n838), .dout(n911));
  jand g00710(.dina(n911), .dinb(n908), .dout(n912));
  jor  g00711(.dina(n912), .dinb(n907), .dout(n913));
  jand g00712(.dina(n913), .dinb(asqrt[59] ), .dout(n914));
  jor  g00713(.dina(n913), .dinb(asqrt[59] ), .dout(n915));
  jxor g00714(.dina(n764), .dinb(n443), .dout(n916));
  jand g00715(.dina(n916), .dinb(asqrt[54] ), .dout(n917));
  jxor g00716(.dina(n917), .dinb(n769), .dout(n918));
  jand g00717(.dina(n918), .dinb(n915), .dout(n919));
  jor  g00718(.dina(n919), .dinb(n914), .dout(n920));
  jand g00719(.dina(n920), .dinb(asqrt[60] ), .dout(n921));
  jor  g00720(.dina(n920), .dinb(asqrt[60] ), .dout(n922));
  jxor g00721(.dina(n772), .dinb(n352), .dout(n923));
  jand g00722(.dina(n923), .dinb(asqrt[54] ), .dout(n924));
  jxor g00723(.dina(n924), .dinb(n777), .dout(n925));
  jnot g00724(.din(n925), .dout(n926));
  jand g00725(.dina(n926), .dinb(n922), .dout(n927));
  jor  g00726(.dina(n927), .dinb(n921), .dout(n928));
  jand g00727(.dina(n928), .dinb(asqrt[61] ), .dout(n929));
  jor  g00728(.dina(n928), .dinb(asqrt[61] ), .dout(n930));
  jxor g00729(.dina(n779), .dinb(n294), .dout(n931));
  jand g00730(.dina(n931), .dinb(asqrt[54] ), .dout(n932));
  jxor g00731(.dina(n932), .dinb(n784), .dout(n933));
  jand g00732(.dina(n933), .dinb(n930), .dout(n934));
  jor  g00733(.dina(n934), .dinb(n929), .dout(n935));
  jand g00734(.dina(n935), .dinb(asqrt[62] ), .dout(n936));
  jnot g00735(.din(n936), .dout(n937));
  jnot g00736(.din(n929), .dout(n938));
  jnot g00737(.din(n921), .dout(n939));
  jnot g00738(.din(n914), .dout(n940));
  jnot g00739(.din(n907), .dout(n941));
  jnot g00740(.din(n900), .dout(n942));
  jnot g00741(.din(n889), .dout(n943));
  jnot g00742(.din(n871), .dout(n944));
  jnot g00743(.din(n868), .dout(n945));
  jor  g00744(.dina(n884), .dinb(n730), .dout(n946));
  jand g00745(.dina(n946), .dinb(n945), .dout(n947));
  jand g00746(.dina(n947), .dinb(n743), .dout(n948));
  jor  g00747(.dina(n884), .dinb(a[108] ), .dout(n949));
  jand g00748(.dina(n949), .dinb(a[109] ), .dout(n950));
  jor  g00749(.dina(n891), .dinb(n950), .dout(n951));
  jor  g00750(.dina(n951), .dinb(n948), .dout(n952));
  jand g00751(.dina(n952), .dinb(n944), .dout(n953));
  jand g00752(.dina(n953), .dinb(n635), .dout(n954));
  jor  g00753(.dina(n896), .dinb(n954), .dout(n955));
  jand g00754(.dina(n955), .dinb(n943), .dout(n956));
  jand g00755(.dina(n956), .dinb(n515), .dout(n957));
  jnot g00756(.din(n904), .dout(n958));
  jor  g00757(.dina(n958), .dinb(n957), .dout(n959));
  jand g00758(.dina(n959), .dinb(n942), .dout(n960));
  jand g00759(.dina(n960), .dinb(n443), .dout(n961));
  jnot g00760(.din(n911), .dout(n962));
  jor  g00761(.dina(n962), .dinb(n961), .dout(n963));
  jand g00762(.dina(n963), .dinb(n941), .dout(n964));
  jand g00763(.dina(n964), .dinb(n352), .dout(n965));
  jnot g00764(.din(n918), .dout(n966));
  jor  g00765(.dina(n966), .dinb(n965), .dout(n967));
  jand g00766(.dina(n967), .dinb(n940), .dout(n968));
  jand g00767(.dina(n968), .dinb(n294), .dout(n969));
  jor  g00768(.dina(n925), .dinb(n969), .dout(n970));
  jand g00769(.dina(n970), .dinb(n939), .dout(n971));
  jand g00770(.dina(n971), .dinb(n239), .dout(n972));
  jnot g00771(.din(n933), .dout(n973));
  jor  g00772(.dina(n973), .dinb(n972), .dout(n974));
  jand g00773(.dina(n974), .dinb(n938), .dout(n975));
  jand g00774(.dina(n975), .dinb(n221), .dout(n976));
  jxor g00775(.dina(n787), .dinb(n239), .dout(n977));
  jand g00776(.dina(n977), .dinb(asqrt[54] ), .dout(n978));
  jxor g00777(.dina(n978), .dinb(n792), .dout(n979));
  jor  g00778(.dina(n979), .dinb(n976), .dout(n980));
  jand g00779(.dina(n980), .dinb(n937), .dout(n981));
  jor  g00780(.dina(n981), .dinb(n864), .dout(n982));
  jor  g00781(.dina(n982), .dinb(n806), .dout(n983));
  jor  g00782(.dina(n983), .dinb(n860), .dout(n984));
  jand g00783(.dina(n984), .dinb(n218), .dout(n985));
  jand g00784(.dina(n884), .dinb(n805), .dout(n986));
  jnot g00785(.din(n986), .dout(n987));
  jor  g00786(.dina(n935), .dinb(asqrt[62] ), .dout(n988));
  jnot g00787(.din(n979), .dout(n989));
  jand g00788(.dina(n989), .dinb(n988), .dout(n990));
  jor  g00789(.dina(n990), .dinb(n936), .dout(n991));
  jor  g00790(.dina(n991), .dinb(n863), .dout(n992));
  jand g00791(.dina(n992), .dinb(n987), .dout(n993));
  jand g00792(.dina(n882), .dinb(n802), .dout(n994));
  jnot g00793(.din(n994), .dout(n995));
  jand g00794(.dina(n809), .dinb(asqrt[63] ), .dout(n996));
  jand g00795(.dina(n996), .dinb(n876), .dout(n997));
  jand g00796(.dina(n997), .dinb(n995), .dout(n998));
  jnot g00797(.din(n998), .dout(n999));
  jand g00798(.dina(n999), .dinb(n993), .dout(n1000));
  jnot g00799(.din(n1000), .dout(n1001));
  jor  g00800(.dina(n1001), .dinb(n985), .dout(asqrt[53] ));
  jnot g00801(.din(n860), .dout(n1003));
  jand g00802(.dina(n991), .dinb(n863), .dout(n1004));
  jand g00803(.dina(n1004), .dinb(n876), .dout(n1005));
  jand g00804(.dina(n1005), .dinb(n1003), .dout(n1006));
  jor  g00805(.dina(n1006), .dinb(asqrt[63] ), .dout(n1007));
  jand g00806(.dina(n1000), .dinb(n1007), .dout(n1008));
  jor  g00807(.dina(n1008), .dinb(n865), .dout(n1009));
  jnot g00808(.din(a[104] ), .dout(n1010));
  jnot g00809(.din(a[105] ), .dout(n1011));
  jand g00810(.dina(n1011), .dinb(n1010), .dout(n1012));
  jand g00811(.dina(n1012), .dinb(n865), .dout(n1013));
  jnot g00812(.din(n1013), .dout(n1014));
  jand g00813(.dina(n1014), .dinb(n1009), .dout(n1015));
  jor  g00814(.dina(n1015), .dinb(n884), .dout(n1016));
  jand g00815(.dina(n1015), .dinb(n884), .dout(n1017));
  jor  g00816(.dina(n1008), .dinb(a[106] ), .dout(n1018));
  jand g00817(.dina(n1018), .dinb(a[107] ), .dout(n1019));
  jand g00818(.dina(asqrt[53] ), .dinb(n867), .dout(n1020));
  jor  g00819(.dina(n1020), .dinb(n1019), .dout(n1021));
  jor  g00820(.dina(n1021), .dinb(n1017), .dout(n1022));
  jand g00821(.dina(n1022), .dinb(n1016), .dout(n1023));
  jor  g00822(.dina(n1023), .dinb(n743), .dout(n1024));
  jand g00823(.dina(n1023), .dinb(n743), .dout(n1025));
  jnot g00824(.din(n867), .dout(n1026));
  jor  g00825(.dina(n1008), .dinb(n1026), .dout(n1027));
  jnot g00826(.din(n992), .dout(n1028));
  jor  g00827(.dina(n997), .dinb(n884), .dout(n1029));
  jor  g00828(.dina(n1029), .dinb(n985), .dout(n1030));
  jor  g00829(.dina(n1030), .dinb(n1028), .dout(n1031));
  jand g00830(.dina(n1031), .dinb(n1027), .dout(n1032));
  jxor g00831(.dina(n1032), .dinb(n730), .dout(n1033));
  jor  g00832(.dina(n1033), .dinb(n1025), .dout(n1034));
  jand g00833(.dina(n1034), .dinb(n1024), .dout(n1035));
  jor  g00834(.dina(n1035), .dinb(n635), .dout(n1036));
  jand g00835(.dina(n1035), .dinb(n635), .dout(n1037));
  jxor g00836(.dina(n870), .dinb(n743), .dout(n1038));
  jor  g00837(.dina(n1038), .dinb(n1008), .dout(n1039));
  jxor g00838(.dina(n1039), .dinb(n886), .dout(n1040));
  jor  g00839(.dina(n1040), .dinb(n1037), .dout(n1041));
  jand g00840(.dina(n1041), .dinb(n1036), .dout(n1042));
  jor  g00841(.dina(n1042), .dinb(n515), .dout(n1043));
  jand g00842(.dina(n1042), .dinb(n515), .dout(n1044));
  jxor g00843(.dina(n888), .dinb(n635), .dout(n1045));
  jor  g00844(.dina(n1045), .dinb(n1008), .dout(n1046));
  jxor g00845(.dina(n1046), .dinb(n897), .dout(n1047));
  jor  g00846(.dina(n1047), .dinb(n1044), .dout(n1048));
  jand g00847(.dina(n1048), .dinb(n1043), .dout(n1049));
  jor  g00848(.dina(n1049), .dinb(n443), .dout(n1050));
  jand g00849(.dina(n1049), .dinb(n443), .dout(n1051));
  jxor g00850(.dina(n899), .dinb(n515), .dout(n1052));
  jor  g00851(.dina(n1052), .dinb(n1008), .dout(n1053));
  jxor g00852(.dina(n1053), .dinb(n958), .dout(n1054));
  jnot g00853(.din(n1054), .dout(n1055));
  jor  g00854(.dina(n1055), .dinb(n1051), .dout(n1056));
  jand g00855(.dina(n1056), .dinb(n1050), .dout(n1057));
  jor  g00856(.dina(n1057), .dinb(n352), .dout(n1058));
  jand g00857(.dina(n1057), .dinb(n352), .dout(n1059));
  jxor g00858(.dina(n906), .dinb(n443), .dout(n1060));
  jor  g00859(.dina(n1060), .dinb(n1008), .dout(n1061));
  jxor g00860(.dina(n1061), .dinb(n962), .dout(n1062));
  jnot g00861(.din(n1062), .dout(n1063));
  jor  g00862(.dina(n1063), .dinb(n1059), .dout(n1064));
  jand g00863(.dina(n1064), .dinb(n1058), .dout(n1065));
  jor  g00864(.dina(n1065), .dinb(n294), .dout(n1066));
  jand g00865(.dina(n1065), .dinb(n294), .dout(n1067));
  jxor g00866(.dina(n913), .dinb(n352), .dout(n1068));
  jor  g00867(.dina(n1068), .dinb(n1008), .dout(n1069));
  jxor g00868(.dina(n1069), .dinb(n966), .dout(n1070));
  jnot g00869(.din(n1070), .dout(n1071));
  jor  g00870(.dina(n1071), .dinb(n1067), .dout(n1072));
  jand g00871(.dina(n1072), .dinb(n1066), .dout(n1073));
  jor  g00872(.dina(n1073), .dinb(n239), .dout(n1074));
  jand g00873(.dina(n1073), .dinb(n239), .dout(n1075));
  jxor g00874(.dina(n920), .dinb(n294), .dout(n1076));
  jor  g00875(.dina(n1076), .dinb(n1008), .dout(n1077));
  jxor g00876(.dina(n1077), .dinb(n926), .dout(n1078));
  jor  g00877(.dina(n1078), .dinb(n1075), .dout(n1079));
  jand g00878(.dina(n1079), .dinb(n1074), .dout(n1080));
  jor  g00879(.dina(n1080), .dinb(n221), .dout(n1081));
  jand g00880(.dina(n1080), .dinb(n221), .dout(n1082));
  jxor g00881(.dina(n928), .dinb(n239), .dout(n1083));
  jor  g00882(.dina(n1083), .dinb(n1008), .dout(n1084));
  jxor g00883(.dina(n1084), .dinb(n973), .dout(n1085));
  jnot g00884(.din(n1085), .dout(n1086));
  jor  g00885(.dina(n1086), .dinb(n1082), .dout(n1087));
  jand g00886(.dina(n1087), .dinb(n1081), .dout(n1088));
  jxor g00887(.dina(n935), .dinb(n221), .dout(n1089));
  jor  g00888(.dina(n1089), .dinb(n1008), .dout(n1090));
  jxor g00889(.dina(n1090), .dinb(n989), .dout(n1091));
  jand g00890(.dina(n1091), .dinb(n1088), .dout(n1092));
  jand g00891(.dina(n1008), .dinb(n981), .dout(n1093));
  jand g00892(.dina(n982), .dinb(asqrt[63] ), .dout(n1094));
  jand g00893(.dina(n1094), .dinb(n992), .dout(n1095));
  jnot g00894(.din(n1095), .dout(n1096));
  jor  g00895(.dina(n1096), .dinb(n1093), .dout(n1097));
  jnot g00896(.din(n1097), .dout(n1098));
  jor  g00897(.dina(n1091), .dinb(n1088), .dout(n1099));
  jand g00898(.dina(asqrt[53] ), .dinb(n1004), .dout(n1100));
  jor  g00899(.dina(n1100), .dinb(n1028), .dout(n1101));
  jor  g00900(.dina(n1101), .dinb(n1099), .dout(n1102));
  jand g00901(.dina(n1102), .dinb(n218), .dout(n1103));
  jand g00902(.dina(n1008), .dinb(n864), .dout(n1104));
  jor  g00903(.dina(n1104), .dinb(n1103), .dout(n1105));
  jor  g00904(.dina(n1105), .dinb(n1098), .dout(n1106));
  jor  g00905(.dina(n1106), .dinb(n1092), .dout(asqrt[52] ));
  jnot g00906(.din(a[102] ), .dout(n1108));
  jnot g00907(.din(a[103] ), .dout(n1109));
  jand g00908(.dina(n1109), .dinb(n1108), .dout(n1110));
  jand g00909(.dina(n1110), .dinb(n1010), .dout(n1111));
  jand g00910(.dina(asqrt[52] ), .dinb(a[104] ), .dout(n1112));
  jor  g00911(.dina(n1112), .dinb(n1111), .dout(n1113));
  jand g00912(.dina(n1113), .dinb(asqrt[53] ), .dout(n1114));
  jor  g00913(.dina(n1113), .dinb(asqrt[53] ), .dout(n1115));
  jand g00914(.dina(asqrt[52] ), .dinb(n1010), .dout(n1116));
  jor  g00915(.dina(n1116), .dinb(n1011), .dout(n1117));
  jnot g00916(.din(n1012), .dout(n1118));
  jnot g00917(.din(n1092), .dout(n1119));
  jnot g00918(.din(n1081), .dout(n1120));
  jnot g00919(.din(n1074), .dout(n1121));
  jnot g00920(.din(n1066), .dout(n1122));
  jnot g00921(.din(n1058), .dout(n1123));
  jnot g00922(.din(n1050), .dout(n1124));
  jnot g00923(.din(n1043), .dout(n1125));
  jnot g00924(.din(n1036), .dout(n1126));
  jnot g00925(.din(n1024), .dout(n1127));
  jnot g00926(.din(n1016), .dout(n1128));
  jand g00927(.dina(asqrt[53] ), .dinb(a[106] ), .dout(n1129));
  jor  g00928(.dina(n1013), .dinb(n1129), .dout(n1130));
  jor  g00929(.dina(n1130), .dinb(asqrt[54] ), .dout(n1131));
  jand g00930(.dina(asqrt[53] ), .dinb(n865), .dout(n1132));
  jor  g00931(.dina(n1132), .dinb(n866), .dout(n1133));
  jand g00932(.dina(n1027), .dinb(n1133), .dout(n1134));
  jand g00933(.dina(n1134), .dinb(n1131), .dout(n1135));
  jor  g00934(.dina(n1135), .dinb(n1128), .dout(n1136));
  jor  g00935(.dina(n1136), .dinb(asqrt[55] ), .dout(n1137));
  jnot g00936(.din(n1033), .dout(n1138));
  jand g00937(.dina(n1138), .dinb(n1137), .dout(n1139));
  jor  g00938(.dina(n1139), .dinb(n1127), .dout(n1140));
  jor  g00939(.dina(n1140), .dinb(asqrt[56] ), .dout(n1141));
  jnot g00940(.din(n1040), .dout(n1142));
  jand g00941(.dina(n1142), .dinb(n1141), .dout(n1143));
  jor  g00942(.dina(n1143), .dinb(n1126), .dout(n1144));
  jor  g00943(.dina(n1144), .dinb(asqrt[57] ), .dout(n1145));
  jnot g00944(.din(n1047), .dout(n1146));
  jand g00945(.dina(n1146), .dinb(n1145), .dout(n1147));
  jor  g00946(.dina(n1147), .dinb(n1125), .dout(n1148));
  jor  g00947(.dina(n1148), .dinb(asqrt[58] ), .dout(n1149));
  jand g00948(.dina(n1054), .dinb(n1149), .dout(n1150));
  jor  g00949(.dina(n1150), .dinb(n1124), .dout(n1151));
  jor  g00950(.dina(n1151), .dinb(asqrt[59] ), .dout(n1152));
  jand g00951(.dina(n1062), .dinb(n1152), .dout(n1153));
  jor  g00952(.dina(n1153), .dinb(n1123), .dout(n1154));
  jor  g00953(.dina(n1154), .dinb(asqrt[60] ), .dout(n1155));
  jand g00954(.dina(n1070), .dinb(n1155), .dout(n1156));
  jor  g00955(.dina(n1156), .dinb(n1122), .dout(n1157));
  jor  g00956(.dina(n1157), .dinb(asqrt[61] ), .dout(n1158));
  jnot g00957(.din(n1078), .dout(n1159));
  jand g00958(.dina(n1159), .dinb(n1158), .dout(n1160));
  jor  g00959(.dina(n1160), .dinb(n1121), .dout(n1161));
  jor  g00960(.dina(n1161), .dinb(asqrt[62] ), .dout(n1162));
  jand g00961(.dina(n1085), .dinb(n1162), .dout(n1163));
  jor  g00962(.dina(n1163), .dinb(n1120), .dout(n1164));
  jnot g00963(.din(n1091), .dout(n1165));
  jand g00964(.dina(n1165), .dinb(n1164), .dout(n1166));
  jnot g00965(.din(n1101), .dout(n1167));
  jand g00966(.dina(n1167), .dinb(n1166), .dout(n1168));
  jor  g00967(.dina(n1168), .dinb(asqrt[63] ), .dout(n1169));
  jnot g00968(.din(n1104), .dout(n1170));
  jand g00969(.dina(n1170), .dinb(n1169), .dout(n1171));
  jand g00970(.dina(n1171), .dinb(n1097), .dout(n1172));
  jand g00971(.dina(n1172), .dinb(n1119), .dout(n1173));
  jor  g00972(.dina(n1173), .dinb(n1118), .dout(n1174));
  jand g00973(.dina(n1174), .dinb(n1117), .dout(n1175));
  jand g00974(.dina(n1175), .dinb(n1115), .dout(n1176));
  jor  g00975(.dina(n1176), .dinb(n1114), .dout(n1177));
  jand g00976(.dina(n1177), .dinb(asqrt[54] ), .dout(n1178));
  jor  g00977(.dina(n1177), .dinb(asqrt[54] ), .dout(n1179));
  jand g00978(.dina(asqrt[52] ), .dinb(n1012), .dout(n1180));
  jand g00979(.dina(n1119), .dinb(asqrt[53] ), .dout(n1181));
  jand g00980(.dina(n1181), .dinb(n1096), .dout(n1182));
  jand g00981(.dina(n1182), .dinb(n1169), .dout(n1183));
  jor  g00982(.dina(n1183), .dinb(n1180), .dout(n1184));
  jxor g00983(.dina(n1184), .dinb(a[106] ), .dout(n1185));
  jnot g00984(.din(n1185), .dout(n1186));
  jand g00985(.dina(n1186), .dinb(n1179), .dout(n1187));
  jor  g00986(.dina(n1187), .dinb(n1178), .dout(n1188));
  jand g00987(.dina(n1188), .dinb(asqrt[55] ), .dout(n1189));
  jor  g00988(.dina(n1188), .dinb(asqrt[55] ), .dout(n1190));
  jxor g00989(.dina(n1015), .dinb(n884), .dout(n1191));
  jand g00990(.dina(n1191), .dinb(asqrt[52] ), .dout(n1192));
  jxor g00991(.dina(n1192), .dinb(n1134), .dout(n1193));
  jand g00992(.dina(n1193), .dinb(n1190), .dout(n1194));
  jor  g00993(.dina(n1194), .dinb(n1189), .dout(n1195));
  jand g00994(.dina(n1195), .dinb(asqrt[56] ), .dout(n1196));
  jor  g00995(.dina(n1195), .dinb(asqrt[56] ), .dout(n1197));
  jxor g00996(.dina(n1023), .dinb(n743), .dout(n1198));
  jand g00997(.dina(n1198), .dinb(asqrt[52] ), .dout(n1199));
  jxor g00998(.dina(n1199), .dinb(n1033), .dout(n1200));
  jnot g00999(.din(n1200), .dout(n1201));
  jand g01000(.dina(n1201), .dinb(n1197), .dout(n1202));
  jor  g01001(.dina(n1202), .dinb(n1196), .dout(n1203));
  jand g01002(.dina(n1203), .dinb(asqrt[57] ), .dout(n1204));
  jor  g01003(.dina(n1203), .dinb(asqrt[57] ), .dout(n1205));
  jxor g01004(.dina(n1035), .dinb(n635), .dout(n1206));
  jand g01005(.dina(n1206), .dinb(asqrt[52] ), .dout(n1207));
  jxor g01006(.dina(n1207), .dinb(n1040), .dout(n1208));
  jnot g01007(.din(n1208), .dout(n1209));
  jand g01008(.dina(n1209), .dinb(n1205), .dout(n1210));
  jor  g01009(.dina(n1210), .dinb(n1204), .dout(n1211));
  jand g01010(.dina(n1211), .dinb(asqrt[58] ), .dout(n1212));
  jor  g01011(.dina(n1211), .dinb(asqrt[58] ), .dout(n1213));
  jxor g01012(.dina(n1042), .dinb(n515), .dout(n1214));
  jand g01013(.dina(n1214), .dinb(asqrt[52] ), .dout(n1215));
  jxor g01014(.dina(n1215), .dinb(n1047), .dout(n1216));
  jnot g01015(.din(n1216), .dout(n1217));
  jand g01016(.dina(n1217), .dinb(n1213), .dout(n1218));
  jor  g01017(.dina(n1218), .dinb(n1212), .dout(n1219));
  jand g01018(.dina(n1219), .dinb(asqrt[59] ), .dout(n1220));
  jor  g01019(.dina(n1219), .dinb(asqrt[59] ), .dout(n1221));
  jxor g01020(.dina(n1049), .dinb(n443), .dout(n1222));
  jand g01021(.dina(n1222), .dinb(asqrt[52] ), .dout(n1223));
  jxor g01022(.dina(n1223), .dinb(n1054), .dout(n1224));
  jand g01023(.dina(n1224), .dinb(n1221), .dout(n1225));
  jor  g01024(.dina(n1225), .dinb(n1220), .dout(n1226));
  jand g01025(.dina(n1226), .dinb(asqrt[60] ), .dout(n1227));
  jor  g01026(.dina(n1226), .dinb(asqrt[60] ), .dout(n1228));
  jxor g01027(.dina(n1057), .dinb(n352), .dout(n1229));
  jand g01028(.dina(n1229), .dinb(asqrt[52] ), .dout(n1230));
  jxor g01029(.dina(n1230), .dinb(n1062), .dout(n1231));
  jand g01030(.dina(n1231), .dinb(n1228), .dout(n1232));
  jor  g01031(.dina(n1232), .dinb(n1227), .dout(n1233));
  jand g01032(.dina(n1233), .dinb(asqrt[61] ), .dout(n1234));
  jor  g01033(.dina(n1233), .dinb(asqrt[61] ), .dout(n1235));
  jxor g01034(.dina(n1065), .dinb(n294), .dout(n1236));
  jand g01035(.dina(n1236), .dinb(asqrt[52] ), .dout(n1237));
  jxor g01036(.dina(n1237), .dinb(n1070), .dout(n1238));
  jand g01037(.dina(n1238), .dinb(n1235), .dout(n1239));
  jor  g01038(.dina(n1239), .dinb(n1234), .dout(n1240));
  jand g01039(.dina(n1240), .dinb(asqrt[62] ), .dout(n1241));
  jor  g01040(.dina(n1240), .dinb(asqrt[62] ), .dout(n1242));
  jxor g01041(.dina(n1073), .dinb(n239), .dout(n1243));
  jand g01042(.dina(n1243), .dinb(asqrt[52] ), .dout(n1244));
  jxor g01043(.dina(n1244), .dinb(n1078), .dout(n1245));
  jnot g01044(.din(n1245), .dout(n1246));
  jand g01045(.dina(n1246), .dinb(n1242), .dout(n1247));
  jor  g01046(.dina(n1247), .dinb(n1241), .dout(n1248));
  jxor g01047(.dina(n1080), .dinb(n221), .dout(n1249));
  jand g01048(.dina(n1249), .dinb(asqrt[52] ), .dout(n1250));
  jxor g01049(.dina(n1250), .dinb(n1086), .dout(n1251));
  jnot g01050(.din(n1251), .dout(n1252));
  jor  g01051(.dina(n1252), .dinb(n1248), .dout(n1253));
  jnot g01052(.din(n1253), .dout(n1254));
  jnot g01053(.din(n1241), .dout(n1256));
  jnot g01054(.din(n1234), .dout(n1257));
  jnot g01055(.din(n1227), .dout(n1258));
  jnot g01056(.din(n1220), .dout(n1259));
  jnot g01057(.din(n1212), .dout(n1260));
  jnot g01058(.din(n1204), .dout(n1261));
  jnot g01059(.din(n1196), .dout(n1262));
  jnot g01060(.din(n1189), .dout(n1263));
  jnot g01061(.din(n1178), .dout(n1264));
  jnot g01062(.din(n1114), .dout(n1265));
  jnot g01063(.din(n1111), .dout(n1266));
  jor  g01064(.dina(n1173), .dinb(n1010), .dout(n1267));
  jand g01065(.dina(n1267), .dinb(n1266), .dout(n1268));
  jand g01066(.dina(n1268), .dinb(n1008), .dout(n1269));
  jor  g01067(.dina(n1173), .dinb(a[104] ), .dout(n1270));
  jand g01068(.dina(n1270), .dinb(a[105] ), .dout(n1271));
  jor  g01069(.dina(n1180), .dinb(n1271), .dout(n1272));
  jor  g01070(.dina(n1272), .dinb(n1269), .dout(n1273));
  jand g01071(.dina(n1273), .dinb(n1265), .dout(n1274));
  jand g01072(.dina(n1274), .dinb(n884), .dout(n1275));
  jor  g01073(.dina(n1185), .dinb(n1275), .dout(n1276));
  jand g01074(.dina(n1276), .dinb(n1264), .dout(n1277));
  jand g01075(.dina(n1277), .dinb(n743), .dout(n1278));
  jnot g01076(.din(n1193), .dout(n1279));
  jor  g01077(.dina(n1279), .dinb(n1278), .dout(n1280));
  jand g01078(.dina(n1280), .dinb(n1263), .dout(n1281));
  jand g01079(.dina(n1281), .dinb(n635), .dout(n1282));
  jor  g01080(.dina(n1200), .dinb(n1282), .dout(n1283));
  jand g01081(.dina(n1283), .dinb(n1262), .dout(n1284));
  jand g01082(.dina(n1284), .dinb(n515), .dout(n1285));
  jor  g01083(.dina(n1208), .dinb(n1285), .dout(n1286));
  jand g01084(.dina(n1286), .dinb(n1261), .dout(n1287));
  jand g01085(.dina(n1287), .dinb(n443), .dout(n1288));
  jor  g01086(.dina(n1216), .dinb(n1288), .dout(n1289));
  jand g01087(.dina(n1289), .dinb(n1260), .dout(n1290));
  jand g01088(.dina(n1290), .dinb(n352), .dout(n1291));
  jnot g01089(.din(n1224), .dout(n1292));
  jor  g01090(.dina(n1292), .dinb(n1291), .dout(n1293));
  jand g01091(.dina(n1293), .dinb(n1259), .dout(n1294));
  jand g01092(.dina(n1294), .dinb(n294), .dout(n1295));
  jnot g01093(.din(n1231), .dout(n1296));
  jor  g01094(.dina(n1296), .dinb(n1295), .dout(n1297));
  jand g01095(.dina(n1297), .dinb(n1258), .dout(n1298));
  jand g01096(.dina(n1298), .dinb(n239), .dout(n1299));
  jnot g01097(.din(n1238), .dout(n1300));
  jor  g01098(.dina(n1300), .dinb(n1299), .dout(n1301));
  jand g01099(.dina(n1301), .dinb(n1257), .dout(n1302));
  jand g01100(.dina(n1302), .dinb(n221), .dout(n1303));
  jor  g01101(.dina(n1245), .dinb(n1303), .dout(n1304));
  jand g01102(.dina(n1304), .dinb(n1256), .dout(n1305));
  jor  g01103(.dina(n1251), .dinb(n1305), .dout(n1306));
  jxor g01104(.dina(n1091), .dinb(n1088), .dout(n1307));
  jnot g01105(.din(n1307), .dout(n1308));
  jand g01106(.dina(n1308), .dinb(asqrt[52] ), .dout(n1309));
  jor  g01107(.dina(n1309), .dinb(n1306), .dout(n1310));
  jand g01108(.dina(n1310), .dinb(n218), .dout(n1311));
  jand g01109(.dina(n1172), .dinb(n1088), .dout(n1312));
  jnot g01110(.din(n1312), .dout(n1313));
  jand g01111(.dina(n1307), .dinb(asqrt[63] ), .dout(n1314));
  jand g01112(.dina(n1314), .dinb(n1313), .dout(n1315));
  jor  g01113(.dina(n1315), .dinb(n1311), .dout(n1316));
  jor  g01114(.dina(n1316), .dinb(n1254), .dout(asqrt[51] ));
  jnot g01115(.din(a[100] ), .dout(n1319));
  jnot g01116(.din(a[101] ), .dout(n1320));
  jand g01117(.dina(n1320), .dinb(n1319), .dout(n1321));
  jand g01118(.dina(n1321), .dinb(n1108), .dout(n1322));
  jnot g01119(.din(n1322), .dout(n1323));
  jand g01120(.dina(n1252), .dinb(n1248), .dout(n1325));
  jnot g01121(.din(n1309), .dout(n1326));
  jand g01122(.dina(n1326), .dinb(n1325), .dout(n1327));
  jor  g01123(.dina(n1327), .dinb(asqrt[63] ), .dout(n1328));
  jnot g01124(.din(n1315), .dout(n1329));
  jand g01125(.dina(n1329), .dinb(n1328), .dout(n1330));
  jand g01126(.dina(n1330), .dinb(n1253), .dout(n1332));
  jor  g01127(.dina(n1332), .dinb(n1108), .dout(n1333));
  jand g01128(.dina(n1333), .dinb(n1323), .dout(n1334));
  jor  g01129(.dina(n1334), .dinb(n1173), .dout(n1335));
  jand g01130(.dina(n1334), .dinb(n1173), .dout(n1336));
  jor  g01131(.dina(n1332), .dinb(a[102] ), .dout(n1337));
  jand g01132(.dina(n1337), .dinb(a[103] ), .dout(n1338));
  jand g01133(.dina(asqrt[51] ), .dinb(n1110), .dout(n1339));
  jor  g01134(.dina(n1339), .dinb(n1338), .dout(n1340));
  jor  g01135(.dina(n1340), .dinb(n1336), .dout(n1341));
  jand g01136(.dina(n1341), .dinb(n1335), .dout(n1342));
  jor  g01137(.dina(n1342), .dinb(n1008), .dout(n1343));
  jand g01138(.dina(n1342), .dinb(n1008), .dout(n1344));
  jnot g01139(.din(n1110), .dout(n1345));
  jor  g01140(.dina(n1332), .dinb(n1345), .dout(n1346));
  jor  g01141(.dina(n1314), .dinb(n1254), .dout(n1347));
  jor  g01142(.dina(n1347), .dinb(n1311), .dout(n1348));
  jor  g01143(.dina(n1348), .dinb(n1173), .dout(n1349));
  jand g01144(.dina(n1349), .dinb(n1346), .dout(n1350));
  jxor g01145(.dina(n1350), .dinb(n1010), .dout(n1351));
  jor  g01146(.dina(n1351), .dinb(n1344), .dout(n1352));
  jand g01147(.dina(n1352), .dinb(n1343), .dout(n1353));
  jor  g01148(.dina(n1353), .dinb(n884), .dout(n1354));
  jand g01149(.dina(n1353), .dinb(n884), .dout(n1355));
  jxor g01150(.dina(n1113), .dinb(n1008), .dout(n1356));
  jor  g01151(.dina(n1356), .dinb(n1332), .dout(n1357));
  jxor g01152(.dina(n1357), .dinb(n1175), .dout(n1358));
  jor  g01153(.dina(n1358), .dinb(n1355), .dout(n1359));
  jand g01154(.dina(n1359), .dinb(n1354), .dout(n1360));
  jor  g01155(.dina(n1360), .dinb(n743), .dout(n1361));
  jand g01156(.dina(n1360), .dinb(n743), .dout(n1362));
  jxor g01157(.dina(n1177), .dinb(n884), .dout(n1363));
  jor  g01158(.dina(n1363), .dinb(n1332), .dout(n1364));
  jxor g01159(.dina(n1364), .dinb(n1186), .dout(n1365));
  jor  g01160(.dina(n1365), .dinb(n1362), .dout(n1366));
  jand g01161(.dina(n1366), .dinb(n1361), .dout(n1367));
  jor  g01162(.dina(n1367), .dinb(n635), .dout(n1368));
  jand g01163(.dina(n1367), .dinb(n635), .dout(n1369));
  jxor g01164(.dina(n1188), .dinb(n743), .dout(n1370));
  jor  g01165(.dina(n1370), .dinb(n1332), .dout(n1371));
  jxor g01166(.dina(n1371), .dinb(n1279), .dout(n1372));
  jnot g01167(.din(n1372), .dout(n1373));
  jor  g01168(.dina(n1373), .dinb(n1369), .dout(n1374));
  jand g01169(.dina(n1374), .dinb(n1368), .dout(n1375));
  jor  g01170(.dina(n1375), .dinb(n515), .dout(n1376));
  jand g01171(.dina(n1375), .dinb(n515), .dout(n1377));
  jxor g01172(.dina(n1195), .dinb(n635), .dout(n1378));
  jor  g01173(.dina(n1378), .dinb(n1332), .dout(n1379));
  jxor g01174(.dina(n1379), .dinb(n1201), .dout(n1380));
  jor  g01175(.dina(n1380), .dinb(n1377), .dout(n1381));
  jand g01176(.dina(n1381), .dinb(n1376), .dout(n1382));
  jor  g01177(.dina(n1382), .dinb(n443), .dout(n1383));
  jand g01178(.dina(n1382), .dinb(n443), .dout(n1384));
  jxor g01179(.dina(n1203), .dinb(n515), .dout(n1385));
  jor  g01180(.dina(n1385), .dinb(n1332), .dout(n1386));
  jxor g01181(.dina(n1386), .dinb(n1209), .dout(n1387));
  jor  g01182(.dina(n1387), .dinb(n1384), .dout(n1388));
  jand g01183(.dina(n1388), .dinb(n1383), .dout(n1389));
  jor  g01184(.dina(n1389), .dinb(n352), .dout(n1390));
  jand g01185(.dina(n1389), .dinb(n352), .dout(n1391));
  jxor g01186(.dina(n1211), .dinb(n443), .dout(n1392));
  jor  g01187(.dina(n1392), .dinb(n1332), .dout(n1393));
  jxor g01188(.dina(n1393), .dinb(n1217), .dout(n1394));
  jor  g01189(.dina(n1394), .dinb(n1391), .dout(n1395));
  jand g01190(.dina(n1395), .dinb(n1390), .dout(n1396));
  jor  g01191(.dina(n1396), .dinb(n294), .dout(n1397));
  jand g01192(.dina(n1396), .dinb(n294), .dout(n1398));
  jxor g01193(.dina(n1219), .dinb(n352), .dout(n1399));
  jor  g01194(.dina(n1399), .dinb(n1332), .dout(n1400));
  jxor g01195(.dina(n1400), .dinb(n1292), .dout(n1401));
  jnot g01196(.din(n1401), .dout(n1402));
  jor  g01197(.dina(n1402), .dinb(n1398), .dout(n1403));
  jand g01198(.dina(n1403), .dinb(n1397), .dout(n1404));
  jor  g01199(.dina(n1404), .dinb(n239), .dout(n1405));
  jand g01200(.dina(n1404), .dinb(n239), .dout(n1406));
  jxor g01201(.dina(n1226), .dinb(n294), .dout(n1407));
  jor  g01202(.dina(n1407), .dinb(n1332), .dout(n1408));
  jxor g01203(.dina(n1408), .dinb(n1296), .dout(n1409));
  jnot g01204(.din(n1409), .dout(n1410));
  jor  g01205(.dina(n1410), .dinb(n1406), .dout(n1411));
  jand g01206(.dina(n1411), .dinb(n1405), .dout(n1412));
  jor  g01207(.dina(n1412), .dinb(n221), .dout(n1413));
  jand g01208(.dina(n1412), .dinb(n221), .dout(n1414));
  jxor g01209(.dina(n1233), .dinb(n239), .dout(n1415));
  jor  g01210(.dina(n1415), .dinb(n1332), .dout(n1416));
  jxor g01211(.dina(n1416), .dinb(n1300), .dout(n1417));
  jnot g01212(.din(n1417), .dout(n1418));
  jor  g01213(.dina(n1418), .dinb(n1414), .dout(n1419));
  jand g01214(.dina(n1419), .dinb(n1413), .dout(n1420));
  jxor g01215(.dina(n1240), .dinb(n221), .dout(n1421));
  jor  g01216(.dina(n1421), .dinb(n1332), .dout(n1422));
  jxor g01217(.dina(n1422), .dinb(n1246), .dout(n1423));
  jand g01218(.dina(n1423), .dinb(n1420), .dout(n1424));
  jand g01219(.dina(n1316), .dinb(n1325), .dout(n1426));
  jor  g01220(.dina(n1423), .dinb(n1420), .dout(n1427));
  jor  g01221(.dina(n1427), .dinb(n1254), .dout(n1428));
  jor  g01222(.dina(n1428), .dinb(n1426), .dout(n1429));
  jand g01223(.dina(n1429), .dinb(n218), .dout(n1430));
  jand g01224(.dina(n1330), .dinb(n1305), .dout(n1431));
  jand g01225(.dina(n1306), .dinb(asqrt[63] ), .dout(n1432));
  jand g01226(.dina(n1432), .dinb(n1253), .dout(n1433));
  jnot g01227(.din(n1433), .dout(n1434));
  jor  g01228(.dina(n1434), .dinb(n1431), .dout(n1435));
  jnot g01229(.din(n1435), .dout(n1436));
  jor  g01230(.dina(n1436), .dinb(n1430), .dout(n1437));
  jor  g01231(.dina(n1437), .dinb(n1424), .dout(asqrt[50] ));
  jnot g01232(.din(a[98] ), .dout(n1440));
  jnot g01233(.din(a[99] ), .dout(n1441));
  jand g01234(.dina(n1441), .dinb(n1440), .dout(n1442));
  jand g01235(.dina(n1442), .dinb(n1319), .dout(n1443));
  jand g01236(.dina(asqrt[50] ), .dinb(a[100] ), .dout(n1444));
  jor  g01237(.dina(n1444), .dinb(n1443), .dout(n1445));
  jand g01238(.dina(n1445), .dinb(asqrt[51] ), .dout(n1446));
  jor  g01239(.dina(n1445), .dinb(asqrt[51] ), .dout(n1447));
  jand g01240(.dina(asqrt[50] ), .dinb(n1319), .dout(n1448));
  jor  g01241(.dina(n1448), .dinb(n1320), .dout(n1449));
  jnot g01242(.din(n1321), .dout(n1450));
  jnot g01243(.din(n1424), .dout(n1451));
  jnot g01244(.din(n1426), .dout(n1453));
  jnot g01245(.din(n1413), .dout(n1454));
  jnot g01246(.din(n1405), .dout(n1455));
  jnot g01247(.din(n1397), .dout(n1456));
  jnot g01248(.din(n1390), .dout(n1457));
  jnot g01249(.din(n1383), .dout(n1458));
  jnot g01250(.din(n1376), .dout(n1459));
  jnot g01251(.din(n1368), .dout(n1460));
  jnot g01252(.din(n1361), .dout(n1461));
  jnot g01253(.din(n1354), .dout(n1462));
  jnot g01254(.din(n1343), .dout(n1463));
  jnot g01255(.din(n1335), .dout(n1464));
  jand g01256(.dina(asqrt[51] ), .dinb(a[102] ), .dout(n1465));
  jor  g01257(.dina(n1465), .dinb(n1322), .dout(n1466));
  jor  g01258(.dina(n1466), .dinb(asqrt[52] ), .dout(n1467));
  jand g01259(.dina(asqrt[51] ), .dinb(n1108), .dout(n1468));
  jor  g01260(.dina(n1468), .dinb(n1109), .dout(n1469));
  jand g01261(.dina(n1346), .dinb(n1469), .dout(n1470));
  jand g01262(.dina(n1470), .dinb(n1467), .dout(n1471));
  jor  g01263(.dina(n1471), .dinb(n1464), .dout(n1472));
  jor  g01264(.dina(n1472), .dinb(asqrt[53] ), .dout(n1473));
  jnot g01265(.din(n1351), .dout(n1474));
  jand g01266(.dina(n1474), .dinb(n1473), .dout(n1475));
  jor  g01267(.dina(n1475), .dinb(n1463), .dout(n1476));
  jor  g01268(.dina(n1476), .dinb(asqrt[54] ), .dout(n1477));
  jnot g01269(.din(n1358), .dout(n1478));
  jand g01270(.dina(n1478), .dinb(n1477), .dout(n1479));
  jor  g01271(.dina(n1479), .dinb(n1462), .dout(n1480));
  jor  g01272(.dina(n1480), .dinb(asqrt[55] ), .dout(n1481));
  jnot g01273(.din(n1365), .dout(n1482));
  jand g01274(.dina(n1482), .dinb(n1481), .dout(n1483));
  jor  g01275(.dina(n1483), .dinb(n1461), .dout(n1484));
  jor  g01276(.dina(n1484), .dinb(asqrt[56] ), .dout(n1485));
  jand g01277(.dina(n1372), .dinb(n1485), .dout(n1486));
  jor  g01278(.dina(n1486), .dinb(n1460), .dout(n1487));
  jor  g01279(.dina(n1487), .dinb(asqrt[57] ), .dout(n1488));
  jnot g01280(.din(n1380), .dout(n1489));
  jand g01281(.dina(n1489), .dinb(n1488), .dout(n1490));
  jor  g01282(.dina(n1490), .dinb(n1459), .dout(n1491));
  jor  g01283(.dina(n1491), .dinb(asqrt[58] ), .dout(n1492));
  jnot g01284(.din(n1387), .dout(n1493));
  jand g01285(.dina(n1493), .dinb(n1492), .dout(n1494));
  jor  g01286(.dina(n1494), .dinb(n1458), .dout(n1495));
  jor  g01287(.dina(n1495), .dinb(asqrt[59] ), .dout(n1496));
  jnot g01288(.din(n1394), .dout(n1497));
  jand g01289(.dina(n1497), .dinb(n1496), .dout(n1498));
  jor  g01290(.dina(n1498), .dinb(n1457), .dout(n1499));
  jor  g01291(.dina(n1499), .dinb(asqrt[60] ), .dout(n1500));
  jand g01292(.dina(n1401), .dinb(n1500), .dout(n1501));
  jor  g01293(.dina(n1501), .dinb(n1456), .dout(n1502));
  jor  g01294(.dina(n1502), .dinb(asqrt[61] ), .dout(n1503));
  jand g01295(.dina(n1409), .dinb(n1503), .dout(n1504));
  jor  g01296(.dina(n1504), .dinb(n1455), .dout(n1505));
  jor  g01297(.dina(n1505), .dinb(asqrt[62] ), .dout(n1506));
  jand g01298(.dina(n1417), .dinb(n1506), .dout(n1507));
  jor  g01299(.dina(n1507), .dinb(n1454), .dout(n1508));
  jnot g01300(.din(n1423), .dout(n1509));
  jand g01301(.dina(n1509), .dinb(n1508), .dout(n1510));
  jand g01302(.dina(n1510), .dinb(n1253), .dout(n1511));
  jand g01303(.dina(n1511), .dinb(n1453), .dout(n1512));
  jor  g01304(.dina(n1512), .dinb(asqrt[63] ), .dout(n1513));
  jand g01305(.dina(n1435), .dinb(n1513), .dout(n1514));
  jand g01306(.dina(n1514), .dinb(n1451), .dout(n1516));
  jor  g01307(.dina(n1516), .dinb(n1450), .dout(n1517));
  jand g01308(.dina(n1517), .dinb(n1449), .dout(n1518));
  jand g01309(.dina(n1518), .dinb(n1447), .dout(n1519));
  jor  g01310(.dina(n1519), .dinb(n1446), .dout(n1520));
  jand g01311(.dina(n1520), .dinb(asqrt[52] ), .dout(n1521));
  jor  g01312(.dina(n1520), .dinb(asqrt[52] ), .dout(n1522));
  jand g01313(.dina(asqrt[50] ), .dinb(n1321), .dout(n1523));
  jand g01314(.dina(n1451), .dinb(asqrt[51] ), .dout(n1524));
  jand g01315(.dina(n1524), .dinb(n1434), .dout(n1525));
  jand g01316(.dina(n1525), .dinb(n1513), .dout(n1526));
  jor  g01317(.dina(n1526), .dinb(n1523), .dout(n1527));
  jxor g01318(.dina(n1527), .dinb(a[102] ), .dout(n1528));
  jnot g01319(.din(n1528), .dout(n1529));
  jand g01320(.dina(n1529), .dinb(n1522), .dout(n1530));
  jor  g01321(.dina(n1530), .dinb(n1521), .dout(n1531));
  jand g01322(.dina(n1531), .dinb(asqrt[53] ), .dout(n1532));
  jor  g01323(.dina(n1531), .dinb(asqrt[53] ), .dout(n1533));
  jxor g01324(.dina(n1334), .dinb(n1173), .dout(n1534));
  jand g01325(.dina(n1534), .dinb(asqrt[50] ), .dout(n1535));
  jxor g01326(.dina(n1535), .dinb(n1470), .dout(n1536));
  jand g01327(.dina(n1536), .dinb(n1533), .dout(n1537));
  jor  g01328(.dina(n1537), .dinb(n1532), .dout(n1538));
  jand g01329(.dina(n1538), .dinb(asqrt[54] ), .dout(n1539));
  jor  g01330(.dina(n1538), .dinb(asqrt[54] ), .dout(n1540));
  jxor g01331(.dina(n1342), .dinb(n1008), .dout(n1541));
  jand g01332(.dina(n1541), .dinb(asqrt[50] ), .dout(n1542));
  jxor g01333(.dina(n1542), .dinb(n1351), .dout(n1543));
  jnot g01334(.din(n1543), .dout(n1544));
  jand g01335(.dina(n1544), .dinb(n1540), .dout(n1545));
  jor  g01336(.dina(n1545), .dinb(n1539), .dout(n1546));
  jand g01337(.dina(n1546), .dinb(asqrt[55] ), .dout(n1547));
  jor  g01338(.dina(n1546), .dinb(asqrt[55] ), .dout(n1548));
  jxor g01339(.dina(n1353), .dinb(n884), .dout(n1549));
  jand g01340(.dina(n1549), .dinb(asqrt[50] ), .dout(n1550));
  jxor g01341(.dina(n1550), .dinb(n1358), .dout(n1551));
  jnot g01342(.din(n1551), .dout(n1552));
  jand g01343(.dina(n1552), .dinb(n1548), .dout(n1553));
  jor  g01344(.dina(n1553), .dinb(n1547), .dout(n1554));
  jand g01345(.dina(n1554), .dinb(asqrt[56] ), .dout(n1555));
  jor  g01346(.dina(n1554), .dinb(asqrt[56] ), .dout(n1556));
  jxor g01347(.dina(n1360), .dinb(n743), .dout(n1557));
  jand g01348(.dina(n1557), .dinb(asqrt[50] ), .dout(n1558));
  jxor g01349(.dina(n1558), .dinb(n1365), .dout(n1559));
  jnot g01350(.din(n1559), .dout(n1560));
  jand g01351(.dina(n1560), .dinb(n1556), .dout(n1561));
  jor  g01352(.dina(n1561), .dinb(n1555), .dout(n1562));
  jand g01353(.dina(n1562), .dinb(asqrt[57] ), .dout(n1563));
  jor  g01354(.dina(n1562), .dinb(asqrt[57] ), .dout(n1564));
  jxor g01355(.dina(n1367), .dinb(n635), .dout(n1565));
  jand g01356(.dina(n1565), .dinb(asqrt[50] ), .dout(n1566));
  jxor g01357(.dina(n1566), .dinb(n1372), .dout(n1567));
  jand g01358(.dina(n1567), .dinb(n1564), .dout(n1568));
  jor  g01359(.dina(n1568), .dinb(n1563), .dout(n1569));
  jand g01360(.dina(n1569), .dinb(asqrt[58] ), .dout(n1570));
  jor  g01361(.dina(n1569), .dinb(asqrt[58] ), .dout(n1571));
  jxor g01362(.dina(n1375), .dinb(n515), .dout(n1572));
  jand g01363(.dina(n1572), .dinb(asqrt[50] ), .dout(n1573));
  jxor g01364(.dina(n1573), .dinb(n1380), .dout(n1574));
  jnot g01365(.din(n1574), .dout(n1575));
  jand g01366(.dina(n1575), .dinb(n1571), .dout(n1576));
  jor  g01367(.dina(n1576), .dinb(n1570), .dout(n1577));
  jand g01368(.dina(n1577), .dinb(asqrt[59] ), .dout(n1578));
  jor  g01369(.dina(n1577), .dinb(asqrt[59] ), .dout(n1579));
  jxor g01370(.dina(n1382), .dinb(n443), .dout(n1580));
  jand g01371(.dina(n1580), .dinb(asqrt[50] ), .dout(n1581));
  jxor g01372(.dina(n1581), .dinb(n1387), .dout(n1582));
  jnot g01373(.din(n1582), .dout(n1583));
  jand g01374(.dina(n1583), .dinb(n1579), .dout(n1584));
  jor  g01375(.dina(n1584), .dinb(n1578), .dout(n1585));
  jand g01376(.dina(n1585), .dinb(asqrt[60] ), .dout(n1586));
  jor  g01377(.dina(n1585), .dinb(asqrt[60] ), .dout(n1587));
  jxor g01378(.dina(n1389), .dinb(n352), .dout(n1588));
  jand g01379(.dina(n1588), .dinb(asqrt[50] ), .dout(n1589));
  jxor g01380(.dina(n1589), .dinb(n1394), .dout(n1590));
  jnot g01381(.din(n1590), .dout(n1591));
  jand g01382(.dina(n1591), .dinb(n1587), .dout(n1592));
  jor  g01383(.dina(n1592), .dinb(n1586), .dout(n1593));
  jand g01384(.dina(n1593), .dinb(asqrt[61] ), .dout(n1594));
  jor  g01385(.dina(n1593), .dinb(asqrt[61] ), .dout(n1595));
  jxor g01386(.dina(n1396), .dinb(n294), .dout(n1596));
  jand g01387(.dina(n1596), .dinb(asqrt[50] ), .dout(n1597));
  jxor g01388(.dina(n1597), .dinb(n1401), .dout(n1598));
  jand g01389(.dina(n1598), .dinb(n1595), .dout(n1599));
  jor  g01390(.dina(n1599), .dinb(n1594), .dout(n1600));
  jand g01391(.dina(n1600), .dinb(asqrt[62] ), .dout(n1601));
  jnot g01392(.din(n1601), .dout(n1602));
  jnot g01393(.din(n1594), .dout(n1603));
  jnot g01394(.din(n1586), .dout(n1604));
  jnot g01395(.din(n1578), .dout(n1605));
  jnot g01396(.din(n1570), .dout(n1606));
  jnot g01397(.din(n1563), .dout(n1607));
  jnot g01398(.din(n1555), .dout(n1608));
  jnot g01399(.din(n1547), .dout(n1609));
  jnot g01400(.din(n1539), .dout(n1610));
  jnot g01401(.din(n1532), .dout(n1611));
  jnot g01402(.din(n1521), .dout(n1612));
  jnot g01403(.din(n1446), .dout(n1613));
  jnot g01404(.din(n1443), .dout(n1614));
  jor  g01405(.dina(n1516), .dinb(n1319), .dout(n1615));
  jand g01406(.dina(n1615), .dinb(n1614), .dout(n1616));
  jand g01407(.dina(n1616), .dinb(n1332), .dout(n1617));
  jor  g01408(.dina(n1516), .dinb(a[100] ), .dout(n1618));
  jand g01409(.dina(n1618), .dinb(a[101] ), .dout(n1619));
  jor  g01410(.dina(n1523), .dinb(n1619), .dout(n1620));
  jor  g01411(.dina(n1620), .dinb(n1617), .dout(n1621));
  jand g01412(.dina(n1621), .dinb(n1613), .dout(n1622));
  jand g01413(.dina(n1622), .dinb(n1173), .dout(n1623));
  jor  g01414(.dina(n1528), .dinb(n1623), .dout(n1624));
  jand g01415(.dina(n1624), .dinb(n1612), .dout(n1625));
  jand g01416(.dina(n1625), .dinb(n1008), .dout(n1626));
  jnot g01417(.din(n1536), .dout(n1627));
  jor  g01418(.dina(n1627), .dinb(n1626), .dout(n1628));
  jand g01419(.dina(n1628), .dinb(n1611), .dout(n1629));
  jand g01420(.dina(n1629), .dinb(n884), .dout(n1630));
  jor  g01421(.dina(n1543), .dinb(n1630), .dout(n1631));
  jand g01422(.dina(n1631), .dinb(n1610), .dout(n1632));
  jand g01423(.dina(n1632), .dinb(n743), .dout(n1633));
  jor  g01424(.dina(n1551), .dinb(n1633), .dout(n1634));
  jand g01425(.dina(n1634), .dinb(n1609), .dout(n1635));
  jand g01426(.dina(n1635), .dinb(n635), .dout(n1636));
  jor  g01427(.dina(n1559), .dinb(n1636), .dout(n1637));
  jand g01428(.dina(n1637), .dinb(n1608), .dout(n1638));
  jand g01429(.dina(n1638), .dinb(n515), .dout(n1639));
  jnot g01430(.din(n1567), .dout(n1640));
  jor  g01431(.dina(n1640), .dinb(n1639), .dout(n1641));
  jand g01432(.dina(n1641), .dinb(n1607), .dout(n1642));
  jand g01433(.dina(n1642), .dinb(n443), .dout(n1643));
  jor  g01434(.dina(n1574), .dinb(n1643), .dout(n1644));
  jand g01435(.dina(n1644), .dinb(n1606), .dout(n1645));
  jand g01436(.dina(n1645), .dinb(n352), .dout(n1646));
  jor  g01437(.dina(n1582), .dinb(n1646), .dout(n1647));
  jand g01438(.dina(n1647), .dinb(n1605), .dout(n1648));
  jand g01439(.dina(n1648), .dinb(n294), .dout(n1649));
  jor  g01440(.dina(n1590), .dinb(n1649), .dout(n1650));
  jand g01441(.dina(n1650), .dinb(n1604), .dout(n1651));
  jand g01442(.dina(n1651), .dinb(n239), .dout(n1652));
  jnot g01443(.din(n1598), .dout(n1653));
  jor  g01444(.dina(n1653), .dinb(n1652), .dout(n1654));
  jand g01445(.dina(n1654), .dinb(n1603), .dout(n1655));
  jand g01446(.dina(n1655), .dinb(n221), .dout(n1656));
  jxor g01447(.dina(n1404), .dinb(n239), .dout(n1657));
  jand g01448(.dina(n1657), .dinb(asqrt[50] ), .dout(n1658));
  jxor g01449(.dina(n1658), .dinb(n1409), .dout(n1659));
  jnot g01450(.din(n1659), .dout(n1660));
  jor  g01451(.dina(n1660), .dinb(n1656), .dout(n1661));
  jand g01452(.dina(n1661), .dinb(n1602), .dout(n1662));
  jxor g01453(.dina(n1412), .dinb(n221), .dout(n1663));
  jand g01454(.dina(n1663), .dinb(asqrt[50] ), .dout(n1664));
  jxor g01455(.dina(n1664), .dinb(n1418), .dout(n1665));
  jor  g01456(.dina(n1665), .dinb(n1662), .dout(n1666));
  jxor g01457(.dina(n1423), .dinb(n1420), .dout(n1667));
  jnot g01458(.din(n1667), .dout(n1668));
  jand g01459(.dina(n1668), .dinb(asqrt[50] ), .dout(n1669));
  jor  g01460(.dina(n1669), .dinb(n1666), .dout(n1670));
  jand g01461(.dina(n1670), .dinb(n218), .dout(n1671));
  jand g01462(.dina(n1516), .dinb(n1423), .dout(n1672));
  jand g01463(.dina(n1665), .dinb(n1662), .dout(n1673));
  jor  g01464(.dina(n1673), .dinb(n1672), .dout(n1674));
  jand g01465(.dina(n1514), .dinb(n1420), .dout(n1675));
  jnot g01466(.din(n1675), .dout(n1676));
  jand g01467(.dina(n1667), .dinb(asqrt[63] ), .dout(n1677));
  jand g01468(.dina(n1677), .dinb(n1676), .dout(n1678));
  jor  g01469(.dina(n1678), .dinb(n1674), .dout(n1679));
  jor  g01470(.dina(n1679), .dinb(n1671), .dout(asqrt[49] ));
  jnot g01471(.din(a[96] ), .dout(n1681));
  jnot g01472(.din(a[97] ), .dout(n1682));
  jand g01473(.dina(n1682), .dinb(n1681), .dout(n1683));
  jand g01474(.dina(n1683), .dinb(n1440), .dout(n1684));
  jnot g01475(.din(n1684), .dout(n1685));
  jor  g01476(.dina(n1600), .dinb(asqrt[62] ), .dout(n1686));
  jand g01477(.dina(n1659), .dinb(n1686), .dout(n1687));
  jor  g01478(.dina(n1687), .dinb(n1601), .dout(n1688));
  jnot g01479(.din(n1665), .dout(n1689));
  jand g01480(.dina(n1689), .dinb(n1688), .dout(n1690));
  jnot g01481(.din(n1669), .dout(n1691));
  jand g01482(.dina(n1691), .dinb(n1690), .dout(n1692));
  jor  g01483(.dina(n1692), .dinb(asqrt[63] ), .dout(n1693));
  jnot g01484(.din(n1672), .dout(n1694));
  jor  g01485(.dina(n1689), .dinb(n1688), .dout(n1695));
  jand g01486(.dina(n1695), .dinb(n1694), .dout(n1696));
  jnot g01487(.din(n1678), .dout(n1697));
  jand g01488(.dina(n1697), .dinb(n1696), .dout(n1698));
  jand g01489(.dina(n1698), .dinb(n1693), .dout(n1699));
  jor  g01490(.dina(n1699), .dinb(n1440), .dout(n1700));
  jand g01491(.dina(n1700), .dinb(n1685), .dout(n1701));
  jor  g01492(.dina(n1701), .dinb(n1516), .dout(n1702));
  jand g01493(.dina(n1701), .dinb(n1516), .dout(n1703));
  jor  g01494(.dina(n1699), .dinb(a[98] ), .dout(n1704));
  jand g01495(.dina(n1704), .dinb(a[99] ), .dout(n1705));
  jand g01496(.dina(asqrt[49] ), .dinb(n1442), .dout(n1706));
  jor  g01497(.dina(n1706), .dinb(n1705), .dout(n1707));
  jor  g01498(.dina(n1707), .dinb(n1703), .dout(n1708));
  jand g01499(.dina(n1708), .dinb(n1702), .dout(n1709));
  jor  g01500(.dina(n1709), .dinb(n1332), .dout(n1710));
  jand g01501(.dina(n1709), .dinb(n1332), .dout(n1711));
  jnot g01502(.din(n1442), .dout(n1712));
  jor  g01503(.dina(n1699), .dinb(n1712), .dout(n1713));
  jor  g01504(.dina(n1673), .dinb(n1516), .dout(n1714));
  jor  g01505(.dina(n1714), .dinb(n1671), .dout(n1715));
  jor  g01506(.dina(n1715), .dinb(n1677), .dout(n1716));
  jand g01507(.dina(n1716), .dinb(n1713), .dout(n1717));
  jxor g01508(.dina(n1717), .dinb(n1319), .dout(n1718));
  jor  g01509(.dina(n1718), .dinb(n1711), .dout(n1719));
  jand g01510(.dina(n1719), .dinb(n1710), .dout(n1720));
  jor  g01511(.dina(n1720), .dinb(n1173), .dout(n1721));
  jand g01512(.dina(n1720), .dinb(n1173), .dout(n1722));
  jxor g01513(.dina(n1445), .dinb(n1332), .dout(n1723));
  jor  g01514(.dina(n1723), .dinb(n1699), .dout(n1724));
  jxor g01515(.dina(n1724), .dinb(n1518), .dout(n1725));
  jor  g01516(.dina(n1725), .dinb(n1722), .dout(n1726));
  jand g01517(.dina(n1726), .dinb(n1721), .dout(n1727));
  jor  g01518(.dina(n1727), .dinb(n1008), .dout(n1728));
  jand g01519(.dina(n1727), .dinb(n1008), .dout(n1729));
  jxor g01520(.dina(n1520), .dinb(n1173), .dout(n1730));
  jor  g01521(.dina(n1730), .dinb(n1699), .dout(n1731));
  jxor g01522(.dina(n1731), .dinb(n1528), .dout(n1732));
  jnot g01523(.din(n1732), .dout(n1733));
  jor  g01524(.dina(n1733), .dinb(n1729), .dout(n1734));
  jand g01525(.dina(n1734), .dinb(n1728), .dout(n1735));
  jor  g01526(.dina(n1735), .dinb(n884), .dout(n1736));
  jand g01527(.dina(n1735), .dinb(n884), .dout(n1737));
  jxor g01528(.dina(n1531), .dinb(n1008), .dout(n1738));
  jor  g01529(.dina(n1738), .dinb(n1699), .dout(n1739));
  jxor g01530(.dina(n1739), .dinb(n1627), .dout(n1740));
  jnot g01531(.din(n1740), .dout(n1741));
  jor  g01532(.dina(n1741), .dinb(n1737), .dout(n1742));
  jand g01533(.dina(n1742), .dinb(n1736), .dout(n1743));
  jor  g01534(.dina(n1743), .dinb(n743), .dout(n1744));
  jand g01535(.dina(n1743), .dinb(n743), .dout(n1745));
  jxor g01536(.dina(n1538), .dinb(n884), .dout(n1746));
  jor  g01537(.dina(n1746), .dinb(n1699), .dout(n1747));
  jxor g01538(.dina(n1747), .dinb(n1544), .dout(n1748));
  jor  g01539(.dina(n1748), .dinb(n1745), .dout(n1749));
  jand g01540(.dina(n1749), .dinb(n1744), .dout(n1750));
  jor  g01541(.dina(n1750), .dinb(n635), .dout(n1751));
  jand g01542(.dina(n1750), .dinb(n635), .dout(n1752));
  jxor g01543(.dina(n1546), .dinb(n743), .dout(n1753));
  jor  g01544(.dina(n1753), .dinb(n1699), .dout(n1754));
  jxor g01545(.dina(n1754), .dinb(n1552), .dout(n1755));
  jor  g01546(.dina(n1755), .dinb(n1752), .dout(n1756));
  jand g01547(.dina(n1756), .dinb(n1751), .dout(n1757));
  jor  g01548(.dina(n1757), .dinb(n515), .dout(n1758));
  jand g01549(.dina(n1757), .dinb(n515), .dout(n1759));
  jxor g01550(.dina(n1554), .dinb(n635), .dout(n1760));
  jor  g01551(.dina(n1760), .dinb(n1699), .dout(n1761));
  jxor g01552(.dina(n1761), .dinb(n1560), .dout(n1762));
  jor  g01553(.dina(n1762), .dinb(n1759), .dout(n1763));
  jand g01554(.dina(n1763), .dinb(n1758), .dout(n1764));
  jor  g01555(.dina(n1764), .dinb(n443), .dout(n1765));
  jand g01556(.dina(n1764), .dinb(n443), .dout(n1766));
  jxor g01557(.dina(n1562), .dinb(n515), .dout(n1767));
  jor  g01558(.dina(n1767), .dinb(n1699), .dout(n1768));
  jxor g01559(.dina(n1768), .dinb(n1640), .dout(n1769));
  jnot g01560(.din(n1769), .dout(n1770));
  jor  g01561(.dina(n1770), .dinb(n1766), .dout(n1771));
  jand g01562(.dina(n1771), .dinb(n1765), .dout(n1772));
  jor  g01563(.dina(n1772), .dinb(n352), .dout(n1773));
  jand g01564(.dina(n1772), .dinb(n352), .dout(n1774));
  jxor g01565(.dina(n1569), .dinb(n443), .dout(n1775));
  jor  g01566(.dina(n1775), .dinb(n1699), .dout(n1776));
  jxor g01567(.dina(n1776), .dinb(n1575), .dout(n1777));
  jor  g01568(.dina(n1777), .dinb(n1774), .dout(n1778));
  jand g01569(.dina(n1778), .dinb(n1773), .dout(n1779));
  jor  g01570(.dina(n1779), .dinb(n294), .dout(n1780));
  jand g01571(.dina(n1779), .dinb(n294), .dout(n1781));
  jxor g01572(.dina(n1577), .dinb(n352), .dout(n1782));
  jor  g01573(.dina(n1782), .dinb(n1699), .dout(n1783));
  jxor g01574(.dina(n1783), .dinb(n1583), .dout(n1784));
  jor  g01575(.dina(n1784), .dinb(n1781), .dout(n1785));
  jand g01576(.dina(n1785), .dinb(n1780), .dout(n1786));
  jor  g01577(.dina(n1786), .dinb(n239), .dout(n1787));
  jand g01578(.dina(n1786), .dinb(n239), .dout(n1788));
  jxor g01579(.dina(n1585), .dinb(n294), .dout(n1789));
  jor  g01580(.dina(n1789), .dinb(n1699), .dout(n1790));
  jxor g01581(.dina(n1790), .dinb(n1591), .dout(n1791));
  jor  g01582(.dina(n1791), .dinb(n1788), .dout(n1792));
  jand g01583(.dina(n1792), .dinb(n1787), .dout(n1793));
  jor  g01584(.dina(n1793), .dinb(n221), .dout(n1794));
  jand g01585(.dina(n1793), .dinb(n221), .dout(n1795));
  jxor g01586(.dina(n1593), .dinb(n239), .dout(n1796));
  jor  g01587(.dina(n1796), .dinb(n1699), .dout(n1797));
  jxor g01588(.dina(n1797), .dinb(n1653), .dout(n1798));
  jnot g01589(.din(n1798), .dout(n1799));
  jor  g01590(.dina(n1799), .dinb(n1795), .dout(n1800));
  jand g01591(.dina(n1800), .dinb(n1794), .dout(n1801));
  jxor g01592(.dina(n1600), .dinb(n221), .dout(n1802));
  jor  g01593(.dina(n1802), .dinb(n1699), .dout(n1803));
  jxor g01594(.dina(n1803), .dinb(n1659), .dout(n1804));
  jand g01595(.dina(n1804), .dinb(n1801), .dout(n1805));
  jand g01596(.dina(n1699), .dinb(n1662), .dout(n1806));
  jand g01597(.dina(n1666), .dinb(asqrt[63] ), .dout(n1807));
  jand g01598(.dina(n1807), .dinb(n1695), .dout(n1808));
  jnot g01599(.din(n1808), .dout(n1809));
  jor  g01600(.dina(n1809), .dinb(n1806), .dout(n1810));
  jnot g01601(.din(n1810), .dout(n1811));
  jor  g01602(.dina(n1804), .dinb(n1801), .dout(n1812));
  jand g01603(.dina(asqrt[49] ), .dinb(n1690), .dout(n1813));
  jor  g01604(.dina(n1813), .dinb(n1812), .dout(n1814));
  jor  g01605(.dina(n1814), .dinb(n1673), .dout(n1815));
  jand g01606(.dina(n1815), .dinb(n218), .dout(n1816));
  jand g01607(.dina(n1699), .dinb(n1665), .dout(n1817));
  jor  g01608(.dina(n1817), .dinb(n1816), .dout(n1818));
  jor  g01609(.dina(n1818), .dinb(n1811), .dout(n1819));
  jor  g01610(.dina(n1819), .dinb(n1805), .dout(asqrt[48] ));
  jnot g01611(.din(n1794), .dout(n1821));
  jnot g01612(.din(n1787), .dout(n1822));
  jnot g01613(.din(n1780), .dout(n1823));
  jnot g01614(.din(n1773), .dout(n1824));
  jnot g01615(.din(n1765), .dout(n1825));
  jnot g01616(.din(n1758), .dout(n1826));
  jnot g01617(.din(n1751), .dout(n1827));
  jnot g01618(.din(n1744), .dout(n1828));
  jnot g01619(.din(n1736), .dout(n1829));
  jnot g01620(.din(n1728), .dout(n1830));
  jnot g01621(.din(n1721), .dout(n1831));
  jnot g01622(.din(n1710), .dout(n1832));
  jnot g01623(.din(n1702), .dout(n1833));
  jand g01624(.dina(asqrt[49] ), .dinb(a[98] ), .dout(n1834));
  jor  g01625(.dina(n1834), .dinb(n1684), .dout(n1835));
  jor  g01626(.dina(n1835), .dinb(asqrt[50] ), .dout(n1836));
  jand g01627(.dina(asqrt[49] ), .dinb(n1440), .dout(n1837));
  jor  g01628(.dina(n1837), .dinb(n1441), .dout(n1838));
  jand g01629(.dina(n1713), .dinb(n1838), .dout(n1839));
  jand g01630(.dina(n1839), .dinb(n1836), .dout(n1840));
  jor  g01631(.dina(n1840), .dinb(n1833), .dout(n1841));
  jor  g01632(.dina(n1841), .dinb(asqrt[51] ), .dout(n1842));
  jnot g01633(.din(n1718), .dout(n1843));
  jand g01634(.dina(n1843), .dinb(n1842), .dout(n1844));
  jor  g01635(.dina(n1844), .dinb(n1832), .dout(n1845));
  jor  g01636(.dina(n1845), .dinb(asqrt[52] ), .dout(n1846));
  jnot g01637(.din(n1725), .dout(n1847));
  jand g01638(.dina(n1847), .dinb(n1846), .dout(n1848));
  jor  g01639(.dina(n1848), .dinb(n1831), .dout(n1849));
  jor  g01640(.dina(n1849), .dinb(asqrt[53] ), .dout(n1850));
  jand g01641(.dina(n1732), .dinb(n1850), .dout(n1851));
  jor  g01642(.dina(n1851), .dinb(n1830), .dout(n1852));
  jor  g01643(.dina(n1852), .dinb(asqrt[54] ), .dout(n1853));
  jand g01644(.dina(n1740), .dinb(n1853), .dout(n1854));
  jor  g01645(.dina(n1854), .dinb(n1829), .dout(n1855));
  jor  g01646(.dina(n1855), .dinb(asqrt[55] ), .dout(n1856));
  jnot g01647(.din(n1748), .dout(n1857));
  jand g01648(.dina(n1857), .dinb(n1856), .dout(n1858));
  jor  g01649(.dina(n1858), .dinb(n1828), .dout(n1859));
  jor  g01650(.dina(n1859), .dinb(asqrt[56] ), .dout(n1860));
  jnot g01651(.din(n1755), .dout(n1861));
  jand g01652(.dina(n1861), .dinb(n1860), .dout(n1862));
  jor  g01653(.dina(n1862), .dinb(n1827), .dout(n1863));
  jor  g01654(.dina(n1863), .dinb(asqrt[57] ), .dout(n1864));
  jnot g01655(.din(n1762), .dout(n1865));
  jand g01656(.dina(n1865), .dinb(n1864), .dout(n1866));
  jor  g01657(.dina(n1866), .dinb(n1826), .dout(n1867));
  jor  g01658(.dina(n1867), .dinb(asqrt[58] ), .dout(n1868));
  jand g01659(.dina(n1769), .dinb(n1868), .dout(n1869));
  jor  g01660(.dina(n1869), .dinb(n1825), .dout(n1870));
  jor  g01661(.dina(n1870), .dinb(asqrt[59] ), .dout(n1871));
  jnot g01662(.din(n1777), .dout(n1872));
  jand g01663(.dina(n1872), .dinb(n1871), .dout(n1873));
  jor  g01664(.dina(n1873), .dinb(n1824), .dout(n1874));
  jor  g01665(.dina(n1874), .dinb(asqrt[60] ), .dout(n1875));
  jnot g01666(.din(n1784), .dout(n1876));
  jand g01667(.dina(n1876), .dinb(n1875), .dout(n1877));
  jor  g01668(.dina(n1877), .dinb(n1823), .dout(n1878));
  jor  g01669(.dina(n1878), .dinb(asqrt[61] ), .dout(n1879));
  jnot g01670(.din(n1791), .dout(n1880));
  jand g01671(.dina(n1880), .dinb(n1879), .dout(n1881));
  jor  g01672(.dina(n1881), .dinb(n1822), .dout(n1882));
  jor  g01673(.dina(n1882), .dinb(asqrt[62] ), .dout(n1883));
  jand g01674(.dina(n1798), .dinb(n1883), .dout(n1884));
  jor  g01675(.dina(n1884), .dinb(n1821), .dout(n1885));
  jnot g01676(.din(n1804), .dout(n1886));
  jand g01677(.dina(n1886), .dinb(n1885), .dout(n1887));
  jand g01678(.dina(n1819), .dinb(n1887), .dout(n1888));
  jxor g01679(.dina(n1793), .dinb(n221), .dout(n1889));
  jand g01680(.dina(n1889), .dinb(asqrt[48] ), .dout(n1890));
  jxor g01681(.dina(n1890), .dinb(n1798), .dout(n1891));
  jnot g01682(.din(n1891), .dout(n1892));
  jand g01683(.dina(asqrt[48] ), .dinb(a[96] ), .dout(n1893));
  jnot g01684(.din(a[94] ), .dout(n1894));
  jnot g01685(.din(a[95] ), .dout(n1895));
  jand g01686(.dina(n1895), .dinb(n1894), .dout(n1896));
  jand g01687(.dina(n1896), .dinb(n1681), .dout(n1897));
  jor  g01688(.dina(n1897), .dinb(n1893), .dout(n1898));
  jand g01689(.dina(n1898), .dinb(asqrt[49] ), .dout(n1899));
  jor  g01690(.dina(n1898), .dinb(asqrt[49] ), .dout(n1900));
  jand g01691(.dina(asqrt[48] ), .dinb(n1681), .dout(n1901));
  jor  g01692(.dina(n1901), .dinb(n1682), .dout(n1902));
  jnot g01693(.din(n1683), .dout(n1903));
  jnot g01694(.din(n1805), .dout(n1904));
  jnot g01695(.din(n1813), .dout(n1905));
  jand g01696(.dina(n1905), .dinb(n1887), .dout(n1906));
  jand g01697(.dina(n1906), .dinb(n1695), .dout(n1907));
  jor  g01698(.dina(n1907), .dinb(asqrt[63] ), .dout(n1908));
  jnot g01699(.din(n1817), .dout(n1909));
  jand g01700(.dina(n1909), .dinb(n1908), .dout(n1910));
  jand g01701(.dina(n1910), .dinb(n1810), .dout(n1911));
  jand g01702(.dina(n1911), .dinb(n1904), .dout(n1912));
  jor  g01703(.dina(n1912), .dinb(n1903), .dout(n1913));
  jand g01704(.dina(n1913), .dinb(n1902), .dout(n1914));
  jand g01705(.dina(n1914), .dinb(n1900), .dout(n1915));
  jor  g01706(.dina(n1915), .dinb(n1899), .dout(n1916));
  jand g01707(.dina(n1916), .dinb(asqrt[50] ), .dout(n1917));
  jor  g01708(.dina(n1916), .dinb(asqrt[50] ), .dout(n1918));
  jand g01709(.dina(asqrt[48] ), .dinb(n1683), .dout(n1919));
  jand g01710(.dina(n1904), .dinb(asqrt[49] ), .dout(n1920));
  jand g01711(.dina(n1920), .dinb(n1809), .dout(n1921));
  jand g01712(.dina(n1921), .dinb(n1908), .dout(n1922));
  jor  g01713(.dina(n1922), .dinb(n1919), .dout(n1923));
  jxor g01714(.dina(n1923), .dinb(a[98] ), .dout(n1924));
  jnot g01715(.din(n1924), .dout(n1925));
  jand g01716(.dina(n1925), .dinb(n1918), .dout(n1926));
  jor  g01717(.dina(n1926), .dinb(n1917), .dout(n1927));
  jand g01718(.dina(n1927), .dinb(asqrt[51] ), .dout(n1928));
  jor  g01719(.dina(n1927), .dinb(asqrt[51] ), .dout(n1929));
  jxor g01720(.dina(n1701), .dinb(n1516), .dout(n1930));
  jand g01721(.dina(n1930), .dinb(asqrt[48] ), .dout(n1931));
  jxor g01722(.dina(n1931), .dinb(n1839), .dout(n1932));
  jand g01723(.dina(n1932), .dinb(n1929), .dout(n1933));
  jor  g01724(.dina(n1933), .dinb(n1928), .dout(n1934));
  jand g01725(.dina(n1934), .dinb(asqrt[52] ), .dout(n1935));
  jor  g01726(.dina(n1934), .dinb(asqrt[52] ), .dout(n1936));
  jxor g01727(.dina(n1709), .dinb(n1332), .dout(n1937));
  jand g01728(.dina(n1937), .dinb(asqrt[48] ), .dout(n1938));
  jxor g01729(.dina(n1938), .dinb(n1718), .dout(n1939));
  jnot g01730(.din(n1939), .dout(n1940));
  jand g01731(.dina(n1940), .dinb(n1936), .dout(n1941));
  jor  g01732(.dina(n1941), .dinb(n1935), .dout(n1942));
  jand g01733(.dina(n1942), .dinb(asqrt[53] ), .dout(n1943));
  jor  g01734(.dina(n1942), .dinb(asqrt[53] ), .dout(n1944));
  jxor g01735(.dina(n1720), .dinb(n1173), .dout(n1945));
  jand g01736(.dina(n1945), .dinb(asqrt[48] ), .dout(n1946));
  jxor g01737(.dina(n1946), .dinb(n1725), .dout(n1947));
  jnot g01738(.din(n1947), .dout(n1948));
  jand g01739(.dina(n1948), .dinb(n1944), .dout(n1949));
  jor  g01740(.dina(n1949), .dinb(n1943), .dout(n1950));
  jand g01741(.dina(n1950), .dinb(asqrt[54] ), .dout(n1951));
  jor  g01742(.dina(n1950), .dinb(asqrt[54] ), .dout(n1952));
  jxor g01743(.dina(n1727), .dinb(n1008), .dout(n1953));
  jand g01744(.dina(n1953), .dinb(asqrt[48] ), .dout(n1954));
  jxor g01745(.dina(n1954), .dinb(n1732), .dout(n1955));
  jand g01746(.dina(n1955), .dinb(n1952), .dout(n1956));
  jor  g01747(.dina(n1956), .dinb(n1951), .dout(n1957));
  jand g01748(.dina(n1957), .dinb(asqrt[55] ), .dout(n1958));
  jor  g01749(.dina(n1957), .dinb(asqrt[55] ), .dout(n1959));
  jxor g01750(.dina(n1735), .dinb(n884), .dout(n1960));
  jand g01751(.dina(n1960), .dinb(asqrt[48] ), .dout(n1961));
  jxor g01752(.dina(n1961), .dinb(n1740), .dout(n1962));
  jand g01753(.dina(n1962), .dinb(n1959), .dout(n1963));
  jor  g01754(.dina(n1963), .dinb(n1958), .dout(n1964));
  jand g01755(.dina(n1964), .dinb(asqrt[56] ), .dout(n1965));
  jor  g01756(.dina(n1964), .dinb(asqrt[56] ), .dout(n1966));
  jxor g01757(.dina(n1743), .dinb(n743), .dout(n1967));
  jand g01758(.dina(n1967), .dinb(asqrt[48] ), .dout(n1968));
  jxor g01759(.dina(n1968), .dinb(n1748), .dout(n1969));
  jnot g01760(.din(n1969), .dout(n1970));
  jand g01761(.dina(n1970), .dinb(n1966), .dout(n1971));
  jor  g01762(.dina(n1971), .dinb(n1965), .dout(n1972));
  jand g01763(.dina(n1972), .dinb(asqrt[57] ), .dout(n1973));
  jor  g01764(.dina(n1972), .dinb(asqrt[57] ), .dout(n1974));
  jxor g01765(.dina(n1750), .dinb(n635), .dout(n1975));
  jand g01766(.dina(n1975), .dinb(asqrt[48] ), .dout(n1976));
  jxor g01767(.dina(n1976), .dinb(n1755), .dout(n1977));
  jnot g01768(.din(n1977), .dout(n1978));
  jand g01769(.dina(n1978), .dinb(n1974), .dout(n1979));
  jor  g01770(.dina(n1979), .dinb(n1973), .dout(n1980));
  jand g01771(.dina(n1980), .dinb(asqrt[58] ), .dout(n1981));
  jor  g01772(.dina(n1980), .dinb(asqrt[58] ), .dout(n1982));
  jxor g01773(.dina(n1757), .dinb(n515), .dout(n1983));
  jand g01774(.dina(n1983), .dinb(asqrt[48] ), .dout(n1984));
  jxor g01775(.dina(n1984), .dinb(n1762), .dout(n1985));
  jnot g01776(.din(n1985), .dout(n1986));
  jand g01777(.dina(n1986), .dinb(n1982), .dout(n1987));
  jor  g01778(.dina(n1987), .dinb(n1981), .dout(n1988));
  jand g01779(.dina(n1988), .dinb(asqrt[59] ), .dout(n1989));
  jor  g01780(.dina(n1988), .dinb(asqrt[59] ), .dout(n1990));
  jxor g01781(.dina(n1764), .dinb(n443), .dout(n1991));
  jand g01782(.dina(n1991), .dinb(asqrt[48] ), .dout(n1992));
  jxor g01783(.dina(n1992), .dinb(n1769), .dout(n1993));
  jand g01784(.dina(n1993), .dinb(n1990), .dout(n1994));
  jor  g01785(.dina(n1994), .dinb(n1989), .dout(n1995));
  jand g01786(.dina(n1995), .dinb(asqrt[60] ), .dout(n1996));
  jor  g01787(.dina(n1995), .dinb(asqrt[60] ), .dout(n1997));
  jxor g01788(.dina(n1772), .dinb(n352), .dout(n1998));
  jand g01789(.dina(n1998), .dinb(asqrt[48] ), .dout(n1999));
  jxor g01790(.dina(n1999), .dinb(n1777), .dout(n2000));
  jnot g01791(.din(n2000), .dout(n2001));
  jand g01792(.dina(n2001), .dinb(n1997), .dout(n2002));
  jor  g01793(.dina(n2002), .dinb(n1996), .dout(n2003));
  jand g01794(.dina(n2003), .dinb(asqrt[61] ), .dout(n2004));
  jor  g01795(.dina(n2003), .dinb(asqrt[61] ), .dout(n2005));
  jxor g01796(.dina(n1779), .dinb(n294), .dout(n2006));
  jand g01797(.dina(n2006), .dinb(asqrt[48] ), .dout(n2007));
  jxor g01798(.dina(n2007), .dinb(n1784), .dout(n2008));
  jnot g01799(.din(n2008), .dout(n2009));
  jand g01800(.dina(n2009), .dinb(n2005), .dout(n2010));
  jor  g01801(.dina(n2010), .dinb(n2004), .dout(n2011));
  jand g01802(.dina(n2011), .dinb(asqrt[62] ), .dout(n2012));
  jnot g01803(.din(n2012), .dout(n2013));
  jnot g01804(.din(n2004), .dout(n2014));
  jnot g01805(.din(n1996), .dout(n2015));
  jnot g01806(.din(n1989), .dout(n2016));
  jnot g01807(.din(n1981), .dout(n2017));
  jnot g01808(.din(n1973), .dout(n2018));
  jnot g01809(.din(n1965), .dout(n2019));
  jnot g01810(.din(n1958), .dout(n2020));
  jnot g01811(.din(n1951), .dout(n2021));
  jnot g01812(.din(n1943), .dout(n2022));
  jnot g01813(.din(n1935), .dout(n2023));
  jnot g01814(.din(n1928), .dout(n2024));
  jnot g01815(.din(n1917), .dout(n2025));
  jnot g01816(.din(n1899), .dout(n2026));
  jor  g01817(.dina(n1912), .dinb(n1681), .dout(n2027));
  jnot g01818(.din(n1897), .dout(n2028));
  jand g01819(.dina(n2028), .dinb(n2027), .dout(n2029));
  jand g01820(.dina(n2029), .dinb(n1699), .dout(n2030));
  jor  g01821(.dina(n1912), .dinb(a[96] ), .dout(n2031));
  jand g01822(.dina(n2031), .dinb(a[97] ), .dout(n2032));
  jor  g01823(.dina(n1919), .dinb(n2032), .dout(n2033));
  jor  g01824(.dina(n2033), .dinb(n2030), .dout(n2034));
  jand g01825(.dina(n2034), .dinb(n2026), .dout(n2035));
  jand g01826(.dina(n2035), .dinb(n1516), .dout(n2036));
  jor  g01827(.dina(n1924), .dinb(n2036), .dout(n2037));
  jand g01828(.dina(n2037), .dinb(n2025), .dout(n2038));
  jand g01829(.dina(n2038), .dinb(n1332), .dout(n2039));
  jnot g01830(.din(n1932), .dout(n2040));
  jor  g01831(.dina(n2040), .dinb(n2039), .dout(n2041));
  jand g01832(.dina(n2041), .dinb(n2024), .dout(n2042));
  jand g01833(.dina(n2042), .dinb(n1173), .dout(n2043));
  jor  g01834(.dina(n1939), .dinb(n2043), .dout(n2044));
  jand g01835(.dina(n2044), .dinb(n2023), .dout(n2045));
  jand g01836(.dina(n2045), .dinb(n1008), .dout(n2046));
  jor  g01837(.dina(n1947), .dinb(n2046), .dout(n2047));
  jand g01838(.dina(n2047), .dinb(n2022), .dout(n2048));
  jand g01839(.dina(n2048), .dinb(n884), .dout(n2049));
  jnot g01840(.din(n1955), .dout(n2050));
  jor  g01841(.dina(n2050), .dinb(n2049), .dout(n2051));
  jand g01842(.dina(n2051), .dinb(n2021), .dout(n2052));
  jand g01843(.dina(n2052), .dinb(n743), .dout(n2053));
  jnot g01844(.din(n1962), .dout(n2054));
  jor  g01845(.dina(n2054), .dinb(n2053), .dout(n2055));
  jand g01846(.dina(n2055), .dinb(n2020), .dout(n2056));
  jand g01847(.dina(n2056), .dinb(n635), .dout(n2057));
  jor  g01848(.dina(n1969), .dinb(n2057), .dout(n2058));
  jand g01849(.dina(n2058), .dinb(n2019), .dout(n2059));
  jand g01850(.dina(n2059), .dinb(n515), .dout(n2060));
  jor  g01851(.dina(n1977), .dinb(n2060), .dout(n2061));
  jand g01852(.dina(n2061), .dinb(n2018), .dout(n2062));
  jand g01853(.dina(n2062), .dinb(n443), .dout(n2063));
  jor  g01854(.dina(n1985), .dinb(n2063), .dout(n2064));
  jand g01855(.dina(n2064), .dinb(n2017), .dout(n2065));
  jand g01856(.dina(n2065), .dinb(n352), .dout(n2066));
  jnot g01857(.din(n1993), .dout(n2067));
  jor  g01858(.dina(n2067), .dinb(n2066), .dout(n2068));
  jand g01859(.dina(n2068), .dinb(n2016), .dout(n2069));
  jand g01860(.dina(n2069), .dinb(n294), .dout(n2070));
  jor  g01861(.dina(n2000), .dinb(n2070), .dout(n2071));
  jand g01862(.dina(n2071), .dinb(n2015), .dout(n2072));
  jand g01863(.dina(n2072), .dinb(n239), .dout(n2073));
  jor  g01864(.dina(n2008), .dinb(n2073), .dout(n2074));
  jand g01865(.dina(n2074), .dinb(n2014), .dout(n2075));
  jand g01866(.dina(n2075), .dinb(n221), .dout(n2076));
  jxor g01867(.dina(n1786), .dinb(n239), .dout(n2077));
  jand g01868(.dina(n2077), .dinb(asqrt[48] ), .dout(n2078));
  jxor g01869(.dina(n2078), .dinb(n1791), .dout(n2079));
  jor  g01870(.dina(n2079), .dinb(n2076), .dout(n2080));
  jand g01871(.dina(n2080), .dinb(n2013), .dout(n2081));
  jor  g01872(.dina(n2081), .dinb(n1892), .dout(n2082));
  jor  g01873(.dina(n2082), .dinb(n1805), .dout(n2083));
  jor  g01874(.dina(n2083), .dinb(n1888), .dout(n2084));
  jand g01875(.dina(n2084), .dinb(n218), .dout(n2085));
  jand g01876(.dina(n1912), .dinb(n1804), .dout(n2086));
  jnot g01877(.din(n2086), .dout(n2087));
  jor  g01878(.dina(n2011), .dinb(asqrt[62] ), .dout(n2088));
  jnot g01879(.din(n2079), .dout(n2089));
  jand g01880(.dina(n2089), .dinb(n2088), .dout(n2090));
  jor  g01881(.dina(n2090), .dinb(n2012), .dout(n2091));
  jor  g01882(.dina(n2091), .dinb(n1891), .dout(n2092));
  jand g01883(.dina(n2092), .dinb(n2087), .dout(n2093));
  jand g01884(.dina(n1911), .dinb(n1801), .dout(n2094));
  jnot g01885(.din(n2094), .dout(n2095));
  jand g01886(.dina(n1812), .dinb(asqrt[63] ), .dout(n2096));
  jand g01887(.dina(n2096), .dinb(n1904), .dout(n2097));
  jand g01888(.dina(n2097), .dinb(n2095), .dout(n2098));
  jnot g01889(.din(n2098), .dout(n2099));
  jand g01890(.dina(n2099), .dinb(n2093), .dout(n2100));
  jnot g01891(.din(n2100), .dout(n2101));
  jor  g01892(.dina(n2101), .dinb(n2085), .dout(asqrt[47] ));
  jnot g01893(.din(n1888), .dout(n2103));
  jand g01894(.dina(n2091), .dinb(n1891), .dout(n2104));
  jand g01895(.dina(n2104), .dinb(n1904), .dout(n2105));
  jand g01896(.dina(n2105), .dinb(n2103), .dout(n2106));
  jor  g01897(.dina(n2106), .dinb(asqrt[63] ), .dout(n2107));
  jand g01898(.dina(n2100), .dinb(n2107), .dout(n2108));
  jor  g01899(.dina(n2108), .dinb(n1894), .dout(n2109));
  jnot g01900(.din(a[92] ), .dout(n2110));
  jnot g01901(.din(a[93] ), .dout(n2111));
  jand g01902(.dina(n2111), .dinb(n2110), .dout(n2112));
  jand g01903(.dina(n2112), .dinb(n1894), .dout(n2113));
  jnot g01904(.din(n2113), .dout(n2114));
  jand g01905(.dina(n2114), .dinb(n2109), .dout(n2115));
  jor  g01906(.dina(n2115), .dinb(n1912), .dout(n2116));
  jand g01907(.dina(n2115), .dinb(n1912), .dout(n2117));
  jor  g01908(.dina(n2108), .dinb(a[94] ), .dout(n2118));
  jand g01909(.dina(n2118), .dinb(a[95] ), .dout(n2119));
  jand g01910(.dina(asqrt[47] ), .dinb(n1896), .dout(n2120));
  jor  g01911(.dina(n2120), .dinb(n2119), .dout(n2121));
  jor  g01912(.dina(n2121), .dinb(n2117), .dout(n2122));
  jand g01913(.dina(n2122), .dinb(n2116), .dout(n2123));
  jor  g01914(.dina(n2123), .dinb(n1699), .dout(n2124));
  jand g01915(.dina(n2123), .dinb(n1699), .dout(n2125));
  jnot g01916(.din(n1896), .dout(n2126));
  jor  g01917(.dina(n2108), .dinb(n2126), .dout(n2127));
  jnot g01918(.din(n2092), .dout(n2128));
  jor  g01919(.dina(n2097), .dinb(n2128), .dout(n2129));
  jor  g01920(.dina(n2129), .dinb(n2085), .dout(n2130));
  jor  g01921(.dina(n2130), .dinb(n1912), .dout(n2131));
  jand g01922(.dina(n2131), .dinb(n2127), .dout(n2132));
  jxor g01923(.dina(n2132), .dinb(n1681), .dout(n2133));
  jor  g01924(.dina(n2133), .dinb(n2125), .dout(n2134));
  jand g01925(.dina(n2134), .dinb(n2124), .dout(n2135));
  jor  g01926(.dina(n2135), .dinb(n1516), .dout(n2136));
  jand g01927(.dina(n2135), .dinb(n1516), .dout(n2137));
  jxor g01928(.dina(n1898), .dinb(n1699), .dout(n2138));
  jor  g01929(.dina(n2138), .dinb(n2108), .dout(n2139));
  jxor g01930(.dina(n2139), .dinb(n2033), .dout(n2140));
  jnot g01931(.din(n2140), .dout(n2141));
  jor  g01932(.dina(n2141), .dinb(n2137), .dout(n2142));
  jand g01933(.dina(n2142), .dinb(n2136), .dout(n2143));
  jor  g01934(.dina(n2143), .dinb(n1332), .dout(n2144));
  jand g01935(.dina(n2143), .dinb(n1332), .dout(n2145));
  jxor g01936(.dina(n1916), .dinb(n1516), .dout(n2146));
  jor  g01937(.dina(n2146), .dinb(n2108), .dout(n2147));
  jxor g01938(.dina(n2147), .dinb(n1925), .dout(n2148));
  jor  g01939(.dina(n2148), .dinb(n2145), .dout(n2149));
  jand g01940(.dina(n2149), .dinb(n2144), .dout(n2150));
  jor  g01941(.dina(n2150), .dinb(n1173), .dout(n2151));
  jand g01942(.dina(n2150), .dinb(n1173), .dout(n2152));
  jxor g01943(.dina(n1927), .dinb(n1332), .dout(n2153));
  jor  g01944(.dina(n2153), .dinb(n2108), .dout(n2154));
  jxor g01945(.dina(n2154), .dinb(n2040), .dout(n2155));
  jnot g01946(.din(n2155), .dout(n2156));
  jor  g01947(.dina(n2156), .dinb(n2152), .dout(n2157));
  jand g01948(.dina(n2157), .dinb(n2151), .dout(n2158));
  jor  g01949(.dina(n2158), .dinb(n1008), .dout(n2159));
  jand g01950(.dina(n2158), .dinb(n1008), .dout(n2160));
  jxor g01951(.dina(n1934), .dinb(n1173), .dout(n2161));
  jor  g01952(.dina(n2161), .dinb(n2108), .dout(n2162));
  jxor g01953(.dina(n2162), .dinb(n1940), .dout(n2163));
  jor  g01954(.dina(n2163), .dinb(n2160), .dout(n2164));
  jand g01955(.dina(n2164), .dinb(n2159), .dout(n2165));
  jor  g01956(.dina(n2165), .dinb(n884), .dout(n2166));
  jand g01957(.dina(n2165), .dinb(n884), .dout(n2167));
  jxor g01958(.dina(n1942), .dinb(n1008), .dout(n2168));
  jor  g01959(.dina(n2168), .dinb(n2108), .dout(n2169));
  jxor g01960(.dina(n2169), .dinb(n1948), .dout(n2170));
  jor  g01961(.dina(n2170), .dinb(n2167), .dout(n2171));
  jand g01962(.dina(n2171), .dinb(n2166), .dout(n2172));
  jor  g01963(.dina(n2172), .dinb(n743), .dout(n2173));
  jand g01964(.dina(n2172), .dinb(n743), .dout(n2174));
  jxor g01965(.dina(n1950), .dinb(n884), .dout(n2175));
  jor  g01966(.dina(n2175), .dinb(n2108), .dout(n2176));
  jxor g01967(.dina(n2176), .dinb(n2050), .dout(n2177));
  jnot g01968(.din(n2177), .dout(n2178));
  jor  g01969(.dina(n2178), .dinb(n2174), .dout(n2179));
  jand g01970(.dina(n2179), .dinb(n2173), .dout(n2180));
  jor  g01971(.dina(n2180), .dinb(n635), .dout(n2181));
  jand g01972(.dina(n2180), .dinb(n635), .dout(n2182));
  jxor g01973(.dina(n1957), .dinb(n743), .dout(n2183));
  jor  g01974(.dina(n2183), .dinb(n2108), .dout(n2184));
  jxor g01975(.dina(n2184), .dinb(n2054), .dout(n2185));
  jnot g01976(.din(n2185), .dout(n2186));
  jor  g01977(.dina(n2186), .dinb(n2182), .dout(n2187));
  jand g01978(.dina(n2187), .dinb(n2181), .dout(n2188));
  jor  g01979(.dina(n2188), .dinb(n515), .dout(n2189));
  jand g01980(.dina(n2188), .dinb(n515), .dout(n2190));
  jxor g01981(.dina(n1964), .dinb(n635), .dout(n2191));
  jor  g01982(.dina(n2191), .dinb(n2108), .dout(n2192));
  jxor g01983(.dina(n2192), .dinb(n1970), .dout(n2193));
  jor  g01984(.dina(n2193), .dinb(n2190), .dout(n2194));
  jand g01985(.dina(n2194), .dinb(n2189), .dout(n2195));
  jor  g01986(.dina(n2195), .dinb(n443), .dout(n2196));
  jand g01987(.dina(n2195), .dinb(n443), .dout(n2197));
  jxor g01988(.dina(n1972), .dinb(n515), .dout(n2198));
  jor  g01989(.dina(n2198), .dinb(n2108), .dout(n2199));
  jxor g01990(.dina(n2199), .dinb(n1978), .dout(n2200));
  jor  g01991(.dina(n2200), .dinb(n2197), .dout(n2201));
  jand g01992(.dina(n2201), .dinb(n2196), .dout(n2202));
  jor  g01993(.dina(n2202), .dinb(n352), .dout(n2203));
  jand g01994(.dina(n2202), .dinb(n352), .dout(n2204));
  jxor g01995(.dina(n1980), .dinb(n443), .dout(n2205));
  jor  g01996(.dina(n2205), .dinb(n2108), .dout(n2206));
  jxor g01997(.dina(n2206), .dinb(n1985), .dout(n2207));
  jnot g01998(.din(n2207), .dout(n2208));
  jor  g01999(.dina(n2208), .dinb(n2204), .dout(n2209));
  jand g02000(.dina(n2209), .dinb(n2203), .dout(n2210));
  jor  g02001(.dina(n2210), .dinb(n294), .dout(n2211));
  jand g02002(.dina(n2210), .dinb(n294), .dout(n2212));
  jxor g02003(.dina(n1988), .dinb(n352), .dout(n2213));
  jor  g02004(.dina(n2213), .dinb(n2108), .dout(n2214));
  jxor g02005(.dina(n2214), .dinb(n2067), .dout(n2215));
  jnot g02006(.din(n2215), .dout(n2216));
  jor  g02007(.dina(n2216), .dinb(n2212), .dout(n2217));
  jand g02008(.dina(n2217), .dinb(n2211), .dout(n2218));
  jor  g02009(.dina(n2218), .dinb(n239), .dout(n2219));
  jand g02010(.dina(n2218), .dinb(n239), .dout(n2220));
  jxor g02011(.dina(n1995), .dinb(n294), .dout(n2221));
  jor  g02012(.dina(n2221), .dinb(n2108), .dout(n2222));
  jxor g02013(.dina(n2222), .dinb(n2001), .dout(n2223));
  jor  g02014(.dina(n2223), .dinb(n2220), .dout(n2224));
  jand g02015(.dina(n2224), .dinb(n2219), .dout(n2225));
  jor  g02016(.dina(n2225), .dinb(n221), .dout(n2226));
  jand g02017(.dina(n2225), .dinb(n221), .dout(n2227));
  jxor g02018(.dina(n2003), .dinb(n239), .dout(n2228));
  jor  g02019(.dina(n2228), .dinb(n2108), .dout(n2229));
  jxor g02020(.dina(n2229), .dinb(n2009), .dout(n2230));
  jor  g02021(.dina(n2230), .dinb(n2227), .dout(n2231));
  jand g02022(.dina(n2231), .dinb(n2226), .dout(n2232));
  jxor g02023(.dina(n2011), .dinb(n221), .dout(n2233));
  jor  g02024(.dina(n2233), .dinb(n2108), .dout(n2234));
  jxor g02025(.dina(n2234), .dinb(n2089), .dout(n2235));
  jand g02026(.dina(n2235), .dinb(n2232), .dout(n2236));
  jor  g02027(.dina(n2235), .dinb(n2232), .dout(n2238));
  jand g02028(.dina(asqrt[47] ), .dinb(n2104), .dout(n2239));
  jor  g02029(.dina(n2239), .dinb(n2128), .dout(n2240));
  jor  g02030(.dina(n2240), .dinb(n2238), .dout(n2241));
  jand g02031(.dina(n2241), .dinb(n218), .dout(n2242));
  jand g02032(.dina(n2108), .dinb(n2081), .dout(n2243));
  jand g02033(.dina(n2082), .dinb(asqrt[63] ), .dout(n2244));
  jand g02034(.dina(n2244), .dinb(n2092), .dout(n2245));
  jnot g02035(.din(n2245), .dout(n2246));
  jor  g02036(.dina(n2246), .dinb(n2243), .dout(n2247));
  jnot g02037(.din(n2247), .dout(n2248));
  jor  g02038(.dina(n2248), .dinb(n2242), .dout(n2249));
  jor  g02039(.dina(n2249), .dinb(n2236), .dout(asqrt[46] ));
  jnot g02040(.din(a[90] ), .dout(n2252));
  jnot g02041(.din(a[91] ), .dout(n2253));
  jand g02042(.dina(n2253), .dinb(n2252), .dout(n2254));
  jand g02043(.dina(n2254), .dinb(n2110), .dout(n2255));
  jand g02044(.dina(asqrt[46] ), .dinb(a[92] ), .dout(n2256));
  jor  g02045(.dina(n2256), .dinb(n2255), .dout(n2257));
  jand g02046(.dina(n2257), .dinb(asqrt[47] ), .dout(n2258));
  jor  g02047(.dina(n2257), .dinb(asqrt[47] ), .dout(n2259));
  jand g02048(.dina(asqrt[46] ), .dinb(n2110), .dout(n2260));
  jor  g02049(.dina(n2260), .dinb(n2111), .dout(n2261));
  jnot g02050(.din(n2112), .dout(n2262));
  jnot g02051(.din(n2236), .dout(n2263));
  jnot g02052(.din(n2226), .dout(n2265));
  jnot g02053(.din(n2219), .dout(n2266));
  jnot g02054(.din(n2211), .dout(n2267));
  jnot g02055(.din(n2203), .dout(n2268));
  jnot g02056(.din(n2196), .dout(n2269));
  jnot g02057(.din(n2189), .dout(n2270));
  jnot g02058(.din(n2181), .dout(n2271));
  jnot g02059(.din(n2173), .dout(n2272));
  jnot g02060(.din(n2166), .dout(n2273));
  jnot g02061(.din(n2159), .dout(n2274));
  jnot g02062(.din(n2151), .dout(n2275));
  jnot g02063(.din(n2144), .dout(n2276));
  jnot g02064(.din(n2136), .dout(n2277));
  jnot g02065(.din(n2124), .dout(n2278));
  jnot g02066(.din(n2116), .dout(n2279));
  jand g02067(.dina(asqrt[47] ), .dinb(a[94] ), .dout(n2280));
  jor  g02068(.dina(n2113), .dinb(n2280), .dout(n2281));
  jor  g02069(.dina(n2281), .dinb(asqrt[48] ), .dout(n2282));
  jand g02070(.dina(asqrt[47] ), .dinb(n1894), .dout(n2283));
  jor  g02071(.dina(n2283), .dinb(n1895), .dout(n2284));
  jand g02072(.dina(n2127), .dinb(n2284), .dout(n2285));
  jand g02073(.dina(n2285), .dinb(n2282), .dout(n2286));
  jor  g02074(.dina(n2286), .dinb(n2279), .dout(n2287));
  jor  g02075(.dina(n2287), .dinb(asqrt[49] ), .dout(n2288));
  jnot g02076(.din(n2133), .dout(n2289));
  jand g02077(.dina(n2289), .dinb(n2288), .dout(n2290));
  jor  g02078(.dina(n2290), .dinb(n2278), .dout(n2291));
  jor  g02079(.dina(n2291), .dinb(asqrt[50] ), .dout(n2292));
  jand g02080(.dina(n2140), .dinb(n2292), .dout(n2293));
  jor  g02081(.dina(n2293), .dinb(n2277), .dout(n2294));
  jor  g02082(.dina(n2294), .dinb(asqrt[51] ), .dout(n2295));
  jnot g02083(.din(n2148), .dout(n2296));
  jand g02084(.dina(n2296), .dinb(n2295), .dout(n2297));
  jor  g02085(.dina(n2297), .dinb(n2276), .dout(n2298));
  jor  g02086(.dina(n2298), .dinb(asqrt[52] ), .dout(n2299));
  jand g02087(.dina(n2155), .dinb(n2299), .dout(n2300));
  jor  g02088(.dina(n2300), .dinb(n2275), .dout(n2301));
  jor  g02089(.dina(n2301), .dinb(asqrt[53] ), .dout(n2302));
  jnot g02090(.din(n2163), .dout(n2303));
  jand g02091(.dina(n2303), .dinb(n2302), .dout(n2304));
  jor  g02092(.dina(n2304), .dinb(n2274), .dout(n2305));
  jor  g02093(.dina(n2305), .dinb(asqrt[54] ), .dout(n2306));
  jnot g02094(.din(n2170), .dout(n2307));
  jand g02095(.dina(n2307), .dinb(n2306), .dout(n2308));
  jor  g02096(.dina(n2308), .dinb(n2273), .dout(n2309));
  jor  g02097(.dina(n2309), .dinb(asqrt[55] ), .dout(n2310));
  jand g02098(.dina(n2177), .dinb(n2310), .dout(n2311));
  jor  g02099(.dina(n2311), .dinb(n2272), .dout(n2312));
  jor  g02100(.dina(n2312), .dinb(asqrt[56] ), .dout(n2313));
  jand g02101(.dina(n2185), .dinb(n2313), .dout(n2314));
  jor  g02102(.dina(n2314), .dinb(n2271), .dout(n2315));
  jor  g02103(.dina(n2315), .dinb(asqrt[57] ), .dout(n2316));
  jnot g02104(.din(n2193), .dout(n2317));
  jand g02105(.dina(n2317), .dinb(n2316), .dout(n2318));
  jor  g02106(.dina(n2318), .dinb(n2270), .dout(n2319));
  jor  g02107(.dina(n2319), .dinb(asqrt[58] ), .dout(n2320));
  jnot g02108(.din(n2200), .dout(n2321));
  jand g02109(.dina(n2321), .dinb(n2320), .dout(n2322));
  jor  g02110(.dina(n2322), .dinb(n2269), .dout(n2323));
  jor  g02111(.dina(n2323), .dinb(asqrt[59] ), .dout(n2324));
  jand g02112(.dina(n2207), .dinb(n2324), .dout(n2325));
  jor  g02113(.dina(n2325), .dinb(n2268), .dout(n2326));
  jor  g02114(.dina(n2326), .dinb(asqrt[60] ), .dout(n2327));
  jand g02115(.dina(n2215), .dinb(n2327), .dout(n2328));
  jor  g02116(.dina(n2328), .dinb(n2267), .dout(n2329));
  jor  g02117(.dina(n2329), .dinb(asqrt[61] ), .dout(n2330));
  jnot g02118(.din(n2223), .dout(n2331));
  jand g02119(.dina(n2331), .dinb(n2330), .dout(n2332));
  jor  g02120(.dina(n2332), .dinb(n2266), .dout(n2333));
  jor  g02121(.dina(n2333), .dinb(asqrt[62] ), .dout(n2334));
  jnot g02122(.din(n2230), .dout(n2335));
  jand g02123(.dina(n2335), .dinb(n2334), .dout(n2336));
  jor  g02124(.dina(n2336), .dinb(n2265), .dout(n2337));
  jnot g02125(.din(n2235), .dout(n2338));
  jand g02126(.dina(n2338), .dinb(n2337), .dout(n2339));
  jnot g02127(.din(n2240), .dout(n2340));
  jand g02128(.dina(n2340), .dinb(n2339), .dout(n2341));
  jor  g02129(.dina(n2341), .dinb(asqrt[63] ), .dout(n2342));
  jand g02130(.dina(n2247), .dinb(n2342), .dout(n2343));
  jand g02131(.dina(n2343), .dinb(n2263), .dout(n2345));
  jor  g02132(.dina(n2345), .dinb(n2262), .dout(n2346));
  jand g02133(.dina(n2346), .dinb(n2261), .dout(n2347));
  jand g02134(.dina(n2347), .dinb(n2259), .dout(n2348));
  jor  g02135(.dina(n2348), .dinb(n2258), .dout(n2349));
  jand g02136(.dina(n2349), .dinb(asqrt[48] ), .dout(n2350));
  jor  g02137(.dina(n2349), .dinb(asqrt[48] ), .dout(n2351));
  jand g02138(.dina(asqrt[46] ), .dinb(n2112), .dout(n2352));
  jand g02139(.dina(n2263), .dinb(asqrt[47] ), .dout(n2353));
  jand g02140(.dina(n2353), .dinb(n2246), .dout(n2354));
  jand g02141(.dina(n2354), .dinb(n2342), .dout(n2355));
  jor  g02142(.dina(n2355), .dinb(n2352), .dout(n2356));
  jxor g02143(.dina(n2356), .dinb(a[94] ), .dout(n2357));
  jnot g02144(.din(n2357), .dout(n2358));
  jand g02145(.dina(n2358), .dinb(n2351), .dout(n2359));
  jor  g02146(.dina(n2359), .dinb(n2350), .dout(n2360));
  jand g02147(.dina(n2360), .dinb(asqrt[49] ), .dout(n2361));
  jor  g02148(.dina(n2360), .dinb(asqrt[49] ), .dout(n2362));
  jxor g02149(.dina(n2115), .dinb(n1912), .dout(n2363));
  jand g02150(.dina(n2363), .dinb(asqrt[46] ), .dout(n2364));
  jxor g02151(.dina(n2364), .dinb(n2285), .dout(n2365));
  jand g02152(.dina(n2365), .dinb(n2362), .dout(n2366));
  jor  g02153(.dina(n2366), .dinb(n2361), .dout(n2367));
  jand g02154(.dina(n2367), .dinb(asqrt[50] ), .dout(n2368));
  jor  g02155(.dina(n2367), .dinb(asqrt[50] ), .dout(n2369));
  jxor g02156(.dina(n2123), .dinb(n1699), .dout(n2370));
  jand g02157(.dina(n2370), .dinb(asqrt[46] ), .dout(n2371));
  jxor g02158(.dina(n2371), .dinb(n2133), .dout(n2372));
  jnot g02159(.din(n2372), .dout(n2373));
  jand g02160(.dina(n2373), .dinb(n2369), .dout(n2374));
  jor  g02161(.dina(n2374), .dinb(n2368), .dout(n2375));
  jand g02162(.dina(n2375), .dinb(asqrt[51] ), .dout(n2376));
  jor  g02163(.dina(n2375), .dinb(asqrt[51] ), .dout(n2377));
  jxor g02164(.dina(n2135), .dinb(n1516), .dout(n2378));
  jand g02165(.dina(n2378), .dinb(asqrt[46] ), .dout(n2379));
  jxor g02166(.dina(n2379), .dinb(n2140), .dout(n2380));
  jand g02167(.dina(n2380), .dinb(n2377), .dout(n2381));
  jor  g02168(.dina(n2381), .dinb(n2376), .dout(n2382));
  jand g02169(.dina(n2382), .dinb(asqrt[52] ), .dout(n2383));
  jor  g02170(.dina(n2382), .dinb(asqrt[52] ), .dout(n2384));
  jxor g02171(.dina(n2143), .dinb(n1332), .dout(n2385));
  jand g02172(.dina(n2385), .dinb(asqrt[46] ), .dout(n2386));
  jxor g02173(.dina(n2386), .dinb(n2148), .dout(n2387));
  jnot g02174(.din(n2387), .dout(n2388));
  jand g02175(.dina(n2388), .dinb(n2384), .dout(n2389));
  jor  g02176(.dina(n2389), .dinb(n2383), .dout(n2390));
  jand g02177(.dina(n2390), .dinb(asqrt[53] ), .dout(n2391));
  jor  g02178(.dina(n2390), .dinb(asqrt[53] ), .dout(n2392));
  jxor g02179(.dina(n2150), .dinb(n1173), .dout(n2393));
  jand g02180(.dina(n2393), .dinb(asqrt[46] ), .dout(n2394));
  jxor g02181(.dina(n2394), .dinb(n2155), .dout(n2395));
  jand g02182(.dina(n2395), .dinb(n2392), .dout(n2396));
  jor  g02183(.dina(n2396), .dinb(n2391), .dout(n2397));
  jand g02184(.dina(n2397), .dinb(asqrt[54] ), .dout(n2398));
  jor  g02185(.dina(n2397), .dinb(asqrt[54] ), .dout(n2399));
  jxor g02186(.dina(n2158), .dinb(n1008), .dout(n2400));
  jand g02187(.dina(n2400), .dinb(asqrt[46] ), .dout(n2401));
  jxor g02188(.dina(n2401), .dinb(n2163), .dout(n2402));
  jnot g02189(.din(n2402), .dout(n2403));
  jand g02190(.dina(n2403), .dinb(n2399), .dout(n2404));
  jor  g02191(.dina(n2404), .dinb(n2398), .dout(n2405));
  jand g02192(.dina(n2405), .dinb(asqrt[55] ), .dout(n2406));
  jor  g02193(.dina(n2405), .dinb(asqrt[55] ), .dout(n2407));
  jxor g02194(.dina(n2165), .dinb(n884), .dout(n2408));
  jand g02195(.dina(n2408), .dinb(asqrt[46] ), .dout(n2409));
  jxor g02196(.dina(n2409), .dinb(n2170), .dout(n2410));
  jnot g02197(.din(n2410), .dout(n2411));
  jand g02198(.dina(n2411), .dinb(n2407), .dout(n2412));
  jor  g02199(.dina(n2412), .dinb(n2406), .dout(n2413));
  jand g02200(.dina(n2413), .dinb(asqrt[56] ), .dout(n2414));
  jor  g02201(.dina(n2413), .dinb(asqrt[56] ), .dout(n2415));
  jxor g02202(.dina(n2172), .dinb(n743), .dout(n2416));
  jand g02203(.dina(n2416), .dinb(asqrt[46] ), .dout(n2417));
  jxor g02204(.dina(n2417), .dinb(n2177), .dout(n2418));
  jand g02205(.dina(n2418), .dinb(n2415), .dout(n2419));
  jor  g02206(.dina(n2419), .dinb(n2414), .dout(n2420));
  jand g02207(.dina(n2420), .dinb(asqrt[57] ), .dout(n2421));
  jor  g02208(.dina(n2420), .dinb(asqrt[57] ), .dout(n2422));
  jxor g02209(.dina(n2180), .dinb(n635), .dout(n2423));
  jand g02210(.dina(n2423), .dinb(asqrt[46] ), .dout(n2424));
  jxor g02211(.dina(n2424), .dinb(n2185), .dout(n2425));
  jand g02212(.dina(n2425), .dinb(n2422), .dout(n2426));
  jor  g02213(.dina(n2426), .dinb(n2421), .dout(n2427));
  jand g02214(.dina(n2427), .dinb(asqrt[58] ), .dout(n2428));
  jor  g02215(.dina(n2427), .dinb(asqrt[58] ), .dout(n2429));
  jxor g02216(.dina(n2188), .dinb(n515), .dout(n2430));
  jand g02217(.dina(n2430), .dinb(asqrt[46] ), .dout(n2431));
  jxor g02218(.dina(n2431), .dinb(n2193), .dout(n2432));
  jnot g02219(.din(n2432), .dout(n2433));
  jand g02220(.dina(n2433), .dinb(n2429), .dout(n2434));
  jor  g02221(.dina(n2434), .dinb(n2428), .dout(n2435));
  jand g02222(.dina(n2435), .dinb(asqrt[59] ), .dout(n2436));
  jor  g02223(.dina(n2435), .dinb(asqrt[59] ), .dout(n2437));
  jxor g02224(.dina(n2195), .dinb(n443), .dout(n2438));
  jand g02225(.dina(n2438), .dinb(asqrt[46] ), .dout(n2439));
  jxor g02226(.dina(n2439), .dinb(n2321), .dout(n2440));
  jand g02227(.dina(n2440), .dinb(n2437), .dout(n2441));
  jor  g02228(.dina(n2441), .dinb(n2436), .dout(n2442));
  jand g02229(.dina(n2442), .dinb(asqrt[60] ), .dout(n2443));
  jor  g02230(.dina(n2442), .dinb(asqrt[60] ), .dout(n2444));
  jxor g02231(.dina(n2202), .dinb(n352), .dout(n2445));
  jand g02232(.dina(n2445), .dinb(asqrt[46] ), .dout(n2446));
  jxor g02233(.dina(n2446), .dinb(n2207), .dout(n2447));
  jand g02234(.dina(n2447), .dinb(n2444), .dout(n2448));
  jor  g02235(.dina(n2448), .dinb(n2443), .dout(n2449));
  jand g02236(.dina(n2449), .dinb(asqrt[61] ), .dout(n2450));
  jor  g02237(.dina(n2449), .dinb(asqrt[61] ), .dout(n2451));
  jxor g02238(.dina(n2210), .dinb(n294), .dout(n2452));
  jand g02239(.dina(n2452), .dinb(asqrt[46] ), .dout(n2453));
  jxor g02240(.dina(n2453), .dinb(n2215), .dout(n2454));
  jand g02241(.dina(n2454), .dinb(n2451), .dout(n2455));
  jor  g02242(.dina(n2455), .dinb(n2450), .dout(n2456));
  jand g02243(.dina(n2456), .dinb(asqrt[62] ), .dout(n2457));
  jor  g02244(.dina(n2456), .dinb(asqrt[62] ), .dout(n2458));
  jxor g02245(.dina(n2218), .dinb(n239), .dout(n2459));
  jand g02246(.dina(n2459), .dinb(asqrt[46] ), .dout(n2460));
  jxor g02247(.dina(n2460), .dinb(n2223), .dout(n2461));
  jnot g02248(.din(n2461), .dout(n2462));
  jand g02249(.dina(n2462), .dinb(n2458), .dout(n2463));
  jor  g02250(.dina(n2463), .dinb(n2457), .dout(n2464));
  jxor g02251(.dina(n2225), .dinb(n221), .dout(n2465));
  jand g02252(.dina(n2465), .dinb(asqrt[46] ), .dout(n2466));
  jxor g02253(.dina(n2466), .dinb(n2230), .dout(n2467));
  jnot g02254(.din(n2467), .dout(n2468));
  jor  g02255(.dina(n2468), .dinb(n2464), .dout(n2469));
  jnot g02256(.din(n2469), .dout(n2470));
  jand g02257(.dina(n2343), .dinb(n2232), .dout(n2471));
  jnot g02258(.din(n2471), .dout(n2472));
  jand g02259(.dina(n2238), .dinb(asqrt[63] ), .dout(n2473));
  jand g02260(.dina(n2473), .dinb(n2263), .dout(n2474));
  jand g02261(.dina(n2474), .dinb(n2472), .dout(n2475));
  jand g02262(.dina(n2249), .dinb(n2339), .dout(n2476));
  jnot g02263(.din(n2457), .dout(n2477));
  jnot g02264(.din(n2450), .dout(n2478));
  jnot g02265(.din(n2443), .dout(n2479));
  jnot g02266(.din(n2436), .dout(n2480));
  jnot g02267(.din(n2428), .dout(n2481));
  jnot g02268(.din(n2421), .dout(n2482));
  jnot g02269(.din(n2414), .dout(n2483));
  jnot g02270(.din(n2406), .dout(n2484));
  jnot g02271(.din(n2398), .dout(n2485));
  jnot g02272(.din(n2391), .dout(n2486));
  jnot g02273(.din(n2383), .dout(n2487));
  jnot g02274(.din(n2376), .dout(n2488));
  jnot g02275(.din(n2368), .dout(n2489));
  jnot g02276(.din(n2361), .dout(n2490));
  jnot g02277(.din(n2350), .dout(n2491));
  jnot g02278(.din(n2258), .dout(n2492));
  jnot g02279(.din(n2255), .dout(n2493));
  jor  g02280(.dina(n2345), .dinb(n2110), .dout(n2494));
  jand g02281(.dina(n2494), .dinb(n2493), .dout(n2495));
  jand g02282(.dina(n2495), .dinb(n2108), .dout(n2496));
  jor  g02283(.dina(n2345), .dinb(a[92] ), .dout(n2497));
  jand g02284(.dina(n2497), .dinb(a[93] ), .dout(n2498));
  jor  g02285(.dina(n2352), .dinb(n2498), .dout(n2499));
  jor  g02286(.dina(n2499), .dinb(n2496), .dout(n2500));
  jand g02287(.dina(n2500), .dinb(n2492), .dout(n2501));
  jand g02288(.dina(n2501), .dinb(n1912), .dout(n2502));
  jor  g02289(.dina(n2357), .dinb(n2502), .dout(n2503));
  jand g02290(.dina(n2503), .dinb(n2491), .dout(n2504));
  jand g02291(.dina(n2504), .dinb(n1699), .dout(n2505));
  jnot g02292(.din(n2365), .dout(n2506));
  jor  g02293(.dina(n2506), .dinb(n2505), .dout(n2507));
  jand g02294(.dina(n2507), .dinb(n2490), .dout(n2508));
  jand g02295(.dina(n2508), .dinb(n1516), .dout(n2509));
  jor  g02296(.dina(n2372), .dinb(n2509), .dout(n2510));
  jand g02297(.dina(n2510), .dinb(n2489), .dout(n2511));
  jand g02298(.dina(n2511), .dinb(n1332), .dout(n2512));
  jnot g02299(.din(n2380), .dout(n2513));
  jor  g02300(.dina(n2513), .dinb(n2512), .dout(n2514));
  jand g02301(.dina(n2514), .dinb(n2488), .dout(n2515));
  jand g02302(.dina(n2515), .dinb(n1173), .dout(n2516));
  jor  g02303(.dina(n2387), .dinb(n2516), .dout(n2517));
  jand g02304(.dina(n2517), .dinb(n2487), .dout(n2518));
  jand g02305(.dina(n2518), .dinb(n1008), .dout(n2519));
  jnot g02306(.din(n2395), .dout(n2520));
  jor  g02307(.dina(n2520), .dinb(n2519), .dout(n2521));
  jand g02308(.dina(n2521), .dinb(n2486), .dout(n2522));
  jand g02309(.dina(n2522), .dinb(n884), .dout(n2523));
  jor  g02310(.dina(n2402), .dinb(n2523), .dout(n2524));
  jand g02311(.dina(n2524), .dinb(n2485), .dout(n2525));
  jand g02312(.dina(n2525), .dinb(n743), .dout(n2526));
  jor  g02313(.dina(n2410), .dinb(n2526), .dout(n2527));
  jand g02314(.dina(n2527), .dinb(n2484), .dout(n2528));
  jand g02315(.dina(n2528), .dinb(n635), .dout(n2529));
  jnot g02316(.din(n2418), .dout(n2530));
  jor  g02317(.dina(n2530), .dinb(n2529), .dout(n2531));
  jand g02318(.dina(n2531), .dinb(n2483), .dout(n2532));
  jand g02319(.dina(n2532), .dinb(n515), .dout(n2533));
  jnot g02320(.din(n2425), .dout(n2534));
  jor  g02321(.dina(n2534), .dinb(n2533), .dout(n2535));
  jand g02322(.dina(n2535), .dinb(n2482), .dout(n2536));
  jand g02323(.dina(n2536), .dinb(n443), .dout(n2537));
  jor  g02324(.dina(n2432), .dinb(n2537), .dout(n2538));
  jand g02325(.dina(n2538), .dinb(n2481), .dout(n2539));
  jand g02326(.dina(n2539), .dinb(n352), .dout(n2540));
  jnot g02327(.din(n2440), .dout(n2541));
  jor  g02328(.dina(n2541), .dinb(n2540), .dout(n2542));
  jand g02329(.dina(n2542), .dinb(n2480), .dout(n2543));
  jand g02330(.dina(n2543), .dinb(n294), .dout(n2544));
  jnot g02331(.din(n2447), .dout(n2545));
  jor  g02332(.dina(n2545), .dinb(n2544), .dout(n2546));
  jand g02333(.dina(n2546), .dinb(n2479), .dout(n2547));
  jand g02334(.dina(n2547), .dinb(n239), .dout(n2548));
  jnot g02335(.din(n2454), .dout(n2549));
  jor  g02336(.dina(n2549), .dinb(n2548), .dout(n2550));
  jand g02337(.dina(n2550), .dinb(n2478), .dout(n2551));
  jand g02338(.dina(n2551), .dinb(n221), .dout(n2552));
  jor  g02339(.dina(n2461), .dinb(n2552), .dout(n2553));
  jand g02340(.dina(n2553), .dinb(n2477), .dout(n2554));
  jor  g02341(.dina(n2467), .dinb(n2554), .dout(n2555));
  jor  g02342(.dina(n2555), .dinb(n2236), .dout(n2556));
  jor  g02343(.dina(n2556), .dinb(n2476), .dout(n2557));
  jand g02344(.dina(n2557), .dinb(n218), .dout(n2558));
  jand g02345(.dina(n2345), .dinb(n2235), .dout(n2559));
  jor  g02346(.dina(n2559), .dinb(n2558), .dout(n2560));
  jor  g02347(.dina(n2560), .dinb(n2475), .dout(n2561));
  jor  g02348(.dina(n2561), .dinb(n2470), .dout(asqrt[45] ));
  jnot g02349(.din(n2475), .dout(n2563));
  jnot g02350(.din(n2476), .dout(n2564));
  jand g02351(.dina(n2468), .dinb(n2464), .dout(n2565));
  jand g02352(.dina(n2565), .dinb(n2263), .dout(n2566));
  jand g02353(.dina(n2566), .dinb(n2564), .dout(n2567));
  jor  g02354(.dina(n2567), .dinb(asqrt[63] ), .dout(n2568));
  jnot g02355(.din(n2559), .dout(n2569));
  jand g02356(.dina(n2569), .dinb(n2568), .dout(n2570));
  jand g02357(.dina(n2570), .dinb(n2563), .dout(n2571));
  jand g02358(.dina(n2571), .dinb(n2469), .dout(n2572));
  jxor g02359(.dina(n2456), .dinb(n221), .dout(n2573));
  jor  g02360(.dina(n2573), .dinb(n2572), .dout(n2574));
  jxor g02361(.dina(n2574), .dinb(n2461), .dout(n2575));
  jnot g02362(.din(n2575), .dout(n2576));
  jor  g02363(.dina(n2572), .dinb(n2252), .dout(n2577));
  jnot g02364(.din(a[88] ), .dout(n2578));
  jnot g02365(.din(a[89] ), .dout(n2579));
  jand g02366(.dina(n2579), .dinb(n2578), .dout(n2580));
  jand g02367(.dina(n2580), .dinb(n2252), .dout(n2581));
  jnot g02368(.din(n2581), .dout(n2582));
  jand g02369(.dina(n2582), .dinb(n2577), .dout(n2583));
  jor  g02370(.dina(n2583), .dinb(n2345), .dout(n2584));
  jand g02371(.dina(n2583), .dinb(n2345), .dout(n2585));
  jor  g02372(.dina(n2572), .dinb(a[90] ), .dout(n2586));
  jand g02373(.dina(n2586), .dinb(a[91] ), .dout(n2587));
  jand g02374(.dina(asqrt[45] ), .dinb(n2254), .dout(n2588));
  jor  g02375(.dina(n2588), .dinb(n2587), .dout(n2589));
  jor  g02376(.dina(n2589), .dinb(n2585), .dout(n2590));
  jand g02377(.dina(n2590), .dinb(n2584), .dout(n2591));
  jor  g02378(.dina(n2591), .dinb(n2108), .dout(n2592));
  jand g02379(.dina(n2591), .dinb(n2108), .dout(n2593));
  jnot g02380(.din(n2254), .dout(n2594));
  jor  g02381(.dina(n2572), .dinb(n2594), .dout(n2595));
  jor  g02382(.dina(n2470), .dinb(n2345), .dout(n2596));
  jor  g02383(.dina(n2596), .dinb(n2474), .dout(n2597));
  jor  g02384(.dina(n2597), .dinb(n2558), .dout(n2598));
  jand g02385(.dina(n2598), .dinb(n2595), .dout(n2599));
  jxor g02386(.dina(n2599), .dinb(n2110), .dout(n2600));
  jor  g02387(.dina(n2600), .dinb(n2593), .dout(n2601));
  jand g02388(.dina(n2601), .dinb(n2592), .dout(n2602));
  jor  g02389(.dina(n2602), .dinb(n1912), .dout(n2603));
  jand g02390(.dina(n2602), .dinb(n1912), .dout(n2604));
  jxor g02391(.dina(n2257), .dinb(n2108), .dout(n2605));
  jor  g02392(.dina(n2605), .dinb(n2572), .dout(n2606));
  jxor g02393(.dina(n2606), .dinb(n2499), .dout(n2607));
  jnot g02394(.din(n2607), .dout(n2608));
  jor  g02395(.dina(n2608), .dinb(n2604), .dout(n2609));
  jand g02396(.dina(n2609), .dinb(n2603), .dout(n2610));
  jor  g02397(.dina(n2610), .dinb(n1699), .dout(n2611));
  jand g02398(.dina(n2610), .dinb(n1699), .dout(n2612));
  jxor g02399(.dina(n2349), .dinb(n1912), .dout(n2613));
  jor  g02400(.dina(n2613), .dinb(n2572), .dout(n2614));
  jxor g02401(.dina(n2614), .dinb(n2358), .dout(n2615));
  jor  g02402(.dina(n2615), .dinb(n2612), .dout(n2616));
  jand g02403(.dina(n2616), .dinb(n2611), .dout(n2617));
  jor  g02404(.dina(n2617), .dinb(n1516), .dout(n2618));
  jand g02405(.dina(n2617), .dinb(n1516), .dout(n2619));
  jxor g02406(.dina(n2360), .dinb(n1699), .dout(n2620));
  jor  g02407(.dina(n2620), .dinb(n2572), .dout(n2621));
  jxor g02408(.dina(n2621), .dinb(n2506), .dout(n2622));
  jnot g02409(.din(n2622), .dout(n2623));
  jor  g02410(.dina(n2623), .dinb(n2619), .dout(n2624));
  jand g02411(.dina(n2624), .dinb(n2618), .dout(n2625));
  jor  g02412(.dina(n2625), .dinb(n1332), .dout(n2626));
  jand g02413(.dina(n2625), .dinb(n1332), .dout(n2627));
  jxor g02414(.dina(n2367), .dinb(n1516), .dout(n2628));
  jor  g02415(.dina(n2628), .dinb(n2572), .dout(n2629));
  jxor g02416(.dina(n2629), .dinb(n2373), .dout(n2630));
  jor  g02417(.dina(n2630), .dinb(n2627), .dout(n2631));
  jand g02418(.dina(n2631), .dinb(n2626), .dout(n2632));
  jor  g02419(.dina(n2632), .dinb(n1173), .dout(n2633));
  jand g02420(.dina(n2632), .dinb(n1173), .dout(n2634));
  jxor g02421(.dina(n2375), .dinb(n1332), .dout(n2635));
  jor  g02422(.dina(n2635), .dinb(n2572), .dout(n2636));
  jxor g02423(.dina(n2636), .dinb(n2513), .dout(n2637));
  jnot g02424(.din(n2637), .dout(n2638));
  jor  g02425(.dina(n2638), .dinb(n2634), .dout(n2639));
  jand g02426(.dina(n2639), .dinb(n2633), .dout(n2640));
  jor  g02427(.dina(n2640), .dinb(n1008), .dout(n2641));
  jand g02428(.dina(n2640), .dinb(n1008), .dout(n2642));
  jxor g02429(.dina(n2382), .dinb(n1173), .dout(n2643));
  jor  g02430(.dina(n2643), .dinb(n2572), .dout(n2644));
  jxor g02431(.dina(n2644), .dinb(n2388), .dout(n2645));
  jor  g02432(.dina(n2645), .dinb(n2642), .dout(n2646));
  jand g02433(.dina(n2646), .dinb(n2641), .dout(n2647));
  jor  g02434(.dina(n2647), .dinb(n884), .dout(n2648));
  jand g02435(.dina(n2647), .dinb(n884), .dout(n2649));
  jxor g02436(.dina(n2390), .dinb(n1008), .dout(n2650));
  jor  g02437(.dina(n2650), .dinb(n2572), .dout(n2651));
  jxor g02438(.dina(n2651), .dinb(n2520), .dout(n2652));
  jnot g02439(.din(n2652), .dout(n2653));
  jor  g02440(.dina(n2653), .dinb(n2649), .dout(n2654));
  jand g02441(.dina(n2654), .dinb(n2648), .dout(n2655));
  jor  g02442(.dina(n2655), .dinb(n743), .dout(n2656));
  jand g02443(.dina(n2655), .dinb(n743), .dout(n2657));
  jxor g02444(.dina(n2397), .dinb(n884), .dout(n2658));
  jor  g02445(.dina(n2658), .dinb(n2572), .dout(n2659));
  jxor g02446(.dina(n2659), .dinb(n2403), .dout(n2660));
  jor  g02447(.dina(n2660), .dinb(n2657), .dout(n2661));
  jand g02448(.dina(n2661), .dinb(n2656), .dout(n2662));
  jor  g02449(.dina(n2662), .dinb(n635), .dout(n2663));
  jand g02450(.dina(n2662), .dinb(n635), .dout(n2664));
  jxor g02451(.dina(n2405), .dinb(n743), .dout(n2665));
  jor  g02452(.dina(n2665), .dinb(n2572), .dout(n2666));
  jxor g02453(.dina(n2666), .dinb(n2411), .dout(n2667));
  jor  g02454(.dina(n2667), .dinb(n2664), .dout(n2668));
  jand g02455(.dina(n2668), .dinb(n2663), .dout(n2669));
  jor  g02456(.dina(n2669), .dinb(n515), .dout(n2670));
  jand g02457(.dina(n2669), .dinb(n515), .dout(n2671));
  jxor g02458(.dina(n2413), .dinb(n635), .dout(n2672));
  jor  g02459(.dina(n2672), .dinb(n2572), .dout(n2673));
  jxor g02460(.dina(n2673), .dinb(n2530), .dout(n2674));
  jnot g02461(.din(n2674), .dout(n2675));
  jor  g02462(.dina(n2675), .dinb(n2671), .dout(n2676));
  jand g02463(.dina(n2676), .dinb(n2670), .dout(n2677));
  jor  g02464(.dina(n2677), .dinb(n443), .dout(n2678));
  jand g02465(.dina(n2677), .dinb(n443), .dout(n2679));
  jxor g02466(.dina(n2420), .dinb(n515), .dout(n2680));
  jor  g02467(.dina(n2680), .dinb(n2572), .dout(n2681));
  jxor g02468(.dina(n2681), .dinb(n2534), .dout(n2682));
  jnot g02469(.din(n2682), .dout(n2683));
  jor  g02470(.dina(n2683), .dinb(n2679), .dout(n2684));
  jand g02471(.dina(n2684), .dinb(n2678), .dout(n2685));
  jor  g02472(.dina(n2685), .dinb(n352), .dout(n2686));
  jand g02473(.dina(n2685), .dinb(n352), .dout(n2687));
  jxor g02474(.dina(n2427), .dinb(n443), .dout(n2688));
  jor  g02475(.dina(n2688), .dinb(n2572), .dout(n2689));
  jxor g02476(.dina(n2689), .dinb(n2433), .dout(n2690));
  jor  g02477(.dina(n2690), .dinb(n2687), .dout(n2691));
  jand g02478(.dina(n2691), .dinb(n2686), .dout(n2692));
  jor  g02479(.dina(n2692), .dinb(n294), .dout(n2693));
  jand g02480(.dina(n2692), .dinb(n294), .dout(n2694));
  jxor g02481(.dina(n2435), .dinb(n352), .dout(n2695));
  jor  g02482(.dina(n2695), .dinb(n2572), .dout(n2696));
  jxor g02483(.dina(n2696), .dinb(n2541), .dout(n2697));
  jnot g02484(.din(n2697), .dout(n2698));
  jor  g02485(.dina(n2698), .dinb(n2694), .dout(n2699));
  jand g02486(.dina(n2699), .dinb(n2693), .dout(n2700));
  jor  g02487(.dina(n2700), .dinb(n239), .dout(n2701));
  jand g02488(.dina(n2700), .dinb(n239), .dout(n2702));
  jxor g02489(.dina(n2442), .dinb(n294), .dout(n2703));
  jor  g02490(.dina(n2703), .dinb(n2572), .dout(n2704));
  jxor g02491(.dina(n2704), .dinb(n2545), .dout(n2705));
  jnot g02492(.din(n2705), .dout(n2706));
  jor  g02493(.dina(n2706), .dinb(n2702), .dout(n2707));
  jand g02494(.dina(n2707), .dinb(n2701), .dout(n2708));
  jor  g02495(.dina(n2708), .dinb(n221), .dout(n2709));
  jand g02496(.dina(n2708), .dinb(n221), .dout(n2710));
  jxor g02497(.dina(n2449), .dinb(n239), .dout(n2711));
  jor  g02498(.dina(n2711), .dinb(n2572), .dout(n2712));
  jxor g02499(.dina(n2712), .dinb(n2549), .dout(n2713));
  jnot g02500(.din(n2713), .dout(n2714));
  jor  g02501(.dina(n2714), .dinb(n2710), .dout(n2715));
  jand g02502(.dina(n2715), .dinb(n2709), .dout(n2716));
  jand g02503(.dina(n2716), .dinb(n2576), .dout(n2717));
  jand g02504(.dina(n2561), .dinb(n2565), .dout(n2719));
  jor  g02505(.dina(n2716), .dinb(n2576), .dout(n2720));
  jor  g02506(.dina(n2720), .dinb(n2470), .dout(n2721));
  jor  g02507(.dina(n2721), .dinb(n2719), .dout(n2722));
  jand g02508(.dina(n2722), .dinb(n218), .dout(n2723));
  jand g02509(.dina(n2571), .dinb(n2554), .dout(n2724));
  jand g02510(.dina(n2555), .dinb(asqrt[63] ), .dout(n2725));
  jand g02511(.dina(n2725), .dinb(n2469), .dout(n2726));
  jnot g02512(.din(n2726), .dout(n2727));
  jor  g02513(.dina(n2727), .dinb(n2724), .dout(n2728));
  jnot g02514(.din(n2728), .dout(n2729));
  jor  g02515(.dina(n2729), .dinb(n2723), .dout(n2730));
  jor  g02516(.dina(n2730), .dinb(n2717), .dout(asqrt[44] ));
  jand g02517(.dina(asqrt[44] ), .dinb(a[88] ), .dout(n2733));
  jnot g02518(.din(a[86] ), .dout(n2734));
  jnot g02519(.din(a[87] ), .dout(n2735));
  jand g02520(.dina(n2735), .dinb(n2734), .dout(n2736));
  jand g02521(.dina(n2736), .dinb(n2578), .dout(n2737));
  jor  g02522(.dina(n2737), .dinb(n2733), .dout(n2738));
  jand g02523(.dina(n2738), .dinb(asqrt[45] ), .dout(n2739));
  jor  g02524(.dina(n2738), .dinb(asqrt[45] ), .dout(n2740));
  jand g02525(.dina(asqrt[44] ), .dinb(n2578), .dout(n2741));
  jor  g02526(.dina(n2741), .dinb(n2579), .dout(n2742));
  jnot g02527(.din(n2580), .dout(n2743));
  jnot g02528(.din(n2717), .dout(n2744));
  jnot g02529(.din(n2719), .dout(n2746));
  jnot g02530(.din(n2709), .dout(n2747));
  jnot g02531(.din(n2701), .dout(n2748));
  jnot g02532(.din(n2693), .dout(n2749));
  jnot g02533(.din(n2686), .dout(n2750));
  jnot g02534(.din(n2678), .dout(n2751));
  jnot g02535(.din(n2670), .dout(n2752));
  jnot g02536(.din(n2663), .dout(n2753));
  jnot g02537(.din(n2656), .dout(n2754));
  jnot g02538(.din(n2648), .dout(n2755));
  jnot g02539(.din(n2641), .dout(n2756));
  jnot g02540(.din(n2633), .dout(n2757));
  jnot g02541(.din(n2626), .dout(n2758));
  jnot g02542(.din(n2618), .dout(n2759));
  jnot g02543(.din(n2611), .dout(n2760));
  jnot g02544(.din(n2603), .dout(n2761));
  jnot g02545(.din(n2592), .dout(n2762));
  jnot g02546(.din(n2584), .dout(n2763));
  jand g02547(.dina(asqrt[45] ), .dinb(a[90] ), .dout(n2764));
  jor  g02548(.dina(n2581), .dinb(n2764), .dout(n2765));
  jor  g02549(.dina(n2765), .dinb(asqrt[46] ), .dout(n2766));
  jand g02550(.dina(asqrt[45] ), .dinb(n2252), .dout(n2767));
  jor  g02551(.dina(n2767), .dinb(n2253), .dout(n2768));
  jand g02552(.dina(n2595), .dinb(n2768), .dout(n2769));
  jand g02553(.dina(n2769), .dinb(n2766), .dout(n2770));
  jor  g02554(.dina(n2770), .dinb(n2763), .dout(n2771));
  jor  g02555(.dina(n2771), .dinb(asqrt[47] ), .dout(n2772));
  jnot g02556(.din(n2600), .dout(n2773));
  jand g02557(.dina(n2773), .dinb(n2772), .dout(n2774));
  jor  g02558(.dina(n2774), .dinb(n2762), .dout(n2775));
  jor  g02559(.dina(n2775), .dinb(asqrt[48] ), .dout(n2776));
  jand g02560(.dina(n2607), .dinb(n2776), .dout(n2777));
  jor  g02561(.dina(n2777), .dinb(n2761), .dout(n2778));
  jor  g02562(.dina(n2778), .dinb(asqrt[49] ), .dout(n2779));
  jnot g02563(.din(n2615), .dout(n2780));
  jand g02564(.dina(n2780), .dinb(n2779), .dout(n2781));
  jor  g02565(.dina(n2781), .dinb(n2760), .dout(n2782));
  jor  g02566(.dina(n2782), .dinb(asqrt[50] ), .dout(n2783));
  jand g02567(.dina(n2622), .dinb(n2783), .dout(n2784));
  jor  g02568(.dina(n2784), .dinb(n2759), .dout(n2785));
  jor  g02569(.dina(n2785), .dinb(asqrt[51] ), .dout(n2786));
  jnot g02570(.din(n2630), .dout(n2787));
  jand g02571(.dina(n2787), .dinb(n2786), .dout(n2788));
  jor  g02572(.dina(n2788), .dinb(n2758), .dout(n2789));
  jor  g02573(.dina(n2789), .dinb(asqrt[52] ), .dout(n2790));
  jand g02574(.dina(n2637), .dinb(n2790), .dout(n2791));
  jor  g02575(.dina(n2791), .dinb(n2757), .dout(n2792));
  jor  g02576(.dina(n2792), .dinb(asqrt[53] ), .dout(n2793));
  jnot g02577(.din(n2645), .dout(n2794));
  jand g02578(.dina(n2794), .dinb(n2793), .dout(n2795));
  jor  g02579(.dina(n2795), .dinb(n2756), .dout(n2796));
  jor  g02580(.dina(n2796), .dinb(asqrt[54] ), .dout(n2797));
  jand g02581(.dina(n2652), .dinb(n2797), .dout(n2798));
  jor  g02582(.dina(n2798), .dinb(n2755), .dout(n2799));
  jor  g02583(.dina(n2799), .dinb(asqrt[55] ), .dout(n2800));
  jnot g02584(.din(n2660), .dout(n2801));
  jand g02585(.dina(n2801), .dinb(n2800), .dout(n2802));
  jor  g02586(.dina(n2802), .dinb(n2754), .dout(n2803));
  jor  g02587(.dina(n2803), .dinb(asqrt[56] ), .dout(n2804));
  jnot g02588(.din(n2667), .dout(n2805));
  jand g02589(.dina(n2805), .dinb(n2804), .dout(n2806));
  jor  g02590(.dina(n2806), .dinb(n2753), .dout(n2807));
  jor  g02591(.dina(n2807), .dinb(asqrt[57] ), .dout(n2808));
  jand g02592(.dina(n2674), .dinb(n2808), .dout(n2809));
  jor  g02593(.dina(n2809), .dinb(n2752), .dout(n2810));
  jor  g02594(.dina(n2810), .dinb(asqrt[58] ), .dout(n2811));
  jand g02595(.dina(n2682), .dinb(n2811), .dout(n2812));
  jor  g02596(.dina(n2812), .dinb(n2751), .dout(n2813));
  jor  g02597(.dina(n2813), .dinb(asqrt[59] ), .dout(n2814));
  jnot g02598(.din(n2690), .dout(n2815));
  jand g02599(.dina(n2815), .dinb(n2814), .dout(n2816));
  jor  g02600(.dina(n2816), .dinb(n2750), .dout(n2817));
  jor  g02601(.dina(n2817), .dinb(asqrt[60] ), .dout(n2818));
  jand g02602(.dina(n2697), .dinb(n2818), .dout(n2819));
  jor  g02603(.dina(n2819), .dinb(n2749), .dout(n2820));
  jor  g02604(.dina(n2820), .dinb(asqrt[61] ), .dout(n2821));
  jand g02605(.dina(n2705), .dinb(n2821), .dout(n2822));
  jor  g02606(.dina(n2822), .dinb(n2748), .dout(n2823));
  jor  g02607(.dina(n2823), .dinb(asqrt[62] ), .dout(n2824));
  jand g02608(.dina(n2713), .dinb(n2824), .dout(n2825));
  jor  g02609(.dina(n2825), .dinb(n2747), .dout(n2826));
  jand g02610(.dina(n2826), .dinb(n2575), .dout(n2827));
  jand g02611(.dina(n2827), .dinb(n2469), .dout(n2828));
  jand g02612(.dina(n2828), .dinb(n2746), .dout(n2829));
  jor  g02613(.dina(n2829), .dinb(asqrt[63] ), .dout(n2830));
  jand g02614(.dina(n2728), .dinb(n2830), .dout(n2831));
  jand g02615(.dina(n2831), .dinb(n2744), .dout(n2833));
  jor  g02616(.dina(n2833), .dinb(n2743), .dout(n2834));
  jand g02617(.dina(n2834), .dinb(n2742), .dout(n2835));
  jand g02618(.dina(n2835), .dinb(n2740), .dout(n2836));
  jor  g02619(.dina(n2836), .dinb(n2739), .dout(n2837));
  jand g02620(.dina(n2837), .dinb(asqrt[46] ), .dout(n2838));
  jor  g02621(.dina(n2837), .dinb(asqrt[46] ), .dout(n2839));
  jand g02622(.dina(asqrt[44] ), .dinb(n2580), .dout(n2840));
  jand g02623(.dina(n2744), .dinb(asqrt[45] ), .dout(n2841));
  jand g02624(.dina(n2841), .dinb(n2727), .dout(n2842));
  jand g02625(.dina(n2842), .dinb(n2830), .dout(n2843));
  jor  g02626(.dina(n2843), .dinb(n2840), .dout(n2844));
  jxor g02627(.dina(n2844), .dinb(a[90] ), .dout(n2845));
  jnot g02628(.din(n2845), .dout(n2846));
  jand g02629(.dina(n2846), .dinb(n2839), .dout(n2847));
  jor  g02630(.dina(n2847), .dinb(n2838), .dout(n2848));
  jand g02631(.dina(n2848), .dinb(asqrt[47] ), .dout(n2849));
  jor  g02632(.dina(n2848), .dinb(asqrt[47] ), .dout(n2850));
  jxor g02633(.dina(n2583), .dinb(n2345), .dout(n2851));
  jand g02634(.dina(n2851), .dinb(asqrt[44] ), .dout(n2852));
  jxor g02635(.dina(n2852), .dinb(n2769), .dout(n2853));
  jand g02636(.dina(n2853), .dinb(n2850), .dout(n2854));
  jor  g02637(.dina(n2854), .dinb(n2849), .dout(n2855));
  jand g02638(.dina(n2855), .dinb(asqrt[48] ), .dout(n2856));
  jor  g02639(.dina(n2855), .dinb(asqrt[48] ), .dout(n2857));
  jxor g02640(.dina(n2591), .dinb(n2108), .dout(n2858));
  jand g02641(.dina(n2858), .dinb(asqrt[44] ), .dout(n2859));
  jxor g02642(.dina(n2859), .dinb(n2600), .dout(n2860));
  jnot g02643(.din(n2860), .dout(n2861));
  jand g02644(.dina(n2861), .dinb(n2857), .dout(n2862));
  jor  g02645(.dina(n2862), .dinb(n2856), .dout(n2863));
  jand g02646(.dina(n2863), .dinb(asqrt[49] ), .dout(n2864));
  jor  g02647(.dina(n2863), .dinb(asqrt[49] ), .dout(n2865));
  jxor g02648(.dina(n2602), .dinb(n1912), .dout(n2866));
  jand g02649(.dina(n2866), .dinb(asqrt[44] ), .dout(n2867));
  jxor g02650(.dina(n2867), .dinb(n2607), .dout(n2868));
  jand g02651(.dina(n2868), .dinb(n2865), .dout(n2869));
  jor  g02652(.dina(n2869), .dinb(n2864), .dout(n2870));
  jand g02653(.dina(n2870), .dinb(asqrt[50] ), .dout(n2871));
  jor  g02654(.dina(n2870), .dinb(asqrt[50] ), .dout(n2872));
  jxor g02655(.dina(n2610), .dinb(n1699), .dout(n2873));
  jand g02656(.dina(n2873), .dinb(asqrt[44] ), .dout(n2874));
  jxor g02657(.dina(n2874), .dinb(n2615), .dout(n2875));
  jnot g02658(.din(n2875), .dout(n2876));
  jand g02659(.dina(n2876), .dinb(n2872), .dout(n2877));
  jor  g02660(.dina(n2877), .dinb(n2871), .dout(n2878));
  jand g02661(.dina(n2878), .dinb(asqrt[51] ), .dout(n2879));
  jor  g02662(.dina(n2878), .dinb(asqrt[51] ), .dout(n2880));
  jxor g02663(.dina(n2617), .dinb(n1516), .dout(n2881));
  jand g02664(.dina(n2881), .dinb(asqrt[44] ), .dout(n2882));
  jxor g02665(.dina(n2882), .dinb(n2622), .dout(n2883));
  jand g02666(.dina(n2883), .dinb(n2880), .dout(n2884));
  jor  g02667(.dina(n2884), .dinb(n2879), .dout(n2885));
  jand g02668(.dina(n2885), .dinb(asqrt[52] ), .dout(n2886));
  jor  g02669(.dina(n2885), .dinb(asqrt[52] ), .dout(n2887));
  jxor g02670(.dina(n2625), .dinb(n1332), .dout(n2888));
  jand g02671(.dina(n2888), .dinb(asqrt[44] ), .dout(n2889));
  jxor g02672(.dina(n2889), .dinb(n2630), .dout(n2890));
  jnot g02673(.din(n2890), .dout(n2891));
  jand g02674(.dina(n2891), .dinb(n2887), .dout(n2892));
  jor  g02675(.dina(n2892), .dinb(n2886), .dout(n2893));
  jand g02676(.dina(n2893), .dinb(asqrt[53] ), .dout(n2894));
  jor  g02677(.dina(n2893), .dinb(asqrt[53] ), .dout(n2895));
  jxor g02678(.dina(n2632), .dinb(n1173), .dout(n2896));
  jand g02679(.dina(n2896), .dinb(asqrt[44] ), .dout(n2897));
  jxor g02680(.dina(n2897), .dinb(n2637), .dout(n2898));
  jand g02681(.dina(n2898), .dinb(n2895), .dout(n2899));
  jor  g02682(.dina(n2899), .dinb(n2894), .dout(n2900));
  jand g02683(.dina(n2900), .dinb(asqrt[54] ), .dout(n2901));
  jor  g02684(.dina(n2900), .dinb(asqrt[54] ), .dout(n2902));
  jxor g02685(.dina(n2640), .dinb(n1008), .dout(n2903));
  jand g02686(.dina(n2903), .dinb(asqrt[44] ), .dout(n2904));
  jxor g02687(.dina(n2904), .dinb(n2645), .dout(n2905));
  jnot g02688(.din(n2905), .dout(n2906));
  jand g02689(.dina(n2906), .dinb(n2902), .dout(n2907));
  jor  g02690(.dina(n2907), .dinb(n2901), .dout(n2908));
  jand g02691(.dina(n2908), .dinb(asqrt[55] ), .dout(n2909));
  jor  g02692(.dina(n2908), .dinb(asqrt[55] ), .dout(n2910));
  jxor g02693(.dina(n2647), .dinb(n884), .dout(n2911));
  jand g02694(.dina(n2911), .dinb(asqrt[44] ), .dout(n2912));
  jxor g02695(.dina(n2912), .dinb(n2652), .dout(n2913));
  jand g02696(.dina(n2913), .dinb(n2910), .dout(n2914));
  jor  g02697(.dina(n2914), .dinb(n2909), .dout(n2915));
  jand g02698(.dina(n2915), .dinb(asqrt[56] ), .dout(n2916));
  jor  g02699(.dina(n2915), .dinb(asqrt[56] ), .dout(n2917));
  jxor g02700(.dina(n2655), .dinb(n743), .dout(n2918));
  jand g02701(.dina(n2918), .dinb(asqrt[44] ), .dout(n2919));
  jxor g02702(.dina(n2919), .dinb(n2660), .dout(n2920));
  jnot g02703(.din(n2920), .dout(n2921));
  jand g02704(.dina(n2921), .dinb(n2917), .dout(n2922));
  jor  g02705(.dina(n2922), .dinb(n2916), .dout(n2923));
  jand g02706(.dina(n2923), .dinb(asqrt[57] ), .dout(n2924));
  jor  g02707(.dina(n2923), .dinb(asqrt[57] ), .dout(n2925));
  jxor g02708(.dina(n2662), .dinb(n635), .dout(n2926));
  jand g02709(.dina(n2926), .dinb(asqrt[44] ), .dout(n2927));
  jxor g02710(.dina(n2927), .dinb(n2667), .dout(n2928));
  jnot g02711(.din(n2928), .dout(n2929));
  jand g02712(.dina(n2929), .dinb(n2925), .dout(n2930));
  jor  g02713(.dina(n2930), .dinb(n2924), .dout(n2931));
  jand g02714(.dina(n2931), .dinb(asqrt[58] ), .dout(n2932));
  jor  g02715(.dina(n2931), .dinb(asqrt[58] ), .dout(n2933));
  jxor g02716(.dina(n2669), .dinb(n515), .dout(n2934));
  jand g02717(.dina(n2934), .dinb(asqrt[44] ), .dout(n2935));
  jxor g02718(.dina(n2935), .dinb(n2674), .dout(n2936));
  jand g02719(.dina(n2936), .dinb(n2933), .dout(n2937));
  jor  g02720(.dina(n2937), .dinb(n2932), .dout(n2938));
  jand g02721(.dina(n2938), .dinb(asqrt[59] ), .dout(n2939));
  jor  g02722(.dina(n2938), .dinb(asqrt[59] ), .dout(n2940));
  jxor g02723(.dina(n2677), .dinb(n443), .dout(n2941));
  jand g02724(.dina(n2941), .dinb(asqrt[44] ), .dout(n2942));
  jxor g02725(.dina(n2942), .dinb(n2682), .dout(n2943));
  jand g02726(.dina(n2943), .dinb(n2940), .dout(n2944));
  jor  g02727(.dina(n2944), .dinb(n2939), .dout(n2945));
  jand g02728(.dina(n2945), .dinb(asqrt[60] ), .dout(n2946));
  jor  g02729(.dina(n2945), .dinb(asqrt[60] ), .dout(n2947));
  jxor g02730(.dina(n2685), .dinb(n352), .dout(n2948));
  jand g02731(.dina(n2948), .dinb(asqrt[44] ), .dout(n2949));
  jxor g02732(.dina(n2949), .dinb(n2690), .dout(n2950));
  jnot g02733(.din(n2950), .dout(n2951));
  jand g02734(.dina(n2951), .dinb(n2947), .dout(n2952));
  jor  g02735(.dina(n2952), .dinb(n2946), .dout(n2953));
  jand g02736(.dina(n2953), .dinb(asqrt[61] ), .dout(n2954));
  jor  g02737(.dina(n2953), .dinb(asqrt[61] ), .dout(n2955));
  jxor g02738(.dina(n2692), .dinb(n294), .dout(n2956));
  jand g02739(.dina(n2956), .dinb(asqrt[44] ), .dout(n2957));
  jxor g02740(.dina(n2957), .dinb(n2697), .dout(n2958));
  jand g02741(.dina(n2958), .dinb(n2955), .dout(n2959));
  jor  g02742(.dina(n2959), .dinb(n2954), .dout(n2960));
  jand g02743(.dina(n2960), .dinb(asqrt[62] ), .dout(n2961));
  jor  g02744(.dina(n2960), .dinb(asqrt[62] ), .dout(n2962));
  jxor g02745(.dina(n2700), .dinb(n239), .dout(n2963));
  jand g02746(.dina(n2963), .dinb(asqrt[44] ), .dout(n2964));
  jxor g02747(.dina(n2964), .dinb(n2705), .dout(n2965));
  jand g02748(.dina(n2965), .dinb(n2962), .dout(n2966));
  jor  g02749(.dina(n2966), .dinb(n2961), .dout(n2967));
  jxor g02750(.dina(n2708), .dinb(n221), .dout(n2968));
  jand g02751(.dina(n2968), .dinb(asqrt[44] ), .dout(n2969));
  jxor g02752(.dina(n2969), .dinb(n2714), .dout(n2970));
  jnot g02753(.din(n2970), .dout(n2971));
  jor  g02754(.dina(n2971), .dinb(n2967), .dout(n2972));
  jnot g02755(.din(n2972), .dout(n2973));
  jand g02756(.dina(n2831), .dinb(n2716), .dout(n2974));
  jnot g02757(.din(n2974), .dout(n2975));
  jand g02758(.dina(n2720), .dinb(asqrt[63] ), .dout(n2976));
  jand g02759(.dina(n2976), .dinb(n2744), .dout(n2977));
  jand g02760(.dina(n2977), .dinb(n2975), .dout(n2978));
  jand g02761(.dina(n2730), .dinb(n2827), .dout(n2979));
  jnot g02762(.din(n2961), .dout(n2980));
  jnot g02763(.din(n2954), .dout(n2981));
  jnot g02764(.din(n2946), .dout(n2982));
  jnot g02765(.din(n2939), .dout(n2983));
  jnot g02766(.din(n2932), .dout(n2984));
  jnot g02767(.din(n2924), .dout(n2985));
  jnot g02768(.din(n2916), .dout(n2986));
  jnot g02769(.din(n2909), .dout(n2987));
  jnot g02770(.din(n2901), .dout(n2988));
  jnot g02771(.din(n2894), .dout(n2989));
  jnot g02772(.din(n2886), .dout(n2990));
  jnot g02773(.din(n2879), .dout(n2991));
  jnot g02774(.din(n2871), .dout(n2992));
  jnot g02775(.din(n2864), .dout(n2993));
  jnot g02776(.din(n2856), .dout(n2994));
  jnot g02777(.din(n2849), .dout(n2995));
  jnot g02778(.din(n2838), .dout(n2996));
  jnot g02779(.din(n2739), .dout(n2997));
  jor  g02780(.dina(n2833), .dinb(n2578), .dout(n2998));
  jnot g02781(.din(n2737), .dout(n2999));
  jand g02782(.dina(n2999), .dinb(n2998), .dout(n3000));
  jand g02783(.dina(n3000), .dinb(n2572), .dout(n3001));
  jor  g02784(.dina(n2833), .dinb(a[88] ), .dout(n3002));
  jand g02785(.dina(n3002), .dinb(a[89] ), .dout(n3003));
  jor  g02786(.dina(n2840), .dinb(n3003), .dout(n3004));
  jor  g02787(.dina(n3004), .dinb(n3001), .dout(n3005));
  jand g02788(.dina(n3005), .dinb(n2997), .dout(n3006));
  jand g02789(.dina(n3006), .dinb(n2345), .dout(n3007));
  jor  g02790(.dina(n2845), .dinb(n3007), .dout(n3008));
  jand g02791(.dina(n3008), .dinb(n2996), .dout(n3009));
  jand g02792(.dina(n3009), .dinb(n2108), .dout(n3010));
  jnot g02793(.din(n2853), .dout(n3011));
  jor  g02794(.dina(n3011), .dinb(n3010), .dout(n3012));
  jand g02795(.dina(n3012), .dinb(n2995), .dout(n3013));
  jand g02796(.dina(n3013), .dinb(n1912), .dout(n3014));
  jor  g02797(.dina(n2860), .dinb(n3014), .dout(n3015));
  jand g02798(.dina(n3015), .dinb(n2994), .dout(n3016));
  jand g02799(.dina(n3016), .dinb(n1699), .dout(n3017));
  jnot g02800(.din(n2868), .dout(n3018));
  jor  g02801(.dina(n3018), .dinb(n3017), .dout(n3019));
  jand g02802(.dina(n3019), .dinb(n2993), .dout(n3020));
  jand g02803(.dina(n3020), .dinb(n1516), .dout(n3021));
  jor  g02804(.dina(n2875), .dinb(n3021), .dout(n3022));
  jand g02805(.dina(n3022), .dinb(n2992), .dout(n3023));
  jand g02806(.dina(n3023), .dinb(n1332), .dout(n3024));
  jnot g02807(.din(n2883), .dout(n3025));
  jor  g02808(.dina(n3025), .dinb(n3024), .dout(n3026));
  jand g02809(.dina(n3026), .dinb(n2991), .dout(n3027));
  jand g02810(.dina(n3027), .dinb(n1173), .dout(n3028));
  jor  g02811(.dina(n2890), .dinb(n3028), .dout(n3029));
  jand g02812(.dina(n3029), .dinb(n2990), .dout(n3030));
  jand g02813(.dina(n3030), .dinb(n1008), .dout(n3031));
  jnot g02814(.din(n2898), .dout(n3032));
  jor  g02815(.dina(n3032), .dinb(n3031), .dout(n3033));
  jand g02816(.dina(n3033), .dinb(n2989), .dout(n3034));
  jand g02817(.dina(n3034), .dinb(n884), .dout(n3035));
  jor  g02818(.dina(n2905), .dinb(n3035), .dout(n3036));
  jand g02819(.dina(n3036), .dinb(n2988), .dout(n3037));
  jand g02820(.dina(n3037), .dinb(n743), .dout(n3038));
  jnot g02821(.din(n2913), .dout(n3039));
  jor  g02822(.dina(n3039), .dinb(n3038), .dout(n3040));
  jand g02823(.dina(n3040), .dinb(n2987), .dout(n3041));
  jand g02824(.dina(n3041), .dinb(n635), .dout(n3042));
  jor  g02825(.dina(n2920), .dinb(n3042), .dout(n3043));
  jand g02826(.dina(n3043), .dinb(n2986), .dout(n3044));
  jand g02827(.dina(n3044), .dinb(n515), .dout(n3045));
  jor  g02828(.dina(n2928), .dinb(n3045), .dout(n3046));
  jand g02829(.dina(n3046), .dinb(n2985), .dout(n3047));
  jand g02830(.dina(n3047), .dinb(n443), .dout(n3048));
  jnot g02831(.din(n2936), .dout(n3049));
  jor  g02832(.dina(n3049), .dinb(n3048), .dout(n3050));
  jand g02833(.dina(n3050), .dinb(n2984), .dout(n3051));
  jand g02834(.dina(n3051), .dinb(n352), .dout(n3052));
  jnot g02835(.din(n2943), .dout(n3053));
  jor  g02836(.dina(n3053), .dinb(n3052), .dout(n3054));
  jand g02837(.dina(n3054), .dinb(n2983), .dout(n3055));
  jand g02838(.dina(n3055), .dinb(n294), .dout(n3056));
  jor  g02839(.dina(n2950), .dinb(n3056), .dout(n3057));
  jand g02840(.dina(n3057), .dinb(n2982), .dout(n3058));
  jand g02841(.dina(n3058), .dinb(n239), .dout(n3059));
  jnot g02842(.din(n2958), .dout(n3060));
  jor  g02843(.dina(n3060), .dinb(n3059), .dout(n3061));
  jand g02844(.dina(n3061), .dinb(n2981), .dout(n3062));
  jand g02845(.dina(n3062), .dinb(n221), .dout(n3063));
  jnot g02846(.din(n2965), .dout(n3064));
  jor  g02847(.dina(n3064), .dinb(n3063), .dout(n3065));
  jand g02848(.dina(n3065), .dinb(n2980), .dout(n3066));
  jor  g02849(.dina(n2970), .dinb(n3066), .dout(n3067));
  jor  g02850(.dina(n3067), .dinb(n2717), .dout(n3068));
  jor  g02851(.dina(n3068), .dinb(n2979), .dout(n3069));
  jand g02852(.dina(n3069), .dinb(n218), .dout(n3070));
  jand g02853(.dina(n2833), .dinb(n2576), .dout(n3071));
  jor  g02854(.dina(n3071), .dinb(n3070), .dout(n3072));
  jor  g02855(.dina(n3072), .dinb(n2978), .dout(n3073));
  jor  g02856(.dina(n3073), .dinb(n2973), .dout(asqrt[43] ));
  jnot g02857(.din(a[84] ), .dout(n3075));
  jnot g02858(.din(a[85] ), .dout(n3076));
  jand g02859(.dina(n3076), .dinb(n3075), .dout(n3077));
  jand g02860(.dina(n3077), .dinb(n2734), .dout(n3078));
  jnot g02861(.din(n3078), .dout(n3079));
  jnot g02862(.din(n2978), .dout(n3080));
  jnot g02863(.din(n2979), .dout(n3081));
  jand g02864(.dina(n2971), .dinb(n2967), .dout(n3082));
  jand g02865(.dina(n3082), .dinb(n2744), .dout(n3083));
  jand g02866(.dina(n3083), .dinb(n3081), .dout(n3084));
  jor  g02867(.dina(n3084), .dinb(asqrt[63] ), .dout(n3085));
  jnot g02868(.din(n3071), .dout(n3086));
  jand g02869(.dina(n3086), .dinb(n3085), .dout(n3087));
  jand g02870(.dina(n3087), .dinb(n3080), .dout(n3088));
  jand g02871(.dina(n3088), .dinb(n2972), .dout(n3089));
  jor  g02872(.dina(n3089), .dinb(n2734), .dout(n3090));
  jand g02873(.dina(n3090), .dinb(n3079), .dout(n3091));
  jor  g02874(.dina(n3091), .dinb(n2833), .dout(n3092));
  jand g02875(.dina(n3091), .dinb(n2833), .dout(n3093));
  jor  g02876(.dina(n3089), .dinb(a[86] ), .dout(n3094));
  jand g02877(.dina(n3094), .dinb(a[87] ), .dout(n3095));
  jand g02878(.dina(asqrt[43] ), .dinb(n2736), .dout(n3096));
  jor  g02879(.dina(n3096), .dinb(n3095), .dout(n3097));
  jor  g02880(.dina(n3097), .dinb(n3093), .dout(n3098));
  jand g02881(.dina(n3098), .dinb(n3092), .dout(n3099));
  jor  g02882(.dina(n3099), .dinb(n2572), .dout(n3100));
  jand g02883(.dina(n3099), .dinb(n2572), .dout(n3101));
  jnot g02884(.din(n2736), .dout(n3102));
  jor  g02885(.dina(n3089), .dinb(n3102), .dout(n3103));
  jor  g02886(.dina(n2977), .dinb(n2973), .dout(n3104));
  jor  g02887(.dina(n3104), .dinb(n3070), .dout(n3105));
  jor  g02888(.dina(n3105), .dinb(n2833), .dout(n3106));
  jand g02889(.dina(n3106), .dinb(n3103), .dout(n3107));
  jxor g02890(.dina(n3107), .dinb(n2578), .dout(n3108));
  jor  g02891(.dina(n3108), .dinb(n3101), .dout(n3109));
  jand g02892(.dina(n3109), .dinb(n3100), .dout(n3110));
  jor  g02893(.dina(n3110), .dinb(n2345), .dout(n3111));
  jand g02894(.dina(n3110), .dinb(n2345), .dout(n3112));
  jxor g02895(.dina(n2738), .dinb(n2572), .dout(n3113));
  jor  g02896(.dina(n3113), .dinb(n3089), .dout(n3114));
  jxor g02897(.dina(n3114), .dinb(n2835), .dout(n3115));
  jor  g02898(.dina(n3115), .dinb(n3112), .dout(n3116));
  jand g02899(.dina(n3116), .dinb(n3111), .dout(n3117));
  jor  g02900(.dina(n3117), .dinb(n2108), .dout(n3118));
  jand g02901(.dina(n3117), .dinb(n2108), .dout(n3119));
  jxor g02902(.dina(n2837), .dinb(n2345), .dout(n3120));
  jor  g02903(.dina(n3120), .dinb(n3089), .dout(n3121));
  jxor g02904(.dina(n3121), .dinb(n2846), .dout(n3122));
  jor  g02905(.dina(n3122), .dinb(n3119), .dout(n3123));
  jand g02906(.dina(n3123), .dinb(n3118), .dout(n3124));
  jor  g02907(.dina(n3124), .dinb(n1912), .dout(n3125));
  jand g02908(.dina(n3124), .dinb(n1912), .dout(n3126));
  jxor g02909(.dina(n2848), .dinb(n2108), .dout(n3127));
  jor  g02910(.dina(n3127), .dinb(n3089), .dout(n3128));
  jxor g02911(.dina(n3128), .dinb(n3011), .dout(n3129));
  jnot g02912(.din(n3129), .dout(n3130));
  jor  g02913(.dina(n3130), .dinb(n3126), .dout(n3131));
  jand g02914(.dina(n3131), .dinb(n3125), .dout(n3132));
  jor  g02915(.dina(n3132), .dinb(n1699), .dout(n3133));
  jand g02916(.dina(n3132), .dinb(n1699), .dout(n3134));
  jxor g02917(.dina(n2855), .dinb(n1912), .dout(n3135));
  jor  g02918(.dina(n3135), .dinb(n3089), .dout(n3136));
  jxor g02919(.dina(n3136), .dinb(n2861), .dout(n3137));
  jor  g02920(.dina(n3137), .dinb(n3134), .dout(n3138));
  jand g02921(.dina(n3138), .dinb(n3133), .dout(n3139));
  jor  g02922(.dina(n3139), .dinb(n1516), .dout(n3140));
  jand g02923(.dina(n3139), .dinb(n1516), .dout(n3141));
  jxor g02924(.dina(n2863), .dinb(n1699), .dout(n3142));
  jor  g02925(.dina(n3142), .dinb(n3089), .dout(n3143));
  jxor g02926(.dina(n3143), .dinb(n3018), .dout(n3144));
  jnot g02927(.din(n3144), .dout(n3145));
  jor  g02928(.dina(n3145), .dinb(n3141), .dout(n3146));
  jand g02929(.dina(n3146), .dinb(n3140), .dout(n3147));
  jor  g02930(.dina(n3147), .dinb(n1332), .dout(n3148));
  jand g02931(.dina(n3147), .dinb(n1332), .dout(n3149));
  jxor g02932(.dina(n2870), .dinb(n1516), .dout(n3150));
  jor  g02933(.dina(n3150), .dinb(n3089), .dout(n3151));
  jxor g02934(.dina(n3151), .dinb(n2876), .dout(n3152));
  jor  g02935(.dina(n3152), .dinb(n3149), .dout(n3153));
  jand g02936(.dina(n3153), .dinb(n3148), .dout(n3154));
  jor  g02937(.dina(n3154), .dinb(n1173), .dout(n3155));
  jand g02938(.dina(n3154), .dinb(n1173), .dout(n3156));
  jxor g02939(.dina(n2878), .dinb(n1332), .dout(n3157));
  jor  g02940(.dina(n3157), .dinb(n3089), .dout(n3158));
  jxor g02941(.dina(n3158), .dinb(n3025), .dout(n3159));
  jnot g02942(.din(n3159), .dout(n3160));
  jor  g02943(.dina(n3160), .dinb(n3156), .dout(n3161));
  jand g02944(.dina(n3161), .dinb(n3155), .dout(n3162));
  jor  g02945(.dina(n3162), .dinb(n1008), .dout(n3163));
  jand g02946(.dina(n3162), .dinb(n1008), .dout(n3164));
  jxor g02947(.dina(n2885), .dinb(n1173), .dout(n3165));
  jor  g02948(.dina(n3165), .dinb(n3089), .dout(n3166));
  jxor g02949(.dina(n3166), .dinb(n2891), .dout(n3167));
  jor  g02950(.dina(n3167), .dinb(n3164), .dout(n3168));
  jand g02951(.dina(n3168), .dinb(n3163), .dout(n3169));
  jor  g02952(.dina(n3169), .dinb(n884), .dout(n3170));
  jand g02953(.dina(n3169), .dinb(n884), .dout(n3171));
  jxor g02954(.dina(n2893), .dinb(n1008), .dout(n3172));
  jor  g02955(.dina(n3172), .dinb(n3089), .dout(n3173));
  jxor g02956(.dina(n3173), .dinb(n3032), .dout(n3174));
  jnot g02957(.din(n3174), .dout(n3175));
  jor  g02958(.dina(n3175), .dinb(n3171), .dout(n3176));
  jand g02959(.dina(n3176), .dinb(n3170), .dout(n3177));
  jor  g02960(.dina(n3177), .dinb(n743), .dout(n3178));
  jand g02961(.dina(n3177), .dinb(n743), .dout(n3179));
  jxor g02962(.dina(n2900), .dinb(n884), .dout(n3180));
  jor  g02963(.dina(n3180), .dinb(n3089), .dout(n3181));
  jxor g02964(.dina(n3181), .dinb(n2906), .dout(n3182));
  jor  g02965(.dina(n3182), .dinb(n3179), .dout(n3183));
  jand g02966(.dina(n3183), .dinb(n3178), .dout(n3184));
  jor  g02967(.dina(n3184), .dinb(n635), .dout(n3185));
  jand g02968(.dina(n3184), .dinb(n635), .dout(n3186));
  jxor g02969(.dina(n2908), .dinb(n743), .dout(n3187));
  jor  g02970(.dina(n3187), .dinb(n3089), .dout(n3188));
  jxor g02971(.dina(n3188), .dinb(n3039), .dout(n3189));
  jnot g02972(.din(n3189), .dout(n3190));
  jor  g02973(.dina(n3190), .dinb(n3186), .dout(n3191));
  jand g02974(.dina(n3191), .dinb(n3185), .dout(n3192));
  jor  g02975(.dina(n3192), .dinb(n515), .dout(n3193));
  jand g02976(.dina(n3192), .dinb(n515), .dout(n3194));
  jxor g02977(.dina(n2915), .dinb(n635), .dout(n3195));
  jor  g02978(.dina(n3195), .dinb(n3089), .dout(n3196));
  jxor g02979(.dina(n3196), .dinb(n2921), .dout(n3197));
  jor  g02980(.dina(n3197), .dinb(n3194), .dout(n3198));
  jand g02981(.dina(n3198), .dinb(n3193), .dout(n3199));
  jor  g02982(.dina(n3199), .dinb(n443), .dout(n3200));
  jand g02983(.dina(n3199), .dinb(n443), .dout(n3201));
  jxor g02984(.dina(n2923), .dinb(n515), .dout(n3202));
  jor  g02985(.dina(n3202), .dinb(n3089), .dout(n3203));
  jxor g02986(.dina(n3203), .dinb(n2929), .dout(n3204));
  jor  g02987(.dina(n3204), .dinb(n3201), .dout(n3205));
  jand g02988(.dina(n3205), .dinb(n3200), .dout(n3206));
  jor  g02989(.dina(n3206), .dinb(n352), .dout(n3207));
  jand g02990(.dina(n3206), .dinb(n352), .dout(n3208));
  jxor g02991(.dina(n2931), .dinb(n443), .dout(n3209));
  jor  g02992(.dina(n3209), .dinb(n3089), .dout(n3210));
  jxor g02993(.dina(n3210), .dinb(n3049), .dout(n3211));
  jnot g02994(.din(n3211), .dout(n3212));
  jor  g02995(.dina(n3212), .dinb(n3208), .dout(n3213));
  jand g02996(.dina(n3213), .dinb(n3207), .dout(n3214));
  jor  g02997(.dina(n3214), .dinb(n294), .dout(n3215));
  jand g02998(.dina(n3214), .dinb(n294), .dout(n3216));
  jxor g02999(.dina(n2938), .dinb(n352), .dout(n3217));
  jor  g03000(.dina(n3217), .dinb(n3089), .dout(n3218));
  jxor g03001(.dina(n3218), .dinb(n3053), .dout(n3219));
  jnot g03002(.din(n3219), .dout(n3220));
  jor  g03003(.dina(n3220), .dinb(n3216), .dout(n3221));
  jand g03004(.dina(n3221), .dinb(n3215), .dout(n3222));
  jor  g03005(.dina(n3222), .dinb(n239), .dout(n3223));
  jand g03006(.dina(n3222), .dinb(n239), .dout(n3224));
  jxor g03007(.dina(n2945), .dinb(n294), .dout(n3225));
  jor  g03008(.dina(n3225), .dinb(n3089), .dout(n3226));
  jxor g03009(.dina(n3226), .dinb(n2951), .dout(n3227));
  jor  g03010(.dina(n3227), .dinb(n3224), .dout(n3228));
  jand g03011(.dina(n3228), .dinb(n3223), .dout(n3229));
  jor  g03012(.dina(n3229), .dinb(n221), .dout(n3230));
  jand g03013(.dina(n3229), .dinb(n221), .dout(n3231));
  jxor g03014(.dina(n2953), .dinb(n239), .dout(n3232));
  jor  g03015(.dina(n3232), .dinb(n3089), .dout(n3233));
  jxor g03016(.dina(n3233), .dinb(n3060), .dout(n3234));
  jnot g03017(.din(n3234), .dout(n3235));
  jor  g03018(.dina(n3235), .dinb(n3231), .dout(n3236));
  jand g03019(.dina(n3236), .dinb(n3230), .dout(n3237));
  jxor g03020(.dina(n2960), .dinb(n221), .dout(n3238));
  jor  g03021(.dina(n3238), .dinb(n3089), .dout(n3239));
  jxor g03022(.dina(n3239), .dinb(n2965), .dout(n3240));
  jand g03023(.dina(n3240), .dinb(n3237), .dout(n3241));
  jand g03024(.dina(n3088), .dinb(n3066), .dout(n3242));
  jand g03025(.dina(n3067), .dinb(asqrt[63] ), .dout(n3243));
  jand g03026(.dina(n3243), .dinb(n2972), .dout(n3244));
  jnot g03027(.din(n3244), .dout(n3245));
  jor  g03028(.dina(n3245), .dinb(n3242), .dout(n3246));
  jnot g03029(.din(n3246), .dout(n3247));
  jor  g03030(.dina(n3240), .dinb(n3237), .dout(n3248));
  jand g03031(.dina(n3073), .dinb(n3082), .dout(n3249));
  jor  g03032(.dina(n3249), .dinb(n2973), .dout(n3250));
  jor  g03033(.dina(n3250), .dinb(n3248), .dout(n3251));
  jand g03034(.dina(n3251), .dinb(n218), .dout(n3252));
  jand g03035(.dina(n3089), .dinb(n2970), .dout(n3253));
  jor  g03036(.dina(n3253), .dinb(n3252), .dout(n3254));
  jor  g03037(.dina(n3254), .dinb(n3247), .dout(n3255));
  jor  g03038(.dina(n3255), .dinb(n3241), .dout(asqrt[42] ));
  jand g03039(.dina(asqrt[42] ), .dinb(a[84] ), .dout(n3257));
  jnot g03040(.din(a[82] ), .dout(n3258));
  jnot g03041(.din(a[83] ), .dout(n3259));
  jand g03042(.dina(n3259), .dinb(n3258), .dout(n3260));
  jand g03043(.dina(n3260), .dinb(n3075), .dout(n3261));
  jor  g03044(.dina(n3261), .dinb(n3257), .dout(n3262));
  jand g03045(.dina(n3262), .dinb(asqrt[43] ), .dout(n3263));
  jor  g03046(.dina(n3262), .dinb(asqrt[43] ), .dout(n3264));
  jand g03047(.dina(asqrt[42] ), .dinb(n3075), .dout(n3265));
  jor  g03048(.dina(n3265), .dinb(n3076), .dout(n3266));
  jnot g03049(.din(n3077), .dout(n3267));
  jnot g03050(.din(n3241), .dout(n3268));
  jnot g03051(.din(n3230), .dout(n3269));
  jnot g03052(.din(n3223), .dout(n3270));
  jnot g03053(.din(n3215), .dout(n3271));
  jnot g03054(.din(n3207), .dout(n3272));
  jnot g03055(.din(n3200), .dout(n3273));
  jnot g03056(.din(n3193), .dout(n3274));
  jnot g03057(.din(n3185), .dout(n3275));
  jnot g03058(.din(n3178), .dout(n3276));
  jnot g03059(.din(n3170), .dout(n3277));
  jnot g03060(.din(n3163), .dout(n3278));
  jnot g03061(.din(n3155), .dout(n3279));
  jnot g03062(.din(n3148), .dout(n3280));
  jnot g03063(.din(n3140), .dout(n3281));
  jnot g03064(.din(n3133), .dout(n3282));
  jnot g03065(.din(n3125), .dout(n3283));
  jnot g03066(.din(n3118), .dout(n3284));
  jnot g03067(.din(n3111), .dout(n3285));
  jnot g03068(.din(n3100), .dout(n3286));
  jnot g03069(.din(n3092), .dout(n3287));
  jand g03070(.dina(asqrt[43] ), .dinb(a[86] ), .dout(n3288));
  jor  g03071(.dina(n3288), .dinb(n3078), .dout(n3289));
  jor  g03072(.dina(n3289), .dinb(asqrt[44] ), .dout(n3290));
  jand g03073(.dina(asqrt[43] ), .dinb(n2734), .dout(n3291));
  jor  g03074(.dina(n3291), .dinb(n2735), .dout(n3292));
  jand g03075(.dina(n3103), .dinb(n3292), .dout(n3293));
  jand g03076(.dina(n3293), .dinb(n3290), .dout(n3294));
  jor  g03077(.dina(n3294), .dinb(n3287), .dout(n3295));
  jor  g03078(.dina(n3295), .dinb(asqrt[45] ), .dout(n3296));
  jnot g03079(.din(n3108), .dout(n3297));
  jand g03080(.dina(n3297), .dinb(n3296), .dout(n3298));
  jor  g03081(.dina(n3298), .dinb(n3286), .dout(n3299));
  jor  g03082(.dina(n3299), .dinb(asqrt[46] ), .dout(n3300));
  jnot g03083(.din(n3115), .dout(n3301));
  jand g03084(.dina(n3301), .dinb(n3300), .dout(n3302));
  jor  g03085(.dina(n3302), .dinb(n3285), .dout(n3303));
  jor  g03086(.dina(n3303), .dinb(asqrt[47] ), .dout(n3304));
  jnot g03087(.din(n3122), .dout(n3305));
  jand g03088(.dina(n3305), .dinb(n3304), .dout(n3306));
  jor  g03089(.dina(n3306), .dinb(n3284), .dout(n3307));
  jor  g03090(.dina(n3307), .dinb(asqrt[48] ), .dout(n3308));
  jand g03091(.dina(n3129), .dinb(n3308), .dout(n3309));
  jor  g03092(.dina(n3309), .dinb(n3283), .dout(n3310));
  jor  g03093(.dina(n3310), .dinb(asqrt[49] ), .dout(n3311));
  jnot g03094(.din(n3137), .dout(n3312));
  jand g03095(.dina(n3312), .dinb(n3311), .dout(n3313));
  jor  g03096(.dina(n3313), .dinb(n3282), .dout(n3314));
  jor  g03097(.dina(n3314), .dinb(asqrt[50] ), .dout(n3315));
  jand g03098(.dina(n3144), .dinb(n3315), .dout(n3316));
  jor  g03099(.dina(n3316), .dinb(n3281), .dout(n3317));
  jor  g03100(.dina(n3317), .dinb(asqrt[51] ), .dout(n3318));
  jnot g03101(.din(n3152), .dout(n3319));
  jand g03102(.dina(n3319), .dinb(n3318), .dout(n3320));
  jor  g03103(.dina(n3320), .dinb(n3280), .dout(n3321));
  jor  g03104(.dina(n3321), .dinb(asqrt[52] ), .dout(n3322));
  jand g03105(.dina(n3159), .dinb(n3322), .dout(n3323));
  jor  g03106(.dina(n3323), .dinb(n3279), .dout(n3324));
  jor  g03107(.dina(n3324), .dinb(asqrt[53] ), .dout(n3325));
  jnot g03108(.din(n3167), .dout(n3326));
  jand g03109(.dina(n3326), .dinb(n3325), .dout(n3327));
  jor  g03110(.dina(n3327), .dinb(n3278), .dout(n3328));
  jor  g03111(.dina(n3328), .dinb(asqrt[54] ), .dout(n3329));
  jand g03112(.dina(n3174), .dinb(n3329), .dout(n3330));
  jor  g03113(.dina(n3330), .dinb(n3277), .dout(n3331));
  jor  g03114(.dina(n3331), .dinb(asqrt[55] ), .dout(n3332));
  jnot g03115(.din(n3182), .dout(n3333));
  jand g03116(.dina(n3333), .dinb(n3332), .dout(n3334));
  jor  g03117(.dina(n3334), .dinb(n3276), .dout(n3335));
  jor  g03118(.dina(n3335), .dinb(asqrt[56] ), .dout(n3336));
  jand g03119(.dina(n3189), .dinb(n3336), .dout(n3337));
  jor  g03120(.dina(n3337), .dinb(n3275), .dout(n3338));
  jor  g03121(.dina(n3338), .dinb(asqrt[57] ), .dout(n3339));
  jnot g03122(.din(n3197), .dout(n3340));
  jand g03123(.dina(n3340), .dinb(n3339), .dout(n3341));
  jor  g03124(.dina(n3341), .dinb(n3274), .dout(n3342));
  jor  g03125(.dina(n3342), .dinb(asqrt[58] ), .dout(n3343));
  jnot g03126(.din(n3204), .dout(n3344));
  jand g03127(.dina(n3344), .dinb(n3343), .dout(n3345));
  jor  g03128(.dina(n3345), .dinb(n3273), .dout(n3346));
  jor  g03129(.dina(n3346), .dinb(asqrt[59] ), .dout(n3347));
  jand g03130(.dina(n3211), .dinb(n3347), .dout(n3348));
  jor  g03131(.dina(n3348), .dinb(n3272), .dout(n3349));
  jor  g03132(.dina(n3349), .dinb(asqrt[60] ), .dout(n3350));
  jand g03133(.dina(n3219), .dinb(n3350), .dout(n3351));
  jor  g03134(.dina(n3351), .dinb(n3271), .dout(n3352));
  jor  g03135(.dina(n3352), .dinb(asqrt[61] ), .dout(n3353));
  jnot g03136(.din(n3227), .dout(n3354));
  jand g03137(.dina(n3354), .dinb(n3353), .dout(n3355));
  jor  g03138(.dina(n3355), .dinb(n3270), .dout(n3356));
  jor  g03139(.dina(n3356), .dinb(asqrt[62] ), .dout(n3357));
  jand g03140(.dina(n3234), .dinb(n3357), .dout(n3358));
  jor  g03141(.dina(n3358), .dinb(n3269), .dout(n3359));
  jnot g03142(.din(n3240), .dout(n3360));
  jand g03143(.dina(n3360), .dinb(n3359), .dout(n3361));
  jnot g03144(.din(n3250), .dout(n3362));
  jand g03145(.dina(n3362), .dinb(n3361), .dout(n3363));
  jor  g03146(.dina(n3363), .dinb(asqrt[63] ), .dout(n3364));
  jnot g03147(.din(n3253), .dout(n3365));
  jand g03148(.dina(n3365), .dinb(n3364), .dout(n3366));
  jand g03149(.dina(n3366), .dinb(n3246), .dout(n3367));
  jand g03150(.dina(n3367), .dinb(n3268), .dout(n3368));
  jor  g03151(.dina(n3368), .dinb(n3267), .dout(n3369));
  jand g03152(.dina(n3369), .dinb(n3266), .dout(n3370));
  jand g03153(.dina(n3370), .dinb(n3264), .dout(n3371));
  jor  g03154(.dina(n3371), .dinb(n3263), .dout(n3372));
  jand g03155(.dina(n3372), .dinb(asqrt[44] ), .dout(n3373));
  jor  g03156(.dina(n3372), .dinb(asqrt[44] ), .dout(n3374));
  jand g03157(.dina(asqrt[42] ), .dinb(n3077), .dout(n3375));
  jand g03158(.dina(n3268), .dinb(asqrt[43] ), .dout(n3376));
  jand g03159(.dina(n3376), .dinb(n3245), .dout(n3377));
  jand g03160(.dina(n3377), .dinb(n3364), .dout(n3378));
  jor  g03161(.dina(n3378), .dinb(n3375), .dout(n3379));
  jxor g03162(.dina(n3379), .dinb(a[86] ), .dout(n3380));
  jnot g03163(.din(n3380), .dout(n3381));
  jand g03164(.dina(n3381), .dinb(n3374), .dout(n3382));
  jor  g03165(.dina(n3382), .dinb(n3373), .dout(n3383));
  jand g03166(.dina(n3383), .dinb(asqrt[45] ), .dout(n3384));
  jor  g03167(.dina(n3383), .dinb(asqrt[45] ), .dout(n3385));
  jxor g03168(.dina(n3091), .dinb(n2833), .dout(n3386));
  jand g03169(.dina(n3386), .dinb(asqrt[42] ), .dout(n3387));
  jxor g03170(.dina(n3387), .dinb(n3293), .dout(n3388));
  jand g03171(.dina(n3388), .dinb(n3385), .dout(n3389));
  jor  g03172(.dina(n3389), .dinb(n3384), .dout(n3390));
  jand g03173(.dina(n3390), .dinb(asqrt[46] ), .dout(n3391));
  jor  g03174(.dina(n3390), .dinb(asqrt[46] ), .dout(n3392));
  jxor g03175(.dina(n3099), .dinb(n2572), .dout(n3393));
  jand g03176(.dina(n3393), .dinb(asqrt[42] ), .dout(n3394));
  jxor g03177(.dina(n3394), .dinb(n3297), .dout(n3395));
  jand g03178(.dina(n3395), .dinb(n3392), .dout(n3396));
  jor  g03179(.dina(n3396), .dinb(n3391), .dout(n3397));
  jand g03180(.dina(n3397), .dinb(asqrt[47] ), .dout(n3398));
  jor  g03181(.dina(n3397), .dinb(asqrt[47] ), .dout(n3399));
  jxor g03182(.dina(n3110), .dinb(n2345), .dout(n3400));
  jand g03183(.dina(n3400), .dinb(asqrt[42] ), .dout(n3401));
  jxor g03184(.dina(n3401), .dinb(n3115), .dout(n3402));
  jnot g03185(.din(n3402), .dout(n3403));
  jand g03186(.dina(n3403), .dinb(n3399), .dout(n3404));
  jor  g03187(.dina(n3404), .dinb(n3398), .dout(n3405));
  jand g03188(.dina(n3405), .dinb(asqrt[48] ), .dout(n3406));
  jor  g03189(.dina(n3405), .dinb(asqrt[48] ), .dout(n3407));
  jxor g03190(.dina(n3117), .dinb(n2108), .dout(n3408));
  jand g03191(.dina(n3408), .dinb(asqrt[42] ), .dout(n3409));
  jxor g03192(.dina(n3409), .dinb(n3122), .dout(n3410));
  jnot g03193(.din(n3410), .dout(n3411));
  jand g03194(.dina(n3411), .dinb(n3407), .dout(n3412));
  jor  g03195(.dina(n3412), .dinb(n3406), .dout(n3413));
  jand g03196(.dina(n3413), .dinb(asqrt[49] ), .dout(n3414));
  jor  g03197(.dina(n3413), .dinb(asqrt[49] ), .dout(n3415));
  jxor g03198(.dina(n3124), .dinb(n1912), .dout(n3416));
  jand g03199(.dina(n3416), .dinb(asqrt[42] ), .dout(n3417));
  jxor g03200(.dina(n3417), .dinb(n3129), .dout(n3418));
  jand g03201(.dina(n3418), .dinb(n3415), .dout(n3419));
  jor  g03202(.dina(n3419), .dinb(n3414), .dout(n3420));
  jand g03203(.dina(n3420), .dinb(asqrt[50] ), .dout(n3421));
  jor  g03204(.dina(n3420), .dinb(asqrt[50] ), .dout(n3422));
  jxor g03205(.dina(n3132), .dinb(n1699), .dout(n3423));
  jand g03206(.dina(n3423), .dinb(asqrt[42] ), .dout(n3424));
  jxor g03207(.dina(n3424), .dinb(n3137), .dout(n3425));
  jnot g03208(.din(n3425), .dout(n3426));
  jand g03209(.dina(n3426), .dinb(n3422), .dout(n3427));
  jor  g03210(.dina(n3427), .dinb(n3421), .dout(n3428));
  jand g03211(.dina(n3428), .dinb(asqrt[51] ), .dout(n3429));
  jor  g03212(.dina(n3428), .dinb(asqrt[51] ), .dout(n3430));
  jxor g03213(.dina(n3139), .dinb(n1516), .dout(n3431));
  jand g03214(.dina(n3431), .dinb(asqrt[42] ), .dout(n3432));
  jxor g03215(.dina(n3432), .dinb(n3144), .dout(n3433));
  jand g03216(.dina(n3433), .dinb(n3430), .dout(n3434));
  jor  g03217(.dina(n3434), .dinb(n3429), .dout(n3435));
  jand g03218(.dina(n3435), .dinb(asqrt[52] ), .dout(n3436));
  jor  g03219(.dina(n3435), .dinb(asqrt[52] ), .dout(n3437));
  jxor g03220(.dina(n3147), .dinb(n1332), .dout(n3438));
  jand g03221(.dina(n3438), .dinb(asqrt[42] ), .dout(n3439));
  jxor g03222(.dina(n3439), .dinb(n3152), .dout(n3440));
  jnot g03223(.din(n3440), .dout(n3441));
  jand g03224(.dina(n3441), .dinb(n3437), .dout(n3442));
  jor  g03225(.dina(n3442), .dinb(n3436), .dout(n3443));
  jand g03226(.dina(n3443), .dinb(asqrt[53] ), .dout(n3444));
  jor  g03227(.dina(n3443), .dinb(asqrt[53] ), .dout(n3445));
  jxor g03228(.dina(n3154), .dinb(n1173), .dout(n3446));
  jand g03229(.dina(n3446), .dinb(asqrt[42] ), .dout(n3447));
  jxor g03230(.dina(n3447), .dinb(n3159), .dout(n3448));
  jand g03231(.dina(n3448), .dinb(n3445), .dout(n3449));
  jor  g03232(.dina(n3449), .dinb(n3444), .dout(n3450));
  jand g03233(.dina(n3450), .dinb(asqrt[54] ), .dout(n3451));
  jor  g03234(.dina(n3450), .dinb(asqrt[54] ), .dout(n3452));
  jxor g03235(.dina(n3162), .dinb(n1008), .dout(n3453));
  jand g03236(.dina(n3453), .dinb(asqrt[42] ), .dout(n3454));
  jxor g03237(.dina(n3454), .dinb(n3167), .dout(n3455));
  jnot g03238(.din(n3455), .dout(n3456));
  jand g03239(.dina(n3456), .dinb(n3452), .dout(n3457));
  jor  g03240(.dina(n3457), .dinb(n3451), .dout(n3458));
  jand g03241(.dina(n3458), .dinb(asqrt[55] ), .dout(n3459));
  jor  g03242(.dina(n3458), .dinb(asqrt[55] ), .dout(n3460));
  jxor g03243(.dina(n3169), .dinb(n884), .dout(n3461));
  jand g03244(.dina(n3461), .dinb(asqrt[42] ), .dout(n3462));
  jxor g03245(.dina(n3462), .dinb(n3174), .dout(n3463));
  jand g03246(.dina(n3463), .dinb(n3460), .dout(n3464));
  jor  g03247(.dina(n3464), .dinb(n3459), .dout(n3465));
  jand g03248(.dina(n3465), .dinb(asqrt[56] ), .dout(n3466));
  jor  g03249(.dina(n3465), .dinb(asqrt[56] ), .dout(n3467));
  jxor g03250(.dina(n3177), .dinb(n743), .dout(n3468));
  jand g03251(.dina(n3468), .dinb(asqrt[42] ), .dout(n3469));
  jxor g03252(.dina(n3469), .dinb(n3182), .dout(n3470));
  jnot g03253(.din(n3470), .dout(n3471));
  jand g03254(.dina(n3471), .dinb(n3467), .dout(n3472));
  jor  g03255(.dina(n3472), .dinb(n3466), .dout(n3473));
  jand g03256(.dina(n3473), .dinb(asqrt[57] ), .dout(n3474));
  jor  g03257(.dina(n3473), .dinb(asqrt[57] ), .dout(n3475));
  jxor g03258(.dina(n3184), .dinb(n635), .dout(n3476));
  jand g03259(.dina(n3476), .dinb(asqrt[42] ), .dout(n3477));
  jxor g03260(.dina(n3477), .dinb(n3189), .dout(n3478));
  jand g03261(.dina(n3478), .dinb(n3475), .dout(n3479));
  jor  g03262(.dina(n3479), .dinb(n3474), .dout(n3480));
  jand g03263(.dina(n3480), .dinb(asqrt[58] ), .dout(n3481));
  jor  g03264(.dina(n3480), .dinb(asqrt[58] ), .dout(n3482));
  jxor g03265(.dina(n3192), .dinb(n515), .dout(n3483));
  jand g03266(.dina(n3483), .dinb(asqrt[42] ), .dout(n3484));
  jxor g03267(.dina(n3484), .dinb(n3197), .dout(n3485));
  jnot g03268(.din(n3485), .dout(n3486));
  jand g03269(.dina(n3486), .dinb(n3482), .dout(n3487));
  jor  g03270(.dina(n3487), .dinb(n3481), .dout(n3488));
  jand g03271(.dina(n3488), .dinb(asqrt[59] ), .dout(n3489));
  jor  g03272(.dina(n3488), .dinb(asqrt[59] ), .dout(n3490));
  jxor g03273(.dina(n3199), .dinb(n443), .dout(n3491));
  jand g03274(.dina(n3491), .dinb(asqrt[42] ), .dout(n3492));
  jxor g03275(.dina(n3492), .dinb(n3204), .dout(n3493));
  jnot g03276(.din(n3493), .dout(n3494));
  jand g03277(.dina(n3494), .dinb(n3490), .dout(n3495));
  jor  g03278(.dina(n3495), .dinb(n3489), .dout(n3496));
  jand g03279(.dina(n3496), .dinb(asqrt[60] ), .dout(n3497));
  jor  g03280(.dina(n3496), .dinb(asqrt[60] ), .dout(n3498));
  jxor g03281(.dina(n3206), .dinb(n352), .dout(n3499));
  jand g03282(.dina(n3499), .dinb(asqrt[42] ), .dout(n3500));
  jxor g03283(.dina(n3500), .dinb(n3211), .dout(n3501));
  jand g03284(.dina(n3501), .dinb(n3498), .dout(n3502));
  jor  g03285(.dina(n3502), .dinb(n3497), .dout(n3503));
  jand g03286(.dina(n3503), .dinb(asqrt[61] ), .dout(n3504));
  jor  g03287(.dina(n3503), .dinb(asqrt[61] ), .dout(n3505));
  jxor g03288(.dina(n3214), .dinb(n294), .dout(n3506));
  jand g03289(.dina(n3506), .dinb(asqrt[42] ), .dout(n3507));
  jxor g03290(.dina(n3507), .dinb(n3219), .dout(n3508));
  jand g03291(.dina(n3508), .dinb(n3505), .dout(n3509));
  jor  g03292(.dina(n3509), .dinb(n3504), .dout(n3510));
  jand g03293(.dina(n3510), .dinb(asqrt[62] ), .dout(n3511));
  jor  g03294(.dina(n3510), .dinb(asqrt[62] ), .dout(n3512));
  jxor g03295(.dina(n3222), .dinb(n239), .dout(n3513));
  jand g03296(.dina(n3513), .dinb(asqrt[42] ), .dout(n3514));
  jxor g03297(.dina(n3514), .dinb(n3227), .dout(n3515));
  jnot g03298(.din(n3515), .dout(n3516));
  jand g03299(.dina(n3516), .dinb(n3512), .dout(n3517));
  jor  g03300(.dina(n3517), .dinb(n3511), .dout(n3518));
  jxor g03301(.dina(n3229), .dinb(n221), .dout(n3519));
  jand g03302(.dina(n3519), .dinb(asqrt[42] ), .dout(n3520));
  jxor g03303(.dina(n3520), .dinb(n3235), .dout(n3521));
  jnot g03304(.din(n3521), .dout(n3522));
  jor  g03305(.dina(n3522), .dinb(n3518), .dout(n3523));
  jnot g03306(.din(n3523), .dout(n3524));
  jnot g03307(.din(n3511), .dout(n3526));
  jnot g03308(.din(n3504), .dout(n3527));
  jnot g03309(.din(n3497), .dout(n3528));
  jnot g03310(.din(n3489), .dout(n3529));
  jnot g03311(.din(n3481), .dout(n3530));
  jnot g03312(.din(n3474), .dout(n3531));
  jnot g03313(.din(n3466), .dout(n3532));
  jnot g03314(.din(n3459), .dout(n3533));
  jnot g03315(.din(n3451), .dout(n3534));
  jnot g03316(.din(n3444), .dout(n3535));
  jnot g03317(.din(n3436), .dout(n3536));
  jnot g03318(.din(n3429), .dout(n3537));
  jnot g03319(.din(n3421), .dout(n3538));
  jnot g03320(.din(n3414), .dout(n3539));
  jnot g03321(.din(n3406), .dout(n3540));
  jnot g03322(.din(n3398), .dout(n3541));
  jnot g03323(.din(n3391), .dout(n3542));
  jnot g03324(.din(n3384), .dout(n3543));
  jnot g03325(.din(n3373), .dout(n3544));
  jnot g03326(.din(n3263), .dout(n3545));
  jor  g03327(.dina(n3368), .dinb(n3075), .dout(n3546));
  jnot g03328(.din(n3261), .dout(n3547));
  jand g03329(.dina(n3547), .dinb(n3546), .dout(n3548));
  jand g03330(.dina(n3548), .dinb(n3089), .dout(n3549));
  jor  g03331(.dina(n3368), .dinb(a[84] ), .dout(n3550));
  jand g03332(.dina(n3550), .dinb(a[85] ), .dout(n3551));
  jor  g03333(.dina(n3375), .dinb(n3551), .dout(n3552));
  jor  g03334(.dina(n3552), .dinb(n3549), .dout(n3553));
  jand g03335(.dina(n3553), .dinb(n3545), .dout(n3554));
  jand g03336(.dina(n3554), .dinb(n2833), .dout(n3555));
  jor  g03337(.dina(n3380), .dinb(n3555), .dout(n3556));
  jand g03338(.dina(n3556), .dinb(n3544), .dout(n3557));
  jand g03339(.dina(n3557), .dinb(n2572), .dout(n3558));
  jnot g03340(.din(n3388), .dout(n3559));
  jor  g03341(.dina(n3559), .dinb(n3558), .dout(n3560));
  jand g03342(.dina(n3560), .dinb(n3543), .dout(n3561));
  jand g03343(.dina(n3561), .dinb(n2345), .dout(n3562));
  jnot g03344(.din(n3395), .dout(n3563));
  jor  g03345(.dina(n3563), .dinb(n3562), .dout(n3564));
  jand g03346(.dina(n3564), .dinb(n3542), .dout(n3565));
  jand g03347(.dina(n3565), .dinb(n2108), .dout(n3566));
  jor  g03348(.dina(n3402), .dinb(n3566), .dout(n3567));
  jand g03349(.dina(n3567), .dinb(n3541), .dout(n3568));
  jand g03350(.dina(n3568), .dinb(n1912), .dout(n3569));
  jor  g03351(.dina(n3410), .dinb(n3569), .dout(n3570));
  jand g03352(.dina(n3570), .dinb(n3540), .dout(n3571));
  jand g03353(.dina(n3571), .dinb(n1699), .dout(n3572));
  jnot g03354(.din(n3418), .dout(n3573));
  jor  g03355(.dina(n3573), .dinb(n3572), .dout(n3574));
  jand g03356(.dina(n3574), .dinb(n3539), .dout(n3575));
  jand g03357(.dina(n3575), .dinb(n1516), .dout(n3576));
  jor  g03358(.dina(n3425), .dinb(n3576), .dout(n3577));
  jand g03359(.dina(n3577), .dinb(n3538), .dout(n3578));
  jand g03360(.dina(n3578), .dinb(n1332), .dout(n3579));
  jnot g03361(.din(n3433), .dout(n3580));
  jor  g03362(.dina(n3580), .dinb(n3579), .dout(n3581));
  jand g03363(.dina(n3581), .dinb(n3537), .dout(n3582));
  jand g03364(.dina(n3582), .dinb(n1173), .dout(n3583));
  jor  g03365(.dina(n3440), .dinb(n3583), .dout(n3584));
  jand g03366(.dina(n3584), .dinb(n3536), .dout(n3585));
  jand g03367(.dina(n3585), .dinb(n1008), .dout(n3586));
  jnot g03368(.din(n3448), .dout(n3587));
  jor  g03369(.dina(n3587), .dinb(n3586), .dout(n3588));
  jand g03370(.dina(n3588), .dinb(n3535), .dout(n3589));
  jand g03371(.dina(n3589), .dinb(n884), .dout(n3590));
  jor  g03372(.dina(n3455), .dinb(n3590), .dout(n3591));
  jand g03373(.dina(n3591), .dinb(n3534), .dout(n3592));
  jand g03374(.dina(n3592), .dinb(n743), .dout(n3593));
  jnot g03375(.din(n3463), .dout(n3594));
  jor  g03376(.dina(n3594), .dinb(n3593), .dout(n3595));
  jand g03377(.dina(n3595), .dinb(n3533), .dout(n3596));
  jand g03378(.dina(n3596), .dinb(n635), .dout(n3597));
  jor  g03379(.dina(n3470), .dinb(n3597), .dout(n3598));
  jand g03380(.dina(n3598), .dinb(n3532), .dout(n3599));
  jand g03381(.dina(n3599), .dinb(n515), .dout(n3600));
  jnot g03382(.din(n3478), .dout(n3601));
  jor  g03383(.dina(n3601), .dinb(n3600), .dout(n3602));
  jand g03384(.dina(n3602), .dinb(n3531), .dout(n3603));
  jand g03385(.dina(n3603), .dinb(n443), .dout(n3604));
  jor  g03386(.dina(n3485), .dinb(n3604), .dout(n3605));
  jand g03387(.dina(n3605), .dinb(n3530), .dout(n3606));
  jand g03388(.dina(n3606), .dinb(n352), .dout(n3607));
  jor  g03389(.dina(n3493), .dinb(n3607), .dout(n3608));
  jand g03390(.dina(n3608), .dinb(n3529), .dout(n3609));
  jand g03391(.dina(n3609), .dinb(n294), .dout(n3610));
  jnot g03392(.din(n3501), .dout(n3611));
  jor  g03393(.dina(n3611), .dinb(n3610), .dout(n3612));
  jand g03394(.dina(n3612), .dinb(n3528), .dout(n3613));
  jand g03395(.dina(n3613), .dinb(n239), .dout(n3614));
  jnot g03396(.din(n3508), .dout(n3615));
  jor  g03397(.dina(n3615), .dinb(n3614), .dout(n3616));
  jand g03398(.dina(n3616), .dinb(n3527), .dout(n3617));
  jand g03399(.dina(n3617), .dinb(n221), .dout(n3618));
  jor  g03400(.dina(n3515), .dinb(n3618), .dout(n3619));
  jand g03401(.dina(n3619), .dinb(n3526), .dout(n3620));
  jor  g03402(.dina(n3521), .dinb(n3620), .dout(n3621));
  jxor g03403(.dina(n3240), .dinb(n3237), .dout(n3622));
  jnot g03404(.din(n3622), .dout(n3623));
  jand g03405(.dina(n3623), .dinb(asqrt[42] ), .dout(n3624));
  jor  g03406(.dina(n3624), .dinb(n3621), .dout(n3625));
  jand g03407(.dina(n3625), .dinb(n218), .dout(n3626));
  jand g03408(.dina(n3367), .dinb(n3237), .dout(n3627));
  jnot g03409(.din(n3627), .dout(n3628));
  jand g03410(.dina(n3622), .dinb(asqrt[63] ), .dout(n3629));
  jand g03411(.dina(n3629), .dinb(n3628), .dout(n3630));
  jor  g03412(.dina(n3630), .dinb(n3626), .dout(n3631));
  jor  g03413(.dina(n3631), .dinb(n3524), .dout(asqrt[41] ));
  jand g03414(.dina(n3522), .dinb(n3518), .dout(n3635));
  jnot g03415(.din(n3624), .dout(n3636));
  jand g03416(.dina(n3636), .dinb(n3635), .dout(n3637));
  jor  g03417(.dina(n3637), .dinb(asqrt[63] ), .dout(n3638));
  jnot g03418(.din(n3630), .dout(n3639));
  jand g03419(.dina(n3639), .dinb(n3638), .dout(n3640));
  jand g03420(.dina(n3640), .dinb(n3523), .dout(n3642));
  jxor g03421(.dina(n3510), .dinb(n221), .dout(n3643));
  jor  g03422(.dina(n3643), .dinb(n3642), .dout(n3644));
  jxor g03423(.dina(n3644), .dinb(n3515), .dout(n3645));
  jnot g03424(.din(n3645), .dout(n3646));
  jor  g03425(.dina(n3642), .dinb(n3258), .dout(n3647));
  jnot g03426(.din(a[80] ), .dout(n3648));
  jnot g03427(.din(a[81] ), .dout(n3649));
  jand g03428(.dina(n3649), .dinb(n3648), .dout(n3650));
  jand g03429(.dina(n3650), .dinb(n3258), .dout(n3651));
  jnot g03430(.din(n3651), .dout(n3652));
  jand g03431(.dina(n3652), .dinb(n3647), .dout(n3653));
  jor  g03432(.dina(n3653), .dinb(n3368), .dout(n3654));
  jand g03433(.dina(n3653), .dinb(n3368), .dout(n3655));
  jor  g03434(.dina(n3642), .dinb(a[82] ), .dout(n3656));
  jand g03435(.dina(n3656), .dinb(a[83] ), .dout(n3657));
  jand g03436(.dina(asqrt[41] ), .dinb(n3260), .dout(n3658));
  jor  g03437(.dina(n3658), .dinb(n3657), .dout(n3659));
  jor  g03438(.dina(n3659), .dinb(n3655), .dout(n3660));
  jand g03439(.dina(n3660), .dinb(n3654), .dout(n3661));
  jor  g03440(.dina(n3661), .dinb(n3089), .dout(n3662));
  jand g03441(.dina(n3661), .dinb(n3089), .dout(n3663));
  jnot g03442(.din(n3260), .dout(n3664));
  jor  g03443(.dina(n3642), .dinb(n3664), .dout(n3665));
  jor  g03444(.dina(n3629), .dinb(n3524), .dout(n3666));
  jor  g03445(.dina(n3666), .dinb(n3626), .dout(n3667));
  jor  g03446(.dina(n3667), .dinb(n3368), .dout(n3668));
  jand g03447(.dina(n3668), .dinb(n3665), .dout(n3669));
  jxor g03448(.dina(n3669), .dinb(n3075), .dout(n3670));
  jor  g03449(.dina(n3670), .dinb(n3663), .dout(n3671));
  jand g03450(.dina(n3671), .dinb(n3662), .dout(n3672));
  jor  g03451(.dina(n3672), .dinb(n2833), .dout(n3673));
  jand g03452(.dina(n3672), .dinb(n2833), .dout(n3674));
  jxor g03453(.dina(n3262), .dinb(n3089), .dout(n3675));
  jor  g03454(.dina(n3675), .dinb(n3642), .dout(n3676));
  jxor g03455(.dina(n3676), .dinb(n3552), .dout(n3677));
  jnot g03456(.din(n3677), .dout(n3678));
  jor  g03457(.dina(n3678), .dinb(n3674), .dout(n3679));
  jand g03458(.dina(n3679), .dinb(n3673), .dout(n3680));
  jor  g03459(.dina(n3680), .dinb(n2572), .dout(n3681));
  jand g03460(.dina(n3680), .dinb(n2572), .dout(n3682));
  jxor g03461(.dina(n3372), .dinb(n2833), .dout(n3683));
  jor  g03462(.dina(n3683), .dinb(n3642), .dout(n3684));
  jxor g03463(.dina(n3684), .dinb(n3381), .dout(n3685));
  jor  g03464(.dina(n3685), .dinb(n3682), .dout(n3686));
  jand g03465(.dina(n3686), .dinb(n3681), .dout(n3687));
  jor  g03466(.dina(n3687), .dinb(n2345), .dout(n3688));
  jand g03467(.dina(n3687), .dinb(n2345), .dout(n3689));
  jxor g03468(.dina(n3383), .dinb(n2572), .dout(n3690));
  jor  g03469(.dina(n3690), .dinb(n3642), .dout(n3691));
  jxor g03470(.dina(n3691), .dinb(n3559), .dout(n3692));
  jnot g03471(.din(n3692), .dout(n3693));
  jor  g03472(.dina(n3693), .dinb(n3689), .dout(n3694));
  jand g03473(.dina(n3694), .dinb(n3688), .dout(n3695));
  jor  g03474(.dina(n3695), .dinb(n2108), .dout(n3696));
  jand g03475(.dina(n3695), .dinb(n2108), .dout(n3697));
  jxor g03476(.dina(n3390), .dinb(n2345), .dout(n3698));
  jor  g03477(.dina(n3698), .dinb(n3642), .dout(n3699));
  jxor g03478(.dina(n3699), .dinb(n3563), .dout(n3700));
  jnot g03479(.din(n3700), .dout(n3701));
  jor  g03480(.dina(n3701), .dinb(n3697), .dout(n3702));
  jand g03481(.dina(n3702), .dinb(n3696), .dout(n3703));
  jor  g03482(.dina(n3703), .dinb(n1912), .dout(n3704));
  jand g03483(.dina(n3703), .dinb(n1912), .dout(n3705));
  jxor g03484(.dina(n3397), .dinb(n2108), .dout(n3706));
  jor  g03485(.dina(n3706), .dinb(n3642), .dout(n3707));
  jxor g03486(.dina(n3707), .dinb(n3403), .dout(n3708));
  jor  g03487(.dina(n3708), .dinb(n3705), .dout(n3709));
  jand g03488(.dina(n3709), .dinb(n3704), .dout(n3710));
  jor  g03489(.dina(n3710), .dinb(n1699), .dout(n3711));
  jand g03490(.dina(n3710), .dinb(n1699), .dout(n3712));
  jxor g03491(.dina(n3405), .dinb(n1912), .dout(n3713));
  jor  g03492(.dina(n3713), .dinb(n3642), .dout(n3714));
  jxor g03493(.dina(n3714), .dinb(n3411), .dout(n3715));
  jor  g03494(.dina(n3715), .dinb(n3712), .dout(n3716));
  jand g03495(.dina(n3716), .dinb(n3711), .dout(n3717));
  jor  g03496(.dina(n3717), .dinb(n1516), .dout(n3718));
  jand g03497(.dina(n3717), .dinb(n1516), .dout(n3719));
  jxor g03498(.dina(n3413), .dinb(n1699), .dout(n3720));
  jor  g03499(.dina(n3720), .dinb(n3642), .dout(n3721));
  jxor g03500(.dina(n3721), .dinb(n3573), .dout(n3722));
  jnot g03501(.din(n3722), .dout(n3723));
  jor  g03502(.dina(n3723), .dinb(n3719), .dout(n3724));
  jand g03503(.dina(n3724), .dinb(n3718), .dout(n3725));
  jor  g03504(.dina(n3725), .dinb(n1332), .dout(n3726));
  jand g03505(.dina(n3725), .dinb(n1332), .dout(n3727));
  jxor g03506(.dina(n3420), .dinb(n1516), .dout(n3728));
  jor  g03507(.dina(n3728), .dinb(n3642), .dout(n3729));
  jxor g03508(.dina(n3729), .dinb(n3426), .dout(n3730));
  jor  g03509(.dina(n3730), .dinb(n3727), .dout(n3731));
  jand g03510(.dina(n3731), .dinb(n3726), .dout(n3732));
  jor  g03511(.dina(n3732), .dinb(n1173), .dout(n3733));
  jand g03512(.dina(n3732), .dinb(n1173), .dout(n3734));
  jxor g03513(.dina(n3428), .dinb(n1332), .dout(n3735));
  jor  g03514(.dina(n3735), .dinb(n3642), .dout(n3736));
  jxor g03515(.dina(n3736), .dinb(n3580), .dout(n3737));
  jnot g03516(.din(n3737), .dout(n3738));
  jor  g03517(.dina(n3738), .dinb(n3734), .dout(n3739));
  jand g03518(.dina(n3739), .dinb(n3733), .dout(n3740));
  jor  g03519(.dina(n3740), .dinb(n1008), .dout(n3741));
  jand g03520(.dina(n3740), .dinb(n1008), .dout(n3742));
  jxor g03521(.dina(n3435), .dinb(n1173), .dout(n3743));
  jor  g03522(.dina(n3743), .dinb(n3642), .dout(n3744));
  jxor g03523(.dina(n3744), .dinb(n3441), .dout(n3745));
  jor  g03524(.dina(n3745), .dinb(n3742), .dout(n3746));
  jand g03525(.dina(n3746), .dinb(n3741), .dout(n3747));
  jor  g03526(.dina(n3747), .dinb(n884), .dout(n3748));
  jand g03527(.dina(n3747), .dinb(n884), .dout(n3749));
  jxor g03528(.dina(n3443), .dinb(n1008), .dout(n3750));
  jor  g03529(.dina(n3750), .dinb(n3642), .dout(n3751));
  jxor g03530(.dina(n3751), .dinb(n3587), .dout(n3752));
  jnot g03531(.din(n3752), .dout(n3753));
  jor  g03532(.dina(n3753), .dinb(n3749), .dout(n3754));
  jand g03533(.dina(n3754), .dinb(n3748), .dout(n3755));
  jor  g03534(.dina(n3755), .dinb(n743), .dout(n3756));
  jand g03535(.dina(n3755), .dinb(n743), .dout(n3757));
  jxor g03536(.dina(n3450), .dinb(n884), .dout(n3758));
  jor  g03537(.dina(n3758), .dinb(n3642), .dout(n3759));
  jxor g03538(.dina(n3759), .dinb(n3456), .dout(n3760));
  jor  g03539(.dina(n3760), .dinb(n3757), .dout(n3761));
  jand g03540(.dina(n3761), .dinb(n3756), .dout(n3762));
  jor  g03541(.dina(n3762), .dinb(n635), .dout(n3763));
  jand g03542(.dina(n3762), .dinb(n635), .dout(n3764));
  jxor g03543(.dina(n3458), .dinb(n743), .dout(n3765));
  jor  g03544(.dina(n3765), .dinb(n3642), .dout(n3766));
  jxor g03545(.dina(n3766), .dinb(n3594), .dout(n3767));
  jnot g03546(.din(n3767), .dout(n3768));
  jor  g03547(.dina(n3768), .dinb(n3764), .dout(n3769));
  jand g03548(.dina(n3769), .dinb(n3763), .dout(n3770));
  jor  g03549(.dina(n3770), .dinb(n515), .dout(n3771));
  jand g03550(.dina(n3770), .dinb(n515), .dout(n3772));
  jxor g03551(.dina(n3465), .dinb(n635), .dout(n3773));
  jor  g03552(.dina(n3773), .dinb(n3642), .dout(n3774));
  jxor g03553(.dina(n3774), .dinb(n3471), .dout(n3775));
  jor  g03554(.dina(n3775), .dinb(n3772), .dout(n3776));
  jand g03555(.dina(n3776), .dinb(n3771), .dout(n3777));
  jor  g03556(.dina(n3777), .dinb(n443), .dout(n3778));
  jand g03557(.dina(n3777), .dinb(n443), .dout(n3779));
  jxor g03558(.dina(n3473), .dinb(n515), .dout(n3780));
  jor  g03559(.dina(n3780), .dinb(n3642), .dout(n3781));
  jxor g03560(.dina(n3781), .dinb(n3601), .dout(n3782));
  jnot g03561(.din(n3782), .dout(n3783));
  jor  g03562(.dina(n3783), .dinb(n3779), .dout(n3784));
  jand g03563(.dina(n3784), .dinb(n3778), .dout(n3785));
  jor  g03564(.dina(n3785), .dinb(n352), .dout(n3786));
  jand g03565(.dina(n3785), .dinb(n352), .dout(n3787));
  jxor g03566(.dina(n3480), .dinb(n443), .dout(n3788));
  jor  g03567(.dina(n3788), .dinb(n3642), .dout(n3789));
  jxor g03568(.dina(n3789), .dinb(n3486), .dout(n3790));
  jor  g03569(.dina(n3790), .dinb(n3787), .dout(n3791));
  jand g03570(.dina(n3791), .dinb(n3786), .dout(n3792));
  jor  g03571(.dina(n3792), .dinb(n294), .dout(n3793));
  jand g03572(.dina(n3792), .dinb(n294), .dout(n3794));
  jxor g03573(.dina(n3488), .dinb(n352), .dout(n3795));
  jor  g03574(.dina(n3795), .dinb(n3642), .dout(n3796));
  jxor g03575(.dina(n3796), .dinb(n3494), .dout(n3797));
  jor  g03576(.dina(n3797), .dinb(n3794), .dout(n3798));
  jand g03577(.dina(n3798), .dinb(n3793), .dout(n3799));
  jor  g03578(.dina(n3799), .dinb(n239), .dout(n3800));
  jand g03579(.dina(n3799), .dinb(n239), .dout(n3801));
  jxor g03580(.dina(n3496), .dinb(n294), .dout(n3802));
  jor  g03581(.dina(n3802), .dinb(n3642), .dout(n3803));
  jxor g03582(.dina(n3803), .dinb(n3611), .dout(n3804));
  jnot g03583(.din(n3804), .dout(n3805));
  jor  g03584(.dina(n3805), .dinb(n3801), .dout(n3806));
  jand g03585(.dina(n3806), .dinb(n3800), .dout(n3807));
  jor  g03586(.dina(n3807), .dinb(n221), .dout(n3808));
  jand g03587(.dina(n3807), .dinb(n221), .dout(n3809));
  jxor g03588(.dina(n3503), .dinb(n239), .dout(n3810));
  jor  g03589(.dina(n3810), .dinb(n3642), .dout(n3811));
  jxor g03590(.dina(n3811), .dinb(n3615), .dout(n3812));
  jnot g03591(.din(n3812), .dout(n3813));
  jor  g03592(.dina(n3813), .dinb(n3809), .dout(n3814));
  jand g03593(.dina(n3814), .dinb(n3808), .dout(n3815));
  jand g03594(.dina(n3815), .dinb(n3646), .dout(n3816));
  jand g03595(.dina(n3640), .dinb(n3620), .dout(n3817));
  jand g03596(.dina(n3621), .dinb(asqrt[63] ), .dout(n3818));
  jand g03597(.dina(n3818), .dinb(n3523), .dout(n3819));
  jnot g03598(.din(n3819), .dout(n3820));
  jor  g03599(.dina(n3820), .dinb(n3817), .dout(n3821));
  jnot g03600(.din(n3821), .dout(n3822));
  jand g03601(.dina(n3631), .dinb(n3635), .dout(n3823));
  jor  g03602(.dina(n3815), .dinb(n3646), .dout(n3824));
  jor  g03603(.dina(n3824), .dinb(n3524), .dout(n3825));
  jor  g03604(.dina(n3825), .dinb(n3823), .dout(n3826));
  jand g03605(.dina(n3826), .dinb(n218), .dout(n3827));
  jand g03606(.dina(n3642), .dinb(n3521), .dout(n3828));
  jor  g03607(.dina(n3828), .dinb(n3827), .dout(n3829));
  jor  g03608(.dina(n3829), .dinb(n3822), .dout(n3830));
  jor  g03609(.dina(n3830), .dinb(n3816), .dout(asqrt[40] ));
  jxor g03610(.dina(n3807), .dinb(n221), .dout(n3832));
  jand g03611(.dina(n3832), .dinb(asqrt[40] ), .dout(n3833));
  jxor g03612(.dina(n3833), .dinb(n3812), .dout(n3834));
  jnot g03613(.din(n3834), .dout(n3835));
  jand g03614(.dina(asqrt[40] ), .dinb(a[80] ), .dout(n3836));
  jnot g03615(.din(a[78] ), .dout(n3837));
  jnot g03616(.din(a[79] ), .dout(n3838));
  jand g03617(.dina(n3838), .dinb(n3837), .dout(n3839));
  jand g03618(.dina(n3839), .dinb(n3648), .dout(n3840));
  jor  g03619(.dina(n3840), .dinb(n3836), .dout(n3841));
  jand g03620(.dina(n3841), .dinb(asqrt[41] ), .dout(n3842));
  jor  g03621(.dina(n3841), .dinb(asqrt[41] ), .dout(n3843));
  jand g03622(.dina(asqrt[40] ), .dinb(n3648), .dout(n3844));
  jor  g03623(.dina(n3844), .dinb(n3649), .dout(n3845));
  jnot g03624(.din(n3650), .dout(n3846));
  jnot g03625(.din(n3816), .dout(n3847));
  jnot g03626(.din(n3823), .dout(n3848));
  jnot g03627(.din(n3808), .dout(n3849));
  jnot g03628(.din(n3800), .dout(n3850));
  jnot g03629(.din(n3793), .dout(n3851));
  jnot g03630(.din(n3786), .dout(n3852));
  jnot g03631(.din(n3778), .dout(n3853));
  jnot g03632(.din(n3771), .dout(n3854));
  jnot g03633(.din(n3763), .dout(n3855));
  jnot g03634(.din(n3756), .dout(n3856));
  jnot g03635(.din(n3748), .dout(n3857));
  jnot g03636(.din(n3741), .dout(n3858));
  jnot g03637(.din(n3733), .dout(n3859));
  jnot g03638(.din(n3726), .dout(n3860));
  jnot g03639(.din(n3718), .dout(n3861));
  jnot g03640(.din(n3711), .dout(n3862));
  jnot g03641(.din(n3704), .dout(n3863));
  jnot g03642(.din(n3696), .dout(n3864));
  jnot g03643(.din(n3688), .dout(n3865));
  jnot g03644(.din(n3681), .dout(n3866));
  jnot g03645(.din(n3673), .dout(n3867));
  jnot g03646(.din(n3662), .dout(n3868));
  jnot g03647(.din(n3654), .dout(n3869));
  jand g03648(.dina(asqrt[41] ), .dinb(a[82] ), .dout(n3870));
  jor  g03649(.dina(n3651), .dinb(n3870), .dout(n3871));
  jor  g03650(.dina(n3871), .dinb(asqrt[42] ), .dout(n3872));
  jand g03651(.dina(asqrt[41] ), .dinb(n3258), .dout(n3873));
  jor  g03652(.dina(n3873), .dinb(n3259), .dout(n3874));
  jand g03653(.dina(n3665), .dinb(n3874), .dout(n3875));
  jand g03654(.dina(n3875), .dinb(n3872), .dout(n3876));
  jor  g03655(.dina(n3876), .dinb(n3869), .dout(n3877));
  jor  g03656(.dina(n3877), .dinb(asqrt[43] ), .dout(n3878));
  jnot g03657(.din(n3670), .dout(n3879));
  jand g03658(.dina(n3879), .dinb(n3878), .dout(n3880));
  jor  g03659(.dina(n3880), .dinb(n3868), .dout(n3881));
  jor  g03660(.dina(n3881), .dinb(asqrt[44] ), .dout(n3882));
  jand g03661(.dina(n3677), .dinb(n3882), .dout(n3883));
  jor  g03662(.dina(n3883), .dinb(n3867), .dout(n3884));
  jor  g03663(.dina(n3884), .dinb(asqrt[45] ), .dout(n3885));
  jnot g03664(.din(n3685), .dout(n3886));
  jand g03665(.dina(n3886), .dinb(n3885), .dout(n3887));
  jor  g03666(.dina(n3887), .dinb(n3866), .dout(n3888));
  jor  g03667(.dina(n3888), .dinb(asqrt[46] ), .dout(n3889));
  jand g03668(.dina(n3692), .dinb(n3889), .dout(n3890));
  jor  g03669(.dina(n3890), .dinb(n3865), .dout(n3891));
  jor  g03670(.dina(n3891), .dinb(asqrt[47] ), .dout(n3892));
  jand g03671(.dina(n3700), .dinb(n3892), .dout(n3893));
  jor  g03672(.dina(n3893), .dinb(n3864), .dout(n3894));
  jor  g03673(.dina(n3894), .dinb(asqrt[48] ), .dout(n3895));
  jnot g03674(.din(n3708), .dout(n3896));
  jand g03675(.dina(n3896), .dinb(n3895), .dout(n3897));
  jor  g03676(.dina(n3897), .dinb(n3863), .dout(n3898));
  jor  g03677(.dina(n3898), .dinb(asqrt[49] ), .dout(n3899));
  jnot g03678(.din(n3715), .dout(n3900));
  jand g03679(.dina(n3900), .dinb(n3899), .dout(n3901));
  jor  g03680(.dina(n3901), .dinb(n3862), .dout(n3902));
  jor  g03681(.dina(n3902), .dinb(asqrt[50] ), .dout(n3903));
  jand g03682(.dina(n3722), .dinb(n3903), .dout(n3904));
  jor  g03683(.dina(n3904), .dinb(n3861), .dout(n3905));
  jor  g03684(.dina(n3905), .dinb(asqrt[51] ), .dout(n3906));
  jnot g03685(.din(n3730), .dout(n3907));
  jand g03686(.dina(n3907), .dinb(n3906), .dout(n3908));
  jor  g03687(.dina(n3908), .dinb(n3860), .dout(n3909));
  jor  g03688(.dina(n3909), .dinb(asqrt[52] ), .dout(n3910));
  jand g03689(.dina(n3737), .dinb(n3910), .dout(n3911));
  jor  g03690(.dina(n3911), .dinb(n3859), .dout(n3912));
  jor  g03691(.dina(n3912), .dinb(asqrt[53] ), .dout(n3913));
  jnot g03692(.din(n3745), .dout(n3914));
  jand g03693(.dina(n3914), .dinb(n3913), .dout(n3915));
  jor  g03694(.dina(n3915), .dinb(n3858), .dout(n3916));
  jor  g03695(.dina(n3916), .dinb(asqrt[54] ), .dout(n3917));
  jand g03696(.dina(n3752), .dinb(n3917), .dout(n3918));
  jor  g03697(.dina(n3918), .dinb(n3857), .dout(n3919));
  jor  g03698(.dina(n3919), .dinb(asqrt[55] ), .dout(n3920));
  jnot g03699(.din(n3760), .dout(n3921));
  jand g03700(.dina(n3921), .dinb(n3920), .dout(n3922));
  jor  g03701(.dina(n3922), .dinb(n3856), .dout(n3923));
  jor  g03702(.dina(n3923), .dinb(asqrt[56] ), .dout(n3924));
  jand g03703(.dina(n3767), .dinb(n3924), .dout(n3925));
  jor  g03704(.dina(n3925), .dinb(n3855), .dout(n3926));
  jor  g03705(.dina(n3926), .dinb(asqrt[57] ), .dout(n3927));
  jnot g03706(.din(n3775), .dout(n3928));
  jand g03707(.dina(n3928), .dinb(n3927), .dout(n3929));
  jor  g03708(.dina(n3929), .dinb(n3854), .dout(n3930));
  jor  g03709(.dina(n3930), .dinb(asqrt[58] ), .dout(n3931));
  jand g03710(.dina(n3782), .dinb(n3931), .dout(n3932));
  jor  g03711(.dina(n3932), .dinb(n3853), .dout(n3933));
  jor  g03712(.dina(n3933), .dinb(asqrt[59] ), .dout(n3934));
  jnot g03713(.din(n3790), .dout(n3935));
  jand g03714(.dina(n3935), .dinb(n3934), .dout(n3936));
  jor  g03715(.dina(n3936), .dinb(n3852), .dout(n3937));
  jor  g03716(.dina(n3937), .dinb(asqrt[60] ), .dout(n3938));
  jnot g03717(.din(n3797), .dout(n3939));
  jand g03718(.dina(n3939), .dinb(n3938), .dout(n3940));
  jor  g03719(.dina(n3940), .dinb(n3851), .dout(n3941));
  jor  g03720(.dina(n3941), .dinb(asqrt[61] ), .dout(n3942));
  jand g03721(.dina(n3804), .dinb(n3942), .dout(n3943));
  jor  g03722(.dina(n3943), .dinb(n3850), .dout(n3944));
  jor  g03723(.dina(n3944), .dinb(asqrt[62] ), .dout(n3945));
  jand g03724(.dina(n3812), .dinb(n3945), .dout(n3946));
  jor  g03725(.dina(n3946), .dinb(n3849), .dout(n3947));
  jand g03726(.dina(n3947), .dinb(n3645), .dout(n3948));
  jand g03727(.dina(n3948), .dinb(n3523), .dout(n3949));
  jand g03728(.dina(n3949), .dinb(n3848), .dout(n3950));
  jor  g03729(.dina(n3950), .dinb(asqrt[63] ), .dout(n3951));
  jnot g03730(.din(n3828), .dout(n3952));
  jand g03731(.dina(n3952), .dinb(n3951), .dout(n3953));
  jand g03732(.dina(n3953), .dinb(n3821), .dout(n3954));
  jand g03733(.dina(n3954), .dinb(n3847), .dout(n3955));
  jor  g03734(.dina(n3955), .dinb(n3846), .dout(n3956));
  jand g03735(.dina(n3956), .dinb(n3845), .dout(n3957));
  jand g03736(.dina(n3957), .dinb(n3843), .dout(n3958));
  jor  g03737(.dina(n3958), .dinb(n3842), .dout(n3959));
  jand g03738(.dina(n3959), .dinb(asqrt[42] ), .dout(n3960));
  jor  g03739(.dina(n3959), .dinb(asqrt[42] ), .dout(n3961));
  jand g03740(.dina(asqrt[40] ), .dinb(n3650), .dout(n3962));
  jand g03741(.dina(n3847), .dinb(asqrt[41] ), .dout(n3963));
  jand g03742(.dina(n3963), .dinb(n3820), .dout(n3964));
  jand g03743(.dina(n3964), .dinb(n3951), .dout(n3965));
  jor  g03744(.dina(n3965), .dinb(n3962), .dout(n3966));
  jxor g03745(.dina(n3966), .dinb(a[82] ), .dout(n3967));
  jnot g03746(.din(n3967), .dout(n3968));
  jand g03747(.dina(n3968), .dinb(n3961), .dout(n3969));
  jor  g03748(.dina(n3969), .dinb(n3960), .dout(n3970));
  jand g03749(.dina(n3970), .dinb(asqrt[43] ), .dout(n3971));
  jor  g03750(.dina(n3970), .dinb(asqrt[43] ), .dout(n3972));
  jxor g03751(.dina(n3653), .dinb(n3368), .dout(n3973));
  jand g03752(.dina(n3973), .dinb(asqrt[40] ), .dout(n3974));
  jxor g03753(.dina(n3974), .dinb(n3875), .dout(n3975));
  jand g03754(.dina(n3975), .dinb(n3972), .dout(n3976));
  jor  g03755(.dina(n3976), .dinb(n3971), .dout(n3977));
  jand g03756(.dina(n3977), .dinb(asqrt[44] ), .dout(n3978));
  jor  g03757(.dina(n3977), .dinb(asqrt[44] ), .dout(n3979));
  jxor g03758(.dina(n3661), .dinb(n3089), .dout(n3980));
  jand g03759(.dina(n3980), .dinb(asqrt[40] ), .dout(n3981));
  jxor g03760(.dina(n3981), .dinb(n3670), .dout(n3982));
  jnot g03761(.din(n3982), .dout(n3983));
  jand g03762(.dina(n3983), .dinb(n3979), .dout(n3984));
  jor  g03763(.dina(n3984), .dinb(n3978), .dout(n3985));
  jand g03764(.dina(n3985), .dinb(asqrt[45] ), .dout(n3986));
  jor  g03765(.dina(n3985), .dinb(asqrt[45] ), .dout(n3987));
  jxor g03766(.dina(n3672), .dinb(n2833), .dout(n3988));
  jand g03767(.dina(n3988), .dinb(asqrt[40] ), .dout(n3989));
  jxor g03768(.dina(n3989), .dinb(n3677), .dout(n3990));
  jand g03769(.dina(n3990), .dinb(n3987), .dout(n3991));
  jor  g03770(.dina(n3991), .dinb(n3986), .dout(n3992));
  jand g03771(.dina(n3992), .dinb(asqrt[46] ), .dout(n3993));
  jor  g03772(.dina(n3992), .dinb(asqrt[46] ), .dout(n3994));
  jxor g03773(.dina(n3680), .dinb(n2572), .dout(n3995));
  jand g03774(.dina(n3995), .dinb(asqrt[40] ), .dout(n3996));
  jxor g03775(.dina(n3996), .dinb(n3685), .dout(n3997));
  jnot g03776(.din(n3997), .dout(n3998));
  jand g03777(.dina(n3998), .dinb(n3994), .dout(n3999));
  jor  g03778(.dina(n3999), .dinb(n3993), .dout(n4000));
  jand g03779(.dina(n4000), .dinb(asqrt[47] ), .dout(n4001));
  jor  g03780(.dina(n4000), .dinb(asqrt[47] ), .dout(n4002));
  jxor g03781(.dina(n3687), .dinb(n2345), .dout(n4003));
  jand g03782(.dina(n4003), .dinb(asqrt[40] ), .dout(n4004));
  jxor g03783(.dina(n4004), .dinb(n3692), .dout(n4005));
  jand g03784(.dina(n4005), .dinb(n4002), .dout(n4006));
  jor  g03785(.dina(n4006), .dinb(n4001), .dout(n4007));
  jand g03786(.dina(n4007), .dinb(asqrt[48] ), .dout(n4008));
  jor  g03787(.dina(n4007), .dinb(asqrt[48] ), .dout(n4009));
  jxor g03788(.dina(n3695), .dinb(n2108), .dout(n4010));
  jand g03789(.dina(n4010), .dinb(asqrt[40] ), .dout(n4011));
  jxor g03790(.dina(n4011), .dinb(n3700), .dout(n4012));
  jand g03791(.dina(n4012), .dinb(n4009), .dout(n4013));
  jor  g03792(.dina(n4013), .dinb(n4008), .dout(n4014));
  jand g03793(.dina(n4014), .dinb(asqrt[49] ), .dout(n4015));
  jor  g03794(.dina(n4014), .dinb(asqrt[49] ), .dout(n4016));
  jxor g03795(.dina(n3703), .dinb(n1912), .dout(n4017));
  jand g03796(.dina(n4017), .dinb(asqrt[40] ), .dout(n4018));
  jxor g03797(.dina(n4018), .dinb(n3708), .dout(n4019));
  jnot g03798(.din(n4019), .dout(n4020));
  jand g03799(.dina(n4020), .dinb(n4016), .dout(n4021));
  jor  g03800(.dina(n4021), .dinb(n4015), .dout(n4022));
  jand g03801(.dina(n4022), .dinb(asqrt[50] ), .dout(n4023));
  jor  g03802(.dina(n4022), .dinb(asqrt[50] ), .dout(n4024));
  jxor g03803(.dina(n3710), .dinb(n1699), .dout(n4025));
  jand g03804(.dina(n4025), .dinb(asqrt[40] ), .dout(n4026));
  jxor g03805(.dina(n4026), .dinb(n3715), .dout(n4027));
  jnot g03806(.din(n4027), .dout(n4028));
  jand g03807(.dina(n4028), .dinb(n4024), .dout(n4029));
  jor  g03808(.dina(n4029), .dinb(n4023), .dout(n4030));
  jand g03809(.dina(n4030), .dinb(asqrt[51] ), .dout(n4031));
  jor  g03810(.dina(n4030), .dinb(asqrt[51] ), .dout(n4032));
  jxor g03811(.dina(n3717), .dinb(n1516), .dout(n4033));
  jand g03812(.dina(n4033), .dinb(asqrt[40] ), .dout(n4034));
  jxor g03813(.dina(n4034), .dinb(n3722), .dout(n4035));
  jand g03814(.dina(n4035), .dinb(n4032), .dout(n4036));
  jor  g03815(.dina(n4036), .dinb(n4031), .dout(n4037));
  jand g03816(.dina(n4037), .dinb(asqrt[52] ), .dout(n4038));
  jor  g03817(.dina(n4037), .dinb(asqrt[52] ), .dout(n4039));
  jxor g03818(.dina(n3725), .dinb(n1332), .dout(n4040));
  jand g03819(.dina(n4040), .dinb(asqrt[40] ), .dout(n4041));
  jxor g03820(.dina(n4041), .dinb(n3730), .dout(n4042));
  jnot g03821(.din(n4042), .dout(n4043));
  jand g03822(.dina(n4043), .dinb(n4039), .dout(n4044));
  jor  g03823(.dina(n4044), .dinb(n4038), .dout(n4045));
  jand g03824(.dina(n4045), .dinb(asqrt[53] ), .dout(n4046));
  jor  g03825(.dina(n4045), .dinb(asqrt[53] ), .dout(n4047));
  jxor g03826(.dina(n3732), .dinb(n1173), .dout(n4048));
  jand g03827(.dina(n4048), .dinb(asqrt[40] ), .dout(n4049));
  jxor g03828(.dina(n4049), .dinb(n3737), .dout(n4050));
  jand g03829(.dina(n4050), .dinb(n4047), .dout(n4051));
  jor  g03830(.dina(n4051), .dinb(n4046), .dout(n4052));
  jand g03831(.dina(n4052), .dinb(asqrt[54] ), .dout(n4053));
  jor  g03832(.dina(n4052), .dinb(asqrt[54] ), .dout(n4054));
  jxor g03833(.dina(n3740), .dinb(n1008), .dout(n4055));
  jand g03834(.dina(n4055), .dinb(asqrt[40] ), .dout(n4056));
  jxor g03835(.dina(n4056), .dinb(n3745), .dout(n4057));
  jnot g03836(.din(n4057), .dout(n4058));
  jand g03837(.dina(n4058), .dinb(n4054), .dout(n4059));
  jor  g03838(.dina(n4059), .dinb(n4053), .dout(n4060));
  jand g03839(.dina(n4060), .dinb(asqrt[55] ), .dout(n4061));
  jor  g03840(.dina(n4060), .dinb(asqrt[55] ), .dout(n4062));
  jxor g03841(.dina(n3747), .dinb(n884), .dout(n4063));
  jand g03842(.dina(n4063), .dinb(asqrt[40] ), .dout(n4064));
  jxor g03843(.dina(n4064), .dinb(n3752), .dout(n4065));
  jand g03844(.dina(n4065), .dinb(n4062), .dout(n4066));
  jor  g03845(.dina(n4066), .dinb(n4061), .dout(n4067));
  jand g03846(.dina(n4067), .dinb(asqrt[56] ), .dout(n4068));
  jor  g03847(.dina(n4067), .dinb(asqrt[56] ), .dout(n4069));
  jxor g03848(.dina(n3755), .dinb(n743), .dout(n4070));
  jand g03849(.dina(n4070), .dinb(asqrt[40] ), .dout(n4071));
  jxor g03850(.dina(n4071), .dinb(n3760), .dout(n4072));
  jnot g03851(.din(n4072), .dout(n4073));
  jand g03852(.dina(n4073), .dinb(n4069), .dout(n4074));
  jor  g03853(.dina(n4074), .dinb(n4068), .dout(n4075));
  jand g03854(.dina(n4075), .dinb(asqrt[57] ), .dout(n4076));
  jor  g03855(.dina(n4075), .dinb(asqrt[57] ), .dout(n4077));
  jxor g03856(.dina(n3762), .dinb(n635), .dout(n4078));
  jand g03857(.dina(n4078), .dinb(asqrt[40] ), .dout(n4079));
  jxor g03858(.dina(n4079), .dinb(n3767), .dout(n4080));
  jand g03859(.dina(n4080), .dinb(n4077), .dout(n4081));
  jor  g03860(.dina(n4081), .dinb(n4076), .dout(n4082));
  jand g03861(.dina(n4082), .dinb(asqrt[58] ), .dout(n4083));
  jor  g03862(.dina(n4082), .dinb(asqrt[58] ), .dout(n4084));
  jxor g03863(.dina(n3770), .dinb(n515), .dout(n4085));
  jand g03864(.dina(n4085), .dinb(asqrt[40] ), .dout(n4086));
  jxor g03865(.dina(n4086), .dinb(n3775), .dout(n4087));
  jnot g03866(.din(n4087), .dout(n4088));
  jand g03867(.dina(n4088), .dinb(n4084), .dout(n4089));
  jor  g03868(.dina(n4089), .dinb(n4083), .dout(n4090));
  jand g03869(.dina(n4090), .dinb(asqrt[59] ), .dout(n4091));
  jor  g03870(.dina(n4090), .dinb(asqrt[59] ), .dout(n4092));
  jxor g03871(.dina(n3777), .dinb(n443), .dout(n4093));
  jand g03872(.dina(n4093), .dinb(asqrt[40] ), .dout(n4094));
  jxor g03873(.dina(n4094), .dinb(n3782), .dout(n4095));
  jand g03874(.dina(n4095), .dinb(n4092), .dout(n4096));
  jor  g03875(.dina(n4096), .dinb(n4091), .dout(n4097));
  jand g03876(.dina(n4097), .dinb(asqrt[60] ), .dout(n4098));
  jor  g03877(.dina(n4097), .dinb(asqrt[60] ), .dout(n4099));
  jxor g03878(.dina(n3785), .dinb(n352), .dout(n4100));
  jand g03879(.dina(n4100), .dinb(asqrt[40] ), .dout(n4101));
  jxor g03880(.dina(n4101), .dinb(n3790), .dout(n4102));
  jnot g03881(.din(n4102), .dout(n4103));
  jand g03882(.dina(n4103), .dinb(n4099), .dout(n4104));
  jor  g03883(.dina(n4104), .dinb(n4098), .dout(n4105));
  jand g03884(.dina(n4105), .dinb(asqrt[61] ), .dout(n4106));
  jor  g03885(.dina(n4105), .dinb(asqrt[61] ), .dout(n4107));
  jxor g03886(.dina(n3792), .dinb(n294), .dout(n4108));
  jand g03887(.dina(n4108), .dinb(asqrt[40] ), .dout(n4109));
  jxor g03888(.dina(n4109), .dinb(n3797), .dout(n4110));
  jnot g03889(.din(n4110), .dout(n4111));
  jand g03890(.dina(n4111), .dinb(n4107), .dout(n4112));
  jor  g03891(.dina(n4112), .dinb(n4106), .dout(n4113));
  jand g03892(.dina(n4113), .dinb(asqrt[62] ), .dout(n4114));
  jnot g03893(.din(n4114), .dout(n4115));
  jnot g03894(.din(n4106), .dout(n4116));
  jnot g03895(.din(n4098), .dout(n4117));
  jnot g03896(.din(n4091), .dout(n4118));
  jnot g03897(.din(n4083), .dout(n4119));
  jnot g03898(.din(n4076), .dout(n4120));
  jnot g03899(.din(n4068), .dout(n4121));
  jnot g03900(.din(n4061), .dout(n4122));
  jnot g03901(.din(n4053), .dout(n4123));
  jnot g03902(.din(n4046), .dout(n4124));
  jnot g03903(.din(n4038), .dout(n4125));
  jnot g03904(.din(n4031), .dout(n4126));
  jnot g03905(.din(n4023), .dout(n4127));
  jnot g03906(.din(n4015), .dout(n4128));
  jnot g03907(.din(n4008), .dout(n4129));
  jnot g03908(.din(n4001), .dout(n4130));
  jnot g03909(.din(n3993), .dout(n4131));
  jnot g03910(.din(n3986), .dout(n4132));
  jnot g03911(.din(n3978), .dout(n4133));
  jnot g03912(.din(n3971), .dout(n4134));
  jnot g03913(.din(n3960), .dout(n4135));
  jnot g03914(.din(n3842), .dout(n4136));
  jor  g03915(.dina(n3955), .dinb(n3648), .dout(n4137));
  jnot g03916(.din(n3840), .dout(n4138));
  jand g03917(.dina(n4138), .dinb(n4137), .dout(n4139));
  jand g03918(.dina(n4139), .dinb(n3642), .dout(n4140));
  jor  g03919(.dina(n3955), .dinb(a[80] ), .dout(n4141));
  jand g03920(.dina(n4141), .dinb(a[81] ), .dout(n4142));
  jor  g03921(.dina(n3962), .dinb(n4142), .dout(n4143));
  jor  g03922(.dina(n4143), .dinb(n4140), .dout(n4144));
  jand g03923(.dina(n4144), .dinb(n4136), .dout(n4145));
  jand g03924(.dina(n4145), .dinb(n3368), .dout(n4146));
  jor  g03925(.dina(n3967), .dinb(n4146), .dout(n4147));
  jand g03926(.dina(n4147), .dinb(n4135), .dout(n4148));
  jand g03927(.dina(n4148), .dinb(n3089), .dout(n4149));
  jnot g03928(.din(n3975), .dout(n4150));
  jor  g03929(.dina(n4150), .dinb(n4149), .dout(n4151));
  jand g03930(.dina(n4151), .dinb(n4134), .dout(n4152));
  jand g03931(.dina(n4152), .dinb(n2833), .dout(n4153));
  jor  g03932(.dina(n3982), .dinb(n4153), .dout(n4154));
  jand g03933(.dina(n4154), .dinb(n4133), .dout(n4155));
  jand g03934(.dina(n4155), .dinb(n2572), .dout(n4156));
  jnot g03935(.din(n3990), .dout(n4157));
  jor  g03936(.dina(n4157), .dinb(n4156), .dout(n4158));
  jand g03937(.dina(n4158), .dinb(n4132), .dout(n4159));
  jand g03938(.dina(n4159), .dinb(n2345), .dout(n4160));
  jor  g03939(.dina(n3997), .dinb(n4160), .dout(n4161));
  jand g03940(.dina(n4161), .dinb(n4131), .dout(n4162));
  jand g03941(.dina(n4162), .dinb(n2108), .dout(n4163));
  jnot g03942(.din(n4005), .dout(n4164));
  jor  g03943(.dina(n4164), .dinb(n4163), .dout(n4165));
  jand g03944(.dina(n4165), .dinb(n4130), .dout(n4166));
  jand g03945(.dina(n4166), .dinb(n1912), .dout(n4167));
  jnot g03946(.din(n4012), .dout(n4168));
  jor  g03947(.dina(n4168), .dinb(n4167), .dout(n4169));
  jand g03948(.dina(n4169), .dinb(n4129), .dout(n4170));
  jand g03949(.dina(n4170), .dinb(n1699), .dout(n4171));
  jor  g03950(.dina(n4019), .dinb(n4171), .dout(n4172));
  jand g03951(.dina(n4172), .dinb(n4128), .dout(n4173));
  jand g03952(.dina(n4173), .dinb(n1516), .dout(n4174));
  jor  g03953(.dina(n4027), .dinb(n4174), .dout(n4175));
  jand g03954(.dina(n4175), .dinb(n4127), .dout(n4176));
  jand g03955(.dina(n4176), .dinb(n1332), .dout(n4177));
  jnot g03956(.din(n4035), .dout(n4178));
  jor  g03957(.dina(n4178), .dinb(n4177), .dout(n4179));
  jand g03958(.dina(n4179), .dinb(n4126), .dout(n4180));
  jand g03959(.dina(n4180), .dinb(n1173), .dout(n4181));
  jor  g03960(.dina(n4042), .dinb(n4181), .dout(n4182));
  jand g03961(.dina(n4182), .dinb(n4125), .dout(n4183));
  jand g03962(.dina(n4183), .dinb(n1008), .dout(n4184));
  jnot g03963(.din(n4050), .dout(n4185));
  jor  g03964(.dina(n4185), .dinb(n4184), .dout(n4186));
  jand g03965(.dina(n4186), .dinb(n4124), .dout(n4187));
  jand g03966(.dina(n4187), .dinb(n884), .dout(n4188));
  jor  g03967(.dina(n4057), .dinb(n4188), .dout(n4189));
  jand g03968(.dina(n4189), .dinb(n4123), .dout(n4190));
  jand g03969(.dina(n4190), .dinb(n743), .dout(n4191));
  jnot g03970(.din(n4065), .dout(n4192));
  jor  g03971(.dina(n4192), .dinb(n4191), .dout(n4193));
  jand g03972(.dina(n4193), .dinb(n4122), .dout(n4194));
  jand g03973(.dina(n4194), .dinb(n635), .dout(n4195));
  jor  g03974(.dina(n4072), .dinb(n4195), .dout(n4196));
  jand g03975(.dina(n4196), .dinb(n4121), .dout(n4197));
  jand g03976(.dina(n4197), .dinb(n515), .dout(n4198));
  jnot g03977(.din(n4080), .dout(n4199));
  jor  g03978(.dina(n4199), .dinb(n4198), .dout(n4200));
  jand g03979(.dina(n4200), .dinb(n4120), .dout(n4201));
  jand g03980(.dina(n4201), .dinb(n443), .dout(n4202));
  jor  g03981(.dina(n4087), .dinb(n4202), .dout(n4203));
  jand g03982(.dina(n4203), .dinb(n4119), .dout(n4204));
  jand g03983(.dina(n4204), .dinb(n352), .dout(n4205));
  jnot g03984(.din(n4095), .dout(n4206));
  jor  g03985(.dina(n4206), .dinb(n4205), .dout(n4207));
  jand g03986(.dina(n4207), .dinb(n4118), .dout(n4208));
  jand g03987(.dina(n4208), .dinb(n294), .dout(n4209));
  jor  g03988(.dina(n4102), .dinb(n4209), .dout(n4210));
  jand g03989(.dina(n4210), .dinb(n4117), .dout(n4211));
  jand g03990(.dina(n4211), .dinb(n239), .dout(n4212));
  jor  g03991(.dina(n4110), .dinb(n4212), .dout(n4213));
  jand g03992(.dina(n4213), .dinb(n4116), .dout(n4214));
  jand g03993(.dina(n4214), .dinb(n221), .dout(n4215));
  jxor g03994(.dina(n3799), .dinb(n239), .dout(n4216));
  jand g03995(.dina(n4216), .dinb(asqrt[40] ), .dout(n4217));
  jxor g03996(.dina(n4217), .dinb(n3804), .dout(n4218));
  jnot g03997(.din(n4218), .dout(n4219));
  jor  g03998(.dina(n4219), .dinb(n4215), .dout(n4220));
  jand g03999(.dina(n4220), .dinb(n4115), .dout(n4221));
  jor  g04000(.dina(n4221), .dinb(n3835), .dout(n4222));
  jxor g04001(.dina(n3815), .dinb(n3646), .dout(n4223));
  jnot g04002(.din(n4223), .dout(n4224));
  jand g04003(.dina(n4224), .dinb(asqrt[40] ), .dout(n4225));
  jor  g04004(.dina(n4225), .dinb(n4222), .dout(n4226));
  jand g04005(.dina(n4226), .dinb(n218), .dout(n4227));
  jand g04006(.dina(n3955), .dinb(n3646), .dout(n4228));
  jand g04007(.dina(n4221), .dinb(n3835), .dout(n4229));
  jor  g04008(.dina(n4229), .dinb(n4228), .dout(n4230));
  jand g04009(.dina(n3954), .dinb(n3815), .dout(n4231));
  jnot g04010(.din(n4231), .dout(n4232));
  jand g04011(.dina(n4223), .dinb(asqrt[63] ), .dout(n4233));
  jand g04012(.dina(n4233), .dinb(n4232), .dout(n4234));
  jor  g04013(.dina(n4234), .dinb(n4230), .dout(n4235));
  jor  g04014(.dina(n4235), .dinb(n4227), .dout(asqrt[39] ));
  jor  g04015(.dina(n4113), .dinb(asqrt[62] ), .dout(n4237));
  jand g04016(.dina(n4218), .dinb(n4237), .dout(n4238));
  jor  g04017(.dina(n4238), .dinb(n4114), .dout(n4239));
  jand g04018(.dina(n4239), .dinb(n3834), .dout(n4240));
  jnot g04019(.din(n4225), .dout(n4241));
  jand g04020(.dina(n4241), .dinb(n4240), .dout(n4242));
  jor  g04021(.dina(n4242), .dinb(asqrt[63] ), .dout(n4243));
  jnot g04022(.din(n4228), .dout(n4244));
  jor  g04023(.dina(n4239), .dinb(n3834), .dout(n4245));
  jand g04024(.dina(n4245), .dinb(n4244), .dout(n4246));
  jnot g04025(.din(n4234), .dout(n4247));
  jand g04026(.dina(n4247), .dinb(n4246), .dout(n4248));
  jand g04027(.dina(n4248), .dinb(n4243), .dout(n4249));
  jxor g04028(.dina(n4113), .dinb(n221), .dout(n4250));
  jor  g04029(.dina(n4250), .dinb(n4249), .dout(n4251));
  jxor g04030(.dina(n4251), .dinb(n4219), .dout(n4252));
  jnot g04031(.din(n4252), .dout(n4253));
  jor  g04032(.dina(n4249), .dinb(n3837), .dout(n4254));
  jnot g04033(.din(a[76] ), .dout(n4255));
  jnot g04034(.din(a[77] ), .dout(n4256));
  jand g04035(.dina(n4256), .dinb(n4255), .dout(n4257));
  jand g04036(.dina(n4257), .dinb(n3837), .dout(n4258));
  jnot g04037(.din(n4258), .dout(n4259));
  jand g04038(.dina(n4259), .dinb(n4254), .dout(n4260));
  jor  g04039(.dina(n4260), .dinb(n3955), .dout(n4261));
  jand g04040(.dina(n4260), .dinb(n3955), .dout(n4262));
  jor  g04041(.dina(n4249), .dinb(a[78] ), .dout(n4263));
  jand g04042(.dina(n4263), .dinb(a[79] ), .dout(n4264));
  jand g04043(.dina(asqrt[39] ), .dinb(n3839), .dout(n4265));
  jor  g04044(.dina(n4265), .dinb(n4264), .dout(n4266));
  jor  g04045(.dina(n4266), .dinb(n4262), .dout(n4267));
  jand g04046(.dina(n4267), .dinb(n4261), .dout(n4268));
  jor  g04047(.dina(n4268), .dinb(n3642), .dout(n4269));
  jand g04048(.dina(n4268), .dinb(n3642), .dout(n4270));
  jnot g04049(.din(n3839), .dout(n4271));
  jor  g04050(.dina(n4249), .dinb(n4271), .dout(n4272));
  jor  g04051(.dina(n4229), .dinb(n3955), .dout(n4273));
  jor  g04052(.dina(n4273), .dinb(n4227), .dout(n4274));
  jor  g04053(.dina(n4274), .dinb(n4233), .dout(n4275));
  jand g04054(.dina(n4275), .dinb(n4272), .dout(n4276));
  jxor g04055(.dina(n4276), .dinb(n3648), .dout(n4277));
  jor  g04056(.dina(n4277), .dinb(n4270), .dout(n4278));
  jand g04057(.dina(n4278), .dinb(n4269), .dout(n4279));
  jor  g04058(.dina(n4279), .dinb(n3368), .dout(n4280));
  jand g04059(.dina(n4279), .dinb(n3368), .dout(n4281));
  jxor g04060(.dina(n3841), .dinb(n3642), .dout(n4282));
  jor  g04061(.dina(n4282), .dinb(n4249), .dout(n4283));
  jxor g04062(.dina(n4283), .dinb(n3957), .dout(n4284));
  jor  g04063(.dina(n4284), .dinb(n4281), .dout(n4285));
  jand g04064(.dina(n4285), .dinb(n4280), .dout(n4286));
  jor  g04065(.dina(n4286), .dinb(n3089), .dout(n4287));
  jand g04066(.dina(n4286), .dinb(n3089), .dout(n4288));
  jxor g04067(.dina(n3959), .dinb(n3368), .dout(n4289));
  jor  g04068(.dina(n4289), .dinb(n4249), .dout(n4290));
  jxor g04069(.dina(n4290), .dinb(n3968), .dout(n4291));
  jor  g04070(.dina(n4291), .dinb(n4288), .dout(n4292));
  jand g04071(.dina(n4292), .dinb(n4287), .dout(n4293));
  jor  g04072(.dina(n4293), .dinb(n2833), .dout(n4294));
  jand g04073(.dina(n4293), .dinb(n2833), .dout(n4295));
  jxor g04074(.dina(n3970), .dinb(n3089), .dout(n4296));
  jor  g04075(.dina(n4296), .dinb(n4249), .dout(n4297));
  jxor g04076(.dina(n4297), .dinb(n4150), .dout(n4298));
  jnot g04077(.din(n4298), .dout(n4299));
  jor  g04078(.dina(n4299), .dinb(n4295), .dout(n4300));
  jand g04079(.dina(n4300), .dinb(n4294), .dout(n4301));
  jor  g04080(.dina(n4301), .dinb(n2572), .dout(n4302));
  jand g04081(.dina(n4301), .dinb(n2572), .dout(n4303));
  jxor g04082(.dina(n3977), .dinb(n2833), .dout(n4304));
  jor  g04083(.dina(n4304), .dinb(n4249), .dout(n4305));
  jxor g04084(.dina(n4305), .dinb(n3983), .dout(n4306));
  jor  g04085(.dina(n4306), .dinb(n4303), .dout(n4307));
  jand g04086(.dina(n4307), .dinb(n4302), .dout(n4308));
  jor  g04087(.dina(n4308), .dinb(n2345), .dout(n4309));
  jand g04088(.dina(n4308), .dinb(n2345), .dout(n4310));
  jxor g04089(.dina(n3985), .dinb(n2572), .dout(n4311));
  jor  g04090(.dina(n4311), .dinb(n4249), .dout(n4312));
  jxor g04091(.dina(n4312), .dinb(n4157), .dout(n4313));
  jnot g04092(.din(n4313), .dout(n4314));
  jor  g04093(.dina(n4314), .dinb(n4310), .dout(n4315));
  jand g04094(.dina(n4315), .dinb(n4309), .dout(n4316));
  jor  g04095(.dina(n4316), .dinb(n2108), .dout(n4317));
  jand g04096(.dina(n4316), .dinb(n2108), .dout(n4318));
  jxor g04097(.dina(n3992), .dinb(n2345), .dout(n4319));
  jor  g04098(.dina(n4319), .dinb(n4249), .dout(n4320));
  jxor g04099(.dina(n4320), .dinb(n3998), .dout(n4321));
  jor  g04100(.dina(n4321), .dinb(n4318), .dout(n4322));
  jand g04101(.dina(n4322), .dinb(n4317), .dout(n4323));
  jor  g04102(.dina(n4323), .dinb(n1912), .dout(n4324));
  jand g04103(.dina(n4323), .dinb(n1912), .dout(n4325));
  jxor g04104(.dina(n4000), .dinb(n2108), .dout(n4326));
  jor  g04105(.dina(n4326), .dinb(n4249), .dout(n4327));
  jxor g04106(.dina(n4327), .dinb(n4164), .dout(n4328));
  jnot g04107(.din(n4328), .dout(n4329));
  jor  g04108(.dina(n4329), .dinb(n4325), .dout(n4330));
  jand g04109(.dina(n4330), .dinb(n4324), .dout(n4331));
  jor  g04110(.dina(n4331), .dinb(n1699), .dout(n4332));
  jand g04111(.dina(n4331), .dinb(n1699), .dout(n4333));
  jxor g04112(.dina(n4007), .dinb(n1912), .dout(n4334));
  jor  g04113(.dina(n4334), .dinb(n4249), .dout(n4335));
  jxor g04114(.dina(n4335), .dinb(n4168), .dout(n4336));
  jnot g04115(.din(n4336), .dout(n4337));
  jor  g04116(.dina(n4337), .dinb(n4333), .dout(n4338));
  jand g04117(.dina(n4338), .dinb(n4332), .dout(n4339));
  jor  g04118(.dina(n4339), .dinb(n1516), .dout(n4340));
  jand g04119(.dina(n4339), .dinb(n1516), .dout(n4341));
  jxor g04120(.dina(n4014), .dinb(n1699), .dout(n4342));
  jor  g04121(.dina(n4342), .dinb(n4249), .dout(n4343));
  jxor g04122(.dina(n4343), .dinb(n4020), .dout(n4344));
  jor  g04123(.dina(n4344), .dinb(n4341), .dout(n4345));
  jand g04124(.dina(n4345), .dinb(n4340), .dout(n4346));
  jor  g04125(.dina(n4346), .dinb(n1332), .dout(n4347));
  jand g04126(.dina(n4346), .dinb(n1332), .dout(n4348));
  jxor g04127(.dina(n4022), .dinb(n1516), .dout(n4349));
  jor  g04128(.dina(n4349), .dinb(n4249), .dout(n4350));
  jxor g04129(.dina(n4350), .dinb(n4028), .dout(n4351));
  jor  g04130(.dina(n4351), .dinb(n4348), .dout(n4352));
  jand g04131(.dina(n4352), .dinb(n4347), .dout(n4353));
  jor  g04132(.dina(n4353), .dinb(n1173), .dout(n4354));
  jand g04133(.dina(n4353), .dinb(n1173), .dout(n4355));
  jxor g04134(.dina(n4030), .dinb(n1332), .dout(n4356));
  jor  g04135(.dina(n4356), .dinb(n4249), .dout(n4357));
  jxor g04136(.dina(n4357), .dinb(n4178), .dout(n4358));
  jnot g04137(.din(n4358), .dout(n4359));
  jor  g04138(.dina(n4359), .dinb(n4355), .dout(n4360));
  jand g04139(.dina(n4360), .dinb(n4354), .dout(n4361));
  jor  g04140(.dina(n4361), .dinb(n1008), .dout(n4362));
  jand g04141(.dina(n4361), .dinb(n1008), .dout(n4363));
  jxor g04142(.dina(n4037), .dinb(n1173), .dout(n4364));
  jor  g04143(.dina(n4364), .dinb(n4249), .dout(n4365));
  jxor g04144(.dina(n4365), .dinb(n4043), .dout(n4366));
  jor  g04145(.dina(n4366), .dinb(n4363), .dout(n4367));
  jand g04146(.dina(n4367), .dinb(n4362), .dout(n4368));
  jor  g04147(.dina(n4368), .dinb(n884), .dout(n4369));
  jand g04148(.dina(n4368), .dinb(n884), .dout(n4370));
  jxor g04149(.dina(n4045), .dinb(n1008), .dout(n4371));
  jor  g04150(.dina(n4371), .dinb(n4249), .dout(n4372));
  jxor g04151(.dina(n4372), .dinb(n4185), .dout(n4373));
  jnot g04152(.din(n4373), .dout(n4374));
  jor  g04153(.dina(n4374), .dinb(n4370), .dout(n4375));
  jand g04154(.dina(n4375), .dinb(n4369), .dout(n4376));
  jor  g04155(.dina(n4376), .dinb(n743), .dout(n4377));
  jand g04156(.dina(n4376), .dinb(n743), .dout(n4378));
  jxor g04157(.dina(n4052), .dinb(n884), .dout(n4379));
  jor  g04158(.dina(n4379), .dinb(n4249), .dout(n4380));
  jxor g04159(.dina(n4380), .dinb(n4058), .dout(n4381));
  jor  g04160(.dina(n4381), .dinb(n4378), .dout(n4382));
  jand g04161(.dina(n4382), .dinb(n4377), .dout(n4383));
  jor  g04162(.dina(n4383), .dinb(n635), .dout(n4384));
  jand g04163(.dina(n4383), .dinb(n635), .dout(n4385));
  jxor g04164(.dina(n4060), .dinb(n743), .dout(n4386));
  jor  g04165(.dina(n4386), .dinb(n4249), .dout(n4387));
  jxor g04166(.dina(n4387), .dinb(n4192), .dout(n4388));
  jnot g04167(.din(n4388), .dout(n4389));
  jor  g04168(.dina(n4389), .dinb(n4385), .dout(n4390));
  jand g04169(.dina(n4390), .dinb(n4384), .dout(n4391));
  jor  g04170(.dina(n4391), .dinb(n515), .dout(n4392));
  jand g04171(.dina(n4391), .dinb(n515), .dout(n4393));
  jxor g04172(.dina(n4067), .dinb(n635), .dout(n4394));
  jor  g04173(.dina(n4394), .dinb(n4249), .dout(n4395));
  jxor g04174(.dina(n4395), .dinb(n4073), .dout(n4396));
  jor  g04175(.dina(n4396), .dinb(n4393), .dout(n4397));
  jand g04176(.dina(n4397), .dinb(n4392), .dout(n4398));
  jor  g04177(.dina(n4398), .dinb(n443), .dout(n4399));
  jand g04178(.dina(n4398), .dinb(n443), .dout(n4400));
  jxor g04179(.dina(n4075), .dinb(n515), .dout(n4401));
  jor  g04180(.dina(n4401), .dinb(n4249), .dout(n4402));
  jxor g04181(.dina(n4402), .dinb(n4199), .dout(n4403));
  jnot g04182(.din(n4403), .dout(n4404));
  jor  g04183(.dina(n4404), .dinb(n4400), .dout(n4405));
  jand g04184(.dina(n4405), .dinb(n4399), .dout(n4406));
  jor  g04185(.dina(n4406), .dinb(n352), .dout(n4407));
  jand g04186(.dina(n4406), .dinb(n352), .dout(n4408));
  jxor g04187(.dina(n4082), .dinb(n443), .dout(n4409));
  jor  g04188(.dina(n4409), .dinb(n4249), .dout(n4410));
  jxor g04189(.dina(n4410), .dinb(n4088), .dout(n4411));
  jor  g04190(.dina(n4411), .dinb(n4408), .dout(n4412));
  jand g04191(.dina(n4412), .dinb(n4407), .dout(n4413));
  jor  g04192(.dina(n4413), .dinb(n294), .dout(n4414));
  jand g04193(.dina(n4413), .dinb(n294), .dout(n4415));
  jxor g04194(.dina(n4090), .dinb(n352), .dout(n4416));
  jor  g04195(.dina(n4416), .dinb(n4249), .dout(n4417));
  jxor g04196(.dina(n4417), .dinb(n4206), .dout(n4418));
  jnot g04197(.din(n4418), .dout(n4419));
  jor  g04198(.dina(n4419), .dinb(n4415), .dout(n4420));
  jand g04199(.dina(n4420), .dinb(n4414), .dout(n4421));
  jor  g04200(.dina(n4421), .dinb(n239), .dout(n4422));
  jand g04201(.dina(n4421), .dinb(n239), .dout(n4423));
  jxor g04202(.dina(n4097), .dinb(n294), .dout(n4424));
  jor  g04203(.dina(n4424), .dinb(n4249), .dout(n4425));
  jxor g04204(.dina(n4425), .dinb(n4103), .dout(n4426));
  jor  g04205(.dina(n4426), .dinb(n4423), .dout(n4427));
  jand g04206(.dina(n4427), .dinb(n4422), .dout(n4428));
  jor  g04207(.dina(n4428), .dinb(n221), .dout(n4429));
  jand g04208(.dina(n4428), .dinb(n221), .dout(n4430));
  jxor g04209(.dina(n4105), .dinb(n239), .dout(n4431));
  jor  g04210(.dina(n4431), .dinb(n4249), .dout(n4432));
  jxor g04211(.dina(n4432), .dinb(n4111), .dout(n4433));
  jor  g04212(.dina(n4433), .dinb(n4430), .dout(n4434));
  jand g04213(.dina(n4434), .dinb(n4429), .dout(n4435));
  jor  g04214(.dina(n4435), .dinb(n4253), .dout(n4436));
  jand g04215(.dina(asqrt[39] ), .dinb(n4240), .dout(n4437));
  jor  g04216(.dina(n4437), .dinb(n4436), .dout(n4438));
  jor  g04217(.dina(n4438), .dinb(n4229), .dout(n4439));
  jand g04218(.dina(n4439), .dinb(n218), .dout(n4440));
  jand g04219(.dina(n4249), .dinb(n3835), .dout(n4441));
  jand g04220(.dina(n4435), .dinb(n4253), .dout(n4442));
  jor  g04221(.dina(n4442), .dinb(n4441), .dout(n4443));
  jand g04222(.dina(n4249), .dinb(n4221), .dout(n4444));
  jand g04223(.dina(n4222), .dinb(asqrt[63] ), .dout(n4445));
  jand g04224(.dina(n4445), .dinb(n4245), .dout(n4446));
  jnot g04225(.din(n4446), .dout(n4447));
  jor  g04226(.dina(n4447), .dinb(n4444), .dout(n4448));
  jnot g04227(.din(n4448), .dout(n4449));
  jor  g04228(.dina(n4449), .dinb(n4443), .dout(n4450));
  jor  g04229(.dina(n4450), .dinb(n4440), .dout(asqrt[38] ));
  jnot g04230(.din(n4433), .dout(n4452));
  jxor g04231(.dina(n4428), .dinb(n221), .dout(n4453));
  jand g04232(.dina(n4453), .dinb(asqrt[38] ), .dout(n4454));
  jxor g04233(.dina(n4454), .dinb(n4452), .dout(n4455));
  jand g04234(.dina(asqrt[38] ), .dinb(a[76] ), .dout(n4456));
  jnot g04235(.din(a[74] ), .dout(n4457));
  jnot g04236(.din(a[75] ), .dout(n4458));
  jand g04237(.dina(n4458), .dinb(n4457), .dout(n4459));
  jand g04238(.dina(n4459), .dinb(n4255), .dout(n4460));
  jor  g04239(.dina(n4460), .dinb(n4456), .dout(n4461));
  jand g04240(.dina(n4461), .dinb(asqrt[39] ), .dout(n4462));
  jor  g04241(.dina(n4461), .dinb(asqrt[39] ), .dout(n4463));
  jand g04242(.dina(asqrt[38] ), .dinb(n4255), .dout(n4464));
  jor  g04243(.dina(n4464), .dinb(n4256), .dout(n4465));
  jnot g04244(.din(n4257), .dout(n4466));
  jnot g04245(.din(n4429), .dout(n4467));
  jnot g04246(.din(n4422), .dout(n4468));
  jnot g04247(.din(n4414), .dout(n4469));
  jnot g04248(.din(n4407), .dout(n4470));
  jnot g04249(.din(n4399), .dout(n4471));
  jnot g04250(.din(n4392), .dout(n4472));
  jnot g04251(.din(n4384), .dout(n4473));
  jnot g04252(.din(n4377), .dout(n4474));
  jnot g04253(.din(n4369), .dout(n4475));
  jnot g04254(.din(n4362), .dout(n4476));
  jnot g04255(.din(n4354), .dout(n4477));
  jnot g04256(.din(n4347), .dout(n4478));
  jnot g04257(.din(n4340), .dout(n4479));
  jnot g04258(.din(n4332), .dout(n4480));
  jnot g04259(.din(n4324), .dout(n4481));
  jnot g04260(.din(n4317), .dout(n4482));
  jnot g04261(.din(n4309), .dout(n4483));
  jnot g04262(.din(n4302), .dout(n4484));
  jnot g04263(.din(n4294), .dout(n4485));
  jnot g04264(.din(n4287), .dout(n4486));
  jnot g04265(.din(n4280), .dout(n4487));
  jnot g04266(.din(n4269), .dout(n4488));
  jnot g04267(.din(n4261), .dout(n4489));
  jand g04268(.dina(asqrt[39] ), .dinb(a[78] ), .dout(n4490));
  jor  g04269(.dina(n4258), .dinb(n4490), .dout(n4491));
  jor  g04270(.dina(n4491), .dinb(asqrt[40] ), .dout(n4492));
  jand g04271(.dina(asqrt[39] ), .dinb(n3837), .dout(n4493));
  jor  g04272(.dina(n4493), .dinb(n3838), .dout(n4494));
  jand g04273(.dina(n4272), .dinb(n4494), .dout(n4495));
  jand g04274(.dina(n4495), .dinb(n4492), .dout(n4496));
  jor  g04275(.dina(n4496), .dinb(n4489), .dout(n4497));
  jor  g04276(.dina(n4497), .dinb(asqrt[41] ), .dout(n4498));
  jnot g04277(.din(n4277), .dout(n4499));
  jand g04278(.dina(n4499), .dinb(n4498), .dout(n4500));
  jor  g04279(.dina(n4500), .dinb(n4488), .dout(n4501));
  jor  g04280(.dina(n4501), .dinb(asqrt[42] ), .dout(n4502));
  jnot g04281(.din(n4284), .dout(n4503));
  jand g04282(.dina(n4503), .dinb(n4502), .dout(n4504));
  jor  g04283(.dina(n4504), .dinb(n4487), .dout(n4505));
  jor  g04284(.dina(n4505), .dinb(asqrt[43] ), .dout(n4506));
  jnot g04285(.din(n4291), .dout(n4507));
  jand g04286(.dina(n4507), .dinb(n4506), .dout(n4508));
  jor  g04287(.dina(n4508), .dinb(n4486), .dout(n4509));
  jor  g04288(.dina(n4509), .dinb(asqrt[44] ), .dout(n4510));
  jand g04289(.dina(n4298), .dinb(n4510), .dout(n4511));
  jor  g04290(.dina(n4511), .dinb(n4485), .dout(n4512));
  jor  g04291(.dina(n4512), .dinb(asqrt[45] ), .dout(n4513));
  jnot g04292(.din(n4306), .dout(n4514));
  jand g04293(.dina(n4514), .dinb(n4513), .dout(n4515));
  jor  g04294(.dina(n4515), .dinb(n4484), .dout(n4516));
  jor  g04295(.dina(n4516), .dinb(asqrt[46] ), .dout(n4517));
  jand g04296(.dina(n4313), .dinb(n4517), .dout(n4518));
  jor  g04297(.dina(n4518), .dinb(n4483), .dout(n4519));
  jor  g04298(.dina(n4519), .dinb(asqrt[47] ), .dout(n4520));
  jnot g04299(.din(n4321), .dout(n4521));
  jand g04300(.dina(n4521), .dinb(n4520), .dout(n4522));
  jor  g04301(.dina(n4522), .dinb(n4482), .dout(n4523));
  jor  g04302(.dina(n4523), .dinb(asqrt[48] ), .dout(n4524));
  jand g04303(.dina(n4328), .dinb(n4524), .dout(n4525));
  jor  g04304(.dina(n4525), .dinb(n4481), .dout(n4526));
  jor  g04305(.dina(n4526), .dinb(asqrt[49] ), .dout(n4527));
  jand g04306(.dina(n4336), .dinb(n4527), .dout(n4528));
  jor  g04307(.dina(n4528), .dinb(n4480), .dout(n4529));
  jor  g04308(.dina(n4529), .dinb(asqrt[50] ), .dout(n4530));
  jnot g04309(.din(n4344), .dout(n4531));
  jand g04310(.dina(n4531), .dinb(n4530), .dout(n4532));
  jor  g04311(.dina(n4532), .dinb(n4479), .dout(n4533));
  jor  g04312(.dina(n4533), .dinb(asqrt[51] ), .dout(n4534));
  jnot g04313(.din(n4351), .dout(n4535));
  jand g04314(.dina(n4535), .dinb(n4534), .dout(n4536));
  jor  g04315(.dina(n4536), .dinb(n4478), .dout(n4537));
  jor  g04316(.dina(n4537), .dinb(asqrt[52] ), .dout(n4538));
  jand g04317(.dina(n4358), .dinb(n4538), .dout(n4539));
  jor  g04318(.dina(n4539), .dinb(n4477), .dout(n4540));
  jor  g04319(.dina(n4540), .dinb(asqrt[53] ), .dout(n4541));
  jnot g04320(.din(n4366), .dout(n4542));
  jand g04321(.dina(n4542), .dinb(n4541), .dout(n4543));
  jor  g04322(.dina(n4543), .dinb(n4476), .dout(n4544));
  jor  g04323(.dina(n4544), .dinb(asqrt[54] ), .dout(n4545));
  jand g04324(.dina(n4373), .dinb(n4545), .dout(n4546));
  jor  g04325(.dina(n4546), .dinb(n4475), .dout(n4547));
  jor  g04326(.dina(n4547), .dinb(asqrt[55] ), .dout(n4548));
  jnot g04327(.din(n4381), .dout(n4549));
  jand g04328(.dina(n4549), .dinb(n4548), .dout(n4550));
  jor  g04329(.dina(n4550), .dinb(n4474), .dout(n4551));
  jor  g04330(.dina(n4551), .dinb(asqrt[56] ), .dout(n4552));
  jand g04331(.dina(n4388), .dinb(n4552), .dout(n4553));
  jor  g04332(.dina(n4553), .dinb(n4473), .dout(n4554));
  jor  g04333(.dina(n4554), .dinb(asqrt[57] ), .dout(n4555));
  jnot g04334(.din(n4396), .dout(n4556));
  jand g04335(.dina(n4556), .dinb(n4555), .dout(n4557));
  jor  g04336(.dina(n4557), .dinb(n4472), .dout(n4558));
  jor  g04337(.dina(n4558), .dinb(asqrt[58] ), .dout(n4559));
  jand g04338(.dina(n4403), .dinb(n4559), .dout(n4560));
  jor  g04339(.dina(n4560), .dinb(n4471), .dout(n4561));
  jor  g04340(.dina(n4561), .dinb(asqrt[59] ), .dout(n4562));
  jnot g04341(.din(n4411), .dout(n4563));
  jand g04342(.dina(n4563), .dinb(n4562), .dout(n4564));
  jor  g04343(.dina(n4564), .dinb(n4470), .dout(n4565));
  jor  g04344(.dina(n4565), .dinb(asqrt[60] ), .dout(n4566));
  jand g04345(.dina(n4418), .dinb(n4566), .dout(n4567));
  jor  g04346(.dina(n4567), .dinb(n4469), .dout(n4568));
  jor  g04347(.dina(n4568), .dinb(asqrt[61] ), .dout(n4569));
  jnot g04348(.din(n4426), .dout(n4570));
  jand g04349(.dina(n4570), .dinb(n4569), .dout(n4571));
  jor  g04350(.dina(n4571), .dinb(n4468), .dout(n4572));
  jor  g04351(.dina(n4572), .dinb(asqrt[62] ), .dout(n4573));
  jand g04352(.dina(n4452), .dinb(n4573), .dout(n4574));
  jor  g04353(.dina(n4574), .dinb(n4467), .dout(n4575));
  jand g04354(.dina(n4575), .dinb(n4252), .dout(n4576));
  jnot g04355(.din(n4437), .dout(n4577));
  jand g04356(.dina(n4577), .dinb(n4576), .dout(n4578));
  jand g04357(.dina(n4578), .dinb(n4245), .dout(n4579));
  jor  g04358(.dina(n4579), .dinb(asqrt[63] ), .dout(n4580));
  jnot g04359(.din(n4450), .dout(n4581));
  jand g04360(.dina(n4581), .dinb(n4580), .dout(n4582));
  jor  g04361(.dina(n4582), .dinb(n4466), .dout(n4583));
  jand g04362(.dina(n4583), .dinb(n4465), .dout(n4584));
  jand g04363(.dina(n4584), .dinb(n4463), .dout(n4585));
  jor  g04364(.dina(n4585), .dinb(n4462), .dout(n4586));
  jand g04365(.dina(n4586), .dinb(asqrt[40] ), .dout(n4587));
  jor  g04366(.dina(n4586), .dinb(asqrt[40] ), .dout(n4588));
  jand g04367(.dina(asqrt[38] ), .dinb(n4257), .dout(n4589));
  jnot g04368(.din(n4442), .dout(n4590));
  jand g04369(.dina(n4447), .dinb(asqrt[39] ), .dout(n4591));
  jand g04370(.dina(n4591), .dinb(n4590), .dout(n4592));
  jand g04371(.dina(n4592), .dinb(n4580), .dout(n4593));
  jor  g04372(.dina(n4593), .dinb(n4589), .dout(n4594));
  jxor g04373(.dina(n4594), .dinb(a[78] ), .dout(n4595));
  jnot g04374(.din(n4595), .dout(n4596));
  jand g04375(.dina(n4596), .dinb(n4588), .dout(n4597));
  jor  g04376(.dina(n4597), .dinb(n4587), .dout(n4598));
  jand g04377(.dina(n4598), .dinb(asqrt[41] ), .dout(n4599));
  jor  g04378(.dina(n4598), .dinb(asqrt[41] ), .dout(n4600));
  jxor g04379(.dina(n4260), .dinb(n3955), .dout(n4601));
  jand g04380(.dina(n4601), .dinb(asqrt[38] ), .dout(n4602));
  jxor g04381(.dina(n4602), .dinb(n4266), .dout(n4603));
  jnot g04382(.din(n4603), .dout(n4604));
  jand g04383(.dina(n4604), .dinb(n4600), .dout(n4605));
  jor  g04384(.dina(n4605), .dinb(n4599), .dout(n4606));
  jand g04385(.dina(n4606), .dinb(asqrt[42] ), .dout(n4607));
  jor  g04386(.dina(n4606), .dinb(asqrt[42] ), .dout(n4608));
  jxor g04387(.dina(n4268), .dinb(n3642), .dout(n4609));
  jand g04388(.dina(n4609), .dinb(asqrt[38] ), .dout(n4610));
  jxor g04389(.dina(n4610), .dinb(n4277), .dout(n4611));
  jnot g04390(.din(n4611), .dout(n4612));
  jand g04391(.dina(n4612), .dinb(n4608), .dout(n4613));
  jor  g04392(.dina(n4613), .dinb(n4607), .dout(n4614));
  jand g04393(.dina(n4614), .dinb(asqrt[43] ), .dout(n4615));
  jor  g04394(.dina(n4614), .dinb(asqrt[43] ), .dout(n4616));
  jxor g04395(.dina(n4279), .dinb(n3368), .dout(n4617));
  jand g04396(.dina(n4617), .dinb(asqrt[38] ), .dout(n4618));
  jxor g04397(.dina(n4618), .dinb(n4284), .dout(n4619));
  jnot g04398(.din(n4619), .dout(n4620));
  jand g04399(.dina(n4620), .dinb(n4616), .dout(n4621));
  jor  g04400(.dina(n4621), .dinb(n4615), .dout(n4622));
  jand g04401(.dina(n4622), .dinb(asqrt[44] ), .dout(n4623));
  jor  g04402(.dina(n4622), .dinb(asqrt[44] ), .dout(n4624));
  jxor g04403(.dina(n4286), .dinb(n3089), .dout(n4625));
  jand g04404(.dina(n4625), .dinb(asqrt[38] ), .dout(n4626));
  jxor g04405(.dina(n4626), .dinb(n4291), .dout(n4627));
  jnot g04406(.din(n4627), .dout(n4628));
  jand g04407(.dina(n4628), .dinb(n4624), .dout(n4629));
  jor  g04408(.dina(n4629), .dinb(n4623), .dout(n4630));
  jand g04409(.dina(n4630), .dinb(asqrt[45] ), .dout(n4631));
  jor  g04410(.dina(n4630), .dinb(asqrt[45] ), .dout(n4632));
  jxor g04411(.dina(n4293), .dinb(n2833), .dout(n4633));
  jand g04412(.dina(n4633), .dinb(asqrt[38] ), .dout(n4634));
  jxor g04413(.dina(n4634), .dinb(n4298), .dout(n4635));
  jand g04414(.dina(n4635), .dinb(n4632), .dout(n4636));
  jor  g04415(.dina(n4636), .dinb(n4631), .dout(n4637));
  jand g04416(.dina(n4637), .dinb(asqrt[46] ), .dout(n4638));
  jor  g04417(.dina(n4637), .dinb(asqrt[46] ), .dout(n4639));
  jxor g04418(.dina(n4301), .dinb(n2572), .dout(n4640));
  jand g04419(.dina(n4640), .dinb(asqrt[38] ), .dout(n4641));
  jxor g04420(.dina(n4641), .dinb(n4306), .dout(n4642));
  jnot g04421(.din(n4642), .dout(n4643));
  jand g04422(.dina(n4643), .dinb(n4639), .dout(n4644));
  jor  g04423(.dina(n4644), .dinb(n4638), .dout(n4645));
  jand g04424(.dina(n4645), .dinb(asqrt[47] ), .dout(n4646));
  jor  g04425(.dina(n4645), .dinb(asqrt[47] ), .dout(n4647));
  jxor g04426(.dina(n4308), .dinb(n2345), .dout(n4648));
  jand g04427(.dina(n4648), .dinb(asqrt[38] ), .dout(n4649));
  jxor g04428(.dina(n4649), .dinb(n4313), .dout(n4650));
  jand g04429(.dina(n4650), .dinb(n4647), .dout(n4651));
  jor  g04430(.dina(n4651), .dinb(n4646), .dout(n4652));
  jand g04431(.dina(n4652), .dinb(asqrt[48] ), .dout(n4653));
  jor  g04432(.dina(n4652), .dinb(asqrt[48] ), .dout(n4654));
  jxor g04433(.dina(n4316), .dinb(n2108), .dout(n4655));
  jand g04434(.dina(n4655), .dinb(asqrt[38] ), .dout(n4656));
  jxor g04435(.dina(n4656), .dinb(n4321), .dout(n4657));
  jnot g04436(.din(n4657), .dout(n4658));
  jand g04437(.dina(n4658), .dinb(n4654), .dout(n4659));
  jor  g04438(.dina(n4659), .dinb(n4653), .dout(n4660));
  jand g04439(.dina(n4660), .dinb(asqrt[49] ), .dout(n4661));
  jor  g04440(.dina(n4660), .dinb(asqrt[49] ), .dout(n4662));
  jxor g04441(.dina(n4323), .dinb(n1912), .dout(n4663));
  jand g04442(.dina(n4663), .dinb(asqrt[38] ), .dout(n4664));
  jxor g04443(.dina(n4664), .dinb(n4328), .dout(n4665));
  jand g04444(.dina(n4665), .dinb(n4662), .dout(n4666));
  jor  g04445(.dina(n4666), .dinb(n4661), .dout(n4667));
  jand g04446(.dina(n4667), .dinb(asqrt[50] ), .dout(n4668));
  jor  g04447(.dina(n4667), .dinb(asqrt[50] ), .dout(n4669));
  jxor g04448(.dina(n4331), .dinb(n1699), .dout(n4670));
  jand g04449(.dina(n4670), .dinb(asqrt[38] ), .dout(n4671));
  jxor g04450(.dina(n4671), .dinb(n4336), .dout(n4672));
  jand g04451(.dina(n4672), .dinb(n4669), .dout(n4673));
  jor  g04452(.dina(n4673), .dinb(n4668), .dout(n4674));
  jand g04453(.dina(n4674), .dinb(asqrt[51] ), .dout(n4675));
  jor  g04454(.dina(n4674), .dinb(asqrt[51] ), .dout(n4676));
  jxor g04455(.dina(n4339), .dinb(n1516), .dout(n4677));
  jand g04456(.dina(n4677), .dinb(asqrt[38] ), .dout(n4678));
  jxor g04457(.dina(n4678), .dinb(n4344), .dout(n4679));
  jnot g04458(.din(n4679), .dout(n4680));
  jand g04459(.dina(n4680), .dinb(n4676), .dout(n4681));
  jor  g04460(.dina(n4681), .dinb(n4675), .dout(n4682));
  jand g04461(.dina(n4682), .dinb(asqrt[52] ), .dout(n4683));
  jor  g04462(.dina(n4682), .dinb(asqrt[52] ), .dout(n4684));
  jxor g04463(.dina(n4346), .dinb(n1332), .dout(n4685));
  jand g04464(.dina(n4685), .dinb(asqrt[38] ), .dout(n4686));
  jxor g04465(.dina(n4686), .dinb(n4351), .dout(n4687));
  jnot g04466(.din(n4687), .dout(n4688));
  jand g04467(.dina(n4688), .dinb(n4684), .dout(n4689));
  jor  g04468(.dina(n4689), .dinb(n4683), .dout(n4690));
  jand g04469(.dina(n4690), .dinb(asqrt[53] ), .dout(n4691));
  jor  g04470(.dina(n4690), .dinb(asqrt[53] ), .dout(n4692));
  jxor g04471(.dina(n4353), .dinb(n1173), .dout(n4693));
  jand g04472(.dina(n4693), .dinb(asqrt[38] ), .dout(n4694));
  jxor g04473(.dina(n4694), .dinb(n4358), .dout(n4695));
  jand g04474(.dina(n4695), .dinb(n4692), .dout(n4696));
  jor  g04475(.dina(n4696), .dinb(n4691), .dout(n4697));
  jand g04476(.dina(n4697), .dinb(asqrt[54] ), .dout(n4698));
  jor  g04477(.dina(n4697), .dinb(asqrt[54] ), .dout(n4699));
  jxor g04478(.dina(n4361), .dinb(n1008), .dout(n4700));
  jand g04479(.dina(n4700), .dinb(asqrt[38] ), .dout(n4701));
  jxor g04480(.dina(n4701), .dinb(n4366), .dout(n4702));
  jnot g04481(.din(n4702), .dout(n4703));
  jand g04482(.dina(n4703), .dinb(n4699), .dout(n4704));
  jor  g04483(.dina(n4704), .dinb(n4698), .dout(n4705));
  jand g04484(.dina(n4705), .dinb(asqrt[55] ), .dout(n4706));
  jor  g04485(.dina(n4705), .dinb(asqrt[55] ), .dout(n4707));
  jxor g04486(.dina(n4368), .dinb(n884), .dout(n4708));
  jand g04487(.dina(n4708), .dinb(asqrt[38] ), .dout(n4709));
  jxor g04488(.dina(n4709), .dinb(n4373), .dout(n4710));
  jand g04489(.dina(n4710), .dinb(n4707), .dout(n4711));
  jor  g04490(.dina(n4711), .dinb(n4706), .dout(n4712));
  jand g04491(.dina(n4712), .dinb(asqrt[56] ), .dout(n4713));
  jor  g04492(.dina(n4712), .dinb(asqrt[56] ), .dout(n4714));
  jxor g04493(.dina(n4376), .dinb(n743), .dout(n4715));
  jand g04494(.dina(n4715), .dinb(asqrt[38] ), .dout(n4716));
  jxor g04495(.dina(n4716), .dinb(n4381), .dout(n4717));
  jnot g04496(.din(n4717), .dout(n4718));
  jand g04497(.dina(n4718), .dinb(n4714), .dout(n4719));
  jor  g04498(.dina(n4719), .dinb(n4713), .dout(n4720));
  jand g04499(.dina(n4720), .dinb(asqrt[57] ), .dout(n4721));
  jor  g04500(.dina(n4720), .dinb(asqrt[57] ), .dout(n4722));
  jxor g04501(.dina(n4383), .dinb(n635), .dout(n4723));
  jand g04502(.dina(n4723), .dinb(asqrt[38] ), .dout(n4724));
  jxor g04503(.dina(n4724), .dinb(n4388), .dout(n4725));
  jand g04504(.dina(n4725), .dinb(n4722), .dout(n4726));
  jor  g04505(.dina(n4726), .dinb(n4721), .dout(n4727));
  jand g04506(.dina(n4727), .dinb(asqrt[58] ), .dout(n4728));
  jor  g04507(.dina(n4727), .dinb(asqrt[58] ), .dout(n4729));
  jxor g04508(.dina(n4391), .dinb(n515), .dout(n4730));
  jand g04509(.dina(n4730), .dinb(asqrt[38] ), .dout(n4731));
  jxor g04510(.dina(n4731), .dinb(n4396), .dout(n4732));
  jnot g04511(.din(n4732), .dout(n4733));
  jand g04512(.dina(n4733), .dinb(n4729), .dout(n4734));
  jor  g04513(.dina(n4734), .dinb(n4728), .dout(n4735));
  jand g04514(.dina(n4735), .dinb(asqrt[59] ), .dout(n4736));
  jor  g04515(.dina(n4735), .dinb(asqrt[59] ), .dout(n4737));
  jxor g04516(.dina(n4398), .dinb(n443), .dout(n4738));
  jand g04517(.dina(n4738), .dinb(asqrt[38] ), .dout(n4739));
  jxor g04518(.dina(n4739), .dinb(n4403), .dout(n4740));
  jand g04519(.dina(n4740), .dinb(n4737), .dout(n4741));
  jor  g04520(.dina(n4741), .dinb(n4736), .dout(n4742));
  jand g04521(.dina(n4742), .dinb(asqrt[60] ), .dout(n4743));
  jor  g04522(.dina(n4742), .dinb(asqrt[60] ), .dout(n4744));
  jxor g04523(.dina(n4406), .dinb(n352), .dout(n4745));
  jand g04524(.dina(n4745), .dinb(asqrt[38] ), .dout(n4746));
  jxor g04525(.dina(n4746), .dinb(n4411), .dout(n4747));
  jnot g04526(.din(n4747), .dout(n4748));
  jand g04527(.dina(n4748), .dinb(n4744), .dout(n4749));
  jor  g04528(.dina(n4749), .dinb(n4743), .dout(n4750));
  jand g04529(.dina(n4750), .dinb(asqrt[61] ), .dout(n4751));
  jor  g04530(.dina(n4750), .dinb(asqrt[61] ), .dout(n4752));
  jxor g04531(.dina(n4413), .dinb(n294), .dout(n4753));
  jand g04532(.dina(n4753), .dinb(asqrt[38] ), .dout(n4754));
  jxor g04533(.dina(n4754), .dinb(n4418), .dout(n4755));
  jand g04534(.dina(n4755), .dinb(n4752), .dout(n4756));
  jor  g04535(.dina(n4756), .dinb(n4751), .dout(n4757));
  jand g04536(.dina(n4757), .dinb(asqrt[62] ), .dout(n4758));
  jor  g04537(.dina(n4757), .dinb(asqrt[62] ), .dout(n4759));
  jxor g04538(.dina(n4421), .dinb(n239), .dout(n4760));
  jand g04539(.dina(n4760), .dinb(asqrt[38] ), .dout(n4761));
  jxor g04540(.dina(n4761), .dinb(n4426), .dout(n4762));
  jnot g04541(.din(n4762), .dout(n4763));
  jand g04542(.dina(n4763), .dinb(n4759), .dout(n4764));
  jor  g04543(.dina(n4764), .dinb(n4758), .dout(n4765));
  jor  g04544(.dina(n4765), .dinb(n4455), .dout(n4766));
  jnot g04545(.din(n4766), .dout(n4767));
  jand g04546(.dina(n4582), .dinb(n4435), .dout(n4768));
  jnot g04547(.din(n4768), .dout(n4769));
  jand g04548(.dina(n4436), .dinb(asqrt[63] ), .dout(n4770));
  jand g04549(.dina(n4770), .dinb(n4590), .dout(n4771));
  jand g04550(.dina(n4771), .dinb(n4769), .dout(n4772));
  jnot g04551(.din(n4455), .dout(n4773));
  jnot g04552(.din(n4758), .dout(n4774));
  jnot g04553(.din(n4751), .dout(n4775));
  jnot g04554(.din(n4743), .dout(n4776));
  jnot g04555(.din(n4736), .dout(n4777));
  jnot g04556(.din(n4728), .dout(n4778));
  jnot g04557(.din(n4721), .dout(n4779));
  jnot g04558(.din(n4713), .dout(n4780));
  jnot g04559(.din(n4706), .dout(n4781));
  jnot g04560(.din(n4698), .dout(n4782));
  jnot g04561(.din(n4691), .dout(n4783));
  jnot g04562(.din(n4683), .dout(n4784));
  jnot g04563(.din(n4675), .dout(n4785));
  jnot g04564(.din(n4668), .dout(n4786));
  jnot g04565(.din(n4661), .dout(n4787));
  jnot g04566(.din(n4653), .dout(n4788));
  jnot g04567(.din(n4646), .dout(n4789));
  jnot g04568(.din(n4638), .dout(n4790));
  jnot g04569(.din(n4631), .dout(n4791));
  jnot g04570(.din(n4623), .dout(n4792));
  jnot g04571(.din(n4615), .dout(n4793));
  jnot g04572(.din(n4607), .dout(n4794));
  jnot g04573(.din(n4599), .dout(n4795));
  jnot g04574(.din(n4587), .dout(n4796));
  jnot g04575(.din(n4462), .dout(n4797));
  jor  g04576(.dina(n4582), .dinb(n4255), .dout(n4798));
  jnot g04577(.din(n4460), .dout(n4799));
  jand g04578(.dina(n4799), .dinb(n4798), .dout(n4800));
  jand g04579(.dina(n4800), .dinb(n4249), .dout(n4801));
  jor  g04580(.dina(n4582), .dinb(a[76] ), .dout(n4802));
  jand g04581(.dina(n4802), .dinb(a[77] ), .dout(n4803));
  jor  g04582(.dina(n4589), .dinb(n4803), .dout(n4804));
  jor  g04583(.dina(n4804), .dinb(n4801), .dout(n4805));
  jand g04584(.dina(n4805), .dinb(n4797), .dout(n4806));
  jand g04585(.dina(n4806), .dinb(n3955), .dout(n4807));
  jor  g04586(.dina(n4595), .dinb(n4807), .dout(n4808));
  jand g04587(.dina(n4808), .dinb(n4796), .dout(n4809));
  jand g04588(.dina(n4809), .dinb(n3642), .dout(n4810));
  jor  g04589(.dina(n4603), .dinb(n4810), .dout(n4811));
  jand g04590(.dina(n4811), .dinb(n4795), .dout(n4812));
  jand g04591(.dina(n4812), .dinb(n3368), .dout(n4813));
  jor  g04592(.dina(n4611), .dinb(n4813), .dout(n4814));
  jand g04593(.dina(n4814), .dinb(n4794), .dout(n4815));
  jand g04594(.dina(n4815), .dinb(n3089), .dout(n4816));
  jor  g04595(.dina(n4619), .dinb(n4816), .dout(n4817));
  jand g04596(.dina(n4817), .dinb(n4793), .dout(n4818));
  jand g04597(.dina(n4818), .dinb(n2833), .dout(n4819));
  jor  g04598(.dina(n4627), .dinb(n4819), .dout(n4820));
  jand g04599(.dina(n4820), .dinb(n4792), .dout(n4821));
  jand g04600(.dina(n4821), .dinb(n2572), .dout(n4822));
  jnot g04601(.din(n4635), .dout(n4823));
  jor  g04602(.dina(n4823), .dinb(n4822), .dout(n4824));
  jand g04603(.dina(n4824), .dinb(n4791), .dout(n4825));
  jand g04604(.dina(n4825), .dinb(n2345), .dout(n4826));
  jor  g04605(.dina(n4642), .dinb(n4826), .dout(n4827));
  jand g04606(.dina(n4827), .dinb(n4790), .dout(n4828));
  jand g04607(.dina(n4828), .dinb(n2108), .dout(n4829));
  jnot g04608(.din(n4650), .dout(n4830));
  jor  g04609(.dina(n4830), .dinb(n4829), .dout(n4831));
  jand g04610(.dina(n4831), .dinb(n4789), .dout(n4832));
  jand g04611(.dina(n4832), .dinb(n1912), .dout(n4833));
  jor  g04612(.dina(n4657), .dinb(n4833), .dout(n4834));
  jand g04613(.dina(n4834), .dinb(n4788), .dout(n4835));
  jand g04614(.dina(n4835), .dinb(n1699), .dout(n4836));
  jnot g04615(.din(n4665), .dout(n4837));
  jor  g04616(.dina(n4837), .dinb(n4836), .dout(n4838));
  jand g04617(.dina(n4838), .dinb(n4787), .dout(n4839));
  jand g04618(.dina(n4839), .dinb(n1516), .dout(n4840));
  jnot g04619(.din(n4672), .dout(n4841));
  jor  g04620(.dina(n4841), .dinb(n4840), .dout(n4842));
  jand g04621(.dina(n4842), .dinb(n4786), .dout(n4843));
  jand g04622(.dina(n4843), .dinb(n1332), .dout(n4844));
  jor  g04623(.dina(n4679), .dinb(n4844), .dout(n4845));
  jand g04624(.dina(n4845), .dinb(n4785), .dout(n4846));
  jand g04625(.dina(n4846), .dinb(n1173), .dout(n4847));
  jor  g04626(.dina(n4687), .dinb(n4847), .dout(n4848));
  jand g04627(.dina(n4848), .dinb(n4784), .dout(n4849));
  jand g04628(.dina(n4849), .dinb(n1008), .dout(n4850));
  jnot g04629(.din(n4695), .dout(n4851));
  jor  g04630(.dina(n4851), .dinb(n4850), .dout(n4852));
  jand g04631(.dina(n4852), .dinb(n4783), .dout(n4853));
  jand g04632(.dina(n4853), .dinb(n884), .dout(n4854));
  jor  g04633(.dina(n4702), .dinb(n4854), .dout(n4855));
  jand g04634(.dina(n4855), .dinb(n4782), .dout(n4856));
  jand g04635(.dina(n4856), .dinb(n743), .dout(n4857));
  jnot g04636(.din(n4710), .dout(n4858));
  jor  g04637(.dina(n4858), .dinb(n4857), .dout(n4859));
  jand g04638(.dina(n4859), .dinb(n4781), .dout(n4860));
  jand g04639(.dina(n4860), .dinb(n635), .dout(n4861));
  jor  g04640(.dina(n4717), .dinb(n4861), .dout(n4862));
  jand g04641(.dina(n4862), .dinb(n4780), .dout(n4863));
  jand g04642(.dina(n4863), .dinb(n515), .dout(n4864));
  jnot g04643(.din(n4725), .dout(n4865));
  jor  g04644(.dina(n4865), .dinb(n4864), .dout(n4866));
  jand g04645(.dina(n4866), .dinb(n4779), .dout(n4867));
  jand g04646(.dina(n4867), .dinb(n443), .dout(n4868));
  jor  g04647(.dina(n4732), .dinb(n4868), .dout(n4869));
  jand g04648(.dina(n4869), .dinb(n4778), .dout(n4870));
  jand g04649(.dina(n4870), .dinb(n352), .dout(n4871));
  jnot g04650(.din(n4740), .dout(n4872));
  jor  g04651(.dina(n4872), .dinb(n4871), .dout(n4873));
  jand g04652(.dina(n4873), .dinb(n4777), .dout(n4874));
  jand g04653(.dina(n4874), .dinb(n294), .dout(n4875));
  jor  g04654(.dina(n4747), .dinb(n4875), .dout(n4876));
  jand g04655(.dina(n4876), .dinb(n4776), .dout(n4877));
  jand g04656(.dina(n4877), .dinb(n239), .dout(n4878));
  jnot g04657(.din(n4755), .dout(n4879));
  jor  g04658(.dina(n4879), .dinb(n4878), .dout(n4880));
  jand g04659(.dina(n4880), .dinb(n4775), .dout(n4881));
  jand g04660(.dina(n4881), .dinb(n221), .dout(n4882));
  jor  g04661(.dina(n4762), .dinb(n4882), .dout(n4883));
  jand g04662(.dina(n4883), .dinb(n4774), .dout(n4884));
  jor  g04663(.dina(n4884), .dinb(n4773), .dout(n4885));
  jand g04664(.dina(asqrt[38] ), .dinb(n4576), .dout(n4886));
  jor  g04665(.dina(n4886), .dinb(n4442), .dout(n4887));
  jor  g04666(.dina(n4887), .dinb(n4885), .dout(n4888));
  jand g04667(.dina(n4888), .dinb(n218), .dout(n4889));
  jand g04668(.dina(n4582), .dinb(n4253), .dout(n4890));
  jor  g04669(.dina(n4890), .dinb(n4889), .dout(n4891));
  jor  g04670(.dina(n4891), .dinb(n4772), .dout(n4892));
  jor  g04671(.dina(n4892), .dinb(n4767), .dout(asqrt[37] ));
  jnot g04672(.din(n4772), .dout(n4894));
  jand g04673(.dina(n4765), .dinb(n4455), .dout(n4895));
  jnot g04674(.din(n4887), .dout(n4896));
  jand g04675(.dina(n4896), .dinb(n4895), .dout(n4897));
  jor  g04676(.dina(n4897), .dinb(asqrt[63] ), .dout(n4898));
  jnot g04677(.din(n4890), .dout(n4899));
  jand g04678(.dina(n4899), .dinb(n4898), .dout(n4900));
  jand g04679(.dina(n4900), .dinb(n4894), .dout(n4901));
  jand g04680(.dina(n4901), .dinb(n4766), .dout(n4902));
  jxor g04681(.dina(n4757), .dinb(n221), .dout(n4903));
  jor  g04682(.dina(n4903), .dinb(n4902), .dout(n4904));
  jxor g04683(.dina(n4904), .dinb(n4762), .dout(n4905));
  jnot g04684(.din(n4905), .dout(n4906));
  jor  g04685(.dina(n4902), .dinb(n4457), .dout(n4907));
  jnot g04686(.din(a[72] ), .dout(n4908));
  jnot g04687(.din(a[73] ), .dout(n4909));
  jand g04688(.dina(n4909), .dinb(n4908), .dout(n4910));
  jand g04689(.dina(n4910), .dinb(n4457), .dout(n4911));
  jnot g04690(.din(n4911), .dout(n4912));
  jand g04691(.dina(n4912), .dinb(n4907), .dout(n4913));
  jor  g04692(.dina(n4913), .dinb(n4582), .dout(n4914));
  jand g04693(.dina(n4913), .dinb(n4582), .dout(n4915));
  jor  g04694(.dina(n4902), .dinb(a[74] ), .dout(n4916));
  jand g04695(.dina(n4916), .dinb(a[75] ), .dout(n4917));
  jand g04696(.dina(asqrt[37] ), .dinb(n4459), .dout(n4918));
  jor  g04697(.dina(n4918), .dinb(n4917), .dout(n4919));
  jor  g04698(.dina(n4919), .dinb(n4915), .dout(n4920));
  jand g04699(.dina(n4920), .dinb(n4914), .dout(n4921));
  jor  g04700(.dina(n4921), .dinb(n4249), .dout(n4922));
  jand g04701(.dina(n4921), .dinb(n4249), .dout(n4923));
  jnot g04702(.din(n4459), .dout(n4924));
  jor  g04703(.dina(n4902), .dinb(n4924), .dout(n4925));
  jor  g04704(.dina(n4767), .dinb(n4582), .dout(n4926));
  jor  g04705(.dina(n4926), .dinb(n4771), .dout(n4927));
  jor  g04706(.dina(n4927), .dinb(n4889), .dout(n4928));
  jand g04707(.dina(n4928), .dinb(n4925), .dout(n4929));
  jxor g04708(.dina(n4929), .dinb(n4255), .dout(n4930));
  jor  g04709(.dina(n4930), .dinb(n4923), .dout(n4931));
  jand g04710(.dina(n4931), .dinb(n4922), .dout(n4932));
  jor  g04711(.dina(n4932), .dinb(n3955), .dout(n4933));
  jand g04712(.dina(n4932), .dinb(n3955), .dout(n4934));
  jxor g04713(.dina(n4461), .dinb(n4249), .dout(n4935));
  jor  g04714(.dina(n4935), .dinb(n4902), .dout(n4936));
  jxor g04715(.dina(n4936), .dinb(n4804), .dout(n4937));
  jnot g04716(.din(n4937), .dout(n4938));
  jor  g04717(.dina(n4938), .dinb(n4934), .dout(n4939));
  jand g04718(.dina(n4939), .dinb(n4933), .dout(n4940));
  jor  g04719(.dina(n4940), .dinb(n3642), .dout(n4941));
  jand g04720(.dina(n4940), .dinb(n3642), .dout(n4942));
  jxor g04721(.dina(n4586), .dinb(n3955), .dout(n4943));
  jor  g04722(.dina(n4943), .dinb(n4902), .dout(n4944));
  jxor g04723(.dina(n4944), .dinb(n4595), .dout(n4945));
  jnot g04724(.din(n4945), .dout(n4946));
  jor  g04725(.dina(n4946), .dinb(n4942), .dout(n4947));
  jand g04726(.dina(n4947), .dinb(n4941), .dout(n4948));
  jor  g04727(.dina(n4948), .dinb(n3368), .dout(n4949));
  jand g04728(.dina(n4948), .dinb(n3368), .dout(n4950));
  jxor g04729(.dina(n4598), .dinb(n3642), .dout(n4951));
  jor  g04730(.dina(n4951), .dinb(n4902), .dout(n4952));
  jxor g04731(.dina(n4952), .dinb(n4604), .dout(n4953));
  jor  g04732(.dina(n4953), .dinb(n4950), .dout(n4954));
  jand g04733(.dina(n4954), .dinb(n4949), .dout(n4955));
  jor  g04734(.dina(n4955), .dinb(n3089), .dout(n4956));
  jand g04735(.dina(n4955), .dinb(n3089), .dout(n4957));
  jxor g04736(.dina(n4606), .dinb(n3368), .dout(n4958));
  jor  g04737(.dina(n4958), .dinb(n4902), .dout(n4959));
  jxor g04738(.dina(n4959), .dinb(n4612), .dout(n4960));
  jor  g04739(.dina(n4960), .dinb(n4957), .dout(n4961));
  jand g04740(.dina(n4961), .dinb(n4956), .dout(n4962));
  jor  g04741(.dina(n4962), .dinb(n2833), .dout(n4963));
  jand g04742(.dina(n4962), .dinb(n2833), .dout(n4964));
  jxor g04743(.dina(n4614), .dinb(n3089), .dout(n4965));
  jor  g04744(.dina(n4965), .dinb(n4902), .dout(n4966));
  jxor g04745(.dina(n4966), .dinb(n4620), .dout(n4967));
  jor  g04746(.dina(n4967), .dinb(n4964), .dout(n4968));
  jand g04747(.dina(n4968), .dinb(n4963), .dout(n4969));
  jor  g04748(.dina(n4969), .dinb(n2572), .dout(n4970));
  jand g04749(.dina(n4969), .dinb(n2572), .dout(n4971));
  jxor g04750(.dina(n4622), .dinb(n2833), .dout(n4972));
  jor  g04751(.dina(n4972), .dinb(n4902), .dout(n4973));
  jxor g04752(.dina(n4973), .dinb(n4628), .dout(n4974));
  jor  g04753(.dina(n4974), .dinb(n4971), .dout(n4975));
  jand g04754(.dina(n4975), .dinb(n4970), .dout(n4976));
  jor  g04755(.dina(n4976), .dinb(n2345), .dout(n4977));
  jand g04756(.dina(n4976), .dinb(n2345), .dout(n4978));
  jxor g04757(.dina(n4630), .dinb(n2572), .dout(n4979));
  jor  g04758(.dina(n4979), .dinb(n4902), .dout(n4980));
  jxor g04759(.dina(n4980), .dinb(n4823), .dout(n4981));
  jnot g04760(.din(n4981), .dout(n4982));
  jor  g04761(.dina(n4982), .dinb(n4978), .dout(n4983));
  jand g04762(.dina(n4983), .dinb(n4977), .dout(n4984));
  jor  g04763(.dina(n4984), .dinb(n2108), .dout(n4985));
  jand g04764(.dina(n4984), .dinb(n2108), .dout(n4986));
  jxor g04765(.dina(n4637), .dinb(n2345), .dout(n4987));
  jor  g04766(.dina(n4987), .dinb(n4902), .dout(n4988));
  jxor g04767(.dina(n4988), .dinb(n4643), .dout(n4989));
  jor  g04768(.dina(n4989), .dinb(n4986), .dout(n4990));
  jand g04769(.dina(n4990), .dinb(n4985), .dout(n4991));
  jor  g04770(.dina(n4991), .dinb(n1912), .dout(n4992));
  jand g04771(.dina(n4991), .dinb(n1912), .dout(n4993));
  jxor g04772(.dina(n4645), .dinb(n2108), .dout(n4994));
  jor  g04773(.dina(n4994), .dinb(n4902), .dout(n4995));
  jxor g04774(.dina(n4995), .dinb(n4830), .dout(n4996));
  jnot g04775(.din(n4996), .dout(n4997));
  jor  g04776(.dina(n4997), .dinb(n4993), .dout(n4998));
  jand g04777(.dina(n4998), .dinb(n4992), .dout(n4999));
  jor  g04778(.dina(n4999), .dinb(n1699), .dout(n5000));
  jand g04779(.dina(n4999), .dinb(n1699), .dout(n5001));
  jxor g04780(.dina(n4652), .dinb(n1912), .dout(n5002));
  jor  g04781(.dina(n5002), .dinb(n4902), .dout(n5003));
  jxor g04782(.dina(n5003), .dinb(n4658), .dout(n5004));
  jor  g04783(.dina(n5004), .dinb(n5001), .dout(n5005));
  jand g04784(.dina(n5005), .dinb(n5000), .dout(n5006));
  jor  g04785(.dina(n5006), .dinb(n1516), .dout(n5007));
  jand g04786(.dina(n5006), .dinb(n1516), .dout(n5008));
  jxor g04787(.dina(n4660), .dinb(n1699), .dout(n5009));
  jor  g04788(.dina(n5009), .dinb(n4902), .dout(n5010));
  jxor g04789(.dina(n5010), .dinb(n4837), .dout(n5011));
  jnot g04790(.din(n5011), .dout(n5012));
  jor  g04791(.dina(n5012), .dinb(n5008), .dout(n5013));
  jand g04792(.dina(n5013), .dinb(n5007), .dout(n5014));
  jor  g04793(.dina(n5014), .dinb(n1332), .dout(n5015));
  jand g04794(.dina(n5014), .dinb(n1332), .dout(n5016));
  jxor g04795(.dina(n4667), .dinb(n1516), .dout(n5017));
  jor  g04796(.dina(n5017), .dinb(n4902), .dout(n5018));
  jxor g04797(.dina(n5018), .dinb(n4841), .dout(n5019));
  jnot g04798(.din(n5019), .dout(n5020));
  jor  g04799(.dina(n5020), .dinb(n5016), .dout(n5021));
  jand g04800(.dina(n5021), .dinb(n5015), .dout(n5022));
  jor  g04801(.dina(n5022), .dinb(n1173), .dout(n5023));
  jand g04802(.dina(n5022), .dinb(n1173), .dout(n5024));
  jxor g04803(.dina(n4674), .dinb(n1332), .dout(n5025));
  jor  g04804(.dina(n5025), .dinb(n4902), .dout(n5026));
  jxor g04805(.dina(n5026), .dinb(n4680), .dout(n5027));
  jor  g04806(.dina(n5027), .dinb(n5024), .dout(n5028));
  jand g04807(.dina(n5028), .dinb(n5023), .dout(n5029));
  jor  g04808(.dina(n5029), .dinb(n1008), .dout(n5030));
  jand g04809(.dina(n5029), .dinb(n1008), .dout(n5031));
  jxor g04810(.dina(n4682), .dinb(n1173), .dout(n5032));
  jor  g04811(.dina(n5032), .dinb(n4902), .dout(n5033));
  jxor g04812(.dina(n5033), .dinb(n4688), .dout(n5034));
  jor  g04813(.dina(n5034), .dinb(n5031), .dout(n5035));
  jand g04814(.dina(n5035), .dinb(n5030), .dout(n5036));
  jor  g04815(.dina(n5036), .dinb(n884), .dout(n5037));
  jand g04816(.dina(n5036), .dinb(n884), .dout(n5038));
  jxor g04817(.dina(n4690), .dinb(n1008), .dout(n5039));
  jor  g04818(.dina(n5039), .dinb(n4902), .dout(n5040));
  jxor g04819(.dina(n5040), .dinb(n4851), .dout(n5041));
  jnot g04820(.din(n5041), .dout(n5042));
  jor  g04821(.dina(n5042), .dinb(n5038), .dout(n5043));
  jand g04822(.dina(n5043), .dinb(n5037), .dout(n5044));
  jor  g04823(.dina(n5044), .dinb(n743), .dout(n5045));
  jand g04824(.dina(n5044), .dinb(n743), .dout(n5046));
  jxor g04825(.dina(n4697), .dinb(n884), .dout(n5047));
  jor  g04826(.dina(n5047), .dinb(n4902), .dout(n5048));
  jxor g04827(.dina(n5048), .dinb(n4703), .dout(n5049));
  jor  g04828(.dina(n5049), .dinb(n5046), .dout(n5050));
  jand g04829(.dina(n5050), .dinb(n5045), .dout(n5051));
  jor  g04830(.dina(n5051), .dinb(n635), .dout(n5052));
  jand g04831(.dina(n5051), .dinb(n635), .dout(n5053));
  jxor g04832(.dina(n4705), .dinb(n743), .dout(n5054));
  jor  g04833(.dina(n5054), .dinb(n4902), .dout(n5055));
  jxor g04834(.dina(n5055), .dinb(n4858), .dout(n5056));
  jnot g04835(.din(n5056), .dout(n5057));
  jor  g04836(.dina(n5057), .dinb(n5053), .dout(n5058));
  jand g04837(.dina(n5058), .dinb(n5052), .dout(n5059));
  jor  g04838(.dina(n5059), .dinb(n515), .dout(n5060));
  jand g04839(.dina(n5059), .dinb(n515), .dout(n5061));
  jxor g04840(.dina(n4712), .dinb(n635), .dout(n5062));
  jor  g04841(.dina(n5062), .dinb(n4902), .dout(n5063));
  jxor g04842(.dina(n5063), .dinb(n4718), .dout(n5064));
  jor  g04843(.dina(n5064), .dinb(n5061), .dout(n5065));
  jand g04844(.dina(n5065), .dinb(n5060), .dout(n5066));
  jor  g04845(.dina(n5066), .dinb(n443), .dout(n5067));
  jand g04846(.dina(n5066), .dinb(n443), .dout(n5068));
  jxor g04847(.dina(n4720), .dinb(n515), .dout(n5069));
  jor  g04848(.dina(n5069), .dinb(n4902), .dout(n5070));
  jxor g04849(.dina(n5070), .dinb(n4865), .dout(n5071));
  jnot g04850(.din(n5071), .dout(n5072));
  jor  g04851(.dina(n5072), .dinb(n5068), .dout(n5073));
  jand g04852(.dina(n5073), .dinb(n5067), .dout(n5074));
  jor  g04853(.dina(n5074), .dinb(n352), .dout(n5075));
  jand g04854(.dina(n5074), .dinb(n352), .dout(n5076));
  jxor g04855(.dina(n4727), .dinb(n443), .dout(n5077));
  jor  g04856(.dina(n5077), .dinb(n4902), .dout(n5078));
  jxor g04857(.dina(n5078), .dinb(n4733), .dout(n5079));
  jor  g04858(.dina(n5079), .dinb(n5076), .dout(n5080));
  jand g04859(.dina(n5080), .dinb(n5075), .dout(n5081));
  jor  g04860(.dina(n5081), .dinb(n294), .dout(n5082));
  jand g04861(.dina(n5081), .dinb(n294), .dout(n5083));
  jxor g04862(.dina(n4735), .dinb(n352), .dout(n5084));
  jor  g04863(.dina(n5084), .dinb(n4902), .dout(n5085));
  jxor g04864(.dina(n5085), .dinb(n4872), .dout(n5086));
  jnot g04865(.din(n5086), .dout(n5087));
  jor  g04866(.dina(n5087), .dinb(n5083), .dout(n5088));
  jand g04867(.dina(n5088), .dinb(n5082), .dout(n5089));
  jor  g04868(.dina(n5089), .dinb(n239), .dout(n5090));
  jand g04869(.dina(n5089), .dinb(n239), .dout(n5091));
  jxor g04870(.dina(n4742), .dinb(n294), .dout(n5092));
  jor  g04871(.dina(n5092), .dinb(n4902), .dout(n5093));
  jxor g04872(.dina(n5093), .dinb(n4748), .dout(n5094));
  jor  g04873(.dina(n5094), .dinb(n5091), .dout(n5095));
  jand g04874(.dina(n5095), .dinb(n5090), .dout(n5096));
  jor  g04875(.dina(n5096), .dinb(n221), .dout(n5097));
  jand g04876(.dina(n5096), .dinb(n221), .dout(n5098));
  jxor g04877(.dina(n4750), .dinb(n239), .dout(n5099));
  jor  g04878(.dina(n5099), .dinb(n4902), .dout(n5100));
  jxor g04879(.dina(n5100), .dinb(n4879), .dout(n5101));
  jnot g04880(.din(n5101), .dout(n5102));
  jor  g04881(.dina(n5102), .dinb(n5098), .dout(n5103));
  jand g04882(.dina(n5103), .dinb(n5097), .dout(n5104));
  jand g04883(.dina(n5104), .dinb(n4906), .dout(n5105));
  jand g04884(.dina(n4892), .dinb(n4895), .dout(n5107));
  jor  g04885(.dina(n5104), .dinb(n4906), .dout(n5108));
  jor  g04886(.dina(n5108), .dinb(n4767), .dout(n5109));
  jor  g04887(.dina(n5109), .dinb(n5107), .dout(n5110));
  jand g04888(.dina(n5110), .dinb(n218), .dout(n5111));
  jand g04889(.dina(n4901), .dinb(n4884), .dout(n5112));
  jand g04890(.dina(n4885), .dinb(asqrt[63] ), .dout(n5113));
  jand g04891(.dina(n5113), .dinb(n4766), .dout(n5114));
  jnot g04892(.din(n5114), .dout(n5115));
  jor  g04893(.dina(n5115), .dinb(n5112), .dout(n5116));
  jnot g04894(.din(n5116), .dout(n5117));
  jor  g04895(.dina(n5117), .dinb(n5111), .dout(n5118));
  jor  g04896(.dina(n5118), .dinb(n5105), .dout(asqrt[36] ));
  jnot g04897(.din(a[70] ), .dout(n5121));
  jnot g04898(.din(a[71] ), .dout(n5122));
  jand g04899(.dina(n5122), .dinb(n5121), .dout(n5123));
  jand g04900(.dina(n5123), .dinb(n4908), .dout(n5124));
  jand g04901(.dina(asqrt[36] ), .dinb(a[72] ), .dout(n5125));
  jor  g04902(.dina(n5125), .dinb(n5124), .dout(n5126));
  jand g04903(.dina(n5126), .dinb(asqrt[37] ), .dout(n5127));
  jor  g04904(.dina(n5126), .dinb(asqrt[37] ), .dout(n5128));
  jand g04905(.dina(asqrt[36] ), .dinb(n4908), .dout(n5129));
  jor  g04906(.dina(n5129), .dinb(n4909), .dout(n5130));
  jnot g04907(.din(n4910), .dout(n5131));
  jnot g04908(.din(n5105), .dout(n5132));
  jnot g04909(.din(n5107), .dout(n5134));
  jnot g04910(.din(n5097), .dout(n5135));
  jnot g04911(.din(n5090), .dout(n5136));
  jnot g04912(.din(n5082), .dout(n5137));
  jnot g04913(.din(n5075), .dout(n5138));
  jnot g04914(.din(n5067), .dout(n5139));
  jnot g04915(.din(n5060), .dout(n5140));
  jnot g04916(.din(n5052), .dout(n5141));
  jnot g04917(.din(n5045), .dout(n5142));
  jnot g04918(.din(n5037), .dout(n5143));
  jnot g04919(.din(n5030), .dout(n5144));
  jnot g04920(.din(n5023), .dout(n5145));
  jnot g04921(.din(n5015), .dout(n5146));
  jnot g04922(.din(n5007), .dout(n5147));
  jnot g04923(.din(n5000), .dout(n5148));
  jnot g04924(.din(n4992), .dout(n5149));
  jnot g04925(.din(n4985), .dout(n5150));
  jnot g04926(.din(n4977), .dout(n5151));
  jnot g04927(.din(n4970), .dout(n5152));
  jnot g04928(.din(n4963), .dout(n5153));
  jnot g04929(.din(n4956), .dout(n5154));
  jnot g04930(.din(n4949), .dout(n5155));
  jnot g04931(.din(n4941), .dout(n5156));
  jnot g04932(.din(n4933), .dout(n5157));
  jnot g04933(.din(n4922), .dout(n5158));
  jnot g04934(.din(n4914), .dout(n5159));
  jand g04935(.dina(asqrt[37] ), .dinb(a[74] ), .dout(n5160));
  jor  g04936(.dina(n4911), .dinb(n5160), .dout(n5161));
  jor  g04937(.dina(n5161), .dinb(asqrt[38] ), .dout(n5162));
  jand g04938(.dina(asqrt[37] ), .dinb(n4457), .dout(n5163));
  jor  g04939(.dina(n5163), .dinb(n4458), .dout(n5164));
  jand g04940(.dina(n4925), .dinb(n5164), .dout(n5165));
  jand g04941(.dina(n5165), .dinb(n5162), .dout(n5166));
  jor  g04942(.dina(n5166), .dinb(n5159), .dout(n5167));
  jor  g04943(.dina(n5167), .dinb(asqrt[39] ), .dout(n5168));
  jnot g04944(.din(n4930), .dout(n5169));
  jand g04945(.dina(n5169), .dinb(n5168), .dout(n5170));
  jor  g04946(.dina(n5170), .dinb(n5158), .dout(n5171));
  jor  g04947(.dina(n5171), .dinb(asqrt[40] ), .dout(n5172));
  jand g04948(.dina(n4937), .dinb(n5172), .dout(n5173));
  jor  g04949(.dina(n5173), .dinb(n5157), .dout(n5174));
  jor  g04950(.dina(n5174), .dinb(asqrt[41] ), .dout(n5175));
  jand g04951(.dina(n4945), .dinb(n5175), .dout(n5176));
  jor  g04952(.dina(n5176), .dinb(n5156), .dout(n5177));
  jor  g04953(.dina(n5177), .dinb(asqrt[42] ), .dout(n5178));
  jnot g04954(.din(n4953), .dout(n5179));
  jand g04955(.dina(n5179), .dinb(n5178), .dout(n5180));
  jor  g04956(.dina(n5180), .dinb(n5155), .dout(n5181));
  jor  g04957(.dina(n5181), .dinb(asqrt[43] ), .dout(n5182));
  jnot g04958(.din(n4960), .dout(n5183));
  jand g04959(.dina(n5183), .dinb(n5182), .dout(n5184));
  jor  g04960(.dina(n5184), .dinb(n5154), .dout(n5185));
  jor  g04961(.dina(n5185), .dinb(asqrt[44] ), .dout(n5186));
  jnot g04962(.din(n4967), .dout(n5187));
  jand g04963(.dina(n5187), .dinb(n5186), .dout(n5188));
  jor  g04964(.dina(n5188), .dinb(n5153), .dout(n5189));
  jor  g04965(.dina(n5189), .dinb(asqrt[45] ), .dout(n5190));
  jnot g04966(.din(n4974), .dout(n5191));
  jand g04967(.dina(n5191), .dinb(n5190), .dout(n5192));
  jor  g04968(.dina(n5192), .dinb(n5152), .dout(n5193));
  jor  g04969(.dina(n5193), .dinb(asqrt[46] ), .dout(n5194));
  jand g04970(.dina(n4981), .dinb(n5194), .dout(n5195));
  jor  g04971(.dina(n5195), .dinb(n5151), .dout(n5196));
  jor  g04972(.dina(n5196), .dinb(asqrt[47] ), .dout(n5197));
  jnot g04973(.din(n4989), .dout(n5198));
  jand g04974(.dina(n5198), .dinb(n5197), .dout(n5199));
  jor  g04975(.dina(n5199), .dinb(n5150), .dout(n5200));
  jor  g04976(.dina(n5200), .dinb(asqrt[48] ), .dout(n5201));
  jand g04977(.dina(n4996), .dinb(n5201), .dout(n5202));
  jor  g04978(.dina(n5202), .dinb(n5149), .dout(n5203));
  jor  g04979(.dina(n5203), .dinb(asqrt[49] ), .dout(n5204));
  jnot g04980(.din(n5004), .dout(n5205));
  jand g04981(.dina(n5205), .dinb(n5204), .dout(n5206));
  jor  g04982(.dina(n5206), .dinb(n5148), .dout(n5207));
  jor  g04983(.dina(n5207), .dinb(asqrt[50] ), .dout(n5208));
  jand g04984(.dina(n5011), .dinb(n5208), .dout(n5209));
  jor  g04985(.dina(n5209), .dinb(n5147), .dout(n5210));
  jor  g04986(.dina(n5210), .dinb(asqrt[51] ), .dout(n5211));
  jand g04987(.dina(n5019), .dinb(n5211), .dout(n5212));
  jor  g04988(.dina(n5212), .dinb(n5146), .dout(n5213));
  jor  g04989(.dina(n5213), .dinb(asqrt[52] ), .dout(n5214));
  jnot g04990(.din(n5027), .dout(n5215));
  jand g04991(.dina(n5215), .dinb(n5214), .dout(n5216));
  jor  g04992(.dina(n5216), .dinb(n5145), .dout(n5217));
  jor  g04993(.dina(n5217), .dinb(asqrt[53] ), .dout(n5218));
  jnot g04994(.din(n5034), .dout(n5219));
  jand g04995(.dina(n5219), .dinb(n5218), .dout(n5220));
  jor  g04996(.dina(n5220), .dinb(n5144), .dout(n5221));
  jor  g04997(.dina(n5221), .dinb(asqrt[54] ), .dout(n5222));
  jand g04998(.dina(n5041), .dinb(n5222), .dout(n5223));
  jor  g04999(.dina(n5223), .dinb(n5143), .dout(n5224));
  jor  g05000(.dina(n5224), .dinb(asqrt[55] ), .dout(n5225));
  jnot g05001(.din(n5049), .dout(n5226));
  jand g05002(.dina(n5226), .dinb(n5225), .dout(n5227));
  jor  g05003(.dina(n5227), .dinb(n5142), .dout(n5228));
  jor  g05004(.dina(n5228), .dinb(asqrt[56] ), .dout(n5229));
  jand g05005(.dina(n5056), .dinb(n5229), .dout(n5230));
  jor  g05006(.dina(n5230), .dinb(n5141), .dout(n5231));
  jor  g05007(.dina(n5231), .dinb(asqrt[57] ), .dout(n5232));
  jnot g05008(.din(n5064), .dout(n5233));
  jand g05009(.dina(n5233), .dinb(n5232), .dout(n5234));
  jor  g05010(.dina(n5234), .dinb(n5140), .dout(n5235));
  jor  g05011(.dina(n5235), .dinb(asqrt[58] ), .dout(n5236));
  jand g05012(.dina(n5071), .dinb(n5236), .dout(n5237));
  jor  g05013(.dina(n5237), .dinb(n5139), .dout(n5238));
  jor  g05014(.dina(n5238), .dinb(asqrt[59] ), .dout(n5239));
  jnot g05015(.din(n5079), .dout(n5240));
  jand g05016(.dina(n5240), .dinb(n5239), .dout(n5241));
  jor  g05017(.dina(n5241), .dinb(n5138), .dout(n5242));
  jor  g05018(.dina(n5242), .dinb(asqrt[60] ), .dout(n5243));
  jand g05019(.dina(n5086), .dinb(n5243), .dout(n5244));
  jor  g05020(.dina(n5244), .dinb(n5137), .dout(n5245));
  jor  g05021(.dina(n5245), .dinb(asqrt[61] ), .dout(n5246));
  jnot g05022(.din(n5094), .dout(n5247));
  jand g05023(.dina(n5247), .dinb(n5246), .dout(n5248));
  jor  g05024(.dina(n5248), .dinb(n5136), .dout(n5249));
  jor  g05025(.dina(n5249), .dinb(asqrt[62] ), .dout(n5250));
  jand g05026(.dina(n5101), .dinb(n5250), .dout(n5251));
  jor  g05027(.dina(n5251), .dinb(n5135), .dout(n5252));
  jand g05028(.dina(n5252), .dinb(n4905), .dout(n5253));
  jand g05029(.dina(n5253), .dinb(n4766), .dout(n5254));
  jand g05030(.dina(n5254), .dinb(n5134), .dout(n5255));
  jor  g05031(.dina(n5255), .dinb(asqrt[63] ), .dout(n5256));
  jand g05032(.dina(n5116), .dinb(n5256), .dout(n5257));
  jand g05033(.dina(n5257), .dinb(n5132), .dout(n5259));
  jor  g05034(.dina(n5259), .dinb(n5131), .dout(n5260));
  jand g05035(.dina(n5260), .dinb(n5130), .dout(n5261));
  jand g05036(.dina(n5261), .dinb(n5128), .dout(n5262));
  jor  g05037(.dina(n5262), .dinb(n5127), .dout(n5263));
  jand g05038(.dina(n5263), .dinb(asqrt[38] ), .dout(n5264));
  jor  g05039(.dina(n5263), .dinb(asqrt[38] ), .dout(n5265));
  jand g05040(.dina(asqrt[36] ), .dinb(n4910), .dout(n5266));
  jand g05041(.dina(n5115), .dinb(n5132), .dout(n5267));
  jand g05042(.dina(n5267), .dinb(n5256), .dout(n5268));
  jand g05043(.dina(n5268), .dinb(asqrt[37] ), .dout(n5269));
  jor  g05044(.dina(n5269), .dinb(n5266), .dout(n5270));
  jxor g05045(.dina(n5270), .dinb(a[74] ), .dout(n5271));
  jnot g05046(.din(n5271), .dout(n5272));
  jand g05047(.dina(n5272), .dinb(n5265), .dout(n5273));
  jor  g05048(.dina(n5273), .dinb(n5264), .dout(n5274));
  jand g05049(.dina(n5274), .dinb(asqrt[39] ), .dout(n5275));
  jor  g05050(.dina(n5274), .dinb(asqrt[39] ), .dout(n5276));
  jxor g05051(.dina(n4913), .dinb(n4582), .dout(n5277));
  jand g05052(.dina(n5277), .dinb(asqrt[36] ), .dout(n5278));
  jxor g05053(.dina(n5278), .dinb(n5165), .dout(n5279));
  jand g05054(.dina(n5279), .dinb(n5276), .dout(n5280));
  jor  g05055(.dina(n5280), .dinb(n5275), .dout(n5281));
  jand g05056(.dina(n5281), .dinb(asqrt[40] ), .dout(n5282));
  jor  g05057(.dina(n5281), .dinb(asqrt[40] ), .dout(n5283));
  jxor g05058(.dina(n4921), .dinb(n4249), .dout(n5284));
  jand g05059(.dina(n5284), .dinb(asqrt[36] ), .dout(n5285));
  jxor g05060(.dina(n5285), .dinb(n4930), .dout(n5286));
  jnot g05061(.din(n5286), .dout(n5287));
  jand g05062(.dina(n5287), .dinb(n5283), .dout(n5288));
  jor  g05063(.dina(n5288), .dinb(n5282), .dout(n5289));
  jand g05064(.dina(n5289), .dinb(asqrt[41] ), .dout(n5290));
  jor  g05065(.dina(n5289), .dinb(asqrt[41] ), .dout(n5291));
  jxor g05066(.dina(n4932), .dinb(n3955), .dout(n5292));
  jand g05067(.dina(n5292), .dinb(asqrt[36] ), .dout(n5293));
  jxor g05068(.dina(n5293), .dinb(n4937), .dout(n5294));
  jand g05069(.dina(n5294), .dinb(n5291), .dout(n5295));
  jor  g05070(.dina(n5295), .dinb(n5290), .dout(n5296));
  jand g05071(.dina(n5296), .dinb(asqrt[42] ), .dout(n5297));
  jor  g05072(.dina(n5296), .dinb(asqrt[42] ), .dout(n5298));
  jxor g05073(.dina(n4940), .dinb(n3642), .dout(n5299));
  jand g05074(.dina(n5299), .dinb(asqrt[36] ), .dout(n5300));
  jxor g05075(.dina(n5300), .dinb(n4945), .dout(n5301));
  jand g05076(.dina(n5301), .dinb(n5298), .dout(n5302));
  jor  g05077(.dina(n5302), .dinb(n5297), .dout(n5303));
  jand g05078(.dina(n5303), .dinb(asqrt[43] ), .dout(n5304));
  jor  g05079(.dina(n5303), .dinb(asqrt[43] ), .dout(n5305));
  jxor g05080(.dina(n4948), .dinb(n3368), .dout(n5306));
  jand g05081(.dina(n5306), .dinb(asqrt[36] ), .dout(n5307));
  jxor g05082(.dina(n5307), .dinb(n5179), .dout(n5308));
  jand g05083(.dina(n5308), .dinb(n5305), .dout(n5309));
  jor  g05084(.dina(n5309), .dinb(n5304), .dout(n5310));
  jand g05085(.dina(n5310), .dinb(asqrt[44] ), .dout(n5311));
  jor  g05086(.dina(n5310), .dinb(asqrt[44] ), .dout(n5312));
  jxor g05087(.dina(n4955), .dinb(n3089), .dout(n5313));
  jand g05088(.dina(n5313), .dinb(asqrt[36] ), .dout(n5314));
  jxor g05089(.dina(n5314), .dinb(n4960), .dout(n5315));
  jnot g05090(.din(n5315), .dout(n5316));
  jand g05091(.dina(n5316), .dinb(n5312), .dout(n5317));
  jor  g05092(.dina(n5317), .dinb(n5311), .dout(n5318));
  jand g05093(.dina(n5318), .dinb(asqrt[45] ), .dout(n5319));
  jor  g05094(.dina(n5318), .dinb(asqrt[45] ), .dout(n5320));
  jxor g05095(.dina(n4962), .dinb(n2833), .dout(n5321));
  jand g05096(.dina(n5321), .dinb(asqrt[36] ), .dout(n5322));
  jxor g05097(.dina(n5322), .dinb(n4967), .dout(n5323));
  jnot g05098(.din(n5323), .dout(n5324));
  jand g05099(.dina(n5324), .dinb(n5320), .dout(n5325));
  jor  g05100(.dina(n5325), .dinb(n5319), .dout(n5326));
  jand g05101(.dina(n5326), .dinb(asqrt[46] ), .dout(n5327));
  jor  g05102(.dina(n5326), .dinb(asqrt[46] ), .dout(n5328));
  jxor g05103(.dina(n4969), .dinb(n2572), .dout(n5329));
  jand g05104(.dina(n5329), .dinb(asqrt[36] ), .dout(n5330));
  jxor g05105(.dina(n5330), .dinb(n4974), .dout(n5331));
  jnot g05106(.din(n5331), .dout(n5332));
  jand g05107(.dina(n5332), .dinb(n5328), .dout(n5333));
  jor  g05108(.dina(n5333), .dinb(n5327), .dout(n5334));
  jand g05109(.dina(n5334), .dinb(asqrt[47] ), .dout(n5335));
  jor  g05110(.dina(n5334), .dinb(asqrt[47] ), .dout(n5336));
  jxor g05111(.dina(n4976), .dinb(n2345), .dout(n5337));
  jand g05112(.dina(n5337), .dinb(asqrt[36] ), .dout(n5338));
  jxor g05113(.dina(n5338), .dinb(n4981), .dout(n5339));
  jand g05114(.dina(n5339), .dinb(n5336), .dout(n5340));
  jor  g05115(.dina(n5340), .dinb(n5335), .dout(n5341));
  jand g05116(.dina(n5341), .dinb(asqrt[48] ), .dout(n5342));
  jor  g05117(.dina(n5341), .dinb(asqrt[48] ), .dout(n5343));
  jxor g05118(.dina(n4984), .dinb(n2108), .dout(n5344));
  jand g05119(.dina(n5344), .dinb(asqrt[36] ), .dout(n5345));
  jxor g05120(.dina(n5345), .dinb(n4989), .dout(n5346));
  jnot g05121(.din(n5346), .dout(n5347));
  jand g05122(.dina(n5347), .dinb(n5343), .dout(n5348));
  jor  g05123(.dina(n5348), .dinb(n5342), .dout(n5349));
  jand g05124(.dina(n5349), .dinb(asqrt[49] ), .dout(n5350));
  jor  g05125(.dina(n5349), .dinb(asqrt[49] ), .dout(n5351));
  jxor g05126(.dina(n4991), .dinb(n1912), .dout(n5352));
  jand g05127(.dina(n5352), .dinb(asqrt[36] ), .dout(n5353));
  jxor g05128(.dina(n5353), .dinb(n4996), .dout(n5354));
  jand g05129(.dina(n5354), .dinb(n5351), .dout(n5355));
  jor  g05130(.dina(n5355), .dinb(n5350), .dout(n5356));
  jand g05131(.dina(n5356), .dinb(asqrt[50] ), .dout(n5357));
  jor  g05132(.dina(n5356), .dinb(asqrt[50] ), .dout(n5358));
  jxor g05133(.dina(n4999), .dinb(n1699), .dout(n5359));
  jand g05134(.dina(n5359), .dinb(asqrt[36] ), .dout(n5360));
  jxor g05135(.dina(n5360), .dinb(n5004), .dout(n5361));
  jnot g05136(.din(n5361), .dout(n5362));
  jand g05137(.dina(n5362), .dinb(n5358), .dout(n5363));
  jor  g05138(.dina(n5363), .dinb(n5357), .dout(n5364));
  jand g05139(.dina(n5364), .dinb(asqrt[51] ), .dout(n5365));
  jor  g05140(.dina(n5364), .dinb(asqrt[51] ), .dout(n5366));
  jxor g05141(.dina(n5006), .dinb(n1516), .dout(n5367));
  jand g05142(.dina(n5367), .dinb(asqrt[36] ), .dout(n5368));
  jxor g05143(.dina(n5368), .dinb(n5011), .dout(n5369));
  jand g05144(.dina(n5369), .dinb(n5366), .dout(n5370));
  jor  g05145(.dina(n5370), .dinb(n5365), .dout(n5371));
  jand g05146(.dina(n5371), .dinb(asqrt[52] ), .dout(n5372));
  jor  g05147(.dina(n5371), .dinb(asqrt[52] ), .dout(n5373));
  jxor g05148(.dina(n5014), .dinb(n1332), .dout(n5374));
  jand g05149(.dina(n5374), .dinb(asqrt[36] ), .dout(n5375));
  jxor g05150(.dina(n5375), .dinb(n5019), .dout(n5376));
  jand g05151(.dina(n5376), .dinb(n5373), .dout(n5377));
  jor  g05152(.dina(n5377), .dinb(n5372), .dout(n5378));
  jand g05153(.dina(n5378), .dinb(asqrt[53] ), .dout(n5379));
  jor  g05154(.dina(n5378), .dinb(asqrt[53] ), .dout(n5380));
  jxor g05155(.dina(n5022), .dinb(n1173), .dout(n5381));
  jand g05156(.dina(n5381), .dinb(asqrt[36] ), .dout(n5382));
  jxor g05157(.dina(n5382), .dinb(n5027), .dout(n5383));
  jnot g05158(.din(n5383), .dout(n5384));
  jand g05159(.dina(n5384), .dinb(n5380), .dout(n5385));
  jor  g05160(.dina(n5385), .dinb(n5379), .dout(n5386));
  jand g05161(.dina(n5386), .dinb(asqrt[54] ), .dout(n5387));
  jor  g05162(.dina(n5386), .dinb(asqrt[54] ), .dout(n5388));
  jxor g05163(.dina(n5029), .dinb(n1008), .dout(n5389));
  jand g05164(.dina(n5389), .dinb(asqrt[36] ), .dout(n5390));
  jxor g05165(.dina(n5390), .dinb(n5034), .dout(n5391));
  jnot g05166(.din(n5391), .dout(n5392));
  jand g05167(.dina(n5392), .dinb(n5388), .dout(n5393));
  jor  g05168(.dina(n5393), .dinb(n5387), .dout(n5394));
  jand g05169(.dina(n5394), .dinb(asqrt[55] ), .dout(n5395));
  jor  g05170(.dina(n5394), .dinb(asqrt[55] ), .dout(n5396));
  jxor g05171(.dina(n5036), .dinb(n884), .dout(n5397));
  jand g05172(.dina(n5397), .dinb(asqrt[36] ), .dout(n5398));
  jxor g05173(.dina(n5398), .dinb(n5041), .dout(n5399));
  jand g05174(.dina(n5399), .dinb(n5396), .dout(n5400));
  jor  g05175(.dina(n5400), .dinb(n5395), .dout(n5401));
  jand g05176(.dina(n5401), .dinb(asqrt[56] ), .dout(n5402));
  jor  g05177(.dina(n5401), .dinb(asqrt[56] ), .dout(n5403));
  jxor g05178(.dina(n5044), .dinb(n743), .dout(n5404));
  jand g05179(.dina(n5404), .dinb(asqrt[36] ), .dout(n5405));
  jxor g05180(.dina(n5405), .dinb(n5049), .dout(n5406));
  jnot g05181(.din(n5406), .dout(n5407));
  jand g05182(.dina(n5407), .dinb(n5403), .dout(n5408));
  jor  g05183(.dina(n5408), .dinb(n5402), .dout(n5409));
  jand g05184(.dina(n5409), .dinb(asqrt[57] ), .dout(n5410));
  jor  g05185(.dina(n5409), .dinb(asqrt[57] ), .dout(n5411));
  jxor g05186(.dina(n5051), .dinb(n635), .dout(n5412));
  jand g05187(.dina(n5412), .dinb(asqrt[36] ), .dout(n5413));
  jxor g05188(.dina(n5413), .dinb(n5056), .dout(n5414));
  jand g05189(.dina(n5414), .dinb(n5411), .dout(n5415));
  jor  g05190(.dina(n5415), .dinb(n5410), .dout(n5416));
  jand g05191(.dina(n5416), .dinb(asqrt[58] ), .dout(n5417));
  jor  g05192(.dina(n5416), .dinb(asqrt[58] ), .dout(n5418));
  jxor g05193(.dina(n5059), .dinb(n515), .dout(n5419));
  jand g05194(.dina(n5419), .dinb(asqrt[36] ), .dout(n5420));
  jxor g05195(.dina(n5420), .dinb(n5064), .dout(n5421));
  jnot g05196(.din(n5421), .dout(n5422));
  jand g05197(.dina(n5422), .dinb(n5418), .dout(n5423));
  jor  g05198(.dina(n5423), .dinb(n5417), .dout(n5424));
  jand g05199(.dina(n5424), .dinb(asqrt[59] ), .dout(n5425));
  jor  g05200(.dina(n5424), .dinb(asqrt[59] ), .dout(n5426));
  jxor g05201(.dina(n5066), .dinb(n443), .dout(n5427));
  jand g05202(.dina(n5427), .dinb(asqrt[36] ), .dout(n5428));
  jxor g05203(.dina(n5428), .dinb(n5072), .dout(n5429));
  jnot g05204(.din(n5429), .dout(n5430));
  jand g05205(.dina(n5430), .dinb(n5426), .dout(n5431));
  jor  g05206(.dina(n5431), .dinb(n5425), .dout(n5432));
  jand g05207(.dina(n5432), .dinb(asqrt[60] ), .dout(n5433));
  jor  g05208(.dina(n5432), .dinb(asqrt[60] ), .dout(n5434));
  jxor g05209(.dina(n5074), .dinb(n352), .dout(n5435));
  jand g05210(.dina(n5435), .dinb(asqrt[36] ), .dout(n5436));
  jxor g05211(.dina(n5436), .dinb(n5079), .dout(n5437));
  jnot g05212(.din(n5437), .dout(n5438));
  jand g05213(.dina(n5438), .dinb(n5434), .dout(n5439));
  jor  g05214(.dina(n5439), .dinb(n5433), .dout(n5440));
  jand g05215(.dina(n5440), .dinb(asqrt[61] ), .dout(n5441));
  jor  g05216(.dina(n5440), .dinb(asqrt[61] ), .dout(n5442));
  jxor g05217(.dina(n5081), .dinb(n294), .dout(n5443));
  jand g05218(.dina(n5443), .dinb(asqrt[36] ), .dout(n5444));
  jxor g05219(.dina(n5444), .dinb(n5086), .dout(n5445));
  jand g05220(.dina(n5445), .dinb(n5442), .dout(n5446));
  jor  g05221(.dina(n5446), .dinb(n5441), .dout(n5447));
  jand g05222(.dina(n5447), .dinb(asqrt[62] ), .dout(n5448));
  jor  g05223(.dina(n5447), .dinb(asqrt[62] ), .dout(n5449));
  jxor g05224(.dina(n5089), .dinb(n239), .dout(n5450));
  jand g05225(.dina(n5450), .dinb(asqrt[36] ), .dout(n5451));
  jxor g05226(.dina(n5451), .dinb(n5094), .dout(n5452));
  jnot g05227(.din(n5452), .dout(n5453));
  jand g05228(.dina(n5453), .dinb(n5449), .dout(n5454));
  jor  g05229(.dina(n5454), .dinb(n5448), .dout(n5455));
  jxor g05230(.dina(n5096), .dinb(n221), .dout(n5456));
  jand g05231(.dina(n5456), .dinb(asqrt[36] ), .dout(n5457));
  jxor g05232(.dina(n5457), .dinb(n5102), .dout(n5458));
  jnot g05233(.din(n5458), .dout(n5459));
  jor  g05234(.dina(n5459), .dinb(n5455), .dout(n5460));
  jnot g05235(.din(n5460), .dout(n5461));
  jand g05236(.dina(n5257), .dinb(n5104), .dout(n5462));
  jnot g05237(.din(n5462), .dout(n5463));
  jand g05238(.dina(n5108), .dinb(asqrt[63] ), .dout(n5464));
  jand g05239(.dina(n5464), .dinb(n5132), .dout(n5465));
  jand g05240(.dina(n5465), .dinb(n5463), .dout(n5466));
  jand g05241(.dina(n5118), .dinb(n5253), .dout(n5467));
  jnot g05242(.din(n5448), .dout(n5468));
  jnot g05243(.din(n5441), .dout(n5469));
  jnot g05244(.din(n5433), .dout(n5470));
  jnot g05245(.din(n5425), .dout(n5471));
  jnot g05246(.din(n5417), .dout(n5472));
  jnot g05247(.din(n5410), .dout(n5473));
  jnot g05248(.din(n5402), .dout(n5474));
  jnot g05249(.din(n5395), .dout(n5475));
  jnot g05250(.din(n5387), .dout(n5476));
  jnot g05251(.din(n5379), .dout(n5477));
  jnot g05252(.din(n5372), .dout(n5478));
  jnot g05253(.din(n5365), .dout(n5479));
  jnot g05254(.din(n5357), .dout(n5480));
  jnot g05255(.din(n5350), .dout(n5481));
  jnot g05256(.din(n5342), .dout(n5482));
  jnot g05257(.din(n5335), .dout(n5483));
  jnot g05258(.din(n5327), .dout(n5484));
  jnot g05259(.din(n5319), .dout(n5485));
  jnot g05260(.din(n5311), .dout(n5486));
  jnot g05261(.din(n5304), .dout(n5487));
  jnot g05262(.din(n5297), .dout(n5488));
  jnot g05263(.din(n5290), .dout(n5489));
  jnot g05264(.din(n5282), .dout(n5490));
  jnot g05265(.din(n5275), .dout(n5491));
  jnot g05266(.din(n5264), .dout(n5492));
  jnot g05267(.din(n5127), .dout(n5493));
  jnot g05268(.din(n5124), .dout(n5494));
  jor  g05269(.dina(n5259), .dinb(n4908), .dout(n5495));
  jand g05270(.dina(n5495), .dinb(n5494), .dout(n5496));
  jand g05271(.dina(n5496), .dinb(n4902), .dout(n5497));
  jor  g05272(.dina(n5259), .dinb(a[72] ), .dout(n5498));
  jand g05273(.dina(n5498), .dinb(a[73] ), .dout(n5499));
  jor  g05274(.dina(n5266), .dinb(n5499), .dout(n5500));
  jor  g05275(.dina(n5500), .dinb(n5497), .dout(n5501));
  jand g05276(.dina(n5501), .dinb(n5493), .dout(n5502));
  jand g05277(.dina(n5502), .dinb(n4582), .dout(n5503));
  jor  g05278(.dina(n5271), .dinb(n5503), .dout(n5504));
  jand g05279(.dina(n5504), .dinb(n5492), .dout(n5505));
  jand g05280(.dina(n5505), .dinb(n4249), .dout(n5506));
  jnot g05281(.din(n5279), .dout(n5507));
  jor  g05282(.dina(n5507), .dinb(n5506), .dout(n5508));
  jand g05283(.dina(n5508), .dinb(n5491), .dout(n5509));
  jand g05284(.dina(n5509), .dinb(n3955), .dout(n5510));
  jor  g05285(.dina(n5286), .dinb(n5510), .dout(n5511));
  jand g05286(.dina(n5511), .dinb(n5490), .dout(n5512));
  jand g05287(.dina(n5512), .dinb(n3642), .dout(n5513));
  jnot g05288(.din(n5294), .dout(n5514));
  jor  g05289(.dina(n5514), .dinb(n5513), .dout(n5515));
  jand g05290(.dina(n5515), .dinb(n5489), .dout(n5516));
  jand g05291(.dina(n5516), .dinb(n3368), .dout(n5517));
  jnot g05292(.din(n5301), .dout(n5518));
  jor  g05293(.dina(n5518), .dinb(n5517), .dout(n5519));
  jand g05294(.dina(n5519), .dinb(n5488), .dout(n5520));
  jand g05295(.dina(n5520), .dinb(n3089), .dout(n5521));
  jnot g05296(.din(n5308), .dout(n5522));
  jor  g05297(.dina(n5522), .dinb(n5521), .dout(n5523));
  jand g05298(.dina(n5523), .dinb(n5487), .dout(n5524));
  jand g05299(.dina(n5524), .dinb(n2833), .dout(n5525));
  jor  g05300(.dina(n5315), .dinb(n5525), .dout(n5526));
  jand g05301(.dina(n5526), .dinb(n5486), .dout(n5527));
  jand g05302(.dina(n5527), .dinb(n2572), .dout(n5528));
  jor  g05303(.dina(n5323), .dinb(n5528), .dout(n5529));
  jand g05304(.dina(n5529), .dinb(n5485), .dout(n5530));
  jand g05305(.dina(n5530), .dinb(n2345), .dout(n5531));
  jor  g05306(.dina(n5331), .dinb(n5531), .dout(n5532));
  jand g05307(.dina(n5532), .dinb(n5484), .dout(n5533));
  jand g05308(.dina(n5533), .dinb(n2108), .dout(n5534));
  jnot g05309(.din(n5339), .dout(n5535));
  jor  g05310(.dina(n5535), .dinb(n5534), .dout(n5536));
  jand g05311(.dina(n5536), .dinb(n5483), .dout(n5537));
  jand g05312(.dina(n5537), .dinb(n1912), .dout(n5538));
  jor  g05313(.dina(n5346), .dinb(n5538), .dout(n5539));
  jand g05314(.dina(n5539), .dinb(n5482), .dout(n5540));
  jand g05315(.dina(n5540), .dinb(n1699), .dout(n5541));
  jnot g05316(.din(n5354), .dout(n5542));
  jor  g05317(.dina(n5542), .dinb(n5541), .dout(n5543));
  jand g05318(.dina(n5543), .dinb(n5481), .dout(n5544));
  jand g05319(.dina(n5544), .dinb(n1516), .dout(n5545));
  jor  g05320(.dina(n5361), .dinb(n5545), .dout(n5546));
  jand g05321(.dina(n5546), .dinb(n5480), .dout(n5547));
  jand g05322(.dina(n5547), .dinb(n1332), .dout(n5548));
  jnot g05323(.din(n5369), .dout(n5549));
  jor  g05324(.dina(n5549), .dinb(n5548), .dout(n5550));
  jand g05325(.dina(n5550), .dinb(n5479), .dout(n5551));
  jand g05326(.dina(n5551), .dinb(n1173), .dout(n5552));
  jnot g05327(.din(n5376), .dout(n5553));
  jor  g05328(.dina(n5553), .dinb(n5552), .dout(n5554));
  jand g05329(.dina(n5554), .dinb(n5478), .dout(n5555));
  jand g05330(.dina(n5555), .dinb(n1008), .dout(n5556));
  jor  g05331(.dina(n5383), .dinb(n5556), .dout(n5557));
  jand g05332(.dina(n5557), .dinb(n5477), .dout(n5558));
  jand g05333(.dina(n5558), .dinb(n884), .dout(n5559));
  jor  g05334(.dina(n5391), .dinb(n5559), .dout(n5560));
  jand g05335(.dina(n5560), .dinb(n5476), .dout(n5561));
  jand g05336(.dina(n5561), .dinb(n743), .dout(n5562));
  jnot g05337(.din(n5399), .dout(n5563));
  jor  g05338(.dina(n5563), .dinb(n5562), .dout(n5564));
  jand g05339(.dina(n5564), .dinb(n5475), .dout(n5565));
  jand g05340(.dina(n5565), .dinb(n635), .dout(n5566));
  jor  g05341(.dina(n5406), .dinb(n5566), .dout(n5567));
  jand g05342(.dina(n5567), .dinb(n5474), .dout(n5568));
  jand g05343(.dina(n5568), .dinb(n515), .dout(n5569));
  jnot g05344(.din(n5414), .dout(n5570));
  jor  g05345(.dina(n5570), .dinb(n5569), .dout(n5571));
  jand g05346(.dina(n5571), .dinb(n5473), .dout(n5572));
  jand g05347(.dina(n5572), .dinb(n443), .dout(n5573));
  jor  g05348(.dina(n5421), .dinb(n5573), .dout(n5574));
  jand g05349(.dina(n5574), .dinb(n5472), .dout(n5575));
  jand g05350(.dina(n5575), .dinb(n352), .dout(n5576));
  jor  g05351(.dina(n5429), .dinb(n5576), .dout(n5577));
  jand g05352(.dina(n5577), .dinb(n5471), .dout(n5578));
  jand g05353(.dina(n5578), .dinb(n294), .dout(n5579));
  jor  g05354(.dina(n5437), .dinb(n5579), .dout(n5580));
  jand g05355(.dina(n5580), .dinb(n5470), .dout(n5581));
  jand g05356(.dina(n5581), .dinb(n239), .dout(n5582));
  jnot g05357(.din(n5445), .dout(n5583));
  jor  g05358(.dina(n5583), .dinb(n5582), .dout(n5584));
  jand g05359(.dina(n5584), .dinb(n5469), .dout(n5585));
  jand g05360(.dina(n5585), .dinb(n221), .dout(n5586));
  jor  g05361(.dina(n5452), .dinb(n5586), .dout(n5587));
  jand g05362(.dina(n5587), .dinb(n5468), .dout(n5588));
  jor  g05363(.dina(n5458), .dinb(n5588), .dout(n5589));
  jor  g05364(.dina(n5589), .dinb(n5105), .dout(n5590));
  jor  g05365(.dina(n5590), .dinb(n5467), .dout(n5591));
  jand g05366(.dina(n5591), .dinb(n218), .dout(n5592));
  jand g05367(.dina(n5259), .dinb(n4906), .dout(n5593));
  jor  g05368(.dina(n5593), .dinb(n5592), .dout(n5594));
  jor  g05369(.dina(n5594), .dinb(n5466), .dout(n5595));
  jor  g05370(.dina(n5595), .dinb(n5461), .dout(asqrt[35] ));
  jnot g05371(.din(n5466), .dout(n5597));
  jnot g05372(.din(n5467), .dout(n5598));
  jand g05373(.dina(n5459), .dinb(n5455), .dout(n5599));
  jand g05374(.dina(n5599), .dinb(n5132), .dout(n5600));
  jand g05375(.dina(n5600), .dinb(n5598), .dout(n5601));
  jor  g05376(.dina(n5601), .dinb(asqrt[63] ), .dout(n5602));
  jnot g05377(.din(n5593), .dout(n5603));
  jand g05378(.dina(n5603), .dinb(n5602), .dout(n5604));
  jand g05379(.dina(n5604), .dinb(n5597), .dout(n5605));
  jand g05380(.dina(n5605), .dinb(n5460), .dout(n5606));
  jxor g05381(.dina(n5447), .dinb(n221), .dout(n5607));
  jor  g05382(.dina(n5607), .dinb(n5606), .dout(n5608));
  jxor g05383(.dina(n5608), .dinb(n5452), .dout(n5609));
  jnot g05384(.din(n5609), .dout(n5610));
  jor  g05385(.dina(n5606), .dinb(n5121), .dout(n5611));
  jnot g05386(.din(a[68] ), .dout(n5612));
  jnot g05387(.din(a[69] ), .dout(n5613));
  jand g05388(.dina(n5613), .dinb(n5612), .dout(n5614));
  jand g05389(.dina(n5614), .dinb(n5121), .dout(n5615));
  jnot g05390(.din(n5615), .dout(n5616));
  jand g05391(.dina(n5616), .dinb(n5611), .dout(n5617));
  jor  g05392(.dina(n5617), .dinb(n5259), .dout(n5618));
  jand g05393(.dina(n5617), .dinb(n5259), .dout(n5619));
  jor  g05394(.dina(n5606), .dinb(a[70] ), .dout(n5620));
  jand g05395(.dina(n5620), .dinb(a[71] ), .dout(n5621));
  jand g05396(.dina(asqrt[35] ), .dinb(n5123), .dout(n5622));
  jor  g05397(.dina(n5622), .dinb(n5621), .dout(n5623));
  jor  g05398(.dina(n5623), .dinb(n5619), .dout(n5624));
  jand g05399(.dina(n5624), .dinb(n5618), .dout(n5625));
  jor  g05400(.dina(n5625), .dinb(n4902), .dout(n5626));
  jand g05401(.dina(n5625), .dinb(n4902), .dout(n5627));
  jnot g05402(.din(n5123), .dout(n5628));
  jor  g05403(.dina(n5606), .dinb(n5628), .dout(n5629));
  jor  g05404(.dina(n5461), .dinb(n5259), .dout(n5630));
  jor  g05405(.dina(n5630), .dinb(n5465), .dout(n5631));
  jor  g05406(.dina(n5631), .dinb(n5592), .dout(n5632));
  jand g05407(.dina(n5632), .dinb(n5629), .dout(n5633));
  jxor g05408(.dina(n5633), .dinb(n4908), .dout(n5634));
  jor  g05409(.dina(n5634), .dinb(n5627), .dout(n5635));
  jand g05410(.dina(n5635), .dinb(n5626), .dout(n5636));
  jor  g05411(.dina(n5636), .dinb(n4582), .dout(n5637));
  jand g05412(.dina(n5636), .dinb(n4582), .dout(n5638));
  jxor g05413(.dina(n5126), .dinb(n4902), .dout(n5639));
  jor  g05414(.dina(n5639), .dinb(n5606), .dout(n5640));
  jxor g05415(.dina(n5640), .dinb(n5500), .dout(n5641));
  jnot g05416(.din(n5641), .dout(n5642));
  jor  g05417(.dina(n5642), .dinb(n5638), .dout(n5643));
  jand g05418(.dina(n5643), .dinb(n5637), .dout(n5644));
  jor  g05419(.dina(n5644), .dinb(n4249), .dout(n5645));
  jand g05420(.dina(n5644), .dinb(n4249), .dout(n5646));
  jxor g05421(.dina(n5263), .dinb(n4582), .dout(n5647));
  jor  g05422(.dina(n5647), .dinb(n5606), .dout(n5648));
  jxor g05423(.dina(n5648), .dinb(n5272), .dout(n5649));
  jor  g05424(.dina(n5649), .dinb(n5646), .dout(n5650));
  jand g05425(.dina(n5650), .dinb(n5645), .dout(n5651));
  jor  g05426(.dina(n5651), .dinb(n3955), .dout(n5652));
  jand g05427(.dina(n5651), .dinb(n3955), .dout(n5653));
  jxor g05428(.dina(n5274), .dinb(n4249), .dout(n5654));
  jor  g05429(.dina(n5654), .dinb(n5606), .dout(n5655));
  jxor g05430(.dina(n5655), .dinb(n5507), .dout(n5656));
  jnot g05431(.din(n5656), .dout(n5657));
  jor  g05432(.dina(n5657), .dinb(n5653), .dout(n5658));
  jand g05433(.dina(n5658), .dinb(n5652), .dout(n5659));
  jor  g05434(.dina(n5659), .dinb(n3642), .dout(n5660));
  jand g05435(.dina(n5659), .dinb(n3642), .dout(n5661));
  jxor g05436(.dina(n5281), .dinb(n3955), .dout(n5662));
  jor  g05437(.dina(n5662), .dinb(n5606), .dout(n5663));
  jxor g05438(.dina(n5663), .dinb(n5287), .dout(n5664));
  jor  g05439(.dina(n5664), .dinb(n5661), .dout(n5665));
  jand g05440(.dina(n5665), .dinb(n5660), .dout(n5666));
  jor  g05441(.dina(n5666), .dinb(n3368), .dout(n5667));
  jand g05442(.dina(n5666), .dinb(n3368), .dout(n5668));
  jxor g05443(.dina(n5289), .dinb(n3642), .dout(n5669));
  jor  g05444(.dina(n5669), .dinb(n5606), .dout(n5670));
  jxor g05445(.dina(n5670), .dinb(n5514), .dout(n5671));
  jnot g05446(.din(n5671), .dout(n5672));
  jor  g05447(.dina(n5672), .dinb(n5668), .dout(n5673));
  jand g05448(.dina(n5673), .dinb(n5667), .dout(n5674));
  jor  g05449(.dina(n5674), .dinb(n3089), .dout(n5675));
  jand g05450(.dina(n5674), .dinb(n3089), .dout(n5676));
  jxor g05451(.dina(n5296), .dinb(n3368), .dout(n5677));
  jor  g05452(.dina(n5677), .dinb(n5606), .dout(n5678));
  jxor g05453(.dina(n5678), .dinb(n5518), .dout(n5679));
  jnot g05454(.din(n5679), .dout(n5680));
  jor  g05455(.dina(n5680), .dinb(n5676), .dout(n5681));
  jand g05456(.dina(n5681), .dinb(n5675), .dout(n5682));
  jor  g05457(.dina(n5682), .dinb(n2833), .dout(n5683));
  jand g05458(.dina(n5682), .dinb(n2833), .dout(n5684));
  jxor g05459(.dina(n5303), .dinb(n3089), .dout(n5685));
  jor  g05460(.dina(n5685), .dinb(n5606), .dout(n5686));
  jxor g05461(.dina(n5686), .dinb(n5522), .dout(n5687));
  jnot g05462(.din(n5687), .dout(n5688));
  jor  g05463(.dina(n5688), .dinb(n5684), .dout(n5689));
  jand g05464(.dina(n5689), .dinb(n5683), .dout(n5690));
  jor  g05465(.dina(n5690), .dinb(n2572), .dout(n5691));
  jand g05466(.dina(n5690), .dinb(n2572), .dout(n5692));
  jxor g05467(.dina(n5310), .dinb(n2833), .dout(n5693));
  jor  g05468(.dina(n5693), .dinb(n5606), .dout(n5694));
  jxor g05469(.dina(n5694), .dinb(n5316), .dout(n5695));
  jor  g05470(.dina(n5695), .dinb(n5692), .dout(n5696));
  jand g05471(.dina(n5696), .dinb(n5691), .dout(n5697));
  jor  g05472(.dina(n5697), .dinb(n2345), .dout(n5698));
  jand g05473(.dina(n5697), .dinb(n2345), .dout(n5699));
  jxor g05474(.dina(n5318), .dinb(n2572), .dout(n5700));
  jor  g05475(.dina(n5700), .dinb(n5606), .dout(n5701));
  jxor g05476(.dina(n5701), .dinb(n5324), .dout(n5702));
  jor  g05477(.dina(n5702), .dinb(n5699), .dout(n5703));
  jand g05478(.dina(n5703), .dinb(n5698), .dout(n5704));
  jor  g05479(.dina(n5704), .dinb(n2108), .dout(n5705));
  jand g05480(.dina(n5704), .dinb(n2108), .dout(n5706));
  jxor g05481(.dina(n5326), .dinb(n2345), .dout(n5707));
  jor  g05482(.dina(n5707), .dinb(n5606), .dout(n5708));
  jxor g05483(.dina(n5708), .dinb(n5332), .dout(n5709));
  jor  g05484(.dina(n5709), .dinb(n5706), .dout(n5710));
  jand g05485(.dina(n5710), .dinb(n5705), .dout(n5711));
  jor  g05486(.dina(n5711), .dinb(n1912), .dout(n5712));
  jand g05487(.dina(n5711), .dinb(n1912), .dout(n5713));
  jxor g05488(.dina(n5334), .dinb(n2108), .dout(n5714));
  jor  g05489(.dina(n5714), .dinb(n5606), .dout(n5715));
  jxor g05490(.dina(n5715), .dinb(n5535), .dout(n5716));
  jnot g05491(.din(n5716), .dout(n5717));
  jor  g05492(.dina(n5717), .dinb(n5713), .dout(n5718));
  jand g05493(.dina(n5718), .dinb(n5712), .dout(n5719));
  jor  g05494(.dina(n5719), .dinb(n1699), .dout(n5720));
  jand g05495(.dina(n5719), .dinb(n1699), .dout(n5721));
  jxor g05496(.dina(n5341), .dinb(n1912), .dout(n5722));
  jor  g05497(.dina(n5722), .dinb(n5606), .dout(n5723));
  jxor g05498(.dina(n5723), .dinb(n5347), .dout(n5724));
  jor  g05499(.dina(n5724), .dinb(n5721), .dout(n5725));
  jand g05500(.dina(n5725), .dinb(n5720), .dout(n5726));
  jor  g05501(.dina(n5726), .dinb(n1516), .dout(n5727));
  jand g05502(.dina(n5726), .dinb(n1516), .dout(n5728));
  jxor g05503(.dina(n5349), .dinb(n1699), .dout(n5729));
  jor  g05504(.dina(n5729), .dinb(n5606), .dout(n5730));
  jxor g05505(.dina(n5730), .dinb(n5542), .dout(n5731));
  jnot g05506(.din(n5731), .dout(n5732));
  jor  g05507(.dina(n5732), .dinb(n5728), .dout(n5733));
  jand g05508(.dina(n5733), .dinb(n5727), .dout(n5734));
  jor  g05509(.dina(n5734), .dinb(n1332), .dout(n5735));
  jand g05510(.dina(n5734), .dinb(n1332), .dout(n5736));
  jxor g05511(.dina(n5356), .dinb(n1516), .dout(n5737));
  jor  g05512(.dina(n5737), .dinb(n5606), .dout(n5738));
  jxor g05513(.dina(n5738), .dinb(n5362), .dout(n5739));
  jor  g05514(.dina(n5739), .dinb(n5736), .dout(n5740));
  jand g05515(.dina(n5740), .dinb(n5735), .dout(n5741));
  jor  g05516(.dina(n5741), .dinb(n1173), .dout(n5742));
  jand g05517(.dina(n5741), .dinb(n1173), .dout(n5743));
  jxor g05518(.dina(n5364), .dinb(n1332), .dout(n5744));
  jor  g05519(.dina(n5744), .dinb(n5606), .dout(n5745));
  jxor g05520(.dina(n5745), .dinb(n5549), .dout(n5746));
  jnot g05521(.din(n5746), .dout(n5747));
  jor  g05522(.dina(n5747), .dinb(n5743), .dout(n5748));
  jand g05523(.dina(n5748), .dinb(n5742), .dout(n5749));
  jor  g05524(.dina(n5749), .dinb(n1008), .dout(n5750));
  jand g05525(.dina(n5749), .dinb(n1008), .dout(n5751));
  jxor g05526(.dina(n5371), .dinb(n1173), .dout(n5752));
  jor  g05527(.dina(n5752), .dinb(n5606), .dout(n5753));
  jxor g05528(.dina(n5753), .dinb(n5553), .dout(n5754));
  jnot g05529(.din(n5754), .dout(n5755));
  jor  g05530(.dina(n5755), .dinb(n5751), .dout(n5756));
  jand g05531(.dina(n5756), .dinb(n5750), .dout(n5757));
  jor  g05532(.dina(n5757), .dinb(n884), .dout(n5758));
  jand g05533(.dina(n5757), .dinb(n884), .dout(n5759));
  jxor g05534(.dina(n5378), .dinb(n1008), .dout(n5760));
  jor  g05535(.dina(n5760), .dinb(n5606), .dout(n5761));
  jxor g05536(.dina(n5761), .dinb(n5384), .dout(n5762));
  jor  g05537(.dina(n5762), .dinb(n5759), .dout(n5763));
  jand g05538(.dina(n5763), .dinb(n5758), .dout(n5764));
  jor  g05539(.dina(n5764), .dinb(n743), .dout(n5765));
  jand g05540(.dina(n5764), .dinb(n743), .dout(n5766));
  jxor g05541(.dina(n5386), .dinb(n884), .dout(n5767));
  jor  g05542(.dina(n5767), .dinb(n5606), .dout(n5768));
  jxor g05543(.dina(n5768), .dinb(n5392), .dout(n5769));
  jor  g05544(.dina(n5769), .dinb(n5766), .dout(n5770));
  jand g05545(.dina(n5770), .dinb(n5765), .dout(n5771));
  jor  g05546(.dina(n5771), .dinb(n635), .dout(n5772));
  jand g05547(.dina(n5771), .dinb(n635), .dout(n5773));
  jxor g05548(.dina(n5394), .dinb(n743), .dout(n5774));
  jor  g05549(.dina(n5774), .dinb(n5606), .dout(n5775));
  jxor g05550(.dina(n5775), .dinb(n5563), .dout(n5776));
  jnot g05551(.din(n5776), .dout(n5777));
  jor  g05552(.dina(n5777), .dinb(n5773), .dout(n5778));
  jand g05553(.dina(n5778), .dinb(n5772), .dout(n5779));
  jor  g05554(.dina(n5779), .dinb(n515), .dout(n5780));
  jand g05555(.dina(n5779), .dinb(n515), .dout(n5781));
  jxor g05556(.dina(n5401), .dinb(n635), .dout(n5782));
  jor  g05557(.dina(n5782), .dinb(n5606), .dout(n5783));
  jxor g05558(.dina(n5783), .dinb(n5407), .dout(n5784));
  jor  g05559(.dina(n5784), .dinb(n5781), .dout(n5785));
  jand g05560(.dina(n5785), .dinb(n5780), .dout(n5786));
  jor  g05561(.dina(n5786), .dinb(n443), .dout(n5787));
  jand g05562(.dina(n5786), .dinb(n443), .dout(n5788));
  jxor g05563(.dina(n5409), .dinb(n515), .dout(n5789));
  jor  g05564(.dina(n5789), .dinb(n5606), .dout(n5790));
  jxor g05565(.dina(n5790), .dinb(n5570), .dout(n5791));
  jnot g05566(.din(n5791), .dout(n5792));
  jor  g05567(.dina(n5792), .dinb(n5788), .dout(n5793));
  jand g05568(.dina(n5793), .dinb(n5787), .dout(n5794));
  jor  g05569(.dina(n5794), .dinb(n352), .dout(n5795));
  jand g05570(.dina(n5794), .dinb(n352), .dout(n5796));
  jxor g05571(.dina(n5416), .dinb(n443), .dout(n5797));
  jor  g05572(.dina(n5797), .dinb(n5606), .dout(n5798));
  jxor g05573(.dina(n5798), .dinb(n5422), .dout(n5799));
  jor  g05574(.dina(n5799), .dinb(n5796), .dout(n5800));
  jand g05575(.dina(n5800), .dinb(n5795), .dout(n5801));
  jor  g05576(.dina(n5801), .dinb(n294), .dout(n5802));
  jand g05577(.dina(n5801), .dinb(n294), .dout(n5803));
  jxor g05578(.dina(n5424), .dinb(n352), .dout(n5804));
  jor  g05579(.dina(n5804), .dinb(n5606), .dout(n5805));
  jxor g05580(.dina(n5805), .dinb(n5430), .dout(n5806));
  jor  g05581(.dina(n5806), .dinb(n5803), .dout(n5807));
  jand g05582(.dina(n5807), .dinb(n5802), .dout(n5808));
  jor  g05583(.dina(n5808), .dinb(n239), .dout(n5809));
  jand g05584(.dina(n5808), .dinb(n239), .dout(n5810));
  jxor g05585(.dina(n5432), .dinb(n294), .dout(n5811));
  jor  g05586(.dina(n5811), .dinb(n5606), .dout(n5812));
  jxor g05587(.dina(n5812), .dinb(n5438), .dout(n5813));
  jor  g05588(.dina(n5813), .dinb(n5810), .dout(n5814));
  jand g05589(.dina(n5814), .dinb(n5809), .dout(n5815));
  jor  g05590(.dina(n5815), .dinb(n221), .dout(n5816));
  jand g05591(.dina(n5815), .dinb(n221), .dout(n5817));
  jxor g05592(.dina(n5440), .dinb(n239), .dout(n5818));
  jor  g05593(.dina(n5818), .dinb(n5606), .dout(n5819));
  jxor g05594(.dina(n5819), .dinb(n5583), .dout(n5820));
  jnot g05595(.din(n5820), .dout(n5821));
  jor  g05596(.dina(n5821), .dinb(n5817), .dout(n5822));
  jand g05597(.dina(n5822), .dinb(n5816), .dout(n5823));
  jand g05598(.dina(n5823), .dinb(n5610), .dout(n5824));
  jor  g05599(.dina(n5823), .dinb(n5610), .dout(n5826));
  jxor g05600(.dina(n5459), .dinb(n5455), .dout(n5827));
  jnot g05601(.din(n5827), .dout(n5828));
  jand g05602(.dina(n5828), .dinb(asqrt[35] ), .dout(n5829));
  jor  g05603(.dina(n5829), .dinb(n5826), .dout(n5830));
  jand g05604(.dina(n5830), .dinb(n218), .dout(n5831));
  jand g05605(.dina(n5605), .dinb(n5588), .dout(n5832));
  jand g05606(.dina(n5827), .dinb(asqrt[63] ), .dout(n5833));
  jnot g05607(.din(n5833), .dout(n5834));
  jor  g05608(.dina(n5834), .dinb(n5832), .dout(n5835));
  jnot g05609(.din(n5835), .dout(n5836));
  jor  g05610(.dina(n5836), .dinb(n5831), .dout(n5837));
  jor  g05611(.dina(n5837), .dinb(n5824), .dout(asqrt[34] ));
  jxor g05612(.dina(n5815), .dinb(n221), .dout(n5840));
  jand g05613(.dina(n5840), .dinb(asqrt[34] ), .dout(n5841));
  jxor g05614(.dina(n5841), .dinb(n5820), .dout(n5842));
  jnot g05615(.din(a[66] ), .dout(n5843));
  jnot g05616(.din(a[67] ), .dout(n5844));
  jand g05617(.dina(n5844), .dinb(n5843), .dout(n5845));
  jand g05618(.dina(n5845), .dinb(n5612), .dout(n5846));
  jand g05619(.dina(asqrt[34] ), .dinb(a[68] ), .dout(n5847));
  jor  g05620(.dina(n5847), .dinb(n5846), .dout(n5848));
  jand g05621(.dina(n5848), .dinb(asqrt[35] ), .dout(n5849));
  jor  g05622(.dina(n5848), .dinb(asqrt[35] ), .dout(n5850));
  jand g05623(.dina(asqrt[34] ), .dinb(n5612), .dout(n5851));
  jor  g05624(.dina(n5851), .dinb(n5613), .dout(n5852));
  jnot g05625(.din(n5614), .dout(n5853));
  jnot g05626(.din(n5824), .dout(n5854));
  jnot g05627(.din(n5816), .dout(n5856));
  jnot g05628(.din(n5809), .dout(n5857));
  jnot g05629(.din(n5802), .dout(n5858));
  jnot g05630(.din(n5795), .dout(n5859));
  jnot g05631(.din(n5787), .dout(n5860));
  jnot g05632(.din(n5780), .dout(n5861));
  jnot g05633(.din(n5772), .dout(n5862));
  jnot g05634(.din(n5765), .dout(n5863));
  jnot g05635(.din(n5758), .dout(n5864));
  jnot g05636(.din(n5750), .dout(n5865));
  jnot g05637(.din(n5742), .dout(n5866));
  jnot g05638(.din(n5735), .dout(n5867));
  jnot g05639(.din(n5727), .dout(n5868));
  jnot g05640(.din(n5720), .dout(n5869));
  jnot g05641(.din(n5712), .dout(n5870));
  jnot g05642(.din(n5705), .dout(n5871));
  jnot g05643(.din(n5698), .dout(n5872));
  jnot g05644(.din(n5691), .dout(n5873));
  jnot g05645(.din(n5683), .dout(n5874));
  jnot g05646(.din(n5675), .dout(n5875));
  jnot g05647(.din(n5667), .dout(n5876));
  jnot g05648(.din(n5660), .dout(n5877));
  jnot g05649(.din(n5652), .dout(n5878));
  jnot g05650(.din(n5645), .dout(n5879));
  jnot g05651(.din(n5637), .dout(n5880));
  jnot g05652(.din(n5626), .dout(n5881));
  jnot g05653(.din(n5618), .dout(n5882));
  jand g05654(.dina(asqrt[35] ), .dinb(a[70] ), .dout(n5883));
  jor  g05655(.dina(n5615), .dinb(n5883), .dout(n5884));
  jor  g05656(.dina(n5884), .dinb(asqrt[36] ), .dout(n5885));
  jand g05657(.dina(asqrt[35] ), .dinb(n5121), .dout(n5886));
  jor  g05658(.dina(n5886), .dinb(n5122), .dout(n5887));
  jand g05659(.dina(n5629), .dinb(n5887), .dout(n5888));
  jand g05660(.dina(n5888), .dinb(n5885), .dout(n5889));
  jor  g05661(.dina(n5889), .dinb(n5882), .dout(n5890));
  jor  g05662(.dina(n5890), .dinb(asqrt[37] ), .dout(n5891));
  jnot g05663(.din(n5634), .dout(n5892));
  jand g05664(.dina(n5892), .dinb(n5891), .dout(n5893));
  jor  g05665(.dina(n5893), .dinb(n5881), .dout(n5894));
  jor  g05666(.dina(n5894), .dinb(asqrt[38] ), .dout(n5895));
  jand g05667(.dina(n5641), .dinb(n5895), .dout(n5896));
  jor  g05668(.dina(n5896), .dinb(n5880), .dout(n5897));
  jor  g05669(.dina(n5897), .dinb(asqrt[39] ), .dout(n5898));
  jnot g05670(.din(n5649), .dout(n5899));
  jand g05671(.dina(n5899), .dinb(n5898), .dout(n5900));
  jor  g05672(.dina(n5900), .dinb(n5879), .dout(n5901));
  jor  g05673(.dina(n5901), .dinb(asqrt[40] ), .dout(n5902));
  jand g05674(.dina(n5656), .dinb(n5902), .dout(n5903));
  jor  g05675(.dina(n5903), .dinb(n5878), .dout(n5904));
  jor  g05676(.dina(n5904), .dinb(asqrt[41] ), .dout(n5905));
  jnot g05677(.din(n5664), .dout(n5906));
  jand g05678(.dina(n5906), .dinb(n5905), .dout(n5907));
  jor  g05679(.dina(n5907), .dinb(n5877), .dout(n5908));
  jor  g05680(.dina(n5908), .dinb(asqrt[42] ), .dout(n5909));
  jand g05681(.dina(n5671), .dinb(n5909), .dout(n5910));
  jor  g05682(.dina(n5910), .dinb(n5876), .dout(n5911));
  jor  g05683(.dina(n5911), .dinb(asqrt[43] ), .dout(n5912));
  jand g05684(.dina(n5679), .dinb(n5912), .dout(n5913));
  jor  g05685(.dina(n5913), .dinb(n5875), .dout(n5914));
  jor  g05686(.dina(n5914), .dinb(asqrt[44] ), .dout(n5915));
  jand g05687(.dina(n5687), .dinb(n5915), .dout(n5916));
  jor  g05688(.dina(n5916), .dinb(n5874), .dout(n5917));
  jor  g05689(.dina(n5917), .dinb(asqrt[45] ), .dout(n5918));
  jnot g05690(.din(n5695), .dout(n5919));
  jand g05691(.dina(n5919), .dinb(n5918), .dout(n5920));
  jor  g05692(.dina(n5920), .dinb(n5873), .dout(n5921));
  jor  g05693(.dina(n5921), .dinb(asqrt[46] ), .dout(n5922));
  jnot g05694(.din(n5702), .dout(n5923));
  jand g05695(.dina(n5923), .dinb(n5922), .dout(n5924));
  jor  g05696(.dina(n5924), .dinb(n5872), .dout(n5925));
  jor  g05697(.dina(n5925), .dinb(asqrt[47] ), .dout(n5926));
  jnot g05698(.din(n5709), .dout(n5927));
  jand g05699(.dina(n5927), .dinb(n5926), .dout(n5928));
  jor  g05700(.dina(n5928), .dinb(n5871), .dout(n5929));
  jor  g05701(.dina(n5929), .dinb(asqrt[48] ), .dout(n5930));
  jand g05702(.dina(n5716), .dinb(n5930), .dout(n5931));
  jor  g05703(.dina(n5931), .dinb(n5870), .dout(n5932));
  jor  g05704(.dina(n5932), .dinb(asqrt[49] ), .dout(n5933));
  jnot g05705(.din(n5724), .dout(n5934));
  jand g05706(.dina(n5934), .dinb(n5933), .dout(n5935));
  jor  g05707(.dina(n5935), .dinb(n5869), .dout(n5936));
  jor  g05708(.dina(n5936), .dinb(asqrt[50] ), .dout(n5937));
  jand g05709(.dina(n5731), .dinb(n5937), .dout(n5938));
  jor  g05710(.dina(n5938), .dinb(n5868), .dout(n5939));
  jor  g05711(.dina(n5939), .dinb(asqrt[51] ), .dout(n5940));
  jnot g05712(.din(n5739), .dout(n5941));
  jand g05713(.dina(n5941), .dinb(n5940), .dout(n5942));
  jor  g05714(.dina(n5942), .dinb(n5867), .dout(n5943));
  jor  g05715(.dina(n5943), .dinb(asqrt[52] ), .dout(n5944));
  jand g05716(.dina(n5746), .dinb(n5944), .dout(n5945));
  jor  g05717(.dina(n5945), .dinb(n5866), .dout(n5946));
  jor  g05718(.dina(n5946), .dinb(asqrt[53] ), .dout(n5947));
  jand g05719(.dina(n5754), .dinb(n5947), .dout(n5948));
  jor  g05720(.dina(n5948), .dinb(n5865), .dout(n5949));
  jor  g05721(.dina(n5949), .dinb(asqrt[54] ), .dout(n5950));
  jnot g05722(.din(n5762), .dout(n5951));
  jand g05723(.dina(n5951), .dinb(n5950), .dout(n5952));
  jor  g05724(.dina(n5952), .dinb(n5864), .dout(n5953));
  jor  g05725(.dina(n5953), .dinb(asqrt[55] ), .dout(n5954));
  jnot g05726(.din(n5769), .dout(n5955));
  jand g05727(.dina(n5955), .dinb(n5954), .dout(n5956));
  jor  g05728(.dina(n5956), .dinb(n5863), .dout(n5957));
  jor  g05729(.dina(n5957), .dinb(asqrt[56] ), .dout(n5958));
  jand g05730(.dina(n5776), .dinb(n5958), .dout(n5959));
  jor  g05731(.dina(n5959), .dinb(n5862), .dout(n5960));
  jor  g05732(.dina(n5960), .dinb(asqrt[57] ), .dout(n5961));
  jnot g05733(.din(n5784), .dout(n5962));
  jand g05734(.dina(n5962), .dinb(n5961), .dout(n5963));
  jor  g05735(.dina(n5963), .dinb(n5861), .dout(n5964));
  jor  g05736(.dina(n5964), .dinb(asqrt[58] ), .dout(n5965));
  jand g05737(.dina(n5791), .dinb(n5965), .dout(n5966));
  jor  g05738(.dina(n5966), .dinb(n5860), .dout(n5967));
  jor  g05739(.dina(n5967), .dinb(asqrt[59] ), .dout(n5968));
  jnot g05740(.din(n5799), .dout(n5969));
  jand g05741(.dina(n5969), .dinb(n5968), .dout(n5970));
  jor  g05742(.dina(n5970), .dinb(n5859), .dout(n5971));
  jor  g05743(.dina(n5971), .dinb(asqrt[60] ), .dout(n5972));
  jnot g05744(.din(n5806), .dout(n5973));
  jand g05745(.dina(n5973), .dinb(n5972), .dout(n5974));
  jor  g05746(.dina(n5974), .dinb(n5858), .dout(n5975));
  jor  g05747(.dina(n5975), .dinb(asqrt[61] ), .dout(n5976));
  jnot g05748(.din(n5813), .dout(n5977));
  jand g05749(.dina(n5977), .dinb(n5976), .dout(n5978));
  jor  g05750(.dina(n5978), .dinb(n5857), .dout(n5979));
  jor  g05751(.dina(n5979), .dinb(asqrt[62] ), .dout(n5980));
  jand g05752(.dina(n5820), .dinb(n5980), .dout(n5981));
  jor  g05753(.dina(n5981), .dinb(n5856), .dout(n5982));
  jand g05754(.dina(n5982), .dinb(n5609), .dout(n5983));
  jnot g05755(.din(n5829), .dout(n5984));
  jand g05756(.dina(n5984), .dinb(n5983), .dout(n5985));
  jor  g05757(.dina(n5985), .dinb(asqrt[63] ), .dout(n5986));
  jand g05758(.dina(n5835), .dinb(n5986), .dout(n5987));
  jand g05759(.dina(n5987), .dinb(n5854), .dout(n5989));
  jor  g05760(.dina(n5989), .dinb(n5853), .dout(n5990));
  jand g05761(.dina(n5990), .dinb(n5852), .dout(n5991));
  jand g05762(.dina(n5991), .dinb(n5850), .dout(n5992));
  jor  g05763(.dina(n5992), .dinb(n5849), .dout(n5993));
  jand g05764(.dina(n5993), .dinb(asqrt[36] ), .dout(n5994));
  jor  g05765(.dina(n5993), .dinb(asqrt[36] ), .dout(n5995));
  jand g05766(.dina(asqrt[34] ), .dinb(n5614), .dout(n5996));
  jand g05767(.dina(n5986), .dinb(asqrt[35] ), .dout(n5997));
  jand g05768(.dina(n5997), .dinb(n5834), .dout(n5998));
  jand g05769(.dina(n5998), .dinb(n5854), .dout(n5999));
  jor  g05770(.dina(n5999), .dinb(n5996), .dout(n6000));
  jxor g05771(.dina(n6000), .dinb(a[70] ), .dout(n6001));
  jnot g05772(.din(n6001), .dout(n6002));
  jand g05773(.dina(n6002), .dinb(n5995), .dout(n6003));
  jor  g05774(.dina(n6003), .dinb(n5994), .dout(n6004));
  jand g05775(.dina(n6004), .dinb(asqrt[37] ), .dout(n6005));
  jor  g05776(.dina(n6004), .dinb(asqrt[37] ), .dout(n6006));
  jxor g05777(.dina(n5617), .dinb(n5259), .dout(n6007));
  jand g05778(.dina(n6007), .dinb(asqrt[34] ), .dout(n6008));
  jxor g05779(.dina(n6008), .dinb(n5888), .dout(n6009));
  jand g05780(.dina(n6009), .dinb(n6006), .dout(n6010));
  jor  g05781(.dina(n6010), .dinb(n6005), .dout(n6011));
  jand g05782(.dina(n6011), .dinb(asqrt[38] ), .dout(n6012));
  jor  g05783(.dina(n6011), .dinb(asqrt[38] ), .dout(n6013));
  jxor g05784(.dina(n5625), .dinb(n4902), .dout(n6014));
  jand g05785(.dina(n6014), .dinb(asqrt[34] ), .dout(n6015));
  jxor g05786(.dina(n6015), .dinb(n5634), .dout(n6016));
  jnot g05787(.din(n6016), .dout(n6017));
  jand g05788(.dina(n6017), .dinb(n6013), .dout(n6018));
  jor  g05789(.dina(n6018), .dinb(n6012), .dout(n6019));
  jand g05790(.dina(n6019), .dinb(asqrt[39] ), .dout(n6020));
  jor  g05791(.dina(n6019), .dinb(asqrt[39] ), .dout(n6021));
  jxor g05792(.dina(n5636), .dinb(n4582), .dout(n6022));
  jand g05793(.dina(n6022), .dinb(asqrt[34] ), .dout(n6023));
  jxor g05794(.dina(n6023), .dinb(n5641), .dout(n6024));
  jand g05795(.dina(n6024), .dinb(n6021), .dout(n6025));
  jor  g05796(.dina(n6025), .dinb(n6020), .dout(n6026));
  jand g05797(.dina(n6026), .dinb(asqrt[40] ), .dout(n6027));
  jor  g05798(.dina(n6026), .dinb(asqrt[40] ), .dout(n6028));
  jxor g05799(.dina(n5644), .dinb(n4249), .dout(n6029));
  jand g05800(.dina(n6029), .dinb(asqrt[34] ), .dout(n6030));
  jxor g05801(.dina(n6030), .dinb(n5649), .dout(n6031));
  jnot g05802(.din(n6031), .dout(n6032));
  jand g05803(.dina(n6032), .dinb(n6028), .dout(n6033));
  jor  g05804(.dina(n6033), .dinb(n6027), .dout(n6034));
  jand g05805(.dina(n6034), .dinb(asqrt[41] ), .dout(n6035));
  jor  g05806(.dina(n6034), .dinb(asqrt[41] ), .dout(n6036));
  jxor g05807(.dina(n5651), .dinb(n3955), .dout(n6037));
  jand g05808(.dina(n6037), .dinb(asqrt[34] ), .dout(n6038));
  jxor g05809(.dina(n6038), .dinb(n5656), .dout(n6039));
  jand g05810(.dina(n6039), .dinb(n6036), .dout(n6040));
  jor  g05811(.dina(n6040), .dinb(n6035), .dout(n6041));
  jand g05812(.dina(n6041), .dinb(asqrt[42] ), .dout(n6042));
  jor  g05813(.dina(n6041), .dinb(asqrt[42] ), .dout(n6043));
  jxor g05814(.dina(n5659), .dinb(n3642), .dout(n6044));
  jand g05815(.dina(n6044), .dinb(asqrt[34] ), .dout(n6045));
  jxor g05816(.dina(n6045), .dinb(n5664), .dout(n6046));
  jnot g05817(.din(n6046), .dout(n6047));
  jand g05818(.dina(n6047), .dinb(n6043), .dout(n6048));
  jor  g05819(.dina(n6048), .dinb(n6042), .dout(n6049));
  jand g05820(.dina(n6049), .dinb(asqrt[43] ), .dout(n6050));
  jor  g05821(.dina(n6049), .dinb(asqrt[43] ), .dout(n6051));
  jxor g05822(.dina(n5666), .dinb(n3368), .dout(n6052));
  jand g05823(.dina(n6052), .dinb(asqrt[34] ), .dout(n6053));
  jxor g05824(.dina(n6053), .dinb(n5671), .dout(n6054));
  jand g05825(.dina(n6054), .dinb(n6051), .dout(n6055));
  jor  g05826(.dina(n6055), .dinb(n6050), .dout(n6056));
  jand g05827(.dina(n6056), .dinb(asqrt[44] ), .dout(n6057));
  jor  g05828(.dina(n6056), .dinb(asqrt[44] ), .dout(n6058));
  jxor g05829(.dina(n5674), .dinb(n3089), .dout(n6059));
  jand g05830(.dina(n6059), .dinb(asqrt[34] ), .dout(n6060));
  jxor g05831(.dina(n6060), .dinb(n5679), .dout(n6061));
  jand g05832(.dina(n6061), .dinb(n6058), .dout(n6062));
  jor  g05833(.dina(n6062), .dinb(n6057), .dout(n6063));
  jand g05834(.dina(n6063), .dinb(asqrt[45] ), .dout(n6064));
  jor  g05835(.dina(n6063), .dinb(asqrt[45] ), .dout(n6065));
  jxor g05836(.dina(n5682), .dinb(n2833), .dout(n6066));
  jand g05837(.dina(n6066), .dinb(asqrt[34] ), .dout(n6067));
  jxor g05838(.dina(n6067), .dinb(n5687), .dout(n6068));
  jand g05839(.dina(n6068), .dinb(n6065), .dout(n6069));
  jor  g05840(.dina(n6069), .dinb(n6064), .dout(n6070));
  jand g05841(.dina(n6070), .dinb(asqrt[46] ), .dout(n6071));
  jor  g05842(.dina(n6070), .dinb(asqrt[46] ), .dout(n6072));
  jxor g05843(.dina(n5690), .dinb(n2572), .dout(n6073));
  jand g05844(.dina(n6073), .dinb(asqrt[34] ), .dout(n6074));
  jxor g05845(.dina(n6074), .dinb(n5695), .dout(n6075));
  jnot g05846(.din(n6075), .dout(n6076));
  jand g05847(.dina(n6076), .dinb(n6072), .dout(n6077));
  jor  g05848(.dina(n6077), .dinb(n6071), .dout(n6078));
  jand g05849(.dina(n6078), .dinb(asqrt[47] ), .dout(n6079));
  jor  g05850(.dina(n6078), .dinb(asqrt[47] ), .dout(n6080));
  jxor g05851(.dina(n5697), .dinb(n2345), .dout(n6081));
  jand g05852(.dina(n6081), .dinb(asqrt[34] ), .dout(n6082));
  jxor g05853(.dina(n6082), .dinb(n5702), .dout(n6083));
  jnot g05854(.din(n6083), .dout(n6084));
  jand g05855(.dina(n6084), .dinb(n6080), .dout(n6085));
  jor  g05856(.dina(n6085), .dinb(n6079), .dout(n6086));
  jand g05857(.dina(n6086), .dinb(asqrt[48] ), .dout(n6087));
  jor  g05858(.dina(n6086), .dinb(asqrt[48] ), .dout(n6088));
  jxor g05859(.dina(n5704), .dinb(n2108), .dout(n6089));
  jand g05860(.dina(n6089), .dinb(asqrt[34] ), .dout(n6090));
  jxor g05861(.dina(n6090), .dinb(n5709), .dout(n6091));
  jnot g05862(.din(n6091), .dout(n6092));
  jand g05863(.dina(n6092), .dinb(n6088), .dout(n6093));
  jor  g05864(.dina(n6093), .dinb(n6087), .dout(n6094));
  jand g05865(.dina(n6094), .dinb(asqrt[49] ), .dout(n6095));
  jor  g05866(.dina(n6094), .dinb(asqrt[49] ), .dout(n6096));
  jxor g05867(.dina(n5711), .dinb(n1912), .dout(n6097));
  jand g05868(.dina(n6097), .dinb(asqrt[34] ), .dout(n6098));
  jxor g05869(.dina(n6098), .dinb(n5716), .dout(n6099));
  jand g05870(.dina(n6099), .dinb(n6096), .dout(n6100));
  jor  g05871(.dina(n6100), .dinb(n6095), .dout(n6101));
  jand g05872(.dina(n6101), .dinb(asqrt[50] ), .dout(n6102));
  jor  g05873(.dina(n6101), .dinb(asqrt[50] ), .dout(n6103));
  jxor g05874(.dina(n5719), .dinb(n1699), .dout(n6104));
  jand g05875(.dina(n6104), .dinb(asqrt[34] ), .dout(n6105));
  jxor g05876(.dina(n6105), .dinb(n5724), .dout(n6106));
  jnot g05877(.din(n6106), .dout(n6107));
  jand g05878(.dina(n6107), .dinb(n6103), .dout(n6108));
  jor  g05879(.dina(n6108), .dinb(n6102), .dout(n6109));
  jand g05880(.dina(n6109), .dinb(asqrt[51] ), .dout(n6110));
  jor  g05881(.dina(n6109), .dinb(asqrt[51] ), .dout(n6111));
  jxor g05882(.dina(n5726), .dinb(n1516), .dout(n6112));
  jand g05883(.dina(n6112), .dinb(asqrt[34] ), .dout(n6113));
  jxor g05884(.dina(n6113), .dinb(n5731), .dout(n6114));
  jand g05885(.dina(n6114), .dinb(n6111), .dout(n6115));
  jor  g05886(.dina(n6115), .dinb(n6110), .dout(n6116));
  jand g05887(.dina(n6116), .dinb(asqrt[52] ), .dout(n6117));
  jor  g05888(.dina(n6116), .dinb(asqrt[52] ), .dout(n6118));
  jxor g05889(.dina(n5734), .dinb(n1332), .dout(n6119));
  jand g05890(.dina(n6119), .dinb(asqrt[34] ), .dout(n6120));
  jxor g05891(.dina(n6120), .dinb(n5739), .dout(n6121));
  jnot g05892(.din(n6121), .dout(n6122));
  jand g05893(.dina(n6122), .dinb(n6118), .dout(n6123));
  jor  g05894(.dina(n6123), .dinb(n6117), .dout(n6124));
  jand g05895(.dina(n6124), .dinb(asqrt[53] ), .dout(n6125));
  jor  g05896(.dina(n6124), .dinb(asqrt[53] ), .dout(n6126));
  jxor g05897(.dina(n5741), .dinb(n1173), .dout(n6127));
  jand g05898(.dina(n6127), .dinb(asqrt[34] ), .dout(n6128));
  jxor g05899(.dina(n6128), .dinb(n5746), .dout(n6129));
  jand g05900(.dina(n6129), .dinb(n6126), .dout(n6130));
  jor  g05901(.dina(n6130), .dinb(n6125), .dout(n6131));
  jand g05902(.dina(n6131), .dinb(asqrt[54] ), .dout(n6132));
  jor  g05903(.dina(n6131), .dinb(asqrt[54] ), .dout(n6133));
  jxor g05904(.dina(n5749), .dinb(n1008), .dout(n6134));
  jand g05905(.dina(n6134), .dinb(asqrt[34] ), .dout(n6135));
  jxor g05906(.dina(n6135), .dinb(n5754), .dout(n6136));
  jand g05907(.dina(n6136), .dinb(n6133), .dout(n6137));
  jor  g05908(.dina(n6137), .dinb(n6132), .dout(n6138));
  jand g05909(.dina(n6138), .dinb(asqrt[55] ), .dout(n6139));
  jor  g05910(.dina(n6138), .dinb(asqrt[55] ), .dout(n6140));
  jxor g05911(.dina(n5757), .dinb(n884), .dout(n6141));
  jand g05912(.dina(n6141), .dinb(asqrt[34] ), .dout(n6142));
  jxor g05913(.dina(n6142), .dinb(n5762), .dout(n6143));
  jnot g05914(.din(n6143), .dout(n6144));
  jand g05915(.dina(n6144), .dinb(n6140), .dout(n6145));
  jor  g05916(.dina(n6145), .dinb(n6139), .dout(n6146));
  jand g05917(.dina(n6146), .dinb(asqrt[56] ), .dout(n6147));
  jor  g05918(.dina(n6146), .dinb(asqrt[56] ), .dout(n6148));
  jxor g05919(.dina(n5764), .dinb(n743), .dout(n6149));
  jand g05920(.dina(n6149), .dinb(asqrt[34] ), .dout(n6150));
  jxor g05921(.dina(n6150), .dinb(n5769), .dout(n6151));
  jnot g05922(.din(n6151), .dout(n6152));
  jand g05923(.dina(n6152), .dinb(n6148), .dout(n6153));
  jor  g05924(.dina(n6153), .dinb(n6147), .dout(n6154));
  jand g05925(.dina(n6154), .dinb(asqrt[57] ), .dout(n6155));
  jor  g05926(.dina(n6154), .dinb(asqrt[57] ), .dout(n6156));
  jxor g05927(.dina(n5771), .dinb(n635), .dout(n6157));
  jand g05928(.dina(n6157), .dinb(asqrt[34] ), .dout(n6158));
  jxor g05929(.dina(n6158), .dinb(n5776), .dout(n6159));
  jand g05930(.dina(n6159), .dinb(n6156), .dout(n6160));
  jor  g05931(.dina(n6160), .dinb(n6155), .dout(n6161));
  jand g05932(.dina(n6161), .dinb(asqrt[58] ), .dout(n6162));
  jor  g05933(.dina(n6161), .dinb(asqrt[58] ), .dout(n6163));
  jxor g05934(.dina(n5779), .dinb(n515), .dout(n6164));
  jand g05935(.dina(n6164), .dinb(asqrt[34] ), .dout(n6165));
  jxor g05936(.dina(n6165), .dinb(n5784), .dout(n6166));
  jnot g05937(.din(n6166), .dout(n6167));
  jand g05938(.dina(n6167), .dinb(n6163), .dout(n6168));
  jor  g05939(.dina(n6168), .dinb(n6162), .dout(n6169));
  jand g05940(.dina(n6169), .dinb(asqrt[59] ), .dout(n6170));
  jor  g05941(.dina(n6169), .dinb(asqrt[59] ), .dout(n6171));
  jxor g05942(.dina(n5786), .dinb(n443), .dout(n6172));
  jand g05943(.dina(n6172), .dinb(asqrt[34] ), .dout(n6173));
  jxor g05944(.dina(n6173), .dinb(n5791), .dout(n6174));
  jand g05945(.dina(n6174), .dinb(n6171), .dout(n6175));
  jor  g05946(.dina(n6175), .dinb(n6170), .dout(n6176));
  jand g05947(.dina(n6176), .dinb(asqrt[60] ), .dout(n6177));
  jor  g05948(.dina(n6176), .dinb(asqrt[60] ), .dout(n6178));
  jxor g05949(.dina(n5794), .dinb(n352), .dout(n6179));
  jand g05950(.dina(n6179), .dinb(asqrt[34] ), .dout(n6180));
  jxor g05951(.dina(n6180), .dinb(n5799), .dout(n6181));
  jnot g05952(.din(n6181), .dout(n6182));
  jand g05953(.dina(n6182), .dinb(n6178), .dout(n6183));
  jor  g05954(.dina(n6183), .dinb(n6177), .dout(n6184));
  jand g05955(.dina(n6184), .dinb(asqrt[61] ), .dout(n6185));
  jor  g05956(.dina(n6184), .dinb(asqrt[61] ), .dout(n6186));
  jxor g05957(.dina(n5801), .dinb(n294), .dout(n6187));
  jand g05958(.dina(n6187), .dinb(asqrt[34] ), .dout(n6188));
  jxor g05959(.dina(n6188), .dinb(n5806), .dout(n6189));
  jnot g05960(.din(n6189), .dout(n6190));
  jand g05961(.dina(n6190), .dinb(n6186), .dout(n6191));
  jor  g05962(.dina(n6191), .dinb(n6185), .dout(n6192));
  jand g05963(.dina(n6192), .dinb(asqrt[62] ), .dout(n6193));
  jor  g05964(.dina(n6192), .dinb(asqrt[62] ), .dout(n6194));
  jxor g05965(.dina(n5808), .dinb(n239), .dout(n6195));
  jand g05966(.dina(n6195), .dinb(asqrt[34] ), .dout(n6196));
  jxor g05967(.dina(n6196), .dinb(n5813), .dout(n6197));
  jnot g05968(.din(n6197), .dout(n6198));
  jand g05969(.dina(n6198), .dinb(n6194), .dout(n6199));
  jor  g05970(.dina(n6199), .dinb(n6193), .dout(n6200));
  jor  g05971(.dina(n6200), .dinb(n5842), .dout(n6201));
  jnot g05972(.din(n6201), .dout(n6202));
  jnot g05973(.din(n5842), .dout(n6204));
  jnot g05974(.din(n6193), .dout(n6205));
  jnot g05975(.din(n6185), .dout(n6206));
  jnot g05976(.din(n6177), .dout(n6207));
  jnot g05977(.din(n6170), .dout(n6208));
  jnot g05978(.din(n6162), .dout(n6209));
  jnot g05979(.din(n6155), .dout(n6210));
  jnot g05980(.din(n6147), .dout(n6211));
  jnot g05981(.din(n6139), .dout(n6212));
  jnot g05982(.din(n6132), .dout(n6213));
  jnot g05983(.din(n6125), .dout(n6214));
  jnot g05984(.din(n6117), .dout(n6215));
  jnot g05985(.din(n6110), .dout(n6216));
  jnot g05986(.din(n6102), .dout(n6217));
  jnot g05987(.din(n6095), .dout(n6218));
  jnot g05988(.din(n6087), .dout(n6219));
  jnot g05989(.din(n6079), .dout(n6220));
  jnot g05990(.din(n6071), .dout(n6221));
  jnot g05991(.din(n6064), .dout(n6222));
  jnot g05992(.din(n6057), .dout(n6223));
  jnot g05993(.din(n6050), .dout(n6224));
  jnot g05994(.din(n6042), .dout(n6225));
  jnot g05995(.din(n6035), .dout(n6226));
  jnot g05996(.din(n6027), .dout(n6227));
  jnot g05997(.din(n6020), .dout(n6228));
  jnot g05998(.din(n6012), .dout(n6229));
  jnot g05999(.din(n6005), .dout(n6230));
  jnot g06000(.din(n5994), .dout(n6231));
  jnot g06001(.din(n5849), .dout(n6232));
  jnot g06002(.din(n5846), .dout(n6233));
  jor  g06003(.dina(n5989), .dinb(n5612), .dout(n6234));
  jand g06004(.dina(n6234), .dinb(n6233), .dout(n6235));
  jand g06005(.dina(n6235), .dinb(n5606), .dout(n6236));
  jor  g06006(.dina(n5989), .dinb(a[68] ), .dout(n6237));
  jand g06007(.dina(n6237), .dinb(a[69] ), .dout(n6238));
  jor  g06008(.dina(n5996), .dinb(n6238), .dout(n6239));
  jor  g06009(.dina(n6239), .dinb(n6236), .dout(n6240));
  jand g06010(.dina(n6240), .dinb(n6232), .dout(n6241));
  jand g06011(.dina(n6241), .dinb(n5259), .dout(n6242));
  jor  g06012(.dina(n6001), .dinb(n6242), .dout(n6243));
  jand g06013(.dina(n6243), .dinb(n6231), .dout(n6244));
  jand g06014(.dina(n6244), .dinb(n4902), .dout(n6245));
  jnot g06015(.din(n6009), .dout(n6246));
  jor  g06016(.dina(n6246), .dinb(n6245), .dout(n6247));
  jand g06017(.dina(n6247), .dinb(n6230), .dout(n6248));
  jand g06018(.dina(n6248), .dinb(n4582), .dout(n6249));
  jor  g06019(.dina(n6016), .dinb(n6249), .dout(n6250));
  jand g06020(.dina(n6250), .dinb(n6229), .dout(n6251));
  jand g06021(.dina(n6251), .dinb(n4249), .dout(n6252));
  jnot g06022(.din(n6024), .dout(n6253));
  jor  g06023(.dina(n6253), .dinb(n6252), .dout(n6254));
  jand g06024(.dina(n6254), .dinb(n6228), .dout(n6255));
  jand g06025(.dina(n6255), .dinb(n3955), .dout(n6256));
  jor  g06026(.dina(n6031), .dinb(n6256), .dout(n6257));
  jand g06027(.dina(n6257), .dinb(n6227), .dout(n6258));
  jand g06028(.dina(n6258), .dinb(n3642), .dout(n6259));
  jnot g06029(.din(n6039), .dout(n6260));
  jor  g06030(.dina(n6260), .dinb(n6259), .dout(n6261));
  jand g06031(.dina(n6261), .dinb(n6226), .dout(n6262));
  jand g06032(.dina(n6262), .dinb(n3368), .dout(n6263));
  jor  g06033(.dina(n6046), .dinb(n6263), .dout(n6264));
  jand g06034(.dina(n6264), .dinb(n6225), .dout(n6265));
  jand g06035(.dina(n6265), .dinb(n3089), .dout(n6266));
  jnot g06036(.din(n6054), .dout(n6267));
  jor  g06037(.dina(n6267), .dinb(n6266), .dout(n6268));
  jand g06038(.dina(n6268), .dinb(n6224), .dout(n6269));
  jand g06039(.dina(n6269), .dinb(n2833), .dout(n6270));
  jnot g06040(.din(n6061), .dout(n6271));
  jor  g06041(.dina(n6271), .dinb(n6270), .dout(n6272));
  jand g06042(.dina(n6272), .dinb(n6223), .dout(n6273));
  jand g06043(.dina(n6273), .dinb(n2572), .dout(n6274));
  jnot g06044(.din(n6068), .dout(n6275));
  jor  g06045(.dina(n6275), .dinb(n6274), .dout(n6276));
  jand g06046(.dina(n6276), .dinb(n6222), .dout(n6277));
  jand g06047(.dina(n6277), .dinb(n2345), .dout(n6278));
  jor  g06048(.dina(n6075), .dinb(n6278), .dout(n6279));
  jand g06049(.dina(n6279), .dinb(n6221), .dout(n6280));
  jand g06050(.dina(n6280), .dinb(n2108), .dout(n6281));
  jor  g06051(.dina(n6083), .dinb(n6281), .dout(n6282));
  jand g06052(.dina(n6282), .dinb(n6220), .dout(n6283));
  jand g06053(.dina(n6283), .dinb(n1912), .dout(n6284));
  jor  g06054(.dina(n6091), .dinb(n6284), .dout(n6285));
  jand g06055(.dina(n6285), .dinb(n6219), .dout(n6286));
  jand g06056(.dina(n6286), .dinb(n1699), .dout(n6287));
  jnot g06057(.din(n6099), .dout(n6288));
  jor  g06058(.dina(n6288), .dinb(n6287), .dout(n6289));
  jand g06059(.dina(n6289), .dinb(n6218), .dout(n6290));
  jand g06060(.dina(n6290), .dinb(n1516), .dout(n6291));
  jor  g06061(.dina(n6106), .dinb(n6291), .dout(n6292));
  jand g06062(.dina(n6292), .dinb(n6217), .dout(n6293));
  jand g06063(.dina(n6293), .dinb(n1332), .dout(n6294));
  jnot g06064(.din(n6114), .dout(n6295));
  jor  g06065(.dina(n6295), .dinb(n6294), .dout(n6296));
  jand g06066(.dina(n6296), .dinb(n6216), .dout(n6297));
  jand g06067(.dina(n6297), .dinb(n1173), .dout(n6298));
  jor  g06068(.dina(n6121), .dinb(n6298), .dout(n6299));
  jand g06069(.dina(n6299), .dinb(n6215), .dout(n6300));
  jand g06070(.dina(n6300), .dinb(n1008), .dout(n6301));
  jnot g06071(.din(n6129), .dout(n6302));
  jor  g06072(.dina(n6302), .dinb(n6301), .dout(n6303));
  jand g06073(.dina(n6303), .dinb(n6214), .dout(n6304));
  jand g06074(.dina(n6304), .dinb(n884), .dout(n6305));
  jnot g06075(.din(n6136), .dout(n6306));
  jor  g06076(.dina(n6306), .dinb(n6305), .dout(n6307));
  jand g06077(.dina(n6307), .dinb(n6213), .dout(n6308));
  jand g06078(.dina(n6308), .dinb(n743), .dout(n6309));
  jor  g06079(.dina(n6143), .dinb(n6309), .dout(n6310));
  jand g06080(.dina(n6310), .dinb(n6212), .dout(n6311));
  jand g06081(.dina(n6311), .dinb(n635), .dout(n6312));
  jor  g06082(.dina(n6151), .dinb(n6312), .dout(n6313));
  jand g06083(.dina(n6313), .dinb(n6211), .dout(n6314));
  jand g06084(.dina(n6314), .dinb(n515), .dout(n6315));
  jnot g06085(.din(n6159), .dout(n6316));
  jor  g06086(.dina(n6316), .dinb(n6315), .dout(n6317));
  jand g06087(.dina(n6317), .dinb(n6210), .dout(n6318));
  jand g06088(.dina(n6318), .dinb(n443), .dout(n6319));
  jor  g06089(.dina(n6166), .dinb(n6319), .dout(n6320));
  jand g06090(.dina(n6320), .dinb(n6209), .dout(n6321));
  jand g06091(.dina(n6321), .dinb(n352), .dout(n6322));
  jnot g06092(.din(n6174), .dout(n6323));
  jor  g06093(.dina(n6323), .dinb(n6322), .dout(n6324));
  jand g06094(.dina(n6324), .dinb(n6208), .dout(n6325));
  jand g06095(.dina(n6325), .dinb(n294), .dout(n6326));
  jor  g06096(.dina(n6181), .dinb(n6326), .dout(n6327));
  jand g06097(.dina(n6327), .dinb(n6207), .dout(n6328));
  jand g06098(.dina(n6328), .dinb(n239), .dout(n6329));
  jor  g06099(.dina(n6189), .dinb(n6329), .dout(n6330));
  jand g06100(.dina(n6330), .dinb(n6206), .dout(n6331));
  jand g06101(.dina(n6331), .dinb(n221), .dout(n6332));
  jor  g06102(.dina(n6197), .dinb(n6332), .dout(n6333));
  jand g06103(.dina(n6333), .dinb(n6205), .dout(n6334));
  jor  g06104(.dina(n6334), .dinb(n6204), .dout(n6335));
  jxor g06105(.dina(n5823), .dinb(n5610), .dout(n6336));
  jnot g06106(.din(n6336), .dout(n6337));
  jand g06107(.dina(n6337), .dinb(asqrt[34] ), .dout(n6338));
  jor  g06108(.dina(n6338), .dinb(n6335), .dout(n6339));
  jand g06109(.dina(n6339), .dinb(n218), .dout(n6340));
  jand g06110(.dina(n5987), .dinb(n5823), .dout(n6341));
  jnot g06111(.din(n6341), .dout(n6342));
  jand g06112(.dina(n6336), .dinb(asqrt[63] ), .dout(n6343));
  jand g06113(.dina(n6343), .dinb(n6342), .dout(n6344));
  jor  g06114(.dina(n6344), .dinb(n6340), .dout(n6345));
  jor  g06115(.dina(n6345), .dinb(n6202), .dout(asqrt[33] ));
  jand g06116(.dina(n6200), .dinb(n5842), .dout(n6348));
  jand g06117(.dina(n6345), .dinb(n6348), .dout(n6349));
  jnot g06118(.din(n6338), .dout(n6351));
  jand g06119(.dina(n6351), .dinb(n6348), .dout(n6352));
  jor  g06120(.dina(n6352), .dinb(asqrt[63] ), .dout(n6353));
  jnot g06121(.din(n6344), .dout(n6354));
  jand g06122(.dina(n6354), .dinb(n6353), .dout(n6355));
  jand g06123(.dina(n6355), .dinb(n6201), .dout(n6357));
  jxor g06124(.dina(n6192), .dinb(n221), .dout(n6358));
  jor  g06125(.dina(n6358), .dinb(n6357), .dout(n6359));
  jxor g06126(.dina(n6359), .dinb(n6197), .dout(n6360));
  jnot g06127(.din(n6360), .dout(n6361));
  jnot g06128(.din(a[64] ), .dout(n6362));
  jnot g06129(.din(a[65] ), .dout(n6363));
  jand g06130(.dina(n6363), .dinb(n6362), .dout(n6364));
  jand g06131(.dina(n6364), .dinb(n5843), .dout(n6365));
  jnot g06132(.din(n6365), .dout(n6366));
  jor  g06133(.dina(n6357), .dinb(n5843), .dout(n6367));
  jand g06134(.dina(n6367), .dinb(n6366), .dout(n6368));
  jor  g06135(.dina(n6368), .dinb(n5989), .dout(n6369));
  jand g06136(.dina(n6368), .dinb(n5989), .dout(n6370));
  jor  g06137(.dina(n6357), .dinb(a[66] ), .dout(n6371));
  jand g06138(.dina(n6371), .dinb(a[67] ), .dout(n6372));
  jand g06139(.dina(asqrt[33] ), .dinb(n5845), .dout(n6373));
  jor  g06140(.dina(n6373), .dinb(n6372), .dout(n6374));
  jor  g06141(.dina(n6374), .dinb(n6370), .dout(n6375));
  jand g06142(.dina(n6375), .dinb(n6369), .dout(n6376));
  jor  g06143(.dina(n6376), .dinb(n5606), .dout(n6377));
  jand g06144(.dina(n6376), .dinb(n5606), .dout(n6378));
  jnot g06145(.din(n5845), .dout(n6379));
  jor  g06146(.dina(n6357), .dinb(n6379), .dout(n6380));
  jor  g06147(.dina(n6343), .dinb(n6202), .dout(n6381));
  jor  g06148(.dina(n6381), .dinb(n6340), .dout(n6382));
  jor  g06149(.dina(n6382), .dinb(n5989), .dout(n6383));
  jand g06150(.dina(n6383), .dinb(n6380), .dout(n6384));
  jxor g06151(.dina(n6384), .dinb(n5612), .dout(n6385));
  jor  g06152(.dina(n6385), .dinb(n6378), .dout(n6386));
  jand g06153(.dina(n6386), .dinb(n6377), .dout(n6387));
  jor  g06154(.dina(n6387), .dinb(n5259), .dout(n6388));
  jand g06155(.dina(n6387), .dinb(n5259), .dout(n6389));
  jxor g06156(.dina(n5848), .dinb(n5606), .dout(n6390));
  jor  g06157(.dina(n6390), .dinb(n6357), .dout(n6391));
  jxor g06158(.dina(n6391), .dinb(n6239), .dout(n6392));
  jnot g06159(.din(n6392), .dout(n6393));
  jor  g06160(.dina(n6393), .dinb(n6389), .dout(n6394));
  jand g06161(.dina(n6394), .dinb(n6388), .dout(n6395));
  jor  g06162(.dina(n6395), .dinb(n4902), .dout(n6396));
  jand g06163(.dina(n6395), .dinb(n4902), .dout(n6397));
  jxor g06164(.dina(n5993), .dinb(n5259), .dout(n6398));
  jor  g06165(.dina(n6398), .dinb(n6357), .dout(n6399));
  jxor g06166(.dina(n6399), .dinb(n6002), .dout(n6400));
  jor  g06167(.dina(n6400), .dinb(n6397), .dout(n6401));
  jand g06168(.dina(n6401), .dinb(n6396), .dout(n6402));
  jor  g06169(.dina(n6402), .dinb(n4582), .dout(n6403));
  jand g06170(.dina(n6402), .dinb(n4582), .dout(n6404));
  jxor g06171(.dina(n6004), .dinb(n4902), .dout(n6405));
  jor  g06172(.dina(n6405), .dinb(n6357), .dout(n6406));
  jxor g06173(.dina(n6406), .dinb(n6246), .dout(n6407));
  jnot g06174(.din(n6407), .dout(n6408));
  jor  g06175(.dina(n6408), .dinb(n6404), .dout(n6409));
  jand g06176(.dina(n6409), .dinb(n6403), .dout(n6410));
  jor  g06177(.dina(n6410), .dinb(n4249), .dout(n6411));
  jand g06178(.dina(n6410), .dinb(n4249), .dout(n6412));
  jxor g06179(.dina(n6011), .dinb(n4582), .dout(n6413));
  jor  g06180(.dina(n6413), .dinb(n6357), .dout(n6414));
  jxor g06181(.dina(n6414), .dinb(n6017), .dout(n6415));
  jor  g06182(.dina(n6415), .dinb(n6412), .dout(n6416));
  jand g06183(.dina(n6416), .dinb(n6411), .dout(n6417));
  jor  g06184(.dina(n6417), .dinb(n3955), .dout(n6418));
  jand g06185(.dina(n6417), .dinb(n3955), .dout(n6419));
  jxor g06186(.dina(n6019), .dinb(n4249), .dout(n6420));
  jor  g06187(.dina(n6420), .dinb(n6357), .dout(n6421));
  jxor g06188(.dina(n6421), .dinb(n6253), .dout(n6422));
  jnot g06189(.din(n6422), .dout(n6423));
  jor  g06190(.dina(n6423), .dinb(n6419), .dout(n6424));
  jand g06191(.dina(n6424), .dinb(n6418), .dout(n6425));
  jor  g06192(.dina(n6425), .dinb(n3642), .dout(n6426));
  jand g06193(.dina(n6425), .dinb(n3642), .dout(n6427));
  jxor g06194(.dina(n6026), .dinb(n3955), .dout(n6428));
  jor  g06195(.dina(n6428), .dinb(n6357), .dout(n6429));
  jxor g06196(.dina(n6429), .dinb(n6032), .dout(n6430));
  jor  g06197(.dina(n6430), .dinb(n6427), .dout(n6431));
  jand g06198(.dina(n6431), .dinb(n6426), .dout(n6432));
  jor  g06199(.dina(n6432), .dinb(n3368), .dout(n6433));
  jand g06200(.dina(n6432), .dinb(n3368), .dout(n6434));
  jxor g06201(.dina(n6034), .dinb(n3642), .dout(n6435));
  jor  g06202(.dina(n6435), .dinb(n6357), .dout(n6436));
  jxor g06203(.dina(n6436), .dinb(n6260), .dout(n6437));
  jnot g06204(.din(n6437), .dout(n6438));
  jor  g06205(.dina(n6438), .dinb(n6434), .dout(n6439));
  jand g06206(.dina(n6439), .dinb(n6433), .dout(n6440));
  jor  g06207(.dina(n6440), .dinb(n3089), .dout(n6441));
  jand g06208(.dina(n6440), .dinb(n3089), .dout(n6442));
  jxor g06209(.dina(n6041), .dinb(n3368), .dout(n6443));
  jor  g06210(.dina(n6443), .dinb(n6357), .dout(n6444));
  jxor g06211(.dina(n6444), .dinb(n6047), .dout(n6445));
  jor  g06212(.dina(n6445), .dinb(n6442), .dout(n6446));
  jand g06213(.dina(n6446), .dinb(n6441), .dout(n6447));
  jor  g06214(.dina(n6447), .dinb(n2833), .dout(n6448));
  jand g06215(.dina(n6447), .dinb(n2833), .dout(n6449));
  jxor g06216(.dina(n6049), .dinb(n3089), .dout(n6450));
  jor  g06217(.dina(n6450), .dinb(n6357), .dout(n6451));
  jxor g06218(.dina(n6451), .dinb(n6267), .dout(n6452));
  jnot g06219(.din(n6452), .dout(n6453));
  jor  g06220(.dina(n6453), .dinb(n6449), .dout(n6454));
  jand g06221(.dina(n6454), .dinb(n6448), .dout(n6455));
  jor  g06222(.dina(n6455), .dinb(n2572), .dout(n6456));
  jand g06223(.dina(n6455), .dinb(n2572), .dout(n6457));
  jxor g06224(.dina(n6056), .dinb(n2833), .dout(n6458));
  jor  g06225(.dina(n6458), .dinb(n6357), .dout(n6459));
  jxor g06226(.dina(n6459), .dinb(n6271), .dout(n6460));
  jnot g06227(.din(n6460), .dout(n6461));
  jor  g06228(.dina(n6461), .dinb(n6457), .dout(n6462));
  jand g06229(.dina(n6462), .dinb(n6456), .dout(n6463));
  jor  g06230(.dina(n6463), .dinb(n2345), .dout(n6464));
  jand g06231(.dina(n6463), .dinb(n2345), .dout(n6465));
  jxor g06232(.dina(n6063), .dinb(n2572), .dout(n6466));
  jor  g06233(.dina(n6466), .dinb(n6357), .dout(n6467));
  jxor g06234(.dina(n6467), .dinb(n6275), .dout(n6468));
  jnot g06235(.din(n6468), .dout(n6469));
  jor  g06236(.dina(n6469), .dinb(n6465), .dout(n6470));
  jand g06237(.dina(n6470), .dinb(n6464), .dout(n6471));
  jor  g06238(.dina(n6471), .dinb(n2108), .dout(n6472));
  jand g06239(.dina(n6471), .dinb(n2108), .dout(n6473));
  jxor g06240(.dina(n6070), .dinb(n2345), .dout(n6474));
  jor  g06241(.dina(n6474), .dinb(n6357), .dout(n6475));
  jxor g06242(.dina(n6475), .dinb(n6076), .dout(n6476));
  jor  g06243(.dina(n6476), .dinb(n6473), .dout(n6477));
  jand g06244(.dina(n6477), .dinb(n6472), .dout(n6478));
  jor  g06245(.dina(n6478), .dinb(n1912), .dout(n6479));
  jand g06246(.dina(n6478), .dinb(n1912), .dout(n6480));
  jxor g06247(.dina(n6078), .dinb(n2108), .dout(n6481));
  jor  g06248(.dina(n6481), .dinb(n6357), .dout(n6482));
  jxor g06249(.dina(n6482), .dinb(n6084), .dout(n6483));
  jor  g06250(.dina(n6483), .dinb(n6480), .dout(n6484));
  jand g06251(.dina(n6484), .dinb(n6479), .dout(n6485));
  jor  g06252(.dina(n6485), .dinb(n1699), .dout(n6486));
  jand g06253(.dina(n6485), .dinb(n1699), .dout(n6487));
  jxor g06254(.dina(n6086), .dinb(n1912), .dout(n6488));
  jor  g06255(.dina(n6488), .dinb(n6357), .dout(n6489));
  jxor g06256(.dina(n6489), .dinb(n6092), .dout(n6490));
  jor  g06257(.dina(n6490), .dinb(n6487), .dout(n6491));
  jand g06258(.dina(n6491), .dinb(n6486), .dout(n6492));
  jor  g06259(.dina(n6492), .dinb(n1516), .dout(n6493));
  jand g06260(.dina(n6492), .dinb(n1516), .dout(n6494));
  jxor g06261(.dina(n6094), .dinb(n1699), .dout(n6495));
  jor  g06262(.dina(n6495), .dinb(n6357), .dout(n6496));
  jxor g06263(.dina(n6496), .dinb(n6288), .dout(n6497));
  jnot g06264(.din(n6497), .dout(n6498));
  jor  g06265(.dina(n6498), .dinb(n6494), .dout(n6499));
  jand g06266(.dina(n6499), .dinb(n6493), .dout(n6500));
  jor  g06267(.dina(n6500), .dinb(n1332), .dout(n6501));
  jand g06268(.dina(n6500), .dinb(n1332), .dout(n6502));
  jxor g06269(.dina(n6101), .dinb(n1516), .dout(n6503));
  jor  g06270(.dina(n6503), .dinb(n6357), .dout(n6504));
  jxor g06271(.dina(n6504), .dinb(n6107), .dout(n6505));
  jor  g06272(.dina(n6505), .dinb(n6502), .dout(n6506));
  jand g06273(.dina(n6506), .dinb(n6501), .dout(n6507));
  jor  g06274(.dina(n6507), .dinb(n1173), .dout(n6508));
  jand g06275(.dina(n6507), .dinb(n1173), .dout(n6509));
  jxor g06276(.dina(n6109), .dinb(n1332), .dout(n6510));
  jor  g06277(.dina(n6510), .dinb(n6357), .dout(n6511));
  jxor g06278(.dina(n6511), .dinb(n6295), .dout(n6512));
  jnot g06279(.din(n6512), .dout(n6513));
  jor  g06280(.dina(n6513), .dinb(n6509), .dout(n6514));
  jand g06281(.dina(n6514), .dinb(n6508), .dout(n6515));
  jor  g06282(.dina(n6515), .dinb(n1008), .dout(n6516));
  jand g06283(.dina(n6515), .dinb(n1008), .dout(n6517));
  jxor g06284(.dina(n6116), .dinb(n1173), .dout(n6518));
  jor  g06285(.dina(n6518), .dinb(n6357), .dout(n6519));
  jxor g06286(.dina(n6519), .dinb(n6122), .dout(n6520));
  jor  g06287(.dina(n6520), .dinb(n6517), .dout(n6521));
  jand g06288(.dina(n6521), .dinb(n6516), .dout(n6522));
  jor  g06289(.dina(n6522), .dinb(n884), .dout(n6523));
  jand g06290(.dina(n6522), .dinb(n884), .dout(n6524));
  jxor g06291(.dina(n6124), .dinb(n1008), .dout(n6525));
  jor  g06292(.dina(n6525), .dinb(n6357), .dout(n6526));
  jxor g06293(.dina(n6526), .dinb(n6302), .dout(n6527));
  jnot g06294(.din(n6527), .dout(n6528));
  jor  g06295(.dina(n6528), .dinb(n6524), .dout(n6529));
  jand g06296(.dina(n6529), .dinb(n6523), .dout(n6530));
  jor  g06297(.dina(n6530), .dinb(n743), .dout(n6531));
  jand g06298(.dina(n6530), .dinb(n743), .dout(n6532));
  jxor g06299(.dina(n6131), .dinb(n884), .dout(n6533));
  jor  g06300(.dina(n6533), .dinb(n6357), .dout(n6534));
  jxor g06301(.dina(n6534), .dinb(n6306), .dout(n6535));
  jnot g06302(.din(n6535), .dout(n6536));
  jor  g06303(.dina(n6536), .dinb(n6532), .dout(n6537));
  jand g06304(.dina(n6537), .dinb(n6531), .dout(n6538));
  jor  g06305(.dina(n6538), .dinb(n635), .dout(n6539));
  jand g06306(.dina(n6538), .dinb(n635), .dout(n6540));
  jxor g06307(.dina(n6138), .dinb(n743), .dout(n6541));
  jor  g06308(.dina(n6541), .dinb(n6357), .dout(n6542));
  jxor g06309(.dina(n6542), .dinb(n6144), .dout(n6543));
  jor  g06310(.dina(n6543), .dinb(n6540), .dout(n6544));
  jand g06311(.dina(n6544), .dinb(n6539), .dout(n6545));
  jor  g06312(.dina(n6545), .dinb(n515), .dout(n6546));
  jand g06313(.dina(n6545), .dinb(n515), .dout(n6547));
  jxor g06314(.dina(n6146), .dinb(n635), .dout(n6548));
  jor  g06315(.dina(n6548), .dinb(n6357), .dout(n6549));
  jxor g06316(.dina(n6549), .dinb(n6152), .dout(n6550));
  jor  g06317(.dina(n6550), .dinb(n6547), .dout(n6551));
  jand g06318(.dina(n6551), .dinb(n6546), .dout(n6552));
  jor  g06319(.dina(n6552), .dinb(n443), .dout(n6553));
  jand g06320(.dina(n6552), .dinb(n443), .dout(n6554));
  jxor g06321(.dina(n6154), .dinb(n515), .dout(n6555));
  jor  g06322(.dina(n6555), .dinb(n6357), .dout(n6556));
  jxor g06323(.dina(n6556), .dinb(n6316), .dout(n6557));
  jnot g06324(.din(n6557), .dout(n6558));
  jor  g06325(.dina(n6558), .dinb(n6554), .dout(n6559));
  jand g06326(.dina(n6559), .dinb(n6553), .dout(n6560));
  jor  g06327(.dina(n6560), .dinb(n352), .dout(n6561));
  jand g06328(.dina(n6560), .dinb(n352), .dout(n6562));
  jxor g06329(.dina(n6161), .dinb(n443), .dout(n6563));
  jor  g06330(.dina(n6563), .dinb(n6357), .dout(n6564));
  jxor g06331(.dina(n6564), .dinb(n6166), .dout(n6565));
  jnot g06332(.din(n6565), .dout(n6566));
  jor  g06333(.dina(n6566), .dinb(n6562), .dout(n6567));
  jand g06334(.dina(n6567), .dinb(n6561), .dout(n6568));
  jor  g06335(.dina(n6568), .dinb(n294), .dout(n6569));
  jand g06336(.dina(n6568), .dinb(n294), .dout(n6570));
  jxor g06337(.dina(n6169), .dinb(n352), .dout(n6571));
  jor  g06338(.dina(n6571), .dinb(n6357), .dout(n6572));
  jxor g06339(.dina(n6572), .dinb(n6323), .dout(n6573));
  jnot g06340(.din(n6573), .dout(n6574));
  jor  g06341(.dina(n6574), .dinb(n6570), .dout(n6575));
  jand g06342(.dina(n6575), .dinb(n6569), .dout(n6576));
  jor  g06343(.dina(n6576), .dinb(n239), .dout(n6577));
  jand g06344(.dina(n6576), .dinb(n239), .dout(n6578));
  jxor g06345(.dina(n6176), .dinb(n294), .dout(n6579));
  jor  g06346(.dina(n6579), .dinb(n6357), .dout(n6580));
  jxor g06347(.dina(n6580), .dinb(n6182), .dout(n6581));
  jor  g06348(.dina(n6581), .dinb(n6578), .dout(n6582));
  jand g06349(.dina(n6582), .dinb(n6577), .dout(n6583));
  jor  g06350(.dina(n6583), .dinb(n221), .dout(n6584));
  jand g06351(.dina(n6583), .dinb(n221), .dout(n6585));
  jxor g06352(.dina(n6184), .dinb(n239), .dout(n6586));
  jor  g06353(.dina(n6586), .dinb(n6357), .dout(n6587));
  jxor g06354(.dina(n6587), .dinb(n6190), .dout(n6588));
  jor  g06355(.dina(n6588), .dinb(n6585), .dout(n6589));
  jand g06356(.dina(n6589), .dinb(n6584), .dout(n6590));
  jor  g06357(.dina(n6590), .dinb(n6361), .dout(n6591));
  jor  g06358(.dina(n6591), .dinb(n6202), .dout(n6592));
  jor  g06359(.dina(n6592), .dinb(n6349), .dout(n6593));
  jand g06360(.dina(n6593), .dinb(n218), .dout(n6594));
  jand g06361(.dina(n6357), .dinb(n6204), .dout(n6595));
  jand g06362(.dina(n6590), .dinb(n6361), .dout(n6596));
  jor  g06363(.dina(n6596), .dinb(n6595), .dout(n6597));
  jand g06364(.dina(n6355), .dinb(n6334), .dout(n6598));
  jand g06365(.dina(n6335), .dinb(asqrt[63] ), .dout(n6599));
  jand g06366(.dina(n6599), .dinb(n6201), .dout(n6600));
  jnot g06367(.din(n6600), .dout(n6601));
  jor  g06368(.dina(n6601), .dinb(n6598), .dout(n6602));
  jnot g06369(.din(n6602), .dout(n6603));
  jor  g06370(.dina(n6603), .dinb(n6597), .dout(n6604));
  jor  g06371(.dina(n6604), .dinb(n6594), .dout(asqrt[32] ));
  jnot g06372(.din(a[62] ), .dout(n6606));
  jnot g06373(.din(a[63] ), .dout(n6607));
  jand g06374(.dina(n6607), .dinb(n6606), .dout(n6608));
  jand g06375(.dina(n6608), .dinb(n6362), .dout(n6609));
  jand g06376(.dina(asqrt[32] ), .dinb(a[64] ), .dout(n6610));
  jor  g06377(.dina(n6610), .dinb(n6609), .dout(n6611));
  jand g06378(.dina(n6611), .dinb(asqrt[33] ), .dout(n6612));
  jor  g06379(.dina(n6611), .dinb(asqrt[33] ), .dout(n6613));
  jand g06380(.dina(asqrt[32] ), .dinb(n6362), .dout(n6614));
  jor  g06381(.dina(n6614), .dinb(n6363), .dout(n6615));
  jnot g06382(.din(n6364), .dout(n6616));
  jnot g06383(.din(n6349), .dout(n6617));
  jnot g06384(.din(n6584), .dout(n6618));
  jnot g06385(.din(n6577), .dout(n6619));
  jnot g06386(.din(n6569), .dout(n6620));
  jnot g06387(.din(n6561), .dout(n6621));
  jnot g06388(.din(n6553), .dout(n6622));
  jnot g06389(.din(n6546), .dout(n6623));
  jnot g06390(.din(n6539), .dout(n6624));
  jnot g06391(.din(n6531), .dout(n6625));
  jnot g06392(.din(n6523), .dout(n6626));
  jnot g06393(.din(n6516), .dout(n6627));
  jnot g06394(.din(n6508), .dout(n6628));
  jnot g06395(.din(n6501), .dout(n6629));
  jnot g06396(.din(n6493), .dout(n6630));
  jnot g06397(.din(n6486), .dout(n6631));
  jnot g06398(.din(n6479), .dout(n6632));
  jnot g06399(.din(n6472), .dout(n6633));
  jnot g06400(.din(n6464), .dout(n6634));
  jnot g06401(.din(n6456), .dout(n6635));
  jnot g06402(.din(n6448), .dout(n6636));
  jnot g06403(.din(n6441), .dout(n6637));
  jnot g06404(.din(n6433), .dout(n6638));
  jnot g06405(.din(n6426), .dout(n6639));
  jnot g06406(.din(n6418), .dout(n6640));
  jnot g06407(.din(n6411), .dout(n6641));
  jnot g06408(.din(n6403), .dout(n6642));
  jnot g06409(.din(n6396), .dout(n6643));
  jnot g06410(.din(n6388), .dout(n6644));
  jnot g06411(.din(n6377), .dout(n6645));
  jnot g06412(.din(n6369), .dout(n6646));
  jand g06413(.dina(asqrt[33] ), .dinb(a[66] ), .dout(n6647));
  jor  g06414(.dina(n6647), .dinb(n6365), .dout(n6648));
  jor  g06415(.dina(n6648), .dinb(asqrt[34] ), .dout(n6649));
  jand g06416(.dina(asqrt[33] ), .dinb(n5843), .dout(n6650));
  jor  g06417(.dina(n6650), .dinb(n5844), .dout(n6651));
  jand g06418(.dina(n6380), .dinb(n6651), .dout(n6652));
  jand g06419(.dina(n6652), .dinb(n6649), .dout(n6653));
  jor  g06420(.dina(n6653), .dinb(n6646), .dout(n6654));
  jor  g06421(.dina(n6654), .dinb(asqrt[35] ), .dout(n6655));
  jnot g06422(.din(n6385), .dout(n6656));
  jand g06423(.dina(n6656), .dinb(n6655), .dout(n6657));
  jor  g06424(.dina(n6657), .dinb(n6645), .dout(n6658));
  jor  g06425(.dina(n6658), .dinb(asqrt[36] ), .dout(n6659));
  jand g06426(.dina(n6392), .dinb(n6659), .dout(n6660));
  jor  g06427(.dina(n6660), .dinb(n6644), .dout(n6661));
  jor  g06428(.dina(n6661), .dinb(asqrt[37] ), .dout(n6662));
  jnot g06429(.din(n6400), .dout(n6663));
  jand g06430(.dina(n6663), .dinb(n6662), .dout(n6664));
  jor  g06431(.dina(n6664), .dinb(n6643), .dout(n6665));
  jor  g06432(.dina(n6665), .dinb(asqrt[38] ), .dout(n6666));
  jand g06433(.dina(n6407), .dinb(n6666), .dout(n6667));
  jor  g06434(.dina(n6667), .dinb(n6642), .dout(n6668));
  jor  g06435(.dina(n6668), .dinb(asqrt[39] ), .dout(n6669));
  jnot g06436(.din(n6415), .dout(n6670));
  jand g06437(.dina(n6670), .dinb(n6669), .dout(n6671));
  jor  g06438(.dina(n6671), .dinb(n6641), .dout(n6672));
  jor  g06439(.dina(n6672), .dinb(asqrt[40] ), .dout(n6673));
  jand g06440(.dina(n6422), .dinb(n6673), .dout(n6674));
  jor  g06441(.dina(n6674), .dinb(n6640), .dout(n6675));
  jor  g06442(.dina(n6675), .dinb(asqrt[41] ), .dout(n6676));
  jnot g06443(.din(n6430), .dout(n6677));
  jand g06444(.dina(n6677), .dinb(n6676), .dout(n6678));
  jor  g06445(.dina(n6678), .dinb(n6639), .dout(n6679));
  jor  g06446(.dina(n6679), .dinb(asqrt[42] ), .dout(n6680));
  jand g06447(.dina(n6437), .dinb(n6680), .dout(n6681));
  jor  g06448(.dina(n6681), .dinb(n6638), .dout(n6682));
  jor  g06449(.dina(n6682), .dinb(asqrt[43] ), .dout(n6683));
  jnot g06450(.din(n6445), .dout(n6684));
  jand g06451(.dina(n6684), .dinb(n6683), .dout(n6685));
  jor  g06452(.dina(n6685), .dinb(n6637), .dout(n6686));
  jor  g06453(.dina(n6686), .dinb(asqrt[44] ), .dout(n6687));
  jand g06454(.dina(n6452), .dinb(n6687), .dout(n6688));
  jor  g06455(.dina(n6688), .dinb(n6636), .dout(n6689));
  jor  g06456(.dina(n6689), .dinb(asqrt[45] ), .dout(n6690));
  jand g06457(.dina(n6460), .dinb(n6690), .dout(n6691));
  jor  g06458(.dina(n6691), .dinb(n6635), .dout(n6692));
  jor  g06459(.dina(n6692), .dinb(asqrt[46] ), .dout(n6693));
  jand g06460(.dina(n6468), .dinb(n6693), .dout(n6694));
  jor  g06461(.dina(n6694), .dinb(n6634), .dout(n6695));
  jor  g06462(.dina(n6695), .dinb(asqrt[47] ), .dout(n6696));
  jnot g06463(.din(n6476), .dout(n6697));
  jand g06464(.dina(n6697), .dinb(n6696), .dout(n6698));
  jor  g06465(.dina(n6698), .dinb(n6633), .dout(n6699));
  jor  g06466(.dina(n6699), .dinb(asqrt[48] ), .dout(n6700));
  jnot g06467(.din(n6483), .dout(n6701));
  jand g06468(.dina(n6701), .dinb(n6700), .dout(n6702));
  jor  g06469(.dina(n6702), .dinb(n6632), .dout(n6703));
  jor  g06470(.dina(n6703), .dinb(asqrt[49] ), .dout(n6704));
  jnot g06471(.din(n6490), .dout(n6705));
  jand g06472(.dina(n6705), .dinb(n6704), .dout(n6706));
  jor  g06473(.dina(n6706), .dinb(n6631), .dout(n6707));
  jor  g06474(.dina(n6707), .dinb(asqrt[50] ), .dout(n6708));
  jand g06475(.dina(n6497), .dinb(n6708), .dout(n6709));
  jor  g06476(.dina(n6709), .dinb(n6630), .dout(n6710));
  jor  g06477(.dina(n6710), .dinb(asqrt[51] ), .dout(n6711));
  jnot g06478(.din(n6505), .dout(n6712));
  jand g06479(.dina(n6712), .dinb(n6711), .dout(n6713));
  jor  g06480(.dina(n6713), .dinb(n6629), .dout(n6714));
  jor  g06481(.dina(n6714), .dinb(asqrt[52] ), .dout(n6715));
  jand g06482(.dina(n6512), .dinb(n6715), .dout(n6716));
  jor  g06483(.dina(n6716), .dinb(n6628), .dout(n6717));
  jor  g06484(.dina(n6717), .dinb(asqrt[53] ), .dout(n6718));
  jnot g06485(.din(n6520), .dout(n6719));
  jand g06486(.dina(n6719), .dinb(n6718), .dout(n6720));
  jor  g06487(.dina(n6720), .dinb(n6627), .dout(n6721));
  jor  g06488(.dina(n6721), .dinb(asqrt[54] ), .dout(n6722));
  jand g06489(.dina(n6527), .dinb(n6722), .dout(n6723));
  jor  g06490(.dina(n6723), .dinb(n6626), .dout(n6724));
  jor  g06491(.dina(n6724), .dinb(asqrt[55] ), .dout(n6725));
  jand g06492(.dina(n6535), .dinb(n6725), .dout(n6726));
  jor  g06493(.dina(n6726), .dinb(n6625), .dout(n6727));
  jor  g06494(.dina(n6727), .dinb(asqrt[56] ), .dout(n6728));
  jnot g06495(.din(n6543), .dout(n6729));
  jand g06496(.dina(n6729), .dinb(n6728), .dout(n6730));
  jor  g06497(.dina(n6730), .dinb(n6624), .dout(n6731));
  jor  g06498(.dina(n6731), .dinb(asqrt[57] ), .dout(n6732));
  jnot g06499(.din(n6550), .dout(n6733));
  jand g06500(.dina(n6733), .dinb(n6732), .dout(n6734));
  jor  g06501(.dina(n6734), .dinb(n6623), .dout(n6735));
  jor  g06502(.dina(n6735), .dinb(asqrt[58] ), .dout(n6736));
  jand g06503(.dina(n6557), .dinb(n6736), .dout(n6737));
  jor  g06504(.dina(n6737), .dinb(n6622), .dout(n6738));
  jor  g06505(.dina(n6738), .dinb(asqrt[59] ), .dout(n6739));
  jand g06506(.dina(n6565), .dinb(n6739), .dout(n6740));
  jor  g06507(.dina(n6740), .dinb(n6621), .dout(n6741));
  jor  g06508(.dina(n6741), .dinb(asqrt[60] ), .dout(n6742));
  jand g06509(.dina(n6573), .dinb(n6742), .dout(n6743));
  jor  g06510(.dina(n6743), .dinb(n6620), .dout(n6744));
  jor  g06511(.dina(n6744), .dinb(asqrt[61] ), .dout(n6745));
  jnot g06512(.din(n6581), .dout(n6746));
  jand g06513(.dina(n6746), .dinb(n6745), .dout(n6747));
  jor  g06514(.dina(n6747), .dinb(n6619), .dout(n6748));
  jor  g06515(.dina(n6748), .dinb(asqrt[62] ), .dout(n6749));
  jnot g06516(.din(n6588), .dout(n6750));
  jand g06517(.dina(n6750), .dinb(n6749), .dout(n6751));
  jor  g06518(.dina(n6751), .dinb(n6618), .dout(n6752));
  jand g06519(.dina(n6752), .dinb(n6360), .dout(n6753));
  jand g06520(.dina(n6753), .dinb(n6201), .dout(n6754));
  jand g06521(.dina(n6754), .dinb(n6617), .dout(n6755));
  jor  g06522(.dina(n6755), .dinb(asqrt[63] ), .dout(n6756));
  jnot g06523(.din(n6604), .dout(n6757));
  jand g06524(.dina(n6757), .dinb(n6756), .dout(n6758));
  jor  g06525(.dina(n6758), .dinb(n6616), .dout(n6759));
  jand g06526(.dina(n6759), .dinb(n6615), .dout(n6760));
  jand g06527(.dina(n6760), .dinb(n6613), .dout(n6761));
  jor  g06528(.dina(n6761), .dinb(n6612), .dout(n6762));
  jand g06529(.dina(n6762), .dinb(asqrt[34] ), .dout(n6763));
  jor  g06530(.dina(n6762), .dinb(asqrt[34] ), .dout(n6764));
  jand g06531(.dina(asqrt[32] ), .dinb(n6364), .dout(n6765));
  jnot g06532(.din(n6596), .dout(n6766));
  jand g06533(.dina(n6601), .dinb(asqrt[33] ), .dout(n6767));
  jand g06534(.dina(n6767), .dinb(n6766), .dout(n6768));
  jand g06535(.dina(n6768), .dinb(n6756), .dout(n6769));
  jor  g06536(.dina(n6769), .dinb(n6765), .dout(n6770));
  jxor g06537(.dina(n6770), .dinb(a[66] ), .dout(n6771));
  jnot g06538(.din(n6771), .dout(n6772));
  jand g06539(.dina(n6772), .dinb(n6764), .dout(n6773));
  jor  g06540(.dina(n6773), .dinb(n6763), .dout(n6774));
  jand g06541(.dina(n6774), .dinb(asqrt[35] ), .dout(n6775));
  jor  g06542(.dina(n6774), .dinb(asqrt[35] ), .dout(n6776));
  jxor g06543(.dina(n6368), .dinb(n5989), .dout(n6777));
  jand g06544(.dina(n6777), .dinb(asqrt[32] ), .dout(n6778));
  jxor g06545(.dina(n6778), .dinb(n6652), .dout(n6779));
  jand g06546(.dina(n6779), .dinb(n6776), .dout(n6780));
  jor  g06547(.dina(n6780), .dinb(n6775), .dout(n6781));
  jand g06548(.dina(n6781), .dinb(asqrt[36] ), .dout(n6782));
  jor  g06549(.dina(n6781), .dinb(asqrt[36] ), .dout(n6783));
  jxor g06550(.dina(n6376), .dinb(n5606), .dout(n6784));
  jand g06551(.dina(n6784), .dinb(asqrt[32] ), .dout(n6785));
  jxor g06552(.dina(n6785), .dinb(n6656), .dout(n6786));
  jand g06553(.dina(n6786), .dinb(n6783), .dout(n6787));
  jor  g06554(.dina(n6787), .dinb(n6782), .dout(n6788));
  jand g06555(.dina(n6788), .dinb(asqrt[37] ), .dout(n6789));
  jor  g06556(.dina(n6788), .dinb(asqrt[37] ), .dout(n6790));
  jxor g06557(.dina(n6387), .dinb(n5259), .dout(n6791));
  jand g06558(.dina(n6791), .dinb(asqrt[32] ), .dout(n6792));
  jxor g06559(.dina(n6792), .dinb(n6392), .dout(n6793));
  jand g06560(.dina(n6793), .dinb(n6790), .dout(n6794));
  jor  g06561(.dina(n6794), .dinb(n6789), .dout(n6795));
  jand g06562(.dina(n6795), .dinb(asqrt[38] ), .dout(n6796));
  jor  g06563(.dina(n6795), .dinb(asqrt[38] ), .dout(n6797));
  jxor g06564(.dina(n6395), .dinb(n4902), .dout(n6798));
  jand g06565(.dina(n6798), .dinb(asqrt[32] ), .dout(n6799));
  jxor g06566(.dina(n6799), .dinb(n6400), .dout(n6800));
  jnot g06567(.din(n6800), .dout(n6801));
  jand g06568(.dina(n6801), .dinb(n6797), .dout(n6802));
  jor  g06569(.dina(n6802), .dinb(n6796), .dout(n6803));
  jand g06570(.dina(n6803), .dinb(asqrt[39] ), .dout(n6804));
  jor  g06571(.dina(n6803), .dinb(asqrt[39] ), .dout(n6805));
  jxor g06572(.dina(n6402), .dinb(n4582), .dout(n6806));
  jand g06573(.dina(n6806), .dinb(asqrt[32] ), .dout(n6807));
  jxor g06574(.dina(n6807), .dinb(n6407), .dout(n6808));
  jand g06575(.dina(n6808), .dinb(n6805), .dout(n6809));
  jor  g06576(.dina(n6809), .dinb(n6804), .dout(n6810));
  jand g06577(.dina(n6810), .dinb(asqrt[40] ), .dout(n6811));
  jor  g06578(.dina(n6810), .dinb(asqrt[40] ), .dout(n6812));
  jxor g06579(.dina(n6410), .dinb(n4249), .dout(n6813));
  jand g06580(.dina(n6813), .dinb(asqrt[32] ), .dout(n6814));
  jxor g06581(.dina(n6814), .dinb(n6415), .dout(n6815));
  jnot g06582(.din(n6815), .dout(n6816));
  jand g06583(.dina(n6816), .dinb(n6812), .dout(n6817));
  jor  g06584(.dina(n6817), .dinb(n6811), .dout(n6818));
  jand g06585(.dina(n6818), .dinb(asqrt[41] ), .dout(n6819));
  jor  g06586(.dina(n6818), .dinb(asqrt[41] ), .dout(n6820));
  jxor g06587(.dina(n6417), .dinb(n3955), .dout(n6821));
  jand g06588(.dina(n6821), .dinb(asqrt[32] ), .dout(n6822));
  jxor g06589(.dina(n6822), .dinb(n6422), .dout(n6823));
  jand g06590(.dina(n6823), .dinb(n6820), .dout(n6824));
  jor  g06591(.dina(n6824), .dinb(n6819), .dout(n6825));
  jand g06592(.dina(n6825), .dinb(asqrt[42] ), .dout(n6826));
  jor  g06593(.dina(n6825), .dinb(asqrt[42] ), .dout(n6827));
  jxor g06594(.dina(n6425), .dinb(n3642), .dout(n6828));
  jand g06595(.dina(n6828), .dinb(asqrt[32] ), .dout(n6829));
  jxor g06596(.dina(n6829), .dinb(n6430), .dout(n6830));
  jnot g06597(.din(n6830), .dout(n6831));
  jand g06598(.dina(n6831), .dinb(n6827), .dout(n6832));
  jor  g06599(.dina(n6832), .dinb(n6826), .dout(n6833));
  jand g06600(.dina(n6833), .dinb(asqrt[43] ), .dout(n6834));
  jor  g06601(.dina(n6833), .dinb(asqrt[43] ), .dout(n6835));
  jxor g06602(.dina(n6432), .dinb(n3368), .dout(n6836));
  jand g06603(.dina(n6836), .dinb(asqrt[32] ), .dout(n6837));
  jxor g06604(.dina(n6837), .dinb(n6437), .dout(n6838));
  jand g06605(.dina(n6838), .dinb(n6835), .dout(n6839));
  jor  g06606(.dina(n6839), .dinb(n6834), .dout(n6840));
  jand g06607(.dina(n6840), .dinb(asqrt[44] ), .dout(n6841));
  jor  g06608(.dina(n6840), .dinb(asqrt[44] ), .dout(n6842));
  jxor g06609(.dina(n6440), .dinb(n3089), .dout(n6843));
  jand g06610(.dina(n6843), .dinb(asqrt[32] ), .dout(n6844));
  jxor g06611(.dina(n6844), .dinb(n6445), .dout(n6845));
  jnot g06612(.din(n6845), .dout(n6846));
  jand g06613(.dina(n6846), .dinb(n6842), .dout(n6847));
  jor  g06614(.dina(n6847), .dinb(n6841), .dout(n6848));
  jand g06615(.dina(n6848), .dinb(asqrt[45] ), .dout(n6849));
  jor  g06616(.dina(n6848), .dinb(asqrt[45] ), .dout(n6850));
  jxor g06617(.dina(n6447), .dinb(n2833), .dout(n6851));
  jand g06618(.dina(n6851), .dinb(asqrt[32] ), .dout(n6852));
  jxor g06619(.dina(n6852), .dinb(n6452), .dout(n6853));
  jand g06620(.dina(n6853), .dinb(n6850), .dout(n6854));
  jor  g06621(.dina(n6854), .dinb(n6849), .dout(n6855));
  jand g06622(.dina(n6855), .dinb(asqrt[46] ), .dout(n6856));
  jor  g06623(.dina(n6855), .dinb(asqrt[46] ), .dout(n6857));
  jxor g06624(.dina(n6455), .dinb(n2572), .dout(n6858));
  jand g06625(.dina(n6858), .dinb(asqrt[32] ), .dout(n6859));
  jxor g06626(.dina(n6859), .dinb(n6460), .dout(n6860));
  jand g06627(.dina(n6860), .dinb(n6857), .dout(n6861));
  jor  g06628(.dina(n6861), .dinb(n6856), .dout(n6862));
  jand g06629(.dina(n6862), .dinb(asqrt[47] ), .dout(n6863));
  jor  g06630(.dina(n6862), .dinb(asqrt[47] ), .dout(n6864));
  jxor g06631(.dina(n6463), .dinb(n2345), .dout(n6865));
  jand g06632(.dina(n6865), .dinb(asqrt[32] ), .dout(n6866));
  jxor g06633(.dina(n6866), .dinb(n6468), .dout(n6867));
  jand g06634(.dina(n6867), .dinb(n6864), .dout(n6868));
  jor  g06635(.dina(n6868), .dinb(n6863), .dout(n6869));
  jand g06636(.dina(n6869), .dinb(asqrt[48] ), .dout(n6870));
  jor  g06637(.dina(n6869), .dinb(asqrt[48] ), .dout(n6871));
  jxor g06638(.dina(n6471), .dinb(n2108), .dout(n6872));
  jand g06639(.dina(n6872), .dinb(asqrt[32] ), .dout(n6873));
  jxor g06640(.dina(n6873), .dinb(n6476), .dout(n6874));
  jnot g06641(.din(n6874), .dout(n6875));
  jand g06642(.dina(n6875), .dinb(n6871), .dout(n6876));
  jor  g06643(.dina(n6876), .dinb(n6870), .dout(n6877));
  jand g06644(.dina(n6877), .dinb(asqrt[49] ), .dout(n6878));
  jor  g06645(.dina(n6877), .dinb(asqrt[49] ), .dout(n6879));
  jxor g06646(.dina(n6478), .dinb(n1912), .dout(n6880));
  jand g06647(.dina(n6880), .dinb(asqrt[32] ), .dout(n6881));
  jxor g06648(.dina(n6881), .dinb(n6483), .dout(n6882));
  jnot g06649(.din(n6882), .dout(n6883));
  jand g06650(.dina(n6883), .dinb(n6879), .dout(n6884));
  jor  g06651(.dina(n6884), .dinb(n6878), .dout(n6885));
  jand g06652(.dina(n6885), .dinb(asqrt[50] ), .dout(n6886));
  jor  g06653(.dina(n6885), .dinb(asqrt[50] ), .dout(n6887));
  jxor g06654(.dina(n6485), .dinb(n1699), .dout(n6888));
  jand g06655(.dina(n6888), .dinb(asqrt[32] ), .dout(n6889));
  jxor g06656(.dina(n6889), .dinb(n6490), .dout(n6890));
  jnot g06657(.din(n6890), .dout(n6891));
  jand g06658(.dina(n6891), .dinb(n6887), .dout(n6892));
  jor  g06659(.dina(n6892), .dinb(n6886), .dout(n6893));
  jand g06660(.dina(n6893), .dinb(asqrt[51] ), .dout(n6894));
  jor  g06661(.dina(n6893), .dinb(asqrt[51] ), .dout(n6895));
  jxor g06662(.dina(n6492), .dinb(n1516), .dout(n6896));
  jand g06663(.dina(n6896), .dinb(asqrt[32] ), .dout(n6897));
  jxor g06664(.dina(n6897), .dinb(n6497), .dout(n6898));
  jand g06665(.dina(n6898), .dinb(n6895), .dout(n6899));
  jor  g06666(.dina(n6899), .dinb(n6894), .dout(n6900));
  jand g06667(.dina(n6900), .dinb(asqrt[52] ), .dout(n6901));
  jor  g06668(.dina(n6900), .dinb(asqrt[52] ), .dout(n6902));
  jxor g06669(.dina(n6500), .dinb(n1332), .dout(n6903));
  jand g06670(.dina(n6903), .dinb(asqrt[32] ), .dout(n6904));
  jxor g06671(.dina(n6904), .dinb(n6505), .dout(n6905));
  jnot g06672(.din(n6905), .dout(n6906));
  jand g06673(.dina(n6906), .dinb(n6902), .dout(n6907));
  jor  g06674(.dina(n6907), .dinb(n6901), .dout(n6908));
  jand g06675(.dina(n6908), .dinb(asqrt[53] ), .dout(n6909));
  jor  g06676(.dina(n6908), .dinb(asqrt[53] ), .dout(n6910));
  jxor g06677(.dina(n6507), .dinb(n1173), .dout(n6911));
  jand g06678(.dina(n6911), .dinb(asqrt[32] ), .dout(n6912));
  jxor g06679(.dina(n6912), .dinb(n6512), .dout(n6913));
  jand g06680(.dina(n6913), .dinb(n6910), .dout(n6914));
  jor  g06681(.dina(n6914), .dinb(n6909), .dout(n6915));
  jand g06682(.dina(n6915), .dinb(asqrt[54] ), .dout(n6916));
  jor  g06683(.dina(n6915), .dinb(asqrt[54] ), .dout(n6917));
  jxor g06684(.dina(n6515), .dinb(n1008), .dout(n6918));
  jand g06685(.dina(n6918), .dinb(asqrt[32] ), .dout(n6919));
  jxor g06686(.dina(n6919), .dinb(n6520), .dout(n6920));
  jnot g06687(.din(n6920), .dout(n6921));
  jand g06688(.dina(n6921), .dinb(n6917), .dout(n6922));
  jor  g06689(.dina(n6922), .dinb(n6916), .dout(n6923));
  jand g06690(.dina(n6923), .dinb(asqrt[55] ), .dout(n6924));
  jor  g06691(.dina(n6923), .dinb(asqrt[55] ), .dout(n6925));
  jxor g06692(.dina(n6522), .dinb(n884), .dout(n6926));
  jand g06693(.dina(n6926), .dinb(asqrt[32] ), .dout(n6927));
  jxor g06694(.dina(n6927), .dinb(n6527), .dout(n6928));
  jand g06695(.dina(n6928), .dinb(n6925), .dout(n6929));
  jor  g06696(.dina(n6929), .dinb(n6924), .dout(n6930));
  jand g06697(.dina(n6930), .dinb(asqrt[56] ), .dout(n6931));
  jor  g06698(.dina(n6930), .dinb(asqrt[56] ), .dout(n6932));
  jxor g06699(.dina(n6530), .dinb(n743), .dout(n6933));
  jand g06700(.dina(n6933), .dinb(asqrt[32] ), .dout(n6934));
  jxor g06701(.dina(n6934), .dinb(n6535), .dout(n6935));
  jand g06702(.dina(n6935), .dinb(n6932), .dout(n6936));
  jor  g06703(.dina(n6936), .dinb(n6931), .dout(n6937));
  jand g06704(.dina(n6937), .dinb(asqrt[57] ), .dout(n6938));
  jor  g06705(.dina(n6937), .dinb(asqrt[57] ), .dout(n6939));
  jxor g06706(.dina(n6538), .dinb(n635), .dout(n6940));
  jand g06707(.dina(n6940), .dinb(asqrt[32] ), .dout(n6941));
  jxor g06708(.dina(n6941), .dinb(n6543), .dout(n6942));
  jnot g06709(.din(n6942), .dout(n6943));
  jand g06710(.dina(n6943), .dinb(n6939), .dout(n6944));
  jor  g06711(.dina(n6944), .dinb(n6938), .dout(n6945));
  jand g06712(.dina(n6945), .dinb(asqrt[58] ), .dout(n6946));
  jor  g06713(.dina(n6945), .dinb(asqrt[58] ), .dout(n6947));
  jxor g06714(.dina(n6545), .dinb(n515), .dout(n6948));
  jand g06715(.dina(n6948), .dinb(asqrt[32] ), .dout(n6949));
  jxor g06716(.dina(n6949), .dinb(n6550), .dout(n6950));
  jnot g06717(.din(n6950), .dout(n6951));
  jand g06718(.dina(n6951), .dinb(n6947), .dout(n6952));
  jor  g06719(.dina(n6952), .dinb(n6946), .dout(n6953));
  jand g06720(.dina(n6953), .dinb(asqrt[59] ), .dout(n6954));
  jor  g06721(.dina(n6953), .dinb(asqrt[59] ), .dout(n6955));
  jxor g06722(.dina(n6552), .dinb(n443), .dout(n6956));
  jand g06723(.dina(n6956), .dinb(asqrt[32] ), .dout(n6957));
  jxor g06724(.dina(n6957), .dinb(n6558), .dout(n6958));
  jnot g06725(.din(n6958), .dout(n6959));
  jand g06726(.dina(n6959), .dinb(n6955), .dout(n6960));
  jor  g06727(.dina(n6960), .dinb(n6954), .dout(n6961));
  jand g06728(.dina(n6961), .dinb(asqrt[60] ), .dout(n6962));
  jor  g06729(.dina(n6961), .dinb(asqrt[60] ), .dout(n6963));
  jxor g06730(.dina(n6560), .dinb(n352), .dout(n6964));
  jand g06731(.dina(n6964), .dinb(asqrt[32] ), .dout(n6965));
  jxor g06732(.dina(n6965), .dinb(n6565), .dout(n6966));
  jand g06733(.dina(n6966), .dinb(n6963), .dout(n6967));
  jor  g06734(.dina(n6967), .dinb(n6962), .dout(n6968));
  jand g06735(.dina(n6968), .dinb(asqrt[61] ), .dout(n6969));
  jor  g06736(.dina(n6968), .dinb(asqrt[61] ), .dout(n6970));
  jxor g06737(.dina(n6568), .dinb(n294), .dout(n6971));
  jand g06738(.dina(n6971), .dinb(asqrt[32] ), .dout(n6972));
  jxor g06739(.dina(n6972), .dinb(n6573), .dout(n6973));
  jand g06740(.dina(n6973), .dinb(n6970), .dout(n6974));
  jor  g06741(.dina(n6974), .dinb(n6969), .dout(n6975));
  jand g06742(.dina(n6975), .dinb(asqrt[62] ), .dout(n6976));
  jor  g06743(.dina(n6975), .dinb(asqrt[62] ), .dout(n6977));
  jxor g06744(.dina(n6576), .dinb(n239), .dout(n6978));
  jand g06745(.dina(n6978), .dinb(asqrt[32] ), .dout(n6979));
  jxor g06746(.dina(n6979), .dinb(n6581), .dout(n6980));
  jnot g06747(.din(n6980), .dout(n6981));
  jand g06748(.dina(n6981), .dinb(n6977), .dout(n6982));
  jor  g06749(.dina(n6982), .dinb(n6976), .dout(n6983));
  jxor g06750(.dina(n6583), .dinb(n221), .dout(n6984));
  jand g06751(.dina(n6984), .dinb(asqrt[32] ), .dout(n6985));
  jxor g06752(.dina(n6985), .dinb(n6588), .dout(n6986));
  jnot g06753(.din(n6986), .dout(n6987));
  jor  g06754(.dina(n6987), .dinb(n6983), .dout(n6988));
  jnot g06755(.din(n6988), .dout(n6989));
  jand g06756(.dina(n6758), .dinb(n6590), .dout(n6990));
  jnot g06757(.din(n6990), .dout(n6991));
  jand g06758(.dina(n6591), .dinb(asqrt[63] ), .dout(n6992));
  jand g06759(.dina(n6992), .dinb(n6766), .dout(n6993));
  jand g06760(.dina(n6993), .dinb(n6991), .dout(n6994));
  jnot g06761(.din(n6976), .dout(n6995));
  jnot g06762(.din(n6969), .dout(n6996));
  jnot g06763(.din(n6962), .dout(n6997));
  jnot g06764(.din(n6954), .dout(n6998));
  jnot g06765(.din(n6946), .dout(n6999));
  jnot g06766(.din(n6938), .dout(n7000));
  jnot g06767(.din(n6931), .dout(n7001));
  jnot g06768(.din(n6924), .dout(n7002));
  jnot g06769(.din(n6916), .dout(n7003));
  jnot g06770(.din(n6909), .dout(n7004));
  jnot g06771(.din(n6901), .dout(n7005));
  jnot g06772(.din(n6894), .dout(n7006));
  jnot g06773(.din(n6886), .dout(n7007));
  jnot g06774(.din(n6878), .dout(n7008));
  jnot g06775(.din(n6870), .dout(n7009));
  jnot g06776(.din(n6863), .dout(n7010));
  jnot g06777(.din(n6856), .dout(n7011));
  jnot g06778(.din(n6849), .dout(n7012));
  jnot g06779(.din(n6841), .dout(n7013));
  jnot g06780(.din(n6834), .dout(n7014));
  jnot g06781(.din(n6826), .dout(n7015));
  jnot g06782(.din(n6819), .dout(n7016));
  jnot g06783(.din(n6811), .dout(n7017));
  jnot g06784(.din(n6804), .dout(n7018));
  jnot g06785(.din(n6796), .dout(n7019));
  jnot g06786(.din(n6789), .dout(n7020));
  jnot g06787(.din(n6782), .dout(n7021));
  jnot g06788(.din(n6775), .dout(n7022));
  jnot g06789(.din(n6763), .dout(n7023));
  jnot g06790(.din(n6612), .dout(n7024));
  jnot g06791(.din(n6609), .dout(n7025));
  jor  g06792(.dina(n6758), .dinb(n6362), .dout(n7026));
  jand g06793(.dina(n7026), .dinb(n7025), .dout(n7027));
  jand g06794(.dina(n7027), .dinb(n6357), .dout(n7028));
  jor  g06795(.dina(n6758), .dinb(a[64] ), .dout(n7029));
  jand g06796(.dina(n7029), .dinb(a[65] ), .dout(n7030));
  jor  g06797(.dina(n6765), .dinb(n7030), .dout(n7031));
  jor  g06798(.dina(n7031), .dinb(n7028), .dout(n7032));
  jand g06799(.dina(n7032), .dinb(n7024), .dout(n7033));
  jand g06800(.dina(n7033), .dinb(n5989), .dout(n7034));
  jor  g06801(.dina(n6771), .dinb(n7034), .dout(n7035));
  jand g06802(.dina(n7035), .dinb(n7023), .dout(n7036));
  jand g06803(.dina(n7036), .dinb(n5606), .dout(n7037));
  jnot g06804(.din(n6779), .dout(n7038));
  jor  g06805(.dina(n7038), .dinb(n7037), .dout(n7039));
  jand g06806(.dina(n7039), .dinb(n7022), .dout(n7040));
  jand g06807(.dina(n7040), .dinb(n5259), .dout(n7041));
  jnot g06808(.din(n6786), .dout(n7042));
  jor  g06809(.dina(n7042), .dinb(n7041), .dout(n7043));
  jand g06810(.dina(n7043), .dinb(n7021), .dout(n7044));
  jand g06811(.dina(n7044), .dinb(n4902), .dout(n7045));
  jnot g06812(.din(n6793), .dout(n7046));
  jor  g06813(.dina(n7046), .dinb(n7045), .dout(n7047));
  jand g06814(.dina(n7047), .dinb(n7020), .dout(n7048));
  jand g06815(.dina(n7048), .dinb(n4582), .dout(n7049));
  jor  g06816(.dina(n6800), .dinb(n7049), .dout(n7050));
  jand g06817(.dina(n7050), .dinb(n7019), .dout(n7051));
  jand g06818(.dina(n7051), .dinb(n4249), .dout(n7052));
  jnot g06819(.din(n6808), .dout(n7053));
  jor  g06820(.dina(n7053), .dinb(n7052), .dout(n7054));
  jand g06821(.dina(n7054), .dinb(n7018), .dout(n7055));
  jand g06822(.dina(n7055), .dinb(n3955), .dout(n7056));
  jor  g06823(.dina(n6815), .dinb(n7056), .dout(n7057));
  jand g06824(.dina(n7057), .dinb(n7017), .dout(n7058));
  jand g06825(.dina(n7058), .dinb(n3642), .dout(n7059));
  jnot g06826(.din(n6823), .dout(n7060));
  jor  g06827(.dina(n7060), .dinb(n7059), .dout(n7061));
  jand g06828(.dina(n7061), .dinb(n7016), .dout(n7062));
  jand g06829(.dina(n7062), .dinb(n3368), .dout(n7063));
  jor  g06830(.dina(n6830), .dinb(n7063), .dout(n7064));
  jand g06831(.dina(n7064), .dinb(n7015), .dout(n7065));
  jand g06832(.dina(n7065), .dinb(n3089), .dout(n7066));
  jnot g06833(.din(n6838), .dout(n7067));
  jor  g06834(.dina(n7067), .dinb(n7066), .dout(n7068));
  jand g06835(.dina(n7068), .dinb(n7014), .dout(n7069));
  jand g06836(.dina(n7069), .dinb(n2833), .dout(n7070));
  jor  g06837(.dina(n6845), .dinb(n7070), .dout(n7071));
  jand g06838(.dina(n7071), .dinb(n7013), .dout(n7072));
  jand g06839(.dina(n7072), .dinb(n2572), .dout(n7073));
  jnot g06840(.din(n6853), .dout(n7074));
  jor  g06841(.dina(n7074), .dinb(n7073), .dout(n7075));
  jand g06842(.dina(n7075), .dinb(n7012), .dout(n7076));
  jand g06843(.dina(n7076), .dinb(n2345), .dout(n7077));
  jnot g06844(.din(n6860), .dout(n7078));
  jor  g06845(.dina(n7078), .dinb(n7077), .dout(n7079));
  jand g06846(.dina(n7079), .dinb(n7011), .dout(n7080));
  jand g06847(.dina(n7080), .dinb(n2108), .dout(n7081));
  jnot g06848(.din(n6867), .dout(n7082));
  jor  g06849(.dina(n7082), .dinb(n7081), .dout(n7083));
  jand g06850(.dina(n7083), .dinb(n7010), .dout(n7084));
  jand g06851(.dina(n7084), .dinb(n1912), .dout(n7085));
  jor  g06852(.dina(n6874), .dinb(n7085), .dout(n7086));
  jand g06853(.dina(n7086), .dinb(n7009), .dout(n7087));
  jand g06854(.dina(n7087), .dinb(n1699), .dout(n7088));
  jor  g06855(.dina(n6882), .dinb(n7088), .dout(n7089));
  jand g06856(.dina(n7089), .dinb(n7008), .dout(n7090));
  jand g06857(.dina(n7090), .dinb(n1516), .dout(n7091));
  jor  g06858(.dina(n6890), .dinb(n7091), .dout(n7092));
  jand g06859(.dina(n7092), .dinb(n7007), .dout(n7093));
  jand g06860(.dina(n7093), .dinb(n1332), .dout(n7094));
  jnot g06861(.din(n6898), .dout(n7095));
  jor  g06862(.dina(n7095), .dinb(n7094), .dout(n7096));
  jand g06863(.dina(n7096), .dinb(n7006), .dout(n7097));
  jand g06864(.dina(n7097), .dinb(n1173), .dout(n7098));
  jor  g06865(.dina(n6905), .dinb(n7098), .dout(n7099));
  jand g06866(.dina(n7099), .dinb(n7005), .dout(n7100));
  jand g06867(.dina(n7100), .dinb(n1008), .dout(n7101));
  jnot g06868(.din(n6913), .dout(n7102));
  jor  g06869(.dina(n7102), .dinb(n7101), .dout(n7103));
  jand g06870(.dina(n7103), .dinb(n7004), .dout(n7104));
  jand g06871(.dina(n7104), .dinb(n884), .dout(n7105));
  jor  g06872(.dina(n6920), .dinb(n7105), .dout(n7106));
  jand g06873(.dina(n7106), .dinb(n7003), .dout(n7107));
  jand g06874(.dina(n7107), .dinb(n743), .dout(n7108));
  jnot g06875(.din(n6928), .dout(n7109));
  jor  g06876(.dina(n7109), .dinb(n7108), .dout(n7110));
  jand g06877(.dina(n7110), .dinb(n7002), .dout(n7111));
  jand g06878(.dina(n7111), .dinb(n635), .dout(n7112));
  jnot g06879(.din(n6935), .dout(n7113));
  jor  g06880(.dina(n7113), .dinb(n7112), .dout(n7114));
  jand g06881(.dina(n7114), .dinb(n7001), .dout(n7115));
  jand g06882(.dina(n7115), .dinb(n515), .dout(n7116));
  jor  g06883(.dina(n6942), .dinb(n7116), .dout(n7117));
  jand g06884(.dina(n7117), .dinb(n7000), .dout(n7118));
  jand g06885(.dina(n7118), .dinb(n443), .dout(n7119));
  jor  g06886(.dina(n6950), .dinb(n7119), .dout(n7120));
  jand g06887(.dina(n7120), .dinb(n6999), .dout(n7121));
  jand g06888(.dina(n7121), .dinb(n352), .dout(n7122));
  jor  g06889(.dina(n6958), .dinb(n7122), .dout(n7123));
  jand g06890(.dina(n7123), .dinb(n6998), .dout(n7124));
  jand g06891(.dina(n7124), .dinb(n294), .dout(n7125));
  jnot g06892(.din(n6966), .dout(n7126));
  jor  g06893(.dina(n7126), .dinb(n7125), .dout(n7127));
  jand g06894(.dina(n7127), .dinb(n6997), .dout(n7128));
  jand g06895(.dina(n7128), .dinb(n239), .dout(n7129));
  jnot g06896(.din(n6973), .dout(n7130));
  jor  g06897(.dina(n7130), .dinb(n7129), .dout(n7131));
  jand g06898(.dina(n7131), .dinb(n6996), .dout(n7132));
  jand g06899(.dina(n7132), .dinb(n221), .dout(n7133));
  jor  g06900(.dina(n6980), .dinb(n7133), .dout(n7134));
  jand g06901(.dina(n7134), .dinb(n6995), .dout(n7135));
  jor  g06902(.dina(n6986), .dinb(n7135), .dout(n7136));
  jand g06903(.dina(asqrt[32] ), .dinb(n6753), .dout(n7137));
  jor  g06904(.dina(n7137), .dinb(n6596), .dout(n7138));
  jor  g06905(.dina(n7138), .dinb(n7136), .dout(n7139));
  jand g06906(.dina(n7139), .dinb(n218), .dout(n7140));
  jand g06907(.dina(n6758), .dinb(n6361), .dout(n7141));
  jor  g06908(.dina(n7141), .dinb(n7140), .dout(n7142));
  jor  g06909(.dina(n7142), .dinb(n6994), .dout(n7143));
  jor  g06910(.dina(n7143), .dinb(n6989), .dout(asqrt[31] ));
  jand g06911(.dina(n6987), .dinb(n6983), .dout(n7145));
  jand g06912(.dina(n7143), .dinb(n7145), .dout(n7146));
  jnot g06913(.din(n6994), .dout(n7147));
  jnot g06914(.din(n7138), .dout(n7148));
  jand g06915(.dina(n7148), .dinb(n7145), .dout(n7149));
  jor  g06916(.dina(n7149), .dinb(asqrt[63] ), .dout(n7150));
  jnot g06917(.din(n7141), .dout(n7151));
  jand g06918(.dina(n7151), .dinb(n7150), .dout(n7152));
  jand g06919(.dina(n7152), .dinb(n7147), .dout(n7153));
  jand g06920(.dina(n7153), .dinb(n6988), .dout(n7154));
  jor  g06921(.dina(n7154), .dinb(n6606), .dout(n7155));
  jnot g06922(.din(a[60] ), .dout(n7156));
  jnot g06923(.din(a[61] ), .dout(n7157));
  jand g06924(.dina(n7157), .dinb(n7156), .dout(n7158));
  jand g06925(.dina(n7158), .dinb(n6606), .dout(n7159));
  jnot g06926(.din(n7159), .dout(n7160));
  jand g06927(.dina(n7160), .dinb(n7155), .dout(n7161));
  jor  g06928(.dina(n7161), .dinb(n6758), .dout(n7162));
  jand g06929(.dina(asqrt[31] ), .dinb(n6608), .dout(n7163));
  jor  g06930(.dina(n7154), .dinb(a[62] ), .dout(n7164));
  jand g06931(.dina(n7164), .dinb(a[63] ), .dout(n7165));
  jor  g06932(.dina(n7165), .dinb(n7163), .dout(n7166));
  jand g06933(.dina(n7161), .dinb(n6758), .dout(n7167));
  jor  g06934(.dina(n7167), .dinb(n7166), .dout(n7168));
  jand g06935(.dina(n7168), .dinb(n7162), .dout(n7169));
  jor  g06936(.dina(n7169), .dinb(n6357), .dout(n7170));
  jand g06937(.dina(n7169), .dinb(n6357), .dout(n7171));
  jnot g06938(.din(n6608), .dout(n7172));
  jor  g06939(.dina(n7154), .dinb(n7172), .dout(n7173));
  jor  g06940(.dina(n6989), .dinb(n6758), .dout(n7174));
  jor  g06941(.dina(n7174), .dinb(n6993), .dout(n7175));
  jor  g06942(.dina(n7175), .dinb(n7140), .dout(n7176));
  jand g06943(.dina(n7176), .dinb(n7173), .dout(n7177));
  jxor g06944(.dina(n7177), .dinb(n6362), .dout(n7178));
  jor  g06945(.dina(n7178), .dinb(n7171), .dout(n7179));
  jand g06946(.dina(n7179), .dinb(n7170), .dout(n7180));
  jor  g06947(.dina(n7180), .dinb(n5989), .dout(n7181));
  jand g06948(.dina(n7180), .dinb(n5989), .dout(n7182));
  jxor g06949(.dina(n6611), .dinb(n6357), .dout(n7183));
  jor  g06950(.dina(n7183), .dinb(n7154), .dout(n7184));
  jxor g06951(.dina(n7184), .dinb(n7031), .dout(n7185));
  jnot g06952(.din(n7185), .dout(n7186));
  jor  g06953(.dina(n7186), .dinb(n7182), .dout(n7187));
  jand g06954(.dina(n7187), .dinb(n7181), .dout(n7188));
  jor  g06955(.dina(n7188), .dinb(n5606), .dout(n7189));
  jand g06956(.dina(n7188), .dinb(n5606), .dout(n7190));
  jxor g06957(.dina(n6762), .dinb(n5989), .dout(n7191));
  jor  g06958(.dina(n7191), .dinb(n7154), .dout(n7192));
  jxor g06959(.dina(n7192), .dinb(n6772), .dout(n7193));
  jor  g06960(.dina(n7193), .dinb(n7190), .dout(n7194));
  jand g06961(.dina(n7194), .dinb(n7189), .dout(n7195));
  jor  g06962(.dina(n7195), .dinb(n5259), .dout(n7196));
  jand g06963(.dina(n7195), .dinb(n5259), .dout(n7197));
  jxor g06964(.dina(n6774), .dinb(n5606), .dout(n7198));
  jor  g06965(.dina(n7198), .dinb(n7154), .dout(n7199));
  jxor g06966(.dina(n7199), .dinb(n7038), .dout(n7200));
  jnot g06967(.din(n7200), .dout(n7201));
  jor  g06968(.dina(n7201), .dinb(n7197), .dout(n7202));
  jand g06969(.dina(n7202), .dinb(n7196), .dout(n7203));
  jor  g06970(.dina(n7203), .dinb(n4902), .dout(n7204));
  jand g06971(.dina(n7203), .dinb(n4902), .dout(n7205));
  jxor g06972(.dina(n6781), .dinb(n5259), .dout(n7206));
  jor  g06973(.dina(n7206), .dinb(n7154), .dout(n7207));
  jxor g06974(.dina(n7207), .dinb(n7042), .dout(n7208));
  jnot g06975(.din(n7208), .dout(n7209));
  jor  g06976(.dina(n7209), .dinb(n7205), .dout(n7210));
  jand g06977(.dina(n7210), .dinb(n7204), .dout(n7211));
  jor  g06978(.dina(n7211), .dinb(n4582), .dout(n7212));
  jand g06979(.dina(n7211), .dinb(n4582), .dout(n7213));
  jxor g06980(.dina(n6788), .dinb(n4902), .dout(n7214));
  jor  g06981(.dina(n7214), .dinb(n7154), .dout(n7215));
  jxor g06982(.dina(n7215), .dinb(n7046), .dout(n7216));
  jnot g06983(.din(n7216), .dout(n7217));
  jor  g06984(.dina(n7217), .dinb(n7213), .dout(n7218));
  jand g06985(.dina(n7218), .dinb(n7212), .dout(n7219));
  jor  g06986(.dina(n7219), .dinb(n4249), .dout(n7220));
  jand g06987(.dina(n7219), .dinb(n4249), .dout(n7221));
  jxor g06988(.dina(n6795), .dinb(n4582), .dout(n7222));
  jor  g06989(.dina(n7222), .dinb(n7154), .dout(n7223));
  jxor g06990(.dina(n7223), .dinb(n6801), .dout(n7224));
  jor  g06991(.dina(n7224), .dinb(n7221), .dout(n7225));
  jand g06992(.dina(n7225), .dinb(n7220), .dout(n7226));
  jor  g06993(.dina(n7226), .dinb(n3955), .dout(n7227));
  jand g06994(.dina(n7226), .dinb(n3955), .dout(n7228));
  jxor g06995(.dina(n6803), .dinb(n4249), .dout(n7229));
  jor  g06996(.dina(n7229), .dinb(n7154), .dout(n7230));
  jxor g06997(.dina(n7230), .dinb(n7053), .dout(n7231));
  jnot g06998(.din(n7231), .dout(n7232));
  jor  g06999(.dina(n7232), .dinb(n7228), .dout(n7233));
  jand g07000(.dina(n7233), .dinb(n7227), .dout(n7234));
  jor  g07001(.dina(n7234), .dinb(n3642), .dout(n7235));
  jand g07002(.dina(n7234), .dinb(n3642), .dout(n7236));
  jxor g07003(.dina(n6810), .dinb(n3955), .dout(n7237));
  jor  g07004(.dina(n7237), .dinb(n7154), .dout(n7238));
  jxor g07005(.dina(n7238), .dinb(n6816), .dout(n7239));
  jor  g07006(.dina(n7239), .dinb(n7236), .dout(n7240));
  jand g07007(.dina(n7240), .dinb(n7235), .dout(n7241));
  jor  g07008(.dina(n7241), .dinb(n3368), .dout(n7242));
  jand g07009(.dina(n7241), .dinb(n3368), .dout(n7243));
  jxor g07010(.dina(n6818), .dinb(n3642), .dout(n7244));
  jor  g07011(.dina(n7244), .dinb(n7154), .dout(n7245));
  jxor g07012(.dina(n7245), .dinb(n7060), .dout(n7246));
  jnot g07013(.din(n7246), .dout(n7247));
  jor  g07014(.dina(n7247), .dinb(n7243), .dout(n7248));
  jand g07015(.dina(n7248), .dinb(n7242), .dout(n7249));
  jor  g07016(.dina(n7249), .dinb(n3089), .dout(n7250));
  jand g07017(.dina(n7249), .dinb(n3089), .dout(n7251));
  jxor g07018(.dina(n6825), .dinb(n3368), .dout(n7252));
  jor  g07019(.dina(n7252), .dinb(n7154), .dout(n7253));
  jxor g07020(.dina(n7253), .dinb(n6831), .dout(n7254));
  jor  g07021(.dina(n7254), .dinb(n7251), .dout(n7255));
  jand g07022(.dina(n7255), .dinb(n7250), .dout(n7256));
  jor  g07023(.dina(n7256), .dinb(n2833), .dout(n7257));
  jand g07024(.dina(n7256), .dinb(n2833), .dout(n7258));
  jxor g07025(.dina(n6833), .dinb(n3089), .dout(n7259));
  jor  g07026(.dina(n7259), .dinb(n7154), .dout(n7260));
  jxor g07027(.dina(n7260), .dinb(n7067), .dout(n7261));
  jnot g07028(.din(n7261), .dout(n7262));
  jor  g07029(.dina(n7262), .dinb(n7258), .dout(n7263));
  jand g07030(.dina(n7263), .dinb(n7257), .dout(n7264));
  jor  g07031(.dina(n7264), .dinb(n2572), .dout(n7265));
  jand g07032(.dina(n7264), .dinb(n2572), .dout(n7266));
  jxor g07033(.dina(n6840), .dinb(n2833), .dout(n7267));
  jor  g07034(.dina(n7267), .dinb(n7154), .dout(n7268));
  jxor g07035(.dina(n7268), .dinb(n6846), .dout(n7269));
  jor  g07036(.dina(n7269), .dinb(n7266), .dout(n7270));
  jand g07037(.dina(n7270), .dinb(n7265), .dout(n7271));
  jor  g07038(.dina(n7271), .dinb(n2345), .dout(n7272));
  jand g07039(.dina(n7271), .dinb(n2345), .dout(n7273));
  jxor g07040(.dina(n6848), .dinb(n2572), .dout(n7274));
  jor  g07041(.dina(n7274), .dinb(n7154), .dout(n7275));
  jxor g07042(.dina(n7275), .dinb(n7074), .dout(n7276));
  jnot g07043(.din(n7276), .dout(n7277));
  jor  g07044(.dina(n7277), .dinb(n7273), .dout(n7278));
  jand g07045(.dina(n7278), .dinb(n7272), .dout(n7279));
  jor  g07046(.dina(n7279), .dinb(n2108), .dout(n7280));
  jand g07047(.dina(n7279), .dinb(n2108), .dout(n7281));
  jxor g07048(.dina(n6855), .dinb(n2345), .dout(n7282));
  jor  g07049(.dina(n7282), .dinb(n7154), .dout(n7283));
  jxor g07050(.dina(n7283), .dinb(n7078), .dout(n7284));
  jnot g07051(.din(n7284), .dout(n7285));
  jor  g07052(.dina(n7285), .dinb(n7281), .dout(n7286));
  jand g07053(.dina(n7286), .dinb(n7280), .dout(n7287));
  jor  g07054(.dina(n7287), .dinb(n1912), .dout(n7288));
  jand g07055(.dina(n7287), .dinb(n1912), .dout(n7289));
  jxor g07056(.dina(n6862), .dinb(n2108), .dout(n7290));
  jor  g07057(.dina(n7290), .dinb(n7154), .dout(n7291));
  jxor g07058(.dina(n7291), .dinb(n7082), .dout(n7292));
  jnot g07059(.din(n7292), .dout(n7293));
  jor  g07060(.dina(n7293), .dinb(n7289), .dout(n7294));
  jand g07061(.dina(n7294), .dinb(n7288), .dout(n7295));
  jor  g07062(.dina(n7295), .dinb(n1699), .dout(n7296));
  jand g07063(.dina(n7295), .dinb(n1699), .dout(n7297));
  jxor g07064(.dina(n6869), .dinb(n1912), .dout(n7298));
  jor  g07065(.dina(n7298), .dinb(n7154), .dout(n7299));
  jxor g07066(.dina(n7299), .dinb(n6875), .dout(n7300));
  jor  g07067(.dina(n7300), .dinb(n7297), .dout(n7301));
  jand g07068(.dina(n7301), .dinb(n7296), .dout(n7302));
  jor  g07069(.dina(n7302), .dinb(n1516), .dout(n7303));
  jand g07070(.dina(n7302), .dinb(n1516), .dout(n7304));
  jxor g07071(.dina(n6877), .dinb(n1699), .dout(n7305));
  jor  g07072(.dina(n7305), .dinb(n7154), .dout(n7306));
  jxor g07073(.dina(n7306), .dinb(n6883), .dout(n7307));
  jor  g07074(.dina(n7307), .dinb(n7304), .dout(n7308));
  jand g07075(.dina(n7308), .dinb(n7303), .dout(n7309));
  jor  g07076(.dina(n7309), .dinb(n1332), .dout(n7310));
  jand g07077(.dina(n7309), .dinb(n1332), .dout(n7311));
  jxor g07078(.dina(n6885), .dinb(n1516), .dout(n7312));
  jor  g07079(.dina(n7312), .dinb(n7154), .dout(n7313));
  jxor g07080(.dina(n7313), .dinb(n6891), .dout(n7314));
  jor  g07081(.dina(n7314), .dinb(n7311), .dout(n7315));
  jand g07082(.dina(n7315), .dinb(n7310), .dout(n7316));
  jor  g07083(.dina(n7316), .dinb(n1173), .dout(n7317));
  jand g07084(.dina(n7316), .dinb(n1173), .dout(n7318));
  jxor g07085(.dina(n6893), .dinb(n1332), .dout(n7319));
  jor  g07086(.dina(n7319), .dinb(n7154), .dout(n7320));
  jxor g07087(.dina(n7320), .dinb(n7095), .dout(n7321));
  jnot g07088(.din(n7321), .dout(n7322));
  jor  g07089(.dina(n7322), .dinb(n7318), .dout(n7323));
  jand g07090(.dina(n7323), .dinb(n7317), .dout(n7324));
  jor  g07091(.dina(n7324), .dinb(n1008), .dout(n7325));
  jand g07092(.dina(n7324), .dinb(n1008), .dout(n7326));
  jxor g07093(.dina(n6900), .dinb(n1173), .dout(n7327));
  jor  g07094(.dina(n7327), .dinb(n7154), .dout(n7328));
  jxor g07095(.dina(n7328), .dinb(n6906), .dout(n7329));
  jor  g07096(.dina(n7329), .dinb(n7326), .dout(n7330));
  jand g07097(.dina(n7330), .dinb(n7325), .dout(n7331));
  jor  g07098(.dina(n7331), .dinb(n884), .dout(n7332));
  jand g07099(.dina(n7331), .dinb(n884), .dout(n7333));
  jxor g07100(.dina(n6908), .dinb(n1008), .dout(n7334));
  jor  g07101(.dina(n7334), .dinb(n7154), .dout(n7335));
  jxor g07102(.dina(n7335), .dinb(n7102), .dout(n7336));
  jnot g07103(.din(n7336), .dout(n7337));
  jor  g07104(.dina(n7337), .dinb(n7333), .dout(n7338));
  jand g07105(.dina(n7338), .dinb(n7332), .dout(n7339));
  jor  g07106(.dina(n7339), .dinb(n743), .dout(n7340));
  jand g07107(.dina(n7339), .dinb(n743), .dout(n7341));
  jxor g07108(.dina(n6915), .dinb(n884), .dout(n7342));
  jor  g07109(.dina(n7342), .dinb(n7154), .dout(n7343));
  jxor g07110(.dina(n7343), .dinb(n6921), .dout(n7344));
  jor  g07111(.dina(n7344), .dinb(n7341), .dout(n7345));
  jand g07112(.dina(n7345), .dinb(n7340), .dout(n7346));
  jor  g07113(.dina(n7346), .dinb(n635), .dout(n7347));
  jand g07114(.dina(n7346), .dinb(n635), .dout(n7348));
  jxor g07115(.dina(n6923), .dinb(n743), .dout(n7349));
  jor  g07116(.dina(n7349), .dinb(n7154), .dout(n7350));
  jxor g07117(.dina(n7350), .dinb(n7109), .dout(n7351));
  jnot g07118(.din(n7351), .dout(n7352));
  jor  g07119(.dina(n7352), .dinb(n7348), .dout(n7353));
  jand g07120(.dina(n7353), .dinb(n7347), .dout(n7354));
  jor  g07121(.dina(n7354), .dinb(n515), .dout(n7355));
  jand g07122(.dina(n7354), .dinb(n515), .dout(n7356));
  jxor g07123(.dina(n6930), .dinb(n635), .dout(n7357));
  jor  g07124(.dina(n7357), .dinb(n7154), .dout(n7358));
  jxor g07125(.dina(n7358), .dinb(n7113), .dout(n7359));
  jnot g07126(.din(n7359), .dout(n7360));
  jor  g07127(.dina(n7360), .dinb(n7356), .dout(n7361));
  jand g07128(.dina(n7361), .dinb(n7355), .dout(n7362));
  jor  g07129(.dina(n7362), .dinb(n443), .dout(n7363));
  jand g07130(.dina(n7362), .dinb(n443), .dout(n7364));
  jxor g07131(.dina(n6937), .dinb(n515), .dout(n7365));
  jor  g07132(.dina(n7365), .dinb(n7154), .dout(n7366));
  jxor g07133(.dina(n7366), .dinb(n6943), .dout(n7367));
  jor  g07134(.dina(n7367), .dinb(n7364), .dout(n7368));
  jand g07135(.dina(n7368), .dinb(n7363), .dout(n7369));
  jor  g07136(.dina(n7369), .dinb(n352), .dout(n7370));
  jand g07137(.dina(n7369), .dinb(n352), .dout(n7371));
  jxor g07138(.dina(n6945), .dinb(n443), .dout(n7372));
  jor  g07139(.dina(n7372), .dinb(n7154), .dout(n7373));
  jxor g07140(.dina(n7373), .dinb(n6951), .dout(n7374));
  jor  g07141(.dina(n7374), .dinb(n7371), .dout(n7375));
  jand g07142(.dina(n7375), .dinb(n7370), .dout(n7376));
  jor  g07143(.dina(n7376), .dinb(n294), .dout(n7377));
  jand g07144(.dina(n7376), .dinb(n294), .dout(n7378));
  jxor g07145(.dina(n6953), .dinb(n352), .dout(n7379));
  jor  g07146(.dina(n7379), .dinb(n7154), .dout(n7380));
  jxor g07147(.dina(n7380), .dinb(n6959), .dout(n7381));
  jor  g07148(.dina(n7381), .dinb(n7378), .dout(n7382));
  jand g07149(.dina(n7382), .dinb(n7377), .dout(n7383));
  jor  g07150(.dina(n7383), .dinb(n239), .dout(n7384));
  jand g07151(.dina(n7383), .dinb(n239), .dout(n7385));
  jxor g07152(.dina(n6961), .dinb(n294), .dout(n7386));
  jor  g07153(.dina(n7386), .dinb(n7154), .dout(n7387));
  jxor g07154(.dina(n7387), .dinb(n7126), .dout(n7388));
  jnot g07155(.din(n7388), .dout(n7389));
  jor  g07156(.dina(n7389), .dinb(n7385), .dout(n7390));
  jand g07157(.dina(n7390), .dinb(n7384), .dout(n7391));
  jor  g07158(.dina(n7391), .dinb(n221), .dout(n7392));
  jand g07159(.dina(n7391), .dinb(n221), .dout(n7393));
  jxor g07160(.dina(n6968), .dinb(n239), .dout(n7394));
  jor  g07161(.dina(n7394), .dinb(n7154), .dout(n7395));
  jxor g07162(.dina(n7395), .dinb(n7130), .dout(n7396));
  jnot g07163(.din(n7396), .dout(n7397));
  jor  g07164(.dina(n7397), .dinb(n7393), .dout(n7398));
  jand g07165(.dina(n7398), .dinb(n7392), .dout(n7399));
  jxor g07166(.dina(n6975), .dinb(n221), .dout(n7400));
  jor  g07167(.dina(n7400), .dinb(n7154), .dout(n7401));
  jxor g07168(.dina(n7401), .dinb(n6981), .dout(n7402));
  jor  g07169(.dina(n7402), .dinb(n7399), .dout(n7403));
  jor  g07170(.dina(n7403), .dinb(n6989), .dout(n7404));
  jor  g07171(.dina(n7404), .dinb(n7146), .dout(n7405));
  jand g07172(.dina(n7405), .dinb(n218), .dout(n7406));
  jand g07173(.dina(n7154), .dinb(n6986), .dout(n7407));
  jand g07174(.dina(n7402), .dinb(n7399), .dout(n7408));
  jor  g07175(.dina(n7408), .dinb(n7407), .dout(n7409));
  jand g07176(.dina(n7153), .dinb(n7135), .dout(n7410));
  jnot g07177(.din(n7410), .dout(n7411));
  jand g07178(.dina(n7136), .dinb(asqrt[63] ), .dout(n7412));
  jand g07179(.dina(n7412), .dinb(n6988), .dout(n7413));
  jand g07180(.dina(n7413), .dinb(n7411), .dout(n7414));
  jor  g07181(.dina(n7414), .dinb(n7409), .dout(n7415));
  jor  g07182(.dina(n7415), .dinb(n7406), .dout(asqrt[30] ));
  jxor g07183(.dina(n7391), .dinb(n221), .dout(n7417));
  jand g07184(.dina(n7417), .dinb(asqrt[30] ), .dout(n7418));
  jxor g07185(.dina(n7418), .dinb(n7396), .dout(n7419));
  jand g07186(.dina(asqrt[30] ), .dinb(a[60] ), .dout(n7420));
  jnot g07187(.din(a[58] ), .dout(n7421));
  jnot g07188(.din(a[59] ), .dout(n7422));
  jand g07189(.dina(n7422), .dinb(n7421), .dout(n7423));
  jand g07190(.dina(n7423), .dinb(n7156), .dout(n7424));
  jor  g07191(.dina(n7424), .dinb(n7420), .dout(n7425));
  jand g07192(.dina(n7425), .dinb(asqrt[31] ), .dout(n7426));
  jor  g07193(.dina(n7425), .dinb(asqrt[31] ), .dout(n7427));
  jand g07194(.dina(asqrt[30] ), .dinb(n7156), .dout(n7428));
  jor  g07195(.dina(n7428), .dinb(n7157), .dout(n7429));
  jnot g07196(.din(n7158), .dout(n7430));
  jnot g07197(.din(n7146), .dout(n7431));
  jnot g07198(.din(n7392), .dout(n7432));
  jnot g07199(.din(n7384), .dout(n7433));
  jnot g07200(.din(n7377), .dout(n7434));
  jnot g07201(.din(n7370), .dout(n7435));
  jnot g07202(.din(n7363), .dout(n7436));
  jnot g07203(.din(n7355), .dout(n7437));
  jnot g07204(.din(n7347), .dout(n7438));
  jnot g07205(.din(n7340), .dout(n7439));
  jnot g07206(.din(n7332), .dout(n7440));
  jnot g07207(.din(n7325), .dout(n7441));
  jnot g07208(.din(n7317), .dout(n7442));
  jnot g07209(.din(n7310), .dout(n7443));
  jnot g07210(.din(n7303), .dout(n7444));
  jnot g07211(.din(n7296), .dout(n7445));
  jnot g07212(.din(n7288), .dout(n7446));
  jnot g07213(.din(n7280), .dout(n7447));
  jnot g07214(.din(n7272), .dout(n7448));
  jnot g07215(.din(n7265), .dout(n7449));
  jnot g07216(.din(n7257), .dout(n7450));
  jnot g07217(.din(n7250), .dout(n7451));
  jnot g07218(.din(n7242), .dout(n7452));
  jnot g07219(.din(n7235), .dout(n7453));
  jnot g07220(.din(n7227), .dout(n7454));
  jnot g07221(.din(n7220), .dout(n7455));
  jnot g07222(.din(n7212), .dout(n7456));
  jnot g07223(.din(n7204), .dout(n7457));
  jnot g07224(.din(n7196), .dout(n7458));
  jnot g07225(.din(n7189), .dout(n7459));
  jnot g07226(.din(n7181), .dout(n7460));
  jnot g07227(.din(n7170), .dout(n7461));
  jnot g07228(.din(n7162), .dout(n7462));
  jand g07229(.dina(asqrt[31] ), .dinb(n6606), .dout(n7463));
  jor  g07230(.dina(n7463), .dinb(n6607), .dout(n7464));
  jand g07231(.dina(n7464), .dinb(n7173), .dout(n7465));
  jand g07232(.dina(asqrt[31] ), .dinb(a[62] ), .dout(n7466));
  jor  g07233(.dina(n7159), .dinb(n7466), .dout(n7467));
  jor  g07234(.dina(n7467), .dinb(asqrt[32] ), .dout(n7468));
  jand g07235(.dina(n7468), .dinb(n7465), .dout(n7469));
  jor  g07236(.dina(n7469), .dinb(n7462), .dout(n7470));
  jor  g07237(.dina(n7470), .dinb(asqrt[33] ), .dout(n7471));
  jnot g07238(.din(n7178), .dout(n7472));
  jand g07239(.dina(n7472), .dinb(n7471), .dout(n7473));
  jor  g07240(.dina(n7473), .dinb(n7461), .dout(n7474));
  jor  g07241(.dina(n7474), .dinb(asqrt[34] ), .dout(n7475));
  jand g07242(.dina(n7185), .dinb(n7475), .dout(n7476));
  jor  g07243(.dina(n7476), .dinb(n7460), .dout(n7477));
  jor  g07244(.dina(n7477), .dinb(asqrt[35] ), .dout(n7478));
  jnot g07245(.din(n7193), .dout(n7479));
  jand g07246(.dina(n7479), .dinb(n7478), .dout(n7480));
  jor  g07247(.dina(n7480), .dinb(n7459), .dout(n7481));
  jor  g07248(.dina(n7481), .dinb(asqrt[36] ), .dout(n7482));
  jand g07249(.dina(n7200), .dinb(n7482), .dout(n7483));
  jor  g07250(.dina(n7483), .dinb(n7458), .dout(n7484));
  jor  g07251(.dina(n7484), .dinb(asqrt[37] ), .dout(n7485));
  jand g07252(.dina(n7208), .dinb(n7485), .dout(n7486));
  jor  g07253(.dina(n7486), .dinb(n7457), .dout(n7487));
  jor  g07254(.dina(n7487), .dinb(asqrt[38] ), .dout(n7488));
  jand g07255(.dina(n7216), .dinb(n7488), .dout(n7489));
  jor  g07256(.dina(n7489), .dinb(n7456), .dout(n7490));
  jor  g07257(.dina(n7490), .dinb(asqrt[39] ), .dout(n7491));
  jnot g07258(.din(n7224), .dout(n7492));
  jand g07259(.dina(n7492), .dinb(n7491), .dout(n7493));
  jor  g07260(.dina(n7493), .dinb(n7455), .dout(n7494));
  jor  g07261(.dina(n7494), .dinb(asqrt[40] ), .dout(n7495));
  jand g07262(.dina(n7231), .dinb(n7495), .dout(n7496));
  jor  g07263(.dina(n7496), .dinb(n7454), .dout(n7497));
  jor  g07264(.dina(n7497), .dinb(asqrt[41] ), .dout(n7498));
  jnot g07265(.din(n7239), .dout(n7499));
  jand g07266(.dina(n7499), .dinb(n7498), .dout(n7500));
  jor  g07267(.dina(n7500), .dinb(n7453), .dout(n7501));
  jor  g07268(.dina(n7501), .dinb(asqrt[42] ), .dout(n7502));
  jand g07269(.dina(n7246), .dinb(n7502), .dout(n7503));
  jor  g07270(.dina(n7503), .dinb(n7452), .dout(n7504));
  jor  g07271(.dina(n7504), .dinb(asqrt[43] ), .dout(n7505));
  jnot g07272(.din(n7254), .dout(n7506));
  jand g07273(.dina(n7506), .dinb(n7505), .dout(n7507));
  jor  g07274(.dina(n7507), .dinb(n7451), .dout(n7508));
  jor  g07275(.dina(n7508), .dinb(asqrt[44] ), .dout(n7509));
  jand g07276(.dina(n7261), .dinb(n7509), .dout(n7510));
  jor  g07277(.dina(n7510), .dinb(n7450), .dout(n7511));
  jor  g07278(.dina(n7511), .dinb(asqrt[45] ), .dout(n7512));
  jnot g07279(.din(n7269), .dout(n7513));
  jand g07280(.dina(n7513), .dinb(n7512), .dout(n7514));
  jor  g07281(.dina(n7514), .dinb(n7449), .dout(n7515));
  jor  g07282(.dina(n7515), .dinb(asqrt[46] ), .dout(n7516));
  jand g07283(.dina(n7276), .dinb(n7516), .dout(n7517));
  jor  g07284(.dina(n7517), .dinb(n7448), .dout(n7518));
  jor  g07285(.dina(n7518), .dinb(asqrt[47] ), .dout(n7519));
  jand g07286(.dina(n7284), .dinb(n7519), .dout(n7520));
  jor  g07287(.dina(n7520), .dinb(n7447), .dout(n7521));
  jor  g07288(.dina(n7521), .dinb(asqrt[48] ), .dout(n7522));
  jand g07289(.dina(n7292), .dinb(n7522), .dout(n7523));
  jor  g07290(.dina(n7523), .dinb(n7446), .dout(n7524));
  jor  g07291(.dina(n7524), .dinb(asqrt[49] ), .dout(n7525));
  jnot g07292(.din(n7300), .dout(n7526));
  jand g07293(.dina(n7526), .dinb(n7525), .dout(n7527));
  jor  g07294(.dina(n7527), .dinb(n7445), .dout(n7528));
  jor  g07295(.dina(n7528), .dinb(asqrt[50] ), .dout(n7529));
  jnot g07296(.din(n7307), .dout(n7530));
  jand g07297(.dina(n7530), .dinb(n7529), .dout(n7531));
  jor  g07298(.dina(n7531), .dinb(n7444), .dout(n7532));
  jor  g07299(.dina(n7532), .dinb(asqrt[51] ), .dout(n7533));
  jnot g07300(.din(n7314), .dout(n7534));
  jand g07301(.dina(n7534), .dinb(n7533), .dout(n7535));
  jor  g07302(.dina(n7535), .dinb(n7443), .dout(n7536));
  jor  g07303(.dina(n7536), .dinb(asqrt[52] ), .dout(n7537));
  jand g07304(.dina(n7321), .dinb(n7537), .dout(n7538));
  jor  g07305(.dina(n7538), .dinb(n7442), .dout(n7539));
  jor  g07306(.dina(n7539), .dinb(asqrt[53] ), .dout(n7540));
  jnot g07307(.din(n7329), .dout(n7541));
  jand g07308(.dina(n7541), .dinb(n7540), .dout(n7542));
  jor  g07309(.dina(n7542), .dinb(n7441), .dout(n7543));
  jor  g07310(.dina(n7543), .dinb(asqrt[54] ), .dout(n7544));
  jand g07311(.dina(n7336), .dinb(n7544), .dout(n7545));
  jor  g07312(.dina(n7545), .dinb(n7440), .dout(n7546));
  jor  g07313(.dina(n7546), .dinb(asqrt[55] ), .dout(n7547));
  jnot g07314(.din(n7344), .dout(n7548));
  jand g07315(.dina(n7548), .dinb(n7547), .dout(n7549));
  jor  g07316(.dina(n7549), .dinb(n7439), .dout(n7550));
  jor  g07317(.dina(n7550), .dinb(asqrt[56] ), .dout(n7551));
  jand g07318(.dina(n7351), .dinb(n7551), .dout(n7552));
  jor  g07319(.dina(n7552), .dinb(n7438), .dout(n7553));
  jor  g07320(.dina(n7553), .dinb(asqrt[57] ), .dout(n7554));
  jand g07321(.dina(n7359), .dinb(n7554), .dout(n7555));
  jor  g07322(.dina(n7555), .dinb(n7437), .dout(n7556));
  jor  g07323(.dina(n7556), .dinb(asqrt[58] ), .dout(n7557));
  jnot g07324(.din(n7367), .dout(n7558));
  jand g07325(.dina(n7558), .dinb(n7557), .dout(n7559));
  jor  g07326(.dina(n7559), .dinb(n7436), .dout(n7560));
  jor  g07327(.dina(n7560), .dinb(asqrt[59] ), .dout(n7561));
  jnot g07328(.din(n7374), .dout(n7562));
  jand g07329(.dina(n7562), .dinb(n7561), .dout(n7563));
  jor  g07330(.dina(n7563), .dinb(n7435), .dout(n7564));
  jor  g07331(.dina(n7564), .dinb(asqrt[60] ), .dout(n7565));
  jnot g07332(.din(n7381), .dout(n7566));
  jand g07333(.dina(n7566), .dinb(n7565), .dout(n7567));
  jor  g07334(.dina(n7567), .dinb(n7434), .dout(n7568));
  jor  g07335(.dina(n7568), .dinb(asqrt[61] ), .dout(n7569));
  jand g07336(.dina(n7388), .dinb(n7569), .dout(n7570));
  jor  g07337(.dina(n7570), .dinb(n7433), .dout(n7571));
  jor  g07338(.dina(n7571), .dinb(asqrt[62] ), .dout(n7572));
  jand g07339(.dina(n7396), .dinb(n7572), .dout(n7573));
  jor  g07340(.dina(n7573), .dinb(n7432), .dout(n7574));
  jnot g07341(.din(n7402), .dout(n7575));
  jand g07342(.dina(n7575), .dinb(n7574), .dout(n7576));
  jand g07343(.dina(n7576), .dinb(n6988), .dout(n7577));
  jand g07344(.dina(n7577), .dinb(n7431), .dout(n7578));
  jor  g07345(.dina(n7578), .dinb(asqrt[63] ), .dout(n7579));
  jnot g07346(.din(n7415), .dout(n7580));
  jand g07347(.dina(n7580), .dinb(n7579), .dout(n7581));
  jor  g07348(.dina(n7581), .dinb(n7430), .dout(n7582));
  jand g07349(.dina(n7582), .dinb(n7429), .dout(n7583));
  jand g07350(.dina(n7583), .dinb(n7427), .dout(n7584));
  jor  g07351(.dina(n7584), .dinb(n7426), .dout(n7585));
  jand g07352(.dina(n7585), .dinb(asqrt[32] ), .dout(n7586));
  jor  g07353(.dina(n7585), .dinb(asqrt[32] ), .dout(n7587));
  jor  g07354(.dina(n7413), .dinb(n7408), .dout(n7588));
  jor  g07355(.dina(n7588), .dinb(n7406), .dout(n7589));
  jor  g07356(.dina(n7589), .dinb(n7154), .dout(n7590));
  jand g07357(.dina(n7590), .dinb(n7582), .dout(n7591));
  jxor g07358(.dina(n7591), .dinb(n6606), .dout(n7592));
  jnot g07359(.din(n7592), .dout(n7593));
  jand g07360(.dina(n7593), .dinb(n7587), .dout(n7594));
  jor  g07361(.dina(n7594), .dinb(n7586), .dout(n7595));
  jand g07362(.dina(n7595), .dinb(asqrt[33] ), .dout(n7596));
  jxor g07363(.dina(n7161), .dinb(n6758), .dout(n7597));
  jand g07364(.dina(n7597), .dinb(asqrt[30] ), .dout(n7598));
  jxor g07365(.dina(n7598), .dinb(n7465), .dout(n7599));
  jor  g07366(.dina(n7595), .dinb(asqrt[33] ), .dout(n7600));
  jand g07367(.dina(n7600), .dinb(n7599), .dout(n7601));
  jor  g07368(.dina(n7601), .dinb(n7596), .dout(n7602));
  jand g07369(.dina(n7602), .dinb(asqrt[34] ), .dout(n7603));
  jor  g07370(.dina(n7602), .dinb(asqrt[34] ), .dout(n7604));
  jxor g07371(.dina(n7169), .dinb(n6357), .dout(n7605));
  jand g07372(.dina(n7605), .dinb(asqrt[30] ), .dout(n7606));
  jxor g07373(.dina(n7606), .dinb(n7178), .dout(n7607));
  jnot g07374(.din(n7607), .dout(n7608));
  jand g07375(.dina(n7608), .dinb(n7604), .dout(n7609));
  jor  g07376(.dina(n7609), .dinb(n7603), .dout(n7610));
  jand g07377(.dina(n7610), .dinb(asqrt[35] ), .dout(n7611));
  jor  g07378(.dina(n7610), .dinb(asqrt[35] ), .dout(n7612));
  jxor g07379(.dina(n7180), .dinb(n5989), .dout(n7613));
  jand g07380(.dina(n7613), .dinb(asqrt[30] ), .dout(n7614));
  jxor g07381(.dina(n7614), .dinb(n7185), .dout(n7615));
  jand g07382(.dina(n7615), .dinb(n7612), .dout(n7616));
  jor  g07383(.dina(n7616), .dinb(n7611), .dout(n7617));
  jand g07384(.dina(n7617), .dinb(asqrt[36] ), .dout(n7618));
  jor  g07385(.dina(n7617), .dinb(asqrt[36] ), .dout(n7619));
  jxor g07386(.dina(n7188), .dinb(n5606), .dout(n7620));
  jand g07387(.dina(n7620), .dinb(asqrt[30] ), .dout(n7621));
  jxor g07388(.dina(n7621), .dinb(n7193), .dout(n7622));
  jnot g07389(.din(n7622), .dout(n7623));
  jand g07390(.dina(n7623), .dinb(n7619), .dout(n7624));
  jor  g07391(.dina(n7624), .dinb(n7618), .dout(n7625));
  jand g07392(.dina(n7625), .dinb(asqrt[37] ), .dout(n7626));
  jor  g07393(.dina(n7625), .dinb(asqrt[37] ), .dout(n7627));
  jxor g07394(.dina(n7195), .dinb(n5259), .dout(n7628));
  jand g07395(.dina(n7628), .dinb(asqrt[30] ), .dout(n7629));
  jxor g07396(.dina(n7629), .dinb(n7200), .dout(n7630));
  jand g07397(.dina(n7630), .dinb(n7627), .dout(n7631));
  jor  g07398(.dina(n7631), .dinb(n7626), .dout(n7632));
  jand g07399(.dina(n7632), .dinb(asqrt[38] ), .dout(n7633));
  jor  g07400(.dina(n7632), .dinb(asqrt[38] ), .dout(n7634));
  jxor g07401(.dina(n7203), .dinb(n4902), .dout(n7635));
  jand g07402(.dina(n7635), .dinb(asqrt[30] ), .dout(n7636));
  jxor g07403(.dina(n7636), .dinb(n7208), .dout(n7637));
  jand g07404(.dina(n7637), .dinb(n7634), .dout(n7638));
  jor  g07405(.dina(n7638), .dinb(n7633), .dout(n7639));
  jand g07406(.dina(n7639), .dinb(asqrt[39] ), .dout(n7640));
  jor  g07407(.dina(n7639), .dinb(asqrt[39] ), .dout(n7641));
  jxor g07408(.dina(n7211), .dinb(n4582), .dout(n7642));
  jand g07409(.dina(n7642), .dinb(asqrt[30] ), .dout(n7643));
  jxor g07410(.dina(n7643), .dinb(n7216), .dout(n7644));
  jand g07411(.dina(n7644), .dinb(n7641), .dout(n7645));
  jor  g07412(.dina(n7645), .dinb(n7640), .dout(n7646));
  jand g07413(.dina(n7646), .dinb(asqrt[40] ), .dout(n7647));
  jor  g07414(.dina(n7646), .dinb(asqrt[40] ), .dout(n7648));
  jxor g07415(.dina(n7219), .dinb(n4249), .dout(n7649));
  jand g07416(.dina(n7649), .dinb(asqrt[30] ), .dout(n7650));
  jxor g07417(.dina(n7650), .dinb(n7224), .dout(n7651));
  jnot g07418(.din(n7651), .dout(n7652));
  jand g07419(.dina(n7652), .dinb(n7648), .dout(n7653));
  jor  g07420(.dina(n7653), .dinb(n7647), .dout(n7654));
  jand g07421(.dina(n7654), .dinb(asqrt[41] ), .dout(n7655));
  jor  g07422(.dina(n7654), .dinb(asqrt[41] ), .dout(n7656));
  jxor g07423(.dina(n7226), .dinb(n3955), .dout(n7657));
  jand g07424(.dina(n7657), .dinb(asqrt[30] ), .dout(n7658));
  jxor g07425(.dina(n7658), .dinb(n7231), .dout(n7659));
  jand g07426(.dina(n7659), .dinb(n7656), .dout(n7660));
  jor  g07427(.dina(n7660), .dinb(n7655), .dout(n7661));
  jand g07428(.dina(n7661), .dinb(asqrt[42] ), .dout(n7662));
  jor  g07429(.dina(n7661), .dinb(asqrt[42] ), .dout(n7663));
  jxor g07430(.dina(n7234), .dinb(n3642), .dout(n7664));
  jand g07431(.dina(n7664), .dinb(asqrt[30] ), .dout(n7665));
  jxor g07432(.dina(n7665), .dinb(n7239), .dout(n7666));
  jnot g07433(.din(n7666), .dout(n7667));
  jand g07434(.dina(n7667), .dinb(n7663), .dout(n7668));
  jor  g07435(.dina(n7668), .dinb(n7662), .dout(n7669));
  jand g07436(.dina(n7669), .dinb(asqrt[43] ), .dout(n7670));
  jor  g07437(.dina(n7669), .dinb(asqrt[43] ), .dout(n7671));
  jxor g07438(.dina(n7241), .dinb(n3368), .dout(n7672));
  jand g07439(.dina(n7672), .dinb(asqrt[30] ), .dout(n7673));
  jxor g07440(.dina(n7673), .dinb(n7246), .dout(n7674));
  jand g07441(.dina(n7674), .dinb(n7671), .dout(n7675));
  jor  g07442(.dina(n7675), .dinb(n7670), .dout(n7676));
  jand g07443(.dina(n7676), .dinb(asqrt[44] ), .dout(n7677));
  jor  g07444(.dina(n7676), .dinb(asqrt[44] ), .dout(n7678));
  jxor g07445(.dina(n7249), .dinb(n3089), .dout(n7679));
  jand g07446(.dina(n7679), .dinb(asqrt[30] ), .dout(n7680));
  jxor g07447(.dina(n7680), .dinb(n7254), .dout(n7681));
  jnot g07448(.din(n7681), .dout(n7682));
  jand g07449(.dina(n7682), .dinb(n7678), .dout(n7683));
  jor  g07450(.dina(n7683), .dinb(n7677), .dout(n7684));
  jand g07451(.dina(n7684), .dinb(asqrt[45] ), .dout(n7685));
  jor  g07452(.dina(n7684), .dinb(asqrt[45] ), .dout(n7686));
  jxor g07453(.dina(n7256), .dinb(n2833), .dout(n7687));
  jand g07454(.dina(n7687), .dinb(asqrt[30] ), .dout(n7688));
  jxor g07455(.dina(n7688), .dinb(n7261), .dout(n7689));
  jand g07456(.dina(n7689), .dinb(n7686), .dout(n7690));
  jor  g07457(.dina(n7690), .dinb(n7685), .dout(n7691));
  jand g07458(.dina(n7691), .dinb(asqrt[46] ), .dout(n7692));
  jor  g07459(.dina(n7691), .dinb(asqrt[46] ), .dout(n7693));
  jxor g07460(.dina(n7264), .dinb(n2572), .dout(n7694));
  jand g07461(.dina(n7694), .dinb(asqrt[30] ), .dout(n7695));
  jxor g07462(.dina(n7695), .dinb(n7269), .dout(n7696));
  jnot g07463(.din(n7696), .dout(n7697));
  jand g07464(.dina(n7697), .dinb(n7693), .dout(n7698));
  jor  g07465(.dina(n7698), .dinb(n7692), .dout(n7699));
  jand g07466(.dina(n7699), .dinb(asqrt[47] ), .dout(n7700));
  jor  g07467(.dina(n7699), .dinb(asqrt[47] ), .dout(n7701));
  jxor g07468(.dina(n7271), .dinb(n2345), .dout(n7702));
  jand g07469(.dina(n7702), .dinb(asqrt[30] ), .dout(n7703));
  jxor g07470(.dina(n7703), .dinb(n7276), .dout(n7704));
  jand g07471(.dina(n7704), .dinb(n7701), .dout(n7705));
  jor  g07472(.dina(n7705), .dinb(n7700), .dout(n7706));
  jand g07473(.dina(n7706), .dinb(asqrt[48] ), .dout(n7707));
  jor  g07474(.dina(n7706), .dinb(asqrt[48] ), .dout(n7708));
  jxor g07475(.dina(n7279), .dinb(n2108), .dout(n7709));
  jand g07476(.dina(n7709), .dinb(asqrt[30] ), .dout(n7710));
  jxor g07477(.dina(n7710), .dinb(n7284), .dout(n7711));
  jand g07478(.dina(n7711), .dinb(n7708), .dout(n7712));
  jor  g07479(.dina(n7712), .dinb(n7707), .dout(n7713));
  jand g07480(.dina(n7713), .dinb(asqrt[49] ), .dout(n7714));
  jor  g07481(.dina(n7713), .dinb(asqrt[49] ), .dout(n7715));
  jxor g07482(.dina(n7287), .dinb(n1912), .dout(n7716));
  jand g07483(.dina(n7716), .dinb(asqrt[30] ), .dout(n7717));
  jxor g07484(.dina(n7717), .dinb(n7292), .dout(n7718));
  jand g07485(.dina(n7718), .dinb(n7715), .dout(n7719));
  jor  g07486(.dina(n7719), .dinb(n7714), .dout(n7720));
  jand g07487(.dina(n7720), .dinb(asqrt[50] ), .dout(n7721));
  jor  g07488(.dina(n7720), .dinb(asqrt[50] ), .dout(n7722));
  jxor g07489(.dina(n7295), .dinb(n1699), .dout(n7723));
  jand g07490(.dina(n7723), .dinb(asqrt[30] ), .dout(n7724));
  jxor g07491(.dina(n7724), .dinb(n7300), .dout(n7725));
  jnot g07492(.din(n7725), .dout(n7726));
  jand g07493(.dina(n7726), .dinb(n7722), .dout(n7727));
  jor  g07494(.dina(n7727), .dinb(n7721), .dout(n7728));
  jand g07495(.dina(n7728), .dinb(asqrt[51] ), .dout(n7729));
  jor  g07496(.dina(n7728), .dinb(asqrt[51] ), .dout(n7730));
  jxor g07497(.dina(n7302), .dinb(n1516), .dout(n7731));
  jand g07498(.dina(n7731), .dinb(asqrt[30] ), .dout(n7732));
  jxor g07499(.dina(n7732), .dinb(n7307), .dout(n7733));
  jnot g07500(.din(n7733), .dout(n7734));
  jand g07501(.dina(n7734), .dinb(n7730), .dout(n7735));
  jor  g07502(.dina(n7735), .dinb(n7729), .dout(n7736));
  jand g07503(.dina(n7736), .dinb(asqrt[52] ), .dout(n7737));
  jor  g07504(.dina(n7736), .dinb(asqrt[52] ), .dout(n7738));
  jxor g07505(.dina(n7309), .dinb(n1332), .dout(n7739));
  jand g07506(.dina(n7739), .dinb(asqrt[30] ), .dout(n7740));
  jxor g07507(.dina(n7740), .dinb(n7314), .dout(n7741));
  jnot g07508(.din(n7741), .dout(n7742));
  jand g07509(.dina(n7742), .dinb(n7738), .dout(n7743));
  jor  g07510(.dina(n7743), .dinb(n7737), .dout(n7744));
  jand g07511(.dina(n7744), .dinb(asqrt[53] ), .dout(n7745));
  jor  g07512(.dina(n7744), .dinb(asqrt[53] ), .dout(n7746));
  jxor g07513(.dina(n7316), .dinb(n1173), .dout(n7747));
  jand g07514(.dina(n7747), .dinb(asqrt[30] ), .dout(n7748));
  jxor g07515(.dina(n7748), .dinb(n7321), .dout(n7749));
  jand g07516(.dina(n7749), .dinb(n7746), .dout(n7750));
  jor  g07517(.dina(n7750), .dinb(n7745), .dout(n7751));
  jand g07518(.dina(n7751), .dinb(asqrt[54] ), .dout(n7752));
  jor  g07519(.dina(n7751), .dinb(asqrt[54] ), .dout(n7753));
  jxor g07520(.dina(n7324), .dinb(n1008), .dout(n7754));
  jand g07521(.dina(n7754), .dinb(asqrt[30] ), .dout(n7755));
  jxor g07522(.dina(n7755), .dinb(n7329), .dout(n7756));
  jnot g07523(.din(n7756), .dout(n7757));
  jand g07524(.dina(n7757), .dinb(n7753), .dout(n7758));
  jor  g07525(.dina(n7758), .dinb(n7752), .dout(n7759));
  jand g07526(.dina(n7759), .dinb(asqrt[55] ), .dout(n7760));
  jor  g07527(.dina(n7759), .dinb(asqrt[55] ), .dout(n7761));
  jxor g07528(.dina(n7331), .dinb(n884), .dout(n7762));
  jand g07529(.dina(n7762), .dinb(asqrt[30] ), .dout(n7763));
  jxor g07530(.dina(n7763), .dinb(n7336), .dout(n7764));
  jand g07531(.dina(n7764), .dinb(n7761), .dout(n7765));
  jor  g07532(.dina(n7765), .dinb(n7760), .dout(n7766));
  jand g07533(.dina(n7766), .dinb(asqrt[56] ), .dout(n7767));
  jor  g07534(.dina(n7766), .dinb(asqrt[56] ), .dout(n7768));
  jxor g07535(.dina(n7339), .dinb(n743), .dout(n7769));
  jand g07536(.dina(n7769), .dinb(asqrt[30] ), .dout(n7770));
  jxor g07537(.dina(n7770), .dinb(n7344), .dout(n7771));
  jnot g07538(.din(n7771), .dout(n7772));
  jand g07539(.dina(n7772), .dinb(n7768), .dout(n7773));
  jor  g07540(.dina(n7773), .dinb(n7767), .dout(n7774));
  jand g07541(.dina(n7774), .dinb(asqrt[57] ), .dout(n7775));
  jor  g07542(.dina(n7774), .dinb(asqrt[57] ), .dout(n7776));
  jxor g07543(.dina(n7346), .dinb(n635), .dout(n7777));
  jand g07544(.dina(n7777), .dinb(asqrt[30] ), .dout(n7778));
  jxor g07545(.dina(n7778), .dinb(n7351), .dout(n7779));
  jand g07546(.dina(n7779), .dinb(n7776), .dout(n7780));
  jor  g07547(.dina(n7780), .dinb(n7775), .dout(n7781));
  jand g07548(.dina(n7781), .dinb(asqrt[58] ), .dout(n7782));
  jor  g07549(.dina(n7781), .dinb(asqrt[58] ), .dout(n7783));
  jxor g07550(.dina(n7354), .dinb(n515), .dout(n7784));
  jand g07551(.dina(n7784), .dinb(asqrt[30] ), .dout(n7785));
  jxor g07552(.dina(n7785), .dinb(n7359), .dout(n7786));
  jand g07553(.dina(n7786), .dinb(n7783), .dout(n7787));
  jor  g07554(.dina(n7787), .dinb(n7782), .dout(n7788));
  jand g07555(.dina(n7788), .dinb(asqrt[59] ), .dout(n7789));
  jor  g07556(.dina(n7788), .dinb(asqrt[59] ), .dout(n7790));
  jxor g07557(.dina(n7362), .dinb(n443), .dout(n7791));
  jand g07558(.dina(n7791), .dinb(asqrt[30] ), .dout(n7792));
  jxor g07559(.dina(n7792), .dinb(n7367), .dout(n7793));
  jnot g07560(.din(n7793), .dout(n7794));
  jand g07561(.dina(n7794), .dinb(n7790), .dout(n7795));
  jor  g07562(.dina(n7795), .dinb(n7789), .dout(n7796));
  jand g07563(.dina(n7796), .dinb(asqrt[60] ), .dout(n7797));
  jor  g07564(.dina(n7796), .dinb(asqrt[60] ), .dout(n7798));
  jxor g07565(.dina(n7369), .dinb(n352), .dout(n7799));
  jand g07566(.dina(n7799), .dinb(asqrt[30] ), .dout(n7800));
  jxor g07567(.dina(n7800), .dinb(n7374), .dout(n7801));
  jnot g07568(.din(n7801), .dout(n7802));
  jand g07569(.dina(n7802), .dinb(n7798), .dout(n7803));
  jor  g07570(.dina(n7803), .dinb(n7797), .dout(n7804));
  jand g07571(.dina(n7804), .dinb(asqrt[61] ), .dout(n7805));
  jor  g07572(.dina(n7804), .dinb(asqrt[61] ), .dout(n7806));
  jxor g07573(.dina(n7376), .dinb(n294), .dout(n7807));
  jand g07574(.dina(n7807), .dinb(asqrt[30] ), .dout(n7808));
  jxor g07575(.dina(n7808), .dinb(n7381), .dout(n7809));
  jnot g07576(.din(n7809), .dout(n7810));
  jand g07577(.dina(n7810), .dinb(n7806), .dout(n7811));
  jor  g07578(.dina(n7811), .dinb(n7805), .dout(n7812));
  jand g07579(.dina(n7812), .dinb(asqrt[62] ), .dout(n7813));
  jor  g07580(.dina(n7812), .dinb(asqrt[62] ), .dout(n7814));
  jxor g07581(.dina(n7383), .dinb(n239), .dout(n7815));
  jand g07582(.dina(n7815), .dinb(asqrt[30] ), .dout(n7816));
  jxor g07583(.dina(n7816), .dinb(n7388), .dout(n7817));
  jand g07584(.dina(n7817), .dinb(n7814), .dout(n7818));
  jor  g07585(.dina(n7818), .dinb(n7813), .dout(n7819));
  jor  g07586(.dina(n7819), .dinb(n7419), .dout(n7820));
  jnot g07587(.din(n7820), .dout(n7821));
  jand g07588(.dina(n7581), .dinb(n7399), .dout(n7822));
  jnot g07589(.din(n7822), .dout(n7823));
  jnot g07590(.din(n7408), .dout(n7824));
  jand g07591(.dina(n7403), .dinb(asqrt[63] ), .dout(n7825));
  jand g07592(.dina(n7825), .dinb(n7824), .dout(n7826));
  jand g07593(.dina(n7826), .dinb(n7823), .dout(n7827));
  jnot g07594(.din(n7419), .dout(n7828));
  jnot g07595(.din(n7813), .dout(n7829));
  jnot g07596(.din(n7805), .dout(n7830));
  jnot g07597(.din(n7797), .dout(n7831));
  jnot g07598(.din(n7789), .dout(n7832));
  jnot g07599(.din(n7782), .dout(n7833));
  jnot g07600(.din(n7775), .dout(n7834));
  jnot g07601(.din(n7767), .dout(n7835));
  jnot g07602(.din(n7760), .dout(n7836));
  jnot g07603(.din(n7752), .dout(n7837));
  jnot g07604(.din(n7745), .dout(n7838));
  jnot g07605(.din(n7737), .dout(n7839));
  jnot g07606(.din(n7729), .dout(n7840));
  jnot g07607(.din(n7721), .dout(n7841));
  jnot g07608(.din(n7714), .dout(n7842));
  jnot g07609(.din(n7707), .dout(n7843));
  jnot g07610(.din(n7700), .dout(n7844));
  jnot g07611(.din(n7692), .dout(n7845));
  jnot g07612(.din(n7685), .dout(n7846));
  jnot g07613(.din(n7677), .dout(n7847));
  jnot g07614(.din(n7670), .dout(n7848));
  jnot g07615(.din(n7662), .dout(n7849));
  jnot g07616(.din(n7655), .dout(n7850));
  jnot g07617(.din(n7647), .dout(n7851));
  jnot g07618(.din(n7640), .dout(n7852));
  jnot g07619(.din(n7633), .dout(n7853));
  jnot g07620(.din(n7626), .dout(n7854));
  jnot g07621(.din(n7618), .dout(n7855));
  jnot g07622(.din(n7611), .dout(n7856));
  jnot g07623(.din(n7603), .dout(n7857));
  jnot g07624(.din(n7596), .dout(n7858));
  jnot g07625(.din(n7599), .dout(n7859));
  jnot g07626(.din(n7586), .dout(n7860));
  jnot g07627(.din(n7426), .dout(n7861));
  jor  g07628(.dina(n7581), .dinb(n7156), .dout(n7862));
  jnot g07629(.din(n7424), .dout(n7863));
  jand g07630(.dina(n7863), .dinb(n7862), .dout(n7864));
  jand g07631(.dina(n7864), .dinb(n7154), .dout(n7865));
  jor  g07632(.dina(n7581), .dinb(a[60] ), .dout(n7866));
  jand g07633(.dina(n7866), .dinb(a[61] ), .dout(n7867));
  jand g07634(.dina(asqrt[30] ), .dinb(n7158), .dout(n7868));
  jor  g07635(.dina(n7868), .dinb(n7867), .dout(n7869));
  jor  g07636(.dina(n7869), .dinb(n7865), .dout(n7870));
  jand g07637(.dina(n7870), .dinb(n7861), .dout(n7871));
  jand g07638(.dina(n7871), .dinb(n6758), .dout(n7872));
  jor  g07639(.dina(n7592), .dinb(n7872), .dout(n7873));
  jand g07640(.dina(n7873), .dinb(n7860), .dout(n7874));
  jand g07641(.dina(n7874), .dinb(n6357), .dout(n7875));
  jor  g07642(.dina(n7875), .dinb(n7859), .dout(n7876));
  jand g07643(.dina(n7876), .dinb(n7858), .dout(n7877));
  jand g07644(.dina(n7877), .dinb(n5989), .dout(n7878));
  jor  g07645(.dina(n7607), .dinb(n7878), .dout(n7879));
  jand g07646(.dina(n7879), .dinb(n7857), .dout(n7880));
  jand g07647(.dina(n7880), .dinb(n5606), .dout(n7881));
  jnot g07648(.din(n7615), .dout(n7882));
  jor  g07649(.dina(n7882), .dinb(n7881), .dout(n7883));
  jand g07650(.dina(n7883), .dinb(n7856), .dout(n7884));
  jand g07651(.dina(n7884), .dinb(n5259), .dout(n7885));
  jor  g07652(.dina(n7622), .dinb(n7885), .dout(n7886));
  jand g07653(.dina(n7886), .dinb(n7855), .dout(n7887));
  jand g07654(.dina(n7887), .dinb(n4902), .dout(n7888));
  jnot g07655(.din(n7630), .dout(n7889));
  jor  g07656(.dina(n7889), .dinb(n7888), .dout(n7890));
  jand g07657(.dina(n7890), .dinb(n7854), .dout(n7891));
  jand g07658(.dina(n7891), .dinb(n4582), .dout(n7892));
  jnot g07659(.din(n7637), .dout(n7893));
  jor  g07660(.dina(n7893), .dinb(n7892), .dout(n7894));
  jand g07661(.dina(n7894), .dinb(n7853), .dout(n7895));
  jand g07662(.dina(n7895), .dinb(n4249), .dout(n7896));
  jnot g07663(.din(n7644), .dout(n7897));
  jor  g07664(.dina(n7897), .dinb(n7896), .dout(n7898));
  jand g07665(.dina(n7898), .dinb(n7852), .dout(n7899));
  jand g07666(.dina(n7899), .dinb(n3955), .dout(n7900));
  jor  g07667(.dina(n7651), .dinb(n7900), .dout(n7901));
  jand g07668(.dina(n7901), .dinb(n7851), .dout(n7902));
  jand g07669(.dina(n7902), .dinb(n3642), .dout(n7903));
  jnot g07670(.din(n7659), .dout(n7904));
  jor  g07671(.dina(n7904), .dinb(n7903), .dout(n7905));
  jand g07672(.dina(n7905), .dinb(n7850), .dout(n7906));
  jand g07673(.dina(n7906), .dinb(n3368), .dout(n7907));
  jor  g07674(.dina(n7666), .dinb(n7907), .dout(n7908));
  jand g07675(.dina(n7908), .dinb(n7849), .dout(n7909));
  jand g07676(.dina(n7909), .dinb(n3089), .dout(n7910));
  jnot g07677(.din(n7674), .dout(n7911));
  jor  g07678(.dina(n7911), .dinb(n7910), .dout(n7912));
  jand g07679(.dina(n7912), .dinb(n7848), .dout(n7913));
  jand g07680(.dina(n7913), .dinb(n2833), .dout(n7914));
  jor  g07681(.dina(n7681), .dinb(n7914), .dout(n7915));
  jand g07682(.dina(n7915), .dinb(n7847), .dout(n7916));
  jand g07683(.dina(n7916), .dinb(n2572), .dout(n7917));
  jnot g07684(.din(n7689), .dout(n7918));
  jor  g07685(.dina(n7918), .dinb(n7917), .dout(n7919));
  jand g07686(.dina(n7919), .dinb(n7846), .dout(n7920));
  jand g07687(.dina(n7920), .dinb(n2345), .dout(n7921));
  jor  g07688(.dina(n7696), .dinb(n7921), .dout(n7922));
  jand g07689(.dina(n7922), .dinb(n7845), .dout(n7923));
  jand g07690(.dina(n7923), .dinb(n2108), .dout(n7924));
  jnot g07691(.din(n7704), .dout(n7925));
  jor  g07692(.dina(n7925), .dinb(n7924), .dout(n7926));
  jand g07693(.dina(n7926), .dinb(n7844), .dout(n7927));
  jand g07694(.dina(n7927), .dinb(n1912), .dout(n7928));
  jnot g07695(.din(n7711), .dout(n7929));
  jor  g07696(.dina(n7929), .dinb(n7928), .dout(n7930));
  jand g07697(.dina(n7930), .dinb(n7843), .dout(n7931));
  jand g07698(.dina(n7931), .dinb(n1699), .dout(n7932));
  jnot g07699(.din(n7718), .dout(n7933));
  jor  g07700(.dina(n7933), .dinb(n7932), .dout(n7934));
  jand g07701(.dina(n7934), .dinb(n7842), .dout(n7935));
  jand g07702(.dina(n7935), .dinb(n1516), .dout(n7936));
  jor  g07703(.dina(n7725), .dinb(n7936), .dout(n7937));
  jand g07704(.dina(n7937), .dinb(n7841), .dout(n7938));
  jand g07705(.dina(n7938), .dinb(n1332), .dout(n7939));
  jor  g07706(.dina(n7733), .dinb(n7939), .dout(n7940));
  jand g07707(.dina(n7940), .dinb(n7840), .dout(n7941));
  jand g07708(.dina(n7941), .dinb(n1173), .dout(n7942));
  jor  g07709(.dina(n7741), .dinb(n7942), .dout(n7943));
  jand g07710(.dina(n7943), .dinb(n7839), .dout(n7944));
  jand g07711(.dina(n7944), .dinb(n1008), .dout(n7945));
  jnot g07712(.din(n7749), .dout(n7946));
  jor  g07713(.dina(n7946), .dinb(n7945), .dout(n7947));
  jand g07714(.dina(n7947), .dinb(n7838), .dout(n7948));
  jand g07715(.dina(n7948), .dinb(n884), .dout(n7949));
  jor  g07716(.dina(n7756), .dinb(n7949), .dout(n7950));
  jand g07717(.dina(n7950), .dinb(n7837), .dout(n7951));
  jand g07718(.dina(n7951), .dinb(n743), .dout(n7952));
  jnot g07719(.din(n7764), .dout(n7953));
  jor  g07720(.dina(n7953), .dinb(n7952), .dout(n7954));
  jand g07721(.dina(n7954), .dinb(n7836), .dout(n7955));
  jand g07722(.dina(n7955), .dinb(n635), .dout(n7956));
  jor  g07723(.dina(n7771), .dinb(n7956), .dout(n7957));
  jand g07724(.dina(n7957), .dinb(n7835), .dout(n7958));
  jand g07725(.dina(n7958), .dinb(n515), .dout(n7959));
  jnot g07726(.din(n7779), .dout(n7960));
  jor  g07727(.dina(n7960), .dinb(n7959), .dout(n7961));
  jand g07728(.dina(n7961), .dinb(n7834), .dout(n7962));
  jand g07729(.dina(n7962), .dinb(n443), .dout(n7963));
  jnot g07730(.din(n7786), .dout(n7964));
  jor  g07731(.dina(n7964), .dinb(n7963), .dout(n7965));
  jand g07732(.dina(n7965), .dinb(n7833), .dout(n7966));
  jand g07733(.dina(n7966), .dinb(n352), .dout(n7967));
  jor  g07734(.dina(n7793), .dinb(n7967), .dout(n7968));
  jand g07735(.dina(n7968), .dinb(n7832), .dout(n7969));
  jand g07736(.dina(n7969), .dinb(n294), .dout(n7970));
  jor  g07737(.dina(n7801), .dinb(n7970), .dout(n7971));
  jand g07738(.dina(n7971), .dinb(n7831), .dout(n7972));
  jand g07739(.dina(n7972), .dinb(n239), .dout(n7973));
  jor  g07740(.dina(n7809), .dinb(n7973), .dout(n7974));
  jand g07741(.dina(n7974), .dinb(n7830), .dout(n7975));
  jand g07742(.dina(n7975), .dinb(n221), .dout(n7976));
  jnot g07743(.din(n7817), .dout(n7977));
  jor  g07744(.dina(n7977), .dinb(n7976), .dout(n7978));
  jand g07745(.dina(n7978), .dinb(n7829), .dout(n7979));
  jor  g07746(.dina(n7979), .dinb(n7828), .dout(n7980));
  jand g07747(.dina(asqrt[30] ), .dinb(n7576), .dout(n7981));
  jor  g07748(.dina(n7981), .dinb(n7408), .dout(n7982));
  jor  g07749(.dina(n7982), .dinb(n7980), .dout(n7983));
  jand g07750(.dina(n7983), .dinb(n218), .dout(n7984));
  jand g07751(.dina(n7581), .dinb(n7402), .dout(n7985));
  jor  g07752(.dina(n7985), .dinb(n7984), .dout(n7986));
  jor  g07753(.dina(n7986), .dinb(n7827), .dout(n7987));
  jor  g07754(.dina(n7987), .dinb(n7821), .dout(asqrt[29] ));
  jand g07755(.dina(n7819), .dinb(n7419), .dout(n7989));
  jand g07756(.dina(n7987), .dinb(n7989), .dout(n7990));
  jnot g07757(.din(a[56] ), .dout(n7991));
  jnot g07758(.din(a[57] ), .dout(n7992));
  jand g07759(.dina(n7992), .dinb(n7991), .dout(n7993));
  jand g07760(.dina(n7993), .dinb(n7421), .dout(n7994));
  jnot g07761(.din(n7994), .dout(n7995));
  jnot g07762(.din(n7827), .dout(n7996));
  jnot g07763(.din(n7982), .dout(n7997));
  jand g07764(.dina(n7997), .dinb(n7989), .dout(n7998));
  jor  g07765(.dina(n7998), .dinb(asqrt[63] ), .dout(n7999));
  jnot g07766(.din(n7985), .dout(n8000));
  jand g07767(.dina(n8000), .dinb(n7999), .dout(n8001));
  jand g07768(.dina(n8001), .dinb(n7996), .dout(n8002));
  jand g07769(.dina(n8002), .dinb(n7820), .dout(n8003));
  jor  g07770(.dina(n8003), .dinb(n7421), .dout(n8004));
  jand g07771(.dina(n8004), .dinb(n7995), .dout(n8005));
  jor  g07772(.dina(n8005), .dinb(n7581), .dout(n8006));
  jand g07773(.dina(n8005), .dinb(n7581), .dout(n8007));
  jor  g07774(.dina(n8003), .dinb(a[58] ), .dout(n8008));
  jand g07775(.dina(n8008), .dinb(a[59] ), .dout(n8009));
  jand g07776(.dina(asqrt[29] ), .dinb(n7423), .dout(n8010));
  jor  g07777(.dina(n8010), .dinb(n8009), .dout(n8011));
  jor  g07778(.dina(n8011), .dinb(n8007), .dout(n8012));
  jand g07779(.dina(n8012), .dinb(n8006), .dout(n8013));
  jor  g07780(.dina(n8013), .dinb(n7154), .dout(n8014));
  jand g07781(.dina(n8013), .dinb(n7154), .dout(n8015));
  jnot g07782(.din(n7423), .dout(n8016));
  jor  g07783(.dina(n8003), .dinb(n8016), .dout(n8017));
  jor  g07784(.dina(n7821), .dinb(n7581), .dout(n8018));
  jor  g07785(.dina(n8018), .dinb(n7826), .dout(n8019));
  jor  g07786(.dina(n8019), .dinb(n7984), .dout(n8020));
  jand g07787(.dina(n8020), .dinb(n8017), .dout(n8021));
  jxor g07788(.dina(n8021), .dinb(n7156), .dout(n8022));
  jor  g07789(.dina(n8022), .dinb(n8015), .dout(n8023));
  jand g07790(.dina(n8023), .dinb(n8014), .dout(n8024));
  jor  g07791(.dina(n8024), .dinb(n6758), .dout(n8025));
  jand g07792(.dina(n8024), .dinb(n6758), .dout(n8026));
  jxor g07793(.dina(n7425), .dinb(n7154), .dout(n8027));
  jor  g07794(.dina(n8027), .dinb(n8003), .dout(n8028));
  jxor g07795(.dina(n8028), .dinb(n7583), .dout(n8029));
  jor  g07796(.dina(n8029), .dinb(n8026), .dout(n8030));
  jand g07797(.dina(n8030), .dinb(n8025), .dout(n8031));
  jor  g07798(.dina(n8031), .dinb(n6357), .dout(n8032));
  jand g07799(.dina(n8031), .dinb(n6357), .dout(n8033));
  jxor g07800(.dina(n7585), .dinb(n6758), .dout(n8034));
  jor  g07801(.dina(n8034), .dinb(n8003), .dout(n8035));
  jxor g07802(.dina(n8035), .dinb(n7593), .dout(n8036));
  jor  g07803(.dina(n8036), .dinb(n8033), .dout(n8037));
  jand g07804(.dina(n8037), .dinb(n8032), .dout(n8038));
  jor  g07805(.dina(n8038), .dinb(n5989), .dout(n8039));
  jxor g07806(.dina(n7595), .dinb(n6357), .dout(n8040));
  jor  g07807(.dina(n8040), .dinb(n8003), .dout(n8041));
  jxor g07808(.dina(n8041), .dinb(n7859), .dout(n8042));
  jnot g07809(.din(n8042), .dout(n8043));
  jand g07810(.dina(n8038), .dinb(n5989), .dout(n8044));
  jor  g07811(.dina(n8044), .dinb(n8043), .dout(n8045));
  jand g07812(.dina(n8045), .dinb(n8039), .dout(n8046));
  jor  g07813(.dina(n8046), .dinb(n5606), .dout(n8047));
  jand g07814(.dina(n8046), .dinb(n5606), .dout(n8048));
  jxor g07815(.dina(n7602), .dinb(n5989), .dout(n8049));
  jor  g07816(.dina(n8049), .dinb(n8003), .dout(n8050));
  jxor g07817(.dina(n8050), .dinb(n7608), .dout(n8051));
  jor  g07818(.dina(n8051), .dinb(n8048), .dout(n8052));
  jand g07819(.dina(n8052), .dinb(n8047), .dout(n8053));
  jor  g07820(.dina(n8053), .dinb(n5259), .dout(n8054));
  jand g07821(.dina(n8053), .dinb(n5259), .dout(n8055));
  jxor g07822(.dina(n7610), .dinb(n5606), .dout(n8056));
  jor  g07823(.dina(n8056), .dinb(n8003), .dout(n8057));
  jxor g07824(.dina(n8057), .dinb(n7882), .dout(n8058));
  jnot g07825(.din(n8058), .dout(n8059));
  jor  g07826(.dina(n8059), .dinb(n8055), .dout(n8060));
  jand g07827(.dina(n8060), .dinb(n8054), .dout(n8061));
  jor  g07828(.dina(n8061), .dinb(n4902), .dout(n8062));
  jand g07829(.dina(n8061), .dinb(n4902), .dout(n8063));
  jxor g07830(.dina(n7617), .dinb(n5259), .dout(n8064));
  jor  g07831(.dina(n8064), .dinb(n8003), .dout(n8065));
  jxor g07832(.dina(n8065), .dinb(n7623), .dout(n8066));
  jor  g07833(.dina(n8066), .dinb(n8063), .dout(n8067));
  jand g07834(.dina(n8067), .dinb(n8062), .dout(n8068));
  jor  g07835(.dina(n8068), .dinb(n4582), .dout(n8069));
  jand g07836(.dina(n8068), .dinb(n4582), .dout(n8070));
  jxor g07837(.dina(n7625), .dinb(n4902), .dout(n8071));
  jor  g07838(.dina(n8071), .dinb(n8003), .dout(n8072));
  jxor g07839(.dina(n8072), .dinb(n7889), .dout(n8073));
  jnot g07840(.din(n8073), .dout(n8074));
  jor  g07841(.dina(n8074), .dinb(n8070), .dout(n8075));
  jand g07842(.dina(n8075), .dinb(n8069), .dout(n8076));
  jor  g07843(.dina(n8076), .dinb(n4249), .dout(n8077));
  jand g07844(.dina(n8076), .dinb(n4249), .dout(n8078));
  jxor g07845(.dina(n7632), .dinb(n4582), .dout(n8079));
  jor  g07846(.dina(n8079), .dinb(n8003), .dout(n8080));
  jxor g07847(.dina(n8080), .dinb(n7893), .dout(n8081));
  jnot g07848(.din(n8081), .dout(n8082));
  jor  g07849(.dina(n8082), .dinb(n8078), .dout(n8083));
  jand g07850(.dina(n8083), .dinb(n8077), .dout(n8084));
  jor  g07851(.dina(n8084), .dinb(n3955), .dout(n8085));
  jand g07852(.dina(n8084), .dinb(n3955), .dout(n8086));
  jxor g07853(.dina(n7639), .dinb(n4249), .dout(n8087));
  jor  g07854(.dina(n8087), .dinb(n8003), .dout(n8088));
  jxor g07855(.dina(n8088), .dinb(n7897), .dout(n8089));
  jnot g07856(.din(n8089), .dout(n8090));
  jor  g07857(.dina(n8090), .dinb(n8086), .dout(n8091));
  jand g07858(.dina(n8091), .dinb(n8085), .dout(n8092));
  jor  g07859(.dina(n8092), .dinb(n3642), .dout(n8093));
  jand g07860(.dina(n8092), .dinb(n3642), .dout(n8094));
  jxor g07861(.dina(n7646), .dinb(n3955), .dout(n8095));
  jor  g07862(.dina(n8095), .dinb(n8003), .dout(n8096));
  jxor g07863(.dina(n8096), .dinb(n7652), .dout(n8097));
  jor  g07864(.dina(n8097), .dinb(n8094), .dout(n8098));
  jand g07865(.dina(n8098), .dinb(n8093), .dout(n8099));
  jor  g07866(.dina(n8099), .dinb(n3368), .dout(n8100));
  jand g07867(.dina(n8099), .dinb(n3368), .dout(n8101));
  jxor g07868(.dina(n7654), .dinb(n3642), .dout(n8102));
  jor  g07869(.dina(n8102), .dinb(n8003), .dout(n8103));
  jxor g07870(.dina(n8103), .dinb(n7904), .dout(n8104));
  jnot g07871(.din(n8104), .dout(n8105));
  jor  g07872(.dina(n8105), .dinb(n8101), .dout(n8106));
  jand g07873(.dina(n8106), .dinb(n8100), .dout(n8107));
  jor  g07874(.dina(n8107), .dinb(n3089), .dout(n8108));
  jand g07875(.dina(n8107), .dinb(n3089), .dout(n8109));
  jxor g07876(.dina(n7661), .dinb(n3368), .dout(n8110));
  jor  g07877(.dina(n8110), .dinb(n8003), .dout(n8111));
  jxor g07878(.dina(n8111), .dinb(n7667), .dout(n8112));
  jor  g07879(.dina(n8112), .dinb(n8109), .dout(n8113));
  jand g07880(.dina(n8113), .dinb(n8108), .dout(n8114));
  jor  g07881(.dina(n8114), .dinb(n2833), .dout(n8115));
  jand g07882(.dina(n8114), .dinb(n2833), .dout(n8116));
  jxor g07883(.dina(n7669), .dinb(n3089), .dout(n8117));
  jor  g07884(.dina(n8117), .dinb(n8003), .dout(n8118));
  jxor g07885(.dina(n8118), .dinb(n7911), .dout(n8119));
  jnot g07886(.din(n8119), .dout(n8120));
  jor  g07887(.dina(n8120), .dinb(n8116), .dout(n8121));
  jand g07888(.dina(n8121), .dinb(n8115), .dout(n8122));
  jor  g07889(.dina(n8122), .dinb(n2572), .dout(n8123));
  jand g07890(.dina(n8122), .dinb(n2572), .dout(n8124));
  jxor g07891(.dina(n7676), .dinb(n2833), .dout(n8125));
  jor  g07892(.dina(n8125), .dinb(n8003), .dout(n8126));
  jxor g07893(.dina(n8126), .dinb(n7682), .dout(n8127));
  jor  g07894(.dina(n8127), .dinb(n8124), .dout(n8128));
  jand g07895(.dina(n8128), .dinb(n8123), .dout(n8129));
  jor  g07896(.dina(n8129), .dinb(n2345), .dout(n8130));
  jand g07897(.dina(n8129), .dinb(n2345), .dout(n8131));
  jxor g07898(.dina(n7684), .dinb(n2572), .dout(n8132));
  jor  g07899(.dina(n8132), .dinb(n8003), .dout(n8133));
  jxor g07900(.dina(n8133), .dinb(n7918), .dout(n8134));
  jnot g07901(.din(n8134), .dout(n8135));
  jor  g07902(.dina(n8135), .dinb(n8131), .dout(n8136));
  jand g07903(.dina(n8136), .dinb(n8130), .dout(n8137));
  jor  g07904(.dina(n8137), .dinb(n2108), .dout(n8138));
  jand g07905(.dina(n8137), .dinb(n2108), .dout(n8139));
  jxor g07906(.dina(n7691), .dinb(n2345), .dout(n8140));
  jor  g07907(.dina(n8140), .dinb(n8003), .dout(n8141));
  jxor g07908(.dina(n8141), .dinb(n7697), .dout(n8142));
  jor  g07909(.dina(n8142), .dinb(n8139), .dout(n8143));
  jand g07910(.dina(n8143), .dinb(n8138), .dout(n8144));
  jor  g07911(.dina(n8144), .dinb(n1912), .dout(n8145));
  jand g07912(.dina(n8144), .dinb(n1912), .dout(n8146));
  jxor g07913(.dina(n7699), .dinb(n2108), .dout(n8147));
  jor  g07914(.dina(n8147), .dinb(n8003), .dout(n8148));
  jxor g07915(.dina(n8148), .dinb(n7925), .dout(n8149));
  jnot g07916(.din(n8149), .dout(n8150));
  jor  g07917(.dina(n8150), .dinb(n8146), .dout(n8151));
  jand g07918(.dina(n8151), .dinb(n8145), .dout(n8152));
  jor  g07919(.dina(n8152), .dinb(n1699), .dout(n8153));
  jand g07920(.dina(n8152), .dinb(n1699), .dout(n8154));
  jxor g07921(.dina(n7706), .dinb(n1912), .dout(n8155));
  jor  g07922(.dina(n8155), .dinb(n8003), .dout(n8156));
  jxor g07923(.dina(n8156), .dinb(n7929), .dout(n8157));
  jnot g07924(.din(n8157), .dout(n8158));
  jor  g07925(.dina(n8158), .dinb(n8154), .dout(n8159));
  jand g07926(.dina(n8159), .dinb(n8153), .dout(n8160));
  jor  g07927(.dina(n8160), .dinb(n1516), .dout(n8161));
  jand g07928(.dina(n8160), .dinb(n1516), .dout(n8162));
  jxor g07929(.dina(n7713), .dinb(n1699), .dout(n8163));
  jor  g07930(.dina(n8163), .dinb(n8003), .dout(n8164));
  jxor g07931(.dina(n8164), .dinb(n7933), .dout(n8165));
  jnot g07932(.din(n8165), .dout(n8166));
  jor  g07933(.dina(n8166), .dinb(n8162), .dout(n8167));
  jand g07934(.dina(n8167), .dinb(n8161), .dout(n8168));
  jor  g07935(.dina(n8168), .dinb(n1332), .dout(n8169));
  jand g07936(.dina(n8168), .dinb(n1332), .dout(n8170));
  jxor g07937(.dina(n7720), .dinb(n1516), .dout(n8171));
  jor  g07938(.dina(n8171), .dinb(n8003), .dout(n8172));
  jxor g07939(.dina(n8172), .dinb(n7726), .dout(n8173));
  jor  g07940(.dina(n8173), .dinb(n8170), .dout(n8174));
  jand g07941(.dina(n8174), .dinb(n8169), .dout(n8175));
  jor  g07942(.dina(n8175), .dinb(n1173), .dout(n8176));
  jand g07943(.dina(n8175), .dinb(n1173), .dout(n8177));
  jxor g07944(.dina(n7728), .dinb(n1332), .dout(n8178));
  jor  g07945(.dina(n8178), .dinb(n8003), .dout(n8179));
  jxor g07946(.dina(n8179), .dinb(n7734), .dout(n8180));
  jor  g07947(.dina(n8180), .dinb(n8177), .dout(n8181));
  jand g07948(.dina(n8181), .dinb(n8176), .dout(n8182));
  jor  g07949(.dina(n8182), .dinb(n1008), .dout(n8183));
  jand g07950(.dina(n8182), .dinb(n1008), .dout(n8184));
  jxor g07951(.dina(n7736), .dinb(n1173), .dout(n8185));
  jor  g07952(.dina(n8185), .dinb(n8003), .dout(n8186));
  jxor g07953(.dina(n8186), .dinb(n7742), .dout(n8187));
  jor  g07954(.dina(n8187), .dinb(n8184), .dout(n8188));
  jand g07955(.dina(n8188), .dinb(n8183), .dout(n8189));
  jor  g07956(.dina(n8189), .dinb(n884), .dout(n8190));
  jand g07957(.dina(n8189), .dinb(n884), .dout(n8191));
  jxor g07958(.dina(n7744), .dinb(n1008), .dout(n8192));
  jor  g07959(.dina(n8192), .dinb(n8003), .dout(n8193));
  jxor g07960(.dina(n8193), .dinb(n7946), .dout(n8194));
  jnot g07961(.din(n8194), .dout(n8195));
  jor  g07962(.dina(n8195), .dinb(n8191), .dout(n8196));
  jand g07963(.dina(n8196), .dinb(n8190), .dout(n8197));
  jor  g07964(.dina(n8197), .dinb(n743), .dout(n8198));
  jand g07965(.dina(n8197), .dinb(n743), .dout(n8199));
  jxor g07966(.dina(n7751), .dinb(n884), .dout(n8200));
  jor  g07967(.dina(n8200), .dinb(n8003), .dout(n8201));
  jxor g07968(.dina(n8201), .dinb(n7757), .dout(n8202));
  jor  g07969(.dina(n8202), .dinb(n8199), .dout(n8203));
  jand g07970(.dina(n8203), .dinb(n8198), .dout(n8204));
  jor  g07971(.dina(n8204), .dinb(n635), .dout(n8205));
  jand g07972(.dina(n8204), .dinb(n635), .dout(n8206));
  jxor g07973(.dina(n7759), .dinb(n743), .dout(n8207));
  jor  g07974(.dina(n8207), .dinb(n8003), .dout(n8208));
  jxor g07975(.dina(n8208), .dinb(n7953), .dout(n8209));
  jnot g07976(.din(n8209), .dout(n8210));
  jor  g07977(.dina(n8210), .dinb(n8206), .dout(n8211));
  jand g07978(.dina(n8211), .dinb(n8205), .dout(n8212));
  jor  g07979(.dina(n8212), .dinb(n515), .dout(n8213));
  jand g07980(.dina(n8212), .dinb(n515), .dout(n8214));
  jxor g07981(.dina(n7766), .dinb(n635), .dout(n8215));
  jor  g07982(.dina(n8215), .dinb(n8003), .dout(n8216));
  jxor g07983(.dina(n8216), .dinb(n7772), .dout(n8217));
  jor  g07984(.dina(n8217), .dinb(n8214), .dout(n8218));
  jand g07985(.dina(n8218), .dinb(n8213), .dout(n8219));
  jor  g07986(.dina(n8219), .dinb(n443), .dout(n8220));
  jand g07987(.dina(n8219), .dinb(n443), .dout(n8221));
  jxor g07988(.dina(n7774), .dinb(n515), .dout(n8222));
  jor  g07989(.dina(n8222), .dinb(n8003), .dout(n8223));
  jxor g07990(.dina(n8223), .dinb(n7960), .dout(n8224));
  jnot g07991(.din(n8224), .dout(n8225));
  jor  g07992(.dina(n8225), .dinb(n8221), .dout(n8226));
  jand g07993(.dina(n8226), .dinb(n8220), .dout(n8227));
  jor  g07994(.dina(n8227), .dinb(n352), .dout(n8228));
  jand g07995(.dina(n8227), .dinb(n352), .dout(n8229));
  jxor g07996(.dina(n7781), .dinb(n443), .dout(n8230));
  jor  g07997(.dina(n8230), .dinb(n8003), .dout(n8231));
  jxor g07998(.dina(n8231), .dinb(n7964), .dout(n8232));
  jnot g07999(.din(n8232), .dout(n8233));
  jor  g08000(.dina(n8233), .dinb(n8229), .dout(n8234));
  jand g08001(.dina(n8234), .dinb(n8228), .dout(n8235));
  jor  g08002(.dina(n8235), .dinb(n294), .dout(n8236));
  jand g08003(.dina(n8235), .dinb(n294), .dout(n8237));
  jxor g08004(.dina(n7788), .dinb(n352), .dout(n8238));
  jor  g08005(.dina(n8238), .dinb(n8003), .dout(n8239));
  jxor g08006(.dina(n8239), .dinb(n7794), .dout(n8240));
  jor  g08007(.dina(n8240), .dinb(n8237), .dout(n8241));
  jand g08008(.dina(n8241), .dinb(n8236), .dout(n8242));
  jor  g08009(.dina(n8242), .dinb(n239), .dout(n8243));
  jand g08010(.dina(n8242), .dinb(n239), .dout(n8244));
  jxor g08011(.dina(n7796), .dinb(n294), .dout(n8245));
  jor  g08012(.dina(n8245), .dinb(n8003), .dout(n8246));
  jxor g08013(.dina(n8246), .dinb(n7802), .dout(n8247));
  jor  g08014(.dina(n8247), .dinb(n8244), .dout(n8248));
  jand g08015(.dina(n8248), .dinb(n8243), .dout(n8249));
  jor  g08016(.dina(n8249), .dinb(n221), .dout(n8250));
  jand g08017(.dina(n8249), .dinb(n221), .dout(n8251));
  jxor g08018(.dina(n7804), .dinb(n239), .dout(n8252));
  jor  g08019(.dina(n8252), .dinb(n8003), .dout(n8253));
  jxor g08020(.dina(n8253), .dinb(n7810), .dout(n8254));
  jor  g08021(.dina(n8254), .dinb(n8251), .dout(n8255));
  jand g08022(.dina(n8255), .dinb(n8250), .dout(n8256));
  jxor g08023(.dina(n7812), .dinb(n221), .dout(n8257));
  jor  g08024(.dina(n8257), .dinb(n8003), .dout(n8258));
  jxor g08025(.dina(n8258), .dinb(n7817), .dout(n8259));
  jor  g08026(.dina(n8259), .dinb(n8256), .dout(n8260));
  jor  g08027(.dina(n8260), .dinb(n7821), .dout(n8261));
  jor  g08028(.dina(n8261), .dinb(n7990), .dout(n8262));
  jand g08029(.dina(n8262), .dinb(n218), .dout(n8263));
  jand g08030(.dina(n8003), .dinb(n7828), .dout(n8264));
  jand g08031(.dina(n8259), .dinb(n8256), .dout(n8265));
  jor  g08032(.dina(n8265), .dinb(n8264), .dout(n8266));
  jand g08033(.dina(n8002), .dinb(n7979), .dout(n8267));
  jnot g08034(.din(n8267), .dout(n8268));
  jand g08035(.dina(n7980), .dinb(asqrt[63] ), .dout(n8269));
  jand g08036(.dina(n8269), .dinb(n7820), .dout(n8270));
  jand g08037(.dina(n8270), .dinb(n8268), .dout(n8271));
  jor  g08038(.dina(n8271), .dinb(n8266), .dout(n8272));
  jor  g08039(.dina(n8272), .dinb(n8263), .dout(asqrt[28] ));
  jnot g08040(.din(n8254), .dout(n8274));
  jxor g08041(.dina(n8249), .dinb(n221), .dout(n8275));
  jand g08042(.dina(n8275), .dinb(asqrt[28] ), .dout(n8276));
  jxor g08043(.dina(n8276), .dinb(n8274), .dout(n8277));
  jand g08044(.dina(asqrt[28] ), .dinb(a[56] ), .dout(n8278));
  jnot g08045(.din(a[54] ), .dout(n8279));
  jnot g08046(.din(a[55] ), .dout(n8280));
  jand g08047(.dina(n8280), .dinb(n8279), .dout(n8281));
  jand g08048(.dina(n8281), .dinb(n7991), .dout(n8282));
  jor  g08049(.dina(n8282), .dinb(n8278), .dout(n8283));
  jand g08050(.dina(n8283), .dinb(asqrt[29] ), .dout(n8284));
  jor  g08051(.dina(n8283), .dinb(asqrt[29] ), .dout(n8285));
  jand g08052(.dina(asqrt[28] ), .dinb(n7991), .dout(n8286));
  jor  g08053(.dina(n8286), .dinb(n7992), .dout(n8287));
  jnot g08054(.din(n7993), .dout(n8288));
  jnot g08055(.din(n7990), .dout(n8289));
  jnot g08056(.din(n8250), .dout(n8290));
  jnot g08057(.din(n8243), .dout(n8291));
  jnot g08058(.din(n8236), .dout(n8292));
  jnot g08059(.din(n8228), .dout(n8293));
  jnot g08060(.din(n8220), .dout(n8294));
  jnot g08061(.din(n8213), .dout(n8295));
  jnot g08062(.din(n8205), .dout(n8296));
  jnot g08063(.din(n8198), .dout(n8297));
  jnot g08064(.din(n8190), .dout(n8298));
  jnot g08065(.din(n8183), .dout(n8299));
  jnot g08066(.din(n8176), .dout(n8300));
  jnot g08067(.din(n8169), .dout(n8301));
  jnot g08068(.din(n8161), .dout(n8302));
  jnot g08069(.din(n8153), .dout(n8303));
  jnot g08070(.din(n8145), .dout(n8304));
  jnot g08071(.din(n8138), .dout(n8305));
  jnot g08072(.din(n8130), .dout(n8306));
  jnot g08073(.din(n8123), .dout(n8307));
  jnot g08074(.din(n8115), .dout(n8308));
  jnot g08075(.din(n8108), .dout(n8309));
  jnot g08076(.din(n8100), .dout(n8310));
  jnot g08077(.din(n8093), .dout(n8311));
  jnot g08078(.din(n8085), .dout(n8312));
  jnot g08079(.din(n8077), .dout(n8313));
  jnot g08080(.din(n8069), .dout(n8314));
  jnot g08081(.din(n8062), .dout(n8315));
  jnot g08082(.din(n8054), .dout(n8316));
  jnot g08083(.din(n8047), .dout(n8317));
  jnot g08084(.din(n8039), .dout(n8318));
  jnot g08085(.din(n8032), .dout(n8319));
  jnot g08086(.din(n8025), .dout(n8320));
  jnot g08087(.din(n8014), .dout(n8321));
  jnot g08088(.din(n8006), .dout(n8322));
  jand g08089(.dina(asqrt[29] ), .dinb(a[58] ), .dout(n8323));
  jor  g08090(.dina(n8323), .dinb(n7994), .dout(n8324));
  jor  g08091(.dina(n8324), .dinb(asqrt[30] ), .dout(n8325));
  jand g08092(.dina(asqrt[29] ), .dinb(n7421), .dout(n8326));
  jor  g08093(.dina(n8326), .dinb(n7422), .dout(n8327));
  jand g08094(.dina(n8017), .dinb(n8327), .dout(n8328));
  jand g08095(.dina(n8328), .dinb(n8325), .dout(n8329));
  jor  g08096(.dina(n8329), .dinb(n8322), .dout(n8330));
  jor  g08097(.dina(n8330), .dinb(asqrt[31] ), .dout(n8331));
  jnot g08098(.din(n8022), .dout(n8332));
  jand g08099(.dina(n8332), .dinb(n8331), .dout(n8333));
  jor  g08100(.dina(n8333), .dinb(n8321), .dout(n8334));
  jor  g08101(.dina(n8334), .dinb(asqrt[32] ), .dout(n8335));
  jnot g08102(.din(n8029), .dout(n8336));
  jand g08103(.dina(n8336), .dinb(n8335), .dout(n8337));
  jor  g08104(.dina(n8337), .dinb(n8320), .dout(n8338));
  jor  g08105(.dina(n8338), .dinb(asqrt[33] ), .dout(n8339));
  jnot g08106(.din(n8036), .dout(n8340));
  jand g08107(.dina(n8340), .dinb(n8339), .dout(n8341));
  jor  g08108(.dina(n8341), .dinb(n8319), .dout(n8342));
  jor  g08109(.dina(n8342), .dinb(asqrt[34] ), .dout(n8343));
  jand g08110(.dina(n8343), .dinb(n8042), .dout(n8344));
  jor  g08111(.dina(n8344), .dinb(n8318), .dout(n8345));
  jor  g08112(.dina(n8345), .dinb(asqrt[35] ), .dout(n8346));
  jnot g08113(.din(n8051), .dout(n8347));
  jand g08114(.dina(n8347), .dinb(n8346), .dout(n8348));
  jor  g08115(.dina(n8348), .dinb(n8317), .dout(n8349));
  jor  g08116(.dina(n8349), .dinb(asqrt[36] ), .dout(n8350));
  jand g08117(.dina(n8058), .dinb(n8350), .dout(n8351));
  jor  g08118(.dina(n8351), .dinb(n8316), .dout(n8352));
  jor  g08119(.dina(n8352), .dinb(asqrt[37] ), .dout(n8353));
  jnot g08120(.din(n8066), .dout(n8354));
  jand g08121(.dina(n8354), .dinb(n8353), .dout(n8355));
  jor  g08122(.dina(n8355), .dinb(n8315), .dout(n8356));
  jor  g08123(.dina(n8356), .dinb(asqrt[38] ), .dout(n8357));
  jand g08124(.dina(n8073), .dinb(n8357), .dout(n8358));
  jor  g08125(.dina(n8358), .dinb(n8314), .dout(n8359));
  jor  g08126(.dina(n8359), .dinb(asqrt[39] ), .dout(n8360));
  jand g08127(.dina(n8081), .dinb(n8360), .dout(n8361));
  jor  g08128(.dina(n8361), .dinb(n8313), .dout(n8362));
  jor  g08129(.dina(n8362), .dinb(asqrt[40] ), .dout(n8363));
  jand g08130(.dina(n8089), .dinb(n8363), .dout(n8364));
  jor  g08131(.dina(n8364), .dinb(n8312), .dout(n8365));
  jor  g08132(.dina(n8365), .dinb(asqrt[41] ), .dout(n8366));
  jnot g08133(.din(n8097), .dout(n8367));
  jand g08134(.dina(n8367), .dinb(n8366), .dout(n8368));
  jor  g08135(.dina(n8368), .dinb(n8311), .dout(n8369));
  jor  g08136(.dina(n8369), .dinb(asqrt[42] ), .dout(n8370));
  jand g08137(.dina(n8104), .dinb(n8370), .dout(n8371));
  jor  g08138(.dina(n8371), .dinb(n8310), .dout(n8372));
  jor  g08139(.dina(n8372), .dinb(asqrt[43] ), .dout(n8373));
  jnot g08140(.din(n8112), .dout(n8374));
  jand g08141(.dina(n8374), .dinb(n8373), .dout(n8375));
  jor  g08142(.dina(n8375), .dinb(n8309), .dout(n8376));
  jor  g08143(.dina(n8376), .dinb(asqrt[44] ), .dout(n8377));
  jand g08144(.dina(n8119), .dinb(n8377), .dout(n8378));
  jor  g08145(.dina(n8378), .dinb(n8308), .dout(n8379));
  jor  g08146(.dina(n8379), .dinb(asqrt[45] ), .dout(n8380));
  jnot g08147(.din(n8127), .dout(n8381));
  jand g08148(.dina(n8381), .dinb(n8380), .dout(n8382));
  jor  g08149(.dina(n8382), .dinb(n8307), .dout(n8383));
  jor  g08150(.dina(n8383), .dinb(asqrt[46] ), .dout(n8384));
  jand g08151(.dina(n8134), .dinb(n8384), .dout(n8385));
  jor  g08152(.dina(n8385), .dinb(n8306), .dout(n8386));
  jor  g08153(.dina(n8386), .dinb(asqrt[47] ), .dout(n8387));
  jnot g08154(.din(n8142), .dout(n8388));
  jand g08155(.dina(n8388), .dinb(n8387), .dout(n8389));
  jor  g08156(.dina(n8389), .dinb(n8305), .dout(n8390));
  jor  g08157(.dina(n8390), .dinb(asqrt[48] ), .dout(n8391));
  jand g08158(.dina(n8149), .dinb(n8391), .dout(n8392));
  jor  g08159(.dina(n8392), .dinb(n8304), .dout(n8393));
  jor  g08160(.dina(n8393), .dinb(asqrt[49] ), .dout(n8394));
  jand g08161(.dina(n8157), .dinb(n8394), .dout(n8395));
  jor  g08162(.dina(n8395), .dinb(n8303), .dout(n8396));
  jor  g08163(.dina(n8396), .dinb(asqrt[50] ), .dout(n8397));
  jand g08164(.dina(n8165), .dinb(n8397), .dout(n8398));
  jor  g08165(.dina(n8398), .dinb(n8302), .dout(n8399));
  jor  g08166(.dina(n8399), .dinb(asqrt[51] ), .dout(n8400));
  jnot g08167(.din(n8173), .dout(n8401));
  jand g08168(.dina(n8401), .dinb(n8400), .dout(n8402));
  jor  g08169(.dina(n8402), .dinb(n8301), .dout(n8403));
  jor  g08170(.dina(n8403), .dinb(asqrt[52] ), .dout(n8404));
  jnot g08171(.din(n8180), .dout(n8405));
  jand g08172(.dina(n8405), .dinb(n8404), .dout(n8406));
  jor  g08173(.dina(n8406), .dinb(n8300), .dout(n8407));
  jor  g08174(.dina(n8407), .dinb(asqrt[53] ), .dout(n8408));
  jnot g08175(.din(n8187), .dout(n8409));
  jand g08176(.dina(n8409), .dinb(n8408), .dout(n8410));
  jor  g08177(.dina(n8410), .dinb(n8299), .dout(n8411));
  jor  g08178(.dina(n8411), .dinb(asqrt[54] ), .dout(n8412));
  jand g08179(.dina(n8194), .dinb(n8412), .dout(n8413));
  jor  g08180(.dina(n8413), .dinb(n8298), .dout(n8414));
  jor  g08181(.dina(n8414), .dinb(asqrt[55] ), .dout(n8415));
  jnot g08182(.din(n8202), .dout(n8416));
  jand g08183(.dina(n8416), .dinb(n8415), .dout(n8417));
  jor  g08184(.dina(n8417), .dinb(n8297), .dout(n8418));
  jor  g08185(.dina(n8418), .dinb(asqrt[56] ), .dout(n8419));
  jand g08186(.dina(n8209), .dinb(n8419), .dout(n8420));
  jor  g08187(.dina(n8420), .dinb(n8296), .dout(n8421));
  jor  g08188(.dina(n8421), .dinb(asqrt[57] ), .dout(n8422));
  jnot g08189(.din(n8217), .dout(n8423));
  jand g08190(.dina(n8423), .dinb(n8422), .dout(n8424));
  jor  g08191(.dina(n8424), .dinb(n8295), .dout(n8425));
  jor  g08192(.dina(n8425), .dinb(asqrt[58] ), .dout(n8426));
  jand g08193(.dina(n8224), .dinb(n8426), .dout(n8427));
  jor  g08194(.dina(n8427), .dinb(n8294), .dout(n8428));
  jor  g08195(.dina(n8428), .dinb(asqrt[59] ), .dout(n8429));
  jand g08196(.dina(n8232), .dinb(n8429), .dout(n8430));
  jor  g08197(.dina(n8430), .dinb(n8293), .dout(n8431));
  jor  g08198(.dina(n8431), .dinb(asqrt[60] ), .dout(n8432));
  jnot g08199(.din(n8240), .dout(n8433));
  jand g08200(.dina(n8433), .dinb(n8432), .dout(n8434));
  jor  g08201(.dina(n8434), .dinb(n8292), .dout(n8435));
  jor  g08202(.dina(n8435), .dinb(asqrt[61] ), .dout(n8436));
  jnot g08203(.din(n8247), .dout(n8437));
  jand g08204(.dina(n8437), .dinb(n8436), .dout(n8438));
  jor  g08205(.dina(n8438), .dinb(n8291), .dout(n8439));
  jor  g08206(.dina(n8439), .dinb(asqrt[62] ), .dout(n8440));
  jand g08207(.dina(n8274), .dinb(n8440), .dout(n8441));
  jor  g08208(.dina(n8441), .dinb(n8290), .dout(n8442));
  jnot g08209(.din(n8259), .dout(n8443));
  jand g08210(.dina(n8443), .dinb(n8442), .dout(n8444));
  jand g08211(.dina(n8444), .dinb(n7820), .dout(n8445));
  jand g08212(.dina(n8445), .dinb(n8289), .dout(n8446));
  jor  g08213(.dina(n8446), .dinb(asqrt[63] ), .dout(n8447));
  jnot g08214(.din(n8272), .dout(n8448));
  jand g08215(.dina(n8448), .dinb(n8447), .dout(n8449));
  jor  g08216(.dina(n8449), .dinb(n8288), .dout(n8450));
  jand g08217(.dina(n8450), .dinb(n8287), .dout(n8451));
  jand g08218(.dina(n8451), .dinb(n8285), .dout(n8452));
  jor  g08219(.dina(n8452), .dinb(n8284), .dout(n8453));
  jand g08220(.dina(n8453), .dinb(asqrt[30] ), .dout(n8454));
  jor  g08221(.dina(n8453), .dinb(asqrt[30] ), .dout(n8455));
  jor  g08222(.dina(n8270), .dinb(n8265), .dout(n8456));
  jor  g08223(.dina(n8456), .dinb(n8263), .dout(n8457));
  jor  g08224(.dina(n8457), .dinb(n8003), .dout(n8458));
  jand g08225(.dina(n8458), .dinb(n8450), .dout(n8459));
  jxor g08226(.dina(n8459), .dinb(n7421), .dout(n8460));
  jnot g08227(.din(n8460), .dout(n8461));
  jand g08228(.dina(n8461), .dinb(n8455), .dout(n8462));
  jor  g08229(.dina(n8462), .dinb(n8454), .dout(n8463));
  jand g08230(.dina(n8463), .dinb(asqrt[31] ), .dout(n8464));
  jor  g08231(.dina(n8463), .dinb(asqrt[31] ), .dout(n8465));
  jxor g08232(.dina(n8005), .dinb(n7581), .dout(n8466));
  jand g08233(.dina(n8466), .dinb(asqrt[28] ), .dout(n8467));
  jxor g08234(.dina(n8467), .dinb(n8328), .dout(n8468));
  jand g08235(.dina(n8468), .dinb(n8465), .dout(n8469));
  jor  g08236(.dina(n8469), .dinb(n8464), .dout(n8470));
  jand g08237(.dina(n8470), .dinb(asqrt[32] ), .dout(n8471));
  jor  g08238(.dina(n8470), .dinb(asqrt[32] ), .dout(n8472));
  jxor g08239(.dina(n8013), .dinb(n7154), .dout(n8473));
  jand g08240(.dina(n8473), .dinb(asqrt[28] ), .dout(n8474));
  jxor g08241(.dina(n8474), .dinb(n8022), .dout(n8475));
  jnot g08242(.din(n8475), .dout(n8476));
  jand g08243(.dina(n8476), .dinb(n8472), .dout(n8477));
  jor  g08244(.dina(n8477), .dinb(n8471), .dout(n8478));
  jand g08245(.dina(n8478), .dinb(asqrt[33] ), .dout(n8479));
  jor  g08246(.dina(n8478), .dinb(asqrt[33] ), .dout(n8480));
  jxor g08247(.dina(n8024), .dinb(n6758), .dout(n8481));
  jand g08248(.dina(n8481), .dinb(asqrt[28] ), .dout(n8482));
  jxor g08249(.dina(n8482), .dinb(n8029), .dout(n8483));
  jnot g08250(.din(n8483), .dout(n8484));
  jand g08251(.dina(n8484), .dinb(n8480), .dout(n8485));
  jor  g08252(.dina(n8485), .dinb(n8479), .dout(n8486));
  jand g08253(.dina(n8486), .dinb(asqrt[34] ), .dout(n8487));
  jor  g08254(.dina(n8486), .dinb(asqrt[34] ), .dout(n8488));
  jxor g08255(.dina(n8031), .dinb(n6357), .dout(n8489));
  jand g08256(.dina(n8489), .dinb(asqrt[28] ), .dout(n8490));
  jxor g08257(.dina(n8490), .dinb(n8036), .dout(n8491));
  jnot g08258(.din(n8491), .dout(n8492));
  jand g08259(.dina(n8492), .dinb(n8488), .dout(n8493));
  jor  g08260(.dina(n8493), .dinb(n8487), .dout(n8494));
  jand g08261(.dina(n8494), .dinb(asqrt[35] ), .dout(n8495));
  jxor g08262(.dina(n8038), .dinb(n5989), .dout(n8496));
  jand g08263(.dina(n8496), .dinb(asqrt[28] ), .dout(n8497));
  jxor g08264(.dina(n8497), .dinb(n8042), .dout(n8498));
  jor  g08265(.dina(n8494), .dinb(asqrt[35] ), .dout(n8499));
  jand g08266(.dina(n8499), .dinb(n8498), .dout(n8500));
  jor  g08267(.dina(n8500), .dinb(n8495), .dout(n8501));
  jand g08268(.dina(n8501), .dinb(asqrt[36] ), .dout(n8502));
  jor  g08269(.dina(n8501), .dinb(asqrt[36] ), .dout(n8503));
  jxor g08270(.dina(n8046), .dinb(n5606), .dout(n8504));
  jand g08271(.dina(n8504), .dinb(asqrt[28] ), .dout(n8505));
  jxor g08272(.dina(n8505), .dinb(n8051), .dout(n8506));
  jnot g08273(.din(n8506), .dout(n8507));
  jand g08274(.dina(n8507), .dinb(n8503), .dout(n8508));
  jor  g08275(.dina(n8508), .dinb(n8502), .dout(n8509));
  jand g08276(.dina(n8509), .dinb(asqrt[37] ), .dout(n8510));
  jor  g08277(.dina(n8509), .dinb(asqrt[37] ), .dout(n8511));
  jxor g08278(.dina(n8053), .dinb(n5259), .dout(n8512));
  jand g08279(.dina(n8512), .dinb(asqrt[28] ), .dout(n8513));
  jxor g08280(.dina(n8513), .dinb(n8058), .dout(n8514));
  jand g08281(.dina(n8514), .dinb(n8511), .dout(n8515));
  jor  g08282(.dina(n8515), .dinb(n8510), .dout(n8516));
  jand g08283(.dina(n8516), .dinb(asqrt[38] ), .dout(n8517));
  jor  g08284(.dina(n8516), .dinb(asqrt[38] ), .dout(n8518));
  jxor g08285(.dina(n8061), .dinb(n4902), .dout(n8519));
  jand g08286(.dina(n8519), .dinb(asqrt[28] ), .dout(n8520));
  jxor g08287(.dina(n8520), .dinb(n8066), .dout(n8521));
  jnot g08288(.din(n8521), .dout(n8522));
  jand g08289(.dina(n8522), .dinb(n8518), .dout(n8523));
  jor  g08290(.dina(n8523), .dinb(n8517), .dout(n8524));
  jand g08291(.dina(n8524), .dinb(asqrt[39] ), .dout(n8525));
  jor  g08292(.dina(n8524), .dinb(asqrt[39] ), .dout(n8526));
  jxor g08293(.dina(n8068), .dinb(n4582), .dout(n8527));
  jand g08294(.dina(n8527), .dinb(asqrt[28] ), .dout(n8528));
  jxor g08295(.dina(n8528), .dinb(n8073), .dout(n8529));
  jand g08296(.dina(n8529), .dinb(n8526), .dout(n8530));
  jor  g08297(.dina(n8530), .dinb(n8525), .dout(n8531));
  jand g08298(.dina(n8531), .dinb(asqrt[40] ), .dout(n8532));
  jor  g08299(.dina(n8531), .dinb(asqrt[40] ), .dout(n8533));
  jxor g08300(.dina(n8076), .dinb(n4249), .dout(n8534));
  jand g08301(.dina(n8534), .dinb(asqrt[28] ), .dout(n8535));
  jxor g08302(.dina(n8535), .dinb(n8081), .dout(n8536));
  jand g08303(.dina(n8536), .dinb(n8533), .dout(n8537));
  jor  g08304(.dina(n8537), .dinb(n8532), .dout(n8538));
  jand g08305(.dina(n8538), .dinb(asqrt[41] ), .dout(n8539));
  jor  g08306(.dina(n8538), .dinb(asqrt[41] ), .dout(n8540));
  jxor g08307(.dina(n8084), .dinb(n3955), .dout(n8541));
  jand g08308(.dina(n8541), .dinb(asqrt[28] ), .dout(n8542));
  jxor g08309(.dina(n8542), .dinb(n8089), .dout(n8543));
  jand g08310(.dina(n8543), .dinb(n8540), .dout(n8544));
  jor  g08311(.dina(n8544), .dinb(n8539), .dout(n8545));
  jand g08312(.dina(n8545), .dinb(asqrt[42] ), .dout(n8546));
  jor  g08313(.dina(n8545), .dinb(asqrt[42] ), .dout(n8547));
  jxor g08314(.dina(n8092), .dinb(n3642), .dout(n8548));
  jand g08315(.dina(n8548), .dinb(asqrt[28] ), .dout(n8549));
  jxor g08316(.dina(n8549), .dinb(n8097), .dout(n8550));
  jnot g08317(.din(n8550), .dout(n8551));
  jand g08318(.dina(n8551), .dinb(n8547), .dout(n8552));
  jor  g08319(.dina(n8552), .dinb(n8546), .dout(n8553));
  jand g08320(.dina(n8553), .dinb(asqrt[43] ), .dout(n8554));
  jor  g08321(.dina(n8553), .dinb(asqrt[43] ), .dout(n8555));
  jxor g08322(.dina(n8099), .dinb(n3368), .dout(n8556));
  jand g08323(.dina(n8556), .dinb(asqrt[28] ), .dout(n8557));
  jxor g08324(.dina(n8557), .dinb(n8104), .dout(n8558));
  jand g08325(.dina(n8558), .dinb(n8555), .dout(n8559));
  jor  g08326(.dina(n8559), .dinb(n8554), .dout(n8560));
  jand g08327(.dina(n8560), .dinb(asqrt[44] ), .dout(n8561));
  jor  g08328(.dina(n8560), .dinb(asqrt[44] ), .dout(n8562));
  jxor g08329(.dina(n8107), .dinb(n3089), .dout(n8563));
  jand g08330(.dina(n8563), .dinb(asqrt[28] ), .dout(n8564));
  jxor g08331(.dina(n8564), .dinb(n8112), .dout(n8565));
  jnot g08332(.din(n8565), .dout(n8566));
  jand g08333(.dina(n8566), .dinb(n8562), .dout(n8567));
  jor  g08334(.dina(n8567), .dinb(n8561), .dout(n8568));
  jand g08335(.dina(n8568), .dinb(asqrt[45] ), .dout(n8569));
  jor  g08336(.dina(n8568), .dinb(asqrt[45] ), .dout(n8570));
  jxor g08337(.dina(n8114), .dinb(n2833), .dout(n8571));
  jand g08338(.dina(n8571), .dinb(asqrt[28] ), .dout(n8572));
  jxor g08339(.dina(n8572), .dinb(n8119), .dout(n8573));
  jand g08340(.dina(n8573), .dinb(n8570), .dout(n8574));
  jor  g08341(.dina(n8574), .dinb(n8569), .dout(n8575));
  jand g08342(.dina(n8575), .dinb(asqrt[46] ), .dout(n8576));
  jor  g08343(.dina(n8575), .dinb(asqrt[46] ), .dout(n8577));
  jxor g08344(.dina(n8122), .dinb(n2572), .dout(n8578));
  jand g08345(.dina(n8578), .dinb(asqrt[28] ), .dout(n8579));
  jxor g08346(.dina(n8579), .dinb(n8127), .dout(n8580));
  jnot g08347(.din(n8580), .dout(n8581));
  jand g08348(.dina(n8581), .dinb(n8577), .dout(n8582));
  jor  g08349(.dina(n8582), .dinb(n8576), .dout(n8583));
  jand g08350(.dina(n8583), .dinb(asqrt[47] ), .dout(n8584));
  jor  g08351(.dina(n8583), .dinb(asqrt[47] ), .dout(n8585));
  jxor g08352(.dina(n8129), .dinb(n2345), .dout(n8586));
  jand g08353(.dina(n8586), .dinb(asqrt[28] ), .dout(n8587));
  jxor g08354(.dina(n8587), .dinb(n8134), .dout(n8588));
  jand g08355(.dina(n8588), .dinb(n8585), .dout(n8589));
  jor  g08356(.dina(n8589), .dinb(n8584), .dout(n8590));
  jand g08357(.dina(n8590), .dinb(asqrt[48] ), .dout(n8591));
  jor  g08358(.dina(n8590), .dinb(asqrt[48] ), .dout(n8592));
  jxor g08359(.dina(n8137), .dinb(n2108), .dout(n8593));
  jand g08360(.dina(n8593), .dinb(asqrt[28] ), .dout(n8594));
  jxor g08361(.dina(n8594), .dinb(n8142), .dout(n8595));
  jnot g08362(.din(n8595), .dout(n8596));
  jand g08363(.dina(n8596), .dinb(n8592), .dout(n8597));
  jor  g08364(.dina(n8597), .dinb(n8591), .dout(n8598));
  jand g08365(.dina(n8598), .dinb(asqrt[49] ), .dout(n8599));
  jor  g08366(.dina(n8598), .dinb(asqrt[49] ), .dout(n8600));
  jxor g08367(.dina(n8144), .dinb(n1912), .dout(n8601));
  jand g08368(.dina(n8601), .dinb(asqrt[28] ), .dout(n8602));
  jxor g08369(.dina(n8602), .dinb(n8149), .dout(n8603));
  jand g08370(.dina(n8603), .dinb(n8600), .dout(n8604));
  jor  g08371(.dina(n8604), .dinb(n8599), .dout(n8605));
  jand g08372(.dina(n8605), .dinb(asqrt[50] ), .dout(n8606));
  jor  g08373(.dina(n8605), .dinb(asqrt[50] ), .dout(n8607));
  jxor g08374(.dina(n8152), .dinb(n1699), .dout(n8608));
  jand g08375(.dina(n8608), .dinb(asqrt[28] ), .dout(n8609));
  jxor g08376(.dina(n8609), .dinb(n8157), .dout(n8610));
  jand g08377(.dina(n8610), .dinb(n8607), .dout(n8611));
  jor  g08378(.dina(n8611), .dinb(n8606), .dout(n8612));
  jand g08379(.dina(n8612), .dinb(asqrt[51] ), .dout(n8613));
  jor  g08380(.dina(n8612), .dinb(asqrt[51] ), .dout(n8614));
  jxor g08381(.dina(n8160), .dinb(n1516), .dout(n8615));
  jand g08382(.dina(n8615), .dinb(asqrt[28] ), .dout(n8616));
  jxor g08383(.dina(n8616), .dinb(n8165), .dout(n8617));
  jand g08384(.dina(n8617), .dinb(n8614), .dout(n8618));
  jor  g08385(.dina(n8618), .dinb(n8613), .dout(n8619));
  jand g08386(.dina(n8619), .dinb(asqrt[52] ), .dout(n8620));
  jor  g08387(.dina(n8619), .dinb(asqrt[52] ), .dout(n8621));
  jxor g08388(.dina(n8168), .dinb(n1332), .dout(n8622));
  jand g08389(.dina(n8622), .dinb(asqrt[28] ), .dout(n8623));
  jxor g08390(.dina(n8623), .dinb(n8173), .dout(n8624));
  jnot g08391(.din(n8624), .dout(n8625));
  jand g08392(.dina(n8625), .dinb(n8621), .dout(n8626));
  jor  g08393(.dina(n8626), .dinb(n8620), .dout(n8627));
  jand g08394(.dina(n8627), .dinb(asqrt[53] ), .dout(n8628));
  jor  g08395(.dina(n8627), .dinb(asqrt[53] ), .dout(n8629));
  jxor g08396(.dina(n8175), .dinb(n1173), .dout(n8630));
  jand g08397(.dina(n8630), .dinb(asqrt[28] ), .dout(n8631));
  jxor g08398(.dina(n8631), .dinb(n8180), .dout(n8632));
  jnot g08399(.din(n8632), .dout(n8633));
  jand g08400(.dina(n8633), .dinb(n8629), .dout(n8634));
  jor  g08401(.dina(n8634), .dinb(n8628), .dout(n8635));
  jand g08402(.dina(n8635), .dinb(asqrt[54] ), .dout(n8636));
  jor  g08403(.dina(n8635), .dinb(asqrt[54] ), .dout(n8637));
  jxor g08404(.dina(n8182), .dinb(n1008), .dout(n8638));
  jand g08405(.dina(n8638), .dinb(asqrt[28] ), .dout(n8639));
  jxor g08406(.dina(n8639), .dinb(n8187), .dout(n8640));
  jnot g08407(.din(n8640), .dout(n8641));
  jand g08408(.dina(n8641), .dinb(n8637), .dout(n8642));
  jor  g08409(.dina(n8642), .dinb(n8636), .dout(n8643));
  jand g08410(.dina(n8643), .dinb(asqrt[55] ), .dout(n8644));
  jor  g08411(.dina(n8643), .dinb(asqrt[55] ), .dout(n8645));
  jxor g08412(.dina(n8189), .dinb(n884), .dout(n8646));
  jand g08413(.dina(n8646), .dinb(asqrt[28] ), .dout(n8647));
  jxor g08414(.dina(n8647), .dinb(n8194), .dout(n8648));
  jand g08415(.dina(n8648), .dinb(n8645), .dout(n8649));
  jor  g08416(.dina(n8649), .dinb(n8644), .dout(n8650));
  jand g08417(.dina(n8650), .dinb(asqrt[56] ), .dout(n8651));
  jor  g08418(.dina(n8650), .dinb(asqrt[56] ), .dout(n8652));
  jxor g08419(.dina(n8197), .dinb(n743), .dout(n8653));
  jand g08420(.dina(n8653), .dinb(asqrt[28] ), .dout(n8654));
  jxor g08421(.dina(n8654), .dinb(n8202), .dout(n8655));
  jnot g08422(.din(n8655), .dout(n8656));
  jand g08423(.dina(n8656), .dinb(n8652), .dout(n8657));
  jor  g08424(.dina(n8657), .dinb(n8651), .dout(n8658));
  jand g08425(.dina(n8658), .dinb(asqrt[57] ), .dout(n8659));
  jor  g08426(.dina(n8658), .dinb(asqrt[57] ), .dout(n8660));
  jxor g08427(.dina(n8204), .dinb(n635), .dout(n8661));
  jand g08428(.dina(n8661), .dinb(asqrt[28] ), .dout(n8662));
  jxor g08429(.dina(n8662), .dinb(n8209), .dout(n8663));
  jand g08430(.dina(n8663), .dinb(n8660), .dout(n8664));
  jor  g08431(.dina(n8664), .dinb(n8659), .dout(n8665));
  jand g08432(.dina(n8665), .dinb(asqrt[58] ), .dout(n8666));
  jor  g08433(.dina(n8665), .dinb(asqrt[58] ), .dout(n8667));
  jxor g08434(.dina(n8212), .dinb(n515), .dout(n8668));
  jand g08435(.dina(n8668), .dinb(asqrt[28] ), .dout(n8669));
  jxor g08436(.dina(n8669), .dinb(n8217), .dout(n8670));
  jnot g08437(.din(n8670), .dout(n8671));
  jand g08438(.dina(n8671), .dinb(n8667), .dout(n8672));
  jor  g08439(.dina(n8672), .dinb(n8666), .dout(n8673));
  jand g08440(.dina(n8673), .dinb(asqrt[59] ), .dout(n8674));
  jor  g08441(.dina(n8673), .dinb(asqrt[59] ), .dout(n8675));
  jxor g08442(.dina(n8219), .dinb(n443), .dout(n8676));
  jand g08443(.dina(n8676), .dinb(asqrt[28] ), .dout(n8677));
  jxor g08444(.dina(n8677), .dinb(n8224), .dout(n8678));
  jand g08445(.dina(n8678), .dinb(n8675), .dout(n8679));
  jor  g08446(.dina(n8679), .dinb(n8674), .dout(n8680));
  jand g08447(.dina(n8680), .dinb(asqrt[60] ), .dout(n8681));
  jor  g08448(.dina(n8680), .dinb(asqrt[60] ), .dout(n8682));
  jxor g08449(.dina(n8227), .dinb(n352), .dout(n8683));
  jand g08450(.dina(n8683), .dinb(asqrt[28] ), .dout(n8684));
  jxor g08451(.dina(n8684), .dinb(n8232), .dout(n8685));
  jand g08452(.dina(n8685), .dinb(n8682), .dout(n8686));
  jor  g08453(.dina(n8686), .dinb(n8681), .dout(n8687));
  jand g08454(.dina(n8687), .dinb(asqrt[61] ), .dout(n8688));
  jor  g08455(.dina(n8687), .dinb(asqrt[61] ), .dout(n8689));
  jxor g08456(.dina(n8235), .dinb(n294), .dout(n8690));
  jand g08457(.dina(n8690), .dinb(asqrt[28] ), .dout(n8691));
  jxor g08458(.dina(n8691), .dinb(n8240), .dout(n8692));
  jnot g08459(.din(n8692), .dout(n8693));
  jand g08460(.dina(n8693), .dinb(n8689), .dout(n8694));
  jor  g08461(.dina(n8694), .dinb(n8688), .dout(n8695));
  jand g08462(.dina(n8695), .dinb(asqrt[62] ), .dout(n8696));
  jor  g08463(.dina(n8695), .dinb(asqrt[62] ), .dout(n8697));
  jxor g08464(.dina(n8242), .dinb(n239), .dout(n8698));
  jand g08465(.dina(n8698), .dinb(asqrt[28] ), .dout(n8699));
  jxor g08466(.dina(n8699), .dinb(n8247), .dout(n8700));
  jnot g08467(.din(n8700), .dout(n8701));
  jand g08468(.dina(n8701), .dinb(n8697), .dout(n8702));
  jor  g08469(.dina(n8702), .dinb(n8696), .dout(n8703));
  jor  g08470(.dina(n8703), .dinb(n8277), .dout(n8704));
  jnot g08471(.din(n8704), .dout(n8705));
  jnot g08472(.din(n8277), .dout(n8707));
  jnot g08473(.din(n8696), .dout(n8708));
  jnot g08474(.din(n8688), .dout(n8709));
  jnot g08475(.din(n8681), .dout(n8710));
  jnot g08476(.din(n8674), .dout(n8711));
  jnot g08477(.din(n8666), .dout(n8712));
  jnot g08478(.din(n8659), .dout(n8713));
  jnot g08479(.din(n8651), .dout(n8714));
  jnot g08480(.din(n8644), .dout(n8715));
  jnot g08481(.din(n8636), .dout(n8716));
  jnot g08482(.din(n8628), .dout(n8717));
  jnot g08483(.din(n8620), .dout(n8718));
  jnot g08484(.din(n8613), .dout(n8719));
  jnot g08485(.din(n8606), .dout(n8720));
  jnot g08486(.din(n8599), .dout(n8721));
  jnot g08487(.din(n8591), .dout(n8722));
  jnot g08488(.din(n8584), .dout(n8723));
  jnot g08489(.din(n8576), .dout(n8724));
  jnot g08490(.din(n8569), .dout(n8725));
  jnot g08491(.din(n8561), .dout(n8726));
  jnot g08492(.din(n8554), .dout(n8727));
  jnot g08493(.din(n8546), .dout(n8728));
  jnot g08494(.din(n8539), .dout(n8729));
  jnot g08495(.din(n8532), .dout(n8730));
  jnot g08496(.din(n8525), .dout(n8731));
  jnot g08497(.din(n8517), .dout(n8732));
  jnot g08498(.din(n8510), .dout(n8733));
  jnot g08499(.din(n8502), .dout(n8734));
  jnot g08500(.din(n8495), .dout(n8735));
  jnot g08501(.din(n8498), .dout(n8736));
  jnot g08502(.din(n8487), .dout(n8737));
  jnot g08503(.din(n8479), .dout(n8738));
  jnot g08504(.din(n8471), .dout(n8739));
  jnot g08505(.din(n8464), .dout(n8740));
  jnot g08506(.din(n8454), .dout(n8741));
  jnot g08507(.din(n8284), .dout(n8742));
  jor  g08508(.dina(n8449), .dinb(n7991), .dout(n8743));
  jnot g08509(.din(n8282), .dout(n8744));
  jand g08510(.dina(n8744), .dinb(n8743), .dout(n8745));
  jand g08511(.dina(n8745), .dinb(n8003), .dout(n8746));
  jor  g08512(.dina(n8449), .dinb(a[56] ), .dout(n8747));
  jand g08513(.dina(n8747), .dinb(a[57] ), .dout(n8748));
  jand g08514(.dina(asqrt[28] ), .dinb(n7993), .dout(n8749));
  jor  g08515(.dina(n8749), .dinb(n8748), .dout(n8750));
  jor  g08516(.dina(n8750), .dinb(n8746), .dout(n8751));
  jand g08517(.dina(n8751), .dinb(n8742), .dout(n8752));
  jand g08518(.dina(n8752), .dinb(n7581), .dout(n8753));
  jor  g08519(.dina(n8460), .dinb(n8753), .dout(n8754));
  jand g08520(.dina(n8754), .dinb(n8741), .dout(n8755));
  jand g08521(.dina(n8755), .dinb(n7154), .dout(n8756));
  jnot g08522(.din(n8468), .dout(n8757));
  jor  g08523(.dina(n8757), .dinb(n8756), .dout(n8758));
  jand g08524(.dina(n8758), .dinb(n8740), .dout(n8759));
  jand g08525(.dina(n8759), .dinb(n6758), .dout(n8760));
  jor  g08526(.dina(n8475), .dinb(n8760), .dout(n8761));
  jand g08527(.dina(n8761), .dinb(n8739), .dout(n8762));
  jand g08528(.dina(n8762), .dinb(n6357), .dout(n8763));
  jor  g08529(.dina(n8483), .dinb(n8763), .dout(n8764));
  jand g08530(.dina(n8764), .dinb(n8738), .dout(n8765));
  jand g08531(.dina(n8765), .dinb(n5989), .dout(n8766));
  jor  g08532(.dina(n8491), .dinb(n8766), .dout(n8767));
  jand g08533(.dina(n8767), .dinb(n8737), .dout(n8768));
  jand g08534(.dina(n8768), .dinb(n5606), .dout(n8769));
  jor  g08535(.dina(n8769), .dinb(n8736), .dout(n8770));
  jand g08536(.dina(n8770), .dinb(n8735), .dout(n8771));
  jand g08537(.dina(n8771), .dinb(n5259), .dout(n8772));
  jor  g08538(.dina(n8506), .dinb(n8772), .dout(n8773));
  jand g08539(.dina(n8773), .dinb(n8734), .dout(n8774));
  jand g08540(.dina(n8774), .dinb(n4902), .dout(n8775));
  jnot g08541(.din(n8514), .dout(n8776));
  jor  g08542(.dina(n8776), .dinb(n8775), .dout(n8777));
  jand g08543(.dina(n8777), .dinb(n8733), .dout(n8778));
  jand g08544(.dina(n8778), .dinb(n4582), .dout(n8779));
  jor  g08545(.dina(n8521), .dinb(n8779), .dout(n8780));
  jand g08546(.dina(n8780), .dinb(n8732), .dout(n8781));
  jand g08547(.dina(n8781), .dinb(n4249), .dout(n8782));
  jnot g08548(.din(n8529), .dout(n8783));
  jor  g08549(.dina(n8783), .dinb(n8782), .dout(n8784));
  jand g08550(.dina(n8784), .dinb(n8731), .dout(n8785));
  jand g08551(.dina(n8785), .dinb(n3955), .dout(n8786));
  jnot g08552(.din(n8536), .dout(n8787));
  jor  g08553(.dina(n8787), .dinb(n8786), .dout(n8788));
  jand g08554(.dina(n8788), .dinb(n8730), .dout(n8789));
  jand g08555(.dina(n8789), .dinb(n3642), .dout(n8790));
  jnot g08556(.din(n8543), .dout(n8791));
  jor  g08557(.dina(n8791), .dinb(n8790), .dout(n8792));
  jand g08558(.dina(n8792), .dinb(n8729), .dout(n8793));
  jand g08559(.dina(n8793), .dinb(n3368), .dout(n8794));
  jor  g08560(.dina(n8550), .dinb(n8794), .dout(n8795));
  jand g08561(.dina(n8795), .dinb(n8728), .dout(n8796));
  jand g08562(.dina(n8796), .dinb(n3089), .dout(n8797));
  jnot g08563(.din(n8558), .dout(n8798));
  jor  g08564(.dina(n8798), .dinb(n8797), .dout(n8799));
  jand g08565(.dina(n8799), .dinb(n8727), .dout(n8800));
  jand g08566(.dina(n8800), .dinb(n2833), .dout(n8801));
  jor  g08567(.dina(n8565), .dinb(n8801), .dout(n8802));
  jand g08568(.dina(n8802), .dinb(n8726), .dout(n8803));
  jand g08569(.dina(n8803), .dinb(n2572), .dout(n8804));
  jnot g08570(.din(n8573), .dout(n8805));
  jor  g08571(.dina(n8805), .dinb(n8804), .dout(n8806));
  jand g08572(.dina(n8806), .dinb(n8725), .dout(n8807));
  jand g08573(.dina(n8807), .dinb(n2345), .dout(n8808));
  jor  g08574(.dina(n8580), .dinb(n8808), .dout(n8809));
  jand g08575(.dina(n8809), .dinb(n8724), .dout(n8810));
  jand g08576(.dina(n8810), .dinb(n2108), .dout(n8811));
  jnot g08577(.din(n8588), .dout(n8812));
  jor  g08578(.dina(n8812), .dinb(n8811), .dout(n8813));
  jand g08579(.dina(n8813), .dinb(n8723), .dout(n8814));
  jand g08580(.dina(n8814), .dinb(n1912), .dout(n8815));
  jor  g08581(.dina(n8595), .dinb(n8815), .dout(n8816));
  jand g08582(.dina(n8816), .dinb(n8722), .dout(n8817));
  jand g08583(.dina(n8817), .dinb(n1699), .dout(n8818));
  jnot g08584(.din(n8603), .dout(n8819));
  jor  g08585(.dina(n8819), .dinb(n8818), .dout(n8820));
  jand g08586(.dina(n8820), .dinb(n8721), .dout(n8821));
  jand g08587(.dina(n8821), .dinb(n1516), .dout(n8822));
  jnot g08588(.din(n8610), .dout(n8823));
  jor  g08589(.dina(n8823), .dinb(n8822), .dout(n8824));
  jand g08590(.dina(n8824), .dinb(n8720), .dout(n8825));
  jand g08591(.dina(n8825), .dinb(n1332), .dout(n8826));
  jnot g08592(.din(n8617), .dout(n8827));
  jor  g08593(.dina(n8827), .dinb(n8826), .dout(n8828));
  jand g08594(.dina(n8828), .dinb(n8719), .dout(n8829));
  jand g08595(.dina(n8829), .dinb(n1173), .dout(n8830));
  jor  g08596(.dina(n8624), .dinb(n8830), .dout(n8831));
  jand g08597(.dina(n8831), .dinb(n8718), .dout(n8832));
  jand g08598(.dina(n8832), .dinb(n1008), .dout(n8833));
  jor  g08599(.dina(n8632), .dinb(n8833), .dout(n8834));
  jand g08600(.dina(n8834), .dinb(n8717), .dout(n8835));
  jand g08601(.dina(n8835), .dinb(n884), .dout(n8836));
  jor  g08602(.dina(n8640), .dinb(n8836), .dout(n8837));
  jand g08603(.dina(n8837), .dinb(n8716), .dout(n8838));
  jand g08604(.dina(n8838), .dinb(n743), .dout(n8839));
  jnot g08605(.din(n8648), .dout(n8840));
  jor  g08606(.dina(n8840), .dinb(n8839), .dout(n8841));
  jand g08607(.dina(n8841), .dinb(n8715), .dout(n8842));
  jand g08608(.dina(n8842), .dinb(n635), .dout(n8843));
  jor  g08609(.dina(n8655), .dinb(n8843), .dout(n8844));
  jand g08610(.dina(n8844), .dinb(n8714), .dout(n8845));
  jand g08611(.dina(n8845), .dinb(n515), .dout(n8846));
  jnot g08612(.din(n8663), .dout(n8847));
  jor  g08613(.dina(n8847), .dinb(n8846), .dout(n8848));
  jand g08614(.dina(n8848), .dinb(n8713), .dout(n8849));
  jand g08615(.dina(n8849), .dinb(n443), .dout(n8850));
  jor  g08616(.dina(n8670), .dinb(n8850), .dout(n8851));
  jand g08617(.dina(n8851), .dinb(n8712), .dout(n8852));
  jand g08618(.dina(n8852), .dinb(n352), .dout(n8853));
  jnot g08619(.din(n8678), .dout(n8854));
  jor  g08620(.dina(n8854), .dinb(n8853), .dout(n8855));
  jand g08621(.dina(n8855), .dinb(n8711), .dout(n8856));
  jand g08622(.dina(n8856), .dinb(n294), .dout(n8857));
  jnot g08623(.din(n8685), .dout(n8858));
  jor  g08624(.dina(n8858), .dinb(n8857), .dout(n8859));
  jand g08625(.dina(n8859), .dinb(n8710), .dout(n8860));
  jand g08626(.dina(n8860), .dinb(n239), .dout(n8861));
  jor  g08627(.dina(n8692), .dinb(n8861), .dout(n8862));
  jand g08628(.dina(n8862), .dinb(n8709), .dout(n8863));
  jand g08629(.dina(n8863), .dinb(n221), .dout(n8864));
  jor  g08630(.dina(n8700), .dinb(n8864), .dout(n8865));
  jand g08631(.dina(n8865), .dinb(n8708), .dout(n8866));
  jor  g08632(.dina(n8866), .dinb(n8707), .dout(n8867));
  jand g08633(.dina(asqrt[28] ), .dinb(n8444), .dout(n8868));
  jor  g08634(.dina(n8868), .dinb(n8867), .dout(n8869));
  jor  g08635(.dina(n8869), .dinb(n8265), .dout(n8870));
  jand g08636(.dina(n8870), .dinb(n218), .dout(n8871));
  jand g08637(.dina(n8449), .dinb(n8256), .dout(n8872));
  jnot g08638(.din(n8872), .dout(n8873));
  jnot g08639(.din(n8265), .dout(n8874));
  jand g08640(.dina(n8260), .dinb(asqrt[63] ), .dout(n8875));
  jand g08641(.dina(n8875), .dinb(n8874), .dout(n8876));
  jand g08642(.dina(n8876), .dinb(n8873), .dout(n8877));
  jor  g08643(.dina(n8877), .dinb(n8871), .dout(n8878));
  jor  g08644(.dina(n8878), .dinb(n8705), .dout(asqrt[27] ));
  jand g08645(.dina(n8703), .dinb(n8277), .dout(n8882));
  jnot g08646(.din(n8868), .dout(n8883));
  jand g08647(.dina(n8883), .dinb(n8882), .dout(n8884));
  jand g08648(.dina(n8884), .dinb(n8874), .dout(n8885));
  jor  g08649(.dina(n8885), .dinb(asqrt[63] ), .dout(n8886));
  jnot g08650(.din(n8877), .dout(n8887));
  jand g08651(.dina(n8887), .dinb(n8886), .dout(n8888));
  jand g08652(.dina(n8888), .dinb(n8704), .dout(n8890));
  jxor g08653(.dina(n8695), .dinb(n221), .dout(n8891));
  jor  g08654(.dina(n8891), .dinb(n8890), .dout(n8892));
  jxor g08655(.dina(n8892), .dinb(n8700), .dout(n8893));
  jnot g08656(.din(n8893), .dout(n8894));
  jnot g08657(.din(a[52] ), .dout(n8895));
  jnot g08658(.din(a[53] ), .dout(n8896));
  jand g08659(.dina(n8896), .dinb(n8895), .dout(n8897));
  jand g08660(.dina(n8897), .dinb(n8279), .dout(n8898));
  jnot g08661(.din(n8898), .dout(n8899));
  jor  g08662(.dina(n8890), .dinb(n8279), .dout(n8900));
  jand g08663(.dina(n8900), .dinb(n8899), .dout(n8901));
  jor  g08664(.dina(n8901), .dinb(n8449), .dout(n8902));
  jand g08665(.dina(n8901), .dinb(n8449), .dout(n8903));
  jor  g08666(.dina(n8890), .dinb(a[54] ), .dout(n8904));
  jand g08667(.dina(n8904), .dinb(a[55] ), .dout(n8905));
  jand g08668(.dina(asqrt[27] ), .dinb(n8281), .dout(n8906));
  jor  g08669(.dina(n8906), .dinb(n8905), .dout(n8907));
  jor  g08670(.dina(n8907), .dinb(n8903), .dout(n8908));
  jand g08671(.dina(n8908), .dinb(n8902), .dout(n8909));
  jor  g08672(.dina(n8909), .dinb(n8003), .dout(n8910));
  jand g08673(.dina(n8909), .dinb(n8003), .dout(n8911));
  jnot g08674(.din(n8281), .dout(n8912));
  jor  g08675(.dina(n8890), .dinb(n8912), .dout(n8913));
  jor  g08676(.dina(n8705), .dinb(n8449), .dout(n8914));
  jor  g08677(.dina(n8914), .dinb(n8876), .dout(n8915));
  jor  g08678(.dina(n8915), .dinb(n8871), .dout(n8916));
  jand g08679(.dina(n8916), .dinb(n8913), .dout(n8917));
  jxor g08680(.dina(n8917), .dinb(n7991), .dout(n8918));
  jor  g08681(.dina(n8918), .dinb(n8911), .dout(n8919));
  jand g08682(.dina(n8919), .dinb(n8910), .dout(n8920));
  jor  g08683(.dina(n8920), .dinb(n7581), .dout(n8921));
  jand g08684(.dina(n8920), .dinb(n7581), .dout(n8922));
  jxor g08685(.dina(n8283), .dinb(n8003), .dout(n8923));
  jor  g08686(.dina(n8923), .dinb(n8890), .dout(n8924));
  jxor g08687(.dina(n8924), .dinb(n8750), .dout(n8925));
  jnot g08688(.din(n8925), .dout(n8926));
  jor  g08689(.dina(n8926), .dinb(n8922), .dout(n8927));
  jand g08690(.dina(n8927), .dinb(n8921), .dout(n8928));
  jor  g08691(.dina(n8928), .dinb(n7154), .dout(n8929));
  jand g08692(.dina(n8928), .dinb(n7154), .dout(n8930));
  jxor g08693(.dina(n8453), .dinb(n7581), .dout(n8931));
  jor  g08694(.dina(n8931), .dinb(n8890), .dout(n8932));
  jxor g08695(.dina(n8932), .dinb(n8461), .dout(n8933));
  jor  g08696(.dina(n8933), .dinb(n8930), .dout(n8934));
  jand g08697(.dina(n8934), .dinb(n8929), .dout(n8935));
  jor  g08698(.dina(n8935), .dinb(n6758), .dout(n8936));
  jand g08699(.dina(n8935), .dinb(n6758), .dout(n8937));
  jxor g08700(.dina(n8463), .dinb(n7154), .dout(n8938));
  jor  g08701(.dina(n8938), .dinb(n8890), .dout(n8939));
  jxor g08702(.dina(n8939), .dinb(n8468), .dout(n8940));
  jor  g08703(.dina(n8940), .dinb(n8937), .dout(n8941));
  jand g08704(.dina(n8941), .dinb(n8936), .dout(n8942));
  jor  g08705(.dina(n8942), .dinb(n6357), .dout(n8943));
  jand g08706(.dina(n8942), .dinb(n6357), .dout(n8944));
  jxor g08707(.dina(n8470), .dinb(n6758), .dout(n8945));
  jor  g08708(.dina(n8945), .dinb(n8890), .dout(n8946));
  jxor g08709(.dina(n8946), .dinb(n8476), .dout(n8947));
  jor  g08710(.dina(n8947), .dinb(n8944), .dout(n8948));
  jand g08711(.dina(n8948), .dinb(n8943), .dout(n8949));
  jor  g08712(.dina(n8949), .dinb(n5989), .dout(n8950));
  jand g08713(.dina(n8949), .dinb(n5989), .dout(n8951));
  jxor g08714(.dina(n8478), .dinb(n6357), .dout(n8952));
  jor  g08715(.dina(n8952), .dinb(n8890), .dout(n8953));
  jxor g08716(.dina(n8953), .dinb(n8484), .dout(n8954));
  jor  g08717(.dina(n8954), .dinb(n8951), .dout(n8955));
  jand g08718(.dina(n8955), .dinb(n8950), .dout(n8956));
  jor  g08719(.dina(n8956), .dinb(n5606), .dout(n8957));
  jand g08720(.dina(n8956), .dinb(n5606), .dout(n8958));
  jxor g08721(.dina(n8486), .dinb(n5989), .dout(n8959));
  jor  g08722(.dina(n8959), .dinb(n8890), .dout(n8960));
  jxor g08723(.dina(n8960), .dinb(n8492), .dout(n8961));
  jor  g08724(.dina(n8961), .dinb(n8958), .dout(n8962));
  jand g08725(.dina(n8962), .dinb(n8957), .dout(n8963));
  jor  g08726(.dina(n8963), .dinb(n5259), .dout(n8964));
  jxor g08727(.dina(n8494), .dinb(n5606), .dout(n8965));
  jor  g08728(.dina(n8965), .dinb(n8890), .dout(n8966));
  jxor g08729(.dina(n8966), .dinb(n8736), .dout(n8967));
  jnot g08730(.din(n8967), .dout(n8968));
  jand g08731(.dina(n8963), .dinb(n5259), .dout(n8969));
  jor  g08732(.dina(n8969), .dinb(n8968), .dout(n8970));
  jand g08733(.dina(n8970), .dinb(n8964), .dout(n8971));
  jor  g08734(.dina(n8971), .dinb(n4902), .dout(n8972));
  jand g08735(.dina(n8971), .dinb(n4902), .dout(n8973));
  jxor g08736(.dina(n8501), .dinb(n5259), .dout(n8974));
  jor  g08737(.dina(n8974), .dinb(n8890), .dout(n8975));
  jxor g08738(.dina(n8975), .dinb(n8507), .dout(n8976));
  jor  g08739(.dina(n8976), .dinb(n8973), .dout(n8977));
  jand g08740(.dina(n8977), .dinb(n8972), .dout(n8978));
  jor  g08741(.dina(n8978), .dinb(n4582), .dout(n8979));
  jand g08742(.dina(n8978), .dinb(n4582), .dout(n8980));
  jxor g08743(.dina(n8509), .dinb(n4902), .dout(n8981));
  jor  g08744(.dina(n8981), .dinb(n8890), .dout(n8982));
  jxor g08745(.dina(n8982), .dinb(n8776), .dout(n8983));
  jnot g08746(.din(n8983), .dout(n8984));
  jor  g08747(.dina(n8984), .dinb(n8980), .dout(n8985));
  jand g08748(.dina(n8985), .dinb(n8979), .dout(n8986));
  jor  g08749(.dina(n8986), .dinb(n4249), .dout(n8987));
  jand g08750(.dina(n8986), .dinb(n4249), .dout(n8988));
  jxor g08751(.dina(n8516), .dinb(n4582), .dout(n8989));
  jor  g08752(.dina(n8989), .dinb(n8890), .dout(n8990));
  jxor g08753(.dina(n8990), .dinb(n8522), .dout(n8991));
  jor  g08754(.dina(n8991), .dinb(n8988), .dout(n8992));
  jand g08755(.dina(n8992), .dinb(n8987), .dout(n8993));
  jor  g08756(.dina(n8993), .dinb(n3955), .dout(n8994));
  jand g08757(.dina(n8993), .dinb(n3955), .dout(n8995));
  jxor g08758(.dina(n8524), .dinb(n4249), .dout(n8996));
  jor  g08759(.dina(n8996), .dinb(n8890), .dout(n8997));
  jxor g08760(.dina(n8997), .dinb(n8783), .dout(n8998));
  jnot g08761(.din(n8998), .dout(n8999));
  jor  g08762(.dina(n8999), .dinb(n8995), .dout(n9000));
  jand g08763(.dina(n9000), .dinb(n8994), .dout(n9001));
  jor  g08764(.dina(n9001), .dinb(n3642), .dout(n9002));
  jand g08765(.dina(n9001), .dinb(n3642), .dout(n9003));
  jxor g08766(.dina(n8531), .dinb(n3955), .dout(n9004));
  jor  g08767(.dina(n9004), .dinb(n8890), .dout(n9005));
  jxor g08768(.dina(n9005), .dinb(n8787), .dout(n9006));
  jnot g08769(.din(n9006), .dout(n9007));
  jor  g08770(.dina(n9007), .dinb(n9003), .dout(n9008));
  jand g08771(.dina(n9008), .dinb(n9002), .dout(n9009));
  jor  g08772(.dina(n9009), .dinb(n3368), .dout(n9010));
  jand g08773(.dina(n9009), .dinb(n3368), .dout(n9011));
  jxor g08774(.dina(n8538), .dinb(n3642), .dout(n9012));
  jor  g08775(.dina(n9012), .dinb(n8890), .dout(n9013));
  jxor g08776(.dina(n9013), .dinb(n8791), .dout(n9014));
  jnot g08777(.din(n9014), .dout(n9015));
  jor  g08778(.dina(n9015), .dinb(n9011), .dout(n9016));
  jand g08779(.dina(n9016), .dinb(n9010), .dout(n9017));
  jor  g08780(.dina(n9017), .dinb(n3089), .dout(n9018));
  jand g08781(.dina(n9017), .dinb(n3089), .dout(n9019));
  jxor g08782(.dina(n8545), .dinb(n3368), .dout(n9020));
  jor  g08783(.dina(n9020), .dinb(n8890), .dout(n9021));
  jxor g08784(.dina(n9021), .dinb(n8551), .dout(n9022));
  jor  g08785(.dina(n9022), .dinb(n9019), .dout(n9023));
  jand g08786(.dina(n9023), .dinb(n9018), .dout(n9024));
  jor  g08787(.dina(n9024), .dinb(n2833), .dout(n9025));
  jand g08788(.dina(n9024), .dinb(n2833), .dout(n9026));
  jxor g08789(.dina(n8553), .dinb(n3089), .dout(n9027));
  jor  g08790(.dina(n9027), .dinb(n8890), .dout(n9028));
  jxor g08791(.dina(n9028), .dinb(n8798), .dout(n9029));
  jnot g08792(.din(n9029), .dout(n9030));
  jor  g08793(.dina(n9030), .dinb(n9026), .dout(n9031));
  jand g08794(.dina(n9031), .dinb(n9025), .dout(n9032));
  jor  g08795(.dina(n9032), .dinb(n2572), .dout(n9033));
  jand g08796(.dina(n9032), .dinb(n2572), .dout(n9034));
  jxor g08797(.dina(n8560), .dinb(n2833), .dout(n9035));
  jor  g08798(.dina(n9035), .dinb(n8890), .dout(n9036));
  jxor g08799(.dina(n9036), .dinb(n8566), .dout(n9037));
  jor  g08800(.dina(n9037), .dinb(n9034), .dout(n9038));
  jand g08801(.dina(n9038), .dinb(n9033), .dout(n9039));
  jor  g08802(.dina(n9039), .dinb(n2345), .dout(n9040));
  jand g08803(.dina(n9039), .dinb(n2345), .dout(n9041));
  jxor g08804(.dina(n8568), .dinb(n2572), .dout(n9042));
  jor  g08805(.dina(n9042), .dinb(n8890), .dout(n9043));
  jxor g08806(.dina(n9043), .dinb(n8805), .dout(n9044));
  jnot g08807(.din(n9044), .dout(n9045));
  jor  g08808(.dina(n9045), .dinb(n9041), .dout(n9046));
  jand g08809(.dina(n9046), .dinb(n9040), .dout(n9047));
  jor  g08810(.dina(n9047), .dinb(n2108), .dout(n9048));
  jand g08811(.dina(n9047), .dinb(n2108), .dout(n9049));
  jxor g08812(.dina(n8575), .dinb(n2345), .dout(n9050));
  jor  g08813(.dina(n9050), .dinb(n8890), .dout(n9051));
  jxor g08814(.dina(n9051), .dinb(n8581), .dout(n9052));
  jor  g08815(.dina(n9052), .dinb(n9049), .dout(n9053));
  jand g08816(.dina(n9053), .dinb(n9048), .dout(n9054));
  jor  g08817(.dina(n9054), .dinb(n1912), .dout(n9055));
  jand g08818(.dina(n9054), .dinb(n1912), .dout(n9056));
  jxor g08819(.dina(n8583), .dinb(n2108), .dout(n9057));
  jor  g08820(.dina(n9057), .dinb(n8890), .dout(n9058));
  jxor g08821(.dina(n9058), .dinb(n8812), .dout(n9059));
  jnot g08822(.din(n9059), .dout(n9060));
  jor  g08823(.dina(n9060), .dinb(n9056), .dout(n9061));
  jand g08824(.dina(n9061), .dinb(n9055), .dout(n9062));
  jor  g08825(.dina(n9062), .dinb(n1699), .dout(n9063));
  jand g08826(.dina(n9062), .dinb(n1699), .dout(n9064));
  jxor g08827(.dina(n8590), .dinb(n1912), .dout(n9065));
  jor  g08828(.dina(n9065), .dinb(n8890), .dout(n9066));
  jxor g08829(.dina(n9066), .dinb(n8596), .dout(n9067));
  jor  g08830(.dina(n9067), .dinb(n9064), .dout(n9068));
  jand g08831(.dina(n9068), .dinb(n9063), .dout(n9069));
  jor  g08832(.dina(n9069), .dinb(n1516), .dout(n9070));
  jand g08833(.dina(n9069), .dinb(n1516), .dout(n9071));
  jxor g08834(.dina(n8598), .dinb(n1699), .dout(n9072));
  jor  g08835(.dina(n9072), .dinb(n8890), .dout(n9073));
  jxor g08836(.dina(n9073), .dinb(n8819), .dout(n9074));
  jnot g08837(.din(n9074), .dout(n9075));
  jor  g08838(.dina(n9075), .dinb(n9071), .dout(n9076));
  jand g08839(.dina(n9076), .dinb(n9070), .dout(n9077));
  jor  g08840(.dina(n9077), .dinb(n1332), .dout(n9078));
  jand g08841(.dina(n9077), .dinb(n1332), .dout(n9079));
  jxor g08842(.dina(n8605), .dinb(n1516), .dout(n9080));
  jor  g08843(.dina(n9080), .dinb(n8890), .dout(n9081));
  jxor g08844(.dina(n9081), .dinb(n8823), .dout(n9082));
  jnot g08845(.din(n9082), .dout(n9083));
  jor  g08846(.dina(n9083), .dinb(n9079), .dout(n9084));
  jand g08847(.dina(n9084), .dinb(n9078), .dout(n9085));
  jor  g08848(.dina(n9085), .dinb(n1173), .dout(n9086));
  jand g08849(.dina(n9085), .dinb(n1173), .dout(n9087));
  jxor g08850(.dina(n8612), .dinb(n1332), .dout(n9088));
  jor  g08851(.dina(n9088), .dinb(n8890), .dout(n9089));
  jxor g08852(.dina(n9089), .dinb(n8827), .dout(n9090));
  jnot g08853(.din(n9090), .dout(n9091));
  jor  g08854(.dina(n9091), .dinb(n9087), .dout(n9092));
  jand g08855(.dina(n9092), .dinb(n9086), .dout(n9093));
  jor  g08856(.dina(n9093), .dinb(n1008), .dout(n9094));
  jand g08857(.dina(n9093), .dinb(n1008), .dout(n9095));
  jxor g08858(.dina(n8619), .dinb(n1173), .dout(n9096));
  jor  g08859(.dina(n9096), .dinb(n8890), .dout(n9097));
  jxor g08860(.dina(n9097), .dinb(n8625), .dout(n9098));
  jor  g08861(.dina(n9098), .dinb(n9095), .dout(n9099));
  jand g08862(.dina(n9099), .dinb(n9094), .dout(n9100));
  jor  g08863(.dina(n9100), .dinb(n884), .dout(n9101));
  jand g08864(.dina(n9100), .dinb(n884), .dout(n9102));
  jxor g08865(.dina(n8627), .dinb(n1008), .dout(n9103));
  jor  g08866(.dina(n9103), .dinb(n8890), .dout(n9104));
  jxor g08867(.dina(n9104), .dinb(n8633), .dout(n9105));
  jor  g08868(.dina(n9105), .dinb(n9102), .dout(n9106));
  jand g08869(.dina(n9106), .dinb(n9101), .dout(n9107));
  jor  g08870(.dina(n9107), .dinb(n743), .dout(n9108));
  jand g08871(.dina(n9107), .dinb(n743), .dout(n9109));
  jxor g08872(.dina(n8635), .dinb(n884), .dout(n9110));
  jor  g08873(.dina(n9110), .dinb(n8890), .dout(n9111));
  jxor g08874(.dina(n9111), .dinb(n8641), .dout(n9112));
  jor  g08875(.dina(n9112), .dinb(n9109), .dout(n9113));
  jand g08876(.dina(n9113), .dinb(n9108), .dout(n9114));
  jor  g08877(.dina(n9114), .dinb(n635), .dout(n9115));
  jand g08878(.dina(n9114), .dinb(n635), .dout(n9116));
  jxor g08879(.dina(n8643), .dinb(n743), .dout(n9117));
  jor  g08880(.dina(n9117), .dinb(n8890), .dout(n9118));
  jxor g08881(.dina(n9118), .dinb(n8840), .dout(n9119));
  jnot g08882(.din(n9119), .dout(n9120));
  jor  g08883(.dina(n9120), .dinb(n9116), .dout(n9121));
  jand g08884(.dina(n9121), .dinb(n9115), .dout(n9122));
  jor  g08885(.dina(n9122), .dinb(n515), .dout(n9123));
  jand g08886(.dina(n9122), .dinb(n515), .dout(n9124));
  jxor g08887(.dina(n8650), .dinb(n635), .dout(n9125));
  jor  g08888(.dina(n9125), .dinb(n8890), .dout(n9126));
  jxor g08889(.dina(n9126), .dinb(n8656), .dout(n9127));
  jor  g08890(.dina(n9127), .dinb(n9124), .dout(n9128));
  jand g08891(.dina(n9128), .dinb(n9123), .dout(n9129));
  jor  g08892(.dina(n9129), .dinb(n443), .dout(n9130));
  jand g08893(.dina(n9129), .dinb(n443), .dout(n9131));
  jxor g08894(.dina(n8658), .dinb(n515), .dout(n9132));
  jor  g08895(.dina(n9132), .dinb(n8890), .dout(n9133));
  jxor g08896(.dina(n9133), .dinb(n8847), .dout(n9134));
  jnot g08897(.din(n9134), .dout(n9135));
  jor  g08898(.dina(n9135), .dinb(n9131), .dout(n9136));
  jand g08899(.dina(n9136), .dinb(n9130), .dout(n9137));
  jor  g08900(.dina(n9137), .dinb(n352), .dout(n9138));
  jand g08901(.dina(n9137), .dinb(n352), .dout(n9139));
  jxor g08902(.dina(n8665), .dinb(n443), .dout(n9140));
  jor  g08903(.dina(n9140), .dinb(n8890), .dout(n9141));
  jxor g08904(.dina(n9141), .dinb(n8671), .dout(n9142));
  jor  g08905(.dina(n9142), .dinb(n9139), .dout(n9143));
  jand g08906(.dina(n9143), .dinb(n9138), .dout(n9144));
  jor  g08907(.dina(n9144), .dinb(n294), .dout(n9145));
  jand g08908(.dina(n9144), .dinb(n294), .dout(n9146));
  jxor g08909(.dina(n8673), .dinb(n352), .dout(n9147));
  jor  g08910(.dina(n9147), .dinb(n8890), .dout(n9148));
  jxor g08911(.dina(n9148), .dinb(n8854), .dout(n9149));
  jnot g08912(.din(n9149), .dout(n9150));
  jor  g08913(.dina(n9150), .dinb(n9146), .dout(n9151));
  jand g08914(.dina(n9151), .dinb(n9145), .dout(n9152));
  jor  g08915(.dina(n9152), .dinb(n239), .dout(n9153));
  jand g08916(.dina(n9152), .dinb(n239), .dout(n9154));
  jxor g08917(.dina(n8680), .dinb(n294), .dout(n9155));
  jor  g08918(.dina(n9155), .dinb(n8890), .dout(n9156));
  jxor g08919(.dina(n9156), .dinb(n8858), .dout(n9157));
  jnot g08920(.din(n9157), .dout(n9158));
  jor  g08921(.dina(n9158), .dinb(n9154), .dout(n9159));
  jand g08922(.dina(n9159), .dinb(n9153), .dout(n9160));
  jor  g08923(.dina(n9160), .dinb(n221), .dout(n9161));
  jand g08924(.dina(n9160), .dinb(n221), .dout(n9162));
  jxor g08925(.dina(n8687), .dinb(n239), .dout(n9163));
  jor  g08926(.dina(n9163), .dinb(n8890), .dout(n9164));
  jxor g08927(.dina(n9164), .dinb(n8693), .dout(n9165));
  jor  g08928(.dina(n9165), .dinb(n9162), .dout(n9166));
  jand g08929(.dina(n9166), .dinb(n9161), .dout(n9167));
  jand g08930(.dina(n9167), .dinb(n8894), .dout(n9168));
  jand g08931(.dina(n8888), .dinb(n8866), .dout(n9169));
  jand g08932(.dina(n8867), .dinb(asqrt[63] ), .dout(n9170));
  jand g08933(.dina(n9170), .dinb(n8704), .dout(n9171));
  jnot g08934(.din(n9171), .dout(n9172));
  jor  g08935(.dina(n9172), .dinb(n9169), .dout(n9173));
  jnot g08936(.din(n9173), .dout(n9174));
  jor  g08937(.dina(n9167), .dinb(n8894), .dout(n9175));
  jand g08938(.dina(n8878), .dinb(n8882), .dout(n9176));
  jor  g08939(.dina(n9176), .dinb(n8705), .dout(n9177));
  jor  g08940(.dina(n9177), .dinb(n9175), .dout(n9178));
  jand g08941(.dina(n9178), .dinb(n218), .dout(n9179));
  jand g08942(.dina(n8890), .dinb(n8707), .dout(n9180));
  jor  g08943(.dina(n9180), .dinb(n9179), .dout(n9181));
  jor  g08944(.dina(n9181), .dinb(n9174), .dout(n9182));
  jor  g08945(.dina(n9182), .dinb(n9168), .dout(asqrt[26] ));
  jnot g08946(.din(n9165), .dout(n9184));
  jxor g08947(.dina(n9160), .dinb(n221), .dout(n9185));
  jand g08948(.dina(n9185), .dinb(asqrt[26] ), .dout(n9186));
  jxor g08949(.dina(n9186), .dinb(n9184), .dout(n9187));
  jnot g08950(.din(a[50] ), .dout(n9188));
  jnot g08951(.din(a[51] ), .dout(n9189));
  jand g08952(.dina(n9189), .dinb(n9188), .dout(n9190));
  jand g08953(.dina(n9190), .dinb(n8895), .dout(n9191));
  jand g08954(.dina(asqrt[26] ), .dinb(a[52] ), .dout(n9192));
  jor  g08955(.dina(n9192), .dinb(n9191), .dout(n9193));
  jand g08956(.dina(n9193), .dinb(asqrt[27] ), .dout(n9194));
  jor  g08957(.dina(n9193), .dinb(asqrt[27] ), .dout(n9195));
  jand g08958(.dina(asqrt[26] ), .dinb(n8895), .dout(n9196));
  jor  g08959(.dina(n9196), .dinb(n8896), .dout(n9197));
  jnot g08960(.din(n8897), .dout(n9198));
  jnot g08961(.din(n9168), .dout(n9199));
  jnot g08962(.din(n9161), .dout(n9200));
  jnot g08963(.din(n9153), .dout(n9201));
  jnot g08964(.din(n9145), .dout(n9202));
  jnot g08965(.din(n9138), .dout(n9203));
  jnot g08966(.din(n9130), .dout(n9204));
  jnot g08967(.din(n9123), .dout(n9205));
  jnot g08968(.din(n9115), .dout(n9206));
  jnot g08969(.din(n9108), .dout(n9207));
  jnot g08970(.din(n9101), .dout(n9208));
  jnot g08971(.din(n9094), .dout(n9209));
  jnot g08972(.din(n9086), .dout(n9210));
  jnot g08973(.din(n9078), .dout(n9211));
  jnot g08974(.din(n9070), .dout(n9212));
  jnot g08975(.din(n9063), .dout(n9213));
  jnot g08976(.din(n9055), .dout(n9214));
  jnot g08977(.din(n9048), .dout(n9215));
  jnot g08978(.din(n9040), .dout(n9216));
  jnot g08979(.din(n9033), .dout(n9217));
  jnot g08980(.din(n9025), .dout(n9218));
  jnot g08981(.din(n9018), .dout(n9219));
  jnot g08982(.din(n9010), .dout(n9220));
  jnot g08983(.din(n9002), .dout(n9221));
  jnot g08984(.din(n8994), .dout(n9222));
  jnot g08985(.din(n8987), .dout(n9223));
  jnot g08986(.din(n8979), .dout(n9224));
  jnot g08987(.din(n8972), .dout(n9225));
  jnot g08988(.din(n8964), .dout(n9226));
  jnot g08989(.din(n8957), .dout(n9227));
  jnot g08990(.din(n8950), .dout(n9228));
  jnot g08991(.din(n8943), .dout(n9229));
  jnot g08992(.din(n8936), .dout(n9230));
  jnot g08993(.din(n8929), .dout(n9231));
  jnot g08994(.din(n8921), .dout(n9232));
  jnot g08995(.din(n8910), .dout(n9233));
  jnot g08996(.din(n8902), .dout(n9234));
  jand g08997(.dina(asqrt[27] ), .dinb(a[54] ), .dout(n9235));
  jor  g08998(.dina(n9235), .dinb(n8898), .dout(n9236));
  jor  g08999(.dina(n9236), .dinb(asqrt[28] ), .dout(n9237));
  jand g09000(.dina(asqrt[27] ), .dinb(n8279), .dout(n9238));
  jor  g09001(.dina(n9238), .dinb(n8280), .dout(n9239));
  jand g09002(.dina(n8913), .dinb(n9239), .dout(n9240));
  jand g09003(.dina(n9240), .dinb(n9237), .dout(n9241));
  jor  g09004(.dina(n9241), .dinb(n9234), .dout(n9242));
  jor  g09005(.dina(n9242), .dinb(asqrt[29] ), .dout(n9243));
  jnot g09006(.din(n8918), .dout(n9244));
  jand g09007(.dina(n9244), .dinb(n9243), .dout(n9245));
  jor  g09008(.dina(n9245), .dinb(n9233), .dout(n9246));
  jor  g09009(.dina(n9246), .dinb(asqrt[30] ), .dout(n9247));
  jand g09010(.dina(n8925), .dinb(n9247), .dout(n9248));
  jor  g09011(.dina(n9248), .dinb(n9232), .dout(n9249));
  jor  g09012(.dina(n9249), .dinb(asqrt[31] ), .dout(n9250));
  jnot g09013(.din(n8933), .dout(n9251));
  jand g09014(.dina(n9251), .dinb(n9250), .dout(n9252));
  jor  g09015(.dina(n9252), .dinb(n9231), .dout(n9253));
  jor  g09016(.dina(n9253), .dinb(asqrt[32] ), .dout(n9254));
  jnot g09017(.din(n8940), .dout(n9255));
  jand g09018(.dina(n9255), .dinb(n9254), .dout(n9256));
  jor  g09019(.dina(n9256), .dinb(n9230), .dout(n9257));
  jor  g09020(.dina(n9257), .dinb(asqrt[33] ), .dout(n9258));
  jnot g09021(.din(n8947), .dout(n9259));
  jand g09022(.dina(n9259), .dinb(n9258), .dout(n9260));
  jor  g09023(.dina(n9260), .dinb(n9229), .dout(n9261));
  jor  g09024(.dina(n9261), .dinb(asqrt[34] ), .dout(n9262));
  jnot g09025(.din(n8954), .dout(n9263));
  jand g09026(.dina(n9263), .dinb(n9262), .dout(n9264));
  jor  g09027(.dina(n9264), .dinb(n9228), .dout(n9265));
  jor  g09028(.dina(n9265), .dinb(asqrt[35] ), .dout(n9266));
  jnot g09029(.din(n8961), .dout(n9267));
  jand g09030(.dina(n9267), .dinb(n9266), .dout(n9268));
  jor  g09031(.dina(n9268), .dinb(n9227), .dout(n9269));
  jor  g09032(.dina(n9269), .dinb(asqrt[36] ), .dout(n9270));
  jand g09033(.dina(n9270), .dinb(n8967), .dout(n9271));
  jor  g09034(.dina(n9271), .dinb(n9226), .dout(n9272));
  jor  g09035(.dina(n9272), .dinb(asqrt[37] ), .dout(n9273));
  jnot g09036(.din(n8976), .dout(n9274));
  jand g09037(.dina(n9274), .dinb(n9273), .dout(n9275));
  jor  g09038(.dina(n9275), .dinb(n9225), .dout(n9276));
  jor  g09039(.dina(n9276), .dinb(asqrt[38] ), .dout(n9277));
  jand g09040(.dina(n8983), .dinb(n9277), .dout(n9278));
  jor  g09041(.dina(n9278), .dinb(n9224), .dout(n9279));
  jor  g09042(.dina(n9279), .dinb(asqrt[39] ), .dout(n9280));
  jnot g09043(.din(n8991), .dout(n9281));
  jand g09044(.dina(n9281), .dinb(n9280), .dout(n9282));
  jor  g09045(.dina(n9282), .dinb(n9223), .dout(n9283));
  jor  g09046(.dina(n9283), .dinb(asqrt[40] ), .dout(n9284));
  jand g09047(.dina(n8998), .dinb(n9284), .dout(n9285));
  jor  g09048(.dina(n9285), .dinb(n9222), .dout(n9286));
  jor  g09049(.dina(n9286), .dinb(asqrt[41] ), .dout(n9287));
  jand g09050(.dina(n9006), .dinb(n9287), .dout(n9288));
  jor  g09051(.dina(n9288), .dinb(n9221), .dout(n9289));
  jor  g09052(.dina(n9289), .dinb(asqrt[42] ), .dout(n9290));
  jand g09053(.dina(n9014), .dinb(n9290), .dout(n9291));
  jor  g09054(.dina(n9291), .dinb(n9220), .dout(n9292));
  jor  g09055(.dina(n9292), .dinb(asqrt[43] ), .dout(n9293));
  jnot g09056(.din(n9022), .dout(n9294));
  jand g09057(.dina(n9294), .dinb(n9293), .dout(n9295));
  jor  g09058(.dina(n9295), .dinb(n9219), .dout(n9296));
  jor  g09059(.dina(n9296), .dinb(asqrt[44] ), .dout(n9297));
  jand g09060(.dina(n9029), .dinb(n9297), .dout(n9298));
  jor  g09061(.dina(n9298), .dinb(n9218), .dout(n9299));
  jor  g09062(.dina(n9299), .dinb(asqrt[45] ), .dout(n9300));
  jnot g09063(.din(n9037), .dout(n9301));
  jand g09064(.dina(n9301), .dinb(n9300), .dout(n9302));
  jor  g09065(.dina(n9302), .dinb(n9217), .dout(n9303));
  jor  g09066(.dina(n9303), .dinb(asqrt[46] ), .dout(n9304));
  jand g09067(.dina(n9044), .dinb(n9304), .dout(n9305));
  jor  g09068(.dina(n9305), .dinb(n9216), .dout(n9306));
  jor  g09069(.dina(n9306), .dinb(asqrt[47] ), .dout(n9307));
  jnot g09070(.din(n9052), .dout(n9308));
  jand g09071(.dina(n9308), .dinb(n9307), .dout(n9309));
  jor  g09072(.dina(n9309), .dinb(n9215), .dout(n9310));
  jor  g09073(.dina(n9310), .dinb(asqrt[48] ), .dout(n9311));
  jand g09074(.dina(n9059), .dinb(n9311), .dout(n9312));
  jor  g09075(.dina(n9312), .dinb(n9214), .dout(n9313));
  jor  g09076(.dina(n9313), .dinb(asqrt[49] ), .dout(n9314));
  jnot g09077(.din(n9067), .dout(n9315));
  jand g09078(.dina(n9315), .dinb(n9314), .dout(n9316));
  jor  g09079(.dina(n9316), .dinb(n9213), .dout(n9317));
  jor  g09080(.dina(n9317), .dinb(asqrt[50] ), .dout(n9318));
  jand g09081(.dina(n9074), .dinb(n9318), .dout(n9319));
  jor  g09082(.dina(n9319), .dinb(n9212), .dout(n9320));
  jor  g09083(.dina(n9320), .dinb(asqrt[51] ), .dout(n9321));
  jand g09084(.dina(n9082), .dinb(n9321), .dout(n9322));
  jor  g09085(.dina(n9322), .dinb(n9211), .dout(n9323));
  jor  g09086(.dina(n9323), .dinb(asqrt[52] ), .dout(n9324));
  jand g09087(.dina(n9090), .dinb(n9324), .dout(n9325));
  jor  g09088(.dina(n9325), .dinb(n9210), .dout(n9326));
  jor  g09089(.dina(n9326), .dinb(asqrt[53] ), .dout(n9327));
  jnot g09090(.din(n9098), .dout(n9328));
  jand g09091(.dina(n9328), .dinb(n9327), .dout(n9329));
  jor  g09092(.dina(n9329), .dinb(n9209), .dout(n9330));
  jor  g09093(.dina(n9330), .dinb(asqrt[54] ), .dout(n9331));
  jnot g09094(.din(n9105), .dout(n9332));
  jand g09095(.dina(n9332), .dinb(n9331), .dout(n9333));
  jor  g09096(.dina(n9333), .dinb(n9208), .dout(n9334));
  jor  g09097(.dina(n9334), .dinb(asqrt[55] ), .dout(n9335));
  jnot g09098(.din(n9112), .dout(n9336));
  jand g09099(.dina(n9336), .dinb(n9335), .dout(n9337));
  jor  g09100(.dina(n9337), .dinb(n9207), .dout(n9338));
  jor  g09101(.dina(n9338), .dinb(asqrt[56] ), .dout(n9339));
  jand g09102(.dina(n9119), .dinb(n9339), .dout(n9340));
  jor  g09103(.dina(n9340), .dinb(n9206), .dout(n9341));
  jor  g09104(.dina(n9341), .dinb(asqrt[57] ), .dout(n9342));
  jnot g09105(.din(n9127), .dout(n9343));
  jand g09106(.dina(n9343), .dinb(n9342), .dout(n9344));
  jor  g09107(.dina(n9344), .dinb(n9205), .dout(n9345));
  jor  g09108(.dina(n9345), .dinb(asqrt[58] ), .dout(n9346));
  jand g09109(.dina(n9134), .dinb(n9346), .dout(n9347));
  jor  g09110(.dina(n9347), .dinb(n9204), .dout(n9348));
  jor  g09111(.dina(n9348), .dinb(asqrt[59] ), .dout(n9349));
  jnot g09112(.din(n9142), .dout(n9350));
  jand g09113(.dina(n9350), .dinb(n9349), .dout(n9351));
  jor  g09114(.dina(n9351), .dinb(n9203), .dout(n9352));
  jor  g09115(.dina(n9352), .dinb(asqrt[60] ), .dout(n9353));
  jand g09116(.dina(n9149), .dinb(n9353), .dout(n9354));
  jor  g09117(.dina(n9354), .dinb(n9202), .dout(n9355));
  jor  g09118(.dina(n9355), .dinb(asqrt[61] ), .dout(n9356));
  jand g09119(.dina(n9157), .dinb(n9356), .dout(n9357));
  jor  g09120(.dina(n9357), .dinb(n9201), .dout(n9358));
  jor  g09121(.dina(n9358), .dinb(asqrt[62] ), .dout(n9359));
  jand g09122(.dina(n9184), .dinb(n9359), .dout(n9360));
  jor  g09123(.dina(n9360), .dinb(n9200), .dout(n9361));
  jand g09124(.dina(n9361), .dinb(n8893), .dout(n9362));
  jnot g09125(.din(n9177), .dout(n9363));
  jand g09126(.dina(n9363), .dinb(n9362), .dout(n9364));
  jor  g09127(.dina(n9364), .dinb(asqrt[63] ), .dout(n9365));
  jnot g09128(.din(n9180), .dout(n9366));
  jand g09129(.dina(n9366), .dinb(n9365), .dout(n9367));
  jand g09130(.dina(n9367), .dinb(n9173), .dout(n9368));
  jand g09131(.dina(n9368), .dinb(n9199), .dout(n9369));
  jor  g09132(.dina(n9369), .dinb(n9198), .dout(n9370));
  jand g09133(.dina(n9370), .dinb(n9197), .dout(n9371));
  jand g09134(.dina(n9371), .dinb(n9195), .dout(n9372));
  jor  g09135(.dina(n9372), .dinb(n9194), .dout(n9373));
  jand g09136(.dina(n9373), .dinb(asqrt[28] ), .dout(n9374));
  jor  g09137(.dina(n9373), .dinb(asqrt[28] ), .dout(n9375));
  jand g09138(.dina(asqrt[26] ), .dinb(n8897), .dout(n9376));
  jand g09139(.dina(n9172), .dinb(n9199), .dout(n9377));
  jand g09140(.dina(n9377), .dinb(n9365), .dout(n9378));
  jand g09141(.dina(n9378), .dinb(asqrt[27] ), .dout(n9379));
  jor  g09142(.dina(n9379), .dinb(n9376), .dout(n9380));
  jxor g09143(.dina(n9380), .dinb(a[54] ), .dout(n9381));
  jnot g09144(.din(n9381), .dout(n9382));
  jand g09145(.dina(n9382), .dinb(n9375), .dout(n9383));
  jor  g09146(.dina(n9383), .dinb(n9374), .dout(n9384));
  jand g09147(.dina(n9384), .dinb(asqrt[29] ), .dout(n9385));
  jor  g09148(.dina(n9384), .dinb(asqrt[29] ), .dout(n9386));
  jxor g09149(.dina(n8901), .dinb(n8449), .dout(n9387));
  jand g09150(.dina(n9387), .dinb(asqrt[26] ), .dout(n9388));
  jxor g09151(.dina(n9388), .dinb(n9240), .dout(n9389));
  jand g09152(.dina(n9389), .dinb(n9386), .dout(n9390));
  jor  g09153(.dina(n9390), .dinb(n9385), .dout(n9391));
  jand g09154(.dina(n9391), .dinb(asqrt[30] ), .dout(n9392));
  jor  g09155(.dina(n9391), .dinb(asqrt[30] ), .dout(n9393));
  jxor g09156(.dina(n8909), .dinb(n8003), .dout(n9394));
  jand g09157(.dina(n9394), .dinb(asqrt[26] ), .dout(n9395));
  jxor g09158(.dina(n9395), .dinb(n8918), .dout(n9396));
  jnot g09159(.din(n9396), .dout(n9397));
  jand g09160(.dina(n9397), .dinb(n9393), .dout(n9398));
  jor  g09161(.dina(n9398), .dinb(n9392), .dout(n9399));
  jand g09162(.dina(n9399), .dinb(asqrt[31] ), .dout(n9400));
  jor  g09163(.dina(n9399), .dinb(asqrt[31] ), .dout(n9401));
  jxor g09164(.dina(n8920), .dinb(n7581), .dout(n9402));
  jand g09165(.dina(n9402), .dinb(asqrt[26] ), .dout(n9403));
  jxor g09166(.dina(n9403), .dinb(n8925), .dout(n9404));
  jand g09167(.dina(n9404), .dinb(n9401), .dout(n9405));
  jor  g09168(.dina(n9405), .dinb(n9400), .dout(n9406));
  jand g09169(.dina(n9406), .dinb(asqrt[32] ), .dout(n9407));
  jor  g09170(.dina(n9406), .dinb(asqrt[32] ), .dout(n9408));
  jxor g09171(.dina(n8928), .dinb(n7154), .dout(n9409));
  jand g09172(.dina(n9409), .dinb(asqrt[26] ), .dout(n9410));
  jxor g09173(.dina(n9410), .dinb(n8933), .dout(n9411));
  jnot g09174(.din(n9411), .dout(n9412));
  jand g09175(.dina(n9412), .dinb(n9408), .dout(n9413));
  jor  g09176(.dina(n9413), .dinb(n9407), .dout(n9414));
  jand g09177(.dina(n9414), .dinb(asqrt[33] ), .dout(n9415));
  jor  g09178(.dina(n9414), .dinb(asqrt[33] ), .dout(n9416));
  jxor g09179(.dina(n8935), .dinb(n6758), .dout(n9417));
  jand g09180(.dina(n9417), .dinb(asqrt[26] ), .dout(n9418));
  jxor g09181(.dina(n9418), .dinb(n8940), .dout(n9419));
  jnot g09182(.din(n9419), .dout(n9420));
  jand g09183(.dina(n9420), .dinb(n9416), .dout(n9421));
  jor  g09184(.dina(n9421), .dinb(n9415), .dout(n9422));
  jand g09185(.dina(n9422), .dinb(asqrt[34] ), .dout(n9423));
  jor  g09186(.dina(n9422), .dinb(asqrt[34] ), .dout(n9424));
  jxor g09187(.dina(n8942), .dinb(n6357), .dout(n9425));
  jand g09188(.dina(n9425), .dinb(asqrt[26] ), .dout(n9426));
  jxor g09189(.dina(n9426), .dinb(n8947), .dout(n9427));
  jnot g09190(.din(n9427), .dout(n9428));
  jand g09191(.dina(n9428), .dinb(n9424), .dout(n9429));
  jor  g09192(.dina(n9429), .dinb(n9423), .dout(n9430));
  jand g09193(.dina(n9430), .dinb(asqrt[35] ), .dout(n9431));
  jor  g09194(.dina(n9430), .dinb(asqrt[35] ), .dout(n9432));
  jxor g09195(.dina(n8949), .dinb(n5989), .dout(n9433));
  jand g09196(.dina(n9433), .dinb(asqrt[26] ), .dout(n9434));
  jxor g09197(.dina(n9434), .dinb(n8954), .dout(n9435));
  jnot g09198(.din(n9435), .dout(n9436));
  jand g09199(.dina(n9436), .dinb(n9432), .dout(n9437));
  jor  g09200(.dina(n9437), .dinb(n9431), .dout(n9438));
  jand g09201(.dina(n9438), .dinb(asqrt[36] ), .dout(n9439));
  jor  g09202(.dina(n9438), .dinb(asqrt[36] ), .dout(n9440));
  jxor g09203(.dina(n8956), .dinb(n5606), .dout(n9441));
  jand g09204(.dina(n9441), .dinb(asqrt[26] ), .dout(n9442));
  jxor g09205(.dina(n9442), .dinb(n8961), .dout(n9443));
  jnot g09206(.din(n9443), .dout(n9444));
  jand g09207(.dina(n9444), .dinb(n9440), .dout(n9445));
  jor  g09208(.dina(n9445), .dinb(n9439), .dout(n9446));
  jand g09209(.dina(n9446), .dinb(asqrt[37] ), .dout(n9447));
  jxor g09210(.dina(n8963), .dinb(n5259), .dout(n9448));
  jand g09211(.dina(n9448), .dinb(asqrt[26] ), .dout(n9449));
  jxor g09212(.dina(n9449), .dinb(n8967), .dout(n9450));
  jor  g09213(.dina(n9446), .dinb(asqrt[37] ), .dout(n9451));
  jand g09214(.dina(n9451), .dinb(n9450), .dout(n9452));
  jor  g09215(.dina(n9452), .dinb(n9447), .dout(n9453));
  jand g09216(.dina(n9453), .dinb(asqrt[38] ), .dout(n9454));
  jor  g09217(.dina(n9453), .dinb(asqrt[38] ), .dout(n9455));
  jxor g09218(.dina(n8971), .dinb(n4902), .dout(n9456));
  jand g09219(.dina(n9456), .dinb(asqrt[26] ), .dout(n9457));
  jxor g09220(.dina(n9457), .dinb(n8976), .dout(n9458));
  jnot g09221(.din(n9458), .dout(n9459));
  jand g09222(.dina(n9459), .dinb(n9455), .dout(n9460));
  jor  g09223(.dina(n9460), .dinb(n9454), .dout(n9461));
  jand g09224(.dina(n9461), .dinb(asqrt[39] ), .dout(n9462));
  jor  g09225(.dina(n9461), .dinb(asqrt[39] ), .dout(n9463));
  jxor g09226(.dina(n8978), .dinb(n4582), .dout(n9464));
  jand g09227(.dina(n9464), .dinb(asqrt[26] ), .dout(n9465));
  jxor g09228(.dina(n9465), .dinb(n8983), .dout(n9466));
  jand g09229(.dina(n9466), .dinb(n9463), .dout(n9467));
  jor  g09230(.dina(n9467), .dinb(n9462), .dout(n9468));
  jand g09231(.dina(n9468), .dinb(asqrt[40] ), .dout(n9469));
  jor  g09232(.dina(n9468), .dinb(asqrt[40] ), .dout(n9470));
  jxor g09233(.dina(n8986), .dinb(n4249), .dout(n9471));
  jand g09234(.dina(n9471), .dinb(asqrt[26] ), .dout(n9472));
  jxor g09235(.dina(n9472), .dinb(n8991), .dout(n9473));
  jnot g09236(.din(n9473), .dout(n9474));
  jand g09237(.dina(n9474), .dinb(n9470), .dout(n9475));
  jor  g09238(.dina(n9475), .dinb(n9469), .dout(n9476));
  jand g09239(.dina(n9476), .dinb(asqrt[41] ), .dout(n9477));
  jor  g09240(.dina(n9476), .dinb(asqrt[41] ), .dout(n9478));
  jxor g09241(.dina(n8993), .dinb(n3955), .dout(n9479));
  jand g09242(.dina(n9479), .dinb(asqrt[26] ), .dout(n9480));
  jxor g09243(.dina(n9480), .dinb(n8998), .dout(n9481));
  jand g09244(.dina(n9481), .dinb(n9478), .dout(n9482));
  jor  g09245(.dina(n9482), .dinb(n9477), .dout(n9483));
  jand g09246(.dina(n9483), .dinb(asqrt[42] ), .dout(n9484));
  jor  g09247(.dina(n9483), .dinb(asqrt[42] ), .dout(n9485));
  jxor g09248(.dina(n9001), .dinb(n3642), .dout(n9486));
  jand g09249(.dina(n9486), .dinb(asqrt[26] ), .dout(n9487));
  jxor g09250(.dina(n9487), .dinb(n9006), .dout(n9488));
  jand g09251(.dina(n9488), .dinb(n9485), .dout(n9489));
  jor  g09252(.dina(n9489), .dinb(n9484), .dout(n9490));
  jand g09253(.dina(n9490), .dinb(asqrt[43] ), .dout(n9491));
  jor  g09254(.dina(n9490), .dinb(asqrt[43] ), .dout(n9492));
  jxor g09255(.dina(n9009), .dinb(n3368), .dout(n9493));
  jand g09256(.dina(n9493), .dinb(asqrt[26] ), .dout(n9494));
  jxor g09257(.dina(n9494), .dinb(n9015), .dout(n9495));
  jnot g09258(.din(n9495), .dout(n9496));
  jand g09259(.dina(n9496), .dinb(n9492), .dout(n9497));
  jor  g09260(.dina(n9497), .dinb(n9491), .dout(n9498));
  jand g09261(.dina(n9498), .dinb(asqrt[44] ), .dout(n9499));
  jor  g09262(.dina(n9498), .dinb(asqrt[44] ), .dout(n9500));
  jxor g09263(.dina(n9017), .dinb(n3089), .dout(n9501));
  jand g09264(.dina(n9501), .dinb(asqrt[26] ), .dout(n9502));
  jxor g09265(.dina(n9502), .dinb(n9022), .dout(n9503));
  jnot g09266(.din(n9503), .dout(n9504));
  jand g09267(.dina(n9504), .dinb(n9500), .dout(n9505));
  jor  g09268(.dina(n9505), .dinb(n9499), .dout(n9506));
  jand g09269(.dina(n9506), .dinb(asqrt[45] ), .dout(n9507));
  jor  g09270(.dina(n9506), .dinb(asqrt[45] ), .dout(n9508));
  jxor g09271(.dina(n9024), .dinb(n2833), .dout(n9509));
  jand g09272(.dina(n9509), .dinb(asqrt[26] ), .dout(n9510));
  jxor g09273(.dina(n9510), .dinb(n9029), .dout(n9511));
  jand g09274(.dina(n9511), .dinb(n9508), .dout(n9512));
  jor  g09275(.dina(n9512), .dinb(n9507), .dout(n9513));
  jand g09276(.dina(n9513), .dinb(asqrt[46] ), .dout(n9514));
  jor  g09277(.dina(n9513), .dinb(asqrt[46] ), .dout(n9515));
  jxor g09278(.dina(n9032), .dinb(n2572), .dout(n9516));
  jand g09279(.dina(n9516), .dinb(asqrt[26] ), .dout(n9517));
  jxor g09280(.dina(n9517), .dinb(n9037), .dout(n9518));
  jnot g09281(.din(n9518), .dout(n9519));
  jand g09282(.dina(n9519), .dinb(n9515), .dout(n9520));
  jor  g09283(.dina(n9520), .dinb(n9514), .dout(n9521));
  jand g09284(.dina(n9521), .dinb(asqrt[47] ), .dout(n9522));
  jor  g09285(.dina(n9521), .dinb(asqrt[47] ), .dout(n9523));
  jxor g09286(.dina(n9039), .dinb(n2345), .dout(n9524));
  jand g09287(.dina(n9524), .dinb(asqrt[26] ), .dout(n9525));
  jxor g09288(.dina(n9525), .dinb(n9044), .dout(n9526));
  jand g09289(.dina(n9526), .dinb(n9523), .dout(n9527));
  jor  g09290(.dina(n9527), .dinb(n9522), .dout(n9528));
  jand g09291(.dina(n9528), .dinb(asqrt[48] ), .dout(n9529));
  jor  g09292(.dina(n9528), .dinb(asqrt[48] ), .dout(n9530));
  jxor g09293(.dina(n9047), .dinb(n2108), .dout(n9531));
  jand g09294(.dina(n9531), .dinb(asqrt[26] ), .dout(n9532));
  jxor g09295(.dina(n9532), .dinb(n9052), .dout(n9533));
  jnot g09296(.din(n9533), .dout(n9534));
  jand g09297(.dina(n9534), .dinb(n9530), .dout(n9535));
  jor  g09298(.dina(n9535), .dinb(n9529), .dout(n9536));
  jand g09299(.dina(n9536), .dinb(asqrt[49] ), .dout(n9537));
  jor  g09300(.dina(n9536), .dinb(asqrt[49] ), .dout(n9538));
  jxor g09301(.dina(n9054), .dinb(n1912), .dout(n9539));
  jand g09302(.dina(n9539), .dinb(asqrt[26] ), .dout(n9540));
  jxor g09303(.dina(n9540), .dinb(n9059), .dout(n9541));
  jand g09304(.dina(n9541), .dinb(n9538), .dout(n9542));
  jor  g09305(.dina(n9542), .dinb(n9537), .dout(n9543));
  jand g09306(.dina(n9543), .dinb(asqrt[50] ), .dout(n9544));
  jor  g09307(.dina(n9543), .dinb(asqrt[50] ), .dout(n9545));
  jxor g09308(.dina(n9062), .dinb(n1699), .dout(n9546));
  jand g09309(.dina(n9546), .dinb(asqrt[26] ), .dout(n9547));
  jxor g09310(.dina(n9547), .dinb(n9067), .dout(n9548));
  jnot g09311(.din(n9548), .dout(n9549));
  jand g09312(.dina(n9549), .dinb(n9545), .dout(n9550));
  jor  g09313(.dina(n9550), .dinb(n9544), .dout(n9551));
  jand g09314(.dina(n9551), .dinb(asqrt[51] ), .dout(n9552));
  jor  g09315(.dina(n9551), .dinb(asqrt[51] ), .dout(n9553));
  jxor g09316(.dina(n9069), .dinb(n1516), .dout(n9554));
  jand g09317(.dina(n9554), .dinb(asqrt[26] ), .dout(n9555));
  jxor g09318(.dina(n9555), .dinb(n9074), .dout(n9556));
  jand g09319(.dina(n9556), .dinb(n9553), .dout(n9557));
  jor  g09320(.dina(n9557), .dinb(n9552), .dout(n9558));
  jand g09321(.dina(n9558), .dinb(asqrt[52] ), .dout(n9559));
  jor  g09322(.dina(n9558), .dinb(asqrt[52] ), .dout(n9560));
  jxor g09323(.dina(n9077), .dinb(n1332), .dout(n9561));
  jand g09324(.dina(n9561), .dinb(asqrt[26] ), .dout(n9562));
  jxor g09325(.dina(n9562), .dinb(n9082), .dout(n9563));
  jand g09326(.dina(n9563), .dinb(n9560), .dout(n9564));
  jor  g09327(.dina(n9564), .dinb(n9559), .dout(n9565));
  jand g09328(.dina(n9565), .dinb(asqrt[53] ), .dout(n9566));
  jor  g09329(.dina(n9565), .dinb(asqrt[53] ), .dout(n9567));
  jxor g09330(.dina(n9085), .dinb(n1173), .dout(n9568));
  jand g09331(.dina(n9568), .dinb(asqrt[26] ), .dout(n9569));
  jxor g09332(.dina(n9569), .dinb(n9090), .dout(n9570));
  jand g09333(.dina(n9570), .dinb(n9567), .dout(n9571));
  jor  g09334(.dina(n9571), .dinb(n9566), .dout(n9572));
  jand g09335(.dina(n9572), .dinb(asqrt[54] ), .dout(n9573));
  jor  g09336(.dina(n9572), .dinb(asqrt[54] ), .dout(n9574));
  jxor g09337(.dina(n9093), .dinb(n1008), .dout(n9575));
  jand g09338(.dina(n9575), .dinb(asqrt[26] ), .dout(n9576));
  jxor g09339(.dina(n9576), .dinb(n9098), .dout(n9577));
  jnot g09340(.din(n9577), .dout(n9578));
  jand g09341(.dina(n9578), .dinb(n9574), .dout(n9579));
  jor  g09342(.dina(n9579), .dinb(n9573), .dout(n9580));
  jand g09343(.dina(n9580), .dinb(asqrt[55] ), .dout(n9581));
  jor  g09344(.dina(n9580), .dinb(asqrt[55] ), .dout(n9582));
  jxor g09345(.dina(n9100), .dinb(n884), .dout(n9583));
  jand g09346(.dina(n9583), .dinb(asqrt[26] ), .dout(n9584));
  jxor g09347(.dina(n9584), .dinb(n9105), .dout(n9585));
  jnot g09348(.din(n9585), .dout(n9586));
  jand g09349(.dina(n9586), .dinb(n9582), .dout(n9587));
  jor  g09350(.dina(n9587), .dinb(n9581), .dout(n9588));
  jand g09351(.dina(n9588), .dinb(asqrt[56] ), .dout(n9589));
  jor  g09352(.dina(n9588), .dinb(asqrt[56] ), .dout(n9590));
  jxor g09353(.dina(n9107), .dinb(n743), .dout(n9591));
  jand g09354(.dina(n9591), .dinb(asqrt[26] ), .dout(n9592));
  jxor g09355(.dina(n9592), .dinb(n9112), .dout(n9593));
  jnot g09356(.din(n9593), .dout(n9594));
  jand g09357(.dina(n9594), .dinb(n9590), .dout(n9595));
  jor  g09358(.dina(n9595), .dinb(n9589), .dout(n9596));
  jand g09359(.dina(n9596), .dinb(asqrt[57] ), .dout(n9597));
  jor  g09360(.dina(n9596), .dinb(asqrt[57] ), .dout(n9598));
  jxor g09361(.dina(n9114), .dinb(n635), .dout(n9599));
  jand g09362(.dina(n9599), .dinb(asqrt[26] ), .dout(n9600));
  jxor g09363(.dina(n9600), .dinb(n9119), .dout(n9601));
  jand g09364(.dina(n9601), .dinb(n9598), .dout(n9602));
  jor  g09365(.dina(n9602), .dinb(n9597), .dout(n9603));
  jand g09366(.dina(n9603), .dinb(asqrt[58] ), .dout(n9604));
  jor  g09367(.dina(n9603), .dinb(asqrt[58] ), .dout(n9605));
  jxor g09368(.dina(n9122), .dinb(n515), .dout(n9606));
  jand g09369(.dina(n9606), .dinb(asqrt[26] ), .dout(n9607));
  jxor g09370(.dina(n9607), .dinb(n9127), .dout(n9608));
  jnot g09371(.din(n9608), .dout(n9609));
  jand g09372(.dina(n9609), .dinb(n9605), .dout(n9610));
  jor  g09373(.dina(n9610), .dinb(n9604), .dout(n9611));
  jand g09374(.dina(n9611), .dinb(asqrt[59] ), .dout(n9612));
  jor  g09375(.dina(n9611), .dinb(asqrt[59] ), .dout(n9613));
  jxor g09376(.dina(n9129), .dinb(n443), .dout(n9614));
  jand g09377(.dina(n9614), .dinb(asqrt[26] ), .dout(n9615));
  jxor g09378(.dina(n9615), .dinb(n9135), .dout(n9616));
  jnot g09379(.din(n9616), .dout(n9617));
  jand g09380(.dina(n9617), .dinb(n9613), .dout(n9618));
  jor  g09381(.dina(n9618), .dinb(n9612), .dout(n9619));
  jand g09382(.dina(n9619), .dinb(asqrt[60] ), .dout(n9620));
  jor  g09383(.dina(n9619), .dinb(asqrt[60] ), .dout(n9621));
  jxor g09384(.dina(n9137), .dinb(n352), .dout(n9622));
  jand g09385(.dina(n9622), .dinb(asqrt[26] ), .dout(n9623));
  jxor g09386(.dina(n9623), .dinb(n9142), .dout(n9624));
  jnot g09387(.din(n9624), .dout(n9625));
  jand g09388(.dina(n9625), .dinb(n9621), .dout(n9626));
  jor  g09389(.dina(n9626), .dinb(n9620), .dout(n9627));
  jand g09390(.dina(n9627), .dinb(asqrt[61] ), .dout(n9628));
  jor  g09391(.dina(n9627), .dinb(asqrt[61] ), .dout(n9629));
  jxor g09392(.dina(n9144), .dinb(n294), .dout(n9630));
  jand g09393(.dina(n9630), .dinb(asqrt[26] ), .dout(n9631));
  jxor g09394(.dina(n9631), .dinb(n9149), .dout(n9632));
  jand g09395(.dina(n9632), .dinb(n9629), .dout(n9633));
  jor  g09396(.dina(n9633), .dinb(n9628), .dout(n9634));
  jand g09397(.dina(n9634), .dinb(asqrt[62] ), .dout(n9635));
  jor  g09398(.dina(n9634), .dinb(asqrt[62] ), .dout(n9636));
  jxor g09399(.dina(n9152), .dinb(n239), .dout(n9637));
  jand g09400(.dina(n9637), .dinb(asqrt[26] ), .dout(n9638));
  jxor g09401(.dina(n9638), .dinb(n9157), .dout(n9639));
  jand g09402(.dina(n9639), .dinb(n9636), .dout(n9640));
  jor  g09403(.dina(n9640), .dinb(n9635), .dout(n9641));
  jor  g09404(.dina(n9641), .dinb(n9187), .dout(n9642));
  jnot g09405(.din(n9642), .dout(n9643));
  jand g09406(.dina(n9368), .dinb(n9167), .dout(n9644));
  jnot g09407(.din(n9644), .dout(n9645));
  jxor g09408(.dina(n9167), .dinb(n8894), .dout(n9646));
  jand g09409(.dina(n9646), .dinb(asqrt[63] ), .dout(n9647));
  jand g09410(.dina(n9647), .dinb(n9645), .dout(n9648));
  jnot g09411(.din(n9187), .dout(n9649));
  jnot g09412(.din(n9635), .dout(n9650));
  jnot g09413(.din(n9628), .dout(n9651));
  jnot g09414(.din(n9620), .dout(n9652));
  jnot g09415(.din(n9612), .dout(n9653));
  jnot g09416(.din(n9604), .dout(n9654));
  jnot g09417(.din(n9597), .dout(n9655));
  jnot g09418(.din(n9589), .dout(n9656));
  jnot g09419(.din(n9581), .dout(n9657));
  jnot g09420(.din(n9573), .dout(n9658));
  jnot g09421(.din(n9566), .dout(n9659));
  jnot g09422(.din(n9559), .dout(n9660));
  jnot g09423(.din(n9552), .dout(n9661));
  jnot g09424(.din(n9544), .dout(n9662));
  jnot g09425(.din(n9537), .dout(n9663));
  jnot g09426(.din(n9529), .dout(n9664));
  jnot g09427(.din(n9522), .dout(n9665));
  jnot g09428(.din(n9514), .dout(n9666));
  jnot g09429(.din(n9507), .dout(n9667));
  jnot g09430(.din(n9499), .dout(n9668));
  jnot g09431(.din(n9491), .dout(n9669));
  jnot g09432(.din(n9484), .dout(n9670));
  jnot g09433(.din(n9477), .dout(n9671));
  jnot g09434(.din(n9469), .dout(n9672));
  jnot g09435(.din(n9462), .dout(n9673));
  jnot g09436(.din(n9454), .dout(n9674));
  jnot g09437(.din(n9447), .dout(n9675));
  jnot g09438(.din(n9450), .dout(n9676));
  jnot g09439(.din(n9439), .dout(n9677));
  jnot g09440(.din(n9431), .dout(n9678));
  jnot g09441(.din(n9423), .dout(n9679));
  jnot g09442(.din(n9415), .dout(n9680));
  jnot g09443(.din(n9407), .dout(n9681));
  jnot g09444(.din(n9400), .dout(n9682));
  jnot g09445(.din(n9392), .dout(n9683));
  jnot g09446(.din(n9385), .dout(n9684));
  jnot g09447(.din(n9374), .dout(n9685));
  jnot g09448(.din(n9194), .dout(n9686));
  jnot g09449(.din(n9191), .dout(n9687));
  jor  g09450(.dina(n9369), .dinb(n8895), .dout(n9688));
  jand g09451(.dina(n9688), .dinb(n9687), .dout(n9689));
  jand g09452(.dina(n9689), .dinb(n8890), .dout(n9690));
  jor  g09453(.dina(n9369), .dinb(a[52] ), .dout(n9691));
  jand g09454(.dina(n9691), .dinb(a[53] ), .dout(n9692));
  jor  g09455(.dina(n9376), .dinb(n9692), .dout(n9693));
  jor  g09456(.dina(n9693), .dinb(n9690), .dout(n9694));
  jand g09457(.dina(n9694), .dinb(n9686), .dout(n9695));
  jand g09458(.dina(n9695), .dinb(n8449), .dout(n9696));
  jor  g09459(.dina(n9381), .dinb(n9696), .dout(n9697));
  jand g09460(.dina(n9697), .dinb(n9685), .dout(n9698));
  jand g09461(.dina(n9698), .dinb(n8003), .dout(n9699));
  jnot g09462(.din(n9389), .dout(n9700));
  jor  g09463(.dina(n9700), .dinb(n9699), .dout(n9701));
  jand g09464(.dina(n9701), .dinb(n9684), .dout(n9702));
  jand g09465(.dina(n9702), .dinb(n7581), .dout(n9703));
  jor  g09466(.dina(n9396), .dinb(n9703), .dout(n9704));
  jand g09467(.dina(n9704), .dinb(n9683), .dout(n9705));
  jand g09468(.dina(n9705), .dinb(n7154), .dout(n9706));
  jnot g09469(.din(n9404), .dout(n9707));
  jor  g09470(.dina(n9707), .dinb(n9706), .dout(n9708));
  jand g09471(.dina(n9708), .dinb(n9682), .dout(n9709));
  jand g09472(.dina(n9709), .dinb(n6758), .dout(n9710));
  jor  g09473(.dina(n9411), .dinb(n9710), .dout(n9711));
  jand g09474(.dina(n9711), .dinb(n9681), .dout(n9712));
  jand g09475(.dina(n9712), .dinb(n6357), .dout(n9713));
  jor  g09476(.dina(n9419), .dinb(n9713), .dout(n9714));
  jand g09477(.dina(n9714), .dinb(n9680), .dout(n9715));
  jand g09478(.dina(n9715), .dinb(n5989), .dout(n9716));
  jor  g09479(.dina(n9427), .dinb(n9716), .dout(n9717));
  jand g09480(.dina(n9717), .dinb(n9679), .dout(n9718));
  jand g09481(.dina(n9718), .dinb(n5606), .dout(n9719));
  jor  g09482(.dina(n9435), .dinb(n9719), .dout(n9720));
  jand g09483(.dina(n9720), .dinb(n9678), .dout(n9721));
  jand g09484(.dina(n9721), .dinb(n5259), .dout(n9722));
  jor  g09485(.dina(n9443), .dinb(n9722), .dout(n9723));
  jand g09486(.dina(n9723), .dinb(n9677), .dout(n9724));
  jand g09487(.dina(n9724), .dinb(n4902), .dout(n9725));
  jor  g09488(.dina(n9725), .dinb(n9676), .dout(n9726));
  jand g09489(.dina(n9726), .dinb(n9675), .dout(n9727));
  jand g09490(.dina(n9727), .dinb(n4582), .dout(n9728));
  jor  g09491(.dina(n9458), .dinb(n9728), .dout(n9729));
  jand g09492(.dina(n9729), .dinb(n9674), .dout(n9730));
  jand g09493(.dina(n9730), .dinb(n4249), .dout(n9731));
  jnot g09494(.din(n9466), .dout(n9732));
  jor  g09495(.dina(n9732), .dinb(n9731), .dout(n9733));
  jand g09496(.dina(n9733), .dinb(n9673), .dout(n9734));
  jand g09497(.dina(n9734), .dinb(n3955), .dout(n9735));
  jor  g09498(.dina(n9473), .dinb(n9735), .dout(n9736));
  jand g09499(.dina(n9736), .dinb(n9672), .dout(n9737));
  jand g09500(.dina(n9737), .dinb(n3642), .dout(n9738));
  jnot g09501(.din(n9481), .dout(n9739));
  jor  g09502(.dina(n9739), .dinb(n9738), .dout(n9740));
  jand g09503(.dina(n9740), .dinb(n9671), .dout(n9741));
  jand g09504(.dina(n9741), .dinb(n3368), .dout(n9742));
  jnot g09505(.din(n9488), .dout(n9743));
  jor  g09506(.dina(n9743), .dinb(n9742), .dout(n9744));
  jand g09507(.dina(n9744), .dinb(n9670), .dout(n9745));
  jand g09508(.dina(n9745), .dinb(n3089), .dout(n9746));
  jor  g09509(.dina(n9495), .dinb(n9746), .dout(n9747));
  jand g09510(.dina(n9747), .dinb(n9669), .dout(n9748));
  jand g09511(.dina(n9748), .dinb(n2833), .dout(n9749));
  jor  g09512(.dina(n9503), .dinb(n9749), .dout(n9750));
  jand g09513(.dina(n9750), .dinb(n9668), .dout(n9751));
  jand g09514(.dina(n9751), .dinb(n2572), .dout(n9752));
  jnot g09515(.din(n9511), .dout(n9753));
  jor  g09516(.dina(n9753), .dinb(n9752), .dout(n9754));
  jand g09517(.dina(n9754), .dinb(n9667), .dout(n9755));
  jand g09518(.dina(n9755), .dinb(n2345), .dout(n9756));
  jor  g09519(.dina(n9518), .dinb(n9756), .dout(n9757));
  jand g09520(.dina(n9757), .dinb(n9666), .dout(n9758));
  jand g09521(.dina(n9758), .dinb(n2108), .dout(n9759));
  jnot g09522(.din(n9526), .dout(n9760));
  jor  g09523(.dina(n9760), .dinb(n9759), .dout(n9761));
  jand g09524(.dina(n9761), .dinb(n9665), .dout(n9762));
  jand g09525(.dina(n9762), .dinb(n1912), .dout(n9763));
  jor  g09526(.dina(n9533), .dinb(n9763), .dout(n9764));
  jand g09527(.dina(n9764), .dinb(n9664), .dout(n9765));
  jand g09528(.dina(n9765), .dinb(n1699), .dout(n9766));
  jnot g09529(.din(n9541), .dout(n9767));
  jor  g09530(.dina(n9767), .dinb(n9766), .dout(n9768));
  jand g09531(.dina(n9768), .dinb(n9663), .dout(n9769));
  jand g09532(.dina(n9769), .dinb(n1516), .dout(n9770));
  jor  g09533(.dina(n9548), .dinb(n9770), .dout(n9771));
  jand g09534(.dina(n9771), .dinb(n9662), .dout(n9772));
  jand g09535(.dina(n9772), .dinb(n1332), .dout(n9773));
  jnot g09536(.din(n9556), .dout(n9774));
  jor  g09537(.dina(n9774), .dinb(n9773), .dout(n9775));
  jand g09538(.dina(n9775), .dinb(n9661), .dout(n9776));
  jand g09539(.dina(n9776), .dinb(n1173), .dout(n9777));
  jnot g09540(.din(n9563), .dout(n9778));
  jor  g09541(.dina(n9778), .dinb(n9777), .dout(n9779));
  jand g09542(.dina(n9779), .dinb(n9660), .dout(n9780));
  jand g09543(.dina(n9780), .dinb(n1008), .dout(n9781));
  jnot g09544(.din(n9570), .dout(n9782));
  jor  g09545(.dina(n9782), .dinb(n9781), .dout(n9783));
  jand g09546(.dina(n9783), .dinb(n9659), .dout(n9784));
  jand g09547(.dina(n9784), .dinb(n884), .dout(n9785));
  jor  g09548(.dina(n9577), .dinb(n9785), .dout(n9786));
  jand g09549(.dina(n9786), .dinb(n9658), .dout(n9787));
  jand g09550(.dina(n9787), .dinb(n743), .dout(n9788));
  jor  g09551(.dina(n9585), .dinb(n9788), .dout(n9789));
  jand g09552(.dina(n9789), .dinb(n9657), .dout(n9790));
  jand g09553(.dina(n9790), .dinb(n635), .dout(n9791));
  jor  g09554(.dina(n9593), .dinb(n9791), .dout(n9792));
  jand g09555(.dina(n9792), .dinb(n9656), .dout(n9793));
  jand g09556(.dina(n9793), .dinb(n515), .dout(n9794));
  jnot g09557(.din(n9601), .dout(n9795));
  jor  g09558(.dina(n9795), .dinb(n9794), .dout(n9796));
  jand g09559(.dina(n9796), .dinb(n9655), .dout(n9797));
  jand g09560(.dina(n9797), .dinb(n443), .dout(n9798));
  jor  g09561(.dina(n9608), .dinb(n9798), .dout(n9799));
  jand g09562(.dina(n9799), .dinb(n9654), .dout(n9800));
  jand g09563(.dina(n9800), .dinb(n352), .dout(n9801));
  jor  g09564(.dina(n9616), .dinb(n9801), .dout(n9802));
  jand g09565(.dina(n9802), .dinb(n9653), .dout(n9803));
  jand g09566(.dina(n9803), .dinb(n294), .dout(n9804));
  jor  g09567(.dina(n9624), .dinb(n9804), .dout(n9805));
  jand g09568(.dina(n9805), .dinb(n9652), .dout(n9806));
  jand g09569(.dina(n9806), .dinb(n239), .dout(n9807));
  jnot g09570(.din(n9632), .dout(n9808));
  jor  g09571(.dina(n9808), .dinb(n9807), .dout(n9809));
  jand g09572(.dina(n9809), .dinb(n9651), .dout(n9810));
  jand g09573(.dina(n9810), .dinb(n221), .dout(n9811));
  jnot g09574(.din(n9639), .dout(n9812));
  jor  g09575(.dina(n9812), .dinb(n9811), .dout(n9813));
  jand g09576(.dina(n9813), .dinb(n9650), .dout(n9814));
  jor  g09577(.dina(n9814), .dinb(n9649), .dout(n9815));
  jor  g09578(.dina(n9646), .dinb(n9369), .dout(n9816));
  jnot g09579(.din(n9816), .dout(n9817));
  jor  g09580(.dina(n9817), .dinb(n9815), .dout(n9818));
  jand g09581(.dina(n9818), .dinb(n218), .dout(n9819));
  jand g09582(.dina(n9369), .dinb(n8894), .dout(n9820));
  jor  g09583(.dina(n9820), .dinb(n9819), .dout(n9821));
  jor  g09584(.dina(n9821), .dinb(n9648), .dout(n9822));
  jor  g09585(.dina(n9822), .dinb(n9643), .dout(asqrt[25] ));
  jand g09586(.dina(n9641), .dinb(n9187), .dout(n9824));
  jand g09587(.dina(n9822), .dinb(n9824), .dout(n9825));
  jnot g09588(.din(n9648), .dout(n9826));
  jand g09589(.dina(n9816), .dinb(n9824), .dout(n9827));
  jor  g09590(.dina(n9827), .dinb(asqrt[63] ), .dout(n9828));
  jnot g09591(.din(n9820), .dout(n9829));
  jand g09592(.dina(n9829), .dinb(n9828), .dout(n9830));
  jand g09593(.dina(n9830), .dinb(n9826), .dout(n9831));
  jand g09594(.dina(n9831), .dinb(n9642), .dout(n9832));
  jor  g09595(.dina(n9832), .dinb(n9188), .dout(n9833));
  jnot g09596(.din(a[48] ), .dout(n9834));
  jnot g09597(.din(a[49] ), .dout(n9835));
  jand g09598(.dina(n9835), .dinb(n9834), .dout(n9836));
  jand g09599(.dina(n9836), .dinb(n9188), .dout(n9837));
  jnot g09600(.din(n9837), .dout(n9838));
  jand g09601(.dina(n9838), .dinb(n9833), .dout(n9839));
  jor  g09602(.dina(n9839), .dinb(n9369), .dout(n9840));
  jand g09603(.dina(n9839), .dinb(n9369), .dout(n9841));
  jor  g09604(.dina(n9832), .dinb(a[50] ), .dout(n9842));
  jand g09605(.dina(n9842), .dinb(a[51] ), .dout(n9843));
  jand g09606(.dina(asqrt[25] ), .dinb(n9190), .dout(n9844));
  jor  g09607(.dina(n9844), .dinb(n9843), .dout(n9845));
  jor  g09608(.dina(n9845), .dinb(n9841), .dout(n9846));
  jand g09609(.dina(n9846), .dinb(n9840), .dout(n9847));
  jor  g09610(.dina(n9847), .dinb(n8890), .dout(n9848));
  jand g09611(.dina(n9847), .dinb(n8890), .dout(n9849));
  jnot g09612(.din(n9190), .dout(n9850));
  jor  g09613(.dina(n9832), .dinb(n9850), .dout(n9851));
  jor  g09614(.dina(n9647), .dinb(n9643), .dout(n9852));
  jor  g09615(.dina(n9852), .dinb(n9819), .dout(n9853));
  jor  g09616(.dina(n9853), .dinb(n9369), .dout(n9854));
  jand g09617(.dina(n9854), .dinb(n9851), .dout(n9855));
  jxor g09618(.dina(n9855), .dinb(n8895), .dout(n9856));
  jor  g09619(.dina(n9856), .dinb(n9849), .dout(n9857));
  jand g09620(.dina(n9857), .dinb(n9848), .dout(n9858));
  jor  g09621(.dina(n9858), .dinb(n8449), .dout(n9859));
  jand g09622(.dina(n9858), .dinb(n8449), .dout(n9860));
  jxor g09623(.dina(n9193), .dinb(n8890), .dout(n9861));
  jor  g09624(.dina(n9861), .dinb(n9832), .dout(n9862));
  jxor g09625(.dina(n9862), .dinb(n9693), .dout(n9863));
  jnot g09626(.din(n9863), .dout(n9864));
  jor  g09627(.dina(n9864), .dinb(n9860), .dout(n9865));
  jand g09628(.dina(n9865), .dinb(n9859), .dout(n9866));
  jor  g09629(.dina(n9866), .dinb(n8003), .dout(n9867));
  jand g09630(.dina(n9866), .dinb(n8003), .dout(n9868));
  jxor g09631(.dina(n9373), .dinb(n8449), .dout(n9869));
  jor  g09632(.dina(n9869), .dinb(n9832), .dout(n9870));
  jxor g09633(.dina(n9870), .dinb(n9382), .dout(n9871));
  jor  g09634(.dina(n9871), .dinb(n9868), .dout(n9872));
  jand g09635(.dina(n9872), .dinb(n9867), .dout(n9873));
  jor  g09636(.dina(n9873), .dinb(n7581), .dout(n9874));
  jand g09637(.dina(n9873), .dinb(n7581), .dout(n9875));
  jxor g09638(.dina(n9384), .dinb(n8003), .dout(n9876));
  jor  g09639(.dina(n9876), .dinb(n9832), .dout(n9877));
  jxor g09640(.dina(n9877), .dinb(n9389), .dout(n9878));
  jor  g09641(.dina(n9878), .dinb(n9875), .dout(n9879));
  jand g09642(.dina(n9879), .dinb(n9874), .dout(n9880));
  jor  g09643(.dina(n9880), .dinb(n7154), .dout(n9881));
  jand g09644(.dina(n9880), .dinb(n7154), .dout(n9882));
  jxor g09645(.dina(n9391), .dinb(n7581), .dout(n9883));
  jor  g09646(.dina(n9883), .dinb(n9832), .dout(n9884));
  jxor g09647(.dina(n9884), .dinb(n9397), .dout(n9885));
  jor  g09648(.dina(n9885), .dinb(n9882), .dout(n9886));
  jand g09649(.dina(n9886), .dinb(n9881), .dout(n9887));
  jor  g09650(.dina(n9887), .dinb(n6758), .dout(n9888));
  jand g09651(.dina(n9887), .dinb(n6758), .dout(n9889));
  jxor g09652(.dina(n9399), .dinb(n7154), .dout(n9890));
  jor  g09653(.dina(n9890), .dinb(n9832), .dout(n9891));
  jxor g09654(.dina(n9891), .dinb(n9707), .dout(n9892));
  jnot g09655(.din(n9892), .dout(n9893));
  jor  g09656(.dina(n9893), .dinb(n9889), .dout(n9894));
  jand g09657(.dina(n9894), .dinb(n9888), .dout(n9895));
  jor  g09658(.dina(n9895), .dinb(n6357), .dout(n9896));
  jand g09659(.dina(n9895), .dinb(n6357), .dout(n9897));
  jxor g09660(.dina(n9406), .dinb(n6758), .dout(n9898));
  jor  g09661(.dina(n9898), .dinb(n9832), .dout(n9899));
  jxor g09662(.dina(n9899), .dinb(n9412), .dout(n9900));
  jor  g09663(.dina(n9900), .dinb(n9897), .dout(n9901));
  jand g09664(.dina(n9901), .dinb(n9896), .dout(n9902));
  jor  g09665(.dina(n9902), .dinb(n5989), .dout(n9903));
  jand g09666(.dina(n9902), .dinb(n5989), .dout(n9904));
  jxor g09667(.dina(n9414), .dinb(n6357), .dout(n9905));
  jor  g09668(.dina(n9905), .dinb(n9832), .dout(n9906));
  jxor g09669(.dina(n9906), .dinb(n9420), .dout(n9907));
  jor  g09670(.dina(n9907), .dinb(n9904), .dout(n9908));
  jand g09671(.dina(n9908), .dinb(n9903), .dout(n9909));
  jor  g09672(.dina(n9909), .dinb(n5606), .dout(n9910));
  jand g09673(.dina(n9909), .dinb(n5606), .dout(n9911));
  jxor g09674(.dina(n9422), .dinb(n5989), .dout(n9912));
  jor  g09675(.dina(n9912), .dinb(n9832), .dout(n9913));
  jxor g09676(.dina(n9913), .dinb(n9428), .dout(n9914));
  jor  g09677(.dina(n9914), .dinb(n9911), .dout(n9915));
  jand g09678(.dina(n9915), .dinb(n9910), .dout(n9916));
  jor  g09679(.dina(n9916), .dinb(n5259), .dout(n9917));
  jand g09680(.dina(n9916), .dinb(n5259), .dout(n9918));
  jxor g09681(.dina(n9430), .dinb(n5606), .dout(n9919));
  jor  g09682(.dina(n9919), .dinb(n9832), .dout(n9920));
  jxor g09683(.dina(n9920), .dinb(n9436), .dout(n9921));
  jor  g09684(.dina(n9921), .dinb(n9918), .dout(n9922));
  jand g09685(.dina(n9922), .dinb(n9917), .dout(n9923));
  jor  g09686(.dina(n9923), .dinb(n4902), .dout(n9924));
  jand g09687(.dina(n9923), .dinb(n4902), .dout(n9925));
  jxor g09688(.dina(n9438), .dinb(n5259), .dout(n9926));
  jor  g09689(.dina(n9926), .dinb(n9832), .dout(n9927));
  jxor g09690(.dina(n9927), .dinb(n9444), .dout(n9928));
  jor  g09691(.dina(n9928), .dinb(n9925), .dout(n9929));
  jand g09692(.dina(n9929), .dinb(n9924), .dout(n9930));
  jor  g09693(.dina(n9930), .dinb(n4582), .dout(n9931));
  jxor g09694(.dina(n9446), .dinb(n4902), .dout(n9932));
  jor  g09695(.dina(n9932), .dinb(n9832), .dout(n9933));
  jxor g09696(.dina(n9933), .dinb(n9676), .dout(n9934));
  jnot g09697(.din(n9934), .dout(n9935));
  jand g09698(.dina(n9930), .dinb(n4582), .dout(n9936));
  jor  g09699(.dina(n9936), .dinb(n9935), .dout(n9937));
  jand g09700(.dina(n9937), .dinb(n9931), .dout(n9938));
  jor  g09701(.dina(n9938), .dinb(n4249), .dout(n9939));
  jand g09702(.dina(n9938), .dinb(n4249), .dout(n9940));
  jxor g09703(.dina(n9453), .dinb(n4582), .dout(n9941));
  jor  g09704(.dina(n9941), .dinb(n9832), .dout(n9942));
  jxor g09705(.dina(n9942), .dinb(n9459), .dout(n9943));
  jor  g09706(.dina(n9943), .dinb(n9940), .dout(n9944));
  jand g09707(.dina(n9944), .dinb(n9939), .dout(n9945));
  jor  g09708(.dina(n9945), .dinb(n3955), .dout(n9946));
  jand g09709(.dina(n9945), .dinb(n3955), .dout(n9947));
  jxor g09710(.dina(n9461), .dinb(n4249), .dout(n9948));
  jor  g09711(.dina(n9948), .dinb(n9832), .dout(n9949));
  jxor g09712(.dina(n9949), .dinb(n9732), .dout(n9950));
  jnot g09713(.din(n9950), .dout(n9951));
  jor  g09714(.dina(n9951), .dinb(n9947), .dout(n9952));
  jand g09715(.dina(n9952), .dinb(n9946), .dout(n9953));
  jor  g09716(.dina(n9953), .dinb(n3642), .dout(n9954));
  jand g09717(.dina(n9953), .dinb(n3642), .dout(n9955));
  jxor g09718(.dina(n9468), .dinb(n3955), .dout(n9956));
  jor  g09719(.dina(n9956), .dinb(n9832), .dout(n9957));
  jxor g09720(.dina(n9957), .dinb(n9474), .dout(n9958));
  jor  g09721(.dina(n9958), .dinb(n9955), .dout(n9959));
  jand g09722(.dina(n9959), .dinb(n9954), .dout(n9960));
  jor  g09723(.dina(n9960), .dinb(n3368), .dout(n9961));
  jand g09724(.dina(n9960), .dinb(n3368), .dout(n9962));
  jxor g09725(.dina(n9476), .dinb(n3642), .dout(n9963));
  jor  g09726(.dina(n9963), .dinb(n9832), .dout(n9964));
  jxor g09727(.dina(n9964), .dinb(n9739), .dout(n9965));
  jnot g09728(.din(n9965), .dout(n9966));
  jor  g09729(.dina(n9966), .dinb(n9962), .dout(n9967));
  jand g09730(.dina(n9967), .dinb(n9961), .dout(n9968));
  jor  g09731(.dina(n9968), .dinb(n3089), .dout(n9969));
  jand g09732(.dina(n9968), .dinb(n3089), .dout(n9970));
  jxor g09733(.dina(n9483), .dinb(n3368), .dout(n9971));
  jor  g09734(.dina(n9971), .dinb(n9832), .dout(n9972));
  jxor g09735(.dina(n9972), .dinb(n9488), .dout(n9973));
  jor  g09736(.dina(n9973), .dinb(n9970), .dout(n9974));
  jand g09737(.dina(n9974), .dinb(n9969), .dout(n9975));
  jor  g09738(.dina(n9975), .dinb(n2833), .dout(n9976));
  jand g09739(.dina(n9975), .dinb(n2833), .dout(n9977));
  jxor g09740(.dina(n9490), .dinb(n3089), .dout(n9978));
  jor  g09741(.dina(n9978), .dinb(n9832), .dout(n9979));
  jxor g09742(.dina(n9979), .dinb(n9496), .dout(n9980));
  jor  g09743(.dina(n9980), .dinb(n9977), .dout(n9981));
  jand g09744(.dina(n9981), .dinb(n9976), .dout(n9982));
  jor  g09745(.dina(n9982), .dinb(n2572), .dout(n9983));
  jand g09746(.dina(n9982), .dinb(n2572), .dout(n9984));
  jxor g09747(.dina(n9498), .dinb(n2833), .dout(n9985));
  jor  g09748(.dina(n9985), .dinb(n9832), .dout(n9986));
  jxor g09749(.dina(n9986), .dinb(n9504), .dout(n9987));
  jor  g09750(.dina(n9987), .dinb(n9984), .dout(n9988));
  jand g09751(.dina(n9988), .dinb(n9983), .dout(n9989));
  jor  g09752(.dina(n9989), .dinb(n2345), .dout(n9990));
  jand g09753(.dina(n9989), .dinb(n2345), .dout(n9991));
  jxor g09754(.dina(n9506), .dinb(n2572), .dout(n9992));
  jor  g09755(.dina(n9992), .dinb(n9832), .dout(n9993));
  jxor g09756(.dina(n9993), .dinb(n9753), .dout(n9994));
  jnot g09757(.din(n9994), .dout(n9995));
  jor  g09758(.dina(n9995), .dinb(n9991), .dout(n9996));
  jand g09759(.dina(n9996), .dinb(n9990), .dout(n9997));
  jor  g09760(.dina(n9997), .dinb(n2108), .dout(n9998));
  jand g09761(.dina(n9997), .dinb(n2108), .dout(n9999));
  jxor g09762(.dina(n9513), .dinb(n2345), .dout(n10000));
  jor  g09763(.dina(n10000), .dinb(n9832), .dout(n10001));
  jxor g09764(.dina(n10001), .dinb(n9519), .dout(n10002));
  jor  g09765(.dina(n10002), .dinb(n9999), .dout(n10003));
  jand g09766(.dina(n10003), .dinb(n9998), .dout(n10004));
  jor  g09767(.dina(n10004), .dinb(n1912), .dout(n10005));
  jand g09768(.dina(n10004), .dinb(n1912), .dout(n10006));
  jxor g09769(.dina(n9521), .dinb(n2108), .dout(n10007));
  jor  g09770(.dina(n10007), .dinb(n9832), .dout(n10008));
  jxor g09771(.dina(n10008), .dinb(n9760), .dout(n10009));
  jnot g09772(.din(n10009), .dout(n10010));
  jor  g09773(.dina(n10010), .dinb(n10006), .dout(n10011));
  jand g09774(.dina(n10011), .dinb(n10005), .dout(n10012));
  jor  g09775(.dina(n10012), .dinb(n1699), .dout(n10013));
  jand g09776(.dina(n10012), .dinb(n1699), .dout(n10014));
  jxor g09777(.dina(n9528), .dinb(n1912), .dout(n10015));
  jor  g09778(.dina(n10015), .dinb(n9832), .dout(n10016));
  jxor g09779(.dina(n10016), .dinb(n9534), .dout(n10017));
  jor  g09780(.dina(n10017), .dinb(n10014), .dout(n10018));
  jand g09781(.dina(n10018), .dinb(n10013), .dout(n10019));
  jor  g09782(.dina(n10019), .dinb(n1516), .dout(n10020));
  jand g09783(.dina(n10019), .dinb(n1516), .dout(n10021));
  jxor g09784(.dina(n9536), .dinb(n1699), .dout(n10022));
  jor  g09785(.dina(n10022), .dinb(n9832), .dout(n10023));
  jxor g09786(.dina(n10023), .dinb(n9767), .dout(n10024));
  jnot g09787(.din(n10024), .dout(n10025));
  jor  g09788(.dina(n10025), .dinb(n10021), .dout(n10026));
  jand g09789(.dina(n10026), .dinb(n10020), .dout(n10027));
  jor  g09790(.dina(n10027), .dinb(n1332), .dout(n10028));
  jand g09791(.dina(n10027), .dinb(n1332), .dout(n10029));
  jxor g09792(.dina(n9543), .dinb(n1516), .dout(n10030));
  jor  g09793(.dina(n10030), .dinb(n9832), .dout(n10031));
  jxor g09794(.dina(n10031), .dinb(n9549), .dout(n10032));
  jor  g09795(.dina(n10032), .dinb(n10029), .dout(n10033));
  jand g09796(.dina(n10033), .dinb(n10028), .dout(n10034));
  jor  g09797(.dina(n10034), .dinb(n1173), .dout(n10035));
  jand g09798(.dina(n10034), .dinb(n1173), .dout(n10036));
  jxor g09799(.dina(n9551), .dinb(n1332), .dout(n10037));
  jor  g09800(.dina(n10037), .dinb(n9832), .dout(n10038));
  jxor g09801(.dina(n10038), .dinb(n9774), .dout(n10039));
  jnot g09802(.din(n10039), .dout(n10040));
  jor  g09803(.dina(n10040), .dinb(n10036), .dout(n10041));
  jand g09804(.dina(n10041), .dinb(n10035), .dout(n10042));
  jor  g09805(.dina(n10042), .dinb(n1008), .dout(n10043));
  jand g09806(.dina(n10042), .dinb(n1008), .dout(n10044));
  jxor g09807(.dina(n9558), .dinb(n1173), .dout(n10045));
  jor  g09808(.dina(n10045), .dinb(n9832), .dout(n10046));
  jxor g09809(.dina(n10046), .dinb(n9778), .dout(n10047));
  jnot g09810(.din(n10047), .dout(n10048));
  jor  g09811(.dina(n10048), .dinb(n10044), .dout(n10049));
  jand g09812(.dina(n10049), .dinb(n10043), .dout(n10050));
  jor  g09813(.dina(n10050), .dinb(n884), .dout(n10051));
  jand g09814(.dina(n10050), .dinb(n884), .dout(n10052));
  jxor g09815(.dina(n9565), .dinb(n1008), .dout(n10053));
  jor  g09816(.dina(n10053), .dinb(n9832), .dout(n10054));
  jxor g09817(.dina(n10054), .dinb(n9782), .dout(n10055));
  jnot g09818(.din(n10055), .dout(n10056));
  jor  g09819(.dina(n10056), .dinb(n10052), .dout(n10057));
  jand g09820(.dina(n10057), .dinb(n10051), .dout(n10058));
  jor  g09821(.dina(n10058), .dinb(n743), .dout(n10059));
  jand g09822(.dina(n10058), .dinb(n743), .dout(n10060));
  jxor g09823(.dina(n9572), .dinb(n884), .dout(n10061));
  jor  g09824(.dina(n10061), .dinb(n9832), .dout(n10062));
  jxor g09825(.dina(n10062), .dinb(n9578), .dout(n10063));
  jor  g09826(.dina(n10063), .dinb(n10060), .dout(n10064));
  jand g09827(.dina(n10064), .dinb(n10059), .dout(n10065));
  jor  g09828(.dina(n10065), .dinb(n635), .dout(n10066));
  jand g09829(.dina(n10065), .dinb(n635), .dout(n10067));
  jxor g09830(.dina(n9580), .dinb(n743), .dout(n10068));
  jor  g09831(.dina(n10068), .dinb(n9832), .dout(n10069));
  jxor g09832(.dina(n10069), .dinb(n9586), .dout(n10070));
  jor  g09833(.dina(n10070), .dinb(n10067), .dout(n10071));
  jand g09834(.dina(n10071), .dinb(n10066), .dout(n10072));
  jor  g09835(.dina(n10072), .dinb(n515), .dout(n10073));
  jand g09836(.dina(n10072), .dinb(n515), .dout(n10074));
  jxor g09837(.dina(n9588), .dinb(n635), .dout(n10075));
  jor  g09838(.dina(n10075), .dinb(n9832), .dout(n10076));
  jxor g09839(.dina(n10076), .dinb(n9594), .dout(n10077));
  jor  g09840(.dina(n10077), .dinb(n10074), .dout(n10078));
  jand g09841(.dina(n10078), .dinb(n10073), .dout(n10079));
  jor  g09842(.dina(n10079), .dinb(n443), .dout(n10080));
  jand g09843(.dina(n10079), .dinb(n443), .dout(n10081));
  jxor g09844(.dina(n9596), .dinb(n515), .dout(n10082));
  jor  g09845(.dina(n10082), .dinb(n9832), .dout(n10083));
  jxor g09846(.dina(n10083), .dinb(n9795), .dout(n10084));
  jnot g09847(.din(n10084), .dout(n10085));
  jor  g09848(.dina(n10085), .dinb(n10081), .dout(n10086));
  jand g09849(.dina(n10086), .dinb(n10080), .dout(n10087));
  jor  g09850(.dina(n10087), .dinb(n352), .dout(n10088));
  jand g09851(.dina(n10087), .dinb(n352), .dout(n10089));
  jxor g09852(.dina(n9603), .dinb(n443), .dout(n10090));
  jor  g09853(.dina(n10090), .dinb(n9832), .dout(n10091));
  jxor g09854(.dina(n10091), .dinb(n9609), .dout(n10092));
  jor  g09855(.dina(n10092), .dinb(n10089), .dout(n10093));
  jand g09856(.dina(n10093), .dinb(n10088), .dout(n10094));
  jor  g09857(.dina(n10094), .dinb(n294), .dout(n10095));
  jand g09858(.dina(n10094), .dinb(n294), .dout(n10096));
  jxor g09859(.dina(n9611), .dinb(n352), .dout(n10097));
  jor  g09860(.dina(n10097), .dinb(n9832), .dout(n10098));
  jxor g09861(.dina(n10098), .dinb(n9617), .dout(n10099));
  jor  g09862(.dina(n10099), .dinb(n10096), .dout(n10100));
  jand g09863(.dina(n10100), .dinb(n10095), .dout(n10101));
  jor  g09864(.dina(n10101), .dinb(n239), .dout(n10102));
  jand g09865(.dina(n10101), .dinb(n239), .dout(n10103));
  jxor g09866(.dina(n9619), .dinb(n294), .dout(n10104));
  jor  g09867(.dina(n10104), .dinb(n9832), .dout(n10105));
  jxor g09868(.dina(n10105), .dinb(n9625), .dout(n10106));
  jor  g09869(.dina(n10106), .dinb(n10103), .dout(n10107));
  jand g09870(.dina(n10107), .dinb(n10102), .dout(n10108));
  jor  g09871(.dina(n10108), .dinb(n221), .dout(n10109));
  jand g09872(.dina(n10108), .dinb(n221), .dout(n10110));
  jxor g09873(.dina(n9627), .dinb(n239), .dout(n10111));
  jor  g09874(.dina(n10111), .dinb(n9832), .dout(n10112));
  jxor g09875(.dina(n10112), .dinb(n9808), .dout(n10113));
  jnot g09876(.din(n10113), .dout(n10114));
  jor  g09877(.dina(n10114), .dinb(n10110), .dout(n10115));
  jand g09878(.dina(n10115), .dinb(n10109), .dout(n10116));
  jxor g09879(.dina(n9634), .dinb(n221), .dout(n10117));
  jor  g09880(.dina(n10117), .dinb(n9832), .dout(n10118));
  jxor g09881(.dina(n10118), .dinb(n9639), .dout(n10119));
  jor  g09882(.dina(n10119), .dinb(n10116), .dout(n10120));
  jor  g09883(.dina(n10120), .dinb(n9643), .dout(n10121));
  jor  g09884(.dina(n10121), .dinb(n9825), .dout(n10122));
  jand g09885(.dina(n10122), .dinb(n218), .dout(n10123));
  jand g09886(.dina(n9832), .dinb(n9649), .dout(n10124));
  jand g09887(.dina(n10119), .dinb(n10116), .dout(n10125));
  jor  g09888(.dina(n10125), .dinb(n10124), .dout(n10126));
  jand g09889(.dina(n9831), .dinb(n9814), .dout(n10127));
  jnot g09890(.din(n10127), .dout(n10128));
  jand g09891(.dina(n9815), .dinb(asqrt[63] ), .dout(n10129));
  jand g09892(.dina(n10129), .dinb(n9642), .dout(n10130));
  jand g09893(.dina(n10130), .dinb(n10128), .dout(n10131));
  jor  g09894(.dina(n10131), .dinb(n10126), .dout(n10132));
  jor  g09895(.dina(n10132), .dinb(n10123), .dout(asqrt[24] ));
  jnot g09896(.din(a[46] ), .dout(n10134));
  jnot g09897(.din(a[47] ), .dout(n10135));
  jand g09898(.dina(n10135), .dinb(n10134), .dout(n10136));
  jand g09899(.dina(n10136), .dinb(n9834), .dout(n10137));
  jand g09900(.dina(asqrt[24] ), .dinb(a[48] ), .dout(n10138));
  jor  g09901(.dina(n10138), .dinb(n10137), .dout(n10139));
  jand g09902(.dina(n10139), .dinb(asqrt[25] ), .dout(n10140));
  jor  g09903(.dina(n10139), .dinb(asqrt[25] ), .dout(n10141));
  jand g09904(.dina(asqrt[24] ), .dinb(n9834), .dout(n10142));
  jor  g09905(.dina(n10142), .dinb(n9835), .dout(n10143));
  jnot g09906(.din(n9836), .dout(n10144));
  jnot g09907(.din(n9825), .dout(n10145));
  jnot g09908(.din(n10109), .dout(n10146));
  jnot g09909(.din(n10102), .dout(n10147));
  jnot g09910(.din(n10095), .dout(n10148));
  jnot g09911(.din(n10088), .dout(n10149));
  jnot g09912(.din(n10080), .dout(n10150));
  jnot g09913(.din(n10073), .dout(n10151));
  jnot g09914(.din(n10066), .dout(n10152));
  jnot g09915(.din(n10059), .dout(n10153));
  jnot g09916(.din(n10051), .dout(n10154));
  jnot g09917(.din(n10043), .dout(n10155));
  jnot g09918(.din(n10035), .dout(n10156));
  jnot g09919(.din(n10028), .dout(n10157));
  jnot g09920(.din(n10020), .dout(n10158));
  jnot g09921(.din(n10013), .dout(n10159));
  jnot g09922(.din(n10005), .dout(n10160));
  jnot g09923(.din(n9998), .dout(n10161));
  jnot g09924(.din(n9990), .dout(n10162));
  jnot g09925(.din(n9983), .dout(n10163));
  jnot g09926(.din(n9976), .dout(n10164));
  jnot g09927(.din(n9969), .dout(n10165));
  jnot g09928(.din(n9961), .dout(n10166));
  jnot g09929(.din(n9954), .dout(n10167));
  jnot g09930(.din(n9946), .dout(n10168));
  jnot g09931(.din(n9939), .dout(n10169));
  jnot g09932(.din(n9931), .dout(n10170));
  jnot g09933(.din(n9924), .dout(n10171));
  jnot g09934(.din(n9917), .dout(n10172));
  jnot g09935(.din(n9910), .dout(n10173));
  jnot g09936(.din(n9903), .dout(n10174));
  jnot g09937(.din(n9896), .dout(n10175));
  jnot g09938(.din(n9888), .dout(n10176));
  jnot g09939(.din(n9881), .dout(n10177));
  jnot g09940(.din(n9874), .dout(n10178));
  jnot g09941(.din(n9867), .dout(n10179));
  jnot g09942(.din(n9859), .dout(n10180));
  jnot g09943(.din(n9848), .dout(n10181));
  jnot g09944(.din(n9840), .dout(n10182));
  jand g09945(.dina(asqrt[25] ), .dinb(a[50] ), .dout(n10183));
  jor  g09946(.dina(n9837), .dinb(n10183), .dout(n10184));
  jor  g09947(.dina(n10184), .dinb(asqrt[26] ), .dout(n10185));
  jand g09948(.dina(asqrt[25] ), .dinb(n9188), .dout(n10186));
  jor  g09949(.dina(n10186), .dinb(n9189), .dout(n10187));
  jand g09950(.dina(n9851), .dinb(n10187), .dout(n10188));
  jand g09951(.dina(n10188), .dinb(n10185), .dout(n10189));
  jor  g09952(.dina(n10189), .dinb(n10182), .dout(n10190));
  jor  g09953(.dina(n10190), .dinb(asqrt[27] ), .dout(n10191));
  jnot g09954(.din(n9856), .dout(n10192));
  jand g09955(.dina(n10192), .dinb(n10191), .dout(n10193));
  jor  g09956(.dina(n10193), .dinb(n10181), .dout(n10194));
  jor  g09957(.dina(n10194), .dinb(asqrt[28] ), .dout(n10195));
  jand g09958(.dina(n9863), .dinb(n10195), .dout(n10196));
  jor  g09959(.dina(n10196), .dinb(n10180), .dout(n10197));
  jor  g09960(.dina(n10197), .dinb(asqrt[29] ), .dout(n10198));
  jnot g09961(.din(n9871), .dout(n10199));
  jand g09962(.dina(n10199), .dinb(n10198), .dout(n10200));
  jor  g09963(.dina(n10200), .dinb(n10179), .dout(n10201));
  jor  g09964(.dina(n10201), .dinb(asqrt[30] ), .dout(n10202));
  jnot g09965(.din(n9878), .dout(n10203));
  jand g09966(.dina(n10203), .dinb(n10202), .dout(n10204));
  jor  g09967(.dina(n10204), .dinb(n10178), .dout(n10205));
  jor  g09968(.dina(n10205), .dinb(asqrt[31] ), .dout(n10206));
  jnot g09969(.din(n9885), .dout(n10207));
  jand g09970(.dina(n10207), .dinb(n10206), .dout(n10208));
  jor  g09971(.dina(n10208), .dinb(n10177), .dout(n10209));
  jor  g09972(.dina(n10209), .dinb(asqrt[32] ), .dout(n10210));
  jand g09973(.dina(n9892), .dinb(n10210), .dout(n10211));
  jor  g09974(.dina(n10211), .dinb(n10176), .dout(n10212));
  jor  g09975(.dina(n10212), .dinb(asqrt[33] ), .dout(n10213));
  jnot g09976(.din(n9900), .dout(n10214));
  jand g09977(.dina(n10214), .dinb(n10213), .dout(n10215));
  jor  g09978(.dina(n10215), .dinb(n10175), .dout(n10216));
  jor  g09979(.dina(n10216), .dinb(asqrt[34] ), .dout(n10217));
  jnot g09980(.din(n9907), .dout(n10218));
  jand g09981(.dina(n10218), .dinb(n10217), .dout(n10219));
  jor  g09982(.dina(n10219), .dinb(n10174), .dout(n10220));
  jor  g09983(.dina(n10220), .dinb(asqrt[35] ), .dout(n10221));
  jnot g09984(.din(n9914), .dout(n10222));
  jand g09985(.dina(n10222), .dinb(n10221), .dout(n10223));
  jor  g09986(.dina(n10223), .dinb(n10173), .dout(n10224));
  jor  g09987(.dina(n10224), .dinb(asqrt[36] ), .dout(n10225));
  jnot g09988(.din(n9921), .dout(n10226));
  jand g09989(.dina(n10226), .dinb(n10225), .dout(n10227));
  jor  g09990(.dina(n10227), .dinb(n10172), .dout(n10228));
  jor  g09991(.dina(n10228), .dinb(asqrt[37] ), .dout(n10229));
  jnot g09992(.din(n9928), .dout(n10230));
  jand g09993(.dina(n10230), .dinb(n10229), .dout(n10231));
  jor  g09994(.dina(n10231), .dinb(n10171), .dout(n10232));
  jor  g09995(.dina(n10232), .dinb(asqrt[38] ), .dout(n10233));
  jand g09996(.dina(n10233), .dinb(n9934), .dout(n10234));
  jor  g09997(.dina(n10234), .dinb(n10170), .dout(n10235));
  jor  g09998(.dina(n10235), .dinb(asqrt[39] ), .dout(n10236));
  jnot g09999(.din(n9943), .dout(n10237));
  jand g10000(.dina(n10237), .dinb(n10236), .dout(n10238));
  jor  g10001(.dina(n10238), .dinb(n10169), .dout(n10239));
  jor  g10002(.dina(n10239), .dinb(asqrt[40] ), .dout(n10240));
  jand g10003(.dina(n9950), .dinb(n10240), .dout(n10241));
  jor  g10004(.dina(n10241), .dinb(n10168), .dout(n10242));
  jor  g10005(.dina(n10242), .dinb(asqrt[41] ), .dout(n10243));
  jnot g10006(.din(n9958), .dout(n10244));
  jand g10007(.dina(n10244), .dinb(n10243), .dout(n10245));
  jor  g10008(.dina(n10245), .dinb(n10167), .dout(n10246));
  jor  g10009(.dina(n10246), .dinb(asqrt[42] ), .dout(n10247));
  jand g10010(.dina(n9965), .dinb(n10247), .dout(n10248));
  jor  g10011(.dina(n10248), .dinb(n10166), .dout(n10249));
  jor  g10012(.dina(n10249), .dinb(asqrt[43] ), .dout(n10250));
  jnot g10013(.din(n9973), .dout(n10251));
  jand g10014(.dina(n10251), .dinb(n10250), .dout(n10252));
  jor  g10015(.dina(n10252), .dinb(n10165), .dout(n10253));
  jor  g10016(.dina(n10253), .dinb(asqrt[44] ), .dout(n10254));
  jnot g10017(.din(n9980), .dout(n10255));
  jand g10018(.dina(n10255), .dinb(n10254), .dout(n10256));
  jor  g10019(.dina(n10256), .dinb(n10164), .dout(n10257));
  jor  g10020(.dina(n10257), .dinb(asqrt[45] ), .dout(n10258));
  jnot g10021(.din(n9987), .dout(n10259));
  jand g10022(.dina(n10259), .dinb(n10258), .dout(n10260));
  jor  g10023(.dina(n10260), .dinb(n10163), .dout(n10261));
  jor  g10024(.dina(n10261), .dinb(asqrt[46] ), .dout(n10262));
  jand g10025(.dina(n9994), .dinb(n10262), .dout(n10263));
  jor  g10026(.dina(n10263), .dinb(n10162), .dout(n10264));
  jor  g10027(.dina(n10264), .dinb(asqrt[47] ), .dout(n10265));
  jnot g10028(.din(n10002), .dout(n10266));
  jand g10029(.dina(n10266), .dinb(n10265), .dout(n10267));
  jor  g10030(.dina(n10267), .dinb(n10161), .dout(n10268));
  jor  g10031(.dina(n10268), .dinb(asqrt[48] ), .dout(n10269));
  jand g10032(.dina(n10009), .dinb(n10269), .dout(n10270));
  jor  g10033(.dina(n10270), .dinb(n10160), .dout(n10271));
  jor  g10034(.dina(n10271), .dinb(asqrt[49] ), .dout(n10272));
  jnot g10035(.din(n10017), .dout(n10273));
  jand g10036(.dina(n10273), .dinb(n10272), .dout(n10274));
  jor  g10037(.dina(n10274), .dinb(n10159), .dout(n10275));
  jor  g10038(.dina(n10275), .dinb(asqrt[50] ), .dout(n10276));
  jand g10039(.dina(n10024), .dinb(n10276), .dout(n10277));
  jor  g10040(.dina(n10277), .dinb(n10158), .dout(n10278));
  jor  g10041(.dina(n10278), .dinb(asqrt[51] ), .dout(n10279));
  jnot g10042(.din(n10032), .dout(n10280));
  jand g10043(.dina(n10280), .dinb(n10279), .dout(n10281));
  jor  g10044(.dina(n10281), .dinb(n10157), .dout(n10282));
  jor  g10045(.dina(n10282), .dinb(asqrt[52] ), .dout(n10283));
  jand g10046(.dina(n10039), .dinb(n10283), .dout(n10284));
  jor  g10047(.dina(n10284), .dinb(n10156), .dout(n10285));
  jor  g10048(.dina(n10285), .dinb(asqrt[53] ), .dout(n10286));
  jand g10049(.dina(n10047), .dinb(n10286), .dout(n10287));
  jor  g10050(.dina(n10287), .dinb(n10155), .dout(n10288));
  jor  g10051(.dina(n10288), .dinb(asqrt[54] ), .dout(n10289));
  jand g10052(.dina(n10055), .dinb(n10289), .dout(n10290));
  jor  g10053(.dina(n10290), .dinb(n10154), .dout(n10291));
  jor  g10054(.dina(n10291), .dinb(asqrt[55] ), .dout(n10292));
  jnot g10055(.din(n10063), .dout(n10293));
  jand g10056(.dina(n10293), .dinb(n10292), .dout(n10294));
  jor  g10057(.dina(n10294), .dinb(n10153), .dout(n10295));
  jor  g10058(.dina(n10295), .dinb(asqrt[56] ), .dout(n10296));
  jnot g10059(.din(n10070), .dout(n10297));
  jand g10060(.dina(n10297), .dinb(n10296), .dout(n10298));
  jor  g10061(.dina(n10298), .dinb(n10152), .dout(n10299));
  jor  g10062(.dina(n10299), .dinb(asqrt[57] ), .dout(n10300));
  jnot g10063(.din(n10077), .dout(n10301));
  jand g10064(.dina(n10301), .dinb(n10300), .dout(n10302));
  jor  g10065(.dina(n10302), .dinb(n10151), .dout(n10303));
  jor  g10066(.dina(n10303), .dinb(asqrt[58] ), .dout(n10304));
  jand g10067(.dina(n10084), .dinb(n10304), .dout(n10305));
  jor  g10068(.dina(n10305), .dinb(n10150), .dout(n10306));
  jor  g10069(.dina(n10306), .dinb(asqrt[59] ), .dout(n10307));
  jnot g10070(.din(n10092), .dout(n10308));
  jand g10071(.dina(n10308), .dinb(n10307), .dout(n10309));
  jor  g10072(.dina(n10309), .dinb(n10149), .dout(n10310));
  jor  g10073(.dina(n10310), .dinb(asqrt[60] ), .dout(n10311));
  jnot g10074(.din(n10099), .dout(n10312));
  jand g10075(.dina(n10312), .dinb(n10311), .dout(n10313));
  jor  g10076(.dina(n10313), .dinb(n10148), .dout(n10314));
  jor  g10077(.dina(n10314), .dinb(asqrt[61] ), .dout(n10315));
  jnot g10078(.din(n10106), .dout(n10316));
  jand g10079(.dina(n10316), .dinb(n10315), .dout(n10317));
  jor  g10080(.dina(n10317), .dinb(n10147), .dout(n10318));
  jor  g10081(.dina(n10318), .dinb(asqrt[62] ), .dout(n10319));
  jand g10082(.dina(n10113), .dinb(n10319), .dout(n10320));
  jor  g10083(.dina(n10320), .dinb(n10146), .dout(n10321));
  jnot g10084(.din(n10119), .dout(n10322));
  jand g10085(.dina(n10322), .dinb(n10321), .dout(n10323));
  jand g10086(.dina(n10323), .dinb(n9642), .dout(n10324));
  jand g10087(.dina(n10324), .dinb(n10145), .dout(n10325));
  jor  g10088(.dina(n10325), .dinb(asqrt[63] ), .dout(n10326));
  jnot g10089(.din(n10132), .dout(n10327));
  jand g10090(.dina(n10327), .dinb(n10326), .dout(n10328));
  jor  g10091(.dina(n10328), .dinb(n10144), .dout(n10329));
  jand g10092(.dina(n10329), .dinb(n10143), .dout(n10330));
  jand g10093(.dina(n10330), .dinb(n10141), .dout(n10331));
  jor  g10094(.dina(n10331), .dinb(n10140), .dout(n10332));
  jand g10095(.dina(n10332), .dinb(asqrt[26] ), .dout(n10333));
  jor  g10096(.dina(n10332), .dinb(asqrt[26] ), .dout(n10334));
  jor  g10097(.dina(n10130), .dinb(n10125), .dout(n10335));
  jor  g10098(.dina(n10335), .dinb(n10123), .dout(n10336));
  jor  g10099(.dina(n10336), .dinb(n9832), .dout(n10337));
  jand g10100(.dina(n10337), .dinb(n10329), .dout(n10338));
  jxor g10101(.dina(n10338), .dinb(n9188), .dout(n10339));
  jnot g10102(.din(n10339), .dout(n10340));
  jand g10103(.dina(n10340), .dinb(n10334), .dout(n10341));
  jor  g10104(.dina(n10341), .dinb(n10333), .dout(n10342));
  jand g10105(.dina(n10342), .dinb(asqrt[27] ), .dout(n10343));
  jor  g10106(.dina(n10342), .dinb(asqrt[27] ), .dout(n10344));
  jxor g10107(.dina(n9839), .dinb(n9369), .dout(n10345));
  jand g10108(.dina(n10345), .dinb(asqrt[24] ), .dout(n10346));
  jxor g10109(.dina(n10346), .dinb(n10188), .dout(n10347));
  jand g10110(.dina(n10347), .dinb(n10344), .dout(n10348));
  jor  g10111(.dina(n10348), .dinb(n10343), .dout(n10349));
  jand g10112(.dina(n10349), .dinb(asqrt[28] ), .dout(n10350));
  jor  g10113(.dina(n10349), .dinb(asqrt[28] ), .dout(n10351));
  jxor g10114(.dina(n9847), .dinb(n8890), .dout(n10352));
  jand g10115(.dina(n10352), .dinb(asqrt[24] ), .dout(n10353));
  jxor g10116(.dina(n10353), .dinb(n9856), .dout(n10354));
  jnot g10117(.din(n10354), .dout(n10355));
  jand g10118(.dina(n10355), .dinb(n10351), .dout(n10356));
  jor  g10119(.dina(n10356), .dinb(n10350), .dout(n10357));
  jand g10120(.dina(n10357), .dinb(asqrt[29] ), .dout(n10358));
  jor  g10121(.dina(n10357), .dinb(asqrt[29] ), .dout(n10359));
  jxor g10122(.dina(n9858), .dinb(n8449), .dout(n10360));
  jand g10123(.dina(n10360), .dinb(asqrt[24] ), .dout(n10361));
  jxor g10124(.dina(n10361), .dinb(n9863), .dout(n10362));
  jand g10125(.dina(n10362), .dinb(n10359), .dout(n10363));
  jor  g10126(.dina(n10363), .dinb(n10358), .dout(n10364));
  jand g10127(.dina(n10364), .dinb(asqrt[30] ), .dout(n10365));
  jor  g10128(.dina(n10364), .dinb(asqrt[30] ), .dout(n10366));
  jxor g10129(.dina(n9866), .dinb(n8003), .dout(n10367));
  jand g10130(.dina(n10367), .dinb(asqrt[24] ), .dout(n10368));
  jxor g10131(.dina(n10368), .dinb(n9871), .dout(n10369));
  jnot g10132(.din(n10369), .dout(n10370));
  jand g10133(.dina(n10370), .dinb(n10366), .dout(n10371));
  jor  g10134(.dina(n10371), .dinb(n10365), .dout(n10372));
  jand g10135(.dina(n10372), .dinb(asqrt[31] ), .dout(n10373));
  jor  g10136(.dina(n10372), .dinb(asqrt[31] ), .dout(n10374));
  jxor g10137(.dina(n9873), .dinb(n7581), .dout(n10375));
  jand g10138(.dina(n10375), .dinb(asqrt[24] ), .dout(n10376));
  jxor g10139(.dina(n10376), .dinb(n9878), .dout(n10377));
  jnot g10140(.din(n10377), .dout(n10378));
  jand g10141(.dina(n10378), .dinb(n10374), .dout(n10379));
  jor  g10142(.dina(n10379), .dinb(n10373), .dout(n10380));
  jand g10143(.dina(n10380), .dinb(asqrt[32] ), .dout(n10381));
  jor  g10144(.dina(n10380), .dinb(asqrt[32] ), .dout(n10382));
  jxor g10145(.dina(n9880), .dinb(n7154), .dout(n10383));
  jand g10146(.dina(n10383), .dinb(asqrt[24] ), .dout(n10384));
  jxor g10147(.dina(n10384), .dinb(n9885), .dout(n10385));
  jnot g10148(.din(n10385), .dout(n10386));
  jand g10149(.dina(n10386), .dinb(n10382), .dout(n10387));
  jor  g10150(.dina(n10387), .dinb(n10381), .dout(n10388));
  jand g10151(.dina(n10388), .dinb(asqrt[33] ), .dout(n10389));
  jor  g10152(.dina(n10388), .dinb(asqrt[33] ), .dout(n10390));
  jxor g10153(.dina(n9887), .dinb(n6758), .dout(n10391));
  jand g10154(.dina(n10391), .dinb(asqrt[24] ), .dout(n10392));
  jxor g10155(.dina(n10392), .dinb(n9892), .dout(n10393));
  jand g10156(.dina(n10393), .dinb(n10390), .dout(n10394));
  jor  g10157(.dina(n10394), .dinb(n10389), .dout(n10395));
  jand g10158(.dina(n10395), .dinb(asqrt[34] ), .dout(n10396));
  jor  g10159(.dina(n10395), .dinb(asqrt[34] ), .dout(n10397));
  jxor g10160(.dina(n9895), .dinb(n6357), .dout(n10398));
  jand g10161(.dina(n10398), .dinb(asqrt[24] ), .dout(n10399));
  jxor g10162(.dina(n10399), .dinb(n9900), .dout(n10400));
  jnot g10163(.din(n10400), .dout(n10401));
  jand g10164(.dina(n10401), .dinb(n10397), .dout(n10402));
  jor  g10165(.dina(n10402), .dinb(n10396), .dout(n10403));
  jand g10166(.dina(n10403), .dinb(asqrt[35] ), .dout(n10404));
  jor  g10167(.dina(n10403), .dinb(asqrt[35] ), .dout(n10405));
  jxor g10168(.dina(n9902), .dinb(n5989), .dout(n10406));
  jand g10169(.dina(n10406), .dinb(asqrt[24] ), .dout(n10407));
  jxor g10170(.dina(n10407), .dinb(n9907), .dout(n10408));
  jnot g10171(.din(n10408), .dout(n10409));
  jand g10172(.dina(n10409), .dinb(n10405), .dout(n10410));
  jor  g10173(.dina(n10410), .dinb(n10404), .dout(n10411));
  jand g10174(.dina(n10411), .dinb(asqrt[36] ), .dout(n10412));
  jor  g10175(.dina(n10411), .dinb(asqrt[36] ), .dout(n10413));
  jxor g10176(.dina(n9909), .dinb(n5606), .dout(n10414));
  jand g10177(.dina(n10414), .dinb(asqrt[24] ), .dout(n10415));
  jxor g10178(.dina(n10415), .dinb(n9914), .dout(n10416));
  jnot g10179(.din(n10416), .dout(n10417));
  jand g10180(.dina(n10417), .dinb(n10413), .dout(n10418));
  jor  g10181(.dina(n10418), .dinb(n10412), .dout(n10419));
  jand g10182(.dina(n10419), .dinb(asqrt[37] ), .dout(n10420));
  jor  g10183(.dina(n10419), .dinb(asqrt[37] ), .dout(n10421));
  jxor g10184(.dina(n9916), .dinb(n5259), .dout(n10422));
  jand g10185(.dina(n10422), .dinb(asqrt[24] ), .dout(n10423));
  jxor g10186(.dina(n10423), .dinb(n9921), .dout(n10424));
  jnot g10187(.din(n10424), .dout(n10425));
  jand g10188(.dina(n10425), .dinb(n10421), .dout(n10426));
  jor  g10189(.dina(n10426), .dinb(n10420), .dout(n10427));
  jand g10190(.dina(n10427), .dinb(asqrt[38] ), .dout(n10428));
  jor  g10191(.dina(n10427), .dinb(asqrt[38] ), .dout(n10429));
  jxor g10192(.dina(n9923), .dinb(n4902), .dout(n10430));
  jand g10193(.dina(n10430), .dinb(asqrt[24] ), .dout(n10431));
  jxor g10194(.dina(n10431), .dinb(n9928), .dout(n10432));
  jnot g10195(.din(n10432), .dout(n10433));
  jand g10196(.dina(n10433), .dinb(n10429), .dout(n10434));
  jor  g10197(.dina(n10434), .dinb(n10428), .dout(n10435));
  jand g10198(.dina(n10435), .dinb(asqrt[39] ), .dout(n10436));
  jxor g10199(.dina(n9930), .dinb(n4582), .dout(n10437));
  jand g10200(.dina(n10437), .dinb(asqrt[24] ), .dout(n10438));
  jxor g10201(.dina(n10438), .dinb(n9934), .dout(n10439));
  jor  g10202(.dina(n10435), .dinb(asqrt[39] ), .dout(n10440));
  jand g10203(.dina(n10440), .dinb(n10439), .dout(n10441));
  jor  g10204(.dina(n10441), .dinb(n10436), .dout(n10442));
  jand g10205(.dina(n10442), .dinb(asqrt[40] ), .dout(n10443));
  jor  g10206(.dina(n10442), .dinb(asqrt[40] ), .dout(n10444));
  jxor g10207(.dina(n9938), .dinb(n4249), .dout(n10445));
  jand g10208(.dina(n10445), .dinb(asqrt[24] ), .dout(n10446));
  jxor g10209(.dina(n10446), .dinb(n9943), .dout(n10447));
  jnot g10210(.din(n10447), .dout(n10448));
  jand g10211(.dina(n10448), .dinb(n10444), .dout(n10449));
  jor  g10212(.dina(n10449), .dinb(n10443), .dout(n10450));
  jand g10213(.dina(n10450), .dinb(asqrt[41] ), .dout(n10451));
  jor  g10214(.dina(n10450), .dinb(asqrt[41] ), .dout(n10452));
  jxor g10215(.dina(n9945), .dinb(n3955), .dout(n10453));
  jand g10216(.dina(n10453), .dinb(asqrt[24] ), .dout(n10454));
  jxor g10217(.dina(n10454), .dinb(n9950), .dout(n10455));
  jand g10218(.dina(n10455), .dinb(n10452), .dout(n10456));
  jor  g10219(.dina(n10456), .dinb(n10451), .dout(n10457));
  jand g10220(.dina(n10457), .dinb(asqrt[42] ), .dout(n10458));
  jor  g10221(.dina(n10457), .dinb(asqrt[42] ), .dout(n10459));
  jxor g10222(.dina(n9953), .dinb(n3642), .dout(n10460));
  jand g10223(.dina(n10460), .dinb(asqrt[24] ), .dout(n10461));
  jxor g10224(.dina(n10461), .dinb(n9958), .dout(n10462));
  jnot g10225(.din(n10462), .dout(n10463));
  jand g10226(.dina(n10463), .dinb(n10459), .dout(n10464));
  jor  g10227(.dina(n10464), .dinb(n10458), .dout(n10465));
  jand g10228(.dina(n10465), .dinb(asqrt[43] ), .dout(n10466));
  jor  g10229(.dina(n10465), .dinb(asqrt[43] ), .dout(n10467));
  jxor g10230(.dina(n9960), .dinb(n3368), .dout(n10468));
  jand g10231(.dina(n10468), .dinb(asqrt[24] ), .dout(n10469));
  jxor g10232(.dina(n10469), .dinb(n9965), .dout(n10470));
  jand g10233(.dina(n10470), .dinb(n10467), .dout(n10471));
  jor  g10234(.dina(n10471), .dinb(n10466), .dout(n10472));
  jand g10235(.dina(n10472), .dinb(asqrt[44] ), .dout(n10473));
  jor  g10236(.dina(n10472), .dinb(asqrt[44] ), .dout(n10474));
  jxor g10237(.dina(n9968), .dinb(n3089), .dout(n10475));
  jand g10238(.dina(n10475), .dinb(asqrt[24] ), .dout(n10476));
  jxor g10239(.dina(n10476), .dinb(n9973), .dout(n10477));
  jnot g10240(.din(n10477), .dout(n10478));
  jand g10241(.dina(n10478), .dinb(n10474), .dout(n10479));
  jor  g10242(.dina(n10479), .dinb(n10473), .dout(n10480));
  jand g10243(.dina(n10480), .dinb(asqrt[45] ), .dout(n10481));
  jor  g10244(.dina(n10480), .dinb(asqrt[45] ), .dout(n10482));
  jxor g10245(.dina(n9975), .dinb(n2833), .dout(n10483));
  jand g10246(.dina(n10483), .dinb(asqrt[24] ), .dout(n10484));
  jxor g10247(.dina(n10484), .dinb(n9980), .dout(n10485));
  jnot g10248(.din(n10485), .dout(n10486));
  jand g10249(.dina(n10486), .dinb(n10482), .dout(n10487));
  jor  g10250(.dina(n10487), .dinb(n10481), .dout(n10488));
  jand g10251(.dina(n10488), .dinb(asqrt[46] ), .dout(n10489));
  jor  g10252(.dina(n10488), .dinb(asqrt[46] ), .dout(n10490));
  jxor g10253(.dina(n9982), .dinb(n2572), .dout(n10491));
  jand g10254(.dina(n10491), .dinb(asqrt[24] ), .dout(n10492));
  jxor g10255(.dina(n10492), .dinb(n9987), .dout(n10493));
  jnot g10256(.din(n10493), .dout(n10494));
  jand g10257(.dina(n10494), .dinb(n10490), .dout(n10495));
  jor  g10258(.dina(n10495), .dinb(n10489), .dout(n10496));
  jand g10259(.dina(n10496), .dinb(asqrt[47] ), .dout(n10497));
  jor  g10260(.dina(n10496), .dinb(asqrt[47] ), .dout(n10498));
  jxor g10261(.dina(n9989), .dinb(n2345), .dout(n10499));
  jand g10262(.dina(n10499), .dinb(asqrt[24] ), .dout(n10500));
  jxor g10263(.dina(n10500), .dinb(n9994), .dout(n10501));
  jand g10264(.dina(n10501), .dinb(n10498), .dout(n10502));
  jor  g10265(.dina(n10502), .dinb(n10497), .dout(n10503));
  jand g10266(.dina(n10503), .dinb(asqrt[48] ), .dout(n10504));
  jor  g10267(.dina(n10503), .dinb(asqrt[48] ), .dout(n10505));
  jxor g10268(.dina(n9997), .dinb(n2108), .dout(n10506));
  jand g10269(.dina(n10506), .dinb(asqrt[24] ), .dout(n10507));
  jxor g10270(.dina(n10507), .dinb(n10002), .dout(n10508));
  jnot g10271(.din(n10508), .dout(n10509));
  jand g10272(.dina(n10509), .dinb(n10505), .dout(n10510));
  jor  g10273(.dina(n10510), .dinb(n10504), .dout(n10511));
  jand g10274(.dina(n10511), .dinb(asqrt[49] ), .dout(n10512));
  jor  g10275(.dina(n10511), .dinb(asqrt[49] ), .dout(n10513));
  jxor g10276(.dina(n10004), .dinb(n1912), .dout(n10514));
  jand g10277(.dina(n10514), .dinb(asqrt[24] ), .dout(n10515));
  jxor g10278(.dina(n10515), .dinb(n10009), .dout(n10516));
  jand g10279(.dina(n10516), .dinb(n10513), .dout(n10517));
  jor  g10280(.dina(n10517), .dinb(n10512), .dout(n10518));
  jand g10281(.dina(n10518), .dinb(asqrt[50] ), .dout(n10519));
  jor  g10282(.dina(n10518), .dinb(asqrt[50] ), .dout(n10520));
  jxor g10283(.dina(n10012), .dinb(n1699), .dout(n10521));
  jand g10284(.dina(n10521), .dinb(asqrt[24] ), .dout(n10522));
  jxor g10285(.dina(n10522), .dinb(n10017), .dout(n10523));
  jnot g10286(.din(n10523), .dout(n10524));
  jand g10287(.dina(n10524), .dinb(n10520), .dout(n10525));
  jor  g10288(.dina(n10525), .dinb(n10519), .dout(n10526));
  jand g10289(.dina(n10526), .dinb(asqrt[51] ), .dout(n10527));
  jor  g10290(.dina(n10526), .dinb(asqrt[51] ), .dout(n10528));
  jxor g10291(.dina(n10019), .dinb(n1516), .dout(n10529));
  jand g10292(.dina(n10529), .dinb(asqrt[24] ), .dout(n10530));
  jxor g10293(.dina(n10530), .dinb(n10024), .dout(n10531));
  jand g10294(.dina(n10531), .dinb(n10528), .dout(n10532));
  jor  g10295(.dina(n10532), .dinb(n10527), .dout(n10533));
  jand g10296(.dina(n10533), .dinb(asqrt[52] ), .dout(n10534));
  jor  g10297(.dina(n10533), .dinb(asqrt[52] ), .dout(n10535));
  jxor g10298(.dina(n10027), .dinb(n1332), .dout(n10536));
  jand g10299(.dina(n10536), .dinb(asqrt[24] ), .dout(n10537));
  jxor g10300(.dina(n10537), .dinb(n10032), .dout(n10538));
  jnot g10301(.din(n10538), .dout(n10539));
  jand g10302(.dina(n10539), .dinb(n10535), .dout(n10540));
  jor  g10303(.dina(n10540), .dinb(n10534), .dout(n10541));
  jand g10304(.dina(n10541), .dinb(asqrt[53] ), .dout(n10542));
  jor  g10305(.dina(n10541), .dinb(asqrt[53] ), .dout(n10543));
  jxor g10306(.dina(n10034), .dinb(n1173), .dout(n10544));
  jand g10307(.dina(n10544), .dinb(asqrt[24] ), .dout(n10545));
  jxor g10308(.dina(n10545), .dinb(n10039), .dout(n10546));
  jand g10309(.dina(n10546), .dinb(n10543), .dout(n10547));
  jor  g10310(.dina(n10547), .dinb(n10542), .dout(n10548));
  jand g10311(.dina(n10548), .dinb(asqrt[54] ), .dout(n10549));
  jor  g10312(.dina(n10548), .dinb(asqrt[54] ), .dout(n10550));
  jxor g10313(.dina(n10042), .dinb(n1008), .dout(n10551));
  jand g10314(.dina(n10551), .dinb(asqrt[24] ), .dout(n10552));
  jxor g10315(.dina(n10552), .dinb(n10047), .dout(n10553));
  jand g10316(.dina(n10553), .dinb(n10550), .dout(n10554));
  jor  g10317(.dina(n10554), .dinb(n10549), .dout(n10555));
  jand g10318(.dina(n10555), .dinb(asqrt[55] ), .dout(n10556));
  jor  g10319(.dina(n10555), .dinb(asqrt[55] ), .dout(n10557));
  jxor g10320(.dina(n10050), .dinb(n884), .dout(n10558));
  jand g10321(.dina(n10558), .dinb(asqrt[24] ), .dout(n10559));
  jxor g10322(.dina(n10559), .dinb(n10055), .dout(n10560));
  jand g10323(.dina(n10560), .dinb(n10557), .dout(n10561));
  jor  g10324(.dina(n10561), .dinb(n10556), .dout(n10562));
  jand g10325(.dina(n10562), .dinb(asqrt[56] ), .dout(n10563));
  jor  g10326(.dina(n10562), .dinb(asqrt[56] ), .dout(n10564));
  jxor g10327(.dina(n10058), .dinb(n743), .dout(n10565));
  jand g10328(.dina(n10565), .dinb(asqrt[24] ), .dout(n10566));
  jxor g10329(.dina(n10566), .dinb(n10063), .dout(n10567));
  jnot g10330(.din(n10567), .dout(n10568));
  jand g10331(.dina(n10568), .dinb(n10564), .dout(n10569));
  jor  g10332(.dina(n10569), .dinb(n10563), .dout(n10570));
  jand g10333(.dina(n10570), .dinb(asqrt[57] ), .dout(n10571));
  jor  g10334(.dina(n10570), .dinb(asqrt[57] ), .dout(n10572));
  jxor g10335(.dina(n10065), .dinb(n635), .dout(n10573));
  jand g10336(.dina(n10573), .dinb(asqrt[24] ), .dout(n10574));
  jxor g10337(.dina(n10574), .dinb(n10070), .dout(n10575));
  jnot g10338(.din(n10575), .dout(n10576));
  jand g10339(.dina(n10576), .dinb(n10572), .dout(n10577));
  jor  g10340(.dina(n10577), .dinb(n10571), .dout(n10578));
  jand g10341(.dina(n10578), .dinb(asqrt[58] ), .dout(n10579));
  jor  g10342(.dina(n10578), .dinb(asqrt[58] ), .dout(n10580));
  jxor g10343(.dina(n10072), .dinb(n515), .dout(n10581));
  jand g10344(.dina(n10581), .dinb(asqrt[24] ), .dout(n10582));
  jxor g10345(.dina(n10582), .dinb(n10077), .dout(n10583));
  jnot g10346(.din(n10583), .dout(n10584));
  jand g10347(.dina(n10584), .dinb(n10580), .dout(n10585));
  jor  g10348(.dina(n10585), .dinb(n10579), .dout(n10586));
  jand g10349(.dina(n10586), .dinb(asqrt[59] ), .dout(n10587));
  jor  g10350(.dina(n10586), .dinb(asqrt[59] ), .dout(n10588));
  jxor g10351(.dina(n10079), .dinb(n443), .dout(n10589));
  jand g10352(.dina(n10589), .dinb(asqrt[24] ), .dout(n10590));
  jxor g10353(.dina(n10590), .dinb(n10084), .dout(n10591));
  jand g10354(.dina(n10591), .dinb(n10588), .dout(n10592));
  jor  g10355(.dina(n10592), .dinb(n10587), .dout(n10593));
  jand g10356(.dina(n10593), .dinb(asqrt[60] ), .dout(n10594));
  jor  g10357(.dina(n10593), .dinb(asqrt[60] ), .dout(n10595));
  jxor g10358(.dina(n10087), .dinb(n352), .dout(n10596));
  jand g10359(.dina(n10596), .dinb(asqrt[24] ), .dout(n10597));
  jxor g10360(.dina(n10597), .dinb(n10092), .dout(n10598));
  jnot g10361(.din(n10598), .dout(n10599));
  jand g10362(.dina(n10599), .dinb(n10595), .dout(n10600));
  jor  g10363(.dina(n10600), .dinb(n10594), .dout(n10601));
  jand g10364(.dina(n10601), .dinb(asqrt[61] ), .dout(n10602));
  jor  g10365(.dina(n10601), .dinb(asqrt[61] ), .dout(n10603));
  jxor g10366(.dina(n10094), .dinb(n294), .dout(n10604));
  jand g10367(.dina(n10604), .dinb(asqrt[24] ), .dout(n10605));
  jxor g10368(.dina(n10605), .dinb(n10099), .dout(n10606));
  jnot g10369(.din(n10606), .dout(n10607));
  jand g10370(.dina(n10607), .dinb(n10603), .dout(n10608));
  jor  g10371(.dina(n10608), .dinb(n10602), .dout(n10609));
  jand g10372(.dina(n10609), .dinb(asqrt[62] ), .dout(n10610));
  jnot g10373(.din(n10610), .dout(n10611));
  jnot g10374(.din(n10602), .dout(n10612));
  jnot g10375(.din(n10594), .dout(n10613));
  jnot g10376(.din(n10587), .dout(n10614));
  jnot g10377(.din(n10579), .dout(n10615));
  jnot g10378(.din(n10571), .dout(n10616));
  jnot g10379(.din(n10563), .dout(n10617));
  jnot g10380(.din(n10556), .dout(n10618));
  jnot g10381(.din(n10549), .dout(n10619));
  jnot g10382(.din(n10542), .dout(n10620));
  jnot g10383(.din(n10534), .dout(n10621));
  jnot g10384(.din(n10527), .dout(n10622));
  jnot g10385(.din(n10519), .dout(n10623));
  jnot g10386(.din(n10512), .dout(n10624));
  jnot g10387(.din(n10504), .dout(n10625));
  jnot g10388(.din(n10497), .dout(n10626));
  jnot g10389(.din(n10489), .dout(n10627));
  jnot g10390(.din(n10481), .dout(n10628));
  jnot g10391(.din(n10473), .dout(n10629));
  jnot g10392(.din(n10466), .dout(n10630));
  jnot g10393(.din(n10458), .dout(n10631));
  jnot g10394(.din(n10451), .dout(n10632));
  jnot g10395(.din(n10443), .dout(n10633));
  jnot g10396(.din(n10436), .dout(n10634));
  jnot g10397(.din(n10439), .dout(n10635));
  jnot g10398(.din(n10428), .dout(n10636));
  jnot g10399(.din(n10420), .dout(n10637));
  jnot g10400(.din(n10412), .dout(n10638));
  jnot g10401(.din(n10404), .dout(n10639));
  jnot g10402(.din(n10396), .dout(n10640));
  jnot g10403(.din(n10389), .dout(n10641));
  jnot g10404(.din(n10381), .dout(n10642));
  jnot g10405(.din(n10373), .dout(n10643));
  jnot g10406(.din(n10365), .dout(n10644));
  jnot g10407(.din(n10358), .dout(n10645));
  jnot g10408(.din(n10350), .dout(n10646));
  jnot g10409(.din(n10343), .dout(n10647));
  jnot g10410(.din(n10333), .dout(n10648));
  jnot g10411(.din(n10140), .dout(n10649));
  jnot g10412(.din(n10137), .dout(n10650));
  jor  g10413(.dina(n10328), .dinb(n9834), .dout(n10651));
  jand g10414(.dina(n10651), .dinb(n10650), .dout(n10652));
  jand g10415(.dina(n10652), .dinb(n9832), .dout(n10653));
  jor  g10416(.dina(n10328), .dinb(a[48] ), .dout(n10654));
  jand g10417(.dina(n10654), .dinb(a[49] ), .dout(n10655));
  jand g10418(.dina(asqrt[24] ), .dinb(n9836), .dout(n10656));
  jor  g10419(.dina(n10656), .dinb(n10655), .dout(n10657));
  jor  g10420(.dina(n10657), .dinb(n10653), .dout(n10658));
  jand g10421(.dina(n10658), .dinb(n10649), .dout(n10659));
  jand g10422(.dina(n10659), .dinb(n9369), .dout(n10660));
  jor  g10423(.dina(n10339), .dinb(n10660), .dout(n10661));
  jand g10424(.dina(n10661), .dinb(n10648), .dout(n10662));
  jand g10425(.dina(n10662), .dinb(n8890), .dout(n10663));
  jnot g10426(.din(n10347), .dout(n10664));
  jor  g10427(.dina(n10664), .dinb(n10663), .dout(n10665));
  jand g10428(.dina(n10665), .dinb(n10647), .dout(n10666));
  jand g10429(.dina(n10666), .dinb(n8449), .dout(n10667));
  jor  g10430(.dina(n10354), .dinb(n10667), .dout(n10668));
  jand g10431(.dina(n10668), .dinb(n10646), .dout(n10669));
  jand g10432(.dina(n10669), .dinb(n8003), .dout(n10670));
  jnot g10433(.din(n10362), .dout(n10671));
  jor  g10434(.dina(n10671), .dinb(n10670), .dout(n10672));
  jand g10435(.dina(n10672), .dinb(n10645), .dout(n10673));
  jand g10436(.dina(n10673), .dinb(n7581), .dout(n10674));
  jor  g10437(.dina(n10369), .dinb(n10674), .dout(n10675));
  jand g10438(.dina(n10675), .dinb(n10644), .dout(n10676));
  jand g10439(.dina(n10676), .dinb(n7154), .dout(n10677));
  jor  g10440(.dina(n10377), .dinb(n10677), .dout(n10678));
  jand g10441(.dina(n10678), .dinb(n10643), .dout(n10679));
  jand g10442(.dina(n10679), .dinb(n6758), .dout(n10680));
  jor  g10443(.dina(n10385), .dinb(n10680), .dout(n10681));
  jand g10444(.dina(n10681), .dinb(n10642), .dout(n10682));
  jand g10445(.dina(n10682), .dinb(n6357), .dout(n10683));
  jnot g10446(.din(n10393), .dout(n10684));
  jor  g10447(.dina(n10684), .dinb(n10683), .dout(n10685));
  jand g10448(.dina(n10685), .dinb(n10641), .dout(n10686));
  jand g10449(.dina(n10686), .dinb(n5989), .dout(n10687));
  jor  g10450(.dina(n10400), .dinb(n10687), .dout(n10688));
  jand g10451(.dina(n10688), .dinb(n10640), .dout(n10689));
  jand g10452(.dina(n10689), .dinb(n5606), .dout(n10690));
  jor  g10453(.dina(n10408), .dinb(n10690), .dout(n10691));
  jand g10454(.dina(n10691), .dinb(n10639), .dout(n10692));
  jand g10455(.dina(n10692), .dinb(n5259), .dout(n10693));
  jor  g10456(.dina(n10416), .dinb(n10693), .dout(n10694));
  jand g10457(.dina(n10694), .dinb(n10638), .dout(n10695));
  jand g10458(.dina(n10695), .dinb(n4902), .dout(n10696));
  jor  g10459(.dina(n10424), .dinb(n10696), .dout(n10697));
  jand g10460(.dina(n10697), .dinb(n10637), .dout(n10698));
  jand g10461(.dina(n10698), .dinb(n4582), .dout(n10699));
  jor  g10462(.dina(n10432), .dinb(n10699), .dout(n10700));
  jand g10463(.dina(n10700), .dinb(n10636), .dout(n10701));
  jand g10464(.dina(n10701), .dinb(n4249), .dout(n10702));
  jor  g10465(.dina(n10702), .dinb(n10635), .dout(n10703));
  jand g10466(.dina(n10703), .dinb(n10634), .dout(n10704));
  jand g10467(.dina(n10704), .dinb(n3955), .dout(n10705));
  jor  g10468(.dina(n10447), .dinb(n10705), .dout(n10706));
  jand g10469(.dina(n10706), .dinb(n10633), .dout(n10707));
  jand g10470(.dina(n10707), .dinb(n3642), .dout(n10708));
  jnot g10471(.din(n10455), .dout(n10709));
  jor  g10472(.dina(n10709), .dinb(n10708), .dout(n10710));
  jand g10473(.dina(n10710), .dinb(n10632), .dout(n10711));
  jand g10474(.dina(n10711), .dinb(n3368), .dout(n10712));
  jor  g10475(.dina(n10462), .dinb(n10712), .dout(n10713));
  jand g10476(.dina(n10713), .dinb(n10631), .dout(n10714));
  jand g10477(.dina(n10714), .dinb(n3089), .dout(n10715));
  jnot g10478(.din(n10470), .dout(n10716));
  jor  g10479(.dina(n10716), .dinb(n10715), .dout(n10717));
  jand g10480(.dina(n10717), .dinb(n10630), .dout(n10718));
  jand g10481(.dina(n10718), .dinb(n2833), .dout(n10719));
  jor  g10482(.dina(n10477), .dinb(n10719), .dout(n10720));
  jand g10483(.dina(n10720), .dinb(n10629), .dout(n10721));
  jand g10484(.dina(n10721), .dinb(n2572), .dout(n10722));
  jor  g10485(.dina(n10485), .dinb(n10722), .dout(n10723));
  jand g10486(.dina(n10723), .dinb(n10628), .dout(n10724));
  jand g10487(.dina(n10724), .dinb(n2345), .dout(n10725));
  jor  g10488(.dina(n10493), .dinb(n10725), .dout(n10726));
  jand g10489(.dina(n10726), .dinb(n10627), .dout(n10727));
  jand g10490(.dina(n10727), .dinb(n2108), .dout(n10728));
  jnot g10491(.din(n10501), .dout(n10729));
  jor  g10492(.dina(n10729), .dinb(n10728), .dout(n10730));
  jand g10493(.dina(n10730), .dinb(n10626), .dout(n10731));
  jand g10494(.dina(n10731), .dinb(n1912), .dout(n10732));
  jor  g10495(.dina(n10508), .dinb(n10732), .dout(n10733));
  jand g10496(.dina(n10733), .dinb(n10625), .dout(n10734));
  jand g10497(.dina(n10734), .dinb(n1699), .dout(n10735));
  jnot g10498(.din(n10516), .dout(n10736));
  jor  g10499(.dina(n10736), .dinb(n10735), .dout(n10737));
  jand g10500(.dina(n10737), .dinb(n10624), .dout(n10738));
  jand g10501(.dina(n10738), .dinb(n1516), .dout(n10739));
  jor  g10502(.dina(n10523), .dinb(n10739), .dout(n10740));
  jand g10503(.dina(n10740), .dinb(n10623), .dout(n10741));
  jand g10504(.dina(n10741), .dinb(n1332), .dout(n10742));
  jnot g10505(.din(n10531), .dout(n10743));
  jor  g10506(.dina(n10743), .dinb(n10742), .dout(n10744));
  jand g10507(.dina(n10744), .dinb(n10622), .dout(n10745));
  jand g10508(.dina(n10745), .dinb(n1173), .dout(n10746));
  jor  g10509(.dina(n10538), .dinb(n10746), .dout(n10747));
  jand g10510(.dina(n10747), .dinb(n10621), .dout(n10748));
  jand g10511(.dina(n10748), .dinb(n1008), .dout(n10749));
  jnot g10512(.din(n10546), .dout(n10750));
  jor  g10513(.dina(n10750), .dinb(n10749), .dout(n10751));
  jand g10514(.dina(n10751), .dinb(n10620), .dout(n10752));
  jand g10515(.dina(n10752), .dinb(n884), .dout(n10753));
  jnot g10516(.din(n10553), .dout(n10754));
  jor  g10517(.dina(n10754), .dinb(n10753), .dout(n10755));
  jand g10518(.dina(n10755), .dinb(n10619), .dout(n10756));
  jand g10519(.dina(n10756), .dinb(n743), .dout(n10757));
  jnot g10520(.din(n10560), .dout(n10758));
  jor  g10521(.dina(n10758), .dinb(n10757), .dout(n10759));
  jand g10522(.dina(n10759), .dinb(n10618), .dout(n10760));
  jand g10523(.dina(n10760), .dinb(n635), .dout(n10761));
  jor  g10524(.dina(n10567), .dinb(n10761), .dout(n10762));
  jand g10525(.dina(n10762), .dinb(n10617), .dout(n10763));
  jand g10526(.dina(n10763), .dinb(n515), .dout(n10764));
  jor  g10527(.dina(n10575), .dinb(n10764), .dout(n10765));
  jand g10528(.dina(n10765), .dinb(n10616), .dout(n10766));
  jand g10529(.dina(n10766), .dinb(n443), .dout(n10767));
  jor  g10530(.dina(n10583), .dinb(n10767), .dout(n10768));
  jand g10531(.dina(n10768), .dinb(n10615), .dout(n10769));
  jand g10532(.dina(n10769), .dinb(n352), .dout(n10770));
  jnot g10533(.din(n10591), .dout(n10771));
  jor  g10534(.dina(n10771), .dinb(n10770), .dout(n10772));
  jand g10535(.dina(n10772), .dinb(n10614), .dout(n10773));
  jand g10536(.dina(n10773), .dinb(n294), .dout(n10774));
  jor  g10537(.dina(n10598), .dinb(n10774), .dout(n10775));
  jand g10538(.dina(n10775), .dinb(n10613), .dout(n10776));
  jand g10539(.dina(n10776), .dinb(n239), .dout(n10777));
  jor  g10540(.dina(n10606), .dinb(n10777), .dout(n10778));
  jand g10541(.dina(n10778), .dinb(n10612), .dout(n10779));
  jand g10542(.dina(n10779), .dinb(n221), .dout(n10780));
  jxor g10543(.dina(n10101), .dinb(n239), .dout(n10781));
  jand g10544(.dina(n10781), .dinb(asqrt[24] ), .dout(n10782));
  jxor g10545(.dina(n10782), .dinb(n10106), .dout(n10783));
  jor  g10546(.dina(n10783), .dinb(n10780), .dout(n10784));
  jand g10547(.dina(n10784), .dinb(n10611), .dout(n10785));
  jxor g10548(.dina(n10108), .dinb(n221), .dout(n10786));
  jand g10549(.dina(n10786), .dinb(asqrt[24] ), .dout(n10787));
  jxor g10550(.dina(n10787), .dinb(n10114), .dout(n10788));
  jor  g10551(.dina(n10788), .dinb(n10785), .dout(n10789));
  jand g10552(.dina(asqrt[24] ), .dinb(n10323), .dout(n10790));
  jor  g10553(.dina(n10790), .dinb(n10125), .dout(n10791));
  jor  g10554(.dina(n10791), .dinb(n10789), .dout(n10792));
  jand g10555(.dina(n10792), .dinb(n218), .dout(n10793));
  jand g10556(.dina(n10328), .dinb(n10119), .dout(n10794));
  jand g10557(.dina(n10788), .dinb(n10785), .dout(n10795));
  jor  g10558(.dina(n10795), .dinb(n10794), .dout(n10796));
  jand g10559(.dina(n10328), .dinb(n10116), .dout(n10797));
  jnot g10560(.din(n10797), .dout(n10798));
  jnot g10561(.din(n10125), .dout(n10799));
  jand g10562(.dina(n10120), .dinb(asqrt[63] ), .dout(n10800));
  jand g10563(.dina(n10800), .dinb(n10799), .dout(n10801));
  jand g10564(.dina(n10801), .dinb(n10798), .dout(n10802));
  jor  g10565(.dina(n10802), .dinb(n10796), .dout(n10803));
  jor  g10566(.dina(n10803), .dinb(n10793), .dout(asqrt[23] ));
  jnot g10567(.din(a[44] ), .dout(n10805));
  jnot g10568(.din(a[45] ), .dout(n10806));
  jand g10569(.dina(n10806), .dinb(n10805), .dout(n10807));
  jand g10570(.dina(n10807), .dinb(n10134), .dout(n10808));
  jnot g10571(.din(n10808), .dout(n10809));
  jor  g10572(.dina(n10609), .dinb(asqrt[62] ), .dout(n10810));
  jnot g10573(.din(n10783), .dout(n10811));
  jand g10574(.dina(n10811), .dinb(n10810), .dout(n10812));
  jor  g10575(.dina(n10812), .dinb(n10610), .dout(n10813));
  jnot g10576(.din(n10788), .dout(n10814));
  jand g10577(.dina(n10814), .dinb(n10813), .dout(n10815));
  jnot g10578(.din(n10791), .dout(n10816));
  jand g10579(.dina(n10816), .dinb(n10815), .dout(n10817));
  jor  g10580(.dina(n10817), .dinb(asqrt[63] ), .dout(n10818));
  jnot g10581(.din(n10794), .dout(n10819));
  jor  g10582(.dina(n10814), .dinb(n10813), .dout(n10820));
  jand g10583(.dina(n10820), .dinb(n10819), .dout(n10821));
  jnot g10584(.din(n10802), .dout(n10822));
  jand g10585(.dina(n10822), .dinb(n10821), .dout(n10823));
  jand g10586(.dina(n10823), .dinb(n10818), .dout(n10824));
  jor  g10587(.dina(n10824), .dinb(n10134), .dout(n10825));
  jand g10588(.dina(n10825), .dinb(n10809), .dout(n10826));
  jor  g10589(.dina(n10826), .dinb(n10328), .dout(n10827));
  jand g10590(.dina(n10826), .dinb(n10328), .dout(n10828));
  jor  g10591(.dina(n10824), .dinb(a[46] ), .dout(n10829));
  jand g10592(.dina(n10829), .dinb(a[47] ), .dout(n10830));
  jand g10593(.dina(asqrt[23] ), .dinb(n10136), .dout(n10831));
  jor  g10594(.dina(n10831), .dinb(n10830), .dout(n10832));
  jor  g10595(.dina(n10832), .dinb(n10828), .dout(n10833));
  jand g10596(.dina(n10833), .dinb(n10827), .dout(n10834));
  jor  g10597(.dina(n10834), .dinb(n9832), .dout(n10835));
  jand g10598(.dina(n10834), .dinb(n9832), .dout(n10836));
  jnot g10599(.din(n10136), .dout(n10837));
  jor  g10600(.dina(n10824), .dinb(n10837), .dout(n10838));
  jor  g10601(.dina(n10801), .dinb(n10328), .dout(n10839));
  jor  g10602(.dina(n10839), .dinb(n10795), .dout(n10840));
  jor  g10603(.dina(n10840), .dinb(n10793), .dout(n10841));
  jand g10604(.dina(n10841), .dinb(n10838), .dout(n10842));
  jxor g10605(.dina(n10842), .dinb(n9834), .dout(n10843));
  jor  g10606(.dina(n10843), .dinb(n10836), .dout(n10844));
  jand g10607(.dina(n10844), .dinb(n10835), .dout(n10845));
  jor  g10608(.dina(n10845), .dinb(n9369), .dout(n10846));
  jand g10609(.dina(n10845), .dinb(n9369), .dout(n10847));
  jxor g10610(.dina(n10139), .dinb(n9832), .dout(n10848));
  jor  g10611(.dina(n10848), .dinb(n10824), .dout(n10849));
  jxor g10612(.dina(n10849), .dinb(n10330), .dout(n10850));
  jor  g10613(.dina(n10850), .dinb(n10847), .dout(n10851));
  jand g10614(.dina(n10851), .dinb(n10846), .dout(n10852));
  jor  g10615(.dina(n10852), .dinb(n8890), .dout(n10853));
  jand g10616(.dina(n10852), .dinb(n8890), .dout(n10854));
  jxor g10617(.dina(n10332), .dinb(n9369), .dout(n10855));
  jor  g10618(.dina(n10855), .dinb(n10824), .dout(n10856));
  jxor g10619(.dina(n10856), .dinb(n10340), .dout(n10857));
  jor  g10620(.dina(n10857), .dinb(n10854), .dout(n10858));
  jand g10621(.dina(n10858), .dinb(n10853), .dout(n10859));
  jor  g10622(.dina(n10859), .dinb(n8449), .dout(n10860));
  jand g10623(.dina(n10859), .dinb(n8449), .dout(n10861));
  jxor g10624(.dina(n10342), .dinb(n8890), .dout(n10862));
  jor  g10625(.dina(n10862), .dinb(n10824), .dout(n10863));
  jxor g10626(.dina(n10863), .dinb(n10664), .dout(n10864));
  jnot g10627(.din(n10864), .dout(n10865));
  jor  g10628(.dina(n10865), .dinb(n10861), .dout(n10866));
  jand g10629(.dina(n10866), .dinb(n10860), .dout(n10867));
  jor  g10630(.dina(n10867), .dinb(n8003), .dout(n10868));
  jand g10631(.dina(n10867), .dinb(n8003), .dout(n10869));
  jxor g10632(.dina(n10349), .dinb(n8449), .dout(n10870));
  jor  g10633(.dina(n10870), .dinb(n10824), .dout(n10871));
  jxor g10634(.dina(n10871), .dinb(n10355), .dout(n10872));
  jor  g10635(.dina(n10872), .dinb(n10869), .dout(n10873));
  jand g10636(.dina(n10873), .dinb(n10868), .dout(n10874));
  jor  g10637(.dina(n10874), .dinb(n7581), .dout(n10875));
  jand g10638(.dina(n10874), .dinb(n7581), .dout(n10876));
  jxor g10639(.dina(n10357), .dinb(n8003), .dout(n10877));
  jor  g10640(.dina(n10877), .dinb(n10824), .dout(n10878));
  jxor g10641(.dina(n10878), .dinb(n10671), .dout(n10879));
  jnot g10642(.din(n10879), .dout(n10880));
  jor  g10643(.dina(n10880), .dinb(n10876), .dout(n10881));
  jand g10644(.dina(n10881), .dinb(n10875), .dout(n10882));
  jor  g10645(.dina(n10882), .dinb(n7154), .dout(n10883));
  jand g10646(.dina(n10882), .dinb(n7154), .dout(n10884));
  jxor g10647(.dina(n10364), .dinb(n7581), .dout(n10885));
  jor  g10648(.dina(n10885), .dinb(n10824), .dout(n10886));
  jxor g10649(.dina(n10886), .dinb(n10370), .dout(n10887));
  jor  g10650(.dina(n10887), .dinb(n10884), .dout(n10888));
  jand g10651(.dina(n10888), .dinb(n10883), .dout(n10889));
  jor  g10652(.dina(n10889), .dinb(n6758), .dout(n10890));
  jand g10653(.dina(n10889), .dinb(n6758), .dout(n10891));
  jxor g10654(.dina(n10372), .dinb(n7154), .dout(n10892));
  jor  g10655(.dina(n10892), .dinb(n10824), .dout(n10893));
  jxor g10656(.dina(n10893), .dinb(n10378), .dout(n10894));
  jor  g10657(.dina(n10894), .dinb(n10891), .dout(n10895));
  jand g10658(.dina(n10895), .dinb(n10890), .dout(n10896));
  jor  g10659(.dina(n10896), .dinb(n6357), .dout(n10897));
  jand g10660(.dina(n10896), .dinb(n6357), .dout(n10898));
  jxor g10661(.dina(n10380), .dinb(n6758), .dout(n10899));
  jor  g10662(.dina(n10899), .dinb(n10824), .dout(n10900));
  jxor g10663(.dina(n10900), .dinb(n10386), .dout(n10901));
  jor  g10664(.dina(n10901), .dinb(n10898), .dout(n10902));
  jand g10665(.dina(n10902), .dinb(n10897), .dout(n10903));
  jor  g10666(.dina(n10903), .dinb(n5989), .dout(n10904));
  jand g10667(.dina(n10903), .dinb(n5989), .dout(n10905));
  jxor g10668(.dina(n10388), .dinb(n6357), .dout(n10906));
  jor  g10669(.dina(n10906), .dinb(n10824), .dout(n10907));
  jxor g10670(.dina(n10907), .dinb(n10684), .dout(n10908));
  jnot g10671(.din(n10908), .dout(n10909));
  jor  g10672(.dina(n10909), .dinb(n10905), .dout(n10910));
  jand g10673(.dina(n10910), .dinb(n10904), .dout(n10911));
  jor  g10674(.dina(n10911), .dinb(n5606), .dout(n10912));
  jand g10675(.dina(n10911), .dinb(n5606), .dout(n10913));
  jxor g10676(.dina(n10395), .dinb(n5989), .dout(n10914));
  jor  g10677(.dina(n10914), .dinb(n10824), .dout(n10915));
  jxor g10678(.dina(n10915), .dinb(n10401), .dout(n10916));
  jor  g10679(.dina(n10916), .dinb(n10913), .dout(n10917));
  jand g10680(.dina(n10917), .dinb(n10912), .dout(n10918));
  jor  g10681(.dina(n10918), .dinb(n5259), .dout(n10919));
  jand g10682(.dina(n10918), .dinb(n5259), .dout(n10920));
  jxor g10683(.dina(n10403), .dinb(n5606), .dout(n10921));
  jor  g10684(.dina(n10921), .dinb(n10824), .dout(n10922));
  jxor g10685(.dina(n10922), .dinb(n10409), .dout(n10923));
  jor  g10686(.dina(n10923), .dinb(n10920), .dout(n10924));
  jand g10687(.dina(n10924), .dinb(n10919), .dout(n10925));
  jor  g10688(.dina(n10925), .dinb(n4902), .dout(n10926));
  jand g10689(.dina(n10925), .dinb(n4902), .dout(n10927));
  jxor g10690(.dina(n10411), .dinb(n5259), .dout(n10928));
  jor  g10691(.dina(n10928), .dinb(n10824), .dout(n10929));
  jxor g10692(.dina(n10929), .dinb(n10417), .dout(n10930));
  jor  g10693(.dina(n10930), .dinb(n10927), .dout(n10931));
  jand g10694(.dina(n10931), .dinb(n10926), .dout(n10932));
  jor  g10695(.dina(n10932), .dinb(n4582), .dout(n10933));
  jand g10696(.dina(n10932), .dinb(n4582), .dout(n10934));
  jxor g10697(.dina(n10419), .dinb(n4902), .dout(n10935));
  jor  g10698(.dina(n10935), .dinb(n10824), .dout(n10936));
  jxor g10699(.dina(n10936), .dinb(n10425), .dout(n10937));
  jor  g10700(.dina(n10937), .dinb(n10934), .dout(n10938));
  jand g10701(.dina(n10938), .dinb(n10933), .dout(n10939));
  jor  g10702(.dina(n10939), .dinb(n4249), .dout(n10940));
  jand g10703(.dina(n10939), .dinb(n4249), .dout(n10941));
  jxor g10704(.dina(n10427), .dinb(n4582), .dout(n10942));
  jor  g10705(.dina(n10942), .dinb(n10824), .dout(n10943));
  jxor g10706(.dina(n10943), .dinb(n10433), .dout(n10944));
  jor  g10707(.dina(n10944), .dinb(n10941), .dout(n10945));
  jand g10708(.dina(n10945), .dinb(n10940), .dout(n10946));
  jor  g10709(.dina(n10946), .dinb(n3955), .dout(n10947));
  jxor g10710(.dina(n10435), .dinb(n4249), .dout(n10948));
  jor  g10711(.dina(n10948), .dinb(n10824), .dout(n10949));
  jxor g10712(.dina(n10949), .dinb(n10635), .dout(n10950));
  jnot g10713(.din(n10950), .dout(n10951));
  jand g10714(.dina(n10946), .dinb(n3955), .dout(n10952));
  jor  g10715(.dina(n10952), .dinb(n10951), .dout(n10953));
  jand g10716(.dina(n10953), .dinb(n10947), .dout(n10954));
  jor  g10717(.dina(n10954), .dinb(n3642), .dout(n10955));
  jand g10718(.dina(n10954), .dinb(n3642), .dout(n10956));
  jxor g10719(.dina(n10442), .dinb(n3955), .dout(n10957));
  jor  g10720(.dina(n10957), .dinb(n10824), .dout(n10958));
  jxor g10721(.dina(n10958), .dinb(n10448), .dout(n10959));
  jor  g10722(.dina(n10959), .dinb(n10956), .dout(n10960));
  jand g10723(.dina(n10960), .dinb(n10955), .dout(n10961));
  jor  g10724(.dina(n10961), .dinb(n3368), .dout(n10962));
  jand g10725(.dina(n10961), .dinb(n3368), .dout(n10963));
  jxor g10726(.dina(n10450), .dinb(n3642), .dout(n10964));
  jor  g10727(.dina(n10964), .dinb(n10824), .dout(n10965));
  jxor g10728(.dina(n10965), .dinb(n10709), .dout(n10966));
  jnot g10729(.din(n10966), .dout(n10967));
  jor  g10730(.dina(n10967), .dinb(n10963), .dout(n10968));
  jand g10731(.dina(n10968), .dinb(n10962), .dout(n10969));
  jor  g10732(.dina(n10969), .dinb(n3089), .dout(n10970));
  jand g10733(.dina(n10969), .dinb(n3089), .dout(n10971));
  jxor g10734(.dina(n10457), .dinb(n3368), .dout(n10972));
  jor  g10735(.dina(n10972), .dinb(n10824), .dout(n10973));
  jxor g10736(.dina(n10973), .dinb(n10463), .dout(n10974));
  jor  g10737(.dina(n10974), .dinb(n10971), .dout(n10975));
  jand g10738(.dina(n10975), .dinb(n10970), .dout(n10976));
  jor  g10739(.dina(n10976), .dinb(n2833), .dout(n10977));
  jand g10740(.dina(n10976), .dinb(n2833), .dout(n10978));
  jxor g10741(.dina(n10465), .dinb(n3089), .dout(n10979));
  jor  g10742(.dina(n10979), .dinb(n10824), .dout(n10980));
  jxor g10743(.dina(n10980), .dinb(n10716), .dout(n10981));
  jnot g10744(.din(n10981), .dout(n10982));
  jor  g10745(.dina(n10982), .dinb(n10978), .dout(n10983));
  jand g10746(.dina(n10983), .dinb(n10977), .dout(n10984));
  jor  g10747(.dina(n10984), .dinb(n2572), .dout(n10985));
  jand g10748(.dina(n10984), .dinb(n2572), .dout(n10986));
  jxor g10749(.dina(n10472), .dinb(n2833), .dout(n10987));
  jor  g10750(.dina(n10987), .dinb(n10824), .dout(n10988));
  jxor g10751(.dina(n10988), .dinb(n10478), .dout(n10989));
  jor  g10752(.dina(n10989), .dinb(n10986), .dout(n10990));
  jand g10753(.dina(n10990), .dinb(n10985), .dout(n10991));
  jor  g10754(.dina(n10991), .dinb(n2345), .dout(n10992));
  jand g10755(.dina(n10991), .dinb(n2345), .dout(n10993));
  jxor g10756(.dina(n10480), .dinb(n2572), .dout(n10994));
  jor  g10757(.dina(n10994), .dinb(n10824), .dout(n10995));
  jxor g10758(.dina(n10995), .dinb(n10486), .dout(n10996));
  jor  g10759(.dina(n10996), .dinb(n10993), .dout(n10997));
  jand g10760(.dina(n10997), .dinb(n10992), .dout(n10998));
  jor  g10761(.dina(n10998), .dinb(n2108), .dout(n10999));
  jand g10762(.dina(n10998), .dinb(n2108), .dout(n11000));
  jxor g10763(.dina(n10488), .dinb(n2345), .dout(n11001));
  jor  g10764(.dina(n11001), .dinb(n10824), .dout(n11002));
  jxor g10765(.dina(n11002), .dinb(n10494), .dout(n11003));
  jor  g10766(.dina(n11003), .dinb(n11000), .dout(n11004));
  jand g10767(.dina(n11004), .dinb(n10999), .dout(n11005));
  jor  g10768(.dina(n11005), .dinb(n1912), .dout(n11006));
  jand g10769(.dina(n11005), .dinb(n1912), .dout(n11007));
  jxor g10770(.dina(n10496), .dinb(n2108), .dout(n11008));
  jor  g10771(.dina(n11008), .dinb(n10824), .dout(n11009));
  jxor g10772(.dina(n11009), .dinb(n10729), .dout(n11010));
  jnot g10773(.din(n11010), .dout(n11011));
  jor  g10774(.dina(n11011), .dinb(n11007), .dout(n11012));
  jand g10775(.dina(n11012), .dinb(n11006), .dout(n11013));
  jor  g10776(.dina(n11013), .dinb(n1699), .dout(n11014));
  jand g10777(.dina(n11013), .dinb(n1699), .dout(n11015));
  jxor g10778(.dina(n10503), .dinb(n1912), .dout(n11016));
  jor  g10779(.dina(n11016), .dinb(n10824), .dout(n11017));
  jxor g10780(.dina(n11017), .dinb(n10509), .dout(n11018));
  jor  g10781(.dina(n11018), .dinb(n11015), .dout(n11019));
  jand g10782(.dina(n11019), .dinb(n11014), .dout(n11020));
  jor  g10783(.dina(n11020), .dinb(n1516), .dout(n11021));
  jand g10784(.dina(n11020), .dinb(n1516), .dout(n11022));
  jxor g10785(.dina(n10511), .dinb(n1699), .dout(n11023));
  jor  g10786(.dina(n11023), .dinb(n10824), .dout(n11024));
  jxor g10787(.dina(n11024), .dinb(n10736), .dout(n11025));
  jnot g10788(.din(n11025), .dout(n11026));
  jor  g10789(.dina(n11026), .dinb(n11022), .dout(n11027));
  jand g10790(.dina(n11027), .dinb(n11021), .dout(n11028));
  jor  g10791(.dina(n11028), .dinb(n1332), .dout(n11029));
  jand g10792(.dina(n11028), .dinb(n1332), .dout(n11030));
  jxor g10793(.dina(n10518), .dinb(n1516), .dout(n11031));
  jor  g10794(.dina(n11031), .dinb(n10824), .dout(n11032));
  jxor g10795(.dina(n11032), .dinb(n10524), .dout(n11033));
  jor  g10796(.dina(n11033), .dinb(n11030), .dout(n11034));
  jand g10797(.dina(n11034), .dinb(n11029), .dout(n11035));
  jor  g10798(.dina(n11035), .dinb(n1173), .dout(n11036));
  jand g10799(.dina(n11035), .dinb(n1173), .dout(n11037));
  jxor g10800(.dina(n10526), .dinb(n1332), .dout(n11038));
  jor  g10801(.dina(n11038), .dinb(n10824), .dout(n11039));
  jxor g10802(.dina(n11039), .dinb(n10743), .dout(n11040));
  jnot g10803(.din(n11040), .dout(n11041));
  jor  g10804(.dina(n11041), .dinb(n11037), .dout(n11042));
  jand g10805(.dina(n11042), .dinb(n11036), .dout(n11043));
  jor  g10806(.dina(n11043), .dinb(n1008), .dout(n11044));
  jand g10807(.dina(n11043), .dinb(n1008), .dout(n11045));
  jxor g10808(.dina(n10533), .dinb(n1173), .dout(n11046));
  jor  g10809(.dina(n11046), .dinb(n10824), .dout(n11047));
  jxor g10810(.dina(n11047), .dinb(n10539), .dout(n11048));
  jor  g10811(.dina(n11048), .dinb(n11045), .dout(n11049));
  jand g10812(.dina(n11049), .dinb(n11044), .dout(n11050));
  jor  g10813(.dina(n11050), .dinb(n884), .dout(n11051));
  jand g10814(.dina(n11050), .dinb(n884), .dout(n11052));
  jxor g10815(.dina(n10541), .dinb(n1008), .dout(n11053));
  jor  g10816(.dina(n11053), .dinb(n10824), .dout(n11054));
  jxor g10817(.dina(n11054), .dinb(n10750), .dout(n11055));
  jnot g10818(.din(n11055), .dout(n11056));
  jor  g10819(.dina(n11056), .dinb(n11052), .dout(n11057));
  jand g10820(.dina(n11057), .dinb(n11051), .dout(n11058));
  jor  g10821(.dina(n11058), .dinb(n743), .dout(n11059));
  jand g10822(.dina(n11058), .dinb(n743), .dout(n11060));
  jxor g10823(.dina(n10548), .dinb(n884), .dout(n11061));
  jor  g10824(.dina(n11061), .dinb(n10824), .dout(n11062));
  jxor g10825(.dina(n11062), .dinb(n10754), .dout(n11063));
  jnot g10826(.din(n11063), .dout(n11064));
  jor  g10827(.dina(n11064), .dinb(n11060), .dout(n11065));
  jand g10828(.dina(n11065), .dinb(n11059), .dout(n11066));
  jor  g10829(.dina(n11066), .dinb(n635), .dout(n11067));
  jand g10830(.dina(n11066), .dinb(n635), .dout(n11068));
  jxor g10831(.dina(n10555), .dinb(n743), .dout(n11069));
  jor  g10832(.dina(n11069), .dinb(n10824), .dout(n11070));
  jxor g10833(.dina(n11070), .dinb(n10758), .dout(n11071));
  jnot g10834(.din(n11071), .dout(n11072));
  jor  g10835(.dina(n11072), .dinb(n11068), .dout(n11073));
  jand g10836(.dina(n11073), .dinb(n11067), .dout(n11074));
  jor  g10837(.dina(n11074), .dinb(n515), .dout(n11075));
  jand g10838(.dina(n11074), .dinb(n515), .dout(n11076));
  jxor g10839(.dina(n10562), .dinb(n635), .dout(n11077));
  jor  g10840(.dina(n11077), .dinb(n10824), .dout(n11078));
  jxor g10841(.dina(n11078), .dinb(n10568), .dout(n11079));
  jor  g10842(.dina(n11079), .dinb(n11076), .dout(n11080));
  jand g10843(.dina(n11080), .dinb(n11075), .dout(n11081));
  jor  g10844(.dina(n11081), .dinb(n443), .dout(n11082));
  jand g10845(.dina(n11081), .dinb(n443), .dout(n11083));
  jxor g10846(.dina(n10570), .dinb(n515), .dout(n11084));
  jor  g10847(.dina(n11084), .dinb(n10824), .dout(n11085));
  jxor g10848(.dina(n11085), .dinb(n10576), .dout(n11086));
  jor  g10849(.dina(n11086), .dinb(n11083), .dout(n11087));
  jand g10850(.dina(n11087), .dinb(n11082), .dout(n11088));
  jor  g10851(.dina(n11088), .dinb(n352), .dout(n11089));
  jand g10852(.dina(n11088), .dinb(n352), .dout(n11090));
  jxor g10853(.dina(n10578), .dinb(n443), .dout(n11091));
  jor  g10854(.dina(n11091), .dinb(n10824), .dout(n11092));
  jxor g10855(.dina(n11092), .dinb(n10584), .dout(n11093));
  jor  g10856(.dina(n11093), .dinb(n11090), .dout(n11094));
  jand g10857(.dina(n11094), .dinb(n11089), .dout(n11095));
  jor  g10858(.dina(n11095), .dinb(n294), .dout(n11096));
  jand g10859(.dina(n11095), .dinb(n294), .dout(n11097));
  jxor g10860(.dina(n10586), .dinb(n352), .dout(n11098));
  jor  g10861(.dina(n11098), .dinb(n10824), .dout(n11099));
  jxor g10862(.dina(n11099), .dinb(n10771), .dout(n11100));
  jnot g10863(.din(n11100), .dout(n11101));
  jor  g10864(.dina(n11101), .dinb(n11097), .dout(n11102));
  jand g10865(.dina(n11102), .dinb(n11096), .dout(n11103));
  jor  g10866(.dina(n11103), .dinb(n239), .dout(n11104));
  jand g10867(.dina(n11103), .dinb(n239), .dout(n11105));
  jxor g10868(.dina(n10593), .dinb(n294), .dout(n11106));
  jor  g10869(.dina(n11106), .dinb(n10824), .dout(n11107));
  jxor g10870(.dina(n11107), .dinb(n10599), .dout(n11108));
  jor  g10871(.dina(n11108), .dinb(n11105), .dout(n11109));
  jand g10872(.dina(n11109), .dinb(n11104), .dout(n11110));
  jor  g10873(.dina(n11110), .dinb(n221), .dout(n11111));
  jand g10874(.dina(n11110), .dinb(n221), .dout(n11112));
  jxor g10875(.dina(n10601), .dinb(n239), .dout(n11113));
  jor  g10876(.dina(n11113), .dinb(n10824), .dout(n11114));
  jxor g10877(.dina(n11114), .dinb(n10607), .dout(n11115));
  jor  g10878(.dina(n11115), .dinb(n11112), .dout(n11116));
  jand g10879(.dina(n11116), .dinb(n11111), .dout(n11117));
  jxor g10880(.dina(n10609), .dinb(n221), .dout(n11118));
  jor  g10881(.dina(n11118), .dinb(n10824), .dout(n11119));
  jxor g10882(.dina(n11119), .dinb(n10811), .dout(n11120));
  jand g10883(.dina(n11120), .dinb(n11117), .dout(n11121));
  jand g10884(.dina(n10824), .dinb(n10785), .dout(n11122));
  jand g10885(.dina(n10789), .dinb(asqrt[63] ), .dout(n11123));
  jand g10886(.dina(n11123), .dinb(n10820), .dout(n11124));
  jnot g10887(.din(n11124), .dout(n11125));
  jor  g10888(.dina(n11125), .dinb(n11122), .dout(n11126));
  jnot g10889(.din(n11126), .dout(n11127));
  jand g10890(.dina(asqrt[23] ), .dinb(n10815), .dout(n11128));
  jor  g10891(.dina(n11120), .dinb(n11117), .dout(n11129));
  jor  g10892(.dina(n11129), .dinb(n10795), .dout(n11130));
  jor  g10893(.dina(n11130), .dinb(n11128), .dout(n11131));
  jand g10894(.dina(n11131), .dinb(n218), .dout(n11132));
  jand g10895(.dina(n10824), .dinb(n10788), .dout(n11133));
  jor  g10896(.dina(n11133), .dinb(n11132), .dout(n11134));
  jor  g10897(.dina(n11134), .dinb(n11127), .dout(n11135));
  jor  g10898(.dina(n11135), .dinb(n11121), .dout(asqrt[22] ));
  jnot g10899(.din(n11115), .dout(n11137));
  jxor g10900(.dina(n11110), .dinb(n221), .dout(n11138));
  jand g10901(.dina(n11138), .dinb(asqrt[22] ), .dout(n11139));
  jxor g10902(.dina(n11139), .dinb(n11137), .dout(n11140));
  jand g10903(.dina(asqrt[22] ), .dinb(a[44] ), .dout(n11141));
  jnot g10904(.din(a[42] ), .dout(n11142));
  jnot g10905(.din(a[43] ), .dout(n11143));
  jand g10906(.dina(n11143), .dinb(n11142), .dout(n11144));
  jand g10907(.dina(n11144), .dinb(n10805), .dout(n11145));
  jor  g10908(.dina(n11145), .dinb(n11141), .dout(n11146));
  jand g10909(.dina(n11146), .dinb(asqrt[23] ), .dout(n11147));
  jor  g10910(.dina(n11146), .dinb(asqrt[23] ), .dout(n11148));
  jand g10911(.dina(asqrt[22] ), .dinb(n10805), .dout(n11149));
  jor  g10912(.dina(n11149), .dinb(n10806), .dout(n11150));
  jnot g10913(.din(n10807), .dout(n11151));
  jnot g10914(.din(n11121), .dout(n11152));
  jnot g10915(.din(n11128), .dout(n11153));
  jnot g10916(.din(n11111), .dout(n11154));
  jnot g10917(.din(n11104), .dout(n11155));
  jnot g10918(.din(n11096), .dout(n11156));
  jnot g10919(.din(n11089), .dout(n11157));
  jnot g10920(.din(n11082), .dout(n11158));
  jnot g10921(.din(n11075), .dout(n11159));
  jnot g10922(.din(n11067), .dout(n11160));
  jnot g10923(.din(n11059), .dout(n11161));
  jnot g10924(.din(n11051), .dout(n11162));
  jnot g10925(.din(n11044), .dout(n11163));
  jnot g10926(.din(n11036), .dout(n11164));
  jnot g10927(.din(n11029), .dout(n11165));
  jnot g10928(.din(n11021), .dout(n11166));
  jnot g10929(.din(n11014), .dout(n11167));
  jnot g10930(.din(n11006), .dout(n11168));
  jnot g10931(.din(n10999), .dout(n11169));
  jnot g10932(.din(n10992), .dout(n11170));
  jnot g10933(.din(n10985), .dout(n11171));
  jnot g10934(.din(n10977), .dout(n11172));
  jnot g10935(.din(n10970), .dout(n11173));
  jnot g10936(.din(n10962), .dout(n11174));
  jnot g10937(.din(n10955), .dout(n11175));
  jnot g10938(.din(n10947), .dout(n11176));
  jnot g10939(.din(n10940), .dout(n11177));
  jnot g10940(.din(n10933), .dout(n11178));
  jnot g10941(.din(n10926), .dout(n11179));
  jnot g10942(.din(n10919), .dout(n11180));
  jnot g10943(.din(n10912), .dout(n11181));
  jnot g10944(.din(n10904), .dout(n11182));
  jnot g10945(.din(n10897), .dout(n11183));
  jnot g10946(.din(n10890), .dout(n11184));
  jnot g10947(.din(n10883), .dout(n11185));
  jnot g10948(.din(n10875), .dout(n11186));
  jnot g10949(.din(n10868), .dout(n11187));
  jnot g10950(.din(n10860), .dout(n11188));
  jnot g10951(.din(n10853), .dout(n11189));
  jnot g10952(.din(n10846), .dout(n11190));
  jnot g10953(.din(n10835), .dout(n11191));
  jnot g10954(.din(n10827), .dout(n11192));
  jand g10955(.dina(asqrt[23] ), .dinb(a[46] ), .dout(n11193));
  jor  g10956(.dina(n11193), .dinb(n10808), .dout(n11194));
  jor  g10957(.dina(n11194), .dinb(asqrt[24] ), .dout(n11195));
  jand g10958(.dina(asqrt[23] ), .dinb(n10134), .dout(n11196));
  jor  g10959(.dina(n11196), .dinb(n10135), .dout(n11197));
  jand g10960(.dina(n10838), .dinb(n11197), .dout(n11198));
  jand g10961(.dina(n11198), .dinb(n11195), .dout(n11199));
  jor  g10962(.dina(n11199), .dinb(n11192), .dout(n11200));
  jor  g10963(.dina(n11200), .dinb(asqrt[25] ), .dout(n11201));
  jnot g10964(.din(n10843), .dout(n11202));
  jand g10965(.dina(n11202), .dinb(n11201), .dout(n11203));
  jor  g10966(.dina(n11203), .dinb(n11191), .dout(n11204));
  jor  g10967(.dina(n11204), .dinb(asqrt[26] ), .dout(n11205));
  jnot g10968(.din(n10850), .dout(n11206));
  jand g10969(.dina(n11206), .dinb(n11205), .dout(n11207));
  jor  g10970(.dina(n11207), .dinb(n11190), .dout(n11208));
  jor  g10971(.dina(n11208), .dinb(asqrt[27] ), .dout(n11209));
  jnot g10972(.din(n10857), .dout(n11210));
  jand g10973(.dina(n11210), .dinb(n11209), .dout(n11211));
  jor  g10974(.dina(n11211), .dinb(n11189), .dout(n11212));
  jor  g10975(.dina(n11212), .dinb(asqrt[28] ), .dout(n11213));
  jand g10976(.dina(n10864), .dinb(n11213), .dout(n11214));
  jor  g10977(.dina(n11214), .dinb(n11188), .dout(n11215));
  jor  g10978(.dina(n11215), .dinb(asqrt[29] ), .dout(n11216));
  jnot g10979(.din(n10872), .dout(n11217));
  jand g10980(.dina(n11217), .dinb(n11216), .dout(n11218));
  jor  g10981(.dina(n11218), .dinb(n11187), .dout(n11219));
  jor  g10982(.dina(n11219), .dinb(asqrt[30] ), .dout(n11220));
  jand g10983(.dina(n10879), .dinb(n11220), .dout(n11221));
  jor  g10984(.dina(n11221), .dinb(n11186), .dout(n11222));
  jor  g10985(.dina(n11222), .dinb(asqrt[31] ), .dout(n11223));
  jnot g10986(.din(n10887), .dout(n11224));
  jand g10987(.dina(n11224), .dinb(n11223), .dout(n11225));
  jor  g10988(.dina(n11225), .dinb(n11185), .dout(n11226));
  jor  g10989(.dina(n11226), .dinb(asqrt[32] ), .dout(n11227));
  jnot g10990(.din(n10894), .dout(n11228));
  jand g10991(.dina(n11228), .dinb(n11227), .dout(n11229));
  jor  g10992(.dina(n11229), .dinb(n11184), .dout(n11230));
  jor  g10993(.dina(n11230), .dinb(asqrt[33] ), .dout(n11231));
  jnot g10994(.din(n10901), .dout(n11232));
  jand g10995(.dina(n11232), .dinb(n11231), .dout(n11233));
  jor  g10996(.dina(n11233), .dinb(n11183), .dout(n11234));
  jor  g10997(.dina(n11234), .dinb(asqrt[34] ), .dout(n11235));
  jand g10998(.dina(n10908), .dinb(n11235), .dout(n11236));
  jor  g10999(.dina(n11236), .dinb(n11182), .dout(n11237));
  jor  g11000(.dina(n11237), .dinb(asqrt[35] ), .dout(n11238));
  jnot g11001(.din(n10916), .dout(n11239));
  jand g11002(.dina(n11239), .dinb(n11238), .dout(n11240));
  jor  g11003(.dina(n11240), .dinb(n11181), .dout(n11241));
  jor  g11004(.dina(n11241), .dinb(asqrt[36] ), .dout(n11242));
  jnot g11005(.din(n10923), .dout(n11243));
  jand g11006(.dina(n11243), .dinb(n11242), .dout(n11244));
  jor  g11007(.dina(n11244), .dinb(n11180), .dout(n11245));
  jor  g11008(.dina(n11245), .dinb(asqrt[37] ), .dout(n11246));
  jnot g11009(.din(n10930), .dout(n11247));
  jand g11010(.dina(n11247), .dinb(n11246), .dout(n11248));
  jor  g11011(.dina(n11248), .dinb(n11179), .dout(n11249));
  jor  g11012(.dina(n11249), .dinb(asqrt[38] ), .dout(n11250));
  jnot g11013(.din(n10937), .dout(n11251));
  jand g11014(.dina(n11251), .dinb(n11250), .dout(n11252));
  jor  g11015(.dina(n11252), .dinb(n11178), .dout(n11253));
  jor  g11016(.dina(n11253), .dinb(asqrt[39] ), .dout(n11254));
  jnot g11017(.din(n10944), .dout(n11255));
  jand g11018(.dina(n11255), .dinb(n11254), .dout(n11256));
  jor  g11019(.dina(n11256), .dinb(n11177), .dout(n11257));
  jor  g11020(.dina(n11257), .dinb(asqrt[40] ), .dout(n11258));
  jand g11021(.dina(n11258), .dinb(n10950), .dout(n11259));
  jor  g11022(.dina(n11259), .dinb(n11176), .dout(n11260));
  jor  g11023(.dina(n11260), .dinb(asqrt[41] ), .dout(n11261));
  jnot g11024(.din(n10959), .dout(n11262));
  jand g11025(.dina(n11262), .dinb(n11261), .dout(n11263));
  jor  g11026(.dina(n11263), .dinb(n11175), .dout(n11264));
  jor  g11027(.dina(n11264), .dinb(asqrt[42] ), .dout(n11265));
  jand g11028(.dina(n10966), .dinb(n11265), .dout(n11266));
  jor  g11029(.dina(n11266), .dinb(n11174), .dout(n11267));
  jor  g11030(.dina(n11267), .dinb(asqrt[43] ), .dout(n11268));
  jnot g11031(.din(n10974), .dout(n11269));
  jand g11032(.dina(n11269), .dinb(n11268), .dout(n11270));
  jor  g11033(.dina(n11270), .dinb(n11173), .dout(n11271));
  jor  g11034(.dina(n11271), .dinb(asqrt[44] ), .dout(n11272));
  jand g11035(.dina(n10981), .dinb(n11272), .dout(n11273));
  jor  g11036(.dina(n11273), .dinb(n11172), .dout(n11274));
  jor  g11037(.dina(n11274), .dinb(asqrt[45] ), .dout(n11275));
  jnot g11038(.din(n10989), .dout(n11276));
  jand g11039(.dina(n11276), .dinb(n11275), .dout(n11277));
  jor  g11040(.dina(n11277), .dinb(n11171), .dout(n11278));
  jor  g11041(.dina(n11278), .dinb(asqrt[46] ), .dout(n11279));
  jnot g11042(.din(n10996), .dout(n11280));
  jand g11043(.dina(n11280), .dinb(n11279), .dout(n11281));
  jor  g11044(.dina(n11281), .dinb(n11170), .dout(n11282));
  jor  g11045(.dina(n11282), .dinb(asqrt[47] ), .dout(n11283));
  jnot g11046(.din(n11003), .dout(n11284));
  jand g11047(.dina(n11284), .dinb(n11283), .dout(n11285));
  jor  g11048(.dina(n11285), .dinb(n11169), .dout(n11286));
  jor  g11049(.dina(n11286), .dinb(asqrt[48] ), .dout(n11287));
  jand g11050(.dina(n11010), .dinb(n11287), .dout(n11288));
  jor  g11051(.dina(n11288), .dinb(n11168), .dout(n11289));
  jor  g11052(.dina(n11289), .dinb(asqrt[49] ), .dout(n11290));
  jnot g11053(.din(n11018), .dout(n11291));
  jand g11054(.dina(n11291), .dinb(n11290), .dout(n11292));
  jor  g11055(.dina(n11292), .dinb(n11167), .dout(n11293));
  jor  g11056(.dina(n11293), .dinb(asqrt[50] ), .dout(n11294));
  jand g11057(.dina(n11025), .dinb(n11294), .dout(n11295));
  jor  g11058(.dina(n11295), .dinb(n11166), .dout(n11296));
  jor  g11059(.dina(n11296), .dinb(asqrt[51] ), .dout(n11297));
  jnot g11060(.din(n11033), .dout(n11298));
  jand g11061(.dina(n11298), .dinb(n11297), .dout(n11299));
  jor  g11062(.dina(n11299), .dinb(n11165), .dout(n11300));
  jor  g11063(.dina(n11300), .dinb(asqrt[52] ), .dout(n11301));
  jand g11064(.dina(n11040), .dinb(n11301), .dout(n11302));
  jor  g11065(.dina(n11302), .dinb(n11164), .dout(n11303));
  jor  g11066(.dina(n11303), .dinb(asqrt[53] ), .dout(n11304));
  jnot g11067(.din(n11048), .dout(n11305));
  jand g11068(.dina(n11305), .dinb(n11304), .dout(n11306));
  jor  g11069(.dina(n11306), .dinb(n11163), .dout(n11307));
  jor  g11070(.dina(n11307), .dinb(asqrt[54] ), .dout(n11308));
  jand g11071(.dina(n11055), .dinb(n11308), .dout(n11309));
  jor  g11072(.dina(n11309), .dinb(n11162), .dout(n11310));
  jor  g11073(.dina(n11310), .dinb(asqrt[55] ), .dout(n11311));
  jand g11074(.dina(n11063), .dinb(n11311), .dout(n11312));
  jor  g11075(.dina(n11312), .dinb(n11161), .dout(n11313));
  jor  g11076(.dina(n11313), .dinb(asqrt[56] ), .dout(n11314));
  jand g11077(.dina(n11071), .dinb(n11314), .dout(n11315));
  jor  g11078(.dina(n11315), .dinb(n11160), .dout(n11316));
  jor  g11079(.dina(n11316), .dinb(asqrt[57] ), .dout(n11317));
  jnot g11080(.din(n11079), .dout(n11318));
  jand g11081(.dina(n11318), .dinb(n11317), .dout(n11319));
  jor  g11082(.dina(n11319), .dinb(n11159), .dout(n11320));
  jor  g11083(.dina(n11320), .dinb(asqrt[58] ), .dout(n11321));
  jnot g11084(.din(n11086), .dout(n11322));
  jand g11085(.dina(n11322), .dinb(n11321), .dout(n11323));
  jor  g11086(.dina(n11323), .dinb(n11158), .dout(n11324));
  jor  g11087(.dina(n11324), .dinb(asqrt[59] ), .dout(n11325));
  jnot g11088(.din(n11093), .dout(n11326));
  jand g11089(.dina(n11326), .dinb(n11325), .dout(n11327));
  jor  g11090(.dina(n11327), .dinb(n11157), .dout(n11328));
  jor  g11091(.dina(n11328), .dinb(asqrt[60] ), .dout(n11329));
  jand g11092(.dina(n11100), .dinb(n11329), .dout(n11330));
  jor  g11093(.dina(n11330), .dinb(n11156), .dout(n11331));
  jor  g11094(.dina(n11331), .dinb(asqrt[61] ), .dout(n11332));
  jnot g11095(.din(n11108), .dout(n11333));
  jand g11096(.dina(n11333), .dinb(n11332), .dout(n11334));
  jor  g11097(.dina(n11334), .dinb(n11155), .dout(n11335));
  jor  g11098(.dina(n11335), .dinb(asqrt[62] ), .dout(n11336));
  jand g11099(.dina(n11137), .dinb(n11336), .dout(n11337));
  jor  g11100(.dina(n11337), .dinb(n11154), .dout(n11338));
  jnot g11101(.din(n11120), .dout(n11339));
  jand g11102(.dina(n11339), .dinb(n11338), .dout(n11340));
  jand g11103(.dina(n11340), .dinb(n10820), .dout(n11341));
  jand g11104(.dina(n11341), .dinb(n11153), .dout(n11342));
  jor  g11105(.dina(n11342), .dinb(asqrt[63] ), .dout(n11343));
  jnot g11106(.din(n11133), .dout(n11344));
  jand g11107(.dina(n11344), .dinb(n11343), .dout(n11345));
  jand g11108(.dina(n11345), .dinb(n11126), .dout(n11346));
  jand g11109(.dina(n11346), .dinb(n11152), .dout(n11347));
  jor  g11110(.dina(n11347), .dinb(n11151), .dout(n11348));
  jand g11111(.dina(n11348), .dinb(n11150), .dout(n11349));
  jand g11112(.dina(n11349), .dinb(n11148), .dout(n11350));
  jor  g11113(.dina(n11350), .dinb(n11147), .dout(n11351));
  jand g11114(.dina(n11351), .dinb(asqrt[24] ), .dout(n11352));
  jor  g11115(.dina(n11351), .dinb(asqrt[24] ), .dout(n11353));
  jand g11116(.dina(asqrt[22] ), .dinb(n10807), .dout(n11354));
  jand g11117(.dina(n11152), .dinb(asqrt[23] ), .dout(n11355));
  jand g11118(.dina(n11355), .dinb(n11125), .dout(n11356));
  jand g11119(.dina(n11356), .dinb(n11343), .dout(n11357));
  jor  g11120(.dina(n11357), .dinb(n11354), .dout(n11358));
  jxor g11121(.dina(n11358), .dinb(a[46] ), .dout(n11359));
  jnot g11122(.din(n11359), .dout(n11360));
  jand g11123(.dina(n11360), .dinb(n11353), .dout(n11361));
  jor  g11124(.dina(n11361), .dinb(n11352), .dout(n11362));
  jand g11125(.dina(n11362), .dinb(asqrt[25] ), .dout(n11363));
  jor  g11126(.dina(n11362), .dinb(asqrt[25] ), .dout(n11364));
  jxor g11127(.dina(n10826), .dinb(n10328), .dout(n11365));
  jand g11128(.dina(n11365), .dinb(asqrt[22] ), .dout(n11366));
  jxor g11129(.dina(n11366), .dinb(n11198), .dout(n11367));
  jand g11130(.dina(n11367), .dinb(n11364), .dout(n11368));
  jor  g11131(.dina(n11368), .dinb(n11363), .dout(n11369));
  jand g11132(.dina(n11369), .dinb(asqrt[26] ), .dout(n11370));
  jor  g11133(.dina(n11369), .dinb(asqrt[26] ), .dout(n11371));
  jxor g11134(.dina(n10834), .dinb(n9832), .dout(n11372));
  jand g11135(.dina(n11372), .dinb(asqrt[22] ), .dout(n11373));
  jxor g11136(.dina(n11373), .dinb(n10843), .dout(n11374));
  jnot g11137(.din(n11374), .dout(n11375));
  jand g11138(.dina(n11375), .dinb(n11371), .dout(n11376));
  jor  g11139(.dina(n11376), .dinb(n11370), .dout(n11377));
  jand g11140(.dina(n11377), .dinb(asqrt[27] ), .dout(n11378));
  jor  g11141(.dina(n11377), .dinb(asqrt[27] ), .dout(n11379));
  jxor g11142(.dina(n10845), .dinb(n9369), .dout(n11380));
  jand g11143(.dina(n11380), .dinb(asqrt[22] ), .dout(n11381));
  jxor g11144(.dina(n11381), .dinb(n10850), .dout(n11382));
  jnot g11145(.din(n11382), .dout(n11383));
  jand g11146(.dina(n11383), .dinb(n11379), .dout(n11384));
  jor  g11147(.dina(n11384), .dinb(n11378), .dout(n11385));
  jand g11148(.dina(n11385), .dinb(asqrt[28] ), .dout(n11386));
  jor  g11149(.dina(n11385), .dinb(asqrt[28] ), .dout(n11387));
  jxor g11150(.dina(n10852), .dinb(n8890), .dout(n11388));
  jand g11151(.dina(n11388), .dinb(asqrt[22] ), .dout(n11389));
  jxor g11152(.dina(n11389), .dinb(n10857), .dout(n11390));
  jnot g11153(.din(n11390), .dout(n11391));
  jand g11154(.dina(n11391), .dinb(n11387), .dout(n11392));
  jor  g11155(.dina(n11392), .dinb(n11386), .dout(n11393));
  jand g11156(.dina(n11393), .dinb(asqrt[29] ), .dout(n11394));
  jor  g11157(.dina(n11393), .dinb(asqrt[29] ), .dout(n11395));
  jxor g11158(.dina(n10859), .dinb(n8449), .dout(n11396));
  jand g11159(.dina(n11396), .dinb(asqrt[22] ), .dout(n11397));
  jxor g11160(.dina(n11397), .dinb(n10864), .dout(n11398));
  jand g11161(.dina(n11398), .dinb(n11395), .dout(n11399));
  jor  g11162(.dina(n11399), .dinb(n11394), .dout(n11400));
  jand g11163(.dina(n11400), .dinb(asqrt[30] ), .dout(n11401));
  jor  g11164(.dina(n11400), .dinb(asqrt[30] ), .dout(n11402));
  jxor g11165(.dina(n10867), .dinb(n8003), .dout(n11403));
  jand g11166(.dina(n11403), .dinb(asqrt[22] ), .dout(n11404));
  jxor g11167(.dina(n11404), .dinb(n10872), .dout(n11405));
  jnot g11168(.din(n11405), .dout(n11406));
  jand g11169(.dina(n11406), .dinb(n11402), .dout(n11407));
  jor  g11170(.dina(n11407), .dinb(n11401), .dout(n11408));
  jand g11171(.dina(n11408), .dinb(asqrt[31] ), .dout(n11409));
  jor  g11172(.dina(n11408), .dinb(asqrt[31] ), .dout(n11410));
  jxor g11173(.dina(n10874), .dinb(n7581), .dout(n11411));
  jand g11174(.dina(n11411), .dinb(asqrt[22] ), .dout(n11412));
  jxor g11175(.dina(n11412), .dinb(n10879), .dout(n11413));
  jand g11176(.dina(n11413), .dinb(n11410), .dout(n11414));
  jor  g11177(.dina(n11414), .dinb(n11409), .dout(n11415));
  jand g11178(.dina(n11415), .dinb(asqrt[32] ), .dout(n11416));
  jor  g11179(.dina(n11415), .dinb(asqrt[32] ), .dout(n11417));
  jxor g11180(.dina(n10882), .dinb(n7154), .dout(n11418));
  jand g11181(.dina(n11418), .dinb(asqrt[22] ), .dout(n11419));
  jxor g11182(.dina(n11419), .dinb(n10887), .dout(n11420));
  jnot g11183(.din(n11420), .dout(n11421));
  jand g11184(.dina(n11421), .dinb(n11417), .dout(n11422));
  jor  g11185(.dina(n11422), .dinb(n11416), .dout(n11423));
  jand g11186(.dina(n11423), .dinb(asqrt[33] ), .dout(n11424));
  jor  g11187(.dina(n11423), .dinb(asqrt[33] ), .dout(n11425));
  jxor g11188(.dina(n10889), .dinb(n6758), .dout(n11426));
  jand g11189(.dina(n11426), .dinb(asqrt[22] ), .dout(n11427));
  jxor g11190(.dina(n11427), .dinb(n10894), .dout(n11428));
  jnot g11191(.din(n11428), .dout(n11429));
  jand g11192(.dina(n11429), .dinb(n11425), .dout(n11430));
  jor  g11193(.dina(n11430), .dinb(n11424), .dout(n11431));
  jand g11194(.dina(n11431), .dinb(asqrt[34] ), .dout(n11432));
  jor  g11195(.dina(n11431), .dinb(asqrt[34] ), .dout(n11433));
  jxor g11196(.dina(n10896), .dinb(n6357), .dout(n11434));
  jand g11197(.dina(n11434), .dinb(asqrt[22] ), .dout(n11435));
  jxor g11198(.dina(n11435), .dinb(n10901), .dout(n11436));
  jnot g11199(.din(n11436), .dout(n11437));
  jand g11200(.dina(n11437), .dinb(n11433), .dout(n11438));
  jor  g11201(.dina(n11438), .dinb(n11432), .dout(n11439));
  jand g11202(.dina(n11439), .dinb(asqrt[35] ), .dout(n11440));
  jor  g11203(.dina(n11439), .dinb(asqrt[35] ), .dout(n11441));
  jxor g11204(.dina(n10903), .dinb(n5989), .dout(n11442));
  jand g11205(.dina(n11442), .dinb(asqrt[22] ), .dout(n11443));
  jxor g11206(.dina(n11443), .dinb(n10908), .dout(n11444));
  jand g11207(.dina(n11444), .dinb(n11441), .dout(n11445));
  jor  g11208(.dina(n11445), .dinb(n11440), .dout(n11446));
  jand g11209(.dina(n11446), .dinb(asqrt[36] ), .dout(n11447));
  jor  g11210(.dina(n11446), .dinb(asqrt[36] ), .dout(n11448));
  jxor g11211(.dina(n10911), .dinb(n5606), .dout(n11449));
  jand g11212(.dina(n11449), .dinb(asqrt[22] ), .dout(n11450));
  jxor g11213(.dina(n11450), .dinb(n10916), .dout(n11451));
  jnot g11214(.din(n11451), .dout(n11452));
  jand g11215(.dina(n11452), .dinb(n11448), .dout(n11453));
  jor  g11216(.dina(n11453), .dinb(n11447), .dout(n11454));
  jand g11217(.dina(n11454), .dinb(asqrt[37] ), .dout(n11455));
  jor  g11218(.dina(n11454), .dinb(asqrt[37] ), .dout(n11456));
  jxor g11219(.dina(n10918), .dinb(n5259), .dout(n11457));
  jand g11220(.dina(n11457), .dinb(asqrt[22] ), .dout(n11458));
  jxor g11221(.dina(n11458), .dinb(n10923), .dout(n11459));
  jnot g11222(.din(n11459), .dout(n11460));
  jand g11223(.dina(n11460), .dinb(n11456), .dout(n11461));
  jor  g11224(.dina(n11461), .dinb(n11455), .dout(n11462));
  jand g11225(.dina(n11462), .dinb(asqrt[38] ), .dout(n11463));
  jor  g11226(.dina(n11462), .dinb(asqrt[38] ), .dout(n11464));
  jxor g11227(.dina(n10925), .dinb(n4902), .dout(n11465));
  jand g11228(.dina(n11465), .dinb(asqrt[22] ), .dout(n11466));
  jxor g11229(.dina(n11466), .dinb(n10930), .dout(n11467));
  jnot g11230(.din(n11467), .dout(n11468));
  jand g11231(.dina(n11468), .dinb(n11464), .dout(n11469));
  jor  g11232(.dina(n11469), .dinb(n11463), .dout(n11470));
  jand g11233(.dina(n11470), .dinb(asqrt[39] ), .dout(n11471));
  jor  g11234(.dina(n11470), .dinb(asqrt[39] ), .dout(n11472));
  jxor g11235(.dina(n10932), .dinb(n4582), .dout(n11473));
  jand g11236(.dina(n11473), .dinb(asqrt[22] ), .dout(n11474));
  jxor g11237(.dina(n11474), .dinb(n10937), .dout(n11475));
  jnot g11238(.din(n11475), .dout(n11476));
  jand g11239(.dina(n11476), .dinb(n11472), .dout(n11477));
  jor  g11240(.dina(n11477), .dinb(n11471), .dout(n11478));
  jand g11241(.dina(n11478), .dinb(asqrt[40] ), .dout(n11479));
  jor  g11242(.dina(n11478), .dinb(asqrt[40] ), .dout(n11480));
  jxor g11243(.dina(n10939), .dinb(n4249), .dout(n11481));
  jand g11244(.dina(n11481), .dinb(asqrt[22] ), .dout(n11482));
  jxor g11245(.dina(n11482), .dinb(n10944), .dout(n11483));
  jnot g11246(.din(n11483), .dout(n11484));
  jand g11247(.dina(n11484), .dinb(n11480), .dout(n11485));
  jor  g11248(.dina(n11485), .dinb(n11479), .dout(n11486));
  jand g11249(.dina(n11486), .dinb(asqrt[41] ), .dout(n11487));
  jxor g11250(.dina(n10946), .dinb(n3955), .dout(n11488));
  jand g11251(.dina(n11488), .dinb(asqrt[22] ), .dout(n11489));
  jxor g11252(.dina(n11489), .dinb(n10950), .dout(n11490));
  jor  g11253(.dina(n11486), .dinb(asqrt[41] ), .dout(n11491));
  jand g11254(.dina(n11491), .dinb(n11490), .dout(n11492));
  jor  g11255(.dina(n11492), .dinb(n11487), .dout(n11493));
  jand g11256(.dina(n11493), .dinb(asqrt[42] ), .dout(n11494));
  jor  g11257(.dina(n11493), .dinb(asqrt[42] ), .dout(n11495));
  jxor g11258(.dina(n10954), .dinb(n3642), .dout(n11496));
  jand g11259(.dina(n11496), .dinb(asqrt[22] ), .dout(n11497));
  jxor g11260(.dina(n11497), .dinb(n10959), .dout(n11498));
  jnot g11261(.din(n11498), .dout(n11499));
  jand g11262(.dina(n11499), .dinb(n11495), .dout(n11500));
  jor  g11263(.dina(n11500), .dinb(n11494), .dout(n11501));
  jand g11264(.dina(n11501), .dinb(asqrt[43] ), .dout(n11502));
  jor  g11265(.dina(n11501), .dinb(asqrt[43] ), .dout(n11503));
  jxor g11266(.dina(n10961), .dinb(n3368), .dout(n11504));
  jand g11267(.dina(n11504), .dinb(asqrt[22] ), .dout(n11505));
  jxor g11268(.dina(n11505), .dinb(n10966), .dout(n11506));
  jand g11269(.dina(n11506), .dinb(n11503), .dout(n11507));
  jor  g11270(.dina(n11507), .dinb(n11502), .dout(n11508));
  jand g11271(.dina(n11508), .dinb(asqrt[44] ), .dout(n11509));
  jor  g11272(.dina(n11508), .dinb(asqrt[44] ), .dout(n11510));
  jxor g11273(.dina(n10969), .dinb(n3089), .dout(n11511));
  jand g11274(.dina(n11511), .dinb(asqrt[22] ), .dout(n11512));
  jxor g11275(.dina(n11512), .dinb(n10974), .dout(n11513));
  jnot g11276(.din(n11513), .dout(n11514));
  jand g11277(.dina(n11514), .dinb(n11510), .dout(n11515));
  jor  g11278(.dina(n11515), .dinb(n11509), .dout(n11516));
  jand g11279(.dina(n11516), .dinb(asqrt[45] ), .dout(n11517));
  jor  g11280(.dina(n11516), .dinb(asqrt[45] ), .dout(n11518));
  jxor g11281(.dina(n10976), .dinb(n2833), .dout(n11519));
  jand g11282(.dina(n11519), .dinb(asqrt[22] ), .dout(n11520));
  jxor g11283(.dina(n11520), .dinb(n10981), .dout(n11521));
  jand g11284(.dina(n11521), .dinb(n11518), .dout(n11522));
  jor  g11285(.dina(n11522), .dinb(n11517), .dout(n11523));
  jand g11286(.dina(n11523), .dinb(asqrt[46] ), .dout(n11524));
  jor  g11287(.dina(n11523), .dinb(asqrt[46] ), .dout(n11525));
  jxor g11288(.dina(n10984), .dinb(n2572), .dout(n11526));
  jand g11289(.dina(n11526), .dinb(asqrt[22] ), .dout(n11527));
  jxor g11290(.dina(n11527), .dinb(n10989), .dout(n11528));
  jnot g11291(.din(n11528), .dout(n11529));
  jand g11292(.dina(n11529), .dinb(n11525), .dout(n11530));
  jor  g11293(.dina(n11530), .dinb(n11524), .dout(n11531));
  jand g11294(.dina(n11531), .dinb(asqrt[47] ), .dout(n11532));
  jor  g11295(.dina(n11531), .dinb(asqrt[47] ), .dout(n11533));
  jxor g11296(.dina(n10991), .dinb(n2345), .dout(n11534));
  jand g11297(.dina(n11534), .dinb(asqrt[22] ), .dout(n11535));
  jxor g11298(.dina(n11535), .dinb(n10996), .dout(n11536));
  jnot g11299(.din(n11536), .dout(n11537));
  jand g11300(.dina(n11537), .dinb(n11533), .dout(n11538));
  jor  g11301(.dina(n11538), .dinb(n11532), .dout(n11539));
  jand g11302(.dina(n11539), .dinb(asqrt[48] ), .dout(n11540));
  jor  g11303(.dina(n11539), .dinb(asqrt[48] ), .dout(n11541));
  jxor g11304(.dina(n10998), .dinb(n2108), .dout(n11542));
  jand g11305(.dina(n11542), .dinb(asqrt[22] ), .dout(n11543));
  jxor g11306(.dina(n11543), .dinb(n11003), .dout(n11544));
  jnot g11307(.din(n11544), .dout(n11545));
  jand g11308(.dina(n11545), .dinb(n11541), .dout(n11546));
  jor  g11309(.dina(n11546), .dinb(n11540), .dout(n11547));
  jand g11310(.dina(n11547), .dinb(asqrt[49] ), .dout(n11548));
  jor  g11311(.dina(n11547), .dinb(asqrt[49] ), .dout(n11549));
  jxor g11312(.dina(n11005), .dinb(n1912), .dout(n11550));
  jand g11313(.dina(n11550), .dinb(asqrt[22] ), .dout(n11551));
  jxor g11314(.dina(n11551), .dinb(n11010), .dout(n11552));
  jand g11315(.dina(n11552), .dinb(n11549), .dout(n11553));
  jor  g11316(.dina(n11553), .dinb(n11548), .dout(n11554));
  jand g11317(.dina(n11554), .dinb(asqrt[50] ), .dout(n11555));
  jor  g11318(.dina(n11554), .dinb(asqrt[50] ), .dout(n11556));
  jxor g11319(.dina(n11013), .dinb(n1699), .dout(n11557));
  jand g11320(.dina(n11557), .dinb(asqrt[22] ), .dout(n11558));
  jxor g11321(.dina(n11558), .dinb(n11018), .dout(n11559));
  jnot g11322(.din(n11559), .dout(n11560));
  jand g11323(.dina(n11560), .dinb(n11556), .dout(n11561));
  jor  g11324(.dina(n11561), .dinb(n11555), .dout(n11562));
  jand g11325(.dina(n11562), .dinb(asqrt[51] ), .dout(n11563));
  jor  g11326(.dina(n11562), .dinb(asqrt[51] ), .dout(n11564));
  jxor g11327(.dina(n11020), .dinb(n1516), .dout(n11565));
  jand g11328(.dina(n11565), .dinb(asqrt[22] ), .dout(n11566));
  jxor g11329(.dina(n11566), .dinb(n11025), .dout(n11567));
  jand g11330(.dina(n11567), .dinb(n11564), .dout(n11568));
  jor  g11331(.dina(n11568), .dinb(n11563), .dout(n11569));
  jand g11332(.dina(n11569), .dinb(asqrt[52] ), .dout(n11570));
  jor  g11333(.dina(n11569), .dinb(asqrt[52] ), .dout(n11571));
  jxor g11334(.dina(n11028), .dinb(n1332), .dout(n11572));
  jand g11335(.dina(n11572), .dinb(asqrt[22] ), .dout(n11573));
  jxor g11336(.dina(n11573), .dinb(n11033), .dout(n11574));
  jnot g11337(.din(n11574), .dout(n11575));
  jand g11338(.dina(n11575), .dinb(n11571), .dout(n11576));
  jor  g11339(.dina(n11576), .dinb(n11570), .dout(n11577));
  jand g11340(.dina(n11577), .dinb(asqrt[53] ), .dout(n11578));
  jor  g11341(.dina(n11577), .dinb(asqrt[53] ), .dout(n11579));
  jxor g11342(.dina(n11035), .dinb(n1173), .dout(n11580));
  jand g11343(.dina(n11580), .dinb(asqrt[22] ), .dout(n11581));
  jxor g11344(.dina(n11581), .dinb(n11040), .dout(n11582));
  jand g11345(.dina(n11582), .dinb(n11579), .dout(n11583));
  jor  g11346(.dina(n11583), .dinb(n11578), .dout(n11584));
  jand g11347(.dina(n11584), .dinb(asqrt[54] ), .dout(n11585));
  jor  g11348(.dina(n11584), .dinb(asqrt[54] ), .dout(n11586));
  jxor g11349(.dina(n11043), .dinb(n1008), .dout(n11587));
  jand g11350(.dina(n11587), .dinb(asqrt[22] ), .dout(n11588));
  jxor g11351(.dina(n11588), .dinb(n11048), .dout(n11589));
  jnot g11352(.din(n11589), .dout(n11590));
  jand g11353(.dina(n11590), .dinb(n11586), .dout(n11591));
  jor  g11354(.dina(n11591), .dinb(n11585), .dout(n11592));
  jand g11355(.dina(n11592), .dinb(asqrt[55] ), .dout(n11593));
  jor  g11356(.dina(n11592), .dinb(asqrt[55] ), .dout(n11594));
  jxor g11357(.dina(n11050), .dinb(n884), .dout(n11595));
  jand g11358(.dina(n11595), .dinb(asqrt[22] ), .dout(n11596));
  jxor g11359(.dina(n11596), .dinb(n11055), .dout(n11597));
  jand g11360(.dina(n11597), .dinb(n11594), .dout(n11598));
  jor  g11361(.dina(n11598), .dinb(n11593), .dout(n11599));
  jand g11362(.dina(n11599), .dinb(asqrt[56] ), .dout(n11600));
  jor  g11363(.dina(n11599), .dinb(asqrt[56] ), .dout(n11601));
  jxor g11364(.dina(n11058), .dinb(n743), .dout(n11602));
  jand g11365(.dina(n11602), .dinb(asqrt[22] ), .dout(n11603));
  jxor g11366(.dina(n11603), .dinb(n11063), .dout(n11604));
  jand g11367(.dina(n11604), .dinb(n11601), .dout(n11605));
  jor  g11368(.dina(n11605), .dinb(n11600), .dout(n11606));
  jand g11369(.dina(n11606), .dinb(asqrt[57] ), .dout(n11607));
  jor  g11370(.dina(n11606), .dinb(asqrt[57] ), .dout(n11608));
  jxor g11371(.dina(n11066), .dinb(n635), .dout(n11609));
  jand g11372(.dina(n11609), .dinb(asqrt[22] ), .dout(n11610));
  jxor g11373(.dina(n11610), .dinb(n11071), .dout(n11611));
  jand g11374(.dina(n11611), .dinb(n11608), .dout(n11612));
  jor  g11375(.dina(n11612), .dinb(n11607), .dout(n11613));
  jand g11376(.dina(n11613), .dinb(asqrt[58] ), .dout(n11614));
  jor  g11377(.dina(n11613), .dinb(asqrt[58] ), .dout(n11615));
  jxor g11378(.dina(n11074), .dinb(n515), .dout(n11616));
  jand g11379(.dina(n11616), .dinb(asqrt[22] ), .dout(n11617));
  jxor g11380(.dina(n11617), .dinb(n11079), .dout(n11618));
  jnot g11381(.din(n11618), .dout(n11619));
  jand g11382(.dina(n11619), .dinb(n11615), .dout(n11620));
  jor  g11383(.dina(n11620), .dinb(n11614), .dout(n11621));
  jand g11384(.dina(n11621), .dinb(asqrt[59] ), .dout(n11622));
  jor  g11385(.dina(n11621), .dinb(asqrt[59] ), .dout(n11623));
  jxor g11386(.dina(n11081), .dinb(n443), .dout(n11624));
  jand g11387(.dina(n11624), .dinb(asqrt[22] ), .dout(n11625));
  jxor g11388(.dina(n11625), .dinb(n11086), .dout(n11626));
  jnot g11389(.din(n11626), .dout(n11627));
  jand g11390(.dina(n11627), .dinb(n11623), .dout(n11628));
  jor  g11391(.dina(n11628), .dinb(n11622), .dout(n11629));
  jand g11392(.dina(n11629), .dinb(asqrt[60] ), .dout(n11630));
  jor  g11393(.dina(n11629), .dinb(asqrt[60] ), .dout(n11631));
  jxor g11394(.dina(n11088), .dinb(n352), .dout(n11632));
  jand g11395(.dina(n11632), .dinb(asqrt[22] ), .dout(n11633));
  jxor g11396(.dina(n11633), .dinb(n11093), .dout(n11634));
  jnot g11397(.din(n11634), .dout(n11635));
  jand g11398(.dina(n11635), .dinb(n11631), .dout(n11636));
  jor  g11399(.dina(n11636), .dinb(n11630), .dout(n11637));
  jand g11400(.dina(n11637), .dinb(asqrt[61] ), .dout(n11638));
  jor  g11401(.dina(n11637), .dinb(asqrt[61] ), .dout(n11639));
  jxor g11402(.dina(n11095), .dinb(n294), .dout(n11640));
  jand g11403(.dina(n11640), .dinb(asqrt[22] ), .dout(n11641));
  jxor g11404(.dina(n11641), .dinb(n11100), .dout(n11642));
  jand g11405(.dina(n11642), .dinb(n11639), .dout(n11643));
  jor  g11406(.dina(n11643), .dinb(n11638), .dout(n11644));
  jand g11407(.dina(n11644), .dinb(asqrt[62] ), .dout(n11645));
  jor  g11408(.dina(n11644), .dinb(asqrt[62] ), .dout(n11646));
  jxor g11409(.dina(n11103), .dinb(n239), .dout(n11647));
  jand g11410(.dina(n11647), .dinb(asqrt[22] ), .dout(n11648));
  jxor g11411(.dina(n11648), .dinb(n11108), .dout(n11649));
  jnot g11412(.din(n11649), .dout(n11650));
  jand g11413(.dina(n11650), .dinb(n11646), .dout(n11651));
  jor  g11414(.dina(n11651), .dinb(n11645), .dout(n11652));
  jor  g11415(.dina(n11652), .dinb(n11140), .dout(n11653));
  jnot g11416(.din(n11653), .dout(n11654));
  jnot g11417(.din(n11140), .dout(n11656));
  jnot g11418(.din(n11645), .dout(n11657));
  jnot g11419(.din(n11638), .dout(n11658));
  jnot g11420(.din(n11630), .dout(n11659));
  jnot g11421(.din(n11622), .dout(n11660));
  jnot g11422(.din(n11614), .dout(n11661));
  jnot g11423(.din(n11607), .dout(n11662));
  jnot g11424(.din(n11600), .dout(n11663));
  jnot g11425(.din(n11593), .dout(n11664));
  jnot g11426(.din(n11585), .dout(n11665));
  jnot g11427(.din(n11578), .dout(n11666));
  jnot g11428(.din(n11570), .dout(n11667));
  jnot g11429(.din(n11563), .dout(n11668));
  jnot g11430(.din(n11555), .dout(n11669));
  jnot g11431(.din(n11548), .dout(n11670));
  jnot g11432(.din(n11540), .dout(n11671));
  jnot g11433(.din(n11532), .dout(n11672));
  jnot g11434(.din(n11524), .dout(n11673));
  jnot g11435(.din(n11517), .dout(n11674));
  jnot g11436(.din(n11509), .dout(n11675));
  jnot g11437(.din(n11502), .dout(n11676));
  jnot g11438(.din(n11494), .dout(n11677));
  jnot g11439(.din(n11487), .dout(n11678));
  jnot g11440(.din(n11490), .dout(n11679));
  jnot g11441(.din(n11479), .dout(n11680));
  jnot g11442(.din(n11471), .dout(n11681));
  jnot g11443(.din(n11463), .dout(n11682));
  jnot g11444(.din(n11455), .dout(n11683));
  jnot g11445(.din(n11447), .dout(n11684));
  jnot g11446(.din(n11440), .dout(n11685));
  jnot g11447(.din(n11432), .dout(n11686));
  jnot g11448(.din(n11424), .dout(n11687));
  jnot g11449(.din(n11416), .dout(n11688));
  jnot g11450(.din(n11409), .dout(n11689));
  jnot g11451(.din(n11401), .dout(n11690));
  jnot g11452(.din(n11394), .dout(n11691));
  jnot g11453(.din(n11386), .dout(n11692));
  jnot g11454(.din(n11378), .dout(n11693));
  jnot g11455(.din(n11370), .dout(n11694));
  jnot g11456(.din(n11363), .dout(n11695));
  jnot g11457(.din(n11352), .dout(n11696));
  jnot g11458(.din(n11147), .dout(n11697));
  jor  g11459(.dina(n11347), .dinb(n10805), .dout(n11698));
  jnot g11460(.din(n11145), .dout(n11699));
  jand g11461(.dina(n11699), .dinb(n11698), .dout(n11700));
  jand g11462(.dina(n11700), .dinb(n10824), .dout(n11701));
  jor  g11463(.dina(n11347), .dinb(a[44] ), .dout(n11702));
  jand g11464(.dina(n11702), .dinb(a[45] ), .dout(n11703));
  jor  g11465(.dina(n11354), .dinb(n11703), .dout(n11704));
  jor  g11466(.dina(n11704), .dinb(n11701), .dout(n11705));
  jand g11467(.dina(n11705), .dinb(n11697), .dout(n11706));
  jand g11468(.dina(n11706), .dinb(n10328), .dout(n11707));
  jor  g11469(.dina(n11359), .dinb(n11707), .dout(n11708));
  jand g11470(.dina(n11708), .dinb(n11696), .dout(n11709));
  jand g11471(.dina(n11709), .dinb(n9832), .dout(n11710));
  jnot g11472(.din(n11367), .dout(n11711));
  jor  g11473(.dina(n11711), .dinb(n11710), .dout(n11712));
  jand g11474(.dina(n11712), .dinb(n11695), .dout(n11713));
  jand g11475(.dina(n11713), .dinb(n9369), .dout(n11714));
  jor  g11476(.dina(n11374), .dinb(n11714), .dout(n11715));
  jand g11477(.dina(n11715), .dinb(n11694), .dout(n11716));
  jand g11478(.dina(n11716), .dinb(n8890), .dout(n11717));
  jor  g11479(.dina(n11382), .dinb(n11717), .dout(n11718));
  jand g11480(.dina(n11718), .dinb(n11693), .dout(n11719));
  jand g11481(.dina(n11719), .dinb(n8449), .dout(n11720));
  jor  g11482(.dina(n11390), .dinb(n11720), .dout(n11721));
  jand g11483(.dina(n11721), .dinb(n11692), .dout(n11722));
  jand g11484(.dina(n11722), .dinb(n8003), .dout(n11723));
  jnot g11485(.din(n11398), .dout(n11724));
  jor  g11486(.dina(n11724), .dinb(n11723), .dout(n11725));
  jand g11487(.dina(n11725), .dinb(n11691), .dout(n11726));
  jand g11488(.dina(n11726), .dinb(n7581), .dout(n11727));
  jor  g11489(.dina(n11405), .dinb(n11727), .dout(n11728));
  jand g11490(.dina(n11728), .dinb(n11690), .dout(n11729));
  jand g11491(.dina(n11729), .dinb(n7154), .dout(n11730));
  jnot g11492(.din(n11413), .dout(n11731));
  jor  g11493(.dina(n11731), .dinb(n11730), .dout(n11732));
  jand g11494(.dina(n11732), .dinb(n11689), .dout(n11733));
  jand g11495(.dina(n11733), .dinb(n6758), .dout(n11734));
  jor  g11496(.dina(n11420), .dinb(n11734), .dout(n11735));
  jand g11497(.dina(n11735), .dinb(n11688), .dout(n11736));
  jand g11498(.dina(n11736), .dinb(n6357), .dout(n11737));
  jor  g11499(.dina(n11428), .dinb(n11737), .dout(n11738));
  jand g11500(.dina(n11738), .dinb(n11687), .dout(n11739));
  jand g11501(.dina(n11739), .dinb(n5989), .dout(n11740));
  jor  g11502(.dina(n11436), .dinb(n11740), .dout(n11741));
  jand g11503(.dina(n11741), .dinb(n11686), .dout(n11742));
  jand g11504(.dina(n11742), .dinb(n5606), .dout(n11743));
  jnot g11505(.din(n11444), .dout(n11744));
  jor  g11506(.dina(n11744), .dinb(n11743), .dout(n11745));
  jand g11507(.dina(n11745), .dinb(n11685), .dout(n11746));
  jand g11508(.dina(n11746), .dinb(n5259), .dout(n11747));
  jor  g11509(.dina(n11451), .dinb(n11747), .dout(n11748));
  jand g11510(.dina(n11748), .dinb(n11684), .dout(n11749));
  jand g11511(.dina(n11749), .dinb(n4902), .dout(n11750));
  jor  g11512(.dina(n11459), .dinb(n11750), .dout(n11751));
  jand g11513(.dina(n11751), .dinb(n11683), .dout(n11752));
  jand g11514(.dina(n11752), .dinb(n4582), .dout(n11753));
  jor  g11515(.dina(n11467), .dinb(n11753), .dout(n11754));
  jand g11516(.dina(n11754), .dinb(n11682), .dout(n11755));
  jand g11517(.dina(n11755), .dinb(n4249), .dout(n11756));
  jor  g11518(.dina(n11475), .dinb(n11756), .dout(n11757));
  jand g11519(.dina(n11757), .dinb(n11681), .dout(n11758));
  jand g11520(.dina(n11758), .dinb(n3955), .dout(n11759));
  jor  g11521(.dina(n11483), .dinb(n11759), .dout(n11760));
  jand g11522(.dina(n11760), .dinb(n11680), .dout(n11761));
  jand g11523(.dina(n11761), .dinb(n3642), .dout(n11762));
  jor  g11524(.dina(n11762), .dinb(n11679), .dout(n11763));
  jand g11525(.dina(n11763), .dinb(n11678), .dout(n11764));
  jand g11526(.dina(n11764), .dinb(n3368), .dout(n11765));
  jor  g11527(.dina(n11498), .dinb(n11765), .dout(n11766));
  jand g11528(.dina(n11766), .dinb(n11677), .dout(n11767));
  jand g11529(.dina(n11767), .dinb(n3089), .dout(n11768));
  jnot g11530(.din(n11506), .dout(n11769));
  jor  g11531(.dina(n11769), .dinb(n11768), .dout(n11770));
  jand g11532(.dina(n11770), .dinb(n11676), .dout(n11771));
  jand g11533(.dina(n11771), .dinb(n2833), .dout(n11772));
  jor  g11534(.dina(n11513), .dinb(n11772), .dout(n11773));
  jand g11535(.dina(n11773), .dinb(n11675), .dout(n11774));
  jand g11536(.dina(n11774), .dinb(n2572), .dout(n11775));
  jnot g11537(.din(n11521), .dout(n11776));
  jor  g11538(.dina(n11776), .dinb(n11775), .dout(n11777));
  jand g11539(.dina(n11777), .dinb(n11674), .dout(n11778));
  jand g11540(.dina(n11778), .dinb(n2345), .dout(n11779));
  jor  g11541(.dina(n11528), .dinb(n11779), .dout(n11780));
  jand g11542(.dina(n11780), .dinb(n11673), .dout(n11781));
  jand g11543(.dina(n11781), .dinb(n2108), .dout(n11782));
  jor  g11544(.dina(n11536), .dinb(n11782), .dout(n11783));
  jand g11545(.dina(n11783), .dinb(n11672), .dout(n11784));
  jand g11546(.dina(n11784), .dinb(n1912), .dout(n11785));
  jor  g11547(.dina(n11544), .dinb(n11785), .dout(n11786));
  jand g11548(.dina(n11786), .dinb(n11671), .dout(n11787));
  jand g11549(.dina(n11787), .dinb(n1699), .dout(n11788));
  jnot g11550(.din(n11552), .dout(n11789));
  jor  g11551(.dina(n11789), .dinb(n11788), .dout(n11790));
  jand g11552(.dina(n11790), .dinb(n11670), .dout(n11791));
  jand g11553(.dina(n11791), .dinb(n1516), .dout(n11792));
  jor  g11554(.dina(n11559), .dinb(n11792), .dout(n11793));
  jand g11555(.dina(n11793), .dinb(n11669), .dout(n11794));
  jand g11556(.dina(n11794), .dinb(n1332), .dout(n11795));
  jnot g11557(.din(n11567), .dout(n11796));
  jor  g11558(.dina(n11796), .dinb(n11795), .dout(n11797));
  jand g11559(.dina(n11797), .dinb(n11668), .dout(n11798));
  jand g11560(.dina(n11798), .dinb(n1173), .dout(n11799));
  jor  g11561(.dina(n11574), .dinb(n11799), .dout(n11800));
  jand g11562(.dina(n11800), .dinb(n11667), .dout(n11801));
  jand g11563(.dina(n11801), .dinb(n1008), .dout(n11802));
  jnot g11564(.din(n11582), .dout(n11803));
  jor  g11565(.dina(n11803), .dinb(n11802), .dout(n11804));
  jand g11566(.dina(n11804), .dinb(n11666), .dout(n11805));
  jand g11567(.dina(n11805), .dinb(n884), .dout(n11806));
  jor  g11568(.dina(n11589), .dinb(n11806), .dout(n11807));
  jand g11569(.dina(n11807), .dinb(n11665), .dout(n11808));
  jand g11570(.dina(n11808), .dinb(n743), .dout(n11809));
  jnot g11571(.din(n11597), .dout(n11810));
  jor  g11572(.dina(n11810), .dinb(n11809), .dout(n11811));
  jand g11573(.dina(n11811), .dinb(n11664), .dout(n11812));
  jand g11574(.dina(n11812), .dinb(n635), .dout(n11813));
  jnot g11575(.din(n11604), .dout(n11814));
  jor  g11576(.dina(n11814), .dinb(n11813), .dout(n11815));
  jand g11577(.dina(n11815), .dinb(n11663), .dout(n11816));
  jand g11578(.dina(n11816), .dinb(n515), .dout(n11817));
  jnot g11579(.din(n11611), .dout(n11818));
  jor  g11580(.dina(n11818), .dinb(n11817), .dout(n11819));
  jand g11581(.dina(n11819), .dinb(n11662), .dout(n11820));
  jand g11582(.dina(n11820), .dinb(n443), .dout(n11821));
  jor  g11583(.dina(n11618), .dinb(n11821), .dout(n11822));
  jand g11584(.dina(n11822), .dinb(n11661), .dout(n11823));
  jand g11585(.dina(n11823), .dinb(n352), .dout(n11824));
  jor  g11586(.dina(n11626), .dinb(n11824), .dout(n11825));
  jand g11587(.dina(n11825), .dinb(n11660), .dout(n11826));
  jand g11588(.dina(n11826), .dinb(n294), .dout(n11827));
  jor  g11589(.dina(n11634), .dinb(n11827), .dout(n11828));
  jand g11590(.dina(n11828), .dinb(n11659), .dout(n11829));
  jand g11591(.dina(n11829), .dinb(n239), .dout(n11830));
  jnot g11592(.din(n11642), .dout(n11831));
  jor  g11593(.dina(n11831), .dinb(n11830), .dout(n11832));
  jand g11594(.dina(n11832), .dinb(n11658), .dout(n11833));
  jand g11595(.dina(n11833), .dinb(n221), .dout(n11834));
  jor  g11596(.dina(n11649), .dinb(n11834), .dout(n11835));
  jand g11597(.dina(n11835), .dinb(n11657), .dout(n11836));
  jor  g11598(.dina(n11836), .dinb(n11656), .dout(n11837));
  jxor g11599(.dina(n11120), .dinb(n11117), .dout(n11838));
  jnot g11600(.din(n11838), .dout(n11839));
  jand g11601(.dina(n11839), .dinb(asqrt[22] ), .dout(n11840));
  jor  g11602(.dina(n11840), .dinb(n11837), .dout(n11841));
  jand g11603(.dina(n11841), .dinb(n218), .dout(n11842));
  jand g11604(.dina(n11346), .dinb(n11117), .dout(n11843));
  jnot g11605(.din(n11843), .dout(n11844));
  jand g11606(.dina(n11838), .dinb(asqrt[63] ), .dout(n11845));
  jand g11607(.dina(n11845), .dinb(n11844), .dout(n11846));
  jor  g11608(.dina(n11846), .dinb(n11842), .dout(n11847));
  jor  g11609(.dina(n11847), .dinb(n11654), .dout(asqrt[21] ));
  jand g11610(.dina(n11652), .dinb(n11140), .dout(n11851));
  jnot g11611(.din(n11840), .dout(n11852));
  jand g11612(.dina(n11852), .dinb(n11851), .dout(n11853));
  jor  g11613(.dina(n11853), .dinb(asqrt[63] ), .dout(n11854));
  jnot g11614(.din(n11846), .dout(n11855));
  jand g11615(.dina(n11855), .dinb(n11854), .dout(n11856));
  jand g11616(.dina(n11856), .dinb(n11653), .dout(n11858));
  jxor g11617(.dina(n11644), .dinb(n221), .dout(n11859));
  jor  g11618(.dina(n11859), .dinb(n11858), .dout(n11860));
  jxor g11619(.dina(n11860), .dinb(n11649), .dout(n11861));
  jnot g11620(.din(n11861), .dout(n11862));
  jor  g11621(.dina(n11858), .dinb(n11142), .dout(n11863));
  jnot g11622(.din(a[40] ), .dout(n11864));
  jnot g11623(.din(a[41] ), .dout(n11865));
  jand g11624(.dina(n11865), .dinb(n11864), .dout(n11866));
  jand g11625(.dina(n11866), .dinb(n11142), .dout(n11867));
  jnot g11626(.din(n11867), .dout(n11868));
  jand g11627(.dina(n11868), .dinb(n11863), .dout(n11869));
  jor  g11628(.dina(n11869), .dinb(n11347), .dout(n11870));
  jand g11629(.dina(n11869), .dinb(n11347), .dout(n11871));
  jor  g11630(.dina(n11858), .dinb(a[42] ), .dout(n11872));
  jand g11631(.dina(n11872), .dinb(a[43] ), .dout(n11873));
  jand g11632(.dina(asqrt[21] ), .dinb(n11144), .dout(n11874));
  jor  g11633(.dina(n11874), .dinb(n11873), .dout(n11875));
  jor  g11634(.dina(n11875), .dinb(n11871), .dout(n11876));
  jand g11635(.dina(n11876), .dinb(n11870), .dout(n11877));
  jor  g11636(.dina(n11877), .dinb(n10824), .dout(n11878));
  jand g11637(.dina(n11877), .dinb(n10824), .dout(n11879));
  jnot g11638(.din(n11144), .dout(n11880));
  jor  g11639(.dina(n11858), .dinb(n11880), .dout(n11881));
  jor  g11640(.dina(n11845), .dinb(n11654), .dout(n11882));
  jor  g11641(.dina(n11882), .dinb(n11842), .dout(n11883));
  jor  g11642(.dina(n11883), .dinb(n11347), .dout(n11884));
  jand g11643(.dina(n11884), .dinb(n11881), .dout(n11885));
  jxor g11644(.dina(n11885), .dinb(n10805), .dout(n11886));
  jor  g11645(.dina(n11886), .dinb(n11879), .dout(n11887));
  jand g11646(.dina(n11887), .dinb(n11878), .dout(n11888));
  jor  g11647(.dina(n11888), .dinb(n10328), .dout(n11889));
  jand g11648(.dina(n11888), .dinb(n10328), .dout(n11890));
  jxor g11649(.dina(n11146), .dinb(n10824), .dout(n11891));
  jor  g11650(.dina(n11891), .dinb(n11858), .dout(n11892));
  jxor g11651(.dina(n11892), .dinb(n11704), .dout(n11893));
  jnot g11652(.din(n11893), .dout(n11894));
  jor  g11653(.dina(n11894), .dinb(n11890), .dout(n11895));
  jand g11654(.dina(n11895), .dinb(n11889), .dout(n11896));
  jor  g11655(.dina(n11896), .dinb(n9832), .dout(n11897));
  jand g11656(.dina(n11896), .dinb(n9832), .dout(n11898));
  jxor g11657(.dina(n11351), .dinb(n10328), .dout(n11899));
  jor  g11658(.dina(n11899), .dinb(n11858), .dout(n11900));
  jxor g11659(.dina(n11900), .dinb(n11360), .dout(n11901));
  jor  g11660(.dina(n11901), .dinb(n11898), .dout(n11902));
  jand g11661(.dina(n11902), .dinb(n11897), .dout(n11903));
  jor  g11662(.dina(n11903), .dinb(n9369), .dout(n11904));
  jand g11663(.dina(n11903), .dinb(n9369), .dout(n11905));
  jxor g11664(.dina(n11362), .dinb(n9832), .dout(n11906));
  jor  g11665(.dina(n11906), .dinb(n11858), .dout(n11907));
  jxor g11666(.dina(n11907), .dinb(n11711), .dout(n11908));
  jnot g11667(.din(n11908), .dout(n11909));
  jor  g11668(.dina(n11909), .dinb(n11905), .dout(n11910));
  jand g11669(.dina(n11910), .dinb(n11904), .dout(n11911));
  jor  g11670(.dina(n11911), .dinb(n8890), .dout(n11912));
  jand g11671(.dina(n11911), .dinb(n8890), .dout(n11913));
  jxor g11672(.dina(n11369), .dinb(n9369), .dout(n11914));
  jor  g11673(.dina(n11914), .dinb(n11858), .dout(n11915));
  jxor g11674(.dina(n11915), .dinb(n11375), .dout(n11916));
  jor  g11675(.dina(n11916), .dinb(n11913), .dout(n11917));
  jand g11676(.dina(n11917), .dinb(n11912), .dout(n11918));
  jor  g11677(.dina(n11918), .dinb(n8449), .dout(n11919));
  jand g11678(.dina(n11918), .dinb(n8449), .dout(n11920));
  jxor g11679(.dina(n11377), .dinb(n8890), .dout(n11921));
  jor  g11680(.dina(n11921), .dinb(n11858), .dout(n11922));
  jxor g11681(.dina(n11922), .dinb(n11383), .dout(n11923));
  jor  g11682(.dina(n11923), .dinb(n11920), .dout(n11924));
  jand g11683(.dina(n11924), .dinb(n11919), .dout(n11925));
  jor  g11684(.dina(n11925), .dinb(n8003), .dout(n11926));
  jand g11685(.dina(n11925), .dinb(n8003), .dout(n11927));
  jxor g11686(.dina(n11385), .dinb(n8449), .dout(n11928));
  jor  g11687(.dina(n11928), .dinb(n11858), .dout(n11929));
  jxor g11688(.dina(n11929), .dinb(n11391), .dout(n11930));
  jor  g11689(.dina(n11930), .dinb(n11927), .dout(n11931));
  jand g11690(.dina(n11931), .dinb(n11926), .dout(n11932));
  jor  g11691(.dina(n11932), .dinb(n7581), .dout(n11933));
  jand g11692(.dina(n11932), .dinb(n7581), .dout(n11934));
  jxor g11693(.dina(n11393), .dinb(n8003), .dout(n11935));
  jor  g11694(.dina(n11935), .dinb(n11858), .dout(n11936));
  jxor g11695(.dina(n11936), .dinb(n11724), .dout(n11937));
  jnot g11696(.din(n11937), .dout(n11938));
  jor  g11697(.dina(n11938), .dinb(n11934), .dout(n11939));
  jand g11698(.dina(n11939), .dinb(n11933), .dout(n11940));
  jor  g11699(.dina(n11940), .dinb(n7154), .dout(n11941));
  jand g11700(.dina(n11940), .dinb(n7154), .dout(n11942));
  jxor g11701(.dina(n11400), .dinb(n7581), .dout(n11943));
  jor  g11702(.dina(n11943), .dinb(n11858), .dout(n11944));
  jxor g11703(.dina(n11944), .dinb(n11406), .dout(n11945));
  jor  g11704(.dina(n11945), .dinb(n11942), .dout(n11946));
  jand g11705(.dina(n11946), .dinb(n11941), .dout(n11947));
  jor  g11706(.dina(n11947), .dinb(n6758), .dout(n11948));
  jand g11707(.dina(n11947), .dinb(n6758), .dout(n11949));
  jxor g11708(.dina(n11408), .dinb(n7154), .dout(n11950));
  jor  g11709(.dina(n11950), .dinb(n11858), .dout(n11951));
  jxor g11710(.dina(n11951), .dinb(n11731), .dout(n11952));
  jnot g11711(.din(n11952), .dout(n11953));
  jor  g11712(.dina(n11953), .dinb(n11949), .dout(n11954));
  jand g11713(.dina(n11954), .dinb(n11948), .dout(n11955));
  jor  g11714(.dina(n11955), .dinb(n6357), .dout(n11956));
  jand g11715(.dina(n11955), .dinb(n6357), .dout(n11957));
  jxor g11716(.dina(n11415), .dinb(n6758), .dout(n11958));
  jor  g11717(.dina(n11958), .dinb(n11858), .dout(n11959));
  jxor g11718(.dina(n11959), .dinb(n11421), .dout(n11960));
  jor  g11719(.dina(n11960), .dinb(n11957), .dout(n11961));
  jand g11720(.dina(n11961), .dinb(n11956), .dout(n11962));
  jor  g11721(.dina(n11962), .dinb(n5989), .dout(n11963));
  jand g11722(.dina(n11962), .dinb(n5989), .dout(n11964));
  jxor g11723(.dina(n11423), .dinb(n6357), .dout(n11965));
  jor  g11724(.dina(n11965), .dinb(n11858), .dout(n11966));
  jxor g11725(.dina(n11966), .dinb(n11429), .dout(n11967));
  jor  g11726(.dina(n11967), .dinb(n11964), .dout(n11968));
  jand g11727(.dina(n11968), .dinb(n11963), .dout(n11969));
  jor  g11728(.dina(n11969), .dinb(n5606), .dout(n11970));
  jand g11729(.dina(n11969), .dinb(n5606), .dout(n11971));
  jxor g11730(.dina(n11431), .dinb(n5989), .dout(n11972));
  jor  g11731(.dina(n11972), .dinb(n11858), .dout(n11973));
  jxor g11732(.dina(n11973), .dinb(n11437), .dout(n11974));
  jor  g11733(.dina(n11974), .dinb(n11971), .dout(n11975));
  jand g11734(.dina(n11975), .dinb(n11970), .dout(n11976));
  jor  g11735(.dina(n11976), .dinb(n5259), .dout(n11977));
  jand g11736(.dina(n11976), .dinb(n5259), .dout(n11978));
  jxor g11737(.dina(n11439), .dinb(n5606), .dout(n11979));
  jor  g11738(.dina(n11979), .dinb(n11858), .dout(n11980));
  jxor g11739(.dina(n11980), .dinb(n11744), .dout(n11981));
  jnot g11740(.din(n11981), .dout(n11982));
  jor  g11741(.dina(n11982), .dinb(n11978), .dout(n11983));
  jand g11742(.dina(n11983), .dinb(n11977), .dout(n11984));
  jor  g11743(.dina(n11984), .dinb(n4902), .dout(n11985));
  jand g11744(.dina(n11984), .dinb(n4902), .dout(n11986));
  jxor g11745(.dina(n11446), .dinb(n5259), .dout(n11987));
  jor  g11746(.dina(n11987), .dinb(n11858), .dout(n11988));
  jxor g11747(.dina(n11988), .dinb(n11452), .dout(n11989));
  jor  g11748(.dina(n11989), .dinb(n11986), .dout(n11990));
  jand g11749(.dina(n11990), .dinb(n11985), .dout(n11991));
  jor  g11750(.dina(n11991), .dinb(n4582), .dout(n11992));
  jand g11751(.dina(n11991), .dinb(n4582), .dout(n11993));
  jxor g11752(.dina(n11454), .dinb(n4902), .dout(n11994));
  jor  g11753(.dina(n11994), .dinb(n11858), .dout(n11995));
  jxor g11754(.dina(n11995), .dinb(n11460), .dout(n11996));
  jor  g11755(.dina(n11996), .dinb(n11993), .dout(n11997));
  jand g11756(.dina(n11997), .dinb(n11992), .dout(n11998));
  jor  g11757(.dina(n11998), .dinb(n4249), .dout(n11999));
  jand g11758(.dina(n11998), .dinb(n4249), .dout(n12000));
  jxor g11759(.dina(n11462), .dinb(n4582), .dout(n12001));
  jor  g11760(.dina(n12001), .dinb(n11858), .dout(n12002));
  jxor g11761(.dina(n12002), .dinb(n11468), .dout(n12003));
  jor  g11762(.dina(n12003), .dinb(n12000), .dout(n12004));
  jand g11763(.dina(n12004), .dinb(n11999), .dout(n12005));
  jor  g11764(.dina(n12005), .dinb(n3955), .dout(n12006));
  jand g11765(.dina(n12005), .dinb(n3955), .dout(n12007));
  jxor g11766(.dina(n11470), .dinb(n4249), .dout(n12008));
  jor  g11767(.dina(n12008), .dinb(n11858), .dout(n12009));
  jxor g11768(.dina(n12009), .dinb(n11476), .dout(n12010));
  jor  g11769(.dina(n12010), .dinb(n12007), .dout(n12011));
  jand g11770(.dina(n12011), .dinb(n12006), .dout(n12012));
  jor  g11771(.dina(n12012), .dinb(n3642), .dout(n12013));
  jand g11772(.dina(n12012), .dinb(n3642), .dout(n12014));
  jxor g11773(.dina(n11478), .dinb(n3955), .dout(n12015));
  jor  g11774(.dina(n12015), .dinb(n11858), .dout(n12016));
  jxor g11775(.dina(n12016), .dinb(n11484), .dout(n12017));
  jor  g11776(.dina(n12017), .dinb(n12014), .dout(n12018));
  jand g11777(.dina(n12018), .dinb(n12013), .dout(n12019));
  jor  g11778(.dina(n12019), .dinb(n3368), .dout(n12020));
  jxor g11779(.dina(n11486), .dinb(n3642), .dout(n12021));
  jor  g11780(.dina(n12021), .dinb(n11858), .dout(n12022));
  jxor g11781(.dina(n12022), .dinb(n11679), .dout(n12023));
  jnot g11782(.din(n12023), .dout(n12024));
  jand g11783(.dina(n12019), .dinb(n3368), .dout(n12025));
  jor  g11784(.dina(n12025), .dinb(n12024), .dout(n12026));
  jand g11785(.dina(n12026), .dinb(n12020), .dout(n12027));
  jor  g11786(.dina(n12027), .dinb(n3089), .dout(n12028));
  jand g11787(.dina(n12027), .dinb(n3089), .dout(n12029));
  jxor g11788(.dina(n11493), .dinb(n3368), .dout(n12030));
  jor  g11789(.dina(n12030), .dinb(n11858), .dout(n12031));
  jxor g11790(.dina(n12031), .dinb(n11499), .dout(n12032));
  jor  g11791(.dina(n12032), .dinb(n12029), .dout(n12033));
  jand g11792(.dina(n12033), .dinb(n12028), .dout(n12034));
  jor  g11793(.dina(n12034), .dinb(n2833), .dout(n12035));
  jand g11794(.dina(n12034), .dinb(n2833), .dout(n12036));
  jxor g11795(.dina(n11501), .dinb(n3089), .dout(n12037));
  jor  g11796(.dina(n12037), .dinb(n11858), .dout(n12038));
  jxor g11797(.dina(n12038), .dinb(n11769), .dout(n12039));
  jnot g11798(.din(n12039), .dout(n12040));
  jor  g11799(.dina(n12040), .dinb(n12036), .dout(n12041));
  jand g11800(.dina(n12041), .dinb(n12035), .dout(n12042));
  jor  g11801(.dina(n12042), .dinb(n2572), .dout(n12043));
  jand g11802(.dina(n12042), .dinb(n2572), .dout(n12044));
  jxor g11803(.dina(n11508), .dinb(n2833), .dout(n12045));
  jor  g11804(.dina(n12045), .dinb(n11858), .dout(n12046));
  jxor g11805(.dina(n12046), .dinb(n11514), .dout(n12047));
  jor  g11806(.dina(n12047), .dinb(n12044), .dout(n12048));
  jand g11807(.dina(n12048), .dinb(n12043), .dout(n12049));
  jor  g11808(.dina(n12049), .dinb(n2345), .dout(n12050));
  jand g11809(.dina(n12049), .dinb(n2345), .dout(n12051));
  jxor g11810(.dina(n11516), .dinb(n2572), .dout(n12052));
  jor  g11811(.dina(n12052), .dinb(n11858), .dout(n12053));
  jxor g11812(.dina(n12053), .dinb(n11776), .dout(n12054));
  jnot g11813(.din(n12054), .dout(n12055));
  jor  g11814(.dina(n12055), .dinb(n12051), .dout(n12056));
  jand g11815(.dina(n12056), .dinb(n12050), .dout(n12057));
  jor  g11816(.dina(n12057), .dinb(n2108), .dout(n12058));
  jand g11817(.dina(n12057), .dinb(n2108), .dout(n12059));
  jxor g11818(.dina(n11523), .dinb(n2345), .dout(n12060));
  jor  g11819(.dina(n12060), .dinb(n11858), .dout(n12061));
  jxor g11820(.dina(n12061), .dinb(n11529), .dout(n12062));
  jor  g11821(.dina(n12062), .dinb(n12059), .dout(n12063));
  jand g11822(.dina(n12063), .dinb(n12058), .dout(n12064));
  jor  g11823(.dina(n12064), .dinb(n1912), .dout(n12065));
  jand g11824(.dina(n12064), .dinb(n1912), .dout(n12066));
  jxor g11825(.dina(n11531), .dinb(n2108), .dout(n12067));
  jor  g11826(.dina(n12067), .dinb(n11858), .dout(n12068));
  jxor g11827(.dina(n12068), .dinb(n11537), .dout(n12069));
  jor  g11828(.dina(n12069), .dinb(n12066), .dout(n12070));
  jand g11829(.dina(n12070), .dinb(n12065), .dout(n12071));
  jor  g11830(.dina(n12071), .dinb(n1699), .dout(n12072));
  jand g11831(.dina(n12071), .dinb(n1699), .dout(n12073));
  jxor g11832(.dina(n11539), .dinb(n1912), .dout(n12074));
  jor  g11833(.dina(n12074), .dinb(n11858), .dout(n12075));
  jxor g11834(.dina(n12075), .dinb(n11545), .dout(n12076));
  jor  g11835(.dina(n12076), .dinb(n12073), .dout(n12077));
  jand g11836(.dina(n12077), .dinb(n12072), .dout(n12078));
  jor  g11837(.dina(n12078), .dinb(n1516), .dout(n12079));
  jand g11838(.dina(n12078), .dinb(n1516), .dout(n12080));
  jxor g11839(.dina(n11547), .dinb(n1699), .dout(n12081));
  jor  g11840(.dina(n12081), .dinb(n11858), .dout(n12082));
  jxor g11841(.dina(n12082), .dinb(n11789), .dout(n12083));
  jnot g11842(.din(n12083), .dout(n12084));
  jor  g11843(.dina(n12084), .dinb(n12080), .dout(n12085));
  jand g11844(.dina(n12085), .dinb(n12079), .dout(n12086));
  jor  g11845(.dina(n12086), .dinb(n1332), .dout(n12087));
  jand g11846(.dina(n12086), .dinb(n1332), .dout(n12088));
  jxor g11847(.dina(n11554), .dinb(n1516), .dout(n12089));
  jor  g11848(.dina(n12089), .dinb(n11858), .dout(n12090));
  jxor g11849(.dina(n12090), .dinb(n11560), .dout(n12091));
  jor  g11850(.dina(n12091), .dinb(n12088), .dout(n12092));
  jand g11851(.dina(n12092), .dinb(n12087), .dout(n12093));
  jor  g11852(.dina(n12093), .dinb(n1173), .dout(n12094));
  jand g11853(.dina(n12093), .dinb(n1173), .dout(n12095));
  jxor g11854(.dina(n11562), .dinb(n1332), .dout(n12096));
  jor  g11855(.dina(n12096), .dinb(n11858), .dout(n12097));
  jxor g11856(.dina(n12097), .dinb(n11796), .dout(n12098));
  jnot g11857(.din(n12098), .dout(n12099));
  jor  g11858(.dina(n12099), .dinb(n12095), .dout(n12100));
  jand g11859(.dina(n12100), .dinb(n12094), .dout(n12101));
  jor  g11860(.dina(n12101), .dinb(n1008), .dout(n12102));
  jand g11861(.dina(n12101), .dinb(n1008), .dout(n12103));
  jxor g11862(.dina(n11569), .dinb(n1173), .dout(n12104));
  jor  g11863(.dina(n12104), .dinb(n11858), .dout(n12105));
  jxor g11864(.dina(n12105), .dinb(n11575), .dout(n12106));
  jor  g11865(.dina(n12106), .dinb(n12103), .dout(n12107));
  jand g11866(.dina(n12107), .dinb(n12102), .dout(n12108));
  jor  g11867(.dina(n12108), .dinb(n884), .dout(n12109));
  jand g11868(.dina(n12108), .dinb(n884), .dout(n12110));
  jxor g11869(.dina(n11577), .dinb(n1008), .dout(n12111));
  jor  g11870(.dina(n12111), .dinb(n11858), .dout(n12112));
  jxor g11871(.dina(n12112), .dinb(n11803), .dout(n12113));
  jnot g11872(.din(n12113), .dout(n12114));
  jor  g11873(.dina(n12114), .dinb(n12110), .dout(n12115));
  jand g11874(.dina(n12115), .dinb(n12109), .dout(n12116));
  jor  g11875(.dina(n12116), .dinb(n743), .dout(n12117));
  jand g11876(.dina(n12116), .dinb(n743), .dout(n12118));
  jxor g11877(.dina(n11584), .dinb(n884), .dout(n12119));
  jor  g11878(.dina(n12119), .dinb(n11858), .dout(n12120));
  jxor g11879(.dina(n12120), .dinb(n11590), .dout(n12121));
  jor  g11880(.dina(n12121), .dinb(n12118), .dout(n12122));
  jand g11881(.dina(n12122), .dinb(n12117), .dout(n12123));
  jor  g11882(.dina(n12123), .dinb(n635), .dout(n12124));
  jand g11883(.dina(n12123), .dinb(n635), .dout(n12125));
  jxor g11884(.dina(n11592), .dinb(n743), .dout(n12126));
  jor  g11885(.dina(n12126), .dinb(n11858), .dout(n12127));
  jxor g11886(.dina(n12127), .dinb(n11810), .dout(n12128));
  jnot g11887(.din(n12128), .dout(n12129));
  jor  g11888(.dina(n12129), .dinb(n12125), .dout(n12130));
  jand g11889(.dina(n12130), .dinb(n12124), .dout(n12131));
  jor  g11890(.dina(n12131), .dinb(n515), .dout(n12132));
  jand g11891(.dina(n12131), .dinb(n515), .dout(n12133));
  jxor g11892(.dina(n11599), .dinb(n635), .dout(n12134));
  jor  g11893(.dina(n12134), .dinb(n11858), .dout(n12135));
  jxor g11894(.dina(n12135), .dinb(n11814), .dout(n12136));
  jnot g11895(.din(n12136), .dout(n12137));
  jor  g11896(.dina(n12137), .dinb(n12133), .dout(n12138));
  jand g11897(.dina(n12138), .dinb(n12132), .dout(n12139));
  jor  g11898(.dina(n12139), .dinb(n443), .dout(n12140));
  jand g11899(.dina(n12139), .dinb(n443), .dout(n12141));
  jxor g11900(.dina(n11606), .dinb(n515), .dout(n12142));
  jor  g11901(.dina(n12142), .dinb(n11858), .dout(n12143));
  jxor g11902(.dina(n12143), .dinb(n11818), .dout(n12144));
  jnot g11903(.din(n12144), .dout(n12145));
  jor  g11904(.dina(n12145), .dinb(n12141), .dout(n12146));
  jand g11905(.dina(n12146), .dinb(n12140), .dout(n12147));
  jor  g11906(.dina(n12147), .dinb(n352), .dout(n12148));
  jand g11907(.dina(n12147), .dinb(n352), .dout(n12149));
  jxor g11908(.dina(n11613), .dinb(n443), .dout(n12150));
  jor  g11909(.dina(n12150), .dinb(n11858), .dout(n12151));
  jxor g11910(.dina(n12151), .dinb(n11619), .dout(n12152));
  jor  g11911(.dina(n12152), .dinb(n12149), .dout(n12153));
  jand g11912(.dina(n12153), .dinb(n12148), .dout(n12154));
  jor  g11913(.dina(n12154), .dinb(n294), .dout(n12155));
  jand g11914(.dina(n12154), .dinb(n294), .dout(n12156));
  jxor g11915(.dina(n11621), .dinb(n352), .dout(n12157));
  jor  g11916(.dina(n12157), .dinb(n11858), .dout(n12158));
  jxor g11917(.dina(n12158), .dinb(n11627), .dout(n12159));
  jor  g11918(.dina(n12159), .dinb(n12156), .dout(n12160));
  jand g11919(.dina(n12160), .dinb(n12155), .dout(n12161));
  jor  g11920(.dina(n12161), .dinb(n239), .dout(n12162));
  jand g11921(.dina(n12161), .dinb(n239), .dout(n12163));
  jxor g11922(.dina(n11629), .dinb(n294), .dout(n12164));
  jor  g11923(.dina(n12164), .dinb(n11858), .dout(n12165));
  jxor g11924(.dina(n12165), .dinb(n11635), .dout(n12166));
  jor  g11925(.dina(n12166), .dinb(n12163), .dout(n12167));
  jand g11926(.dina(n12167), .dinb(n12162), .dout(n12168));
  jor  g11927(.dina(n12168), .dinb(n221), .dout(n12169));
  jand g11928(.dina(n12168), .dinb(n221), .dout(n12170));
  jxor g11929(.dina(n11637), .dinb(n239), .dout(n12171));
  jor  g11930(.dina(n12171), .dinb(n11858), .dout(n12172));
  jxor g11931(.dina(n12172), .dinb(n11831), .dout(n12173));
  jnot g11932(.din(n12173), .dout(n12174));
  jor  g11933(.dina(n12174), .dinb(n12170), .dout(n12175));
  jand g11934(.dina(n12175), .dinb(n12169), .dout(n12176));
  jand g11935(.dina(n12176), .dinb(n11862), .dout(n12177));
  jand g11936(.dina(n11847), .dinb(n11851), .dout(n12179));
  jor  g11937(.dina(n12176), .dinb(n11862), .dout(n12180));
  jor  g11938(.dina(n12180), .dinb(n11654), .dout(n12181));
  jor  g11939(.dina(n12181), .dinb(n12179), .dout(n12182));
  jand g11940(.dina(n12182), .dinb(n218), .dout(n12183));
  jand g11941(.dina(n11856), .dinb(n11836), .dout(n12184));
  jand g11942(.dina(n11837), .dinb(asqrt[63] ), .dout(n12185));
  jand g11943(.dina(n12185), .dinb(n11653), .dout(n12186));
  jnot g11944(.din(n12186), .dout(n12187));
  jor  g11945(.dina(n12187), .dinb(n12184), .dout(n12188));
  jnot g11946(.din(n12188), .dout(n12189));
  jor  g11947(.dina(n12189), .dinb(n12183), .dout(n12190));
  jor  g11948(.dina(n12190), .dinb(n12177), .dout(asqrt[20] ));
  jxor g11949(.dina(n12168), .dinb(n221), .dout(n12193));
  jand g11950(.dina(n12193), .dinb(asqrt[20] ), .dout(n12194));
  jxor g11951(.dina(n12194), .dinb(n12173), .dout(n12195));
  jnot g11952(.din(a[38] ), .dout(n12196));
  jnot g11953(.din(a[39] ), .dout(n12197));
  jand g11954(.dina(n12197), .dinb(n12196), .dout(n12198));
  jand g11955(.dina(n12198), .dinb(n11864), .dout(n12199));
  jand g11956(.dina(asqrt[20] ), .dinb(a[40] ), .dout(n12200));
  jor  g11957(.dina(n12200), .dinb(n12199), .dout(n12201));
  jand g11958(.dina(n12201), .dinb(asqrt[21] ), .dout(n12202));
  jor  g11959(.dina(n12201), .dinb(asqrt[21] ), .dout(n12203));
  jand g11960(.dina(asqrt[20] ), .dinb(n11864), .dout(n12204));
  jor  g11961(.dina(n12204), .dinb(n11865), .dout(n12205));
  jnot g11962(.din(n11866), .dout(n12206));
  jnot g11963(.din(n12177), .dout(n12207));
  jnot g11964(.din(n12179), .dout(n12209));
  jnot g11965(.din(n12169), .dout(n12210));
  jnot g11966(.din(n12162), .dout(n12211));
  jnot g11967(.din(n12155), .dout(n12212));
  jnot g11968(.din(n12148), .dout(n12213));
  jnot g11969(.din(n12140), .dout(n12214));
  jnot g11970(.din(n12132), .dout(n12215));
  jnot g11971(.din(n12124), .dout(n12216));
  jnot g11972(.din(n12117), .dout(n12217));
  jnot g11973(.din(n12109), .dout(n12218));
  jnot g11974(.din(n12102), .dout(n12219));
  jnot g11975(.din(n12094), .dout(n12220));
  jnot g11976(.din(n12087), .dout(n12221));
  jnot g11977(.din(n12079), .dout(n12222));
  jnot g11978(.din(n12072), .dout(n12223));
  jnot g11979(.din(n12065), .dout(n12224));
  jnot g11980(.din(n12058), .dout(n12225));
  jnot g11981(.din(n12050), .dout(n12226));
  jnot g11982(.din(n12043), .dout(n12227));
  jnot g11983(.din(n12035), .dout(n12228));
  jnot g11984(.din(n12028), .dout(n12229));
  jnot g11985(.din(n12020), .dout(n12230));
  jnot g11986(.din(n12013), .dout(n12231));
  jnot g11987(.din(n12006), .dout(n12232));
  jnot g11988(.din(n11999), .dout(n12233));
  jnot g11989(.din(n11992), .dout(n12234));
  jnot g11990(.din(n11985), .dout(n12235));
  jnot g11991(.din(n11977), .dout(n12236));
  jnot g11992(.din(n11970), .dout(n12237));
  jnot g11993(.din(n11963), .dout(n12238));
  jnot g11994(.din(n11956), .dout(n12239));
  jnot g11995(.din(n11948), .dout(n12240));
  jnot g11996(.din(n11941), .dout(n12241));
  jnot g11997(.din(n11933), .dout(n12242));
  jnot g11998(.din(n11926), .dout(n12243));
  jnot g11999(.din(n11919), .dout(n12244));
  jnot g12000(.din(n11912), .dout(n12245));
  jnot g12001(.din(n11904), .dout(n12246));
  jnot g12002(.din(n11897), .dout(n12247));
  jnot g12003(.din(n11889), .dout(n12248));
  jnot g12004(.din(n11878), .dout(n12249));
  jnot g12005(.din(n11870), .dout(n12250));
  jand g12006(.dina(asqrt[21] ), .dinb(a[42] ), .dout(n12251));
  jor  g12007(.dina(n11867), .dinb(n12251), .dout(n12252));
  jor  g12008(.dina(n12252), .dinb(asqrt[22] ), .dout(n12253));
  jand g12009(.dina(asqrt[21] ), .dinb(n11142), .dout(n12254));
  jor  g12010(.dina(n12254), .dinb(n11143), .dout(n12255));
  jand g12011(.dina(n11881), .dinb(n12255), .dout(n12256));
  jand g12012(.dina(n12256), .dinb(n12253), .dout(n12257));
  jor  g12013(.dina(n12257), .dinb(n12250), .dout(n12258));
  jor  g12014(.dina(n12258), .dinb(asqrt[23] ), .dout(n12259));
  jnot g12015(.din(n11886), .dout(n12260));
  jand g12016(.dina(n12260), .dinb(n12259), .dout(n12261));
  jor  g12017(.dina(n12261), .dinb(n12249), .dout(n12262));
  jor  g12018(.dina(n12262), .dinb(asqrt[24] ), .dout(n12263));
  jand g12019(.dina(n11893), .dinb(n12263), .dout(n12264));
  jor  g12020(.dina(n12264), .dinb(n12248), .dout(n12265));
  jor  g12021(.dina(n12265), .dinb(asqrt[25] ), .dout(n12266));
  jnot g12022(.din(n11901), .dout(n12267));
  jand g12023(.dina(n12267), .dinb(n12266), .dout(n12268));
  jor  g12024(.dina(n12268), .dinb(n12247), .dout(n12269));
  jor  g12025(.dina(n12269), .dinb(asqrt[26] ), .dout(n12270));
  jand g12026(.dina(n11908), .dinb(n12270), .dout(n12271));
  jor  g12027(.dina(n12271), .dinb(n12246), .dout(n12272));
  jor  g12028(.dina(n12272), .dinb(asqrt[27] ), .dout(n12273));
  jnot g12029(.din(n11916), .dout(n12274));
  jand g12030(.dina(n12274), .dinb(n12273), .dout(n12275));
  jor  g12031(.dina(n12275), .dinb(n12245), .dout(n12276));
  jor  g12032(.dina(n12276), .dinb(asqrt[28] ), .dout(n12277));
  jnot g12033(.din(n11923), .dout(n12278));
  jand g12034(.dina(n12278), .dinb(n12277), .dout(n12279));
  jor  g12035(.dina(n12279), .dinb(n12244), .dout(n12280));
  jor  g12036(.dina(n12280), .dinb(asqrt[29] ), .dout(n12281));
  jnot g12037(.din(n11930), .dout(n12282));
  jand g12038(.dina(n12282), .dinb(n12281), .dout(n12283));
  jor  g12039(.dina(n12283), .dinb(n12243), .dout(n12284));
  jor  g12040(.dina(n12284), .dinb(asqrt[30] ), .dout(n12285));
  jand g12041(.dina(n11937), .dinb(n12285), .dout(n12286));
  jor  g12042(.dina(n12286), .dinb(n12242), .dout(n12287));
  jor  g12043(.dina(n12287), .dinb(asqrt[31] ), .dout(n12288));
  jnot g12044(.din(n11945), .dout(n12289));
  jand g12045(.dina(n12289), .dinb(n12288), .dout(n12290));
  jor  g12046(.dina(n12290), .dinb(n12241), .dout(n12291));
  jor  g12047(.dina(n12291), .dinb(asqrt[32] ), .dout(n12292));
  jand g12048(.dina(n11952), .dinb(n12292), .dout(n12293));
  jor  g12049(.dina(n12293), .dinb(n12240), .dout(n12294));
  jor  g12050(.dina(n12294), .dinb(asqrt[33] ), .dout(n12295));
  jnot g12051(.din(n11960), .dout(n12296));
  jand g12052(.dina(n12296), .dinb(n12295), .dout(n12297));
  jor  g12053(.dina(n12297), .dinb(n12239), .dout(n12298));
  jor  g12054(.dina(n12298), .dinb(asqrt[34] ), .dout(n12299));
  jnot g12055(.din(n11967), .dout(n12300));
  jand g12056(.dina(n12300), .dinb(n12299), .dout(n12301));
  jor  g12057(.dina(n12301), .dinb(n12238), .dout(n12302));
  jor  g12058(.dina(n12302), .dinb(asqrt[35] ), .dout(n12303));
  jnot g12059(.din(n11974), .dout(n12304));
  jand g12060(.dina(n12304), .dinb(n12303), .dout(n12305));
  jor  g12061(.dina(n12305), .dinb(n12237), .dout(n12306));
  jor  g12062(.dina(n12306), .dinb(asqrt[36] ), .dout(n12307));
  jand g12063(.dina(n11981), .dinb(n12307), .dout(n12308));
  jor  g12064(.dina(n12308), .dinb(n12236), .dout(n12309));
  jor  g12065(.dina(n12309), .dinb(asqrt[37] ), .dout(n12310));
  jnot g12066(.din(n11989), .dout(n12311));
  jand g12067(.dina(n12311), .dinb(n12310), .dout(n12312));
  jor  g12068(.dina(n12312), .dinb(n12235), .dout(n12313));
  jor  g12069(.dina(n12313), .dinb(asqrt[38] ), .dout(n12314));
  jnot g12070(.din(n11996), .dout(n12315));
  jand g12071(.dina(n12315), .dinb(n12314), .dout(n12316));
  jor  g12072(.dina(n12316), .dinb(n12234), .dout(n12317));
  jor  g12073(.dina(n12317), .dinb(asqrt[39] ), .dout(n12318));
  jnot g12074(.din(n12003), .dout(n12319));
  jand g12075(.dina(n12319), .dinb(n12318), .dout(n12320));
  jor  g12076(.dina(n12320), .dinb(n12233), .dout(n12321));
  jor  g12077(.dina(n12321), .dinb(asqrt[40] ), .dout(n12322));
  jnot g12078(.din(n12010), .dout(n12323));
  jand g12079(.dina(n12323), .dinb(n12322), .dout(n12324));
  jor  g12080(.dina(n12324), .dinb(n12232), .dout(n12325));
  jor  g12081(.dina(n12325), .dinb(asqrt[41] ), .dout(n12326));
  jnot g12082(.din(n12017), .dout(n12327));
  jand g12083(.dina(n12327), .dinb(n12326), .dout(n12328));
  jor  g12084(.dina(n12328), .dinb(n12231), .dout(n12329));
  jor  g12085(.dina(n12329), .dinb(asqrt[42] ), .dout(n12330));
  jand g12086(.dina(n12330), .dinb(n12023), .dout(n12331));
  jor  g12087(.dina(n12331), .dinb(n12230), .dout(n12332));
  jor  g12088(.dina(n12332), .dinb(asqrt[43] ), .dout(n12333));
  jnot g12089(.din(n12032), .dout(n12334));
  jand g12090(.dina(n12334), .dinb(n12333), .dout(n12335));
  jor  g12091(.dina(n12335), .dinb(n12229), .dout(n12336));
  jor  g12092(.dina(n12336), .dinb(asqrt[44] ), .dout(n12337));
  jand g12093(.dina(n12039), .dinb(n12337), .dout(n12338));
  jor  g12094(.dina(n12338), .dinb(n12228), .dout(n12339));
  jor  g12095(.dina(n12339), .dinb(asqrt[45] ), .dout(n12340));
  jnot g12096(.din(n12047), .dout(n12341));
  jand g12097(.dina(n12341), .dinb(n12340), .dout(n12342));
  jor  g12098(.dina(n12342), .dinb(n12227), .dout(n12343));
  jor  g12099(.dina(n12343), .dinb(asqrt[46] ), .dout(n12344));
  jand g12100(.dina(n12054), .dinb(n12344), .dout(n12345));
  jor  g12101(.dina(n12345), .dinb(n12226), .dout(n12346));
  jor  g12102(.dina(n12346), .dinb(asqrt[47] ), .dout(n12347));
  jnot g12103(.din(n12062), .dout(n12348));
  jand g12104(.dina(n12348), .dinb(n12347), .dout(n12349));
  jor  g12105(.dina(n12349), .dinb(n12225), .dout(n12350));
  jor  g12106(.dina(n12350), .dinb(asqrt[48] ), .dout(n12351));
  jnot g12107(.din(n12069), .dout(n12352));
  jand g12108(.dina(n12352), .dinb(n12351), .dout(n12353));
  jor  g12109(.dina(n12353), .dinb(n12224), .dout(n12354));
  jor  g12110(.dina(n12354), .dinb(asqrt[49] ), .dout(n12355));
  jnot g12111(.din(n12076), .dout(n12356));
  jand g12112(.dina(n12356), .dinb(n12355), .dout(n12357));
  jor  g12113(.dina(n12357), .dinb(n12223), .dout(n12358));
  jor  g12114(.dina(n12358), .dinb(asqrt[50] ), .dout(n12359));
  jand g12115(.dina(n12083), .dinb(n12359), .dout(n12360));
  jor  g12116(.dina(n12360), .dinb(n12222), .dout(n12361));
  jor  g12117(.dina(n12361), .dinb(asqrt[51] ), .dout(n12362));
  jnot g12118(.din(n12091), .dout(n12363));
  jand g12119(.dina(n12363), .dinb(n12362), .dout(n12364));
  jor  g12120(.dina(n12364), .dinb(n12221), .dout(n12365));
  jor  g12121(.dina(n12365), .dinb(asqrt[52] ), .dout(n12366));
  jand g12122(.dina(n12098), .dinb(n12366), .dout(n12367));
  jor  g12123(.dina(n12367), .dinb(n12220), .dout(n12368));
  jor  g12124(.dina(n12368), .dinb(asqrt[53] ), .dout(n12369));
  jnot g12125(.din(n12106), .dout(n12370));
  jand g12126(.dina(n12370), .dinb(n12369), .dout(n12371));
  jor  g12127(.dina(n12371), .dinb(n12219), .dout(n12372));
  jor  g12128(.dina(n12372), .dinb(asqrt[54] ), .dout(n12373));
  jand g12129(.dina(n12113), .dinb(n12373), .dout(n12374));
  jor  g12130(.dina(n12374), .dinb(n12218), .dout(n12375));
  jor  g12131(.dina(n12375), .dinb(asqrt[55] ), .dout(n12376));
  jnot g12132(.din(n12121), .dout(n12377));
  jand g12133(.dina(n12377), .dinb(n12376), .dout(n12378));
  jor  g12134(.dina(n12378), .dinb(n12217), .dout(n12379));
  jor  g12135(.dina(n12379), .dinb(asqrt[56] ), .dout(n12380));
  jand g12136(.dina(n12128), .dinb(n12380), .dout(n12381));
  jor  g12137(.dina(n12381), .dinb(n12216), .dout(n12382));
  jor  g12138(.dina(n12382), .dinb(asqrt[57] ), .dout(n12383));
  jand g12139(.dina(n12136), .dinb(n12383), .dout(n12384));
  jor  g12140(.dina(n12384), .dinb(n12215), .dout(n12385));
  jor  g12141(.dina(n12385), .dinb(asqrt[58] ), .dout(n12386));
  jand g12142(.dina(n12144), .dinb(n12386), .dout(n12387));
  jor  g12143(.dina(n12387), .dinb(n12214), .dout(n12388));
  jor  g12144(.dina(n12388), .dinb(asqrt[59] ), .dout(n12389));
  jnot g12145(.din(n12152), .dout(n12390));
  jand g12146(.dina(n12390), .dinb(n12389), .dout(n12391));
  jor  g12147(.dina(n12391), .dinb(n12213), .dout(n12392));
  jor  g12148(.dina(n12392), .dinb(asqrt[60] ), .dout(n12393));
  jnot g12149(.din(n12159), .dout(n12394));
  jand g12150(.dina(n12394), .dinb(n12393), .dout(n12395));
  jor  g12151(.dina(n12395), .dinb(n12212), .dout(n12396));
  jor  g12152(.dina(n12396), .dinb(asqrt[61] ), .dout(n12397));
  jnot g12153(.din(n12166), .dout(n12398));
  jand g12154(.dina(n12398), .dinb(n12397), .dout(n12399));
  jor  g12155(.dina(n12399), .dinb(n12211), .dout(n12400));
  jor  g12156(.dina(n12400), .dinb(asqrt[62] ), .dout(n12401));
  jand g12157(.dina(n12173), .dinb(n12401), .dout(n12402));
  jor  g12158(.dina(n12402), .dinb(n12210), .dout(n12403));
  jand g12159(.dina(n12403), .dinb(n11861), .dout(n12404));
  jand g12160(.dina(n12404), .dinb(n11653), .dout(n12405));
  jand g12161(.dina(n12405), .dinb(n12209), .dout(n12406));
  jor  g12162(.dina(n12406), .dinb(asqrt[63] ), .dout(n12407));
  jand g12163(.dina(n12188), .dinb(n12407), .dout(n12408));
  jand g12164(.dina(n12408), .dinb(n12207), .dout(n12410));
  jor  g12165(.dina(n12410), .dinb(n12206), .dout(n12411));
  jand g12166(.dina(n12411), .dinb(n12205), .dout(n12412));
  jand g12167(.dina(n12412), .dinb(n12203), .dout(n12413));
  jor  g12168(.dina(n12413), .dinb(n12202), .dout(n12414));
  jand g12169(.dina(n12414), .dinb(asqrt[22] ), .dout(n12415));
  jor  g12170(.dina(n12414), .dinb(asqrt[22] ), .dout(n12416));
  jand g12171(.dina(asqrt[20] ), .dinb(n11866), .dout(n12417));
  jand g12172(.dina(n12187), .dinb(n12207), .dout(n12418));
  jand g12173(.dina(n12418), .dinb(n12407), .dout(n12419));
  jand g12174(.dina(n12419), .dinb(asqrt[21] ), .dout(n12420));
  jor  g12175(.dina(n12420), .dinb(n12417), .dout(n12421));
  jxor g12176(.dina(n12421), .dinb(a[42] ), .dout(n12422));
  jnot g12177(.din(n12422), .dout(n12423));
  jand g12178(.dina(n12423), .dinb(n12416), .dout(n12424));
  jor  g12179(.dina(n12424), .dinb(n12415), .dout(n12425));
  jand g12180(.dina(n12425), .dinb(asqrt[23] ), .dout(n12426));
  jor  g12181(.dina(n12425), .dinb(asqrt[23] ), .dout(n12427));
  jxor g12182(.dina(n11869), .dinb(n11347), .dout(n12428));
  jand g12183(.dina(n12428), .dinb(asqrt[20] ), .dout(n12429));
  jxor g12184(.dina(n12429), .dinb(n12256), .dout(n12430));
  jand g12185(.dina(n12430), .dinb(n12427), .dout(n12431));
  jor  g12186(.dina(n12431), .dinb(n12426), .dout(n12432));
  jand g12187(.dina(n12432), .dinb(asqrt[24] ), .dout(n12433));
  jor  g12188(.dina(n12432), .dinb(asqrt[24] ), .dout(n12434));
  jxor g12189(.dina(n11877), .dinb(n10824), .dout(n12435));
  jand g12190(.dina(n12435), .dinb(asqrt[20] ), .dout(n12436));
  jxor g12191(.dina(n12436), .dinb(n11886), .dout(n12437));
  jnot g12192(.din(n12437), .dout(n12438));
  jand g12193(.dina(n12438), .dinb(n12434), .dout(n12439));
  jor  g12194(.dina(n12439), .dinb(n12433), .dout(n12440));
  jand g12195(.dina(n12440), .dinb(asqrt[25] ), .dout(n12441));
  jor  g12196(.dina(n12440), .dinb(asqrt[25] ), .dout(n12442));
  jxor g12197(.dina(n11888), .dinb(n10328), .dout(n12443));
  jand g12198(.dina(n12443), .dinb(asqrt[20] ), .dout(n12444));
  jxor g12199(.dina(n12444), .dinb(n11893), .dout(n12445));
  jand g12200(.dina(n12445), .dinb(n12442), .dout(n12446));
  jor  g12201(.dina(n12446), .dinb(n12441), .dout(n12447));
  jand g12202(.dina(n12447), .dinb(asqrt[26] ), .dout(n12448));
  jor  g12203(.dina(n12447), .dinb(asqrt[26] ), .dout(n12449));
  jxor g12204(.dina(n11896), .dinb(n9832), .dout(n12450));
  jand g12205(.dina(n12450), .dinb(asqrt[20] ), .dout(n12451));
  jxor g12206(.dina(n12451), .dinb(n11901), .dout(n12452));
  jnot g12207(.din(n12452), .dout(n12453));
  jand g12208(.dina(n12453), .dinb(n12449), .dout(n12454));
  jor  g12209(.dina(n12454), .dinb(n12448), .dout(n12455));
  jand g12210(.dina(n12455), .dinb(asqrt[27] ), .dout(n12456));
  jor  g12211(.dina(n12455), .dinb(asqrt[27] ), .dout(n12457));
  jxor g12212(.dina(n11903), .dinb(n9369), .dout(n12458));
  jand g12213(.dina(n12458), .dinb(asqrt[20] ), .dout(n12459));
  jxor g12214(.dina(n12459), .dinb(n11908), .dout(n12460));
  jand g12215(.dina(n12460), .dinb(n12457), .dout(n12461));
  jor  g12216(.dina(n12461), .dinb(n12456), .dout(n12462));
  jand g12217(.dina(n12462), .dinb(asqrt[28] ), .dout(n12463));
  jor  g12218(.dina(n12462), .dinb(asqrt[28] ), .dout(n12464));
  jxor g12219(.dina(n11911), .dinb(n8890), .dout(n12465));
  jand g12220(.dina(n12465), .dinb(asqrt[20] ), .dout(n12466));
  jxor g12221(.dina(n12466), .dinb(n11916), .dout(n12467));
  jnot g12222(.din(n12467), .dout(n12468));
  jand g12223(.dina(n12468), .dinb(n12464), .dout(n12469));
  jor  g12224(.dina(n12469), .dinb(n12463), .dout(n12470));
  jand g12225(.dina(n12470), .dinb(asqrt[29] ), .dout(n12471));
  jor  g12226(.dina(n12470), .dinb(asqrt[29] ), .dout(n12472));
  jxor g12227(.dina(n11918), .dinb(n8449), .dout(n12473));
  jand g12228(.dina(n12473), .dinb(asqrt[20] ), .dout(n12474));
  jxor g12229(.dina(n12474), .dinb(n11923), .dout(n12475));
  jnot g12230(.din(n12475), .dout(n12476));
  jand g12231(.dina(n12476), .dinb(n12472), .dout(n12477));
  jor  g12232(.dina(n12477), .dinb(n12471), .dout(n12478));
  jand g12233(.dina(n12478), .dinb(asqrt[30] ), .dout(n12479));
  jor  g12234(.dina(n12478), .dinb(asqrt[30] ), .dout(n12480));
  jxor g12235(.dina(n11925), .dinb(n8003), .dout(n12481));
  jand g12236(.dina(n12481), .dinb(asqrt[20] ), .dout(n12482));
  jxor g12237(.dina(n12482), .dinb(n11930), .dout(n12483));
  jnot g12238(.din(n12483), .dout(n12484));
  jand g12239(.dina(n12484), .dinb(n12480), .dout(n12485));
  jor  g12240(.dina(n12485), .dinb(n12479), .dout(n12486));
  jand g12241(.dina(n12486), .dinb(asqrt[31] ), .dout(n12487));
  jor  g12242(.dina(n12486), .dinb(asqrt[31] ), .dout(n12488));
  jxor g12243(.dina(n11932), .dinb(n7581), .dout(n12489));
  jand g12244(.dina(n12489), .dinb(asqrt[20] ), .dout(n12490));
  jxor g12245(.dina(n12490), .dinb(n11937), .dout(n12491));
  jand g12246(.dina(n12491), .dinb(n12488), .dout(n12492));
  jor  g12247(.dina(n12492), .dinb(n12487), .dout(n12493));
  jand g12248(.dina(n12493), .dinb(asqrt[32] ), .dout(n12494));
  jor  g12249(.dina(n12493), .dinb(asqrt[32] ), .dout(n12495));
  jxor g12250(.dina(n11940), .dinb(n7154), .dout(n12496));
  jand g12251(.dina(n12496), .dinb(asqrt[20] ), .dout(n12497));
  jxor g12252(.dina(n12497), .dinb(n11945), .dout(n12498));
  jnot g12253(.din(n12498), .dout(n12499));
  jand g12254(.dina(n12499), .dinb(n12495), .dout(n12500));
  jor  g12255(.dina(n12500), .dinb(n12494), .dout(n12501));
  jand g12256(.dina(n12501), .dinb(asqrt[33] ), .dout(n12502));
  jor  g12257(.dina(n12501), .dinb(asqrt[33] ), .dout(n12503));
  jxor g12258(.dina(n11947), .dinb(n6758), .dout(n12504));
  jand g12259(.dina(n12504), .dinb(asqrt[20] ), .dout(n12505));
  jxor g12260(.dina(n12505), .dinb(n11952), .dout(n12506));
  jand g12261(.dina(n12506), .dinb(n12503), .dout(n12507));
  jor  g12262(.dina(n12507), .dinb(n12502), .dout(n12508));
  jand g12263(.dina(n12508), .dinb(asqrt[34] ), .dout(n12509));
  jor  g12264(.dina(n12508), .dinb(asqrt[34] ), .dout(n12510));
  jxor g12265(.dina(n11955), .dinb(n6357), .dout(n12511));
  jand g12266(.dina(n12511), .dinb(asqrt[20] ), .dout(n12512));
  jxor g12267(.dina(n12512), .dinb(n11960), .dout(n12513));
  jnot g12268(.din(n12513), .dout(n12514));
  jand g12269(.dina(n12514), .dinb(n12510), .dout(n12515));
  jor  g12270(.dina(n12515), .dinb(n12509), .dout(n12516));
  jand g12271(.dina(n12516), .dinb(asqrt[35] ), .dout(n12517));
  jor  g12272(.dina(n12516), .dinb(asqrt[35] ), .dout(n12518));
  jxor g12273(.dina(n11962), .dinb(n5989), .dout(n12519));
  jand g12274(.dina(n12519), .dinb(asqrt[20] ), .dout(n12520));
  jxor g12275(.dina(n12520), .dinb(n11967), .dout(n12521));
  jnot g12276(.din(n12521), .dout(n12522));
  jand g12277(.dina(n12522), .dinb(n12518), .dout(n12523));
  jor  g12278(.dina(n12523), .dinb(n12517), .dout(n12524));
  jand g12279(.dina(n12524), .dinb(asqrt[36] ), .dout(n12525));
  jor  g12280(.dina(n12524), .dinb(asqrt[36] ), .dout(n12526));
  jxor g12281(.dina(n11969), .dinb(n5606), .dout(n12527));
  jand g12282(.dina(n12527), .dinb(asqrt[20] ), .dout(n12528));
  jxor g12283(.dina(n12528), .dinb(n11974), .dout(n12529));
  jnot g12284(.din(n12529), .dout(n12530));
  jand g12285(.dina(n12530), .dinb(n12526), .dout(n12531));
  jor  g12286(.dina(n12531), .dinb(n12525), .dout(n12532));
  jand g12287(.dina(n12532), .dinb(asqrt[37] ), .dout(n12533));
  jor  g12288(.dina(n12532), .dinb(asqrt[37] ), .dout(n12534));
  jxor g12289(.dina(n11976), .dinb(n5259), .dout(n12535));
  jand g12290(.dina(n12535), .dinb(asqrt[20] ), .dout(n12536));
  jxor g12291(.dina(n12536), .dinb(n11981), .dout(n12537));
  jand g12292(.dina(n12537), .dinb(n12534), .dout(n12538));
  jor  g12293(.dina(n12538), .dinb(n12533), .dout(n12539));
  jand g12294(.dina(n12539), .dinb(asqrt[38] ), .dout(n12540));
  jor  g12295(.dina(n12539), .dinb(asqrt[38] ), .dout(n12541));
  jxor g12296(.dina(n11984), .dinb(n4902), .dout(n12542));
  jand g12297(.dina(n12542), .dinb(asqrt[20] ), .dout(n12543));
  jxor g12298(.dina(n12543), .dinb(n11989), .dout(n12544));
  jnot g12299(.din(n12544), .dout(n12545));
  jand g12300(.dina(n12545), .dinb(n12541), .dout(n12546));
  jor  g12301(.dina(n12546), .dinb(n12540), .dout(n12547));
  jand g12302(.dina(n12547), .dinb(asqrt[39] ), .dout(n12548));
  jor  g12303(.dina(n12547), .dinb(asqrt[39] ), .dout(n12549));
  jxor g12304(.dina(n11991), .dinb(n4582), .dout(n12550));
  jand g12305(.dina(n12550), .dinb(asqrt[20] ), .dout(n12551));
  jxor g12306(.dina(n12551), .dinb(n11996), .dout(n12552));
  jnot g12307(.din(n12552), .dout(n12553));
  jand g12308(.dina(n12553), .dinb(n12549), .dout(n12554));
  jor  g12309(.dina(n12554), .dinb(n12548), .dout(n12555));
  jand g12310(.dina(n12555), .dinb(asqrt[40] ), .dout(n12556));
  jor  g12311(.dina(n12555), .dinb(asqrt[40] ), .dout(n12557));
  jxor g12312(.dina(n11998), .dinb(n4249), .dout(n12558));
  jand g12313(.dina(n12558), .dinb(asqrt[20] ), .dout(n12559));
  jxor g12314(.dina(n12559), .dinb(n12003), .dout(n12560));
  jnot g12315(.din(n12560), .dout(n12561));
  jand g12316(.dina(n12561), .dinb(n12557), .dout(n12562));
  jor  g12317(.dina(n12562), .dinb(n12556), .dout(n12563));
  jand g12318(.dina(n12563), .dinb(asqrt[41] ), .dout(n12564));
  jor  g12319(.dina(n12563), .dinb(asqrt[41] ), .dout(n12565));
  jxor g12320(.dina(n12005), .dinb(n3955), .dout(n12566));
  jand g12321(.dina(n12566), .dinb(asqrt[20] ), .dout(n12567));
  jxor g12322(.dina(n12567), .dinb(n12010), .dout(n12568));
  jnot g12323(.din(n12568), .dout(n12569));
  jand g12324(.dina(n12569), .dinb(n12565), .dout(n12570));
  jor  g12325(.dina(n12570), .dinb(n12564), .dout(n12571));
  jand g12326(.dina(n12571), .dinb(asqrt[42] ), .dout(n12572));
  jor  g12327(.dina(n12571), .dinb(asqrt[42] ), .dout(n12573));
  jxor g12328(.dina(n12012), .dinb(n3642), .dout(n12574));
  jand g12329(.dina(n12574), .dinb(asqrt[20] ), .dout(n12575));
  jxor g12330(.dina(n12575), .dinb(n12017), .dout(n12576));
  jnot g12331(.din(n12576), .dout(n12577));
  jand g12332(.dina(n12577), .dinb(n12573), .dout(n12578));
  jor  g12333(.dina(n12578), .dinb(n12572), .dout(n12579));
  jand g12334(.dina(n12579), .dinb(asqrt[43] ), .dout(n12580));
  jxor g12335(.dina(n12019), .dinb(n3368), .dout(n12581));
  jand g12336(.dina(n12581), .dinb(asqrt[20] ), .dout(n12582));
  jxor g12337(.dina(n12582), .dinb(n12023), .dout(n12583));
  jor  g12338(.dina(n12579), .dinb(asqrt[43] ), .dout(n12584));
  jand g12339(.dina(n12584), .dinb(n12583), .dout(n12585));
  jor  g12340(.dina(n12585), .dinb(n12580), .dout(n12586));
  jand g12341(.dina(n12586), .dinb(asqrt[44] ), .dout(n12587));
  jor  g12342(.dina(n12586), .dinb(asqrt[44] ), .dout(n12588));
  jxor g12343(.dina(n12027), .dinb(n3089), .dout(n12589));
  jand g12344(.dina(n12589), .dinb(asqrt[20] ), .dout(n12590));
  jxor g12345(.dina(n12590), .dinb(n12032), .dout(n12591));
  jnot g12346(.din(n12591), .dout(n12592));
  jand g12347(.dina(n12592), .dinb(n12588), .dout(n12593));
  jor  g12348(.dina(n12593), .dinb(n12587), .dout(n12594));
  jand g12349(.dina(n12594), .dinb(asqrt[45] ), .dout(n12595));
  jor  g12350(.dina(n12594), .dinb(asqrt[45] ), .dout(n12596));
  jxor g12351(.dina(n12034), .dinb(n2833), .dout(n12597));
  jand g12352(.dina(n12597), .dinb(asqrt[20] ), .dout(n12598));
  jxor g12353(.dina(n12598), .dinb(n12039), .dout(n12599));
  jand g12354(.dina(n12599), .dinb(n12596), .dout(n12600));
  jor  g12355(.dina(n12600), .dinb(n12595), .dout(n12601));
  jand g12356(.dina(n12601), .dinb(asqrt[46] ), .dout(n12602));
  jor  g12357(.dina(n12601), .dinb(asqrt[46] ), .dout(n12603));
  jxor g12358(.dina(n12042), .dinb(n2572), .dout(n12604));
  jand g12359(.dina(n12604), .dinb(asqrt[20] ), .dout(n12605));
  jxor g12360(.dina(n12605), .dinb(n12047), .dout(n12606));
  jnot g12361(.din(n12606), .dout(n12607));
  jand g12362(.dina(n12607), .dinb(n12603), .dout(n12608));
  jor  g12363(.dina(n12608), .dinb(n12602), .dout(n12609));
  jand g12364(.dina(n12609), .dinb(asqrt[47] ), .dout(n12610));
  jor  g12365(.dina(n12609), .dinb(asqrt[47] ), .dout(n12611));
  jxor g12366(.dina(n12049), .dinb(n2345), .dout(n12612));
  jand g12367(.dina(n12612), .dinb(asqrt[20] ), .dout(n12613));
  jxor g12368(.dina(n12613), .dinb(n12054), .dout(n12614));
  jand g12369(.dina(n12614), .dinb(n12611), .dout(n12615));
  jor  g12370(.dina(n12615), .dinb(n12610), .dout(n12616));
  jand g12371(.dina(n12616), .dinb(asqrt[48] ), .dout(n12617));
  jor  g12372(.dina(n12616), .dinb(asqrt[48] ), .dout(n12618));
  jxor g12373(.dina(n12057), .dinb(n2108), .dout(n12619));
  jand g12374(.dina(n12619), .dinb(asqrt[20] ), .dout(n12620));
  jxor g12375(.dina(n12620), .dinb(n12062), .dout(n12621));
  jnot g12376(.din(n12621), .dout(n12622));
  jand g12377(.dina(n12622), .dinb(n12618), .dout(n12623));
  jor  g12378(.dina(n12623), .dinb(n12617), .dout(n12624));
  jand g12379(.dina(n12624), .dinb(asqrt[49] ), .dout(n12625));
  jor  g12380(.dina(n12624), .dinb(asqrt[49] ), .dout(n12626));
  jxor g12381(.dina(n12064), .dinb(n1912), .dout(n12627));
  jand g12382(.dina(n12627), .dinb(asqrt[20] ), .dout(n12628));
  jxor g12383(.dina(n12628), .dinb(n12069), .dout(n12629));
  jnot g12384(.din(n12629), .dout(n12630));
  jand g12385(.dina(n12630), .dinb(n12626), .dout(n12631));
  jor  g12386(.dina(n12631), .dinb(n12625), .dout(n12632));
  jand g12387(.dina(n12632), .dinb(asqrt[50] ), .dout(n12633));
  jor  g12388(.dina(n12632), .dinb(asqrt[50] ), .dout(n12634));
  jxor g12389(.dina(n12071), .dinb(n1699), .dout(n12635));
  jand g12390(.dina(n12635), .dinb(asqrt[20] ), .dout(n12636));
  jxor g12391(.dina(n12636), .dinb(n12076), .dout(n12637));
  jnot g12392(.din(n12637), .dout(n12638));
  jand g12393(.dina(n12638), .dinb(n12634), .dout(n12639));
  jor  g12394(.dina(n12639), .dinb(n12633), .dout(n12640));
  jand g12395(.dina(n12640), .dinb(asqrt[51] ), .dout(n12641));
  jor  g12396(.dina(n12640), .dinb(asqrt[51] ), .dout(n12642));
  jxor g12397(.dina(n12078), .dinb(n1516), .dout(n12643));
  jand g12398(.dina(n12643), .dinb(asqrt[20] ), .dout(n12644));
  jxor g12399(.dina(n12644), .dinb(n12083), .dout(n12645));
  jand g12400(.dina(n12645), .dinb(n12642), .dout(n12646));
  jor  g12401(.dina(n12646), .dinb(n12641), .dout(n12647));
  jand g12402(.dina(n12647), .dinb(asqrt[52] ), .dout(n12648));
  jor  g12403(.dina(n12647), .dinb(asqrt[52] ), .dout(n12649));
  jxor g12404(.dina(n12086), .dinb(n1332), .dout(n12650));
  jand g12405(.dina(n12650), .dinb(asqrt[20] ), .dout(n12651));
  jxor g12406(.dina(n12651), .dinb(n12091), .dout(n12652));
  jnot g12407(.din(n12652), .dout(n12653));
  jand g12408(.dina(n12653), .dinb(n12649), .dout(n12654));
  jor  g12409(.dina(n12654), .dinb(n12648), .dout(n12655));
  jand g12410(.dina(n12655), .dinb(asqrt[53] ), .dout(n12656));
  jor  g12411(.dina(n12655), .dinb(asqrt[53] ), .dout(n12657));
  jxor g12412(.dina(n12093), .dinb(n1173), .dout(n12658));
  jand g12413(.dina(n12658), .dinb(asqrt[20] ), .dout(n12659));
  jxor g12414(.dina(n12659), .dinb(n12098), .dout(n12660));
  jand g12415(.dina(n12660), .dinb(n12657), .dout(n12661));
  jor  g12416(.dina(n12661), .dinb(n12656), .dout(n12662));
  jand g12417(.dina(n12662), .dinb(asqrt[54] ), .dout(n12663));
  jor  g12418(.dina(n12662), .dinb(asqrt[54] ), .dout(n12664));
  jxor g12419(.dina(n12101), .dinb(n1008), .dout(n12665));
  jand g12420(.dina(n12665), .dinb(asqrt[20] ), .dout(n12666));
  jxor g12421(.dina(n12666), .dinb(n12106), .dout(n12667));
  jnot g12422(.din(n12667), .dout(n12668));
  jand g12423(.dina(n12668), .dinb(n12664), .dout(n12669));
  jor  g12424(.dina(n12669), .dinb(n12663), .dout(n12670));
  jand g12425(.dina(n12670), .dinb(asqrt[55] ), .dout(n12671));
  jor  g12426(.dina(n12670), .dinb(asqrt[55] ), .dout(n12672));
  jxor g12427(.dina(n12108), .dinb(n884), .dout(n12673));
  jand g12428(.dina(n12673), .dinb(asqrt[20] ), .dout(n12674));
  jxor g12429(.dina(n12674), .dinb(n12113), .dout(n12675));
  jand g12430(.dina(n12675), .dinb(n12672), .dout(n12676));
  jor  g12431(.dina(n12676), .dinb(n12671), .dout(n12677));
  jand g12432(.dina(n12677), .dinb(asqrt[56] ), .dout(n12678));
  jor  g12433(.dina(n12677), .dinb(asqrt[56] ), .dout(n12679));
  jxor g12434(.dina(n12116), .dinb(n743), .dout(n12680));
  jand g12435(.dina(n12680), .dinb(asqrt[20] ), .dout(n12681));
  jxor g12436(.dina(n12681), .dinb(n12121), .dout(n12682));
  jnot g12437(.din(n12682), .dout(n12683));
  jand g12438(.dina(n12683), .dinb(n12679), .dout(n12684));
  jor  g12439(.dina(n12684), .dinb(n12678), .dout(n12685));
  jand g12440(.dina(n12685), .dinb(asqrt[57] ), .dout(n12686));
  jor  g12441(.dina(n12685), .dinb(asqrt[57] ), .dout(n12687));
  jxor g12442(.dina(n12123), .dinb(n635), .dout(n12688));
  jand g12443(.dina(n12688), .dinb(asqrt[20] ), .dout(n12689));
  jxor g12444(.dina(n12689), .dinb(n12128), .dout(n12690));
  jand g12445(.dina(n12690), .dinb(n12687), .dout(n12691));
  jor  g12446(.dina(n12691), .dinb(n12686), .dout(n12692));
  jand g12447(.dina(n12692), .dinb(asqrt[58] ), .dout(n12693));
  jor  g12448(.dina(n12692), .dinb(asqrt[58] ), .dout(n12694));
  jxor g12449(.dina(n12131), .dinb(n515), .dout(n12695));
  jand g12450(.dina(n12695), .dinb(asqrt[20] ), .dout(n12696));
  jxor g12451(.dina(n12696), .dinb(n12136), .dout(n12697));
  jand g12452(.dina(n12697), .dinb(n12694), .dout(n12698));
  jor  g12453(.dina(n12698), .dinb(n12693), .dout(n12699));
  jand g12454(.dina(n12699), .dinb(asqrt[59] ), .dout(n12700));
  jor  g12455(.dina(n12699), .dinb(asqrt[59] ), .dout(n12701));
  jxor g12456(.dina(n12139), .dinb(n443), .dout(n12702));
  jand g12457(.dina(n12702), .dinb(asqrt[20] ), .dout(n12703));
  jxor g12458(.dina(n12703), .dinb(n12144), .dout(n12704));
  jand g12459(.dina(n12704), .dinb(n12701), .dout(n12705));
  jor  g12460(.dina(n12705), .dinb(n12700), .dout(n12706));
  jand g12461(.dina(n12706), .dinb(asqrt[60] ), .dout(n12707));
  jor  g12462(.dina(n12706), .dinb(asqrt[60] ), .dout(n12708));
  jxor g12463(.dina(n12147), .dinb(n352), .dout(n12709));
  jand g12464(.dina(n12709), .dinb(asqrt[20] ), .dout(n12710));
  jxor g12465(.dina(n12710), .dinb(n12152), .dout(n12711));
  jnot g12466(.din(n12711), .dout(n12712));
  jand g12467(.dina(n12712), .dinb(n12708), .dout(n12713));
  jor  g12468(.dina(n12713), .dinb(n12707), .dout(n12714));
  jand g12469(.dina(n12714), .dinb(asqrt[61] ), .dout(n12715));
  jor  g12470(.dina(n12714), .dinb(asqrt[61] ), .dout(n12716));
  jxor g12471(.dina(n12154), .dinb(n294), .dout(n12717));
  jand g12472(.dina(n12717), .dinb(asqrt[20] ), .dout(n12718));
  jxor g12473(.dina(n12718), .dinb(n12159), .dout(n12719));
  jnot g12474(.din(n12719), .dout(n12720));
  jand g12475(.dina(n12720), .dinb(n12716), .dout(n12721));
  jor  g12476(.dina(n12721), .dinb(n12715), .dout(n12722));
  jand g12477(.dina(n12722), .dinb(asqrt[62] ), .dout(n12723));
  jor  g12478(.dina(n12722), .dinb(asqrt[62] ), .dout(n12724));
  jxor g12479(.dina(n12161), .dinb(n239), .dout(n12725));
  jand g12480(.dina(n12725), .dinb(asqrt[20] ), .dout(n12726));
  jxor g12481(.dina(n12726), .dinb(n12166), .dout(n12727));
  jnot g12482(.din(n12727), .dout(n12728));
  jand g12483(.dina(n12728), .dinb(n12724), .dout(n12729));
  jor  g12484(.dina(n12729), .dinb(n12723), .dout(n12730));
  jor  g12485(.dina(n12730), .dinb(n12195), .dout(n12731));
  jnot g12486(.din(n12731), .dout(n12732));
  jand g12487(.dina(n12408), .dinb(n12176), .dout(n12733));
  jnot g12488(.din(n12733), .dout(n12734));
  jand g12489(.dina(n12180), .dinb(asqrt[63] ), .dout(n12735));
  jand g12490(.dina(n12735), .dinb(n12207), .dout(n12736));
  jand g12491(.dina(n12736), .dinb(n12734), .dout(n12737));
  jand g12492(.dina(n12190), .dinb(n12404), .dout(n12738));
  jnot g12493(.din(n12195), .dout(n12739));
  jnot g12494(.din(n12723), .dout(n12740));
  jnot g12495(.din(n12715), .dout(n12741));
  jnot g12496(.din(n12707), .dout(n12742));
  jnot g12497(.din(n12700), .dout(n12743));
  jnot g12498(.din(n12693), .dout(n12744));
  jnot g12499(.din(n12686), .dout(n12745));
  jnot g12500(.din(n12678), .dout(n12746));
  jnot g12501(.din(n12671), .dout(n12747));
  jnot g12502(.din(n12663), .dout(n12748));
  jnot g12503(.din(n12656), .dout(n12749));
  jnot g12504(.din(n12648), .dout(n12750));
  jnot g12505(.din(n12641), .dout(n12751));
  jnot g12506(.din(n12633), .dout(n12752));
  jnot g12507(.din(n12625), .dout(n12753));
  jnot g12508(.din(n12617), .dout(n12754));
  jnot g12509(.din(n12610), .dout(n12755));
  jnot g12510(.din(n12602), .dout(n12756));
  jnot g12511(.din(n12595), .dout(n12757));
  jnot g12512(.din(n12587), .dout(n12758));
  jnot g12513(.din(n12580), .dout(n12759));
  jnot g12514(.din(n12583), .dout(n12760));
  jnot g12515(.din(n12572), .dout(n12761));
  jnot g12516(.din(n12564), .dout(n12762));
  jnot g12517(.din(n12556), .dout(n12763));
  jnot g12518(.din(n12548), .dout(n12764));
  jnot g12519(.din(n12540), .dout(n12765));
  jnot g12520(.din(n12533), .dout(n12766));
  jnot g12521(.din(n12525), .dout(n12767));
  jnot g12522(.din(n12517), .dout(n12768));
  jnot g12523(.din(n12509), .dout(n12769));
  jnot g12524(.din(n12502), .dout(n12770));
  jnot g12525(.din(n12494), .dout(n12771));
  jnot g12526(.din(n12487), .dout(n12772));
  jnot g12527(.din(n12479), .dout(n12773));
  jnot g12528(.din(n12471), .dout(n12774));
  jnot g12529(.din(n12463), .dout(n12775));
  jnot g12530(.din(n12456), .dout(n12776));
  jnot g12531(.din(n12448), .dout(n12777));
  jnot g12532(.din(n12441), .dout(n12778));
  jnot g12533(.din(n12433), .dout(n12779));
  jnot g12534(.din(n12426), .dout(n12780));
  jnot g12535(.din(n12415), .dout(n12781));
  jnot g12536(.din(n12202), .dout(n12782));
  jnot g12537(.din(n12199), .dout(n12783));
  jor  g12538(.dina(n12410), .dinb(n11864), .dout(n12784));
  jand g12539(.dina(n12784), .dinb(n12783), .dout(n12785));
  jand g12540(.dina(n12785), .dinb(n11858), .dout(n12786));
  jor  g12541(.dina(n12410), .dinb(a[40] ), .dout(n12787));
  jand g12542(.dina(n12787), .dinb(a[41] ), .dout(n12788));
  jor  g12543(.dina(n12417), .dinb(n12788), .dout(n12789));
  jor  g12544(.dina(n12789), .dinb(n12786), .dout(n12790));
  jand g12545(.dina(n12790), .dinb(n12782), .dout(n12791));
  jand g12546(.dina(n12791), .dinb(n11347), .dout(n12792));
  jor  g12547(.dina(n12422), .dinb(n12792), .dout(n12793));
  jand g12548(.dina(n12793), .dinb(n12781), .dout(n12794));
  jand g12549(.dina(n12794), .dinb(n10824), .dout(n12795));
  jnot g12550(.din(n12430), .dout(n12796));
  jor  g12551(.dina(n12796), .dinb(n12795), .dout(n12797));
  jand g12552(.dina(n12797), .dinb(n12780), .dout(n12798));
  jand g12553(.dina(n12798), .dinb(n10328), .dout(n12799));
  jor  g12554(.dina(n12437), .dinb(n12799), .dout(n12800));
  jand g12555(.dina(n12800), .dinb(n12779), .dout(n12801));
  jand g12556(.dina(n12801), .dinb(n9832), .dout(n12802));
  jnot g12557(.din(n12445), .dout(n12803));
  jor  g12558(.dina(n12803), .dinb(n12802), .dout(n12804));
  jand g12559(.dina(n12804), .dinb(n12778), .dout(n12805));
  jand g12560(.dina(n12805), .dinb(n9369), .dout(n12806));
  jor  g12561(.dina(n12452), .dinb(n12806), .dout(n12807));
  jand g12562(.dina(n12807), .dinb(n12777), .dout(n12808));
  jand g12563(.dina(n12808), .dinb(n8890), .dout(n12809));
  jnot g12564(.din(n12460), .dout(n12810));
  jor  g12565(.dina(n12810), .dinb(n12809), .dout(n12811));
  jand g12566(.dina(n12811), .dinb(n12776), .dout(n12812));
  jand g12567(.dina(n12812), .dinb(n8449), .dout(n12813));
  jor  g12568(.dina(n12467), .dinb(n12813), .dout(n12814));
  jand g12569(.dina(n12814), .dinb(n12775), .dout(n12815));
  jand g12570(.dina(n12815), .dinb(n8003), .dout(n12816));
  jor  g12571(.dina(n12475), .dinb(n12816), .dout(n12817));
  jand g12572(.dina(n12817), .dinb(n12774), .dout(n12818));
  jand g12573(.dina(n12818), .dinb(n7581), .dout(n12819));
  jor  g12574(.dina(n12483), .dinb(n12819), .dout(n12820));
  jand g12575(.dina(n12820), .dinb(n12773), .dout(n12821));
  jand g12576(.dina(n12821), .dinb(n7154), .dout(n12822));
  jnot g12577(.din(n12491), .dout(n12823));
  jor  g12578(.dina(n12823), .dinb(n12822), .dout(n12824));
  jand g12579(.dina(n12824), .dinb(n12772), .dout(n12825));
  jand g12580(.dina(n12825), .dinb(n6758), .dout(n12826));
  jor  g12581(.dina(n12498), .dinb(n12826), .dout(n12827));
  jand g12582(.dina(n12827), .dinb(n12771), .dout(n12828));
  jand g12583(.dina(n12828), .dinb(n6357), .dout(n12829));
  jnot g12584(.din(n12506), .dout(n12830));
  jor  g12585(.dina(n12830), .dinb(n12829), .dout(n12831));
  jand g12586(.dina(n12831), .dinb(n12770), .dout(n12832));
  jand g12587(.dina(n12832), .dinb(n5989), .dout(n12833));
  jor  g12588(.dina(n12513), .dinb(n12833), .dout(n12834));
  jand g12589(.dina(n12834), .dinb(n12769), .dout(n12835));
  jand g12590(.dina(n12835), .dinb(n5606), .dout(n12836));
  jor  g12591(.dina(n12521), .dinb(n12836), .dout(n12837));
  jand g12592(.dina(n12837), .dinb(n12768), .dout(n12838));
  jand g12593(.dina(n12838), .dinb(n5259), .dout(n12839));
  jor  g12594(.dina(n12529), .dinb(n12839), .dout(n12840));
  jand g12595(.dina(n12840), .dinb(n12767), .dout(n12841));
  jand g12596(.dina(n12841), .dinb(n4902), .dout(n12842));
  jnot g12597(.din(n12537), .dout(n12843));
  jor  g12598(.dina(n12843), .dinb(n12842), .dout(n12844));
  jand g12599(.dina(n12844), .dinb(n12766), .dout(n12845));
  jand g12600(.dina(n12845), .dinb(n4582), .dout(n12846));
  jor  g12601(.dina(n12544), .dinb(n12846), .dout(n12847));
  jand g12602(.dina(n12847), .dinb(n12765), .dout(n12848));
  jand g12603(.dina(n12848), .dinb(n4249), .dout(n12849));
  jor  g12604(.dina(n12552), .dinb(n12849), .dout(n12850));
  jand g12605(.dina(n12850), .dinb(n12764), .dout(n12851));
  jand g12606(.dina(n12851), .dinb(n3955), .dout(n12852));
  jor  g12607(.dina(n12560), .dinb(n12852), .dout(n12853));
  jand g12608(.dina(n12853), .dinb(n12763), .dout(n12854));
  jand g12609(.dina(n12854), .dinb(n3642), .dout(n12855));
  jor  g12610(.dina(n12568), .dinb(n12855), .dout(n12856));
  jand g12611(.dina(n12856), .dinb(n12762), .dout(n12857));
  jand g12612(.dina(n12857), .dinb(n3368), .dout(n12858));
  jor  g12613(.dina(n12576), .dinb(n12858), .dout(n12859));
  jand g12614(.dina(n12859), .dinb(n12761), .dout(n12860));
  jand g12615(.dina(n12860), .dinb(n3089), .dout(n12861));
  jor  g12616(.dina(n12861), .dinb(n12760), .dout(n12862));
  jand g12617(.dina(n12862), .dinb(n12759), .dout(n12863));
  jand g12618(.dina(n12863), .dinb(n2833), .dout(n12864));
  jor  g12619(.dina(n12591), .dinb(n12864), .dout(n12865));
  jand g12620(.dina(n12865), .dinb(n12758), .dout(n12866));
  jand g12621(.dina(n12866), .dinb(n2572), .dout(n12867));
  jnot g12622(.din(n12599), .dout(n12868));
  jor  g12623(.dina(n12868), .dinb(n12867), .dout(n12869));
  jand g12624(.dina(n12869), .dinb(n12757), .dout(n12870));
  jand g12625(.dina(n12870), .dinb(n2345), .dout(n12871));
  jor  g12626(.dina(n12606), .dinb(n12871), .dout(n12872));
  jand g12627(.dina(n12872), .dinb(n12756), .dout(n12873));
  jand g12628(.dina(n12873), .dinb(n2108), .dout(n12874));
  jnot g12629(.din(n12614), .dout(n12875));
  jor  g12630(.dina(n12875), .dinb(n12874), .dout(n12876));
  jand g12631(.dina(n12876), .dinb(n12755), .dout(n12877));
  jand g12632(.dina(n12877), .dinb(n1912), .dout(n12878));
  jor  g12633(.dina(n12621), .dinb(n12878), .dout(n12879));
  jand g12634(.dina(n12879), .dinb(n12754), .dout(n12880));
  jand g12635(.dina(n12880), .dinb(n1699), .dout(n12881));
  jor  g12636(.dina(n12629), .dinb(n12881), .dout(n12882));
  jand g12637(.dina(n12882), .dinb(n12753), .dout(n12883));
  jand g12638(.dina(n12883), .dinb(n1516), .dout(n12884));
  jor  g12639(.dina(n12637), .dinb(n12884), .dout(n12885));
  jand g12640(.dina(n12885), .dinb(n12752), .dout(n12886));
  jand g12641(.dina(n12886), .dinb(n1332), .dout(n12887));
  jnot g12642(.din(n12645), .dout(n12888));
  jor  g12643(.dina(n12888), .dinb(n12887), .dout(n12889));
  jand g12644(.dina(n12889), .dinb(n12751), .dout(n12890));
  jand g12645(.dina(n12890), .dinb(n1173), .dout(n12891));
  jor  g12646(.dina(n12652), .dinb(n12891), .dout(n12892));
  jand g12647(.dina(n12892), .dinb(n12750), .dout(n12893));
  jand g12648(.dina(n12893), .dinb(n1008), .dout(n12894));
  jnot g12649(.din(n12660), .dout(n12895));
  jor  g12650(.dina(n12895), .dinb(n12894), .dout(n12896));
  jand g12651(.dina(n12896), .dinb(n12749), .dout(n12897));
  jand g12652(.dina(n12897), .dinb(n884), .dout(n12898));
  jor  g12653(.dina(n12667), .dinb(n12898), .dout(n12899));
  jand g12654(.dina(n12899), .dinb(n12748), .dout(n12900));
  jand g12655(.dina(n12900), .dinb(n743), .dout(n12901));
  jnot g12656(.din(n12675), .dout(n12902));
  jor  g12657(.dina(n12902), .dinb(n12901), .dout(n12903));
  jand g12658(.dina(n12903), .dinb(n12747), .dout(n12904));
  jand g12659(.dina(n12904), .dinb(n635), .dout(n12905));
  jor  g12660(.dina(n12682), .dinb(n12905), .dout(n12906));
  jand g12661(.dina(n12906), .dinb(n12746), .dout(n12907));
  jand g12662(.dina(n12907), .dinb(n515), .dout(n12908));
  jnot g12663(.din(n12690), .dout(n12909));
  jor  g12664(.dina(n12909), .dinb(n12908), .dout(n12910));
  jand g12665(.dina(n12910), .dinb(n12745), .dout(n12911));
  jand g12666(.dina(n12911), .dinb(n443), .dout(n12912));
  jnot g12667(.din(n12697), .dout(n12913));
  jor  g12668(.dina(n12913), .dinb(n12912), .dout(n12914));
  jand g12669(.dina(n12914), .dinb(n12744), .dout(n12915));
  jand g12670(.dina(n12915), .dinb(n352), .dout(n12916));
  jnot g12671(.din(n12704), .dout(n12917));
  jor  g12672(.dina(n12917), .dinb(n12916), .dout(n12918));
  jand g12673(.dina(n12918), .dinb(n12743), .dout(n12919));
  jand g12674(.dina(n12919), .dinb(n294), .dout(n12920));
  jor  g12675(.dina(n12711), .dinb(n12920), .dout(n12921));
  jand g12676(.dina(n12921), .dinb(n12742), .dout(n12922));
  jand g12677(.dina(n12922), .dinb(n239), .dout(n12923));
  jor  g12678(.dina(n12719), .dinb(n12923), .dout(n12924));
  jand g12679(.dina(n12924), .dinb(n12741), .dout(n12925));
  jand g12680(.dina(n12925), .dinb(n221), .dout(n12926));
  jor  g12681(.dina(n12727), .dinb(n12926), .dout(n12927));
  jand g12682(.dina(n12927), .dinb(n12740), .dout(n12928));
  jor  g12683(.dina(n12928), .dinb(n12739), .dout(n12929));
  jor  g12684(.dina(n12929), .dinb(n12177), .dout(n12930));
  jor  g12685(.dina(n12930), .dinb(n12738), .dout(n12931));
  jand g12686(.dina(n12931), .dinb(n218), .dout(n12932));
  jand g12687(.dina(n12410), .dinb(n11862), .dout(n12933));
  jor  g12688(.dina(n12933), .dinb(n12932), .dout(n12934));
  jor  g12689(.dina(n12934), .dinb(n12737), .dout(n12935));
  jor  g12690(.dina(n12935), .dinb(n12732), .dout(asqrt[19] ));
  jand g12691(.dina(n12730), .dinb(n12195), .dout(n12937));
  jand g12692(.dina(n12935), .dinb(n12937), .dout(n12938));
  jnot g12693(.din(n12737), .dout(n12939));
  jnot g12694(.din(n12738), .dout(n12940));
  jand g12695(.dina(n12937), .dinb(n12207), .dout(n12941));
  jand g12696(.dina(n12941), .dinb(n12940), .dout(n12942));
  jor  g12697(.dina(n12942), .dinb(asqrt[63] ), .dout(n12943));
  jnot g12698(.din(n12933), .dout(n12944));
  jand g12699(.dina(n12944), .dinb(n12943), .dout(n12945));
  jand g12700(.dina(n12945), .dinb(n12939), .dout(n12946));
  jand g12701(.dina(n12946), .dinb(n12731), .dout(n12947));
  jxor g12702(.dina(n12722), .dinb(n221), .dout(n12948));
  jor  g12703(.dina(n12948), .dinb(n12947), .dout(n12949));
  jxor g12704(.dina(n12949), .dinb(n12727), .dout(n12950));
  jnot g12705(.din(n12950), .dout(n12951));
  jor  g12706(.dina(n12947), .dinb(n12196), .dout(n12952));
  jnot g12707(.din(a[36] ), .dout(n12953));
  jnot g12708(.din(a[37] ), .dout(n12954));
  jand g12709(.dina(n12954), .dinb(n12953), .dout(n12955));
  jand g12710(.dina(n12955), .dinb(n12196), .dout(n12956));
  jnot g12711(.din(n12956), .dout(n12957));
  jand g12712(.dina(n12957), .dinb(n12952), .dout(n12958));
  jor  g12713(.dina(n12958), .dinb(n12410), .dout(n12959));
  jand g12714(.dina(n12958), .dinb(n12410), .dout(n12960));
  jor  g12715(.dina(n12947), .dinb(a[38] ), .dout(n12961));
  jand g12716(.dina(n12961), .dinb(a[39] ), .dout(n12962));
  jand g12717(.dina(asqrt[19] ), .dinb(n12198), .dout(n12963));
  jor  g12718(.dina(n12963), .dinb(n12962), .dout(n12964));
  jor  g12719(.dina(n12964), .dinb(n12960), .dout(n12965));
  jand g12720(.dina(n12965), .dinb(n12959), .dout(n12966));
  jor  g12721(.dina(n12966), .dinb(n11858), .dout(n12967));
  jand g12722(.dina(n12966), .dinb(n11858), .dout(n12968));
  jnot g12723(.din(n12198), .dout(n12969));
  jor  g12724(.dina(n12947), .dinb(n12969), .dout(n12970));
  jor  g12725(.dina(n12732), .dinb(n12410), .dout(n12971));
  jor  g12726(.dina(n12971), .dinb(n12736), .dout(n12972));
  jor  g12727(.dina(n12972), .dinb(n12932), .dout(n12973));
  jand g12728(.dina(n12973), .dinb(n12970), .dout(n12974));
  jxor g12729(.dina(n12974), .dinb(n11864), .dout(n12975));
  jor  g12730(.dina(n12975), .dinb(n12968), .dout(n12976));
  jand g12731(.dina(n12976), .dinb(n12967), .dout(n12977));
  jor  g12732(.dina(n12977), .dinb(n11347), .dout(n12978));
  jand g12733(.dina(n12977), .dinb(n11347), .dout(n12979));
  jxor g12734(.dina(n12201), .dinb(n11858), .dout(n12980));
  jor  g12735(.dina(n12980), .dinb(n12947), .dout(n12981));
  jxor g12736(.dina(n12981), .dinb(n12789), .dout(n12982));
  jnot g12737(.din(n12982), .dout(n12983));
  jor  g12738(.dina(n12983), .dinb(n12979), .dout(n12984));
  jand g12739(.dina(n12984), .dinb(n12978), .dout(n12985));
  jor  g12740(.dina(n12985), .dinb(n10824), .dout(n12986));
  jand g12741(.dina(n12985), .dinb(n10824), .dout(n12987));
  jxor g12742(.dina(n12414), .dinb(n11347), .dout(n12988));
  jor  g12743(.dina(n12988), .dinb(n12947), .dout(n12989));
  jxor g12744(.dina(n12989), .dinb(n12423), .dout(n12990));
  jor  g12745(.dina(n12990), .dinb(n12987), .dout(n12991));
  jand g12746(.dina(n12991), .dinb(n12986), .dout(n12992));
  jor  g12747(.dina(n12992), .dinb(n10328), .dout(n12993));
  jand g12748(.dina(n12992), .dinb(n10328), .dout(n12994));
  jxor g12749(.dina(n12425), .dinb(n10824), .dout(n12995));
  jor  g12750(.dina(n12995), .dinb(n12947), .dout(n12996));
  jxor g12751(.dina(n12996), .dinb(n12796), .dout(n12997));
  jnot g12752(.din(n12997), .dout(n12998));
  jor  g12753(.dina(n12998), .dinb(n12994), .dout(n12999));
  jand g12754(.dina(n12999), .dinb(n12993), .dout(n13000));
  jor  g12755(.dina(n13000), .dinb(n9832), .dout(n13001));
  jand g12756(.dina(n13000), .dinb(n9832), .dout(n13002));
  jxor g12757(.dina(n12432), .dinb(n10328), .dout(n13003));
  jor  g12758(.dina(n13003), .dinb(n12947), .dout(n13004));
  jxor g12759(.dina(n13004), .dinb(n12438), .dout(n13005));
  jor  g12760(.dina(n13005), .dinb(n13002), .dout(n13006));
  jand g12761(.dina(n13006), .dinb(n13001), .dout(n13007));
  jor  g12762(.dina(n13007), .dinb(n9369), .dout(n13008));
  jand g12763(.dina(n13007), .dinb(n9369), .dout(n13009));
  jxor g12764(.dina(n12440), .dinb(n9832), .dout(n13010));
  jor  g12765(.dina(n13010), .dinb(n12947), .dout(n13011));
  jxor g12766(.dina(n13011), .dinb(n12803), .dout(n13012));
  jnot g12767(.din(n13012), .dout(n13013));
  jor  g12768(.dina(n13013), .dinb(n13009), .dout(n13014));
  jand g12769(.dina(n13014), .dinb(n13008), .dout(n13015));
  jor  g12770(.dina(n13015), .dinb(n8890), .dout(n13016));
  jand g12771(.dina(n13015), .dinb(n8890), .dout(n13017));
  jxor g12772(.dina(n12447), .dinb(n9369), .dout(n13018));
  jor  g12773(.dina(n13018), .dinb(n12947), .dout(n13019));
  jxor g12774(.dina(n13019), .dinb(n12453), .dout(n13020));
  jor  g12775(.dina(n13020), .dinb(n13017), .dout(n13021));
  jand g12776(.dina(n13021), .dinb(n13016), .dout(n13022));
  jor  g12777(.dina(n13022), .dinb(n8449), .dout(n13023));
  jand g12778(.dina(n13022), .dinb(n8449), .dout(n13024));
  jxor g12779(.dina(n12455), .dinb(n8890), .dout(n13025));
  jor  g12780(.dina(n13025), .dinb(n12947), .dout(n13026));
  jxor g12781(.dina(n13026), .dinb(n12810), .dout(n13027));
  jnot g12782(.din(n13027), .dout(n13028));
  jor  g12783(.dina(n13028), .dinb(n13024), .dout(n13029));
  jand g12784(.dina(n13029), .dinb(n13023), .dout(n13030));
  jor  g12785(.dina(n13030), .dinb(n8003), .dout(n13031));
  jand g12786(.dina(n13030), .dinb(n8003), .dout(n13032));
  jxor g12787(.dina(n12462), .dinb(n8449), .dout(n13033));
  jor  g12788(.dina(n13033), .dinb(n12947), .dout(n13034));
  jxor g12789(.dina(n13034), .dinb(n12468), .dout(n13035));
  jor  g12790(.dina(n13035), .dinb(n13032), .dout(n13036));
  jand g12791(.dina(n13036), .dinb(n13031), .dout(n13037));
  jor  g12792(.dina(n13037), .dinb(n7581), .dout(n13038));
  jand g12793(.dina(n13037), .dinb(n7581), .dout(n13039));
  jxor g12794(.dina(n12470), .dinb(n8003), .dout(n13040));
  jor  g12795(.dina(n13040), .dinb(n12947), .dout(n13041));
  jxor g12796(.dina(n13041), .dinb(n12476), .dout(n13042));
  jor  g12797(.dina(n13042), .dinb(n13039), .dout(n13043));
  jand g12798(.dina(n13043), .dinb(n13038), .dout(n13044));
  jor  g12799(.dina(n13044), .dinb(n7154), .dout(n13045));
  jand g12800(.dina(n13044), .dinb(n7154), .dout(n13046));
  jxor g12801(.dina(n12478), .dinb(n7581), .dout(n13047));
  jor  g12802(.dina(n13047), .dinb(n12947), .dout(n13048));
  jxor g12803(.dina(n13048), .dinb(n12484), .dout(n13049));
  jor  g12804(.dina(n13049), .dinb(n13046), .dout(n13050));
  jand g12805(.dina(n13050), .dinb(n13045), .dout(n13051));
  jor  g12806(.dina(n13051), .dinb(n6758), .dout(n13052));
  jand g12807(.dina(n13051), .dinb(n6758), .dout(n13053));
  jxor g12808(.dina(n12486), .dinb(n7154), .dout(n13054));
  jor  g12809(.dina(n13054), .dinb(n12947), .dout(n13055));
  jxor g12810(.dina(n13055), .dinb(n12823), .dout(n13056));
  jnot g12811(.din(n13056), .dout(n13057));
  jor  g12812(.dina(n13057), .dinb(n13053), .dout(n13058));
  jand g12813(.dina(n13058), .dinb(n13052), .dout(n13059));
  jor  g12814(.dina(n13059), .dinb(n6357), .dout(n13060));
  jand g12815(.dina(n13059), .dinb(n6357), .dout(n13061));
  jxor g12816(.dina(n12493), .dinb(n6758), .dout(n13062));
  jor  g12817(.dina(n13062), .dinb(n12947), .dout(n13063));
  jxor g12818(.dina(n13063), .dinb(n12499), .dout(n13064));
  jor  g12819(.dina(n13064), .dinb(n13061), .dout(n13065));
  jand g12820(.dina(n13065), .dinb(n13060), .dout(n13066));
  jor  g12821(.dina(n13066), .dinb(n5989), .dout(n13067));
  jand g12822(.dina(n13066), .dinb(n5989), .dout(n13068));
  jxor g12823(.dina(n12501), .dinb(n6357), .dout(n13069));
  jor  g12824(.dina(n13069), .dinb(n12947), .dout(n13070));
  jxor g12825(.dina(n13070), .dinb(n12830), .dout(n13071));
  jnot g12826(.din(n13071), .dout(n13072));
  jor  g12827(.dina(n13072), .dinb(n13068), .dout(n13073));
  jand g12828(.dina(n13073), .dinb(n13067), .dout(n13074));
  jor  g12829(.dina(n13074), .dinb(n5606), .dout(n13075));
  jand g12830(.dina(n13074), .dinb(n5606), .dout(n13076));
  jxor g12831(.dina(n12508), .dinb(n5989), .dout(n13077));
  jor  g12832(.dina(n13077), .dinb(n12947), .dout(n13078));
  jxor g12833(.dina(n13078), .dinb(n12514), .dout(n13079));
  jor  g12834(.dina(n13079), .dinb(n13076), .dout(n13080));
  jand g12835(.dina(n13080), .dinb(n13075), .dout(n13081));
  jor  g12836(.dina(n13081), .dinb(n5259), .dout(n13082));
  jand g12837(.dina(n13081), .dinb(n5259), .dout(n13083));
  jxor g12838(.dina(n12516), .dinb(n5606), .dout(n13084));
  jor  g12839(.dina(n13084), .dinb(n12947), .dout(n13085));
  jxor g12840(.dina(n13085), .dinb(n12522), .dout(n13086));
  jor  g12841(.dina(n13086), .dinb(n13083), .dout(n13087));
  jand g12842(.dina(n13087), .dinb(n13082), .dout(n13088));
  jor  g12843(.dina(n13088), .dinb(n4902), .dout(n13089));
  jand g12844(.dina(n13088), .dinb(n4902), .dout(n13090));
  jxor g12845(.dina(n12524), .dinb(n5259), .dout(n13091));
  jor  g12846(.dina(n13091), .dinb(n12947), .dout(n13092));
  jxor g12847(.dina(n13092), .dinb(n12530), .dout(n13093));
  jor  g12848(.dina(n13093), .dinb(n13090), .dout(n13094));
  jand g12849(.dina(n13094), .dinb(n13089), .dout(n13095));
  jor  g12850(.dina(n13095), .dinb(n4582), .dout(n13096));
  jand g12851(.dina(n13095), .dinb(n4582), .dout(n13097));
  jxor g12852(.dina(n12532), .dinb(n4902), .dout(n13098));
  jor  g12853(.dina(n13098), .dinb(n12947), .dout(n13099));
  jxor g12854(.dina(n13099), .dinb(n12843), .dout(n13100));
  jnot g12855(.din(n13100), .dout(n13101));
  jor  g12856(.dina(n13101), .dinb(n13097), .dout(n13102));
  jand g12857(.dina(n13102), .dinb(n13096), .dout(n13103));
  jor  g12858(.dina(n13103), .dinb(n4249), .dout(n13104));
  jand g12859(.dina(n13103), .dinb(n4249), .dout(n13105));
  jxor g12860(.dina(n12539), .dinb(n4582), .dout(n13106));
  jor  g12861(.dina(n13106), .dinb(n12947), .dout(n13107));
  jxor g12862(.dina(n13107), .dinb(n12545), .dout(n13108));
  jor  g12863(.dina(n13108), .dinb(n13105), .dout(n13109));
  jand g12864(.dina(n13109), .dinb(n13104), .dout(n13110));
  jor  g12865(.dina(n13110), .dinb(n3955), .dout(n13111));
  jand g12866(.dina(n13110), .dinb(n3955), .dout(n13112));
  jxor g12867(.dina(n12547), .dinb(n4249), .dout(n13113));
  jor  g12868(.dina(n13113), .dinb(n12947), .dout(n13114));
  jxor g12869(.dina(n13114), .dinb(n12553), .dout(n13115));
  jor  g12870(.dina(n13115), .dinb(n13112), .dout(n13116));
  jand g12871(.dina(n13116), .dinb(n13111), .dout(n13117));
  jor  g12872(.dina(n13117), .dinb(n3642), .dout(n13118));
  jand g12873(.dina(n13117), .dinb(n3642), .dout(n13119));
  jxor g12874(.dina(n12555), .dinb(n3955), .dout(n13120));
  jor  g12875(.dina(n13120), .dinb(n12947), .dout(n13121));
  jxor g12876(.dina(n13121), .dinb(n12561), .dout(n13122));
  jor  g12877(.dina(n13122), .dinb(n13119), .dout(n13123));
  jand g12878(.dina(n13123), .dinb(n13118), .dout(n13124));
  jor  g12879(.dina(n13124), .dinb(n3368), .dout(n13125));
  jand g12880(.dina(n13124), .dinb(n3368), .dout(n13126));
  jxor g12881(.dina(n12563), .dinb(n3642), .dout(n13127));
  jor  g12882(.dina(n13127), .dinb(n12947), .dout(n13128));
  jxor g12883(.dina(n13128), .dinb(n12569), .dout(n13129));
  jor  g12884(.dina(n13129), .dinb(n13126), .dout(n13130));
  jand g12885(.dina(n13130), .dinb(n13125), .dout(n13131));
  jor  g12886(.dina(n13131), .dinb(n3089), .dout(n13132));
  jand g12887(.dina(n13131), .dinb(n3089), .dout(n13133));
  jxor g12888(.dina(n12571), .dinb(n3368), .dout(n13134));
  jor  g12889(.dina(n13134), .dinb(n12947), .dout(n13135));
  jxor g12890(.dina(n13135), .dinb(n12576), .dout(n13136));
  jnot g12891(.din(n13136), .dout(n13137));
  jor  g12892(.dina(n13137), .dinb(n13133), .dout(n13138));
  jand g12893(.dina(n13138), .dinb(n13132), .dout(n13139));
  jor  g12894(.dina(n13139), .dinb(n2833), .dout(n13140));
  jxor g12895(.dina(n12579), .dinb(n3089), .dout(n13141));
  jor  g12896(.dina(n13141), .dinb(n12947), .dout(n13142));
  jxor g12897(.dina(n13142), .dinb(n12760), .dout(n13143));
  jnot g12898(.din(n13143), .dout(n13144));
  jand g12899(.dina(n13139), .dinb(n2833), .dout(n13145));
  jor  g12900(.dina(n13145), .dinb(n13144), .dout(n13146));
  jand g12901(.dina(n13146), .dinb(n13140), .dout(n13147));
  jor  g12902(.dina(n13147), .dinb(n2572), .dout(n13148));
  jand g12903(.dina(n13147), .dinb(n2572), .dout(n13149));
  jxor g12904(.dina(n12586), .dinb(n2833), .dout(n13150));
  jor  g12905(.dina(n13150), .dinb(n12947), .dout(n13151));
  jxor g12906(.dina(n13151), .dinb(n12592), .dout(n13152));
  jor  g12907(.dina(n13152), .dinb(n13149), .dout(n13153));
  jand g12908(.dina(n13153), .dinb(n13148), .dout(n13154));
  jor  g12909(.dina(n13154), .dinb(n2345), .dout(n13155));
  jand g12910(.dina(n13154), .dinb(n2345), .dout(n13156));
  jxor g12911(.dina(n12594), .dinb(n2572), .dout(n13157));
  jor  g12912(.dina(n13157), .dinb(n12947), .dout(n13158));
  jxor g12913(.dina(n13158), .dinb(n12868), .dout(n13159));
  jnot g12914(.din(n13159), .dout(n13160));
  jor  g12915(.dina(n13160), .dinb(n13156), .dout(n13161));
  jand g12916(.dina(n13161), .dinb(n13155), .dout(n13162));
  jor  g12917(.dina(n13162), .dinb(n2108), .dout(n13163));
  jand g12918(.dina(n13162), .dinb(n2108), .dout(n13164));
  jxor g12919(.dina(n12601), .dinb(n2345), .dout(n13165));
  jor  g12920(.dina(n13165), .dinb(n12947), .dout(n13166));
  jxor g12921(.dina(n13166), .dinb(n12607), .dout(n13167));
  jor  g12922(.dina(n13167), .dinb(n13164), .dout(n13168));
  jand g12923(.dina(n13168), .dinb(n13163), .dout(n13169));
  jor  g12924(.dina(n13169), .dinb(n1912), .dout(n13170));
  jand g12925(.dina(n13169), .dinb(n1912), .dout(n13171));
  jxor g12926(.dina(n12609), .dinb(n2108), .dout(n13172));
  jor  g12927(.dina(n13172), .dinb(n12947), .dout(n13173));
  jxor g12928(.dina(n13173), .dinb(n12875), .dout(n13174));
  jnot g12929(.din(n13174), .dout(n13175));
  jor  g12930(.dina(n13175), .dinb(n13171), .dout(n13176));
  jand g12931(.dina(n13176), .dinb(n13170), .dout(n13177));
  jor  g12932(.dina(n13177), .dinb(n1699), .dout(n13178));
  jand g12933(.dina(n13177), .dinb(n1699), .dout(n13179));
  jxor g12934(.dina(n12616), .dinb(n1912), .dout(n13180));
  jor  g12935(.dina(n13180), .dinb(n12947), .dout(n13181));
  jxor g12936(.dina(n13181), .dinb(n12622), .dout(n13182));
  jor  g12937(.dina(n13182), .dinb(n13179), .dout(n13183));
  jand g12938(.dina(n13183), .dinb(n13178), .dout(n13184));
  jor  g12939(.dina(n13184), .dinb(n1516), .dout(n13185));
  jand g12940(.dina(n13184), .dinb(n1516), .dout(n13186));
  jxor g12941(.dina(n12624), .dinb(n1699), .dout(n13187));
  jor  g12942(.dina(n13187), .dinb(n12947), .dout(n13188));
  jxor g12943(.dina(n13188), .dinb(n12630), .dout(n13189));
  jor  g12944(.dina(n13189), .dinb(n13186), .dout(n13190));
  jand g12945(.dina(n13190), .dinb(n13185), .dout(n13191));
  jor  g12946(.dina(n13191), .dinb(n1332), .dout(n13192));
  jand g12947(.dina(n13191), .dinb(n1332), .dout(n13193));
  jxor g12948(.dina(n12632), .dinb(n1516), .dout(n13194));
  jor  g12949(.dina(n13194), .dinb(n12947), .dout(n13195));
  jxor g12950(.dina(n13195), .dinb(n12638), .dout(n13196));
  jor  g12951(.dina(n13196), .dinb(n13193), .dout(n13197));
  jand g12952(.dina(n13197), .dinb(n13192), .dout(n13198));
  jor  g12953(.dina(n13198), .dinb(n1173), .dout(n13199));
  jand g12954(.dina(n13198), .dinb(n1173), .dout(n13200));
  jxor g12955(.dina(n12640), .dinb(n1332), .dout(n13201));
  jor  g12956(.dina(n13201), .dinb(n12947), .dout(n13202));
  jxor g12957(.dina(n13202), .dinb(n12888), .dout(n13203));
  jnot g12958(.din(n13203), .dout(n13204));
  jor  g12959(.dina(n13204), .dinb(n13200), .dout(n13205));
  jand g12960(.dina(n13205), .dinb(n13199), .dout(n13206));
  jor  g12961(.dina(n13206), .dinb(n1008), .dout(n13207));
  jand g12962(.dina(n13206), .dinb(n1008), .dout(n13208));
  jxor g12963(.dina(n12647), .dinb(n1173), .dout(n13209));
  jor  g12964(.dina(n13209), .dinb(n12947), .dout(n13210));
  jxor g12965(.dina(n13210), .dinb(n12653), .dout(n13211));
  jor  g12966(.dina(n13211), .dinb(n13208), .dout(n13212));
  jand g12967(.dina(n13212), .dinb(n13207), .dout(n13213));
  jor  g12968(.dina(n13213), .dinb(n884), .dout(n13214));
  jand g12969(.dina(n13213), .dinb(n884), .dout(n13215));
  jxor g12970(.dina(n12655), .dinb(n1008), .dout(n13216));
  jor  g12971(.dina(n13216), .dinb(n12947), .dout(n13217));
  jxor g12972(.dina(n13217), .dinb(n12895), .dout(n13218));
  jnot g12973(.din(n13218), .dout(n13219));
  jor  g12974(.dina(n13219), .dinb(n13215), .dout(n13220));
  jand g12975(.dina(n13220), .dinb(n13214), .dout(n13221));
  jor  g12976(.dina(n13221), .dinb(n743), .dout(n13222));
  jand g12977(.dina(n13221), .dinb(n743), .dout(n13223));
  jxor g12978(.dina(n12662), .dinb(n884), .dout(n13224));
  jor  g12979(.dina(n13224), .dinb(n12947), .dout(n13225));
  jxor g12980(.dina(n13225), .dinb(n12668), .dout(n13226));
  jor  g12981(.dina(n13226), .dinb(n13223), .dout(n13227));
  jand g12982(.dina(n13227), .dinb(n13222), .dout(n13228));
  jor  g12983(.dina(n13228), .dinb(n635), .dout(n13229));
  jand g12984(.dina(n13228), .dinb(n635), .dout(n13230));
  jxor g12985(.dina(n12670), .dinb(n743), .dout(n13231));
  jor  g12986(.dina(n13231), .dinb(n12947), .dout(n13232));
  jxor g12987(.dina(n13232), .dinb(n12902), .dout(n13233));
  jnot g12988(.din(n13233), .dout(n13234));
  jor  g12989(.dina(n13234), .dinb(n13230), .dout(n13235));
  jand g12990(.dina(n13235), .dinb(n13229), .dout(n13236));
  jor  g12991(.dina(n13236), .dinb(n515), .dout(n13237));
  jand g12992(.dina(n13236), .dinb(n515), .dout(n13238));
  jxor g12993(.dina(n12677), .dinb(n635), .dout(n13239));
  jor  g12994(.dina(n13239), .dinb(n12947), .dout(n13240));
  jxor g12995(.dina(n13240), .dinb(n12683), .dout(n13241));
  jor  g12996(.dina(n13241), .dinb(n13238), .dout(n13242));
  jand g12997(.dina(n13242), .dinb(n13237), .dout(n13243));
  jor  g12998(.dina(n13243), .dinb(n443), .dout(n13244));
  jand g12999(.dina(n13243), .dinb(n443), .dout(n13245));
  jxor g13000(.dina(n12685), .dinb(n515), .dout(n13246));
  jor  g13001(.dina(n13246), .dinb(n12947), .dout(n13247));
  jxor g13002(.dina(n13247), .dinb(n12909), .dout(n13248));
  jnot g13003(.din(n13248), .dout(n13249));
  jor  g13004(.dina(n13249), .dinb(n13245), .dout(n13250));
  jand g13005(.dina(n13250), .dinb(n13244), .dout(n13251));
  jor  g13006(.dina(n13251), .dinb(n352), .dout(n13252));
  jand g13007(.dina(n13251), .dinb(n352), .dout(n13253));
  jxor g13008(.dina(n12692), .dinb(n443), .dout(n13254));
  jor  g13009(.dina(n13254), .dinb(n12947), .dout(n13255));
  jxor g13010(.dina(n13255), .dinb(n12913), .dout(n13256));
  jnot g13011(.din(n13256), .dout(n13257));
  jor  g13012(.dina(n13257), .dinb(n13253), .dout(n13258));
  jand g13013(.dina(n13258), .dinb(n13252), .dout(n13259));
  jor  g13014(.dina(n13259), .dinb(n294), .dout(n13260));
  jand g13015(.dina(n13259), .dinb(n294), .dout(n13261));
  jxor g13016(.dina(n12699), .dinb(n352), .dout(n13262));
  jor  g13017(.dina(n13262), .dinb(n12947), .dout(n13263));
  jxor g13018(.dina(n13263), .dinb(n12917), .dout(n13264));
  jnot g13019(.din(n13264), .dout(n13265));
  jor  g13020(.dina(n13265), .dinb(n13261), .dout(n13266));
  jand g13021(.dina(n13266), .dinb(n13260), .dout(n13267));
  jor  g13022(.dina(n13267), .dinb(n239), .dout(n13268));
  jand g13023(.dina(n13267), .dinb(n239), .dout(n13269));
  jxor g13024(.dina(n12706), .dinb(n294), .dout(n13270));
  jor  g13025(.dina(n13270), .dinb(n12947), .dout(n13271));
  jxor g13026(.dina(n13271), .dinb(n12712), .dout(n13272));
  jor  g13027(.dina(n13272), .dinb(n13269), .dout(n13273));
  jand g13028(.dina(n13273), .dinb(n13268), .dout(n13274));
  jor  g13029(.dina(n13274), .dinb(n221), .dout(n13275));
  jand g13030(.dina(n13274), .dinb(n221), .dout(n13276));
  jxor g13031(.dina(n12714), .dinb(n239), .dout(n13277));
  jor  g13032(.dina(n13277), .dinb(n12947), .dout(n13278));
  jxor g13033(.dina(n13278), .dinb(n12720), .dout(n13279));
  jor  g13034(.dina(n13279), .dinb(n13276), .dout(n13280));
  jand g13035(.dina(n13280), .dinb(n13275), .dout(n13281));
  jor  g13036(.dina(n13281), .dinb(n12951), .dout(n13282));
  jor  g13037(.dina(n13282), .dinb(n12732), .dout(n13283));
  jor  g13038(.dina(n13283), .dinb(n12938), .dout(n13284));
  jand g13039(.dina(n13284), .dinb(n218), .dout(n13285));
  jand g13040(.dina(n12947), .dinb(n12739), .dout(n13286));
  jand g13041(.dina(n13281), .dinb(n12951), .dout(n13287));
  jor  g13042(.dina(n13287), .dinb(n13286), .dout(n13288));
  jand g13043(.dina(n12946), .dinb(n12928), .dout(n13289));
  jnot g13044(.din(n13289), .dout(n13290));
  jand g13045(.dina(n12929), .dinb(asqrt[63] ), .dout(n13291));
  jand g13046(.dina(n13291), .dinb(n12731), .dout(n13292));
  jand g13047(.dina(n13292), .dinb(n13290), .dout(n13293));
  jor  g13048(.dina(n13293), .dinb(n13288), .dout(n13294));
  jor  g13049(.dina(n13294), .dinb(n13285), .dout(asqrt[18] ));
  jnot g13050(.din(a[34] ), .dout(n13296));
  jnot g13051(.din(a[35] ), .dout(n13297));
  jand g13052(.dina(n13297), .dinb(n13296), .dout(n13298));
  jand g13053(.dina(n13298), .dinb(n12953), .dout(n13299));
  jand g13054(.dina(asqrt[18] ), .dinb(a[36] ), .dout(n13300));
  jor  g13055(.dina(n13300), .dinb(n13299), .dout(n13301));
  jand g13056(.dina(n13301), .dinb(asqrt[19] ), .dout(n13302));
  jor  g13057(.dina(n13301), .dinb(asqrt[19] ), .dout(n13303));
  jand g13058(.dina(asqrt[18] ), .dinb(n12953), .dout(n13304));
  jor  g13059(.dina(n13304), .dinb(n12954), .dout(n13305));
  jnot g13060(.din(n12955), .dout(n13306));
  jnot g13061(.din(n12938), .dout(n13307));
  jnot g13062(.din(n13275), .dout(n13308));
  jnot g13063(.din(n13268), .dout(n13309));
  jnot g13064(.din(n13260), .dout(n13310));
  jnot g13065(.din(n13252), .dout(n13311));
  jnot g13066(.din(n13244), .dout(n13312));
  jnot g13067(.din(n13237), .dout(n13313));
  jnot g13068(.din(n13229), .dout(n13314));
  jnot g13069(.din(n13222), .dout(n13315));
  jnot g13070(.din(n13214), .dout(n13316));
  jnot g13071(.din(n13207), .dout(n13317));
  jnot g13072(.din(n13199), .dout(n13318));
  jnot g13073(.din(n13192), .dout(n13319));
  jnot g13074(.din(n13185), .dout(n13320));
  jnot g13075(.din(n13178), .dout(n13321));
  jnot g13076(.din(n13170), .dout(n13322));
  jnot g13077(.din(n13163), .dout(n13323));
  jnot g13078(.din(n13155), .dout(n13324));
  jnot g13079(.din(n13148), .dout(n13325));
  jnot g13080(.din(n13140), .dout(n13326));
  jnot g13081(.din(n13132), .dout(n13327));
  jnot g13082(.din(n13125), .dout(n13328));
  jnot g13083(.din(n13118), .dout(n13329));
  jnot g13084(.din(n13111), .dout(n13330));
  jnot g13085(.din(n13104), .dout(n13331));
  jnot g13086(.din(n13096), .dout(n13332));
  jnot g13087(.din(n13089), .dout(n13333));
  jnot g13088(.din(n13082), .dout(n13334));
  jnot g13089(.din(n13075), .dout(n13335));
  jnot g13090(.din(n13067), .dout(n13336));
  jnot g13091(.din(n13060), .dout(n13337));
  jnot g13092(.din(n13052), .dout(n13338));
  jnot g13093(.din(n13045), .dout(n13339));
  jnot g13094(.din(n13038), .dout(n13340));
  jnot g13095(.din(n13031), .dout(n13341));
  jnot g13096(.din(n13023), .dout(n13342));
  jnot g13097(.din(n13016), .dout(n13343));
  jnot g13098(.din(n13008), .dout(n13344));
  jnot g13099(.din(n13001), .dout(n13345));
  jnot g13100(.din(n12993), .dout(n13346));
  jnot g13101(.din(n12986), .dout(n13347));
  jnot g13102(.din(n12978), .dout(n13348));
  jnot g13103(.din(n12967), .dout(n13349));
  jnot g13104(.din(n12959), .dout(n13350));
  jand g13105(.dina(asqrt[19] ), .dinb(a[38] ), .dout(n13351));
  jor  g13106(.dina(n12956), .dinb(n13351), .dout(n13352));
  jor  g13107(.dina(n13352), .dinb(asqrt[20] ), .dout(n13353));
  jand g13108(.dina(asqrt[19] ), .dinb(n12196), .dout(n13354));
  jor  g13109(.dina(n13354), .dinb(n12197), .dout(n13355));
  jand g13110(.dina(n12970), .dinb(n13355), .dout(n13356));
  jand g13111(.dina(n13356), .dinb(n13353), .dout(n13357));
  jor  g13112(.dina(n13357), .dinb(n13350), .dout(n13358));
  jor  g13113(.dina(n13358), .dinb(asqrt[21] ), .dout(n13359));
  jnot g13114(.din(n12975), .dout(n13360));
  jand g13115(.dina(n13360), .dinb(n13359), .dout(n13361));
  jor  g13116(.dina(n13361), .dinb(n13349), .dout(n13362));
  jor  g13117(.dina(n13362), .dinb(asqrt[22] ), .dout(n13363));
  jand g13118(.dina(n12982), .dinb(n13363), .dout(n13364));
  jor  g13119(.dina(n13364), .dinb(n13348), .dout(n13365));
  jor  g13120(.dina(n13365), .dinb(asqrt[23] ), .dout(n13366));
  jnot g13121(.din(n12990), .dout(n13367));
  jand g13122(.dina(n13367), .dinb(n13366), .dout(n13368));
  jor  g13123(.dina(n13368), .dinb(n13347), .dout(n13369));
  jor  g13124(.dina(n13369), .dinb(asqrt[24] ), .dout(n13370));
  jand g13125(.dina(n12997), .dinb(n13370), .dout(n13371));
  jor  g13126(.dina(n13371), .dinb(n13346), .dout(n13372));
  jor  g13127(.dina(n13372), .dinb(asqrt[25] ), .dout(n13373));
  jnot g13128(.din(n13005), .dout(n13374));
  jand g13129(.dina(n13374), .dinb(n13373), .dout(n13375));
  jor  g13130(.dina(n13375), .dinb(n13345), .dout(n13376));
  jor  g13131(.dina(n13376), .dinb(asqrt[26] ), .dout(n13377));
  jand g13132(.dina(n13012), .dinb(n13377), .dout(n13378));
  jor  g13133(.dina(n13378), .dinb(n13344), .dout(n13379));
  jor  g13134(.dina(n13379), .dinb(asqrt[27] ), .dout(n13380));
  jnot g13135(.din(n13020), .dout(n13381));
  jand g13136(.dina(n13381), .dinb(n13380), .dout(n13382));
  jor  g13137(.dina(n13382), .dinb(n13343), .dout(n13383));
  jor  g13138(.dina(n13383), .dinb(asqrt[28] ), .dout(n13384));
  jand g13139(.dina(n13027), .dinb(n13384), .dout(n13385));
  jor  g13140(.dina(n13385), .dinb(n13342), .dout(n13386));
  jor  g13141(.dina(n13386), .dinb(asqrt[29] ), .dout(n13387));
  jnot g13142(.din(n13035), .dout(n13388));
  jand g13143(.dina(n13388), .dinb(n13387), .dout(n13389));
  jor  g13144(.dina(n13389), .dinb(n13341), .dout(n13390));
  jor  g13145(.dina(n13390), .dinb(asqrt[30] ), .dout(n13391));
  jnot g13146(.din(n13042), .dout(n13392));
  jand g13147(.dina(n13392), .dinb(n13391), .dout(n13393));
  jor  g13148(.dina(n13393), .dinb(n13340), .dout(n13394));
  jor  g13149(.dina(n13394), .dinb(asqrt[31] ), .dout(n13395));
  jnot g13150(.din(n13049), .dout(n13396));
  jand g13151(.dina(n13396), .dinb(n13395), .dout(n13397));
  jor  g13152(.dina(n13397), .dinb(n13339), .dout(n13398));
  jor  g13153(.dina(n13398), .dinb(asqrt[32] ), .dout(n13399));
  jand g13154(.dina(n13056), .dinb(n13399), .dout(n13400));
  jor  g13155(.dina(n13400), .dinb(n13338), .dout(n13401));
  jor  g13156(.dina(n13401), .dinb(asqrt[33] ), .dout(n13402));
  jnot g13157(.din(n13064), .dout(n13403));
  jand g13158(.dina(n13403), .dinb(n13402), .dout(n13404));
  jor  g13159(.dina(n13404), .dinb(n13337), .dout(n13405));
  jor  g13160(.dina(n13405), .dinb(asqrt[34] ), .dout(n13406));
  jand g13161(.dina(n13071), .dinb(n13406), .dout(n13407));
  jor  g13162(.dina(n13407), .dinb(n13336), .dout(n13408));
  jor  g13163(.dina(n13408), .dinb(asqrt[35] ), .dout(n13409));
  jnot g13164(.din(n13079), .dout(n13410));
  jand g13165(.dina(n13410), .dinb(n13409), .dout(n13411));
  jor  g13166(.dina(n13411), .dinb(n13335), .dout(n13412));
  jor  g13167(.dina(n13412), .dinb(asqrt[36] ), .dout(n13413));
  jnot g13168(.din(n13086), .dout(n13414));
  jand g13169(.dina(n13414), .dinb(n13413), .dout(n13415));
  jor  g13170(.dina(n13415), .dinb(n13334), .dout(n13416));
  jor  g13171(.dina(n13416), .dinb(asqrt[37] ), .dout(n13417));
  jnot g13172(.din(n13093), .dout(n13418));
  jand g13173(.dina(n13418), .dinb(n13417), .dout(n13419));
  jor  g13174(.dina(n13419), .dinb(n13333), .dout(n13420));
  jor  g13175(.dina(n13420), .dinb(asqrt[38] ), .dout(n13421));
  jand g13176(.dina(n13100), .dinb(n13421), .dout(n13422));
  jor  g13177(.dina(n13422), .dinb(n13332), .dout(n13423));
  jor  g13178(.dina(n13423), .dinb(asqrt[39] ), .dout(n13424));
  jnot g13179(.din(n13108), .dout(n13425));
  jand g13180(.dina(n13425), .dinb(n13424), .dout(n13426));
  jor  g13181(.dina(n13426), .dinb(n13331), .dout(n13427));
  jor  g13182(.dina(n13427), .dinb(asqrt[40] ), .dout(n13428));
  jnot g13183(.din(n13115), .dout(n13429));
  jand g13184(.dina(n13429), .dinb(n13428), .dout(n13430));
  jor  g13185(.dina(n13430), .dinb(n13330), .dout(n13431));
  jor  g13186(.dina(n13431), .dinb(asqrt[41] ), .dout(n13432));
  jnot g13187(.din(n13122), .dout(n13433));
  jand g13188(.dina(n13433), .dinb(n13432), .dout(n13434));
  jor  g13189(.dina(n13434), .dinb(n13329), .dout(n13435));
  jor  g13190(.dina(n13435), .dinb(asqrt[42] ), .dout(n13436));
  jnot g13191(.din(n13129), .dout(n13437));
  jand g13192(.dina(n13437), .dinb(n13436), .dout(n13438));
  jor  g13193(.dina(n13438), .dinb(n13328), .dout(n13439));
  jor  g13194(.dina(n13439), .dinb(asqrt[43] ), .dout(n13440));
  jand g13195(.dina(n13136), .dinb(n13440), .dout(n13441));
  jor  g13196(.dina(n13441), .dinb(n13327), .dout(n13442));
  jor  g13197(.dina(n13442), .dinb(asqrt[44] ), .dout(n13443));
  jand g13198(.dina(n13443), .dinb(n13143), .dout(n13444));
  jor  g13199(.dina(n13444), .dinb(n13326), .dout(n13445));
  jor  g13200(.dina(n13445), .dinb(asqrt[45] ), .dout(n13446));
  jnot g13201(.din(n13152), .dout(n13447));
  jand g13202(.dina(n13447), .dinb(n13446), .dout(n13448));
  jor  g13203(.dina(n13448), .dinb(n13325), .dout(n13449));
  jor  g13204(.dina(n13449), .dinb(asqrt[46] ), .dout(n13450));
  jand g13205(.dina(n13159), .dinb(n13450), .dout(n13451));
  jor  g13206(.dina(n13451), .dinb(n13324), .dout(n13452));
  jor  g13207(.dina(n13452), .dinb(asqrt[47] ), .dout(n13453));
  jnot g13208(.din(n13167), .dout(n13454));
  jand g13209(.dina(n13454), .dinb(n13453), .dout(n13455));
  jor  g13210(.dina(n13455), .dinb(n13323), .dout(n13456));
  jor  g13211(.dina(n13456), .dinb(asqrt[48] ), .dout(n13457));
  jand g13212(.dina(n13174), .dinb(n13457), .dout(n13458));
  jor  g13213(.dina(n13458), .dinb(n13322), .dout(n13459));
  jor  g13214(.dina(n13459), .dinb(asqrt[49] ), .dout(n13460));
  jnot g13215(.din(n13182), .dout(n13461));
  jand g13216(.dina(n13461), .dinb(n13460), .dout(n13462));
  jor  g13217(.dina(n13462), .dinb(n13321), .dout(n13463));
  jor  g13218(.dina(n13463), .dinb(asqrt[50] ), .dout(n13464));
  jnot g13219(.din(n13189), .dout(n13465));
  jand g13220(.dina(n13465), .dinb(n13464), .dout(n13466));
  jor  g13221(.dina(n13466), .dinb(n13320), .dout(n13467));
  jor  g13222(.dina(n13467), .dinb(asqrt[51] ), .dout(n13468));
  jnot g13223(.din(n13196), .dout(n13469));
  jand g13224(.dina(n13469), .dinb(n13468), .dout(n13470));
  jor  g13225(.dina(n13470), .dinb(n13319), .dout(n13471));
  jor  g13226(.dina(n13471), .dinb(asqrt[52] ), .dout(n13472));
  jand g13227(.dina(n13203), .dinb(n13472), .dout(n13473));
  jor  g13228(.dina(n13473), .dinb(n13318), .dout(n13474));
  jor  g13229(.dina(n13474), .dinb(asqrt[53] ), .dout(n13475));
  jnot g13230(.din(n13211), .dout(n13476));
  jand g13231(.dina(n13476), .dinb(n13475), .dout(n13477));
  jor  g13232(.dina(n13477), .dinb(n13317), .dout(n13478));
  jor  g13233(.dina(n13478), .dinb(asqrt[54] ), .dout(n13479));
  jand g13234(.dina(n13218), .dinb(n13479), .dout(n13480));
  jor  g13235(.dina(n13480), .dinb(n13316), .dout(n13481));
  jor  g13236(.dina(n13481), .dinb(asqrt[55] ), .dout(n13482));
  jnot g13237(.din(n13226), .dout(n13483));
  jand g13238(.dina(n13483), .dinb(n13482), .dout(n13484));
  jor  g13239(.dina(n13484), .dinb(n13315), .dout(n13485));
  jor  g13240(.dina(n13485), .dinb(asqrt[56] ), .dout(n13486));
  jand g13241(.dina(n13233), .dinb(n13486), .dout(n13487));
  jor  g13242(.dina(n13487), .dinb(n13314), .dout(n13488));
  jor  g13243(.dina(n13488), .dinb(asqrt[57] ), .dout(n13489));
  jnot g13244(.din(n13241), .dout(n13490));
  jand g13245(.dina(n13490), .dinb(n13489), .dout(n13491));
  jor  g13246(.dina(n13491), .dinb(n13313), .dout(n13492));
  jor  g13247(.dina(n13492), .dinb(asqrt[58] ), .dout(n13493));
  jand g13248(.dina(n13248), .dinb(n13493), .dout(n13494));
  jor  g13249(.dina(n13494), .dinb(n13312), .dout(n13495));
  jor  g13250(.dina(n13495), .dinb(asqrt[59] ), .dout(n13496));
  jand g13251(.dina(n13256), .dinb(n13496), .dout(n13497));
  jor  g13252(.dina(n13497), .dinb(n13311), .dout(n13498));
  jor  g13253(.dina(n13498), .dinb(asqrt[60] ), .dout(n13499));
  jand g13254(.dina(n13264), .dinb(n13499), .dout(n13500));
  jor  g13255(.dina(n13500), .dinb(n13310), .dout(n13501));
  jor  g13256(.dina(n13501), .dinb(asqrt[61] ), .dout(n13502));
  jnot g13257(.din(n13272), .dout(n13503));
  jand g13258(.dina(n13503), .dinb(n13502), .dout(n13504));
  jor  g13259(.dina(n13504), .dinb(n13309), .dout(n13505));
  jor  g13260(.dina(n13505), .dinb(asqrt[62] ), .dout(n13506));
  jnot g13261(.din(n13279), .dout(n13507));
  jand g13262(.dina(n13507), .dinb(n13506), .dout(n13508));
  jor  g13263(.dina(n13508), .dinb(n13308), .dout(n13509));
  jand g13264(.dina(n13509), .dinb(n12950), .dout(n13510));
  jand g13265(.dina(n13510), .dinb(n12731), .dout(n13511));
  jand g13266(.dina(n13511), .dinb(n13307), .dout(n13512));
  jor  g13267(.dina(n13512), .dinb(asqrt[63] ), .dout(n13513));
  jnot g13268(.din(n13294), .dout(n13514));
  jand g13269(.dina(n13514), .dinb(n13513), .dout(n13515));
  jor  g13270(.dina(n13515), .dinb(n13306), .dout(n13516));
  jand g13271(.dina(n13516), .dinb(n13305), .dout(n13517));
  jand g13272(.dina(n13517), .dinb(n13303), .dout(n13518));
  jor  g13273(.dina(n13518), .dinb(n13302), .dout(n13519));
  jand g13274(.dina(n13519), .dinb(asqrt[20] ), .dout(n13520));
  jor  g13275(.dina(n13519), .dinb(asqrt[20] ), .dout(n13521));
  jor  g13276(.dina(n13292), .dinb(n13287), .dout(n13522));
  jor  g13277(.dina(n13522), .dinb(n13285), .dout(n13523));
  jor  g13278(.dina(n13523), .dinb(n12947), .dout(n13524));
  jand g13279(.dina(n13524), .dinb(n13516), .dout(n13525));
  jxor g13280(.dina(n13525), .dinb(n12196), .dout(n13526));
  jnot g13281(.din(n13526), .dout(n13527));
  jand g13282(.dina(n13527), .dinb(n13521), .dout(n13528));
  jor  g13283(.dina(n13528), .dinb(n13520), .dout(n13529));
  jand g13284(.dina(n13529), .dinb(asqrt[21] ), .dout(n13530));
  jor  g13285(.dina(n13529), .dinb(asqrt[21] ), .dout(n13531));
  jxor g13286(.dina(n12958), .dinb(n12410), .dout(n13532));
  jand g13287(.dina(n13532), .dinb(asqrt[18] ), .dout(n13533));
  jxor g13288(.dina(n13533), .dinb(n12964), .dout(n13534));
  jnot g13289(.din(n13534), .dout(n13535));
  jand g13290(.dina(n13535), .dinb(n13531), .dout(n13536));
  jor  g13291(.dina(n13536), .dinb(n13530), .dout(n13537));
  jand g13292(.dina(n13537), .dinb(asqrt[22] ), .dout(n13538));
  jor  g13293(.dina(n13537), .dinb(asqrt[22] ), .dout(n13539));
  jxor g13294(.dina(n12966), .dinb(n11858), .dout(n13540));
  jand g13295(.dina(n13540), .dinb(asqrt[18] ), .dout(n13541));
  jxor g13296(.dina(n13541), .dinb(n12975), .dout(n13542));
  jnot g13297(.din(n13542), .dout(n13543));
  jand g13298(.dina(n13543), .dinb(n13539), .dout(n13544));
  jor  g13299(.dina(n13544), .dinb(n13538), .dout(n13545));
  jand g13300(.dina(n13545), .dinb(asqrt[23] ), .dout(n13546));
  jor  g13301(.dina(n13545), .dinb(asqrt[23] ), .dout(n13547));
  jxor g13302(.dina(n12977), .dinb(n11347), .dout(n13548));
  jand g13303(.dina(n13548), .dinb(asqrt[18] ), .dout(n13549));
  jxor g13304(.dina(n13549), .dinb(n12982), .dout(n13550));
  jand g13305(.dina(n13550), .dinb(n13547), .dout(n13551));
  jor  g13306(.dina(n13551), .dinb(n13546), .dout(n13552));
  jand g13307(.dina(n13552), .dinb(asqrt[24] ), .dout(n13553));
  jor  g13308(.dina(n13552), .dinb(asqrt[24] ), .dout(n13554));
  jxor g13309(.dina(n12985), .dinb(n10824), .dout(n13555));
  jand g13310(.dina(n13555), .dinb(asqrt[18] ), .dout(n13556));
  jxor g13311(.dina(n13556), .dinb(n12990), .dout(n13557));
  jnot g13312(.din(n13557), .dout(n13558));
  jand g13313(.dina(n13558), .dinb(n13554), .dout(n13559));
  jor  g13314(.dina(n13559), .dinb(n13553), .dout(n13560));
  jand g13315(.dina(n13560), .dinb(asqrt[25] ), .dout(n13561));
  jor  g13316(.dina(n13560), .dinb(asqrt[25] ), .dout(n13562));
  jxor g13317(.dina(n12992), .dinb(n10328), .dout(n13563));
  jand g13318(.dina(n13563), .dinb(asqrt[18] ), .dout(n13564));
  jxor g13319(.dina(n13564), .dinb(n12997), .dout(n13565));
  jand g13320(.dina(n13565), .dinb(n13562), .dout(n13566));
  jor  g13321(.dina(n13566), .dinb(n13561), .dout(n13567));
  jand g13322(.dina(n13567), .dinb(asqrt[26] ), .dout(n13568));
  jor  g13323(.dina(n13567), .dinb(asqrt[26] ), .dout(n13569));
  jxor g13324(.dina(n13000), .dinb(n9832), .dout(n13570));
  jand g13325(.dina(n13570), .dinb(asqrt[18] ), .dout(n13571));
  jxor g13326(.dina(n13571), .dinb(n13005), .dout(n13572));
  jnot g13327(.din(n13572), .dout(n13573));
  jand g13328(.dina(n13573), .dinb(n13569), .dout(n13574));
  jor  g13329(.dina(n13574), .dinb(n13568), .dout(n13575));
  jand g13330(.dina(n13575), .dinb(asqrt[27] ), .dout(n13576));
  jor  g13331(.dina(n13575), .dinb(asqrt[27] ), .dout(n13577));
  jxor g13332(.dina(n13007), .dinb(n9369), .dout(n13578));
  jand g13333(.dina(n13578), .dinb(asqrt[18] ), .dout(n13579));
  jxor g13334(.dina(n13579), .dinb(n13012), .dout(n13580));
  jand g13335(.dina(n13580), .dinb(n13577), .dout(n13581));
  jor  g13336(.dina(n13581), .dinb(n13576), .dout(n13582));
  jand g13337(.dina(n13582), .dinb(asqrt[28] ), .dout(n13583));
  jor  g13338(.dina(n13582), .dinb(asqrt[28] ), .dout(n13584));
  jxor g13339(.dina(n13015), .dinb(n8890), .dout(n13585));
  jand g13340(.dina(n13585), .dinb(asqrt[18] ), .dout(n13586));
  jxor g13341(.dina(n13586), .dinb(n13020), .dout(n13587));
  jnot g13342(.din(n13587), .dout(n13588));
  jand g13343(.dina(n13588), .dinb(n13584), .dout(n13589));
  jor  g13344(.dina(n13589), .dinb(n13583), .dout(n13590));
  jand g13345(.dina(n13590), .dinb(asqrt[29] ), .dout(n13591));
  jor  g13346(.dina(n13590), .dinb(asqrt[29] ), .dout(n13592));
  jxor g13347(.dina(n13022), .dinb(n8449), .dout(n13593));
  jand g13348(.dina(n13593), .dinb(asqrt[18] ), .dout(n13594));
  jxor g13349(.dina(n13594), .dinb(n13027), .dout(n13595));
  jand g13350(.dina(n13595), .dinb(n13592), .dout(n13596));
  jor  g13351(.dina(n13596), .dinb(n13591), .dout(n13597));
  jand g13352(.dina(n13597), .dinb(asqrt[30] ), .dout(n13598));
  jor  g13353(.dina(n13597), .dinb(asqrt[30] ), .dout(n13599));
  jxor g13354(.dina(n13030), .dinb(n8003), .dout(n13600));
  jand g13355(.dina(n13600), .dinb(asqrt[18] ), .dout(n13601));
  jxor g13356(.dina(n13601), .dinb(n13035), .dout(n13602));
  jnot g13357(.din(n13602), .dout(n13603));
  jand g13358(.dina(n13603), .dinb(n13599), .dout(n13604));
  jor  g13359(.dina(n13604), .dinb(n13598), .dout(n13605));
  jand g13360(.dina(n13605), .dinb(asqrt[31] ), .dout(n13606));
  jor  g13361(.dina(n13605), .dinb(asqrt[31] ), .dout(n13607));
  jxor g13362(.dina(n13037), .dinb(n7581), .dout(n13608));
  jand g13363(.dina(n13608), .dinb(asqrt[18] ), .dout(n13609));
  jxor g13364(.dina(n13609), .dinb(n13042), .dout(n13610));
  jnot g13365(.din(n13610), .dout(n13611));
  jand g13366(.dina(n13611), .dinb(n13607), .dout(n13612));
  jor  g13367(.dina(n13612), .dinb(n13606), .dout(n13613));
  jand g13368(.dina(n13613), .dinb(asqrt[32] ), .dout(n13614));
  jor  g13369(.dina(n13613), .dinb(asqrt[32] ), .dout(n13615));
  jxor g13370(.dina(n13044), .dinb(n7154), .dout(n13616));
  jand g13371(.dina(n13616), .dinb(asqrt[18] ), .dout(n13617));
  jxor g13372(.dina(n13617), .dinb(n13049), .dout(n13618));
  jnot g13373(.din(n13618), .dout(n13619));
  jand g13374(.dina(n13619), .dinb(n13615), .dout(n13620));
  jor  g13375(.dina(n13620), .dinb(n13614), .dout(n13621));
  jand g13376(.dina(n13621), .dinb(asqrt[33] ), .dout(n13622));
  jor  g13377(.dina(n13621), .dinb(asqrt[33] ), .dout(n13623));
  jxor g13378(.dina(n13051), .dinb(n6758), .dout(n13624));
  jand g13379(.dina(n13624), .dinb(asqrt[18] ), .dout(n13625));
  jxor g13380(.dina(n13625), .dinb(n13056), .dout(n13626));
  jand g13381(.dina(n13626), .dinb(n13623), .dout(n13627));
  jor  g13382(.dina(n13627), .dinb(n13622), .dout(n13628));
  jand g13383(.dina(n13628), .dinb(asqrt[34] ), .dout(n13629));
  jor  g13384(.dina(n13628), .dinb(asqrt[34] ), .dout(n13630));
  jxor g13385(.dina(n13059), .dinb(n6357), .dout(n13631));
  jand g13386(.dina(n13631), .dinb(asqrt[18] ), .dout(n13632));
  jxor g13387(.dina(n13632), .dinb(n13064), .dout(n13633));
  jnot g13388(.din(n13633), .dout(n13634));
  jand g13389(.dina(n13634), .dinb(n13630), .dout(n13635));
  jor  g13390(.dina(n13635), .dinb(n13629), .dout(n13636));
  jand g13391(.dina(n13636), .dinb(asqrt[35] ), .dout(n13637));
  jor  g13392(.dina(n13636), .dinb(asqrt[35] ), .dout(n13638));
  jxor g13393(.dina(n13066), .dinb(n5989), .dout(n13639));
  jand g13394(.dina(n13639), .dinb(asqrt[18] ), .dout(n13640));
  jxor g13395(.dina(n13640), .dinb(n13071), .dout(n13641));
  jand g13396(.dina(n13641), .dinb(n13638), .dout(n13642));
  jor  g13397(.dina(n13642), .dinb(n13637), .dout(n13643));
  jand g13398(.dina(n13643), .dinb(asqrt[36] ), .dout(n13644));
  jor  g13399(.dina(n13643), .dinb(asqrt[36] ), .dout(n13645));
  jxor g13400(.dina(n13074), .dinb(n5606), .dout(n13646));
  jand g13401(.dina(n13646), .dinb(asqrt[18] ), .dout(n13647));
  jxor g13402(.dina(n13647), .dinb(n13079), .dout(n13648));
  jnot g13403(.din(n13648), .dout(n13649));
  jand g13404(.dina(n13649), .dinb(n13645), .dout(n13650));
  jor  g13405(.dina(n13650), .dinb(n13644), .dout(n13651));
  jand g13406(.dina(n13651), .dinb(asqrt[37] ), .dout(n13652));
  jor  g13407(.dina(n13651), .dinb(asqrt[37] ), .dout(n13653));
  jxor g13408(.dina(n13081), .dinb(n5259), .dout(n13654));
  jand g13409(.dina(n13654), .dinb(asqrt[18] ), .dout(n13655));
  jxor g13410(.dina(n13655), .dinb(n13086), .dout(n13656));
  jnot g13411(.din(n13656), .dout(n13657));
  jand g13412(.dina(n13657), .dinb(n13653), .dout(n13658));
  jor  g13413(.dina(n13658), .dinb(n13652), .dout(n13659));
  jand g13414(.dina(n13659), .dinb(asqrt[38] ), .dout(n13660));
  jor  g13415(.dina(n13659), .dinb(asqrt[38] ), .dout(n13661));
  jxor g13416(.dina(n13088), .dinb(n4902), .dout(n13662));
  jand g13417(.dina(n13662), .dinb(asqrt[18] ), .dout(n13663));
  jxor g13418(.dina(n13663), .dinb(n13093), .dout(n13664));
  jnot g13419(.din(n13664), .dout(n13665));
  jand g13420(.dina(n13665), .dinb(n13661), .dout(n13666));
  jor  g13421(.dina(n13666), .dinb(n13660), .dout(n13667));
  jand g13422(.dina(n13667), .dinb(asqrt[39] ), .dout(n13668));
  jor  g13423(.dina(n13667), .dinb(asqrt[39] ), .dout(n13669));
  jxor g13424(.dina(n13095), .dinb(n4582), .dout(n13670));
  jand g13425(.dina(n13670), .dinb(asqrt[18] ), .dout(n13671));
  jxor g13426(.dina(n13671), .dinb(n13100), .dout(n13672));
  jand g13427(.dina(n13672), .dinb(n13669), .dout(n13673));
  jor  g13428(.dina(n13673), .dinb(n13668), .dout(n13674));
  jand g13429(.dina(n13674), .dinb(asqrt[40] ), .dout(n13675));
  jor  g13430(.dina(n13674), .dinb(asqrt[40] ), .dout(n13676));
  jxor g13431(.dina(n13103), .dinb(n4249), .dout(n13677));
  jand g13432(.dina(n13677), .dinb(asqrt[18] ), .dout(n13678));
  jxor g13433(.dina(n13678), .dinb(n13108), .dout(n13679));
  jnot g13434(.din(n13679), .dout(n13680));
  jand g13435(.dina(n13680), .dinb(n13676), .dout(n13681));
  jor  g13436(.dina(n13681), .dinb(n13675), .dout(n13682));
  jand g13437(.dina(n13682), .dinb(asqrt[41] ), .dout(n13683));
  jor  g13438(.dina(n13682), .dinb(asqrt[41] ), .dout(n13684));
  jxor g13439(.dina(n13110), .dinb(n3955), .dout(n13685));
  jand g13440(.dina(n13685), .dinb(asqrt[18] ), .dout(n13686));
  jxor g13441(.dina(n13686), .dinb(n13115), .dout(n13687));
  jnot g13442(.din(n13687), .dout(n13688));
  jand g13443(.dina(n13688), .dinb(n13684), .dout(n13689));
  jor  g13444(.dina(n13689), .dinb(n13683), .dout(n13690));
  jand g13445(.dina(n13690), .dinb(asqrt[42] ), .dout(n13691));
  jor  g13446(.dina(n13690), .dinb(asqrt[42] ), .dout(n13692));
  jxor g13447(.dina(n13117), .dinb(n3642), .dout(n13693));
  jand g13448(.dina(n13693), .dinb(asqrt[18] ), .dout(n13694));
  jxor g13449(.dina(n13694), .dinb(n13122), .dout(n13695));
  jnot g13450(.din(n13695), .dout(n13696));
  jand g13451(.dina(n13696), .dinb(n13692), .dout(n13697));
  jor  g13452(.dina(n13697), .dinb(n13691), .dout(n13698));
  jand g13453(.dina(n13698), .dinb(asqrt[43] ), .dout(n13699));
  jor  g13454(.dina(n13698), .dinb(asqrt[43] ), .dout(n13700));
  jxor g13455(.dina(n13124), .dinb(n3368), .dout(n13701));
  jand g13456(.dina(n13701), .dinb(asqrt[18] ), .dout(n13702));
  jxor g13457(.dina(n13702), .dinb(n13129), .dout(n13703));
  jnot g13458(.din(n13703), .dout(n13704));
  jand g13459(.dina(n13704), .dinb(n13700), .dout(n13705));
  jor  g13460(.dina(n13705), .dinb(n13699), .dout(n13706));
  jand g13461(.dina(n13706), .dinb(asqrt[44] ), .dout(n13707));
  jor  g13462(.dina(n13706), .dinb(asqrt[44] ), .dout(n13708));
  jxor g13463(.dina(n13131), .dinb(n3089), .dout(n13709));
  jand g13464(.dina(n13709), .dinb(asqrt[18] ), .dout(n13710));
  jxor g13465(.dina(n13710), .dinb(n13136), .dout(n13711));
  jand g13466(.dina(n13711), .dinb(n13708), .dout(n13712));
  jor  g13467(.dina(n13712), .dinb(n13707), .dout(n13713));
  jand g13468(.dina(n13713), .dinb(asqrt[45] ), .dout(n13714));
  jxor g13469(.dina(n13139), .dinb(n2833), .dout(n13715));
  jand g13470(.dina(n13715), .dinb(asqrt[18] ), .dout(n13716));
  jxor g13471(.dina(n13716), .dinb(n13143), .dout(n13717));
  jor  g13472(.dina(n13713), .dinb(asqrt[45] ), .dout(n13718));
  jand g13473(.dina(n13718), .dinb(n13717), .dout(n13719));
  jor  g13474(.dina(n13719), .dinb(n13714), .dout(n13720));
  jand g13475(.dina(n13720), .dinb(asqrt[46] ), .dout(n13721));
  jor  g13476(.dina(n13720), .dinb(asqrt[46] ), .dout(n13722));
  jxor g13477(.dina(n13147), .dinb(n2572), .dout(n13723));
  jand g13478(.dina(n13723), .dinb(asqrt[18] ), .dout(n13724));
  jxor g13479(.dina(n13724), .dinb(n13152), .dout(n13725));
  jnot g13480(.din(n13725), .dout(n13726));
  jand g13481(.dina(n13726), .dinb(n13722), .dout(n13727));
  jor  g13482(.dina(n13727), .dinb(n13721), .dout(n13728));
  jand g13483(.dina(n13728), .dinb(asqrt[47] ), .dout(n13729));
  jor  g13484(.dina(n13728), .dinb(asqrt[47] ), .dout(n13730));
  jxor g13485(.dina(n13154), .dinb(n2345), .dout(n13731));
  jand g13486(.dina(n13731), .dinb(asqrt[18] ), .dout(n13732));
  jxor g13487(.dina(n13732), .dinb(n13159), .dout(n13733));
  jand g13488(.dina(n13733), .dinb(n13730), .dout(n13734));
  jor  g13489(.dina(n13734), .dinb(n13729), .dout(n13735));
  jand g13490(.dina(n13735), .dinb(asqrt[48] ), .dout(n13736));
  jor  g13491(.dina(n13735), .dinb(asqrt[48] ), .dout(n13737));
  jxor g13492(.dina(n13162), .dinb(n2108), .dout(n13738));
  jand g13493(.dina(n13738), .dinb(asqrt[18] ), .dout(n13739));
  jxor g13494(.dina(n13739), .dinb(n13167), .dout(n13740));
  jnot g13495(.din(n13740), .dout(n13741));
  jand g13496(.dina(n13741), .dinb(n13737), .dout(n13742));
  jor  g13497(.dina(n13742), .dinb(n13736), .dout(n13743));
  jand g13498(.dina(n13743), .dinb(asqrt[49] ), .dout(n13744));
  jor  g13499(.dina(n13743), .dinb(asqrt[49] ), .dout(n13745));
  jxor g13500(.dina(n13169), .dinb(n1912), .dout(n13746));
  jand g13501(.dina(n13746), .dinb(asqrt[18] ), .dout(n13747));
  jxor g13502(.dina(n13747), .dinb(n13174), .dout(n13748));
  jand g13503(.dina(n13748), .dinb(n13745), .dout(n13749));
  jor  g13504(.dina(n13749), .dinb(n13744), .dout(n13750));
  jand g13505(.dina(n13750), .dinb(asqrt[50] ), .dout(n13751));
  jor  g13506(.dina(n13750), .dinb(asqrt[50] ), .dout(n13752));
  jxor g13507(.dina(n13177), .dinb(n1699), .dout(n13753));
  jand g13508(.dina(n13753), .dinb(asqrt[18] ), .dout(n13754));
  jxor g13509(.dina(n13754), .dinb(n13182), .dout(n13755));
  jnot g13510(.din(n13755), .dout(n13756));
  jand g13511(.dina(n13756), .dinb(n13752), .dout(n13757));
  jor  g13512(.dina(n13757), .dinb(n13751), .dout(n13758));
  jand g13513(.dina(n13758), .dinb(asqrt[51] ), .dout(n13759));
  jor  g13514(.dina(n13758), .dinb(asqrt[51] ), .dout(n13760));
  jxor g13515(.dina(n13184), .dinb(n1516), .dout(n13761));
  jand g13516(.dina(n13761), .dinb(asqrt[18] ), .dout(n13762));
  jxor g13517(.dina(n13762), .dinb(n13189), .dout(n13763));
  jnot g13518(.din(n13763), .dout(n13764));
  jand g13519(.dina(n13764), .dinb(n13760), .dout(n13765));
  jor  g13520(.dina(n13765), .dinb(n13759), .dout(n13766));
  jand g13521(.dina(n13766), .dinb(asqrt[52] ), .dout(n13767));
  jor  g13522(.dina(n13766), .dinb(asqrt[52] ), .dout(n13768));
  jxor g13523(.dina(n13191), .dinb(n1332), .dout(n13769));
  jand g13524(.dina(n13769), .dinb(asqrt[18] ), .dout(n13770));
  jxor g13525(.dina(n13770), .dinb(n13196), .dout(n13771));
  jnot g13526(.din(n13771), .dout(n13772));
  jand g13527(.dina(n13772), .dinb(n13768), .dout(n13773));
  jor  g13528(.dina(n13773), .dinb(n13767), .dout(n13774));
  jand g13529(.dina(n13774), .dinb(asqrt[53] ), .dout(n13775));
  jor  g13530(.dina(n13774), .dinb(asqrt[53] ), .dout(n13776));
  jxor g13531(.dina(n13198), .dinb(n1173), .dout(n13777));
  jand g13532(.dina(n13777), .dinb(asqrt[18] ), .dout(n13778));
  jxor g13533(.dina(n13778), .dinb(n13203), .dout(n13779));
  jand g13534(.dina(n13779), .dinb(n13776), .dout(n13780));
  jor  g13535(.dina(n13780), .dinb(n13775), .dout(n13781));
  jand g13536(.dina(n13781), .dinb(asqrt[54] ), .dout(n13782));
  jor  g13537(.dina(n13781), .dinb(asqrt[54] ), .dout(n13783));
  jxor g13538(.dina(n13206), .dinb(n1008), .dout(n13784));
  jand g13539(.dina(n13784), .dinb(asqrt[18] ), .dout(n13785));
  jxor g13540(.dina(n13785), .dinb(n13211), .dout(n13786));
  jnot g13541(.din(n13786), .dout(n13787));
  jand g13542(.dina(n13787), .dinb(n13783), .dout(n13788));
  jor  g13543(.dina(n13788), .dinb(n13782), .dout(n13789));
  jand g13544(.dina(n13789), .dinb(asqrt[55] ), .dout(n13790));
  jor  g13545(.dina(n13789), .dinb(asqrt[55] ), .dout(n13791));
  jxor g13546(.dina(n13213), .dinb(n884), .dout(n13792));
  jand g13547(.dina(n13792), .dinb(asqrt[18] ), .dout(n13793));
  jxor g13548(.dina(n13793), .dinb(n13218), .dout(n13794));
  jand g13549(.dina(n13794), .dinb(n13791), .dout(n13795));
  jor  g13550(.dina(n13795), .dinb(n13790), .dout(n13796));
  jand g13551(.dina(n13796), .dinb(asqrt[56] ), .dout(n13797));
  jor  g13552(.dina(n13796), .dinb(asqrt[56] ), .dout(n13798));
  jxor g13553(.dina(n13221), .dinb(n743), .dout(n13799));
  jand g13554(.dina(n13799), .dinb(asqrt[18] ), .dout(n13800));
  jxor g13555(.dina(n13800), .dinb(n13226), .dout(n13801));
  jnot g13556(.din(n13801), .dout(n13802));
  jand g13557(.dina(n13802), .dinb(n13798), .dout(n13803));
  jor  g13558(.dina(n13803), .dinb(n13797), .dout(n13804));
  jand g13559(.dina(n13804), .dinb(asqrt[57] ), .dout(n13805));
  jor  g13560(.dina(n13804), .dinb(asqrt[57] ), .dout(n13806));
  jxor g13561(.dina(n13228), .dinb(n635), .dout(n13807));
  jand g13562(.dina(n13807), .dinb(asqrt[18] ), .dout(n13808));
  jxor g13563(.dina(n13808), .dinb(n13233), .dout(n13809));
  jand g13564(.dina(n13809), .dinb(n13806), .dout(n13810));
  jor  g13565(.dina(n13810), .dinb(n13805), .dout(n13811));
  jand g13566(.dina(n13811), .dinb(asqrt[58] ), .dout(n13812));
  jor  g13567(.dina(n13811), .dinb(asqrt[58] ), .dout(n13813));
  jxor g13568(.dina(n13236), .dinb(n515), .dout(n13814));
  jand g13569(.dina(n13814), .dinb(asqrt[18] ), .dout(n13815));
  jxor g13570(.dina(n13815), .dinb(n13241), .dout(n13816));
  jnot g13571(.din(n13816), .dout(n13817));
  jand g13572(.dina(n13817), .dinb(n13813), .dout(n13818));
  jor  g13573(.dina(n13818), .dinb(n13812), .dout(n13819));
  jand g13574(.dina(n13819), .dinb(asqrt[59] ), .dout(n13820));
  jor  g13575(.dina(n13819), .dinb(asqrt[59] ), .dout(n13821));
  jxor g13576(.dina(n13243), .dinb(n443), .dout(n13822));
  jand g13577(.dina(n13822), .dinb(asqrt[18] ), .dout(n13823));
  jxor g13578(.dina(n13823), .dinb(n13248), .dout(n13824));
  jand g13579(.dina(n13824), .dinb(n13821), .dout(n13825));
  jor  g13580(.dina(n13825), .dinb(n13820), .dout(n13826));
  jand g13581(.dina(n13826), .dinb(asqrt[60] ), .dout(n13827));
  jor  g13582(.dina(n13826), .dinb(asqrt[60] ), .dout(n13828));
  jxor g13583(.dina(n13251), .dinb(n352), .dout(n13829));
  jand g13584(.dina(n13829), .dinb(asqrt[18] ), .dout(n13830));
  jxor g13585(.dina(n13830), .dinb(n13256), .dout(n13831));
  jand g13586(.dina(n13831), .dinb(n13828), .dout(n13832));
  jor  g13587(.dina(n13832), .dinb(n13827), .dout(n13833));
  jand g13588(.dina(n13833), .dinb(asqrt[61] ), .dout(n13834));
  jor  g13589(.dina(n13833), .dinb(asqrt[61] ), .dout(n13835));
  jxor g13590(.dina(n13259), .dinb(n294), .dout(n13836));
  jand g13591(.dina(n13836), .dinb(asqrt[18] ), .dout(n13837));
  jxor g13592(.dina(n13837), .dinb(n13264), .dout(n13838));
  jand g13593(.dina(n13838), .dinb(n13835), .dout(n13839));
  jor  g13594(.dina(n13839), .dinb(n13834), .dout(n13840));
  jand g13595(.dina(n13840), .dinb(asqrt[62] ), .dout(n13841));
  jor  g13596(.dina(n13840), .dinb(asqrt[62] ), .dout(n13842));
  jxor g13597(.dina(n13267), .dinb(n239), .dout(n13843));
  jand g13598(.dina(n13843), .dinb(asqrt[18] ), .dout(n13844));
  jxor g13599(.dina(n13844), .dinb(n13272), .dout(n13845));
  jnot g13600(.din(n13845), .dout(n13846));
  jand g13601(.dina(n13846), .dinb(n13842), .dout(n13847));
  jor  g13602(.dina(n13847), .dinb(n13841), .dout(n13848));
  jxor g13603(.dina(n13274), .dinb(n221), .dout(n13849));
  jand g13604(.dina(n13849), .dinb(asqrt[18] ), .dout(n13850));
  jxor g13605(.dina(n13850), .dinb(n13279), .dout(n13851));
  jnot g13606(.din(n13851), .dout(n13852));
  jor  g13607(.dina(n13852), .dinb(n13848), .dout(n13853));
  jnot g13608(.din(n13853), .dout(n13854));
  jand g13609(.dina(n13515), .dinb(n13281), .dout(n13855));
  jnot g13610(.din(n13855), .dout(n13856));
  jnot g13611(.din(n13287), .dout(n13857));
  jand g13612(.dina(n13282), .dinb(asqrt[63] ), .dout(n13858));
  jand g13613(.dina(n13858), .dinb(n13857), .dout(n13859));
  jand g13614(.dina(n13859), .dinb(n13856), .dout(n13860));
  jnot g13615(.din(n13841), .dout(n13861));
  jnot g13616(.din(n13834), .dout(n13862));
  jnot g13617(.din(n13827), .dout(n13863));
  jnot g13618(.din(n13820), .dout(n13864));
  jnot g13619(.din(n13812), .dout(n13865));
  jnot g13620(.din(n13805), .dout(n13866));
  jnot g13621(.din(n13797), .dout(n13867));
  jnot g13622(.din(n13790), .dout(n13868));
  jnot g13623(.din(n13782), .dout(n13869));
  jnot g13624(.din(n13775), .dout(n13870));
  jnot g13625(.din(n13767), .dout(n13871));
  jnot g13626(.din(n13759), .dout(n13872));
  jnot g13627(.din(n13751), .dout(n13873));
  jnot g13628(.din(n13744), .dout(n13874));
  jnot g13629(.din(n13736), .dout(n13875));
  jnot g13630(.din(n13729), .dout(n13876));
  jnot g13631(.din(n13721), .dout(n13877));
  jnot g13632(.din(n13714), .dout(n13878));
  jnot g13633(.din(n13717), .dout(n13879));
  jnot g13634(.din(n13707), .dout(n13880));
  jnot g13635(.din(n13699), .dout(n13881));
  jnot g13636(.din(n13691), .dout(n13882));
  jnot g13637(.din(n13683), .dout(n13883));
  jnot g13638(.din(n13675), .dout(n13884));
  jnot g13639(.din(n13668), .dout(n13885));
  jnot g13640(.din(n13660), .dout(n13886));
  jnot g13641(.din(n13652), .dout(n13887));
  jnot g13642(.din(n13644), .dout(n13888));
  jnot g13643(.din(n13637), .dout(n13889));
  jnot g13644(.din(n13629), .dout(n13890));
  jnot g13645(.din(n13622), .dout(n13891));
  jnot g13646(.din(n13614), .dout(n13892));
  jnot g13647(.din(n13606), .dout(n13893));
  jnot g13648(.din(n13598), .dout(n13894));
  jnot g13649(.din(n13591), .dout(n13895));
  jnot g13650(.din(n13583), .dout(n13896));
  jnot g13651(.din(n13576), .dout(n13897));
  jnot g13652(.din(n13568), .dout(n13898));
  jnot g13653(.din(n13561), .dout(n13899));
  jnot g13654(.din(n13553), .dout(n13900));
  jnot g13655(.din(n13546), .dout(n13901));
  jnot g13656(.din(n13538), .dout(n13902));
  jnot g13657(.din(n13530), .dout(n13903));
  jnot g13658(.din(n13520), .dout(n13904));
  jnot g13659(.din(n13302), .dout(n13905));
  jnot g13660(.din(n13299), .dout(n13906));
  jor  g13661(.dina(n13515), .dinb(n12953), .dout(n13907));
  jand g13662(.dina(n13907), .dinb(n13906), .dout(n13908));
  jand g13663(.dina(n13908), .dinb(n12947), .dout(n13909));
  jor  g13664(.dina(n13515), .dinb(a[36] ), .dout(n13910));
  jand g13665(.dina(n13910), .dinb(a[37] ), .dout(n13911));
  jand g13666(.dina(asqrt[18] ), .dinb(n12955), .dout(n13912));
  jor  g13667(.dina(n13912), .dinb(n13911), .dout(n13913));
  jor  g13668(.dina(n13913), .dinb(n13909), .dout(n13914));
  jand g13669(.dina(n13914), .dinb(n13905), .dout(n13915));
  jand g13670(.dina(n13915), .dinb(n12410), .dout(n13916));
  jor  g13671(.dina(n13526), .dinb(n13916), .dout(n13917));
  jand g13672(.dina(n13917), .dinb(n13904), .dout(n13918));
  jand g13673(.dina(n13918), .dinb(n11858), .dout(n13919));
  jor  g13674(.dina(n13534), .dinb(n13919), .dout(n13920));
  jand g13675(.dina(n13920), .dinb(n13903), .dout(n13921));
  jand g13676(.dina(n13921), .dinb(n11347), .dout(n13922));
  jor  g13677(.dina(n13542), .dinb(n13922), .dout(n13923));
  jand g13678(.dina(n13923), .dinb(n13902), .dout(n13924));
  jand g13679(.dina(n13924), .dinb(n10824), .dout(n13925));
  jnot g13680(.din(n13550), .dout(n13926));
  jor  g13681(.dina(n13926), .dinb(n13925), .dout(n13927));
  jand g13682(.dina(n13927), .dinb(n13901), .dout(n13928));
  jand g13683(.dina(n13928), .dinb(n10328), .dout(n13929));
  jor  g13684(.dina(n13557), .dinb(n13929), .dout(n13930));
  jand g13685(.dina(n13930), .dinb(n13900), .dout(n13931));
  jand g13686(.dina(n13931), .dinb(n9832), .dout(n13932));
  jnot g13687(.din(n13565), .dout(n13933));
  jor  g13688(.dina(n13933), .dinb(n13932), .dout(n13934));
  jand g13689(.dina(n13934), .dinb(n13899), .dout(n13935));
  jand g13690(.dina(n13935), .dinb(n9369), .dout(n13936));
  jor  g13691(.dina(n13572), .dinb(n13936), .dout(n13937));
  jand g13692(.dina(n13937), .dinb(n13898), .dout(n13938));
  jand g13693(.dina(n13938), .dinb(n8890), .dout(n13939));
  jnot g13694(.din(n13580), .dout(n13940));
  jor  g13695(.dina(n13940), .dinb(n13939), .dout(n13941));
  jand g13696(.dina(n13941), .dinb(n13897), .dout(n13942));
  jand g13697(.dina(n13942), .dinb(n8449), .dout(n13943));
  jor  g13698(.dina(n13587), .dinb(n13943), .dout(n13944));
  jand g13699(.dina(n13944), .dinb(n13896), .dout(n13945));
  jand g13700(.dina(n13945), .dinb(n8003), .dout(n13946));
  jnot g13701(.din(n13595), .dout(n13947));
  jor  g13702(.dina(n13947), .dinb(n13946), .dout(n13948));
  jand g13703(.dina(n13948), .dinb(n13895), .dout(n13949));
  jand g13704(.dina(n13949), .dinb(n7581), .dout(n13950));
  jor  g13705(.dina(n13602), .dinb(n13950), .dout(n13951));
  jand g13706(.dina(n13951), .dinb(n13894), .dout(n13952));
  jand g13707(.dina(n13952), .dinb(n7154), .dout(n13953));
  jor  g13708(.dina(n13610), .dinb(n13953), .dout(n13954));
  jand g13709(.dina(n13954), .dinb(n13893), .dout(n13955));
  jand g13710(.dina(n13955), .dinb(n6758), .dout(n13956));
  jor  g13711(.dina(n13618), .dinb(n13956), .dout(n13957));
  jand g13712(.dina(n13957), .dinb(n13892), .dout(n13958));
  jand g13713(.dina(n13958), .dinb(n6357), .dout(n13959));
  jnot g13714(.din(n13626), .dout(n13960));
  jor  g13715(.dina(n13960), .dinb(n13959), .dout(n13961));
  jand g13716(.dina(n13961), .dinb(n13891), .dout(n13962));
  jand g13717(.dina(n13962), .dinb(n5989), .dout(n13963));
  jor  g13718(.dina(n13633), .dinb(n13963), .dout(n13964));
  jand g13719(.dina(n13964), .dinb(n13890), .dout(n13965));
  jand g13720(.dina(n13965), .dinb(n5606), .dout(n13966));
  jnot g13721(.din(n13641), .dout(n13967));
  jor  g13722(.dina(n13967), .dinb(n13966), .dout(n13968));
  jand g13723(.dina(n13968), .dinb(n13889), .dout(n13969));
  jand g13724(.dina(n13969), .dinb(n5259), .dout(n13970));
  jor  g13725(.dina(n13648), .dinb(n13970), .dout(n13971));
  jand g13726(.dina(n13971), .dinb(n13888), .dout(n13972));
  jand g13727(.dina(n13972), .dinb(n4902), .dout(n13973));
  jor  g13728(.dina(n13656), .dinb(n13973), .dout(n13974));
  jand g13729(.dina(n13974), .dinb(n13887), .dout(n13975));
  jand g13730(.dina(n13975), .dinb(n4582), .dout(n13976));
  jor  g13731(.dina(n13664), .dinb(n13976), .dout(n13977));
  jand g13732(.dina(n13977), .dinb(n13886), .dout(n13978));
  jand g13733(.dina(n13978), .dinb(n4249), .dout(n13979));
  jnot g13734(.din(n13672), .dout(n13980));
  jor  g13735(.dina(n13980), .dinb(n13979), .dout(n13981));
  jand g13736(.dina(n13981), .dinb(n13885), .dout(n13982));
  jand g13737(.dina(n13982), .dinb(n3955), .dout(n13983));
  jor  g13738(.dina(n13679), .dinb(n13983), .dout(n13984));
  jand g13739(.dina(n13984), .dinb(n13884), .dout(n13985));
  jand g13740(.dina(n13985), .dinb(n3642), .dout(n13986));
  jor  g13741(.dina(n13687), .dinb(n13986), .dout(n13987));
  jand g13742(.dina(n13987), .dinb(n13883), .dout(n13988));
  jand g13743(.dina(n13988), .dinb(n3368), .dout(n13989));
  jor  g13744(.dina(n13695), .dinb(n13989), .dout(n13990));
  jand g13745(.dina(n13990), .dinb(n13882), .dout(n13991));
  jand g13746(.dina(n13991), .dinb(n3089), .dout(n13992));
  jor  g13747(.dina(n13703), .dinb(n13992), .dout(n13993));
  jand g13748(.dina(n13993), .dinb(n13881), .dout(n13994));
  jand g13749(.dina(n13994), .dinb(n2833), .dout(n13995));
  jnot g13750(.din(n13711), .dout(n13996));
  jor  g13751(.dina(n13996), .dinb(n13995), .dout(n13997));
  jand g13752(.dina(n13997), .dinb(n13880), .dout(n13998));
  jand g13753(.dina(n13998), .dinb(n2572), .dout(n13999));
  jor  g13754(.dina(n13999), .dinb(n13879), .dout(n14000));
  jand g13755(.dina(n14000), .dinb(n13878), .dout(n14001));
  jand g13756(.dina(n14001), .dinb(n2345), .dout(n14002));
  jor  g13757(.dina(n13725), .dinb(n14002), .dout(n14003));
  jand g13758(.dina(n14003), .dinb(n13877), .dout(n14004));
  jand g13759(.dina(n14004), .dinb(n2108), .dout(n14005));
  jnot g13760(.din(n13733), .dout(n14006));
  jor  g13761(.dina(n14006), .dinb(n14005), .dout(n14007));
  jand g13762(.dina(n14007), .dinb(n13876), .dout(n14008));
  jand g13763(.dina(n14008), .dinb(n1912), .dout(n14009));
  jor  g13764(.dina(n13740), .dinb(n14009), .dout(n14010));
  jand g13765(.dina(n14010), .dinb(n13875), .dout(n14011));
  jand g13766(.dina(n14011), .dinb(n1699), .dout(n14012));
  jnot g13767(.din(n13748), .dout(n14013));
  jor  g13768(.dina(n14013), .dinb(n14012), .dout(n14014));
  jand g13769(.dina(n14014), .dinb(n13874), .dout(n14015));
  jand g13770(.dina(n14015), .dinb(n1516), .dout(n14016));
  jor  g13771(.dina(n13755), .dinb(n14016), .dout(n14017));
  jand g13772(.dina(n14017), .dinb(n13873), .dout(n14018));
  jand g13773(.dina(n14018), .dinb(n1332), .dout(n14019));
  jor  g13774(.dina(n13763), .dinb(n14019), .dout(n14020));
  jand g13775(.dina(n14020), .dinb(n13872), .dout(n14021));
  jand g13776(.dina(n14021), .dinb(n1173), .dout(n14022));
  jor  g13777(.dina(n13771), .dinb(n14022), .dout(n14023));
  jand g13778(.dina(n14023), .dinb(n13871), .dout(n14024));
  jand g13779(.dina(n14024), .dinb(n1008), .dout(n14025));
  jnot g13780(.din(n13779), .dout(n14026));
  jor  g13781(.dina(n14026), .dinb(n14025), .dout(n14027));
  jand g13782(.dina(n14027), .dinb(n13870), .dout(n14028));
  jand g13783(.dina(n14028), .dinb(n884), .dout(n14029));
  jor  g13784(.dina(n13786), .dinb(n14029), .dout(n14030));
  jand g13785(.dina(n14030), .dinb(n13869), .dout(n14031));
  jand g13786(.dina(n14031), .dinb(n743), .dout(n14032));
  jnot g13787(.din(n13794), .dout(n14033));
  jor  g13788(.dina(n14033), .dinb(n14032), .dout(n14034));
  jand g13789(.dina(n14034), .dinb(n13868), .dout(n14035));
  jand g13790(.dina(n14035), .dinb(n635), .dout(n14036));
  jor  g13791(.dina(n13801), .dinb(n14036), .dout(n14037));
  jand g13792(.dina(n14037), .dinb(n13867), .dout(n14038));
  jand g13793(.dina(n14038), .dinb(n515), .dout(n14039));
  jnot g13794(.din(n13809), .dout(n14040));
  jor  g13795(.dina(n14040), .dinb(n14039), .dout(n14041));
  jand g13796(.dina(n14041), .dinb(n13866), .dout(n14042));
  jand g13797(.dina(n14042), .dinb(n443), .dout(n14043));
  jor  g13798(.dina(n13816), .dinb(n14043), .dout(n14044));
  jand g13799(.dina(n14044), .dinb(n13865), .dout(n14045));
  jand g13800(.dina(n14045), .dinb(n352), .dout(n14046));
  jnot g13801(.din(n13824), .dout(n14047));
  jor  g13802(.dina(n14047), .dinb(n14046), .dout(n14048));
  jand g13803(.dina(n14048), .dinb(n13864), .dout(n14049));
  jand g13804(.dina(n14049), .dinb(n294), .dout(n14050));
  jnot g13805(.din(n13831), .dout(n14051));
  jor  g13806(.dina(n14051), .dinb(n14050), .dout(n14052));
  jand g13807(.dina(n14052), .dinb(n13863), .dout(n14053));
  jand g13808(.dina(n14053), .dinb(n239), .dout(n14054));
  jnot g13809(.din(n13838), .dout(n14055));
  jor  g13810(.dina(n14055), .dinb(n14054), .dout(n14056));
  jand g13811(.dina(n14056), .dinb(n13862), .dout(n14057));
  jand g13812(.dina(n14057), .dinb(n221), .dout(n14058));
  jor  g13813(.dina(n13845), .dinb(n14058), .dout(n14059));
  jand g13814(.dina(n14059), .dinb(n13861), .dout(n14060));
  jor  g13815(.dina(n13851), .dinb(n14060), .dout(n14061));
  jand g13816(.dina(asqrt[18] ), .dinb(n13510), .dout(n14062));
  jor  g13817(.dina(n14062), .dinb(n13287), .dout(n14063));
  jor  g13818(.dina(n14063), .dinb(n14061), .dout(n14064));
  jand g13819(.dina(n14064), .dinb(n218), .dout(n14065));
  jand g13820(.dina(n13515), .dinb(n12951), .dout(n14066));
  jor  g13821(.dina(n14066), .dinb(n14065), .dout(n14067));
  jor  g13822(.dina(n14067), .dinb(n13860), .dout(n14068));
  jor  g13823(.dina(n14068), .dinb(n13854), .dout(asqrt[17] ));
  jnot g13824(.din(n13860), .dout(n14070));
  jand g13825(.dina(n13852), .dinb(n13848), .dout(n14071));
  jnot g13826(.din(n14063), .dout(n14072));
  jand g13827(.dina(n14072), .dinb(n14071), .dout(n14073));
  jor  g13828(.dina(n14073), .dinb(asqrt[63] ), .dout(n14074));
  jnot g13829(.din(n14066), .dout(n14075));
  jand g13830(.dina(n14075), .dinb(n14074), .dout(n14076));
  jand g13831(.dina(n14076), .dinb(n14070), .dout(n14077));
  jand g13832(.dina(n14077), .dinb(n13853), .dout(n14078));
  jor  g13833(.dina(n14078), .dinb(n13296), .dout(n14079));
  jnot g13834(.din(a[32] ), .dout(n14080));
  jnot g13835(.din(a[33] ), .dout(n14081));
  jand g13836(.dina(n14081), .dinb(n14080), .dout(n14082));
  jand g13837(.dina(n14082), .dinb(n13296), .dout(n14083));
  jnot g13838(.din(n14083), .dout(n14084));
  jand g13839(.dina(n14084), .dinb(n14079), .dout(n14085));
  jor  g13840(.dina(n14085), .dinb(n13515), .dout(n14086));
  jand g13841(.dina(n14085), .dinb(n13515), .dout(n14087));
  jor  g13842(.dina(n14078), .dinb(a[34] ), .dout(n14088));
  jand g13843(.dina(n14088), .dinb(a[35] ), .dout(n14089));
  jand g13844(.dina(asqrt[17] ), .dinb(n13298), .dout(n14090));
  jor  g13845(.dina(n14090), .dinb(n14089), .dout(n14091));
  jor  g13846(.dina(n14091), .dinb(n14087), .dout(n14092));
  jand g13847(.dina(n14092), .dinb(n14086), .dout(n14093));
  jor  g13848(.dina(n14093), .dinb(n12947), .dout(n14094));
  jand g13849(.dina(n14093), .dinb(n12947), .dout(n14095));
  jnot g13850(.din(n13298), .dout(n14096));
  jor  g13851(.dina(n14078), .dinb(n14096), .dout(n14097));
  jor  g13852(.dina(n13854), .dinb(n13515), .dout(n14098));
  jor  g13853(.dina(n14098), .dinb(n14065), .dout(n14099));
  jor  g13854(.dina(n14099), .dinb(n13859), .dout(n14100));
  jand g13855(.dina(n14100), .dinb(n14097), .dout(n14101));
  jxor g13856(.dina(n14101), .dinb(n12953), .dout(n14102));
  jor  g13857(.dina(n14102), .dinb(n14095), .dout(n14103));
  jand g13858(.dina(n14103), .dinb(n14094), .dout(n14104));
  jor  g13859(.dina(n14104), .dinb(n12410), .dout(n14105));
  jand g13860(.dina(n14104), .dinb(n12410), .dout(n14106));
  jxor g13861(.dina(n13301), .dinb(n12947), .dout(n14107));
  jor  g13862(.dina(n14107), .dinb(n14078), .dout(n14108));
  jxor g13863(.dina(n14108), .dinb(n13913), .dout(n14109));
  jnot g13864(.din(n14109), .dout(n14110));
  jor  g13865(.dina(n14110), .dinb(n14106), .dout(n14111));
  jand g13866(.dina(n14111), .dinb(n14105), .dout(n14112));
  jor  g13867(.dina(n14112), .dinb(n11858), .dout(n14113));
  jand g13868(.dina(n14112), .dinb(n11858), .dout(n14114));
  jxor g13869(.dina(n13519), .dinb(n12410), .dout(n14115));
  jor  g13870(.dina(n14115), .dinb(n14078), .dout(n14116));
  jxor g13871(.dina(n14116), .dinb(n13527), .dout(n14117));
  jor  g13872(.dina(n14117), .dinb(n14114), .dout(n14118));
  jand g13873(.dina(n14118), .dinb(n14113), .dout(n14119));
  jor  g13874(.dina(n14119), .dinb(n11347), .dout(n14120));
  jand g13875(.dina(n14119), .dinb(n11347), .dout(n14121));
  jxor g13876(.dina(n13529), .dinb(n11858), .dout(n14122));
  jor  g13877(.dina(n14122), .dinb(n14078), .dout(n14123));
  jxor g13878(.dina(n14123), .dinb(n13535), .dout(n14124));
  jor  g13879(.dina(n14124), .dinb(n14121), .dout(n14125));
  jand g13880(.dina(n14125), .dinb(n14120), .dout(n14126));
  jor  g13881(.dina(n14126), .dinb(n10824), .dout(n14127));
  jand g13882(.dina(n14126), .dinb(n10824), .dout(n14128));
  jxor g13883(.dina(n13537), .dinb(n11347), .dout(n14129));
  jor  g13884(.dina(n14129), .dinb(n14078), .dout(n14130));
  jxor g13885(.dina(n14130), .dinb(n13543), .dout(n14131));
  jor  g13886(.dina(n14131), .dinb(n14128), .dout(n14132));
  jand g13887(.dina(n14132), .dinb(n14127), .dout(n14133));
  jor  g13888(.dina(n14133), .dinb(n10328), .dout(n14134));
  jand g13889(.dina(n14133), .dinb(n10328), .dout(n14135));
  jxor g13890(.dina(n13545), .dinb(n10824), .dout(n14136));
  jor  g13891(.dina(n14136), .dinb(n14078), .dout(n14137));
  jxor g13892(.dina(n14137), .dinb(n13926), .dout(n14138));
  jnot g13893(.din(n14138), .dout(n14139));
  jor  g13894(.dina(n14139), .dinb(n14135), .dout(n14140));
  jand g13895(.dina(n14140), .dinb(n14134), .dout(n14141));
  jor  g13896(.dina(n14141), .dinb(n9832), .dout(n14142));
  jand g13897(.dina(n14141), .dinb(n9832), .dout(n14143));
  jxor g13898(.dina(n13552), .dinb(n10328), .dout(n14144));
  jor  g13899(.dina(n14144), .dinb(n14078), .dout(n14145));
  jxor g13900(.dina(n14145), .dinb(n13558), .dout(n14146));
  jor  g13901(.dina(n14146), .dinb(n14143), .dout(n14147));
  jand g13902(.dina(n14147), .dinb(n14142), .dout(n14148));
  jor  g13903(.dina(n14148), .dinb(n9369), .dout(n14149));
  jand g13904(.dina(n14148), .dinb(n9369), .dout(n14150));
  jxor g13905(.dina(n13560), .dinb(n9832), .dout(n14151));
  jor  g13906(.dina(n14151), .dinb(n14078), .dout(n14152));
  jxor g13907(.dina(n14152), .dinb(n13933), .dout(n14153));
  jnot g13908(.din(n14153), .dout(n14154));
  jor  g13909(.dina(n14154), .dinb(n14150), .dout(n14155));
  jand g13910(.dina(n14155), .dinb(n14149), .dout(n14156));
  jor  g13911(.dina(n14156), .dinb(n8890), .dout(n14157));
  jand g13912(.dina(n14156), .dinb(n8890), .dout(n14158));
  jxor g13913(.dina(n13567), .dinb(n9369), .dout(n14159));
  jor  g13914(.dina(n14159), .dinb(n14078), .dout(n14160));
  jxor g13915(.dina(n14160), .dinb(n13573), .dout(n14161));
  jor  g13916(.dina(n14161), .dinb(n14158), .dout(n14162));
  jand g13917(.dina(n14162), .dinb(n14157), .dout(n14163));
  jor  g13918(.dina(n14163), .dinb(n8449), .dout(n14164));
  jand g13919(.dina(n14163), .dinb(n8449), .dout(n14165));
  jxor g13920(.dina(n13575), .dinb(n8890), .dout(n14166));
  jor  g13921(.dina(n14166), .dinb(n14078), .dout(n14167));
  jxor g13922(.dina(n14167), .dinb(n13940), .dout(n14168));
  jnot g13923(.din(n14168), .dout(n14169));
  jor  g13924(.dina(n14169), .dinb(n14165), .dout(n14170));
  jand g13925(.dina(n14170), .dinb(n14164), .dout(n14171));
  jor  g13926(.dina(n14171), .dinb(n8003), .dout(n14172));
  jand g13927(.dina(n14171), .dinb(n8003), .dout(n14173));
  jxor g13928(.dina(n13582), .dinb(n8449), .dout(n14174));
  jor  g13929(.dina(n14174), .dinb(n14078), .dout(n14175));
  jxor g13930(.dina(n14175), .dinb(n13588), .dout(n14176));
  jor  g13931(.dina(n14176), .dinb(n14173), .dout(n14177));
  jand g13932(.dina(n14177), .dinb(n14172), .dout(n14178));
  jor  g13933(.dina(n14178), .dinb(n7581), .dout(n14179));
  jand g13934(.dina(n14178), .dinb(n7581), .dout(n14180));
  jxor g13935(.dina(n13590), .dinb(n8003), .dout(n14181));
  jor  g13936(.dina(n14181), .dinb(n14078), .dout(n14182));
  jxor g13937(.dina(n14182), .dinb(n13947), .dout(n14183));
  jnot g13938(.din(n14183), .dout(n14184));
  jor  g13939(.dina(n14184), .dinb(n14180), .dout(n14185));
  jand g13940(.dina(n14185), .dinb(n14179), .dout(n14186));
  jor  g13941(.dina(n14186), .dinb(n7154), .dout(n14187));
  jand g13942(.dina(n14186), .dinb(n7154), .dout(n14188));
  jxor g13943(.dina(n13597), .dinb(n7581), .dout(n14189));
  jor  g13944(.dina(n14189), .dinb(n14078), .dout(n14190));
  jxor g13945(.dina(n14190), .dinb(n13603), .dout(n14191));
  jor  g13946(.dina(n14191), .dinb(n14188), .dout(n14192));
  jand g13947(.dina(n14192), .dinb(n14187), .dout(n14193));
  jor  g13948(.dina(n14193), .dinb(n6758), .dout(n14194));
  jand g13949(.dina(n14193), .dinb(n6758), .dout(n14195));
  jxor g13950(.dina(n13605), .dinb(n7154), .dout(n14196));
  jor  g13951(.dina(n14196), .dinb(n14078), .dout(n14197));
  jxor g13952(.dina(n14197), .dinb(n13611), .dout(n14198));
  jor  g13953(.dina(n14198), .dinb(n14195), .dout(n14199));
  jand g13954(.dina(n14199), .dinb(n14194), .dout(n14200));
  jor  g13955(.dina(n14200), .dinb(n6357), .dout(n14201));
  jand g13956(.dina(n14200), .dinb(n6357), .dout(n14202));
  jxor g13957(.dina(n13613), .dinb(n6758), .dout(n14203));
  jor  g13958(.dina(n14203), .dinb(n14078), .dout(n14204));
  jxor g13959(.dina(n14204), .dinb(n13619), .dout(n14205));
  jor  g13960(.dina(n14205), .dinb(n14202), .dout(n14206));
  jand g13961(.dina(n14206), .dinb(n14201), .dout(n14207));
  jor  g13962(.dina(n14207), .dinb(n5989), .dout(n14208));
  jand g13963(.dina(n14207), .dinb(n5989), .dout(n14209));
  jxor g13964(.dina(n13621), .dinb(n6357), .dout(n14210));
  jor  g13965(.dina(n14210), .dinb(n14078), .dout(n14211));
  jxor g13966(.dina(n14211), .dinb(n13960), .dout(n14212));
  jnot g13967(.din(n14212), .dout(n14213));
  jor  g13968(.dina(n14213), .dinb(n14209), .dout(n14214));
  jand g13969(.dina(n14214), .dinb(n14208), .dout(n14215));
  jor  g13970(.dina(n14215), .dinb(n5606), .dout(n14216));
  jand g13971(.dina(n14215), .dinb(n5606), .dout(n14217));
  jxor g13972(.dina(n13628), .dinb(n5989), .dout(n14218));
  jor  g13973(.dina(n14218), .dinb(n14078), .dout(n14219));
  jxor g13974(.dina(n14219), .dinb(n13634), .dout(n14220));
  jor  g13975(.dina(n14220), .dinb(n14217), .dout(n14221));
  jand g13976(.dina(n14221), .dinb(n14216), .dout(n14222));
  jor  g13977(.dina(n14222), .dinb(n5259), .dout(n14223));
  jand g13978(.dina(n14222), .dinb(n5259), .dout(n14224));
  jxor g13979(.dina(n13636), .dinb(n5606), .dout(n14225));
  jor  g13980(.dina(n14225), .dinb(n14078), .dout(n14226));
  jxor g13981(.dina(n14226), .dinb(n13967), .dout(n14227));
  jnot g13982(.din(n14227), .dout(n14228));
  jor  g13983(.dina(n14228), .dinb(n14224), .dout(n14229));
  jand g13984(.dina(n14229), .dinb(n14223), .dout(n14230));
  jor  g13985(.dina(n14230), .dinb(n4902), .dout(n14231));
  jand g13986(.dina(n14230), .dinb(n4902), .dout(n14232));
  jxor g13987(.dina(n13643), .dinb(n5259), .dout(n14233));
  jor  g13988(.dina(n14233), .dinb(n14078), .dout(n14234));
  jxor g13989(.dina(n14234), .dinb(n13649), .dout(n14235));
  jor  g13990(.dina(n14235), .dinb(n14232), .dout(n14236));
  jand g13991(.dina(n14236), .dinb(n14231), .dout(n14237));
  jor  g13992(.dina(n14237), .dinb(n4582), .dout(n14238));
  jand g13993(.dina(n14237), .dinb(n4582), .dout(n14239));
  jxor g13994(.dina(n13651), .dinb(n4902), .dout(n14240));
  jor  g13995(.dina(n14240), .dinb(n14078), .dout(n14241));
  jxor g13996(.dina(n14241), .dinb(n13657), .dout(n14242));
  jor  g13997(.dina(n14242), .dinb(n14239), .dout(n14243));
  jand g13998(.dina(n14243), .dinb(n14238), .dout(n14244));
  jor  g13999(.dina(n14244), .dinb(n4249), .dout(n14245));
  jand g14000(.dina(n14244), .dinb(n4249), .dout(n14246));
  jxor g14001(.dina(n13659), .dinb(n4582), .dout(n14247));
  jor  g14002(.dina(n14247), .dinb(n14078), .dout(n14248));
  jxor g14003(.dina(n14248), .dinb(n13665), .dout(n14249));
  jor  g14004(.dina(n14249), .dinb(n14246), .dout(n14250));
  jand g14005(.dina(n14250), .dinb(n14245), .dout(n14251));
  jor  g14006(.dina(n14251), .dinb(n3955), .dout(n14252));
  jand g14007(.dina(n14251), .dinb(n3955), .dout(n14253));
  jxor g14008(.dina(n13667), .dinb(n4249), .dout(n14254));
  jor  g14009(.dina(n14254), .dinb(n14078), .dout(n14255));
  jxor g14010(.dina(n14255), .dinb(n13980), .dout(n14256));
  jnot g14011(.din(n14256), .dout(n14257));
  jor  g14012(.dina(n14257), .dinb(n14253), .dout(n14258));
  jand g14013(.dina(n14258), .dinb(n14252), .dout(n14259));
  jor  g14014(.dina(n14259), .dinb(n3642), .dout(n14260));
  jand g14015(.dina(n14259), .dinb(n3642), .dout(n14261));
  jxor g14016(.dina(n13674), .dinb(n3955), .dout(n14262));
  jor  g14017(.dina(n14262), .dinb(n14078), .dout(n14263));
  jxor g14018(.dina(n14263), .dinb(n13680), .dout(n14264));
  jor  g14019(.dina(n14264), .dinb(n14261), .dout(n14265));
  jand g14020(.dina(n14265), .dinb(n14260), .dout(n14266));
  jor  g14021(.dina(n14266), .dinb(n3368), .dout(n14267));
  jand g14022(.dina(n14266), .dinb(n3368), .dout(n14268));
  jxor g14023(.dina(n13682), .dinb(n3642), .dout(n14269));
  jor  g14024(.dina(n14269), .dinb(n14078), .dout(n14270));
  jxor g14025(.dina(n14270), .dinb(n13688), .dout(n14271));
  jor  g14026(.dina(n14271), .dinb(n14268), .dout(n14272));
  jand g14027(.dina(n14272), .dinb(n14267), .dout(n14273));
  jor  g14028(.dina(n14273), .dinb(n3089), .dout(n14274));
  jand g14029(.dina(n14273), .dinb(n3089), .dout(n14275));
  jxor g14030(.dina(n13690), .dinb(n3368), .dout(n14276));
  jor  g14031(.dina(n14276), .dinb(n14078), .dout(n14277));
  jxor g14032(.dina(n14277), .dinb(n13696), .dout(n14278));
  jor  g14033(.dina(n14278), .dinb(n14275), .dout(n14279));
  jand g14034(.dina(n14279), .dinb(n14274), .dout(n14280));
  jor  g14035(.dina(n14280), .dinb(n2833), .dout(n14281));
  jand g14036(.dina(n14280), .dinb(n2833), .dout(n14282));
  jxor g14037(.dina(n13698), .dinb(n3089), .dout(n14283));
  jor  g14038(.dina(n14283), .dinb(n14078), .dout(n14284));
  jxor g14039(.dina(n14284), .dinb(n13704), .dout(n14285));
  jor  g14040(.dina(n14285), .dinb(n14282), .dout(n14286));
  jand g14041(.dina(n14286), .dinb(n14281), .dout(n14287));
  jor  g14042(.dina(n14287), .dinb(n2572), .dout(n14288));
  jand g14043(.dina(n14287), .dinb(n2572), .dout(n14289));
  jxor g14044(.dina(n13706), .dinb(n2833), .dout(n14290));
  jor  g14045(.dina(n14290), .dinb(n14078), .dout(n14291));
  jxor g14046(.dina(n14291), .dinb(n13996), .dout(n14292));
  jnot g14047(.din(n14292), .dout(n14293));
  jor  g14048(.dina(n14293), .dinb(n14289), .dout(n14294));
  jand g14049(.dina(n14294), .dinb(n14288), .dout(n14295));
  jor  g14050(.dina(n14295), .dinb(n2345), .dout(n14296));
  jxor g14051(.dina(n13713), .dinb(n2572), .dout(n14297));
  jor  g14052(.dina(n14297), .dinb(n14078), .dout(n14298));
  jxor g14053(.dina(n14298), .dinb(n13879), .dout(n14299));
  jnot g14054(.din(n14299), .dout(n14300));
  jand g14055(.dina(n14295), .dinb(n2345), .dout(n14301));
  jor  g14056(.dina(n14301), .dinb(n14300), .dout(n14302));
  jand g14057(.dina(n14302), .dinb(n14296), .dout(n14303));
  jor  g14058(.dina(n14303), .dinb(n2108), .dout(n14304));
  jand g14059(.dina(n14303), .dinb(n2108), .dout(n14305));
  jxor g14060(.dina(n13720), .dinb(n2345), .dout(n14306));
  jor  g14061(.dina(n14306), .dinb(n14078), .dout(n14307));
  jxor g14062(.dina(n14307), .dinb(n13726), .dout(n14308));
  jor  g14063(.dina(n14308), .dinb(n14305), .dout(n14309));
  jand g14064(.dina(n14309), .dinb(n14304), .dout(n14310));
  jor  g14065(.dina(n14310), .dinb(n1912), .dout(n14311));
  jand g14066(.dina(n14310), .dinb(n1912), .dout(n14312));
  jxor g14067(.dina(n13728), .dinb(n2108), .dout(n14313));
  jor  g14068(.dina(n14313), .dinb(n14078), .dout(n14314));
  jxor g14069(.dina(n14314), .dinb(n14006), .dout(n14315));
  jnot g14070(.din(n14315), .dout(n14316));
  jor  g14071(.dina(n14316), .dinb(n14312), .dout(n14317));
  jand g14072(.dina(n14317), .dinb(n14311), .dout(n14318));
  jor  g14073(.dina(n14318), .dinb(n1699), .dout(n14319));
  jand g14074(.dina(n14318), .dinb(n1699), .dout(n14320));
  jxor g14075(.dina(n13735), .dinb(n1912), .dout(n14321));
  jor  g14076(.dina(n14321), .dinb(n14078), .dout(n14322));
  jxor g14077(.dina(n14322), .dinb(n13741), .dout(n14323));
  jor  g14078(.dina(n14323), .dinb(n14320), .dout(n14324));
  jand g14079(.dina(n14324), .dinb(n14319), .dout(n14325));
  jor  g14080(.dina(n14325), .dinb(n1516), .dout(n14326));
  jand g14081(.dina(n14325), .dinb(n1516), .dout(n14327));
  jxor g14082(.dina(n13743), .dinb(n1699), .dout(n14328));
  jor  g14083(.dina(n14328), .dinb(n14078), .dout(n14329));
  jxor g14084(.dina(n14329), .dinb(n14013), .dout(n14330));
  jnot g14085(.din(n14330), .dout(n14331));
  jor  g14086(.dina(n14331), .dinb(n14327), .dout(n14332));
  jand g14087(.dina(n14332), .dinb(n14326), .dout(n14333));
  jor  g14088(.dina(n14333), .dinb(n1332), .dout(n14334));
  jand g14089(.dina(n14333), .dinb(n1332), .dout(n14335));
  jxor g14090(.dina(n13750), .dinb(n1516), .dout(n14336));
  jor  g14091(.dina(n14336), .dinb(n14078), .dout(n14337));
  jxor g14092(.dina(n14337), .dinb(n13756), .dout(n14338));
  jor  g14093(.dina(n14338), .dinb(n14335), .dout(n14339));
  jand g14094(.dina(n14339), .dinb(n14334), .dout(n14340));
  jor  g14095(.dina(n14340), .dinb(n1173), .dout(n14341));
  jand g14096(.dina(n14340), .dinb(n1173), .dout(n14342));
  jxor g14097(.dina(n13758), .dinb(n1332), .dout(n14343));
  jor  g14098(.dina(n14343), .dinb(n14078), .dout(n14344));
  jxor g14099(.dina(n14344), .dinb(n13764), .dout(n14345));
  jor  g14100(.dina(n14345), .dinb(n14342), .dout(n14346));
  jand g14101(.dina(n14346), .dinb(n14341), .dout(n14347));
  jor  g14102(.dina(n14347), .dinb(n1008), .dout(n14348));
  jand g14103(.dina(n14347), .dinb(n1008), .dout(n14349));
  jxor g14104(.dina(n13766), .dinb(n1173), .dout(n14350));
  jor  g14105(.dina(n14350), .dinb(n14078), .dout(n14351));
  jxor g14106(.dina(n14351), .dinb(n13772), .dout(n14352));
  jor  g14107(.dina(n14352), .dinb(n14349), .dout(n14353));
  jand g14108(.dina(n14353), .dinb(n14348), .dout(n14354));
  jor  g14109(.dina(n14354), .dinb(n884), .dout(n14355));
  jand g14110(.dina(n14354), .dinb(n884), .dout(n14356));
  jxor g14111(.dina(n13774), .dinb(n1008), .dout(n14357));
  jor  g14112(.dina(n14357), .dinb(n14078), .dout(n14358));
  jxor g14113(.dina(n14358), .dinb(n14026), .dout(n14359));
  jnot g14114(.din(n14359), .dout(n14360));
  jor  g14115(.dina(n14360), .dinb(n14356), .dout(n14361));
  jand g14116(.dina(n14361), .dinb(n14355), .dout(n14362));
  jor  g14117(.dina(n14362), .dinb(n743), .dout(n14363));
  jand g14118(.dina(n14362), .dinb(n743), .dout(n14364));
  jxor g14119(.dina(n13781), .dinb(n884), .dout(n14365));
  jor  g14120(.dina(n14365), .dinb(n14078), .dout(n14366));
  jxor g14121(.dina(n14366), .dinb(n13787), .dout(n14367));
  jor  g14122(.dina(n14367), .dinb(n14364), .dout(n14368));
  jand g14123(.dina(n14368), .dinb(n14363), .dout(n14369));
  jor  g14124(.dina(n14369), .dinb(n635), .dout(n14370));
  jand g14125(.dina(n14369), .dinb(n635), .dout(n14371));
  jxor g14126(.dina(n13789), .dinb(n743), .dout(n14372));
  jor  g14127(.dina(n14372), .dinb(n14078), .dout(n14373));
  jxor g14128(.dina(n14373), .dinb(n14033), .dout(n14374));
  jnot g14129(.din(n14374), .dout(n14375));
  jor  g14130(.dina(n14375), .dinb(n14371), .dout(n14376));
  jand g14131(.dina(n14376), .dinb(n14370), .dout(n14377));
  jor  g14132(.dina(n14377), .dinb(n515), .dout(n14378));
  jand g14133(.dina(n14377), .dinb(n515), .dout(n14379));
  jxor g14134(.dina(n13796), .dinb(n635), .dout(n14380));
  jor  g14135(.dina(n14380), .dinb(n14078), .dout(n14381));
  jxor g14136(.dina(n14381), .dinb(n13802), .dout(n14382));
  jor  g14137(.dina(n14382), .dinb(n14379), .dout(n14383));
  jand g14138(.dina(n14383), .dinb(n14378), .dout(n14384));
  jor  g14139(.dina(n14384), .dinb(n443), .dout(n14385));
  jand g14140(.dina(n14384), .dinb(n443), .dout(n14386));
  jxor g14141(.dina(n13804), .dinb(n515), .dout(n14387));
  jor  g14142(.dina(n14387), .dinb(n14078), .dout(n14388));
  jxor g14143(.dina(n14388), .dinb(n14040), .dout(n14389));
  jnot g14144(.din(n14389), .dout(n14390));
  jor  g14145(.dina(n14390), .dinb(n14386), .dout(n14391));
  jand g14146(.dina(n14391), .dinb(n14385), .dout(n14392));
  jor  g14147(.dina(n14392), .dinb(n352), .dout(n14393));
  jand g14148(.dina(n14392), .dinb(n352), .dout(n14394));
  jxor g14149(.dina(n13811), .dinb(n443), .dout(n14395));
  jor  g14150(.dina(n14395), .dinb(n14078), .dout(n14396));
  jxor g14151(.dina(n14396), .dinb(n13817), .dout(n14397));
  jor  g14152(.dina(n14397), .dinb(n14394), .dout(n14398));
  jand g14153(.dina(n14398), .dinb(n14393), .dout(n14399));
  jor  g14154(.dina(n14399), .dinb(n294), .dout(n14400));
  jand g14155(.dina(n14399), .dinb(n294), .dout(n14401));
  jxor g14156(.dina(n13819), .dinb(n352), .dout(n14402));
  jor  g14157(.dina(n14402), .dinb(n14078), .dout(n14403));
  jxor g14158(.dina(n14403), .dinb(n14047), .dout(n14404));
  jnot g14159(.din(n14404), .dout(n14405));
  jor  g14160(.dina(n14405), .dinb(n14401), .dout(n14406));
  jand g14161(.dina(n14406), .dinb(n14400), .dout(n14407));
  jor  g14162(.dina(n14407), .dinb(n239), .dout(n14408));
  jand g14163(.dina(n14407), .dinb(n239), .dout(n14409));
  jxor g14164(.dina(n13826), .dinb(n294), .dout(n14410));
  jor  g14165(.dina(n14410), .dinb(n14078), .dout(n14411));
  jxor g14166(.dina(n14411), .dinb(n14051), .dout(n14412));
  jnot g14167(.din(n14412), .dout(n14413));
  jor  g14168(.dina(n14413), .dinb(n14409), .dout(n14414));
  jand g14169(.dina(n14414), .dinb(n14408), .dout(n14415));
  jor  g14170(.dina(n14415), .dinb(n221), .dout(n14416));
  jand g14171(.dina(n14415), .dinb(n221), .dout(n14417));
  jxor g14172(.dina(n13833), .dinb(n239), .dout(n14418));
  jor  g14173(.dina(n14418), .dinb(n14078), .dout(n14419));
  jxor g14174(.dina(n14419), .dinb(n14055), .dout(n14420));
  jnot g14175(.din(n14420), .dout(n14421));
  jor  g14176(.dina(n14421), .dinb(n14417), .dout(n14422));
  jand g14177(.dina(n14422), .dinb(n14416), .dout(n14423));
  jxor g14178(.dina(n13840), .dinb(n221), .dout(n14424));
  jor  g14179(.dina(n14424), .dinb(n14078), .dout(n14425));
  jxor g14180(.dina(n14425), .dinb(n13846), .dout(n14426));
  jand g14181(.dina(n14426), .dinb(n14423), .dout(n14427));
  jor  g14182(.dina(n14426), .dinb(n14423), .dout(n14429));
  jxor g14183(.dina(n13852), .dinb(n13848), .dout(n14430));
  jnot g14184(.din(n14430), .dout(n14431));
  jand g14185(.dina(n14431), .dinb(asqrt[17] ), .dout(n14432));
  jor  g14186(.dina(n14432), .dinb(n14429), .dout(n14433));
  jand g14187(.dina(n14433), .dinb(n218), .dout(n14434));
  jand g14188(.dina(n14077), .dinb(n14060), .dout(n14435));
  jand g14189(.dina(n14430), .dinb(asqrt[63] ), .dout(n14436));
  jnot g14190(.din(n14436), .dout(n14437));
  jor  g14191(.dina(n14437), .dinb(n14435), .dout(n14438));
  jnot g14192(.din(n14438), .dout(n14439));
  jor  g14193(.dina(n14439), .dinb(n14434), .dout(n14440));
  jor  g14194(.dina(n14440), .dinb(n14427), .dout(asqrt[16] ));
  jnot g14195(.din(a[30] ), .dout(n14443));
  jnot g14196(.din(a[31] ), .dout(n14444));
  jand g14197(.dina(n14444), .dinb(n14443), .dout(n14445));
  jand g14198(.dina(n14445), .dinb(n14080), .dout(n14446));
  jand g14199(.dina(asqrt[16] ), .dinb(a[32] ), .dout(n14447));
  jor  g14200(.dina(n14447), .dinb(n14446), .dout(n14448));
  jand g14201(.dina(n14448), .dinb(asqrt[17] ), .dout(n14449));
  jor  g14202(.dina(n14448), .dinb(asqrt[17] ), .dout(n14450));
  jand g14203(.dina(asqrt[16] ), .dinb(n14080), .dout(n14451));
  jor  g14204(.dina(n14451), .dinb(n14081), .dout(n14452));
  jnot g14205(.din(n14082), .dout(n14453));
  jnot g14206(.din(n14427), .dout(n14454));
  jnot g14207(.din(n14416), .dout(n14456));
  jnot g14208(.din(n14408), .dout(n14457));
  jnot g14209(.din(n14400), .dout(n14458));
  jnot g14210(.din(n14393), .dout(n14459));
  jnot g14211(.din(n14385), .dout(n14460));
  jnot g14212(.din(n14378), .dout(n14461));
  jnot g14213(.din(n14370), .dout(n14462));
  jnot g14214(.din(n14363), .dout(n14463));
  jnot g14215(.din(n14355), .dout(n14464));
  jnot g14216(.din(n14348), .dout(n14465));
  jnot g14217(.din(n14341), .dout(n14466));
  jnot g14218(.din(n14334), .dout(n14467));
  jnot g14219(.din(n14326), .dout(n14468));
  jnot g14220(.din(n14319), .dout(n14469));
  jnot g14221(.din(n14311), .dout(n14470));
  jnot g14222(.din(n14304), .dout(n14471));
  jnot g14223(.din(n14296), .dout(n14472));
  jnot g14224(.din(n14288), .dout(n14473));
  jnot g14225(.din(n14281), .dout(n14474));
  jnot g14226(.din(n14274), .dout(n14475));
  jnot g14227(.din(n14267), .dout(n14476));
  jnot g14228(.din(n14260), .dout(n14477));
  jnot g14229(.din(n14252), .dout(n14478));
  jnot g14230(.din(n14245), .dout(n14479));
  jnot g14231(.din(n14238), .dout(n14480));
  jnot g14232(.din(n14231), .dout(n14481));
  jnot g14233(.din(n14223), .dout(n14482));
  jnot g14234(.din(n14216), .dout(n14483));
  jnot g14235(.din(n14208), .dout(n14484));
  jnot g14236(.din(n14201), .dout(n14485));
  jnot g14237(.din(n14194), .dout(n14486));
  jnot g14238(.din(n14187), .dout(n14487));
  jnot g14239(.din(n14179), .dout(n14488));
  jnot g14240(.din(n14172), .dout(n14489));
  jnot g14241(.din(n14164), .dout(n14490));
  jnot g14242(.din(n14157), .dout(n14491));
  jnot g14243(.din(n14149), .dout(n14492));
  jnot g14244(.din(n14142), .dout(n14493));
  jnot g14245(.din(n14134), .dout(n14494));
  jnot g14246(.din(n14127), .dout(n14495));
  jnot g14247(.din(n14120), .dout(n14496));
  jnot g14248(.din(n14113), .dout(n14497));
  jnot g14249(.din(n14105), .dout(n14498));
  jnot g14250(.din(n14094), .dout(n14499));
  jnot g14251(.din(n14086), .dout(n14500));
  jand g14252(.dina(asqrt[17] ), .dinb(a[34] ), .dout(n14501));
  jor  g14253(.dina(n14083), .dinb(n14501), .dout(n14502));
  jor  g14254(.dina(n14502), .dinb(asqrt[18] ), .dout(n14503));
  jand g14255(.dina(asqrt[17] ), .dinb(n13296), .dout(n14504));
  jor  g14256(.dina(n14504), .dinb(n13297), .dout(n14505));
  jand g14257(.dina(n14097), .dinb(n14505), .dout(n14506));
  jand g14258(.dina(n14506), .dinb(n14503), .dout(n14507));
  jor  g14259(.dina(n14507), .dinb(n14500), .dout(n14508));
  jor  g14260(.dina(n14508), .dinb(asqrt[19] ), .dout(n14509));
  jnot g14261(.din(n14102), .dout(n14510));
  jand g14262(.dina(n14510), .dinb(n14509), .dout(n14511));
  jor  g14263(.dina(n14511), .dinb(n14499), .dout(n14512));
  jor  g14264(.dina(n14512), .dinb(asqrt[20] ), .dout(n14513));
  jand g14265(.dina(n14109), .dinb(n14513), .dout(n14514));
  jor  g14266(.dina(n14514), .dinb(n14498), .dout(n14515));
  jor  g14267(.dina(n14515), .dinb(asqrt[21] ), .dout(n14516));
  jnot g14268(.din(n14117), .dout(n14517));
  jand g14269(.dina(n14517), .dinb(n14516), .dout(n14518));
  jor  g14270(.dina(n14518), .dinb(n14497), .dout(n14519));
  jor  g14271(.dina(n14519), .dinb(asqrt[22] ), .dout(n14520));
  jnot g14272(.din(n14124), .dout(n14521));
  jand g14273(.dina(n14521), .dinb(n14520), .dout(n14522));
  jor  g14274(.dina(n14522), .dinb(n14496), .dout(n14523));
  jor  g14275(.dina(n14523), .dinb(asqrt[23] ), .dout(n14524));
  jnot g14276(.din(n14131), .dout(n14525));
  jand g14277(.dina(n14525), .dinb(n14524), .dout(n14526));
  jor  g14278(.dina(n14526), .dinb(n14495), .dout(n14527));
  jor  g14279(.dina(n14527), .dinb(asqrt[24] ), .dout(n14528));
  jand g14280(.dina(n14138), .dinb(n14528), .dout(n14529));
  jor  g14281(.dina(n14529), .dinb(n14494), .dout(n14530));
  jor  g14282(.dina(n14530), .dinb(asqrt[25] ), .dout(n14531));
  jnot g14283(.din(n14146), .dout(n14532));
  jand g14284(.dina(n14532), .dinb(n14531), .dout(n14533));
  jor  g14285(.dina(n14533), .dinb(n14493), .dout(n14534));
  jor  g14286(.dina(n14534), .dinb(asqrt[26] ), .dout(n14535));
  jand g14287(.dina(n14153), .dinb(n14535), .dout(n14536));
  jor  g14288(.dina(n14536), .dinb(n14492), .dout(n14537));
  jor  g14289(.dina(n14537), .dinb(asqrt[27] ), .dout(n14538));
  jnot g14290(.din(n14161), .dout(n14539));
  jand g14291(.dina(n14539), .dinb(n14538), .dout(n14540));
  jor  g14292(.dina(n14540), .dinb(n14491), .dout(n14541));
  jor  g14293(.dina(n14541), .dinb(asqrt[28] ), .dout(n14542));
  jand g14294(.dina(n14168), .dinb(n14542), .dout(n14543));
  jor  g14295(.dina(n14543), .dinb(n14490), .dout(n14544));
  jor  g14296(.dina(n14544), .dinb(asqrt[29] ), .dout(n14545));
  jnot g14297(.din(n14176), .dout(n14546));
  jand g14298(.dina(n14546), .dinb(n14545), .dout(n14547));
  jor  g14299(.dina(n14547), .dinb(n14489), .dout(n14548));
  jor  g14300(.dina(n14548), .dinb(asqrt[30] ), .dout(n14549));
  jand g14301(.dina(n14183), .dinb(n14549), .dout(n14550));
  jor  g14302(.dina(n14550), .dinb(n14488), .dout(n14551));
  jor  g14303(.dina(n14551), .dinb(asqrt[31] ), .dout(n14552));
  jnot g14304(.din(n14191), .dout(n14553));
  jand g14305(.dina(n14553), .dinb(n14552), .dout(n14554));
  jor  g14306(.dina(n14554), .dinb(n14487), .dout(n14555));
  jor  g14307(.dina(n14555), .dinb(asqrt[32] ), .dout(n14556));
  jnot g14308(.din(n14198), .dout(n14557));
  jand g14309(.dina(n14557), .dinb(n14556), .dout(n14558));
  jor  g14310(.dina(n14558), .dinb(n14486), .dout(n14559));
  jor  g14311(.dina(n14559), .dinb(asqrt[33] ), .dout(n14560));
  jnot g14312(.din(n14205), .dout(n14561));
  jand g14313(.dina(n14561), .dinb(n14560), .dout(n14562));
  jor  g14314(.dina(n14562), .dinb(n14485), .dout(n14563));
  jor  g14315(.dina(n14563), .dinb(asqrt[34] ), .dout(n14564));
  jand g14316(.dina(n14212), .dinb(n14564), .dout(n14565));
  jor  g14317(.dina(n14565), .dinb(n14484), .dout(n14566));
  jor  g14318(.dina(n14566), .dinb(asqrt[35] ), .dout(n14567));
  jnot g14319(.din(n14220), .dout(n14568));
  jand g14320(.dina(n14568), .dinb(n14567), .dout(n14569));
  jor  g14321(.dina(n14569), .dinb(n14483), .dout(n14570));
  jor  g14322(.dina(n14570), .dinb(asqrt[36] ), .dout(n14571));
  jand g14323(.dina(n14227), .dinb(n14571), .dout(n14572));
  jor  g14324(.dina(n14572), .dinb(n14482), .dout(n14573));
  jor  g14325(.dina(n14573), .dinb(asqrt[37] ), .dout(n14574));
  jnot g14326(.din(n14235), .dout(n14575));
  jand g14327(.dina(n14575), .dinb(n14574), .dout(n14576));
  jor  g14328(.dina(n14576), .dinb(n14481), .dout(n14577));
  jor  g14329(.dina(n14577), .dinb(asqrt[38] ), .dout(n14578));
  jnot g14330(.din(n14242), .dout(n14579));
  jand g14331(.dina(n14579), .dinb(n14578), .dout(n14580));
  jor  g14332(.dina(n14580), .dinb(n14480), .dout(n14581));
  jor  g14333(.dina(n14581), .dinb(asqrt[39] ), .dout(n14582));
  jnot g14334(.din(n14249), .dout(n14583));
  jand g14335(.dina(n14583), .dinb(n14582), .dout(n14584));
  jor  g14336(.dina(n14584), .dinb(n14479), .dout(n14585));
  jor  g14337(.dina(n14585), .dinb(asqrt[40] ), .dout(n14586));
  jand g14338(.dina(n14256), .dinb(n14586), .dout(n14587));
  jor  g14339(.dina(n14587), .dinb(n14478), .dout(n14588));
  jor  g14340(.dina(n14588), .dinb(asqrt[41] ), .dout(n14589));
  jnot g14341(.din(n14264), .dout(n14590));
  jand g14342(.dina(n14590), .dinb(n14589), .dout(n14591));
  jor  g14343(.dina(n14591), .dinb(n14477), .dout(n14592));
  jor  g14344(.dina(n14592), .dinb(asqrt[42] ), .dout(n14593));
  jnot g14345(.din(n14271), .dout(n14594));
  jand g14346(.dina(n14594), .dinb(n14593), .dout(n14595));
  jor  g14347(.dina(n14595), .dinb(n14476), .dout(n14596));
  jor  g14348(.dina(n14596), .dinb(asqrt[43] ), .dout(n14597));
  jnot g14349(.din(n14278), .dout(n14598));
  jand g14350(.dina(n14598), .dinb(n14597), .dout(n14599));
  jor  g14351(.dina(n14599), .dinb(n14475), .dout(n14600));
  jor  g14352(.dina(n14600), .dinb(asqrt[44] ), .dout(n14601));
  jnot g14353(.din(n14285), .dout(n14602));
  jand g14354(.dina(n14602), .dinb(n14601), .dout(n14603));
  jor  g14355(.dina(n14603), .dinb(n14474), .dout(n14604));
  jor  g14356(.dina(n14604), .dinb(asqrt[45] ), .dout(n14605));
  jand g14357(.dina(n14292), .dinb(n14605), .dout(n14606));
  jor  g14358(.dina(n14606), .dinb(n14473), .dout(n14607));
  jor  g14359(.dina(n14607), .dinb(asqrt[46] ), .dout(n14608));
  jand g14360(.dina(n14608), .dinb(n14299), .dout(n14609));
  jor  g14361(.dina(n14609), .dinb(n14472), .dout(n14610));
  jor  g14362(.dina(n14610), .dinb(asqrt[47] ), .dout(n14611));
  jnot g14363(.din(n14308), .dout(n14612));
  jand g14364(.dina(n14612), .dinb(n14611), .dout(n14613));
  jor  g14365(.dina(n14613), .dinb(n14471), .dout(n14614));
  jor  g14366(.dina(n14614), .dinb(asqrt[48] ), .dout(n14615));
  jand g14367(.dina(n14315), .dinb(n14615), .dout(n14616));
  jor  g14368(.dina(n14616), .dinb(n14470), .dout(n14617));
  jor  g14369(.dina(n14617), .dinb(asqrt[49] ), .dout(n14618));
  jnot g14370(.din(n14323), .dout(n14619));
  jand g14371(.dina(n14619), .dinb(n14618), .dout(n14620));
  jor  g14372(.dina(n14620), .dinb(n14469), .dout(n14621));
  jor  g14373(.dina(n14621), .dinb(asqrt[50] ), .dout(n14622));
  jand g14374(.dina(n14330), .dinb(n14622), .dout(n14623));
  jor  g14375(.dina(n14623), .dinb(n14468), .dout(n14624));
  jor  g14376(.dina(n14624), .dinb(asqrt[51] ), .dout(n14625));
  jnot g14377(.din(n14338), .dout(n14626));
  jand g14378(.dina(n14626), .dinb(n14625), .dout(n14627));
  jor  g14379(.dina(n14627), .dinb(n14467), .dout(n14628));
  jor  g14380(.dina(n14628), .dinb(asqrt[52] ), .dout(n14629));
  jnot g14381(.din(n14345), .dout(n14630));
  jand g14382(.dina(n14630), .dinb(n14629), .dout(n14631));
  jor  g14383(.dina(n14631), .dinb(n14466), .dout(n14632));
  jor  g14384(.dina(n14632), .dinb(asqrt[53] ), .dout(n14633));
  jnot g14385(.din(n14352), .dout(n14634));
  jand g14386(.dina(n14634), .dinb(n14633), .dout(n14635));
  jor  g14387(.dina(n14635), .dinb(n14465), .dout(n14636));
  jor  g14388(.dina(n14636), .dinb(asqrt[54] ), .dout(n14637));
  jand g14389(.dina(n14359), .dinb(n14637), .dout(n14638));
  jor  g14390(.dina(n14638), .dinb(n14464), .dout(n14639));
  jor  g14391(.dina(n14639), .dinb(asqrt[55] ), .dout(n14640));
  jnot g14392(.din(n14367), .dout(n14641));
  jand g14393(.dina(n14641), .dinb(n14640), .dout(n14642));
  jor  g14394(.dina(n14642), .dinb(n14463), .dout(n14643));
  jor  g14395(.dina(n14643), .dinb(asqrt[56] ), .dout(n14644));
  jand g14396(.dina(n14374), .dinb(n14644), .dout(n14645));
  jor  g14397(.dina(n14645), .dinb(n14462), .dout(n14646));
  jor  g14398(.dina(n14646), .dinb(asqrt[57] ), .dout(n14647));
  jnot g14399(.din(n14382), .dout(n14648));
  jand g14400(.dina(n14648), .dinb(n14647), .dout(n14649));
  jor  g14401(.dina(n14649), .dinb(n14461), .dout(n14650));
  jor  g14402(.dina(n14650), .dinb(asqrt[58] ), .dout(n14651));
  jand g14403(.dina(n14389), .dinb(n14651), .dout(n14652));
  jor  g14404(.dina(n14652), .dinb(n14460), .dout(n14653));
  jor  g14405(.dina(n14653), .dinb(asqrt[59] ), .dout(n14654));
  jnot g14406(.din(n14397), .dout(n14655));
  jand g14407(.dina(n14655), .dinb(n14654), .dout(n14656));
  jor  g14408(.dina(n14656), .dinb(n14459), .dout(n14657));
  jor  g14409(.dina(n14657), .dinb(asqrt[60] ), .dout(n14658));
  jand g14410(.dina(n14404), .dinb(n14658), .dout(n14659));
  jor  g14411(.dina(n14659), .dinb(n14458), .dout(n14660));
  jor  g14412(.dina(n14660), .dinb(asqrt[61] ), .dout(n14661));
  jand g14413(.dina(n14412), .dinb(n14661), .dout(n14662));
  jor  g14414(.dina(n14662), .dinb(n14457), .dout(n14663));
  jor  g14415(.dina(n14663), .dinb(asqrt[62] ), .dout(n14664));
  jand g14416(.dina(n14420), .dinb(n14664), .dout(n14665));
  jor  g14417(.dina(n14665), .dinb(n14456), .dout(n14666));
  jnot g14418(.din(n14426), .dout(n14667));
  jand g14419(.dina(n14667), .dinb(n14666), .dout(n14668));
  jnot g14420(.din(n14432), .dout(n14669));
  jand g14421(.dina(n14669), .dinb(n14668), .dout(n14670));
  jor  g14422(.dina(n14670), .dinb(asqrt[63] ), .dout(n14671));
  jand g14423(.dina(n14438), .dinb(n14671), .dout(n14672));
  jand g14424(.dina(n14672), .dinb(n14454), .dout(n14674));
  jor  g14425(.dina(n14674), .dinb(n14453), .dout(n14675));
  jand g14426(.dina(n14675), .dinb(n14452), .dout(n14676));
  jand g14427(.dina(n14676), .dinb(n14450), .dout(n14677));
  jor  g14428(.dina(n14677), .dinb(n14449), .dout(n14678));
  jand g14429(.dina(n14678), .dinb(asqrt[18] ), .dout(n14679));
  jor  g14430(.dina(n14678), .dinb(asqrt[18] ), .dout(n14680));
  jand g14431(.dina(asqrt[16] ), .dinb(n14082), .dout(n14681));
  jand g14432(.dina(n14437), .dinb(n14454), .dout(n14682));
  jand g14433(.dina(n14682), .dinb(n14671), .dout(n14683));
  jand g14434(.dina(n14683), .dinb(asqrt[17] ), .dout(n14684));
  jor  g14435(.dina(n14684), .dinb(n14681), .dout(n14685));
  jxor g14436(.dina(n14685), .dinb(a[34] ), .dout(n14686));
  jnot g14437(.din(n14686), .dout(n14687));
  jand g14438(.dina(n14687), .dinb(n14680), .dout(n14688));
  jor  g14439(.dina(n14688), .dinb(n14679), .dout(n14689));
  jand g14440(.dina(n14689), .dinb(asqrt[19] ), .dout(n14690));
  jor  g14441(.dina(n14689), .dinb(asqrt[19] ), .dout(n14691));
  jxor g14442(.dina(n14085), .dinb(n13515), .dout(n14692));
  jand g14443(.dina(n14692), .dinb(asqrt[16] ), .dout(n14693));
  jxor g14444(.dina(n14693), .dinb(n14506), .dout(n14694));
  jand g14445(.dina(n14694), .dinb(n14691), .dout(n14695));
  jor  g14446(.dina(n14695), .dinb(n14690), .dout(n14696));
  jand g14447(.dina(n14696), .dinb(asqrt[20] ), .dout(n14697));
  jor  g14448(.dina(n14696), .dinb(asqrt[20] ), .dout(n14698));
  jxor g14449(.dina(n14093), .dinb(n12947), .dout(n14699));
  jand g14450(.dina(n14699), .dinb(asqrt[16] ), .dout(n14700));
  jxor g14451(.dina(n14700), .dinb(n14102), .dout(n14701));
  jnot g14452(.din(n14701), .dout(n14702));
  jand g14453(.dina(n14702), .dinb(n14698), .dout(n14703));
  jor  g14454(.dina(n14703), .dinb(n14697), .dout(n14704));
  jand g14455(.dina(n14704), .dinb(asqrt[21] ), .dout(n14705));
  jor  g14456(.dina(n14704), .dinb(asqrt[21] ), .dout(n14706));
  jxor g14457(.dina(n14104), .dinb(n12410), .dout(n14707));
  jand g14458(.dina(n14707), .dinb(asqrt[16] ), .dout(n14708));
  jxor g14459(.dina(n14708), .dinb(n14109), .dout(n14709));
  jand g14460(.dina(n14709), .dinb(n14706), .dout(n14710));
  jor  g14461(.dina(n14710), .dinb(n14705), .dout(n14711));
  jand g14462(.dina(n14711), .dinb(asqrt[22] ), .dout(n14712));
  jor  g14463(.dina(n14711), .dinb(asqrt[22] ), .dout(n14713));
  jxor g14464(.dina(n14112), .dinb(n11858), .dout(n14714));
  jand g14465(.dina(n14714), .dinb(asqrt[16] ), .dout(n14715));
  jxor g14466(.dina(n14715), .dinb(n14117), .dout(n14716));
  jnot g14467(.din(n14716), .dout(n14717));
  jand g14468(.dina(n14717), .dinb(n14713), .dout(n14718));
  jor  g14469(.dina(n14718), .dinb(n14712), .dout(n14719));
  jand g14470(.dina(n14719), .dinb(asqrt[23] ), .dout(n14720));
  jor  g14471(.dina(n14719), .dinb(asqrt[23] ), .dout(n14721));
  jxor g14472(.dina(n14119), .dinb(n11347), .dout(n14722));
  jand g14473(.dina(n14722), .dinb(asqrt[16] ), .dout(n14723));
  jxor g14474(.dina(n14723), .dinb(n14124), .dout(n14724));
  jnot g14475(.din(n14724), .dout(n14725));
  jand g14476(.dina(n14725), .dinb(n14721), .dout(n14726));
  jor  g14477(.dina(n14726), .dinb(n14720), .dout(n14727));
  jand g14478(.dina(n14727), .dinb(asqrt[24] ), .dout(n14728));
  jor  g14479(.dina(n14727), .dinb(asqrt[24] ), .dout(n14729));
  jxor g14480(.dina(n14126), .dinb(n10824), .dout(n14730));
  jand g14481(.dina(n14730), .dinb(asqrt[16] ), .dout(n14731));
  jxor g14482(.dina(n14731), .dinb(n14131), .dout(n14732));
  jnot g14483(.din(n14732), .dout(n14733));
  jand g14484(.dina(n14733), .dinb(n14729), .dout(n14734));
  jor  g14485(.dina(n14734), .dinb(n14728), .dout(n14735));
  jand g14486(.dina(n14735), .dinb(asqrt[25] ), .dout(n14736));
  jor  g14487(.dina(n14735), .dinb(asqrt[25] ), .dout(n14737));
  jxor g14488(.dina(n14133), .dinb(n10328), .dout(n14738));
  jand g14489(.dina(n14738), .dinb(asqrt[16] ), .dout(n14739));
  jxor g14490(.dina(n14739), .dinb(n14138), .dout(n14740));
  jand g14491(.dina(n14740), .dinb(n14737), .dout(n14741));
  jor  g14492(.dina(n14741), .dinb(n14736), .dout(n14742));
  jand g14493(.dina(n14742), .dinb(asqrt[26] ), .dout(n14743));
  jor  g14494(.dina(n14742), .dinb(asqrt[26] ), .dout(n14744));
  jxor g14495(.dina(n14141), .dinb(n9832), .dout(n14745));
  jand g14496(.dina(n14745), .dinb(asqrt[16] ), .dout(n14746));
  jxor g14497(.dina(n14746), .dinb(n14146), .dout(n14747));
  jnot g14498(.din(n14747), .dout(n14748));
  jand g14499(.dina(n14748), .dinb(n14744), .dout(n14749));
  jor  g14500(.dina(n14749), .dinb(n14743), .dout(n14750));
  jand g14501(.dina(n14750), .dinb(asqrt[27] ), .dout(n14751));
  jor  g14502(.dina(n14750), .dinb(asqrt[27] ), .dout(n14752));
  jxor g14503(.dina(n14148), .dinb(n9369), .dout(n14753));
  jand g14504(.dina(n14753), .dinb(asqrt[16] ), .dout(n14754));
  jxor g14505(.dina(n14754), .dinb(n14153), .dout(n14755));
  jand g14506(.dina(n14755), .dinb(n14752), .dout(n14756));
  jor  g14507(.dina(n14756), .dinb(n14751), .dout(n14757));
  jand g14508(.dina(n14757), .dinb(asqrt[28] ), .dout(n14758));
  jor  g14509(.dina(n14757), .dinb(asqrt[28] ), .dout(n14759));
  jxor g14510(.dina(n14156), .dinb(n8890), .dout(n14760));
  jand g14511(.dina(n14760), .dinb(asqrt[16] ), .dout(n14761));
  jxor g14512(.dina(n14761), .dinb(n14161), .dout(n14762));
  jnot g14513(.din(n14762), .dout(n14763));
  jand g14514(.dina(n14763), .dinb(n14759), .dout(n14764));
  jor  g14515(.dina(n14764), .dinb(n14758), .dout(n14765));
  jand g14516(.dina(n14765), .dinb(asqrt[29] ), .dout(n14766));
  jor  g14517(.dina(n14765), .dinb(asqrt[29] ), .dout(n14767));
  jxor g14518(.dina(n14163), .dinb(n8449), .dout(n14768));
  jand g14519(.dina(n14768), .dinb(asqrt[16] ), .dout(n14769));
  jxor g14520(.dina(n14769), .dinb(n14168), .dout(n14770));
  jand g14521(.dina(n14770), .dinb(n14767), .dout(n14771));
  jor  g14522(.dina(n14771), .dinb(n14766), .dout(n14772));
  jand g14523(.dina(n14772), .dinb(asqrt[30] ), .dout(n14773));
  jor  g14524(.dina(n14772), .dinb(asqrt[30] ), .dout(n14774));
  jxor g14525(.dina(n14171), .dinb(n8003), .dout(n14775));
  jand g14526(.dina(n14775), .dinb(asqrt[16] ), .dout(n14776));
  jxor g14527(.dina(n14776), .dinb(n14176), .dout(n14777));
  jnot g14528(.din(n14777), .dout(n14778));
  jand g14529(.dina(n14778), .dinb(n14774), .dout(n14779));
  jor  g14530(.dina(n14779), .dinb(n14773), .dout(n14780));
  jand g14531(.dina(n14780), .dinb(asqrt[31] ), .dout(n14781));
  jor  g14532(.dina(n14780), .dinb(asqrt[31] ), .dout(n14782));
  jxor g14533(.dina(n14178), .dinb(n7581), .dout(n14783));
  jand g14534(.dina(n14783), .dinb(asqrt[16] ), .dout(n14784));
  jxor g14535(.dina(n14784), .dinb(n14183), .dout(n14785));
  jand g14536(.dina(n14785), .dinb(n14782), .dout(n14786));
  jor  g14537(.dina(n14786), .dinb(n14781), .dout(n14787));
  jand g14538(.dina(n14787), .dinb(asqrt[32] ), .dout(n14788));
  jor  g14539(.dina(n14787), .dinb(asqrt[32] ), .dout(n14789));
  jxor g14540(.dina(n14186), .dinb(n7154), .dout(n14790));
  jand g14541(.dina(n14790), .dinb(asqrt[16] ), .dout(n14791));
  jxor g14542(.dina(n14791), .dinb(n14191), .dout(n14792));
  jnot g14543(.din(n14792), .dout(n14793));
  jand g14544(.dina(n14793), .dinb(n14789), .dout(n14794));
  jor  g14545(.dina(n14794), .dinb(n14788), .dout(n14795));
  jand g14546(.dina(n14795), .dinb(asqrt[33] ), .dout(n14796));
  jor  g14547(.dina(n14795), .dinb(asqrt[33] ), .dout(n14797));
  jxor g14548(.dina(n14193), .dinb(n6758), .dout(n14798));
  jand g14549(.dina(n14798), .dinb(asqrt[16] ), .dout(n14799));
  jxor g14550(.dina(n14799), .dinb(n14198), .dout(n14800));
  jnot g14551(.din(n14800), .dout(n14801));
  jand g14552(.dina(n14801), .dinb(n14797), .dout(n14802));
  jor  g14553(.dina(n14802), .dinb(n14796), .dout(n14803));
  jand g14554(.dina(n14803), .dinb(asqrt[34] ), .dout(n14804));
  jor  g14555(.dina(n14803), .dinb(asqrt[34] ), .dout(n14805));
  jxor g14556(.dina(n14200), .dinb(n6357), .dout(n14806));
  jand g14557(.dina(n14806), .dinb(asqrt[16] ), .dout(n14807));
  jxor g14558(.dina(n14807), .dinb(n14205), .dout(n14808));
  jnot g14559(.din(n14808), .dout(n14809));
  jand g14560(.dina(n14809), .dinb(n14805), .dout(n14810));
  jor  g14561(.dina(n14810), .dinb(n14804), .dout(n14811));
  jand g14562(.dina(n14811), .dinb(asqrt[35] ), .dout(n14812));
  jor  g14563(.dina(n14811), .dinb(asqrt[35] ), .dout(n14813));
  jxor g14564(.dina(n14207), .dinb(n5989), .dout(n14814));
  jand g14565(.dina(n14814), .dinb(asqrt[16] ), .dout(n14815));
  jxor g14566(.dina(n14815), .dinb(n14212), .dout(n14816));
  jand g14567(.dina(n14816), .dinb(n14813), .dout(n14817));
  jor  g14568(.dina(n14817), .dinb(n14812), .dout(n14818));
  jand g14569(.dina(n14818), .dinb(asqrt[36] ), .dout(n14819));
  jor  g14570(.dina(n14818), .dinb(asqrt[36] ), .dout(n14820));
  jxor g14571(.dina(n14215), .dinb(n5606), .dout(n14821));
  jand g14572(.dina(n14821), .dinb(asqrt[16] ), .dout(n14822));
  jxor g14573(.dina(n14822), .dinb(n14220), .dout(n14823));
  jnot g14574(.din(n14823), .dout(n14824));
  jand g14575(.dina(n14824), .dinb(n14820), .dout(n14825));
  jor  g14576(.dina(n14825), .dinb(n14819), .dout(n14826));
  jand g14577(.dina(n14826), .dinb(asqrt[37] ), .dout(n14827));
  jor  g14578(.dina(n14826), .dinb(asqrt[37] ), .dout(n14828));
  jxor g14579(.dina(n14222), .dinb(n5259), .dout(n14829));
  jand g14580(.dina(n14829), .dinb(asqrt[16] ), .dout(n14830));
  jxor g14581(.dina(n14830), .dinb(n14227), .dout(n14831));
  jand g14582(.dina(n14831), .dinb(n14828), .dout(n14832));
  jor  g14583(.dina(n14832), .dinb(n14827), .dout(n14833));
  jand g14584(.dina(n14833), .dinb(asqrt[38] ), .dout(n14834));
  jor  g14585(.dina(n14833), .dinb(asqrt[38] ), .dout(n14835));
  jxor g14586(.dina(n14230), .dinb(n4902), .dout(n14836));
  jand g14587(.dina(n14836), .dinb(asqrt[16] ), .dout(n14837));
  jxor g14588(.dina(n14837), .dinb(n14235), .dout(n14838));
  jnot g14589(.din(n14838), .dout(n14839));
  jand g14590(.dina(n14839), .dinb(n14835), .dout(n14840));
  jor  g14591(.dina(n14840), .dinb(n14834), .dout(n14841));
  jand g14592(.dina(n14841), .dinb(asqrt[39] ), .dout(n14842));
  jor  g14593(.dina(n14841), .dinb(asqrt[39] ), .dout(n14843));
  jxor g14594(.dina(n14237), .dinb(n4582), .dout(n14844));
  jand g14595(.dina(n14844), .dinb(asqrt[16] ), .dout(n14845));
  jxor g14596(.dina(n14845), .dinb(n14242), .dout(n14846));
  jnot g14597(.din(n14846), .dout(n14847));
  jand g14598(.dina(n14847), .dinb(n14843), .dout(n14848));
  jor  g14599(.dina(n14848), .dinb(n14842), .dout(n14849));
  jand g14600(.dina(n14849), .dinb(asqrt[40] ), .dout(n14850));
  jor  g14601(.dina(n14849), .dinb(asqrt[40] ), .dout(n14851));
  jxor g14602(.dina(n14244), .dinb(n4249), .dout(n14852));
  jand g14603(.dina(n14852), .dinb(asqrt[16] ), .dout(n14853));
  jxor g14604(.dina(n14853), .dinb(n14249), .dout(n14854));
  jnot g14605(.din(n14854), .dout(n14855));
  jand g14606(.dina(n14855), .dinb(n14851), .dout(n14856));
  jor  g14607(.dina(n14856), .dinb(n14850), .dout(n14857));
  jand g14608(.dina(n14857), .dinb(asqrt[41] ), .dout(n14858));
  jor  g14609(.dina(n14857), .dinb(asqrt[41] ), .dout(n14859));
  jxor g14610(.dina(n14251), .dinb(n3955), .dout(n14860));
  jand g14611(.dina(n14860), .dinb(asqrt[16] ), .dout(n14861));
  jxor g14612(.dina(n14861), .dinb(n14256), .dout(n14862));
  jand g14613(.dina(n14862), .dinb(n14859), .dout(n14863));
  jor  g14614(.dina(n14863), .dinb(n14858), .dout(n14864));
  jand g14615(.dina(n14864), .dinb(asqrt[42] ), .dout(n14865));
  jor  g14616(.dina(n14864), .dinb(asqrt[42] ), .dout(n14866));
  jxor g14617(.dina(n14259), .dinb(n3642), .dout(n14867));
  jand g14618(.dina(n14867), .dinb(asqrt[16] ), .dout(n14868));
  jxor g14619(.dina(n14868), .dinb(n14264), .dout(n14869));
  jnot g14620(.din(n14869), .dout(n14870));
  jand g14621(.dina(n14870), .dinb(n14866), .dout(n14871));
  jor  g14622(.dina(n14871), .dinb(n14865), .dout(n14872));
  jand g14623(.dina(n14872), .dinb(asqrt[43] ), .dout(n14873));
  jor  g14624(.dina(n14872), .dinb(asqrt[43] ), .dout(n14874));
  jxor g14625(.dina(n14266), .dinb(n3368), .dout(n14875));
  jand g14626(.dina(n14875), .dinb(asqrt[16] ), .dout(n14876));
  jxor g14627(.dina(n14876), .dinb(n14594), .dout(n14877));
  jand g14628(.dina(n14877), .dinb(n14874), .dout(n14878));
  jor  g14629(.dina(n14878), .dinb(n14873), .dout(n14879));
  jand g14630(.dina(n14879), .dinb(asqrt[44] ), .dout(n14880));
  jor  g14631(.dina(n14879), .dinb(asqrt[44] ), .dout(n14881));
  jxor g14632(.dina(n14273), .dinb(n3089), .dout(n14882));
  jand g14633(.dina(n14882), .dinb(asqrt[16] ), .dout(n14883));
  jxor g14634(.dina(n14883), .dinb(n14278), .dout(n14884));
  jnot g14635(.din(n14884), .dout(n14885));
  jand g14636(.dina(n14885), .dinb(n14881), .dout(n14886));
  jor  g14637(.dina(n14886), .dinb(n14880), .dout(n14887));
  jand g14638(.dina(n14887), .dinb(asqrt[45] ), .dout(n14888));
  jor  g14639(.dina(n14887), .dinb(asqrt[45] ), .dout(n14889));
  jxor g14640(.dina(n14280), .dinb(n2833), .dout(n14890));
  jand g14641(.dina(n14890), .dinb(asqrt[16] ), .dout(n14891));
  jxor g14642(.dina(n14891), .dinb(n14285), .dout(n14892));
  jnot g14643(.din(n14892), .dout(n14893));
  jand g14644(.dina(n14893), .dinb(n14889), .dout(n14894));
  jor  g14645(.dina(n14894), .dinb(n14888), .dout(n14895));
  jand g14646(.dina(n14895), .dinb(asqrt[46] ), .dout(n14896));
  jor  g14647(.dina(n14895), .dinb(asqrt[46] ), .dout(n14897));
  jxor g14648(.dina(n14287), .dinb(n2572), .dout(n14898));
  jand g14649(.dina(n14898), .dinb(asqrt[16] ), .dout(n14899));
  jxor g14650(.dina(n14899), .dinb(n14292), .dout(n14900));
  jand g14651(.dina(n14900), .dinb(n14897), .dout(n14901));
  jor  g14652(.dina(n14901), .dinb(n14896), .dout(n14902));
  jand g14653(.dina(n14902), .dinb(asqrt[47] ), .dout(n14903));
  jxor g14654(.dina(n14295), .dinb(n2345), .dout(n14904));
  jand g14655(.dina(n14904), .dinb(asqrt[16] ), .dout(n14905));
  jxor g14656(.dina(n14905), .dinb(n14299), .dout(n14906));
  jor  g14657(.dina(n14902), .dinb(asqrt[47] ), .dout(n14907));
  jand g14658(.dina(n14907), .dinb(n14906), .dout(n14908));
  jor  g14659(.dina(n14908), .dinb(n14903), .dout(n14909));
  jand g14660(.dina(n14909), .dinb(asqrt[48] ), .dout(n14910));
  jor  g14661(.dina(n14909), .dinb(asqrt[48] ), .dout(n14911));
  jxor g14662(.dina(n14303), .dinb(n2108), .dout(n14912));
  jand g14663(.dina(n14912), .dinb(asqrt[16] ), .dout(n14913));
  jxor g14664(.dina(n14913), .dinb(n14308), .dout(n14914));
  jnot g14665(.din(n14914), .dout(n14915));
  jand g14666(.dina(n14915), .dinb(n14911), .dout(n14916));
  jor  g14667(.dina(n14916), .dinb(n14910), .dout(n14917));
  jand g14668(.dina(n14917), .dinb(asqrt[49] ), .dout(n14918));
  jor  g14669(.dina(n14917), .dinb(asqrt[49] ), .dout(n14919));
  jxor g14670(.dina(n14310), .dinb(n1912), .dout(n14920));
  jand g14671(.dina(n14920), .dinb(asqrt[16] ), .dout(n14921));
  jxor g14672(.dina(n14921), .dinb(n14315), .dout(n14922));
  jand g14673(.dina(n14922), .dinb(n14919), .dout(n14923));
  jor  g14674(.dina(n14923), .dinb(n14918), .dout(n14924));
  jand g14675(.dina(n14924), .dinb(asqrt[50] ), .dout(n14925));
  jor  g14676(.dina(n14924), .dinb(asqrt[50] ), .dout(n14926));
  jxor g14677(.dina(n14318), .dinb(n1699), .dout(n14927));
  jand g14678(.dina(n14927), .dinb(asqrt[16] ), .dout(n14928));
  jxor g14679(.dina(n14928), .dinb(n14323), .dout(n14929));
  jnot g14680(.din(n14929), .dout(n14930));
  jand g14681(.dina(n14930), .dinb(n14926), .dout(n14931));
  jor  g14682(.dina(n14931), .dinb(n14925), .dout(n14932));
  jand g14683(.dina(n14932), .dinb(asqrt[51] ), .dout(n14933));
  jor  g14684(.dina(n14932), .dinb(asqrt[51] ), .dout(n14934));
  jxor g14685(.dina(n14325), .dinb(n1516), .dout(n14935));
  jand g14686(.dina(n14935), .dinb(asqrt[16] ), .dout(n14936));
  jxor g14687(.dina(n14936), .dinb(n14330), .dout(n14937));
  jand g14688(.dina(n14937), .dinb(n14934), .dout(n14938));
  jor  g14689(.dina(n14938), .dinb(n14933), .dout(n14939));
  jand g14690(.dina(n14939), .dinb(asqrt[52] ), .dout(n14940));
  jor  g14691(.dina(n14939), .dinb(asqrt[52] ), .dout(n14941));
  jxor g14692(.dina(n14333), .dinb(n1332), .dout(n14942));
  jand g14693(.dina(n14942), .dinb(asqrt[16] ), .dout(n14943));
  jxor g14694(.dina(n14943), .dinb(n14338), .dout(n14944));
  jnot g14695(.din(n14944), .dout(n14945));
  jand g14696(.dina(n14945), .dinb(n14941), .dout(n14946));
  jor  g14697(.dina(n14946), .dinb(n14940), .dout(n14947));
  jand g14698(.dina(n14947), .dinb(asqrt[53] ), .dout(n14948));
  jor  g14699(.dina(n14947), .dinb(asqrt[53] ), .dout(n14949));
  jxor g14700(.dina(n14340), .dinb(n1173), .dout(n14950));
  jand g14701(.dina(n14950), .dinb(asqrt[16] ), .dout(n14951));
  jxor g14702(.dina(n14951), .dinb(n14345), .dout(n14952));
  jnot g14703(.din(n14952), .dout(n14953));
  jand g14704(.dina(n14953), .dinb(n14949), .dout(n14954));
  jor  g14705(.dina(n14954), .dinb(n14948), .dout(n14955));
  jand g14706(.dina(n14955), .dinb(asqrt[54] ), .dout(n14956));
  jor  g14707(.dina(n14955), .dinb(asqrt[54] ), .dout(n14957));
  jxor g14708(.dina(n14347), .dinb(n1008), .dout(n14958));
  jand g14709(.dina(n14958), .dinb(asqrt[16] ), .dout(n14959));
  jxor g14710(.dina(n14959), .dinb(n14352), .dout(n14960));
  jnot g14711(.din(n14960), .dout(n14961));
  jand g14712(.dina(n14961), .dinb(n14957), .dout(n14962));
  jor  g14713(.dina(n14962), .dinb(n14956), .dout(n14963));
  jand g14714(.dina(n14963), .dinb(asqrt[55] ), .dout(n14964));
  jor  g14715(.dina(n14963), .dinb(asqrt[55] ), .dout(n14965));
  jxor g14716(.dina(n14354), .dinb(n884), .dout(n14966));
  jand g14717(.dina(n14966), .dinb(asqrt[16] ), .dout(n14967));
  jxor g14718(.dina(n14967), .dinb(n14359), .dout(n14968));
  jand g14719(.dina(n14968), .dinb(n14965), .dout(n14969));
  jor  g14720(.dina(n14969), .dinb(n14964), .dout(n14970));
  jand g14721(.dina(n14970), .dinb(asqrt[56] ), .dout(n14971));
  jor  g14722(.dina(n14970), .dinb(asqrt[56] ), .dout(n14972));
  jxor g14723(.dina(n14362), .dinb(n743), .dout(n14973));
  jand g14724(.dina(n14973), .dinb(asqrt[16] ), .dout(n14974));
  jxor g14725(.dina(n14974), .dinb(n14367), .dout(n14975));
  jnot g14726(.din(n14975), .dout(n14976));
  jand g14727(.dina(n14976), .dinb(n14972), .dout(n14977));
  jor  g14728(.dina(n14977), .dinb(n14971), .dout(n14978));
  jand g14729(.dina(n14978), .dinb(asqrt[57] ), .dout(n14979));
  jor  g14730(.dina(n14978), .dinb(asqrt[57] ), .dout(n14980));
  jxor g14731(.dina(n14369), .dinb(n635), .dout(n14981));
  jand g14732(.dina(n14981), .dinb(asqrt[16] ), .dout(n14982));
  jxor g14733(.dina(n14982), .dinb(n14374), .dout(n14983));
  jand g14734(.dina(n14983), .dinb(n14980), .dout(n14984));
  jor  g14735(.dina(n14984), .dinb(n14979), .dout(n14985));
  jand g14736(.dina(n14985), .dinb(asqrt[58] ), .dout(n14986));
  jor  g14737(.dina(n14985), .dinb(asqrt[58] ), .dout(n14987));
  jxor g14738(.dina(n14377), .dinb(n515), .dout(n14988));
  jand g14739(.dina(n14988), .dinb(asqrt[16] ), .dout(n14989));
  jxor g14740(.dina(n14989), .dinb(n14382), .dout(n14990));
  jnot g14741(.din(n14990), .dout(n14991));
  jand g14742(.dina(n14991), .dinb(n14987), .dout(n14992));
  jor  g14743(.dina(n14992), .dinb(n14986), .dout(n14993));
  jand g14744(.dina(n14993), .dinb(asqrt[59] ), .dout(n14994));
  jor  g14745(.dina(n14993), .dinb(asqrt[59] ), .dout(n14995));
  jxor g14746(.dina(n14384), .dinb(n443), .dout(n14996));
  jand g14747(.dina(n14996), .dinb(asqrt[16] ), .dout(n14997));
  jxor g14748(.dina(n14997), .dinb(n14389), .dout(n14998));
  jand g14749(.dina(n14998), .dinb(n14995), .dout(n14999));
  jor  g14750(.dina(n14999), .dinb(n14994), .dout(n15000));
  jand g14751(.dina(n15000), .dinb(asqrt[60] ), .dout(n15001));
  jor  g14752(.dina(n15000), .dinb(asqrt[60] ), .dout(n15002));
  jxor g14753(.dina(n14392), .dinb(n352), .dout(n15003));
  jand g14754(.dina(n15003), .dinb(asqrt[16] ), .dout(n15004));
  jxor g14755(.dina(n15004), .dinb(n14397), .dout(n15005));
  jnot g14756(.din(n15005), .dout(n15006));
  jand g14757(.dina(n15006), .dinb(n15002), .dout(n15007));
  jor  g14758(.dina(n15007), .dinb(n15001), .dout(n15008));
  jand g14759(.dina(n15008), .dinb(asqrt[61] ), .dout(n15009));
  jor  g14760(.dina(n15008), .dinb(asqrt[61] ), .dout(n15010));
  jxor g14761(.dina(n14399), .dinb(n294), .dout(n15011));
  jand g14762(.dina(n15011), .dinb(asqrt[16] ), .dout(n15012));
  jxor g14763(.dina(n15012), .dinb(n14404), .dout(n15013));
  jand g14764(.dina(n15013), .dinb(n15010), .dout(n15014));
  jor  g14765(.dina(n15014), .dinb(n15009), .dout(n15015));
  jand g14766(.dina(n15015), .dinb(asqrt[62] ), .dout(n15016));
  jnot g14767(.din(n15016), .dout(n15017));
  jnot g14768(.din(n15009), .dout(n15018));
  jnot g14769(.din(n15001), .dout(n15019));
  jnot g14770(.din(n14994), .dout(n15020));
  jnot g14771(.din(n14986), .dout(n15021));
  jnot g14772(.din(n14979), .dout(n15022));
  jnot g14773(.din(n14971), .dout(n15023));
  jnot g14774(.din(n14964), .dout(n15024));
  jnot g14775(.din(n14956), .dout(n15025));
  jnot g14776(.din(n14948), .dout(n15026));
  jnot g14777(.din(n14940), .dout(n15027));
  jnot g14778(.din(n14933), .dout(n15028));
  jnot g14779(.din(n14925), .dout(n15029));
  jnot g14780(.din(n14918), .dout(n15030));
  jnot g14781(.din(n14910), .dout(n15031));
  jnot g14782(.din(n14903), .dout(n15032));
  jnot g14783(.din(n14906), .dout(n15033));
  jnot g14784(.din(n14896), .dout(n15034));
  jnot g14785(.din(n14888), .dout(n15035));
  jnot g14786(.din(n14880), .dout(n15036));
  jnot g14787(.din(n14873), .dout(n15037));
  jnot g14788(.din(n14865), .dout(n15038));
  jnot g14789(.din(n14858), .dout(n15039));
  jnot g14790(.din(n14850), .dout(n15040));
  jnot g14791(.din(n14842), .dout(n15041));
  jnot g14792(.din(n14834), .dout(n15042));
  jnot g14793(.din(n14827), .dout(n15043));
  jnot g14794(.din(n14819), .dout(n15044));
  jnot g14795(.din(n14812), .dout(n15045));
  jnot g14796(.din(n14804), .dout(n15046));
  jnot g14797(.din(n14796), .dout(n15047));
  jnot g14798(.din(n14788), .dout(n15048));
  jnot g14799(.din(n14781), .dout(n15049));
  jnot g14800(.din(n14773), .dout(n15050));
  jnot g14801(.din(n14766), .dout(n15051));
  jnot g14802(.din(n14758), .dout(n15052));
  jnot g14803(.din(n14751), .dout(n15053));
  jnot g14804(.din(n14743), .dout(n15054));
  jnot g14805(.din(n14736), .dout(n15055));
  jnot g14806(.din(n14728), .dout(n15056));
  jnot g14807(.din(n14720), .dout(n15057));
  jnot g14808(.din(n14712), .dout(n15058));
  jnot g14809(.din(n14705), .dout(n15059));
  jnot g14810(.din(n14697), .dout(n15060));
  jnot g14811(.din(n14690), .dout(n15061));
  jnot g14812(.din(n14679), .dout(n15062));
  jnot g14813(.din(n14449), .dout(n15063));
  jnot g14814(.din(n14446), .dout(n15064));
  jor  g14815(.dina(n14674), .dinb(n14080), .dout(n15065));
  jand g14816(.dina(n15065), .dinb(n15064), .dout(n15066));
  jand g14817(.dina(n15066), .dinb(n14078), .dout(n15067));
  jor  g14818(.dina(n14674), .dinb(a[32] ), .dout(n15068));
  jand g14819(.dina(n15068), .dinb(a[33] ), .dout(n15069));
  jor  g14820(.dina(n14681), .dinb(n15069), .dout(n15070));
  jor  g14821(.dina(n15070), .dinb(n15067), .dout(n15071));
  jand g14822(.dina(n15071), .dinb(n15063), .dout(n15072));
  jand g14823(.dina(n15072), .dinb(n13515), .dout(n15073));
  jor  g14824(.dina(n14686), .dinb(n15073), .dout(n15074));
  jand g14825(.dina(n15074), .dinb(n15062), .dout(n15075));
  jand g14826(.dina(n15075), .dinb(n12947), .dout(n15076));
  jnot g14827(.din(n14694), .dout(n15077));
  jor  g14828(.dina(n15077), .dinb(n15076), .dout(n15078));
  jand g14829(.dina(n15078), .dinb(n15061), .dout(n15079));
  jand g14830(.dina(n15079), .dinb(n12410), .dout(n15080));
  jor  g14831(.dina(n14701), .dinb(n15080), .dout(n15081));
  jand g14832(.dina(n15081), .dinb(n15060), .dout(n15082));
  jand g14833(.dina(n15082), .dinb(n11858), .dout(n15083));
  jnot g14834(.din(n14709), .dout(n15084));
  jor  g14835(.dina(n15084), .dinb(n15083), .dout(n15085));
  jand g14836(.dina(n15085), .dinb(n15059), .dout(n15086));
  jand g14837(.dina(n15086), .dinb(n11347), .dout(n15087));
  jor  g14838(.dina(n14716), .dinb(n15087), .dout(n15088));
  jand g14839(.dina(n15088), .dinb(n15058), .dout(n15089));
  jand g14840(.dina(n15089), .dinb(n10824), .dout(n15090));
  jor  g14841(.dina(n14724), .dinb(n15090), .dout(n15091));
  jand g14842(.dina(n15091), .dinb(n15057), .dout(n15092));
  jand g14843(.dina(n15092), .dinb(n10328), .dout(n15093));
  jor  g14844(.dina(n14732), .dinb(n15093), .dout(n15094));
  jand g14845(.dina(n15094), .dinb(n15056), .dout(n15095));
  jand g14846(.dina(n15095), .dinb(n9832), .dout(n15096));
  jnot g14847(.din(n14740), .dout(n15097));
  jor  g14848(.dina(n15097), .dinb(n15096), .dout(n15098));
  jand g14849(.dina(n15098), .dinb(n15055), .dout(n15099));
  jand g14850(.dina(n15099), .dinb(n9369), .dout(n15100));
  jor  g14851(.dina(n14747), .dinb(n15100), .dout(n15101));
  jand g14852(.dina(n15101), .dinb(n15054), .dout(n15102));
  jand g14853(.dina(n15102), .dinb(n8890), .dout(n15103));
  jnot g14854(.din(n14755), .dout(n15104));
  jor  g14855(.dina(n15104), .dinb(n15103), .dout(n15105));
  jand g14856(.dina(n15105), .dinb(n15053), .dout(n15106));
  jand g14857(.dina(n15106), .dinb(n8449), .dout(n15107));
  jor  g14858(.dina(n14762), .dinb(n15107), .dout(n15108));
  jand g14859(.dina(n15108), .dinb(n15052), .dout(n15109));
  jand g14860(.dina(n15109), .dinb(n8003), .dout(n15110));
  jnot g14861(.din(n14770), .dout(n15111));
  jor  g14862(.dina(n15111), .dinb(n15110), .dout(n15112));
  jand g14863(.dina(n15112), .dinb(n15051), .dout(n15113));
  jand g14864(.dina(n15113), .dinb(n7581), .dout(n15114));
  jor  g14865(.dina(n14777), .dinb(n15114), .dout(n15115));
  jand g14866(.dina(n15115), .dinb(n15050), .dout(n15116));
  jand g14867(.dina(n15116), .dinb(n7154), .dout(n15117));
  jnot g14868(.din(n14785), .dout(n15118));
  jor  g14869(.dina(n15118), .dinb(n15117), .dout(n15119));
  jand g14870(.dina(n15119), .dinb(n15049), .dout(n15120));
  jand g14871(.dina(n15120), .dinb(n6758), .dout(n15121));
  jor  g14872(.dina(n14792), .dinb(n15121), .dout(n15122));
  jand g14873(.dina(n15122), .dinb(n15048), .dout(n15123));
  jand g14874(.dina(n15123), .dinb(n6357), .dout(n15124));
  jor  g14875(.dina(n14800), .dinb(n15124), .dout(n15125));
  jand g14876(.dina(n15125), .dinb(n15047), .dout(n15126));
  jand g14877(.dina(n15126), .dinb(n5989), .dout(n15127));
  jor  g14878(.dina(n14808), .dinb(n15127), .dout(n15128));
  jand g14879(.dina(n15128), .dinb(n15046), .dout(n15129));
  jand g14880(.dina(n15129), .dinb(n5606), .dout(n15130));
  jnot g14881(.din(n14816), .dout(n15131));
  jor  g14882(.dina(n15131), .dinb(n15130), .dout(n15132));
  jand g14883(.dina(n15132), .dinb(n15045), .dout(n15133));
  jand g14884(.dina(n15133), .dinb(n5259), .dout(n15134));
  jor  g14885(.dina(n14823), .dinb(n15134), .dout(n15135));
  jand g14886(.dina(n15135), .dinb(n15044), .dout(n15136));
  jand g14887(.dina(n15136), .dinb(n4902), .dout(n15137));
  jnot g14888(.din(n14831), .dout(n15138));
  jor  g14889(.dina(n15138), .dinb(n15137), .dout(n15139));
  jand g14890(.dina(n15139), .dinb(n15043), .dout(n15140));
  jand g14891(.dina(n15140), .dinb(n4582), .dout(n15141));
  jor  g14892(.dina(n14838), .dinb(n15141), .dout(n15142));
  jand g14893(.dina(n15142), .dinb(n15042), .dout(n15143));
  jand g14894(.dina(n15143), .dinb(n4249), .dout(n15144));
  jor  g14895(.dina(n14846), .dinb(n15144), .dout(n15145));
  jand g14896(.dina(n15145), .dinb(n15041), .dout(n15146));
  jand g14897(.dina(n15146), .dinb(n3955), .dout(n15147));
  jor  g14898(.dina(n14854), .dinb(n15147), .dout(n15148));
  jand g14899(.dina(n15148), .dinb(n15040), .dout(n15149));
  jand g14900(.dina(n15149), .dinb(n3642), .dout(n15150));
  jnot g14901(.din(n14862), .dout(n15151));
  jor  g14902(.dina(n15151), .dinb(n15150), .dout(n15152));
  jand g14903(.dina(n15152), .dinb(n15039), .dout(n15153));
  jand g14904(.dina(n15153), .dinb(n3368), .dout(n15154));
  jor  g14905(.dina(n14869), .dinb(n15154), .dout(n15155));
  jand g14906(.dina(n15155), .dinb(n15038), .dout(n15156));
  jand g14907(.dina(n15156), .dinb(n3089), .dout(n15157));
  jnot g14908(.din(n14877), .dout(n15158));
  jor  g14909(.dina(n15158), .dinb(n15157), .dout(n15159));
  jand g14910(.dina(n15159), .dinb(n15037), .dout(n15160));
  jand g14911(.dina(n15160), .dinb(n2833), .dout(n15161));
  jor  g14912(.dina(n14884), .dinb(n15161), .dout(n15162));
  jand g14913(.dina(n15162), .dinb(n15036), .dout(n15163));
  jand g14914(.dina(n15163), .dinb(n2572), .dout(n15164));
  jor  g14915(.dina(n14892), .dinb(n15164), .dout(n15165));
  jand g14916(.dina(n15165), .dinb(n15035), .dout(n15166));
  jand g14917(.dina(n15166), .dinb(n2345), .dout(n15167));
  jnot g14918(.din(n14900), .dout(n15168));
  jor  g14919(.dina(n15168), .dinb(n15167), .dout(n15169));
  jand g14920(.dina(n15169), .dinb(n15034), .dout(n15170));
  jand g14921(.dina(n15170), .dinb(n2108), .dout(n15171));
  jor  g14922(.dina(n15171), .dinb(n15033), .dout(n15172));
  jand g14923(.dina(n15172), .dinb(n15032), .dout(n15173));
  jand g14924(.dina(n15173), .dinb(n1912), .dout(n15174));
  jor  g14925(.dina(n14914), .dinb(n15174), .dout(n15175));
  jand g14926(.dina(n15175), .dinb(n15031), .dout(n15176));
  jand g14927(.dina(n15176), .dinb(n1699), .dout(n15177));
  jnot g14928(.din(n14922), .dout(n15178));
  jor  g14929(.dina(n15178), .dinb(n15177), .dout(n15179));
  jand g14930(.dina(n15179), .dinb(n15030), .dout(n15180));
  jand g14931(.dina(n15180), .dinb(n1516), .dout(n15181));
  jor  g14932(.dina(n14929), .dinb(n15181), .dout(n15182));
  jand g14933(.dina(n15182), .dinb(n15029), .dout(n15183));
  jand g14934(.dina(n15183), .dinb(n1332), .dout(n15184));
  jnot g14935(.din(n14937), .dout(n15185));
  jor  g14936(.dina(n15185), .dinb(n15184), .dout(n15186));
  jand g14937(.dina(n15186), .dinb(n15028), .dout(n15187));
  jand g14938(.dina(n15187), .dinb(n1173), .dout(n15188));
  jor  g14939(.dina(n14944), .dinb(n15188), .dout(n15189));
  jand g14940(.dina(n15189), .dinb(n15027), .dout(n15190));
  jand g14941(.dina(n15190), .dinb(n1008), .dout(n15191));
  jor  g14942(.dina(n14952), .dinb(n15191), .dout(n15192));
  jand g14943(.dina(n15192), .dinb(n15026), .dout(n15193));
  jand g14944(.dina(n15193), .dinb(n884), .dout(n15194));
  jor  g14945(.dina(n14960), .dinb(n15194), .dout(n15195));
  jand g14946(.dina(n15195), .dinb(n15025), .dout(n15196));
  jand g14947(.dina(n15196), .dinb(n743), .dout(n15197));
  jnot g14948(.din(n14968), .dout(n15198));
  jor  g14949(.dina(n15198), .dinb(n15197), .dout(n15199));
  jand g14950(.dina(n15199), .dinb(n15024), .dout(n15200));
  jand g14951(.dina(n15200), .dinb(n635), .dout(n15201));
  jor  g14952(.dina(n14975), .dinb(n15201), .dout(n15202));
  jand g14953(.dina(n15202), .dinb(n15023), .dout(n15203));
  jand g14954(.dina(n15203), .dinb(n515), .dout(n15204));
  jnot g14955(.din(n14983), .dout(n15205));
  jor  g14956(.dina(n15205), .dinb(n15204), .dout(n15206));
  jand g14957(.dina(n15206), .dinb(n15022), .dout(n15207));
  jand g14958(.dina(n15207), .dinb(n443), .dout(n15208));
  jor  g14959(.dina(n14990), .dinb(n15208), .dout(n15209));
  jand g14960(.dina(n15209), .dinb(n15021), .dout(n15210));
  jand g14961(.dina(n15210), .dinb(n352), .dout(n15211));
  jnot g14962(.din(n14998), .dout(n15212));
  jor  g14963(.dina(n15212), .dinb(n15211), .dout(n15213));
  jand g14964(.dina(n15213), .dinb(n15020), .dout(n15214));
  jand g14965(.dina(n15214), .dinb(n294), .dout(n15215));
  jor  g14966(.dina(n15005), .dinb(n15215), .dout(n15216));
  jand g14967(.dina(n15216), .dinb(n15019), .dout(n15217));
  jand g14968(.dina(n15217), .dinb(n239), .dout(n15218));
  jnot g14969(.din(n15013), .dout(n15219));
  jor  g14970(.dina(n15219), .dinb(n15218), .dout(n15220));
  jand g14971(.dina(n15220), .dinb(n15018), .dout(n15221));
  jand g14972(.dina(n15221), .dinb(n221), .dout(n15222));
  jxor g14973(.dina(n14407), .dinb(n239), .dout(n15223));
  jand g14974(.dina(n15223), .dinb(asqrt[16] ), .dout(n15224));
  jxor g14975(.dina(n15224), .dinb(n14412), .dout(n15225));
  jnot g14976(.din(n15225), .dout(n15226));
  jor  g14977(.dina(n15226), .dinb(n15222), .dout(n15227));
  jand g14978(.dina(n15227), .dinb(n15017), .dout(n15228));
  jxor g14979(.dina(n14415), .dinb(n221), .dout(n15229));
  jand g14980(.dina(n15229), .dinb(asqrt[16] ), .dout(n15230));
  jxor g14981(.dina(n15230), .dinb(n14421), .dout(n15231));
  jor  g14982(.dina(n15231), .dinb(n15228), .dout(n15232));
  jxor g14983(.dina(n14426), .dinb(n14423), .dout(n15233));
  jnot g14984(.din(n15233), .dout(n15234));
  jand g14985(.dina(n15234), .dinb(asqrt[16] ), .dout(n15235));
  jor  g14986(.dina(n15235), .dinb(n15232), .dout(n15236));
  jand g14987(.dina(n15236), .dinb(n218), .dout(n15237));
  jand g14988(.dina(n14674), .dinb(n14426), .dout(n15238));
  jand g14989(.dina(n15231), .dinb(n15228), .dout(n15239));
  jor  g14990(.dina(n15239), .dinb(n15238), .dout(n15240));
  jand g14991(.dina(n14672), .dinb(n14423), .dout(n15241));
  jnot g14992(.din(n15241), .dout(n15242));
  jand g14993(.dina(n15233), .dinb(asqrt[63] ), .dout(n15243));
  jand g14994(.dina(n15243), .dinb(n15242), .dout(n15244));
  jor  g14995(.dina(n15244), .dinb(n15240), .dout(n15245));
  jor  g14996(.dina(n15245), .dinb(n15237), .dout(asqrt[15] ));
  jor  g14997(.dina(n15015), .dinb(asqrt[62] ), .dout(n15247));
  jand g14998(.dina(n15225), .dinb(n15247), .dout(n15248));
  jor  g14999(.dina(n15248), .dinb(n15016), .dout(n15249));
  jnot g15000(.din(n15231), .dout(n15250));
  jand g15001(.dina(n15250), .dinb(n15249), .dout(n15251));
  jnot g15002(.din(n15235), .dout(n15252));
  jand g15003(.dina(n15252), .dinb(n15251), .dout(n15253));
  jor  g15004(.dina(n15253), .dinb(asqrt[63] ), .dout(n15254));
  jnot g15005(.din(n15238), .dout(n15255));
  jor  g15006(.dina(n15250), .dinb(n15249), .dout(n15256));
  jand g15007(.dina(n15256), .dinb(n15255), .dout(n15257));
  jnot g15008(.din(n15244), .dout(n15258));
  jand g15009(.dina(n15258), .dinb(n15257), .dout(n15259));
  jand g15010(.dina(n15259), .dinb(n15254), .dout(n15260));
  jxor g15011(.dina(n15015), .dinb(n221), .dout(n15261));
  jor  g15012(.dina(n15261), .dinb(n15260), .dout(n15262));
  jxor g15013(.dina(n15262), .dinb(n15226), .dout(n15263));
  jnot g15014(.din(n15263), .dout(n15264));
  jnot g15015(.din(a[28] ), .dout(n15265));
  jnot g15016(.din(a[29] ), .dout(n15266));
  jand g15017(.dina(n15266), .dinb(n15265), .dout(n15267));
  jand g15018(.dina(n15267), .dinb(n14443), .dout(n15268));
  jnot g15019(.din(n15268), .dout(n15269));
  jor  g15020(.dina(n15260), .dinb(n14443), .dout(n15270));
  jand g15021(.dina(n15270), .dinb(n15269), .dout(n15271));
  jor  g15022(.dina(n15271), .dinb(n14674), .dout(n15272));
  jand g15023(.dina(n15271), .dinb(n14674), .dout(n15273));
  jor  g15024(.dina(n15260), .dinb(a[30] ), .dout(n15274));
  jand g15025(.dina(n15274), .dinb(a[31] ), .dout(n15275));
  jand g15026(.dina(asqrt[15] ), .dinb(n14445), .dout(n15276));
  jor  g15027(.dina(n15276), .dinb(n15275), .dout(n15277));
  jor  g15028(.dina(n15277), .dinb(n15273), .dout(n15278));
  jand g15029(.dina(n15278), .dinb(n15272), .dout(n15279));
  jor  g15030(.dina(n15279), .dinb(n14078), .dout(n15280));
  jand g15031(.dina(n15279), .dinb(n14078), .dout(n15281));
  jnot g15032(.din(n14445), .dout(n15282));
  jor  g15033(.dina(n15260), .dinb(n15282), .dout(n15283));
  jor  g15034(.dina(n15239), .dinb(n14674), .dout(n15284));
  jor  g15035(.dina(n15284), .dinb(n15237), .dout(n15285));
  jor  g15036(.dina(n15285), .dinb(n15243), .dout(n15286));
  jand g15037(.dina(n15286), .dinb(n15283), .dout(n15287));
  jxor g15038(.dina(n15287), .dinb(n14080), .dout(n15288));
  jor  g15039(.dina(n15288), .dinb(n15281), .dout(n15289));
  jand g15040(.dina(n15289), .dinb(n15280), .dout(n15290));
  jor  g15041(.dina(n15290), .dinb(n13515), .dout(n15291));
  jand g15042(.dina(n15290), .dinb(n13515), .dout(n15292));
  jxor g15043(.dina(n14448), .dinb(n14078), .dout(n15293));
  jor  g15044(.dina(n15293), .dinb(n15260), .dout(n15294));
  jxor g15045(.dina(n15294), .dinb(n15070), .dout(n15295));
  jnot g15046(.din(n15295), .dout(n15296));
  jor  g15047(.dina(n15296), .dinb(n15292), .dout(n15297));
  jand g15048(.dina(n15297), .dinb(n15291), .dout(n15298));
  jor  g15049(.dina(n15298), .dinb(n12947), .dout(n15299));
  jand g15050(.dina(n15298), .dinb(n12947), .dout(n15300));
  jxor g15051(.dina(n14678), .dinb(n13515), .dout(n15301));
  jor  g15052(.dina(n15301), .dinb(n15260), .dout(n15302));
  jxor g15053(.dina(n15302), .dinb(n14687), .dout(n15303));
  jor  g15054(.dina(n15303), .dinb(n15300), .dout(n15304));
  jand g15055(.dina(n15304), .dinb(n15299), .dout(n15305));
  jor  g15056(.dina(n15305), .dinb(n12410), .dout(n15306));
  jand g15057(.dina(n15305), .dinb(n12410), .dout(n15307));
  jxor g15058(.dina(n14689), .dinb(n12947), .dout(n15308));
  jor  g15059(.dina(n15308), .dinb(n15260), .dout(n15309));
  jxor g15060(.dina(n15309), .dinb(n15077), .dout(n15310));
  jnot g15061(.din(n15310), .dout(n15311));
  jor  g15062(.dina(n15311), .dinb(n15307), .dout(n15312));
  jand g15063(.dina(n15312), .dinb(n15306), .dout(n15313));
  jor  g15064(.dina(n15313), .dinb(n11858), .dout(n15314));
  jand g15065(.dina(n15313), .dinb(n11858), .dout(n15315));
  jxor g15066(.dina(n14696), .dinb(n12410), .dout(n15316));
  jor  g15067(.dina(n15316), .dinb(n15260), .dout(n15317));
  jxor g15068(.dina(n15317), .dinb(n14702), .dout(n15318));
  jor  g15069(.dina(n15318), .dinb(n15315), .dout(n15319));
  jand g15070(.dina(n15319), .dinb(n15314), .dout(n15320));
  jor  g15071(.dina(n15320), .dinb(n11347), .dout(n15321));
  jand g15072(.dina(n15320), .dinb(n11347), .dout(n15322));
  jxor g15073(.dina(n14704), .dinb(n11858), .dout(n15323));
  jor  g15074(.dina(n15323), .dinb(n15260), .dout(n15324));
  jxor g15075(.dina(n15324), .dinb(n15084), .dout(n15325));
  jnot g15076(.din(n15325), .dout(n15326));
  jor  g15077(.dina(n15326), .dinb(n15322), .dout(n15327));
  jand g15078(.dina(n15327), .dinb(n15321), .dout(n15328));
  jor  g15079(.dina(n15328), .dinb(n10824), .dout(n15329));
  jand g15080(.dina(n15328), .dinb(n10824), .dout(n15330));
  jxor g15081(.dina(n14711), .dinb(n11347), .dout(n15331));
  jor  g15082(.dina(n15331), .dinb(n15260), .dout(n15332));
  jxor g15083(.dina(n15332), .dinb(n14717), .dout(n15333));
  jor  g15084(.dina(n15333), .dinb(n15330), .dout(n15334));
  jand g15085(.dina(n15334), .dinb(n15329), .dout(n15335));
  jor  g15086(.dina(n15335), .dinb(n10328), .dout(n15336));
  jand g15087(.dina(n15335), .dinb(n10328), .dout(n15337));
  jxor g15088(.dina(n14719), .dinb(n10824), .dout(n15338));
  jor  g15089(.dina(n15338), .dinb(n15260), .dout(n15339));
  jxor g15090(.dina(n15339), .dinb(n14725), .dout(n15340));
  jor  g15091(.dina(n15340), .dinb(n15337), .dout(n15341));
  jand g15092(.dina(n15341), .dinb(n15336), .dout(n15342));
  jor  g15093(.dina(n15342), .dinb(n9832), .dout(n15343));
  jand g15094(.dina(n15342), .dinb(n9832), .dout(n15344));
  jxor g15095(.dina(n14727), .dinb(n10328), .dout(n15345));
  jor  g15096(.dina(n15345), .dinb(n15260), .dout(n15346));
  jxor g15097(.dina(n15346), .dinb(n14733), .dout(n15347));
  jor  g15098(.dina(n15347), .dinb(n15344), .dout(n15348));
  jand g15099(.dina(n15348), .dinb(n15343), .dout(n15349));
  jor  g15100(.dina(n15349), .dinb(n9369), .dout(n15350));
  jand g15101(.dina(n15349), .dinb(n9369), .dout(n15351));
  jxor g15102(.dina(n14735), .dinb(n9832), .dout(n15352));
  jor  g15103(.dina(n15352), .dinb(n15260), .dout(n15353));
  jxor g15104(.dina(n15353), .dinb(n15097), .dout(n15354));
  jnot g15105(.din(n15354), .dout(n15355));
  jor  g15106(.dina(n15355), .dinb(n15351), .dout(n15356));
  jand g15107(.dina(n15356), .dinb(n15350), .dout(n15357));
  jor  g15108(.dina(n15357), .dinb(n8890), .dout(n15358));
  jand g15109(.dina(n15357), .dinb(n8890), .dout(n15359));
  jxor g15110(.dina(n14742), .dinb(n9369), .dout(n15360));
  jor  g15111(.dina(n15360), .dinb(n15260), .dout(n15361));
  jxor g15112(.dina(n15361), .dinb(n14748), .dout(n15362));
  jor  g15113(.dina(n15362), .dinb(n15359), .dout(n15363));
  jand g15114(.dina(n15363), .dinb(n15358), .dout(n15364));
  jor  g15115(.dina(n15364), .dinb(n8449), .dout(n15365));
  jand g15116(.dina(n15364), .dinb(n8449), .dout(n15366));
  jxor g15117(.dina(n14750), .dinb(n8890), .dout(n15367));
  jor  g15118(.dina(n15367), .dinb(n15260), .dout(n15368));
  jxor g15119(.dina(n15368), .dinb(n15104), .dout(n15369));
  jnot g15120(.din(n15369), .dout(n15370));
  jor  g15121(.dina(n15370), .dinb(n15366), .dout(n15371));
  jand g15122(.dina(n15371), .dinb(n15365), .dout(n15372));
  jor  g15123(.dina(n15372), .dinb(n8003), .dout(n15373));
  jand g15124(.dina(n15372), .dinb(n8003), .dout(n15374));
  jxor g15125(.dina(n14757), .dinb(n8449), .dout(n15375));
  jor  g15126(.dina(n15375), .dinb(n15260), .dout(n15376));
  jxor g15127(.dina(n15376), .dinb(n14763), .dout(n15377));
  jor  g15128(.dina(n15377), .dinb(n15374), .dout(n15378));
  jand g15129(.dina(n15378), .dinb(n15373), .dout(n15379));
  jor  g15130(.dina(n15379), .dinb(n7581), .dout(n15380));
  jand g15131(.dina(n15379), .dinb(n7581), .dout(n15381));
  jxor g15132(.dina(n14765), .dinb(n8003), .dout(n15382));
  jor  g15133(.dina(n15382), .dinb(n15260), .dout(n15383));
  jxor g15134(.dina(n15383), .dinb(n15111), .dout(n15384));
  jnot g15135(.din(n15384), .dout(n15385));
  jor  g15136(.dina(n15385), .dinb(n15381), .dout(n15386));
  jand g15137(.dina(n15386), .dinb(n15380), .dout(n15387));
  jor  g15138(.dina(n15387), .dinb(n7154), .dout(n15388));
  jand g15139(.dina(n15387), .dinb(n7154), .dout(n15389));
  jxor g15140(.dina(n14772), .dinb(n7581), .dout(n15390));
  jor  g15141(.dina(n15390), .dinb(n15260), .dout(n15391));
  jxor g15142(.dina(n15391), .dinb(n14778), .dout(n15392));
  jor  g15143(.dina(n15392), .dinb(n15389), .dout(n15393));
  jand g15144(.dina(n15393), .dinb(n15388), .dout(n15394));
  jor  g15145(.dina(n15394), .dinb(n6758), .dout(n15395));
  jand g15146(.dina(n15394), .dinb(n6758), .dout(n15396));
  jxor g15147(.dina(n14780), .dinb(n7154), .dout(n15397));
  jor  g15148(.dina(n15397), .dinb(n15260), .dout(n15398));
  jxor g15149(.dina(n15398), .dinb(n15118), .dout(n15399));
  jnot g15150(.din(n15399), .dout(n15400));
  jor  g15151(.dina(n15400), .dinb(n15396), .dout(n15401));
  jand g15152(.dina(n15401), .dinb(n15395), .dout(n15402));
  jor  g15153(.dina(n15402), .dinb(n6357), .dout(n15403));
  jand g15154(.dina(n15402), .dinb(n6357), .dout(n15404));
  jxor g15155(.dina(n14787), .dinb(n6758), .dout(n15405));
  jor  g15156(.dina(n15405), .dinb(n15260), .dout(n15406));
  jxor g15157(.dina(n15406), .dinb(n14793), .dout(n15407));
  jor  g15158(.dina(n15407), .dinb(n15404), .dout(n15408));
  jand g15159(.dina(n15408), .dinb(n15403), .dout(n15409));
  jor  g15160(.dina(n15409), .dinb(n5989), .dout(n15410));
  jand g15161(.dina(n15409), .dinb(n5989), .dout(n15411));
  jxor g15162(.dina(n14795), .dinb(n6357), .dout(n15412));
  jor  g15163(.dina(n15412), .dinb(n15260), .dout(n15413));
  jxor g15164(.dina(n15413), .dinb(n14801), .dout(n15414));
  jor  g15165(.dina(n15414), .dinb(n15411), .dout(n15415));
  jand g15166(.dina(n15415), .dinb(n15410), .dout(n15416));
  jor  g15167(.dina(n15416), .dinb(n5606), .dout(n15417));
  jand g15168(.dina(n15416), .dinb(n5606), .dout(n15418));
  jxor g15169(.dina(n14803), .dinb(n5989), .dout(n15419));
  jor  g15170(.dina(n15419), .dinb(n15260), .dout(n15420));
  jxor g15171(.dina(n15420), .dinb(n14809), .dout(n15421));
  jor  g15172(.dina(n15421), .dinb(n15418), .dout(n15422));
  jand g15173(.dina(n15422), .dinb(n15417), .dout(n15423));
  jor  g15174(.dina(n15423), .dinb(n5259), .dout(n15424));
  jand g15175(.dina(n15423), .dinb(n5259), .dout(n15425));
  jxor g15176(.dina(n14811), .dinb(n5606), .dout(n15426));
  jor  g15177(.dina(n15426), .dinb(n15260), .dout(n15427));
  jxor g15178(.dina(n15427), .dinb(n15131), .dout(n15428));
  jnot g15179(.din(n15428), .dout(n15429));
  jor  g15180(.dina(n15429), .dinb(n15425), .dout(n15430));
  jand g15181(.dina(n15430), .dinb(n15424), .dout(n15431));
  jor  g15182(.dina(n15431), .dinb(n4902), .dout(n15432));
  jand g15183(.dina(n15431), .dinb(n4902), .dout(n15433));
  jxor g15184(.dina(n14818), .dinb(n5259), .dout(n15434));
  jor  g15185(.dina(n15434), .dinb(n15260), .dout(n15435));
  jxor g15186(.dina(n15435), .dinb(n14824), .dout(n15436));
  jor  g15187(.dina(n15436), .dinb(n15433), .dout(n15437));
  jand g15188(.dina(n15437), .dinb(n15432), .dout(n15438));
  jor  g15189(.dina(n15438), .dinb(n4582), .dout(n15439));
  jand g15190(.dina(n15438), .dinb(n4582), .dout(n15440));
  jxor g15191(.dina(n14826), .dinb(n4902), .dout(n15441));
  jor  g15192(.dina(n15441), .dinb(n15260), .dout(n15442));
  jxor g15193(.dina(n15442), .dinb(n15138), .dout(n15443));
  jnot g15194(.din(n15443), .dout(n15444));
  jor  g15195(.dina(n15444), .dinb(n15440), .dout(n15445));
  jand g15196(.dina(n15445), .dinb(n15439), .dout(n15446));
  jor  g15197(.dina(n15446), .dinb(n4249), .dout(n15447));
  jand g15198(.dina(n15446), .dinb(n4249), .dout(n15448));
  jxor g15199(.dina(n14833), .dinb(n4582), .dout(n15449));
  jor  g15200(.dina(n15449), .dinb(n15260), .dout(n15450));
  jxor g15201(.dina(n15450), .dinb(n14839), .dout(n15451));
  jor  g15202(.dina(n15451), .dinb(n15448), .dout(n15452));
  jand g15203(.dina(n15452), .dinb(n15447), .dout(n15453));
  jor  g15204(.dina(n15453), .dinb(n3955), .dout(n15454));
  jand g15205(.dina(n15453), .dinb(n3955), .dout(n15455));
  jxor g15206(.dina(n14841), .dinb(n4249), .dout(n15456));
  jor  g15207(.dina(n15456), .dinb(n15260), .dout(n15457));
  jxor g15208(.dina(n15457), .dinb(n14847), .dout(n15458));
  jor  g15209(.dina(n15458), .dinb(n15455), .dout(n15459));
  jand g15210(.dina(n15459), .dinb(n15454), .dout(n15460));
  jor  g15211(.dina(n15460), .dinb(n3642), .dout(n15461));
  jand g15212(.dina(n15460), .dinb(n3642), .dout(n15462));
  jxor g15213(.dina(n14849), .dinb(n3955), .dout(n15463));
  jor  g15214(.dina(n15463), .dinb(n15260), .dout(n15464));
  jxor g15215(.dina(n15464), .dinb(n14855), .dout(n15465));
  jor  g15216(.dina(n15465), .dinb(n15462), .dout(n15466));
  jand g15217(.dina(n15466), .dinb(n15461), .dout(n15467));
  jor  g15218(.dina(n15467), .dinb(n3368), .dout(n15468));
  jand g15219(.dina(n15467), .dinb(n3368), .dout(n15469));
  jxor g15220(.dina(n14857), .dinb(n3642), .dout(n15470));
  jor  g15221(.dina(n15470), .dinb(n15260), .dout(n15471));
  jxor g15222(.dina(n15471), .dinb(n15151), .dout(n15472));
  jnot g15223(.din(n15472), .dout(n15473));
  jor  g15224(.dina(n15473), .dinb(n15469), .dout(n15474));
  jand g15225(.dina(n15474), .dinb(n15468), .dout(n15475));
  jor  g15226(.dina(n15475), .dinb(n3089), .dout(n15476));
  jand g15227(.dina(n15475), .dinb(n3089), .dout(n15477));
  jxor g15228(.dina(n14864), .dinb(n3368), .dout(n15478));
  jor  g15229(.dina(n15478), .dinb(n15260), .dout(n15479));
  jxor g15230(.dina(n15479), .dinb(n14870), .dout(n15480));
  jor  g15231(.dina(n15480), .dinb(n15477), .dout(n15481));
  jand g15232(.dina(n15481), .dinb(n15476), .dout(n15482));
  jor  g15233(.dina(n15482), .dinb(n2833), .dout(n15483));
  jand g15234(.dina(n15482), .dinb(n2833), .dout(n15484));
  jxor g15235(.dina(n14872), .dinb(n3089), .dout(n15485));
  jor  g15236(.dina(n15485), .dinb(n15260), .dout(n15486));
  jxor g15237(.dina(n15486), .dinb(n15158), .dout(n15487));
  jnot g15238(.din(n15487), .dout(n15488));
  jor  g15239(.dina(n15488), .dinb(n15484), .dout(n15489));
  jand g15240(.dina(n15489), .dinb(n15483), .dout(n15490));
  jor  g15241(.dina(n15490), .dinb(n2572), .dout(n15491));
  jand g15242(.dina(n15490), .dinb(n2572), .dout(n15492));
  jxor g15243(.dina(n14879), .dinb(n2833), .dout(n15493));
  jor  g15244(.dina(n15493), .dinb(n15260), .dout(n15494));
  jxor g15245(.dina(n15494), .dinb(n14885), .dout(n15495));
  jor  g15246(.dina(n15495), .dinb(n15492), .dout(n15496));
  jand g15247(.dina(n15496), .dinb(n15491), .dout(n15497));
  jor  g15248(.dina(n15497), .dinb(n2345), .dout(n15498));
  jand g15249(.dina(n15497), .dinb(n2345), .dout(n15499));
  jxor g15250(.dina(n14887), .dinb(n2572), .dout(n15500));
  jor  g15251(.dina(n15500), .dinb(n15260), .dout(n15501));
  jxor g15252(.dina(n15501), .dinb(n14893), .dout(n15502));
  jor  g15253(.dina(n15502), .dinb(n15499), .dout(n15503));
  jand g15254(.dina(n15503), .dinb(n15498), .dout(n15504));
  jor  g15255(.dina(n15504), .dinb(n2108), .dout(n15505));
  jand g15256(.dina(n15504), .dinb(n2108), .dout(n15506));
  jxor g15257(.dina(n14895), .dinb(n2345), .dout(n15507));
  jor  g15258(.dina(n15507), .dinb(n15260), .dout(n15508));
  jxor g15259(.dina(n15508), .dinb(n15168), .dout(n15509));
  jnot g15260(.din(n15509), .dout(n15510));
  jor  g15261(.dina(n15510), .dinb(n15506), .dout(n15511));
  jand g15262(.dina(n15511), .dinb(n15505), .dout(n15512));
  jor  g15263(.dina(n15512), .dinb(n1912), .dout(n15513));
  jxor g15264(.dina(n14902), .dinb(n2108), .dout(n15514));
  jor  g15265(.dina(n15514), .dinb(n15260), .dout(n15515));
  jxor g15266(.dina(n15515), .dinb(n15033), .dout(n15516));
  jnot g15267(.din(n15516), .dout(n15517));
  jand g15268(.dina(n15512), .dinb(n1912), .dout(n15518));
  jor  g15269(.dina(n15518), .dinb(n15517), .dout(n15519));
  jand g15270(.dina(n15519), .dinb(n15513), .dout(n15520));
  jor  g15271(.dina(n15520), .dinb(n1699), .dout(n15521));
  jand g15272(.dina(n15520), .dinb(n1699), .dout(n15522));
  jxor g15273(.dina(n14909), .dinb(n1912), .dout(n15523));
  jor  g15274(.dina(n15523), .dinb(n15260), .dout(n15524));
  jxor g15275(.dina(n15524), .dinb(n14915), .dout(n15525));
  jor  g15276(.dina(n15525), .dinb(n15522), .dout(n15526));
  jand g15277(.dina(n15526), .dinb(n15521), .dout(n15527));
  jor  g15278(.dina(n15527), .dinb(n1516), .dout(n15528));
  jand g15279(.dina(n15527), .dinb(n1516), .dout(n15529));
  jxor g15280(.dina(n14917), .dinb(n1699), .dout(n15530));
  jor  g15281(.dina(n15530), .dinb(n15260), .dout(n15531));
  jxor g15282(.dina(n15531), .dinb(n15178), .dout(n15532));
  jnot g15283(.din(n15532), .dout(n15533));
  jor  g15284(.dina(n15533), .dinb(n15529), .dout(n15534));
  jand g15285(.dina(n15534), .dinb(n15528), .dout(n15535));
  jor  g15286(.dina(n15535), .dinb(n1332), .dout(n15536));
  jand g15287(.dina(n15535), .dinb(n1332), .dout(n15537));
  jxor g15288(.dina(n14924), .dinb(n1516), .dout(n15538));
  jor  g15289(.dina(n15538), .dinb(n15260), .dout(n15539));
  jxor g15290(.dina(n15539), .dinb(n14930), .dout(n15540));
  jor  g15291(.dina(n15540), .dinb(n15537), .dout(n15541));
  jand g15292(.dina(n15541), .dinb(n15536), .dout(n15542));
  jor  g15293(.dina(n15542), .dinb(n1173), .dout(n15543));
  jand g15294(.dina(n15542), .dinb(n1173), .dout(n15544));
  jxor g15295(.dina(n14932), .dinb(n1332), .dout(n15545));
  jor  g15296(.dina(n15545), .dinb(n15260), .dout(n15546));
  jxor g15297(.dina(n15546), .dinb(n15185), .dout(n15547));
  jnot g15298(.din(n15547), .dout(n15548));
  jor  g15299(.dina(n15548), .dinb(n15544), .dout(n15549));
  jand g15300(.dina(n15549), .dinb(n15543), .dout(n15550));
  jor  g15301(.dina(n15550), .dinb(n1008), .dout(n15551));
  jand g15302(.dina(n15550), .dinb(n1008), .dout(n15552));
  jxor g15303(.dina(n14939), .dinb(n1173), .dout(n15553));
  jor  g15304(.dina(n15553), .dinb(n15260), .dout(n15554));
  jxor g15305(.dina(n15554), .dinb(n14945), .dout(n15555));
  jor  g15306(.dina(n15555), .dinb(n15552), .dout(n15556));
  jand g15307(.dina(n15556), .dinb(n15551), .dout(n15557));
  jor  g15308(.dina(n15557), .dinb(n884), .dout(n15558));
  jand g15309(.dina(n15557), .dinb(n884), .dout(n15559));
  jxor g15310(.dina(n14947), .dinb(n1008), .dout(n15560));
  jor  g15311(.dina(n15560), .dinb(n15260), .dout(n15561));
  jxor g15312(.dina(n15561), .dinb(n14953), .dout(n15562));
  jor  g15313(.dina(n15562), .dinb(n15559), .dout(n15563));
  jand g15314(.dina(n15563), .dinb(n15558), .dout(n15564));
  jor  g15315(.dina(n15564), .dinb(n743), .dout(n15565));
  jand g15316(.dina(n15564), .dinb(n743), .dout(n15566));
  jxor g15317(.dina(n14955), .dinb(n884), .dout(n15567));
  jor  g15318(.dina(n15567), .dinb(n15260), .dout(n15568));
  jxor g15319(.dina(n15568), .dinb(n14961), .dout(n15569));
  jor  g15320(.dina(n15569), .dinb(n15566), .dout(n15570));
  jand g15321(.dina(n15570), .dinb(n15565), .dout(n15571));
  jor  g15322(.dina(n15571), .dinb(n635), .dout(n15572));
  jand g15323(.dina(n15571), .dinb(n635), .dout(n15573));
  jxor g15324(.dina(n14963), .dinb(n743), .dout(n15574));
  jor  g15325(.dina(n15574), .dinb(n15260), .dout(n15575));
  jxor g15326(.dina(n15575), .dinb(n15198), .dout(n15576));
  jnot g15327(.din(n15576), .dout(n15577));
  jor  g15328(.dina(n15577), .dinb(n15573), .dout(n15578));
  jand g15329(.dina(n15578), .dinb(n15572), .dout(n15579));
  jor  g15330(.dina(n15579), .dinb(n515), .dout(n15580));
  jand g15331(.dina(n15579), .dinb(n515), .dout(n15581));
  jxor g15332(.dina(n14970), .dinb(n635), .dout(n15582));
  jor  g15333(.dina(n15582), .dinb(n15260), .dout(n15583));
  jxor g15334(.dina(n15583), .dinb(n14976), .dout(n15584));
  jor  g15335(.dina(n15584), .dinb(n15581), .dout(n15585));
  jand g15336(.dina(n15585), .dinb(n15580), .dout(n15586));
  jor  g15337(.dina(n15586), .dinb(n443), .dout(n15587));
  jand g15338(.dina(n15586), .dinb(n443), .dout(n15588));
  jxor g15339(.dina(n14978), .dinb(n515), .dout(n15589));
  jor  g15340(.dina(n15589), .dinb(n15260), .dout(n15590));
  jxor g15341(.dina(n15590), .dinb(n15205), .dout(n15591));
  jnot g15342(.din(n15591), .dout(n15592));
  jor  g15343(.dina(n15592), .dinb(n15588), .dout(n15593));
  jand g15344(.dina(n15593), .dinb(n15587), .dout(n15594));
  jor  g15345(.dina(n15594), .dinb(n352), .dout(n15595));
  jand g15346(.dina(n15594), .dinb(n352), .dout(n15596));
  jxor g15347(.dina(n14985), .dinb(n443), .dout(n15597));
  jor  g15348(.dina(n15597), .dinb(n15260), .dout(n15598));
  jxor g15349(.dina(n15598), .dinb(n14991), .dout(n15599));
  jor  g15350(.dina(n15599), .dinb(n15596), .dout(n15600));
  jand g15351(.dina(n15600), .dinb(n15595), .dout(n15601));
  jor  g15352(.dina(n15601), .dinb(n294), .dout(n15602));
  jand g15353(.dina(n15601), .dinb(n294), .dout(n15603));
  jxor g15354(.dina(n14993), .dinb(n352), .dout(n15604));
  jor  g15355(.dina(n15604), .dinb(n15260), .dout(n15605));
  jxor g15356(.dina(n15605), .dinb(n15212), .dout(n15606));
  jnot g15357(.din(n15606), .dout(n15607));
  jor  g15358(.dina(n15607), .dinb(n15603), .dout(n15608));
  jand g15359(.dina(n15608), .dinb(n15602), .dout(n15609));
  jor  g15360(.dina(n15609), .dinb(n239), .dout(n15610));
  jand g15361(.dina(n15609), .dinb(n239), .dout(n15611));
  jxor g15362(.dina(n15000), .dinb(n294), .dout(n15612));
  jor  g15363(.dina(n15612), .dinb(n15260), .dout(n15613));
  jxor g15364(.dina(n15613), .dinb(n15006), .dout(n15614));
  jor  g15365(.dina(n15614), .dinb(n15611), .dout(n15615));
  jand g15366(.dina(n15615), .dinb(n15610), .dout(n15616));
  jor  g15367(.dina(n15616), .dinb(n221), .dout(n15617));
  jand g15368(.dina(n15616), .dinb(n221), .dout(n15618));
  jxor g15369(.dina(n15008), .dinb(n239), .dout(n15619));
  jor  g15370(.dina(n15619), .dinb(n15260), .dout(n15620));
  jxor g15371(.dina(n15620), .dinb(n15219), .dout(n15621));
  jnot g15372(.din(n15621), .dout(n15622));
  jor  g15373(.dina(n15622), .dinb(n15618), .dout(n15623));
  jand g15374(.dina(n15623), .dinb(n15617), .dout(n15624));
  jor  g15375(.dina(n15624), .dinb(n15264), .dout(n15625));
  jand g15376(.dina(asqrt[15] ), .dinb(n15251), .dout(n15626));
  jor  g15377(.dina(n15626), .dinb(n15625), .dout(n15627));
  jor  g15378(.dina(n15627), .dinb(n15239), .dout(n15628));
  jand g15379(.dina(n15628), .dinb(n218), .dout(n15629));
  jand g15380(.dina(n15260), .dinb(n15231), .dout(n15630));
  jand g15381(.dina(n15624), .dinb(n15264), .dout(n15631));
  jor  g15382(.dina(n15631), .dinb(n15630), .dout(n15632));
  jand g15383(.dina(n15260), .dinb(n15228), .dout(n15633));
  jand g15384(.dina(n15232), .dinb(asqrt[63] ), .dout(n15634));
  jand g15385(.dina(n15634), .dinb(n15256), .dout(n15635));
  jnot g15386(.din(n15635), .dout(n15636));
  jor  g15387(.dina(n15636), .dinb(n15633), .dout(n15637));
  jnot g15388(.din(n15637), .dout(n15638));
  jor  g15389(.dina(n15638), .dinb(n15632), .dout(n15639));
  jor  g15390(.dina(n15639), .dinb(n15629), .dout(asqrt[14] ));
  jand g15391(.dina(asqrt[14] ), .dinb(a[28] ), .dout(n15641));
  jnot g15392(.din(a[26] ), .dout(n15642));
  jnot g15393(.din(a[27] ), .dout(n15643));
  jand g15394(.dina(n15643), .dinb(n15642), .dout(n15644));
  jand g15395(.dina(n15644), .dinb(n15265), .dout(n15645));
  jor  g15396(.dina(n15645), .dinb(n15641), .dout(n15646));
  jand g15397(.dina(n15646), .dinb(asqrt[15] ), .dout(n15647));
  jor  g15398(.dina(n15646), .dinb(asqrt[15] ), .dout(n15648));
  jand g15399(.dina(asqrt[14] ), .dinb(n15265), .dout(n15649));
  jor  g15400(.dina(n15649), .dinb(n15266), .dout(n15650));
  jnot g15401(.din(n15267), .dout(n15651));
  jnot g15402(.din(n15617), .dout(n15652));
  jnot g15403(.din(n15610), .dout(n15653));
  jnot g15404(.din(n15602), .dout(n15654));
  jnot g15405(.din(n15595), .dout(n15655));
  jnot g15406(.din(n15587), .dout(n15656));
  jnot g15407(.din(n15580), .dout(n15657));
  jnot g15408(.din(n15572), .dout(n15658));
  jnot g15409(.din(n15565), .dout(n15659));
  jnot g15410(.din(n15558), .dout(n15660));
  jnot g15411(.din(n15551), .dout(n15661));
  jnot g15412(.din(n15543), .dout(n15662));
  jnot g15413(.din(n15536), .dout(n15663));
  jnot g15414(.din(n15528), .dout(n15664));
  jnot g15415(.din(n15521), .dout(n15665));
  jnot g15416(.din(n15513), .dout(n15666));
  jnot g15417(.din(n15505), .dout(n15667));
  jnot g15418(.din(n15498), .dout(n15668));
  jnot g15419(.din(n15491), .dout(n15669));
  jnot g15420(.din(n15483), .dout(n15670));
  jnot g15421(.din(n15476), .dout(n15671));
  jnot g15422(.din(n15468), .dout(n15672));
  jnot g15423(.din(n15461), .dout(n15673));
  jnot g15424(.din(n15454), .dout(n15674));
  jnot g15425(.din(n15447), .dout(n15675));
  jnot g15426(.din(n15439), .dout(n15676));
  jnot g15427(.din(n15432), .dout(n15677));
  jnot g15428(.din(n15424), .dout(n15678));
  jnot g15429(.din(n15417), .dout(n15679));
  jnot g15430(.din(n15410), .dout(n15680));
  jnot g15431(.din(n15403), .dout(n15681));
  jnot g15432(.din(n15395), .dout(n15682));
  jnot g15433(.din(n15388), .dout(n15683));
  jnot g15434(.din(n15380), .dout(n15684));
  jnot g15435(.din(n15373), .dout(n15685));
  jnot g15436(.din(n15365), .dout(n15686));
  jnot g15437(.din(n15358), .dout(n15687));
  jnot g15438(.din(n15350), .dout(n15688));
  jnot g15439(.din(n15343), .dout(n15689));
  jnot g15440(.din(n15336), .dout(n15690));
  jnot g15441(.din(n15329), .dout(n15691));
  jnot g15442(.din(n15321), .dout(n15692));
  jnot g15443(.din(n15314), .dout(n15693));
  jnot g15444(.din(n15306), .dout(n15694));
  jnot g15445(.din(n15299), .dout(n15695));
  jnot g15446(.din(n15291), .dout(n15696));
  jnot g15447(.din(n15280), .dout(n15697));
  jnot g15448(.din(n15272), .dout(n15698));
  jand g15449(.dina(asqrt[15] ), .dinb(a[30] ), .dout(n15699));
  jor  g15450(.dina(n15699), .dinb(n15268), .dout(n15700));
  jor  g15451(.dina(n15700), .dinb(asqrt[16] ), .dout(n15701));
  jand g15452(.dina(asqrt[15] ), .dinb(n14443), .dout(n15702));
  jor  g15453(.dina(n15702), .dinb(n14444), .dout(n15703));
  jand g15454(.dina(n15283), .dinb(n15703), .dout(n15704));
  jand g15455(.dina(n15704), .dinb(n15701), .dout(n15705));
  jor  g15456(.dina(n15705), .dinb(n15698), .dout(n15706));
  jor  g15457(.dina(n15706), .dinb(asqrt[17] ), .dout(n15707));
  jnot g15458(.din(n15288), .dout(n15708));
  jand g15459(.dina(n15708), .dinb(n15707), .dout(n15709));
  jor  g15460(.dina(n15709), .dinb(n15697), .dout(n15710));
  jor  g15461(.dina(n15710), .dinb(asqrt[18] ), .dout(n15711));
  jand g15462(.dina(n15295), .dinb(n15711), .dout(n15712));
  jor  g15463(.dina(n15712), .dinb(n15696), .dout(n15713));
  jor  g15464(.dina(n15713), .dinb(asqrt[19] ), .dout(n15714));
  jnot g15465(.din(n15303), .dout(n15715));
  jand g15466(.dina(n15715), .dinb(n15714), .dout(n15716));
  jor  g15467(.dina(n15716), .dinb(n15695), .dout(n15717));
  jor  g15468(.dina(n15717), .dinb(asqrt[20] ), .dout(n15718));
  jand g15469(.dina(n15310), .dinb(n15718), .dout(n15719));
  jor  g15470(.dina(n15719), .dinb(n15694), .dout(n15720));
  jor  g15471(.dina(n15720), .dinb(asqrt[21] ), .dout(n15721));
  jnot g15472(.din(n15318), .dout(n15722));
  jand g15473(.dina(n15722), .dinb(n15721), .dout(n15723));
  jor  g15474(.dina(n15723), .dinb(n15693), .dout(n15724));
  jor  g15475(.dina(n15724), .dinb(asqrt[22] ), .dout(n15725));
  jand g15476(.dina(n15325), .dinb(n15725), .dout(n15726));
  jor  g15477(.dina(n15726), .dinb(n15692), .dout(n15727));
  jor  g15478(.dina(n15727), .dinb(asqrt[23] ), .dout(n15728));
  jnot g15479(.din(n15333), .dout(n15729));
  jand g15480(.dina(n15729), .dinb(n15728), .dout(n15730));
  jor  g15481(.dina(n15730), .dinb(n15691), .dout(n15731));
  jor  g15482(.dina(n15731), .dinb(asqrt[24] ), .dout(n15732));
  jnot g15483(.din(n15340), .dout(n15733));
  jand g15484(.dina(n15733), .dinb(n15732), .dout(n15734));
  jor  g15485(.dina(n15734), .dinb(n15690), .dout(n15735));
  jor  g15486(.dina(n15735), .dinb(asqrt[25] ), .dout(n15736));
  jnot g15487(.din(n15347), .dout(n15737));
  jand g15488(.dina(n15737), .dinb(n15736), .dout(n15738));
  jor  g15489(.dina(n15738), .dinb(n15689), .dout(n15739));
  jor  g15490(.dina(n15739), .dinb(asqrt[26] ), .dout(n15740));
  jand g15491(.dina(n15354), .dinb(n15740), .dout(n15741));
  jor  g15492(.dina(n15741), .dinb(n15688), .dout(n15742));
  jor  g15493(.dina(n15742), .dinb(asqrt[27] ), .dout(n15743));
  jnot g15494(.din(n15362), .dout(n15744));
  jand g15495(.dina(n15744), .dinb(n15743), .dout(n15745));
  jor  g15496(.dina(n15745), .dinb(n15687), .dout(n15746));
  jor  g15497(.dina(n15746), .dinb(asqrt[28] ), .dout(n15747));
  jand g15498(.dina(n15369), .dinb(n15747), .dout(n15748));
  jor  g15499(.dina(n15748), .dinb(n15686), .dout(n15749));
  jor  g15500(.dina(n15749), .dinb(asqrt[29] ), .dout(n15750));
  jnot g15501(.din(n15377), .dout(n15751));
  jand g15502(.dina(n15751), .dinb(n15750), .dout(n15752));
  jor  g15503(.dina(n15752), .dinb(n15685), .dout(n15753));
  jor  g15504(.dina(n15753), .dinb(asqrt[30] ), .dout(n15754));
  jand g15505(.dina(n15384), .dinb(n15754), .dout(n15755));
  jor  g15506(.dina(n15755), .dinb(n15684), .dout(n15756));
  jor  g15507(.dina(n15756), .dinb(asqrt[31] ), .dout(n15757));
  jnot g15508(.din(n15392), .dout(n15758));
  jand g15509(.dina(n15758), .dinb(n15757), .dout(n15759));
  jor  g15510(.dina(n15759), .dinb(n15683), .dout(n15760));
  jor  g15511(.dina(n15760), .dinb(asqrt[32] ), .dout(n15761));
  jand g15512(.dina(n15399), .dinb(n15761), .dout(n15762));
  jor  g15513(.dina(n15762), .dinb(n15682), .dout(n15763));
  jor  g15514(.dina(n15763), .dinb(asqrt[33] ), .dout(n15764));
  jnot g15515(.din(n15407), .dout(n15765));
  jand g15516(.dina(n15765), .dinb(n15764), .dout(n15766));
  jor  g15517(.dina(n15766), .dinb(n15681), .dout(n15767));
  jor  g15518(.dina(n15767), .dinb(asqrt[34] ), .dout(n15768));
  jnot g15519(.din(n15414), .dout(n15769));
  jand g15520(.dina(n15769), .dinb(n15768), .dout(n15770));
  jor  g15521(.dina(n15770), .dinb(n15680), .dout(n15771));
  jor  g15522(.dina(n15771), .dinb(asqrt[35] ), .dout(n15772));
  jnot g15523(.din(n15421), .dout(n15773));
  jand g15524(.dina(n15773), .dinb(n15772), .dout(n15774));
  jor  g15525(.dina(n15774), .dinb(n15679), .dout(n15775));
  jor  g15526(.dina(n15775), .dinb(asqrt[36] ), .dout(n15776));
  jand g15527(.dina(n15428), .dinb(n15776), .dout(n15777));
  jor  g15528(.dina(n15777), .dinb(n15678), .dout(n15778));
  jor  g15529(.dina(n15778), .dinb(asqrt[37] ), .dout(n15779));
  jnot g15530(.din(n15436), .dout(n15780));
  jand g15531(.dina(n15780), .dinb(n15779), .dout(n15781));
  jor  g15532(.dina(n15781), .dinb(n15677), .dout(n15782));
  jor  g15533(.dina(n15782), .dinb(asqrt[38] ), .dout(n15783));
  jand g15534(.dina(n15443), .dinb(n15783), .dout(n15784));
  jor  g15535(.dina(n15784), .dinb(n15676), .dout(n15785));
  jor  g15536(.dina(n15785), .dinb(asqrt[39] ), .dout(n15786));
  jnot g15537(.din(n15451), .dout(n15787));
  jand g15538(.dina(n15787), .dinb(n15786), .dout(n15788));
  jor  g15539(.dina(n15788), .dinb(n15675), .dout(n15789));
  jor  g15540(.dina(n15789), .dinb(asqrt[40] ), .dout(n15790));
  jnot g15541(.din(n15458), .dout(n15791));
  jand g15542(.dina(n15791), .dinb(n15790), .dout(n15792));
  jor  g15543(.dina(n15792), .dinb(n15674), .dout(n15793));
  jor  g15544(.dina(n15793), .dinb(asqrt[41] ), .dout(n15794));
  jnot g15545(.din(n15465), .dout(n15795));
  jand g15546(.dina(n15795), .dinb(n15794), .dout(n15796));
  jor  g15547(.dina(n15796), .dinb(n15673), .dout(n15797));
  jor  g15548(.dina(n15797), .dinb(asqrt[42] ), .dout(n15798));
  jand g15549(.dina(n15472), .dinb(n15798), .dout(n15799));
  jor  g15550(.dina(n15799), .dinb(n15672), .dout(n15800));
  jor  g15551(.dina(n15800), .dinb(asqrt[43] ), .dout(n15801));
  jnot g15552(.din(n15480), .dout(n15802));
  jand g15553(.dina(n15802), .dinb(n15801), .dout(n15803));
  jor  g15554(.dina(n15803), .dinb(n15671), .dout(n15804));
  jor  g15555(.dina(n15804), .dinb(asqrt[44] ), .dout(n15805));
  jand g15556(.dina(n15487), .dinb(n15805), .dout(n15806));
  jor  g15557(.dina(n15806), .dinb(n15670), .dout(n15807));
  jor  g15558(.dina(n15807), .dinb(asqrt[45] ), .dout(n15808));
  jnot g15559(.din(n15495), .dout(n15809));
  jand g15560(.dina(n15809), .dinb(n15808), .dout(n15810));
  jor  g15561(.dina(n15810), .dinb(n15669), .dout(n15811));
  jor  g15562(.dina(n15811), .dinb(asqrt[46] ), .dout(n15812));
  jnot g15563(.din(n15502), .dout(n15813));
  jand g15564(.dina(n15813), .dinb(n15812), .dout(n15814));
  jor  g15565(.dina(n15814), .dinb(n15668), .dout(n15815));
  jor  g15566(.dina(n15815), .dinb(asqrt[47] ), .dout(n15816));
  jand g15567(.dina(n15509), .dinb(n15816), .dout(n15817));
  jor  g15568(.dina(n15817), .dinb(n15667), .dout(n15818));
  jor  g15569(.dina(n15818), .dinb(asqrt[48] ), .dout(n15819));
  jand g15570(.dina(n15819), .dinb(n15516), .dout(n15820));
  jor  g15571(.dina(n15820), .dinb(n15666), .dout(n15821));
  jor  g15572(.dina(n15821), .dinb(asqrt[49] ), .dout(n15822));
  jnot g15573(.din(n15525), .dout(n15823));
  jand g15574(.dina(n15823), .dinb(n15822), .dout(n15824));
  jor  g15575(.dina(n15824), .dinb(n15665), .dout(n15825));
  jor  g15576(.dina(n15825), .dinb(asqrt[50] ), .dout(n15826));
  jand g15577(.dina(n15532), .dinb(n15826), .dout(n15827));
  jor  g15578(.dina(n15827), .dinb(n15664), .dout(n15828));
  jor  g15579(.dina(n15828), .dinb(asqrt[51] ), .dout(n15829));
  jnot g15580(.din(n15540), .dout(n15830));
  jand g15581(.dina(n15830), .dinb(n15829), .dout(n15831));
  jor  g15582(.dina(n15831), .dinb(n15663), .dout(n15832));
  jor  g15583(.dina(n15832), .dinb(asqrt[52] ), .dout(n15833));
  jand g15584(.dina(n15547), .dinb(n15833), .dout(n15834));
  jor  g15585(.dina(n15834), .dinb(n15662), .dout(n15835));
  jor  g15586(.dina(n15835), .dinb(asqrt[53] ), .dout(n15836));
  jnot g15587(.din(n15555), .dout(n15837));
  jand g15588(.dina(n15837), .dinb(n15836), .dout(n15838));
  jor  g15589(.dina(n15838), .dinb(n15661), .dout(n15839));
  jor  g15590(.dina(n15839), .dinb(asqrt[54] ), .dout(n15840));
  jnot g15591(.din(n15562), .dout(n15841));
  jand g15592(.dina(n15841), .dinb(n15840), .dout(n15842));
  jor  g15593(.dina(n15842), .dinb(n15660), .dout(n15843));
  jor  g15594(.dina(n15843), .dinb(asqrt[55] ), .dout(n15844));
  jnot g15595(.din(n15569), .dout(n15845));
  jand g15596(.dina(n15845), .dinb(n15844), .dout(n15846));
  jor  g15597(.dina(n15846), .dinb(n15659), .dout(n15847));
  jor  g15598(.dina(n15847), .dinb(asqrt[56] ), .dout(n15848));
  jand g15599(.dina(n15576), .dinb(n15848), .dout(n15849));
  jor  g15600(.dina(n15849), .dinb(n15658), .dout(n15850));
  jor  g15601(.dina(n15850), .dinb(asqrt[57] ), .dout(n15851));
  jnot g15602(.din(n15584), .dout(n15852));
  jand g15603(.dina(n15852), .dinb(n15851), .dout(n15853));
  jor  g15604(.dina(n15853), .dinb(n15657), .dout(n15854));
  jor  g15605(.dina(n15854), .dinb(asqrt[58] ), .dout(n15855));
  jand g15606(.dina(n15591), .dinb(n15855), .dout(n15856));
  jor  g15607(.dina(n15856), .dinb(n15656), .dout(n15857));
  jor  g15608(.dina(n15857), .dinb(asqrt[59] ), .dout(n15858));
  jnot g15609(.din(n15599), .dout(n15859));
  jand g15610(.dina(n15859), .dinb(n15858), .dout(n15860));
  jor  g15611(.dina(n15860), .dinb(n15655), .dout(n15861));
  jor  g15612(.dina(n15861), .dinb(asqrt[60] ), .dout(n15862));
  jand g15613(.dina(n15606), .dinb(n15862), .dout(n15863));
  jor  g15614(.dina(n15863), .dinb(n15654), .dout(n15864));
  jor  g15615(.dina(n15864), .dinb(asqrt[61] ), .dout(n15865));
  jnot g15616(.din(n15614), .dout(n15866));
  jand g15617(.dina(n15866), .dinb(n15865), .dout(n15867));
  jor  g15618(.dina(n15867), .dinb(n15653), .dout(n15868));
  jor  g15619(.dina(n15868), .dinb(asqrt[62] ), .dout(n15869));
  jand g15620(.dina(n15621), .dinb(n15869), .dout(n15870));
  jor  g15621(.dina(n15870), .dinb(n15652), .dout(n15871));
  jand g15622(.dina(n15871), .dinb(n15263), .dout(n15872));
  jnot g15623(.din(n15626), .dout(n15873));
  jand g15624(.dina(n15873), .dinb(n15872), .dout(n15874));
  jand g15625(.dina(n15874), .dinb(n15256), .dout(n15875));
  jor  g15626(.dina(n15875), .dinb(asqrt[63] ), .dout(n15876));
  jnot g15627(.din(n15639), .dout(n15877));
  jand g15628(.dina(n15877), .dinb(n15876), .dout(n15878));
  jor  g15629(.dina(n15878), .dinb(n15651), .dout(n15879));
  jand g15630(.dina(n15879), .dinb(n15650), .dout(n15880));
  jand g15631(.dina(n15880), .dinb(n15648), .dout(n15881));
  jor  g15632(.dina(n15881), .dinb(n15647), .dout(n15882));
  jand g15633(.dina(n15882), .dinb(asqrt[16] ), .dout(n15883));
  jor  g15634(.dina(n15882), .dinb(asqrt[16] ), .dout(n15884));
  jand g15635(.dina(asqrt[14] ), .dinb(n15267), .dout(n15885));
  jnot g15636(.din(n15631), .dout(n15886));
  jand g15637(.dina(n15636), .dinb(asqrt[15] ), .dout(n15887));
  jand g15638(.dina(n15887), .dinb(n15886), .dout(n15888));
  jand g15639(.dina(n15888), .dinb(n15876), .dout(n15889));
  jor  g15640(.dina(n15889), .dinb(n15885), .dout(n15890));
  jxor g15641(.dina(n15890), .dinb(a[30] ), .dout(n15891));
  jnot g15642(.din(n15891), .dout(n15892));
  jand g15643(.dina(n15892), .dinb(n15884), .dout(n15893));
  jor  g15644(.dina(n15893), .dinb(n15883), .dout(n15894));
  jand g15645(.dina(n15894), .dinb(asqrt[17] ), .dout(n15895));
  jor  g15646(.dina(n15894), .dinb(asqrt[17] ), .dout(n15896));
  jxor g15647(.dina(n15271), .dinb(n14674), .dout(n15897));
  jand g15648(.dina(n15897), .dinb(asqrt[14] ), .dout(n15898));
  jxor g15649(.dina(n15898), .dinb(n15704), .dout(n15899));
  jand g15650(.dina(n15899), .dinb(n15896), .dout(n15900));
  jor  g15651(.dina(n15900), .dinb(n15895), .dout(n15901));
  jand g15652(.dina(n15901), .dinb(asqrt[18] ), .dout(n15902));
  jor  g15653(.dina(n15901), .dinb(asqrt[18] ), .dout(n15903));
  jxor g15654(.dina(n15279), .dinb(n14078), .dout(n15904));
  jand g15655(.dina(n15904), .dinb(asqrt[14] ), .dout(n15905));
  jxor g15656(.dina(n15905), .dinb(n15708), .dout(n15906));
  jand g15657(.dina(n15906), .dinb(n15903), .dout(n15907));
  jor  g15658(.dina(n15907), .dinb(n15902), .dout(n15908));
  jand g15659(.dina(n15908), .dinb(asqrt[19] ), .dout(n15909));
  jor  g15660(.dina(n15908), .dinb(asqrt[19] ), .dout(n15910));
  jxor g15661(.dina(n15290), .dinb(n13515), .dout(n15911));
  jand g15662(.dina(n15911), .dinb(asqrt[14] ), .dout(n15912));
  jxor g15663(.dina(n15912), .dinb(n15295), .dout(n15913));
  jand g15664(.dina(n15913), .dinb(n15910), .dout(n15914));
  jor  g15665(.dina(n15914), .dinb(n15909), .dout(n15915));
  jand g15666(.dina(n15915), .dinb(asqrt[20] ), .dout(n15916));
  jor  g15667(.dina(n15915), .dinb(asqrt[20] ), .dout(n15917));
  jxor g15668(.dina(n15298), .dinb(n12947), .dout(n15918));
  jand g15669(.dina(n15918), .dinb(asqrt[14] ), .dout(n15919));
  jxor g15670(.dina(n15919), .dinb(n15303), .dout(n15920));
  jnot g15671(.din(n15920), .dout(n15921));
  jand g15672(.dina(n15921), .dinb(n15917), .dout(n15922));
  jor  g15673(.dina(n15922), .dinb(n15916), .dout(n15923));
  jand g15674(.dina(n15923), .dinb(asqrt[21] ), .dout(n15924));
  jor  g15675(.dina(n15923), .dinb(asqrt[21] ), .dout(n15925));
  jxor g15676(.dina(n15305), .dinb(n12410), .dout(n15926));
  jand g15677(.dina(n15926), .dinb(asqrt[14] ), .dout(n15927));
  jxor g15678(.dina(n15927), .dinb(n15310), .dout(n15928));
  jand g15679(.dina(n15928), .dinb(n15925), .dout(n15929));
  jor  g15680(.dina(n15929), .dinb(n15924), .dout(n15930));
  jand g15681(.dina(n15930), .dinb(asqrt[22] ), .dout(n15931));
  jor  g15682(.dina(n15930), .dinb(asqrt[22] ), .dout(n15932));
  jxor g15683(.dina(n15313), .dinb(n11858), .dout(n15933));
  jand g15684(.dina(n15933), .dinb(asqrt[14] ), .dout(n15934));
  jxor g15685(.dina(n15934), .dinb(n15318), .dout(n15935));
  jnot g15686(.din(n15935), .dout(n15936));
  jand g15687(.dina(n15936), .dinb(n15932), .dout(n15937));
  jor  g15688(.dina(n15937), .dinb(n15931), .dout(n15938));
  jand g15689(.dina(n15938), .dinb(asqrt[23] ), .dout(n15939));
  jor  g15690(.dina(n15938), .dinb(asqrt[23] ), .dout(n15940));
  jxor g15691(.dina(n15320), .dinb(n11347), .dout(n15941));
  jand g15692(.dina(n15941), .dinb(asqrt[14] ), .dout(n15942));
  jxor g15693(.dina(n15942), .dinb(n15325), .dout(n15943));
  jand g15694(.dina(n15943), .dinb(n15940), .dout(n15944));
  jor  g15695(.dina(n15944), .dinb(n15939), .dout(n15945));
  jand g15696(.dina(n15945), .dinb(asqrt[24] ), .dout(n15946));
  jor  g15697(.dina(n15945), .dinb(asqrt[24] ), .dout(n15947));
  jxor g15698(.dina(n15328), .dinb(n10824), .dout(n15948));
  jand g15699(.dina(n15948), .dinb(asqrt[14] ), .dout(n15949));
  jxor g15700(.dina(n15949), .dinb(n15333), .dout(n15950));
  jnot g15701(.din(n15950), .dout(n15951));
  jand g15702(.dina(n15951), .dinb(n15947), .dout(n15952));
  jor  g15703(.dina(n15952), .dinb(n15946), .dout(n15953));
  jand g15704(.dina(n15953), .dinb(asqrt[25] ), .dout(n15954));
  jor  g15705(.dina(n15953), .dinb(asqrt[25] ), .dout(n15955));
  jxor g15706(.dina(n15335), .dinb(n10328), .dout(n15956));
  jand g15707(.dina(n15956), .dinb(asqrt[14] ), .dout(n15957));
  jxor g15708(.dina(n15957), .dinb(n15340), .dout(n15958));
  jnot g15709(.din(n15958), .dout(n15959));
  jand g15710(.dina(n15959), .dinb(n15955), .dout(n15960));
  jor  g15711(.dina(n15960), .dinb(n15954), .dout(n15961));
  jand g15712(.dina(n15961), .dinb(asqrt[26] ), .dout(n15962));
  jor  g15713(.dina(n15961), .dinb(asqrt[26] ), .dout(n15963));
  jxor g15714(.dina(n15342), .dinb(n9832), .dout(n15964));
  jand g15715(.dina(n15964), .dinb(asqrt[14] ), .dout(n15965));
  jxor g15716(.dina(n15965), .dinb(n15347), .dout(n15966));
  jnot g15717(.din(n15966), .dout(n15967));
  jand g15718(.dina(n15967), .dinb(n15963), .dout(n15968));
  jor  g15719(.dina(n15968), .dinb(n15962), .dout(n15969));
  jand g15720(.dina(n15969), .dinb(asqrt[27] ), .dout(n15970));
  jor  g15721(.dina(n15969), .dinb(asqrt[27] ), .dout(n15971));
  jxor g15722(.dina(n15349), .dinb(n9369), .dout(n15972));
  jand g15723(.dina(n15972), .dinb(asqrt[14] ), .dout(n15973));
  jxor g15724(.dina(n15973), .dinb(n15354), .dout(n15974));
  jand g15725(.dina(n15974), .dinb(n15971), .dout(n15975));
  jor  g15726(.dina(n15975), .dinb(n15970), .dout(n15976));
  jand g15727(.dina(n15976), .dinb(asqrt[28] ), .dout(n15977));
  jor  g15728(.dina(n15976), .dinb(asqrt[28] ), .dout(n15978));
  jxor g15729(.dina(n15357), .dinb(n8890), .dout(n15979));
  jand g15730(.dina(n15979), .dinb(asqrt[14] ), .dout(n15980));
  jxor g15731(.dina(n15980), .dinb(n15362), .dout(n15981));
  jnot g15732(.din(n15981), .dout(n15982));
  jand g15733(.dina(n15982), .dinb(n15978), .dout(n15983));
  jor  g15734(.dina(n15983), .dinb(n15977), .dout(n15984));
  jand g15735(.dina(n15984), .dinb(asqrt[29] ), .dout(n15985));
  jor  g15736(.dina(n15984), .dinb(asqrt[29] ), .dout(n15986));
  jxor g15737(.dina(n15364), .dinb(n8449), .dout(n15987));
  jand g15738(.dina(n15987), .dinb(asqrt[14] ), .dout(n15988));
  jxor g15739(.dina(n15988), .dinb(n15369), .dout(n15989));
  jand g15740(.dina(n15989), .dinb(n15986), .dout(n15990));
  jor  g15741(.dina(n15990), .dinb(n15985), .dout(n15991));
  jand g15742(.dina(n15991), .dinb(asqrt[30] ), .dout(n15992));
  jor  g15743(.dina(n15991), .dinb(asqrt[30] ), .dout(n15993));
  jxor g15744(.dina(n15372), .dinb(n8003), .dout(n15994));
  jand g15745(.dina(n15994), .dinb(asqrt[14] ), .dout(n15995));
  jxor g15746(.dina(n15995), .dinb(n15377), .dout(n15996));
  jnot g15747(.din(n15996), .dout(n15997));
  jand g15748(.dina(n15997), .dinb(n15993), .dout(n15998));
  jor  g15749(.dina(n15998), .dinb(n15992), .dout(n15999));
  jand g15750(.dina(n15999), .dinb(asqrt[31] ), .dout(n16000));
  jor  g15751(.dina(n15999), .dinb(asqrt[31] ), .dout(n16001));
  jxor g15752(.dina(n15379), .dinb(n7581), .dout(n16002));
  jand g15753(.dina(n16002), .dinb(asqrt[14] ), .dout(n16003));
  jxor g15754(.dina(n16003), .dinb(n15384), .dout(n16004));
  jand g15755(.dina(n16004), .dinb(n16001), .dout(n16005));
  jor  g15756(.dina(n16005), .dinb(n16000), .dout(n16006));
  jand g15757(.dina(n16006), .dinb(asqrt[32] ), .dout(n16007));
  jor  g15758(.dina(n16006), .dinb(asqrt[32] ), .dout(n16008));
  jxor g15759(.dina(n15387), .dinb(n7154), .dout(n16009));
  jand g15760(.dina(n16009), .dinb(asqrt[14] ), .dout(n16010));
  jxor g15761(.dina(n16010), .dinb(n15392), .dout(n16011));
  jnot g15762(.din(n16011), .dout(n16012));
  jand g15763(.dina(n16012), .dinb(n16008), .dout(n16013));
  jor  g15764(.dina(n16013), .dinb(n16007), .dout(n16014));
  jand g15765(.dina(n16014), .dinb(asqrt[33] ), .dout(n16015));
  jor  g15766(.dina(n16014), .dinb(asqrt[33] ), .dout(n16016));
  jxor g15767(.dina(n15394), .dinb(n6758), .dout(n16017));
  jand g15768(.dina(n16017), .dinb(asqrt[14] ), .dout(n16018));
  jxor g15769(.dina(n16018), .dinb(n15399), .dout(n16019));
  jand g15770(.dina(n16019), .dinb(n16016), .dout(n16020));
  jor  g15771(.dina(n16020), .dinb(n16015), .dout(n16021));
  jand g15772(.dina(n16021), .dinb(asqrt[34] ), .dout(n16022));
  jor  g15773(.dina(n16021), .dinb(asqrt[34] ), .dout(n16023));
  jxor g15774(.dina(n15402), .dinb(n6357), .dout(n16024));
  jand g15775(.dina(n16024), .dinb(asqrt[14] ), .dout(n16025));
  jxor g15776(.dina(n16025), .dinb(n15407), .dout(n16026));
  jnot g15777(.din(n16026), .dout(n16027));
  jand g15778(.dina(n16027), .dinb(n16023), .dout(n16028));
  jor  g15779(.dina(n16028), .dinb(n16022), .dout(n16029));
  jand g15780(.dina(n16029), .dinb(asqrt[35] ), .dout(n16030));
  jor  g15781(.dina(n16029), .dinb(asqrt[35] ), .dout(n16031));
  jxor g15782(.dina(n15409), .dinb(n5989), .dout(n16032));
  jand g15783(.dina(n16032), .dinb(asqrt[14] ), .dout(n16033));
  jxor g15784(.dina(n16033), .dinb(n15414), .dout(n16034));
  jnot g15785(.din(n16034), .dout(n16035));
  jand g15786(.dina(n16035), .dinb(n16031), .dout(n16036));
  jor  g15787(.dina(n16036), .dinb(n16030), .dout(n16037));
  jand g15788(.dina(n16037), .dinb(asqrt[36] ), .dout(n16038));
  jor  g15789(.dina(n16037), .dinb(asqrt[36] ), .dout(n16039));
  jxor g15790(.dina(n15416), .dinb(n5606), .dout(n16040));
  jand g15791(.dina(n16040), .dinb(asqrt[14] ), .dout(n16041));
  jxor g15792(.dina(n16041), .dinb(n15421), .dout(n16042));
  jnot g15793(.din(n16042), .dout(n16043));
  jand g15794(.dina(n16043), .dinb(n16039), .dout(n16044));
  jor  g15795(.dina(n16044), .dinb(n16038), .dout(n16045));
  jand g15796(.dina(n16045), .dinb(asqrt[37] ), .dout(n16046));
  jor  g15797(.dina(n16045), .dinb(asqrt[37] ), .dout(n16047));
  jxor g15798(.dina(n15423), .dinb(n5259), .dout(n16048));
  jand g15799(.dina(n16048), .dinb(asqrt[14] ), .dout(n16049));
  jxor g15800(.dina(n16049), .dinb(n15428), .dout(n16050));
  jand g15801(.dina(n16050), .dinb(n16047), .dout(n16051));
  jor  g15802(.dina(n16051), .dinb(n16046), .dout(n16052));
  jand g15803(.dina(n16052), .dinb(asqrt[38] ), .dout(n16053));
  jor  g15804(.dina(n16052), .dinb(asqrt[38] ), .dout(n16054));
  jxor g15805(.dina(n15431), .dinb(n4902), .dout(n16055));
  jand g15806(.dina(n16055), .dinb(asqrt[14] ), .dout(n16056));
  jxor g15807(.dina(n16056), .dinb(n15436), .dout(n16057));
  jnot g15808(.din(n16057), .dout(n16058));
  jand g15809(.dina(n16058), .dinb(n16054), .dout(n16059));
  jor  g15810(.dina(n16059), .dinb(n16053), .dout(n16060));
  jand g15811(.dina(n16060), .dinb(asqrt[39] ), .dout(n16061));
  jor  g15812(.dina(n16060), .dinb(asqrt[39] ), .dout(n16062));
  jxor g15813(.dina(n15438), .dinb(n4582), .dout(n16063));
  jand g15814(.dina(n16063), .dinb(asqrt[14] ), .dout(n16064));
  jxor g15815(.dina(n16064), .dinb(n15443), .dout(n16065));
  jand g15816(.dina(n16065), .dinb(n16062), .dout(n16066));
  jor  g15817(.dina(n16066), .dinb(n16061), .dout(n16067));
  jand g15818(.dina(n16067), .dinb(asqrt[40] ), .dout(n16068));
  jor  g15819(.dina(n16067), .dinb(asqrt[40] ), .dout(n16069));
  jxor g15820(.dina(n15446), .dinb(n4249), .dout(n16070));
  jand g15821(.dina(n16070), .dinb(asqrt[14] ), .dout(n16071));
  jxor g15822(.dina(n16071), .dinb(n15451), .dout(n16072));
  jnot g15823(.din(n16072), .dout(n16073));
  jand g15824(.dina(n16073), .dinb(n16069), .dout(n16074));
  jor  g15825(.dina(n16074), .dinb(n16068), .dout(n16075));
  jand g15826(.dina(n16075), .dinb(asqrt[41] ), .dout(n16076));
  jor  g15827(.dina(n16075), .dinb(asqrt[41] ), .dout(n16077));
  jxor g15828(.dina(n15453), .dinb(n3955), .dout(n16078));
  jand g15829(.dina(n16078), .dinb(asqrt[14] ), .dout(n16079));
  jxor g15830(.dina(n16079), .dinb(n15458), .dout(n16080));
  jnot g15831(.din(n16080), .dout(n16081));
  jand g15832(.dina(n16081), .dinb(n16077), .dout(n16082));
  jor  g15833(.dina(n16082), .dinb(n16076), .dout(n16083));
  jand g15834(.dina(n16083), .dinb(asqrt[42] ), .dout(n16084));
  jor  g15835(.dina(n16083), .dinb(asqrt[42] ), .dout(n16085));
  jxor g15836(.dina(n15460), .dinb(n3642), .dout(n16086));
  jand g15837(.dina(n16086), .dinb(asqrt[14] ), .dout(n16087));
  jxor g15838(.dina(n16087), .dinb(n15465), .dout(n16088));
  jnot g15839(.din(n16088), .dout(n16089));
  jand g15840(.dina(n16089), .dinb(n16085), .dout(n16090));
  jor  g15841(.dina(n16090), .dinb(n16084), .dout(n16091));
  jand g15842(.dina(n16091), .dinb(asqrt[43] ), .dout(n16092));
  jor  g15843(.dina(n16091), .dinb(asqrt[43] ), .dout(n16093));
  jxor g15844(.dina(n15467), .dinb(n3368), .dout(n16094));
  jand g15845(.dina(n16094), .dinb(asqrt[14] ), .dout(n16095));
  jxor g15846(.dina(n16095), .dinb(n15472), .dout(n16096));
  jand g15847(.dina(n16096), .dinb(n16093), .dout(n16097));
  jor  g15848(.dina(n16097), .dinb(n16092), .dout(n16098));
  jand g15849(.dina(n16098), .dinb(asqrt[44] ), .dout(n16099));
  jor  g15850(.dina(n16098), .dinb(asqrt[44] ), .dout(n16100));
  jxor g15851(.dina(n15475), .dinb(n3089), .dout(n16101));
  jand g15852(.dina(n16101), .dinb(asqrt[14] ), .dout(n16102));
  jxor g15853(.dina(n16102), .dinb(n15480), .dout(n16103));
  jnot g15854(.din(n16103), .dout(n16104));
  jand g15855(.dina(n16104), .dinb(n16100), .dout(n16105));
  jor  g15856(.dina(n16105), .dinb(n16099), .dout(n16106));
  jand g15857(.dina(n16106), .dinb(asqrt[45] ), .dout(n16107));
  jor  g15858(.dina(n16106), .dinb(asqrt[45] ), .dout(n16108));
  jxor g15859(.dina(n15482), .dinb(n2833), .dout(n16109));
  jand g15860(.dina(n16109), .dinb(asqrt[14] ), .dout(n16110));
  jxor g15861(.dina(n16110), .dinb(n15487), .dout(n16111));
  jand g15862(.dina(n16111), .dinb(n16108), .dout(n16112));
  jor  g15863(.dina(n16112), .dinb(n16107), .dout(n16113));
  jand g15864(.dina(n16113), .dinb(asqrt[46] ), .dout(n16114));
  jor  g15865(.dina(n16113), .dinb(asqrt[46] ), .dout(n16115));
  jxor g15866(.dina(n15490), .dinb(n2572), .dout(n16116));
  jand g15867(.dina(n16116), .dinb(asqrt[14] ), .dout(n16117));
  jxor g15868(.dina(n16117), .dinb(n15495), .dout(n16118));
  jnot g15869(.din(n16118), .dout(n16119));
  jand g15870(.dina(n16119), .dinb(n16115), .dout(n16120));
  jor  g15871(.dina(n16120), .dinb(n16114), .dout(n16121));
  jand g15872(.dina(n16121), .dinb(asqrt[47] ), .dout(n16122));
  jor  g15873(.dina(n16121), .dinb(asqrt[47] ), .dout(n16123));
  jxor g15874(.dina(n15497), .dinb(n2345), .dout(n16124));
  jand g15875(.dina(n16124), .dinb(asqrt[14] ), .dout(n16125));
  jxor g15876(.dina(n16125), .dinb(n15502), .dout(n16126));
  jnot g15877(.din(n16126), .dout(n16127));
  jand g15878(.dina(n16127), .dinb(n16123), .dout(n16128));
  jor  g15879(.dina(n16128), .dinb(n16122), .dout(n16129));
  jand g15880(.dina(n16129), .dinb(asqrt[48] ), .dout(n16130));
  jor  g15881(.dina(n16129), .dinb(asqrt[48] ), .dout(n16131));
  jxor g15882(.dina(n15504), .dinb(n2108), .dout(n16132));
  jand g15883(.dina(n16132), .dinb(asqrt[14] ), .dout(n16133));
  jxor g15884(.dina(n16133), .dinb(n15509), .dout(n16134));
  jand g15885(.dina(n16134), .dinb(n16131), .dout(n16135));
  jor  g15886(.dina(n16135), .dinb(n16130), .dout(n16136));
  jand g15887(.dina(n16136), .dinb(asqrt[49] ), .dout(n16137));
  jxor g15888(.dina(n15512), .dinb(n1912), .dout(n16138));
  jand g15889(.dina(n16138), .dinb(asqrt[14] ), .dout(n16139));
  jxor g15890(.dina(n16139), .dinb(n15516), .dout(n16140));
  jor  g15891(.dina(n16136), .dinb(asqrt[49] ), .dout(n16141));
  jand g15892(.dina(n16141), .dinb(n16140), .dout(n16142));
  jor  g15893(.dina(n16142), .dinb(n16137), .dout(n16143));
  jand g15894(.dina(n16143), .dinb(asqrt[50] ), .dout(n16144));
  jor  g15895(.dina(n16143), .dinb(asqrt[50] ), .dout(n16145));
  jxor g15896(.dina(n15520), .dinb(n1699), .dout(n16146));
  jand g15897(.dina(n16146), .dinb(asqrt[14] ), .dout(n16147));
  jxor g15898(.dina(n16147), .dinb(n15525), .dout(n16148));
  jnot g15899(.din(n16148), .dout(n16149));
  jand g15900(.dina(n16149), .dinb(n16145), .dout(n16150));
  jor  g15901(.dina(n16150), .dinb(n16144), .dout(n16151));
  jand g15902(.dina(n16151), .dinb(asqrt[51] ), .dout(n16152));
  jor  g15903(.dina(n16151), .dinb(asqrt[51] ), .dout(n16153));
  jxor g15904(.dina(n15527), .dinb(n1516), .dout(n16154));
  jand g15905(.dina(n16154), .dinb(asqrt[14] ), .dout(n16155));
  jxor g15906(.dina(n16155), .dinb(n15532), .dout(n16156));
  jand g15907(.dina(n16156), .dinb(n16153), .dout(n16157));
  jor  g15908(.dina(n16157), .dinb(n16152), .dout(n16158));
  jand g15909(.dina(n16158), .dinb(asqrt[52] ), .dout(n16159));
  jor  g15910(.dina(n16158), .dinb(asqrt[52] ), .dout(n16160));
  jxor g15911(.dina(n15535), .dinb(n1332), .dout(n16161));
  jand g15912(.dina(n16161), .dinb(asqrt[14] ), .dout(n16162));
  jxor g15913(.dina(n16162), .dinb(n15540), .dout(n16163));
  jnot g15914(.din(n16163), .dout(n16164));
  jand g15915(.dina(n16164), .dinb(n16160), .dout(n16165));
  jor  g15916(.dina(n16165), .dinb(n16159), .dout(n16166));
  jand g15917(.dina(n16166), .dinb(asqrt[53] ), .dout(n16167));
  jor  g15918(.dina(n16166), .dinb(asqrt[53] ), .dout(n16168));
  jxor g15919(.dina(n15542), .dinb(n1173), .dout(n16169));
  jand g15920(.dina(n16169), .dinb(asqrt[14] ), .dout(n16170));
  jxor g15921(.dina(n16170), .dinb(n15547), .dout(n16171));
  jand g15922(.dina(n16171), .dinb(n16168), .dout(n16172));
  jor  g15923(.dina(n16172), .dinb(n16167), .dout(n16173));
  jand g15924(.dina(n16173), .dinb(asqrt[54] ), .dout(n16174));
  jor  g15925(.dina(n16173), .dinb(asqrt[54] ), .dout(n16175));
  jxor g15926(.dina(n15550), .dinb(n1008), .dout(n16176));
  jand g15927(.dina(n16176), .dinb(asqrt[14] ), .dout(n16177));
  jxor g15928(.dina(n16177), .dinb(n15555), .dout(n16178));
  jnot g15929(.din(n16178), .dout(n16179));
  jand g15930(.dina(n16179), .dinb(n16175), .dout(n16180));
  jor  g15931(.dina(n16180), .dinb(n16174), .dout(n16181));
  jand g15932(.dina(n16181), .dinb(asqrt[55] ), .dout(n16182));
  jor  g15933(.dina(n16181), .dinb(asqrt[55] ), .dout(n16183));
  jxor g15934(.dina(n15557), .dinb(n884), .dout(n16184));
  jand g15935(.dina(n16184), .dinb(asqrt[14] ), .dout(n16185));
  jxor g15936(.dina(n16185), .dinb(n15562), .dout(n16186));
  jnot g15937(.din(n16186), .dout(n16187));
  jand g15938(.dina(n16187), .dinb(n16183), .dout(n16188));
  jor  g15939(.dina(n16188), .dinb(n16182), .dout(n16189));
  jand g15940(.dina(n16189), .dinb(asqrt[56] ), .dout(n16190));
  jor  g15941(.dina(n16189), .dinb(asqrt[56] ), .dout(n16191));
  jxor g15942(.dina(n15564), .dinb(n743), .dout(n16192));
  jand g15943(.dina(n16192), .dinb(asqrt[14] ), .dout(n16193));
  jxor g15944(.dina(n16193), .dinb(n15569), .dout(n16194));
  jnot g15945(.din(n16194), .dout(n16195));
  jand g15946(.dina(n16195), .dinb(n16191), .dout(n16196));
  jor  g15947(.dina(n16196), .dinb(n16190), .dout(n16197));
  jand g15948(.dina(n16197), .dinb(asqrt[57] ), .dout(n16198));
  jor  g15949(.dina(n16197), .dinb(asqrt[57] ), .dout(n16199));
  jxor g15950(.dina(n15571), .dinb(n635), .dout(n16200));
  jand g15951(.dina(n16200), .dinb(asqrt[14] ), .dout(n16201));
  jxor g15952(.dina(n16201), .dinb(n15576), .dout(n16202));
  jand g15953(.dina(n16202), .dinb(n16199), .dout(n16203));
  jor  g15954(.dina(n16203), .dinb(n16198), .dout(n16204));
  jand g15955(.dina(n16204), .dinb(asqrt[58] ), .dout(n16205));
  jor  g15956(.dina(n16204), .dinb(asqrt[58] ), .dout(n16206));
  jxor g15957(.dina(n15579), .dinb(n515), .dout(n16207));
  jand g15958(.dina(n16207), .dinb(asqrt[14] ), .dout(n16208));
  jxor g15959(.dina(n16208), .dinb(n15584), .dout(n16209));
  jnot g15960(.din(n16209), .dout(n16210));
  jand g15961(.dina(n16210), .dinb(n16206), .dout(n16211));
  jor  g15962(.dina(n16211), .dinb(n16205), .dout(n16212));
  jand g15963(.dina(n16212), .dinb(asqrt[59] ), .dout(n16213));
  jor  g15964(.dina(n16212), .dinb(asqrt[59] ), .dout(n16214));
  jxor g15965(.dina(n15586), .dinb(n443), .dout(n16215));
  jand g15966(.dina(n16215), .dinb(asqrt[14] ), .dout(n16216));
  jxor g15967(.dina(n16216), .dinb(n15591), .dout(n16217));
  jand g15968(.dina(n16217), .dinb(n16214), .dout(n16218));
  jor  g15969(.dina(n16218), .dinb(n16213), .dout(n16219));
  jand g15970(.dina(n16219), .dinb(asqrt[60] ), .dout(n16220));
  jor  g15971(.dina(n16219), .dinb(asqrt[60] ), .dout(n16221));
  jxor g15972(.dina(n15594), .dinb(n352), .dout(n16222));
  jand g15973(.dina(n16222), .dinb(asqrt[14] ), .dout(n16223));
  jxor g15974(.dina(n16223), .dinb(n15599), .dout(n16224));
  jnot g15975(.din(n16224), .dout(n16225));
  jand g15976(.dina(n16225), .dinb(n16221), .dout(n16226));
  jor  g15977(.dina(n16226), .dinb(n16220), .dout(n16227));
  jand g15978(.dina(n16227), .dinb(asqrt[61] ), .dout(n16228));
  jor  g15979(.dina(n16227), .dinb(asqrt[61] ), .dout(n16229));
  jxor g15980(.dina(n15601), .dinb(n294), .dout(n16230));
  jand g15981(.dina(n16230), .dinb(asqrt[14] ), .dout(n16231));
  jxor g15982(.dina(n16231), .dinb(n15606), .dout(n16232));
  jand g15983(.dina(n16232), .dinb(n16229), .dout(n16233));
  jor  g15984(.dina(n16233), .dinb(n16228), .dout(n16234));
  jand g15985(.dina(n16234), .dinb(asqrt[62] ), .dout(n16235));
  jnot g15986(.din(n16235), .dout(n16236));
  jnot g15987(.din(n16228), .dout(n16237));
  jnot g15988(.din(n16220), .dout(n16238));
  jnot g15989(.din(n16213), .dout(n16239));
  jnot g15990(.din(n16205), .dout(n16240));
  jnot g15991(.din(n16198), .dout(n16241));
  jnot g15992(.din(n16190), .dout(n16242));
  jnot g15993(.din(n16182), .dout(n16243));
  jnot g15994(.din(n16174), .dout(n16244));
  jnot g15995(.din(n16167), .dout(n16245));
  jnot g15996(.din(n16159), .dout(n16246));
  jnot g15997(.din(n16152), .dout(n16247));
  jnot g15998(.din(n16144), .dout(n16248));
  jnot g15999(.din(n16137), .dout(n16249));
  jnot g16000(.din(n16140), .dout(n16250));
  jnot g16001(.din(n16130), .dout(n16251));
  jnot g16002(.din(n16122), .dout(n16252));
  jnot g16003(.din(n16114), .dout(n16253));
  jnot g16004(.din(n16107), .dout(n16254));
  jnot g16005(.din(n16099), .dout(n16255));
  jnot g16006(.din(n16092), .dout(n16256));
  jnot g16007(.din(n16084), .dout(n16257));
  jnot g16008(.din(n16076), .dout(n16258));
  jnot g16009(.din(n16068), .dout(n16259));
  jnot g16010(.din(n16061), .dout(n16260));
  jnot g16011(.din(n16053), .dout(n16261));
  jnot g16012(.din(n16046), .dout(n16262));
  jnot g16013(.din(n16038), .dout(n16263));
  jnot g16014(.din(n16030), .dout(n16264));
  jnot g16015(.din(n16022), .dout(n16265));
  jnot g16016(.din(n16015), .dout(n16266));
  jnot g16017(.din(n16007), .dout(n16267));
  jnot g16018(.din(n16000), .dout(n16268));
  jnot g16019(.din(n15992), .dout(n16269));
  jnot g16020(.din(n15985), .dout(n16270));
  jnot g16021(.din(n15977), .dout(n16271));
  jnot g16022(.din(n15970), .dout(n16272));
  jnot g16023(.din(n15962), .dout(n16273));
  jnot g16024(.din(n15954), .dout(n16274));
  jnot g16025(.din(n15946), .dout(n16275));
  jnot g16026(.din(n15939), .dout(n16276));
  jnot g16027(.din(n15931), .dout(n16277));
  jnot g16028(.din(n15924), .dout(n16278));
  jnot g16029(.din(n15916), .dout(n16279));
  jnot g16030(.din(n15909), .dout(n16280));
  jnot g16031(.din(n15902), .dout(n16281));
  jnot g16032(.din(n15895), .dout(n16282));
  jnot g16033(.din(n15883), .dout(n16283));
  jnot g16034(.din(n15647), .dout(n16284));
  jor  g16035(.dina(n15878), .dinb(n15265), .dout(n16285));
  jnot g16036(.din(n15645), .dout(n16286));
  jand g16037(.dina(n16286), .dinb(n16285), .dout(n16287));
  jand g16038(.dina(n16287), .dinb(n15260), .dout(n16288));
  jor  g16039(.dina(n15878), .dinb(a[28] ), .dout(n16289));
  jand g16040(.dina(n16289), .dinb(a[29] ), .dout(n16290));
  jor  g16041(.dina(n15885), .dinb(n16290), .dout(n16291));
  jor  g16042(.dina(n16291), .dinb(n16288), .dout(n16292));
  jand g16043(.dina(n16292), .dinb(n16284), .dout(n16293));
  jand g16044(.dina(n16293), .dinb(n14674), .dout(n16294));
  jor  g16045(.dina(n15891), .dinb(n16294), .dout(n16295));
  jand g16046(.dina(n16295), .dinb(n16283), .dout(n16296));
  jand g16047(.dina(n16296), .dinb(n14078), .dout(n16297));
  jnot g16048(.din(n15899), .dout(n16298));
  jor  g16049(.dina(n16298), .dinb(n16297), .dout(n16299));
  jand g16050(.dina(n16299), .dinb(n16282), .dout(n16300));
  jand g16051(.dina(n16300), .dinb(n13515), .dout(n16301));
  jnot g16052(.din(n15906), .dout(n16302));
  jor  g16053(.dina(n16302), .dinb(n16301), .dout(n16303));
  jand g16054(.dina(n16303), .dinb(n16281), .dout(n16304));
  jand g16055(.dina(n16304), .dinb(n12947), .dout(n16305));
  jnot g16056(.din(n15913), .dout(n16306));
  jor  g16057(.dina(n16306), .dinb(n16305), .dout(n16307));
  jand g16058(.dina(n16307), .dinb(n16280), .dout(n16308));
  jand g16059(.dina(n16308), .dinb(n12410), .dout(n16309));
  jor  g16060(.dina(n15920), .dinb(n16309), .dout(n16310));
  jand g16061(.dina(n16310), .dinb(n16279), .dout(n16311));
  jand g16062(.dina(n16311), .dinb(n11858), .dout(n16312));
  jnot g16063(.din(n15928), .dout(n16313));
  jor  g16064(.dina(n16313), .dinb(n16312), .dout(n16314));
  jand g16065(.dina(n16314), .dinb(n16278), .dout(n16315));
  jand g16066(.dina(n16315), .dinb(n11347), .dout(n16316));
  jor  g16067(.dina(n15935), .dinb(n16316), .dout(n16317));
  jand g16068(.dina(n16317), .dinb(n16277), .dout(n16318));
  jand g16069(.dina(n16318), .dinb(n10824), .dout(n16319));
  jnot g16070(.din(n15943), .dout(n16320));
  jor  g16071(.dina(n16320), .dinb(n16319), .dout(n16321));
  jand g16072(.dina(n16321), .dinb(n16276), .dout(n16322));
  jand g16073(.dina(n16322), .dinb(n10328), .dout(n16323));
  jor  g16074(.dina(n15950), .dinb(n16323), .dout(n16324));
  jand g16075(.dina(n16324), .dinb(n16275), .dout(n16325));
  jand g16076(.dina(n16325), .dinb(n9832), .dout(n16326));
  jor  g16077(.dina(n15958), .dinb(n16326), .dout(n16327));
  jand g16078(.dina(n16327), .dinb(n16274), .dout(n16328));
  jand g16079(.dina(n16328), .dinb(n9369), .dout(n16329));
  jor  g16080(.dina(n15966), .dinb(n16329), .dout(n16330));
  jand g16081(.dina(n16330), .dinb(n16273), .dout(n16331));
  jand g16082(.dina(n16331), .dinb(n8890), .dout(n16332));
  jnot g16083(.din(n15974), .dout(n16333));
  jor  g16084(.dina(n16333), .dinb(n16332), .dout(n16334));
  jand g16085(.dina(n16334), .dinb(n16272), .dout(n16335));
  jand g16086(.dina(n16335), .dinb(n8449), .dout(n16336));
  jor  g16087(.dina(n15981), .dinb(n16336), .dout(n16337));
  jand g16088(.dina(n16337), .dinb(n16271), .dout(n16338));
  jand g16089(.dina(n16338), .dinb(n8003), .dout(n16339));
  jnot g16090(.din(n15989), .dout(n16340));
  jor  g16091(.dina(n16340), .dinb(n16339), .dout(n16341));
  jand g16092(.dina(n16341), .dinb(n16270), .dout(n16342));
  jand g16093(.dina(n16342), .dinb(n7581), .dout(n16343));
  jor  g16094(.dina(n15996), .dinb(n16343), .dout(n16344));
  jand g16095(.dina(n16344), .dinb(n16269), .dout(n16345));
  jand g16096(.dina(n16345), .dinb(n7154), .dout(n16346));
  jnot g16097(.din(n16004), .dout(n16347));
  jor  g16098(.dina(n16347), .dinb(n16346), .dout(n16348));
  jand g16099(.dina(n16348), .dinb(n16268), .dout(n16349));
  jand g16100(.dina(n16349), .dinb(n6758), .dout(n16350));
  jor  g16101(.dina(n16011), .dinb(n16350), .dout(n16351));
  jand g16102(.dina(n16351), .dinb(n16267), .dout(n16352));
  jand g16103(.dina(n16352), .dinb(n6357), .dout(n16353));
  jnot g16104(.din(n16019), .dout(n16354));
  jor  g16105(.dina(n16354), .dinb(n16353), .dout(n16355));
  jand g16106(.dina(n16355), .dinb(n16266), .dout(n16356));
  jand g16107(.dina(n16356), .dinb(n5989), .dout(n16357));
  jor  g16108(.dina(n16026), .dinb(n16357), .dout(n16358));
  jand g16109(.dina(n16358), .dinb(n16265), .dout(n16359));
  jand g16110(.dina(n16359), .dinb(n5606), .dout(n16360));
  jor  g16111(.dina(n16034), .dinb(n16360), .dout(n16361));
  jand g16112(.dina(n16361), .dinb(n16264), .dout(n16362));
  jand g16113(.dina(n16362), .dinb(n5259), .dout(n16363));
  jor  g16114(.dina(n16042), .dinb(n16363), .dout(n16364));
  jand g16115(.dina(n16364), .dinb(n16263), .dout(n16365));
  jand g16116(.dina(n16365), .dinb(n4902), .dout(n16366));
  jnot g16117(.din(n16050), .dout(n16367));
  jor  g16118(.dina(n16367), .dinb(n16366), .dout(n16368));
  jand g16119(.dina(n16368), .dinb(n16262), .dout(n16369));
  jand g16120(.dina(n16369), .dinb(n4582), .dout(n16370));
  jor  g16121(.dina(n16057), .dinb(n16370), .dout(n16371));
  jand g16122(.dina(n16371), .dinb(n16261), .dout(n16372));
  jand g16123(.dina(n16372), .dinb(n4249), .dout(n16373));
  jnot g16124(.din(n16065), .dout(n16374));
  jor  g16125(.dina(n16374), .dinb(n16373), .dout(n16375));
  jand g16126(.dina(n16375), .dinb(n16260), .dout(n16376));
  jand g16127(.dina(n16376), .dinb(n3955), .dout(n16377));
  jor  g16128(.dina(n16072), .dinb(n16377), .dout(n16378));
  jand g16129(.dina(n16378), .dinb(n16259), .dout(n16379));
  jand g16130(.dina(n16379), .dinb(n3642), .dout(n16380));
  jor  g16131(.dina(n16080), .dinb(n16380), .dout(n16381));
  jand g16132(.dina(n16381), .dinb(n16258), .dout(n16382));
  jand g16133(.dina(n16382), .dinb(n3368), .dout(n16383));
  jor  g16134(.dina(n16088), .dinb(n16383), .dout(n16384));
  jand g16135(.dina(n16384), .dinb(n16257), .dout(n16385));
  jand g16136(.dina(n16385), .dinb(n3089), .dout(n16386));
  jnot g16137(.din(n16096), .dout(n16387));
  jor  g16138(.dina(n16387), .dinb(n16386), .dout(n16388));
  jand g16139(.dina(n16388), .dinb(n16256), .dout(n16389));
  jand g16140(.dina(n16389), .dinb(n2833), .dout(n16390));
  jor  g16141(.dina(n16103), .dinb(n16390), .dout(n16391));
  jand g16142(.dina(n16391), .dinb(n16255), .dout(n16392));
  jand g16143(.dina(n16392), .dinb(n2572), .dout(n16393));
  jnot g16144(.din(n16111), .dout(n16394));
  jor  g16145(.dina(n16394), .dinb(n16393), .dout(n16395));
  jand g16146(.dina(n16395), .dinb(n16254), .dout(n16396));
  jand g16147(.dina(n16396), .dinb(n2345), .dout(n16397));
  jor  g16148(.dina(n16118), .dinb(n16397), .dout(n16398));
  jand g16149(.dina(n16398), .dinb(n16253), .dout(n16399));
  jand g16150(.dina(n16399), .dinb(n2108), .dout(n16400));
  jor  g16151(.dina(n16126), .dinb(n16400), .dout(n16401));
  jand g16152(.dina(n16401), .dinb(n16252), .dout(n16402));
  jand g16153(.dina(n16402), .dinb(n1912), .dout(n16403));
  jnot g16154(.din(n16134), .dout(n16404));
  jor  g16155(.dina(n16404), .dinb(n16403), .dout(n16405));
  jand g16156(.dina(n16405), .dinb(n16251), .dout(n16406));
  jand g16157(.dina(n16406), .dinb(n1699), .dout(n16407));
  jor  g16158(.dina(n16407), .dinb(n16250), .dout(n16408));
  jand g16159(.dina(n16408), .dinb(n16249), .dout(n16409));
  jand g16160(.dina(n16409), .dinb(n1516), .dout(n16410));
  jor  g16161(.dina(n16148), .dinb(n16410), .dout(n16411));
  jand g16162(.dina(n16411), .dinb(n16248), .dout(n16412));
  jand g16163(.dina(n16412), .dinb(n1332), .dout(n16413));
  jnot g16164(.din(n16156), .dout(n16414));
  jor  g16165(.dina(n16414), .dinb(n16413), .dout(n16415));
  jand g16166(.dina(n16415), .dinb(n16247), .dout(n16416));
  jand g16167(.dina(n16416), .dinb(n1173), .dout(n16417));
  jor  g16168(.dina(n16163), .dinb(n16417), .dout(n16418));
  jand g16169(.dina(n16418), .dinb(n16246), .dout(n16419));
  jand g16170(.dina(n16419), .dinb(n1008), .dout(n16420));
  jnot g16171(.din(n16171), .dout(n16421));
  jor  g16172(.dina(n16421), .dinb(n16420), .dout(n16422));
  jand g16173(.dina(n16422), .dinb(n16245), .dout(n16423));
  jand g16174(.dina(n16423), .dinb(n884), .dout(n16424));
  jor  g16175(.dina(n16178), .dinb(n16424), .dout(n16425));
  jand g16176(.dina(n16425), .dinb(n16244), .dout(n16426));
  jand g16177(.dina(n16426), .dinb(n743), .dout(n16427));
  jor  g16178(.dina(n16186), .dinb(n16427), .dout(n16428));
  jand g16179(.dina(n16428), .dinb(n16243), .dout(n16429));
  jand g16180(.dina(n16429), .dinb(n635), .dout(n16430));
  jor  g16181(.dina(n16194), .dinb(n16430), .dout(n16431));
  jand g16182(.dina(n16431), .dinb(n16242), .dout(n16432));
  jand g16183(.dina(n16432), .dinb(n515), .dout(n16433));
  jnot g16184(.din(n16202), .dout(n16434));
  jor  g16185(.dina(n16434), .dinb(n16433), .dout(n16435));
  jand g16186(.dina(n16435), .dinb(n16241), .dout(n16436));
  jand g16187(.dina(n16436), .dinb(n443), .dout(n16437));
  jor  g16188(.dina(n16209), .dinb(n16437), .dout(n16438));
  jand g16189(.dina(n16438), .dinb(n16240), .dout(n16439));
  jand g16190(.dina(n16439), .dinb(n352), .dout(n16440));
  jnot g16191(.din(n16217), .dout(n16441));
  jor  g16192(.dina(n16441), .dinb(n16440), .dout(n16442));
  jand g16193(.dina(n16442), .dinb(n16239), .dout(n16443));
  jand g16194(.dina(n16443), .dinb(n294), .dout(n16444));
  jor  g16195(.dina(n16224), .dinb(n16444), .dout(n16445));
  jand g16196(.dina(n16445), .dinb(n16238), .dout(n16446));
  jand g16197(.dina(n16446), .dinb(n239), .dout(n16447));
  jnot g16198(.din(n16232), .dout(n16448));
  jor  g16199(.dina(n16448), .dinb(n16447), .dout(n16449));
  jand g16200(.dina(n16449), .dinb(n16237), .dout(n16450));
  jand g16201(.dina(n16450), .dinb(n221), .dout(n16451));
  jxor g16202(.dina(n15609), .dinb(n239), .dout(n16452));
  jand g16203(.dina(n16452), .dinb(asqrt[14] ), .dout(n16453));
  jxor g16204(.dina(n16453), .dinb(n15614), .dout(n16454));
  jor  g16205(.dina(n16454), .dinb(n16451), .dout(n16455));
  jand g16206(.dina(n16455), .dinb(n16236), .dout(n16456));
  jxor g16207(.dina(n15616), .dinb(n221), .dout(n16457));
  jand g16208(.dina(n16457), .dinb(asqrt[14] ), .dout(n16458));
  jxor g16209(.dina(n16458), .dinb(n15622), .dout(n16459));
  jor  g16210(.dina(n16459), .dinb(n16456), .dout(n16460));
  jand g16211(.dina(asqrt[14] ), .dinb(n15872), .dout(n16461));
  jor  g16212(.dina(n16461), .dinb(n15631), .dout(n16462));
  jor  g16213(.dina(n16462), .dinb(n16460), .dout(n16463));
  jand g16214(.dina(n16463), .dinb(n218), .dout(n16464));
  jand g16215(.dina(n15878), .dinb(n15264), .dout(n16465));
  jand g16216(.dina(n16459), .dinb(n16456), .dout(n16466));
  jor  g16217(.dina(n16466), .dinb(n16465), .dout(n16467));
  jand g16218(.dina(n15878), .dinb(n15624), .dout(n16468));
  jnot g16219(.din(n16468), .dout(n16469));
  jand g16220(.dina(n15625), .dinb(asqrt[63] ), .dout(n16470));
  jand g16221(.dina(n16470), .dinb(n15886), .dout(n16471));
  jand g16222(.dina(n16471), .dinb(n16469), .dout(n16472));
  jor  g16223(.dina(n16472), .dinb(n16467), .dout(n16473));
  jor  g16224(.dina(n16473), .dinb(n16464), .dout(asqrt[13] ));
  jor  g16225(.dina(n16234), .dinb(asqrt[62] ), .dout(n16475));
  jnot g16226(.din(n16454), .dout(n16476));
  jand g16227(.dina(n16476), .dinb(n16475), .dout(n16477));
  jor  g16228(.dina(n16477), .dinb(n16235), .dout(n16478));
  jnot g16229(.din(n16459), .dout(n16479));
  jand g16230(.dina(n16479), .dinb(n16478), .dout(n16480));
  jnot g16231(.din(n16462), .dout(n16481));
  jand g16232(.dina(n16481), .dinb(n16480), .dout(n16482));
  jor  g16233(.dina(n16482), .dinb(asqrt[63] ), .dout(n16483));
  jnot g16234(.din(n16465), .dout(n16484));
  jor  g16235(.dina(n16479), .dinb(n16478), .dout(n16485));
  jand g16236(.dina(n16485), .dinb(n16484), .dout(n16486));
  jnot g16237(.din(n16472), .dout(n16487));
  jand g16238(.dina(n16487), .dinb(n16486), .dout(n16488));
  jand g16239(.dina(n16488), .dinb(n16483), .dout(n16489));
  jxor g16240(.dina(n16234), .dinb(n221), .dout(n16490));
  jor  g16241(.dina(n16490), .dinb(n16489), .dout(n16491));
  jxor g16242(.dina(n16491), .dinb(n16454), .dout(n16492));
  jnot g16243(.din(n16492), .dout(n16493));
  jnot g16244(.din(a[24] ), .dout(n16494));
  jnot g16245(.din(a[25] ), .dout(n16495));
  jand g16246(.dina(n16495), .dinb(n16494), .dout(n16496));
  jand g16247(.dina(n16496), .dinb(n15642), .dout(n16497));
  jnot g16248(.din(n16497), .dout(n16498));
  jor  g16249(.dina(n16489), .dinb(n15642), .dout(n16499));
  jand g16250(.dina(n16499), .dinb(n16498), .dout(n16500));
  jor  g16251(.dina(n16500), .dinb(n15878), .dout(n16501));
  jand g16252(.dina(n16500), .dinb(n15878), .dout(n16502));
  jor  g16253(.dina(n16489), .dinb(a[26] ), .dout(n16503));
  jand g16254(.dina(n16503), .dinb(a[27] ), .dout(n16504));
  jand g16255(.dina(asqrt[13] ), .dinb(n15644), .dout(n16505));
  jor  g16256(.dina(n16505), .dinb(n16504), .dout(n16506));
  jor  g16257(.dina(n16506), .dinb(n16502), .dout(n16507));
  jand g16258(.dina(n16507), .dinb(n16501), .dout(n16508));
  jor  g16259(.dina(n16508), .dinb(n15260), .dout(n16509));
  jand g16260(.dina(n16508), .dinb(n15260), .dout(n16510));
  jnot g16261(.din(n15644), .dout(n16511));
  jor  g16262(.dina(n16489), .dinb(n16511), .dout(n16512));
  jor  g16263(.dina(n16471), .dinb(n15878), .dout(n16513));
  jor  g16264(.dina(n16513), .dinb(n16464), .dout(n16514));
  jor  g16265(.dina(n16514), .dinb(n16466), .dout(n16515));
  jand g16266(.dina(n16515), .dinb(n16512), .dout(n16516));
  jxor g16267(.dina(n16516), .dinb(n15265), .dout(n16517));
  jor  g16268(.dina(n16517), .dinb(n16510), .dout(n16518));
  jand g16269(.dina(n16518), .dinb(n16509), .dout(n16519));
  jor  g16270(.dina(n16519), .dinb(n14674), .dout(n16520));
  jand g16271(.dina(n16519), .dinb(n14674), .dout(n16521));
  jxor g16272(.dina(n15646), .dinb(n15260), .dout(n16522));
  jor  g16273(.dina(n16522), .dinb(n16489), .dout(n16523));
  jxor g16274(.dina(n16523), .dinb(n16291), .dout(n16524));
  jnot g16275(.din(n16524), .dout(n16525));
  jor  g16276(.dina(n16525), .dinb(n16521), .dout(n16526));
  jand g16277(.dina(n16526), .dinb(n16520), .dout(n16527));
  jor  g16278(.dina(n16527), .dinb(n14078), .dout(n16528));
  jand g16279(.dina(n16527), .dinb(n14078), .dout(n16529));
  jxor g16280(.dina(n15882), .dinb(n14674), .dout(n16530));
  jor  g16281(.dina(n16530), .dinb(n16489), .dout(n16531));
  jxor g16282(.dina(n16531), .dinb(n15892), .dout(n16532));
  jor  g16283(.dina(n16532), .dinb(n16529), .dout(n16533));
  jand g16284(.dina(n16533), .dinb(n16528), .dout(n16534));
  jor  g16285(.dina(n16534), .dinb(n13515), .dout(n16535));
  jand g16286(.dina(n16534), .dinb(n13515), .dout(n16536));
  jxor g16287(.dina(n15894), .dinb(n14078), .dout(n16537));
  jor  g16288(.dina(n16537), .dinb(n16489), .dout(n16538));
  jxor g16289(.dina(n16538), .dinb(n15899), .dout(n16539));
  jor  g16290(.dina(n16539), .dinb(n16536), .dout(n16540));
  jand g16291(.dina(n16540), .dinb(n16535), .dout(n16541));
  jor  g16292(.dina(n16541), .dinb(n12947), .dout(n16542));
  jand g16293(.dina(n16541), .dinb(n12947), .dout(n16543));
  jxor g16294(.dina(n15901), .dinb(n13515), .dout(n16544));
  jor  g16295(.dina(n16544), .dinb(n16489), .dout(n16545));
  jxor g16296(.dina(n16545), .dinb(n16302), .dout(n16546));
  jnot g16297(.din(n16546), .dout(n16547));
  jor  g16298(.dina(n16547), .dinb(n16543), .dout(n16548));
  jand g16299(.dina(n16548), .dinb(n16542), .dout(n16549));
  jor  g16300(.dina(n16549), .dinb(n12410), .dout(n16550));
  jand g16301(.dina(n16549), .dinb(n12410), .dout(n16551));
  jxor g16302(.dina(n15908), .dinb(n12947), .dout(n16552));
  jor  g16303(.dina(n16552), .dinb(n16489), .dout(n16553));
  jxor g16304(.dina(n16553), .dinb(n16306), .dout(n16554));
  jnot g16305(.din(n16554), .dout(n16555));
  jor  g16306(.dina(n16555), .dinb(n16551), .dout(n16556));
  jand g16307(.dina(n16556), .dinb(n16550), .dout(n16557));
  jor  g16308(.dina(n16557), .dinb(n11858), .dout(n16558));
  jand g16309(.dina(n16557), .dinb(n11858), .dout(n16559));
  jxor g16310(.dina(n15915), .dinb(n12410), .dout(n16560));
  jor  g16311(.dina(n16560), .dinb(n16489), .dout(n16561));
  jxor g16312(.dina(n16561), .dinb(n15921), .dout(n16562));
  jor  g16313(.dina(n16562), .dinb(n16559), .dout(n16563));
  jand g16314(.dina(n16563), .dinb(n16558), .dout(n16564));
  jor  g16315(.dina(n16564), .dinb(n11347), .dout(n16565));
  jand g16316(.dina(n16564), .dinb(n11347), .dout(n16566));
  jxor g16317(.dina(n15923), .dinb(n11858), .dout(n16567));
  jor  g16318(.dina(n16567), .dinb(n16489), .dout(n16568));
  jxor g16319(.dina(n16568), .dinb(n16313), .dout(n16569));
  jnot g16320(.din(n16569), .dout(n16570));
  jor  g16321(.dina(n16570), .dinb(n16566), .dout(n16571));
  jand g16322(.dina(n16571), .dinb(n16565), .dout(n16572));
  jor  g16323(.dina(n16572), .dinb(n10824), .dout(n16573));
  jand g16324(.dina(n16572), .dinb(n10824), .dout(n16574));
  jxor g16325(.dina(n15930), .dinb(n11347), .dout(n16575));
  jor  g16326(.dina(n16575), .dinb(n16489), .dout(n16576));
  jxor g16327(.dina(n16576), .dinb(n15936), .dout(n16577));
  jor  g16328(.dina(n16577), .dinb(n16574), .dout(n16578));
  jand g16329(.dina(n16578), .dinb(n16573), .dout(n16579));
  jor  g16330(.dina(n16579), .dinb(n10328), .dout(n16580));
  jand g16331(.dina(n16579), .dinb(n10328), .dout(n16581));
  jxor g16332(.dina(n15938), .dinb(n10824), .dout(n16582));
  jor  g16333(.dina(n16582), .dinb(n16489), .dout(n16583));
  jxor g16334(.dina(n16583), .dinb(n16320), .dout(n16584));
  jnot g16335(.din(n16584), .dout(n16585));
  jor  g16336(.dina(n16585), .dinb(n16581), .dout(n16586));
  jand g16337(.dina(n16586), .dinb(n16580), .dout(n16587));
  jor  g16338(.dina(n16587), .dinb(n9832), .dout(n16588));
  jand g16339(.dina(n16587), .dinb(n9832), .dout(n16589));
  jxor g16340(.dina(n15945), .dinb(n10328), .dout(n16590));
  jor  g16341(.dina(n16590), .dinb(n16489), .dout(n16591));
  jxor g16342(.dina(n16591), .dinb(n15951), .dout(n16592));
  jor  g16343(.dina(n16592), .dinb(n16589), .dout(n16593));
  jand g16344(.dina(n16593), .dinb(n16588), .dout(n16594));
  jor  g16345(.dina(n16594), .dinb(n9369), .dout(n16595));
  jand g16346(.dina(n16594), .dinb(n9369), .dout(n16596));
  jxor g16347(.dina(n15953), .dinb(n9832), .dout(n16597));
  jor  g16348(.dina(n16597), .dinb(n16489), .dout(n16598));
  jxor g16349(.dina(n16598), .dinb(n15959), .dout(n16599));
  jor  g16350(.dina(n16599), .dinb(n16596), .dout(n16600));
  jand g16351(.dina(n16600), .dinb(n16595), .dout(n16601));
  jor  g16352(.dina(n16601), .dinb(n8890), .dout(n16602));
  jand g16353(.dina(n16601), .dinb(n8890), .dout(n16603));
  jxor g16354(.dina(n15961), .dinb(n9369), .dout(n16604));
  jor  g16355(.dina(n16604), .dinb(n16489), .dout(n16605));
  jxor g16356(.dina(n16605), .dinb(n15967), .dout(n16606));
  jor  g16357(.dina(n16606), .dinb(n16603), .dout(n16607));
  jand g16358(.dina(n16607), .dinb(n16602), .dout(n16608));
  jor  g16359(.dina(n16608), .dinb(n8449), .dout(n16609));
  jand g16360(.dina(n16608), .dinb(n8449), .dout(n16610));
  jxor g16361(.dina(n15969), .dinb(n8890), .dout(n16611));
  jor  g16362(.dina(n16611), .dinb(n16489), .dout(n16612));
  jxor g16363(.dina(n16612), .dinb(n16333), .dout(n16613));
  jnot g16364(.din(n16613), .dout(n16614));
  jor  g16365(.dina(n16614), .dinb(n16610), .dout(n16615));
  jand g16366(.dina(n16615), .dinb(n16609), .dout(n16616));
  jor  g16367(.dina(n16616), .dinb(n8003), .dout(n16617));
  jand g16368(.dina(n16616), .dinb(n8003), .dout(n16618));
  jxor g16369(.dina(n15976), .dinb(n8449), .dout(n16619));
  jor  g16370(.dina(n16619), .dinb(n16489), .dout(n16620));
  jxor g16371(.dina(n16620), .dinb(n15982), .dout(n16621));
  jor  g16372(.dina(n16621), .dinb(n16618), .dout(n16622));
  jand g16373(.dina(n16622), .dinb(n16617), .dout(n16623));
  jor  g16374(.dina(n16623), .dinb(n7581), .dout(n16624));
  jand g16375(.dina(n16623), .dinb(n7581), .dout(n16625));
  jxor g16376(.dina(n15984), .dinb(n8003), .dout(n16626));
  jor  g16377(.dina(n16626), .dinb(n16489), .dout(n16627));
  jxor g16378(.dina(n16627), .dinb(n16340), .dout(n16628));
  jnot g16379(.din(n16628), .dout(n16629));
  jor  g16380(.dina(n16629), .dinb(n16625), .dout(n16630));
  jand g16381(.dina(n16630), .dinb(n16624), .dout(n16631));
  jor  g16382(.dina(n16631), .dinb(n7154), .dout(n16632));
  jand g16383(.dina(n16631), .dinb(n7154), .dout(n16633));
  jxor g16384(.dina(n15991), .dinb(n7581), .dout(n16634));
  jor  g16385(.dina(n16634), .dinb(n16489), .dout(n16635));
  jxor g16386(.dina(n16635), .dinb(n15997), .dout(n16636));
  jor  g16387(.dina(n16636), .dinb(n16633), .dout(n16637));
  jand g16388(.dina(n16637), .dinb(n16632), .dout(n16638));
  jor  g16389(.dina(n16638), .dinb(n6758), .dout(n16639));
  jand g16390(.dina(n16638), .dinb(n6758), .dout(n16640));
  jxor g16391(.dina(n15999), .dinb(n7154), .dout(n16641));
  jor  g16392(.dina(n16641), .dinb(n16489), .dout(n16642));
  jxor g16393(.dina(n16642), .dinb(n16347), .dout(n16643));
  jnot g16394(.din(n16643), .dout(n16644));
  jor  g16395(.dina(n16644), .dinb(n16640), .dout(n16645));
  jand g16396(.dina(n16645), .dinb(n16639), .dout(n16646));
  jor  g16397(.dina(n16646), .dinb(n6357), .dout(n16647));
  jand g16398(.dina(n16646), .dinb(n6357), .dout(n16648));
  jxor g16399(.dina(n16006), .dinb(n6758), .dout(n16649));
  jor  g16400(.dina(n16649), .dinb(n16489), .dout(n16650));
  jxor g16401(.dina(n16650), .dinb(n16012), .dout(n16651));
  jor  g16402(.dina(n16651), .dinb(n16648), .dout(n16652));
  jand g16403(.dina(n16652), .dinb(n16647), .dout(n16653));
  jor  g16404(.dina(n16653), .dinb(n5989), .dout(n16654));
  jand g16405(.dina(n16653), .dinb(n5989), .dout(n16655));
  jxor g16406(.dina(n16014), .dinb(n6357), .dout(n16656));
  jor  g16407(.dina(n16656), .dinb(n16489), .dout(n16657));
  jxor g16408(.dina(n16657), .dinb(n16354), .dout(n16658));
  jnot g16409(.din(n16658), .dout(n16659));
  jor  g16410(.dina(n16659), .dinb(n16655), .dout(n16660));
  jand g16411(.dina(n16660), .dinb(n16654), .dout(n16661));
  jor  g16412(.dina(n16661), .dinb(n5606), .dout(n16662));
  jand g16413(.dina(n16661), .dinb(n5606), .dout(n16663));
  jxor g16414(.dina(n16021), .dinb(n5989), .dout(n16664));
  jor  g16415(.dina(n16664), .dinb(n16489), .dout(n16665));
  jxor g16416(.dina(n16665), .dinb(n16027), .dout(n16666));
  jor  g16417(.dina(n16666), .dinb(n16663), .dout(n16667));
  jand g16418(.dina(n16667), .dinb(n16662), .dout(n16668));
  jor  g16419(.dina(n16668), .dinb(n5259), .dout(n16669));
  jand g16420(.dina(n16668), .dinb(n5259), .dout(n16670));
  jxor g16421(.dina(n16029), .dinb(n5606), .dout(n16671));
  jor  g16422(.dina(n16671), .dinb(n16489), .dout(n16672));
  jxor g16423(.dina(n16672), .dinb(n16035), .dout(n16673));
  jor  g16424(.dina(n16673), .dinb(n16670), .dout(n16674));
  jand g16425(.dina(n16674), .dinb(n16669), .dout(n16675));
  jor  g16426(.dina(n16675), .dinb(n4902), .dout(n16676));
  jand g16427(.dina(n16675), .dinb(n4902), .dout(n16677));
  jxor g16428(.dina(n16037), .dinb(n5259), .dout(n16678));
  jor  g16429(.dina(n16678), .dinb(n16489), .dout(n16679));
  jxor g16430(.dina(n16679), .dinb(n16043), .dout(n16680));
  jor  g16431(.dina(n16680), .dinb(n16677), .dout(n16681));
  jand g16432(.dina(n16681), .dinb(n16676), .dout(n16682));
  jor  g16433(.dina(n16682), .dinb(n4582), .dout(n16683));
  jand g16434(.dina(n16682), .dinb(n4582), .dout(n16684));
  jxor g16435(.dina(n16045), .dinb(n4902), .dout(n16685));
  jor  g16436(.dina(n16685), .dinb(n16489), .dout(n16686));
  jxor g16437(.dina(n16686), .dinb(n16367), .dout(n16687));
  jnot g16438(.din(n16687), .dout(n16688));
  jor  g16439(.dina(n16688), .dinb(n16684), .dout(n16689));
  jand g16440(.dina(n16689), .dinb(n16683), .dout(n16690));
  jor  g16441(.dina(n16690), .dinb(n4249), .dout(n16691));
  jand g16442(.dina(n16690), .dinb(n4249), .dout(n16692));
  jxor g16443(.dina(n16052), .dinb(n4582), .dout(n16693));
  jor  g16444(.dina(n16693), .dinb(n16489), .dout(n16694));
  jxor g16445(.dina(n16694), .dinb(n16058), .dout(n16695));
  jor  g16446(.dina(n16695), .dinb(n16692), .dout(n16696));
  jand g16447(.dina(n16696), .dinb(n16691), .dout(n16697));
  jor  g16448(.dina(n16697), .dinb(n3955), .dout(n16698));
  jand g16449(.dina(n16697), .dinb(n3955), .dout(n16699));
  jxor g16450(.dina(n16060), .dinb(n4249), .dout(n16700));
  jor  g16451(.dina(n16700), .dinb(n16489), .dout(n16701));
  jxor g16452(.dina(n16701), .dinb(n16374), .dout(n16702));
  jnot g16453(.din(n16702), .dout(n16703));
  jor  g16454(.dina(n16703), .dinb(n16699), .dout(n16704));
  jand g16455(.dina(n16704), .dinb(n16698), .dout(n16705));
  jor  g16456(.dina(n16705), .dinb(n3642), .dout(n16706));
  jand g16457(.dina(n16705), .dinb(n3642), .dout(n16707));
  jxor g16458(.dina(n16067), .dinb(n3955), .dout(n16708));
  jor  g16459(.dina(n16708), .dinb(n16489), .dout(n16709));
  jxor g16460(.dina(n16709), .dinb(n16073), .dout(n16710));
  jor  g16461(.dina(n16710), .dinb(n16707), .dout(n16711));
  jand g16462(.dina(n16711), .dinb(n16706), .dout(n16712));
  jor  g16463(.dina(n16712), .dinb(n3368), .dout(n16713));
  jand g16464(.dina(n16712), .dinb(n3368), .dout(n16714));
  jxor g16465(.dina(n16075), .dinb(n3642), .dout(n16715));
  jor  g16466(.dina(n16715), .dinb(n16489), .dout(n16716));
  jxor g16467(.dina(n16716), .dinb(n16081), .dout(n16717));
  jor  g16468(.dina(n16717), .dinb(n16714), .dout(n16718));
  jand g16469(.dina(n16718), .dinb(n16713), .dout(n16719));
  jor  g16470(.dina(n16719), .dinb(n3089), .dout(n16720));
  jand g16471(.dina(n16719), .dinb(n3089), .dout(n16721));
  jxor g16472(.dina(n16083), .dinb(n3368), .dout(n16722));
  jor  g16473(.dina(n16722), .dinb(n16489), .dout(n16723));
  jxor g16474(.dina(n16723), .dinb(n16089), .dout(n16724));
  jor  g16475(.dina(n16724), .dinb(n16721), .dout(n16725));
  jand g16476(.dina(n16725), .dinb(n16720), .dout(n16726));
  jor  g16477(.dina(n16726), .dinb(n2833), .dout(n16727));
  jand g16478(.dina(n16726), .dinb(n2833), .dout(n16728));
  jxor g16479(.dina(n16091), .dinb(n3089), .dout(n16729));
  jor  g16480(.dina(n16729), .dinb(n16489), .dout(n16730));
  jxor g16481(.dina(n16730), .dinb(n16387), .dout(n16731));
  jnot g16482(.din(n16731), .dout(n16732));
  jor  g16483(.dina(n16732), .dinb(n16728), .dout(n16733));
  jand g16484(.dina(n16733), .dinb(n16727), .dout(n16734));
  jor  g16485(.dina(n16734), .dinb(n2572), .dout(n16735));
  jand g16486(.dina(n16734), .dinb(n2572), .dout(n16736));
  jxor g16487(.dina(n16098), .dinb(n2833), .dout(n16737));
  jor  g16488(.dina(n16737), .dinb(n16489), .dout(n16738));
  jxor g16489(.dina(n16738), .dinb(n16104), .dout(n16739));
  jor  g16490(.dina(n16739), .dinb(n16736), .dout(n16740));
  jand g16491(.dina(n16740), .dinb(n16735), .dout(n16741));
  jor  g16492(.dina(n16741), .dinb(n2345), .dout(n16742));
  jand g16493(.dina(n16741), .dinb(n2345), .dout(n16743));
  jxor g16494(.dina(n16106), .dinb(n2572), .dout(n16744));
  jor  g16495(.dina(n16744), .dinb(n16489), .dout(n16745));
  jxor g16496(.dina(n16745), .dinb(n16394), .dout(n16746));
  jnot g16497(.din(n16746), .dout(n16747));
  jor  g16498(.dina(n16747), .dinb(n16743), .dout(n16748));
  jand g16499(.dina(n16748), .dinb(n16742), .dout(n16749));
  jor  g16500(.dina(n16749), .dinb(n2108), .dout(n16750));
  jand g16501(.dina(n16749), .dinb(n2108), .dout(n16751));
  jxor g16502(.dina(n16113), .dinb(n2345), .dout(n16752));
  jor  g16503(.dina(n16752), .dinb(n16489), .dout(n16753));
  jxor g16504(.dina(n16753), .dinb(n16119), .dout(n16754));
  jor  g16505(.dina(n16754), .dinb(n16751), .dout(n16755));
  jand g16506(.dina(n16755), .dinb(n16750), .dout(n16756));
  jor  g16507(.dina(n16756), .dinb(n1912), .dout(n16757));
  jand g16508(.dina(n16756), .dinb(n1912), .dout(n16758));
  jxor g16509(.dina(n16121), .dinb(n2108), .dout(n16759));
  jor  g16510(.dina(n16759), .dinb(n16489), .dout(n16760));
  jxor g16511(.dina(n16760), .dinb(n16127), .dout(n16761));
  jor  g16512(.dina(n16761), .dinb(n16758), .dout(n16762));
  jand g16513(.dina(n16762), .dinb(n16757), .dout(n16763));
  jor  g16514(.dina(n16763), .dinb(n1699), .dout(n16764));
  jand g16515(.dina(n16763), .dinb(n1699), .dout(n16765));
  jxor g16516(.dina(n16129), .dinb(n1912), .dout(n16766));
  jor  g16517(.dina(n16766), .dinb(n16489), .dout(n16767));
  jxor g16518(.dina(n16767), .dinb(n16404), .dout(n16768));
  jnot g16519(.din(n16768), .dout(n16769));
  jor  g16520(.dina(n16769), .dinb(n16765), .dout(n16770));
  jand g16521(.dina(n16770), .dinb(n16764), .dout(n16771));
  jor  g16522(.dina(n16771), .dinb(n1516), .dout(n16772));
  jxor g16523(.dina(n16136), .dinb(n1699), .dout(n16773));
  jor  g16524(.dina(n16773), .dinb(n16489), .dout(n16774));
  jxor g16525(.dina(n16774), .dinb(n16250), .dout(n16775));
  jnot g16526(.din(n16775), .dout(n16776));
  jand g16527(.dina(n16771), .dinb(n1516), .dout(n16777));
  jor  g16528(.dina(n16777), .dinb(n16776), .dout(n16778));
  jand g16529(.dina(n16778), .dinb(n16772), .dout(n16779));
  jor  g16530(.dina(n16779), .dinb(n1332), .dout(n16780));
  jand g16531(.dina(n16779), .dinb(n1332), .dout(n16781));
  jxor g16532(.dina(n16143), .dinb(n1516), .dout(n16782));
  jor  g16533(.dina(n16782), .dinb(n16489), .dout(n16783));
  jxor g16534(.dina(n16783), .dinb(n16149), .dout(n16784));
  jor  g16535(.dina(n16784), .dinb(n16781), .dout(n16785));
  jand g16536(.dina(n16785), .dinb(n16780), .dout(n16786));
  jor  g16537(.dina(n16786), .dinb(n1173), .dout(n16787));
  jand g16538(.dina(n16786), .dinb(n1173), .dout(n16788));
  jxor g16539(.dina(n16151), .dinb(n1332), .dout(n16789));
  jor  g16540(.dina(n16789), .dinb(n16489), .dout(n16790));
  jxor g16541(.dina(n16790), .dinb(n16414), .dout(n16791));
  jnot g16542(.din(n16791), .dout(n16792));
  jor  g16543(.dina(n16792), .dinb(n16788), .dout(n16793));
  jand g16544(.dina(n16793), .dinb(n16787), .dout(n16794));
  jor  g16545(.dina(n16794), .dinb(n1008), .dout(n16795));
  jand g16546(.dina(n16794), .dinb(n1008), .dout(n16796));
  jxor g16547(.dina(n16158), .dinb(n1173), .dout(n16797));
  jor  g16548(.dina(n16797), .dinb(n16489), .dout(n16798));
  jxor g16549(.dina(n16798), .dinb(n16164), .dout(n16799));
  jor  g16550(.dina(n16799), .dinb(n16796), .dout(n16800));
  jand g16551(.dina(n16800), .dinb(n16795), .dout(n16801));
  jor  g16552(.dina(n16801), .dinb(n884), .dout(n16802));
  jand g16553(.dina(n16801), .dinb(n884), .dout(n16803));
  jxor g16554(.dina(n16166), .dinb(n1008), .dout(n16804));
  jor  g16555(.dina(n16804), .dinb(n16489), .dout(n16805));
  jxor g16556(.dina(n16805), .dinb(n16421), .dout(n16806));
  jnot g16557(.din(n16806), .dout(n16807));
  jor  g16558(.dina(n16807), .dinb(n16803), .dout(n16808));
  jand g16559(.dina(n16808), .dinb(n16802), .dout(n16809));
  jor  g16560(.dina(n16809), .dinb(n743), .dout(n16810));
  jand g16561(.dina(n16809), .dinb(n743), .dout(n16811));
  jxor g16562(.dina(n16173), .dinb(n884), .dout(n16812));
  jor  g16563(.dina(n16812), .dinb(n16489), .dout(n16813));
  jxor g16564(.dina(n16813), .dinb(n16179), .dout(n16814));
  jor  g16565(.dina(n16814), .dinb(n16811), .dout(n16815));
  jand g16566(.dina(n16815), .dinb(n16810), .dout(n16816));
  jor  g16567(.dina(n16816), .dinb(n635), .dout(n16817));
  jand g16568(.dina(n16816), .dinb(n635), .dout(n16818));
  jxor g16569(.dina(n16181), .dinb(n743), .dout(n16819));
  jor  g16570(.dina(n16819), .dinb(n16489), .dout(n16820));
  jxor g16571(.dina(n16820), .dinb(n16187), .dout(n16821));
  jor  g16572(.dina(n16821), .dinb(n16818), .dout(n16822));
  jand g16573(.dina(n16822), .dinb(n16817), .dout(n16823));
  jor  g16574(.dina(n16823), .dinb(n515), .dout(n16824));
  jand g16575(.dina(n16823), .dinb(n515), .dout(n16825));
  jxor g16576(.dina(n16189), .dinb(n635), .dout(n16826));
  jor  g16577(.dina(n16826), .dinb(n16489), .dout(n16827));
  jxor g16578(.dina(n16827), .dinb(n16195), .dout(n16828));
  jor  g16579(.dina(n16828), .dinb(n16825), .dout(n16829));
  jand g16580(.dina(n16829), .dinb(n16824), .dout(n16830));
  jor  g16581(.dina(n16830), .dinb(n443), .dout(n16831));
  jand g16582(.dina(n16830), .dinb(n443), .dout(n16832));
  jxor g16583(.dina(n16197), .dinb(n515), .dout(n16833));
  jor  g16584(.dina(n16833), .dinb(n16489), .dout(n16834));
  jxor g16585(.dina(n16834), .dinb(n16434), .dout(n16835));
  jnot g16586(.din(n16835), .dout(n16836));
  jor  g16587(.dina(n16836), .dinb(n16832), .dout(n16837));
  jand g16588(.dina(n16837), .dinb(n16831), .dout(n16838));
  jor  g16589(.dina(n16838), .dinb(n352), .dout(n16839));
  jand g16590(.dina(n16838), .dinb(n352), .dout(n16840));
  jxor g16591(.dina(n16204), .dinb(n443), .dout(n16841));
  jor  g16592(.dina(n16841), .dinb(n16489), .dout(n16842));
  jxor g16593(.dina(n16842), .dinb(n16210), .dout(n16843));
  jor  g16594(.dina(n16843), .dinb(n16840), .dout(n16844));
  jand g16595(.dina(n16844), .dinb(n16839), .dout(n16845));
  jor  g16596(.dina(n16845), .dinb(n294), .dout(n16846));
  jand g16597(.dina(n16845), .dinb(n294), .dout(n16847));
  jxor g16598(.dina(n16212), .dinb(n352), .dout(n16848));
  jor  g16599(.dina(n16848), .dinb(n16489), .dout(n16849));
  jxor g16600(.dina(n16849), .dinb(n16441), .dout(n16850));
  jnot g16601(.din(n16850), .dout(n16851));
  jor  g16602(.dina(n16851), .dinb(n16847), .dout(n16852));
  jand g16603(.dina(n16852), .dinb(n16846), .dout(n16853));
  jor  g16604(.dina(n16853), .dinb(n239), .dout(n16854));
  jand g16605(.dina(n16853), .dinb(n239), .dout(n16855));
  jxor g16606(.dina(n16219), .dinb(n294), .dout(n16856));
  jor  g16607(.dina(n16856), .dinb(n16489), .dout(n16857));
  jxor g16608(.dina(n16857), .dinb(n16225), .dout(n16858));
  jor  g16609(.dina(n16858), .dinb(n16855), .dout(n16859));
  jand g16610(.dina(n16859), .dinb(n16854), .dout(n16860));
  jor  g16611(.dina(n16860), .dinb(n221), .dout(n16861));
  jand g16612(.dina(n16860), .dinb(n221), .dout(n16862));
  jxor g16613(.dina(n16227), .dinb(n239), .dout(n16863));
  jor  g16614(.dina(n16863), .dinb(n16489), .dout(n16864));
  jxor g16615(.dina(n16864), .dinb(n16448), .dout(n16865));
  jnot g16616(.din(n16865), .dout(n16866));
  jor  g16617(.dina(n16866), .dinb(n16862), .dout(n16867));
  jand g16618(.dina(n16867), .dinb(n16861), .dout(n16868));
  jand g16619(.dina(n16868), .dinb(n16493), .dout(n16869));
  jor  g16620(.dina(n16868), .dinb(n16493), .dout(n16871));
  jand g16621(.dina(asqrt[13] ), .dinb(n16480), .dout(n16872));
  jor  g16622(.dina(n16872), .dinb(n16871), .dout(n16873));
  jor  g16623(.dina(n16873), .dinb(n16466), .dout(n16874));
  jand g16624(.dina(n16874), .dinb(n218), .dout(n16875));
  jand g16625(.dina(n16489), .dinb(n16456), .dout(n16876));
  jand g16626(.dina(n16460), .dinb(asqrt[63] ), .dout(n16877));
  jand g16627(.dina(n16877), .dinb(n16485), .dout(n16878));
  jnot g16628(.din(n16878), .dout(n16879));
  jor  g16629(.dina(n16879), .dinb(n16876), .dout(n16880));
  jnot g16630(.din(n16880), .dout(n16881));
  jor  g16631(.dina(n16881), .dinb(n16875), .dout(n16882));
  jor  g16632(.dina(n16882), .dinb(n16869), .dout(asqrt[12] ));
  jnot g16633(.din(a[22] ), .dout(n16885));
  jnot g16634(.din(a[23] ), .dout(n16886));
  jand g16635(.dina(n16886), .dinb(n16885), .dout(n16887));
  jand g16636(.dina(n16887), .dinb(n16494), .dout(n16888));
  jand g16637(.dina(asqrt[12] ), .dinb(a[24] ), .dout(n16889));
  jor  g16638(.dina(n16889), .dinb(n16888), .dout(n16890));
  jand g16639(.dina(n16890), .dinb(asqrt[13] ), .dout(n16891));
  jor  g16640(.dina(n16890), .dinb(asqrt[13] ), .dout(n16892));
  jand g16641(.dina(asqrt[12] ), .dinb(n16494), .dout(n16893));
  jor  g16642(.dina(n16893), .dinb(n16495), .dout(n16894));
  jnot g16643(.din(n16496), .dout(n16895));
  jnot g16644(.din(n16869), .dout(n16896));
  jnot g16645(.din(n16861), .dout(n16898));
  jnot g16646(.din(n16854), .dout(n16899));
  jnot g16647(.din(n16846), .dout(n16900));
  jnot g16648(.din(n16839), .dout(n16901));
  jnot g16649(.din(n16831), .dout(n16902));
  jnot g16650(.din(n16824), .dout(n16903));
  jnot g16651(.din(n16817), .dout(n16904));
  jnot g16652(.din(n16810), .dout(n16905));
  jnot g16653(.din(n16802), .dout(n16906));
  jnot g16654(.din(n16795), .dout(n16907));
  jnot g16655(.din(n16787), .dout(n16908));
  jnot g16656(.din(n16780), .dout(n16909));
  jnot g16657(.din(n16772), .dout(n16910));
  jnot g16658(.din(n16764), .dout(n16911));
  jnot g16659(.din(n16757), .dout(n16912));
  jnot g16660(.din(n16750), .dout(n16913));
  jnot g16661(.din(n16742), .dout(n16914));
  jnot g16662(.din(n16735), .dout(n16915));
  jnot g16663(.din(n16727), .dout(n16916));
  jnot g16664(.din(n16720), .dout(n16917));
  jnot g16665(.din(n16713), .dout(n16918));
  jnot g16666(.din(n16706), .dout(n16919));
  jnot g16667(.din(n16698), .dout(n16920));
  jnot g16668(.din(n16691), .dout(n16921));
  jnot g16669(.din(n16683), .dout(n16922));
  jnot g16670(.din(n16676), .dout(n16923));
  jnot g16671(.din(n16669), .dout(n16924));
  jnot g16672(.din(n16662), .dout(n16925));
  jnot g16673(.din(n16654), .dout(n16926));
  jnot g16674(.din(n16647), .dout(n16927));
  jnot g16675(.din(n16639), .dout(n16928));
  jnot g16676(.din(n16632), .dout(n16929));
  jnot g16677(.din(n16624), .dout(n16930));
  jnot g16678(.din(n16617), .dout(n16931));
  jnot g16679(.din(n16609), .dout(n16932));
  jnot g16680(.din(n16602), .dout(n16933));
  jnot g16681(.din(n16595), .dout(n16934));
  jnot g16682(.din(n16588), .dout(n16935));
  jnot g16683(.din(n16580), .dout(n16936));
  jnot g16684(.din(n16573), .dout(n16937));
  jnot g16685(.din(n16565), .dout(n16938));
  jnot g16686(.din(n16558), .dout(n16939));
  jnot g16687(.din(n16550), .dout(n16940));
  jnot g16688(.din(n16542), .dout(n16941));
  jnot g16689(.din(n16535), .dout(n16942));
  jnot g16690(.din(n16528), .dout(n16943));
  jnot g16691(.din(n16520), .dout(n16944));
  jnot g16692(.din(n16509), .dout(n16945));
  jnot g16693(.din(n16501), .dout(n16946));
  jand g16694(.dina(asqrt[13] ), .dinb(a[26] ), .dout(n16947));
  jor  g16695(.dina(n16947), .dinb(n16497), .dout(n16948));
  jor  g16696(.dina(n16948), .dinb(asqrt[14] ), .dout(n16949));
  jand g16697(.dina(asqrt[13] ), .dinb(n15642), .dout(n16950));
  jor  g16698(.dina(n16950), .dinb(n15643), .dout(n16951));
  jand g16699(.dina(n16512), .dinb(n16951), .dout(n16952));
  jand g16700(.dina(n16952), .dinb(n16949), .dout(n16953));
  jor  g16701(.dina(n16953), .dinb(n16946), .dout(n16954));
  jor  g16702(.dina(n16954), .dinb(asqrt[15] ), .dout(n16955));
  jnot g16703(.din(n16517), .dout(n16956));
  jand g16704(.dina(n16956), .dinb(n16955), .dout(n16957));
  jor  g16705(.dina(n16957), .dinb(n16945), .dout(n16958));
  jor  g16706(.dina(n16958), .dinb(asqrt[16] ), .dout(n16959));
  jand g16707(.dina(n16524), .dinb(n16959), .dout(n16960));
  jor  g16708(.dina(n16960), .dinb(n16944), .dout(n16961));
  jor  g16709(.dina(n16961), .dinb(asqrt[17] ), .dout(n16962));
  jnot g16710(.din(n16532), .dout(n16963));
  jand g16711(.dina(n16963), .dinb(n16962), .dout(n16964));
  jor  g16712(.dina(n16964), .dinb(n16943), .dout(n16965));
  jor  g16713(.dina(n16965), .dinb(asqrt[18] ), .dout(n16966));
  jnot g16714(.din(n16539), .dout(n16967));
  jand g16715(.dina(n16967), .dinb(n16966), .dout(n16968));
  jor  g16716(.dina(n16968), .dinb(n16942), .dout(n16969));
  jor  g16717(.dina(n16969), .dinb(asqrt[19] ), .dout(n16970));
  jand g16718(.dina(n16546), .dinb(n16970), .dout(n16971));
  jor  g16719(.dina(n16971), .dinb(n16941), .dout(n16972));
  jor  g16720(.dina(n16972), .dinb(asqrt[20] ), .dout(n16973));
  jand g16721(.dina(n16554), .dinb(n16973), .dout(n16974));
  jor  g16722(.dina(n16974), .dinb(n16940), .dout(n16975));
  jor  g16723(.dina(n16975), .dinb(asqrt[21] ), .dout(n16976));
  jnot g16724(.din(n16562), .dout(n16977));
  jand g16725(.dina(n16977), .dinb(n16976), .dout(n16978));
  jor  g16726(.dina(n16978), .dinb(n16939), .dout(n16979));
  jor  g16727(.dina(n16979), .dinb(asqrt[22] ), .dout(n16980));
  jand g16728(.dina(n16569), .dinb(n16980), .dout(n16981));
  jor  g16729(.dina(n16981), .dinb(n16938), .dout(n16982));
  jor  g16730(.dina(n16982), .dinb(asqrt[23] ), .dout(n16983));
  jnot g16731(.din(n16577), .dout(n16984));
  jand g16732(.dina(n16984), .dinb(n16983), .dout(n16985));
  jor  g16733(.dina(n16985), .dinb(n16937), .dout(n16986));
  jor  g16734(.dina(n16986), .dinb(asqrt[24] ), .dout(n16987));
  jand g16735(.dina(n16584), .dinb(n16987), .dout(n16988));
  jor  g16736(.dina(n16988), .dinb(n16936), .dout(n16989));
  jor  g16737(.dina(n16989), .dinb(asqrt[25] ), .dout(n16990));
  jnot g16738(.din(n16592), .dout(n16991));
  jand g16739(.dina(n16991), .dinb(n16990), .dout(n16992));
  jor  g16740(.dina(n16992), .dinb(n16935), .dout(n16993));
  jor  g16741(.dina(n16993), .dinb(asqrt[26] ), .dout(n16994));
  jnot g16742(.din(n16599), .dout(n16995));
  jand g16743(.dina(n16995), .dinb(n16994), .dout(n16996));
  jor  g16744(.dina(n16996), .dinb(n16934), .dout(n16997));
  jor  g16745(.dina(n16997), .dinb(asqrt[27] ), .dout(n16998));
  jnot g16746(.din(n16606), .dout(n16999));
  jand g16747(.dina(n16999), .dinb(n16998), .dout(n17000));
  jor  g16748(.dina(n17000), .dinb(n16933), .dout(n17001));
  jor  g16749(.dina(n17001), .dinb(asqrt[28] ), .dout(n17002));
  jand g16750(.dina(n16613), .dinb(n17002), .dout(n17003));
  jor  g16751(.dina(n17003), .dinb(n16932), .dout(n17004));
  jor  g16752(.dina(n17004), .dinb(asqrt[29] ), .dout(n17005));
  jnot g16753(.din(n16621), .dout(n17006));
  jand g16754(.dina(n17006), .dinb(n17005), .dout(n17007));
  jor  g16755(.dina(n17007), .dinb(n16931), .dout(n17008));
  jor  g16756(.dina(n17008), .dinb(asqrt[30] ), .dout(n17009));
  jand g16757(.dina(n16628), .dinb(n17009), .dout(n17010));
  jor  g16758(.dina(n17010), .dinb(n16930), .dout(n17011));
  jor  g16759(.dina(n17011), .dinb(asqrt[31] ), .dout(n17012));
  jnot g16760(.din(n16636), .dout(n17013));
  jand g16761(.dina(n17013), .dinb(n17012), .dout(n17014));
  jor  g16762(.dina(n17014), .dinb(n16929), .dout(n17015));
  jor  g16763(.dina(n17015), .dinb(asqrt[32] ), .dout(n17016));
  jand g16764(.dina(n16643), .dinb(n17016), .dout(n17017));
  jor  g16765(.dina(n17017), .dinb(n16928), .dout(n17018));
  jor  g16766(.dina(n17018), .dinb(asqrt[33] ), .dout(n17019));
  jnot g16767(.din(n16651), .dout(n17020));
  jand g16768(.dina(n17020), .dinb(n17019), .dout(n17021));
  jor  g16769(.dina(n17021), .dinb(n16927), .dout(n17022));
  jor  g16770(.dina(n17022), .dinb(asqrt[34] ), .dout(n17023));
  jand g16771(.dina(n16658), .dinb(n17023), .dout(n17024));
  jor  g16772(.dina(n17024), .dinb(n16926), .dout(n17025));
  jor  g16773(.dina(n17025), .dinb(asqrt[35] ), .dout(n17026));
  jnot g16774(.din(n16666), .dout(n17027));
  jand g16775(.dina(n17027), .dinb(n17026), .dout(n17028));
  jor  g16776(.dina(n17028), .dinb(n16925), .dout(n17029));
  jor  g16777(.dina(n17029), .dinb(asqrt[36] ), .dout(n17030));
  jnot g16778(.din(n16673), .dout(n17031));
  jand g16779(.dina(n17031), .dinb(n17030), .dout(n17032));
  jor  g16780(.dina(n17032), .dinb(n16924), .dout(n17033));
  jor  g16781(.dina(n17033), .dinb(asqrt[37] ), .dout(n17034));
  jnot g16782(.din(n16680), .dout(n17035));
  jand g16783(.dina(n17035), .dinb(n17034), .dout(n17036));
  jor  g16784(.dina(n17036), .dinb(n16923), .dout(n17037));
  jor  g16785(.dina(n17037), .dinb(asqrt[38] ), .dout(n17038));
  jand g16786(.dina(n16687), .dinb(n17038), .dout(n17039));
  jor  g16787(.dina(n17039), .dinb(n16922), .dout(n17040));
  jor  g16788(.dina(n17040), .dinb(asqrt[39] ), .dout(n17041));
  jnot g16789(.din(n16695), .dout(n17042));
  jand g16790(.dina(n17042), .dinb(n17041), .dout(n17043));
  jor  g16791(.dina(n17043), .dinb(n16921), .dout(n17044));
  jor  g16792(.dina(n17044), .dinb(asqrt[40] ), .dout(n17045));
  jand g16793(.dina(n16702), .dinb(n17045), .dout(n17046));
  jor  g16794(.dina(n17046), .dinb(n16920), .dout(n17047));
  jor  g16795(.dina(n17047), .dinb(asqrt[41] ), .dout(n17048));
  jnot g16796(.din(n16710), .dout(n17049));
  jand g16797(.dina(n17049), .dinb(n17048), .dout(n17050));
  jor  g16798(.dina(n17050), .dinb(n16919), .dout(n17051));
  jor  g16799(.dina(n17051), .dinb(asqrt[42] ), .dout(n17052));
  jnot g16800(.din(n16717), .dout(n17053));
  jand g16801(.dina(n17053), .dinb(n17052), .dout(n17054));
  jor  g16802(.dina(n17054), .dinb(n16918), .dout(n17055));
  jor  g16803(.dina(n17055), .dinb(asqrt[43] ), .dout(n17056));
  jnot g16804(.din(n16724), .dout(n17057));
  jand g16805(.dina(n17057), .dinb(n17056), .dout(n17058));
  jor  g16806(.dina(n17058), .dinb(n16917), .dout(n17059));
  jor  g16807(.dina(n17059), .dinb(asqrt[44] ), .dout(n17060));
  jand g16808(.dina(n16731), .dinb(n17060), .dout(n17061));
  jor  g16809(.dina(n17061), .dinb(n16916), .dout(n17062));
  jor  g16810(.dina(n17062), .dinb(asqrt[45] ), .dout(n17063));
  jnot g16811(.din(n16739), .dout(n17064));
  jand g16812(.dina(n17064), .dinb(n17063), .dout(n17065));
  jor  g16813(.dina(n17065), .dinb(n16915), .dout(n17066));
  jor  g16814(.dina(n17066), .dinb(asqrt[46] ), .dout(n17067));
  jand g16815(.dina(n16746), .dinb(n17067), .dout(n17068));
  jor  g16816(.dina(n17068), .dinb(n16914), .dout(n17069));
  jor  g16817(.dina(n17069), .dinb(asqrt[47] ), .dout(n17070));
  jnot g16818(.din(n16754), .dout(n17071));
  jand g16819(.dina(n17071), .dinb(n17070), .dout(n17072));
  jor  g16820(.dina(n17072), .dinb(n16913), .dout(n17073));
  jor  g16821(.dina(n17073), .dinb(asqrt[48] ), .dout(n17074));
  jnot g16822(.din(n16761), .dout(n17075));
  jand g16823(.dina(n17075), .dinb(n17074), .dout(n17076));
  jor  g16824(.dina(n17076), .dinb(n16912), .dout(n17077));
  jor  g16825(.dina(n17077), .dinb(asqrt[49] ), .dout(n17078));
  jand g16826(.dina(n16768), .dinb(n17078), .dout(n17079));
  jor  g16827(.dina(n17079), .dinb(n16911), .dout(n17080));
  jor  g16828(.dina(n17080), .dinb(asqrt[50] ), .dout(n17081));
  jand g16829(.dina(n17081), .dinb(n16775), .dout(n17082));
  jor  g16830(.dina(n17082), .dinb(n16910), .dout(n17083));
  jor  g16831(.dina(n17083), .dinb(asqrt[51] ), .dout(n17084));
  jnot g16832(.din(n16784), .dout(n17085));
  jand g16833(.dina(n17085), .dinb(n17084), .dout(n17086));
  jor  g16834(.dina(n17086), .dinb(n16909), .dout(n17087));
  jor  g16835(.dina(n17087), .dinb(asqrt[52] ), .dout(n17088));
  jand g16836(.dina(n16791), .dinb(n17088), .dout(n17089));
  jor  g16837(.dina(n17089), .dinb(n16908), .dout(n17090));
  jor  g16838(.dina(n17090), .dinb(asqrt[53] ), .dout(n17091));
  jnot g16839(.din(n16799), .dout(n17092));
  jand g16840(.dina(n17092), .dinb(n17091), .dout(n17093));
  jor  g16841(.dina(n17093), .dinb(n16907), .dout(n17094));
  jor  g16842(.dina(n17094), .dinb(asqrt[54] ), .dout(n17095));
  jand g16843(.dina(n16806), .dinb(n17095), .dout(n17096));
  jor  g16844(.dina(n17096), .dinb(n16906), .dout(n17097));
  jor  g16845(.dina(n17097), .dinb(asqrt[55] ), .dout(n17098));
  jnot g16846(.din(n16814), .dout(n17099));
  jand g16847(.dina(n17099), .dinb(n17098), .dout(n17100));
  jor  g16848(.dina(n17100), .dinb(n16905), .dout(n17101));
  jor  g16849(.dina(n17101), .dinb(asqrt[56] ), .dout(n17102));
  jnot g16850(.din(n16821), .dout(n17103));
  jand g16851(.dina(n17103), .dinb(n17102), .dout(n17104));
  jor  g16852(.dina(n17104), .dinb(n16904), .dout(n17105));
  jor  g16853(.dina(n17105), .dinb(asqrt[57] ), .dout(n17106));
  jnot g16854(.din(n16828), .dout(n17107));
  jand g16855(.dina(n17107), .dinb(n17106), .dout(n17108));
  jor  g16856(.dina(n17108), .dinb(n16903), .dout(n17109));
  jor  g16857(.dina(n17109), .dinb(asqrt[58] ), .dout(n17110));
  jand g16858(.dina(n16835), .dinb(n17110), .dout(n17111));
  jor  g16859(.dina(n17111), .dinb(n16902), .dout(n17112));
  jor  g16860(.dina(n17112), .dinb(asqrt[59] ), .dout(n17113));
  jnot g16861(.din(n16843), .dout(n17114));
  jand g16862(.dina(n17114), .dinb(n17113), .dout(n17115));
  jor  g16863(.dina(n17115), .dinb(n16901), .dout(n17116));
  jor  g16864(.dina(n17116), .dinb(asqrt[60] ), .dout(n17117));
  jand g16865(.dina(n16850), .dinb(n17117), .dout(n17118));
  jor  g16866(.dina(n17118), .dinb(n16900), .dout(n17119));
  jor  g16867(.dina(n17119), .dinb(asqrt[61] ), .dout(n17120));
  jnot g16868(.din(n16858), .dout(n17121));
  jand g16869(.dina(n17121), .dinb(n17120), .dout(n17122));
  jor  g16870(.dina(n17122), .dinb(n16899), .dout(n17123));
  jor  g16871(.dina(n17123), .dinb(asqrt[62] ), .dout(n17124));
  jand g16872(.dina(n16865), .dinb(n17124), .dout(n17125));
  jor  g16873(.dina(n17125), .dinb(n16898), .dout(n17126));
  jand g16874(.dina(n17126), .dinb(n16492), .dout(n17127));
  jnot g16875(.din(n16872), .dout(n17128));
  jand g16876(.dina(n17128), .dinb(n17127), .dout(n17129));
  jand g16877(.dina(n17129), .dinb(n16485), .dout(n17130));
  jor  g16878(.dina(n17130), .dinb(asqrt[63] ), .dout(n17131));
  jand g16879(.dina(n16880), .dinb(n17131), .dout(n17132));
  jand g16880(.dina(n17132), .dinb(n16896), .dout(n17134));
  jor  g16881(.dina(n17134), .dinb(n16895), .dout(n17135));
  jand g16882(.dina(n17135), .dinb(n16894), .dout(n17136));
  jand g16883(.dina(n17136), .dinb(n16892), .dout(n17137));
  jor  g16884(.dina(n17137), .dinb(n16891), .dout(n17138));
  jand g16885(.dina(n17138), .dinb(asqrt[14] ), .dout(n17139));
  jor  g16886(.dina(n17138), .dinb(asqrt[14] ), .dout(n17140));
  jand g16887(.dina(asqrt[12] ), .dinb(n16496), .dout(n17141));
  jand g16888(.dina(n16896), .dinb(asqrt[13] ), .dout(n17142));
  jand g16889(.dina(n17142), .dinb(n17131), .dout(n17143));
  jand g16890(.dina(n17143), .dinb(n16879), .dout(n17144));
  jor  g16891(.dina(n17144), .dinb(n17141), .dout(n17145));
  jxor g16892(.dina(n17145), .dinb(a[26] ), .dout(n17146));
  jnot g16893(.din(n17146), .dout(n17147));
  jand g16894(.dina(n17147), .dinb(n17140), .dout(n17148));
  jor  g16895(.dina(n17148), .dinb(n17139), .dout(n17149));
  jand g16896(.dina(n17149), .dinb(asqrt[15] ), .dout(n17150));
  jor  g16897(.dina(n17149), .dinb(asqrt[15] ), .dout(n17151));
  jxor g16898(.dina(n16500), .dinb(n15878), .dout(n17152));
  jand g16899(.dina(n17152), .dinb(asqrt[12] ), .dout(n17153));
  jxor g16900(.dina(n17153), .dinb(n16952), .dout(n17154));
  jand g16901(.dina(n17154), .dinb(n17151), .dout(n17155));
  jor  g16902(.dina(n17155), .dinb(n17150), .dout(n17156));
  jand g16903(.dina(n17156), .dinb(asqrt[16] ), .dout(n17157));
  jor  g16904(.dina(n17156), .dinb(asqrt[16] ), .dout(n17158));
  jxor g16905(.dina(n16508), .dinb(n15260), .dout(n17159));
  jand g16906(.dina(n17159), .dinb(asqrt[12] ), .dout(n17160));
  jxor g16907(.dina(n17160), .dinb(n16517), .dout(n17161));
  jnot g16908(.din(n17161), .dout(n17162));
  jand g16909(.dina(n17162), .dinb(n17158), .dout(n17163));
  jor  g16910(.dina(n17163), .dinb(n17157), .dout(n17164));
  jand g16911(.dina(n17164), .dinb(asqrt[17] ), .dout(n17165));
  jor  g16912(.dina(n17164), .dinb(asqrt[17] ), .dout(n17166));
  jxor g16913(.dina(n16519), .dinb(n14674), .dout(n17167));
  jand g16914(.dina(n17167), .dinb(asqrt[12] ), .dout(n17168));
  jxor g16915(.dina(n17168), .dinb(n16524), .dout(n17169));
  jand g16916(.dina(n17169), .dinb(n17166), .dout(n17170));
  jor  g16917(.dina(n17170), .dinb(n17165), .dout(n17171));
  jand g16918(.dina(n17171), .dinb(asqrt[18] ), .dout(n17172));
  jor  g16919(.dina(n17171), .dinb(asqrt[18] ), .dout(n17173));
  jxor g16920(.dina(n16527), .dinb(n14078), .dout(n17174));
  jand g16921(.dina(n17174), .dinb(asqrt[12] ), .dout(n17175));
  jxor g16922(.dina(n17175), .dinb(n16532), .dout(n17176));
  jnot g16923(.din(n17176), .dout(n17177));
  jand g16924(.dina(n17177), .dinb(n17173), .dout(n17178));
  jor  g16925(.dina(n17178), .dinb(n17172), .dout(n17179));
  jand g16926(.dina(n17179), .dinb(asqrt[19] ), .dout(n17180));
  jor  g16927(.dina(n17179), .dinb(asqrt[19] ), .dout(n17181));
  jxor g16928(.dina(n16534), .dinb(n13515), .dout(n17182));
  jand g16929(.dina(n17182), .dinb(asqrt[12] ), .dout(n17183));
  jxor g16930(.dina(n17183), .dinb(n16539), .dout(n17184));
  jnot g16931(.din(n17184), .dout(n17185));
  jand g16932(.dina(n17185), .dinb(n17181), .dout(n17186));
  jor  g16933(.dina(n17186), .dinb(n17180), .dout(n17187));
  jand g16934(.dina(n17187), .dinb(asqrt[20] ), .dout(n17188));
  jor  g16935(.dina(n17187), .dinb(asqrt[20] ), .dout(n17189));
  jxor g16936(.dina(n16541), .dinb(n12947), .dout(n17190));
  jand g16937(.dina(n17190), .dinb(asqrt[12] ), .dout(n17191));
  jxor g16938(.dina(n17191), .dinb(n16546), .dout(n17192));
  jand g16939(.dina(n17192), .dinb(n17189), .dout(n17193));
  jor  g16940(.dina(n17193), .dinb(n17188), .dout(n17194));
  jand g16941(.dina(n17194), .dinb(asqrt[21] ), .dout(n17195));
  jor  g16942(.dina(n17194), .dinb(asqrt[21] ), .dout(n17196));
  jxor g16943(.dina(n16549), .dinb(n12410), .dout(n17197));
  jand g16944(.dina(n17197), .dinb(asqrt[12] ), .dout(n17198));
  jxor g16945(.dina(n17198), .dinb(n16554), .dout(n17199));
  jand g16946(.dina(n17199), .dinb(n17196), .dout(n17200));
  jor  g16947(.dina(n17200), .dinb(n17195), .dout(n17201));
  jand g16948(.dina(n17201), .dinb(asqrt[22] ), .dout(n17202));
  jor  g16949(.dina(n17201), .dinb(asqrt[22] ), .dout(n17203));
  jxor g16950(.dina(n16557), .dinb(n11858), .dout(n17204));
  jand g16951(.dina(n17204), .dinb(asqrt[12] ), .dout(n17205));
  jxor g16952(.dina(n17205), .dinb(n16562), .dout(n17206));
  jnot g16953(.din(n17206), .dout(n17207));
  jand g16954(.dina(n17207), .dinb(n17203), .dout(n17208));
  jor  g16955(.dina(n17208), .dinb(n17202), .dout(n17209));
  jand g16956(.dina(n17209), .dinb(asqrt[23] ), .dout(n17210));
  jor  g16957(.dina(n17209), .dinb(asqrt[23] ), .dout(n17211));
  jxor g16958(.dina(n16564), .dinb(n11347), .dout(n17212));
  jand g16959(.dina(n17212), .dinb(asqrt[12] ), .dout(n17213));
  jxor g16960(.dina(n17213), .dinb(n16569), .dout(n17214));
  jand g16961(.dina(n17214), .dinb(n17211), .dout(n17215));
  jor  g16962(.dina(n17215), .dinb(n17210), .dout(n17216));
  jand g16963(.dina(n17216), .dinb(asqrt[24] ), .dout(n17217));
  jor  g16964(.dina(n17216), .dinb(asqrt[24] ), .dout(n17218));
  jxor g16965(.dina(n16572), .dinb(n10824), .dout(n17219));
  jand g16966(.dina(n17219), .dinb(asqrt[12] ), .dout(n17220));
  jxor g16967(.dina(n17220), .dinb(n16577), .dout(n17221));
  jnot g16968(.din(n17221), .dout(n17222));
  jand g16969(.dina(n17222), .dinb(n17218), .dout(n17223));
  jor  g16970(.dina(n17223), .dinb(n17217), .dout(n17224));
  jand g16971(.dina(n17224), .dinb(asqrt[25] ), .dout(n17225));
  jor  g16972(.dina(n17224), .dinb(asqrt[25] ), .dout(n17226));
  jxor g16973(.dina(n16579), .dinb(n10328), .dout(n17227));
  jand g16974(.dina(n17227), .dinb(asqrt[12] ), .dout(n17228));
  jxor g16975(.dina(n17228), .dinb(n16584), .dout(n17229));
  jand g16976(.dina(n17229), .dinb(n17226), .dout(n17230));
  jor  g16977(.dina(n17230), .dinb(n17225), .dout(n17231));
  jand g16978(.dina(n17231), .dinb(asqrt[26] ), .dout(n17232));
  jor  g16979(.dina(n17231), .dinb(asqrt[26] ), .dout(n17233));
  jxor g16980(.dina(n16587), .dinb(n9832), .dout(n17234));
  jand g16981(.dina(n17234), .dinb(asqrt[12] ), .dout(n17235));
  jxor g16982(.dina(n17235), .dinb(n16592), .dout(n17236));
  jnot g16983(.din(n17236), .dout(n17237));
  jand g16984(.dina(n17237), .dinb(n17233), .dout(n17238));
  jor  g16985(.dina(n17238), .dinb(n17232), .dout(n17239));
  jand g16986(.dina(n17239), .dinb(asqrt[27] ), .dout(n17240));
  jor  g16987(.dina(n17239), .dinb(asqrt[27] ), .dout(n17241));
  jxor g16988(.dina(n16594), .dinb(n9369), .dout(n17242));
  jand g16989(.dina(n17242), .dinb(asqrt[12] ), .dout(n17243));
  jxor g16990(.dina(n17243), .dinb(n16599), .dout(n17244));
  jnot g16991(.din(n17244), .dout(n17245));
  jand g16992(.dina(n17245), .dinb(n17241), .dout(n17246));
  jor  g16993(.dina(n17246), .dinb(n17240), .dout(n17247));
  jand g16994(.dina(n17247), .dinb(asqrt[28] ), .dout(n17248));
  jor  g16995(.dina(n17247), .dinb(asqrt[28] ), .dout(n17249));
  jxor g16996(.dina(n16601), .dinb(n8890), .dout(n17250));
  jand g16997(.dina(n17250), .dinb(asqrt[12] ), .dout(n17251));
  jxor g16998(.dina(n17251), .dinb(n16606), .dout(n17252));
  jnot g16999(.din(n17252), .dout(n17253));
  jand g17000(.dina(n17253), .dinb(n17249), .dout(n17254));
  jor  g17001(.dina(n17254), .dinb(n17248), .dout(n17255));
  jand g17002(.dina(n17255), .dinb(asqrt[29] ), .dout(n17256));
  jor  g17003(.dina(n17255), .dinb(asqrt[29] ), .dout(n17257));
  jxor g17004(.dina(n16608), .dinb(n8449), .dout(n17258));
  jand g17005(.dina(n17258), .dinb(asqrt[12] ), .dout(n17259));
  jxor g17006(.dina(n17259), .dinb(n16613), .dout(n17260));
  jand g17007(.dina(n17260), .dinb(n17257), .dout(n17261));
  jor  g17008(.dina(n17261), .dinb(n17256), .dout(n17262));
  jand g17009(.dina(n17262), .dinb(asqrt[30] ), .dout(n17263));
  jor  g17010(.dina(n17262), .dinb(asqrt[30] ), .dout(n17264));
  jxor g17011(.dina(n16616), .dinb(n8003), .dout(n17265));
  jand g17012(.dina(n17265), .dinb(asqrt[12] ), .dout(n17266));
  jxor g17013(.dina(n17266), .dinb(n16621), .dout(n17267));
  jnot g17014(.din(n17267), .dout(n17268));
  jand g17015(.dina(n17268), .dinb(n17264), .dout(n17269));
  jor  g17016(.dina(n17269), .dinb(n17263), .dout(n17270));
  jand g17017(.dina(n17270), .dinb(asqrt[31] ), .dout(n17271));
  jor  g17018(.dina(n17270), .dinb(asqrt[31] ), .dout(n17272));
  jxor g17019(.dina(n16623), .dinb(n7581), .dout(n17273));
  jand g17020(.dina(n17273), .dinb(asqrt[12] ), .dout(n17274));
  jxor g17021(.dina(n17274), .dinb(n16628), .dout(n17275));
  jand g17022(.dina(n17275), .dinb(n17272), .dout(n17276));
  jor  g17023(.dina(n17276), .dinb(n17271), .dout(n17277));
  jand g17024(.dina(n17277), .dinb(asqrt[32] ), .dout(n17278));
  jor  g17025(.dina(n17277), .dinb(asqrt[32] ), .dout(n17279));
  jxor g17026(.dina(n16631), .dinb(n7154), .dout(n17280));
  jand g17027(.dina(n17280), .dinb(asqrt[12] ), .dout(n17281));
  jxor g17028(.dina(n17281), .dinb(n16636), .dout(n17282));
  jnot g17029(.din(n17282), .dout(n17283));
  jand g17030(.dina(n17283), .dinb(n17279), .dout(n17284));
  jor  g17031(.dina(n17284), .dinb(n17278), .dout(n17285));
  jand g17032(.dina(n17285), .dinb(asqrt[33] ), .dout(n17286));
  jor  g17033(.dina(n17285), .dinb(asqrt[33] ), .dout(n17287));
  jxor g17034(.dina(n16638), .dinb(n6758), .dout(n17288));
  jand g17035(.dina(n17288), .dinb(asqrt[12] ), .dout(n17289));
  jxor g17036(.dina(n17289), .dinb(n16643), .dout(n17290));
  jand g17037(.dina(n17290), .dinb(n17287), .dout(n17291));
  jor  g17038(.dina(n17291), .dinb(n17286), .dout(n17292));
  jand g17039(.dina(n17292), .dinb(asqrt[34] ), .dout(n17293));
  jor  g17040(.dina(n17292), .dinb(asqrt[34] ), .dout(n17294));
  jxor g17041(.dina(n16646), .dinb(n6357), .dout(n17295));
  jand g17042(.dina(n17295), .dinb(asqrt[12] ), .dout(n17296));
  jxor g17043(.dina(n17296), .dinb(n16651), .dout(n17297));
  jnot g17044(.din(n17297), .dout(n17298));
  jand g17045(.dina(n17298), .dinb(n17294), .dout(n17299));
  jor  g17046(.dina(n17299), .dinb(n17293), .dout(n17300));
  jand g17047(.dina(n17300), .dinb(asqrt[35] ), .dout(n17301));
  jor  g17048(.dina(n17300), .dinb(asqrt[35] ), .dout(n17302));
  jxor g17049(.dina(n16653), .dinb(n5989), .dout(n17303));
  jand g17050(.dina(n17303), .dinb(asqrt[12] ), .dout(n17304));
  jxor g17051(.dina(n17304), .dinb(n16658), .dout(n17305));
  jand g17052(.dina(n17305), .dinb(n17302), .dout(n17306));
  jor  g17053(.dina(n17306), .dinb(n17301), .dout(n17307));
  jand g17054(.dina(n17307), .dinb(asqrt[36] ), .dout(n17308));
  jor  g17055(.dina(n17307), .dinb(asqrt[36] ), .dout(n17309));
  jxor g17056(.dina(n16661), .dinb(n5606), .dout(n17310));
  jand g17057(.dina(n17310), .dinb(asqrt[12] ), .dout(n17311));
  jxor g17058(.dina(n17311), .dinb(n16666), .dout(n17312));
  jnot g17059(.din(n17312), .dout(n17313));
  jand g17060(.dina(n17313), .dinb(n17309), .dout(n17314));
  jor  g17061(.dina(n17314), .dinb(n17308), .dout(n17315));
  jand g17062(.dina(n17315), .dinb(asqrt[37] ), .dout(n17316));
  jor  g17063(.dina(n17315), .dinb(asqrt[37] ), .dout(n17317));
  jxor g17064(.dina(n16668), .dinb(n5259), .dout(n17318));
  jand g17065(.dina(n17318), .dinb(asqrt[12] ), .dout(n17319));
  jxor g17066(.dina(n17319), .dinb(n16673), .dout(n17320));
  jnot g17067(.din(n17320), .dout(n17321));
  jand g17068(.dina(n17321), .dinb(n17317), .dout(n17322));
  jor  g17069(.dina(n17322), .dinb(n17316), .dout(n17323));
  jand g17070(.dina(n17323), .dinb(asqrt[38] ), .dout(n17324));
  jor  g17071(.dina(n17323), .dinb(asqrt[38] ), .dout(n17325));
  jxor g17072(.dina(n16675), .dinb(n4902), .dout(n17326));
  jand g17073(.dina(n17326), .dinb(asqrt[12] ), .dout(n17327));
  jxor g17074(.dina(n17327), .dinb(n16680), .dout(n17328));
  jnot g17075(.din(n17328), .dout(n17329));
  jand g17076(.dina(n17329), .dinb(n17325), .dout(n17330));
  jor  g17077(.dina(n17330), .dinb(n17324), .dout(n17331));
  jand g17078(.dina(n17331), .dinb(asqrt[39] ), .dout(n17332));
  jor  g17079(.dina(n17331), .dinb(asqrt[39] ), .dout(n17333));
  jxor g17080(.dina(n16682), .dinb(n4582), .dout(n17334));
  jand g17081(.dina(n17334), .dinb(asqrt[12] ), .dout(n17335));
  jxor g17082(.dina(n17335), .dinb(n16687), .dout(n17336));
  jand g17083(.dina(n17336), .dinb(n17333), .dout(n17337));
  jor  g17084(.dina(n17337), .dinb(n17332), .dout(n17338));
  jand g17085(.dina(n17338), .dinb(asqrt[40] ), .dout(n17339));
  jor  g17086(.dina(n17338), .dinb(asqrt[40] ), .dout(n17340));
  jxor g17087(.dina(n16690), .dinb(n4249), .dout(n17341));
  jand g17088(.dina(n17341), .dinb(asqrt[12] ), .dout(n17342));
  jxor g17089(.dina(n17342), .dinb(n16695), .dout(n17343));
  jnot g17090(.din(n17343), .dout(n17344));
  jand g17091(.dina(n17344), .dinb(n17340), .dout(n17345));
  jor  g17092(.dina(n17345), .dinb(n17339), .dout(n17346));
  jand g17093(.dina(n17346), .dinb(asqrt[41] ), .dout(n17347));
  jor  g17094(.dina(n17346), .dinb(asqrt[41] ), .dout(n17348));
  jxor g17095(.dina(n16697), .dinb(n3955), .dout(n17349));
  jand g17096(.dina(n17349), .dinb(asqrt[12] ), .dout(n17350));
  jxor g17097(.dina(n17350), .dinb(n16702), .dout(n17351));
  jand g17098(.dina(n17351), .dinb(n17348), .dout(n17352));
  jor  g17099(.dina(n17352), .dinb(n17347), .dout(n17353));
  jand g17100(.dina(n17353), .dinb(asqrt[42] ), .dout(n17354));
  jor  g17101(.dina(n17353), .dinb(asqrt[42] ), .dout(n17355));
  jxor g17102(.dina(n16705), .dinb(n3642), .dout(n17356));
  jand g17103(.dina(n17356), .dinb(asqrt[12] ), .dout(n17357));
  jxor g17104(.dina(n17357), .dinb(n16710), .dout(n17358));
  jnot g17105(.din(n17358), .dout(n17359));
  jand g17106(.dina(n17359), .dinb(n17355), .dout(n17360));
  jor  g17107(.dina(n17360), .dinb(n17354), .dout(n17361));
  jand g17108(.dina(n17361), .dinb(asqrt[43] ), .dout(n17362));
  jor  g17109(.dina(n17361), .dinb(asqrt[43] ), .dout(n17363));
  jxor g17110(.dina(n16712), .dinb(n3368), .dout(n17364));
  jand g17111(.dina(n17364), .dinb(asqrt[12] ), .dout(n17365));
  jxor g17112(.dina(n17365), .dinb(n16717), .dout(n17366));
  jnot g17113(.din(n17366), .dout(n17367));
  jand g17114(.dina(n17367), .dinb(n17363), .dout(n17368));
  jor  g17115(.dina(n17368), .dinb(n17362), .dout(n17369));
  jand g17116(.dina(n17369), .dinb(asqrt[44] ), .dout(n17370));
  jor  g17117(.dina(n17369), .dinb(asqrt[44] ), .dout(n17371));
  jxor g17118(.dina(n16719), .dinb(n3089), .dout(n17372));
  jand g17119(.dina(n17372), .dinb(asqrt[12] ), .dout(n17373));
  jxor g17120(.dina(n17373), .dinb(n16724), .dout(n17374));
  jnot g17121(.din(n17374), .dout(n17375));
  jand g17122(.dina(n17375), .dinb(n17371), .dout(n17376));
  jor  g17123(.dina(n17376), .dinb(n17370), .dout(n17377));
  jand g17124(.dina(n17377), .dinb(asqrt[45] ), .dout(n17378));
  jor  g17125(.dina(n17377), .dinb(asqrt[45] ), .dout(n17379));
  jxor g17126(.dina(n16726), .dinb(n2833), .dout(n17380));
  jand g17127(.dina(n17380), .dinb(asqrt[12] ), .dout(n17381));
  jxor g17128(.dina(n17381), .dinb(n16731), .dout(n17382));
  jand g17129(.dina(n17382), .dinb(n17379), .dout(n17383));
  jor  g17130(.dina(n17383), .dinb(n17378), .dout(n17384));
  jand g17131(.dina(n17384), .dinb(asqrt[46] ), .dout(n17385));
  jor  g17132(.dina(n17384), .dinb(asqrt[46] ), .dout(n17386));
  jxor g17133(.dina(n16734), .dinb(n2572), .dout(n17387));
  jand g17134(.dina(n17387), .dinb(asqrt[12] ), .dout(n17388));
  jxor g17135(.dina(n17388), .dinb(n16739), .dout(n17389));
  jnot g17136(.din(n17389), .dout(n17390));
  jand g17137(.dina(n17390), .dinb(n17386), .dout(n17391));
  jor  g17138(.dina(n17391), .dinb(n17385), .dout(n17392));
  jand g17139(.dina(n17392), .dinb(asqrt[47] ), .dout(n17393));
  jor  g17140(.dina(n17392), .dinb(asqrt[47] ), .dout(n17394));
  jxor g17141(.dina(n16741), .dinb(n2345), .dout(n17395));
  jand g17142(.dina(n17395), .dinb(asqrt[12] ), .dout(n17396));
  jxor g17143(.dina(n17396), .dinb(n16746), .dout(n17397));
  jand g17144(.dina(n17397), .dinb(n17394), .dout(n17398));
  jor  g17145(.dina(n17398), .dinb(n17393), .dout(n17399));
  jand g17146(.dina(n17399), .dinb(asqrt[48] ), .dout(n17400));
  jor  g17147(.dina(n17399), .dinb(asqrt[48] ), .dout(n17401));
  jxor g17148(.dina(n16749), .dinb(n2108), .dout(n17402));
  jand g17149(.dina(n17402), .dinb(asqrt[12] ), .dout(n17403));
  jxor g17150(.dina(n17403), .dinb(n16754), .dout(n17404));
  jnot g17151(.din(n17404), .dout(n17405));
  jand g17152(.dina(n17405), .dinb(n17401), .dout(n17406));
  jor  g17153(.dina(n17406), .dinb(n17400), .dout(n17407));
  jand g17154(.dina(n17407), .dinb(asqrt[49] ), .dout(n17408));
  jor  g17155(.dina(n17407), .dinb(asqrt[49] ), .dout(n17409));
  jxor g17156(.dina(n16756), .dinb(n1912), .dout(n17410));
  jand g17157(.dina(n17410), .dinb(asqrt[12] ), .dout(n17411));
  jxor g17158(.dina(n17411), .dinb(n16761), .dout(n17412));
  jnot g17159(.din(n17412), .dout(n17413));
  jand g17160(.dina(n17413), .dinb(n17409), .dout(n17414));
  jor  g17161(.dina(n17414), .dinb(n17408), .dout(n17415));
  jand g17162(.dina(n17415), .dinb(asqrt[50] ), .dout(n17416));
  jor  g17163(.dina(n17415), .dinb(asqrt[50] ), .dout(n17417));
  jxor g17164(.dina(n16763), .dinb(n1699), .dout(n17418));
  jand g17165(.dina(n17418), .dinb(asqrt[12] ), .dout(n17419));
  jxor g17166(.dina(n17419), .dinb(n16768), .dout(n17420));
  jand g17167(.dina(n17420), .dinb(n17417), .dout(n17421));
  jor  g17168(.dina(n17421), .dinb(n17416), .dout(n17422));
  jand g17169(.dina(n17422), .dinb(asqrt[51] ), .dout(n17423));
  jxor g17170(.dina(n16771), .dinb(n1516), .dout(n17424));
  jand g17171(.dina(n17424), .dinb(asqrt[12] ), .dout(n17425));
  jxor g17172(.dina(n17425), .dinb(n16775), .dout(n17426));
  jor  g17173(.dina(n17422), .dinb(asqrt[51] ), .dout(n17427));
  jand g17174(.dina(n17427), .dinb(n17426), .dout(n17428));
  jor  g17175(.dina(n17428), .dinb(n17423), .dout(n17429));
  jand g17176(.dina(n17429), .dinb(asqrt[52] ), .dout(n17430));
  jor  g17177(.dina(n17429), .dinb(asqrt[52] ), .dout(n17431));
  jxor g17178(.dina(n16779), .dinb(n1332), .dout(n17432));
  jand g17179(.dina(n17432), .dinb(asqrt[12] ), .dout(n17433));
  jxor g17180(.dina(n17433), .dinb(n16784), .dout(n17434));
  jnot g17181(.din(n17434), .dout(n17435));
  jand g17182(.dina(n17435), .dinb(n17431), .dout(n17436));
  jor  g17183(.dina(n17436), .dinb(n17430), .dout(n17437));
  jand g17184(.dina(n17437), .dinb(asqrt[53] ), .dout(n17438));
  jor  g17185(.dina(n17437), .dinb(asqrt[53] ), .dout(n17439));
  jxor g17186(.dina(n16786), .dinb(n1173), .dout(n17440));
  jand g17187(.dina(n17440), .dinb(asqrt[12] ), .dout(n17441));
  jxor g17188(.dina(n17441), .dinb(n16791), .dout(n17442));
  jand g17189(.dina(n17442), .dinb(n17439), .dout(n17443));
  jor  g17190(.dina(n17443), .dinb(n17438), .dout(n17444));
  jand g17191(.dina(n17444), .dinb(asqrt[54] ), .dout(n17445));
  jor  g17192(.dina(n17444), .dinb(asqrt[54] ), .dout(n17446));
  jxor g17193(.dina(n16794), .dinb(n1008), .dout(n17447));
  jand g17194(.dina(n17447), .dinb(asqrt[12] ), .dout(n17448));
  jxor g17195(.dina(n17448), .dinb(n16799), .dout(n17449));
  jnot g17196(.din(n17449), .dout(n17450));
  jand g17197(.dina(n17450), .dinb(n17446), .dout(n17451));
  jor  g17198(.dina(n17451), .dinb(n17445), .dout(n17452));
  jand g17199(.dina(n17452), .dinb(asqrt[55] ), .dout(n17453));
  jor  g17200(.dina(n17452), .dinb(asqrt[55] ), .dout(n17454));
  jxor g17201(.dina(n16801), .dinb(n884), .dout(n17455));
  jand g17202(.dina(n17455), .dinb(asqrt[12] ), .dout(n17456));
  jxor g17203(.dina(n17456), .dinb(n16806), .dout(n17457));
  jand g17204(.dina(n17457), .dinb(n17454), .dout(n17458));
  jor  g17205(.dina(n17458), .dinb(n17453), .dout(n17459));
  jand g17206(.dina(n17459), .dinb(asqrt[56] ), .dout(n17460));
  jor  g17207(.dina(n17459), .dinb(asqrt[56] ), .dout(n17461));
  jxor g17208(.dina(n16809), .dinb(n743), .dout(n17462));
  jand g17209(.dina(n17462), .dinb(asqrt[12] ), .dout(n17463));
  jxor g17210(.dina(n17463), .dinb(n16814), .dout(n17464));
  jnot g17211(.din(n17464), .dout(n17465));
  jand g17212(.dina(n17465), .dinb(n17461), .dout(n17466));
  jor  g17213(.dina(n17466), .dinb(n17460), .dout(n17467));
  jand g17214(.dina(n17467), .dinb(asqrt[57] ), .dout(n17468));
  jor  g17215(.dina(n17467), .dinb(asqrt[57] ), .dout(n17469));
  jxor g17216(.dina(n16816), .dinb(n635), .dout(n17470));
  jand g17217(.dina(n17470), .dinb(asqrt[12] ), .dout(n17471));
  jxor g17218(.dina(n17471), .dinb(n16821), .dout(n17472));
  jnot g17219(.din(n17472), .dout(n17473));
  jand g17220(.dina(n17473), .dinb(n17469), .dout(n17474));
  jor  g17221(.dina(n17474), .dinb(n17468), .dout(n17475));
  jand g17222(.dina(n17475), .dinb(asqrt[58] ), .dout(n17476));
  jor  g17223(.dina(n17475), .dinb(asqrt[58] ), .dout(n17477));
  jxor g17224(.dina(n16823), .dinb(n515), .dout(n17478));
  jand g17225(.dina(n17478), .dinb(asqrt[12] ), .dout(n17479));
  jxor g17226(.dina(n17479), .dinb(n16828), .dout(n17480));
  jnot g17227(.din(n17480), .dout(n17481));
  jand g17228(.dina(n17481), .dinb(n17477), .dout(n17482));
  jor  g17229(.dina(n17482), .dinb(n17476), .dout(n17483));
  jand g17230(.dina(n17483), .dinb(asqrt[59] ), .dout(n17484));
  jor  g17231(.dina(n17483), .dinb(asqrt[59] ), .dout(n17485));
  jxor g17232(.dina(n16830), .dinb(n443), .dout(n17486));
  jand g17233(.dina(n17486), .dinb(asqrt[12] ), .dout(n17487));
  jxor g17234(.dina(n17487), .dinb(n16835), .dout(n17488));
  jand g17235(.dina(n17488), .dinb(n17485), .dout(n17489));
  jor  g17236(.dina(n17489), .dinb(n17484), .dout(n17490));
  jand g17237(.dina(n17490), .dinb(asqrt[60] ), .dout(n17491));
  jor  g17238(.dina(n17490), .dinb(asqrt[60] ), .dout(n17492));
  jxor g17239(.dina(n16838), .dinb(n352), .dout(n17493));
  jand g17240(.dina(n17493), .dinb(asqrt[12] ), .dout(n17494));
  jxor g17241(.dina(n17494), .dinb(n16843), .dout(n17495));
  jnot g17242(.din(n17495), .dout(n17496));
  jand g17243(.dina(n17496), .dinb(n17492), .dout(n17497));
  jor  g17244(.dina(n17497), .dinb(n17491), .dout(n17498));
  jand g17245(.dina(n17498), .dinb(asqrt[61] ), .dout(n17499));
  jor  g17246(.dina(n17498), .dinb(asqrt[61] ), .dout(n17500));
  jxor g17247(.dina(n16845), .dinb(n294), .dout(n17501));
  jand g17248(.dina(n17501), .dinb(asqrt[12] ), .dout(n17502));
  jxor g17249(.dina(n17502), .dinb(n16850), .dout(n17503));
  jand g17250(.dina(n17503), .dinb(n17500), .dout(n17504));
  jor  g17251(.dina(n17504), .dinb(n17499), .dout(n17505));
  jand g17252(.dina(n17505), .dinb(asqrt[62] ), .dout(n17506));
  jor  g17253(.dina(n17505), .dinb(asqrt[62] ), .dout(n17507));
  jxor g17254(.dina(n16853), .dinb(n239), .dout(n17508));
  jand g17255(.dina(n17508), .dinb(asqrt[12] ), .dout(n17509));
  jxor g17256(.dina(n17509), .dinb(n16858), .dout(n17510));
  jnot g17257(.din(n17510), .dout(n17511));
  jand g17258(.dina(n17511), .dinb(n17507), .dout(n17512));
  jor  g17259(.dina(n17512), .dinb(n17506), .dout(n17513));
  jxor g17260(.dina(n16860), .dinb(n221), .dout(n17514));
  jand g17261(.dina(n17514), .dinb(asqrt[12] ), .dout(n17515));
  jxor g17262(.dina(n17515), .dinb(n16866), .dout(n17516));
  jnot g17263(.din(n17516), .dout(n17517));
  jor  g17264(.dina(n17517), .dinb(n17513), .dout(n17518));
  jnot g17265(.din(n17518), .dout(n17519));
  jand g17266(.dina(n17132), .dinb(n16868), .dout(n17520));
  jnot g17267(.din(n17520), .dout(n17521));
  jand g17268(.dina(n16871), .dinb(asqrt[63] ), .dout(n17522));
  jand g17269(.dina(n17522), .dinb(n16896), .dout(n17523));
  jand g17270(.dina(n17523), .dinb(n17521), .dout(n17524));
  jand g17271(.dina(n16882), .dinb(n17127), .dout(n17525));
  jnot g17272(.din(n17506), .dout(n17526));
  jnot g17273(.din(n17499), .dout(n17527));
  jnot g17274(.din(n17491), .dout(n17528));
  jnot g17275(.din(n17484), .dout(n17529));
  jnot g17276(.din(n17476), .dout(n17530));
  jnot g17277(.din(n17468), .dout(n17531));
  jnot g17278(.din(n17460), .dout(n17532));
  jnot g17279(.din(n17453), .dout(n17533));
  jnot g17280(.din(n17445), .dout(n17534));
  jnot g17281(.din(n17438), .dout(n17535));
  jnot g17282(.din(n17430), .dout(n17536));
  jnot g17283(.din(n17423), .dout(n17537));
  jnot g17284(.din(n17426), .dout(n17538));
  jnot g17285(.din(n17416), .dout(n17539));
  jnot g17286(.din(n17408), .dout(n17540));
  jnot g17287(.din(n17400), .dout(n17541));
  jnot g17288(.din(n17393), .dout(n17542));
  jnot g17289(.din(n17385), .dout(n17543));
  jnot g17290(.din(n17378), .dout(n17544));
  jnot g17291(.din(n17370), .dout(n17545));
  jnot g17292(.din(n17362), .dout(n17546));
  jnot g17293(.din(n17354), .dout(n17547));
  jnot g17294(.din(n17347), .dout(n17548));
  jnot g17295(.din(n17339), .dout(n17549));
  jnot g17296(.din(n17332), .dout(n17550));
  jnot g17297(.din(n17324), .dout(n17551));
  jnot g17298(.din(n17316), .dout(n17552));
  jnot g17299(.din(n17308), .dout(n17553));
  jnot g17300(.din(n17301), .dout(n17554));
  jnot g17301(.din(n17293), .dout(n17555));
  jnot g17302(.din(n17286), .dout(n17556));
  jnot g17303(.din(n17278), .dout(n17557));
  jnot g17304(.din(n17271), .dout(n17558));
  jnot g17305(.din(n17263), .dout(n17559));
  jnot g17306(.din(n17256), .dout(n17560));
  jnot g17307(.din(n17248), .dout(n17561));
  jnot g17308(.din(n17240), .dout(n17562));
  jnot g17309(.din(n17232), .dout(n17563));
  jnot g17310(.din(n17225), .dout(n17564));
  jnot g17311(.din(n17217), .dout(n17565));
  jnot g17312(.din(n17210), .dout(n17566));
  jnot g17313(.din(n17202), .dout(n17567));
  jnot g17314(.din(n17195), .dout(n17568));
  jnot g17315(.din(n17188), .dout(n17569));
  jnot g17316(.din(n17180), .dout(n17570));
  jnot g17317(.din(n17172), .dout(n17571));
  jnot g17318(.din(n17165), .dout(n17572));
  jnot g17319(.din(n17157), .dout(n17573));
  jnot g17320(.din(n17150), .dout(n17574));
  jnot g17321(.din(n17139), .dout(n17575));
  jnot g17322(.din(n16891), .dout(n17576));
  jnot g17323(.din(n16888), .dout(n17577));
  jor  g17324(.dina(n17134), .dinb(n16494), .dout(n17578));
  jand g17325(.dina(n17578), .dinb(n17577), .dout(n17579));
  jand g17326(.dina(n17579), .dinb(n16489), .dout(n17580));
  jor  g17327(.dina(n17134), .dinb(a[24] ), .dout(n17581));
  jand g17328(.dina(n17581), .dinb(a[25] ), .dout(n17582));
  jor  g17329(.dina(n17141), .dinb(n17582), .dout(n17583));
  jor  g17330(.dina(n17583), .dinb(n17580), .dout(n17584));
  jand g17331(.dina(n17584), .dinb(n17576), .dout(n17585));
  jand g17332(.dina(n17585), .dinb(n15878), .dout(n17586));
  jor  g17333(.dina(n17146), .dinb(n17586), .dout(n17587));
  jand g17334(.dina(n17587), .dinb(n17575), .dout(n17588));
  jand g17335(.dina(n17588), .dinb(n15260), .dout(n17589));
  jnot g17336(.din(n17154), .dout(n17590));
  jor  g17337(.dina(n17590), .dinb(n17589), .dout(n17591));
  jand g17338(.dina(n17591), .dinb(n17574), .dout(n17592));
  jand g17339(.dina(n17592), .dinb(n14674), .dout(n17593));
  jor  g17340(.dina(n17161), .dinb(n17593), .dout(n17594));
  jand g17341(.dina(n17594), .dinb(n17573), .dout(n17595));
  jand g17342(.dina(n17595), .dinb(n14078), .dout(n17596));
  jnot g17343(.din(n17169), .dout(n17597));
  jor  g17344(.dina(n17597), .dinb(n17596), .dout(n17598));
  jand g17345(.dina(n17598), .dinb(n17572), .dout(n17599));
  jand g17346(.dina(n17599), .dinb(n13515), .dout(n17600));
  jor  g17347(.dina(n17176), .dinb(n17600), .dout(n17601));
  jand g17348(.dina(n17601), .dinb(n17571), .dout(n17602));
  jand g17349(.dina(n17602), .dinb(n12947), .dout(n17603));
  jor  g17350(.dina(n17184), .dinb(n17603), .dout(n17604));
  jand g17351(.dina(n17604), .dinb(n17570), .dout(n17605));
  jand g17352(.dina(n17605), .dinb(n12410), .dout(n17606));
  jnot g17353(.din(n17192), .dout(n17607));
  jor  g17354(.dina(n17607), .dinb(n17606), .dout(n17608));
  jand g17355(.dina(n17608), .dinb(n17569), .dout(n17609));
  jand g17356(.dina(n17609), .dinb(n11858), .dout(n17610));
  jnot g17357(.din(n17199), .dout(n17611));
  jor  g17358(.dina(n17611), .dinb(n17610), .dout(n17612));
  jand g17359(.dina(n17612), .dinb(n17568), .dout(n17613));
  jand g17360(.dina(n17613), .dinb(n11347), .dout(n17614));
  jor  g17361(.dina(n17206), .dinb(n17614), .dout(n17615));
  jand g17362(.dina(n17615), .dinb(n17567), .dout(n17616));
  jand g17363(.dina(n17616), .dinb(n10824), .dout(n17617));
  jnot g17364(.din(n17214), .dout(n17618));
  jor  g17365(.dina(n17618), .dinb(n17617), .dout(n17619));
  jand g17366(.dina(n17619), .dinb(n17566), .dout(n17620));
  jand g17367(.dina(n17620), .dinb(n10328), .dout(n17621));
  jor  g17368(.dina(n17221), .dinb(n17621), .dout(n17622));
  jand g17369(.dina(n17622), .dinb(n17565), .dout(n17623));
  jand g17370(.dina(n17623), .dinb(n9832), .dout(n17624));
  jnot g17371(.din(n17229), .dout(n17625));
  jor  g17372(.dina(n17625), .dinb(n17624), .dout(n17626));
  jand g17373(.dina(n17626), .dinb(n17564), .dout(n17627));
  jand g17374(.dina(n17627), .dinb(n9369), .dout(n17628));
  jor  g17375(.dina(n17236), .dinb(n17628), .dout(n17629));
  jand g17376(.dina(n17629), .dinb(n17563), .dout(n17630));
  jand g17377(.dina(n17630), .dinb(n8890), .dout(n17631));
  jor  g17378(.dina(n17244), .dinb(n17631), .dout(n17632));
  jand g17379(.dina(n17632), .dinb(n17562), .dout(n17633));
  jand g17380(.dina(n17633), .dinb(n8449), .dout(n17634));
  jor  g17381(.dina(n17252), .dinb(n17634), .dout(n17635));
  jand g17382(.dina(n17635), .dinb(n17561), .dout(n17636));
  jand g17383(.dina(n17636), .dinb(n8003), .dout(n17637));
  jnot g17384(.din(n17260), .dout(n17638));
  jor  g17385(.dina(n17638), .dinb(n17637), .dout(n17639));
  jand g17386(.dina(n17639), .dinb(n17560), .dout(n17640));
  jand g17387(.dina(n17640), .dinb(n7581), .dout(n17641));
  jor  g17388(.dina(n17267), .dinb(n17641), .dout(n17642));
  jand g17389(.dina(n17642), .dinb(n17559), .dout(n17643));
  jand g17390(.dina(n17643), .dinb(n7154), .dout(n17644));
  jnot g17391(.din(n17275), .dout(n17645));
  jor  g17392(.dina(n17645), .dinb(n17644), .dout(n17646));
  jand g17393(.dina(n17646), .dinb(n17558), .dout(n17647));
  jand g17394(.dina(n17647), .dinb(n6758), .dout(n17648));
  jor  g17395(.dina(n17282), .dinb(n17648), .dout(n17649));
  jand g17396(.dina(n17649), .dinb(n17557), .dout(n17650));
  jand g17397(.dina(n17650), .dinb(n6357), .dout(n17651));
  jnot g17398(.din(n17290), .dout(n17652));
  jor  g17399(.dina(n17652), .dinb(n17651), .dout(n17653));
  jand g17400(.dina(n17653), .dinb(n17556), .dout(n17654));
  jand g17401(.dina(n17654), .dinb(n5989), .dout(n17655));
  jor  g17402(.dina(n17297), .dinb(n17655), .dout(n17656));
  jand g17403(.dina(n17656), .dinb(n17555), .dout(n17657));
  jand g17404(.dina(n17657), .dinb(n5606), .dout(n17658));
  jnot g17405(.din(n17305), .dout(n17659));
  jor  g17406(.dina(n17659), .dinb(n17658), .dout(n17660));
  jand g17407(.dina(n17660), .dinb(n17554), .dout(n17661));
  jand g17408(.dina(n17661), .dinb(n5259), .dout(n17662));
  jor  g17409(.dina(n17312), .dinb(n17662), .dout(n17663));
  jand g17410(.dina(n17663), .dinb(n17553), .dout(n17664));
  jand g17411(.dina(n17664), .dinb(n4902), .dout(n17665));
  jor  g17412(.dina(n17320), .dinb(n17665), .dout(n17666));
  jand g17413(.dina(n17666), .dinb(n17552), .dout(n17667));
  jand g17414(.dina(n17667), .dinb(n4582), .dout(n17668));
  jor  g17415(.dina(n17328), .dinb(n17668), .dout(n17669));
  jand g17416(.dina(n17669), .dinb(n17551), .dout(n17670));
  jand g17417(.dina(n17670), .dinb(n4249), .dout(n17671));
  jnot g17418(.din(n17336), .dout(n17672));
  jor  g17419(.dina(n17672), .dinb(n17671), .dout(n17673));
  jand g17420(.dina(n17673), .dinb(n17550), .dout(n17674));
  jand g17421(.dina(n17674), .dinb(n3955), .dout(n17675));
  jor  g17422(.dina(n17343), .dinb(n17675), .dout(n17676));
  jand g17423(.dina(n17676), .dinb(n17549), .dout(n17677));
  jand g17424(.dina(n17677), .dinb(n3642), .dout(n17678));
  jnot g17425(.din(n17351), .dout(n17679));
  jor  g17426(.dina(n17679), .dinb(n17678), .dout(n17680));
  jand g17427(.dina(n17680), .dinb(n17548), .dout(n17681));
  jand g17428(.dina(n17681), .dinb(n3368), .dout(n17682));
  jor  g17429(.dina(n17358), .dinb(n17682), .dout(n17683));
  jand g17430(.dina(n17683), .dinb(n17547), .dout(n17684));
  jand g17431(.dina(n17684), .dinb(n3089), .dout(n17685));
  jor  g17432(.dina(n17366), .dinb(n17685), .dout(n17686));
  jand g17433(.dina(n17686), .dinb(n17546), .dout(n17687));
  jand g17434(.dina(n17687), .dinb(n2833), .dout(n17688));
  jor  g17435(.dina(n17374), .dinb(n17688), .dout(n17689));
  jand g17436(.dina(n17689), .dinb(n17545), .dout(n17690));
  jand g17437(.dina(n17690), .dinb(n2572), .dout(n17691));
  jnot g17438(.din(n17382), .dout(n17692));
  jor  g17439(.dina(n17692), .dinb(n17691), .dout(n17693));
  jand g17440(.dina(n17693), .dinb(n17544), .dout(n17694));
  jand g17441(.dina(n17694), .dinb(n2345), .dout(n17695));
  jor  g17442(.dina(n17389), .dinb(n17695), .dout(n17696));
  jand g17443(.dina(n17696), .dinb(n17543), .dout(n17697));
  jand g17444(.dina(n17697), .dinb(n2108), .dout(n17698));
  jnot g17445(.din(n17397), .dout(n17699));
  jor  g17446(.dina(n17699), .dinb(n17698), .dout(n17700));
  jand g17447(.dina(n17700), .dinb(n17542), .dout(n17701));
  jand g17448(.dina(n17701), .dinb(n1912), .dout(n17702));
  jor  g17449(.dina(n17404), .dinb(n17702), .dout(n17703));
  jand g17450(.dina(n17703), .dinb(n17541), .dout(n17704));
  jand g17451(.dina(n17704), .dinb(n1699), .dout(n17705));
  jor  g17452(.dina(n17412), .dinb(n17705), .dout(n17706));
  jand g17453(.dina(n17706), .dinb(n17540), .dout(n17707));
  jand g17454(.dina(n17707), .dinb(n1516), .dout(n17708));
  jnot g17455(.din(n17420), .dout(n17709));
  jor  g17456(.dina(n17709), .dinb(n17708), .dout(n17710));
  jand g17457(.dina(n17710), .dinb(n17539), .dout(n17711));
  jand g17458(.dina(n17711), .dinb(n1332), .dout(n17712));
  jor  g17459(.dina(n17712), .dinb(n17538), .dout(n17713));
  jand g17460(.dina(n17713), .dinb(n17537), .dout(n17714));
  jand g17461(.dina(n17714), .dinb(n1173), .dout(n17715));
  jor  g17462(.dina(n17434), .dinb(n17715), .dout(n17716));
  jand g17463(.dina(n17716), .dinb(n17536), .dout(n17717));
  jand g17464(.dina(n17717), .dinb(n1008), .dout(n17718));
  jnot g17465(.din(n17442), .dout(n17719));
  jor  g17466(.dina(n17719), .dinb(n17718), .dout(n17720));
  jand g17467(.dina(n17720), .dinb(n17535), .dout(n17721));
  jand g17468(.dina(n17721), .dinb(n884), .dout(n17722));
  jor  g17469(.dina(n17449), .dinb(n17722), .dout(n17723));
  jand g17470(.dina(n17723), .dinb(n17534), .dout(n17724));
  jand g17471(.dina(n17724), .dinb(n743), .dout(n17725));
  jnot g17472(.din(n17457), .dout(n17726));
  jor  g17473(.dina(n17726), .dinb(n17725), .dout(n17727));
  jand g17474(.dina(n17727), .dinb(n17533), .dout(n17728));
  jand g17475(.dina(n17728), .dinb(n635), .dout(n17729));
  jor  g17476(.dina(n17464), .dinb(n17729), .dout(n17730));
  jand g17477(.dina(n17730), .dinb(n17532), .dout(n17731));
  jand g17478(.dina(n17731), .dinb(n515), .dout(n17732));
  jor  g17479(.dina(n17472), .dinb(n17732), .dout(n17733));
  jand g17480(.dina(n17733), .dinb(n17531), .dout(n17734));
  jand g17481(.dina(n17734), .dinb(n443), .dout(n17735));
  jor  g17482(.dina(n17480), .dinb(n17735), .dout(n17736));
  jand g17483(.dina(n17736), .dinb(n17530), .dout(n17737));
  jand g17484(.dina(n17737), .dinb(n352), .dout(n17738));
  jnot g17485(.din(n17488), .dout(n17739));
  jor  g17486(.dina(n17739), .dinb(n17738), .dout(n17740));
  jand g17487(.dina(n17740), .dinb(n17529), .dout(n17741));
  jand g17488(.dina(n17741), .dinb(n294), .dout(n17742));
  jor  g17489(.dina(n17495), .dinb(n17742), .dout(n17743));
  jand g17490(.dina(n17743), .dinb(n17528), .dout(n17744));
  jand g17491(.dina(n17744), .dinb(n239), .dout(n17745));
  jnot g17492(.din(n17503), .dout(n17746));
  jor  g17493(.dina(n17746), .dinb(n17745), .dout(n17747));
  jand g17494(.dina(n17747), .dinb(n17527), .dout(n17748));
  jand g17495(.dina(n17748), .dinb(n221), .dout(n17749));
  jor  g17496(.dina(n17510), .dinb(n17749), .dout(n17750));
  jand g17497(.dina(n17750), .dinb(n17526), .dout(n17751));
  jor  g17498(.dina(n17516), .dinb(n17751), .dout(n17752));
  jor  g17499(.dina(n17752), .dinb(n16869), .dout(n17753));
  jor  g17500(.dina(n17753), .dinb(n17525), .dout(n17754));
  jand g17501(.dina(n17754), .dinb(n218), .dout(n17755));
  jand g17502(.dina(n17134), .dinb(n16493), .dout(n17756));
  jor  g17503(.dina(n17756), .dinb(n17755), .dout(n17757));
  jor  g17504(.dina(n17757), .dinb(n17524), .dout(n17758));
  jor  g17505(.dina(n17758), .dinb(n17519), .dout(asqrt[11] ));
  jnot g17506(.din(n17524), .dout(n17760));
  jnot g17507(.din(n17525), .dout(n17761));
  jand g17508(.dina(n17517), .dinb(n17513), .dout(n17762));
  jand g17509(.dina(n17762), .dinb(n16896), .dout(n17763));
  jand g17510(.dina(n17763), .dinb(n17761), .dout(n17764));
  jor  g17511(.dina(n17764), .dinb(asqrt[63] ), .dout(n17765));
  jnot g17512(.din(n17756), .dout(n17766));
  jand g17513(.dina(n17766), .dinb(n17765), .dout(n17767));
  jand g17514(.dina(n17767), .dinb(n17760), .dout(n17768));
  jand g17515(.dina(n17768), .dinb(n17518), .dout(n17769));
  jxor g17516(.dina(n17505), .dinb(n221), .dout(n17770));
  jor  g17517(.dina(n17770), .dinb(n17769), .dout(n17771));
  jxor g17518(.dina(n17771), .dinb(n17510), .dout(n17772));
  jnot g17519(.din(n17772), .dout(n17773));
  jnot g17520(.din(a[20] ), .dout(n17774));
  jnot g17521(.din(a[21] ), .dout(n17775));
  jand g17522(.dina(n17775), .dinb(n17774), .dout(n17776));
  jand g17523(.dina(n17776), .dinb(n16885), .dout(n17777));
  jnot g17524(.din(n17777), .dout(n17778));
  jor  g17525(.dina(n17769), .dinb(n16885), .dout(n17779));
  jand g17526(.dina(n17779), .dinb(n17778), .dout(n17780));
  jor  g17527(.dina(n17780), .dinb(n17134), .dout(n17781));
  jand g17528(.dina(n17780), .dinb(n17134), .dout(n17782));
  jor  g17529(.dina(n17769), .dinb(a[22] ), .dout(n17783));
  jand g17530(.dina(n17783), .dinb(a[23] ), .dout(n17784));
  jand g17531(.dina(asqrt[11] ), .dinb(n16887), .dout(n17785));
  jor  g17532(.dina(n17785), .dinb(n17784), .dout(n17786));
  jor  g17533(.dina(n17786), .dinb(n17782), .dout(n17787));
  jand g17534(.dina(n17787), .dinb(n17781), .dout(n17788));
  jor  g17535(.dina(n17788), .dinb(n16489), .dout(n17789));
  jand g17536(.dina(n17788), .dinb(n16489), .dout(n17790));
  jnot g17537(.din(n16887), .dout(n17791));
  jor  g17538(.dina(n17769), .dinb(n17791), .dout(n17792));
  jor  g17539(.dina(n17519), .dinb(n17134), .dout(n17793));
  jor  g17540(.dina(n17793), .dinb(n17523), .dout(n17794));
  jor  g17541(.dina(n17794), .dinb(n17755), .dout(n17795));
  jand g17542(.dina(n17795), .dinb(n17792), .dout(n17796));
  jxor g17543(.dina(n17796), .dinb(n16494), .dout(n17797));
  jor  g17544(.dina(n17797), .dinb(n17790), .dout(n17798));
  jand g17545(.dina(n17798), .dinb(n17789), .dout(n17799));
  jor  g17546(.dina(n17799), .dinb(n15878), .dout(n17800));
  jand g17547(.dina(n17799), .dinb(n15878), .dout(n17801));
  jxor g17548(.dina(n16890), .dinb(n16489), .dout(n17802));
  jor  g17549(.dina(n17802), .dinb(n17769), .dout(n17803));
  jxor g17550(.dina(n17803), .dinb(n17583), .dout(n17804));
  jnot g17551(.din(n17804), .dout(n17805));
  jor  g17552(.dina(n17805), .dinb(n17801), .dout(n17806));
  jand g17553(.dina(n17806), .dinb(n17800), .dout(n17807));
  jor  g17554(.dina(n17807), .dinb(n15260), .dout(n17808));
  jand g17555(.dina(n17807), .dinb(n15260), .dout(n17809));
  jxor g17556(.dina(n17138), .dinb(n15878), .dout(n17810));
  jor  g17557(.dina(n17810), .dinb(n17769), .dout(n17811));
  jxor g17558(.dina(n17811), .dinb(n17147), .dout(n17812));
  jor  g17559(.dina(n17812), .dinb(n17809), .dout(n17813));
  jand g17560(.dina(n17813), .dinb(n17808), .dout(n17814));
  jor  g17561(.dina(n17814), .dinb(n14674), .dout(n17815));
  jand g17562(.dina(n17814), .dinb(n14674), .dout(n17816));
  jxor g17563(.dina(n17149), .dinb(n15260), .dout(n17817));
  jor  g17564(.dina(n17817), .dinb(n17769), .dout(n17818));
  jxor g17565(.dina(n17818), .dinb(n17590), .dout(n17819));
  jnot g17566(.din(n17819), .dout(n17820));
  jor  g17567(.dina(n17820), .dinb(n17816), .dout(n17821));
  jand g17568(.dina(n17821), .dinb(n17815), .dout(n17822));
  jor  g17569(.dina(n17822), .dinb(n14078), .dout(n17823));
  jand g17570(.dina(n17822), .dinb(n14078), .dout(n17824));
  jxor g17571(.dina(n17156), .dinb(n14674), .dout(n17825));
  jor  g17572(.dina(n17825), .dinb(n17769), .dout(n17826));
  jxor g17573(.dina(n17826), .dinb(n17162), .dout(n17827));
  jor  g17574(.dina(n17827), .dinb(n17824), .dout(n17828));
  jand g17575(.dina(n17828), .dinb(n17823), .dout(n17829));
  jor  g17576(.dina(n17829), .dinb(n13515), .dout(n17830));
  jand g17577(.dina(n17829), .dinb(n13515), .dout(n17831));
  jxor g17578(.dina(n17164), .dinb(n14078), .dout(n17832));
  jor  g17579(.dina(n17832), .dinb(n17769), .dout(n17833));
  jxor g17580(.dina(n17833), .dinb(n17597), .dout(n17834));
  jnot g17581(.din(n17834), .dout(n17835));
  jor  g17582(.dina(n17835), .dinb(n17831), .dout(n17836));
  jand g17583(.dina(n17836), .dinb(n17830), .dout(n17837));
  jor  g17584(.dina(n17837), .dinb(n12947), .dout(n17838));
  jand g17585(.dina(n17837), .dinb(n12947), .dout(n17839));
  jxor g17586(.dina(n17171), .dinb(n13515), .dout(n17840));
  jor  g17587(.dina(n17840), .dinb(n17769), .dout(n17841));
  jxor g17588(.dina(n17841), .dinb(n17177), .dout(n17842));
  jor  g17589(.dina(n17842), .dinb(n17839), .dout(n17843));
  jand g17590(.dina(n17843), .dinb(n17838), .dout(n17844));
  jor  g17591(.dina(n17844), .dinb(n12410), .dout(n17845));
  jand g17592(.dina(n17844), .dinb(n12410), .dout(n17846));
  jxor g17593(.dina(n17179), .dinb(n12947), .dout(n17847));
  jor  g17594(.dina(n17847), .dinb(n17769), .dout(n17848));
  jxor g17595(.dina(n17848), .dinb(n17185), .dout(n17849));
  jor  g17596(.dina(n17849), .dinb(n17846), .dout(n17850));
  jand g17597(.dina(n17850), .dinb(n17845), .dout(n17851));
  jor  g17598(.dina(n17851), .dinb(n11858), .dout(n17852));
  jand g17599(.dina(n17851), .dinb(n11858), .dout(n17853));
  jxor g17600(.dina(n17187), .dinb(n12410), .dout(n17854));
  jor  g17601(.dina(n17854), .dinb(n17769), .dout(n17855));
  jxor g17602(.dina(n17855), .dinb(n17607), .dout(n17856));
  jnot g17603(.din(n17856), .dout(n17857));
  jor  g17604(.dina(n17857), .dinb(n17853), .dout(n17858));
  jand g17605(.dina(n17858), .dinb(n17852), .dout(n17859));
  jor  g17606(.dina(n17859), .dinb(n11347), .dout(n17860));
  jand g17607(.dina(n17859), .dinb(n11347), .dout(n17861));
  jxor g17608(.dina(n17194), .dinb(n11858), .dout(n17862));
  jor  g17609(.dina(n17862), .dinb(n17769), .dout(n17863));
  jxor g17610(.dina(n17863), .dinb(n17611), .dout(n17864));
  jnot g17611(.din(n17864), .dout(n17865));
  jor  g17612(.dina(n17865), .dinb(n17861), .dout(n17866));
  jand g17613(.dina(n17866), .dinb(n17860), .dout(n17867));
  jor  g17614(.dina(n17867), .dinb(n10824), .dout(n17868));
  jand g17615(.dina(n17867), .dinb(n10824), .dout(n17869));
  jxor g17616(.dina(n17201), .dinb(n11347), .dout(n17870));
  jor  g17617(.dina(n17870), .dinb(n17769), .dout(n17871));
  jxor g17618(.dina(n17871), .dinb(n17207), .dout(n17872));
  jor  g17619(.dina(n17872), .dinb(n17869), .dout(n17873));
  jand g17620(.dina(n17873), .dinb(n17868), .dout(n17874));
  jor  g17621(.dina(n17874), .dinb(n10328), .dout(n17875));
  jand g17622(.dina(n17874), .dinb(n10328), .dout(n17876));
  jxor g17623(.dina(n17209), .dinb(n10824), .dout(n17877));
  jor  g17624(.dina(n17877), .dinb(n17769), .dout(n17878));
  jxor g17625(.dina(n17878), .dinb(n17618), .dout(n17879));
  jnot g17626(.din(n17879), .dout(n17880));
  jor  g17627(.dina(n17880), .dinb(n17876), .dout(n17881));
  jand g17628(.dina(n17881), .dinb(n17875), .dout(n17882));
  jor  g17629(.dina(n17882), .dinb(n9832), .dout(n17883));
  jand g17630(.dina(n17882), .dinb(n9832), .dout(n17884));
  jxor g17631(.dina(n17216), .dinb(n10328), .dout(n17885));
  jor  g17632(.dina(n17885), .dinb(n17769), .dout(n17886));
  jxor g17633(.dina(n17886), .dinb(n17222), .dout(n17887));
  jor  g17634(.dina(n17887), .dinb(n17884), .dout(n17888));
  jand g17635(.dina(n17888), .dinb(n17883), .dout(n17889));
  jor  g17636(.dina(n17889), .dinb(n9369), .dout(n17890));
  jand g17637(.dina(n17889), .dinb(n9369), .dout(n17891));
  jxor g17638(.dina(n17224), .dinb(n9832), .dout(n17892));
  jor  g17639(.dina(n17892), .dinb(n17769), .dout(n17893));
  jxor g17640(.dina(n17893), .dinb(n17625), .dout(n17894));
  jnot g17641(.din(n17894), .dout(n17895));
  jor  g17642(.dina(n17895), .dinb(n17891), .dout(n17896));
  jand g17643(.dina(n17896), .dinb(n17890), .dout(n17897));
  jor  g17644(.dina(n17897), .dinb(n8890), .dout(n17898));
  jand g17645(.dina(n17897), .dinb(n8890), .dout(n17899));
  jxor g17646(.dina(n17231), .dinb(n9369), .dout(n17900));
  jor  g17647(.dina(n17900), .dinb(n17769), .dout(n17901));
  jxor g17648(.dina(n17901), .dinb(n17237), .dout(n17902));
  jor  g17649(.dina(n17902), .dinb(n17899), .dout(n17903));
  jand g17650(.dina(n17903), .dinb(n17898), .dout(n17904));
  jor  g17651(.dina(n17904), .dinb(n8449), .dout(n17905));
  jand g17652(.dina(n17904), .dinb(n8449), .dout(n17906));
  jxor g17653(.dina(n17239), .dinb(n8890), .dout(n17907));
  jor  g17654(.dina(n17907), .dinb(n17769), .dout(n17908));
  jxor g17655(.dina(n17908), .dinb(n17245), .dout(n17909));
  jor  g17656(.dina(n17909), .dinb(n17906), .dout(n17910));
  jand g17657(.dina(n17910), .dinb(n17905), .dout(n17911));
  jor  g17658(.dina(n17911), .dinb(n8003), .dout(n17912));
  jand g17659(.dina(n17911), .dinb(n8003), .dout(n17913));
  jxor g17660(.dina(n17247), .dinb(n8449), .dout(n17914));
  jor  g17661(.dina(n17914), .dinb(n17769), .dout(n17915));
  jxor g17662(.dina(n17915), .dinb(n17253), .dout(n17916));
  jor  g17663(.dina(n17916), .dinb(n17913), .dout(n17917));
  jand g17664(.dina(n17917), .dinb(n17912), .dout(n17918));
  jor  g17665(.dina(n17918), .dinb(n7581), .dout(n17919));
  jand g17666(.dina(n17918), .dinb(n7581), .dout(n17920));
  jxor g17667(.dina(n17255), .dinb(n8003), .dout(n17921));
  jor  g17668(.dina(n17921), .dinb(n17769), .dout(n17922));
  jxor g17669(.dina(n17922), .dinb(n17638), .dout(n17923));
  jnot g17670(.din(n17923), .dout(n17924));
  jor  g17671(.dina(n17924), .dinb(n17920), .dout(n17925));
  jand g17672(.dina(n17925), .dinb(n17919), .dout(n17926));
  jor  g17673(.dina(n17926), .dinb(n7154), .dout(n17927));
  jand g17674(.dina(n17926), .dinb(n7154), .dout(n17928));
  jxor g17675(.dina(n17262), .dinb(n7581), .dout(n17929));
  jor  g17676(.dina(n17929), .dinb(n17769), .dout(n17930));
  jxor g17677(.dina(n17930), .dinb(n17268), .dout(n17931));
  jor  g17678(.dina(n17931), .dinb(n17928), .dout(n17932));
  jand g17679(.dina(n17932), .dinb(n17927), .dout(n17933));
  jor  g17680(.dina(n17933), .dinb(n6758), .dout(n17934));
  jand g17681(.dina(n17933), .dinb(n6758), .dout(n17935));
  jxor g17682(.dina(n17270), .dinb(n7154), .dout(n17936));
  jor  g17683(.dina(n17936), .dinb(n17769), .dout(n17937));
  jxor g17684(.dina(n17937), .dinb(n17645), .dout(n17938));
  jnot g17685(.din(n17938), .dout(n17939));
  jor  g17686(.dina(n17939), .dinb(n17935), .dout(n17940));
  jand g17687(.dina(n17940), .dinb(n17934), .dout(n17941));
  jor  g17688(.dina(n17941), .dinb(n6357), .dout(n17942));
  jand g17689(.dina(n17941), .dinb(n6357), .dout(n17943));
  jxor g17690(.dina(n17277), .dinb(n6758), .dout(n17944));
  jor  g17691(.dina(n17944), .dinb(n17769), .dout(n17945));
  jxor g17692(.dina(n17945), .dinb(n17283), .dout(n17946));
  jor  g17693(.dina(n17946), .dinb(n17943), .dout(n17947));
  jand g17694(.dina(n17947), .dinb(n17942), .dout(n17948));
  jor  g17695(.dina(n17948), .dinb(n5989), .dout(n17949));
  jand g17696(.dina(n17948), .dinb(n5989), .dout(n17950));
  jxor g17697(.dina(n17285), .dinb(n6357), .dout(n17951));
  jor  g17698(.dina(n17951), .dinb(n17769), .dout(n17952));
  jxor g17699(.dina(n17952), .dinb(n17652), .dout(n17953));
  jnot g17700(.din(n17953), .dout(n17954));
  jor  g17701(.dina(n17954), .dinb(n17950), .dout(n17955));
  jand g17702(.dina(n17955), .dinb(n17949), .dout(n17956));
  jor  g17703(.dina(n17956), .dinb(n5606), .dout(n17957));
  jand g17704(.dina(n17956), .dinb(n5606), .dout(n17958));
  jxor g17705(.dina(n17292), .dinb(n5989), .dout(n17959));
  jor  g17706(.dina(n17959), .dinb(n17769), .dout(n17960));
  jxor g17707(.dina(n17960), .dinb(n17298), .dout(n17961));
  jor  g17708(.dina(n17961), .dinb(n17958), .dout(n17962));
  jand g17709(.dina(n17962), .dinb(n17957), .dout(n17963));
  jor  g17710(.dina(n17963), .dinb(n5259), .dout(n17964));
  jand g17711(.dina(n17963), .dinb(n5259), .dout(n17965));
  jxor g17712(.dina(n17300), .dinb(n5606), .dout(n17966));
  jor  g17713(.dina(n17966), .dinb(n17769), .dout(n17967));
  jxor g17714(.dina(n17967), .dinb(n17659), .dout(n17968));
  jnot g17715(.din(n17968), .dout(n17969));
  jor  g17716(.dina(n17969), .dinb(n17965), .dout(n17970));
  jand g17717(.dina(n17970), .dinb(n17964), .dout(n17971));
  jor  g17718(.dina(n17971), .dinb(n4902), .dout(n17972));
  jand g17719(.dina(n17971), .dinb(n4902), .dout(n17973));
  jxor g17720(.dina(n17307), .dinb(n5259), .dout(n17974));
  jor  g17721(.dina(n17974), .dinb(n17769), .dout(n17975));
  jxor g17722(.dina(n17975), .dinb(n17313), .dout(n17976));
  jor  g17723(.dina(n17976), .dinb(n17973), .dout(n17977));
  jand g17724(.dina(n17977), .dinb(n17972), .dout(n17978));
  jor  g17725(.dina(n17978), .dinb(n4582), .dout(n17979));
  jand g17726(.dina(n17978), .dinb(n4582), .dout(n17980));
  jxor g17727(.dina(n17315), .dinb(n4902), .dout(n17981));
  jor  g17728(.dina(n17981), .dinb(n17769), .dout(n17982));
  jxor g17729(.dina(n17982), .dinb(n17321), .dout(n17983));
  jor  g17730(.dina(n17983), .dinb(n17980), .dout(n17984));
  jand g17731(.dina(n17984), .dinb(n17979), .dout(n17985));
  jor  g17732(.dina(n17985), .dinb(n4249), .dout(n17986));
  jand g17733(.dina(n17985), .dinb(n4249), .dout(n17987));
  jxor g17734(.dina(n17323), .dinb(n4582), .dout(n17988));
  jor  g17735(.dina(n17988), .dinb(n17769), .dout(n17989));
  jxor g17736(.dina(n17989), .dinb(n17329), .dout(n17990));
  jor  g17737(.dina(n17990), .dinb(n17987), .dout(n17991));
  jand g17738(.dina(n17991), .dinb(n17986), .dout(n17992));
  jor  g17739(.dina(n17992), .dinb(n3955), .dout(n17993));
  jand g17740(.dina(n17992), .dinb(n3955), .dout(n17994));
  jxor g17741(.dina(n17331), .dinb(n4249), .dout(n17995));
  jor  g17742(.dina(n17995), .dinb(n17769), .dout(n17996));
  jxor g17743(.dina(n17996), .dinb(n17672), .dout(n17997));
  jnot g17744(.din(n17997), .dout(n17998));
  jor  g17745(.dina(n17998), .dinb(n17994), .dout(n17999));
  jand g17746(.dina(n17999), .dinb(n17993), .dout(n18000));
  jor  g17747(.dina(n18000), .dinb(n3642), .dout(n18001));
  jand g17748(.dina(n18000), .dinb(n3642), .dout(n18002));
  jxor g17749(.dina(n17338), .dinb(n3955), .dout(n18003));
  jor  g17750(.dina(n18003), .dinb(n17769), .dout(n18004));
  jxor g17751(.dina(n18004), .dinb(n17344), .dout(n18005));
  jor  g17752(.dina(n18005), .dinb(n18002), .dout(n18006));
  jand g17753(.dina(n18006), .dinb(n18001), .dout(n18007));
  jor  g17754(.dina(n18007), .dinb(n3368), .dout(n18008));
  jand g17755(.dina(n18007), .dinb(n3368), .dout(n18009));
  jxor g17756(.dina(n17346), .dinb(n3642), .dout(n18010));
  jor  g17757(.dina(n18010), .dinb(n17769), .dout(n18011));
  jxor g17758(.dina(n18011), .dinb(n17679), .dout(n18012));
  jnot g17759(.din(n18012), .dout(n18013));
  jor  g17760(.dina(n18013), .dinb(n18009), .dout(n18014));
  jand g17761(.dina(n18014), .dinb(n18008), .dout(n18015));
  jor  g17762(.dina(n18015), .dinb(n3089), .dout(n18016));
  jand g17763(.dina(n18015), .dinb(n3089), .dout(n18017));
  jxor g17764(.dina(n17353), .dinb(n3368), .dout(n18018));
  jor  g17765(.dina(n18018), .dinb(n17769), .dout(n18019));
  jxor g17766(.dina(n18019), .dinb(n17359), .dout(n18020));
  jor  g17767(.dina(n18020), .dinb(n18017), .dout(n18021));
  jand g17768(.dina(n18021), .dinb(n18016), .dout(n18022));
  jor  g17769(.dina(n18022), .dinb(n2833), .dout(n18023));
  jand g17770(.dina(n18022), .dinb(n2833), .dout(n18024));
  jxor g17771(.dina(n17361), .dinb(n3089), .dout(n18025));
  jor  g17772(.dina(n18025), .dinb(n17769), .dout(n18026));
  jxor g17773(.dina(n18026), .dinb(n17367), .dout(n18027));
  jor  g17774(.dina(n18027), .dinb(n18024), .dout(n18028));
  jand g17775(.dina(n18028), .dinb(n18023), .dout(n18029));
  jor  g17776(.dina(n18029), .dinb(n2572), .dout(n18030));
  jand g17777(.dina(n18029), .dinb(n2572), .dout(n18031));
  jxor g17778(.dina(n17369), .dinb(n2833), .dout(n18032));
  jor  g17779(.dina(n18032), .dinb(n17769), .dout(n18033));
  jxor g17780(.dina(n18033), .dinb(n17375), .dout(n18034));
  jor  g17781(.dina(n18034), .dinb(n18031), .dout(n18035));
  jand g17782(.dina(n18035), .dinb(n18030), .dout(n18036));
  jor  g17783(.dina(n18036), .dinb(n2345), .dout(n18037));
  jand g17784(.dina(n18036), .dinb(n2345), .dout(n18038));
  jxor g17785(.dina(n17377), .dinb(n2572), .dout(n18039));
  jor  g17786(.dina(n18039), .dinb(n17769), .dout(n18040));
  jxor g17787(.dina(n18040), .dinb(n17692), .dout(n18041));
  jnot g17788(.din(n18041), .dout(n18042));
  jor  g17789(.dina(n18042), .dinb(n18038), .dout(n18043));
  jand g17790(.dina(n18043), .dinb(n18037), .dout(n18044));
  jor  g17791(.dina(n18044), .dinb(n2108), .dout(n18045));
  jand g17792(.dina(n18044), .dinb(n2108), .dout(n18046));
  jxor g17793(.dina(n17384), .dinb(n2345), .dout(n18047));
  jor  g17794(.dina(n18047), .dinb(n17769), .dout(n18048));
  jxor g17795(.dina(n18048), .dinb(n17390), .dout(n18049));
  jor  g17796(.dina(n18049), .dinb(n18046), .dout(n18050));
  jand g17797(.dina(n18050), .dinb(n18045), .dout(n18051));
  jor  g17798(.dina(n18051), .dinb(n1912), .dout(n18052));
  jand g17799(.dina(n18051), .dinb(n1912), .dout(n18053));
  jxor g17800(.dina(n17392), .dinb(n2108), .dout(n18054));
  jor  g17801(.dina(n18054), .dinb(n17769), .dout(n18055));
  jxor g17802(.dina(n18055), .dinb(n17699), .dout(n18056));
  jnot g17803(.din(n18056), .dout(n18057));
  jor  g17804(.dina(n18057), .dinb(n18053), .dout(n18058));
  jand g17805(.dina(n18058), .dinb(n18052), .dout(n18059));
  jor  g17806(.dina(n18059), .dinb(n1699), .dout(n18060));
  jand g17807(.dina(n18059), .dinb(n1699), .dout(n18061));
  jxor g17808(.dina(n17399), .dinb(n1912), .dout(n18062));
  jor  g17809(.dina(n18062), .dinb(n17769), .dout(n18063));
  jxor g17810(.dina(n18063), .dinb(n17405), .dout(n18064));
  jor  g17811(.dina(n18064), .dinb(n18061), .dout(n18065));
  jand g17812(.dina(n18065), .dinb(n18060), .dout(n18066));
  jor  g17813(.dina(n18066), .dinb(n1516), .dout(n18067));
  jand g17814(.dina(n18066), .dinb(n1516), .dout(n18068));
  jxor g17815(.dina(n17407), .dinb(n1699), .dout(n18069));
  jor  g17816(.dina(n18069), .dinb(n17769), .dout(n18070));
  jxor g17817(.dina(n18070), .dinb(n17413), .dout(n18071));
  jor  g17818(.dina(n18071), .dinb(n18068), .dout(n18072));
  jand g17819(.dina(n18072), .dinb(n18067), .dout(n18073));
  jor  g17820(.dina(n18073), .dinb(n1332), .dout(n18074));
  jand g17821(.dina(n18073), .dinb(n1332), .dout(n18075));
  jxor g17822(.dina(n17415), .dinb(n1516), .dout(n18076));
  jor  g17823(.dina(n18076), .dinb(n17769), .dout(n18077));
  jxor g17824(.dina(n18077), .dinb(n17709), .dout(n18078));
  jnot g17825(.din(n18078), .dout(n18079));
  jor  g17826(.dina(n18079), .dinb(n18075), .dout(n18080));
  jand g17827(.dina(n18080), .dinb(n18074), .dout(n18081));
  jor  g17828(.dina(n18081), .dinb(n1173), .dout(n18082));
  jxor g17829(.dina(n17422), .dinb(n1332), .dout(n18083));
  jor  g17830(.dina(n18083), .dinb(n17769), .dout(n18084));
  jxor g17831(.dina(n18084), .dinb(n17538), .dout(n18085));
  jnot g17832(.din(n18085), .dout(n18086));
  jand g17833(.dina(n18081), .dinb(n1173), .dout(n18087));
  jor  g17834(.dina(n18087), .dinb(n18086), .dout(n18088));
  jand g17835(.dina(n18088), .dinb(n18082), .dout(n18089));
  jor  g17836(.dina(n18089), .dinb(n1008), .dout(n18090));
  jand g17837(.dina(n18089), .dinb(n1008), .dout(n18091));
  jxor g17838(.dina(n17429), .dinb(n1173), .dout(n18092));
  jor  g17839(.dina(n18092), .dinb(n17769), .dout(n18093));
  jxor g17840(.dina(n18093), .dinb(n17435), .dout(n18094));
  jor  g17841(.dina(n18094), .dinb(n18091), .dout(n18095));
  jand g17842(.dina(n18095), .dinb(n18090), .dout(n18096));
  jor  g17843(.dina(n18096), .dinb(n884), .dout(n18097));
  jand g17844(.dina(n18096), .dinb(n884), .dout(n18098));
  jxor g17845(.dina(n17437), .dinb(n1008), .dout(n18099));
  jor  g17846(.dina(n18099), .dinb(n17769), .dout(n18100));
  jxor g17847(.dina(n18100), .dinb(n17719), .dout(n18101));
  jnot g17848(.din(n18101), .dout(n18102));
  jor  g17849(.dina(n18102), .dinb(n18098), .dout(n18103));
  jand g17850(.dina(n18103), .dinb(n18097), .dout(n18104));
  jor  g17851(.dina(n18104), .dinb(n743), .dout(n18105));
  jand g17852(.dina(n18104), .dinb(n743), .dout(n18106));
  jxor g17853(.dina(n17444), .dinb(n884), .dout(n18107));
  jor  g17854(.dina(n18107), .dinb(n17769), .dout(n18108));
  jxor g17855(.dina(n18108), .dinb(n17450), .dout(n18109));
  jor  g17856(.dina(n18109), .dinb(n18106), .dout(n18110));
  jand g17857(.dina(n18110), .dinb(n18105), .dout(n18111));
  jor  g17858(.dina(n18111), .dinb(n635), .dout(n18112));
  jand g17859(.dina(n18111), .dinb(n635), .dout(n18113));
  jxor g17860(.dina(n17452), .dinb(n743), .dout(n18114));
  jor  g17861(.dina(n18114), .dinb(n17769), .dout(n18115));
  jxor g17862(.dina(n18115), .dinb(n17726), .dout(n18116));
  jnot g17863(.din(n18116), .dout(n18117));
  jor  g17864(.dina(n18117), .dinb(n18113), .dout(n18118));
  jand g17865(.dina(n18118), .dinb(n18112), .dout(n18119));
  jor  g17866(.dina(n18119), .dinb(n515), .dout(n18120));
  jand g17867(.dina(n18119), .dinb(n515), .dout(n18121));
  jxor g17868(.dina(n17459), .dinb(n635), .dout(n18122));
  jor  g17869(.dina(n18122), .dinb(n17769), .dout(n18123));
  jxor g17870(.dina(n18123), .dinb(n17465), .dout(n18124));
  jor  g17871(.dina(n18124), .dinb(n18121), .dout(n18125));
  jand g17872(.dina(n18125), .dinb(n18120), .dout(n18126));
  jor  g17873(.dina(n18126), .dinb(n443), .dout(n18127));
  jand g17874(.dina(n18126), .dinb(n443), .dout(n18128));
  jxor g17875(.dina(n17467), .dinb(n515), .dout(n18129));
  jor  g17876(.dina(n18129), .dinb(n17769), .dout(n18130));
  jxor g17877(.dina(n18130), .dinb(n17473), .dout(n18131));
  jor  g17878(.dina(n18131), .dinb(n18128), .dout(n18132));
  jand g17879(.dina(n18132), .dinb(n18127), .dout(n18133));
  jor  g17880(.dina(n18133), .dinb(n352), .dout(n18134));
  jand g17881(.dina(n18133), .dinb(n352), .dout(n18135));
  jxor g17882(.dina(n17475), .dinb(n443), .dout(n18136));
  jor  g17883(.dina(n18136), .dinb(n17769), .dout(n18137));
  jxor g17884(.dina(n18137), .dinb(n17481), .dout(n18138));
  jor  g17885(.dina(n18138), .dinb(n18135), .dout(n18139));
  jand g17886(.dina(n18139), .dinb(n18134), .dout(n18140));
  jor  g17887(.dina(n18140), .dinb(n294), .dout(n18141));
  jand g17888(.dina(n18140), .dinb(n294), .dout(n18142));
  jxor g17889(.dina(n17483), .dinb(n352), .dout(n18143));
  jor  g17890(.dina(n18143), .dinb(n17769), .dout(n18144));
  jxor g17891(.dina(n18144), .dinb(n17739), .dout(n18145));
  jnot g17892(.din(n18145), .dout(n18146));
  jor  g17893(.dina(n18146), .dinb(n18142), .dout(n18147));
  jand g17894(.dina(n18147), .dinb(n18141), .dout(n18148));
  jor  g17895(.dina(n18148), .dinb(n239), .dout(n18149));
  jand g17896(.dina(n18148), .dinb(n239), .dout(n18150));
  jxor g17897(.dina(n17490), .dinb(n294), .dout(n18151));
  jor  g17898(.dina(n18151), .dinb(n17769), .dout(n18152));
  jxor g17899(.dina(n18152), .dinb(n17496), .dout(n18153));
  jor  g17900(.dina(n18153), .dinb(n18150), .dout(n18154));
  jand g17901(.dina(n18154), .dinb(n18149), .dout(n18155));
  jor  g17902(.dina(n18155), .dinb(n221), .dout(n18156));
  jand g17903(.dina(n18155), .dinb(n221), .dout(n18157));
  jxor g17904(.dina(n17498), .dinb(n239), .dout(n18158));
  jor  g17905(.dina(n18158), .dinb(n17769), .dout(n18159));
  jxor g17906(.dina(n18159), .dinb(n17746), .dout(n18160));
  jnot g17907(.din(n18160), .dout(n18161));
  jor  g17908(.dina(n18161), .dinb(n18157), .dout(n18162));
  jand g17909(.dina(n18162), .dinb(n18156), .dout(n18163));
  jand g17910(.dina(n18163), .dinb(n17773), .dout(n18164));
  jand g17911(.dina(n17768), .dinb(n17751), .dout(n18165));
  jand g17912(.dina(n17752), .dinb(asqrt[63] ), .dout(n18166));
  jand g17913(.dina(n18166), .dinb(n17518), .dout(n18167));
  jnot g17914(.din(n18167), .dout(n18168));
  jor  g17915(.dina(n18168), .dinb(n18165), .dout(n18169));
  jnot g17916(.din(n18169), .dout(n18170));
  jand g17917(.dina(n17758), .dinb(n17762), .dout(n18171));
  jor  g17918(.dina(n18163), .dinb(n17773), .dout(n18172));
  jor  g17919(.dina(n18172), .dinb(n17519), .dout(n18173));
  jor  g17920(.dina(n18173), .dinb(n18171), .dout(n18174));
  jand g17921(.dina(n18174), .dinb(n218), .dout(n18175));
  jand g17922(.dina(n17769), .dinb(n17516), .dout(n18176));
  jor  g17923(.dina(n18176), .dinb(n18175), .dout(n18177));
  jor  g17924(.dina(n18177), .dinb(n18170), .dout(n18178));
  jor  g17925(.dina(n18178), .dinb(n18164), .dout(asqrt[10] ));
  jxor g17926(.dina(n18155), .dinb(n221), .dout(n18180));
  jand g17927(.dina(n18180), .dinb(asqrt[10] ), .dout(n18181));
  jxor g17928(.dina(n18181), .dinb(n18160), .dout(n18182));
  jnot g17929(.din(n18182), .dout(n18183));
  jand g17930(.dina(asqrt[10] ), .dinb(a[20] ), .dout(n18184));
  jnot g17931(.din(a[18] ), .dout(n18185));
  jnot g17932(.din(a[19] ), .dout(n18186));
  jand g17933(.dina(n18186), .dinb(n18185), .dout(n18187));
  jand g17934(.dina(n18187), .dinb(n17774), .dout(n18188));
  jor  g17935(.dina(n18188), .dinb(n18184), .dout(n18189));
  jand g17936(.dina(n18189), .dinb(asqrt[11] ), .dout(n18190));
  jor  g17937(.dina(n18189), .dinb(asqrt[11] ), .dout(n18191));
  jand g17938(.dina(asqrt[10] ), .dinb(n17774), .dout(n18192));
  jor  g17939(.dina(n18192), .dinb(n17775), .dout(n18193));
  jnot g17940(.din(n17776), .dout(n18194));
  jnot g17941(.din(n18164), .dout(n18195));
  jnot g17942(.din(n18171), .dout(n18196));
  jnot g17943(.din(n18156), .dout(n18197));
  jnot g17944(.din(n18149), .dout(n18198));
  jnot g17945(.din(n18141), .dout(n18199));
  jnot g17946(.din(n18134), .dout(n18200));
  jnot g17947(.din(n18127), .dout(n18201));
  jnot g17948(.din(n18120), .dout(n18202));
  jnot g17949(.din(n18112), .dout(n18203));
  jnot g17950(.din(n18105), .dout(n18204));
  jnot g17951(.din(n18097), .dout(n18205));
  jnot g17952(.din(n18090), .dout(n18206));
  jnot g17953(.din(n18082), .dout(n18207));
  jnot g17954(.din(n18074), .dout(n18208));
  jnot g17955(.din(n18067), .dout(n18209));
  jnot g17956(.din(n18060), .dout(n18210));
  jnot g17957(.din(n18052), .dout(n18211));
  jnot g17958(.din(n18045), .dout(n18212));
  jnot g17959(.din(n18037), .dout(n18213));
  jnot g17960(.din(n18030), .dout(n18214));
  jnot g17961(.din(n18023), .dout(n18215));
  jnot g17962(.din(n18016), .dout(n18216));
  jnot g17963(.din(n18008), .dout(n18217));
  jnot g17964(.din(n18001), .dout(n18218));
  jnot g17965(.din(n17993), .dout(n18219));
  jnot g17966(.din(n17986), .dout(n18220));
  jnot g17967(.din(n17979), .dout(n18221));
  jnot g17968(.din(n17972), .dout(n18222));
  jnot g17969(.din(n17964), .dout(n18223));
  jnot g17970(.din(n17957), .dout(n18224));
  jnot g17971(.din(n17949), .dout(n18225));
  jnot g17972(.din(n17942), .dout(n18226));
  jnot g17973(.din(n17934), .dout(n18227));
  jnot g17974(.din(n17927), .dout(n18228));
  jnot g17975(.din(n17919), .dout(n18229));
  jnot g17976(.din(n17912), .dout(n18230));
  jnot g17977(.din(n17905), .dout(n18231));
  jnot g17978(.din(n17898), .dout(n18232));
  jnot g17979(.din(n17890), .dout(n18233));
  jnot g17980(.din(n17883), .dout(n18234));
  jnot g17981(.din(n17875), .dout(n18235));
  jnot g17982(.din(n17868), .dout(n18236));
  jnot g17983(.din(n17860), .dout(n18237));
  jnot g17984(.din(n17852), .dout(n18238));
  jnot g17985(.din(n17845), .dout(n18239));
  jnot g17986(.din(n17838), .dout(n18240));
  jnot g17987(.din(n17830), .dout(n18241));
  jnot g17988(.din(n17823), .dout(n18242));
  jnot g17989(.din(n17815), .dout(n18243));
  jnot g17990(.din(n17808), .dout(n18244));
  jnot g17991(.din(n17800), .dout(n18245));
  jnot g17992(.din(n17789), .dout(n18246));
  jnot g17993(.din(n17781), .dout(n18247));
  jand g17994(.dina(asqrt[11] ), .dinb(a[22] ), .dout(n18248));
  jor  g17995(.dina(n18248), .dinb(n17777), .dout(n18249));
  jor  g17996(.dina(n18249), .dinb(asqrt[12] ), .dout(n18250));
  jand g17997(.dina(asqrt[11] ), .dinb(n16885), .dout(n18251));
  jor  g17998(.dina(n18251), .dinb(n16886), .dout(n18252));
  jand g17999(.dina(n17792), .dinb(n18252), .dout(n18253));
  jand g18000(.dina(n18253), .dinb(n18250), .dout(n18254));
  jor  g18001(.dina(n18254), .dinb(n18247), .dout(n18255));
  jor  g18002(.dina(n18255), .dinb(asqrt[13] ), .dout(n18256));
  jnot g18003(.din(n17797), .dout(n18257));
  jand g18004(.dina(n18257), .dinb(n18256), .dout(n18258));
  jor  g18005(.dina(n18258), .dinb(n18246), .dout(n18259));
  jor  g18006(.dina(n18259), .dinb(asqrt[14] ), .dout(n18260));
  jand g18007(.dina(n17804), .dinb(n18260), .dout(n18261));
  jor  g18008(.dina(n18261), .dinb(n18245), .dout(n18262));
  jor  g18009(.dina(n18262), .dinb(asqrt[15] ), .dout(n18263));
  jnot g18010(.din(n17812), .dout(n18264));
  jand g18011(.dina(n18264), .dinb(n18263), .dout(n18265));
  jor  g18012(.dina(n18265), .dinb(n18244), .dout(n18266));
  jor  g18013(.dina(n18266), .dinb(asqrt[16] ), .dout(n18267));
  jand g18014(.dina(n17819), .dinb(n18267), .dout(n18268));
  jor  g18015(.dina(n18268), .dinb(n18243), .dout(n18269));
  jor  g18016(.dina(n18269), .dinb(asqrt[17] ), .dout(n18270));
  jnot g18017(.din(n17827), .dout(n18271));
  jand g18018(.dina(n18271), .dinb(n18270), .dout(n18272));
  jor  g18019(.dina(n18272), .dinb(n18242), .dout(n18273));
  jor  g18020(.dina(n18273), .dinb(asqrt[18] ), .dout(n18274));
  jand g18021(.dina(n17834), .dinb(n18274), .dout(n18275));
  jor  g18022(.dina(n18275), .dinb(n18241), .dout(n18276));
  jor  g18023(.dina(n18276), .dinb(asqrt[19] ), .dout(n18277));
  jnot g18024(.din(n17842), .dout(n18278));
  jand g18025(.dina(n18278), .dinb(n18277), .dout(n18279));
  jor  g18026(.dina(n18279), .dinb(n18240), .dout(n18280));
  jor  g18027(.dina(n18280), .dinb(asqrt[20] ), .dout(n18281));
  jnot g18028(.din(n17849), .dout(n18282));
  jand g18029(.dina(n18282), .dinb(n18281), .dout(n18283));
  jor  g18030(.dina(n18283), .dinb(n18239), .dout(n18284));
  jor  g18031(.dina(n18284), .dinb(asqrt[21] ), .dout(n18285));
  jand g18032(.dina(n17856), .dinb(n18285), .dout(n18286));
  jor  g18033(.dina(n18286), .dinb(n18238), .dout(n18287));
  jor  g18034(.dina(n18287), .dinb(asqrt[22] ), .dout(n18288));
  jand g18035(.dina(n17864), .dinb(n18288), .dout(n18289));
  jor  g18036(.dina(n18289), .dinb(n18237), .dout(n18290));
  jor  g18037(.dina(n18290), .dinb(asqrt[23] ), .dout(n18291));
  jnot g18038(.din(n17872), .dout(n18292));
  jand g18039(.dina(n18292), .dinb(n18291), .dout(n18293));
  jor  g18040(.dina(n18293), .dinb(n18236), .dout(n18294));
  jor  g18041(.dina(n18294), .dinb(asqrt[24] ), .dout(n18295));
  jand g18042(.dina(n17879), .dinb(n18295), .dout(n18296));
  jor  g18043(.dina(n18296), .dinb(n18235), .dout(n18297));
  jor  g18044(.dina(n18297), .dinb(asqrt[25] ), .dout(n18298));
  jnot g18045(.din(n17887), .dout(n18299));
  jand g18046(.dina(n18299), .dinb(n18298), .dout(n18300));
  jor  g18047(.dina(n18300), .dinb(n18234), .dout(n18301));
  jor  g18048(.dina(n18301), .dinb(asqrt[26] ), .dout(n18302));
  jand g18049(.dina(n17894), .dinb(n18302), .dout(n18303));
  jor  g18050(.dina(n18303), .dinb(n18233), .dout(n18304));
  jor  g18051(.dina(n18304), .dinb(asqrt[27] ), .dout(n18305));
  jnot g18052(.din(n17902), .dout(n18306));
  jand g18053(.dina(n18306), .dinb(n18305), .dout(n18307));
  jor  g18054(.dina(n18307), .dinb(n18232), .dout(n18308));
  jor  g18055(.dina(n18308), .dinb(asqrt[28] ), .dout(n18309));
  jnot g18056(.din(n17909), .dout(n18310));
  jand g18057(.dina(n18310), .dinb(n18309), .dout(n18311));
  jor  g18058(.dina(n18311), .dinb(n18231), .dout(n18312));
  jor  g18059(.dina(n18312), .dinb(asqrt[29] ), .dout(n18313));
  jnot g18060(.din(n17916), .dout(n18314));
  jand g18061(.dina(n18314), .dinb(n18313), .dout(n18315));
  jor  g18062(.dina(n18315), .dinb(n18230), .dout(n18316));
  jor  g18063(.dina(n18316), .dinb(asqrt[30] ), .dout(n18317));
  jand g18064(.dina(n17923), .dinb(n18317), .dout(n18318));
  jor  g18065(.dina(n18318), .dinb(n18229), .dout(n18319));
  jor  g18066(.dina(n18319), .dinb(asqrt[31] ), .dout(n18320));
  jnot g18067(.din(n17931), .dout(n18321));
  jand g18068(.dina(n18321), .dinb(n18320), .dout(n18322));
  jor  g18069(.dina(n18322), .dinb(n18228), .dout(n18323));
  jor  g18070(.dina(n18323), .dinb(asqrt[32] ), .dout(n18324));
  jand g18071(.dina(n17938), .dinb(n18324), .dout(n18325));
  jor  g18072(.dina(n18325), .dinb(n18227), .dout(n18326));
  jor  g18073(.dina(n18326), .dinb(asqrt[33] ), .dout(n18327));
  jnot g18074(.din(n17946), .dout(n18328));
  jand g18075(.dina(n18328), .dinb(n18327), .dout(n18329));
  jor  g18076(.dina(n18329), .dinb(n18226), .dout(n18330));
  jor  g18077(.dina(n18330), .dinb(asqrt[34] ), .dout(n18331));
  jand g18078(.dina(n17953), .dinb(n18331), .dout(n18332));
  jor  g18079(.dina(n18332), .dinb(n18225), .dout(n18333));
  jor  g18080(.dina(n18333), .dinb(asqrt[35] ), .dout(n18334));
  jnot g18081(.din(n17961), .dout(n18335));
  jand g18082(.dina(n18335), .dinb(n18334), .dout(n18336));
  jor  g18083(.dina(n18336), .dinb(n18224), .dout(n18337));
  jor  g18084(.dina(n18337), .dinb(asqrt[36] ), .dout(n18338));
  jand g18085(.dina(n17968), .dinb(n18338), .dout(n18339));
  jor  g18086(.dina(n18339), .dinb(n18223), .dout(n18340));
  jor  g18087(.dina(n18340), .dinb(asqrt[37] ), .dout(n18341));
  jnot g18088(.din(n17976), .dout(n18342));
  jand g18089(.dina(n18342), .dinb(n18341), .dout(n18343));
  jor  g18090(.dina(n18343), .dinb(n18222), .dout(n18344));
  jor  g18091(.dina(n18344), .dinb(asqrt[38] ), .dout(n18345));
  jnot g18092(.din(n17983), .dout(n18346));
  jand g18093(.dina(n18346), .dinb(n18345), .dout(n18347));
  jor  g18094(.dina(n18347), .dinb(n18221), .dout(n18348));
  jor  g18095(.dina(n18348), .dinb(asqrt[39] ), .dout(n18349));
  jnot g18096(.din(n17990), .dout(n18350));
  jand g18097(.dina(n18350), .dinb(n18349), .dout(n18351));
  jor  g18098(.dina(n18351), .dinb(n18220), .dout(n18352));
  jor  g18099(.dina(n18352), .dinb(asqrt[40] ), .dout(n18353));
  jand g18100(.dina(n17997), .dinb(n18353), .dout(n18354));
  jor  g18101(.dina(n18354), .dinb(n18219), .dout(n18355));
  jor  g18102(.dina(n18355), .dinb(asqrt[41] ), .dout(n18356));
  jnot g18103(.din(n18005), .dout(n18357));
  jand g18104(.dina(n18357), .dinb(n18356), .dout(n18358));
  jor  g18105(.dina(n18358), .dinb(n18218), .dout(n18359));
  jor  g18106(.dina(n18359), .dinb(asqrt[42] ), .dout(n18360));
  jand g18107(.dina(n18012), .dinb(n18360), .dout(n18361));
  jor  g18108(.dina(n18361), .dinb(n18217), .dout(n18362));
  jor  g18109(.dina(n18362), .dinb(asqrt[43] ), .dout(n18363));
  jnot g18110(.din(n18020), .dout(n18364));
  jand g18111(.dina(n18364), .dinb(n18363), .dout(n18365));
  jor  g18112(.dina(n18365), .dinb(n18216), .dout(n18366));
  jor  g18113(.dina(n18366), .dinb(asqrt[44] ), .dout(n18367));
  jnot g18114(.din(n18027), .dout(n18368));
  jand g18115(.dina(n18368), .dinb(n18367), .dout(n18369));
  jor  g18116(.dina(n18369), .dinb(n18215), .dout(n18370));
  jor  g18117(.dina(n18370), .dinb(asqrt[45] ), .dout(n18371));
  jnot g18118(.din(n18034), .dout(n18372));
  jand g18119(.dina(n18372), .dinb(n18371), .dout(n18373));
  jor  g18120(.dina(n18373), .dinb(n18214), .dout(n18374));
  jor  g18121(.dina(n18374), .dinb(asqrt[46] ), .dout(n18375));
  jand g18122(.dina(n18041), .dinb(n18375), .dout(n18376));
  jor  g18123(.dina(n18376), .dinb(n18213), .dout(n18377));
  jor  g18124(.dina(n18377), .dinb(asqrt[47] ), .dout(n18378));
  jnot g18125(.din(n18049), .dout(n18379));
  jand g18126(.dina(n18379), .dinb(n18378), .dout(n18380));
  jor  g18127(.dina(n18380), .dinb(n18212), .dout(n18381));
  jor  g18128(.dina(n18381), .dinb(asqrt[48] ), .dout(n18382));
  jand g18129(.dina(n18056), .dinb(n18382), .dout(n18383));
  jor  g18130(.dina(n18383), .dinb(n18211), .dout(n18384));
  jor  g18131(.dina(n18384), .dinb(asqrt[49] ), .dout(n18385));
  jnot g18132(.din(n18064), .dout(n18386));
  jand g18133(.dina(n18386), .dinb(n18385), .dout(n18387));
  jor  g18134(.dina(n18387), .dinb(n18210), .dout(n18388));
  jor  g18135(.dina(n18388), .dinb(asqrt[50] ), .dout(n18389));
  jnot g18136(.din(n18071), .dout(n18390));
  jand g18137(.dina(n18390), .dinb(n18389), .dout(n18391));
  jor  g18138(.dina(n18391), .dinb(n18209), .dout(n18392));
  jor  g18139(.dina(n18392), .dinb(asqrt[51] ), .dout(n18393));
  jand g18140(.dina(n18078), .dinb(n18393), .dout(n18394));
  jor  g18141(.dina(n18394), .dinb(n18208), .dout(n18395));
  jor  g18142(.dina(n18395), .dinb(asqrt[52] ), .dout(n18396));
  jand g18143(.dina(n18396), .dinb(n18085), .dout(n18397));
  jor  g18144(.dina(n18397), .dinb(n18207), .dout(n18398));
  jor  g18145(.dina(n18398), .dinb(asqrt[53] ), .dout(n18399));
  jnot g18146(.din(n18094), .dout(n18400));
  jand g18147(.dina(n18400), .dinb(n18399), .dout(n18401));
  jor  g18148(.dina(n18401), .dinb(n18206), .dout(n18402));
  jor  g18149(.dina(n18402), .dinb(asqrt[54] ), .dout(n18403));
  jand g18150(.dina(n18101), .dinb(n18403), .dout(n18404));
  jor  g18151(.dina(n18404), .dinb(n18205), .dout(n18405));
  jor  g18152(.dina(n18405), .dinb(asqrt[55] ), .dout(n18406));
  jnot g18153(.din(n18109), .dout(n18407));
  jand g18154(.dina(n18407), .dinb(n18406), .dout(n18408));
  jor  g18155(.dina(n18408), .dinb(n18204), .dout(n18409));
  jor  g18156(.dina(n18409), .dinb(asqrt[56] ), .dout(n18410));
  jand g18157(.dina(n18116), .dinb(n18410), .dout(n18411));
  jor  g18158(.dina(n18411), .dinb(n18203), .dout(n18412));
  jor  g18159(.dina(n18412), .dinb(asqrt[57] ), .dout(n18413));
  jnot g18160(.din(n18124), .dout(n18414));
  jand g18161(.dina(n18414), .dinb(n18413), .dout(n18415));
  jor  g18162(.dina(n18415), .dinb(n18202), .dout(n18416));
  jor  g18163(.dina(n18416), .dinb(asqrt[58] ), .dout(n18417));
  jnot g18164(.din(n18131), .dout(n18418));
  jand g18165(.dina(n18418), .dinb(n18417), .dout(n18419));
  jor  g18166(.dina(n18419), .dinb(n18201), .dout(n18420));
  jor  g18167(.dina(n18420), .dinb(asqrt[59] ), .dout(n18421));
  jnot g18168(.din(n18138), .dout(n18422));
  jand g18169(.dina(n18422), .dinb(n18421), .dout(n18423));
  jor  g18170(.dina(n18423), .dinb(n18200), .dout(n18424));
  jor  g18171(.dina(n18424), .dinb(asqrt[60] ), .dout(n18425));
  jand g18172(.dina(n18145), .dinb(n18425), .dout(n18426));
  jor  g18173(.dina(n18426), .dinb(n18199), .dout(n18427));
  jor  g18174(.dina(n18427), .dinb(asqrt[61] ), .dout(n18428));
  jnot g18175(.din(n18153), .dout(n18429));
  jand g18176(.dina(n18429), .dinb(n18428), .dout(n18430));
  jor  g18177(.dina(n18430), .dinb(n18198), .dout(n18431));
  jor  g18178(.dina(n18431), .dinb(asqrt[62] ), .dout(n18432));
  jand g18179(.dina(n18160), .dinb(n18432), .dout(n18433));
  jor  g18180(.dina(n18433), .dinb(n18197), .dout(n18434));
  jand g18181(.dina(n18434), .dinb(n17772), .dout(n18435));
  jand g18182(.dina(n18435), .dinb(n17518), .dout(n18436));
  jand g18183(.dina(n18436), .dinb(n18196), .dout(n18437));
  jor  g18184(.dina(n18437), .dinb(asqrt[63] ), .dout(n18438));
  jnot g18185(.din(n18176), .dout(n18439));
  jand g18186(.dina(n18439), .dinb(n18438), .dout(n18440));
  jand g18187(.dina(n18440), .dinb(n18169), .dout(n18441));
  jand g18188(.dina(n18441), .dinb(n18195), .dout(n18442));
  jor  g18189(.dina(n18442), .dinb(n18194), .dout(n18443));
  jand g18190(.dina(n18443), .dinb(n18193), .dout(n18444));
  jand g18191(.dina(n18444), .dinb(n18191), .dout(n18445));
  jor  g18192(.dina(n18445), .dinb(n18190), .dout(n18446));
  jand g18193(.dina(n18446), .dinb(asqrt[12] ), .dout(n18447));
  jor  g18194(.dina(n18446), .dinb(asqrt[12] ), .dout(n18448));
  jand g18195(.dina(asqrt[10] ), .dinb(n17776), .dout(n18449));
  jand g18196(.dina(n18195), .dinb(asqrt[11] ), .dout(n18450));
  jand g18197(.dina(n18450), .dinb(n18438), .dout(n18451));
  jand g18198(.dina(n18451), .dinb(n18168), .dout(n18452));
  jor  g18199(.dina(n18452), .dinb(n18449), .dout(n18453));
  jxor g18200(.dina(n18453), .dinb(a[22] ), .dout(n18454));
  jnot g18201(.din(n18454), .dout(n18455));
  jand g18202(.dina(n18455), .dinb(n18448), .dout(n18456));
  jor  g18203(.dina(n18456), .dinb(n18447), .dout(n18457));
  jand g18204(.dina(n18457), .dinb(asqrt[13] ), .dout(n18458));
  jor  g18205(.dina(n18457), .dinb(asqrt[13] ), .dout(n18459));
  jxor g18206(.dina(n17780), .dinb(n17134), .dout(n18460));
  jand g18207(.dina(n18460), .dinb(asqrt[10] ), .dout(n18461));
  jxor g18208(.dina(n18461), .dinb(n18253), .dout(n18462));
  jand g18209(.dina(n18462), .dinb(n18459), .dout(n18463));
  jor  g18210(.dina(n18463), .dinb(n18458), .dout(n18464));
  jand g18211(.dina(n18464), .dinb(asqrt[14] ), .dout(n18465));
  jor  g18212(.dina(n18464), .dinb(asqrt[14] ), .dout(n18466));
  jxor g18213(.dina(n17788), .dinb(n16489), .dout(n18467));
  jand g18214(.dina(n18467), .dinb(asqrt[10] ), .dout(n18468));
  jxor g18215(.dina(n18468), .dinb(n17797), .dout(n18469));
  jnot g18216(.din(n18469), .dout(n18470));
  jand g18217(.dina(n18470), .dinb(n18466), .dout(n18471));
  jor  g18218(.dina(n18471), .dinb(n18465), .dout(n18472));
  jand g18219(.dina(n18472), .dinb(asqrt[15] ), .dout(n18473));
  jor  g18220(.dina(n18472), .dinb(asqrt[15] ), .dout(n18474));
  jxor g18221(.dina(n17799), .dinb(n15878), .dout(n18475));
  jand g18222(.dina(n18475), .dinb(asqrt[10] ), .dout(n18476));
  jxor g18223(.dina(n18476), .dinb(n17804), .dout(n18477));
  jand g18224(.dina(n18477), .dinb(n18474), .dout(n18478));
  jor  g18225(.dina(n18478), .dinb(n18473), .dout(n18479));
  jand g18226(.dina(n18479), .dinb(asqrt[16] ), .dout(n18480));
  jor  g18227(.dina(n18479), .dinb(asqrt[16] ), .dout(n18481));
  jxor g18228(.dina(n17807), .dinb(n15260), .dout(n18482));
  jand g18229(.dina(n18482), .dinb(asqrt[10] ), .dout(n18483));
  jxor g18230(.dina(n18483), .dinb(n17812), .dout(n18484));
  jnot g18231(.din(n18484), .dout(n18485));
  jand g18232(.dina(n18485), .dinb(n18481), .dout(n18486));
  jor  g18233(.dina(n18486), .dinb(n18480), .dout(n18487));
  jand g18234(.dina(n18487), .dinb(asqrt[17] ), .dout(n18488));
  jor  g18235(.dina(n18487), .dinb(asqrt[17] ), .dout(n18489));
  jxor g18236(.dina(n17814), .dinb(n14674), .dout(n18490));
  jand g18237(.dina(n18490), .dinb(asqrt[10] ), .dout(n18491));
  jxor g18238(.dina(n18491), .dinb(n17819), .dout(n18492));
  jand g18239(.dina(n18492), .dinb(n18489), .dout(n18493));
  jor  g18240(.dina(n18493), .dinb(n18488), .dout(n18494));
  jand g18241(.dina(n18494), .dinb(asqrt[18] ), .dout(n18495));
  jor  g18242(.dina(n18494), .dinb(asqrt[18] ), .dout(n18496));
  jxor g18243(.dina(n17822), .dinb(n14078), .dout(n18497));
  jand g18244(.dina(n18497), .dinb(asqrt[10] ), .dout(n18498));
  jxor g18245(.dina(n18498), .dinb(n17827), .dout(n18499));
  jnot g18246(.din(n18499), .dout(n18500));
  jand g18247(.dina(n18500), .dinb(n18496), .dout(n18501));
  jor  g18248(.dina(n18501), .dinb(n18495), .dout(n18502));
  jand g18249(.dina(n18502), .dinb(asqrt[19] ), .dout(n18503));
  jor  g18250(.dina(n18502), .dinb(asqrt[19] ), .dout(n18504));
  jxor g18251(.dina(n17829), .dinb(n13515), .dout(n18505));
  jand g18252(.dina(n18505), .dinb(asqrt[10] ), .dout(n18506));
  jxor g18253(.dina(n18506), .dinb(n17834), .dout(n18507));
  jand g18254(.dina(n18507), .dinb(n18504), .dout(n18508));
  jor  g18255(.dina(n18508), .dinb(n18503), .dout(n18509));
  jand g18256(.dina(n18509), .dinb(asqrt[20] ), .dout(n18510));
  jor  g18257(.dina(n18509), .dinb(asqrt[20] ), .dout(n18511));
  jxor g18258(.dina(n17837), .dinb(n12947), .dout(n18512));
  jand g18259(.dina(n18512), .dinb(asqrt[10] ), .dout(n18513));
  jxor g18260(.dina(n18513), .dinb(n17842), .dout(n18514));
  jnot g18261(.din(n18514), .dout(n18515));
  jand g18262(.dina(n18515), .dinb(n18511), .dout(n18516));
  jor  g18263(.dina(n18516), .dinb(n18510), .dout(n18517));
  jand g18264(.dina(n18517), .dinb(asqrt[21] ), .dout(n18518));
  jor  g18265(.dina(n18517), .dinb(asqrt[21] ), .dout(n18519));
  jxor g18266(.dina(n17844), .dinb(n12410), .dout(n18520));
  jand g18267(.dina(n18520), .dinb(asqrt[10] ), .dout(n18521));
  jxor g18268(.dina(n18521), .dinb(n17849), .dout(n18522));
  jnot g18269(.din(n18522), .dout(n18523));
  jand g18270(.dina(n18523), .dinb(n18519), .dout(n18524));
  jor  g18271(.dina(n18524), .dinb(n18518), .dout(n18525));
  jand g18272(.dina(n18525), .dinb(asqrt[22] ), .dout(n18526));
  jor  g18273(.dina(n18525), .dinb(asqrt[22] ), .dout(n18527));
  jxor g18274(.dina(n17851), .dinb(n11858), .dout(n18528));
  jand g18275(.dina(n18528), .dinb(asqrt[10] ), .dout(n18529));
  jxor g18276(.dina(n18529), .dinb(n17856), .dout(n18530));
  jand g18277(.dina(n18530), .dinb(n18527), .dout(n18531));
  jor  g18278(.dina(n18531), .dinb(n18526), .dout(n18532));
  jand g18279(.dina(n18532), .dinb(asqrt[23] ), .dout(n18533));
  jor  g18280(.dina(n18532), .dinb(asqrt[23] ), .dout(n18534));
  jxor g18281(.dina(n17859), .dinb(n11347), .dout(n18535));
  jand g18282(.dina(n18535), .dinb(asqrt[10] ), .dout(n18536));
  jxor g18283(.dina(n18536), .dinb(n17864), .dout(n18537));
  jand g18284(.dina(n18537), .dinb(n18534), .dout(n18538));
  jor  g18285(.dina(n18538), .dinb(n18533), .dout(n18539));
  jand g18286(.dina(n18539), .dinb(asqrt[24] ), .dout(n18540));
  jor  g18287(.dina(n18539), .dinb(asqrt[24] ), .dout(n18541));
  jxor g18288(.dina(n17867), .dinb(n10824), .dout(n18542));
  jand g18289(.dina(n18542), .dinb(asqrt[10] ), .dout(n18543));
  jxor g18290(.dina(n18543), .dinb(n17872), .dout(n18544));
  jnot g18291(.din(n18544), .dout(n18545));
  jand g18292(.dina(n18545), .dinb(n18541), .dout(n18546));
  jor  g18293(.dina(n18546), .dinb(n18540), .dout(n18547));
  jand g18294(.dina(n18547), .dinb(asqrt[25] ), .dout(n18548));
  jor  g18295(.dina(n18547), .dinb(asqrt[25] ), .dout(n18549));
  jxor g18296(.dina(n17874), .dinb(n10328), .dout(n18550));
  jand g18297(.dina(n18550), .dinb(asqrt[10] ), .dout(n18551));
  jxor g18298(.dina(n18551), .dinb(n17879), .dout(n18552));
  jand g18299(.dina(n18552), .dinb(n18549), .dout(n18553));
  jor  g18300(.dina(n18553), .dinb(n18548), .dout(n18554));
  jand g18301(.dina(n18554), .dinb(asqrt[26] ), .dout(n18555));
  jor  g18302(.dina(n18554), .dinb(asqrt[26] ), .dout(n18556));
  jxor g18303(.dina(n17882), .dinb(n9832), .dout(n18557));
  jand g18304(.dina(n18557), .dinb(asqrt[10] ), .dout(n18558));
  jxor g18305(.dina(n18558), .dinb(n17887), .dout(n18559));
  jnot g18306(.din(n18559), .dout(n18560));
  jand g18307(.dina(n18560), .dinb(n18556), .dout(n18561));
  jor  g18308(.dina(n18561), .dinb(n18555), .dout(n18562));
  jand g18309(.dina(n18562), .dinb(asqrt[27] ), .dout(n18563));
  jor  g18310(.dina(n18562), .dinb(asqrt[27] ), .dout(n18564));
  jxor g18311(.dina(n17889), .dinb(n9369), .dout(n18565));
  jand g18312(.dina(n18565), .dinb(asqrt[10] ), .dout(n18566));
  jxor g18313(.dina(n18566), .dinb(n17894), .dout(n18567));
  jand g18314(.dina(n18567), .dinb(n18564), .dout(n18568));
  jor  g18315(.dina(n18568), .dinb(n18563), .dout(n18569));
  jand g18316(.dina(n18569), .dinb(asqrt[28] ), .dout(n18570));
  jor  g18317(.dina(n18569), .dinb(asqrt[28] ), .dout(n18571));
  jxor g18318(.dina(n17897), .dinb(n8890), .dout(n18572));
  jand g18319(.dina(n18572), .dinb(asqrt[10] ), .dout(n18573));
  jxor g18320(.dina(n18573), .dinb(n17902), .dout(n18574));
  jnot g18321(.din(n18574), .dout(n18575));
  jand g18322(.dina(n18575), .dinb(n18571), .dout(n18576));
  jor  g18323(.dina(n18576), .dinb(n18570), .dout(n18577));
  jand g18324(.dina(n18577), .dinb(asqrt[29] ), .dout(n18578));
  jor  g18325(.dina(n18577), .dinb(asqrt[29] ), .dout(n18579));
  jxor g18326(.dina(n17904), .dinb(n8449), .dout(n18580));
  jand g18327(.dina(n18580), .dinb(asqrt[10] ), .dout(n18581));
  jxor g18328(.dina(n18581), .dinb(n17909), .dout(n18582));
  jnot g18329(.din(n18582), .dout(n18583));
  jand g18330(.dina(n18583), .dinb(n18579), .dout(n18584));
  jor  g18331(.dina(n18584), .dinb(n18578), .dout(n18585));
  jand g18332(.dina(n18585), .dinb(asqrt[30] ), .dout(n18586));
  jor  g18333(.dina(n18585), .dinb(asqrt[30] ), .dout(n18587));
  jxor g18334(.dina(n17911), .dinb(n8003), .dout(n18588));
  jand g18335(.dina(n18588), .dinb(asqrt[10] ), .dout(n18589));
  jxor g18336(.dina(n18589), .dinb(n17916), .dout(n18590));
  jnot g18337(.din(n18590), .dout(n18591));
  jand g18338(.dina(n18591), .dinb(n18587), .dout(n18592));
  jor  g18339(.dina(n18592), .dinb(n18586), .dout(n18593));
  jand g18340(.dina(n18593), .dinb(asqrt[31] ), .dout(n18594));
  jor  g18341(.dina(n18593), .dinb(asqrt[31] ), .dout(n18595));
  jxor g18342(.dina(n17918), .dinb(n7581), .dout(n18596));
  jand g18343(.dina(n18596), .dinb(asqrt[10] ), .dout(n18597));
  jxor g18344(.dina(n18597), .dinb(n17923), .dout(n18598));
  jand g18345(.dina(n18598), .dinb(n18595), .dout(n18599));
  jor  g18346(.dina(n18599), .dinb(n18594), .dout(n18600));
  jand g18347(.dina(n18600), .dinb(asqrt[32] ), .dout(n18601));
  jor  g18348(.dina(n18600), .dinb(asqrt[32] ), .dout(n18602));
  jxor g18349(.dina(n17926), .dinb(n7154), .dout(n18603));
  jand g18350(.dina(n18603), .dinb(asqrt[10] ), .dout(n18604));
  jxor g18351(.dina(n18604), .dinb(n17931), .dout(n18605));
  jnot g18352(.din(n18605), .dout(n18606));
  jand g18353(.dina(n18606), .dinb(n18602), .dout(n18607));
  jor  g18354(.dina(n18607), .dinb(n18601), .dout(n18608));
  jand g18355(.dina(n18608), .dinb(asqrt[33] ), .dout(n18609));
  jor  g18356(.dina(n18608), .dinb(asqrt[33] ), .dout(n18610));
  jxor g18357(.dina(n17933), .dinb(n6758), .dout(n18611));
  jand g18358(.dina(n18611), .dinb(asqrt[10] ), .dout(n18612));
  jxor g18359(.dina(n18612), .dinb(n17938), .dout(n18613));
  jand g18360(.dina(n18613), .dinb(n18610), .dout(n18614));
  jor  g18361(.dina(n18614), .dinb(n18609), .dout(n18615));
  jand g18362(.dina(n18615), .dinb(asqrt[34] ), .dout(n18616));
  jor  g18363(.dina(n18615), .dinb(asqrt[34] ), .dout(n18617));
  jxor g18364(.dina(n17941), .dinb(n6357), .dout(n18618));
  jand g18365(.dina(n18618), .dinb(asqrt[10] ), .dout(n18619));
  jxor g18366(.dina(n18619), .dinb(n17946), .dout(n18620));
  jnot g18367(.din(n18620), .dout(n18621));
  jand g18368(.dina(n18621), .dinb(n18617), .dout(n18622));
  jor  g18369(.dina(n18622), .dinb(n18616), .dout(n18623));
  jand g18370(.dina(n18623), .dinb(asqrt[35] ), .dout(n18624));
  jor  g18371(.dina(n18623), .dinb(asqrt[35] ), .dout(n18625));
  jxor g18372(.dina(n17948), .dinb(n5989), .dout(n18626));
  jand g18373(.dina(n18626), .dinb(asqrt[10] ), .dout(n18627));
  jxor g18374(.dina(n18627), .dinb(n17953), .dout(n18628));
  jand g18375(.dina(n18628), .dinb(n18625), .dout(n18629));
  jor  g18376(.dina(n18629), .dinb(n18624), .dout(n18630));
  jand g18377(.dina(n18630), .dinb(asqrt[36] ), .dout(n18631));
  jor  g18378(.dina(n18630), .dinb(asqrt[36] ), .dout(n18632));
  jxor g18379(.dina(n17956), .dinb(n5606), .dout(n18633));
  jand g18380(.dina(n18633), .dinb(asqrt[10] ), .dout(n18634));
  jxor g18381(.dina(n18634), .dinb(n17961), .dout(n18635));
  jnot g18382(.din(n18635), .dout(n18636));
  jand g18383(.dina(n18636), .dinb(n18632), .dout(n18637));
  jor  g18384(.dina(n18637), .dinb(n18631), .dout(n18638));
  jand g18385(.dina(n18638), .dinb(asqrt[37] ), .dout(n18639));
  jor  g18386(.dina(n18638), .dinb(asqrt[37] ), .dout(n18640));
  jxor g18387(.dina(n17963), .dinb(n5259), .dout(n18641));
  jand g18388(.dina(n18641), .dinb(asqrt[10] ), .dout(n18642));
  jxor g18389(.dina(n18642), .dinb(n17968), .dout(n18643));
  jand g18390(.dina(n18643), .dinb(n18640), .dout(n18644));
  jor  g18391(.dina(n18644), .dinb(n18639), .dout(n18645));
  jand g18392(.dina(n18645), .dinb(asqrt[38] ), .dout(n18646));
  jor  g18393(.dina(n18645), .dinb(asqrt[38] ), .dout(n18647));
  jxor g18394(.dina(n17971), .dinb(n4902), .dout(n18648));
  jand g18395(.dina(n18648), .dinb(asqrt[10] ), .dout(n18649));
  jxor g18396(.dina(n18649), .dinb(n17976), .dout(n18650));
  jnot g18397(.din(n18650), .dout(n18651));
  jand g18398(.dina(n18651), .dinb(n18647), .dout(n18652));
  jor  g18399(.dina(n18652), .dinb(n18646), .dout(n18653));
  jand g18400(.dina(n18653), .dinb(asqrt[39] ), .dout(n18654));
  jor  g18401(.dina(n18653), .dinb(asqrt[39] ), .dout(n18655));
  jxor g18402(.dina(n17978), .dinb(n4582), .dout(n18656));
  jand g18403(.dina(n18656), .dinb(asqrt[10] ), .dout(n18657));
  jxor g18404(.dina(n18657), .dinb(n17983), .dout(n18658));
  jnot g18405(.din(n18658), .dout(n18659));
  jand g18406(.dina(n18659), .dinb(n18655), .dout(n18660));
  jor  g18407(.dina(n18660), .dinb(n18654), .dout(n18661));
  jand g18408(.dina(n18661), .dinb(asqrt[40] ), .dout(n18662));
  jor  g18409(.dina(n18661), .dinb(asqrt[40] ), .dout(n18663));
  jxor g18410(.dina(n17985), .dinb(n4249), .dout(n18664));
  jand g18411(.dina(n18664), .dinb(asqrt[10] ), .dout(n18665));
  jxor g18412(.dina(n18665), .dinb(n17990), .dout(n18666));
  jnot g18413(.din(n18666), .dout(n18667));
  jand g18414(.dina(n18667), .dinb(n18663), .dout(n18668));
  jor  g18415(.dina(n18668), .dinb(n18662), .dout(n18669));
  jand g18416(.dina(n18669), .dinb(asqrt[41] ), .dout(n18670));
  jor  g18417(.dina(n18669), .dinb(asqrt[41] ), .dout(n18671));
  jxor g18418(.dina(n17992), .dinb(n3955), .dout(n18672));
  jand g18419(.dina(n18672), .dinb(asqrt[10] ), .dout(n18673));
  jxor g18420(.dina(n18673), .dinb(n17997), .dout(n18674));
  jand g18421(.dina(n18674), .dinb(n18671), .dout(n18675));
  jor  g18422(.dina(n18675), .dinb(n18670), .dout(n18676));
  jand g18423(.dina(n18676), .dinb(asqrt[42] ), .dout(n18677));
  jor  g18424(.dina(n18676), .dinb(asqrt[42] ), .dout(n18678));
  jxor g18425(.dina(n18000), .dinb(n3642), .dout(n18679));
  jand g18426(.dina(n18679), .dinb(asqrt[10] ), .dout(n18680));
  jxor g18427(.dina(n18680), .dinb(n18005), .dout(n18681));
  jnot g18428(.din(n18681), .dout(n18682));
  jand g18429(.dina(n18682), .dinb(n18678), .dout(n18683));
  jor  g18430(.dina(n18683), .dinb(n18677), .dout(n18684));
  jand g18431(.dina(n18684), .dinb(asqrt[43] ), .dout(n18685));
  jor  g18432(.dina(n18684), .dinb(asqrt[43] ), .dout(n18686));
  jxor g18433(.dina(n18007), .dinb(n3368), .dout(n18687));
  jand g18434(.dina(n18687), .dinb(asqrt[10] ), .dout(n18688));
  jxor g18435(.dina(n18688), .dinb(n18013), .dout(n18689));
  jnot g18436(.din(n18689), .dout(n18690));
  jand g18437(.dina(n18690), .dinb(n18686), .dout(n18691));
  jor  g18438(.dina(n18691), .dinb(n18685), .dout(n18692));
  jand g18439(.dina(n18692), .dinb(asqrt[44] ), .dout(n18693));
  jor  g18440(.dina(n18692), .dinb(asqrt[44] ), .dout(n18694));
  jxor g18441(.dina(n18015), .dinb(n3089), .dout(n18695));
  jand g18442(.dina(n18695), .dinb(asqrt[10] ), .dout(n18696));
  jxor g18443(.dina(n18696), .dinb(n18020), .dout(n18697));
  jnot g18444(.din(n18697), .dout(n18698));
  jand g18445(.dina(n18698), .dinb(n18694), .dout(n18699));
  jor  g18446(.dina(n18699), .dinb(n18693), .dout(n18700));
  jand g18447(.dina(n18700), .dinb(asqrt[45] ), .dout(n18701));
  jor  g18448(.dina(n18700), .dinb(asqrt[45] ), .dout(n18702));
  jxor g18449(.dina(n18022), .dinb(n2833), .dout(n18703));
  jand g18450(.dina(n18703), .dinb(asqrt[10] ), .dout(n18704));
  jxor g18451(.dina(n18704), .dinb(n18027), .dout(n18705));
  jnot g18452(.din(n18705), .dout(n18706));
  jand g18453(.dina(n18706), .dinb(n18702), .dout(n18707));
  jor  g18454(.dina(n18707), .dinb(n18701), .dout(n18708));
  jand g18455(.dina(n18708), .dinb(asqrt[46] ), .dout(n18709));
  jor  g18456(.dina(n18708), .dinb(asqrt[46] ), .dout(n18710));
  jxor g18457(.dina(n18029), .dinb(n2572), .dout(n18711));
  jand g18458(.dina(n18711), .dinb(asqrt[10] ), .dout(n18712));
  jxor g18459(.dina(n18712), .dinb(n18034), .dout(n18713));
  jnot g18460(.din(n18713), .dout(n18714));
  jand g18461(.dina(n18714), .dinb(n18710), .dout(n18715));
  jor  g18462(.dina(n18715), .dinb(n18709), .dout(n18716));
  jand g18463(.dina(n18716), .dinb(asqrt[47] ), .dout(n18717));
  jor  g18464(.dina(n18716), .dinb(asqrt[47] ), .dout(n18718));
  jxor g18465(.dina(n18036), .dinb(n2345), .dout(n18719));
  jand g18466(.dina(n18719), .dinb(asqrt[10] ), .dout(n18720));
  jxor g18467(.dina(n18720), .dinb(n18041), .dout(n18721));
  jand g18468(.dina(n18721), .dinb(n18718), .dout(n18722));
  jor  g18469(.dina(n18722), .dinb(n18717), .dout(n18723));
  jand g18470(.dina(n18723), .dinb(asqrt[48] ), .dout(n18724));
  jor  g18471(.dina(n18723), .dinb(asqrt[48] ), .dout(n18725));
  jxor g18472(.dina(n18044), .dinb(n2108), .dout(n18726));
  jand g18473(.dina(n18726), .dinb(asqrt[10] ), .dout(n18727));
  jxor g18474(.dina(n18727), .dinb(n18049), .dout(n18728));
  jnot g18475(.din(n18728), .dout(n18729));
  jand g18476(.dina(n18729), .dinb(n18725), .dout(n18730));
  jor  g18477(.dina(n18730), .dinb(n18724), .dout(n18731));
  jand g18478(.dina(n18731), .dinb(asqrt[49] ), .dout(n18732));
  jor  g18479(.dina(n18731), .dinb(asqrt[49] ), .dout(n18733));
  jxor g18480(.dina(n18051), .dinb(n1912), .dout(n18734));
  jand g18481(.dina(n18734), .dinb(asqrt[10] ), .dout(n18735));
  jxor g18482(.dina(n18735), .dinb(n18056), .dout(n18736));
  jand g18483(.dina(n18736), .dinb(n18733), .dout(n18737));
  jor  g18484(.dina(n18737), .dinb(n18732), .dout(n18738));
  jand g18485(.dina(n18738), .dinb(asqrt[50] ), .dout(n18739));
  jor  g18486(.dina(n18738), .dinb(asqrt[50] ), .dout(n18740));
  jxor g18487(.dina(n18059), .dinb(n1699), .dout(n18741));
  jand g18488(.dina(n18741), .dinb(asqrt[10] ), .dout(n18742));
  jxor g18489(.dina(n18742), .dinb(n18064), .dout(n18743));
  jnot g18490(.din(n18743), .dout(n18744));
  jand g18491(.dina(n18744), .dinb(n18740), .dout(n18745));
  jor  g18492(.dina(n18745), .dinb(n18739), .dout(n18746));
  jand g18493(.dina(n18746), .dinb(asqrt[51] ), .dout(n18747));
  jor  g18494(.dina(n18746), .dinb(asqrt[51] ), .dout(n18748));
  jxor g18495(.dina(n18066), .dinb(n1516), .dout(n18749));
  jand g18496(.dina(n18749), .dinb(asqrt[10] ), .dout(n18750));
  jxor g18497(.dina(n18750), .dinb(n18071), .dout(n18751));
  jnot g18498(.din(n18751), .dout(n18752));
  jand g18499(.dina(n18752), .dinb(n18748), .dout(n18753));
  jor  g18500(.dina(n18753), .dinb(n18747), .dout(n18754));
  jand g18501(.dina(n18754), .dinb(asqrt[52] ), .dout(n18755));
  jor  g18502(.dina(n18754), .dinb(asqrt[52] ), .dout(n18756));
  jxor g18503(.dina(n18073), .dinb(n1332), .dout(n18757));
  jand g18504(.dina(n18757), .dinb(asqrt[10] ), .dout(n18758));
  jxor g18505(.dina(n18758), .dinb(n18078), .dout(n18759));
  jand g18506(.dina(n18759), .dinb(n18756), .dout(n18760));
  jor  g18507(.dina(n18760), .dinb(n18755), .dout(n18761));
  jand g18508(.dina(n18761), .dinb(asqrt[53] ), .dout(n18762));
  jxor g18509(.dina(n18081), .dinb(n1173), .dout(n18763));
  jand g18510(.dina(n18763), .dinb(asqrt[10] ), .dout(n18764));
  jxor g18511(.dina(n18764), .dinb(n18085), .dout(n18765));
  jor  g18512(.dina(n18761), .dinb(asqrt[53] ), .dout(n18766));
  jand g18513(.dina(n18766), .dinb(n18765), .dout(n18767));
  jor  g18514(.dina(n18767), .dinb(n18762), .dout(n18768));
  jand g18515(.dina(n18768), .dinb(asqrt[54] ), .dout(n18769));
  jor  g18516(.dina(n18768), .dinb(asqrt[54] ), .dout(n18770));
  jxor g18517(.dina(n18089), .dinb(n1008), .dout(n18771));
  jand g18518(.dina(n18771), .dinb(asqrt[10] ), .dout(n18772));
  jxor g18519(.dina(n18772), .dinb(n18094), .dout(n18773));
  jnot g18520(.din(n18773), .dout(n18774));
  jand g18521(.dina(n18774), .dinb(n18770), .dout(n18775));
  jor  g18522(.dina(n18775), .dinb(n18769), .dout(n18776));
  jand g18523(.dina(n18776), .dinb(asqrt[55] ), .dout(n18777));
  jor  g18524(.dina(n18776), .dinb(asqrt[55] ), .dout(n18778));
  jxor g18525(.dina(n18096), .dinb(n884), .dout(n18779));
  jand g18526(.dina(n18779), .dinb(asqrt[10] ), .dout(n18780));
  jxor g18527(.dina(n18780), .dinb(n18101), .dout(n18781));
  jand g18528(.dina(n18781), .dinb(n18778), .dout(n18782));
  jor  g18529(.dina(n18782), .dinb(n18777), .dout(n18783));
  jand g18530(.dina(n18783), .dinb(asqrt[56] ), .dout(n18784));
  jor  g18531(.dina(n18783), .dinb(asqrt[56] ), .dout(n18785));
  jxor g18532(.dina(n18104), .dinb(n743), .dout(n18786));
  jand g18533(.dina(n18786), .dinb(asqrt[10] ), .dout(n18787));
  jxor g18534(.dina(n18787), .dinb(n18109), .dout(n18788));
  jnot g18535(.din(n18788), .dout(n18789));
  jand g18536(.dina(n18789), .dinb(n18785), .dout(n18790));
  jor  g18537(.dina(n18790), .dinb(n18784), .dout(n18791));
  jand g18538(.dina(n18791), .dinb(asqrt[57] ), .dout(n18792));
  jor  g18539(.dina(n18791), .dinb(asqrt[57] ), .dout(n18793));
  jxor g18540(.dina(n18111), .dinb(n635), .dout(n18794));
  jand g18541(.dina(n18794), .dinb(asqrt[10] ), .dout(n18795));
  jxor g18542(.dina(n18795), .dinb(n18116), .dout(n18796));
  jand g18543(.dina(n18796), .dinb(n18793), .dout(n18797));
  jor  g18544(.dina(n18797), .dinb(n18792), .dout(n18798));
  jand g18545(.dina(n18798), .dinb(asqrt[58] ), .dout(n18799));
  jor  g18546(.dina(n18798), .dinb(asqrt[58] ), .dout(n18800));
  jxor g18547(.dina(n18119), .dinb(n515), .dout(n18801));
  jand g18548(.dina(n18801), .dinb(asqrt[10] ), .dout(n18802));
  jxor g18549(.dina(n18802), .dinb(n18124), .dout(n18803));
  jnot g18550(.din(n18803), .dout(n18804));
  jand g18551(.dina(n18804), .dinb(n18800), .dout(n18805));
  jor  g18552(.dina(n18805), .dinb(n18799), .dout(n18806));
  jand g18553(.dina(n18806), .dinb(asqrt[59] ), .dout(n18807));
  jor  g18554(.dina(n18806), .dinb(asqrt[59] ), .dout(n18808));
  jxor g18555(.dina(n18126), .dinb(n443), .dout(n18809));
  jand g18556(.dina(n18809), .dinb(asqrt[10] ), .dout(n18810));
  jxor g18557(.dina(n18810), .dinb(n18131), .dout(n18811));
  jnot g18558(.din(n18811), .dout(n18812));
  jand g18559(.dina(n18812), .dinb(n18808), .dout(n18813));
  jor  g18560(.dina(n18813), .dinb(n18807), .dout(n18814));
  jand g18561(.dina(n18814), .dinb(asqrt[60] ), .dout(n18815));
  jor  g18562(.dina(n18814), .dinb(asqrt[60] ), .dout(n18816));
  jxor g18563(.dina(n18133), .dinb(n352), .dout(n18817));
  jand g18564(.dina(n18817), .dinb(asqrt[10] ), .dout(n18818));
  jxor g18565(.dina(n18818), .dinb(n18138), .dout(n18819));
  jnot g18566(.din(n18819), .dout(n18820));
  jand g18567(.dina(n18820), .dinb(n18816), .dout(n18821));
  jor  g18568(.dina(n18821), .dinb(n18815), .dout(n18822));
  jand g18569(.dina(n18822), .dinb(asqrt[61] ), .dout(n18823));
  jor  g18570(.dina(n18822), .dinb(asqrt[61] ), .dout(n18824));
  jxor g18571(.dina(n18140), .dinb(n294), .dout(n18825));
  jand g18572(.dina(n18825), .dinb(asqrt[10] ), .dout(n18826));
  jxor g18573(.dina(n18826), .dinb(n18145), .dout(n18827));
  jand g18574(.dina(n18827), .dinb(n18824), .dout(n18828));
  jor  g18575(.dina(n18828), .dinb(n18823), .dout(n18829));
  jand g18576(.dina(n18829), .dinb(asqrt[62] ), .dout(n18830));
  jnot g18577(.din(n18830), .dout(n18831));
  jnot g18578(.din(n18823), .dout(n18832));
  jnot g18579(.din(n18815), .dout(n18833));
  jnot g18580(.din(n18807), .dout(n18834));
  jnot g18581(.din(n18799), .dout(n18835));
  jnot g18582(.din(n18792), .dout(n18836));
  jnot g18583(.din(n18784), .dout(n18837));
  jnot g18584(.din(n18777), .dout(n18838));
  jnot g18585(.din(n18769), .dout(n18839));
  jnot g18586(.din(n18762), .dout(n18840));
  jnot g18587(.din(n18765), .dout(n18841));
  jnot g18588(.din(n18755), .dout(n18842));
  jnot g18589(.din(n18747), .dout(n18843));
  jnot g18590(.din(n18739), .dout(n18844));
  jnot g18591(.din(n18732), .dout(n18845));
  jnot g18592(.din(n18724), .dout(n18846));
  jnot g18593(.din(n18717), .dout(n18847));
  jnot g18594(.din(n18709), .dout(n18848));
  jnot g18595(.din(n18701), .dout(n18849));
  jnot g18596(.din(n18693), .dout(n18850));
  jnot g18597(.din(n18685), .dout(n18851));
  jnot g18598(.din(n18677), .dout(n18852));
  jnot g18599(.din(n18670), .dout(n18853));
  jnot g18600(.din(n18662), .dout(n18854));
  jnot g18601(.din(n18654), .dout(n18855));
  jnot g18602(.din(n18646), .dout(n18856));
  jnot g18603(.din(n18639), .dout(n18857));
  jnot g18604(.din(n18631), .dout(n18858));
  jnot g18605(.din(n18624), .dout(n18859));
  jnot g18606(.din(n18616), .dout(n18860));
  jnot g18607(.din(n18609), .dout(n18861));
  jnot g18608(.din(n18601), .dout(n18862));
  jnot g18609(.din(n18594), .dout(n18863));
  jnot g18610(.din(n18586), .dout(n18864));
  jnot g18611(.din(n18578), .dout(n18865));
  jnot g18612(.din(n18570), .dout(n18866));
  jnot g18613(.din(n18563), .dout(n18867));
  jnot g18614(.din(n18555), .dout(n18868));
  jnot g18615(.din(n18548), .dout(n18869));
  jnot g18616(.din(n18540), .dout(n18870));
  jnot g18617(.din(n18533), .dout(n18871));
  jnot g18618(.din(n18526), .dout(n18872));
  jnot g18619(.din(n18518), .dout(n18873));
  jnot g18620(.din(n18510), .dout(n18874));
  jnot g18621(.din(n18503), .dout(n18875));
  jnot g18622(.din(n18495), .dout(n18876));
  jnot g18623(.din(n18488), .dout(n18877));
  jnot g18624(.din(n18480), .dout(n18878));
  jnot g18625(.din(n18473), .dout(n18879));
  jnot g18626(.din(n18465), .dout(n18880));
  jnot g18627(.din(n18458), .dout(n18881));
  jnot g18628(.din(n18447), .dout(n18882));
  jnot g18629(.din(n18190), .dout(n18883));
  jor  g18630(.dina(n18442), .dinb(n17774), .dout(n18884));
  jnot g18631(.din(n18188), .dout(n18885));
  jand g18632(.dina(n18885), .dinb(n18884), .dout(n18886));
  jand g18633(.dina(n18886), .dinb(n17769), .dout(n18887));
  jor  g18634(.dina(n18442), .dinb(a[20] ), .dout(n18888));
  jand g18635(.dina(n18888), .dinb(a[21] ), .dout(n18889));
  jor  g18636(.dina(n18449), .dinb(n18889), .dout(n18890));
  jor  g18637(.dina(n18890), .dinb(n18887), .dout(n18891));
  jand g18638(.dina(n18891), .dinb(n18883), .dout(n18892));
  jand g18639(.dina(n18892), .dinb(n17134), .dout(n18893));
  jor  g18640(.dina(n18454), .dinb(n18893), .dout(n18894));
  jand g18641(.dina(n18894), .dinb(n18882), .dout(n18895));
  jand g18642(.dina(n18895), .dinb(n16489), .dout(n18896));
  jnot g18643(.din(n18462), .dout(n18897));
  jor  g18644(.dina(n18897), .dinb(n18896), .dout(n18898));
  jand g18645(.dina(n18898), .dinb(n18881), .dout(n18899));
  jand g18646(.dina(n18899), .dinb(n15878), .dout(n18900));
  jor  g18647(.dina(n18469), .dinb(n18900), .dout(n18901));
  jand g18648(.dina(n18901), .dinb(n18880), .dout(n18902));
  jand g18649(.dina(n18902), .dinb(n15260), .dout(n18903));
  jnot g18650(.din(n18477), .dout(n18904));
  jor  g18651(.dina(n18904), .dinb(n18903), .dout(n18905));
  jand g18652(.dina(n18905), .dinb(n18879), .dout(n18906));
  jand g18653(.dina(n18906), .dinb(n14674), .dout(n18907));
  jor  g18654(.dina(n18484), .dinb(n18907), .dout(n18908));
  jand g18655(.dina(n18908), .dinb(n18878), .dout(n18909));
  jand g18656(.dina(n18909), .dinb(n14078), .dout(n18910));
  jnot g18657(.din(n18492), .dout(n18911));
  jor  g18658(.dina(n18911), .dinb(n18910), .dout(n18912));
  jand g18659(.dina(n18912), .dinb(n18877), .dout(n18913));
  jand g18660(.dina(n18913), .dinb(n13515), .dout(n18914));
  jor  g18661(.dina(n18499), .dinb(n18914), .dout(n18915));
  jand g18662(.dina(n18915), .dinb(n18876), .dout(n18916));
  jand g18663(.dina(n18916), .dinb(n12947), .dout(n18917));
  jnot g18664(.din(n18507), .dout(n18918));
  jor  g18665(.dina(n18918), .dinb(n18917), .dout(n18919));
  jand g18666(.dina(n18919), .dinb(n18875), .dout(n18920));
  jand g18667(.dina(n18920), .dinb(n12410), .dout(n18921));
  jor  g18668(.dina(n18514), .dinb(n18921), .dout(n18922));
  jand g18669(.dina(n18922), .dinb(n18874), .dout(n18923));
  jand g18670(.dina(n18923), .dinb(n11858), .dout(n18924));
  jor  g18671(.dina(n18522), .dinb(n18924), .dout(n18925));
  jand g18672(.dina(n18925), .dinb(n18873), .dout(n18926));
  jand g18673(.dina(n18926), .dinb(n11347), .dout(n18927));
  jnot g18674(.din(n18530), .dout(n18928));
  jor  g18675(.dina(n18928), .dinb(n18927), .dout(n18929));
  jand g18676(.dina(n18929), .dinb(n18872), .dout(n18930));
  jand g18677(.dina(n18930), .dinb(n10824), .dout(n18931));
  jnot g18678(.din(n18537), .dout(n18932));
  jor  g18679(.dina(n18932), .dinb(n18931), .dout(n18933));
  jand g18680(.dina(n18933), .dinb(n18871), .dout(n18934));
  jand g18681(.dina(n18934), .dinb(n10328), .dout(n18935));
  jor  g18682(.dina(n18544), .dinb(n18935), .dout(n18936));
  jand g18683(.dina(n18936), .dinb(n18870), .dout(n18937));
  jand g18684(.dina(n18937), .dinb(n9832), .dout(n18938));
  jnot g18685(.din(n18552), .dout(n18939));
  jor  g18686(.dina(n18939), .dinb(n18938), .dout(n18940));
  jand g18687(.dina(n18940), .dinb(n18869), .dout(n18941));
  jand g18688(.dina(n18941), .dinb(n9369), .dout(n18942));
  jor  g18689(.dina(n18559), .dinb(n18942), .dout(n18943));
  jand g18690(.dina(n18943), .dinb(n18868), .dout(n18944));
  jand g18691(.dina(n18944), .dinb(n8890), .dout(n18945));
  jnot g18692(.din(n18567), .dout(n18946));
  jor  g18693(.dina(n18946), .dinb(n18945), .dout(n18947));
  jand g18694(.dina(n18947), .dinb(n18867), .dout(n18948));
  jand g18695(.dina(n18948), .dinb(n8449), .dout(n18949));
  jor  g18696(.dina(n18574), .dinb(n18949), .dout(n18950));
  jand g18697(.dina(n18950), .dinb(n18866), .dout(n18951));
  jand g18698(.dina(n18951), .dinb(n8003), .dout(n18952));
  jor  g18699(.dina(n18582), .dinb(n18952), .dout(n18953));
  jand g18700(.dina(n18953), .dinb(n18865), .dout(n18954));
  jand g18701(.dina(n18954), .dinb(n7581), .dout(n18955));
  jor  g18702(.dina(n18590), .dinb(n18955), .dout(n18956));
  jand g18703(.dina(n18956), .dinb(n18864), .dout(n18957));
  jand g18704(.dina(n18957), .dinb(n7154), .dout(n18958));
  jnot g18705(.din(n18598), .dout(n18959));
  jor  g18706(.dina(n18959), .dinb(n18958), .dout(n18960));
  jand g18707(.dina(n18960), .dinb(n18863), .dout(n18961));
  jand g18708(.dina(n18961), .dinb(n6758), .dout(n18962));
  jor  g18709(.dina(n18605), .dinb(n18962), .dout(n18963));
  jand g18710(.dina(n18963), .dinb(n18862), .dout(n18964));
  jand g18711(.dina(n18964), .dinb(n6357), .dout(n18965));
  jnot g18712(.din(n18613), .dout(n18966));
  jor  g18713(.dina(n18966), .dinb(n18965), .dout(n18967));
  jand g18714(.dina(n18967), .dinb(n18861), .dout(n18968));
  jand g18715(.dina(n18968), .dinb(n5989), .dout(n18969));
  jor  g18716(.dina(n18620), .dinb(n18969), .dout(n18970));
  jand g18717(.dina(n18970), .dinb(n18860), .dout(n18971));
  jand g18718(.dina(n18971), .dinb(n5606), .dout(n18972));
  jnot g18719(.din(n18628), .dout(n18973));
  jor  g18720(.dina(n18973), .dinb(n18972), .dout(n18974));
  jand g18721(.dina(n18974), .dinb(n18859), .dout(n18975));
  jand g18722(.dina(n18975), .dinb(n5259), .dout(n18976));
  jor  g18723(.dina(n18635), .dinb(n18976), .dout(n18977));
  jand g18724(.dina(n18977), .dinb(n18858), .dout(n18978));
  jand g18725(.dina(n18978), .dinb(n4902), .dout(n18979));
  jnot g18726(.din(n18643), .dout(n18980));
  jor  g18727(.dina(n18980), .dinb(n18979), .dout(n18981));
  jand g18728(.dina(n18981), .dinb(n18857), .dout(n18982));
  jand g18729(.dina(n18982), .dinb(n4582), .dout(n18983));
  jor  g18730(.dina(n18650), .dinb(n18983), .dout(n18984));
  jand g18731(.dina(n18984), .dinb(n18856), .dout(n18985));
  jand g18732(.dina(n18985), .dinb(n4249), .dout(n18986));
  jor  g18733(.dina(n18658), .dinb(n18986), .dout(n18987));
  jand g18734(.dina(n18987), .dinb(n18855), .dout(n18988));
  jand g18735(.dina(n18988), .dinb(n3955), .dout(n18989));
  jor  g18736(.dina(n18666), .dinb(n18989), .dout(n18990));
  jand g18737(.dina(n18990), .dinb(n18854), .dout(n18991));
  jand g18738(.dina(n18991), .dinb(n3642), .dout(n18992));
  jnot g18739(.din(n18674), .dout(n18993));
  jor  g18740(.dina(n18993), .dinb(n18992), .dout(n18994));
  jand g18741(.dina(n18994), .dinb(n18853), .dout(n18995));
  jand g18742(.dina(n18995), .dinb(n3368), .dout(n18996));
  jor  g18743(.dina(n18681), .dinb(n18996), .dout(n18997));
  jand g18744(.dina(n18997), .dinb(n18852), .dout(n18998));
  jand g18745(.dina(n18998), .dinb(n3089), .dout(n18999));
  jor  g18746(.dina(n18689), .dinb(n18999), .dout(n19000));
  jand g18747(.dina(n19000), .dinb(n18851), .dout(n19001));
  jand g18748(.dina(n19001), .dinb(n2833), .dout(n19002));
  jor  g18749(.dina(n18697), .dinb(n19002), .dout(n19003));
  jand g18750(.dina(n19003), .dinb(n18850), .dout(n19004));
  jand g18751(.dina(n19004), .dinb(n2572), .dout(n19005));
  jor  g18752(.dina(n18705), .dinb(n19005), .dout(n19006));
  jand g18753(.dina(n19006), .dinb(n18849), .dout(n19007));
  jand g18754(.dina(n19007), .dinb(n2345), .dout(n19008));
  jor  g18755(.dina(n18713), .dinb(n19008), .dout(n19009));
  jand g18756(.dina(n19009), .dinb(n18848), .dout(n19010));
  jand g18757(.dina(n19010), .dinb(n2108), .dout(n19011));
  jnot g18758(.din(n18721), .dout(n19012));
  jor  g18759(.dina(n19012), .dinb(n19011), .dout(n19013));
  jand g18760(.dina(n19013), .dinb(n18847), .dout(n19014));
  jand g18761(.dina(n19014), .dinb(n1912), .dout(n19015));
  jor  g18762(.dina(n18728), .dinb(n19015), .dout(n19016));
  jand g18763(.dina(n19016), .dinb(n18846), .dout(n19017));
  jand g18764(.dina(n19017), .dinb(n1699), .dout(n19018));
  jnot g18765(.din(n18736), .dout(n19019));
  jor  g18766(.dina(n19019), .dinb(n19018), .dout(n19020));
  jand g18767(.dina(n19020), .dinb(n18845), .dout(n19021));
  jand g18768(.dina(n19021), .dinb(n1516), .dout(n19022));
  jor  g18769(.dina(n18743), .dinb(n19022), .dout(n19023));
  jand g18770(.dina(n19023), .dinb(n18844), .dout(n19024));
  jand g18771(.dina(n19024), .dinb(n1332), .dout(n19025));
  jor  g18772(.dina(n18751), .dinb(n19025), .dout(n19026));
  jand g18773(.dina(n19026), .dinb(n18843), .dout(n19027));
  jand g18774(.dina(n19027), .dinb(n1173), .dout(n19028));
  jnot g18775(.din(n18759), .dout(n19029));
  jor  g18776(.dina(n19029), .dinb(n19028), .dout(n19030));
  jand g18777(.dina(n19030), .dinb(n18842), .dout(n19031));
  jand g18778(.dina(n19031), .dinb(n1008), .dout(n19032));
  jor  g18779(.dina(n19032), .dinb(n18841), .dout(n19033));
  jand g18780(.dina(n19033), .dinb(n18840), .dout(n19034));
  jand g18781(.dina(n19034), .dinb(n884), .dout(n19035));
  jor  g18782(.dina(n18773), .dinb(n19035), .dout(n19036));
  jand g18783(.dina(n19036), .dinb(n18839), .dout(n19037));
  jand g18784(.dina(n19037), .dinb(n743), .dout(n19038));
  jnot g18785(.din(n18781), .dout(n19039));
  jor  g18786(.dina(n19039), .dinb(n19038), .dout(n19040));
  jand g18787(.dina(n19040), .dinb(n18838), .dout(n19041));
  jand g18788(.dina(n19041), .dinb(n635), .dout(n19042));
  jor  g18789(.dina(n18788), .dinb(n19042), .dout(n19043));
  jand g18790(.dina(n19043), .dinb(n18837), .dout(n19044));
  jand g18791(.dina(n19044), .dinb(n515), .dout(n19045));
  jnot g18792(.din(n18796), .dout(n19046));
  jor  g18793(.dina(n19046), .dinb(n19045), .dout(n19047));
  jand g18794(.dina(n19047), .dinb(n18836), .dout(n19048));
  jand g18795(.dina(n19048), .dinb(n443), .dout(n19049));
  jor  g18796(.dina(n18803), .dinb(n19049), .dout(n19050));
  jand g18797(.dina(n19050), .dinb(n18835), .dout(n19051));
  jand g18798(.dina(n19051), .dinb(n352), .dout(n19052));
  jor  g18799(.dina(n18811), .dinb(n19052), .dout(n19053));
  jand g18800(.dina(n19053), .dinb(n18834), .dout(n19054));
  jand g18801(.dina(n19054), .dinb(n294), .dout(n19055));
  jor  g18802(.dina(n18819), .dinb(n19055), .dout(n19056));
  jand g18803(.dina(n19056), .dinb(n18833), .dout(n19057));
  jand g18804(.dina(n19057), .dinb(n239), .dout(n19058));
  jnot g18805(.din(n18827), .dout(n19059));
  jor  g18806(.dina(n19059), .dinb(n19058), .dout(n19060));
  jand g18807(.dina(n19060), .dinb(n18832), .dout(n19061));
  jand g18808(.dina(n19061), .dinb(n221), .dout(n19062));
  jxor g18809(.dina(n18148), .dinb(n239), .dout(n19063));
  jand g18810(.dina(n19063), .dinb(asqrt[10] ), .dout(n19064));
  jxor g18811(.dina(n19064), .dinb(n18153), .dout(n19065));
  jor  g18812(.dina(n19065), .dinb(n19062), .dout(n19066));
  jand g18813(.dina(n19066), .dinb(n18831), .dout(n19067));
  jor  g18814(.dina(n19067), .dinb(n18183), .dout(n19068));
  jand g18815(.dina(n18178), .dinb(n18435), .dout(n19069));
  jor  g18816(.dina(n19069), .dinb(n18164), .dout(n19070));
  jor  g18817(.dina(n19070), .dinb(n19068), .dout(n19071));
  jand g18818(.dina(n19071), .dinb(n218), .dout(n19072));
  jand g18819(.dina(n18442), .dinb(n17773), .dout(n19073));
  jand g18820(.dina(n19067), .dinb(n18183), .dout(n19074));
  jor  g18821(.dina(n19074), .dinb(n19073), .dout(n19075));
  jand g18822(.dina(n18441), .dinb(n18163), .dout(n19076));
  jnot g18823(.din(n19076), .dout(n19077));
  jand g18824(.dina(n18172), .dinb(asqrt[63] ), .dout(n19078));
  jand g18825(.dina(n19078), .dinb(n18195), .dout(n19079));
  jand g18826(.dina(n19079), .dinb(n19077), .dout(n19080));
  jor  g18827(.dina(n19080), .dinb(n19075), .dout(n19081));
  jor  g18828(.dina(n19081), .dinb(n19072), .dout(asqrt[9] ));
  jor  g18829(.dina(n18829), .dinb(asqrt[62] ), .dout(n19083));
  jnot g18830(.din(n19065), .dout(n19084));
  jand g18831(.dina(n19084), .dinb(n19083), .dout(n19085));
  jor  g18832(.dina(n19085), .dinb(n18830), .dout(n19086));
  jand g18833(.dina(n19086), .dinb(n18182), .dout(n19087));
  jnot g18834(.din(n19070), .dout(n19088));
  jand g18835(.dina(n19088), .dinb(n19087), .dout(n19089));
  jor  g18836(.dina(n19089), .dinb(asqrt[63] ), .dout(n19090));
  jnot g18837(.din(n19073), .dout(n19091));
  jor  g18838(.dina(n19086), .dinb(n18182), .dout(n19092));
  jand g18839(.dina(n19092), .dinb(n19091), .dout(n19093));
  jnot g18840(.din(n19080), .dout(n19094));
  jand g18841(.dina(n19094), .dinb(n19093), .dout(n19095));
  jand g18842(.dina(n19095), .dinb(n19090), .dout(n19096));
  jxor g18843(.dina(n18829), .dinb(n221), .dout(n19097));
  jor  g18844(.dina(n19097), .dinb(n19096), .dout(n19098));
  jxor g18845(.dina(n19098), .dinb(n19065), .dout(n19099));
  jnot g18846(.din(n19099), .dout(n19100));
  jnot g18847(.din(a[16] ), .dout(n19101));
  jnot g18848(.din(a[17] ), .dout(n19102));
  jand g18849(.dina(n19102), .dinb(n19101), .dout(n19103));
  jand g18850(.dina(n19103), .dinb(n18185), .dout(n19104));
  jnot g18851(.din(n19104), .dout(n19105));
  jor  g18852(.dina(n19096), .dinb(n18185), .dout(n19106));
  jand g18853(.dina(n19106), .dinb(n19105), .dout(n19107));
  jor  g18854(.dina(n19107), .dinb(n18442), .dout(n19108));
  jand g18855(.dina(n19107), .dinb(n18442), .dout(n19109));
  jor  g18856(.dina(n19096), .dinb(a[18] ), .dout(n19110));
  jand g18857(.dina(n19110), .dinb(a[19] ), .dout(n19111));
  jand g18858(.dina(asqrt[9] ), .dinb(n18187), .dout(n19112));
  jor  g18859(.dina(n19112), .dinb(n19111), .dout(n19113));
  jor  g18860(.dina(n19113), .dinb(n19109), .dout(n19114));
  jand g18861(.dina(n19114), .dinb(n19108), .dout(n19115));
  jor  g18862(.dina(n19115), .dinb(n17769), .dout(n19116));
  jand g18863(.dina(n19115), .dinb(n17769), .dout(n19117));
  jnot g18864(.din(n18187), .dout(n19118));
  jor  g18865(.dina(n19096), .dinb(n19118), .dout(n19119));
  jor  g18866(.dina(n19079), .dinb(n18442), .dout(n19120));
  jor  g18867(.dina(n19120), .dinb(n19074), .dout(n19121));
  jor  g18868(.dina(n19121), .dinb(n19072), .dout(n19122));
  jand g18869(.dina(n19122), .dinb(n19119), .dout(n19123));
  jxor g18870(.dina(n19123), .dinb(n17774), .dout(n19124));
  jor  g18871(.dina(n19124), .dinb(n19117), .dout(n19125));
  jand g18872(.dina(n19125), .dinb(n19116), .dout(n19126));
  jor  g18873(.dina(n19126), .dinb(n17134), .dout(n19127));
  jand g18874(.dina(n19126), .dinb(n17134), .dout(n19128));
  jxor g18875(.dina(n18189), .dinb(n17769), .dout(n19129));
  jor  g18876(.dina(n19129), .dinb(n19096), .dout(n19130));
  jxor g18877(.dina(n19130), .dinb(n18890), .dout(n19131));
  jnot g18878(.din(n19131), .dout(n19132));
  jor  g18879(.dina(n19132), .dinb(n19128), .dout(n19133));
  jand g18880(.dina(n19133), .dinb(n19127), .dout(n19134));
  jor  g18881(.dina(n19134), .dinb(n16489), .dout(n19135));
  jand g18882(.dina(n19134), .dinb(n16489), .dout(n19136));
  jxor g18883(.dina(n18446), .dinb(n17134), .dout(n19137));
  jor  g18884(.dina(n19137), .dinb(n19096), .dout(n19138));
  jxor g18885(.dina(n19138), .dinb(n18455), .dout(n19139));
  jor  g18886(.dina(n19139), .dinb(n19136), .dout(n19140));
  jand g18887(.dina(n19140), .dinb(n19135), .dout(n19141));
  jor  g18888(.dina(n19141), .dinb(n15878), .dout(n19142));
  jand g18889(.dina(n19141), .dinb(n15878), .dout(n19143));
  jxor g18890(.dina(n18457), .dinb(n16489), .dout(n19144));
  jor  g18891(.dina(n19144), .dinb(n19096), .dout(n19145));
  jxor g18892(.dina(n19145), .dinb(n18897), .dout(n19146));
  jnot g18893(.din(n19146), .dout(n19147));
  jor  g18894(.dina(n19147), .dinb(n19143), .dout(n19148));
  jand g18895(.dina(n19148), .dinb(n19142), .dout(n19149));
  jor  g18896(.dina(n19149), .dinb(n15260), .dout(n19150));
  jand g18897(.dina(n19149), .dinb(n15260), .dout(n19151));
  jxor g18898(.dina(n18464), .dinb(n15878), .dout(n19152));
  jor  g18899(.dina(n19152), .dinb(n19096), .dout(n19153));
  jxor g18900(.dina(n19153), .dinb(n18470), .dout(n19154));
  jor  g18901(.dina(n19154), .dinb(n19151), .dout(n19155));
  jand g18902(.dina(n19155), .dinb(n19150), .dout(n19156));
  jor  g18903(.dina(n19156), .dinb(n14674), .dout(n19157));
  jand g18904(.dina(n19156), .dinb(n14674), .dout(n19158));
  jxor g18905(.dina(n18472), .dinb(n15260), .dout(n19159));
  jor  g18906(.dina(n19159), .dinb(n19096), .dout(n19160));
  jxor g18907(.dina(n19160), .dinb(n18904), .dout(n19161));
  jnot g18908(.din(n19161), .dout(n19162));
  jor  g18909(.dina(n19162), .dinb(n19158), .dout(n19163));
  jand g18910(.dina(n19163), .dinb(n19157), .dout(n19164));
  jor  g18911(.dina(n19164), .dinb(n14078), .dout(n19165));
  jand g18912(.dina(n19164), .dinb(n14078), .dout(n19166));
  jxor g18913(.dina(n18479), .dinb(n14674), .dout(n19167));
  jor  g18914(.dina(n19167), .dinb(n19096), .dout(n19168));
  jxor g18915(.dina(n19168), .dinb(n18485), .dout(n19169));
  jor  g18916(.dina(n19169), .dinb(n19166), .dout(n19170));
  jand g18917(.dina(n19170), .dinb(n19165), .dout(n19171));
  jor  g18918(.dina(n19171), .dinb(n13515), .dout(n19172));
  jand g18919(.dina(n19171), .dinb(n13515), .dout(n19173));
  jxor g18920(.dina(n18487), .dinb(n14078), .dout(n19174));
  jor  g18921(.dina(n19174), .dinb(n19096), .dout(n19175));
  jxor g18922(.dina(n19175), .dinb(n18911), .dout(n19176));
  jnot g18923(.din(n19176), .dout(n19177));
  jor  g18924(.dina(n19177), .dinb(n19173), .dout(n19178));
  jand g18925(.dina(n19178), .dinb(n19172), .dout(n19179));
  jor  g18926(.dina(n19179), .dinb(n12947), .dout(n19180));
  jand g18927(.dina(n19179), .dinb(n12947), .dout(n19181));
  jxor g18928(.dina(n18494), .dinb(n13515), .dout(n19182));
  jor  g18929(.dina(n19182), .dinb(n19096), .dout(n19183));
  jxor g18930(.dina(n19183), .dinb(n18500), .dout(n19184));
  jor  g18931(.dina(n19184), .dinb(n19181), .dout(n19185));
  jand g18932(.dina(n19185), .dinb(n19180), .dout(n19186));
  jor  g18933(.dina(n19186), .dinb(n12410), .dout(n19187));
  jand g18934(.dina(n19186), .dinb(n12410), .dout(n19188));
  jxor g18935(.dina(n18502), .dinb(n12947), .dout(n19189));
  jor  g18936(.dina(n19189), .dinb(n19096), .dout(n19190));
  jxor g18937(.dina(n19190), .dinb(n18918), .dout(n19191));
  jnot g18938(.din(n19191), .dout(n19192));
  jor  g18939(.dina(n19192), .dinb(n19188), .dout(n19193));
  jand g18940(.dina(n19193), .dinb(n19187), .dout(n19194));
  jor  g18941(.dina(n19194), .dinb(n11858), .dout(n19195));
  jand g18942(.dina(n19194), .dinb(n11858), .dout(n19196));
  jxor g18943(.dina(n18509), .dinb(n12410), .dout(n19197));
  jor  g18944(.dina(n19197), .dinb(n19096), .dout(n19198));
  jxor g18945(.dina(n19198), .dinb(n18515), .dout(n19199));
  jor  g18946(.dina(n19199), .dinb(n19196), .dout(n19200));
  jand g18947(.dina(n19200), .dinb(n19195), .dout(n19201));
  jor  g18948(.dina(n19201), .dinb(n11347), .dout(n19202));
  jand g18949(.dina(n19201), .dinb(n11347), .dout(n19203));
  jxor g18950(.dina(n18517), .dinb(n11858), .dout(n19204));
  jor  g18951(.dina(n19204), .dinb(n19096), .dout(n19205));
  jxor g18952(.dina(n19205), .dinb(n18523), .dout(n19206));
  jor  g18953(.dina(n19206), .dinb(n19203), .dout(n19207));
  jand g18954(.dina(n19207), .dinb(n19202), .dout(n19208));
  jor  g18955(.dina(n19208), .dinb(n10824), .dout(n19209));
  jand g18956(.dina(n19208), .dinb(n10824), .dout(n19210));
  jxor g18957(.dina(n18525), .dinb(n11347), .dout(n19211));
  jor  g18958(.dina(n19211), .dinb(n19096), .dout(n19212));
  jxor g18959(.dina(n19212), .dinb(n18928), .dout(n19213));
  jnot g18960(.din(n19213), .dout(n19214));
  jor  g18961(.dina(n19214), .dinb(n19210), .dout(n19215));
  jand g18962(.dina(n19215), .dinb(n19209), .dout(n19216));
  jor  g18963(.dina(n19216), .dinb(n10328), .dout(n19217));
  jand g18964(.dina(n19216), .dinb(n10328), .dout(n19218));
  jxor g18965(.dina(n18532), .dinb(n10824), .dout(n19219));
  jor  g18966(.dina(n19219), .dinb(n19096), .dout(n19220));
  jxor g18967(.dina(n19220), .dinb(n18932), .dout(n19221));
  jnot g18968(.din(n19221), .dout(n19222));
  jor  g18969(.dina(n19222), .dinb(n19218), .dout(n19223));
  jand g18970(.dina(n19223), .dinb(n19217), .dout(n19224));
  jor  g18971(.dina(n19224), .dinb(n9832), .dout(n19225));
  jand g18972(.dina(n19224), .dinb(n9832), .dout(n19226));
  jxor g18973(.dina(n18539), .dinb(n10328), .dout(n19227));
  jor  g18974(.dina(n19227), .dinb(n19096), .dout(n19228));
  jxor g18975(.dina(n19228), .dinb(n18545), .dout(n19229));
  jor  g18976(.dina(n19229), .dinb(n19226), .dout(n19230));
  jand g18977(.dina(n19230), .dinb(n19225), .dout(n19231));
  jor  g18978(.dina(n19231), .dinb(n9369), .dout(n19232));
  jand g18979(.dina(n19231), .dinb(n9369), .dout(n19233));
  jxor g18980(.dina(n18547), .dinb(n9832), .dout(n19234));
  jor  g18981(.dina(n19234), .dinb(n19096), .dout(n19235));
  jxor g18982(.dina(n19235), .dinb(n18939), .dout(n19236));
  jnot g18983(.din(n19236), .dout(n19237));
  jor  g18984(.dina(n19237), .dinb(n19233), .dout(n19238));
  jand g18985(.dina(n19238), .dinb(n19232), .dout(n19239));
  jor  g18986(.dina(n19239), .dinb(n8890), .dout(n19240));
  jand g18987(.dina(n19239), .dinb(n8890), .dout(n19241));
  jxor g18988(.dina(n18554), .dinb(n9369), .dout(n19242));
  jor  g18989(.dina(n19242), .dinb(n19096), .dout(n19243));
  jxor g18990(.dina(n19243), .dinb(n18560), .dout(n19244));
  jor  g18991(.dina(n19244), .dinb(n19241), .dout(n19245));
  jand g18992(.dina(n19245), .dinb(n19240), .dout(n19246));
  jor  g18993(.dina(n19246), .dinb(n8449), .dout(n19247));
  jand g18994(.dina(n19246), .dinb(n8449), .dout(n19248));
  jxor g18995(.dina(n18562), .dinb(n8890), .dout(n19249));
  jor  g18996(.dina(n19249), .dinb(n19096), .dout(n19250));
  jxor g18997(.dina(n19250), .dinb(n18946), .dout(n19251));
  jnot g18998(.din(n19251), .dout(n19252));
  jor  g18999(.dina(n19252), .dinb(n19248), .dout(n19253));
  jand g19000(.dina(n19253), .dinb(n19247), .dout(n19254));
  jor  g19001(.dina(n19254), .dinb(n8003), .dout(n19255));
  jand g19002(.dina(n19254), .dinb(n8003), .dout(n19256));
  jxor g19003(.dina(n18569), .dinb(n8449), .dout(n19257));
  jor  g19004(.dina(n19257), .dinb(n19096), .dout(n19258));
  jxor g19005(.dina(n19258), .dinb(n18575), .dout(n19259));
  jor  g19006(.dina(n19259), .dinb(n19256), .dout(n19260));
  jand g19007(.dina(n19260), .dinb(n19255), .dout(n19261));
  jor  g19008(.dina(n19261), .dinb(n7581), .dout(n19262));
  jand g19009(.dina(n19261), .dinb(n7581), .dout(n19263));
  jxor g19010(.dina(n18577), .dinb(n8003), .dout(n19264));
  jor  g19011(.dina(n19264), .dinb(n19096), .dout(n19265));
  jxor g19012(.dina(n19265), .dinb(n18583), .dout(n19266));
  jor  g19013(.dina(n19266), .dinb(n19263), .dout(n19267));
  jand g19014(.dina(n19267), .dinb(n19262), .dout(n19268));
  jor  g19015(.dina(n19268), .dinb(n7154), .dout(n19269));
  jand g19016(.dina(n19268), .dinb(n7154), .dout(n19270));
  jxor g19017(.dina(n18585), .dinb(n7581), .dout(n19271));
  jor  g19018(.dina(n19271), .dinb(n19096), .dout(n19272));
  jxor g19019(.dina(n19272), .dinb(n18591), .dout(n19273));
  jor  g19020(.dina(n19273), .dinb(n19270), .dout(n19274));
  jand g19021(.dina(n19274), .dinb(n19269), .dout(n19275));
  jor  g19022(.dina(n19275), .dinb(n6758), .dout(n19276));
  jand g19023(.dina(n19275), .dinb(n6758), .dout(n19277));
  jxor g19024(.dina(n18593), .dinb(n7154), .dout(n19278));
  jor  g19025(.dina(n19278), .dinb(n19096), .dout(n19279));
  jxor g19026(.dina(n19279), .dinb(n18959), .dout(n19280));
  jnot g19027(.din(n19280), .dout(n19281));
  jor  g19028(.dina(n19281), .dinb(n19277), .dout(n19282));
  jand g19029(.dina(n19282), .dinb(n19276), .dout(n19283));
  jor  g19030(.dina(n19283), .dinb(n6357), .dout(n19284));
  jand g19031(.dina(n19283), .dinb(n6357), .dout(n19285));
  jxor g19032(.dina(n18600), .dinb(n6758), .dout(n19286));
  jor  g19033(.dina(n19286), .dinb(n19096), .dout(n19287));
  jxor g19034(.dina(n19287), .dinb(n18606), .dout(n19288));
  jor  g19035(.dina(n19288), .dinb(n19285), .dout(n19289));
  jand g19036(.dina(n19289), .dinb(n19284), .dout(n19290));
  jor  g19037(.dina(n19290), .dinb(n5989), .dout(n19291));
  jand g19038(.dina(n19290), .dinb(n5989), .dout(n19292));
  jxor g19039(.dina(n18608), .dinb(n6357), .dout(n19293));
  jor  g19040(.dina(n19293), .dinb(n19096), .dout(n19294));
  jxor g19041(.dina(n19294), .dinb(n18966), .dout(n19295));
  jnot g19042(.din(n19295), .dout(n19296));
  jor  g19043(.dina(n19296), .dinb(n19292), .dout(n19297));
  jand g19044(.dina(n19297), .dinb(n19291), .dout(n19298));
  jor  g19045(.dina(n19298), .dinb(n5606), .dout(n19299));
  jand g19046(.dina(n19298), .dinb(n5606), .dout(n19300));
  jxor g19047(.dina(n18615), .dinb(n5989), .dout(n19301));
  jor  g19048(.dina(n19301), .dinb(n19096), .dout(n19302));
  jxor g19049(.dina(n19302), .dinb(n18621), .dout(n19303));
  jor  g19050(.dina(n19303), .dinb(n19300), .dout(n19304));
  jand g19051(.dina(n19304), .dinb(n19299), .dout(n19305));
  jor  g19052(.dina(n19305), .dinb(n5259), .dout(n19306));
  jand g19053(.dina(n19305), .dinb(n5259), .dout(n19307));
  jxor g19054(.dina(n18623), .dinb(n5606), .dout(n19308));
  jor  g19055(.dina(n19308), .dinb(n19096), .dout(n19309));
  jxor g19056(.dina(n19309), .dinb(n18973), .dout(n19310));
  jnot g19057(.din(n19310), .dout(n19311));
  jor  g19058(.dina(n19311), .dinb(n19307), .dout(n19312));
  jand g19059(.dina(n19312), .dinb(n19306), .dout(n19313));
  jor  g19060(.dina(n19313), .dinb(n4902), .dout(n19314));
  jand g19061(.dina(n19313), .dinb(n4902), .dout(n19315));
  jxor g19062(.dina(n18630), .dinb(n5259), .dout(n19316));
  jor  g19063(.dina(n19316), .dinb(n19096), .dout(n19317));
  jxor g19064(.dina(n19317), .dinb(n18636), .dout(n19318));
  jor  g19065(.dina(n19318), .dinb(n19315), .dout(n19319));
  jand g19066(.dina(n19319), .dinb(n19314), .dout(n19320));
  jor  g19067(.dina(n19320), .dinb(n4582), .dout(n19321));
  jand g19068(.dina(n19320), .dinb(n4582), .dout(n19322));
  jxor g19069(.dina(n18638), .dinb(n4902), .dout(n19323));
  jor  g19070(.dina(n19323), .dinb(n19096), .dout(n19324));
  jxor g19071(.dina(n19324), .dinb(n18980), .dout(n19325));
  jnot g19072(.din(n19325), .dout(n19326));
  jor  g19073(.dina(n19326), .dinb(n19322), .dout(n19327));
  jand g19074(.dina(n19327), .dinb(n19321), .dout(n19328));
  jor  g19075(.dina(n19328), .dinb(n4249), .dout(n19329));
  jand g19076(.dina(n19328), .dinb(n4249), .dout(n19330));
  jxor g19077(.dina(n18645), .dinb(n4582), .dout(n19331));
  jor  g19078(.dina(n19331), .dinb(n19096), .dout(n19332));
  jxor g19079(.dina(n19332), .dinb(n18651), .dout(n19333));
  jor  g19080(.dina(n19333), .dinb(n19330), .dout(n19334));
  jand g19081(.dina(n19334), .dinb(n19329), .dout(n19335));
  jor  g19082(.dina(n19335), .dinb(n3955), .dout(n19336));
  jand g19083(.dina(n19335), .dinb(n3955), .dout(n19337));
  jxor g19084(.dina(n18653), .dinb(n4249), .dout(n19338));
  jor  g19085(.dina(n19338), .dinb(n19096), .dout(n19339));
  jxor g19086(.dina(n19339), .dinb(n18659), .dout(n19340));
  jor  g19087(.dina(n19340), .dinb(n19337), .dout(n19341));
  jand g19088(.dina(n19341), .dinb(n19336), .dout(n19342));
  jor  g19089(.dina(n19342), .dinb(n3642), .dout(n19343));
  jand g19090(.dina(n19342), .dinb(n3642), .dout(n19344));
  jxor g19091(.dina(n18661), .dinb(n3955), .dout(n19345));
  jor  g19092(.dina(n19345), .dinb(n19096), .dout(n19346));
  jxor g19093(.dina(n19346), .dinb(n18667), .dout(n19347));
  jor  g19094(.dina(n19347), .dinb(n19344), .dout(n19348));
  jand g19095(.dina(n19348), .dinb(n19343), .dout(n19349));
  jor  g19096(.dina(n19349), .dinb(n3368), .dout(n19350));
  jand g19097(.dina(n19349), .dinb(n3368), .dout(n19351));
  jxor g19098(.dina(n18669), .dinb(n3642), .dout(n19352));
  jor  g19099(.dina(n19352), .dinb(n19096), .dout(n19353));
  jxor g19100(.dina(n19353), .dinb(n18993), .dout(n19354));
  jnot g19101(.din(n19354), .dout(n19355));
  jor  g19102(.dina(n19355), .dinb(n19351), .dout(n19356));
  jand g19103(.dina(n19356), .dinb(n19350), .dout(n19357));
  jor  g19104(.dina(n19357), .dinb(n3089), .dout(n19358));
  jand g19105(.dina(n19357), .dinb(n3089), .dout(n19359));
  jxor g19106(.dina(n18676), .dinb(n3368), .dout(n19360));
  jor  g19107(.dina(n19360), .dinb(n19096), .dout(n19361));
  jxor g19108(.dina(n19361), .dinb(n18682), .dout(n19362));
  jor  g19109(.dina(n19362), .dinb(n19359), .dout(n19363));
  jand g19110(.dina(n19363), .dinb(n19358), .dout(n19364));
  jor  g19111(.dina(n19364), .dinb(n2833), .dout(n19365));
  jand g19112(.dina(n19364), .dinb(n2833), .dout(n19366));
  jxor g19113(.dina(n18684), .dinb(n3089), .dout(n19367));
  jor  g19114(.dina(n19367), .dinb(n19096), .dout(n19368));
  jxor g19115(.dina(n19368), .dinb(n18690), .dout(n19369));
  jor  g19116(.dina(n19369), .dinb(n19366), .dout(n19370));
  jand g19117(.dina(n19370), .dinb(n19365), .dout(n19371));
  jor  g19118(.dina(n19371), .dinb(n2572), .dout(n19372));
  jand g19119(.dina(n19371), .dinb(n2572), .dout(n19373));
  jxor g19120(.dina(n18692), .dinb(n2833), .dout(n19374));
  jor  g19121(.dina(n19374), .dinb(n19096), .dout(n19375));
  jxor g19122(.dina(n19375), .dinb(n18698), .dout(n19376));
  jor  g19123(.dina(n19376), .dinb(n19373), .dout(n19377));
  jand g19124(.dina(n19377), .dinb(n19372), .dout(n19378));
  jor  g19125(.dina(n19378), .dinb(n2345), .dout(n19379));
  jand g19126(.dina(n19378), .dinb(n2345), .dout(n19380));
  jxor g19127(.dina(n18700), .dinb(n2572), .dout(n19381));
  jor  g19128(.dina(n19381), .dinb(n19096), .dout(n19382));
  jxor g19129(.dina(n19382), .dinb(n18706), .dout(n19383));
  jor  g19130(.dina(n19383), .dinb(n19380), .dout(n19384));
  jand g19131(.dina(n19384), .dinb(n19379), .dout(n19385));
  jor  g19132(.dina(n19385), .dinb(n2108), .dout(n19386));
  jand g19133(.dina(n19385), .dinb(n2108), .dout(n19387));
  jxor g19134(.dina(n18708), .dinb(n2345), .dout(n19388));
  jor  g19135(.dina(n19388), .dinb(n19096), .dout(n19389));
  jxor g19136(.dina(n19389), .dinb(n18714), .dout(n19390));
  jor  g19137(.dina(n19390), .dinb(n19387), .dout(n19391));
  jand g19138(.dina(n19391), .dinb(n19386), .dout(n19392));
  jor  g19139(.dina(n19392), .dinb(n1912), .dout(n19393));
  jand g19140(.dina(n19392), .dinb(n1912), .dout(n19394));
  jxor g19141(.dina(n18716), .dinb(n2108), .dout(n19395));
  jor  g19142(.dina(n19395), .dinb(n19096), .dout(n19396));
  jxor g19143(.dina(n19396), .dinb(n19012), .dout(n19397));
  jnot g19144(.din(n19397), .dout(n19398));
  jor  g19145(.dina(n19398), .dinb(n19394), .dout(n19399));
  jand g19146(.dina(n19399), .dinb(n19393), .dout(n19400));
  jor  g19147(.dina(n19400), .dinb(n1699), .dout(n19401));
  jand g19148(.dina(n19400), .dinb(n1699), .dout(n19402));
  jxor g19149(.dina(n18723), .dinb(n1912), .dout(n19403));
  jor  g19150(.dina(n19403), .dinb(n19096), .dout(n19404));
  jxor g19151(.dina(n19404), .dinb(n18729), .dout(n19405));
  jor  g19152(.dina(n19405), .dinb(n19402), .dout(n19406));
  jand g19153(.dina(n19406), .dinb(n19401), .dout(n19407));
  jor  g19154(.dina(n19407), .dinb(n1516), .dout(n19408));
  jand g19155(.dina(n19407), .dinb(n1516), .dout(n19409));
  jxor g19156(.dina(n18731), .dinb(n1699), .dout(n19410));
  jor  g19157(.dina(n19410), .dinb(n19096), .dout(n19411));
  jxor g19158(.dina(n19411), .dinb(n19019), .dout(n19412));
  jnot g19159(.din(n19412), .dout(n19413));
  jor  g19160(.dina(n19413), .dinb(n19409), .dout(n19414));
  jand g19161(.dina(n19414), .dinb(n19408), .dout(n19415));
  jor  g19162(.dina(n19415), .dinb(n1332), .dout(n19416));
  jand g19163(.dina(n19415), .dinb(n1332), .dout(n19417));
  jxor g19164(.dina(n18738), .dinb(n1516), .dout(n19418));
  jor  g19165(.dina(n19418), .dinb(n19096), .dout(n19419));
  jxor g19166(.dina(n19419), .dinb(n18744), .dout(n19420));
  jor  g19167(.dina(n19420), .dinb(n19417), .dout(n19421));
  jand g19168(.dina(n19421), .dinb(n19416), .dout(n19422));
  jor  g19169(.dina(n19422), .dinb(n1173), .dout(n19423));
  jand g19170(.dina(n19422), .dinb(n1173), .dout(n19424));
  jxor g19171(.dina(n18746), .dinb(n1332), .dout(n19425));
  jor  g19172(.dina(n19425), .dinb(n19096), .dout(n19426));
  jxor g19173(.dina(n19426), .dinb(n18752), .dout(n19427));
  jor  g19174(.dina(n19427), .dinb(n19424), .dout(n19428));
  jand g19175(.dina(n19428), .dinb(n19423), .dout(n19429));
  jor  g19176(.dina(n19429), .dinb(n1008), .dout(n19430));
  jand g19177(.dina(n19429), .dinb(n1008), .dout(n19431));
  jxor g19178(.dina(n18754), .dinb(n1173), .dout(n19432));
  jor  g19179(.dina(n19432), .dinb(n19096), .dout(n19433));
  jxor g19180(.dina(n19433), .dinb(n19029), .dout(n19434));
  jnot g19181(.din(n19434), .dout(n19435));
  jor  g19182(.dina(n19435), .dinb(n19431), .dout(n19436));
  jand g19183(.dina(n19436), .dinb(n19430), .dout(n19437));
  jor  g19184(.dina(n19437), .dinb(n884), .dout(n19438));
  jxor g19185(.dina(n18761), .dinb(n1008), .dout(n19439));
  jor  g19186(.dina(n19439), .dinb(n19096), .dout(n19440));
  jxor g19187(.dina(n19440), .dinb(n18841), .dout(n19441));
  jnot g19188(.din(n19441), .dout(n19442));
  jand g19189(.dina(n19437), .dinb(n884), .dout(n19443));
  jor  g19190(.dina(n19443), .dinb(n19442), .dout(n19444));
  jand g19191(.dina(n19444), .dinb(n19438), .dout(n19445));
  jor  g19192(.dina(n19445), .dinb(n743), .dout(n19446));
  jand g19193(.dina(n19445), .dinb(n743), .dout(n19447));
  jxor g19194(.dina(n18768), .dinb(n884), .dout(n19448));
  jor  g19195(.dina(n19448), .dinb(n19096), .dout(n19449));
  jxor g19196(.dina(n19449), .dinb(n18774), .dout(n19450));
  jor  g19197(.dina(n19450), .dinb(n19447), .dout(n19451));
  jand g19198(.dina(n19451), .dinb(n19446), .dout(n19452));
  jor  g19199(.dina(n19452), .dinb(n635), .dout(n19453));
  jand g19200(.dina(n19452), .dinb(n635), .dout(n19454));
  jxor g19201(.dina(n18776), .dinb(n743), .dout(n19455));
  jor  g19202(.dina(n19455), .dinb(n19096), .dout(n19456));
  jxor g19203(.dina(n19456), .dinb(n19039), .dout(n19457));
  jnot g19204(.din(n19457), .dout(n19458));
  jor  g19205(.dina(n19458), .dinb(n19454), .dout(n19459));
  jand g19206(.dina(n19459), .dinb(n19453), .dout(n19460));
  jor  g19207(.dina(n19460), .dinb(n515), .dout(n19461));
  jand g19208(.dina(n19460), .dinb(n515), .dout(n19462));
  jxor g19209(.dina(n18783), .dinb(n635), .dout(n19463));
  jor  g19210(.dina(n19463), .dinb(n19096), .dout(n19464));
  jxor g19211(.dina(n19464), .dinb(n18789), .dout(n19465));
  jor  g19212(.dina(n19465), .dinb(n19462), .dout(n19466));
  jand g19213(.dina(n19466), .dinb(n19461), .dout(n19467));
  jor  g19214(.dina(n19467), .dinb(n443), .dout(n19468));
  jand g19215(.dina(n19467), .dinb(n443), .dout(n19469));
  jxor g19216(.dina(n18791), .dinb(n515), .dout(n19470));
  jor  g19217(.dina(n19470), .dinb(n19096), .dout(n19471));
  jxor g19218(.dina(n19471), .dinb(n19046), .dout(n19472));
  jnot g19219(.din(n19472), .dout(n19473));
  jor  g19220(.dina(n19473), .dinb(n19469), .dout(n19474));
  jand g19221(.dina(n19474), .dinb(n19468), .dout(n19475));
  jor  g19222(.dina(n19475), .dinb(n352), .dout(n19476));
  jand g19223(.dina(n19475), .dinb(n352), .dout(n19477));
  jxor g19224(.dina(n18798), .dinb(n443), .dout(n19478));
  jor  g19225(.dina(n19478), .dinb(n19096), .dout(n19479));
  jxor g19226(.dina(n19479), .dinb(n18803), .dout(n19480));
  jnot g19227(.din(n19480), .dout(n19481));
  jor  g19228(.dina(n19481), .dinb(n19477), .dout(n19482));
  jand g19229(.dina(n19482), .dinb(n19476), .dout(n19483));
  jor  g19230(.dina(n19483), .dinb(n294), .dout(n19484));
  jand g19231(.dina(n19483), .dinb(n294), .dout(n19485));
  jxor g19232(.dina(n18806), .dinb(n352), .dout(n19486));
  jor  g19233(.dina(n19486), .dinb(n19096), .dout(n19487));
  jxor g19234(.dina(n19487), .dinb(n18812), .dout(n19488));
  jor  g19235(.dina(n19488), .dinb(n19485), .dout(n19489));
  jand g19236(.dina(n19489), .dinb(n19484), .dout(n19490));
  jor  g19237(.dina(n19490), .dinb(n239), .dout(n19491));
  jand g19238(.dina(n19490), .dinb(n239), .dout(n19492));
  jxor g19239(.dina(n18814), .dinb(n294), .dout(n19493));
  jor  g19240(.dina(n19493), .dinb(n19096), .dout(n19494));
  jxor g19241(.dina(n19494), .dinb(n18820), .dout(n19495));
  jor  g19242(.dina(n19495), .dinb(n19492), .dout(n19496));
  jand g19243(.dina(n19496), .dinb(n19491), .dout(n19497));
  jor  g19244(.dina(n19497), .dinb(n221), .dout(n19498));
  jand g19245(.dina(n19497), .dinb(n221), .dout(n19499));
  jxor g19246(.dina(n18822), .dinb(n239), .dout(n19500));
  jor  g19247(.dina(n19500), .dinb(n19096), .dout(n19501));
  jxor g19248(.dina(n19501), .dinb(n19059), .dout(n19502));
  jnot g19249(.din(n19502), .dout(n19503));
  jor  g19250(.dina(n19503), .dinb(n19499), .dout(n19504));
  jand g19251(.dina(n19504), .dinb(n19498), .dout(n19505));
  jor  g19252(.dina(n19505), .dinb(n19100), .dout(n19506));
  jand g19253(.dina(asqrt[9] ), .dinb(n19087), .dout(n19507));
  jor  g19254(.dina(n19507), .dinb(n19074), .dout(n19508));
  jor  g19255(.dina(n19508), .dinb(n19506), .dout(n19509));
  jand g19256(.dina(n19509), .dinb(n218), .dout(n19510));
  jand g19257(.dina(n19505), .dinb(n19100), .dout(n19511));
  jand g19258(.dina(asqrt[9] ), .dinb(n18182), .dout(n19512));
  jor  g19259(.dina(n19512), .dinb(n19086), .dout(n19513));
  jand g19260(.dina(n19513), .dinb(n19068), .dout(n19514));
  jand g19261(.dina(n19514), .dinb(asqrt[63] ), .dout(n19515));
  jor  g19262(.dina(n19515), .dinb(n19511), .dout(n19516));
  jor  g19263(.dina(n19516), .dinb(n19510), .dout(asqrt[8] ));
  jxor g19264(.dina(n19497), .dinb(n221), .dout(n19520));
  jand g19265(.dina(n19520), .dinb(asqrt[8] ), .dout(n19521));
  jxor g19266(.dina(n19521), .dinb(n19502), .dout(n19522));
  jnot g19267(.din(n19522), .dout(n19523));
  jnot g19268(.din(a[14] ), .dout(n19524));
  jnot g19269(.din(a[15] ), .dout(n19525));
  jand g19270(.dina(n19525), .dinb(n19524), .dout(n19526));
  jand g19271(.dina(n19526), .dinb(n19101), .dout(n19527));
  jand g19272(.dina(asqrt[8] ), .dinb(a[16] ), .dout(n19528));
  jor  g19273(.dina(n19528), .dinb(n19527), .dout(n19529));
  jand g19274(.dina(n19529), .dinb(asqrt[9] ), .dout(n19530));
  jor  g19275(.dina(n19529), .dinb(asqrt[9] ), .dout(n19531));
  jand g19276(.dina(asqrt[8] ), .dinb(n19101), .dout(n19532));
  jor  g19277(.dina(n19532), .dinb(n19102), .dout(n19533));
  jnot g19278(.din(n19103), .dout(n19534));
  jnot g19279(.din(n19498), .dout(n19535));
  jnot g19280(.din(n19491), .dout(n19536));
  jnot g19281(.din(n19484), .dout(n19537));
  jnot g19282(.din(n19476), .dout(n19538));
  jnot g19283(.din(n19468), .dout(n19539));
  jnot g19284(.din(n19461), .dout(n19540));
  jnot g19285(.din(n19453), .dout(n19541));
  jnot g19286(.din(n19446), .dout(n19542));
  jnot g19287(.din(n19438), .dout(n19543));
  jnot g19288(.din(n19430), .dout(n19544));
  jnot g19289(.din(n19423), .dout(n19545));
  jnot g19290(.din(n19416), .dout(n19546));
  jnot g19291(.din(n19408), .dout(n19547));
  jnot g19292(.din(n19401), .dout(n19548));
  jnot g19293(.din(n19393), .dout(n19549));
  jnot g19294(.din(n19386), .dout(n19550));
  jnot g19295(.din(n19379), .dout(n19551));
  jnot g19296(.din(n19372), .dout(n19552));
  jnot g19297(.din(n19365), .dout(n19553));
  jnot g19298(.din(n19358), .dout(n19554));
  jnot g19299(.din(n19350), .dout(n19555));
  jnot g19300(.din(n19343), .dout(n19556));
  jnot g19301(.din(n19336), .dout(n19557));
  jnot g19302(.din(n19329), .dout(n19558));
  jnot g19303(.din(n19321), .dout(n19559));
  jnot g19304(.din(n19314), .dout(n19560));
  jnot g19305(.din(n19306), .dout(n19561));
  jnot g19306(.din(n19299), .dout(n19562));
  jnot g19307(.din(n19291), .dout(n19563));
  jnot g19308(.din(n19284), .dout(n19564));
  jnot g19309(.din(n19276), .dout(n19565));
  jnot g19310(.din(n19269), .dout(n19566));
  jnot g19311(.din(n19262), .dout(n19567));
  jnot g19312(.din(n19255), .dout(n19568));
  jnot g19313(.din(n19247), .dout(n19569));
  jnot g19314(.din(n19240), .dout(n19570));
  jnot g19315(.din(n19232), .dout(n19571));
  jnot g19316(.din(n19225), .dout(n19572));
  jnot g19317(.din(n19217), .dout(n19573));
  jnot g19318(.din(n19209), .dout(n19574));
  jnot g19319(.din(n19202), .dout(n19575));
  jnot g19320(.din(n19195), .dout(n19576));
  jnot g19321(.din(n19187), .dout(n19577));
  jnot g19322(.din(n19180), .dout(n19578));
  jnot g19323(.din(n19172), .dout(n19579));
  jnot g19324(.din(n19165), .dout(n19580));
  jnot g19325(.din(n19157), .dout(n19581));
  jnot g19326(.din(n19150), .dout(n19582));
  jnot g19327(.din(n19142), .dout(n19583));
  jnot g19328(.din(n19135), .dout(n19584));
  jnot g19329(.din(n19127), .dout(n19585));
  jnot g19330(.din(n19116), .dout(n19586));
  jnot g19331(.din(n19108), .dout(n19587));
  jand g19332(.dina(asqrt[9] ), .dinb(a[18] ), .dout(n19588));
  jor  g19333(.dina(n19588), .dinb(n19104), .dout(n19589));
  jor  g19334(.dina(n19589), .dinb(asqrt[10] ), .dout(n19590));
  jand g19335(.dina(asqrt[9] ), .dinb(n18185), .dout(n19591));
  jor  g19336(.dina(n19591), .dinb(n18186), .dout(n19592));
  jand g19337(.dina(n19119), .dinb(n19592), .dout(n19593));
  jand g19338(.dina(n19593), .dinb(n19590), .dout(n19594));
  jor  g19339(.dina(n19594), .dinb(n19587), .dout(n19595));
  jor  g19340(.dina(n19595), .dinb(asqrt[11] ), .dout(n19596));
  jnot g19341(.din(n19124), .dout(n19597));
  jand g19342(.dina(n19597), .dinb(n19596), .dout(n19598));
  jor  g19343(.dina(n19598), .dinb(n19586), .dout(n19599));
  jor  g19344(.dina(n19599), .dinb(asqrt[12] ), .dout(n19600));
  jand g19345(.dina(n19131), .dinb(n19600), .dout(n19601));
  jor  g19346(.dina(n19601), .dinb(n19585), .dout(n19602));
  jor  g19347(.dina(n19602), .dinb(asqrt[13] ), .dout(n19603));
  jnot g19348(.din(n19139), .dout(n19604));
  jand g19349(.dina(n19604), .dinb(n19603), .dout(n19605));
  jor  g19350(.dina(n19605), .dinb(n19584), .dout(n19606));
  jor  g19351(.dina(n19606), .dinb(asqrt[14] ), .dout(n19607));
  jand g19352(.dina(n19146), .dinb(n19607), .dout(n19608));
  jor  g19353(.dina(n19608), .dinb(n19583), .dout(n19609));
  jor  g19354(.dina(n19609), .dinb(asqrt[15] ), .dout(n19610));
  jnot g19355(.din(n19154), .dout(n19611));
  jand g19356(.dina(n19611), .dinb(n19610), .dout(n19612));
  jor  g19357(.dina(n19612), .dinb(n19582), .dout(n19613));
  jor  g19358(.dina(n19613), .dinb(asqrt[16] ), .dout(n19614));
  jand g19359(.dina(n19161), .dinb(n19614), .dout(n19615));
  jor  g19360(.dina(n19615), .dinb(n19581), .dout(n19616));
  jor  g19361(.dina(n19616), .dinb(asqrt[17] ), .dout(n19617));
  jnot g19362(.din(n19169), .dout(n19618));
  jand g19363(.dina(n19618), .dinb(n19617), .dout(n19619));
  jor  g19364(.dina(n19619), .dinb(n19580), .dout(n19620));
  jor  g19365(.dina(n19620), .dinb(asqrt[18] ), .dout(n19621));
  jand g19366(.dina(n19176), .dinb(n19621), .dout(n19622));
  jor  g19367(.dina(n19622), .dinb(n19579), .dout(n19623));
  jor  g19368(.dina(n19623), .dinb(asqrt[19] ), .dout(n19624));
  jnot g19369(.din(n19184), .dout(n19625));
  jand g19370(.dina(n19625), .dinb(n19624), .dout(n19626));
  jor  g19371(.dina(n19626), .dinb(n19578), .dout(n19627));
  jor  g19372(.dina(n19627), .dinb(asqrt[20] ), .dout(n19628));
  jand g19373(.dina(n19191), .dinb(n19628), .dout(n19629));
  jor  g19374(.dina(n19629), .dinb(n19577), .dout(n19630));
  jor  g19375(.dina(n19630), .dinb(asqrt[21] ), .dout(n19631));
  jnot g19376(.din(n19199), .dout(n19632));
  jand g19377(.dina(n19632), .dinb(n19631), .dout(n19633));
  jor  g19378(.dina(n19633), .dinb(n19576), .dout(n19634));
  jor  g19379(.dina(n19634), .dinb(asqrt[22] ), .dout(n19635));
  jnot g19380(.din(n19206), .dout(n19636));
  jand g19381(.dina(n19636), .dinb(n19635), .dout(n19637));
  jor  g19382(.dina(n19637), .dinb(n19575), .dout(n19638));
  jor  g19383(.dina(n19638), .dinb(asqrt[23] ), .dout(n19639));
  jand g19384(.dina(n19213), .dinb(n19639), .dout(n19640));
  jor  g19385(.dina(n19640), .dinb(n19574), .dout(n19641));
  jor  g19386(.dina(n19641), .dinb(asqrt[24] ), .dout(n19642));
  jand g19387(.dina(n19221), .dinb(n19642), .dout(n19643));
  jor  g19388(.dina(n19643), .dinb(n19573), .dout(n19644));
  jor  g19389(.dina(n19644), .dinb(asqrt[25] ), .dout(n19645));
  jnot g19390(.din(n19229), .dout(n19646));
  jand g19391(.dina(n19646), .dinb(n19645), .dout(n19647));
  jor  g19392(.dina(n19647), .dinb(n19572), .dout(n19648));
  jor  g19393(.dina(n19648), .dinb(asqrt[26] ), .dout(n19649));
  jand g19394(.dina(n19236), .dinb(n19649), .dout(n19650));
  jor  g19395(.dina(n19650), .dinb(n19571), .dout(n19651));
  jor  g19396(.dina(n19651), .dinb(asqrt[27] ), .dout(n19652));
  jnot g19397(.din(n19244), .dout(n19653));
  jand g19398(.dina(n19653), .dinb(n19652), .dout(n19654));
  jor  g19399(.dina(n19654), .dinb(n19570), .dout(n19655));
  jor  g19400(.dina(n19655), .dinb(asqrt[28] ), .dout(n19656));
  jand g19401(.dina(n19251), .dinb(n19656), .dout(n19657));
  jor  g19402(.dina(n19657), .dinb(n19569), .dout(n19658));
  jor  g19403(.dina(n19658), .dinb(asqrt[29] ), .dout(n19659));
  jnot g19404(.din(n19259), .dout(n19660));
  jand g19405(.dina(n19660), .dinb(n19659), .dout(n19661));
  jor  g19406(.dina(n19661), .dinb(n19568), .dout(n19662));
  jor  g19407(.dina(n19662), .dinb(asqrt[30] ), .dout(n19663));
  jnot g19408(.din(n19266), .dout(n19664));
  jand g19409(.dina(n19664), .dinb(n19663), .dout(n19665));
  jor  g19410(.dina(n19665), .dinb(n19567), .dout(n19666));
  jor  g19411(.dina(n19666), .dinb(asqrt[31] ), .dout(n19667));
  jnot g19412(.din(n19273), .dout(n19668));
  jand g19413(.dina(n19668), .dinb(n19667), .dout(n19669));
  jor  g19414(.dina(n19669), .dinb(n19566), .dout(n19670));
  jor  g19415(.dina(n19670), .dinb(asqrt[32] ), .dout(n19671));
  jand g19416(.dina(n19280), .dinb(n19671), .dout(n19672));
  jor  g19417(.dina(n19672), .dinb(n19565), .dout(n19673));
  jor  g19418(.dina(n19673), .dinb(asqrt[33] ), .dout(n19674));
  jnot g19419(.din(n19288), .dout(n19675));
  jand g19420(.dina(n19675), .dinb(n19674), .dout(n19676));
  jor  g19421(.dina(n19676), .dinb(n19564), .dout(n19677));
  jor  g19422(.dina(n19677), .dinb(asqrt[34] ), .dout(n19678));
  jand g19423(.dina(n19295), .dinb(n19678), .dout(n19679));
  jor  g19424(.dina(n19679), .dinb(n19563), .dout(n19680));
  jor  g19425(.dina(n19680), .dinb(asqrt[35] ), .dout(n19681));
  jnot g19426(.din(n19303), .dout(n19682));
  jand g19427(.dina(n19682), .dinb(n19681), .dout(n19683));
  jor  g19428(.dina(n19683), .dinb(n19562), .dout(n19684));
  jor  g19429(.dina(n19684), .dinb(asqrt[36] ), .dout(n19685));
  jand g19430(.dina(n19310), .dinb(n19685), .dout(n19686));
  jor  g19431(.dina(n19686), .dinb(n19561), .dout(n19687));
  jor  g19432(.dina(n19687), .dinb(asqrt[37] ), .dout(n19688));
  jnot g19433(.din(n19318), .dout(n19689));
  jand g19434(.dina(n19689), .dinb(n19688), .dout(n19690));
  jor  g19435(.dina(n19690), .dinb(n19560), .dout(n19691));
  jor  g19436(.dina(n19691), .dinb(asqrt[38] ), .dout(n19692));
  jand g19437(.dina(n19325), .dinb(n19692), .dout(n19693));
  jor  g19438(.dina(n19693), .dinb(n19559), .dout(n19694));
  jor  g19439(.dina(n19694), .dinb(asqrt[39] ), .dout(n19695));
  jnot g19440(.din(n19333), .dout(n19696));
  jand g19441(.dina(n19696), .dinb(n19695), .dout(n19697));
  jor  g19442(.dina(n19697), .dinb(n19558), .dout(n19698));
  jor  g19443(.dina(n19698), .dinb(asqrt[40] ), .dout(n19699));
  jnot g19444(.din(n19340), .dout(n19700));
  jand g19445(.dina(n19700), .dinb(n19699), .dout(n19701));
  jor  g19446(.dina(n19701), .dinb(n19557), .dout(n19702));
  jor  g19447(.dina(n19702), .dinb(asqrt[41] ), .dout(n19703));
  jnot g19448(.din(n19347), .dout(n19704));
  jand g19449(.dina(n19704), .dinb(n19703), .dout(n19705));
  jor  g19450(.dina(n19705), .dinb(n19556), .dout(n19706));
  jor  g19451(.dina(n19706), .dinb(asqrt[42] ), .dout(n19707));
  jand g19452(.dina(n19354), .dinb(n19707), .dout(n19708));
  jor  g19453(.dina(n19708), .dinb(n19555), .dout(n19709));
  jor  g19454(.dina(n19709), .dinb(asqrt[43] ), .dout(n19710));
  jnot g19455(.din(n19362), .dout(n19711));
  jand g19456(.dina(n19711), .dinb(n19710), .dout(n19712));
  jor  g19457(.dina(n19712), .dinb(n19554), .dout(n19713));
  jor  g19458(.dina(n19713), .dinb(asqrt[44] ), .dout(n19714));
  jnot g19459(.din(n19369), .dout(n19715));
  jand g19460(.dina(n19715), .dinb(n19714), .dout(n19716));
  jor  g19461(.dina(n19716), .dinb(n19553), .dout(n19717));
  jor  g19462(.dina(n19717), .dinb(asqrt[45] ), .dout(n19718));
  jnot g19463(.din(n19376), .dout(n19719));
  jand g19464(.dina(n19719), .dinb(n19718), .dout(n19720));
  jor  g19465(.dina(n19720), .dinb(n19552), .dout(n19721));
  jor  g19466(.dina(n19721), .dinb(asqrt[46] ), .dout(n19722));
  jnot g19467(.din(n19383), .dout(n19723));
  jand g19468(.dina(n19723), .dinb(n19722), .dout(n19724));
  jor  g19469(.dina(n19724), .dinb(n19551), .dout(n19725));
  jor  g19470(.dina(n19725), .dinb(asqrt[47] ), .dout(n19726));
  jnot g19471(.din(n19390), .dout(n19727));
  jand g19472(.dina(n19727), .dinb(n19726), .dout(n19728));
  jor  g19473(.dina(n19728), .dinb(n19550), .dout(n19729));
  jor  g19474(.dina(n19729), .dinb(asqrt[48] ), .dout(n19730));
  jand g19475(.dina(n19397), .dinb(n19730), .dout(n19731));
  jor  g19476(.dina(n19731), .dinb(n19549), .dout(n19732));
  jor  g19477(.dina(n19732), .dinb(asqrt[49] ), .dout(n19733));
  jnot g19478(.din(n19405), .dout(n19734));
  jand g19479(.dina(n19734), .dinb(n19733), .dout(n19735));
  jor  g19480(.dina(n19735), .dinb(n19548), .dout(n19736));
  jor  g19481(.dina(n19736), .dinb(asqrt[50] ), .dout(n19737));
  jand g19482(.dina(n19412), .dinb(n19737), .dout(n19738));
  jor  g19483(.dina(n19738), .dinb(n19547), .dout(n19739));
  jor  g19484(.dina(n19739), .dinb(asqrt[51] ), .dout(n19740));
  jnot g19485(.din(n19420), .dout(n19741));
  jand g19486(.dina(n19741), .dinb(n19740), .dout(n19742));
  jor  g19487(.dina(n19742), .dinb(n19546), .dout(n19743));
  jor  g19488(.dina(n19743), .dinb(asqrt[52] ), .dout(n19744));
  jnot g19489(.din(n19427), .dout(n19745));
  jand g19490(.dina(n19745), .dinb(n19744), .dout(n19746));
  jor  g19491(.dina(n19746), .dinb(n19545), .dout(n19747));
  jor  g19492(.dina(n19747), .dinb(asqrt[53] ), .dout(n19748));
  jand g19493(.dina(n19434), .dinb(n19748), .dout(n19749));
  jor  g19494(.dina(n19749), .dinb(n19544), .dout(n19750));
  jor  g19495(.dina(n19750), .dinb(asqrt[54] ), .dout(n19751));
  jand g19496(.dina(n19751), .dinb(n19441), .dout(n19752));
  jor  g19497(.dina(n19752), .dinb(n19543), .dout(n19753));
  jor  g19498(.dina(n19753), .dinb(asqrt[55] ), .dout(n19754));
  jnot g19499(.din(n19450), .dout(n19755));
  jand g19500(.dina(n19755), .dinb(n19754), .dout(n19756));
  jor  g19501(.dina(n19756), .dinb(n19542), .dout(n19757));
  jor  g19502(.dina(n19757), .dinb(asqrt[56] ), .dout(n19758));
  jand g19503(.dina(n19457), .dinb(n19758), .dout(n19759));
  jor  g19504(.dina(n19759), .dinb(n19541), .dout(n19760));
  jor  g19505(.dina(n19760), .dinb(asqrt[57] ), .dout(n19761));
  jnot g19506(.din(n19465), .dout(n19762));
  jand g19507(.dina(n19762), .dinb(n19761), .dout(n19763));
  jor  g19508(.dina(n19763), .dinb(n19540), .dout(n19764));
  jor  g19509(.dina(n19764), .dinb(asqrt[58] ), .dout(n19765));
  jand g19510(.dina(n19472), .dinb(n19765), .dout(n19766));
  jor  g19511(.dina(n19766), .dinb(n19539), .dout(n19767));
  jor  g19512(.dina(n19767), .dinb(asqrt[59] ), .dout(n19768));
  jand g19513(.dina(n19480), .dinb(n19768), .dout(n19769));
  jor  g19514(.dina(n19769), .dinb(n19538), .dout(n19770));
  jor  g19515(.dina(n19770), .dinb(asqrt[60] ), .dout(n19771));
  jnot g19516(.din(n19488), .dout(n19772));
  jand g19517(.dina(n19772), .dinb(n19771), .dout(n19773));
  jor  g19518(.dina(n19773), .dinb(n19537), .dout(n19774));
  jor  g19519(.dina(n19774), .dinb(asqrt[61] ), .dout(n19775));
  jnot g19520(.din(n19495), .dout(n19776));
  jand g19521(.dina(n19776), .dinb(n19775), .dout(n19777));
  jor  g19522(.dina(n19777), .dinb(n19536), .dout(n19778));
  jor  g19523(.dina(n19778), .dinb(asqrt[62] ), .dout(n19779));
  jand g19524(.dina(n19502), .dinb(n19779), .dout(n19780));
  jor  g19525(.dina(n19780), .dinb(n19535), .dout(n19781));
  jand g19526(.dina(n19781), .dinb(n19099), .dout(n19782));
  jnot g19527(.din(n19508), .dout(n19783));
  jand g19528(.dina(n19783), .dinb(n19782), .dout(n19784));
  jor  g19529(.dina(n19784), .dinb(asqrt[63] ), .dout(n19785));
  jor  g19530(.dina(n19781), .dinb(n19099), .dout(n19786));
  jnot g19531(.din(n19515), .dout(n19787));
  jand g19532(.dina(n19787), .dinb(n19786), .dout(n19788));
  jand g19533(.dina(n19788), .dinb(n19785), .dout(n19791));
  jor  g19534(.dina(n19791), .dinb(n19534), .dout(n19792));
  jand g19535(.dina(n19792), .dinb(n19533), .dout(n19793));
  jand g19536(.dina(n19793), .dinb(n19531), .dout(n19794));
  jor  g19537(.dina(n19794), .dinb(n19530), .dout(n19795));
  jand g19538(.dina(n19795), .dinb(asqrt[10] ), .dout(n19796));
  jor  g19539(.dina(n19795), .dinb(asqrt[10] ), .dout(n19797));
  jand g19540(.dina(asqrt[8] ), .dinb(n19103), .dout(n19798));
  jand g19541(.dina(n19788), .dinb(asqrt[9] ), .dout(n19799));
  jand g19542(.dina(n19799), .dinb(n19785), .dout(n19800));
  jor  g19543(.dina(n19800), .dinb(n19798), .dout(n19801));
  jxor g19544(.dina(n19801), .dinb(a[18] ), .dout(n19802));
  jnot g19545(.din(n19802), .dout(n19803));
  jand g19546(.dina(n19803), .dinb(n19797), .dout(n19804));
  jor  g19547(.dina(n19804), .dinb(n19796), .dout(n19805));
  jand g19548(.dina(n19805), .dinb(asqrt[11] ), .dout(n19806));
  jor  g19549(.dina(n19805), .dinb(asqrt[11] ), .dout(n19807));
  jxor g19550(.dina(n19107), .dinb(n18442), .dout(n19808));
  jand g19551(.dina(n19808), .dinb(asqrt[8] ), .dout(n19809));
  jxor g19552(.dina(n19809), .dinb(n19113), .dout(n19810));
  jnot g19553(.din(n19810), .dout(n19811));
  jand g19554(.dina(n19811), .dinb(n19807), .dout(n19812));
  jor  g19555(.dina(n19812), .dinb(n19806), .dout(n19813));
  jand g19556(.dina(n19813), .dinb(asqrt[12] ), .dout(n19814));
  jor  g19557(.dina(n19813), .dinb(asqrt[12] ), .dout(n19815));
  jxor g19558(.dina(n19115), .dinb(n17769), .dout(n19816));
  jand g19559(.dina(n19816), .dinb(asqrt[8] ), .dout(n19817));
  jxor g19560(.dina(n19817), .dinb(n19124), .dout(n19818));
  jnot g19561(.din(n19818), .dout(n19819));
  jand g19562(.dina(n19819), .dinb(n19815), .dout(n19820));
  jor  g19563(.dina(n19820), .dinb(n19814), .dout(n19821));
  jand g19564(.dina(n19821), .dinb(asqrt[13] ), .dout(n19822));
  jor  g19565(.dina(n19821), .dinb(asqrt[13] ), .dout(n19823));
  jxor g19566(.dina(n19126), .dinb(n17134), .dout(n19824));
  jand g19567(.dina(n19824), .dinb(asqrt[8] ), .dout(n19825));
  jxor g19568(.dina(n19825), .dinb(n19131), .dout(n19826));
  jand g19569(.dina(n19826), .dinb(n19823), .dout(n19827));
  jor  g19570(.dina(n19827), .dinb(n19822), .dout(n19828));
  jand g19571(.dina(n19828), .dinb(asqrt[14] ), .dout(n19829));
  jor  g19572(.dina(n19828), .dinb(asqrt[14] ), .dout(n19830));
  jxor g19573(.dina(n19134), .dinb(n16489), .dout(n19831));
  jand g19574(.dina(n19831), .dinb(asqrt[8] ), .dout(n19832));
  jxor g19575(.dina(n19832), .dinb(n19139), .dout(n19833));
  jnot g19576(.din(n19833), .dout(n19834));
  jand g19577(.dina(n19834), .dinb(n19830), .dout(n19835));
  jor  g19578(.dina(n19835), .dinb(n19829), .dout(n19836));
  jand g19579(.dina(n19836), .dinb(asqrt[15] ), .dout(n19837));
  jor  g19580(.dina(n19836), .dinb(asqrt[15] ), .dout(n19838));
  jxor g19581(.dina(n19141), .dinb(n15878), .dout(n19839));
  jand g19582(.dina(n19839), .dinb(asqrt[8] ), .dout(n19840));
  jxor g19583(.dina(n19840), .dinb(n19146), .dout(n19841));
  jand g19584(.dina(n19841), .dinb(n19838), .dout(n19842));
  jor  g19585(.dina(n19842), .dinb(n19837), .dout(n19843));
  jand g19586(.dina(n19843), .dinb(asqrt[16] ), .dout(n19844));
  jor  g19587(.dina(n19843), .dinb(asqrt[16] ), .dout(n19845));
  jxor g19588(.dina(n19149), .dinb(n15260), .dout(n19846));
  jand g19589(.dina(n19846), .dinb(asqrt[8] ), .dout(n19847));
  jxor g19590(.dina(n19847), .dinb(n19154), .dout(n19848));
  jnot g19591(.din(n19848), .dout(n19849));
  jand g19592(.dina(n19849), .dinb(n19845), .dout(n19850));
  jor  g19593(.dina(n19850), .dinb(n19844), .dout(n19851));
  jand g19594(.dina(n19851), .dinb(asqrt[17] ), .dout(n19852));
  jor  g19595(.dina(n19851), .dinb(asqrt[17] ), .dout(n19853));
  jxor g19596(.dina(n19156), .dinb(n14674), .dout(n19854));
  jand g19597(.dina(n19854), .dinb(asqrt[8] ), .dout(n19855));
  jxor g19598(.dina(n19855), .dinb(n19161), .dout(n19856));
  jand g19599(.dina(n19856), .dinb(n19853), .dout(n19857));
  jor  g19600(.dina(n19857), .dinb(n19852), .dout(n19858));
  jand g19601(.dina(n19858), .dinb(asqrt[18] ), .dout(n19859));
  jor  g19602(.dina(n19858), .dinb(asqrt[18] ), .dout(n19860));
  jxor g19603(.dina(n19164), .dinb(n14078), .dout(n19861));
  jand g19604(.dina(n19861), .dinb(asqrt[8] ), .dout(n19862));
  jxor g19605(.dina(n19862), .dinb(n19169), .dout(n19863));
  jnot g19606(.din(n19863), .dout(n19864));
  jand g19607(.dina(n19864), .dinb(n19860), .dout(n19865));
  jor  g19608(.dina(n19865), .dinb(n19859), .dout(n19866));
  jand g19609(.dina(n19866), .dinb(asqrt[19] ), .dout(n19867));
  jor  g19610(.dina(n19866), .dinb(asqrt[19] ), .dout(n19868));
  jxor g19611(.dina(n19171), .dinb(n13515), .dout(n19869));
  jand g19612(.dina(n19869), .dinb(asqrt[8] ), .dout(n19870));
  jxor g19613(.dina(n19870), .dinb(n19176), .dout(n19871));
  jand g19614(.dina(n19871), .dinb(n19868), .dout(n19872));
  jor  g19615(.dina(n19872), .dinb(n19867), .dout(n19873));
  jand g19616(.dina(n19873), .dinb(asqrt[20] ), .dout(n19874));
  jor  g19617(.dina(n19873), .dinb(asqrt[20] ), .dout(n19875));
  jxor g19618(.dina(n19179), .dinb(n12947), .dout(n19876));
  jand g19619(.dina(n19876), .dinb(asqrt[8] ), .dout(n19877));
  jxor g19620(.dina(n19877), .dinb(n19184), .dout(n19878));
  jnot g19621(.din(n19878), .dout(n19879));
  jand g19622(.dina(n19879), .dinb(n19875), .dout(n19880));
  jor  g19623(.dina(n19880), .dinb(n19874), .dout(n19881));
  jand g19624(.dina(n19881), .dinb(asqrt[21] ), .dout(n19882));
  jor  g19625(.dina(n19881), .dinb(asqrt[21] ), .dout(n19883));
  jxor g19626(.dina(n19186), .dinb(n12410), .dout(n19884));
  jand g19627(.dina(n19884), .dinb(asqrt[8] ), .dout(n19885));
  jxor g19628(.dina(n19885), .dinb(n19191), .dout(n19886));
  jand g19629(.dina(n19886), .dinb(n19883), .dout(n19887));
  jor  g19630(.dina(n19887), .dinb(n19882), .dout(n19888));
  jand g19631(.dina(n19888), .dinb(asqrt[22] ), .dout(n19889));
  jor  g19632(.dina(n19888), .dinb(asqrt[22] ), .dout(n19890));
  jxor g19633(.dina(n19194), .dinb(n11858), .dout(n19891));
  jand g19634(.dina(n19891), .dinb(asqrt[8] ), .dout(n19892));
  jxor g19635(.dina(n19892), .dinb(n19199), .dout(n19893));
  jnot g19636(.din(n19893), .dout(n19894));
  jand g19637(.dina(n19894), .dinb(n19890), .dout(n19895));
  jor  g19638(.dina(n19895), .dinb(n19889), .dout(n19896));
  jand g19639(.dina(n19896), .dinb(asqrt[23] ), .dout(n19897));
  jor  g19640(.dina(n19896), .dinb(asqrt[23] ), .dout(n19898));
  jxor g19641(.dina(n19201), .dinb(n11347), .dout(n19899));
  jand g19642(.dina(n19899), .dinb(asqrt[8] ), .dout(n19900));
  jxor g19643(.dina(n19900), .dinb(n19206), .dout(n19901));
  jnot g19644(.din(n19901), .dout(n19902));
  jand g19645(.dina(n19902), .dinb(n19898), .dout(n19903));
  jor  g19646(.dina(n19903), .dinb(n19897), .dout(n19904));
  jand g19647(.dina(n19904), .dinb(asqrt[24] ), .dout(n19905));
  jor  g19648(.dina(n19904), .dinb(asqrt[24] ), .dout(n19906));
  jxor g19649(.dina(n19208), .dinb(n10824), .dout(n19907));
  jand g19650(.dina(n19907), .dinb(asqrt[8] ), .dout(n19908));
  jxor g19651(.dina(n19908), .dinb(n19213), .dout(n19909));
  jand g19652(.dina(n19909), .dinb(n19906), .dout(n19910));
  jor  g19653(.dina(n19910), .dinb(n19905), .dout(n19911));
  jand g19654(.dina(n19911), .dinb(asqrt[25] ), .dout(n19912));
  jor  g19655(.dina(n19911), .dinb(asqrt[25] ), .dout(n19913));
  jxor g19656(.dina(n19216), .dinb(n10328), .dout(n19914));
  jand g19657(.dina(n19914), .dinb(asqrt[8] ), .dout(n19915));
  jxor g19658(.dina(n19915), .dinb(n19221), .dout(n19916));
  jand g19659(.dina(n19916), .dinb(n19913), .dout(n19917));
  jor  g19660(.dina(n19917), .dinb(n19912), .dout(n19918));
  jand g19661(.dina(n19918), .dinb(asqrt[26] ), .dout(n19919));
  jor  g19662(.dina(n19918), .dinb(asqrt[26] ), .dout(n19920));
  jxor g19663(.dina(n19224), .dinb(n9832), .dout(n19921));
  jand g19664(.dina(n19921), .dinb(asqrt[8] ), .dout(n19922));
  jxor g19665(.dina(n19922), .dinb(n19229), .dout(n19923));
  jnot g19666(.din(n19923), .dout(n19924));
  jand g19667(.dina(n19924), .dinb(n19920), .dout(n19925));
  jor  g19668(.dina(n19925), .dinb(n19919), .dout(n19926));
  jand g19669(.dina(n19926), .dinb(asqrt[27] ), .dout(n19927));
  jor  g19670(.dina(n19926), .dinb(asqrt[27] ), .dout(n19928));
  jxor g19671(.dina(n19231), .dinb(n9369), .dout(n19929));
  jand g19672(.dina(n19929), .dinb(asqrt[8] ), .dout(n19930));
  jxor g19673(.dina(n19930), .dinb(n19236), .dout(n19931));
  jand g19674(.dina(n19931), .dinb(n19928), .dout(n19932));
  jor  g19675(.dina(n19932), .dinb(n19927), .dout(n19933));
  jand g19676(.dina(n19933), .dinb(asqrt[28] ), .dout(n19934));
  jor  g19677(.dina(n19933), .dinb(asqrt[28] ), .dout(n19935));
  jxor g19678(.dina(n19239), .dinb(n8890), .dout(n19936));
  jand g19679(.dina(n19936), .dinb(asqrt[8] ), .dout(n19937));
  jxor g19680(.dina(n19937), .dinb(n19244), .dout(n19938));
  jnot g19681(.din(n19938), .dout(n19939));
  jand g19682(.dina(n19939), .dinb(n19935), .dout(n19940));
  jor  g19683(.dina(n19940), .dinb(n19934), .dout(n19941));
  jand g19684(.dina(n19941), .dinb(asqrt[29] ), .dout(n19942));
  jor  g19685(.dina(n19941), .dinb(asqrt[29] ), .dout(n19943));
  jxor g19686(.dina(n19246), .dinb(n8449), .dout(n19944));
  jand g19687(.dina(n19944), .dinb(asqrt[8] ), .dout(n19945));
  jxor g19688(.dina(n19945), .dinb(n19251), .dout(n19946));
  jand g19689(.dina(n19946), .dinb(n19943), .dout(n19947));
  jor  g19690(.dina(n19947), .dinb(n19942), .dout(n19948));
  jand g19691(.dina(n19948), .dinb(asqrt[30] ), .dout(n19949));
  jor  g19692(.dina(n19948), .dinb(asqrt[30] ), .dout(n19950));
  jxor g19693(.dina(n19254), .dinb(n8003), .dout(n19951));
  jand g19694(.dina(n19951), .dinb(asqrt[8] ), .dout(n19952));
  jxor g19695(.dina(n19952), .dinb(n19259), .dout(n19953));
  jnot g19696(.din(n19953), .dout(n19954));
  jand g19697(.dina(n19954), .dinb(n19950), .dout(n19955));
  jor  g19698(.dina(n19955), .dinb(n19949), .dout(n19956));
  jand g19699(.dina(n19956), .dinb(asqrt[31] ), .dout(n19957));
  jor  g19700(.dina(n19956), .dinb(asqrt[31] ), .dout(n19958));
  jxor g19701(.dina(n19261), .dinb(n7581), .dout(n19959));
  jand g19702(.dina(n19959), .dinb(asqrt[8] ), .dout(n19960));
  jxor g19703(.dina(n19960), .dinb(n19266), .dout(n19961));
  jnot g19704(.din(n19961), .dout(n19962));
  jand g19705(.dina(n19962), .dinb(n19958), .dout(n19963));
  jor  g19706(.dina(n19963), .dinb(n19957), .dout(n19964));
  jand g19707(.dina(n19964), .dinb(asqrt[32] ), .dout(n19965));
  jor  g19708(.dina(n19964), .dinb(asqrt[32] ), .dout(n19966));
  jxor g19709(.dina(n19268), .dinb(n7154), .dout(n19967));
  jand g19710(.dina(n19967), .dinb(asqrt[8] ), .dout(n19968));
  jxor g19711(.dina(n19968), .dinb(n19273), .dout(n19969));
  jnot g19712(.din(n19969), .dout(n19970));
  jand g19713(.dina(n19970), .dinb(n19966), .dout(n19971));
  jor  g19714(.dina(n19971), .dinb(n19965), .dout(n19972));
  jand g19715(.dina(n19972), .dinb(asqrt[33] ), .dout(n19973));
  jor  g19716(.dina(n19972), .dinb(asqrt[33] ), .dout(n19974));
  jxor g19717(.dina(n19275), .dinb(n6758), .dout(n19975));
  jand g19718(.dina(n19975), .dinb(asqrt[8] ), .dout(n19976));
  jxor g19719(.dina(n19976), .dinb(n19280), .dout(n19977));
  jand g19720(.dina(n19977), .dinb(n19974), .dout(n19978));
  jor  g19721(.dina(n19978), .dinb(n19973), .dout(n19979));
  jand g19722(.dina(n19979), .dinb(asqrt[34] ), .dout(n19980));
  jor  g19723(.dina(n19979), .dinb(asqrt[34] ), .dout(n19981));
  jxor g19724(.dina(n19283), .dinb(n6357), .dout(n19982));
  jand g19725(.dina(n19982), .dinb(asqrt[8] ), .dout(n19983));
  jxor g19726(.dina(n19983), .dinb(n19288), .dout(n19984));
  jnot g19727(.din(n19984), .dout(n19985));
  jand g19728(.dina(n19985), .dinb(n19981), .dout(n19986));
  jor  g19729(.dina(n19986), .dinb(n19980), .dout(n19987));
  jand g19730(.dina(n19987), .dinb(asqrt[35] ), .dout(n19988));
  jor  g19731(.dina(n19987), .dinb(asqrt[35] ), .dout(n19989));
  jxor g19732(.dina(n19290), .dinb(n5989), .dout(n19990));
  jand g19733(.dina(n19990), .dinb(asqrt[8] ), .dout(n19991));
  jxor g19734(.dina(n19991), .dinb(n19295), .dout(n19992));
  jand g19735(.dina(n19992), .dinb(n19989), .dout(n19993));
  jor  g19736(.dina(n19993), .dinb(n19988), .dout(n19994));
  jand g19737(.dina(n19994), .dinb(asqrt[36] ), .dout(n19995));
  jor  g19738(.dina(n19994), .dinb(asqrt[36] ), .dout(n19996));
  jxor g19739(.dina(n19298), .dinb(n5606), .dout(n19997));
  jand g19740(.dina(n19997), .dinb(asqrt[8] ), .dout(n19998));
  jxor g19741(.dina(n19998), .dinb(n19303), .dout(n19999));
  jnot g19742(.din(n19999), .dout(n20000));
  jand g19743(.dina(n20000), .dinb(n19996), .dout(n20001));
  jor  g19744(.dina(n20001), .dinb(n19995), .dout(n20002));
  jand g19745(.dina(n20002), .dinb(asqrt[37] ), .dout(n20003));
  jor  g19746(.dina(n20002), .dinb(asqrt[37] ), .dout(n20004));
  jxor g19747(.dina(n19305), .dinb(n5259), .dout(n20005));
  jand g19748(.dina(n20005), .dinb(asqrt[8] ), .dout(n20006));
  jxor g19749(.dina(n20006), .dinb(n19310), .dout(n20007));
  jand g19750(.dina(n20007), .dinb(n20004), .dout(n20008));
  jor  g19751(.dina(n20008), .dinb(n20003), .dout(n20009));
  jand g19752(.dina(n20009), .dinb(asqrt[38] ), .dout(n20010));
  jor  g19753(.dina(n20009), .dinb(asqrt[38] ), .dout(n20011));
  jxor g19754(.dina(n19313), .dinb(n4902), .dout(n20012));
  jand g19755(.dina(n20012), .dinb(asqrt[8] ), .dout(n20013));
  jxor g19756(.dina(n20013), .dinb(n19318), .dout(n20014));
  jnot g19757(.din(n20014), .dout(n20015));
  jand g19758(.dina(n20015), .dinb(n20011), .dout(n20016));
  jor  g19759(.dina(n20016), .dinb(n20010), .dout(n20017));
  jand g19760(.dina(n20017), .dinb(asqrt[39] ), .dout(n20018));
  jor  g19761(.dina(n20017), .dinb(asqrt[39] ), .dout(n20019));
  jxor g19762(.dina(n19320), .dinb(n4582), .dout(n20020));
  jand g19763(.dina(n20020), .dinb(asqrt[8] ), .dout(n20021));
  jxor g19764(.dina(n20021), .dinb(n19325), .dout(n20022));
  jand g19765(.dina(n20022), .dinb(n20019), .dout(n20023));
  jor  g19766(.dina(n20023), .dinb(n20018), .dout(n20024));
  jand g19767(.dina(n20024), .dinb(asqrt[40] ), .dout(n20025));
  jor  g19768(.dina(n20024), .dinb(asqrt[40] ), .dout(n20026));
  jxor g19769(.dina(n19328), .dinb(n4249), .dout(n20027));
  jand g19770(.dina(n20027), .dinb(asqrt[8] ), .dout(n20028));
  jxor g19771(.dina(n20028), .dinb(n19333), .dout(n20029));
  jnot g19772(.din(n20029), .dout(n20030));
  jand g19773(.dina(n20030), .dinb(n20026), .dout(n20031));
  jor  g19774(.dina(n20031), .dinb(n20025), .dout(n20032));
  jand g19775(.dina(n20032), .dinb(asqrt[41] ), .dout(n20033));
  jor  g19776(.dina(n20032), .dinb(asqrt[41] ), .dout(n20034));
  jxor g19777(.dina(n19335), .dinb(n3955), .dout(n20035));
  jand g19778(.dina(n20035), .dinb(asqrt[8] ), .dout(n20036));
  jxor g19779(.dina(n20036), .dinb(n19340), .dout(n20037));
  jnot g19780(.din(n20037), .dout(n20038));
  jand g19781(.dina(n20038), .dinb(n20034), .dout(n20039));
  jor  g19782(.dina(n20039), .dinb(n20033), .dout(n20040));
  jand g19783(.dina(n20040), .dinb(asqrt[42] ), .dout(n20041));
  jor  g19784(.dina(n20040), .dinb(asqrt[42] ), .dout(n20042));
  jxor g19785(.dina(n19342), .dinb(n3642), .dout(n20043));
  jand g19786(.dina(n20043), .dinb(asqrt[8] ), .dout(n20044));
  jxor g19787(.dina(n20044), .dinb(n19347), .dout(n20045));
  jnot g19788(.din(n20045), .dout(n20046));
  jand g19789(.dina(n20046), .dinb(n20042), .dout(n20047));
  jor  g19790(.dina(n20047), .dinb(n20041), .dout(n20048));
  jand g19791(.dina(n20048), .dinb(asqrt[43] ), .dout(n20049));
  jor  g19792(.dina(n20048), .dinb(asqrt[43] ), .dout(n20050));
  jxor g19793(.dina(n19349), .dinb(n3368), .dout(n20051));
  jand g19794(.dina(n20051), .dinb(asqrt[8] ), .dout(n20052));
  jxor g19795(.dina(n20052), .dinb(n19354), .dout(n20053));
  jand g19796(.dina(n20053), .dinb(n20050), .dout(n20054));
  jor  g19797(.dina(n20054), .dinb(n20049), .dout(n20055));
  jand g19798(.dina(n20055), .dinb(asqrt[44] ), .dout(n20056));
  jor  g19799(.dina(n20055), .dinb(asqrt[44] ), .dout(n20057));
  jxor g19800(.dina(n19357), .dinb(n3089), .dout(n20058));
  jand g19801(.dina(n20058), .dinb(asqrt[8] ), .dout(n20059));
  jxor g19802(.dina(n20059), .dinb(n19362), .dout(n20060));
  jnot g19803(.din(n20060), .dout(n20061));
  jand g19804(.dina(n20061), .dinb(n20057), .dout(n20062));
  jor  g19805(.dina(n20062), .dinb(n20056), .dout(n20063));
  jand g19806(.dina(n20063), .dinb(asqrt[45] ), .dout(n20064));
  jor  g19807(.dina(n20063), .dinb(asqrt[45] ), .dout(n20065));
  jxor g19808(.dina(n19364), .dinb(n2833), .dout(n20066));
  jand g19809(.dina(n20066), .dinb(asqrt[8] ), .dout(n20067));
  jxor g19810(.dina(n20067), .dinb(n19369), .dout(n20068));
  jnot g19811(.din(n20068), .dout(n20069));
  jand g19812(.dina(n20069), .dinb(n20065), .dout(n20070));
  jor  g19813(.dina(n20070), .dinb(n20064), .dout(n20071));
  jand g19814(.dina(n20071), .dinb(asqrt[46] ), .dout(n20072));
  jor  g19815(.dina(n20071), .dinb(asqrt[46] ), .dout(n20073));
  jxor g19816(.dina(n19371), .dinb(n2572), .dout(n20074));
  jand g19817(.dina(n20074), .dinb(asqrt[8] ), .dout(n20075));
  jxor g19818(.dina(n20075), .dinb(n19376), .dout(n20076));
  jnot g19819(.din(n20076), .dout(n20077));
  jand g19820(.dina(n20077), .dinb(n20073), .dout(n20078));
  jor  g19821(.dina(n20078), .dinb(n20072), .dout(n20079));
  jand g19822(.dina(n20079), .dinb(asqrt[47] ), .dout(n20080));
  jor  g19823(.dina(n20079), .dinb(asqrt[47] ), .dout(n20081));
  jxor g19824(.dina(n19378), .dinb(n2345), .dout(n20082));
  jand g19825(.dina(n20082), .dinb(asqrt[8] ), .dout(n20083));
  jxor g19826(.dina(n20083), .dinb(n19383), .dout(n20084));
  jnot g19827(.din(n20084), .dout(n20085));
  jand g19828(.dina(n20085), .dinb(n20081), .dout(n20086));
  jor  g19829(.dina(n20086), .dinb(n20080), .dout(n20087));
  jand g19830(.dina(n20087), .dinb(asqrt[48] ), .dout(n20088));
  jor  g19831(.dina(n20087), .dinb(asqrt[48] ), .dout(n20089));
  jxor g19832(.dina(n19385), .dinb(n2108), .dout(n20090));
  jand g19833(.dina(n20090), .dinb(asqrt[8] ), .dout(n20091));
  jxor g19834(.dina(n20091), .dinb(n19390), .dout(n20092));
  jnot g19835(.din(n20092), .dout(n20093));
  jand g19836(.dina(n20093), .dinb(n20089), .dout(n20094));
  jor  g19837(.dina(n20094), .dinb(n20088), .dout(n20095));
  jand g19838(.dina(n20095), .dinb(asqrt[49] ), .dout(n20096));
  jor  g19839(.dina(n20095), .dinb(asqrt[49] ), .dout(n20097));
  jxor g19840(.dina(n19392), .dinb(n1912), .dout(n20098));
  jand g19841(.dina(n20098), .dinb(asqrt[8] ), .dout(n20099));
  jxor g19842(.dina(n20099), .dinb(n19397), .dout(n20100));
  jand g19843(.dina(n20100), .dinb(n20097), .dout(n20101));
  jor  g19844(.dina(n20101), .dinb(n20096), .dout(n20102));
  jand g19845(.dina(n20102), .dinb(asqrt[50] ), .dout(n20103));
  jor  g19846(.dina(n20102), .dinb(asqrt[50] ), .dout(n20104));
  jxor g19847(.dina(n19400), .dinb(n1699), .dout(n20105));
  jand g19848(.dina(n20105), .dinb(asqrt[8] ), .dout(n20106));
  jxor g19849(.dina(n20106), .dinb(n19405), .dout(n20107));
  jnot g19850(.din(n20107), .dout(n20108));
  jand g19851(.dina(n20108), .dinb(n20104), .dout(n20109));
  jor  g19852(.dina(n20109), .dinb(n20103), .dout(n20110));
  jand g19853(.dina(n20110), .dinb(asqrt[51] ), .dout(n20111));
  jor  g19854(.dina(n20110), .dinb(asqrt[51] ), .dout(n20112));
  jxor g19855(.dina(n19407), .dinb(n1516), .dout(n20113));
  jand g19856(.dina(n20113), .dinb(asqrt[8] ), .dout(n20114));
  jxor g19857(.dina(n20114), .dinb(n19412), .dout(n20115));
  jand g19858(.dina(n20115), .dinb(n20112), .dout(n20116));
  jor  g19859(.dina(n20116), .dinb(n20111), .dout(n20117));
  jand g19860(.dina(n20117), .dinb(asqrt[52] ), .dout(n20118));
  jor  g19861(.dina(n20117), .dinb(asqrt[52] ), .dout(n20119));
  jxor g19862(.dina(n19415), .dinb(n1332), .dout(n20120));
  jand g19863(.dina(n20120), .dinb(asqrt[8] ), .dout(n20121));
  jxor g19864(.dina(n20121), .dinb(n19420), .dout(n20122));
  jnot g19865(.din(n20122), .dout(n20123));
  jand g19866(.dina(n20123), .dinb(n20119), .dout(n20124));
  jor  g19867(.dina(n20124), .dinb(n20118), .dout(n20125));
  jand g19868(.dina(n20125), .dinb(asqrt[53] ), .dout(n20126));
  jor  g19869(.dina(n20125), .dinb(asqrt[53] ), .dout(n20127));
  jxor g19870(.dina(n19422), .dinb(n1173), .dout(n20128));
  jand g19871(.dina(n20128), .dinb(asqrt[8] ), .dout(n20129));
  jxor g19872(.dina(n20129), .dinb(n19427), .dout(n20130));
  jnot g19873(.din(n20130), .dout(n20131));
  jand g19874(.dina(n20131), .dinb(n20127), .dout(n20132));
  jor  g19875(.dina(n20132), .dinb(n20126), .dout(n20133));
  jand g19876(.dina(n20133), .dinb(asqrt[54] ), .dout(n20134));
  jor  g19877(.dina(n20133), .dinb(asqrt[54] ), .dout(n20135));
  jxor g19878(.dina(n19429), .dinb(n1008), .dout(n20136));
  jand g19879(.dina(n20136), .dinb(asqrt[8] ), .dout(n20137));
  jxor g19880(.dina(n20137), .dinb(n19434), .dout(n20138));
  jand g19881(.dina(n20138), .dinb(n20135), .dout(n20139));
  jor  g19882(.dina(n20139), .dinb(n20134), .dout(n20140));
  jand g19883(.dina(n20140), .dinb(asqrt[55] ), .dout(n20141));
  jxor g19884(.dina(n19437), .dinb(n884), .dout(n20142));
  jand g19885(.dina(n20142), .dinb(asqrt[8] ), .dout(n20143));
  jxor g19886(.dina(n20143), .dinb(n19441), .dout(n20144));
  jor  g19887(.dina(n20140), .dinb(asqrt[55] ), .dout(n20145));
  jand g19888(.dina(n20145), .dinb(n20144), .dout(n20146));
  jor  g19889(.dina(n20146), .dinb(n20141), .dout(n20147));
  jand g19890(.dina(n20147), .dinb(asqrt[56] ), .dout(n20148));
  jor  g19891(.dina(n20147), .dinb(asqrt[56] ), .dout(n20149));
  jxor g19892(.dina(n19445), .dinb(n743), .dout(n20150));
  jand g19893(.dina(n20150), .dinb(asqrt[8] ), .dout(n20151));
  jxor g19894(.dina(n20151), .dinb(n19450), .dout(n20152));
  jnot g19895(.din(n20152), .dout(n20153));
  jand g19896(.dina(n20153), .dinb(n20149), .dout(n20154));
  jor  g19897(.dina(n20154), .dinb(n20148), .dout(n20155));
  jand g19898(.dina(n20155), .dinb(asqrt[57] ), .dout(n20156));
  jor  g19899(.dina(n20155), .dinb(asqrt[57] ), .dout(n20157));
  jxor g19900(.dina(n19452), .dinb(n635), .dout(n20158));
  jand g19901(.dina(n20158), .dinb(asqrt[8] ), .dout(n20159));
  jxor g19902(.dina(n20159), .dinb(n19457), .dout(n20160));
  jand g19903(.dina(n20160), .dinb(n20157), .dout(n20161));
  jor  g19904(.dina(n20161), .dinb(n20156), .dout(n20162));
  jand g19905(.dina(n20162), .dinb(asqrt[58] ), .dout(n20163));
  jor  g19906(.dina(n20162), .dinb(asqrt[58] ), .dout(n20164));
  jxor g19907(.dina(n19460), .dinb(n515), .dout(n20165));
  jand g19908(.dina(n20165), .dinb(asqrt[8] ), .dout(n20166));
  jxor g19909(.dina(n20166), .dinb(n19465), .dout(n20167));
  jnot g19910(.din(n20167), .dout(n20168));
  jand g19911(.dina(n20168), .dinb(n20164), .dout(n20169));
  jor  g19912(.dina(n20169), .dinb(n20163), .dout(n20170));
  jand g19913(.dina(n20170), .dinb(asqrt[59] ), .dout(n20171));
  jor  g19914(.dina(n20170), .dinb(asqrt[59] ), .dout(n20172));
  jxor g19915(.dina(n19467), .dinb(n443), .dout(n20173));
  jand g19916(.dina(n20173), .dinb(asqrt[8] ), .dout(n20174));
  jxor g19917(.dina(n20174), .dinb(n19473), .dout(n20175));
  jnot g19918(.din(n20175), .dout(n20176));
  jand g19919(.dina(n20176), .dinb(n20172), .dout(n20177));
  jor  g19920(.dina(n20177), .dinb(n20171), .dout(n20178));
  jand g19921(.dina(n20178), .dinb(asqrt[60] ), .dout(n20179));
  jor  g19922(.dina(n20178), .dinb(asqrt[60] ), .dout(n20180));
  jxor g19923(.dina(n19475), .dinb(n352), .dout(n20181));
  jand g19924(.dina(n20181), .dinb(asqrt[8] ), .dout(n20182));
  jxor g19925(.dina(n20182), .dinb(n19480), .dout(n20183));
  jand g19926(.dina(n20183), .dinb(n20180), .dout(n20184));
  jor  g19927(.dina(n20184), .dinb(n20179), .dout(n20185));
  jand g19928(.dina(n20185), .dinb(asqrt[61] ), .dout(n20186));
  jor  g19929(.dina(n20185), .dinb(asqrt[61] ), .dout(n20187));
  jxor g19930(.dina(n19483), .dinb(n294), .dout(n20188));
  jand g19931(.dina(n20188), .dinb(asqrt[8] ), .dout(n20189));
  jxor g19932(.dina(n20189), .dinb(n19488), .dout(n20190));
  jnot g19933(.din(n20190), .dout(n20191));
  jand g19934(.dina(n20191), .dinb(n20187), .dout(n20192));
  jor  g19935(.dina(n20192), .dinb(n20186), .dout(n20193));
  jand g19936(.dina(n20193), .dinb(asqrt[62] ), .dout(n20194));
  jnot g19937(.din(n20194), .dout(n20195));
  jnot g19938(.din(n20186), .dout(n20196));
  jnot g19939(.din(n20179), .dout(n20197));
  jnot g19940(.din(n20171), .dout(n20198));
  jnot g19941(.din(n20163), .dout(n20199));
  jnot g19942(.din(n20156), .dout(n20200));
  jnot g19943(.din(n20148), .dout(n20201));
  jnot g19944(.din(n20141), .dout(n20202));
  jnot g19945(.din(n20144), .dout(n20203));
  jnot g19946(.din(n20134), .dout(n20204));
  jnot g19947(.din(n20126), .dout(n20205));
  jnot g19948(.din(n20118), .dout(n20206));
  jnot g19949(.din(n20111), .dout(n20207));
  jnot g19950(.din(n20103), .dout(n20208));
  jnot g19951(.din(n20096), .dout(n20209));
  jnot g19952(.din(n20088), .dout(n20210));
  jnot g19953(.din(n20080), .dout(n20211));
  jnot g19954(.din(n20072), .dout(n20212));
  jnot g19955(.din(n20064), .dout(n20213));
  jnot g19956(.din(n20056), .dout(n20214));
  jnot g19957(.din(n20049), .dout(n20215));
  jnot g19958(.din(n20041), .dout(n20216));
  jnot g19959(.din(n20033), .dout(n20217));
  jnot g19960(.din(n20025), .dout(n20218));
  jnot g19961(.din(n20018), .dout(n20219));
  jnot g19962(.din(n20010), .dout(n20220));
  jnot g19963(.din(n20003), .dout(n20221));
  jnot g19964(.din(n19995), .dout(n20222));
  jnot g19965(.din(n19988), .dout(n20223));
  jnot g19966(.din(n19980), .dout(n20224));
  jnot g19967(.din(n19973), .dout(n20225));
  jnot g19968(.din(n19965), .dout(n20226));
  jnot g19969(.din(n19957), .dout(n20227));
  jnot g19970(.din(n19949), .dout(n20228));
  jnot g19971(.din(n19942), .dout(n20229));
  jnot g19972(.din(n19934), .dout(n20230));
  jnot g19973(.din(n19927), .dout(n20231));
  jnot g19974(.din(n19919), .dout(n20232));
  jnot g19975(.din(n19912), .dout(n20233));
  jnot g19976(.din(n19905), .dout(n20234));
  jnot g19977(.din(n19897), .dout(n20235));
  jnot g19978(.din(n19889), .dout(n20236));
  jnot g19979(.din(n19882), .dout(n20237));
  jnot g19980(.din(n19874), .dout(n20238));
  jnot g19981(.din(n19867), .dout(n20239));
  jnot g19982(.din(n19859), .dout(n20240));
  jnot g19983(.din(n19852), .dout(n20241));
  jnot g19984(.din(n19844), .dout(n20242));
  jnot g19985(.din(n19837), .dout(n20243));
  jnot g19986(.din(n19829), .dout(n20244));
  jnot g19987(.din(n19822), .dout(n20245));
  jnot g19988(.din(n19814), .dout(n20246));
  jnot g19989(.din(n19806), .dout(n20247));
  jnot g19990(.din(n19796), .dout(n20248));
  jnot g19991(.din(n19530), .dout(n20249));
  jnot g19992(.din(n19527), .dout(n20250));
  jor  g19993(.dina(n19791), .dinb(n19101), .dout(n20251));
  jand g19994(.dina(n20251), .dinb(n20250), .dout(n20252));
  jand g19995(.dina(n20252), .dinb(n19096), .dout(n20253));
  jor  g19996(.dina(n19791), .dinb(a[16] ), .dout(n20254));
  jand g19997(.dina(n20254), .dinb(a[17] ), .dout(n20255));
  jor  g19998(.dina(n19798), .dinb(n20255), .dout(n20256));
  jor  g19999(.dina(n20256), .dinb(n20253), .dout(n20257));
  jand g20000(.dina(n20257), .dinb(n20249), .dout(n20258));
  jand g20001(.dina(n20258), .dinb(n18442), .dout(n20259));
  jor  g20002(.dina(n19802), .dinb(n20259), .dout(n20260));
  jand g20003(.dina(n20260), .dinb(n20248), .dout(n20261));
  jand g20004(.dina(n20261), .dinb(n17769), .dout(n20262));
  jor  g20005(.dina(n19810), .dinb(n20262), .dout(n20263));
  jand g20006(.dina(n20263), .dinb(n20247), .dout(n20264));
  jand g20007(.dina(n20264), .dinb(n17134), .dout(n20265));
  jor  g20008(.dina(n19818), .dinb(n20265), .dout(n20266));
  jand g20009(.dina(n20266), .dinb(n20246), .dout(n20267));
  jand g20010(.dina(n20267), .dinb(n16489), .dout(n20268));
  jnot g20011(.din(n19826), .dout(n20269));
  jor  g20012(.dina(n20269), .dinb(n20268), .dout(n20270));
  jand g20013(.dina(n20270), .dinb(n20245), .dout(n20271));
  jand g20014(.dina(n20271), .dinb(n15878), .dout(n20272));
  jor  g20015(.dina(n19833), .dinb(n20272), .dout(n20273));
  jand g20016(.dina(n20273), .dinb(n20244), .dout(n20274));
  jand g20017(.dina(n20274), .dinb(n15260), .dout(n20275));
  jnot g20018(.din(n19841), .dout(n20276));
  jor  g20019(.dina(n20276), .dinb(n20275), .dout(n20277));
  jand g20020(.dina(n20277), .dinb(n20243), .dout(n20278));
  jand g20021(.dina(n20278), .dinb(n14674), .dout(n20279));
  jor  g20022(.dina(n19848), .dinb(n20279), .dout(n20280));
  jand g20023(.dina(n20280), .dinb(n20242), .dout(n20281));
  jand g20024(.dina(n20281), .dinb(n14078), .dout(n20282));
  jnot g20025(.din(n19856), .dout(n20283));
  jor  g20026(.dina(n20283), .dinb(n20282), .dout(n20284));
  jand g20027(.dina(n20284), .dinb(n20241), .dout(n20285));
  jand g20028(.dina(n20285), .dinb(n13515), .dout(n20286));
  jor  g20029(.dina(n19863), .dinb(n20286), .dout(n20287));
  jand g20030(.dina(n20287), .dinb(n20240), .dout(n20288));
  jand g20031(.dina(n20288), .dinb(n12947), .dout(n20289));
  jnot g20032(.din(n19871), .dout(n20290));
  jor  g20033(.dina(n20290), .dinb(n20289), .dout(n20291));
  jand g20034(.dina(n20291), .dinb(n20239), .dout(n20292));
  jand g20035(.dina(n20292), .dinb(n12410), .dout(n20293));
  jor  g20036(.dina(n19878), .dinb(n20293), .dout(n20294));
  jand g20037(.dina(n20294), .dinb(n20238), .dout(n20295));
  jand g20038(.dina(n20295), .dinb(n11858), .dout(n20296));
  jnot g20039(.din(n19886), .dout(n20297));
  jor  g20040(.dina(n20297), .dinb(n20296), .dout(n20298));
  jand g20041(.dina(n20298), .dinb(n20237), .dout(n20299));
  jand g20042(.dina(n20299), .dinb(n11347), .dout(n20300));
  jor  g20043(.dina(n19893), .dinb(n20300), .dout(n20301));
  jand g20044(.dina(n20301), .dinb(n20236), .dout(n20302));
  jand g20045(.dina(n20302), .dinb(n10824), .dout(n20303));
  jor  g20046(.dina(n19901), .dinb(n20303), .dout(n20304));
  jand g20047(.dina(n20304), .dinb(n20235), .dout(n20305));
  jand g20048(.dina(n20305), .dinb(n10328), .dout(n20306));
  jnot g20049(.din(n19909), .dout(n20307));
  jor  g20050(.dina(n20307), .dinb(n20306), .dout(n20308));
  jand g20051(.dina(n20308), .dinb(n20234), .dout(n20309));
  jand g20052(.dina(n20309), .dinb(n9832), .dout(n20310));
  jnot g20053(.din(n19916), .dout(n20311));
  jor  g20054(.dina(n20311), .dinb(n20310), .dout(n20312));
  jand g20055(.dina(n20312), .dinb(n20233), .dout(n20313));
  jand g20056(.dina(n20313), .dinb(n9369), .dout(n20314));
  jor  g20057(.dina(n19923), .dinb(n20314), .dout(n20315));
  jand g20058(.dina(n20315), .dinb(n20232), .dout(n20316));
  jand g20059(.dina(n20316), .dinb(n8890), .dout(n20317));
  jnot g20060(.din(n19931), .dout(n20318));
  jor  g20061(.dina(n20318), .dinb(n20317), .dout(n20319));
  jand g20062(.dina(n20319), .dinb(n20231), .dout(n20320));
  jand g20063(.dina(n20320), .dinb(n8449), .dout(n20321));
  jor  g20064(.dina(n19938), .dinb(n20321), .dout(n20322));
  jand g20065(.dina(n20322), .dinb(n20230), .dout(n20323));
  jand g20066(.dina(n20323), .dinb(n8003), .dout(n20324));
  jnot g20067(.din(n19946), .dout(n20325));
  jor  g20068(.dina(n20325), .dinb(n20324), .dout(n20326));
  jand g20069(.dina(n20326), .dinb(n20229), .dout(n20327));
  jand g20070(.dina(n20327), .dinb(n7581), .dout(n20328));
  jor  g20071(.dina(n19953), .dinb(n20328), .dout(n20329));
  jand g20072(.dina(n20329), .dinb(n20228), .dout(n20330));
  jand g20073(.dina(n20330), .dinb(n7154), .dout(n20331));
  jor  g20074(.dina(n19961), .dinb(n20331), .dout(n20332));
  jand g20075(.dina(n20332), .dinb(n20227), .dout(n20333));
  jand g20076(.dina(n20333), .dinb(n6758), .dout(n20334));
  jor  g20077(.dina(n19969), .dinb(n20334), .dout(n20335));
  jand g20078(.dina(n20335), .dinb(n20226), .dout(n20336));
  jand g20079(.dina(n20336), .dinb(n6357), .dout(n20337));
  jnot g20080(.din(n19977), .dout(n20338));
  jor  g20081(.dina(n20338), .dinb(n20337), .dout(n20339));
  jand g20082(.dina(n20339), .dinb(n20225), .dout(n20340));
  jand g20083(.dina(n20340), .dinb(n5989), .dout(n20341));
  jor  g20084(.dina(n19984), .dinb(n20341), .dout(n20342));
  jand g20085(.dina(n20342), .dinb(n20224), .dout(n20343));
  jand g20086(.dina(n20343), .dinb(n5606), .dout(n20344));
  jnot g20087(.din(n19992), .dout(n20345));
  jor  g20088(.dina(n20345), .dinb(n20344), .dout(n20346));
  jand g20089(.dina(n20346), .dinb(n20223), .dout(n20347));
  jand g20090(.dina(n20347), .dinb(n5259), .dout(n20348));
  jor  g20091(.dina(n19999), .dinb(n20348), .dout(n20349));
  jand g20092(.dina(n20349), .dinb(n20222), .dout(n20350));
  jand g20093(.dina(n20350), .dinb(n4902), .dout(n20351));
  jnot g20094(.din(n20007), .dout(n20352));
  jor  g20095(.dina(n20352), .dinb(n20351), .dout(n20353));
  jand g20096(.dina(n20353), .dinb(n20221), .dout(n20354));
  jand g20097(.dina(n20354), .dinb(n4582), .dout(n20355));
  jor  g20098(.dina(n20014), .dinb(n20355), .dout(n20356));
  jand g20099(.dina(n20356), .dinb(n20220), .dout(n20357));
  jand g20100(.dina(n20357), .dinb(n4249), .dout(n20358));
  jnot g20101(.din(n20022), .dout(n20359));
  jor  g20102(.dina(n20359), .dinb(n20358), .dout(n20360));
  jand g20103(.dina(n20360), .dinb(n20219), .dout(n20361));
  jand g20104(.dina(n20361), .dinb(n3955), .dout(n20362));
  jor  g20105(.dina(n20029), .dinb(n20362), .dout(n20363));
  jand g20106(.dina(n20363), .dinb(n20218), .dout(n20364));
  jand g20107(.dina(n20364), .dinb(n3642), .dout(n20365));
  jor  g20108(.dina(n20037), .dinb(n20365), .dout(n20366));
  jand g20109(.dina(n20366), .dinb(n20217), .dout(n20367));
  jand g20110(.dina(n20367), .dinb(n3368), .dout(n20368));
  jor  g20111(.dina(n20045), .dinb(n20368), .dout(n20369));
  jand g20112(.dina(n20369), .dinb(n20216), .dout(n20370));
  jand g20113(.dina(n20370), .dinb(n3089), .dout(n20371));
  jnot g20114(.din(n20053), .dout(n20372));
  jor  g20115(.dina(n20372), .dinb(n20371), .dout(n20373));
  jand g20116(.dina(n20373), .dinb(n20215), .dout(n20374));
  jand g20117(.dina(n20374), .dinb(n2833), .dout(n20375));
  jor  g20118(.dina(n20060), .dinb(n20375), .dout(n20376));
  jand g20119(.dina(n20376), .dinb(n20214), .dout(n20377));
  jand g20120(.dina(n20377), .dinb(n2572), .dout(n20378));
  jor  g20121(.dina(n20068), .dinb(n20378), .dout(n20379));
  jand g20122(.dina(n20379), .dinb(n20213), .dout(n20380));
  jand g20123(.dina(n20380), .dinb(n2345), .dout(n20381));
  jor  g20124(.dina(n20076), .dinb(n20381), .dout(n20382));
  jand g20125(.dina(n20382), .dinb(n20212), .dout(n20383));
  jand g20126(.dina(n20383), .dinb(n2108), .dout(n20384));
  jor  g20127(.dina(n20084), .dinb(n20384), .dout(n20385));
  jand g20128(.dina(n20385), .dinb(n20211), .dout(n20386));
  jand g20129(.dina(n20386), .dinb(n1912), .dout(n20387));
  jor  g20130(.dina(n20092), .dinb(n20387), .dout(n20388));
  jand g20131(.dina(n20388), .dinb(n20210), .dout(n20389));
  jand g20132(.dina(n20389), .dinb(n1699), .dout(n20390));
  jnot g20133(.din(n20100), .dout(n20391));
  jor  g20134(.dina(n20391), .dinb(n20390), .dout(n20392));
  jand g20135(.dina(n20392), .dinb(n20209), .dout(n20393));
  jand g20136(.dina(n20393), .dinb(n1516), .dout(n20394));
  jor  g20137(.dina(n20107), .dinb(n20394), .dout(n20395));
  jand g20138(.dina(n20395), .dinb(n20208), .dout(n20396));
  jand g20139(.dina(n20396), .dinb(n1332), .dout(n20397));
  jnot g20140(.din(n20115), .dout(n20398));
  jor  g20141(.dina(n20398), .dinb(n20397), .dout(n20399));
  jand g20142(.dina(n20399), .dinb(n20207), .dout(n20400));
  jand g20143(.dina(n20400), .dinb(n1173), .dout(n20401));
  jor  g20144(.dina(n20122), .dinb(n20401), .dout(n20402));
  jand g20145(.dina(n20402), .dinb(n20206), .dout(n20403));
  jand g20146(.dina(n20403), .dinb(n1008), .dout(n20404));
  jor  g20147(.dina(n20130), .dinb(n20404), .dout(n20405));
  jand g20148(.dina(n20405), .dinb(n20205), .dout(n20406));
  jand g20149(.dina(n20406), .dinb(n884), .dout(n20407));
  jnot g20150(.din(n20138), .dout(n20408));
  jor  g20151(.dina(n20408), .dinb(n20407), .dout(n20409));
  jand g20152(.dina(n20409), .dinb(n20204), .dout(n20410));
  jand g20153(.dina(n20410), .dinb(n743), .dout(n20411));
  jor  g20154(.dina(n20411), .dinb(n20203), .dout(n20412));
  jand g20155(.dina(n20412), .dinb(n20202), .dout(n20413));
  jand g20156(.dina(n20413), .dinb(n635), .dout(n20414));
  jor  g20157(.dina(n20152), .dinb(n20414), .dout(n20415));
  jand g20158(.dina(n20415), .dinb(n20201), .dout(n20416));
  jand g20159(.dina(n20416), .dinb(n515), .dout(n20417));
  jnot g20160(.din(n20160), .dout(n20418));
  jor  g20161(.dina(n20418), .dinb(n20417), .dout(n20419));
  jand g20162(.dina(n20419), .dinb(n20200), .dout(n20420));
  jand g20163(.dina(n20420), .dinb(n443), .dout(n20421));
  jor  g20164(.dina(n20167), .dinb(n20421), .dout(n20422));
  jand g20165(.dina(n20422), .dinb(n20199), .dout(n20423));
  jand g20166(.dina(n20423), .dinb(n352), .dout(n20424));
  jor  g20167(.dina(n20175), .dinb(n20424), .dout(n20425));
  jand g20168(.dina(n20425), .dinb(n20198), .dout(n20426));
  jand g20169(.dina(n20426), .dinb(n294), .dout(n20427));
  jnot g20170(.din(n20183), .dout(n20428));
  jor  g20171(.dina(n20428), .dinb(n20427), .dout(n20429));
  jand g20172(.dina(n20429), .dinb(n20197), .dout(n20430));
  jand g20173(.dina(n20430), .dinb(n239), .dout(n20431));
  jor  g20174(.dina(n20190), .dinb(n20431), .dout(n20432));
  jand g20175(.dina(n20432), .dinb(n20196), .dout(n20433));
  jand g20176(.dina(n20433), .dinb(n221), .dout(n20434));
  jxor g20177(.dina(n19490), .dinb(n239), .dout(n20435));
  jand g20178(.dina(n20435), .dinb(asqrt[8] ), .dout(n20436));
  jxor g20179(.dina(n20436), .dinb(n19495), .dout(n20437));
  jor  g20180(.dina(n20437), .dinb(n20434), .dout(n20438));
  jand g20181(.dina(n20438), .dinb(n20195), .dout(n20439));
  jor  g20182(.dina(n20439), .dinb(n19523), .dout(n20440));
  jand g20183(.dina(asqrt[8] ), .dinb(n19782), .dout(n20441));
  jor  g20184(.dina(n20441), .dinb(n19511), .dout(n20442));
  jor  g20185(.dina(n20442), .dinb(n20440), .dout(n20443));
  jand g20186(.dina(n20443), .dinb(n218), .dout(n20444));
  jand g20187(.dina(n19791), .dinb(n19100), .dout(n20445));
  jand g20188(.dina(n20439), .dinb(n19523), .dout(n20446));
  jor  g20189(.dina(n20446), .dinb(n20445), .dout(n20447));
  jand g20190(.dina(n19791), .dinb(n19505), .dout(n20448));
  jnot g20191(.din(n20448), .dout(n20449));
  jand g20192(.dina(n19786), .dinb(asqrt[63] ), .dout(n20450));
  jand g20193(.dina(n20450), .dinb(n19506), .dout(n20451));
  jand g20194(.dina(n20451), .dinb(n20449), .dout(n20452));
  jor  g20195(.dina(n20452), .dinb(n20447), .dout(n20453));
  jor  g20196(.dina(n20453), .dinb(n20444), .dout(asqrt[7] ));
  jor  g20197(.dina(n20193), .dinb(asqrt[62] ), .dout(n20455));
  jnot g20198(.din(n20437), .dout(n20456));
  jand g20199(.dina(n20456), .dinb(n20455), .dout(n20457));
  jor  g20200(.dina(n20457), .dinb(n20194), .dout(n20458));
  jand g20201(.dina(n20458), .dinb(n19522), .dout(n20459));
  jnot g20202(.din(n20442), .dout(n20460));
  jand g20203(.dina(n20460), .dinb(n20459), .dout(n20461));
  jor  g20204(.dina(n20461), .dinb(asqrt[63] ), .dout(n20462));
  jnot g20205(.din(n20445), .dout(n20463));
  jor  g20206(.dina(n20458), .dinb(n19522), .dout(n20464));
  jand g20207(.dina(n20464), .dinb(n20463), .dout(n20465));
  jnot g20208(.din(n20452), .dout(n20466));
  jand g20209(.dina(n20466), .dinb(n20465), .dout(n20467));
  jand g20210(.dina(n20467), .dinb(n20462), .dout(n20468));
  jxor g20211(.dina(n20193), .dinb(n221), .dout(n20469));
  jor  g20212(.dina(n20469), .dinb(n20468), .dout(n20470));
  jxor g20213(.dina(n20470), .dinb(n20437), .dout(n20471));
  jnot g20214(.din(n20471), .dout(n20472));
  jnot g20215(.din(a[12] ), .dout(n20473));
  jnot g20216(.din(a[13] ), .dout(n20474));
  jand g20217(.dina(n20474), .dinb(n20473), .dout(n20475));
  jand g20218(.dina(n20475), .dinb(n19524), .dout(n20476));
  jnot g20219(.din(n20476), .dout(n20477));
  jor  g20220(.dina(n20468), .dinb(n19524), .dout(n20478));
  jand g20221(.dina(n20478), .dinb(n20477), .dout(n20479));
  jor  g20222(.dina(n20479), .dinb(n19791), .dout(n20480));
  jand g20223(.dina(n20479), .dinb(n19791), .dout(n20481));
  jor  g20224(.dina(n20468), .dinb(a[14] ), .dout(n20482));
  jand g20225(.dina(n20482), .dinb(a[15] ), .dout(n20483));
  jand g20226(.dina(asqrt[7] ), .dinb(n19526), .dout(n20484));
  jor  g20227(.dina(n20484), .dinb(n20483), .dout(n20485));
  jor  g20228(.dina(n20485), .dinb(n20481), .dout(n20486));
  jand g20229(.dina(n20486), .dinb(n20480), .dout(n20487));
  jor  g20230(.dina(n20487), .dinb(n19096), .dout(n20488));
  jand g20231(.dina(n20487), .dinb(n19096), .dout(n20489));
  jnot g20232(.din(n19526), .dout(n20490));
  jor  g20233(.dina(n20468), .dinb(n20490), .dout(n20491));
  jor  g20234(.dina(n20451), .dinb(n20446), .dout(n20492));
  jor  g20235(.dina(n20492), .dinb(n20444), .dout(n20493));
  jor  g20236(.dina(n20493), .dinb(n19791), .dout(n20494));
  jand g20237(.dina(n20494), .dinb(n20491), .dout(n20495));
  jxor g20238(.dina(n20495), .dinb(n19101), .dout(n20496));
  jor  g20239(.dina(n20496), .dinb(n20489), .dout(n20497));
  jand g20240(.dina(n20497), .dinb(n20488), .dout(n20498));
  jor  g20241(.dina(n20498), .dinb(n18442), .dout(n20499));
  jand g20242(.dina(n20498), .dinb(n18442), .dout(n20500));
  jxor g20243(.dina(n19529), .dinb(n19096), .dout(n20501));
  jor  g20244(.dina(n20501), .dinb(n20468), .dout(n20502));
  jxor g20245(.dina(n20502), .dinb(n20256), .dout(n20503));
  jnot g20246(.din(n20503), .dout(n20504));
  jor  g20247(.dina(n20504), .dinb(n20500), .dout(n20505));
  jand g20248(.dina(n20505), .dinb(n20499), .dout(n20506));
  jor  g20249(.dina(n20506), .dinb(n17769), .dout(n20507));
  jand g20250(.dina(n20506), .dinb(n17769), .dout(n20508));
  jxor g20251(.dina(n19795), .dinb(n18442), .dout(n20509));
  jor  g20252(.dina(n20509), .dinb(n20468), .dout(n20510));
  jxor g20253(.dina(n20510), .dinb(n19803), .dout(n20511));
  jor  g20254(.dina(n20511), .dinb(n20508), .dout(n20512));
  jand g20255(.dina(n20512), .dinb(n20507), .dout(n20513));
  jor  g20256(.dina(n20513), .dinb(n17134), .dout(n20514));
  jand g20257(.dina(n20513), .dinb(n17134), .dout(n20515));
  jxor g20258(.dina(n19805), .dinb(n17769), .dout(n20516));
  jor  g20259(.dina(n20516), .dinb(n20468), .dout(n20517));
  jxor g20260(.dina(n20517), .dinb(n19811), .dout(n20518));
  jor  g20261(.dina(n20518), .dinb(n20515), .dout(n20519));
  jand g20262(.dina(n20519), .dinb(n20514), .dout(n20520));
  jor  g20263(.dina(n20520), .dinb(n16489), .dout(n20521));
  jand g20264(.dina(n20520), .dinb(n16489), .dout(n20522));
  jxor g20265(.dina(n19813), .dinb(n17134), .dout(n20523));
  jor  g20266(.dina(n20523), .dinb(n20468), .dout(n20524));
  jxor g20267(.dina(n20524), .dinb(n19819), .dout(n20525));
  jor  g20268(.dina(n20525), .dinb(n20522), .dout(n20526));
  jand g20269(.dina(n20526), .dinb(n20521), .dout(n20527));
  jor  g20270(.dina(n20527), .dinb(n15878), .dout(n20528));
  jand g20271(.dina(n20527), .dinb(n15878), .dout(n20529));
  jxor g20272(.dina(n19821), .dinb(n16489), .dout(n20530));
  jor  g20273(.dina(n20530), .dinb(n20468), .dout(n20531));
  jxor g20274(.dina(n20531), .dinb(n20269), .dout(n20532));
  jnot g20275(.din(n20532), .dout(n20533));
  jor  g20276(.dina(n20533), .dinb(n20529), .dout(n20534));
  jand g20277(.dina(n20534), .dinb(n20528), .dout(n20535));
  jor  g20278(.dina(n20535), .dinb(n15260), .dout(n20536));
  jand g20279(.dina(n20535), .dinb(n15260), .dout(n20537));
  jxor g20280(.dina(n19828), .dinb(n15878), .dout(n20538));
  jor  g20281(.dina(n20538), .dinb(n20468), .dout(n20539));
  jxor g20282(.dina(n20539), .dinb(n19834), .dout(n20540));
  jor  g20283(.dina(n20540), .dinb(n20537), .dout(n20541));
  jand g20284(.dina(n20541), .dinb(n20536), .dout(n20542));
  jor  g20285(.dina(n20542), .dinb(n14674), .dout(n20543));
  jand g20286(.dina(n20542), .dinb(n14674), .dout(n20544));
  jxor g20287(.dina(n19836), .dinb(n15260), .dout(n20545));
  jor  g20288(.dina(n20545), .dinb(n20468), .dout(n20546));
  jxor g20289(.dina(n20546), .dinb(n20276), .dout(n20547));
  jnot g20290(.din(n20547), .dout(n20548));
  jor  g20291(.dina(n20548), .dinb(n20544), .dout(n20549));
  jand g20292(.dina(n20549), .dinb(n20543), .dout(n20550));
  jor  g20293(.dina(n20550), .dinb(n14078), .dout(n20551));
  jand g20294(.dina(n20550), .dinb(n14078), .dout(n20552));
  jxor g20295(.dina(n19843), .dinb(n14674), .dout(n20553));
  jor  g20296(.dina(n20553), .dinb(n20468), .dout(n20554));
  jxor g20297(.dina(n20554), .dinb(n19849), .dout(n20555));
  jor  g20298(.dina(n20555), .dinb(n20552), .dout(n20556));
  jand g20299(.dina(n20556), .dinb(n20551), .dout(n20557));
  jor  g20300(.dina(n20557), .dinb(n13515), .dout(n20558));
  jand g20301(.dina(n20557), .dinb(n13515), .dout(n20559));
  jxor g20302(.dina(n19851), .dinb(n14078), .dout(n20560));
  jor  g20303(.dina(n20560), .dinb(n20468), .dout(n20561));
  jxor g20304(.dina(n20561), .dinb(n20283), .dout(n20562));
  jnot g20305(.din(n20562), .dout(n20563));
  jor  g20306(.dina(n20563), .dinb(n20559), .dout(n20564));
  jand g20307(.dina(n20564), .dinb(n20558), .dout(n20565));
  jor  g20308(.dina(n20565), .dinb(n12947), .dout(n20566));
  jand g20309(.dina(n20565), .dinb(n12947), .dout(n20567));
  jxor g20310(.dina(n19858), .dinb(n13515), .dout(n20568));
  jor  g20311(.dina(n20568), .dinb(n20468), .dout(n20569));
  jxor g20312(.dina(n20569), .dinb(n19864), .dout(n20570));
  jor  g20313(.dina(n20570), .dinb(n20567), .dout(n20571));
  jand g20314(.dina(n20571), .dinb(n20566), .dout(n20572));
  jor  g20315(.dina(n20572), .dinb(n12410), .dout(n20573));
  jand g20316(.dina(n20572), .dinb(n12410), .dout(n20574));
  jxor g20317(.dina(n19866), .dinb(n12947), .dout(n20575));
  jor  g20318(.dina(n20575), .dinb(n20468), .dout(n20576));
  jxor g20319(.dina(n20576), .dinb(n20290), .dout(n20577));
  jnot g20320(.din(n20577), .dout(n20578));
  jor  g20321(.dina(n20578), .dinb(n20574), .dout(n20579));
  jand g20322(.dina(n20579), .dinb(n20573), .dout(n20580));
  jor  g20323(.dina(n20580), .dinb(n11858), .dout(n20581));
  jand g20324(.dina(n20580), .dinb(n11858), .dout(n20582));
  jxor g20325(.dina(n19873), .dinb(n12410), .dout(n20583));
  jor  g20326(.dina(n20583), .dinb(n20468), .dout(n20584));
  jxor g20327(.dina(n20584), .dinb(n19879), .dout(n20585));
  jor  g20328(.dina(n20585), .dinb(n20582), .dout(n20586));
  jand g20329(.dina(n20586), .dinb(n20581), .dout(n20587));
  jor  g20330(.dina(n20587), .dinb(n11347), .dout(n20588));
  jand g20331(.dina(n20587), .dinb(n11347), .dout(n20589));
  jxor g20332(.dina(n19881), .dinb(n11858), .dout(n20590));
  jor  g20333(.dina(n20590), .dinb(n20468), .dout(n20591));
  jxor g20334(.dina(n20591), .dinb(n20297), .dout(n20592));
  jnot g20335(.din(n20592), .dout(n20593));
  jor  g20336(.dina(n20593), .dinb(n20589), .dout(n20594));
  jand g20337(.dina(n20594), .dinb(n20588), .dout(n20595));
  jor  g20338(.dina(n20595), .dinb(n10824), .dout(n20596));
  jand g20339(.dina(n20595), .dinb(n10824), .dout(n20597));
  jxor g20340(.dina(n19888), .dinb(n11347), .dout(n20598));
  jor  g20341(.dina(n20598), .dinb(n20468), .dout(n20599));
  jxor g20342(.dina(n20599), .dinb(n19894), .dout(n20600));
  jor  g20343(.dina(n20600), .dinb(n20597), .dout(n20601));
  jand g20344(.dina(n20601), .dinb(n20596), .dout(n20602));
  jor  g20345(.dina(n20602), .dinb(n10328), .dout(n20603));
  jand g20346(.dina(n20602), .dinb(n10328), .dout(n20604));
  jxor g20347(.dina(n19896), .dinb(n10824), .dout(n20605));
  jor  g20348(.dina(n20605), .dinb(n20468), .dout(n20606));
  jxor g20349(.dina(n20606), .dinb(n19902), .dout(n20607));
  jor  g20350(.dina(n20607), .dinb(n20604), .dout(n20608));
  jand g20351(.dina(n20608), .dinb(n20603), .dout(n20609));
  jor  g20352(.dina(n20609), .dinb(n9832), .dout(n20610));
  jand g20353(.dina(n20609), .dinb(n9832), .dout(n20611));
  jxor g20354(.dina(n19904), .dinb(n10328), .dout(n20612));
  jor  g20355(.dina(n20612), .dinb(n20468), .dout(n20613));
  jxor g20356(.dina(n20613), .dinb(n20307), .dout(n20614));
  jnot g20357(.din(n20614), .dout(n20615));
  jor  g20358(.dina(n20615), .dinb(n20611), .dout(n20616));
  jand g20359(.dina(n20616), .dinb(n20610), .dout(n20617));
  jor  g20360(.dina(n20617), .dinb(n9369), .dout(n20618));
  jand g20361(.dina(n20617), .dinb(n9369), .dout(n20619));
  jxor g20362(.dina(n19911), .dinb(n9832), .dout(n20620));
  jor  g20363(.dina(n20620), .dinb(n20468), .dout(n20621));
  jxor g20364(.dina(n20621), .dinb(n20311), .dout(n20622));
  jnot g20365(.din(n20622), .dout(n20623));
  jor  g20366(.dina(n20623), .dinb(n20619), .dout(n20624));
  jand g20367(.dina(n20624), .dinb(n20618), .dout(n20625));
  jor  g20368(.dina(n20625), .dinb(n8890), .dout(n20626));
  jand g20369(.dina(n20625), .dinb(n8890), .dout(n20627));
  jxor g20370(.dina(n19918), .dinb(n9369), .dout(n20628));
  jor  g20371(.dina(n20628), .dinb(n20468), .dout(n20629));
  jxor g20372(.dina(n20629), .dinb(n19924), .dout(n20630));
  jor  g20373(.dina(n20630), .dinb(n20627), .dout(n20631));
  jand g20374(.dina(n20631), .dinb(n20626), .dout(n20632));
  jor  g20375(.dina(n20632), .dinb(n8449), .dout(n20633));
  jand g20376(.dina(n20632), .dinb(n8449), .dout(n20634));
  jxor g20377(.dina(n19926), .dinb(n8890), .dout(n20635));
  jor  g20378(.dina(n20635), .dinb(n20468), .dout(n20636));
  jxor g20379(.dina(n20636), .dinb(n20318), .dout(n20637));
  jnot g20380(.din(n20637), .dout(n20638));
  jor  g20381(.dina(n20638), .dinb(n20634), .dout(n20639));
  jand g20382(.dina(n20639), .dinb(n20633), .dout(n20640));
  jor  g20383(.dina(n20640), .dinb(n8003), .dout(n20641));
  jand g20384(.dina(n20640), .dinb(n8003), .dout(n20642));
  jxor g20385(.dina(n19933), .dinb(n8449), .dout(n20643));
  jor  g20386(.dina(n20643), .dinb(n20468), .dout(n20644));
  jxor g20387(.dina(n20644), .dinb(n19939), .dout(n20645));
  jor  g20388(.dina(n20645), .dinb(n20642), .dout(n20646));
  jand g20389(.dina(n20646), .dinb(n20641), .dout(n20647));
  jor  g20390(.dina(n20647), .dinb(n7581), .dout(n20648));
  jand g20391(.dina(n20647), .dinb(n7581), .dout(n20649));
  jxor g20392(.dina(n19941), .dinb(n8003), .dout(n20650));
  jor  g20393(.dina(n20650), .dinb(n20468), .dout(n20651));
  jxor g20394(.dina(n20651), .dinb(n20325), .dout(n20652));
  jnot g20395(.din(n20652), .dout(n20653));
  jor  g20396(.dina(n20653), .dinb(n20649), .dout(n20654));
  jand g20397(.dina(n20654), .dinb(n20648), .dout(n20655));
  jor  g20398(.dina(n20655), .dinb(n7154), .dout(n20656));
  jand g20399(.dina(n20655), .dinb(n7154), .dout(n20657));
  jxor g20400(.dina(n19948), .dinb(n7581), .dout(n20658));
  jor  g20401(.dina(n20658), .dinb(n20468), .dout(n20659));
  jxor g20402(.dina(n20659), .dinb(n19954), .dout(n20660));
  jor  g20403(.dina(n20660), .dinb(n20657), .dout(n20661));
  jand g20404(.dina(n20661), .dinb(n20656), .dout(n20662));
  jor  g20405(.dina(n20662), .dinb(n6758), .dout(n20663));
  jand g20406(.dina(n20662), .dinb(n6758), .dout(n20664));
  jxor g20407(.dina(n19956), .dinb(n7154), .dout(n20665));
  jor  g20408(.dina(n20665), .dinb(n20468), .dout(n20666));
  jxor g20409(.dina(n20666), .dinb(n19962), .dout(n20667));
  jor  g20410(.dina(n20667), .dinb(n20664), .dout(n20668));
  jand g20411(.dina(n20668), .dinb(n20663), .dout(n20669));
  jor  g20412(.dina(n20669), .dinb(n6357), .dout(n20670));
  jand g20413(.dina(n20669), .dinb(n6357), .dout(n20671));
  jxor g20414(.dina(n19964), .dinb(n6758), .dout(n20672));
  jor  g20415(.dina(n20672), .dinb(n20468), .dout(n20673));
  jxor g20416(.dina(n20673), .dinb(n19970), .dout(n20674));
  jor  g20417(.dina(n20674), .dinb(n20671), .dout(n20675));
  jand g20418(.dina(n20675), .dinb(n20670), .dout(n20676));
  jor  g20419(.dina(n20676), .dinb(n5989), .dout(n20677));
  jand g20420(.dina(n20676), .dinb(n5989), .dout(n20678));
  jxor g20421(.dina(n19972), .dinb(n6357), .dout(n20679));
  jor  g20422(.dina(n20679), .dinb(n20468), .dout(n20680));
  jxor g20423(.dina(n20680), .dinb(n20338), .dout(n20681));
  jnot g20424(.din(n20681), .dout(n20682));
  jor  g20425(.dina(n20682), .dinb(n20678), .dout(n20683));
  jand g20426(.dina(n20683), .dinb(n20677), .dout(n20684));
  jor  g20427(.dina(n20684), .dinb(n5606), .dout(n20685));
  jand g20428(.dina(n20684), .dinb(n5606), .dout(n20686));
  jxor g20429(.dina(n19979), .dinb(n5989), .dout(n20687));
  jor  g20430(.dina(n20687), .dinb(n20468), .dout(n20688));
  jxor g20431(.dina(n20688), .dinb(n19985), .dout(n20689));
  jor  g20432(.dina(n20689), .dinb(n20686), .dout(n20690));
  jand g20433(.dina(n20690), .dinb(n20685), .dout(n20691));
  jor  g20434(.dina(n20691), .dinb(n5259), .dout(n20692));
  jand g20435(.dina(n20691), .dinb(n5259), .dout(n20693));
  jxor g20436(.dina(n19987), .dinb(n5606), .dout(n20694));
  jor  g20437(.dina(n20694), .dinb(n20468), .dout(n20695));
  jxor g20438(.dina(n20695), .dinb(n20345), .dout(n20696));
  jnot g20439(.din(n20696), .dout(n20697));
  jor  g20440(.dina(n20697), .dinb(n20693), .dout(n20698));
  jand g20441(.dina(n20698), .dinb(n20692), .dout(n20699));
  jor  g20442(.dina(n20699), .dinb(n4902), .dout(n20700));
  jand g20443(.dina(n20699), .dinb(n4902), .dout(n20701));
  jxor g20444(.dina(n19994), .dinb(n5259), .dout(n20702));
  jor  g20445(.dina(n20702), .dinb(n20468), .dout(n20703));
  jxor g20446(.dina(n20703), .dinb(n20000), .dout(n20704));
  jor  g20447(.dina(n20704), .dinb(n20701), .dout(n20705));
  jand g20448(.dina(n20705), .dinb(n20700), .dout(n20706));
  jor  g20449(.dina(n20706), .dinb(n4582), .dout(n20707));
  jand g20450(.dina(n20706), .dinb(n4582), .dout(n20708));
  jxor g20451(.dina(n20002), .dinb(n4902), .dout(n20709));
  jor  g20452(.dina(n20709), .dinb(n20468), .dout(n20710));
  jxor g20453(.dina(n20710), .dinb(n20352), .dout(n20711));
  jnot g20454(.din(n20711), .dout(n20712));
  jor  g20455(.dina(n20712), .dinb(n20708), .dout(n20713));
  jand g20456(.dina(n20713), .dinb(n20707), .dout(n20714));
  jor  g20457(.dina(n20714), .dinb(n4249), .dout(n20715));
  jand g20458(.dina(n20714), .dinb(n4249), .dout(n20716));
  jxor g20459(.dina(n20009), .dinb(n4582), .dout(n20717));
  jor  g20460(.dina(n20717), .dinb(n20468), .dout(n20718));
  jxor g20461(.dina(n20718), .dinb(n20015), .dout(n20719));
  jor  g20462(.dina(n20719), .dinb(n20716), .dout(n20720));
  jand g20463(.dina(n20720), .dinb(n20715), .dout(n20721));
  jor  g20464(.dina(n20721), .dinb(n3955), .dout(n20722));
  jand g20465(.dina(n20721), .dinb(n3955), .dout(n20723));
  jxor g20466(.dina(n20017), .dinb(n4249), .dout(n20724));
  jor  g20467(.dina(n20724), .dinb(n20468), .dout(n20725));
  jxor g20468(.dina(n20725), .dinb(n20359), .dout(n20726));
  jnot g20469(.din(n20726), .dout(n20727));
  jor  g20470(.dina(n20727), .dinb(n20723), .dout(n20728));
  jand g20471(.dina(n20728), .dinb(n20722), .dout(n20729));
  jor  g20472(.dina(n20729), .dinb(n3642), .dout(n20730));
  jand g20473(.dina(n20729), .dinb(n3642), .dout(n20731));
  jxor g20474(.dina(n20024), .dinb(n3955), .dout(n20732));
  jor  g20475(.dina(n20732), .dinb(n20468), .dout(n20733));
  jxor g20476(.dina(n20733), .dinb(n20030), .dout(n20734));
  jor  g20477(.dina(n20734), .dinb(n20731), .dout(n20735));
  jand g20478(.dina(n20735), .dinb(n20730), .dout(n20736));
  jor  g20479(.dina(n20736), .dinb(n3368), .dout(n20737));
  jand g20480(.dina(n20736), .dinb(n3368), .dout(n20738));
  jxor g20481(.dina(n20032), .dinb(n3642), .dout(n20739));
  jor  g20482(.dina(n20739), .dinb(n20468), .dout(n20740));
  jxor g20483(.dina(n20740), .dinb(n20038), .dout(n20741));
  jor  g20484(.dina(n20741), .dinb(n20738), .dout(n20742));
  jand g20485(.dina(n20742), .dinb(n20737), .dout(n20743));
  jor  g20486(.dina(n20743), .dinb(n3089), .dout(n20744));
  jand g20487(.dina(n20743), .dinb(n3089), .dout(n20745));
  jxor g20488(.dina(n20040), .dinb(n3368), .dout(n20746));
  jor  g20489(.dina(n20746), .dinb(n20468), .dout(n20747));
  jxor g20490(.dina(n20747), .dinb(n20046), .dout(n20748));
  jor  g20491(.dina(n20748), .dinb(n20745), .dout(n20749));
  jand g20492(.dina(n20749), .dinb(n20744), .dout(n20750));
  jor  g20493(.dina(n20750), .dinb(n2833), .dout(n20751));
  jand g20494(.dina(n20750), .dinb(n2833), .dout(n20752));
  jxor g20495(.dina(n20048), .dinb(n3089), .dout(n20753));
  jor  g20496(.dina(n20753), .dinb(n20468), .dout(n20754));
  jxor g20497(.dina(n20754), .dinb(n20372), .dout(n20755));
  jnot g20498(.din(n20755), .dout(n20756));
  jor  g20499(.dina(n20756), .dinb(n20752), .dout(n20757));
  jand g20500(.dina(n20757), .dinb(n20751), .dout(n20758));
  jor  g20501(.dina(n20758), .dinb(n2572), .dout(n20759));
  jand g20502(.dina(n20758), .dinb(n2572), .dout(n20760));
  jxor g20503(.dina(n20055), .dinb(n2833), .dout(n20761));
  jor  g20504(.dina(n20761), .dinb(n20468), .dout(n20762));
  jxor g20505(.dina(n20762), .dinb(n20061), .dout(n20763));
  jor  g20506(.dina(n20763), .dinb(n20760), .dout(n20764));
  jand g20507(.dina(n20764), .dinb(n20759), .dout(n20765));
  jor  g20508(.dina(n20765), .dinb(n2345), .dout(n20766));
  jand g20509(.dina(n20765), .dinb(n2345), .dout(n20767));
  jxor g20510(.dina(n20063), .dinb(n2572), .dout(n20768));
  jor  g20511(.dina(n20768), .dinb(n20468), .dout(n20769));
  jxor g20512(.dina(n20769), .dinb(n20069), .dout(n20770));
  jor  g20513(.dina(n20770), .dinb(n20767), .dout(n20771));
  jand g20514(.dina(n20771), .dinb(n20766), .dout(n20772));
  jor  g20515(.dina(n20772), .dinb(n2108), .dout(n20773));
  jand g20516(.dina(n20772), .dinb(n2108), .dout(n20774));
  jxor g20517(.dina(n20071), .dinb(n2345), .dout(n20775));
  jor  g20518(.dina(n20775), .dinb(n20468), .dout(n20776));
  jxor g20519(.dina(n20776), .dinb(n20077), .dout(n20777));
  jor  g20520(.dina(n20777), .dinb(n20774), .dout(n20778));
  jand g20521(.dina(n20778), .dinb(n20773), .dout(n20779));
  jor  g20522(.dina(n20779), .dinb(n1912), .dout(n20780));
  jand g20523(.dina(n20779), .dinb(n1912), .dout(n20781));
  jxor g20524(.dina(n20079), .dinb(n2108), .dout(n20782));
  jor  g20525(.dina(n20782), .dinb(n20468), .dout(n20783));
  jxor g20526(.dina(n20783), .dinb(n20085), .dout(n20784));
  jor  g20527(.dina(n20784), .dinb(n20781), .dout(n20785));
  jand g20528(.dina(n20785), .dinb(n20780), .dout(n20786));
  jor  g20529(.dina(n20786), .dinb(n1699), .dout(n20787));
  jand g20530(.dina(n20786), .dinb(n1699), .dout(n20788));
  jxor g20531(.dina(n20087), .dinb(n1912), .dout(n20789));
  jor  g20532(.dina(n20789), .dinb(n20468), .dout(n20790));
  jxor g20533(.dina(n20790), .dinb(n20093), .dout(n20791));
  jor  g20534(.dina(n20791), .dinb(n20788), .dout(n20792));
  jand g20535(.dina(n20792), .dinb(n20787), .dout(n20793));
  jor  g20536(.dina(n20793), .dinb(n1516), .dout(n20794));
  jand g20537(.dina(n20793), .dinb(n1516), .dout(n20795));
  jxor g20538(.dina(n20095), .dinb(n1699), .dout(n20796));
  jor  g20539(.dina(n20796), .dinb(n20468), .dout(n20797));
  jxor g20540(.dina(n20797), .dinb(n20391), .dout(n20798));
  jnot g20541(.din(n20798), .dout(n20799));
  jor  g20542(.dina(n20799), .dinb(n20795), .dout(n20800));
  jand g20543(.dina(n20800), .dinb(n20794), .dout(n20801));
  jor  g20544(.dina(n20801), .dinb(n1332), .dout(n20802));
  jand g20545(.dina(n20801), .dinb(n1332), .dout(n20803));
  jxor g20546(.dina(n20102), .dinb(n1516), .dout(n20804));
  jor  g20547(.dina(n20804), .dinb(n20468), .dout(n20805));
  jxor g20548(.dina(n20805), .dinb(n20108), .dout(n20806));
  jor  g20549(.dina(n20806), .dinb(n20803), .dout(n20807));
  jand g20550(.dina(n20807), .dinb(n20802), .dout(n20808));
  jor  g20551(.dina(n20808), .dinb(n1173), .dout(n20809));
  jand g20552(.dina(n20808), .dinb(n1173), .dout(n20810));
  jxor g20553(.dina(n20110), .dinb(n1332), .dout(n20811));
  jor  g20554(.dina(n20811), .dinb(n20468), .dout(n20812));
  jxor g20555(.dina(n20812), .dinb(n20398), .dout(n20813));
  jnot g20556(.din(n20813), .dout(n20814));
  jor  g20557(.dina(n20814), .dinb(n20810), .dout(n20815));
  jand g20558(.dina(n20815), .dinb(n20809), .dout(n20816));
  jor  g20559(.dina(n20816), .dinb(n1008), .dout(n20817));
  jand g20560(.dina(n20816), .dinb(n1008), .dout(n20818));
  jxor g20561(.dina(n20117), .dinb(n1173), .dout(n20819));
  jor  g20562(.dina(n20819), .dinb(n20468), .dout(n20820));
  jxor g20563(.dina(n20820), .dinb(n20123), .dout(n20821));
  jor  g20564(.dina(n20821), .dinb(n20818), .dout(n20822));
  jand g20565(.dina(n20822), .dinb(n20817), .dout(n20823));
  jor  g20566(.dina(n20823), .dinb(n884), .dout(n20824));
  jand g20567(.dina(n20823), .dinb(n884), .dout(n20825));
  jxor g20568(.dina(n20125), .dinb(n1008), .dout(n20826));
  jor  g20569(.dina(n20826), .dinb(n20468), .dout(n20827));
  jxor g20570(.dina(n20827), .dinb(n20131), .dout(n20828));
  jor  g20571(.dina(n20828), .dinb(n20825), .dout(n20829));
  jand g20572(.dina(n20829), .dinb(n20824), .dout(n20830));
  jor  g20573(.dina(n20830), .dinb(n743), .dout(n20831));
  jand g20574(.dina(n20830), .dinb(n743), .dout(n20832));
  jxor g20575(.dina(n20133), .dinb(n884), .dout(n20833));
  jor  g20576(.dina(n20833), .dinb(n20468), .dout(n20834));
  jxor g20577(.dina(n20834), .dinb(n20408), .dout(n20835));
  jnot g20578(.din(n20835), .dout(n20836));
  jor  g20579(.dina(n20836), .dinb(n20832), .dout(n20837));
  jand g20580(.dina(n20837), .dinb(n20831), .dout(n20838));
  jor  g20581(.dina(n20838), .dinb(n635), .dout(n20839));
  jxor g20582(.dina(n20140), .dinb(n743), .dout(n20840));
  jor  g20583(.dina(n20840), .dinb(n20468), .dout(n20841));
  jxor g20584(.dina(n20841), .dinb(n20203), .dout(n20842));
  jnot g20585(.din(n20842), .dout(n20843));
  jand g20586(.dina(n20838), .dinb(n635), .dout(n20844));
  jor  g20587(.dina(n20844), .dinb(n20843), .dout(n20845));
  jand g20588(.dina(n20845), .dinb(n20839), .dout(n20846));
  jor  g20589(.dina(n20846), .dinb(n515), .dout(n20847));
  jand g20590(.dina(n20846), .dinb(n515), .dout(n20848));
  jxor g20591(.dina(n20147), .dinb(n635), .dout(n20849));
  jor  g20592(.dina(n20849), .dinb(n20468), .dout(n20850));
  jxor g20593(.dina(n20850), .dinb(n20153), .dout(n20851));
  jor  g20594(.dina(n20851), .dinb(n20848), .dout(n20852));
  jand g20595(.dina(n20852), .dinb(n20847), .dout(n20853));
  jor  g20596(.dina(n20853), .dinb(n443), .dout(n20854));
  jand g20597(.dina(n20853), .dinb(n443), .dout(n20855));
  jxor g20598(.dina(n20155), .dinb(n515), .dout(n20856));
  jor  g20599(.dina(n20856), .dinb(n20468), .dout(n20857));
  jxor g20600(.dina(n20857), .dinb(n20418), .dout(n20858));
  jnot g20601(.din(n20858), .dout(n20859));
  jor  g20602(.dina(n20859), .dinb(n20855), .dout(n20860));
  jand g20603(.dina(n20860), .dinb(n20854), .dout(n20861));
  jor  g20604(.dina(n20861), .dinb(n352), .dout(n20862));
  jand g20605(.dina(n20861), .dinb(n352), .dout(n20863));
  jxor g20606(.dina(n20162), .dinb(n443), .dout(n20864));
  jor  g20607(.dina(n20864), .dinb(n20468), .dout(n20865));
  jxor g20608(.dina(n20865), .dinb(n20168), .dout(n20866));
  jor  g20609(.dina(n20866), .dinb(n20863), .dout(n20867));
  jand g20610(.dina(n20867), .dinb(n20862), .dout(n20868));
  jor  g20611(.dina(n20868), .dinb(n294), .dout(n20869));
  jand g20612(.dina(n20868), .dinb(n294), .dout(n20870));
  jxor g20613(.dina(n20170), .dinb(n352), .dout(n20871));
  jor  g20614(.dina(n20871), .dinb(n20468), .dout(n20872));
  jxor g20615(.dina(n20872), .dinb(n20176), .dout(n20873));
  jor  g20616(.dina(n20873), .dinb(n20870), .dout(n20874));
  jand g20617(.dina(n20874), .dinb(n20869), .dout(n20875));
  jor  g20618(.dina(n20875), .dinb(n239), .dout(n20876));
  jand g20619(.dina(n20875), .dinb(n239), .dout(n20877));
  jxor g20620(.dina(n20178), .dinb(n294), .dout(n20878));
  jor  g20621(.dina(n20878), .dinb(n20468), .dout(n20879));
  jxor g20622(.dina(n20879), .dinb(n20428), .dout(n20880));
  jnot g20623(.din(n20880), .dout(n20881));
  jor  g20624(.dina(n20881), .dinb(n20877), .dout(n20882));
  jand g20625(.dina(n20882), .dinb(n20876), .dout(n20883));
  jor  g20626(.dina(n20883), .dinb(n221), .dout(n20884));
  jand g20627(.dina(n20883), .dinb(n221), .dout(n20885));
  jxor g20628(.dina(n20185), .dinb(n239), .dout(n20886));
  jor  g20629(.dina(n20886), .dinb(n20468), .dout(n20887));
  jxor g20630(.dina(n20887), .dinb(n20191), .dout(n20888));
  jor  g20631(.dina(n20888), .dinb(n20885), .dout(n20889));
  jand g20632(.dina(n20889), .dinb(n20884), .dout(n20890));
  jor  g20633(.dina(n20890), .dinb(n20472), .dout(n20891));
  jand g20634(.dina(asqrt[7] ), .dinb(n20459), .dout(n20892));
  jor  g20635(.dina(n20892), .dinb(n20446), .dout(n20893));
  jor  g20636(.dina(n20893), .dinb(n20891), .dout(n20894));
  jand g20637(.dina(n20894), .dinb(n218), .dout(n20895));
  jand g20638(.dina(n20468), .dinb(n19523), .dout(n20896));
  jand g20639(.dina(n20890), .dinb(n20472), .dout(n20897));
  jor  g20640(.dina(n20897), .dinb(n20896), .dout(n20898));
  jand g20641(.dina(n20468), .dinb(n20439), .dout(n20899));
  jand g20642(.dina(n20440), .dinb(asqrt[63] ), .dout(n20900));
  jand g20643(.dina(n20900), .dinb(n20464), .dout(n20901));
  jnot g20644(.din(n20901), .dout(n20902));
  jor  g20645(.dina(n20902), .dinb(n20899), .dout(n20903));
  jnot g20646(.din(n20903), .dout(n20904));
  jor  g20647(.dina(n20904), .dinb(n20898), .dout(n20905));
  jor  g20648(.dina(n20905), .dinb(n20895), .dout(asqrt[6] ));
  jnot g20649(.din(a[10] ), .dout(n20907));
  jnot g20650(.din(a[11] ), .dout(n20908));
  jand g20651(.dina(n20908), .dinb(n20907), .dout(n20909));
  jand g20652(.dina(n20909), .dinb(n20473), .dout(n20910));
  jand g20653(.dina(asqrt[6] ), .dinb(a[12] ), .dout(n20911));
  jor  g20654(.dina(n20911), .dinb(n20910), .dout(n20912));
  jand g20655(.dina(n20912), .dinb(asqrt[7] ), .dout(n20913));
  jor  g20656(.dina(n20912), .dinb(asqrt[7] ), .dout(n20914));
  jand g20657(.dina(asqrt[6] ), .dinb(n20473), .dout(n20915));
  jor  g20658(.dina(n20915), .dinb(n20474), .dout(n20916));
  jnot g20659(.din(n20475), .dout(n20917));
  jnot g20660(.din(n20884), .dout(n20918));
  jnot g20661(.din(n20876), .dout(n20919));
  jnot g20662(.din(n20869), .dout(n20920));
  jnot g20663(.din(n20862), .dout(n20921));
  jnot g20664(.din(n20854), .dout(n20922));
  jnot g20665(.din(n20847), .dout(n20923));
  jnot g20666(.din(n20839), .dout(n20924));
  jnot g20667(.din(n20831), .dout(n20925));
  jnot g20668(.din(n20824), .dout(n20926));
  jnot g20669(.din(n20817), .dout(n20927));
  jnot g20670(.din(n20809), .dout(n20928));
  jnot g20671(.din(n20802), .dout(n20929));
  jnot g20672(.din(n20794), .dout(n20930));
  jnot g20673(.din(n20787), .dout(n20931));
  jnot g20674(.din(n20780), .dout(n20932));
  jnot g20675(.din(n20773), .dout(n20933));
  jnot g20676(.din(n20766), .dout(n20934));
  jnot g20677(.din(n20759), .dout(n20935));
  jnot g20678(.din(n20751), .dout(n20936));
  jnot g20679(.din(n20744), .dout(n20937));
  jnot g20680(.din(n20737), .dout(n20938));
  jnot g20681(.din(n20730), .dout(n20939));
  jnot g20682(.din(n20722), .dout(n20940));
  jnot g20683(.din(n20715), .dout(n20941));
  jnot g20684(.din(n20707), .dout(n20942));
  jnot g20685(.din(n20700), .dout(n20943));
  jnot g20686(.din(n20692), .dout(n20944));
  jnot g20687(.din(n20685), .dout(n20945));
  jnot g20688(.din(n20677), .dout(n20946));
  jnot g20689(.din(n20670), .dout(n20947));
  jnot g20690(.din(n20663), .dout(n20948));
  jnot g20691(.din(n20656), .dout(n20949));
  jnot g20692(.din(n20648), .dout(n20950));
  jnot g20693(.din(n20641), .dout(n20951));
  jnot g20694(.din(n20633), .dout(n20952));
  jnot g20695(.din(n20626), .dout(n20953));
  jnot g20696(.din(n20618), .dout(n20954));
  jnot g20697(.din(n20610), .dout(n20955));
  jnot g20698(.din(n20603), .dout(n20956));
  jnot g20699(.din(n20596), .dout(n20957));
  jnot g20700(.din(n20588), .dout(n20958));
  jnot g20701(.din(n20581), .dout(n20959));
  jnot g20702(.din(n20573), .dout(n20960));
  jnot g20703(.din(n20566), .dout(n20961));
  jnot g20704(.din(n20558), .dout(n20962));
  jnot g20705(.din(n20551), .dout(n20963));
  jnot g20706(.din(n20543), .dout(n20964));
  jnot g20707(.din(n20536), .dout(n20965));
  jnot g20708(.din(n20528), .dout(n20966));
  jnot g20709(.din(n20521), .dout(n20967));
  jnot g20710(.din(n20514), .dout(n20968));
  jnot g20711(.din(n20507), .dout(n20969));
  jnot g20712(.din(n20499), .dout(n20970));
  jnot g20713(.din(n20488), .dout(n20971));
  jnot g20714(.din(n20480), .dout(n20972));
  jand g20715(.dina(asqrt[7] ), .dinb(a[14] ), .dout(n20973));
  jor  g20716(.dina(n20973), .dinb(n20476), .dout(n20974));
  jor  g20717(.dina(n20974), .dinb(asqrt[8] ), .dout(n20975));
  jand g20718(.dina(asqrt[7] ), .dinb(n19524), .dout(n20976));
  jor  g20719(.dina(n20976), .dinb(n19525), .dout(n20977));
  jand g20720(.dina(n20491), .dinb(n20977), .dout(n20978));
  jand g20721(.dina(n20978), .dinb(n20975), .dout(n20979));
  jor  g20722(.dina(n20979), .dinb(n20972), .dout(n20980));
  jor  g20723(.dina(n20980), .dinb(asqrt[9] ), .dout(n20981));
  jnot g20724(.din(n20496), .dout(n20982));
  jand g20725(.dina(n20982), .dinb(n20981), .dout(n20983));
  jor  g20726(.dina(n20983), .dinb(n20971), .dout(n20984));
  jor  g20727(.dina(n20984), .dinb(asqrt[10] ), .dout(n20985));
  jand g20728(.dina(n20503), .dinb(n20985), .dout(n20986));
  jor  g20729(.dina(n20986), .dinb(n20970), .dout(n20987));
  jor  g20730(.dina(n20987), .dinb(asqrt[11] ), .dout(n20988));
  jnot g20731(.din(n20511), .dout(n20989));
  jand g20732(.dina(n20989), .dinb(n20988), .dout(n20990));
  jor  g20733(.dina(n20990), .dinb(n20969), .dout(n20991));
  jor  g20734(.dina(n20991), .dinb(asqrt[12] ), .dout(n20992));
  jnot g20735(.din(n20518), .dout(n20993));
  jand g20736(.dina(n20993), .dinb(n20992), .dout(n20994));
  jor  g20737(.dina(n20994), .dinb(n20968), .dout(n20995));
  jor  g20738(.dina(n20995), .dinb(asqrt[13] ), .dout(n20996));
  jnot g20739(.din(n20525), .dout(n20997));
  jand g20740(.dina(n20997), .dinb(n20996), .dout(n20998));
  jor  g20741(.dina(n20998), .dinb(n20967), .dout(n20999));
  jor  g20742(.dina(n20999), .dinb(asqrt[14] ), .dout(n21000));
  jand g20743(.dina(n20532), .dinb(n21000), .dout(n21001));
  jor  g20744(.dina(n21001), .dinb(n20966), .dout(n21002));
  jor  g20745(.dina(n21002), .dinb(asqrt[15] ), .dout(n21003));
  jnot g20746(.din(n20540), .dout(n21004));
  jand g20747(.dina(n21004), .dinb(n21003), .dout(n21005));
  jor  g20748(.dina(n21005), .dinb(n20965), .dout(n21006));
  jor  g20749(.dina(n21006), .dinb(asqrt[16] ), .dout(n21007));
  jand g20750(.dina(n20547), .dinb(n21007), .dout(n21008));
  jor  g20751(.dina(n21008), .dinb(n20964), .dout(n21009));
  jor  g20752(.dina(n21009), .dinb(asqrt[17] ), .dout(n21010));
  jnot g20753(.din(n20555), .dout(n21011));
  jand g20754(.dina(n21011), .dinb(n21010), .dout(n21012));
  jor  g20755(.dina(n21012), .dinb(n20963), .dout(n21013));
  jor  g20756(.dina(n21013), .dinb(asqrt[18] ), .dout(n21014));
  jand g20757(.dina(n20562), .dinb(n21014), .dout(n21015));
  jor  g20758(.dina(n21015), .dinb(n20962), .dout(n21016));
  jor  g20759(.dina(n21016), .dinb(asqrt[19] ), .dout(n21017));
  jnot g20760(.din(n20570), .dout(n21018));
  jand g20761(.dina(n21018), .dinb(n21017), .dout(n21019));
  jor  g20762(.dina(n21019), .dinb(n20961), .dout(n21020));
  jor  g20763(.dina(n21020), .dinb(asqrt[20] ), .dout(n21021));
  jand g20764(.dina(n20577), .dinb(n21021), .dout(n21022));
  jor  g20765(.dina(n21022), .dinb(n20960), .dout(n21023));
  jor  g20766(.dina(n21023), .dinb(asqrt[21] ), .dout(n21024));
  jnot g20767(.din(n20585), .dout(n21025));
  jand g20768(.dina(n21025), .dinb(n21024), .dout(n21026));
  jor  g20769(.dina(n21026), .dinb(n20959), .dout(n21027));
  jor  g20770(.dina(n21027), .dinb(asqrt[22] ), .dout(n21028));
  jand g20771(.dina(n20592), .dinb(n21028), .dout(n21029));
  jor  g20772(.dina(n21029), .dinb(n20958), .dout(n21030));
  jor  g20773(.dina(n21030), .dinb(asqrt[23] ), .dout(n21031));
  jnot g20774(.din(n20600), .dout(n21032));
  jand g20775(.dina(n21032), .dinb(n21031), .dout(n21033));
  jor  g20776(.dina(n21033), .dinb(n20957), .dout(n21034));
  jor  g20777(.dina(n21034), .dinb(asqrt[24] ), .dout(n21035));
  jnot g20778(.din(n20607), .dout(n21036));
  jand g20779(.dina(n21036), .dinb(n21035), .dout(n21037));
  jor  g20780(.dina(n21037), .dinb(n20956), .dout(n21038));
  jor  g20781(.dina(n21038), .dinb(asqrt[25] ), .dout(n21039));
  jand g20782(.dina(n20614), .dinb(n21039), .dout(n21040));
  jor  g20783(.dina(n21040), .dinb(n20955), .dout(n21041));
  jor  g20784(.dina(n21041), .dinb(asqrt[26] ), .dout(n21042));
  jand g20785(.dina(n20622), .dinb(n21042), .dout(n21043));
  jor  g20786(.dina(n21043), .dinb(n20954), .dout(n21044));
  jor  g20787(.dina(n21044), .dinb(asqrt[27] ), .dout(n21045));
  jnot g20788(.din(n20630), .dout(n21046));
  jand g20789(.dina(n21046), .dinb(n21045), .dout(n21047));
  jor  g20790(.dina(n21047), .dinb(n20953), .dout(n21048));
  jor  g20791(.dina(n21048), .dinb(asqrt[28] ), .dout(n21049));
  jand g20792(.dina(n20637), .dinb(n21049), .dout(n21050));
  jor  g20793(.dina(n21050), .dinb(n20952), .dout(n21051));
  jor  g20794(.dina(n21051), .dinb(asqrt[29] ), .dout(n21052));
  jnot g20795(.din(n20645), .dout(n21053));
  jand g20796(.dina(n21053), .dinb(n21052), .dout(n21054));
  jor  g20797(.dina(n21054), .dinb(n20951), .dout(n21055));
  jor  g20798(.dina(n21055), .dinb(asqrt[30] ), .dout(n21056));
  jand g20799(.dina(n20652), .dinb(n21056), .dout(n21057));
  jor  g20800(.dina(n21057), .dinb(n20950), .dout(n21058));
  jor  g20801(.dina(n21058), .dinb(asqrt[31] ), .dout(n21059));
  jnot g20802(.din(n20660), .dout(n21060));
  jand g20803(.dina(n21060), .dinb(n21059), .dout(n21061));
  jor  g20804(.dina(n21061), .dinb(n20949), .dout(n21062));
  jor  g20805(.dina(n21062), .dinb(asqrt[32] ), .dout(n21063));
  jnot g20806(.din(n20667), .dout(n21064));
  jand g20807(.dina(n21064), .dinb(n21063), .dout(n21065));
  jor  g20808(.dina(n21065), .dinb(n20948), .dout(n21066));
  jor  g20809(.dina(n21066), .dinb(asqrt[33] ), .dout(n21067));
  jnot g20810(.din(n20674), .dout(n21068));
  jand g20811(.dina(n21068), .dinb(n21067), .dout(n21069));
  jor  g20812(.dina(n21069), .dinb(n20947), .dout(n21070));
  jor  g20813(.dina(n21070), .dinb(asqrt[34] ), .dout(n21071));
  jand g20814(.dina(n20681), .dinb(n21071), .dout(n21072));
  jor  g20815(.dina(n21072), .dinb(n20946), .dout(n21073));
  jor  g20816(.dina(n21073), .dinb(asqrt[35] ), .dout(n21074));
  jnot g20817(.din(n20689), .dout(n21075));
  jand g20818(.dina(n21075), .dinb(n21074), .dout(n21076));
  jor  g20819(.dina(n21076), .dinb(n20945), .dout(n21077));
  jor  g20820(.dina(n21077), .dinb(asqrt[36] ), .dout(n21078));
  jand g20821(.dina(n20696), .dinb(n21078), .dout(n21079));
  jor  g20822(.dina(n21079), .dinb(n20944), .dout(n21080));
  jor  g20823(.dina(n21080), .dinb(asqrt[37] ), .dout(n21081));
  jnot g20824(.din(n20704), .dout(n21082));
  jand g20825(.dina(n21082), .dinb(n21081), .dout(n21083));
  jor  g20826(.dina(n21083), .dinb(n20943), .dout(n21084));
  jor  g20827(.dina(n21084), .dinb(asqrt[38] ), .dout(n21085));
  jand g20828(.dina(n20711), .dinb(n21085), .dout(n21086));
  jor  g20829(.dina(n21086), .dinb(n20942), .dout(n21087));
  jor  g20830(.dina(n21087), .dinb(asqrt[39] ), .dout(n21088));
  jnot g20831(.din(n20719), .dout(n21089));
  jand g20832(.dina(n21089), .dinb(n21088), .dout(n21090));
  jor  g20833(.dina(n21090), .dinb(n20941), .dout(n21091));
  jor  g20834(.dina(n21091), .dinb(asqrt[40] ), .dout(n21092));
  jand g20835(.dina(n20726), .dinb(n21092), .dout(n21093));
  jor  g20836(.dina(n21093), .dinb(n20940), .dout(n21094));
  jor  g20837(.dina(n21094), .dinb(asqrt[41] ), .dout(n21095));
  jnot g20838(.din(n20734), .dout(n21096));
  jand g20839(.dina(n21096), .dinb(n21095), .dout(n21097));
  jor  g20840(.dina(n21097), .dinb(n20939), .dout(n21098));
  jor  g20841(.dina(n21098), .dinb(asqrt[42] ), .dout(n21099));
  jnot g20842(.din(n20741), .dout(n21100));
  jand g20843(.dina(n21100), .dinb(n21099), .dout(n21101));
  jor  g20844(.dina(n21101), .dinb(n20938), .dout(n21102));
  jor  g20845(.dina(n21102), .dinb(asqrt[43] ), .dout(n21103));
  jnot g20846(.din(n20748), .dout(n21104));
  jand g20847(.dina(n21104), .dinb(n21103), .dout(n21105));
  jor  g20848(.dina(n21105), .dinb(n20937), .dout(n21106));
  jor  g20849(.dina(n21106), .dinb(asqrt[44] ), .dout(n21107));
  jand g20850(.dina(n20755), .dinb(n21107), .dout(n21108));
  jor  g20851(.dina(n21108), .dinb(n20936), .dout(n21109));
  jor  g20852(.dina(n21109), .dinb(asqrt[45] ), .dout(n21110));
  jnot g20853(.din(n20763), .dout(n21111));
  jand g20854(.dina(n21111), .dinb(n21110), .dout(n21112));
  jor  g20855(.dina(n21112), .dinb(n20935), .dout(n21113));
  jor  g20856(.dina(n21113), .dinb(asqrt[46] ), .dout(n21114));
  jnot g20857(.din(n20770), .dout(n21115));
  jand g20858(.dina(n21115), .dinb(n21114), .dout(n21116));
  jor  g20859(.dina(n21116), .dinb(n20934), .dout(n21117));
  jor  g20860(.dina(n21117), .dinb(asqrt[47] ), .dout(n21118));
  jnot g20861(.din(n20777), .dout(n21119));
  jand g20862(.dina(n21119), .dinb(n21118), .dout(n21120));
  jor  g20863(.dina(n21120), .dinb(n20933), .dout(n21121));
  jor  g20864(.dina(n21121), .dinb(asqrt[48] ), .dout(n21122));
  jnot g20865(.din(n20784), .dout(n21123));
  jand g20866(.dina(n21123), .dinb(n21122), .dout(n21124));
  jor  g20867(.dina(n21124), .dinb(n20932), .dout(n21125));
  jor  g20868(.dina(n21125), .dinb(asqrt[49] ), .dout(n21126));
  jnot g20869(.din(n20791), .dout(n21127));
  jand g20870(.dina(n21127), .dinb(n21126), .dout(n21128));
  jor  g20871(.dina(n21128), .dinb(n20931), .dout(n21129));
  jor  g20872(.dina(n21129), .dinb(asqrt[50] ), .dout(n21130));
  jand g20873(.dina(n20798), .dinb(n21130), .dout(n21131));
  jor  g20874(.dina(n21131), .dinb(n20930), .dout(n21132));
  jor  g20875(.dina(n21132), .dinb(asqrt[51] ), .dout(n21133));
  jnot g20876(.din(n20806), .dout(n21134));
  jand g20877(.dina(n21134), .dinb(n21133), .dout(n21135));
  jor  g20878(.dina(n21135), .dinb(n20929), .dout(n21136));
  jor  g20879(.dina(n21136), .dinb(asqrt[52] ), .dout(n21137));
  jand g20880(.dina(n20813), .dinb(n21137), .dout(n21138));
  jor  g20881(.dina(n21138), .dinb(n20928), .dout(n21139));
  jor  g20882(.dina(n21139), .dinb(asqrt[53] ), .dout(n21140));
  jnot g20883(.din(n20821), .dout(n21141));
  jand g20884(.dina(n21141), .dinb(n21140), .dout(n21142));
  jor  g20885(.dina(n21142), .dinb(n20927), .dout(n21143));
  jor  g20886(.dina(n21143), .dinb(asqrt[54] ), .dout(n21144));
  jnot g20887(.din(n20828), .dout(n21145));
  jand g20888(.dina(n21145), .dinb(n21144), .dout(n21146));
  jor  g20889(.dina(n21146), .dinb(n20926), .dout(n21147));
  jor  g20890(.dina(n21147), .dinb(asqrt[55] ), .dout(n21148));
  jand g20891(.dina(n20835), .dinb(n21148), .dout(n21149));
  jor  g20892(.dina(n21149), .dinb(n20925), .dout(n21150));
  jor  g20893(.dina(n21150), .dinb(asqrt[56] ), .dout(n21151));
  jand g20894(.dina(n21151), .dinb(n20842), .dout(n21152));
  jor  g20895(.dina(n21152), .dinb(n20924), .dout(n21153));
  jor  g20896(.dina(n21153), .dinb(asqrt[57] ), .dout(n21154));
  jnot g20897(.din(n20851), .dout(n21155));
  jand g20898(.dina(n21155), .dinb(n21154), .dout(n21156));
  jor  g20899(.dina(n21156), .dinb(n20923), .dout(n21157));
  jor  g20900(.dina(n21157), .dinb(asqrt[58] ), .dout(n21158));
  jand g20901(.dina(n20858), .dinb(n21158), .dout(n21159));
  jor  g20902(.dina(n21159), .dinb(n20922), .dout(n21160));
  jor  g20903(.dina(n21160), .dinb(asqrt[59] ), .dout(n21161));
  jnot g20904(.din(n20866), .dout(n21162));
  jand g20905(.dina(n21162), .dinb(n21161), .dout(n21163));
  jor  g20906(.dina(n21163), .dinb(n20921), .dout(n21164));
  jor  g20907(.dina(n21164), .dinb(asqrt[60] ), .dout(n21165));
  jnot g20908(.din(n20873), .dout(n21166));
  jand g20909(.dina(n21166), .dinb(n21165), .dout(n21167));
  jor  g20910(.dina(n21167), .dinb(n20920), .dout(n21168));
  jor  g20911(.dina(n21168), .dinb(asqrt[61] ), .dout(n21169));
  jand g20912(.dina(n20880), .dinb(n21169), .dout(n21170));
  jor  g20913(.dina(n21170), .dinb(n20919), .dout(n21171));
  jor  g20914(.dina(n21171), .dinb(asqrt[62] ), .dout(n21172));
  jnot g20915(.din(n20888), .dout(n21173));
  jand g20916(.dina(n21173), .dinb(n21172), .dout(n21174));
  jor  g20917(.dina(n21174), .dinb(n20918), .dout(n21175));
  jand g20918(.dina(n21175), .dinb(n20471), .dout(n21176));
  jnot g20919(.din(n20893), .dout(n21177));
  jand g20920(.dina(n21177), .dinb(n21176), .dout(n21178));
  jor  g20921(.dina(n21178), .dinb(asqrt[63] ), .dout(n21179));
  jnot g20922(.din(n20896), .dout(n21180));
  jor  g20923(.dina(n21175), .dinb(n20471), .dout(n21181));
  jand g20924(.dina(n21181), .dinb(n21180), .dout(n21182));
  jand g20925(.dina(n20903), .dinb(n21182), .dout(n21183));
  jand g20926(.dina(n21183), .dinb(n21179), .dout(n21184));
  jor  g20927(.dina(n21184), .dinb(n20917), .dout(n21185));
  jand g20928(.dina(n21185), .dinb(n20916), .dout(n21186));
  jand g20929(.dina(n21186), .dinb(n20914), .dout(n21187));
  jor  g20930(.dina(n21187), .dinb(n20913), .dout(n21188));
  jand g20931(.dina(n21188), .dinb(asqrt[8] ), .dout(n21189));
  jor  g20932(.dina(n21188), .dinb(asqrt[8] ), .dout(n21190));
  jand g20933(.dina(asqrt[6] ), .dinb(n20475), .dout(n21191));
  jand g20934(.dina(n20902), .dinb(asqrt[7] ), .dout(n21192));
  jand g20935(.dina(n21192), .dinb(n21181), .dout(n21193));
  jand g20936(.dina(n21193), .dinb(n21179), .dout(n21194));
  jor  g20937(.dina(n21194), .dinb(n21191), .dout(n21195));
  jxor g20938(.dina(n21195), .dinb(a[14] ), .dout(n21196));
  jnot g20939(.din(n21196), .dout(n21197));
  jand g20940(.dina(n21197), .dinb(n21190), .dout(n21198));
  jor  g20941(.dina(n21198), .dinb(n21189), .dout(n21199));
  jand g20942(.dina(n21199), .dinb(asqrt[9] ), .dout(n21200));
  jor  g20943(.dina(n21199), .dinb(asqrt[9] ), .dout(n21201));
  jxor g20944(.dina(n20479), .dinb(n19791), .dout(n21202));
  jand g20945(.dina(n21202), .dinb(asqrt[6] ), .dout(n21203));
  jxor g20946(.dina(n21203), .dinb(n20978), .dout(n21204));
  jand g20947(.dina(n21204), .dinb(n21201), .dout(n21205));
  jor  g20948(.dina(n21205), .dinb(n21200), .dout(n21206));
  jand g20949(.dina(n21206), .dinb(asqrt[10] ), .dout(n21207));
  jor  g20950(.dina(n21206), .dinb(asqrt[10] ), .dout(n21208));
  jxor g20951(.dina(n20487), .dinb(n19096), .dout(n21209));
  jand g20952(.dina(n21209), .dinb(asqrt[6] ), .dout(n21210));
  jxor g20953(.dina(n21210), .dinb(n20496), .dout(n21211));
  jnot g20954(.din(n21211), .dout(n21212));
  jand g20955(.dina(n21212), .dinb(n21208), .dout(n21213));
  jor  g20956(.dina(n21213), .dinb(n21207), .dout(n21214));
  jand g20957(.dina(n21214), .dinb(asqrt[11] ), .dout(n21215));
  jor  g20958(.dina(n21214), .dinb(asqrt[11] ), .dout(n21216));
  jxor g20959(.dina(n20498), .dinb(n18442), .dout(n21217));
  jand g20960(.dina(n21217), .dinb(asqrt[6] ), .dout(n21218));
  jxor g20961(.dina(n21218), .dinb(n20503), .dout(n21219));
  jand g20962(.dina(n21219), .dinb(n21216), .dout(n21220));
  jor  g20963(.dina(n21220), .dinb(n21215), .dout(n21221));
  jand g20964(.dina(n21221), .dinb(asqrt[12] ), .dout(n21222));
  jor  g20965(.dina(n21221), .dinb(asqrt[12] ), .dout(n21223));
  jxor g20966(.dina(n20506), .dinb(n17769), .dout(n21224));
  jand g20967(.dina(n21224), .dinb(asqrt[6] ), .dout(n21225));
  jxor g20968(.dina(n21225), .dinb(n20511), .dout(n21226));
  jnot g20969(.din(n21226), .dout(n21227));
  jand g20970(.dina(n21227), .dinb(n21223), .dout(n21228));
  jor  g20971(.dina(n21228), .dinb(n21222), .dout(n21229));
  jand g20972(.dina(n21229), .dinb(asqrt[13] ), .dout(n21230));
  jor  g20973(.dina(n21229), .dinb(asqrt[13] ), .dout(n21231));
  jxor g20974(.dina(n20513), .dinb(n17134), .dout(n21232));
  jand g20975(.dina(n21232), .dinb(asqrt[6] ), .dout(n21233));
  jxor g20976(.dina(n21233), .dinb(n20518), .dout(n21234));
  jnot g20977(.din(n21234), .dout(n21235));
  jand g20978(.dina(n21235), .dinb(n21231), .dout(n21236));
  jor  g20979(.dina(n21236), .dinb(n21230), .dout(n21237));
  jand g20980(.dina(n21237), .dinb(asqrt[14] ), .dout(n21238));
  jor  g20981(.dina(n21237), .dinb(asqrt[14] ), .dout(n21239));
  jxor g20982(.dina(n20520), .dinb(n16489), .dout(n21240));
  jand g20983(.dina(n21240), .dinb(asqrt[6] ), .dout(n21241));
  jxor g20984(.dina(n21241), .dinb(n20525), .dout(n21242));
  jnot g20985(.din(n21242), .dout(n21243));
  jand g20986(.dina(n21243), .dinb(n21239), .dout(n21244));
  jor  g20987(.dina(n21244), .dinb(n21238), .dout(n21245));
  jand g20988(.dina(n21245), .dinb(asqrt[15] ), .dout(n21246));
  jor  g20989(.dina(n21245), .dinb(asqrt[15] ), .dout(n21247));
  jxor g20990(.dina(n20527), .dinb(n15878), .dout(n21248));
  jand g20991(.dina(n21248), .dinb(asqrt[6] ), .dout(n21249));
  jxor g20992(.dina(n21249), .dinb(n20532), .dout(n21250));
  jand g20993(.dina(n21250), .dinb(n21247), .dout(n21251));
  jor  g20994(.dina(n21251), .dinb(n21246), .dout(n21252));
  jand g20995(.dina(n21252), .dinb(asqrt[16] ), .dout(n21253));
  jor  g20996(.dina(n21252), .dinb(asqrt[16] ), .dout(n21254));
  jxor g20997(.dina(n20535), .dinb(n15260), .dout(n21255));
  jand g20998(.dina(n21255), .dinb(asqrt[6] ), .dout(n21256));
  jxor g20999(.dina(n21256), .dinb(n20540), .dout(n21257));
  jnot g21000(.din(n21257), .dout(n21258));
  jand g21001(.dina(n21258), .dinb(n21254), .dout(n21259));
  jor  g21002(.dina(n21259), .dinb(n21253), .dout(n21260));
  jand g21003(.dina(n21260), .dinb(asqrt[17] ), .dout(n21261));
  jor  g21004(.dina(n21260), .dinb(asqrt[17] ), .dout(n21262));
  jxor g21005(.dina(n20542), .dinb(n14674), .dout(n21263));
  jand g21006(.dina(n21263), .dinb(asqrt[6] ), .dout(n21264));
  jxor g21007(.dina(n21264), .dinb(n20548), .dout(n21265));
  jnot g21008(.din(n21265), .dout(n21266));
  jand g21009(.dina(n21266), .dinb(n21262), .dout(n21267));
  jor  g21010(.dina(n21267), .dinb(n21261), .dout(n21268));
  jand g21011(.dina(n21268), .dinb(asqrt[18] ), .dout(n21269));
  jor  g21012(.dina(n21268), .dinb(asqrt[18] ), .dout(n21270));
  jxor g21013(.dina(n20550), .dinb(n14078), .dout(n21271));
  jand g21014(.dina(n21271), .dinb(asqrt[6] ), .dout(n21272));
  jxor g21015(.dina(n21272), .dinb(n20555), .dout(n21273));
  jnot g21016(.din(n21273), .dout(n21274));
  jand g21017(.dina(n21274), .dinb(n21270), .dout(n21275));
  jor  g21018(.dina(n21275), .dinb(n21269), .dout(n21276));
  jand g21019(.dina(n21276), .dinb(asqrt[19] ), .dout(n21277));
  jor  g21020(.dina(n21276), .dinb(asqrt[19] ), .dout(n21278));
  jxor g21021(.dina(n20557), .dinb(n13515), .dout(n21279));
  jand g21022(.dina(n21279), .dinb(asqrt[6] ), .dout(n21280));
  jxor g21023(.dina(n21280), .dinb(n20562), .dout(n21281));
  jand g21024(.dina(n21281), .dinb(n21278), .dout(n21282));
  jor  g21025(.dina(n21282), .dinb(n21277), .dout(n21283));
  jand g21026(.dina(n21283), .dinb(asqrt[20] ), .dout(n21284));
  jor  g21027(.dina(n21283), .dinb(asqrt[20] ), .dout(n21285));
  jxor g21028(.dina(n20565), .dinb(n12947), .dout(n21286));
  jand g21029(.dina(n21286), .dinb(asqrt[6] ), .dout(n21287));
  jxor g21030(.dina(n21287), .dinb(n20570), .dout(n21288));
  jnot g21031(.din(n21288), .dout(n21289));
  jand g21032(.dina(n21289), .dinb(n21285), .dout(n21290));
  jor  g21033(.dina(n21290), .dinb(n21284), .dout(n21291));
  jand g21034(.dina(n21291), .dinb(asqrt[21] ), .dout(n21292));
  jor  g21035(.dina(n21291), .dinb(asqrt[21] ), .dout(n21293));
  jxor g21036(.dina(n20572), .dinb(n12410), .dout(n21294));
  jand g21037(.dina(n21294), .dinb(asqrt[6] ), .dout(n21295));
  jxor g21038(.dina(n21295), .dinb(n20577), .dout(n21296));
  jand g21039(.dina(n21296), .dinb(n21293), .dout(n21297));
  jor  g21040(.dina(n21297), .dinb(n21292), .dout(n21298));
  jand g21041(.dina(n21298), .dinb(asqrt[22] ), .dout(n21299));
  jor  g21042(.dina(n21298), .dinb(asqrt[22] ), .dout(n21300));
  jxor g21043(.dina(n20580), .dinb(n11858), .dout(n21301));
  jand g21044(.dina(n21301), .dinb(asqrt[6] ), .dout(n21302));
  jxor g21045(.dina(n21302), .dinb(n20585), .dout(n21303));
  jnot g21046(.din(n21303), .dout(n21304));
  jand g21047(.dina(n21304), .dinb(n21300), .dout(n21305));
  jor  g21048(.dina(n21305), .dinb(n21299), .dout(n21306));
  jand g21049(.dina(n21306), .dinb(asqrt[23] ), .dout(n21307));
  jor  g21050(.dina(n21306), .dinb(asqrt[23] ), .dout(n21308));
  jxor g21051(.dina(n20587), .dinb(n11347), .dout(n21309));
  jand g21052(.dina(n21309), .dinb(asqrt[6] ), .dout(n21310));
  jxor g21053(.dina(n21310), .dinb(n20592), .dout(n21311));
  jand g21054(.dina(n21311), .dinb(n21308), .dout(n21312));
  jor  g21055(.dina(n21312), .dinb(n21307), .dout(n21313));
  jand g21056(.dina(n21313), .dinb(asqrt[24] ), .dout(n21314));
  jor  g21057(.dina(n21313), .dinb(asqrt[24] ), .dout(n21315));
  jxor g21058(.dina(n20595), .dinb(n10824), .dout(n21316));
  jand g21059(.dina(n21316), .dinb(asqrt[6] ), .dout(n21317));
  jxor g21060(.dina(n21317), .dinb(n20600), .dout(n21318));
  jnot g21061(.din(n21318), .dout(n21319));
  jand g21062(.dina(n21319), .dinb(n21315), .dout(n21320));
  jor  g21063(.dina(n21320), .dinb(n21314), .dout(n21321));
  jand g21064(.dina(n21321), .dinb(asqrt[25] ), .dout(n21322));
  jor  g21065(.dina(n21321), .dinb(asqrt[25] ), .dout(n21323));
  jxor g21066(.dina(n20602), .dinb(n10328), .dout(n21324));
  jand g21067(.dina(n21324), .dinb(asqrt[6] ), .dout(n21325));
  jxor g21068(.dina(n21325), .dinb(n20607), .dout(n21326));
  jnot g21069(.din(n21326), .dout(n21327));
  jand g21070(.dina(n21327), .dinb(n21323), .dout(n21328));
  jor  g21071(.dina(n21328), .dinb(n21322), .dout(n21329));
  jand g21072(.dina(n21329), .dinb(asqrt[26] ), .dout(n21330));
  jor  g21073(.dina(n21329), .dinb(asqrt[26] ), .dout(n21331));
  jxor g21074(.dina(n20609), .dinb(n9832), .dout(n21332));
  jand g21075(.dina(n21332), .dinb(asqrt[6] ), .dout(n21333));
  jxor g21076(.dina(n21333), .dinb(n20614), .dout(n21334));
  jand g21077(.dina(n21334), .dinb(n21331), .dout(n21335));
  jor  g21078(.dina(n21335), .dinb(n21330), .dout(n21336));
  jand g21079(.dina(n21336), .dinb(asqrt[27] ), .dout(n21337));
  jor  g21080(.dina(n21336), .dinb(asqrt[27] ), .dout(n21338));
  jxor g21081(.dina(n20617), .dinb(n9369), .dout(n21339));
  jand g21082(.dina(n21339), .dinb(asqrt[6] ), .dout(n21340));
  jxor g21083(.dina(n21340), .dinb(n20622), .dout(n21341));
  jand g21084(.dina(n21341), .dinb(n21338), .dout(n21342));
  jor  g21085(.dina(n21342), .dinb(n21337), .dout(n21343));
  jand g21086(.dina(n21343), .dinb(asqrt[28] ), .dout(n21344));
  jor  g21087(.dina(n21343), .dinb(asqrt[28] ), .dout(n21345));
  jxor g21088(.dina(n20625), .dinb(n8890), .dout(n21346));
  jand g21089(.dina(n21346), .dinb(asqrt[6] ), .dout(n21347));
  jxor g21090(.dina(n21347), .dinb(n20630), .dout(n21348));
  jnot g21091(.din(n21348), .dout(n21349));
  jand g21092(.dina(n21349), .dinb(n21345), .dout(n21350));
  jor  g21093(.dina(n21350), .dinb(n21344), .dout(n21351));
  jand g21094(.dina(n21351), .dinb(asqrt[29] ), .dout(n21352));
  jor  g21095(.dina(n21351), .dinb(asqrt[29] ), .dout(n21353));
  jxor g21096(.dina(n20632), .dinb(n8449), .dout(n21354));
  jand g21097(.dina(n21354), .dinb(asqrt[6] ), .dout(n21355));
  jxor g21098(.dina(n21355), .dinb(n20637), .dout(n21356));
  jand g21099(.dina(n21356), .dinb(n21353), .dout(n21357));
  jor  g21100(.dina(n21357), .dinb(n21352), .dout(n21358));
  jand g21101(.dina(n21358), .dinb(asqrt[30] ), .dout(n21359));
  jor  g21102(.dina(n21358), .dinb(asqrt[30] ), .dout(n21360));
  jxor g21103(.dina(n20640), .dinb(n8003), .dout(n21361));
  jand g21104(.dina(n21361), .dinb(asqrt[6] ), .dout(n21362));
  jxor g21105(.dina(n21362), .dinb(n20645), .dout(n21363));
  jnot g21106(.din(n21363), .dout(n21364));
  jand g21107(.dina(n21364), .dinb(n21360), .dout(n21365));
  jor  g21108(.dina(n21365), .dinb(n21359), .dout(n21366));
  jand g21109(.dina(n21366), .dinb(asqrt[31] ), .dout(n21367));
  jor  g21110(.dina(n21366), .dinb(asqrt[31] ), .dout(n21368));
  jxor g21111(.dina(n20647), .dinb(n7581), .dout(n21369));
  jand g21112(.dina(n21369), .dinb(asqrt[6] ), .dout(n21370));
  jxor g21113(.dina(n21370), .dinb(n20652), .dout(n21371));
  jand g21114(.dina(n21371), .dinb(n21368), .dout(n21372));
  jor  g21115(.dina(n21372), .dinb(n21367), .dout(n21373));
  jand g21116(.dina(n21373), .dinb(asqrt[32] ), .dout(n21374));
  jor  g21117(.dina(n21373), .dinb(asqrt[32] ), .dout(n21375));
  jxor g21118(.dina(n20655), .dinb(n7154), .dout(n21376));
  jand g21119(.dina(n21376), .dinb(asqrt[6] ), .dout(n21377));
  jxor g21120(.dina(n21377), .dinb(n20660), .dout(n21378));
  jnot g21121(.din(n21378), .dout(n21379));
  jand g21122(.dina(n21379), .dinb(n21375), .dout(n21380));
  jor  g21123(.dina(n21380), .dinb(n21374), .dout(n21381));
  jand g21124(.dina(n21381), .dinb(asqrt[33] ), .dout(n21382));
  jor  g21125(.dina(n21381), .dinb(asqrt[33] ), .dout(n21383));
  jxor g21126(.dina(n20662), .dinb(n6758), .dout(n21384));
  jand g21127(.dina(n21384), .dinb(asqrt[6] ), .dout(n21385));
  jxor g21128(.dina(n21385), .dinb(n20667), .dout(n21386));
  jnot g21129(.din(n21386), .dout(n21387));
  jand g21130(.dina(n21387), .dinb(n21383), .dout(n21388));
  jor  g21131(.dina(n21388), .dinb(n21382), .dout(n21389));
  jand g21132(.dina(n21389), .dinb(asqrt[34] ), .dout(n21390));
  jor  g21133(.dina(n21389), .dinb(asqrt[34] ), .dout(n21391));
  jxor g21134(.dina(n20669), .dinb(n6357), .dout(n21392));
  jand g21135(.dina(n21392), .dinb(asqrt[6] ), .dout(n21393));
  jxor g21136(.dina(n21393), .dinb(n20674), .dout(n21394));
  jnot g21137(.din(n21394), .dout(n21395));
  jand g21138(.dina(n21395), .dinb(n21391), .dout(n21396));
  jor  g21139(.dina(n21396), .dinb(n21390), .dout(n21397));
  jand g21140(.dina(n21397), .dinb(asqrt[35] ), .dout(n21398));
  jor  g21141(.dina(n21397), .dinb(asqrt[35] ), .dout(n21399));
  jxor g21142(.dina(n20676), .dinb(n5989), .dout(n21400));
  jand g21143(.dina(n21400), .dinb(asqrt[6] ), .dout(n21401));
  jxor g21144(.dina(n21401), .dinb(n20681), .dout(n21402));
  jand g21145(.dina(n21402), .dinb(n21399), .dout(n21403));
  jor  g21146(.dina(n21403), .dinb(n21398), .dout(n21404));
  jand g21147(.dina(n21404), .dinb(asqrt[36] ), .dout(n21405));
  jor  g21148(.dina(n21404), .dinb(asqrt[36] ), .dout(n21406));
  jxor g21149(.dina(n20684), .dinb(n5606), .dout(n21407));
  jand g21150(.dina(n21407), .dinb(asqrt[6] ), .dout(n21408));
  jxor g21151(.dina(n21408), .dinb(n20689), .dout(n21409));
  jnot g21152(.din(n21409), .dout(n21410));
  jand g21153(.dina(n21410), .dinb(n21406), .dout(n21411));
  jor  g21154(.dina(n21411), .dinb(n21405), .dout(n21412));
  jand g21155(.dina(n21412), .dinb(asqrt[37] ), .dout(n21413));
  jor  g21156(.dina(n21412), .dinb(asqrt[37] ), .dout(n21414));
  jxor g21157(.dina(n20691), .dinb(n5259), .dout(n21415));
  jand g21158(.dina(n21415), .dinb(asqrt[6] ), .dout(n21416));
  jxor g21159(.dina(n21416), .dinb(n20696), .dout(n21417));
  jand g21160(.dina(n21417), .dinb(n21414), .dout(n21418));
  jor  g21161(.dina(n21418), .dinb(n21413), .dout(n21419));
  jand g21162(.dina(n21419), .dinb(asqrt[38] ), .dout(n21420));
  jor  g21163(.dina(n21419), .dinb(asqrt[38] ), .dout(n21421));
  jxor g21164(.dina(n20699), .dinb(n4902), .dout(n21422));
  jand g21165(.dina(n21422), .dinb(asqrt[6] ), .dout(n21423));
  jxor g21166(.dina(n21423), .dinb(n20704), .dout(n21424));
  jnot g21167(.din(n21424), .dout(n21425));
  jand g21168(.dina(n21425), .dinb(n21421), .dout(n21426));
  jor  g21169(.dina(n21426), .dinb(n21420), .dout(n21427));
  jand g21170(.dina(n21427), .dinb(asqrt[39] ), .dout(n21428));
  jor  g21171(.dina(n21427), .dinb(asqrt[39] ), .dout(n21429));
  jxor g21172(.dina(n20706), .dinb(n4582), .dout(n21430));
  jand g21173(.dina(n21430), .dinb(asqrt[6] ), .dout(n21431));
  jxor g21174(.dina(n21431), .dinb(n20711), .dout(n21432));
  jand g21175(.dina(n21432), .dinb(n21429), .dout(n21433));
  jor  g21176(.dina(n21433), .dinb(n21428), .dout(n21434));
  jand g21177(.dina(n21434), .dinb(asqrt[40] ), .dout(n21435));
  jor  g21178(.dina(n21434), .dinb(asqrt[40] ), .dout(n21436));
  jxor g21179(.dina(n20714), .dinb(n4249), .dout(n21437));
  jand g21180(.dina(n21437), .dinb(asqrt[6] ), .dout(n21438));
  jxor g21181(.dina(n21438), .dinb(n20719), .dout(n21439));
  jnot g21182(.din(n21439), .dout(n21440));
  jand g21183(.dina(n21440), .dinb(n21436), .dout(n21441));
  jor  g21184(.dina(n21441), .dinb(n21435), .dout(n21442));
  jand g21185(.dina(n21442), .dinb(asqrt[41] ), .dout(n21443));
  jor  g21186(.dina(n21442), .dinb(asqrt[41] ), .dout(n21444));
  jxor g21187(.dina(n20721), .dinb(n3955), .dout(n21445));
  jand g21188(.dina(n21445), .dinb(asqrt[6] ), .dout(n21446));
  jxor g21189(.dina(n21446), .dinb(n20726), .dout(n21447));
  jand g21190(.dina(n21447), .dinb(n21444), .dout(n21448));
  jor  g21191(.dina(n21448), .dinb(n21443), .dout(n21449));
  jand g21192(.dina(n21449), .dinb(asqrt[42] ), .dout(n21450));
  jor  g21193(.dina(n21449), .dinb(asqrt[42] ), .dout(n21451));
  jxor g21194(.dina(n20729), .dinb(n3642), .dout(n21452));
  jand g21195(.dina(n21452), .dinb(asqrt[6] ), .dout(n21453));
  jxor g21196(.dina(n21453), .dinb(n20734), .dout(n21454));
  jnot g21197(.din(n21454), .dout(n21455));
  jand g21198(.dina(n21455), .dinb(n21451), .dout(n21456));
  jor  g21199(.dina(n21456), .dinb(n21450), .dout(n21457));
  jand g21200(.dina(n21457), .dinb(asqrt[43] ), .dout(n21458));
  jor  g21201(.dina(n21457), .dinb(asqrt[43] ), .dout(n21459));
  jxor g21202(.dina(n20736), .dinb(n3368), .dout(n21460));
  jand g21203(.dina(n21460), .dinb(asqrt[6] ), .dout(n21461));
  jxor g21204(.dina(n21461), .dinb(n20741), .dout(n21462));
  jnot g21205(.din(n21462), .dout(n21463));
  jand g21206(.dina(n21463), .dinb(n21459), .dout(n21464));
  jor  g21207(.dina(n21464), .dinb(n21458), .dout(n21465));
  jand g21208(.dina(n21465), .dinb(asqrt[44] ), .dout(n21466));
  jor  g21209(.dina(n21465), .dinb(asqrt[44] ), .dout(n21467));
  jxor g21210(.dina(n20743), .dinb(n3089), .dout(n21468));
  jand g21211(.dina(n21468), .dinb(asqrt[6] ), .dout(n21469));
  jxor g21212(.dina(n21469), .dinb(n20748), .dout(n21470));
  jnot g21213(.din(n21470), .dout(n21471));
  jand g21214(.dina(n21471), .dinb(n21467), .dout(n21472));
  jor  g21215(.dina(n21472), .dinb(n21466), .dout(n21473));
  jand g21216(.dina(n21473), .dinb(asqrt[45] ), .dout(n21474));
  jor  g21217(.dina(n21473), .dinb(asqrt[45] ), .dout(n21475));
  jxor g21218(.dina(n20750), .dinb(n2833), .dout(n21476));
  jand g21219(.dina(n21476), .dinb(asqrt[6] ), .dout(n21477));
  jxor g21220(.dina(n21477), .dinb(n20755), .dout(n21478));
  jand g21221(.dina(n21478), .dinb(n21475), .dout(n21479));
  jor  g21222(.dina(n21479), .dinb(n21474), .dout(n21480));
  jand g21223(.dina(n21480), .dinb(asqrt[46] ), .dout(n21481));
  jor  g21224(.dina(n21480), .dinb(asqrt[46] ), .dout(n21482));
  jxor g21225(.dina(n20758), .dinb(n2572), .dout(n21483));
  jand g21226(.dina(n21483), .dinb(asqrt[6] ), .dout(n21484));
  jxor g21227(.dina(n21484), .dinb(n20763), .dout(n21485));
  jnot g21228(.din(n21485), .dout(n21486));
  jand g21229(.dina(n21486), .dinb(n21482), .dout(n21487));
  jor  g21230(.dina(n21487), .dinb(n21481), .dout(n21488));
  jand g21231(.dina(n21488), .dinb(asqrt[47] ), .dout(n21489));
  jor  g21232(.dina(n21488), .dinb(asqrt[47] ), .dout(n21490));
  jxor g21233(.dina(n20765), .dinb(n2345), .dout(n21491));
  jand g21234(.dina(n21491), .dinb(asqrt[6] ), .dout(n21492));
  jxor g21235(.dina(n21492), .dinb(n20770), .dout(n21493));
  jnot g21236(.din(n21493), .dout(n21494));
  jand g21237(.dina(n21494), .dinb(n21490), .dout(n21495));
  jor  g21238(.dina(n21495), .dinb(n21489), .dout(n21496));
  jand g21239(.dina(n21496), .dinb(asqrt[48] ), .dout(n21497));
  jor  g21240(.dina(n21496), .dinb(asqrt[48] ), .dout(n21498));
  jxor g21241(.dina(n20772), .dinb(n2108), .dout(n21499));
  jand g21242(.dina(n21499), .dinb(asqrt[6] ), .dout(n21500));
  jxor g21243(.dina(n21500), .dinb(n20777), .dout(n21501));
  jnot g21244(.din(n21501), .dout(n21502));
  jand g21245(.dina(n21502), .dinb(n21498), .dout(n21503));
  jor  g21246(.dina(n21503), .dinb(n21497), .dout(n21504));
  jand g21247(.dina(n21504), .dinb(asqrt[49] ), .dout(n21505));
  jor  g21248(.dina(n21504), .dinb(asqrt[49] ), .dout(n21506));
  jxor g21249(.dina(n20779), .dinb(n1912), .dout(n21507));
  jand g21250(.dina(n21507), .dinb(asqrt[6] ), .dout(n21508));
  jxor g21251(.dina(n21508), .dinb(n20784), .dout(n21509));
  jnot g21252(.din(n21509), .dout(n21510));
  jand g21253(.dina(n21510), .dinb(n21506), .dout(n21511));
  jor  g21254(.dina(n21511), .dinb(n21505), .dout(n21512));
  jand g21255(.dina(n21512), .dinb(asqrt[50] ), .dout(n21513));
  jor  g21256(.dina(n21512), .dinb(asqrt[50] ), .dout(n21514));
  jxor g21257(.dina(n20786), .dinb(n1699), .dout(n21515));
  jand g21258(.dina(n21515), .dinb(asqrt[6] ), .dout(n21516));
  jxor g21259(.dina(n21516), .dinb(n20791), .dout(n21517));
  jnot g21260(.din(n21517), .dout(n21518));
  jand g21261(.dina(n21518), .dinb(n21514), .dout(n21519));
  jor  g21262(.dina(n21519), .dinb(n21513), .dout(n21520));
  jand g21263(.dina(n21520), .dinb(asqrt[51] ), .dout(n21521));
  jor  g21264(.dina(n21520), .dinb(asqrt[51] ), .dout(n21522));
  jxor g21265(.dina(n20793), .dinb(n1516), .dout(n21523));
  jand g21266(.dina(n21523), .dinb(asqrt[6] ), .dout(n21524));
  jxor g21267(.dina(n21524), .dinb(n20798), .dout(n21525));
  jand g21268(.dina(n21525), .dinb(n21522), .dout(n21526));
  jor  g21269(.dina(n21526), .dinb(n21521), .dout(n21527));
  jand g21270(.dina(n21527), .dinb(asqrt[52] ), .dout(n21528));
  jor  g21271(.dina(n21527), .dinb(asqrt[52] ), .dout(n21529));
  jxor g21272(.dina(n20801), .dinb(n1332), .dout(n21530));
  jand g21273(.dina(n21530), .dinb(asqrt[6] ), .dout(n21531));
  jxor g21274(.dina(n21531), .dinb(n20806), .dout(n21532));
  jnot g21275(.din(n21532), .dout(n21533));
  jand g21276(.dina(n21533), .dinb(n21529), .dout(n21534));
  jor  g21277(.dina(n21534), .dinb(n21528), .dout(n21535));
  jand g21278(.dina(n21535), .dinb(asqrt[53] ), .dout(n21536));
  jor  g21279(.dina(n21535), .dinb(asqrt[53] ), .dout(n21537));
  jxor g21280(.dina(n20808), .dinb(n1173), .dout(n21538));
  jand g21281(.dina(n21538), .dinb(asqrt[6] ), .dout(n21539));
  jxor g21282(.dina(n21539), .dinb(n20813), .dout(n21540));
  jand g21283(.dina(n21540), .dinb(n21537), .dout(n21541));
  jor  g21284(.dina(n21541), .dinb(n21536), .dout(n21542));
  jand g21285(.dina(n21542), .dinb(asqrt[54] ), .dout(n21543));
  jor  g21286(.dina(n21542), .dinb(asqrt[54] ), .dout(n21544));
  jxor g21287(.dina(n20816), .dinb(n1008), .dout(n21545));
  jand g21288(.dina(n21545), .dinb(asqrt[6] ), .dout(n21546));
  jxor g21289(.dina(n21546), .dinb(n20821), .dout(n21547));
  jnot g21290(.din(n21547), .dout(n21548));
  jand g21291(.dina(n21548), .dinb(n21544), .dout(n21549));
  jor  g21292(.dina(n21549), .dinb(n21543), .dout(n21550));
  jand g21293(.dina(n21550), .dinb(asqrt[55] ), .dout(n21551));
  jor  g21294(.dina(n21550), .dinb(asqrt[55] ), .dout(n21552));
  jxor g21295(.dina(n20823), .dinb(n884), .dout(n21553));
  jand g21296(.dina(n21553), .dinb(asqrt[6] ), .dout(n21554));
  jxor g21297(.dina(n21554), .dinb(n20828), .dout(n21555));
  jnot g21298(.din(n21555), .dout(n21556));
  jand g21299(.dina(n21556), .dinb(n21552), .dout(n21557));
  jor  g21300(.dina(n21557), .dinb(n21551), .dout(n21558));
  jand g21301(.dina(n21558), .dinb(asqrt[56] ), .dout(n21559));
  jor  g21302(.dina(n21558), .dinb(asqrt[56] ), .dout(n21560));
  jxor g21303(.dina(n20830), .dinb(n743), .dout(n21561));
  jand g21304(.dina(n21561), .dinb(asqrt[6] ), .dout(n21562));
  jxor g21305(.dina(n21562), .dinb(n20835), .dout(n21563));
  jand g21306(.dina(n21563), .dinb(n21560), .dout(n21564));
  jor  g21307(.dina(n21564), .dinb(n21559), .dout(n21565));
  jand g21308(.dina(n21565), .dinb(asqrt[57] ), .dout(n21566));
  jor  g21309(.dina(n21565), .dinb(asqrt[57] ), .dout(n21567));
  jxor g21310(.dina(n20838), .dinb(n635), .dout(n21568));
  jand g21311(.dina(n21568), .dinb(asqrt[6] ), .dout(n21569));
  jxor g21312(.dina(n21569), .dinb(n20842), .dout(n21570));
  jand g21313(.dina(n21570), .dinb(n21567), .dout(n21571));
  jor  g21314(.dina(n21571), .dinb(n21566), .dout(n21572));
  jand g21315(.dina(n21572), .dinb(asqrt[58] ), .dout(n21573));
  jor  g21316(.dina(n21572), .dinb(asqrt[58] ), .dout(n21574));
  jxor g21317(.dina(n20846), .dinb(n515), .dout(n21575));
  jand g21318(.dina(n21575), .dinb(asqrt[6] ), .dout(n21576));
  jxor g21319(.dina(n21576), .dinb(n20851), .dout(n21577));
  jnot g21320(.din(n21577), .dout(n21578));
  jand g21321(.dina(n21578), .dinb(n21574), .dout(n21579));
  jor  g21322(.dina(n21579), .dinb(n21573), .dout(n21580));
  jand g21323(.dina(n21580), .dinb(asqrt[59] ), .dout(n21581));
  jor  g21324(.dina(n21580), .dinb(asqrt[59] ), .dout(n21582));
  jxor g21325(.dina(n20853), .dinb(n443), .dout(n21583));
  jand g21326(.dina(n21583), .dinb(asqrt[6] ), .dout(n21584));
  jxor g21327(.dina(n21584), .dinb(n20859), .dout(n21585));
  jnot g21328(.din(n21585), .dout(n21586));
  jand g21329(.dina(n21586), .dinb(n21582), .dout(n21587));
  jor  g21330(.dina(n21587), .dinb(n21581), .dout(n21588));
  jand g21331(.dina(n21588), .dinb(asqrt[60] ), .dout(n21589));
  jor  g21332(.dina(n21588), .dinb(asqrt[60] ), .dout(n21590));
  jxor g21333(.dina(n20861), .dinb(n352), .dout(n21591));
  jand g21334(.dina(n21591), .dinb(asqrt[6] ), .dout(n21592));
  jxor g21335(.dina(n21592), .dinb(n20866), .dout(n21593));
  jnot g21336(.din(n21593), .dout(n21594));
  jand g21337(.dina(n21594), .dinb(n21590), .dout(n21595));
  jor  g21338(.dina(n21595), .dinb(n21589), .dout(n21596));
  jand g21339(.dina(n21596), .dinb(asqrt[61] ), .dout(n21597));
  jor  g21340(.dina(n21596), .dinb(asqrt[61] ), .dout(n21598));
  jxor g21341(.dina(n20868), .dinb(n294), .dout(n21599));
  jand g21342(.dina(n21599), .dinb(asqrt[6] ), .dout(n21600));
  jxor g21343(.dina(n21600), .dinb(n20873), .dout(n21601));
  jnot g21344(.din(n21601), .dout(n21602));
  jand g21345(.dina(n21602), .dinb(n21598), .dout(n21603));
  jor  g21346(.dina(n21603), .dinb(n21597), .dout(n21604));
  jand g21347(.dina(n21604), .dinb(asqrt[62] ), .dout(n21605));
  jor  g21348(.dina(n21604), .dinb(asqrt[62] ), .dout(n21606));
  jxor g21349(.dina(n20875), .dinb(n239), .dout(n21607));
  jand g21350(.dina(n21607), .dinb(asqrt[6] ), .dout(n21608));
  jxor g21351(.dina(n21608), .dinb(n20880), .dout(n21609));
  jand g21352(.dina(n21609), .dinb(n21606), .dout(n21610));
  jor  g21353(.dina(n21610), .dinb(n21605), .dout(n21611));
  jxor g21354(.dina(n20883), .dinb(n221), .dout(n21612));
  jand g21355(.dina(n21612), .dinb(asqrt[6] ), .dout(n21613));
  jxor g21356(.dina(n21613), .dinb(n20888), .dout(n21614));
  jnot g21357(.din(n21614), .dout(n21615));
  jor  g21358(.dina(n21615), .dinb(n21611), .dout(n21616));
  jnot g21359(.din(n21616), .dout(n21617));
  jand g21360(.dina(asqrt[6] ), .dinb(n21176), .dout(n21618));
  jnot g21361(.din(n21605), .dout(n21619));
  jnot g21362(.din(n21597), .dout(n21620));
  jnot g21363(.din(n21589), .dout(n21621));
  jnot g21364(.din(n21581), .dout(n21622));
  jnot g21365(.din(n21573), .dout(n21623));
  jnot g21366(.din(n21566), .dout(n21624));
  jnot g21367(.din(n21559), .dout(n21625));
  jnot g21368(.din(n21551), .dout(n21626));
  jnot g21369(.din(n21543), .dout(n21627));
  jnot g21370(.din(n21536), .dout(n21628));
  jnot g21371(.din(n21528), .dout(n21629));
  jnot g21372(.din(n21521), .dout(n21630));
  jnot g21373(.din(n21513), .dout(n21631));
  jnot g21374(.din(n21505), .dout(n21632));
  jnot g21375(.din(n21497), .dout(n21633));
  jnot g21376(.din(n21489), .dout(n21634));
  jnot g21377(.din(n21481), .dout(n21635));
  jnot g21378(.din(n21474), .dout(n21636));
  jnot g21379(.din(n21466), .dout(n21637));
  jnot g21380(.din(n21458), .dout(n21638));
  jnot g21381(.din(n21450), .dout(n21639));
  jnot g21382(.din(n21443), .dout(n21640));
  jnot g21383(.din(n21435), .dout(n21641));
  jnot g21384(.din(n21428), .dout(n21642));
  jnot g21385(.din(n21420), .dout(n21643));
  jnot g21386(.din(n21413), .dout(n21644));
  jnot g21387(.din(n21405), .dout(n21645));
  jnot g21388(.din(n21398), .dout(n21646));
  jnot g21389(.din(n21390), .dout(n21647));
  jnot g21390(.din(n21382), .dout(n21648));
  jnot g21391(.din(n21374), .dout(n21649));
  jnot g21392(.din(n21367), .dout(n21650));
  jnot g21393(.din(n21359), .dout(n21651));
  jnot g21394(.din(n21352), .dout(n21652));
  jnot g21395(.din(n21344), .dout(n21653));
  jnot g21396(.din(n21337), .dout(n21654));
  jnot g21397(.din(n21330), .dout(n21655));
  jnot g21398(.din(n21322), .dout(n21656));
  jnot g21399(.din(n21314), .dout(n21657));
  jnot g21400(.din(n21307), .dout(n21658));
  jnot g21401(.din(n21299), .dout(n21659));
  jnot g21402(.din(n21292), .dout(n21660));
  jnot g21403(.din(n21284), .dout(n21661));
  jnot g21404(.din(n21277), .dout(n21662));
  jnot g21405(.din(n21269), .dout(n21663));
  jnot g21406(.din(n21261), .dout(n21664));
  jnot g21407(.din(n21253), .dout(n21665));
  jnot g21408(.din(n21246), .dout(n21666));
  jnot g21409(.din(n21238), .dout(n21667));
  jnot g21410(.din(n21230), .dout(n21668));
  jnot g21411(.din(n21222), .dout(n21669));
  jnot g21412(.din(n21215), .dout(n21670));
  jnot g21413(.din(n21207), .dout(n21671));
  jnot g21414(.din(n21200), .dout(n21672));
  jnot g21415(.din(n21189), .dout(n21673));
  jnot g21416(.din(n20913), .dout(n21674));
  jnot g21417(.din(n20910), .dout(n21675));
  jor  g21418(.dina(n21184), .dinb(n20473), .dout(n21676));
  jand g21419(.dina(n21676), .dinb(n21675), .dout(n21677));
  jand g21420(.dina(n21677), .dinb(n20468), .dout(n21678));
  jor  g21421(.dina(n21184), .dinb(a[12] ), .dout(n21679));
  jand g21422(.dina(n21679), .dinb(a[13] ), .dout(n21680));
  jor  g21423(.dina(n21191), .dinb(n21680), .dout(n21681));
  jor  g21424(.dina(n21681), .dinb(n21678), .dout(n21682));
  jand g21425(.dina(n21682), .dinb(n21674), .dout(n21683));
  jand g21426(.dina(n21683), .dinb(n19791), .dout(n21684));
  jor  g21427(.dina(n21196), .dinb(n21684), .dout(n21685));
  jand g21428(.dina(n21685), .dinb(n21673), .dout(n21686));
  jand g21429(.dina(n21686), .dinb(n19096), .dout(n21687));
  jnot g21430(.din(n21204), .dout(n21688));
  jor  g21431(.dina(n21688), .dinb(n21687), .dout(n21689));
  jand g21432(.dina(n21689), .dinb(n21672), .dout(n21690));
  jand g21433(.dina(n21690), .dinb(n18442), .dout(n21691));
  jor  g21434(.dina(n21211), .dinb(n21691), .dout(n21692));
  jand g21435(.dina(n21692), .dinb(n21671), .dout(n21693));
  jand g21436(.dina(n21693), .dinb(n17769), .dout(n21694));
  jnot g21437(.din(n21219), .dout(n21695));
  jor  g21438(.dina(n21695), .dinb(n21694), .dout(n21696));
  jand g21439(.dina(n21696), .dinb(n21670), .dout(n21697));
  jand g21440(.dina(n21697), .dinb(n17134), .dout(n21698));
  jor  g21441(.dina(n21226), .dinb(n21698), .dout(n21699));
  jand g21442(.dina(n21699), .dinb(n21669), .dout(n21700));
  jand g21443(.dina(n21700), .dinb(n16489), .dout(n21701));
  jor  g21444(.dina(n21234), .dinb(n21701), .dout(n21702));
  jand g21445(.dina(n21702), .dinb(n21668), .dout(n21703));
  jand g21446(.dina(n21703), .dinb(n15878), .dout(n21704));
  jor  g21447(.dina(n21242), .dinb(n21704), .dout(n21705));
  jand g21448(.dina(n21705), .dinb(n21667), .dout(n21706));
  jand g21449(.dina(n21706), .dinb(n15260), .dout(n21707));
  jnot g21450(.din(n21250), .dout(n21708));
  jor  g21451(.dina(n21708), .dinb(n21707), .dout(n21709));
  jand g21452(.dina(n21709), .dinb(n21666), .dout(n21710));
  jand g21453(.dina(n21710), .dinb(n14674), .dout(n21711));
  jor  g21454(.dina(n21257), .dinb(n21711), .dout(n21712));
  jand g21455(.dina(n21712), .dinb(n21665), .dout(n21713));
  jand g21456(.dina(n21713), .dinb(n14078), .dout(n21714));
  jor  g21457(.dina(n21265), .dinb(n21714), .dout(n21715));
  jand g21458(.dina(n21715), .dinb(n21664), .dout(n21716));
  jand g21459(.dina(n21716), .dinb(n13515), .dout(n21717));
  jor  g21460(.dina(n21273), .dinb(n21717), .dout(n21718));
  jand g21461(.dina(n21718), .dinb(n21663), .dout(n21719));
  jand g21462(.dina(n21719), .dinb(n12947), .dout(n21720));
  jnot g21463(.din(n21281), .dout(n21721));
  jor  g21464(.dina(n21721), .dinb(n21720), .dout(n21722));
  jand g21465(.dina(n21722), .dinb(n21662), .dout(n21723));
  jand g21466(.dina(n21723), .dinb(n12410), .dout(n21724));
  jor  g21467(.dina(n21288), .dinb(n21724), .dout(n21725));
  jand g21468(.dina(n21725), .dinb(n21661), .dout(n21726));
  jand g21469(.dina(n21726), .dinb(n11858), .dout(n21727));
  jnot g21470(.din(n21296), .dout(n21728));
  jor  g21471(.dina(n21728), .dinb(n21727), .dout(n21729));
  jand g21472(.dina(n21729), .dinb(n21660), .dout(n21730));
  jand g21473(.dina(n21730), .dinb(n11347), .dout(n21731));
  jor  g21474(.dina(n21303), .dinb(n21731), .dout(n21732));
  jand g21475(.dina(n21732), .dinb(n21659), .dout(n21733));
  jand g21476(.dina(n21733), .dinb(n10824), .dout(n21734));
  jnot g21477(.din(n21311), .dout(n21735));
  jor  g21478(.dina(n21735), .dinb(n21734), .dout(n21736));
  jand g21479(.dina(n21736), .dinb(n21658), .dout(n21737));
  jand g21480(.dina(n21737), .dinb(n10328), .dout(n21738));
  jor  g21481(.dina(n21318), .dinb(n21738), .dout(n21739));
  jand g21482(.dina(n21739), .dinb(n21657), .dout(n21740));
  jand g21483(.dina(n21740), .dinb(n9832), .dout(n21741));
  jor  g21484(.dina(n21326), .dinb(n21741), .dout(n21742));
  jand g21485(.dina(n21742), .dinb(n21656), .dout(n21743));
  jand g21486(.dina(n21743), .dinb(n9369), .dout(n21744));
  jnot g21487(.din(n21334), .dout(n21745));
  jor  g21488(.dina(n21745), .dinb(n21744), .dout(n21746));
  jand g21489(.dina(n21746), .dinb(n21655), .dout(n21747));
  jand g21490(.dina(n21747), .dinb(n8890), .dout(n21748));
  jnot g21491(.din(n21341), .dout(n21749));
  jor  g21492(.dina(n21749), .dinb(n21748), .dout(n21750));
  jand g21493(.dina(n21750), .dinb(n21654), .dout(n21751));
  jand g21494(.dina(n21751), .dinb(n8449), .dout(n21752));
  jor  g21495(.dina(n21348), .dinb(n21752), .dout(n21753));
  jand g21496(.dina(n21753), .dinb(n21653), .dout(n21754));
  jand g21497(.dina(n21754), .dinb(n8003), .dout(n21755));
  jnot g21498(.din(n21356), .dout(n21756));
  jor  g21499(.dina(n21756), .dinb(n21755), .dout(n21757));
  jand g21500(.dina(n21757), .dinb(n21652), .dout(n21758));
  jand g21501(.dina(n21758), .dinb(n7581), .dout(n21759));
  jor  g21502(.dina(n21363), .dinb(n21759), .dout(n21760));
  jand g21503(.dina(n21760), .dinb(n21651), .dout(n21761));
  jand g21504(.dina(n21761), .dinb(n7154), .dout(n21762));
  jnot g21505(.din(n21371), .dout(n21763));
  jor  g21506(.dina(n21763), .dinb(n21762), .dout(n21764));
  jand g21507(.dina(n21764), .dinb(n21650), .dout(n21765));
  jand g21508(.dina(n21765), .dinb(n6758), .dout(n21766));
  jor  g21509(.dina(n21378), .dinb(n21766), .dout(n21767));
  jand g21510(.dina(n21767), .dinb(n21649), .dout(n21768));
  jand g21511(.dina(n21768), .dinb(n6357), .dout(n21769));
  jor  g21512(.dina(n21386), .dinb(n21769), .dout(n21770));
  jand g21513(.dina(n21770), .dinb(n21648), .dout(n21771));
  jand g21514(.dina(n21771), .dinb(n5989), .dout(n21772));
  jor  g21515(.dina(n21394), .dinb(n21772), .dout(n21773));
  jand g21516(.dina(n21773), .dinb(n21647), .dout(n21774));
  jand g21517(.dina(n21774), .dinb(n5606), .dout(n21775));
  jnot g21518(.din(n21402), .dout(n21776));
  jor  g21519(.dina(n21776), .dinb(n21775), .dout(n21777));
  jand g21520(.dina(n21777), .dinb(n21646), .dout(n21778));
  jand g21521(.dina(n21778), .dinb(n5259), .dout(n21779));
  jor  g21522(.dina(n21409), .dinb(n21779), .dout(n21780));
  jand g21523(.dina(n21780), .dinb(n21645), .dout(n21781));
  jand g21524(.dina(n21781), .dinb(n4902), .dout(n21782));
  jnot g21525(.din(n21417), .dout(n21783));
  jor  g21526(.dina(n21783), .dinb(n21782), .dout(n21784));
  jand g21527(.dina(n21784), .dinb(n21644), .dout(n21785));
  jand g21528(.dina(n21785), .dinb(n4582), .dout(n21786));
  jor  g21529(.dina(n21424), .dinb(n21786), .dout(n21787));
  jand g21530(.dina(n21787), .dinb(n21643), .dout(n21788));
  jand g21531(.dina(n21788), .dinb(n4249), .dout(n21789));
  jnot g21532(.din(n21432), .dout(n21790));
  jor  g21533(.dina(n21790), .dinb(n21789), .dout(n21791));
  jand g21534(.dina(n21791), .dinb(n21642), .dout(n21792));
  jand g21535(.dina(n21792), .dinb(n3955), .dout(n21793));
  jor  g21536(.dina(n21439), .dinb(n21793), .dout(n21794));
  jand g21537(.dina(n21794), .dinb(n21641), .dout(n21795));
  jand g21538(.dina(n21795), .dinb(n3642), .dout(n21796));
  jnot g21539(.din(n21447), .dout(n21797));
  jor  g21540(.dina(n21797), .dinb(n21796), .dout(n21798));
  jand g21541(.dina(n21798), .dinb(n21640), .dout(n21799));
  jand g21542(.dina(n21799), .dinb(n3368), .dout(n21800));
  jor  g21543(.dina(n21454), .dinb(n21800), .dout(n21801));
  jand g21544(.dina(n21801), .dinb(n21639), .dout(n21802));
  jand g21545(.dina(n21802), .dinb(n3089), .dout(n21803));
  jor  g21546(.dina(n21462), .dinb(n21803), .dout(n21804));
  jand g21547(.dina(n21804), .dinb(n21638), .dout(n21805));
  jand g21548(.dina(n21805), .dinb(n2833), .dout(n21806));
  jor  g21549(.dina(n21470), .dinb(n21806), .dout(n21807));
  jand g21550(.dina(n21807), .dinb(n21637), .dout(n21808));
  jand g21551(.dina(n21808), .dinb(n2572), .dout(n21809));
  jnot g21552(.din(n21478), .dout(n21810));
  jor  g21553(.dina(n21810), .dinb(n21809), .dout(n21811));
  jand g21554(.dina(n21811), .dinb(n21636), .dout(n21812));
  jand g21555(.dina(n21812), .dinb(n2345), .dout(n21813));
  jor  g21556(.dina(n21485), .dinb(n21813), .dout(n21814));
  jand g21557(.dina(n21814), .dinb(n21635), .dout(n21815));
  jand g21558(.dina(n21815), .dinb(n2108), .dout(n21816));
  jor  g21559(.dina(n21493), .dinb(n21816), .dout(n21817));
  jand g21560(.dina(n21817), .dinb(n21634), .dout(n21818));
  jand g21561(.dina(n21818), .dinb(n1912), .dout(n21819));
  jor  g21562(.dina(n21501), .dinb(n21819), .dout(n21820));
  jand g21563(.dina(n21820), .dinb(n21633), .dout(n21821));
  jand g21564(.dina(n21821), .dinb(n1699), .dout(n21822));
  jor  g21565(.dina(n21509), .dinb(n21822), .dout(n21823));
  jand g21566(.dina(n21823), .dinb(n21632), .dout(n21824));
  jand g21567(.dina(n21824), .dinb(n1516), .dout(n21825));
  jor  g21568(.dina(n21517), .dinb(n21825), .dout(n21826));
  jand g21569(.dina(n21826), .dinb(n21631), .dout(n21827));
  jand g21570(.dina(n21827), .dinb(n1332), .dout(n21828));
  jnot g21571(.din(n21525), .dout(n21829));
  jor  g21572(.dina(n21829), .dinb(n21828), .dout(n21830));
  jand g21573(.dina(n21830), .dinb(n21630), .dout(n21831));
  jand g21574(.dina(n21831), .dinb(n1173), .dout(n21832));
  jor  g21575(.dina(n21532), .dinb(n21832), .dout(n21833));
  jand g21576(.dina(n21833), .dinb(n21629), .dout(n21834));
  jand g21577(.dina(n21834), .dinb(n1008), .dout(n21835));
  jnot g21578(.din(n21540), .dout(n21836));
  jor  g21579(.dina(n21836), .dinb(n21835), .dout(n21837));
  jand g21580(.dina(n21837), .dinb(n21628), .dout(n21838));
  jand g21581(.dina(n21838), .dinb(n884), .dout(n21839));
  jor  g21582(.dina(n21547), .dinb(n21839), .dout(n21840));
  jand g21583(.dina(n21840), .dinb(n21627), .dout(n21841));
  jand g21584(.dina(n21841), .dinb(n743), .dout(n21842));
  jor  g21585(.dina(n21555), .dinb(n21842), .dout(n21843));
  jand g21586(.dina(n21843), .dinb(n21626), .dout(n21844));
  jand g21587(.dina(n21844), .dinb(n635), .dout(n21845));
  jnot g21588(.din(n21563), .dout(n21846));
  jor  g21589(.dina(n21846), .dinb(n21845), .dout(n21847));
  jand g21590(.dina(n21847), .dinb(n21625), .dout(n21848));
  jand g21591(.dina(n21848), .dinb(n515), .dout(n21849));
  jnot g21592(.din(n21570), .dout(n21850));
  jor  g21593(.dina(n21850), .dinb(n21849), .dout(n21851));
  jand g21594(.dina(n21851), .dinb(n21624), .dout(n21852));
  jand g21595(.dina(n21852), .dinb(n443), .dout(n21853));
  jor  g21596(.dina(n21577), .dinb(n21853), .dout(n21854));
  jand g21597(.dina(n21854), .dinb(n21623), .dout(n21855));
  jand g21598(.dina(n21855), .dinb(n352), .dout(n21856));
  jor  g21599(.dina(n21585), .dinb(n21856), .dout(n21857));
  jand g21600(.dina(n21857), .dinb(n21622), .dout(n21858));
  jand g21601(.dina(n21858), .dinb(n294), .dout(n21859));
  jor  g21602(.dina(n21593), .dinb(n21859), .dout(n21860));
  jand g21603(.dina(n21860), .dinb(n21621), .dout(n21861));
  jand g21604(.dina(n21861), .dinb(n239), .dout(n21862));
  jor  g21605(.dina(n21601), .dinb(n21862), .dout(n21863));
  jand g21606(.dina(n21863), .dinb(n21620), .dout(n21864));
  jand g21607(.dina(n21864), .dinb(n221), .dout(n21865));
  jnot g21608(.din(n21609), .dout(n21866));
  jor  g21609(.dina(n21866), .dinb(n21865), .dout(n21867));
  jand g21610(.dina(n21867), .dinb(n21619), .dout(n21868));
  jor  g21611(.dina(n21614), .dinb(n21868), .dout(n21869));
  jor  g21612(.dina(n21869), .dinb(n20897), .dout(n21870));
  jor  g21613(.dina(n21870), .dinb(n21618), .dout(n21871));
  jand g21614(.dina(n21871), .dinb(n218), .dout(n21872));
  jand g21615(.dina(n21184), .dinb(n20890), .dout(n21873));
  jnot g21616(.din(n21873), .dout(n21874));
  jand g21617(.dina(n20891), .dinb(asqrt[63] ), .dout(n21875));
  jand g21618(.dina(n21875), .dinb(n21181), .dout(n21876));
  jand g21619(.dina(n21876), .dinb(n21874), .dout(n21877));
  jor  g21620(.dina(n21877), .dinb(n21872), .dout(n21878));
  jor  g21621(.dina(n21878), .dinb(n21617), .dout(asqrt[5] ));
  jnot g21622(.din(n21618), .dout(n21880));
  jand g21623(.dina(n21615), .dinb(n21611), .dout(n21881));
  jand g21624(.dina(n21881), .dinb(n21181), .dout(n21882));
  jand g21625(.dina(n21882), .dinb(n21880), .dout(n21883));
  jor  g21626(.dina(n21883), .dinb(asqrt[63] ), .dout(n21884));
  jnot g21627(.din(n21877), .dout(n21885));
  jand g21628(.dina(n21885), .dinb(n21884), .dout(n21886));
  jand g21629(.dina(n21886), .dinb(n21616), .dout(n21887));
  jor  g21630(.dina(n21887), .dinb(n20907), .dout(n21888));
  jnot g21631(.din(a[8] ), .dout(n21889));
  jnot g21632(.din(a[9] ), .dout(n21890));
  jand g21633(.dina(n21890), .dinb(n21889), .dout(n21891));
  jand g21634(.dina(n21891), .dinb(n20907), .dout(n21892));
  jnot g21635(.din(n21892), .dout(n21893));
  jand g21636(.dina(n21893), .dinb(n21888), .dout(n21894));
  jor  g21637(.dina(n21894), .dinb(n21184), .dout(n21895));
  jand g21638(.dina(n21894), .dinb(n21184), .dout(n21896));
  jor  g21639(.dina(n21887), .dinb(a[10] ), .dout(n21897));
  jand g21640(.dina(n21897), .dinb(a[11] ), .dout(n21898));
  jand g21641(.dina(asqrt[5] ), .dinb(n20909), .dout(n21899));
  jor  g21642(.dina(n21899), .dinb(n21898), .dout(n21900));
  jor  g21643(.dina(n21900), .dinb(n21896), .dout(n21901));
  jand g21644(.dina(n21901), .dinb(n21895), .dout(n21902));
  jor  g21645(.dina(n21902), .dinb(n20468), .dout(n21903));
  jand g21646(.dina(n21902), .dinb(n20468), .dout(n21904));
  jnot g21647(.din(n20909), .dout(n21905));
  jor  g21648(.dina(n21887), .dinb(n21905), .dout(n21906));
  jor  g21649(.dina(asqrt[5] ), .dinb(n21184), .dout(n21907));
  jand g21650(.dina(n21907), .dinb(n21906), .dout(n21908));
  jxor g21651(.dina(n21908), .dinb(n20473), .dout(n21909));
  jor  g21652(.dina(n21909), .dinb(n21904), .dout(n21910));
  jand g21653(.dina(n21910), .dinb(n21903), .dout(n21911));
  jor  g21654(.dina(n21911), .dinb(n19791), .dout(n21912));
  jand g21655(.dina(n21911), .dinb(n19791), .dout(n21913));
  jxor g21656(.dina(n20912), .dinb(n20468), .dout(n21914));
  jor  g21657(.dina(n21914), .dinb(n21887), .dout(n21915));
  jxor g21658(.dina(n21915), .dinb(n21681), .dout(n21916));
  jnot g21659(.din(n21916), .dout(n21917));
  jor  g21660(.dina(n21917), .dinb(n21913), .dout(n21918));
  jand g21661(.dina(n21918), .dinb(n21912), .dout(n21919));
  jor  g21662(.dina(n21919), .dinb(n19096), .dout(n21920));
  jand g21663(.dina(n21919), .dinb(n19096), .dout(n21921));
  jxor g21664(.dina(n21188), .dinb(n19791), .dout(n21922));
  jor  g21665(.dina(n21922), .dinb(n21887), .dout(n21923));
  jxor g21666(.dina(n21923), .dinb(n21197), .dout(n21924));
  jor  g21667(.dina(n21924), .dinb(n21921), .dout(n21925));
  jand g21668(.dina(n21925), .dinb(n21920), .dout(n21926));
  jor  g21669(.dina(n21926), .dinb(n18442), .dout(n21927));
  jand g21670(.dina(n21926), .dinb(n18442), .dout(n21928));
  jxor g21671(.dina(n21199), .dinb(n19096), .dout(n21929));
  jor  g21672(.dina(n21929), .dinb(n21887), .dout(n21930));
  jxor g21673(.dina(n21930), .dinb(n21688), .dout(n21931));
  jnot g21674(.din(n21931), .dout(n21932));
  jor  g21675(.dina(n21932), .dinb(n21928), .dout(n21933));
  jand g21676(.dina(n21933), .dinb(n21927), .dout(n21934));
  jor  g21677(.dina(n21934), .dinb(n17769), .dout(n21935));
  jand g21678(.dina(n21934), .dinb(n17769), .dout(n21936));
  jxor g21679(.dina(n21206), .dinb(n18442), .dout(n21937));
  jor  g21680(.dina(n21937), .dinb(n21887), .dout(n21938));
  jxor g21681(.dina(n21938), .dinb(n21212), .dout(n21939));
  jor  g21682(.dina(n21939), .dinb(n21936), .dout(n21940));
  jand g21683(.dina(n21940), .dinb(n21935), .dout(n21941));
  jor  g21684(.dina(n21941), .dinb(n17134), .dout(n21942));
  jand g21685(.dina(n21941), .dinb(n17134), .dout(n21943));
  jxor g21686(.dina(n21214), .dinb(n17769), .dout(n21944));
  jor  g21687(.dina(n21944), .dinb(n21887), .dout(n21945));
  jxor g21688(.dina(n21945), .dinb(n21695), .dout(n21946));
  jnot g21689(.din(n21946), .dout(n21947));
  jor  g21690(.dina(n21947), .dinb(n21943), .dout(n21948));
  jand g21691(.dina(n21948), .dinb(n21942), .dout(n21949));
  jor  g21692(.dina(n21949), .dinb(n16489), .dout(n21950));
  jand g21693(.dina(n21949), .dinb(n16489), .dout(n21951));
  jxor g21694(.dina(n21221), .dinb(n17134), .dout(n21952));
  jor  g21695(.dina(n21952), .dinb(n21887), .dout(n21953));
  jxor g21696(.dina(n21953), .dinb(n21227), .dout(n21954));
  jor  g21697(.dina(n21954), .dinb(n21951), .dout(n21955));
  jand g21698(.dina(n21955), .dinb(n21950), .dout(n21956));
  jor  g21699(.dina(n21956), .dinb(n15878), .dout(n21957));
  jand g21700(.dina(n21956), .dinb(n15878), .dout(n21958));
  jxor g21701(.dina(n21229), .dinb(n16489), .dout(n21959));
  jor  g21702(.dina(n21959), .dinb(n21887), .dout(n21960));
  jxor g21703(.dina(n21960), .dinb(n21235), .dout(n21961));
  jor  g21704(.dina(n21961), .dinb(n21958), .dout(n21962));
  jand g21705(.dina(n21962), .dinb(n21957), .dout(n21963));
  jor  g21706(.dina(n21963), .dinb(n15260), .dout(n21964));
  jand g21707(.dina(n21963), .dinb(n15260), .dout(n21965));
  jxor g21708(.dina(n21237), .dinb(n15878), .dout(n21966));
  jor  g21709(.dina(n21966), .dinb(n21887), .dout(n21967));
  jxor g21710(.dina(n21967), .dinb(n21243), .dout(n21968));
  jor  g21711(.dina(n21968), .dinb(n21965), .dout(n21969));
  jand g21712(.dina(n21969), .dinb(n21964), .dout(n21970));
  jor  g21713(.dina(n21970), .dinb(n14674), .dout(n21971));
  jand g21714(.dina(n21970), .dinb(n14674), .dout(n21972));
  jxor g21715(.dina(n21245), .dinb(n15260), .dout(n21973));
  jor  g21716(.dina(n21973), .dinb(n21887), .dout(n21974));
  jxor g21717(.dina(n21974), .dinb(n21708), .dout(n21975));
  jnot g21718(.din(n21975), .dout(n21976));
  jor  g21719(.dina(n21976), .dinb(n21972), .dout(n21977));
  jand g21720(.dina(n21977), .dinb(n21971), .dout(n21978));
  jor  g21721(.dina(n21978), .dinb(n14078), .dout(n21979));
  jand g21722(.dina(n21978), .dinb(n14078), .dout(n21980));
  jxor g21723(.dina(n21252), .dinb(n14674), .dout(n21981));
  jor  g21724(.dina(n21981), .dinb(n21887), .dout(n21982));
  jxor g21725(.dina(n21982), .dinb(n21258), .dout(n21983));
  jor  g21726(.dina(n21983), .dinb(n21980), .dout(n21984));
  jand g21727(.dina(n21984), .dinb(n21979), .dout(n21985));
  jor  g21728(.dina(n21985), .dinb(n13515), .dout(n21986));
  jand g21729(.dina(n21985), .dinb(n13515), .dout(n21987));
  jxor g21730(.dina(n21260), .dinb(n14078), .dout(n21988));
  jor  g21731(.dina(n21988), .dinb(n21887), .dout(n21989));
  jxor g21732(.dina(n21989), .dinb(n21266), .dout(n21990));
  jor  g21733(.dina(n21990), .dinb(n21987), .dout(n21991));
  jand g21734(.dina(n21991), .dinb(n21986), .dout(n21992));
  jor  g21735(.dina(n21992), .dinb(n12947), .dout(n21993));
  jand g21736(.dina(n21992), .dinb(n12947), .dout(n21994));
  jxor g21737(.dina(n21268), .dinb(n13515), .dout(n21995));
  jor  g21738(.dina(n21995), .dinb(n21887), .dout(n21996));
  jxor g21739(.dina(n21996), .dinb(n21274), .dout(n21997));
  jor  g21740(.dina(n21997), .dinb(n21994), .dout(n21998));
  jand g21741(.dina(n21998), .dinb(n21993), .dout(n21999));
  jor  g21742(.dina(n21999), .dinb(n12410), .dout(n22000));
  jand g21743(.dina(n21999), .dinb(n12410), .dout(n22001));
  jxor g21744(.dina(n21276), .dinb(n12947), .dout(n22002));
  jor  g21745(.dina(n22002), .dinb(n21887), .dout(n22003));
  jxor g21746(.dina(n22003), .dinb(n21721), .dout(n22004));
  jnot g21747(.din(n22004), .dout(n22005));
  jor  g21748(.dina(n22005), .dinb(n22001), .dout(n22006));
  jand g21749(.dina(n22006), .dinb(n22000), .dout(n22007));
  jor  g21750(.dina(n22007), .dinb(n11858), .dout(n22008));
  jand g21751(.dina(n22007), .dinb(n11858), .dout(n22009));
  jxor g21752(.dina(n21283), .dinb(n12410), .dout(n22010));
  jor  g21753(.dina(n22010), .dinb(n21887), .dout(n22011));
  jxor g21754(.dina(n22011), .dinb(n21289), .dout(n22012));
  jor  g21755(.dina(n22012), .dinb(n22009), .dout(n22013));
  jand g21756(.dina(n22013), .dinb(n22008), .dout(n22014));
  jor  g21757(.dina(n22014), .dinb(n11347), .dout(n22015));
  jand g21758(.dina(n22014), .dinb(n11347), .dout(n22016));
  jxor g21759(.dina(n21291), .dinb(n11858), .dout(n22017));
  jor  g21760(.dina(n22017), .dinb(n21887), .dout(n22018));
  jxor g21761(.dina(n22018), .dinb(n21728), .dout(n22019));
  jnot g21762(.din(n22019), .dout(n22020));
  jor  g21763(.dina(n22020), .dinb(n22016), .dout(n22021));
  jand g21764(.dina(n22021), .dinb(n22015), .dout(n22022));
  jor  g21765(.dina(n22022), .dinb(n10824), .dout(n22023));
  jand g21766(.dina(n22022), .dinb(n10824), .dout(n22024));
  jxor g21767(.dina(n21298), .dinb(n11347), .dout(n22025));
  jor  g21768(.dina(n22025), .dinb(n21887), .dout(n22026));
  jxor g21769(.dina(n22026), .dinb(n21304), .dout(n22027));
  jor  g21770(.dina(n22027), .dinb(n22024), .dout(n22028));
  jand g21771(.dina(n22028), .dinb(n22023), .dout(n22029));
  jor  g21772(.dina(n22029), .dinb(n10328), .dout(n22030));
  jand g21773(.dina(n22029), .dinb(n10328), .dout(n22031));
  jxor g21774(.dina(n21306), .dinb(n10824), .dout(n22032));
  jor  g21775(.dina(n22032), .dinb(n21887), .dout(n22033));
  jxor g21776(.dina(n22033), .dinb(n21735), .dout(n22034));
  jnot g21777(.din(n22034), .dout(n22035));
  jor  g21778(.dina(n22035), .dinb(n22031), .dout(n22036));
  jand g21779(.dina(n22036), .dinb(n22030), .dout(n22037));
  jor  g21780(.dina(n22037), .dinb(n9832), .dout(n22038));
  jand g21781(.dina(n22037), .dinb(n9832), .dout(n22039));
  jxor g21782(.dina(n21313), .dinb(n10328), .dout(n22040));
  jor  g21783(.dina(n22040), .dinb(n21887), .dout(n22041));
  jxor g21784(.dina(n22041), .dinb(n21319), .dout(n22042));
  jor  g21785(.dina(n22042), .dinb(n22039), .dout(n22043));
  jand g21786(.dina(n22043), .dinb(n22038), .dout(n22044));
  jor  g21787(.dina(n22044), .dinb(n9369), .dout(n22045));
  jand g21788(.dina(n22044), .dinb(n9369), .dout(n22046));
  jxor g21789(.dina(n21321), .dinb(n9832), .dout(n22047));
  jor  g21790(.dina(n22047), .dinb(n21887), .dout(n22048));
  jxor g21791(.dina(n22048), .dinb(n21327), .dout(n22049));
  jor  g21792(.dina(n22049), .dinb(n22046), .dout(n22050));
  jand g21793(.dina(n22050), .dinb(n22045), .dout(n22051));
  jor  g21794(.dina(n22051), .dinb(n8890), .dout(n22052));
  jand g21795(.dina(n22051), .dinb(n8890), .dout(n22053));
  jxor g21796(.dina(n21329), .dinb(n9369), .dout(n22054));
  jor  g21797(.dina(n22054), .dinb(n21887), .dout(n22055));
  jxor g21798(.dina(n22055), .dinb(n21745), .dout(n22056));
  jnot g21799(.din(n22056), .dout(n22057));
  jor  g21800(.dina(n22057), .dinb(n22053), .dout(n22058));
  jand g21801(.dina(n22058), .dinb(n22052), .dout(n22059));
  jor  g21802(.dina(n22059), .dinb(n8449), .dout(n22060));
  jand g21803(.dina(n22059), .dinb(n8449), .dout(n22061));
  jxor g21804(.dina(n21336), .dinb(n8890), .dout(n22062));
  jor  g21805(.dina(n22062), .dinb(n21887), .dout(n22063));
  jxor g21806(.dina(n22063), .dinb(n21749), .dout(n22064));
  jnot g21807(.din(n22064), .dout(n22065));
  jor  g21808(.dina(n22065), .dinb(n22061), .dout(n22066));
  jand g21809(.dina(n22066), .dinb(n22060), .dout(n22067));
  jor  g21810(.dina(n22067), .dinb(n8003), .dout(n22068));
  jand g21811(.dina(n22067), .dinb(n8003), .dout(n22069));
  jxor g21812(.dina(n21343), .dinb(n8449), .dout(n22070));
  jor  g21813(.dina(n22070), .dinb(n21887), .dout(n22071));
  jxor g21814(.dina(n22071), .dinb(n21349), .dout(n22072));
  jor  g21815(.dina(n22072), .dinb(n22069), .dout(n22073));
  jand g21816(.dina(n22073), .dinb(n22068), .dout(n22074));
  jor  g21817(.dina(n22074), .dinb(n7581), .dout(n22075));
  jand g21818(.dina(n22074), .dinb(n7581), .dout(n22076));
  jxor g21819(.dina(n21351), .dinb(n8003), .dout(n22077));
  jor  g21820(.dina(n22077), .dinb(n21887), .dout(n22078));
  jxor g21821(.dina(n22078), .dinb(n21756), .dout(n22079));
  jnot g21822(.din(n22079), .dout(n22080));
  jor  g21823(.dina(n22080), .dinb(n22076), .dout(n22081));
  jand g21824(.dina(n22081), .dinb(n22075), .dout(n22082));
  jor  g21825(.dina(n22082), .dinb(n7154), .dout(n22083));
  jand g21826(.dina(n22082), .dinb(n7154), .dout(n22084));
  jxor g21827(.dina(n21358), .dinb(n7581), .dout(n22085));
  jor  g21828(.dina(n22085), .dinb(n21887), .dout(n22086));
  jxor g21829(.dina(n22086), .dinb(n21364), .dout(n22087));
  jor  g21830(.dina(n22087), .dinb(n22084), .dout(n22088));
  jand g21831(.dina(n22088), .dinb(n22083), .dout(n22089));
  jor  g21832(.dina(n22089), .dinb(n6758), .dout(n22090));
  jand g21833(.dina(n22089), .dinb(n6758), .dout(n22091));
  jxor g21834(.dina(n21366), .dinb(n7154), .dout(n22092));
  jor  g21835(.dina(n22092), .dinb(n21887), .dout(n22093));
  jxor g21836(.dina(n22093), .dinb(n21763), .dout(n22094));
  jnot g21837(.din(n22094), .dout(n22095));
  jor  g21838(.dina(n22095), .dinb(n22091), .dout(n22096));
  jand g21839(.dina(n22096), .dinb(n22090), .dout(n22097));
  jor  g21840(.dina(n22097), .dinb(n6357), .dout(n22098));
  jand g21841(.dina(n22097), .dinb(n6357), .dout(n22099));
  jxor g21842(.dina(n21373), .dinb(n6758), .dout(n22100));
  jor  g21843(.dina(n22100), .dinb(n21887), .dout(n22101));
  jxor g21844(.dina(n22101), .dinb(n21379), .dout(n22102));
  jor  g21845(.dina(n22102), .dinb(n22099), .dout(n22103));
  jand g21846(.dina(n22103), .dinb(n22098), .dout(n22104));
  jor  g21847(.dina(n22104), .dinb(n5989), .dout(n22105));
  jand g21848(.dina(n22104), .dinb(n5989), .dout(n22106));
  jxor g21849(.dina(n21381), .dinb(n6357), .dout(n22107));
  jor  g21850(.dina(n22107), .dinb(n21887), .dout(n22108));
  jxor g21851(.dina(n22108), .dinb(n21387), .dout(n22109));
  jor  g21852(.dina(n22109), .dinb(n22106), .dout(n22110));
  jand g21853(.dina(n22110), .dinb(n22105), .dout(n22111));
  jor  g21854(.dina(n22111), .dinb(n5606), .dout(n22112));
  jand g21855(.dina(n22111), .dinb(n5606), .dout(n22113));
  jxor g21856(.dina(n21389), .dinb(n5989), .dout(n22114));
  jor  g21857(.dina(n22114), .dinb(n21887), .dout(n22115));
  jxor g21858(.dina(n22115), .dinb(n21395), .dout(n22116));
  jor  g21859(.dina(n22116), .dinb(n22113), .dout(n22117));
  jand g21860(.dina(n22117), .dinb(n22112), .dout(n22118));
  jor  g21861(.dina(n22118), .dinb(n5259), .dout(n22119));
  jand g21862(.dina(n22118), .dinb(n5259), .dout(n22120));
  jxor g21863(.dina(n21397), .dinb(n5606), .dout(n22121));
  jor  g21864(.dina(n22121), .dinb(n21887), .dout(n22122));
  jxor g21865(.dina(n22122), .dinb(n21776), .dout(n22123));
  jnot g21866(.din(n22123), .dout(n22124));
  jor  g21867(.dina(n22124), .dinb(n22120), .dout(n22125));
  jand g21868(.dina(n22125), .dinb(n22119), .dout(n22126));
  jor  g21869(.dina(n22126), .dinb(n4902), .dout(n22127));
  jand g21870(.dina(n22126), .dinb(n4902), .dout(n22128));
  jxor g21871(.dina(n21404), .dinb(n5259), .dout(n22129));
  jor  g21872(.dina(n22129), .dinb(n21887), .dout(n22130));
  jxor g21873(.dina(n22130), .dinb(n21410), .dout(n22131));
  jor  g21874(.dina(n22131), .dinb(n22128), .dout(n22132));
  jand g21875(.dina(n22132), .dinb(n22127), .dout(n22133));
  jor  g21876(.dina(n22133), .dinb(n4582), .dout(n22134));
  jand g21877(.dina(n22133), .dinb(n4582), .dout(n22135));
  jxor g21878(.dina(n21412), .dinb(n4902), .dout(n22136));
  jor  g21879(.dina(n22136), .dinb(n21887), .dout(n22137));
  jxor g21880(.dina(n22137), .dinb(n21783), .dout(n22138));
  jnot g21881(.din(n22138), .dout(n22139));
  jor  g21882(.dina(n22139), .dinb(n22135), .dout(n22140));
  jand g21883(.dina(n22140), .dinb(n22134), .dout(n22141));
  jor  g21884(.dina(n22141), .dinb(n4249), .dout(n22142));
  jand g21885(.dina(n22141), .dinb(n4249), .dout(n22143));
  jxor g21886(.dina(n21419), .dinb(n4582), .dout(n22144));
  jor  g21887(.dina(n22144), .dinb(n21887), .dout(n22145));
  jxor g21888(.dina(n22145), .dinb(n21425), .dout(n22146));
  jor  g21889(.dina(n22146), .dinb(n22143), .dout(n22147));
  jand g21890(.dina(n22147), .dinb(n22142), .dout(n22148));
  jor  g21891(.dina(n22148), .dinb(n3955), .dout(n22149));
  jand g21892(.dina(n22148), .dinb(n3955), .dout(n22150));
  jxor g21893(.dina(n21427), .dinb(n4249), .dout(n22151));
  jor  g21894(.dina(n22151), .dinb(n21887), .dout(n22152));
  jxor g21895(.dina(n22152), .dinb(n21790), .dout(n22153));
  jnot g21896(.din(n22153), .dout(n22154));
  jor  g21897(.dina(n22154), .dinb(n22150), .dout(n22155));
  jand g21898(.dina(n22155), .dinb(n22149), .dout(n22156));
  jor  g21899(.dina(n22156), .dinb(n3642), .dout(n22157));
  jand g21900(.dina(n22156), .dinb(n3642), .dout(n22158));
  jxor g21901(.dina(n21434), .dinb(n3955), .dout(n22159));
  jor  g21902(.dina(n22159), .dinb(n21887), .dout(n22160));
  jxor g21903(.dina(n22160), .dinb(n21440), .dout(n22161));
  jor  g21904(.dina(n22161), .dinb(n22158), .dout(n22162));
  jand g21905(.dina(n22162), .dinb(n22157), .dout(n22163));
  jor  g21906(.dina(n22163), .dinb(n3368), .dout(n22164));
  jand g21907(.dina(n22163), .dinb(n3368), .dout(n22165));
  jxor g21908(.dina(n21442), .dinb(n3642), .dout(n22166));
  jor  g21909(.dina(n22166), .dinb(n21887), .dout(n22167));
  jxor g21910(.dina(n22167), .dinb(n21797), .dout(n22168));
  jnot g21911(.din(n22168), .dout(n22169));
  jor  g21912(.dina(n22169), .dinb(n22165), .dout(n22170));
  jand g21913(.dina(n22170), .dinb(n22164), .dout(n22171));
  jor  g21914(.dina(n22171), .dinb(n3089), .dout(n22172));
  jand g21915(.dina(n22171), .dinb(n3089), .dout(n22173));
  jxor g21916(.dina(n21449), .dinb(n3368), .dout(n22174));
  jor  g21917(.dina(n22174), .dinb(n21887), .dout(n22175));
  jxor g21918(.dina(n22175), .dinb(n21455), .dout(n22176));
  jor  g21919(.dina(n22176), .dinb(n22173), .dout(n22177));
  jand g21920(.dina(n22177), .dinb(n22172), .dout(n22178));
  jor  g21921(.dina(n22178), .dinb(n2833), .dout(n22179));
  jand g21922(.dina(n22178), .dinb(n2833), .dout(n22180));
  jxor g21923(.dina(n21457), .dinb(n3089), .dout(n22181));
  jor  g21924(.dina(n22181), .dinb(n21887), .dout(n22182));
  jxor g21925(.dina(n22182), .dinb(n21463), .dout(n22183));
  jor  g21926(.dina(n22183), .dinb(n22180), .dout(n22184));
  jand g21927(.dina(n22184), .dinb(n22179), .dout(n22185));
  jor  g21928(.dina(n22185), .dinb(n2572), .dout(n22186));
  jand g21929(.dina(n22185), .dinb(n2572), .dout(n22187));
  jxor g21930(.dina(n21465), .dinb(n2833), .dout(n22188));
  jor  g21931(.dina(n22188), .dinb(n21887), .dout(n22189));
  jxor g21932(.dina(n22189), .dinb(n21471), .dout(n22190));
  jor  g21933(.dina(n22190), .dinb(n22187), .dout(n22191));
  jand g21934(.dina(n22191), .dinb(n22186), .dout(n22192));
  jor  g21935(.dina(n22192), .dinb(n2345), .dout(n22193));
  jand g21936(.dina(n22192), .dinb(n2345), .dout(n22194));
  jxor g21937(.dina(n21473), .dinb(n2572), .dout(n22195));
  jor  g21938(.dina(n22195), .dinb(n21887), .dout(n22196));
  jxor g21939(.dina(n22196), .dinb(n21810), .dout(n22197));
  jnot g21940(.din(n22197), .dout(n22198));
  jor  g21941(.dina(n22198), .dinb(n22194), .dout(n22199));
  jand g21942(.dina(n22199), .dinb(n22193), .dout(n22200));
  jor  g21943(.dina(n22200), .dinb(n2108), .dout(n22201));
  jand g21944(.dina(n22200), .dinb(n2108), .dout(n22202));
  jxor g21945(.dina(n21480), .dinb(n2345), .dout(n22203));
  jor  g21946(.dina(n22203), .dinb(n21887), .dout(n22204));
  jxor g21947(.dina(n22204), .dinb(n21486), .dout(n22205));
  jor  g21948(.dina(n22205), .dinb(n22202), .dout(n22206));
  jand g21949(.dina(n22206), .dinb(n22201), .dout(n22207));
  jor  g21950(.dina(n22207), .dinb(n1912), .dout(n22208));
  jand g21951(.dina(n22207), .dinb(n1912), .dout(n22209));
  jxor g21952(.dina(n21488), .dinb(n2108), .dout(n22210));
  jor  g21953(.dina(n22210), .dinb(n21887), .dout(n22211));
  jxor g21954(.dina(n22211), .dinb(n21494), .dout(n22212));
  jor  g21955(.dina(n22212), .dinb(n22209), .dout(n22213));
  jand g21956(.dina(n22213), .dinb(n22208), .dout(n22214));
  jor  g21957(.dina(n22214), .dinb(n1699), .dout(n22215));
  jand g21958(.dina(n22214), .dinb(n1699), .dout(n22216));
  jxor g21959(.dina(n21496), .dinb(n1912), .dout(n22217));
  jor  g21960(.dina(n22217), .dinb(n21887), .dout(n22218));
  jxor g21961(.dina(n22218), .dinb(n21502), .dout(n22219));
  jor  g21962(.dina(n22219), .dinb(n22216), .dout(n22220));
  jand g21963(.dina(n22220), .dinb(n22215), .dout(n22221));
  jor  g21964(.dina(n22221), .dinb(n1516), .dout(n22222));
  jand g21965(.dina(n22221), .dinb(n1516), .dout(n22223));
  jxor g21966(.dina(n21504), .dinb(n1699), .dout(n22224));
  jor  g21967(.dina(n22224), .dinb(n21887), .dout(n22225));
  jxor g21968(.dina(n22225), .dinb(n21510), .dout(n22226));
  jor  g21969(.dina(n22226), .dinb(n22223), .dout(n22227));
  jand g21970(.dina(n22227), .dinb(n22222), .dout(n22228));
  jor  g21971(.dina(n22228), .dinb(n1332), .dout(n22229));
  jand g21972(.dina(n22228), .dinb(n1332), .dout(n22230));
  jxor g21973(.dina(n21512), .dinb(n1516), .dout(n22231));
  jor  g21974(.dina(n22231), .dinb(n21887), .dout(n22232));
  jxor g21975(.dina(n22232), .dinb(n21518), .dout(n22233));
  jor  g21976(.dina(n22233), .dinb(n22230), .dout(n22234));
  jand g21977(.dina(n22234), .dinb(n22229), .dout(n22235));
  jor  g21978(.dina(n22235), .dinb(n1173), .dout(n22236));
  jand g21979(.dina(n22235), .dinb(n1173), .dout(n22237));
  jxor g21980(.dina(n21520), .dinb(n1332), .dout(n22238));
  jor  g21981(.dina(n22238), .dinb(n21887), .dout(n22239));
  jxor g21982(.dina(n22239), .dinb(n21829), .dout(n22240));
  jnot g21983(.din(n22240), .dout(n22241));
  jor  g21984(.dina(n22241), .dinb(n22237), .dout(n22242));
  jand g21985(.dina(n22242), .dinb(n22236), .dout(n22243));
  jor  g21986(.dina(n22243), .dinb(n1008), .dout(n22244));
  jand g21987(.dina(n22243), .dinb(n1008), .dout(n22245));
  jxor g21988(.dina(n21527), .dinb(n1173), .dout(n22246));
  jor  g21989(.dina(n22246), .dinb(n21887), .dout(n22247));
  jxor g21990(.dina(n22247), .dinb(n21533), .dout(n22248));
  jor  g21991(.dina(n22248), .dinb(n22245), .dout(n22249));
  jand g21992(.dina(n22249), .dinb(n22244), .dout(n22250));
  jor  g21993(.dina(n22250), .dinb(n884), .dout(n22251));
  jand g21994(.dina(n22250), .dinb(n884), .dout(n22252));
  jxor g21995(.dina(n21535), .dinb(n1008), .dout(n22253));
  jor  g21996(.dina(n22253), .dinb(n21887), .dout(n22254));
  jxor g21997(.dina(n22254), .dinb(n21836), .dout(n22255));
  jnot g21998(.din(n22255), .dout(n22256));
  jor  g21999(.dina(n22256), .dinb(n22252), .dout(n22257));
  jand g22000(.dina(n22257), .dinb(n22251), .dout(n22258));
  jor  g22001(.dina(n22258), .dinb(n743), .dout(n22259));
  jand g22002(.dina(n22258), .dinb(n743), .dout(n22260));
  jxor g22003(.dina(n21542), .dinb(n884), .dout(n22261));
  jor  g22004(.dina(n22261), .dinb(n21887), .dout(n22262));
  jxor g22005(.dina(n22262), .dinb(n21548), .dout(n22263));
  jor  g22006(.dina(n22263), .dinb(n22260), .dout(n22264));
  jand g22007(.dina(n22264), .dinb(n22259), .dout(n22265));
  jor  g22008(.dina(n22265), .dinb(n635), .dout(n22266));
  jand g22009(.dina(n22265), .dinb(n635), .dout(n22267));
  jxor g22010(.dina(n21550), .dinb(n743), .dout(n22268));
  jor  g22011(.dina(n22268), .dinb(n21887), .dout(n22269));
  jxor g22012(.dina(n22269), .dinb(n21556), .dout(n22270));
  jor  g22013(.dina(n22270), .dinb(n22267), .dout(n22271));
  jand g22014(.dina(n22271), .dinb(n22266), .dout(n22272));
  jor  g22015(.dina(n22272), .dinb(n515), .dout(n22273));
  jand g22016(.dina(n22272), .dinb(n515), .dout(n22274));
  jxor g22017(.dina(n21558), .dinb(n635), .dout(n22275));
  jor  g22018(.dina(n22275), .dinb(n21887), .dout(n22276));
  jxor g22019(.dina(n22276), .dinb(n21846), .dout(n22277));
  jnot g22020(.din(n22277), .dout(n22278));
  jor  g22021(.dina(n22278), .dinb(n22274), .dout(n22279));
  jand g22022(.dina(n22279), .dinb(n22273), .dout(n22280));
  jor  g22023(.dina(n22280), .dinb(n443), .dout(n22281));
  jand g22024(.dina(n22280), .dinb(n443), .dout(n22282));
  jxor g22025(.dina(n21565), .dinb(n515), .dout(n22283));
  jor  g22026(.dina(n22283), .dinb(n21887), .dout(n22284));
  jxor g22027(.dina(n22284), .dinb(n21850), .dout(n22285));
  jnot g22028(.din(n22285), .dout(n22286));
  jor  g22029(.dina(n22286), .dinb(n22282), .dout(n22287));
  jand g22030(.dina(n22287), .dinb(n22281), .dout(n22288));
  jor  g22031(.dina(n22288), .dinb(n352), .dout(n22289));
  jand g22032(.dina(n22288), .dinb(n352), .dout(n22290));
  jxor g22033(.dina(n21572), .dinb(n443), .dout(n22291));
  jor  g22034(.dina(n22291), .dinb(n21887), .dout(n22292));
  jxor g22035(.dina(n22292), .dinb(n21578), .dout(n22293));
  jor  g22036(.dina(n22293), .dinb(n22290), .dout(n22294));
  jand g22037(.dina(n22294), .dinb(n22289), .dout(n22295));
  jor  g22038(.dina(n22295), .dinb(n294), .dout(n22296));
  jand g22039(.dina(n22295), .dinb(n294), .dout(n22297));
  jxor g22040(.dina(n21580), .dinb(n352), .dout(n22298));
  jor  g22041(.dina(n22298), .dinb(n21887), .dout(n22299));
  jxor g22042(.dina(n22299), .dinb(n21586), .dout(n22300));
  jor  g22043(.dina(n22300), .dinb(n22297), .dout(n22301));
  jand g22044(.dina(n22301), .dinb(n22296), .dout(n22302));
  jor  g22045(.dina(n22302), .dinb(n239), .dout(n22303));
  jand g22046(.dina(n22302), .dinb(n239), .dout(n22304));
  jxor g22047(.dina(n21588), .dinb(n294), .dout(n22305));
  jor  g22048(.dina(n22305), .dinb(n21887), .dout(n22306));
  jxor g22049(.dina(n22306), .dinb(n21594), .dout(n22307));
  jor  g22050(.dina(n22307), .dinb(n22304), .dout(n22308));
  jand g22051(.dina(n22308), .dinb(n22303), .dout(n22309));
  jor  g22052(.dina(n22309), .dinb(n221), .dout(n22310));
  jand g22053(.dina(n22309), .dinb(n221), .dout(n22311));
  jxor g22054(.dina(n21596), .dinb(n239), .dout(n22312));
  jor  g22055(.dina(n22312), .dinb(n21887), .dout(n22313));
  jxor g22056(.dina(n22313), .dinb(n21601), .dout(n22314));
  jnot g22057(.din(n22314), .dout(n22315));
  jor  g22058(.dina(n22315), .dinb(n22311), .dout(n22316));
  jand g22059(.dina(n22316), .dinb(n22310), .dout(n22317));
  jxor g22060(.dina(n21604), .dinb(n221), .dout(n22318));
  jor  g22061(.dina(n22318), .dinb(n21887), .dout(n22319));
  jxor g22062(.dina(n22319), .dinb(n21609), .dout(n22320));
  jand g22063(.dina(n22320), .dinb(n22317), .dout(n22321));
  jor  g22064(.dina(n22320), .dinb(n22317), .dout(n22322));
  jxor g22065(.dina(n21615), .dinb(n21611), .dout(n22323));
  jnot g22066(.din(n22323), .dout(n22324));
  jand g22067(.dina(n22324), .dinb(asqrt[5] ), .dout(n22325));
  jor  g22068(.dina(n22325), .dinb(n22322), .dout(n22326));
  jand g22069(.dina(n22326), .dinb(n218), .dout(n22327));
  jand g22070(.dina(n21887), .dinb(n21868), .dout(n22328));
  jor  g22071(.dina(n22328), .dinb(n22324), .dout(n22329));
  jor  g22072(.dina(n22329), .dinb(n218), .dout(n22330));
  jnot g22073(.din(n22330), .dout(n22331));
  jor  g22074(.dina(n22331), .dinb(n22327), .dout(n22332));
  jor  g22075(.dina(n22332), .dinb(n22321), .dout(asqrt[4] ));
  jnot g22076(.din(a[6] ), .dout(n22334));
  jnot g22077(.din(a[7] ), .dout(n22335));
  jand g22078(.dina(n22335), .dinb(n22334), .dout(n22336));
  jand g22079(.dina(n22336), .dinb(n21889), .dout(n22337));
  jand g22080(.dina(asqrt[4] ), .dinb(a[8] ), .dout(n22338));
  jor  g22081(.dina(n22338), .dinb(n22337), .dout(n22339));
  jand g22082(.dina(n22339), .dinb(asqrt[5] ), .dout(n22340));
  jor  g22083(.dina(n22339), .dinb(asqrt[5] ), .dout(n22341));
  jand g22084(.dina(asqrt[4] ), .dinb(n21889), .dout(n22342));
  jor  g22085(.dina(n22342), .dinb(n21890), .dout(n22343));
  jnot g22086(.din(n21891), .dout(n22344));
  jnot g22087(.din(n22321), .dout(n22345));
  jnot g22088(.din(n22310), .dout(n22346));
  jnot g22089(.din(n22303), .dout(n22347));
  jnot g22090(.din(n22296), .dout(n22348));
  jnot g22091(.din(n22289), .dout(n22349));
  jnot g22092(.din(n22281), .dout(n22350));
  jnot g22093(.din(n22273), .dout(n22351));
  jnot g22094(.din(n22266), .dout(n22352));
  jnot g22095(.din(n22259), .dout(n22353));
  jnot g22096(.din(n22251), .dout(n22354));
  jnot g22097(.din(n22244), .dout(n22355));
  jnot g22098(.din(n22236), .dout(n22356));
  jnot g22099(.din(n22229), .dout(n22357));
  jnot g22100(.din(n22222), .dout(n22358));
  jnot g22101(.din(n22215), .dout(n22359));
  jnot g22102(.din(n22208), .dout(n22360));
  jnot g22103(.din(n22201), .dout(n22361));
  jnot g22104(.din(n22193), .dout(n22362));
  jnot g22105(.din(n22186), .dout(n22363));
  jnot g22106(.din(n22179), .dout(n22364));
  jnot g22107(.din(n22172), .dout(n22365));
  jnot g22108(.din(n22164), .dout(n22366));
  jnot g22109(.din(n22157), .dout(n22367));
  jnot g22110(.din(n22149), .dout(n22368));
  jnot g22111(.din(n22142), .dout(n22369));
  jnot g22112(.din(n22134), .dout(n22370));
  jnot g22113(.din(n22127), .dout(n22371));
  jnot g22114(.din(n22119), .dout(n22372));
  jnot g22115(.din(n22112), .dout(n22373));
  jnot g22116(.din(n22105), .dout(n22374));
  jnot g22117(.din(n22098), .dout(n22375));
  jnot g22118(.din(n22090), .dout(n22376));
  jnot g22119(.din(n22083), .dout(n22377));
  jnot g22120(.din(n22075), .dout(n22378));
  jnot g22121(.din(n22068), .dout(n22379));
  jnot g22122(.din(n22060), .dout(n22380));
  jnot g22123(.din(n22052), .dout(n22381));
  jnot g22124(.din(n22045), .dout(n22382));
  jnot g22125(.din(n22038), .dout(n22383));
  jnot g22126(.din(n22030), .dout(n22384));
  jnot g22127(.din(n22023), .dout(n22385));
  jnot g22128(.din(n22015), .dout(n22386));
  jnot g22129(.din(n22008), .dout(n22387));
  jnot g22130(.din(n22000), .dout(n22388));
  jnot g22131(.din(n21993), .dout(n22389));
  jnot g22132(.din(n21986), .dout(n22390));
  jnot g22133(.din(n21979), .dout(n22391));
  jnot g22134(.din(n21971), .dout(n22392));
  jnot g22135(.din(n21964), .dout(n22393));
  jnot g22136(.din(n21957), .dout(n22394));
  jnot g22137(.din(n21950), .dout(n22395));
  jnot g22138(.din(n21942), .dout(n22396));
  jnot g22139(.din(n21935), .dout(n22397));
  jnot g22140(.din(n21927), .dout(n22398));
  jnot g22141(.din(n21920), .dout(n22399));
  jnot g22142(.din(n21912), .dout(n22400));
  jnot g22143(.din(n21903), .dout(n22401));
  jnot g22144(.din(n21895), .dout(n22402));
  jand g22145(.dina(asqrt[5] ), .dinb(a[10] ), .dout(n22403));
  jor  g22146(.dina(n21892), .dinb(n22403), .dout(n22404));
  jor  g22147(.dina(n22404), .dinb(asqrt[6] ), .dout(n22405));
  jand g22148(.dina(asqrt[5] ), .dinb(n20907), .dout(n22406));
  jor  g22149(.dina(n22406), .dinb(n20908), .dout(n22407));
  jand g22150(.dina(n21906), .dinb(n22407), .dout(n22408));
  jand g22151(.dina(n22408), .dinb(n22405), .dout(n22409));
  jor  g22152(.dina(n22409), .dinb(n22402), .dout(n22410));
  jor  g22153(.dina(n22410), .dinb(asqrt[7] ), .dout(n22411));
  jnot g22154(.din(n21909), .dout(n22412));
  jand g22155(.dina(n22412), .dinb(n22411), .dout(n22413));
  jor  g22156(.dina(n22413), .dinb(n22401), .dout(n22414));
  jor  g22157(.dina(n22414), .dinb(asqrt[8] ), .dout(n22415));
  jand g22158(.dina(n21916), .dinb(n22415), .dout(n22416));
  jor  g22159(.dina(n22416), .dinb(n22400), .dout(n22417));
  jor  g22160(.dina(n22417), .dinb(asqrt[9] ), .dout(n22418));
  jnot g22161(.din(n21924), .dout(n22419));
  jand g22162(.dina(n22419), .dinb(n22418), .dout(n22420));
  jor  g22163(.dina(n22420), .dinb(n22399), .dout(n22421));
  jor  g22164(.dina(n22421), .dinb(asqrt[10] ), .dout(n22422));
  jand g22165(.dina(n21931), .dinb(n22422), .dout(n22423));
  jor  g22166(.dina(n22423), .dinb(n22398), .dout(n22424));
  jor  g22167(.dina(n22424), .dinb(asqrt[11] ), .dout(n22425));
  jnot g22168(.din(n21939), .dout(n22426));
  jand g22169(.dina(n22426), .dinb(n22425), .dout(n22427));
  jor  g22170(.dina(n22427), .dinb(n22397), .dout(n22428));
  jor  g22171(.dina(n22428), .dinb(asqrt[12] ), .dout(n22429));
  jand g22172(.dina(n21946), .dinb(n22429), .dout(n22430));
  jor  g22173(.dina(n22430), .dinb(n22396), .dout(n22431));
  jor  g22174(.dina(n22431), .dinb(asqrt[13] ), .dout(n22432));
  jnot g22175(.din(n21954), .dout(n22433));
  jand g22176(.dina(n22433), .dinb(n22432), .dout(n22434));
  jor  g22177(.dina(n22434), .dinb(n22395), .dout(n22435));
  jor  g22178(.dina(n22435), .dinb(asqrt[14] ), .dout(n22436));
  jnot g22179(.din(n21961), .dout(n22437));
  jand g22180(.dina(n22437), .dinb(n22436), .dout(n22438));
  jor  g22181(.dina(n22438), .dinb(n22394), .dout(n22439));
  jor  g22182(.dina(n22439), .dinb(asqrt[15] ), .dout(n22440));
  jnot g22183(.din(n21968), .dout(n22441));
  jand g22184(.dina(n22441), .dinb(n22440), .dout(n22442));
  jor  g22185(.dina(n22442), .dinb(n22393), .dout(n22443));
  jor  g22186(.dina(n22443), .dinb(asqrt[16] ), .dout(n22444));
  jand g22187(.dina(n21975), .dinb(n22444), .dout(n22445));
  jor  g22188(.dina(n22445), .dinb(n22392), .dout(n22446));
  jor  g22189(.dina(n22446), .dinb(asqrt[17] ), .dout(n22447));
  jnot g22190(.din(n21983), .dout(n22448));
  jand g22191(.dina(n22448), .dinb(n22447), .dout(n22449));
  jor  g22192(.dina(n22449), .dinb(n22391), .dout(n22450));
  jor  g22193(.dina(n22450), .dinb(asqrt[18] ), .dout(n22451));
  jnot g22194(.din(n21990), .dout(n22452));
  jand g22195(.dina(n22452), .dinb(n22451), .dout(n22453));
  jor  g22196(.dina(n22453), .dinb(n22390), .dout(n22454));
  jor  g22197(.dina(n22454), .dinb(asqrt[19] ), .dout(n22455));
  jnot g22198(.din(n21997), .dout(n22456));
  jand g22199(.dina(n22456), .dinb(n22455), .dout(n22457));
  jor  g22200(.dina(n22457), .dinb(n22389), .dout(n22458));
  jor  g22201(.dina(n22458), .dinb(asqrt[20] ), .dout(n22459));
  jand g22202(.dina(n22004), .dinb(n22459), .dout(n22460));
  jor  g22203(.dina(n22460), .dinb(n22388), .dout(n22461));
  jor  g22204(.dina(n22461), .dinb(asqrt[21] ), .dout(n22462));
  jnot g22205(.din(n22012), .dout(n22463));
  jand g22206(.dina(n22463), .dinb(n22462), .dout(n22464));
  jor  g22207(.dina(n22464), .dinb(n22387), .dout(n22465));
  jor  g22208(.dina(n22465), .dinb(asqrt[22] ), .dout(n22466));
  jand g22209(.dina(n22019), .dinb(n22466), .dout(n22467));
  jor  g22210(.dina(n22467), .dinb(n22386), .dout(n22468));
  jor  g22211(.dina(n22468), .dinb(asqrt[23] ), .dout(n22469));
  jnot g22212(.din(n22027), .dout(n22470));
  jand g22213(.dina(n22470), .dinb(n22469), .dout(n22471));
  jor  g22214(.dina(n22471), .dinb(n22385), .dout(n22472));
  jor  g22215(.dina(n22472), .dinb(asqrt[24] ), .dout(n22473));
  jand g22216(.dina(n22034), .dinb(n22473), .dout(n22474));
  jor  g22217(.dina(n22474), .dinb(n22384), .dout(n22475));
  jor  g22218(.dina(n22475), .dinb(asqrt[25] ), .dout(n22476));
  jnot g22219(.din(n22042), .dout(n22477));
  jand g22220(.dina(n22477), .dinb(n22476), .dout(n22478));
  jor  g22221(.dina(n22478), .dinb(n22383), .dout(n22479));
  jor  g22222(.dina(n22479), .dinb(asqrt[26] ), .dout(n22480));
  jnot g22223(.din(n22049), .dout(n22481));
  jand g22224(.dina(n22481), .dinb(n22480), .dout(n22482));
  jor  g22225(.dina(n22482), .dinb(n22382), .dout(n22483));
  jor  g22226(.dina(n22483), .dinb(asqrt[27] ), .dout(n22484));
  jand g22227(.dina(n22056), .dinb(n22484), .dout(n22485));
  jor  g22228(.dina(n22485), .dinb(n22381), .dout(n22486));
  jor  g22229(.dina(n22486), .dinb(asqrt[28] ), .dout(n22487));
  jand g22230(.dina(n22064), .dinb(n22487), .dout(n22488));
  jor  g22231(.dina(n22488), .dinb(n22380), .dout(n22489));
  jor  g22232(.dina(n22489), .dinb(asqrt[29] ), .dout(n22490));
  jnot g22233(.din(n22072), .dout(n22491));
  jand g22234(.dina(n22491), .dinb(n22490), .dout(n22492));
  jor  g22235(.dina(n22492), .dinb(n22379), .dout(n22493));
  jor  g22236(.dina(n22493), .dinb(asqrt[30] ), .dout(n22494));
  jand g22237(.dina(n22079), .dinb(n22494), .dout(n22495));
  jor  g22238(.dina(n22495), .dinb(n22378), .dout(n22496));
  jor  g22239(.dina(n22496), .dinb(asqrt[31] ), .dout(n22497));
  jnot g22240(.din(n22087), .dout(n22498));
  jand g22241(.dina(n22498), .dinb(n22497), .dout(n22499));
  jor  g22242(.dina(n22499), .dinb(n22377), .dout(n22500));
  jor  g22243(.dina(n22500), .dinb(asqrt[32] ), .dout(n22501));
  jand g22244(.dina(n22094), .dinb(n22501), .dout(n22502));
  jor  g22245(.dina(n22502), .dinb(n22376), .dout(n22503));
  jor  g22246(.dina(n22503), .dinb(asqrt[33] ), .dout(n22504));
  jnot g22247(.din(n22102), .dout(n22505));
  jand g22248(.dina(n22505), .dinb(n22504), .dout(n22506));
  jor  g22249(.dina(n22506), .dinb(n22375), .dout(n22507));
  jor  g22250(.dina(n22507), .dinb(asqrt[34] ), .dout(n22508));
  jnot g22251(.din(n22109), .dout(n22509));
  jand g22252(.dina(n22509), .dinb(n22508), .dout(n22510));
  jor  g22253(.dina(n22510), .dinb(n22374), .dout(n22511));
  jor  g22254(.dina(n22511), .dinb(asqrt[35] ), .dout(n22512));
  jnot g22255(.din(n22116), .dout(n22513));
  jand g22256(.dina(n22513), .dinb(n22512), .dout(n22514));
  jor  g22257(.dina(n22514), .dinb(n22373), .dout(n22515));
  jor  g22258(.dina(n22515), .dinb(asqrt[36] ), .dout(n22516));
  jand g22259(.dina(n22123), .dinb(n22516), .dout(n22517));
  jor  g22260(.dina(n22517), .dinb(n22372), .dout(n22518));
  jor  g22261(.dina(n22518), .dinb(asqrt[37] ), .dout(n22519));
  jnot g22262(.din(n22131), .dout(n22520));
  jand g22263(.dina(n22520), .dinb(n22519), .dout(n22521));
  jor  g22264(.dina(n22521), .dinb(n22371), .dout(n22522));
  jor  g22265(.dina(n22522), .dinb(asqrt[38] ), .dout(n22523));
  jand g22266(.dina(n22138), .dinb(n22523), .dout(n22524));
  jor  g22267(.dina(n22524), .dinb(n22370), .dout(n22525));
  jor  g22268(.dina(n22525), .dinb(asqrt[39] ), .dout(n22526));
  jnot g22269(.din(n22146), .dout(n22527));
  jand g22270(.dina(n22527), .dinb(n22526), .dout(n22528));
  jor  g22271(.dina(n22528), .dinb(n22369), .dout(n22529));
  jor  g22272(.dina(n22529), .dinb(asqrt[40] ), .dout(n22530));
  jand g22273(.dina(n22153), .dinb(n22530), .dout(n22531));
  jor  g22274(.dina(n22531), .dinb(n22368), .dout(n22532));
  jor  g22275(.dina(n22532), .dinb(asqrt[41] ), .dout(n22533));
  jnot g22276(.din(n22161), .dout(n22534));
  jand g22277(.dina(n22534), .dinb(n22533), .dout(n22535));
  jor  g22278(.dina(n22535), .dinb(n22367), .dout(n22536));
  jor  g22279(.dina(n22536), .dinb(asqrt[42] ), .dout(n22537));
  jand g22280(.dina(n22168), .dinb(n22537), .dout(n22538));
  jor  g22281(.dina(n22538), .dinb(n22366), .dout(n22539));
  jor  g22282(.dina(n22539), .dinb(asqrt[43] ), .dout(n22540));
  jnot g22283(.din(n22176), .dout(n22541));
  jand g22284(.dina(n22541), .dinb(n22540), .dout(n22542));
  jor  g22285(.dina(n22542), .dinb(n22365), .dout(n22543));
  jor  g22286(.dina(n22543), .dinb(asqrt[44] ), .dout(n22544));
  jnot g22287(.din(n22183), .dout(n22545));
  jand g22288(.dina(n22545), .dinb(n22544), .dout(n22546));
  jor  g22289(.dina(n22546), .dinb(n22364), .dout(n22547));
  jor  g22290(.dina(n22547), .dinb(asqrt[45] ), .dout(n22548));
  jnot g22291(.din(n22190), .dout(n22549));
  jand g22292(.dina(n22549), .dinb(n22548), .dout(n22550));
  jor  g22293(.dina(n22550), .dinb(n22363), .dout(n22551));
  jor  g22294(.dina(n22551), .dinb(asqrt[46] ), .dout(n22552));
  jand g22295(.dina(n22197), .dinb(n22552), .dout(n22553));
  jor  g22296(.dina(n22553), .dinb(n22362), .dout(n22554));
  jor  g22297(.dina(n22554), .dinb(asqrt[47] ), .dout(n22555));
  jnot g22298(.din(n22205), .dout(n22556));
  jand g22299(.dina(n22556), .dinb(n22555), .dout(n22557));
  jor  g22300(.dina(n22557), .dinb(n22361), .dout(n22558));
  jor  g22301(.dina(n22558), .dinb(asqrt[48] ), .dout(n22559));
  jnot g22302(.din(n22212), .dout(n22560));
  jand g22303(.dina(n22560), .dinb(n22559), .dout(n22561));
  jor  g22304(.dina(n22561), .dinb(n22360), .dout(n22562));
  jor  g22305(.dina(n22562), .dinb(asqrt[49] ), .dout(n22563));
  jnot g22306(.din(n22219), .dout(n22564));
  jand g22307(.dina(n22564), .dinb(n22563), .dout(n22565));
  jor  g22308(.dina(n22565), .dinb(n22359), .dout(n22566));
  jor  g22309(.dina(n22566), .dinb(asqrt[50] ), .dout(n22567));
  jnot g22310(.din(n22226), .dout(n22568));
  jand g22311(.dina(n22568), .dinb(n22567), .dout(n22569));
  jor  g22312(.dina(n22569), .dinb(n22358), .dout(n22570));
  jor  g22313(.dina(n22570), .dinb(asqrt[51] ), .dout(n22571));
  jnot g22314(.din(n22233), .dout(n22572));
  jand g22315(.dina(n22572), .dinb(n22571), .dout(n22573));
  jor  g22316(.dina(n22573), .dinb(n22357), .dout(n22574));
  jor  g22317(.dina(n22574), .dinb(asqrt[52] ), .dout(n22575));
  jand g22318(.dina(n22240), .dinb(n22575), .dout(n22576));
  jor  g22319(.dina(n22576), .dinb(n22356), .dout(n22577));
  jor  g22320(.dina(n22577), .dinb(asqrt[53] ), .dout(n22578));
  jnot g22321(.din(n22248), .dout(n22579));
  jand g22322(.dina(n22579), .dinb(n22578), .dout(n22580));
  jor  g22323(.dina(n22580), .dinb(n22355), .dout(n22581));
  jor  g22324(.dina(n22581), .dinb(asqrt[54] ), .dout(n22582));
  jand g22325(.dina(n22255), .dinb(n22582), .dout(n22583));
  jor  g22326(.dina(n22583), .dinb(n22354), .dout(n22584));
  jor  g22327(.dina(n22584), .dinb(asqrt[55] ), .dout(n22585));
  jnot g22328(.din(n22263), .dout(n22586));
  jand g22329(.dina(n22586), .dinb(n22585), .dout(n22587));
  jor  g22330(.dina(n22587), .dinb(n22353), .dout(n22588));
  jor  g22331(.dina(n22588), .dinb(asqrt[56] ), .dout(n22589));
  jnot g22332(.din(n22270), .dout(n22590));
  jand g22333(.dina(n22590), .dinb(n22589), .dout(n22591));
  jor  g22334(.dina(n22591), .dinb(n22352), .dout(n22592));
  jor  g22335(.dina(n22592), .dinb(asqrt[57] ), .dout(n22593));
  jand g22336(.dina(n22277), .dinb(n22593), .dout(n22594));
  jor  g22337(.dina(n22594), .dinb(n22351), .dout(n22595));
  jor  g22338(.dina(n22595), .dinb(asqrt[58] ), .dout(n22596));
  jand g22339(.dina(n22285), .dinb(n22596), .dout(n22597));
  jor  g22340(.dina(n22597), .dinb(n22350), .dout(n22598));
  jor  g22341(.dina(n22598), .dinb(asqrt[59] ), .dout(n22599));
  jnot g22342(.din(n22293), .dout(n22600));
  jand g22343(.dina(n22600), .dinb(n22599), .dout(n22601));
  jor  g22344(.dina(n22601), .dinb(n22349), .dout(n22602));
  jor  g22345(.dina(n22602), .dinb(asqrt[60] ), .dout(n22603));
  jnot g22346(.din(n22300), .dout(n22604));
  jand g22347(.dina(n22604), .dinb(n22603), .dout(n22605));
  jor  g22348(.dina(n22605), .dinb(n22348), .dout(n22606));
  jor  g22349(.dina(n22606), .dinb(asqrt[61] ), .dout(n22607));
  jnot g22350(.din(n22307), .dout(n22608));
  jand g22351(.dina(n22608), .dinb(n22607), .dout(n22609));
  jor  g22352(.dina(n22609), .dinb(n22347), .dout(n22610));
  jor  g22353(.dina(n22610), .dinb(asqrt[62] ), .dout(n22611));
  jand g22354(.dina(n22314), .dinb(n22611), .dout(n22612));
  jor  g22355(.dina(n22612), .dinb(n22346), .dout(n22613));
  jnot g22356(.din(n22320), .dout(n22614));
  jand g22357(.dina(n22614), .dinb(n22613), .dout(n22615));
  jnot g22358(.din(n22325), .dout(n22616));
  jand g22359(.dina(n22616), .dinb(n22615), .dout(n22617));
  jor  g22360(.dina(n22617), .dinb(asqrt[63] ), .dout(n22618));
  jand g22361(.dina(n22330), .dinb(n22618), .dout(n22619));
  jand g22362(.dina(n22619), .dinb(n22345), .dout(n22620));
  jor  g22363(.dina(n22620), .dinb(n22344), .dout(n22621));
  jand g22364(.dina(n22621), .dinb(n22343), .dout(n22622));
  jand g22365(.dina(n22622), .dinb(n22341), .dout(n22623));
  jor  g22366(.dina(n22623), .dinb(n22340), .dout(n22624));
  jand g22367(.dina(n22624), .dinb(asqrt[6] ), .dout(n22625));
  jor  g22368(.dina(n22624), .dinb(asqrt[6] ), .dout(n22626));
  jor  g22369(.dina(asqrt[4] ), .dinb(n21887), .dout(n22627));
  jand g22370(.dina(n22627), .dinb(n22621), .dout(n22628));
  jxor g22371(.dina(n22628), .dinb(n20907), .dout(n22629));
  jnot g22372(.din(n22629), .dout(n22630));
  jand g22373(.dina(n22630), .dinb(n22626), .dout(n22631));
  jor  g22374(.dina(n22631), .dinb(n22625), .dout(n22632));
  jand g22375(.dina(n22632), .dinb(asqrt[7] ), .dout(n22633));
  jor  g22376(.dina(n22632), .dinb(asqrt[7] ), .dout(n22634));
  jxor g22377(.dina(n21894), .dinb(n21184), .dout(n22635));
  jand g22378(.dina(n22635), .dinb(asqrt[4] ), .dout(n22636));
  jxor g22379(.dina(n22636), .dinb(n22408), .dout(n22637));
  jand g22380(.dina(n22637), .dinb(n22634), .dout(n22638));
  jor  g22381(.dina(n22638), .dinb(n22633), .dout(n22639));
  jand g22382(.dina(n22639), .dinb(asqrt[8] ), .dout(n22640));
  jor  g22383(.dina(n22639), .dinb(asqrt[8] ), .dout(n22641));
  jxor g22384(.dina(n21902), .dinb(n20468), .dout(n22642));
  jand g22385(.dina(n22642), .dinb(asqrt[4] ), .dout(n22643));
  jxor g22386(.dina(n22643), .dinb(n22412), .dout(n22644));
  jand g22387(.dina(n22644), .dinb(n22641), .dout(n22645));
  jor  g22388(.dina(n22645), .dinb(n22640), .dout(n22646));
  jand g22389(.dina(n22646), .dinb(asqrt[9] ), .dout(n22647));
  jor  g22390(.dina(n22646), .dinb(asqrt[9] ), .dout(n22648));
  jxor g22391(.dina(n21911), .dinb(n19791), .dout(n22649));
  jand g22392(.dina(n22649), .dinb(asqrt[4] ), .dout(n22650));
  jxor g22393(.dina(n22650), .dinb(n21916), .dout(n22651));
  jand g22394(.dina(n22651), .dinb(n22648), .dout(n22652));
  jor  g22395(.dina(n22652), .dinb(n22647), .dout(n22653));
  jand g22396(.dina(n22653), .dinb(asqrt[10] ), .dout(n22654));
  jor  g22397(.dina(n22653), .dinb(asqrt[10] ), .dout(n22655));
  jxor g22398(.dina(n21919), .dinb(n19096), .dout(n22656));
  jand g22399(.dina(n22656), .dinb(asqrt[4] ), .dout(n22657));
  jxor g22400(.dina(n22657), .dinb(n21924), .dout(n22658));
  jnot g22401(.din(n22658), .dout(n22659));
  jand g22402(.dina(n22659), .dinb(n22655), .dout(n22660));
  jor  g22403(.dina(n22660), .dinb(n22654), .dout(n22661));
  jand g22404(.dina(n22661), .dinb(asqrt[11] ), .dout(n22662));
  jor  g22405(.dina(n22661), .dinb(asqrt[11] ), .dout(n22663));
  jxor g22406(.dina(n21926), .dinb(n18442), .dout(n22664));
  jand g22407(.dina(n22664), .dinb(asqrt[4] ), .dout(n22665));
  jxor g22408(.dina(n22665), .dinb(n21931), .dout(n22666));
  jand g22409(.dina(n22666), .dinb(n22663), .dout(n22667));
  jor  g22410(.dina(n22667), .dinb(n22662), .dout(n22668));
  jand g22411(.dina(n22668), .dinb(asqrt[12] ), .dout(n22669));
  jor  g22412(.dina(n22668), .dinb(asqrt[12] ), .dout(n22670));
  jxor g22413(.dina(n21934), .dinb(n17769), .dout(n22671));
  jand g22414(.dina(n22671), .dinb(asqrt[4] ), .dout(n22672));
  jxor g22415(.dina(n22672), .dinb(n21939), .dout(n22673));
  jnot g22416(.din(n22673), .dout(n22674));
  jand g22417(.dina(n22674), .dinb(n22670), .dout(n22675));
  jor  g22418(.dina(n22675), .dinb(n22669), .dout(n22676));
  jand g22419(.dina(n22676), .dinb(asqrt[13] ), .dout(n22677));
  jor  g22420(.dina(n22676), .dinb(asqrt[13] ), .dout(n22678));
  jxor g22421(.dina(n21941), .dinb(n17134), .dout(n22679));
  jand g22422(.dina(n22679), .dinb(asqrt[4] ), .dout(n22680));
  jxor g22423(.dina(n22680), .dinb(n21946), .dout(n22681));
  jand g22424(.dina(n22681), .dinb(n22678), .dout(n22682));
  jor  g22425(.dina(n22682), .dinb(n22677), .dout(n22683));
  jand g22426(.dina(n22683), .dinb(asqrt[14] ), .dout(n22684));
  jor  g22427(.dina(n22683), .dinb(asqrt[14] ), .dout(n22685));
  jxor g22428(.dina(n21949), .dinb(n16489), .dout(n22686));
  jand g22429(.dina(n22686), .dinb(asqrt[4] ), .dout(n22687));
  jxor g22430(.dina(n22687), .dinb(n21954), .dout(n22688));
  jnot g22431(.din(n22688), .dout(n22689));
  jand g22432(.dina(n22689), .dinb(n22685), .dout(n22690));
  jor  g22433(.dina(n22690), .dinb(n22684), .dout(n22691));
  jand g22434(.dina(n22691), .dinb(asqrt[15] ), .dout(n22692));
  jor  g22435(.dina(n22691), .dinb(asqrt[15] ), .dout(n22693));
  jxor g22436(.dina(n21956), .dinb(n15878), .dout(n22694));
  jand g22437(.dina(n22694), .dinb(asqrt[4] ), .dout(n22695));
  jxor g22438(.dina(n22695), .dinb(n21961), .dout(n22696));
  jnot g22439(.din(n22696), .dout(n22697));
  jand g22440(.dina(n22697), .dinb(n22693), .dout(n22698));
  jor  g22441(.dina(n22698), .dinb(n22692), .dout(n22699));
  jand g22442(.dina(n22699), .dinb(asqrt[16] ), .dout(n22700));
  jor  g22443(.dina(n22699), .dinb(asqrt[16] ), .dout(n22701));
  jxor g22444(.dina(n21963), .dinb(n15260), .dout(n22702));
  jand g22445(.dina(n22702), .dinb(asqrt[4] ), .dout(n22703));
  jxor g22446(.dina(n22703), .dinb(n21968), .dout(n22704));
  jnot g22447(.din(n22704), .dout(n22705));
  jand g22448(.dina(n22705), .dinb(n22701), .dout(n22706));
  jor  g22449(.dina(n22706), .dinb(n22700), .dout(n22707));
  jand g22450(.dina(n22707), .dinb(asqrt[17] ), .dout(n22708));
  jor  g22451(.dina(n22707), .dinb(asqrt[17] ), .dout(n22709));
  jxor g22452(.dina(n21970), .dinb(n14674), .dout(n22710));
  jand g22453(.dina(n22710), .dinb(asqrt[4] ), .dout(n22711));
  jxor g22454(.dina(n22711), .dinb(n21975), .dout(n22712));
  jand g22455(.dina(n22712), .dinb(n22709), .dout(n22713));
  jor  g22456(.dina(n22713), .dinb(n22708), .dout(n22714));
  jand g22457(.dina(n22714), .dinb(asqrt[18] ), .dout(n22715));
  jor  g22458(.dina(n22714), .dinb(asqrt[18] ), .dout(n22716));
  jxor g22459(.dina(n21978), .dinb(n14078), .dout(n22717));
  jand g22460(.dina(n22717), .dinb(asqrt[4] ), .dout(n22718));
  jxor g22461(.dina(n22718), .dinb(n21983), .dout(n22719));
  jnot g22462(.din(n22719), .dout(n22720));
  jand g22463(.dina(n22720), .dinb(n22716), .dout(n22721));
  jor  g22464(.dina(n22721), .dinb(n22715), .dout(n22722));
  jand g22465(.dina(n22722), .dinb(asqrt[19] ), .dout(n22723));
  jor  g22466(.dina(n22722), .dinb(asqrt[19] ), .dout(n22724));
  jxor g22467(.dina(n21985), .dinb(n13515), .dout(n22725));
  jand g22468(.dina(n22725), .dinb(asqrt[4] ), .dout(n22726));
  jxor g22469(.dina(n22726), .dinb(n21990), .dout(n22727));
  jnot g22470(.din(n22727), .dout(n22728));
  jand g22471(.dina(n22728), .dinb(n22724), .dout(n22729));
  jor  g22472(.dina(n22729), .dinb(n22723), .dout(n22730));
  jand g22473(.dina(n22730), .dinb(asqrt[20] ), .dout(n22731));
  jor  g22474(.dina(n22730), .dinb(asqrt[20] ), .dout(n22732));
  jxor g22475(.dina(n21992), .dinb(n12947), .dout(n22733));
  jand g22476(.dina(n22733), .dinb(asqrt[4] ), .dout(n22734));
  jxor g22477(.dina(n22734), .dinb(n21997), .dout(n22735));
  jnot g22478(.din(n22735), .dout(n22736));
  jand g22479(.dina(n22736), .dinb(n22732), .dout(n22737));
  jor  g22480(.dina(n22737), .dinb(n22731), .dout(n22738));
  jand g22481(.dina(n22738), .dinb(asqrt[21] ), .dout(n22739));
  jor  g22482(.dina(n22738), .dinb(asqrt[21] ), .dout(n22740));
  jxor g22483(.dina(n21999), .dinb(n12410), .dout(n22741));
  jand g22484(.dina(n22741), .dinb(asqrt[4] ), .dout(n22742));
  jxor g22485(.dina(n22742), .dinb(n22004), .dout(n22743));
  jand g22486(.dina(n22743), .dinb(n22740), .dout(n22744));
  jor  g22487(.dina(n22744), .dinb(n22739), .dout(n22745));
  jand g22488(.dina(n22745), .dinb(asqrt[22] ), .dout(n22746));
  jor  g22489(.dina(n22745), .dinb(asqrt[22] ), .dout(n22747));
  jxor g22490(.dina(n22007), .dinb(n11858), .dout(n22748));
  jand g22491(.dina(n22748), .dinb(asqrt[4] ), .dout(n22749));
  jxor g22492(.dina(n22749), .dinb(n22012), .dout(n22750));
  jnot g22493(.din(n22750), .dout(n22751));
  jand g22494(.dina(n22751), .dinb(n22747), .dout(n22752));
  jor  g22495(.dina(n22752), .dinb(n22746), .dout(n22753));
  jand g22496(.dina(n22753), .dinb(asqrt[23] ), .dout(n22754));
  jor  g22497(.dina(n22753), .dinb(asqrt[23] ), .dout(n22755));
  jxor g22498(.dina(n22014), .dinb(n11347), .dout(n22756));
  jand g22499(.dina(n22756), .dinb(asqrt[4] ), .dout(n22757));
  jxor g22500(.dina(n22757), .dinb(n22019), .dout(n22758));
  jand g22501(.dina(n22758), .dinb(n22755), .dout(n22759));
  jor  g22502(.dina(n22759), .dinb(n22754), .dout(n22760));
  jand g22503(.dina(n22760), .dinb(asqrt[24] ), .dout(n22761));
  jor  g22504(.dina(n22760), .dinb(asqrt[24] ), .dout(n22762));
  jxor g22505(.dina(n22022), .dinb(n10824), .dout(n22763));
  jand g22506(.dina(n22763), .dinb(asqrt[4] ), .dout(n22764));
  jxor g22507(.dina(n22764), .dinb(n22027), .dout(n22765));
  jnot g22508(.din(n22765), .dout(n22766));
  jand g22509(.dina(n22766), .dinb(n22762), .dout(n22767));
  jor  g22510(.dina(n22767), .dinb(n22761), .dout(n22768));
  jand g22511(.dina(n22768), .dinb(asqrt[25] ), .dout(n22769));
  jor  g22512(.dina(n22768), .dinb(asqrt[25] ), .dout(n22770));
  jxor g22513(.dina(n22029), .dinb(n10328), .dout(n22771));
  jand g22514(.dina(n22771), .dinb(asqrt[4] ), .dout(n22772));
  jxor g22515(.dina(n22772), .dinb(n22034), .dout(n22773));
  jand g22516(.dina(n22773), .dinb(n22770), .dout(n22774));
  jor  g22517(.dina(n22774), .dinb(n22769), .dout(n22775));
  jand g22518(.dina(n22775), .dinb(asqrt[26] ), .dout(n22776));
  jor  g22519(.dina(n22775), .dinb(asqrt[26] ), .dout(n22777));
  jxor g22520(.dina(n22037), .dinb(n9832), .dout(n22778));
  jand g22521(.dina(n22778), .dinb(asqrt[4] ), .dout(n22779));
  jxor g22522(.dina(n22779), .dinb(n22042), .dout(n22780));
  jnot g22523(.din(n22780), .dout(n22781));
  jand g22524(.dina(n22781), .dinb(n22777), .dout(n22782));
  jor  g22525(.dina(n22782), .dinb(n22776), .dout(n22783));
  jand g22526(.dina(n22783), .dinb(asqrt[27] ), .dout(n22784));
  jor  g22527(.dina(n22783), .dinb(asqrt[27] ), .dout(n22785));
  jxor g22528(.dina(n22044), .dinb(n9369), .dout(n22786));
  jand g22529(.dina(n22786), .dinb(asqrt[4] ), .dout(n22787));
  jxor g22530(.dina(n22787), .dinb(n22049), .dout(n22788));
  jnot g22531(.din(n22788), .dout(n22789));
  jand g22532(.dina(n22789), .dinb(n22785), .dout(n22790));
  jor  g22533(.dina(n22790), .dinb(n22784), .dout(n22791));
  jand g22534(.dina(n22791), .dinb(asqrt[28] ), .dout(n22792));
  jor  g22535(.dina(n22791), .dinb(asqrt[28] ), .dout(n22793));
  jxor g22536(.dina(n22051), .dinb(n8890), .dout(n22794));
  jand g22537(.dina(n22794), .dinb(asqrt[4] ), .dout(n22795));
  jxor g22538(.dina(n22795), .dinb(n22056), .dout(n22796));
  jand g22539(.dina(n22796), .dinb(n22793), .dout(n22797));
  jor  g22540(.dina(n22797), .dinb(n22792), .dout(n22798));
  jand g22541(.dina(n22798), .dinb(asqrt[29] ), .dout(n22799));
  jor  g22542(.dina(n22798), .dinb(asqrt[29] ), .dout(n22800));
  jxor g22543(.dina(n22059), .dinb(n8449), .dout(n22801));
  jand g22544(.dina(n22801), .dinb(asqrt[4] ), .dout(n22802));
  jxor g22545(.dina(n22802), .dinb(n22064), .dout(n22803));
  jand g22546(.dina(n22803), .dinb(n22800), .dout(n22804));
  jor  g22547(.dina(n22804), .dinb(n22799), .dout(n22805));
  jand g22548(.dina(n22805), .dinb(asqrt[30] ), .dout(n22806));
  jor  g22549(.dina(n22805), .dinb(asqrt[30] ), .dout(n22807));
  jxor g22550(.dina(n22067), .dinb(n8003), .dout(n22808));
  jand g22551(.dina(n22808), .dinb(asqrt[4] ), .dout(n22809));
  jxor g22552(.dina(n22809), .dinb(n22072), .dout(n22810));
  jnot g22553(.din(n22810), .dout(n22811));
  jand g22554(.dina(n22811), .dinb(n22807), .dout(n22812));
  jor  g22555(.dina(n22812), .dinb(n22806), .dout(n22813));
  jand g22556(.dina(n22813), .dinb(asqrt[31] ), .dout(n22814));
  jor  g22557(.dina(n22813), .dinb(asqrt[31] ), .dout(n22815));
  jxor g22558(.dina(n22074), .dinb(n7581), .dout(n22816));
  jand g22559(.dina(n22816), .dinb(asqrt[4] ), .dout(n22817));
  jxor g22560(.dina(n22817), .dinb(n22079), .dout(n22818));
  jand g22561(.dina(n22818), .dinb(n22815), .dout(n22819));
  jor  g22562(.dina(n22819), .dinb(n22814), .dout(n22820));
  jand g22563(.dina(n22820), .dinb(asqrt[32] ), .dout(n22821));
  jor  g22564(.dina(n22820), .dinb(asqrt[32] ), .dout(n22822));
  jxor g22565(.dina(n22082), .dinb(n7154), .dout(n22823));
  jand g22566(.dina(n22823), .dinb(asqrt[4] ), .dout(n22824));
  jxor g22567(.dina(n22824), .dinb(n22087), .dout(n22825));
  jnot g22568(.din(n22825), .dout(n22826));
  jand g22569(.dina(n22826), .dinb(n22822), .dout(n22827));
  jor  g22570(.dina(n22827), .dinb(n22821), .dout(n22828));
  jand g22571(.dina(n22828), .dinb(asqrt[33] ), .dout(n22829));
  jor  g22572(.dina(n22828), .dinb(asqrt[33] ), .dout(n22830));
  jxor g22573(.dina(n22089), .dinb(n6758), .dout(n22831));
  jand g22574(.dina(n22831), .dinb(asqrt[4] ), .dout(n22832));
  jxor g22575(.dina(n22832), .dinb(n22094), .dout(n22833));
  jand g22576(.dina(n22833), .dinb(n22830), .dout(n22834));
  jor  g22577(.dina(n22834), .dinb(n22829), .dout(n22835));
  jand g22578(.dina(n22835), .dinb(asqrt[34] ), .dout(n22836));
  jor  g22579(.dina(n22835), .dinb(asqrt[34] ), .dout(n22837));
  jxor g22580(.dina(n22097), .dinb(n6357), .dout(n22838));
  jand g22581(.dina(n22838), .dinb(asqrt[4] ), .dout(n22839));
  jxor g22582(.dina(n22839), .dinb(n22102), .dout(n22840));
  jnot g22583(.din(n22840), .dout(n22841));
  jand g22584(.dina(n22841), .dinb(n22837), .dout(n22842));
  jor  g22585(.dina(n22842), .dinb(n22836), .dout(n22843));
  jand g22586(.dina(n22843), .dinb(asqrt[35] ), .dout(n22844));
  jor  g22587(.dina(n22843), .dinb(asqrt[35] ), .dout(n22845));
  jxor g22588(.dina(n22104), .dinb(n5989), .dout(n22846));
  jand g22589(.dina(n22846), .dinb(asqrt[4] ), .dout(n22847));
  jxor g22590(.dina(n22847), .dinb(n22109), .dout(n22848));
  jnot g22591(.din(n22848), .dout(n22849));
  jand g22592(.dina(n22849), .dinb(n22845), .dout(n22850));
  jor  g22593(.dina(n22850), .dinb(n22844), .dout(n22851));
  jand g22594(.dina(n22851), .dinb(asqrt[36] ), .dout(n22852));
  jor  g22595(.dina(n22851), .dinb(asqrt[36] ), .dout(n22853));
  jxor g22596(.dina(n22111), .dinb(n5606), .dout(n22854));
  jand g22597(.dina(n22854), .dinb(asqrt[4] ), .dout(n22855));
  jxor g22598(.dina(n22855), .dinb(n22116), .dout(n22856));
  jnot g22599(.din(n22856), .dout(n22857));
  jand g22600(.dina(n22857), .dinb(n22853), .dout(n22858));
  jor  g22601(.dina(n22858), .dinb(n22852), .dout(n22859));
  jand g22602(.dina(n22859), .dinb(asqrt[37] ), .dout(n22860));
  jor  g22603(.dina(n22859), .dinb(asqrt[37] ), .dout(n22861));
  jxor g22604(.dina(n22118), .dinb(n5259), .dout(n22862));
  jand g22605(.dina(n22862), .dinb(asqrt[4] ), .dout(n22863));
  jxor g22606(.dina(n22863), .dinb(n22123), .dout(n22864));
  jand g22607(.dina(n22864), .dinb(n22861), .dout(n22865));
  jor  g22608(.dina(n22865), .dinb(n22860), .dout(n22866));
  jand g22609(.dina(n22866), .dinb(asqrt[38] ), .dout(n22867));
  jor  g22610(.dina(n22866), .dinb(asqrt[38] ), .dout(n22868));
  jxor g22611(.dina(n22126), .dinb(n4902), .dout(n22869));
  jand g22612(.dina(n22869), .dinb(asqrt[4] ), .dout(n22870));
  jxor g22613(.dina(n22870), .dinb(n22131), .dout(n22871));
  jnot g22614(.din(n22871), .dout(n22872));
  jand g22615(.dina(n22872), .dinb(n22868), .dout(n22873));
  jor  g22616(.dina(n22873), .dinb(n22867), .dout(n22874));
  jand g22617(.dina(n22874), .dinb(asqrt[39] ), .dout(n22875));
  jor  g22618(.dina(n22874), .dinb(asqrt[39] ), .dout(n22876));
  jxor g22619(.dina(n22133), .dinb(n4582), .dout(n22877));
  jand g22620(.dina(n22877), .dinb(asqrt[4] ), .dout(n22878));
  jxor g22621(.dina(n22878), .dinb(n22138), .dout(n22879));
  jand g22622(.dina(n22879), .dinb(n22876), .dout(n22880));
  jor  g22623(.dina(n22880), .dinb(n22875), .dout(n22881));
  jand g22624(.dina(n22881), .dinb(asqrt[40] ), .dout(n22882));
  jor  g22625(.dina(n22881), .dinb(asqrt[40] ), .dout(n22883));
  jxor g22626(.dina(n22141), .dinb(n4249), .dout(n22884));
  jand g22627(.dina(n22884), .dinb(asqrt[4] ), .dout(n22885));
  jxor g22628(.dina(n22885), .dinb(n22146), .dout(n22886));
  jnot g22629(.din(n22886), .dout(n22887));
  jand g22630(.dina(n22887), .dinb(n22883), .dout(n22888));
  jor  g22631(.dina(n22888), .dinb(n22882), .dout(n22889));
  jand g22632(.dina(n22889), .dinb(asqrt[41] ), .dout(n22890));
  jor  g22633(.dina(n22889), .dinb(asqrt[41] ), .dout(n22891));
  jxor g22634(.dina(n22148), .dinb(n3955), .dout(n22892));
  jand g22635(.dina(n22892), .dinb(asqrt[4] ), .dout(n22893));
  jxor g22636(.dina(n22893), .dinb(n22153), .dout(n22894));
  jand g22637(.dina(n22894), .dinb(n22891), .dout(n22895));
  jor  g22638(.dina(n22895), .dinb(n22890), .dout(n22896));
  jand g22639(.dina(n22896), .dinb(asqrt[42] ), .dout(n22897));
  jor  g22640(.dina(n22896), .dinb(asqrt[42] ), .dout(n22898));
  jxor g22641(.dina(n22156), .dinb(n3642), .dout(n22899));
  jand g22642(.dina(n22899), .dinb(asqrt[4] ), .dout(n22900));
  jxor g22643(.dina(n22900), .dinb(n22161), .dout(n22901));
  jnot g22644(.din(n22901), .dout(n22902));
  jand g22645(.dina(n22902), .dinb(n22898), .dout(n22903));
  jor  g22646(.dina(n22903), .dinb(n22897), .dout(n22904));
  jand g22647(.dina(n22904), .dinb(asqrt[43] ), .dout(n22905));
  jor  g22648(.dina(n22904), .dinb(asqrt[43] ), .dout(n22906));
  jxor g22649(.dina(n22163), .dinb(n3368), .dout(n22907));
  jand g22650(.dina(n22907), .dinb(asqrt[4] ), .dout(n22908));
  jxor g22651(.dina(n22908), .dinb(n22168), .dout(n22909));
  jand g22652(.dina(n22909), .dinb(n22906), .dout(n22910));
  jor  g22653(.dina(n22910), .dinb(n22905), .dout(n22911));
  jand g22654(.dina(n22911), .dinb(asqrt[44] ), .dout(n22912));
  jor  g22655(.dina(n22911), .dinb(asqrt[44] ), .dout(n22913));
  jxor g22656(.dina(n22171), .dinb(n3089), .dout(n22914));
  jand g22657(.dina(n22914), .dinb(asqrt[4] ), .dout(n22915));
  jxor g22658(.dina(n22915), .dinb(n22176), .dout(n22916));
  jnot g22659(.din(n22916), .dout(n22917));
  jand g22660(.dina(n22917), .dinb(n22913), .dout(n22918));
  jor  g22661(.dina(n22918), .dinb(n22912), .dout(n22919));
  jand g22662(.dina(n22919), .dinb(asqrt[45] ), .dout(n22920));
  jor  g22663(.dina(n22919), .dinb(asqrt[45] ), .dout(n22921));
  jxor g22664(.dina(n22178), .dinb(n2833), .dout(n22922));
  jand g22665(.dina(n22922), .dinb(asqrt[4] ), .dout(n22923));
  jxor g22666(.dina(n22923), .dinb(n22183), .dout(n22924));
  jnot g22667(.din(n22924), .dout(n22925));
  jand g22668(.dina(n22925), .dinb(n22921), .dout(n22926));
  jor  g22669(.dina(n22926), .dinb(n22920), .dout(n22927));
  jand g22670(.dina(n22927), .dinb(asqrt[46] ), .dout(n22928));
  jor  g22671(.dina(n22927), .dinb(asqrt[46] ), .dout(n22929));
  jxor g22672(.dina(n22185), .dinb(n2572), .dout(n22930));
  jand g22673(.dina(n22930), .dinb(asqrt[4] ), .dout(n22931));
  jxor g22674(.dina(n22931), .dinb(n22190), .dout(n22932));
  jnot g22675(.din(n22932), .dout(n22933));
  jand g22676(.dina(n22933), .dinb(n22929), .dout(n22934));
  jor  g22677(.dina(n22934), .dinb(n22928), .dout(n22935));
  jand g22678(.dina(n22935), .dinb(asqrt[47] ), .dout(n22936));
  jor  g22679(.dina(n22935), .dinb(asqrt[47] ), .dout(n22937));
  jxor g22680(.dina(n22192), .dinb(n2345), .dout(n22938));
  jand g22681(.dina(n22938), .dinb(asqrt[4] ), .dout(n22939));
  jxor g22682(.dina(n22939), .dinb(n22197), .dout(n22940));
  jand g22683(.dina(n22940), .dinb(n22937), .dout(n22941));
  jor  g22684(.dina(n22941), .dinb(n22936), .dout(n22942));
  jand g22685(.dina(n22942), .dinb(asqrt[48] ), .dout(n22943));
  jor  g22686(.dina(n22942), .dinb(asqrt[48] ), .dout(n22944));
  jxor g22687(.dina(n22200), .dinb(n2108), .dout(n22945));
  jand g22688(.dina(n22945), .dinb(asqrt[4] ), .dout(n22946));
  jxor g22689(.dina(n22946), .dinb(n22205), .dout(n22947));
  jnot g22690(.din(n22947), .dout(n22948));
  jand g22691(.dina(n22948), .dinb(n22944), .dout(n22949));
  jor  g22692(.dina(n22949), .dinb(n22943), .dout(n22950));
  jand g22693(.dina(n22950), .dinb(asqrt[49] ), .dout(n22951));
  jor  g22694(.dina(n22950), .dinb(asqrt[49] ), .dout(n22952));
  jxor g22695(.dina(n22207), .dinb(n1912), .dout(n22953));
  jand g22696(.dina(n22953), .dinb(asqrt[4] ), .dout(n22954));
  jxor g22697(.dina(n22954), .dinb(n22212), .dout(n22955));
  jnot g22698(.din(n22955), .dout(n22956));
  jand g22699(.dina(n22956), .dinb(n22952), .dout(n22957));
  jor  g22700(.dina(n22957), .dinb(n22951), .dout(n22958));
  jand g22701(.dina(n22958), .dinb(asqrt[50] ), .dout(n22959));
  jor  g22702(.dina(n22958), .dinb(asqrt[50] ), .dout(n22960));
  jxor g22703(.dina(n22214), .dinb(n1699), .dout(n22961));
  jand g22704(.dina(n22961), .dinb(asqrt[4] ), .dout(n22962));
  jxor g22705(.dina(n22962), .dinb(n22219), .dout(n22963));
  jnot g22706(.din(n22963), .dout(n22964));
  jand g22707(.dina(n22964), .dinb(n22960), .dout(n22965));
  jor  g22708(.dina(n22965), .dinb(n22959), .dout(n22966));
  jand g22709(.dina(n22966), .dinb(asqrt[51] ), .dout(n22967));
  jor  g22710(.dina(n22966), .dinb(asqrt[51] ), .dout(n22968));
  jxor g22711(.dina(n22221), .dinb(n1516), .dout(n22969));
  jand g22712(.dina(n22969), .dinb(asqrt[4] ), .dout(n22970));
  jxor g22713(.dina(n22970), .dinb(n22226), .dout(n22971));
  jnot g22714(.din(n22971), .dout(n22972));
  jand g22715(.dina(n22972), .dinb(n22968), .dout(n22973));
  jor  g22716(.dina(n22973), .dinb(n22967), .dout(n22974));
  jand g22717(.dina(n22974), .dinb(asqrt[52] ), .dout(n22975));
  jor  g22718(.dina(n22974), .dinb(asqrt[52] ), .dout(n22976));
  jxor g22719(.dina(n22228), .dinb(n1332), .dout(n22977));
  jand g22720(.dina(n22977), .dinb(asqrt[4] ), .dout(n22978));
  jxor g22721(.dina(n22978), .dinb(n22233), .dout(n22979));
  jnot g22722(.din(n22979), .dout(n22980));
  jand g22723(.dina(n22980), .dinb(n22976), .dout(n22981));
  jor  g22724(.dina(n22981), .dinb(n22975), .dout(n22982));
  jand g22725(.dina(n22982), .dinb(asqrt[53] ), .dout(n22983));
  jor  g22726(.dina(n22982), .dinb(asqrt[53] ), .dout(n22984));
  jxor g22727(.dina(n22235), .dinb(n1173), .dout(n22985));
  jand g22728(.dina(n22985), .dinb(asqrt[4] ), .dout(n22986));
  jxor g22729(.dina(n22986), .dinb(n22240), .dout(n22987));
  jand g22730(.dina(n22987), .dinb(n22984), .dout(n22988));
  jor  g22731(.dina(n22988), .dinb(n22983), .dout(n22989));
  jand g22732(.dina(n22989), .dinb(asqrt[54] ), .dout(n22990));
  jor  g22733(.dina(n22989), .dinb(asqrt[54] ), .dout(n22991));
  jxor g22734(.dina(n22243), .dinb(n1008), .dout(n22992));
  jand g22735(.dina(n22992), .dinb(asqrt[4] ), .dout(n22993));
  jxor g22736(.dina(n22993), .dinb(n22248), .dout(n22994));
  jnot g22737(.din(n22994), .dout(n22995));
  jand g22738(.dina(n22995), .dinb(n22991), .dout(n22996));
  jor  g22739(.dina(n22996), .dinb(n22990), .dout(n22997));
  jand g22740(.dina(n22997), .dinb(asqrt[55] ), .dout(n22998));
  jor  g22741(.dina(n22997), .dinb(asqrt[55] ), .dout(n22999));
  jxor g22742(.dina(n22250), .dinb(n884), .dout(n23000));
  jand g22743(.dina(n23000), .dinb(asqrt[4] ), .dout(n23001));
  jxor g22744(.dina(n23001), .dinb(n22255), .dout(n23002));
  jand g22745(.dina(n23002), .dinb(n22999), .dout(n23003));
  jor  g22746(.dina(n23003), .dinb(n22998), .dout(n23004));
  jand g22747(.dina(n23004), .dinb(asqrt[56] ), .dout(n23005));
  jor  g22748(.dina(n23004), .dinb(asqrt[56] ), .dout(n23006));
  jxor g22749(.dina(n22258), .dinb(n743), .dout(n23007));
  jand g22750(.dina(n23007), .dinb(asqrt[4] ), .dout(n23008));
  jxor g22751(.dina(n23008), .dinb(n22263), .dout(n23009));
  jnot g22752(.din(n23009), .dout(n23010));
  jand g22753(.dina(n23010), .dinb(n23006), .dout(n23011));
  jor  g22754(.dina(n23011), .dinb(n23005), .dout(n23012));
  jand g22755(.dina(n23012), .dinb(asqrt[57] ), .dout(n23013));
  jor  g22756(.dina(n23012), .dinb(asqrt[57] ), .dout(n23014));
  jxor g22757(.dina(n22265), .dinb(n635), .dout(n23015));
  jand g22758(.dina(n23015), .dinb(asqrt[4] ), .dout(n23016));
  jxor g22759(.dina(n23016), .dinb(n22270), .dout(n23017));
  jnot g22760(.din(n23017), .dout(n23018));
  jand g22761(.dina(n23018), .dinb(n23014), .dout(n23019));
  jor  g22762(.dina(n23019), .dinb(n23013), .dout(n23020));
  jand g22763(.dina(n23020), .dinb(asqrt[58] ), .dout(n23021));
  jor  g22764(.dina(n23020), .dinb(asqrt[58] ), .dout(n23022));
  jxor g22765(.dina(n22272), .dinb(n515), .dout(n23023));
  jand g22766(.dina(n23023), .dinb(asqrt[4] ), .dout(n23024));
  jxor g22767(.dina(n23024), .dinb(n22277), .dout(n23025));
  jand g22768(.dina(n23025), .dinb(n23022), .dout(n23026));
  jor  g22769(.dina(n23026), .dinb(n23021), .dout(n23027));
  jand g22770(.dina(n23027), .dinb(asqrt[59] ), .dout(n23028));
  jor  g22771(.dina(n23027), .dinb(asqrt[59] ), .dout(n23029));
  jxor g22772(.dina(n22280), .dinb(n443), .dout(n23030));
  jand g22773(.dina(n23030), .dinb(asqrt[4] ), .dout(n23031));
  jxor g22774(.dina(n23031), .dinb(n22285), .dout(n23032));
  jand g22775(.dina(n23032), .dinb(n23029), .dout(n23033));
  jor  g22776(.dina(n23033), .dinb(n23028), .dout(n23034));
  jand g22777(.dina(n23034), .dinb(asqrt[60] ), .dout(n23035));
  jor  g22778(.dina(n23034), .dinb(asqrt[60] ), .dout(n23036));
  jxor g22779(.dina(n22288), .dinb(n352), .dout(n23037));
  jand g22780(.dina(n23037), .dinb(asqrt[4] ), .dout(n23038));
  jxor g22781(.dina(n23038), .dinb(n22293), .dout(n23039));
  jnot g22782(.din(n23039), .dout(n23040));
  jand g22783(.dina(n23040), .dinb(n23036), .dout(n23041));
  jor  g22784(.dina(n23041), .dinb(n23035), .dout(n23042));
  jand g22785(.dina(n23042), .dinb(asqrt[61] ), .dout(n23043));
  jor  g22786(.dina(n23042), .dinb(asqrt[61] ), .dout(n23044));
  jxor g22787(.dina(n22295), .dinb(n294), .dout(n23045));
  jand g22788(.dina(n23045), .dinb(asqrt[4] ), .dout(n23046));
  jxor g22789(.dina(n23046), .dinb(n22300), .dout(n23047));
  jnot g22790(.din(n23047), .dout(n23048));
  jand g22791(.dina(n23048), .dinb(n23044), .dout(n23049));
  jor  g22792(.dina(n23049), .dinb(n23043), .dout(n23050));
  jand g22793(.dina(n23050), .dinb(asqrt[62] ), .dout(n23051));
  jor  g22794(.dina(n23050), .dinb(asqrt[62] ), .dout(n23052));
  jxor g22795(.dina(n22302), .dinb(n239), .dout(n23053));
  jand g22796(.dina(n23053), .dinb(asqrt[4] ), .dout(n23054));
  jxor g22797(.dina(n23054), .dinb(n22307), .dout(n23055));
  jnot g22798(.din(n23055), .dout(n23056));
  jand g22799(.dina(n23056), .dinb(n23052), .dout(n23057));
  jor  g22800(.dina(n23057), .dinb(n23051), .dout(n23058));
  jxor g22801(.dina(n22309), .dinb(n221), .dout(n23059));
  jand g22802(.dina(n23059), .dinb(asqrt[4] ), .dout(n23060));
  jxor g22803(.dina(n23060), .dinb(n22315), .dout(n23061));
  jnot g22804(.din(n23061), .dout(n23062));
  jor  g22805(.dina(n23062), .dinb(n23058), .dout(n23063));
  jnot g22806(.din(n23063), .dout(n23064));
  jand g22807(.dina(n22332), .dinb(n22615), .dout(n23065));
  jnot g22808(.din(n23051), .dout(n23066));
  jnot g22809(.din(n23043), .dout(n23067));
  jnot g22810(.din(n23035), .dout(n23068));
  jnot g22811(.din(n23028), .dout(n23069));
  jnot g22812(.din(n23021), .dout(n23070));
  jnot g22813(.din(n23013), .dout(n23071));
  jnot g22814(.din(n23005), .dout(n23072));
  jnot g22815(.din(n22998), .dout(n23073));
  jnot g22816(.din(n22990), .dout(n23074));
  jnot g22817(.din(n22983), .dout(n23075));
  jnot g22818(.din(n22975), .dout(n23076));
  jnot g22819(.din(n22967), .dout(n23077));
  jnot g22820(.din(n22959), .dout(n23078));
  jnot g22821(.din(n22951), .dout(n23079));
  jnot g22822(.din(n22943), .dout(n23080));
  jnot g22823(.din(n22936), .dout(n23081));
  jnot g22824(.din(n22928), .dout(n23082));
  jnot g22825(.din(n22920), .dout(n23083));
  jnot g22826(.din(n22912), .dout(n23084));
  jnot g22827(.din(n22905), .dout(n23085));
  jnot g22828(.din(n22897), .dout(n23086));
  jnot g22829(.din(n22890), .dout(n23087));
  jnot g22830(.din(n22882), .dout(n23088));
  jnot g22831(.din(n22875), .dout(n23089));
  jnot g22832(.din(n22867), .dout(n23090));
  jnot g22833(.din(n22860), .dout(n23091));
  jnot g22834(.din(n22852), .dout(n23092));
  jnot g22835(.din(n22844), .dout(n23093));
  jnot g22836(.din(n22836), .dout(n23094));
  jnot g22837(.din(n22829), .dout(n23095));
  jnot g22838(.din(n22821), .dout(n23096));
  jnot g22839(.din(n22814), .dout(n23097));
  jnot g22840(.din(n22806), .dout(n23098));
  jnot g22841(.din(n22799), .dout(n23099));
  jnot g22842(.din(n22792), .dout(n23100));
  jnot g22843(.din(n22784), .dout(n23101));
  jnot g22844(.din(n22776), .dout(n23102));
  jnot g22845(.din(n22769), .dout(n23103));
  jnot g22846(.din(n22761), .dout(n23104));
  jnot g22847(.din(n22754), .dout(n23105));
  jnot g22848(.din(n22746), .dout(n23106));
  jnot g22849(.din(n22739), .dout(n23107));
  jnot g22850(.din(n22731), .dout(n23108));
  jnot g22851(.din(n22723), .dout(n23109));
  jnot g22852(.din(n22715), .dout(n23110));
  jnot g22853(.din(n22708), .dout(n23111));
  jnot g22854(.din(n22700), .dout(n23112));
  jnot g22855(.din(n22692), .dout(n23113));
  jnot g22856(.din(n22684), .dout(n23114));
  jnot g22857(.din(n22677), .dout(n23115));
  jnot g22858(.din(n22669), .dout(n23116));
  jnot g22859(.din(n22662), .dout(n23117));
  jnot g22860(.din(n22654), .dout(n23118));
  jnot g22861(.din(n22647), .dout(n23119));
  jnot g22862(.din(n22640), .dout(n23120));
  jnot g22863(.din(n22633), .dout(n23121));
  jnot g22864(.din(n22625), .dout(n23122));
  jnot g22865(.din(n22340), .dout(n23123));
  jnot g22866(.din(n22337), .dout(n23124));
  jor  g22867(.dina(n22620), .dinb(n21889), .dout(n23125));
  jand g22868(.dina(n23125), .dinb(n23124), .dout(n23126));
  jand g22869(.dina(n23126), .dinb(n21887), .dout(n23127));
  jor  g22870(.dina(n22620), .dinb(a[8] ), .dout(n23128));
  jand g22871(.dina(n23128), .dinb(a[9] ), .dout(n23129));
  jand g22872(.dina(asqrt[4] ), .dinb(n21891), .dout(n23130));
  jor  g22873(.dina(n23130), .dinb(n23129), .dout(n23131));
  jor  g22874(.dina(n23131), .dinb(n23127), .dout(n23132));
  jand g22875(.dina(n23132), .dinb(n23123), .dout(n23133));
  jand g22876(.dina(n23133), .dinb(n21184), .dout(n23134));
  jor  g22877(.dina(n22629), .dinb(n23134), .dout(n23135));
  jand g22878(.dina(n23135), .dinb(n23122), .dout(n23136));
  jand g22879(.dina(n23136), .dinb(n20468), .dout(n23137));
  jnot g22880(.din(n22637), .dout(n23138));
  jor  g22881(.dina(n23138), .dinb(n23137), .dout(n23139));
  jand g22882(.dina(n23139), .dinb(n23121), .dout(n23140));
  jand g22883(.dina(n23140), .dinb(n19791), .dout(n23141));
  jnot g22884(.din(n22644), .dout(n23142));
  jor  g22885(.dina(n23142), .dinb(n23141), .dout(n23143));
  jand g22886(.dina(n23143), .dinb(n23120), .dout(n23144));
  jand g22887(.dina(n23144), .dinb(n19096), .dout(n23145));
  jnot g22888(.din(n22651), .dout(n23146));
  jor  g22889(.dina(n23146), .dinb(n23145), .dout(n23147));
  jand g22890(.dina(n23147), .dinb(n23119), .dout(n23148));
  jand g22891(.dina(n23148), .dinb(n18442), .dout(n23149));
  jor  g22892(.dina(n22658), .dinb(n23149), .dout(n23150));
  jand g22893(.dina(n23150), .dinb(n23118), .dout(n23151));
  jand g22894(.dina(n23151), .dinb(n17769), .dout(n23152));
  jnot g22895(.din(n22666), .dout(n23153));
  jor  g22896(.dina(n23153), .dinb(n23152), .dout(n23154));
  jand g22897(.dina(n23154), .dinb(n23117), .dout(n23155));
  jand g22898(.dina(n23155), .dinb(n17134), .dout(n23156));
  jor  g22899(.dina(n22673), .dinb(n23156), .dout(n23157));
  jand g22900(.dina(n23157), .dinb(n23116), .dout(n23158));
  jand g22901(.dina(n23158), .dinb(n16489), .dout(n23159));
  jnot g22902(.din(n22681), .dout(n23160));
  jor  g22903(.dina(n23160), .dinb(n23159), .dout(n23161));
  jand g22904(.dina(n23161), .dinb(n23115), .dout(n23162));
  jand g22905(.dina(n23162), .dinb(n15878), .dout(n23163));
  jor  g22906(.dina(n22688), .dinb(n23163), .dout(n23164));
  jand g22907(.dina(n23164), .dinb(n23114), .dout(n23165));
  jand g22908(.dina(n23165), .dinb(n15260), .dout(n23166));
  jor  g22909(.dina(n22696), .dinb(n23166), .dout(n23167));
  jand g22910(.dina(n23167), .dinb(n23113), .dout(n23168));
  jand g22911(.dina(n23168), .dinb(n14674), .dout(n23169));
  jor  g22912(.dina(n22704), .dinb(n23169), .dout(n23170));
  jand g22913(.dina(n23170), .dinb(n23112), .dout(n23171));
  jand g22914(.dina(n23171), .dinb(n14078), .dout(n23172));
  jnot g22915(.din(n22712), .dout(n23173));
  jor  g22916(.dina(n23173), .dinb(n23172), .dout(n23174));
  jand g22917(.dina(n23174), .dinb(n23111), .dout(n23175));
  jand g22918(.dina(n23175), .dinb(n13515), .dout(n23176));
  jor  g22919(.dina(n22719), .dinb(n23176), .dout(n23177));
  jand g22920(.dina(n23177), .dinb(n23110), .dout(n23178));
  jand g22921(.dina(n23178), .dinb(n12947), .dout(n23179));
  jor  g22922(.dina(n22727), .dinb(n23179), .dout(n23180));
  jand g22923(.dina(n23180), .dinb(n23109), .dout(n23181));
  jand g22924(.dina(n23181), .dinb(n12410), .dout(n23182));
  jor  g22925(.dina(n22735), .dinb(n23182), .dout(n23183));
  jand g22926(.dina(n23183), .dinb(n23108), .dout(n23184));
  jand g22927(.dina(n23184), .dinb(n11858), .dout(n23185));
  jnot g22928(.din(n22743), .dout(n23186));
  jor  g22929(.dina(n23186), .dinb(n23185), .dout(n23187));
  jand g22930(.dina(n23187), .dinb(n23107), .dout(n23188));
  jand g22931(.dina(n23188), .dinb(n11347), .dout(n23189));
  jor  g22932(.dina(n22750), .dinb(n23189), .dout(n23190));
  jand g22933(.dina(n23190), .dinb(n23106), .dout(n23191));
  jand g22934(.dina(n23191), .dinb(n10824), .dout(n23192));
  jnot g22935(.din(n22758), .dout(n23193));
  jor  g22936(.dina(n23193), .dinb(n23192), .dout(n23194));
  jand g22937(.dina(n23194), .dinb(n23105), .dout(n23195));
  jand g22938(.dina(n23195), .dinb(n10328), .dout(n23196));
  jor  g22939(.dina(n22765), .dinb(n23196), .dout(n23197));
  jand g22940(.dina(n23197), .dinb(n23104), .dout(n23198));
  jand g22941(.dina(n23198), .dinb(n9832), .dout(n23199));
  jnot g22942(.din(n22773), .dout(n23200));
  jor  g22943(.dina(n23200), .dinb(n23199), .dout(n23201));
  jand g22944(.dina(n23201), .dinb(n23103), .dout(n23202));
  jand g22945(.dina(n23202), .dinb(n9369), .dout(n23203));
  jor  g22946(.dina(n22780), .dinb(n23203), .dout(n23204));
  jand g22947(.dina(n23204), .dinb(n23102), .dout(n23205));
  jand g22948(.dina(n23205), .dinb(n8890), .dout(n23206));
  jor  g22949(.dina(n22788), .dinb(n23206), .dout(n23207));
  jand g22950(.dina(n23207), .dinb(n23101), .dout(n23208));
  jand g22951(.dina(n23208), .dinb(n8449), .dout(n23209));
  jnot g22952(.din(n22796), .dout(n23210));
  jor  g22953(.dina(n23210), .dinb(n23209), .dout(n23211));
  jand g22954(.dina(n23211), .dinb(n23100), .dout(n23212));
  jand g22955(.dina(n23212), .dinb(n8003), .dout(n23213));
  jnot g22956(.din(n22803), .dout(n23214));
  jor  g22957(.dina(n23214), .dinb(n23213), .dout(n23215));
  jand g22958(.dina(n23215), .dinb(n23099), .dout(n23216));
  jand g22959(.dina(n23216), .dinb(n7581), .dout(n23217));
  jor  g22960(.dina(n22810), .dinb(n23217), .dout(n23218));
  jand g22961(.dina(n23218), .dinb(n23098), .dout(n23219));
  jand g22962(.dina(n23219), .dinb(n7154), .dout(n23220));
  jnot g22963(.din(n22818), .dout(n23221));
  jor  g22964(.dina(n23221), .dinb(n23220), .dout(n23222));
  jand g22965(.dina(n23222), .dinb(n23097), .dout(n23223));
  jand g22966(.dina(n23223), .dinb(n6758), .dout(n23224));
  jor  g22967(.dina(n22825), .dinb(n23224), .dout(n23225));
  jand g22968(.dina(n23225), .dinb(n23096), .dout(n23226));
  jand g22969(.dina(n23226), .dinb(n6357), .dout(n23227));
  jnot g22970(.din(n22833), .dout(n23228));
  jor  g22971(.dina(n23228), .dinb(n23227), .dout(n23229));
  jand g22972(.dina(n23229), .dinb(n23095), .dout(n23230));
  jand g22973(.dina(n23230), .dinb(n5989), .dout(n23231));
  jor  g22974(.dina(n22840), .dinb(n23231), .dout(n23232));
  jand g22975(.dina(n23232), .dinb(n23094), .dout(n23233));
  jand g22976(.dina(n23233), .dinb(n5606), .dout(n23234));
  jor  g22977(.dina(n22848), .dinb(n23234), .dout(n23235));
  jand g22978(.dina(n23235), .dinb(n23093), .dout(n23236));
  jand g22979(.dina(n23236), .dinb(n5259), .dout(n23237));
  jor  g22980(.dina(n22856), .dinb(n23237), .dout(n23238));
  jand g22981(.dina(n23238), .dinb(n23092), .dout(n23239));
  jand g22982(.dina(n23239), .dinb(n4902), .dout(n23240));
  jnot g22983(.din(n22864), .dout(n23241));
  jor  g22984(.dina(n23241), .dinb(n23240), .dout(n23242));
  jand g22985(.dina(n23242), .dinb(n23091), .dout(n23243));
  jand g22986(.dina(n23243), .dinb(n4582), .dout(n23244));
  jor  g22987(.dina(n22871), .dinb(n23244), .dout(n23245));
  jand g22988(.dina(n23245), .dinb(n23090), .dout(n23246));
  jand g22989(.dina(n23246), .dinb(n4249), .dout(n23247));
  jnot g22990(.din(n22879), .dout(n23248));
  jor  g22991(.dina(n23248), .dinb(n23247), .dout(n23249));
  jand g22992(.dina(n23249), .dinb(n23089), .dout(n23250));
  jand g22993(.dina(n23250), .dinb(n3955), .dout(n23251));
  jor  g22994(.dina(n22886), .dinb(n23251), .dout(n23252));
  jand g22995(.dina(n23252), .dinb(n23088), .dout(n23253));
  jand g22996(.dina(n23253), .dinb(n3642), .dout(n23254));
  jnot g22997(.din(n22894), .dout(n23255));
  jor  g22998(.dina(n23255), .dinb(n23254), .dout(n23256));
  jand g22999(.dina(n23256), .dinb(n23087), .dout(n23257));
  jand g23000(.dina(n23257), .dinb(n3368), .dout(n23258));
  jor  g23001(.dina(n22901), .dinb(n23258), .dout(n23259));
  jand g23002(.dina(n23259), .dinb(n23086), .dout(n23260));
  jand g23003(.dina(n23260), .dinb(n3089), .dout(n23261));
  jnot g23004(.din(n22909), .dout(n23262));
  jor  g23005(.dina(n23262), .dinb(n23261), .dout(n23263));
  jand g23006(.dina(n23263), .dinb(n23085), .dout(n23264));
  jand g23007(.dina(n23264), .dinb(n2833), .dout(n23265));
  jor  g23008(.dina(n22916), .dinb(n23265), .dout(n23266));
  jand g23009(.dina(n23266), .dinb(n23084), .dout(n23267));
  jand g23010(.dina(n23267), .dinb(n2572), .dout(n23268));
  jor  g23011(.dina(n22924), .dinb(n23268), .dout(n23269));
  jand g23012(.dina(n23269), .dinb(n23083), .dout(n23270));
  jand g23013(.dina(n23270), .dinb(n2345), .dout(n23271));
  jor  g23014(.dina(n22932), .dinb(n23271), .dout(n23272));
  jand g23015(.dina(n23272), .dinb(n23082), .dout(n23273));
  jand g23016(.dina(n23273), .dinb(n2108), .dout(n23274));
  jnot g23017(.din(n22940), .dout(n23275));
  jor  g23018(.dina(n23275), .dinb(n23274), .dout(n23276));
  jand g23019(.dina(n23276), .dinb(n23081), .dout(n23277));
  jand g23020(.dina(n23277), .dinb(n1912), .dout(n23278));
  jor  g23021(.dina(n22947), .dinb(n23278), .dout(n23279));
  jand g23022(.dina(n23279), .dinb(n23080), .dout(n23280));
  jand g23023(.dina(n23280), .dinb(n1699), .dout(n23281));
  jor  g23024(.dina(n22955), .dinb(n23281), .dout(n23282));
  jand g23025(.dina(n23282), .dinb(n23079), .dout(n23283));
  jand g23026(.dina(n23283), .dinb(n1516), .dout(n23284));
  jor  g23027(.dina(n22963), .dinb(n23284), .dout(n23285));
  jand g23028(.dina(n23285), .dinb(n23078), .dout(n23286));
  jand g23029(.dina(n23286), .dinb(n1332), .dout(n23287));
  jor  g23030(.dina(n22971), .dinb(n23287), .dout(n23288));
  jand g23031(.dina(n23288), .dinb(n23077), .dout(n23289));
  jand g23032(.dina(n23289), .dinb(n1173), .dout(n23290));
  jor  g23033(.dina(n22979), .dinb(n23290), .dout(n23291));
  jand g23034(.dina(n23291), .dinb(n23076), .dout(n23292));
  jand g23035(.dina(n23292), .dinb(n1008), .dout(n23293));
  jnot g23036(.din(n22987), .dout(n23294));
  jor  g23037(.dina(n23294), .dinb(n23293), .dout(n23295));
  jand g23038(.dina(n23295), .dinb(n23075), .dout(n23296));
  jand g23039(.dina(n23296), .dinb(n884), .dout(n23297));
  jor  g23040(.dina(n22994), .dinb(n23297), .dout(n23298));
  jand g23041(.dina(n23298), .dinb(n23074), .dout(n23299));
  jand g23042(.dina(n23299), .dinb(n743), .dout(n23300));
  jnot g23043(.din(n23002), .dout(n23301));
  jor  g23044(.dina(n23301), .dinb(n23300), .dout(n23302));
  jand g23045(.dina(n23302), .dinb(n23073), .dout(n23303));
  jand g23046(.dina(n23303), .dinb(n635), .dout(n23304));
  jor  g23047(.dina(n23009), .dinb(n23304), .dout(n23305));
  jand g23048(.dina(n23305), .dinb(n23072), .dout(n23306));
  jand g23049(.dina(n23306), .dinb(n515), .dout(n23307));
  jor  g23050(.dina(n23017), .dinb(n23307), .dout(n23308));
  jand g23051(.dina(n23308), .dinb(n23071), .dout(n23309));
  jand g23052(.dina(n23309), .dinb(n443), .dout(n23310));
  jnot g23053(.din(n23025), .dout(n23311));
  jor  g23054(.dina(n23311), .dinb(n23310), .dout(n23312));
  jand g23055(.dina(n23312), .dinb(n23070), .dout(n23313));
  jand g23056(.dina(n23313), .dinb(n352), .dout(n23314));
  jnot g23057(.din(n23032), .dout(n23315));
  jor  g23058(.dina(n23315), .dinb(n23314), .dout(n23316));
  jand g23059(.dina(n23316), .dinb(n23069), .dout(n23317));
  jand g23060(.dina(n23317), .dinb(n294), .dout(n23318));
  jor  g23061(.dina(n23039), .dinb(n23318), .dout(n23319));
  jand g23062(.dina(n23319), .dinb(n23068), .dout(n23320));
  jand g23063(.dina(n23320), .dinb(n239), .dout(n23321));
  jor  g23064(.dina(n23047), .dinb(n23321), .dout(n23322));
  jand g23065(.dina(n23322), .dinb(n23067), .dout(n23323));
  jand g23066(.dina(n23323), .dinb(n221), .dout(n23324));
  jor  g23067(.dina(n23055), .dinb(n23324), .dout(n23325));
  jand g23068(.dina(n23325), .dinb(n23066), .dout(n23326));
  jor  g23069(.dina(n23061), .dinb(n23326), .dout(n23327));
  jor  g23070(.dina(n23327), .dinb(n22321), .dout(n23328));
  jor  g23071(.dina(n23328), .dinb(n23065), .dout(n23329));
  jand g23072(.dina(n23329), .dinb(n218), .dout(n23330));
  jand g23073(.dina(n22619), .dinb(n22317), .dout(n23331));
  jnot g23074(.din(n23331), .dout(n23332));
  jxor g23075(.dina(n22320), .dinb(n22317), .dout(n23333));
  jand g23076(.dina(n23333), .dinb(n23332), .dout(n23334));
  jand g23077(.dina(n23334), .dinb(asqrt[63] ), .dout(n23335));
  jor  g23078(.dina(n23335), .dinb(n23330), .dout(n23336));
  jor  g23079(.dina(n23336), .dinb(n23064), .dout(asqrt[3] ));
  jnot g23080(.din(n23065), .dout(n23338));
  jand g23081(.dina(n23062), .dinb(n23058), .dout(n23339));
  jand g23082(.dina(n23339), .dinb(n22345), .dout(n23340));
  jand g23083(.dina(n23340), .dinb(n23338), .dout(n23341));
  jor  g23084(.dina(n23341), .dinb(asqrt[63] ), .dout(n23342));
  jnot g23085(.din(n23335), .dout(n23343));
  jand g23086(.dina(n23343), .dinb(n23342), .dout(n23344));
  jand g23087(.dina(n23344), .dinb(n23063), .dout(n23345));
  jxor g23088(.dina(n23050), .dinb(n221), .dout(n23346));
  jor  g23089(.dina(n23346), .dinb(n23345), .dout(n23347));
  jxor g23090(.dina(n23347), .dinb(n23055), .dout(n23348));
  jnot g23091(.din(n23348), .dout(n23349));
  jor  g23092(.dina(n23345), .dinb(n22334), .dout(n23350));
  jnot g23093(.din(a[4] ), .dout(n23351));
  jnot g23094(.din(a[5] ), .dout(n23352));
  jand g23095(.dina(n23352), .dinb(n23351), .dout(n23353));
  jand g23096(.dina(n23353), .dinb(n22334), .dout(n23354));
  jnot g23097(.din(n23354), .dout(n23355));
  jand g23098(.dina(n23355), .dinb(n23350), .dout(n23356));
  jor  g23099(.dina(n23356), .dinb(n22620), .dout(n23357));
  jand g23100(.dina(n23356), .dinb(n22620), .dout(n23358));
  jor  g23101(.dina(n23345), .dinb(a[6] ), .dout(n23359));
  jand g23102(.dina(n23359), .dinb(a[7] ), .dout(n23360));
  jand g23103(.dina(asqrt[3] ), .dinb(n22336), .dout(n23361));
  jor  g23104(.dina(n23361), .dinb(n23360), .dout(n23362));
  jor  g23105(.dina(n23362), .dinb(n23358), .dout(n23363));
  jand g23106(.dina(n23363), .dinb(n23357), .dout(n23364));
  jor  g23107(.dina(n23364), .dinb(n21887), .dout(n23365));
  jand g23108(.dina(n23364), .dinb(n21887), .dout(n23366));
  jnot g23109(.din(n22336), .dout(n23367));
  jor  g23110(.dina(n23345), .dinb(n23367), .dout(n23368));
  jor  g23111(.dina(asqrt[3] ), .dinb(n22620), .dout(n23369));
  jand g23112(.dina(n23369), .dinb(n23368), .dout(n23370));
  jxor g23113(.dina(n23370), .dinb(n21889), .dout(n23371));
  jor  g23114(.dina(n23371), .dinb(n23366), .dout(n23372));
  jand g23115(.dina(n23372), .dinb(n23365), .dout(n23373));
  jor  g23116(.dina(n23373), .dinb(n21184), .dout(n23374));
  jand g23117(.dina(n23373), .dinb(n21184), .dout(n23375));
  jxor g23118(.dina(n22339), .dinb(n21887), .dout(n23376));
  jor  g23119(.dina(n23376), .dinb(n23345), .dout(n23377));
  jxor g23120(.dina(n23377), .dinb(n22622), .dout(n23378));
  jor  g23121(.dina(n23378), .dinb(n23375), .dout(n23379));
  jand g23122(.dina(n23379), .dinb(n23374), .dout(n23380));
  jor  g23123(.dina(n23380), .dinb(n20468), .dout(n23381));
  jand g23124(.dina(n23380), .dinb(n20468), .dout(n23382));
  jxor g23125(.dina(n22624), .dinb(n21184), .dout(n23383));
  jor  g23126(.dina(n23383), .dinb(n23345), .dout(n23384));
  jxor g23127(.dina(n23384), .dinb(n22630), .dout(n23385));
  jor  g23128(.dina(n23385), .dinb(n23382), .dout(n23386));
  jand g23129(.dina(n23386), .dinb(n23381), .dout(n23387));
  jor  g23130(.dina(n23387), .dinb(n19791), .dout(n23388));
  jand g23131(.dina(n23387), .dinb(n19791), .dout(n23389));
  jxor g23132(.dina(n22632), .dinb(n20468), .dout(n23390));
  jor  g23133(.dina(n23390), .dinb(n23345), .dout(n23391));
  jxor g23134(.dina(n23391), .dinb(n23138), .dout(n23392));
  jnot g23135(.din(n23392), .dout(n23393));
  jor  g23136(.dina(n23393), .dinb(n23389), .dout(n23394));
  jand g23137(.dina(n23394), .dinb(n23388), .dout(n23395));
  jor  g23138(.dina(n23395), .dinb(n19096), .dout(n23396));
  jand g23139(.dina(n23395), .dinb(n19096), .dout(n23397));
  jxor g23140(.dina(n22639), .dinb(n19791), .dout(n23398));
  jor  g23141(.dina(n23398), .dinb(n23345), .dout(n23399));
  jxor g23142(.dina(n23399), .dinb(n23142), .dout(n23400));
  jnot g23143(.din(n23400), .dout(n23401));
  jor  g23144(.dina(n23401), .dinb(n23397), .dout(n23402));
  jand g23145(.dina(n23402), .dinb(n23396), .dout(n23403));
  jor  g23146(.dina(n23403), .dinb(n18442), .dout(n23404));
  jand g23147(.dina(n23403), .dinb(n18442), .dout(n23405));
  jxor g23148(.dina(n22646), .dinb(n19096), .dout(n23406));
  jor  g23149(.dina(n23406), .dinb(n23345), .dout(n23407));
  jxor g23150(.dina(n23407), .dinb(n23146), .dout(n23408));
  jnot g23151(.din(n23408), .dout(n23409));
  jor  g23152(.dina(n23409), .dinb(n23405), .dout(n23410));
  jand g23153(.dina(n23410), .dinb(n23404), .dout(n23411));
  jor  g23154(.dina(n23411), .dinb(n17769), .dout(n23412));
  jand g23155(.dina(n23411), .dinb(n17769), .dout(n23413));
  jxor g23156(.dina(n22653), .dinb(n18442), .dout(n23414));
  jor  g23157(.dina(n23414), .dinb(n23345), .dout(n23415));
  jxor g23158(.dina(n23415), .dinb(n22659), .dout(n23416));
  jor  g23159(.dina(n23416), .dinb(n23413), .dout(n23417));
  jand g23160(.dina(n23417), .dinb(n23412), .dout(n23418));
  jor  g23161(.dina(n23418), .dinb(n17134), .dout(n23419));
  jand g23162(.dina(n23418), .dinb(n17134), .dout(n23420));
  jxor g23163(.dina(n22661), .dinb(n17769), .dout(n23421));
  jor  g23164(.dina(n23421), .dinb(n23345), .dout(n23422));
  jxor g23165(.dina(n23422), .dinb(n23153), .dout(n23423));
  jnot g23166(.din(n23423), .dout(n23424));
  jor  g23167(.dina(n23424), .dinb(n23420), .dout(n23425));
  jand g23168(.dina(n23425), .dinb(n23419), .dout(n23426));
  jor  g23169(.dina(n23426), .dinb(n16489), .dout(n23427));
  jand g23170(.dina(n23426), .dinb(n16489), .dout(n23428));
  jxor g23171(.dina(n22668), .dinb(n17134), .dout(n23429));
  jor  g23172(.dina(n23429), .dinb(n23345), .dout(n23430));
  jxor g23173(.dina(n23430), .dinb(n22674), .dout(n23431));
  jor  g23174(.dina(n23431), .dinb(n23428), .dout(n23432));
  jand g23175(.dina(n23432), .dinb(n23427), .dout(n23433));
  jor  g23176(.dina(n23433), .dinb(n15878), .dout(n23434));
  jand g23177(.dina(n23433), .dinb(n15878), .dout(n23435));
  jxor g23178(.dina(n22676), .dinb(n16489), .dout(n23436));
  jor  g23179(.dina(n23436), .dinb(n23345), .dout(n23437));
  jxor g23180(.dina(n23437), .dinb(n23160), .dout(n23438));
  jnot g23181(.din(n23438), .dout(n23439));
  jor  g23182(.dina(n23439), .dinb(n23435), .dout(n23440));
  jand g23183(.dina(n23440), .dinb(n23434), .dout(n23441));
  jor  g23184(.dina(n23441), .dinb(n15260), .dout(n23442));
  jand g23185(.dina(n23441), .dinb(n15260), .dout(n23443));
  jxor g23186(.dina(n22683), .dinb(n15878), .dout(n23444));
  jor  g23187(.dina(n23444), .dinb(n23345), .dout(n23445));
  jxor g23188(.dina(n23445), .dinb(n22689), .dout(n23446));
  jor  g23189(.dina(n23446), .dinb(n23443), .dout(n23447));
  jand g23190(.dina(n23447), .dinb(n23442), .dout(n23448));
  jor  g23191(.dina(n23448), .dinb(n14674), .dout(n23449));
  jand g23192(.dina(n23448), .dinb(n14674), .dout(n23450));
  jxor g23193(.dina(n22691), .dinb(n15260), .dout(n23451));
  jor  g23194(.dina(n23451), .dinb(n23345), .dout(n23452));
  jxor g23195(.dina(n23452), .dinb(n22697), .dout(n23453));
  jor  g23196(.dina(n23453), .dinb(n23450), .dout(n23454));
  jand g23197(.dina(n23454), .dinb(n23449), .dout(n23455));
  jor  g23198(.dina(n23455), .dinb(n14078), .dout(n23456));
  jand g23199(.dina(n23455), .dinb(n14078), .dout(n23457));
  jxor g23200(.dina(n22699), .dinb(n14674), .dout(n23458));
  jor  g23201(.dina(n23458), .dinb(n23345), .dout(n23459));
  jxor g23202(.dina(n23459), .dinb(n22705), .dout(n23460));
  jor  g23203(.dina(n23460), .dinb(n23457), .dout(n23461));
  jand g23204(.dina(n23461), .dinb(n23456), .dout(n23462));
  jor  g23205(.dina(n23462), .dinb(n13515), .dout(n23463));
  jand g23206(.dina(n23462), .dinb(n13515), .dout(n23464));
  jxor g23207(.dina(n22707), .dinb(n14078), .dout(n23465));
  jor  g23208(.dina(n23465), .dinb(n23345), .dout(n23466));
  jxor g23209(.dina(n23466), .dinb(n23173), .dout(n23467));
  jnot g23210(.din(n23467), .dout(n23468));
  jor  g23211(.dina(n23468), .dinb(n23464), .dout(n23469));
  jand g23212(.dina(n23469), .dinb(n23463), .dout(n23470));
  jor  g23213(.dina(n23470), .dinb(n12947), .dout(n23471));
  jand g23214(.dina(n23470), .dinb(n12947), .dout(n23472));
  jxor g23215(.dina(n22714), .dinb(n13515), .dout(n23473));
  jor  g23216(.dina(n23473), .dinb(n23345), .dout(n23474));
  jxor g23217(.dina(n23474), .dinb(n22720), .dout(n23475));
  jor  g23218(.dina(n23475), .dinb(n23472), .dout(n23476));
  jand g23219(.dina(n23476), .dinb(n23471), .dout(n23477));
  jor  g23220(.dina(n23477), .dinb(n12410), .dout(n23478));
  jand g23221(.dina(n23477), .dinb(n12410), .dout(n23479));
  jxor g23222(.dina(n22722), .dinb(n12947), .dout(n23480));
  jor  g23223(.dina(n23480), .dinb(n23345), .dout(n23481));
  jxor g23224(.dina(n23481), .dinb(n22728), .dout(n23482));
  jor  g23225(.dina(n23482), .dinb(n23479), .dout(n23483));
  jand g23226(.dina(n23483), .dinb(n23478), .dout(n23484));
  jor  g23227(.dina(n23484), .dinb(n11858), .dout(n23485));
  jand g23228(.dina(n23484), .dinb(n11858), .dout(n23486));
  jxor g23229(.dina(n22730), .dinb(n12410), .dout(n23487));
  jor  g23230(.dina(n23487), .dinb(n23345), .dout(n23488));
  jxor g23231(.dina(n23488), .dinb(n22736), .dout(n23489));
  jor  g23232(.dina(n23489), .dinb(n23486), .dout(n23490));
  jand g23233(.dina(n23490), .dinb(n23485), .dout(n23491));
  jor  g23234(.dina(n23491), .dinb(n11347), .dout(n23492));
  jand g23235(.dina(n23491), .dinb(n11347), .dout(n23493));
  jxor g23236(.dina(n22738), .dinb(n11858), .dout(n23494));
  jor  g23237(.dina(n23494), .dinb(n23345), .dout(n23495));
  jxor g23238(.dina(n23495), .dinb(n23186), .dout(n23496));
  jnot g23239(.din(n23496), .dout(n23497));
  jor  g23240(.dina(n23497), .dinb(n23493), .dout(n23498));
  jand g23241(.dina(n23498), .dinb(n23492), .dout(n23499));
  jor  g23242(.dina(n23499), .dinb(n10824), .dout(n23500));
  jand g23243(.dina(n23499), .dinb(n10824), .dout(n23501));
  jxor g23244(.dina(n22745), .dinb(n11347), .dout(n23502));
  jor  g23245(.dina(n23502), .dinb(n23345), .dout(n23503));
  jxor g23246(.dina(n23503), .dinb(n22751), .dout(n23504));
  jor  g23247(.dina(n23504), .dinb(n23501), .dout(n23505));
  jand g23248(.dina(n23505), .dinb(n23500), .dout(n23506));
  jor  g23249(.dina(n23506), .dinb(n10328), .dout(n23507));
  jand g23250(.dina(n23506), .dinb(n10328), .dout(n23508));
  jxor g23251(.dina(n22753), .dinb(n10824), .dout(n23509));
  jor  g23252(.dina(n23509), .dinb(n23345), .dout(n23510));
  jxor g23253(.dina(n23510), .dinb(n23193), .dout(n23511));
  jnot g23254(.din(n23511), .dout(n23512));
  jor  g23255(.dina(n23512), .dinb(n23508), .dout(n23513));
  jand g23256(.dina(n23513), .dinb(n23507), .dout(n23514));
  jor  g23257(.dina(n23514), .dinb(n9832), .dout(n23515));
  jand g23258(.dina(n23514), .dinb(n9832), .dout(n23516));
  jxor g23259(.dina(n22760), .dinb(n10328), .dout(n23517));
  jor  g23260(.dina(n23517), .dinb(n23345), .dout(n23518));
  jxor g23261(.dina(n23518), .dinb(n22766), .dout(n23519));
  jor  g23262(.dina(n23519), .dinb(n23516), .dout(n23520));
  jand g23263(.dina(n23520), .dinb(n23515), .dout(n23521));
  jor  g23264(.dina(n23521), .dinb(n9369), .dout(n23522));
  jand g23265(.dina(n23521), .dinb(n9369), .dout(n23523));
  jxor g23266(.dina(n22768), .dinb(n9832), .dout(n23524));
  jor  g23267(.dina(n23524), .dinb(n23345), .dout(n23525));
  jxor g23268(.dina(n23525), .dinb(n23200), .dout(n23526));
  jnot g23269(.din(n23526), .dout(n23527));
  jor  g23270(.dina(n23527), .dinb(n23523), .dout(n23528));
  jand g23271(.dina(n23528), .dinb(n23522), .dout(n23529));
  jor  g23272(.dina(n23529), .dinb(n8890), .dout(n23530));
  jand g23273(.dina(n23529), .dinb(n8890), .dout(n23531));
  jxor g23274(.dina(n22775), .dinb(n9369), .dout(n23532));
  jor  g23275(.dina(n23532), .dinb(n23345), .dout(n23533));
  jxor g23276(.dina(n23533), .dinb(n22781), .dout(n23534));
  jor  g23277(.dina(n23534), .dinb(n23531), .dout(n23535));
  jand g23278(.dina(n23535), .dinb(n23530), .dout(n23536));
  jor  g23279(.dina(n23536), .dinb(n8449), .dout(n23537));
  jand g23280(.dina(n23536), .dinb(n8449), .dout(n23538));
  jxor g23281(.dina(n22783), .dinb(n8890), .dout(n23539));
  jor  g23282(.dina(n23539), .dinb(n23345), .dout(n23540));
  jxor g23283(.dina(n23540), .dinb(n22789), .dout(n23541));
  jor  g23284(.dina(n23541), .dinb(n23538), .dout(n23542));
  jand g23285(.dina(n23542), .dinb(n23537), .dout(n23543));
  jor  g23286(.dina(n23543), .dinb(n8003), .dout(n23544));
  jand g23287(.dina(n23543), .dinb(n8003), .dout(n23545));
  jxor g23288(.dina(n22791), .dinb(n8449), .dout(n23546));
  jor  g23289(.dina(n23546), .dinb(n23345), .dout(n23547));
  jxor g23290(.dina(n23547), .dinb(n23210), .dout(n23548));
  jnot g23291(.din(n23548), .dout(n23549));
  jor  g23292(.dina(n23549), .dinb(n23545), .dout(n23550));
  jand g23293(.dina(n23550), .dinb(n23544), .dout(n23551));
  jor  g23294(.dina(n23551), .dinb(n7581), .dout(n23552));
  jand g23295(.dina(n23551), .dinb(n7581), .dout(n23553));
  jxor g23296(.dina(n22798), .dinb(n8003), .dout(n23554));
  jor  g23297(.dina(n23554), .dinb(n23345), .dout(n23555));
  jxor g23298(.dina(n23555), .dinb(n23214), .dout(n23556));
  jnot g23299(.din(n23556), .dout(n23557));
  jor  g23300(.dina(n23557), .dinb(n23553), .dout(n23558));
  jand g23301(.dina(n23558), .dinb(n23552), .dout(n23559));
  jor  g23302(.dina(n23559), .dinb(n7154), .dout(n23560));
  jand g23303(.dina(n23559), .dinb(n7154), .dout(n23561));
  jxor g23304(.dina(n22805), .dinb(n7581), .dout(n23562));
  jor  g23305(.dina(n23562), .dinb(n23345), .dout(n23563));
  jxor g23306(.dina(n23563), .dinb(n22811), .dout(n23564));
  jor  g23307(.dina(n23564), .dinb(n23561), .dout(n23565));
  jand g23308(.dina(n23565), .dinb(n23560), .dout(n23566));
  jor  g23309(.dina(n23566), .dinb(n6758), .dout(n23567));
  jand g23310(.dina(n23566), .dinb(n6758), .dout(n23568));
  jxor g23311(.dina(n22813), .dinb(n7154), .dout(n23569));
  jor  g23312(.dina(n23569), .dinb(n23345), .dout(n23570));
  jxor g23313(.dina(n23570), .dinb(n23221), .dout(n23571));
  jnot g23314(.din(n23571), .dout(n23572));
  jor  g23315(.dina(n23572), .dinb(n23568), .dout(n23573));
  jand g23316(.dina(n23573), .dinb(n23567), .dout(n23574));
  jor  g23317(.dina(n23574), .dinb(n6357), .dout(n23575));
  jand g23318(.dina(n23574), .dinb(n6357), .dout(n23576));
  jxor g23319(.dina(n22820), .dinb(n6758), .dout(n23577));
  jor  g23320(.dina(n23577), .dinb(n23345), .dout(n23578));
  jxor g23321(.dina(n23578), .dinb(n22826), .dout(n23579));
  jor  g23322(.dina(n23579), .dinb(n23576), .dout(n23580));
  jand g23323(.dina(n23580), .dinb(n23575), .dout(n23581));
  jor  g23324(.dina(n23581), .dinb(n5989), .dout(n23582));
  jand g23325(.dina(n23581), .dinb(n5989), .dout(n23583));
  jxor g23326(.dina(n22828), .dinb(n6357), .dout(n23584));
  jor  g23327(.dina(n23584), .dinb(n23345), .dout(n23585));
  jxor g23328(.dina(n23585), .dinb(n23228), .dout(n23586));
  jnot g23329(.din(n23586), .dout(n23587));
  jor  g23330(.dina(n23587), .dinb(n23583), .dout(n23588));
  jand g23331(.dina(n23588), .dinb(n23582), .dout(n23589));
  jor  g23332(.dina(n23589), .dinb(n5606), .dout(n23590));
  jand g23333(.dina(n23589), .dinb(n5606), .dout(n23591));
  jxor g23334(.dina(n22835), .dinb(n5989), .dout(n23592));
  jor  g23335(.dina(n23592), .dinb(n23345), .dout(n23593));
  jxor g23336(.dina(n23593), .dinb(n22841), .dout(n23594));
  jor  g23337(.dina(n23594), .dinb(n23591), .dout(n23595));
  jand g23338(.dina(n23595), .dinb(n23590), .dout(n23596));
  jor  g23339(.dina(n23596), .dinb(n5259), .dout(n23597));
  jand g23340(.dina(n23596), .dinb(n5259), .dout(n23598));
  jxor g23341(.dina(n22843), .dinb(n5606), .dout(n23599));
  jor  g23342(.dina(n23599), .dinb(n23345), .dout(n23600));
  jxor g23343(.dina(n23600), .dinb(n22849), .dout(n23601));
  jor  g23344(.dina(n23601), .dinb(n23598), .dout(n23602));
  jand g23345(.dina(n23602), .dinb(n23597), .dout(n23603));
  jor  g23346(.dina(n23603), .dinb(n4902), .dout(n23604));
  jand g23347(.dina(n23603), .dinb(n4902), .dout(n23605));
  jxor g23348(.dina(n22851), .dinb(n5259), .dout(n23606));
  jor  g23349(.dina(n23606), .dinb(n23345), .dout(n23607));
  jxor g23350(.dina(n23607), .dinb(n22857), .dout(n23608));
  jor  g23351(.dina(n23608), .dinb(n23605), .dout(n23609));
  jand g23352(.dina(n23609), .dinb(n23604), .dout(n23610));
  jor  g23353(.dina(n23610), .dinb(n4582), .dout(n23611));
  jand g23354(.dina(n23610), .dinb(n4582), .dout(n23612));
  jxor g23355(.dina(n22859), .dinb(n4902), .dout(n23613));
  jor  g23356(.dina(n23613), .dinb(n23345), .dout(n23614));
  jxor g23357(.dina(n23614), .dinb(n23241), .dout(n23615));
  jnot g23358(.din(n23615), .dout(n23616));
  jor  g23359(.dina(n23616), .dinb(n23612), .dout(n23617));
  jand g23360(.dina(n23617), .dinb(n23611), .dout(n23618));
  jor  g23361(.dina(n23618), .dinb(n4249), .dout(n23619));
  jand g23362(.dina(n23618), .dinb(n4249), .dout(n23620));
  jxor g23363(.dina(n22866), .dinb(n4582), .dout(n23621));
  jor  g23364(.dina(n23621), .dinb(n23345), .dout(n23622));
  jxor g23365(.dina(n23622), .dinb(n22872), .dout(n23623));
  jor  g23366(.dina(n23623), .dinb(n23620), .dout(n23624));
  jand g23367(.dina(n23624), .dinb(n23619), .dout(n23625));
  jor  g23368(.dina(n23625), .dinb(n3955), .dout(n23626));
  jand g23369(.dina(n23625), .dinb(n3955), .dout(n23627));
  jxor g23370(.dina(n22874), .dinb(n4249), .dout(n23628));
  jor  g23371(.dina(n23628), .dinb(n23345), .dout(n23629));
  jxor g23372(.dina(n23629), .dinb(n23248), .dout(n23630));
  jnot g23373(.din(n23630), .dout(n23631));
  jor  g23374(.dina(n23631), .dinb(n23627), .dout(n23632));
  jand g23375(.dina(n23632), .dinb(n23626), .dout(n23633));
  jor  g23376(.dina(n23633), .dinb(n3642), .dout(n23634));
  jand g23377(.dina(n23633), .dinb(n3642), .dout(n23635));
  jxor g23378(.dina(n22881), .dinb(n3955), .dout(n23636));
  jor  g23379(.dina(n23636), .dinb(n23345), .dout(n23637));
  jxor g23380(.dina(n23637), .dinb(n22887), .dout(n23638));
  jor  g23381(.dina(n23638), .dinb(n23635), .dout(n23639));
  jand g23382(.dina(n23639), .dinb(n23634), .dout(n23640));
  jor  g23383(.dina(n23640), .dinb(n3368), .dout(n23641));
  jand g23384(.dina(n23640), .dinb(n3368), .dout(n23642));
  jxor g23385(.dina(n22889), .dinb(n3642), .dout(n23643));
  jor  g23386(.dina(n23643), .dinb(n23345), .dout(n23644));
  jxor g23387(.dina(n23644), .dinb(n23255), .dout(n23645));
  jnot g23388(.din(n23645), .dout(n23646));
  jor  g23389(.dina(n23646), .dinb(n23642), .dout(n23647));
  jand g23390(.dina(n23647), .dinb(n23641), .dout(n23648));
  jor  g23391(.dina(n23648), .dinb(n3089), .dout(n23649));
  jand g23392(.dina(n23648), .dinb(n3089), .dout(n23650));
  jxor g23393(.dina(n22896), .dinb(n3368), .dout(n23651));
  jor  g23394(.dina(n23651), .dinb(n23345), .dout(n23652));
  jxor g23395(.dina(n23652), .dinb(n22902), .dout(n23653));
  jor  g23396(.dina(n23653), .dinb(n23650), .dout(n23654));
  jand g23397(.dina(n23654), .dinb(n23649), .dout(n23655));
  jor  g23398(.dina(n23655), .dinb(n2833), .dout(n23656));
  jand g23399(.dina(n23655), .dinb(n2833), .dout(n23657));
  jxor g23400(.dina(n22904), .dinb(n3089), .dout(n23658));
  jor  g23401(.dina(n23658), .dinb(n23345), .dout(n23659));
  jxor g23402(.dina(n23659), .dinb(n23262), .dout(n23660));
  jnot g23403(.din(n23660), .dout(n23661));
  jor  g23404(.dina(n23661), .dinb(n23657), .dout(n23662));
  jand g23405(.dina(n23662), .dinb(n23656), .dout(n23663));
  jor  g23406(.dina(n23663), .dinb(n2572), .dout(n23664));
  jand g23407(.dina(n23663), .dinb(n2572), .dout(n23665));
  jxor g23408(.dina(n22911), .dinb(n2833), .dout(n23666));
  jor  g23409(.dina(n23666), .dinb(n23345), .dout(n23667));
  jxor g23410(.dina(n23667), .dinb(n22917), .dout(n23668));
  jor  g23411(.dina(n23668), .dinb(n23665), .dout(n23669));
  jand g23412(.dina(n23669), .dinb(n23664), .dout(n23670));
  jor  g23413(.dina(n23670), .dinb(n2345), .dout(n23671));
  jand g23414(.dina(n23670), .dinb(n2345), .dout(n23672));
  jxor g23415(.dina(n22919), .dinb(n2572), .dout(n23673));
  jor  g23416(.dina(n23673), .dinb(n23345), .dout(n23674));
  jxor g23417(.dina(n23674), .dinb(n22925), .dout(n23675));
  jor  g23418(.dina(n23675), .dinb(n23672), .dout(n23676));
  jand g23419(.dina(n23676), .dinb(n23671), .dout(n23677));
  jor  g23420(.dina(n23677), .dinb(n2108), .dout(n23678));
  jand g23421(.dina(n23677), .dinb(n2108), .dout(n23679));
  jxor g23422(.dina(n22927), .dinb(n2345), .dout(n23680));
  jor  g23423(.dina(n23680), .dinb(n23345), .dout(n23681));
  jxor g23424(.dina(n23681), .dinb(n22933), .dout(n23682));
  jor  g23425(.dina(n23682), .dinb(n23679), .dout(n23683));
  jand g23426(.dina(n23683), .dinb(n23678), .dout(n23684));
  jor  g23427(.dina(n23684), .dinb(n1912), .dout(n23685));
  jand g23428(.dina(n23684), .dinb(n1912), .dout(n23686));
  jxor g23429(.dina(n22935), .dinb(n2108), .dout(n23687));
  jor  g23430(.dina(n23687), .dinb(n23345), .dout(n23688));
  jxor g23431(.dina(n23688), .dinb(n23275), .dout(n23689));
  jnot g23432(.din(n23689), .dout(n23690));
  jor  g23433(.dina(n23690), .dinb(n23686), .dout(n23691));
  jand g23434(.dina(n23691), .dinb(n23685), .dout(n23692));
  jor  g23435(.dina(n23692), .dinb(n1699), .dout(n23693));
  jand g23436(.dina(n23692), .dinb(n1699), .dout(n23694));
  jxor g23437(.dina(n22942), .dinb(n1912), .dout(n23695));
  jor  g23438(.dina(n23695), .dinb(n23345), .dout(n23696));
  jxor g23439(.dina(n23696), .dinb(n22948), .dout(n23697));
  jor  g23440(.dina(n23697), .dinb(n23694), .dout(n23698));
  jand g23441(.dina(n23698), .dinb(n23693), .dout(n23699));
  jor  g23442(.dina(n23699), .dinb(n1516), .dout(n23700));
  jand g23443(.dina(n23699), .dinb(n1516), .dout(n23701));
  jxor g23444(.dina(n22950), .dinb(n1699), .dout(n23702));
  jor  g23445(.dina(n23702), .dinb(n23345), .dout(n23703));
  jxor g23446(.dina(n23703), .dinb(n22956), .dout(n23704));
  jor  g23447(.dina(n23704), .dinb(n23701), .dout(n23705));
  jand g23448(.dina(n23705), .dinb(n23700), .dout(n23706));
  jor  g23449(.dina(n23706), .dinb(n1332), .dout(n23707));
  jand g23450(.dina(n23706), .dinb(n1332), .dout(n23708));
  jxor g23451(.dina(n22958), .dinb(n1516), .dout(n23709));
  jor  g23452(.dina(n23709), .dinb(n23345), .dout(n23710));
  jxor g23453(.dina(n23710), .dinb(n22964), .dout(n23711));
  jor  g23454(.dina(n23711), .dinb(n23708), .dout(n23712));
  jand g23455(.dina(n23712), .dinb(n23707), .dout(n23713));
  jor  g23456(.dina(n23713), .dinb(n1173), .dout(n23714));
  jand g23457(.dina(n23713), .dinb(n1173), .dout(n23715));
  jxor g23458(.dina(n22966), .dinb(n1332), .dout(n23716));
  jor  g23459(.dina(n23716), .dinb(n23345), .dout(n23717));
  jxor g23460(.dina(n23717), .dinb(n22972), .dout(n23718));
  jor  g23461(.dina(n23718), .dinb(n23715), .dout(n23719));
  jand g23462(.dina(n23719), .dinb(n23714), .dout(n23720));
  jor  g23463(.dina(n23720), .dinb(n1008), .dout(n23721));
  jand g23464(.dina(n23720), .dinb(n1008), .dout(n23722));
  jxor g23465(.dina(n22974), .dinb(n1173), .dout(n23723));
  jor  g23466(.dina(n23723), .dinb(n23345), .dout(n23724));
  jxor g23467(.dina(n23724), .dinb(n22980), .dout(n23725));
  jor  g23468(.dina(n23725), .dinb(n23722), .dout(n23726));
  jand g23469(.dina(n23726), .dinb(n23721), .dout(n23727));
  jor  g23470(.dina(n23727), .dinb(n884), .dout(n23728));
  jand g23471(.dina(n23727), .dinb(n884), .dout(n23729));
  jxor g23472(.dina(n22982), .dinb(n1008), .dout(n23730));
  jor  g23473(.dina(n23730), .dinb(n23345), .dout(n23731));
  jxor g23474(.dina(n23731), .dinb(n23294), .dout(n23732));
  jnot g23475(.din(n23732), .dout(n23733));
  jor  g23476(.dina(n23733), .dinb(n23729), .dout(n23734));
  jand g23477(.dina(n23734), .dinb(n23728), .dout(n23735));
  jor  g23478(.dina(n23735), .dinb(n743), .dout(n23736));
  jand g23479(.dina(n23735), .dinb(n743), .dout(n23737));
  jxor g23480(.dina(n22989), .dinb(n884), .dout(n23738));
  jor  g23481(.dina(n23738), .dinb(n23345), .dout(n23739));
  jxor g23482(.dina(n23739), .dinb(n22995), .dout(n23740));
  jor  g23483(.dina(n23740), .dinb(n23737), .dout(n23741));
  jand g23484(.dina(n23741), .dinb(n23736), .dout(n23742));
  jor  g23485(.dina(n23742), .dinb(n635), .dout(n23743));
  jand g23486(.dina(n23742), .dinb(n635), .dout(n23744));
  jxor g23487(.dina(n22997), .dinb(n743), .dout(n23745));
  jor  g23488(.dina(n23745), .dinb(n23345), .dout(n23746));
  jxor g23489(.dina(n23746), .dinb(n23301), .dout(n23747));
  jnot g23490(.din(n23747), .dout(n23748));
  jor  g23491(.dina(n23748), .dinb(n23744), .dout(n23749));
  jand g23492(.dina(n23749), .dinb(n23743), .dout(n23750));
  jor  g23493(.dina(n23750), .dinb(n515), .dout(n23751));
  jand g23494(.dina(n23750), .dinb(n515), .dout(n23752));
  jxor g23495(.dina(n23004), .dinb(n635), .dout(n23753));
  jor  g23496(.dina(n23753), .dinb(n23345), .dout(n23754));
  jxor g23497(.dina(n23754), .dinb(n23010), .dout(n23755));
  jor  g23498(.dina(n23755), .dinb(n23752), .dout(n23756));
  jand g23499(.dina(n23756), .dinb(n23751), .dout(n23757));
  jor  g23500(.dina(n23757), .dinb(n443), .dout(n23758));
  jand g23501(.dina(n23757), .dinb(n443), .dout(n23759));
  jxor g23502(.dina(n23012), .dinb(n515), .dout(n23760));
  jor  g23503(.dina(n23760), .dinb(n23345), .dout(n23761));
  jxor g23504(.dina(n23761), .dinb(n23018), .dout(n23762));
  jor  g23505(.dina(n23762), .dinb(n23759), .dout(n23763));
  jand g23506(.dina(n23763), .dinb(n23758), .dout(n23764));
  jor  g23507(.dina(n23764), .dinb(n352), .dout(n23765));
  jand g23508(.dina(n23764), .dinb(n352), .dout(n23766));
  jxor g23509(.dina(n23020), .dinb(n443), .dout(n23767));
  jor  g23510(.dina(n23767), .dinb(n23345), .dout(n23768));
  jxor g23511(.dina(n23768), .dinb(n23311), .dout(n23769));
  jnot g23512(.din(n23769), .dout(n23770));
  jor  g23513(.dina(n23770), .dinb(n23766), .dout(n23771));
  jand g23514(.dina(n23771), .dinb(n23765), .dout(n23772));
  jor  g23515(.dina(n23772), .dinb(n294), .dout(n23773));
  jand g23516(.dina(n23772), .dinb(n294), .dout(n23774));
  jxor g23517(.dina(n23027), .dinb(n352), .dout(n23775));
  jor  g23518(.dina(n23775), .dinb(n23345), .dout(n23776));
  jxor g23519(.dina(n23776), .dinb(n23315), .dout(n23777));
  jnot g23520(.din(n23777), .dout(n23778));
  jor  g23521(.dina(n23778), .dinb(n23774), .dout(n23779));
  jand g23522(.dina(n23779), .dinb(n23773), .dout(n23780));
  jor  g23523(.dina(n23780), .dinb(n239), .dout(n23781));
  jand g23524(.dina(n23780), .dinb(n239), .dout(n23782));
  jxor g23525(.dina(n23034), .dinb(n294), .dout(n23783));
  jor  g23526(.dina(n23783), .dinb(n23345), .dout(n23784));
  jxor g23527(.dina(n23784), .dinb(n23040), .dout(n23785));
  jor  g23528(.dina(n23785), .dinb(n23782), .dout(n23786));
  jand g23529(.dina(n23786), .dinb(n23781), .dout(n23787));
  jor  g23530(.dina(n23787), .dinb(n221), .dout(n23788));
  jand g23531(.dina(n23787), .dinb(n221), .dout(n23789));
  jxor g23532(.dina(n23042), .dinb(n239), .dout(n23790));
  jor  g23533(.dina(n23790), .dinb(n23345), .dout(n23791));
  jxor g23534(.dina(n23791), .dinb(n23048), .dout(n23792));
  jor  g23535(.dina(n23792), .dinb(n23789), .dout(n23793));
  jand g23536(.dina(n23793), .dinb(n23788), .dout(n23794));
  jand g23537(.dina(n23794), .dinb(n23349), .dout(n23795));
  jand g23538(.dina(n23336), .dinb(n23339), .dout(n23796));
  jor  g23539(.dina(n23794), .dinb(n23349), .dout(n23797));
  jor  g23540(.dina(n23797), .dinb(n23064), .dout(n23798));
  jor  g23541(.dina(n23798), .dinb(n23796), .dout(n23799));
  jand g23542(.dina(n23799), .dinb(n218), .dout(n23800));
  jand g23543(.dina(n23344), .dinb(n23326), .dout(n23801));
  jnot g23544(.din(n23801), .dout(n23802));
  jand g23545(.dina(n23063), .dinb(asqrt[63] ), .dout(n23803));
  jand g23546(.dina(n23803), .dinb(n23327), .dout(n23804));
  jand g23547(.dina(n23804), .dinb(n23802), .dout(n23805));
  jor  g23548(.dina(n23805), .dinb(n23800), .dout(n23806));
  jor  g23549(.dina(n23806), .dinb(n23795), .dout(asqrt[2] ));
  jand g23550(.dina(asqrt[2] ), .dinb(a[4] ), .dout(n23808));
  jor  g23551(.dina(a[3] ), .dinb(a[2] ), .dout(n23809));
  jnot g23552(.din(n23809), .dout(n23810));
  jand g23553(.dina(n23810), .dinb(n23351), .dout(n23811));
  jor  g23554(.dina(n23811), .dinb(n23808), .dout(n23812));
  jand g23555(.dina(n23812), .dinb(asqrt[3] ), .dout(n23813));
  jor  g23556(.dina(n23812), .dinb(asqrt[3] ), .dout(n23814));
  jand g23557(.dina(asqrt[2] ), .dinb(n23351), .dout(n23815));
  jor  g23558(.dina(n23815), .dinb(n23352), .dout(n23816));
  jnot g23559(.din(n23353), .dout(n23817));
  jnot g23560(.din(n23795), .dout(n23818));
  jnot g23561(.din(n23796), .dout(n23819));
  jnot g23562(.din(n23788), .dout(n23820));
  jnot g23563(.din(n23781), .dout(n23821));
  jnot g23564(.din(n23773), .dout(n23822));
  jnot g23565(.din(n23765), .dout(n23823));
  jnot g23566(.din(n23758), .dout(n23824));
  jnot g23567(.din(n23751), .dout(n23825));
  jnot g23568(.din(n23743), .dout(n23826));
  jnot g23569(.din(n23736), .dout(n23827));
  jnot g23570(.din(n23728), .dout(n23828));
  jnot g23571(.din(n23721), .dout(n23829));
  jnot g23572(.din(n23714), .dout(n23830));
  jnot g23573(.din(n23707), .dout(n23831));
  jnot g23574(.din(n23700), .dout(n23832));
  jnot g23575(.din(n23693), .dout(n23833));
  jnot g23576(.din(n23685), .dout(n23834));
  jnot g23577(.din(n23678), .dout(n23835));
  jnot g23578(.din(n23671), .dout(n23836));
  jnot g23579(.din(n23664), .dout(n23837));
  jnot g23580(.din(n23656), .dout(n23838));
  jnot g23581(.din(n23649), .dout(n23839));
  jnot g23582(.din(n23641), .dout(n23840));
  jnot g23583(.din(n23634), .dout(n23841));
  jnot g23584(.din(n23626), .dout(n23842));
  jnot g23585(.din(n23619), .dout(n23843));
  jnot g23586(.din(n23611), .dout(n23844));
  jnot g23587(.din(n23604), .dout(n23845));
  jnot g23588(.din(n23597), .dout(n23846));
  jnot g23589(.din(n23590), .dout(n23847));
  jnot g23590(.din(n23582), .dout(n23848));
  jnot g23591(.din(n23575), .dout(n23849));
  jnot g23592(.din(n23567), .dout(n23850));
  jnot g23593(.din(n23560), .dout(n23851));
  jnot g23594(.din(n23552), .dout(n23852));
  jnot g23595(.din(n23544), .dout(n23853));
  jnot g23596(.din(n23537), .dout(n23854));
  jnot g23597(.din(n23530), .dout(n23855));
  jnot g23598(.din(n23522), .dout(n23856));
  jnot g23599(.din(n23515), .dout(n23857));
  jnot g23600(.din(n23507), .dout(n23858));
  jnot g23601(.din(n23500), .dout(n23859));
  jnot g23602(.din(n23492), .dout(n23860));
  jnot g23603(.din(n23485), .dout(n23861));
  jnot g23604(.din(n23478), .dout(n23862));
  jnot g23605(.din(n23471), .dout(n23863));
  jnot g23606(.din(n23463), .dout(n23864));
  jnot g23607(.din(n23456), .dout(n23865));
  jnot g23608(.din(n23449), .dout(n23866));
  jnot g23609(.din(n23442), .dout(n23867));
  jnot g23610(.din(n23434), .dout(n23868));
  jnot g23611(.din(n23427), .dout(n23869));
  jnot g23612(.din(n23419), .dout(n23870));
  jnot g23613(.din(n23412), .dout(n23871));
  jnot g23614(.din(n23404), .dout(n23872));
  jnot g23615(.din(n23396), .dout(n23873));
  jnot g23616(.din(n23388), .dout(n23874));
  jnot g23617(.din(n23381), .dout(n23875));
  jnot g23618(.din(n23374), .dout(n23876));
  jnot g23619(.din(n23365), .dout(n23877));
  jnot g23620(.din(n23357), .dout(n23878));
  jand g23621(.dina(asqrt[3] ), .dinb(a[6] ), .dout(n23879));
  jor  g23622(.dina(n23354), .dinb(n23879), .dout(n23880));
  jor  g23623(.dina(n23880), .dinb(asqrt[4] ), .dout(n23881));
  jand g23624(.dina(asqrt[3] ), .dinb(n22334), .dout(n23882));
  jor  g23625(.dina(n23882), .dinb(n22335), .dout(n23883));
  jand g23626(.dina(n23368), .dinb(n23883), .dout(n23884));
  jand g23627(.dina(n23884), .dinb(n23881), .dout(n23885));
  jor  g23628(.dina(n23885), .dinb(n23878), .dout(n23886));
  jor  g23629(.dina(n23886), .dinb(asqrt[5] ), .dout(n23887));
  jnot g23630(.din(n23371), .dout(n23888));
  jand g23631(.dina(n23888), .dinb(n23887), .dout(n23889));
  jor  g23632(.dina(n23889), .dinb(n23877), .dout(n23890));
  jor  g23633(.dina(n23890), .dinb(asqrt[6] ), .dout(n23891));
  jnot g23634(.din(n23378), .dout(n23892));
  jand g23635(.dina(n23892), .dinb(n23891), .dout(n23893));
  jor  g23636(.dina(n23893), .dinb(n23876), .dout(n23894));
  jor  g23637(.dina(n23894), .dinb(asqrt[7] ), .dout(n23895));
  jnot g23638(.din(n23385), .dout(n23896));
  jand g23639(.dina(n23896), .dinb(n23895), .dout(n23897));
  jor  g23640(.dina(n23897), .dinb(n23875), .dout(n23898));
  jor  g23641(.dina(n23898), .dinb(asqrt[8] ), .dout(n23899));
  jand g23642(.dina(n23392), .dinb(n23899), .dout(n23900));
  jor  g23643(.dina(n23900), .dinb(n23874), .dout(n23901));
  jor  g23644(.dina(n23901), .dinb(asqrt[9] ), .dout(n23902));
  jand g23645(.dina(n23400), .dinb(n23902), .dout(n23903));
  jor  g23646(.dina(n23903), .dinb(n23873), .dout(n23904));
  jor  g23647(.dina(n23904), .dinb(asqrt[10] ), .dout(n23905));
  jand g23648(.dina(n23408), .dinb(n23905), .dout(n23906));
  jor  g23649(.dina(n23906), .dinb(n23872), .dout(n23907));
  jor  g23650(.dina(n23907), .dinb(asqrt[11] ), .dout(n23908));
  jnot g23651(.din(n23416), .dout(n23909));
  jand g23652(.dina(n23909), .dinb(n23908), .dout(n23910));
  jor  g23653(.dina(n23910), .dinb(n23871), .dout(n23911));
  jor  g23654(.dina(n23911), .dinb(asqrt[12] ), .dout(n23912));
  jand g23655(.dina(n23423), .dinb(n23912), .dout(n23913));
  jor  g23656(.dina(n23913), .dinb(n23870), .dout(n23914));
  jor  g23657(.dina(n23914), .dinb(asqrt[13] ), .dout(n23915));
  jnot g23658(.din(n23431), .dout(n23916));
  jand g23659(.dina(n23916), .dinb(n23915), .dout(n23917));
  jor  g23660(.dina(n23917), .dinb(n23869), .dout(n23918));
  jor  g23661(.dina(n23918), .dinb(asqrt[14] ), .dout(n23919));
  jand g23662(.dina(n23438), .dinb(n23919), .dout(n23920));
  jor  g23663(.dina(n23920), .dinb(n23868), .dout(n23921));
  jor  g23664(.dina(n23921), .dinb(asqrt[15] ), .dout(n23922));
  jnot g23665(.din(n23446), .dout(n23923));
  jand g23666(.dina(n23923), .dinb(n23922), .dout(n23924));
  jor  g23667(.dina(n23924), .dinb(n23867), .dout(n23925));
  jor  g23668(.dina(n23925), .dinb(asqrt[16] ), .dout(n23926));
  jnot g23669(.din(n23453), .dout(n23927));
  jand g23670(.dina(n23927), .dinb(n23926), .dout(n23928));
  jor  g23671(.dina(n23928), .dinb(n23866), .dout(n23929));
  jor  g23672(.dina(n23929), .dinb(asqrt[17] ), .dout(n23930));
  jnot g23673(.din(n23460), .dout(n23931));
  jand g23674(.dina(n23931), .dinb(n23930), .dout(n23932));
  jor  g23675(.dina(n23932), .dinb(n23865), .dout(n23933));
  jor  g23676(.dina(n23933), .dinb(asqrt[18] ), .dout(n23934));
  jand g23677(.dina(n23467), .dinb(n23934), .dout(n23935));
  jor  g23678(.dina(n23935), .dinb(n23864), .dout(n23936));
  jor  g23679(.dina(n23936), .dinb(asqrt[19] ), .dout(n23937));
  jnot g23680(.din(n23475), .dout(n23938));
  jand g23681(.dina(n23938), .dinb(n23937), .dout(n23939));
  jor  g23682(.dina(n23939), .dinb(n23863), .dout(n23940));
  jor  g23683(.dina(n23940), .dinb(asqrt[20] ), .dout(n23941));
  jnot g23684(.din(n23482), .dout(n23942));
  jand g23685(.dina(n23942), .dinb(n23941), .dout(n23943));
  jor  g23686(.dina(n23943), .dinb(n23862), .dout(n23944));
  jor  g23687(.dina(n23944), .dinb(asqrt[21] ), .dout(n23945));
  jnot g23688(.din(n23489), .dout(n23946));
  jand g23689(.dina(n23946), .dinb(n23945), .dout(n23947));
  jor  g23690(.dina(n23947), .dinb(n23861), .dout(n23948));
  jor  g23691(.dina(n23948), .dinb(asqrt[22] ), .dout(n23949));
  jand g23692(.dina(n23496), .dinb(n23949), .dout(n23950));
  jor  g23693(.dina(n23950), .dinb(n23860), .dout(n23951));
  jor  g23694(.dina(n23951), .dinb(asqrt[23] ), .dout(n23952));
  jnot g23695(.din(n23504), .dout(n23953));
  jand g23696(.dina(n23953), .dinb(n23952), .dout(n23954));
  jor  g23697(.dina(n23954), .dinb(n23859), .dout(n23955));
  jor  g23698(.dina(n23955), .dinb(asqrt[24] ), .dout(n23956));
  jand g23699(.dina(n23511), .dinb(n23956), .dout(n23957));
  jor  g23700(.dina(n23957), .dinb(n23858), .dout(n23958));
  jor  g23701(.dina(n23958), .dinb(asqrt[25] ), .dout(n23959));
  jnot g23702(.din(n23519), .dout(n23960));
  jand g23703(.dina(n23960), .dinb(n23959), .dout(n23961));
  jor  g23704(.dina(n23961), .dinb(n23857), .dout(n23962));
  jor  g23705(.dina(n23962), .dinb(asqrt[26] ), .dout(n23963));
  jand g23706(.dina(n23526), .dinb(n23963), .dout(n23964));
  jor  g23707(.dina(n23964), .dinb(n23856), .dout(n23965));
  jor  g23708(.dina(n23965), .dinb(asqrt[27] ), .dout(n23966));
  jnot g23709(.din(n23534), .dout(n23967));
  jand g23710(.dina(n23967), .dinb(n23966), .dout(n23968));
  jor  g23711(.dina(n23968), .dinb(n23855), .dout(n23969));
  jor  g23712(.dina(n23969), .dinb(asqrt[28] ), .dout(n23970));
  jnot g23713(.din(n23541), .dout(n23971));
  jand g23714(.dina(n23971), .dinb(n23970), .dout(n23972));
  jor  g23715(.dina(n23972), .dinb(n23854), .dout(n23973));
  jor  g23716(.dina(n23973), .dinb(asqrt[29] ), .dout(n23974));
  jand g23717(.dina(n23548), .dinb(n23974), .dout(n23975));
  jor  g23718(.dina(n23975), .dinb(n23853), .dout(n23976));
  jor  g23719(.dina(n23976), .dinb(asqrt[30] ), .dout(n23977));
  jand g23720(.dina(n23556), .dinb(n23977), .dout(n23978));
  jor  g23721(.dina(n23978), .dinb(n23852), .dout(n23979));
  jor  g23722(.dina(n23979), .dinb(asqrt[31] ), .dout(n23980));
  jnot g23723(.din(n23564), .dout(n23981));
  jand g23724(.dina(n23981), .dinb(n23980), .dout(n23982));
  jor  g23725(.dina(n23982), .dinb(n23851), .dout(n23983));
  jor  g23726(.dina(n23983), .dinb(asqrt[32] ), .dout(n23984));
  jand g23727(.dina(n23571), .dinb(n23984), .dout(n23985));
  jor  g23728(.dina(n23985), .dinb(n23850), .dout(n23986));
  jor  g23729(.dina(n23986), .dinb(asqrt[33] ), .dout(n23987));
  jnot g23730(.din(n23579), .dout(n23988));
  jand g23731(.dina(n23988), .dinb(n23987), .dout(n23989));
  jor  g23732(.dina(n23989), .dinb(n23849), .dout(n23990));
  jor  g23733(.dina(n23990), .dinb(asqrt[34] ), .dout(n23991));
  jand g23734(.dina(n23586), .dinb(n23991), .dout(n23992));
  jor  g23735(.dina(n23992), .dinb(n23848), .dout(n23993));
  jor  g23736(.dina(n23993), .dinb(asqrt[35] ), .dout(n23994));
  jnot g23737(.din(n23594), .dout(n23995));
  jand g23738(.dina(n23995), .dinb(n23994), .dout(n23996));
  jor  g23739(.dina(n23996), .dinb(n23847), .dout(n23997));
  jor  g23740(.dina(n23997), .dinb(asqrt[36] ), .dout(n23998));
  jnot g23741(.din(n23601), .dout(n23999));
  jand g23742(.dina(n23999), .dinb(n23998), .dout(n24000));
  jor  g23743(.dina(n24000), .dinb(n23846), .dout(n24001));
  jor  g23744(.dina(n24001), .dinb(asqrt[37] ), .dout(n24002));
  jnot g23745(.din(n23608), .dout(n24003));
  jand g23746(.dina(n24003), .dinb(n24002), .dout(n24004));
  jor  g23747(.dina(n24004), .dinb(n23845), .dout(n24005));
  jor  g23748(.dina(n24005), .dinb(asqrt[38] ), .dout(n24006));
  jand g23749(.dina(n23615), .dinb(n24006), .dout(n24007));
  jor  g23750(.dina(n24007), .dinb(n23844), .dout(n24008));
  jor  g23751(.dina(n24008), .dinb(asqrt[39] ), .dout(n24009));
  jnot g23752(.din(n23623), .dout(n24010));
  jand g23753(.dina(n24010), .dinb(n24009), .dout(n24011));
  jor  g23754(.dina(n24011), .dinb(n23843), .dout(n24012));
  jor  g23755(.dina(n24012), .dinb(asqrt[40] ), .dout(n24013));
  jand g23756(.dina(n23630), .dinb(n24013), .dout(n24014));
  jor  g23757(.dina(n24014), .dinb(n23842), .dout(n24015));
  jor  g23758(.dina(n24015), .dinb(asqrt[41] ), .dout(n24016));
  jnot g23759(.din(n23638), .dout(n24017));
  jand g23760(.dina(n24017), .dinb(n24016), .dout(n24018));
  jor  g23761(.dina(n24018), .dinb(n23841), .dout(n24019));
  jor  g23762(.dina(n24019), .dinb(asqrt[42] ), .dout(n24020));
  jand g23763(.dina(n23645), .dinb(n24020), .dout(n24021));
  jor  g23764(.dina(n24021), .dinb(n23840), .dout(n24022));
  jor  g23765(.dina(n24022), .dinb(asqrt[43] ), .dout(n24023));
  jnot g23766(.din(n23653), .dout(n24024));
  jand g23767(.dina(n24024), .dinb(n24023), .dout(n24025));
  jor  g23768(.dina(n24025), .dinb(n23839), .dout(n24026));
  jor  g23769(.dina(n24026), .dinb(asqrt[44] ), .dout(n24027));
  jand g23770(.dina(n23660), .dinb(n24027), .dout(n24028));
  jor  g23771(.dina(n24028), .dinb(n23838), .dout(n24029));
  jor  g23772(.dina(n24029), .dinb(asqrt[45] ), .dout(n24030));
  jnot g23773(.din(n23668), .dout(n24031));
  jand g23774(.dina(n24031), .dinb(n24030), .dout(n24032));
  jor  g23775(.dina(n24032), .dinb(n23837), .dout(n24033));
  jor  g23776(.dina(n24033), .dinb(asqrt[46] ), .dout(n24034));
  jnot g23777(.din(n23675), .dout(n24035));
  jand g23778(.dina(n24035), .dinb(n24034), .dout(n24036));
  jor  g23779(.dina(n24036), .dinb(n23836), .dout(n24037));
  jor  g23780(.dina(n24037), .dinb(asqrt[47] ), .dout(n24038));
  jnot g23781(.din(n23682), .dout(n24039));
  jand g23782(.dina(n24039), .dinb(n24038), .dout(n24040));
  jor  g23783(.dina(n24040), .dinb(n23835), .dout(n24041));
  jor  g23784(.dina(n24041), .dinb(asqrt[48] ), .dout(n24042));
  jand g23785(.dina(n23689), .dinb(n24042), .dout(n24043));
  jor  g23786(.dina(n24043), .dinb(n23834), .dout(n24044));
  jor  g23787(.dina(n24044), .dinb(asqrt[49] ), .dout(n24045));
  jnot g23788(.din(n23697), .dout(n24046));
  jand g23789(.dina(n24046), .dinb(n24045), .dout(n24047));
  jor  g23790(.dina(n24047), .dinb(n23833), .dout(n24048));
  jor  g23791(.dina(n24048), .dinb(asqrt[50] ), .dout(n24049));
  jnot g23792(.din(n23704), .dout(n24050));
  jand g23793(.dina(n24050), .dinb(n24049), .dout(n24051));
  jor  g23794(.dina(n24051), .dinb(n23832), .dout(n24052));
  jor  g23795(.dina(n24052), .dinb(asqrt[51] ), .dout(n24053));
  jnot g23796(.din(n23711), .dout(n24054));
  jand g23797(.dina(n24054), .dinb(n24053), .dout(n24055));
  jor  g23798(.dina(n24055), .dinb(n23831), .dout(n24056));
  jor  g23799(.dina(n24056), .dinb(asqrt[52] ), .dout(n24057));
  jnot g23800(.din(n23718), .dout(n24058));
  jand g23801(.dina(n24058), .dinb(n24057), .dout(n24059));
  jor  g23802(.dina(n24059), .dinb(n23830), .dout(n24060));
  jor  g23803(.dina(n24060), .dinb(asqrt[53] ), .dout(n24061));
  jnot g23804(.din(n23725), .dout(n24062));
  jand g23805(.dina(n24062), .dinb(n24061), .dout(n24063));
  jor  g23806(.dina(n24063), .dinb(n23829), .dout(n24064));
  jor  g23807(.dina(n24064), .dinb(asqrt[54] ), .dout(n24065));
  jand g23808(.dina(n23732), .dinb(n24065), .dout(n24066));
  jor  g23809(.dina(n24066), .dinb(n23828), .dout(n24067));
  jor  g23810(.dina(n24067), .dinb(asqrt[55] ), .dout(n24068));
  jnot g23811(.din(n23740), .dout(n24069));
  jand g23812(.dina(n24069), .dinb(n24068), .dout(n24070));
  jor  g23813(.dina(n24070), .dinb(n23827), .dout(n24071));
  jor  g23814(.dina(n24071), .dinb(asqrt[56] ), .dout(n24072));
  jand g23815(.dina(n23747), .dinb(n24072), .dout(n24073));
  jor  g23816(.dina(n24073), .dinb(n23826), .dout(n24074));
  jor  g23817(.dina(n24074), .dinb(asqrt[57] ), .dout(n24075));
  jnot g23818(.din(n23755), .dout(n24076));
  jand g23819(.dina(n24076), .dinb(n24075), .dout(n24077));
  jor  g23820(.dina(n24077), .dinb(n23825), .dout(n24078));
  jor  g23821(.dina(n24078), .dinb(asqrt[58] ), .dout(n24079));
  jnot g23822(.din(n23762), .dout(n24080));
  jand g23823(.dina(n24080), .dinb(n24079), .dout(n24081));
  jor  g23824(.dina(n24081), .dinb(n23824), .dout(n24082));
  jor  g23825(.dina(n24082), .dinb(asqrt[59] ), .dout(n24083));
  jand g23826(.dina(n23769), .dinb(n24083), .dout(n24084));
  jor  g23827(.dina(n24084), .dinb(n23823), .dout(n24085));
  jor  g23828(.dina(n24085), .dinb(asqrt[60] ), .dout(n24086));
  jand g23829(.dina(n23777), .dinb(n24086), .dout(n24087));
  jor  g23830(.dina(n24087), .dinb(n23822), .dout(n24088));
  jor  g23831(.dina(n24088), .dinb(asqrt[61] ), .dout(n24089));
  jnot g23832(.din(n23785), .dout(n24090));
  jand g23833(.dina(n24090), .dinb(n24089), .dout(n24091));
  jor  g23834(.dina(n24091), .dinb(n23821), .dout(n24092));
  jor  g23835(.dina(n24092), .dinb(asqrt[62] ), .dout(n24093));
  jnot g23836(.din(n23792), .dout(n24094));
  jand g23837(.dina(n24094), .dinb(n24093), .dout(n24095));
  jor  g23838(.dina(n24095), .dinb(n23820), .dout(n24096));
  jand g23839(.dina(n24096), .dinb(n23348), .dout(n24097));
  jand g23840(.dina(n24097), .dinb(n23063), .dout(n24098));
  jand g23841(.dina(n24098), .dinb(n23819), .dout(n24099));
  jor  g23842(.dina(n24099), .dinb(asqrt[63] ), .dout(n24100));
  jnot g23843(.din(n23805), .dout(n24101));
  jand g23844(.dina(n24101), .dinb(n24100), .dout(n24102));
  jand g23845(.dina(n24102), .dinb(n23818), .dout(n24103));
  jor  g23846(.dina(n24103), .dinb(n23817), .dout(n24104));
  jand g23847(.dina(n24104), .dinb(n23816), .dout(n24105));
  jand g23848(.dina(n24105), .dinb(n23814), .dout(n24106));
  jor  g23849(.dina(n24106), .dinb(n23813), .dout(n24107));
  jand g23850(.dina(n24107), .dinb(asqrt[4] ), .dout(n24108));
  jor  g23851(.dina(n24107), .dinb(asqrt[4] ), .dout(n24109));
  jor  g23852(.dina(asqrt[2] ), .dinb(n23345), .dout(n24110));
  jand g23853(.dina(n24110), .dinb(n24104), .dout(n24111));
  jxor g23854(.dina(n24111), .dinb(n22334), .dout(n24112));
  jnot g23855(.din(n24112), .dout(n24113));
  jand g23856(.dina(n24113), .dinb(n24109), .dout(n24114));
  jor  g23857(.dina(n24114), .dinb(n24108), .dout(n24115));
  jand g23858(.dina(n24115), .dinb(asqrt[5] ), .dout(n24116));
  jor  g23859(.dina(n24115), .dinb(asqrt[5] ), .dout(n24117));
  jxor g23860(.dina(n23356), .dinb(n22620), .dout(n24118));
  jand g23861(.dina(n24118), .dinb(asqrt[2] ), .dout(n24119));
  jxor g23862(.dina(n24119), .dinb(n23884), .dout(n24120));
  jand g23863(.dina(n24120), .dinb(n24117), .dout(n24121));
  jor  g23864(.dina(n24121), .dinb(n24116), .dout(n24122));
  jand g23865(.dina(n24122), .dinb(asqrt[6] ), .dout(n24123));
  jor  g23866(.dina(n24122), .dinb(asqrt[6] ), .dout(n24124));
  jxor g23867(.dina(n23364), .dinb(n21887), .dout(n24125));
  jand g23868(.dina(n24125), .dinb(asqrt[2] ), .dout(n24126));
  jxor g23869(.dina(n24126), .dinb(n23888), .dout(n24127));
  jand g23870(.dina(n24127), .dinb(n24124), .dout(n24128));
  jor  g23871(.dina(n24128), .dinb(n24123), .dout(n24129));
  jand g23872(.dina(n24129), .dinb(asqrt[7] ), .dout(n24130));
  jor  g23873(.dina(n24129), .dinb(asqrt[7] ), .dout(n24131));
  jxor g23874(.dina(n23373), .dinb(n21184), .dout(n24132));
  jand g23875(.dina(n24132), .dinb(asqrt[2] ), .dout(n24133));
  jxor g23876(.dina(n24133), .dinb(n23378), .dout(n24134));
  jnot g23877(.din(n24134), .dout(n24135));
  jand g23878(.dina(n24135), .dinb(n24131), .dout(n24136));
  jor  g23879(.dina(n24136), .dinb(n24130), .dout(n24137));
  jand g23880(.dina(n24137), .dinb(asqrt[8] ), .dout(n24138));
  jor  g23881(.dina(n24137), .dinb(asqrt[8] ), .dout(n24139));
  jxor g23882(.dina(n23380), .dinb(n20468), .dout(n24140));
  jand g23883(.dina(n24140), .dinb(asqrt[2] ), .dout(n24141));
  jxor g23884(.dina(n24141), .dinb(n23385), .dout(n24142));
  jnot g23885(.din(n24142), .dout(n24143));
  jand g23886(.dina(n24143), .dinb(n24139), .dout(n24144));
  jor  g23887(.dina(n24144), .dinb(n24138), .dout(n24145));
  jand g23888(.dina(n24145), .dinb(asqrt[9] ), .dout(n24146));
  jor  g23889(.dina(n24145), .dinb(asqrt[9] ), .dout(n24147));
  jxor g23890(.dina(n23387), .dinb(n19791), .dout(n24148));
  jand g23891(.dina(n24148), .dinb(asqrt[2] ), .dout(n24149));
  jxor g23892(.dina(n24149), .dinb(n23392), .dout(n24150));
  jand g23893(.dina(n24150), .dinb(n24147), .dout(n24151));
  jor  g23894(.dina(n24151), .dinb(n24146), .dout(n24152));
  jand g23895(.dina(n24152), .dinb(asqrt[10] ), .dout(n24153));
  jor  g23896(.dina(n24152), .dinb(asqrt[10] ), .dout(n24154));
  jxor g23897(.dina(n23395), .dinb(n19096), .dout(n24155));
  jand g23898(.dina(n24155), .dinb(asqrt[2] ), .dout(n24156));
  jxor g23899(.dina(n24156), .dinb(n23400), .dout(n24157));
  jand g23900(.dina(n24157), .dinb(n24154), .dout(n24158));
  jor  g23901(.dina(n24158), .dinb(n24153), .dout(n24159));
  jand g23902(.dina(n24159), .dinb(asqrt[11] ), .dout(n24160));
  jor  g23903(.dina(n24159), .dinb(asqrt[11] ), .dout(n24161));
  jxor g23904(.dina(n23403), .dinb(n18442), .dout(n24162));
  jand g23905(.dina(n24162), .dinb(asqrt[2] ), .dout(n24163));
  jxor g23906(.dina(n24163), .dinb(n23408), .dout(n24164));
  jand g23907(.dina(n24164), .dinb(n24161), .dout(n24165));
  jor  g23908(.dina(n24165), .dinb(n24160), .dout(n24166));
  jand g23909(.dina(n24166), .dinb(asqrt[12] ), .dout(n24167));
  jor  g23910(.dina(n24166), .dinb(asqrt[12] ), .dout(n24168));
  jxor g23911(.dina(n23411), .dinb(n17769), .dout(n24169));
  jand g23912(.dina(n24169), .dinb(asqrt[2] ), .dout(n24170));
  jxor g23913(.dina(n24170), .dinb(n23416), .dout(n24171));
  jnot g23914(.din(n24171), .dout(n24172));
  jand g23915(.dina(n24172), .dinb(n24168), .dout(n24173));
  jor  g23916(.dina(n24173), .dinb(n24167), .dout(n24174));
  jand g23917(.dina(n24174), .dinb(asqrt[13] ), .dout(n24175));
  jor  g23918(.dina(n24174), .dinb(asqrt[13] ), .dout(n24176));
  jxor g23919(.dina(n23418), .dinb(n17134), .dout(n24177));
  jand g23920(.dina(n24177), .dinb(asqrt[2] ), .dout(n24178));
  jxor g23921(.dina(n24178), .dinb(n23423), .dout(n24179));
  jand g23922(.dina(n24179), .dinb(n24176), .dout(n24180));
  jor  g23923(.dina(n24180), .dinb(n24175), .dout(n24181));
  jand g23924(.dina(n24181), .dinb(asqrt[14] ), .dout(n24182));
  jor  g23925(.dina(n24181), .dinb(asqrt[14] ), .dout(n24183));
  jxor g23926(.dina(n23426), .dinb(n16489), .dout(n24184));
  jand g23927(.dina(n24184), .dinb(asqrt[2] ), .dout(n24185));
  jxor g23928(.dina(n24185), .dinb(n23431), .dout(n24186));
  jnot g23929(.din(n24186), .dout(n24187));
  jand g23930(.dina(n24187), .dinb(n24183), .dout(n24188));
  jor  g23931(.dina(n24188), .dinb(n24182), .dout(n24189));
  jand g23932(.dina(n24189), .dinb(asqrt[15] ), .dout(n24190));
  jor  g23933(.dina(n24189), .dinb(asqrt[15] ), .dout(n24191));
  jxor g23934(.dina(n23433), .dinb(n15878), .dout(n24192));
  jand g23935(.dina(n24192), .dinb(asqrt[2] ), .dout(n24193));
  jxor g23936(.dina(n24193), .dinb(n23438), .dout(n24194));
  jand g23937(.dina(n24194), .dinb(n24191), .dout(n24195));
  jor  g23938(.dina(n24195), .dinb(n24190), .dout(n24196));
  jand g23939(.dina(n24196), .dinb(asqrt[16] ), .dout(n24197));
  jor  g23940(.dina(n24196), .dinb(asqrt[16] ), .dout(n24198));
  jxor g23941(.dina(n23441), .dinb(n15260), .dout(n24199));
  jand g23942(.dina(n24199), .dinb(asqrt[2] ), .dout(n24200));
  jxor g23943(.dina(n24200), .dinb(n23446), .dout(n24201));
  jnot g23944(.din(n24201), .dout(n24202));
  jand g23945(.dina(n24202), .dinb(n24198), .dout(n24203));
  jor  g23946(.dina(n24203), .dinb(n24197), .dout(n24204));
  jand g23947(.dina(n24204), .dinb(asqrt[17] ), .dout(n24205));
  jor  g23948(.dina(n24204), .dinb(asqrt[17] ), .dout(n24206));
  jxor g23949(.dina(n23448), .dinb(n14674), .dout(n24207));
  jand g23950(.dina(n24207), .dinb(asqrt[2] ), .dout(n24208));
  jxor g23951(.dina(n24208), .dinb(n23453), .dout(n24209));
  jnot g23952(.din(n24209), .dout(n24210));
  jand g23953(.dina(n24210), .dinb(n24206), .dout(n24211));
  jor  g23954(.dina(n24211), .dinb(n24205), .dout(n24212));
  jand g23955(.dina(n24212), .dinb(asqrt[18] ), .dout(n24213));
  jor  g23956(.dina(n24212), .dinb(asqrt[18] ), .dout(n24214));
  jxor g23957(.dina(n23455), .dinb(n14078), .dout(n24215));
  jand g23958(.dina(n24215), .dinb(asqrt[2] ), .dout(n24216));
  jxor g23959(.dina(n24216), .dinb(n23460), .dout(n24217));
  jnot g23960(.din(n24217), .dout(n24218));
  jand g23961(.dina(n24218), .dinb(n24214), .dout(n24219));
  jor  g23962(.dina(n24219), .dinb(n24213), .dout(n24220));
  jand g23963(.dina(n24220), .dinb(asqrt[19] ), .dout(n24221));
  jor  g23964(.dina(n24220), .dinb(asqrt[19] ), .dout(n24222));
  jxor g23965(.dina(n23462), .dinb(n13515), .dout(n24223));
  jand g23966(.dina(n24223), .dinb(asqrt[2] ), .dout(n24224));
  jxor g23967(.dina(n24224), .dinb(n23467), .dout(n24225));
  jand g23968(.dina(n24225), .dinb(n24222), .dout(n24226));
  jor  g23969(.dina(n24226), .dinb(n24221), .dout(n24227));
  jand g23970(.dina(n24227), .dinb(asqrt[20] ), .dout(n24228));
  jor  g23971(.dina(n24227), .dinb(asqrt[20] ), .dout(n24229));
  jxor g23972(.dina(n23470), .dinb(n12947), .dout(n24230));
  jand g23973(.dina(n24230), .dinb(asqrt[2] ), .dout(n24231));
  jxor g23974(.dina(n24231), .dinb(n23475), .dout(n24232));
  jnot g23975(.din(n24232), .dout(n24233));
  jand g23976(.dina(n24233), .dinb(n24229), .dout(n24234));
  jor  g23977(.dina(n24234), .dinb(n24228), .dout(n24235));
  jand g23978(.dina(n24235), .dinb(asqrt[21] ), .dout(n24236));
  jor  g23979(.dina(n24235), .dinb(asqrt[21] ), .dout(n24237));
  jxor g23980(.dina(n23477), .dinb(n12410), .dout(n24238));
  jand g23981(.dina(n24238), .dinb(asqrt[2] ), .dout(n24239));
  jxor g23982(.dina(n24239), .dinb(n23482), .dout(n24240));
  jnot g23983(.din(n24240), .dout(n24241));
  jand g23984(.dina(n24241), .dinb(n24237), .dout(n24242));
  jor  g23985(.dina(n24242), .dinb(n24236), .dout(n24243));
  jand g23986(.dina(n24243), .dinb(asqrt[22] ), .dout(n24244));
  jor  g23987(.dina(n24243), .dinb(asqrt[22] ), .dout(n24245));
  jxor g23988(.dina(n23484), .dinb(n11858), .dout(n24246));
  jand g23989(.dina(n24246), .dinb(asqrt[2] ), .dout(n24247));
  jxor g23990(.dina(n24247), .dinb(n23489), .dout(n24248));
  jnot g23991(.din(n24248), .dout(n24249));
  jand g23992(.dina(n24249), .dinb(n24245), .dout(n24250));
  jor  g23993(.dina(n24250), .dinb(n24244), .dout(n24251));
  jand g23994(.dina(n24251), .dinb(asqrt[23] ), .dout(n24252));
  jor  g23995(.dina(n24251), .dinb(asqrt[23] ), .dout(n24253));
  jxor g23996(.dina(n23491), .dinb(n11347), .dout(n24254));
  jand g23997(.dina(n24254), .dinb(asqrt[2] ), .dout(n24255));
  jxor g23998(.dina(n24255), .dinb(n23496), .dout(n24256));
  jand g23999(.dina(n24256), .dinb(n24253), .dout(n24257));
  jor  g24000(.dina(n24257), .dinb(n24252), .dout(n24258));
  jand g24001(.dina(n24258), .dinb(asqrt[24] ), .dout(n24259));
  jor  g24002(.dina(n24258), .dinb(asqrt[24] ), .dout(n24260));
  jxor g24003(.dina(n23499), .dinb(n10824), .dout(n24261));
  jand g24004(.dina(n24261), .dinb(asqrt[2] ), .dout(n24262));
  jxor g24005(.dina(n24262), .dinb(n23504), .dout(n24263));
  jnot g24006(.din(n24263), .dout(n24264));
  jand g24007(.dina(n24264), .dinb(n24260), .dout(n24265));
  jor  g24008(.dina(n24265), .dinb(n24259), .dout(n24266));
  jand g24009(.dina(n24266), .dinb(asqrt[25] ), .dout(n24267));
  jor  g24010(.dina(n24266), .dinb(asqrt[25] ), .dout(n24268));
  jxor g24011(.dina(n23506), .dinb(n10328), .dout(n24269));
  jand g24012(.dina(n24269), .dinb(asqrt[2] ), .dout(n24270));
  jxor g24013(.dina(n24270), .dinb(n23511), .dout(n24271));
  jand g24014(.dina(n24271), .dinb(n24268), .dout(n24272));
  jor  g24015(.dina(n24272), .dinb(n24267), .dout(n24273));
  jand g24016(.dina(n24273), .dinb(asqrt[26] ), .dout(n24274));
  jor  g24017(.dina(n24273), .dinb(asqrt[26] ), .dout(n24275));
  jxor g24018(.dina(n23514), .dinb(n9832), .dout(n24276));
  jand g24019(.dina(n24276), .dinb(asqrt[2] ), .dout(n24277));
  jxor g24020(.dina(n24277), .dinb(n23519), .dout(n24278));
  jnot g24021(.din(n24278), .dout(n24279));
  jand g24022(.dina(n24279), .dinb(n24275), .dout(n24280));
  jor  g24023(.dina(n24280), .dinb(n24274), .dout(n24281));
  jand g24024(.dina(n24281), .dinb(asqrt[27] ), .dout(n24282));
  jor  g24025(.dina(n24281), .dinb(asqrt[27] ), .dout(n24283));
  jxor g24026(.dina(n23521), .dinb(n9369), .dout(n24284));
  jand g24027(.dina(n24284), .dinb(asqrt[2] ), .dout(n24285));
  jxor g24028(.dina(n24285), .dinb(n23526), .dout(n24286));
  jand g24029(.dina(n24286), .dinb(n24283), .dout(n24287));
  jor  g24030(.dina(n24287), .dinb(n24282), .dout(n24288));
  jand g24031(.dina(n24288), .dinb(asqrt[28] ), .dout(n24289));
  jor  g24032(.dina(n24288), .dinb(asqrt[28] ), .dout(n24290));
  jxor g24033(.dina(n23529), .dinb(n8890), .dout(n24291));
  jand g24034(.dina(n24291), .dinb(asqrt[2] ), .dout(n24292));
  jxor g24035(.dina(n24292), .dinb(n23534), .dout(n24293));
  jnot g24036(.din(n24293), .dout(n24294));
  jand g24037(.dina(n24294), .dinb(n24290), .dout(n24295));
  jor  g24038(.dina(n24295), .dinb(n24289), .dout(n24296));
  jand g24039(.dina(n24296), .dinb(asqrt[29] ), .dout(n24297));
  jor  g24040(.dina(n24296), .dinb(asqrt[29] ), .dout(n24298));
  jxor g24041(.dina(n23536), .dinb(n8449), .dout(n24299));
  jand g24042(.dina(n24299), .dinb(asqrt[2] ), .dout(n24300));
  jxor g24043(.dina(n24300), .dinb(n23541), .dout(n24301));
  jnot g24044(.din(n24301), .dout(n24302));
  jand g24045(.dina(n24302), .dinb(n24298), .dout(n24303));
  jor  g24046(.dina(n24303), .dinb(n24297), .dout(n24304));
  jand g24047(.dina(n24304), .dinb(asqrt[30] ), .dout(n24305));
  jor  g24048(.dina(n24304), .dinb(asqrt[30] ), .dout(n24306));
  jxor g24049(.dina(n23543), .dinb(n8003), .dout(n24307));
  jand g24050(.dina(n24307), .dinb(asqrt[2] ), .dout(n24308));
  jxor g24051(.dina(n24308), .dinb(n23548), .dout(n24309));
  jand g24052(.dina(n24309), .dinb(n24306), .dout(n24310));
  jor  g24053(.dina(n24310), .dinb(n24305), .dout(n24311));
  jand g24054(.dina(n24311), .dinb(asqrt[31] ), .dout(n24312));
  jor  g24055(.dina(n24311), .dinb(asqrt[31] ), .dout(n24313));
  jxor g24056(.dina(n23551), .dinb(n7581), .dout(n24314));
  jand g24057(.dina(n24314), .dinb(asqrt[2] ), .dout(n24315));
  jxor g24058(.dina(n24315), .dinb(n23556), .dout(n24316));
  jand g24059(.dina(n24316), .dinb(n24313), .dout(n24317));
  jor  g24060(.dina(n24317), .dinb(n24312), .dout(n24318));
  jand g24061(.dina(n24318), .dinb(asqrt[32] ), .dout(n24319));
  jor  g24062(.dina(n24318), .dinb(asqrt[32] ), .dout(n24320));
  jxor g24063(.dina(n23559), .dinb(n7154), .dout(n24321));
  jand g24064(.dina(n24321), .dinb(asqrt[2] ), .dout(n24322));
  jxor g24065(.dina(n24322), .dinb(n23564), .dout(n24323));
  jnot g24066(.din(n24323), .dout(n24324));
  jand g24067(.dina(n24324), .dinb(n24320), .dout(n24325));
  jor  g24068(.dina(n24325), .dinb(n24319), .dout(n24326));
  jand g24069(.dina(n24326), .dinb(asqrt[33] ), .dout(n24327));
  jor  g24070(.dina(n24326), .dinb(asqrt[33] ), .dout(n24328));
  jxor g24071(.dina(n23566), .dinb(n6758), .dout(n24329));
  jand g24072(.dina(n24329), .dinb(asqrt[2] ), .dout(n24330));
  jxor g24073(.dina(n24330), .dinb(n23571), .dout(n24331));
  jand g24074(.dina(n24331), .dinb(n24328), .dout(n24332));
  jor  g24075(.dina(n24332), .dinb(n24327), .dout(n24333));
  jand g24076(.dina(n24333), .dinb(asqrt[34] ), .dout(n24334));
  jor  g24077(.dina(n24333), .dinb(asqrt[34] ), .dout(n24335));
  jxor g24078(.dina(n23574), .dinb(n6357), .dout(n24336));
  jand g24079(.dina(n24336), .dinb(asqrt[2] ), .dout(n24337));
  jxor g24080(.dina(n24337), .dinb(n23579), .dout(n24338));
  jnot g24081(.din(n24338), .dout(n24339));
  jand g24082(.dina(n24339), .dinb(n24335), .dout(n24340));
  jor  g24083(.dina(n24340), .dinb(n24334), .dout(n24341));
  jand g24084(.dina(n24341), .dinb(asqrt[35] ), .dout(n24342));
  jor  g24085(.dina(n24341), .dinb(asqrt[35] ), .dout(n24343));
  jxor g24086(.dina(n23581), .dinb(n5989), .dout(n24344));
  jand g24087(.dina(n24344), .dinb(asqrt[2] ), .dout(n24345));
  jxor g24088(.dina(n24345), .dinb(n23586), .dout(n24346));
  jand g24089(.dina(n24346), .dinb(n24343), .dout(n24347));
  jor  g24090(.dina(n24347), .dinb(n24342), .dout(n24348));
  jand g24091(.dina(n24348), .dinb(asqrt[36] ), .dout(n24349));
  jor  g24092(.dina(n24348), .dinb(asqrt[36] ), .dout(n24350));
  jxor g24093(.dina(n23589), .dinb(n5606), .dout(n24351));
  jand g24094(.dina(n24351), .dinb(asqrt[2] ), .dout(n24352));
  jxor g24095(.dina(n24352), .dinb(n23594), .dout(n24353));
  jnot g24096(.din(n24353), .dout(n24354));
  jand g24097(.dina(n24354), .dinb(n24350), .dout(n24355));
  jor  g24098(.dina(n24355), .dinb(n24349), .dout(n24356));
  jand g24099(.dina(n24356), .dinb(asqrt[37] ), .dout(n24357));
  jor  g24100(.dina(n24356), .dinb(asqrt[37] ), .dout(n24358));
  jxor g24101(.dina(n23596), .dinb(n5259), .dout(n24359));
  jand g24102(.dina(n24359), .dinb(asqrt[2] ), .dout(n24360));
  jxor g24103(.dina(n24360), .dinb(n23601), .dout(n24361));
  jnot g24104(.din(n24361), .dout(n24362));
  jand g24105(.dina(n24362), .dinb(n24358), .dout(n24363));
  jor  g24106(.dina(n24363), .dinb(n24357), .dout(n24364));
  jand g24107(.dina(n24364), .dinb(asqrt[38] ), .dout(n24365));
  jor  g24108(.dina(n24364), .dinb(asqrt[38] ), .dout(n24366));
  jxor g24109(.dina(n23603), .dinb(n4902), .dout(n24367));
  jand g24110(.dina(n24367), .dinb(asqrt[2] ), .dout(n24368));
  jxor g24111(.dina(n24368), .dinb(n23608), .dout(n24369));
  jnot g24112(.din(n24369), .dout(n24370));
  jand g24113(.dina(n24370), .dinb(n24366), .dout(n24371));
  jor  g24114(.dina(n24371), .dinb(n24365), .dout(n24372));
  jand g24115(.dina(n24372), .dinb(asqrt[39] ), .dout(n24373));
  jor  g24116(.dina(n24372), .dinb(asqrt[39] ), .dout(n24374));
  jxor g24117(.dina(n23610), .dinb(n4582), .dout(n24375));
  jand g24118(.dina(n24375), .dinb(asqrt[2] ), .dout(n24376));
  jxor g24119(.dina(n24376), .dinb(n23615), .dout(n24377));
  jand g24120(.dina(n24377), .dinb(n24374), .dout(n24378));
  jor  g24121(.dina(n24378), .dinb(n24373), .dout(n24379));
  jand g24122(.dina(n24379), .dinb(asqrt[40] ), .dout(n24380));
  jor  g24123(.dina(n24379), .dinb(asqrt[40] ), .dout(n24381));
  jxor g24124(.dina(n23618), .dinb(n4249), .dout(n24382));
  jand g24125(.dina(n24382), .dinb(asqrt[2] ), .dout(n24383));
  jxor g24126(.dina(n24383), .dinb(n23623), .dout(n24384));
  jnot g24127(.din(n24384), .dout(n24385));
  jand g24128(.dina(n24385), .dinb(n24381), .dout(n24386));
  jor  g24129(.dina(n24386), .dinb(n24380), .dout(n24387));
  jand g24130(.dina(n24387), .dinb(asqrt[41] ), .dout(n24388));
  jor  g24131(.dina(n24387), .dinb(asqrt[41] ), .dout(n24389));
  jxor g24132(.dina(n23625), .dinb(n3955), .dout(n24390));
  jand g24133(.dina(n24390), .dinb(asqrt[2] ), .dout(n24391));
  jxor g24134(.dina(n24391), .dinb(n23630), .dout(n24392));
  jand g24135(.dina(n24392), .dinb(n24389), .dout(n24393));
  jor  g24136(.dina(n24393), .dinb(n24388), .dout(n24394));
  jand g24137(.dina(n24394), .dinb(asqrt[42] ), .dout(n24395));
  jor  g24138(.dina(n24394), .dinb(asqrt[42] ), .dout(n24396));
  jxor g24139(.dina(n23633), .dinb(n3642), .dout(n24397));
  jand g24140(.dina(n24397), .dinb(asqrt[2] ), .dout(n24398));
  jxor g24141(.dina(n24398), .dinb(n23638), .dout(n24399));
  jnot g24142(.din(n24399), .dout(n24400));
  jand g24143(.dina(n24400), .dinb(n24396), .dout(n24401));
  jor  g24144(.dina(n24401), .dinb(n24395), .dout(n24402));
  jand g24145(.dina(n24402), .dinb(asqrt[43] ), .dout(n24403));
  jor  g24146(.dina(n24402), .dinb(asqrt[43] ), .dout(n24404));
  jxor g24147(.dina(n23640), .dinb(n3368), .dout(n24405));
  jand g24148(.dina(n24405), .dinb(asqrt[2] ), .dout(n24406));
  jxor g24149(.dina(n24406), .dinb(n23645), .dout(n24407));
  jand g24150(.dina(n24407), .dinb(n24404), .dout(n24408));
  jor  g24151(.dina(n24408), .dinb(n24403), .dout(n24409));
  jand g24152(.dina(n24409), .dinb(asqrt[44] ), .dout(n24410));
  jor  g24153(.dina(n24409), .dinb(asqrt[44] ), .dout(n24411));
  jxor g24154(.dina(n23648), .dinb(n3089), .dout(n24412));
  jand g24155(.dina(n24412), .dinb(asqrt[2] ), .dout(n24413));
  jxor g24156(.dina(n24413), .dinb(n23653), .dout(n24414));
  jnot g24157(.din(n24414), .dout(n24415));
  jand g24158(.dina(n24415), .dinb(n24411), .dout(n24416));
  jor  g24159(.dina(n24416), .dinb(n24410), .dout(n24417));
  jand g24160(.dina(n24417), .dinb(asqrt[45] ), .dout(n24418));
  jor  g24161(.dina(n24417), .dinb(asqrt[45] ), .dout(n24419));
  jxor g24162(.dina(n23655), .dinb(n2833), .dout(n24420));
  jand g24163(.dina(n24420), .dinb(asqrt[2] ), .dout(n24421));
  jxor g24164(.dina(n24421), .dinb(n23660), .dout(n24422));
  jand g24165(.dina(n24422), .dinb(n24419), .dout(n24423));
  jor  g24166(.dina(n24423), .dinb(n24418), .dout(n24424));
  jand g24167(.dina(n24424), .dinb(asqrt[46] ), .dout(n24425));
  jor  g24168(.dina(n24424), .dinb(asqrt[46] ), .dout(n24426));
  jxor g24169(.dina(n23663), .dinb(n2572), .dout(n24427));
  jand g24170(.dina(n24427), .dinb(asqrt[2] ), .dout(n24428));
  jxor g24171(.dina(n24428), .dinb(n23668), .dout(n24429));
  jnot g24172(.din(n24429), .dout(n24430));
  jand g24173(.dina(n24430), .dinb(n24426), .dout(n24431));
  jor  g24174(.dina(n24431), .dinb(n24425), .dout(n24432));
  jand g24175(.dina(n24432), .dinb(asqrt[47] ), .dout(n24433));
  jor  g24176(.dina(n24432), .dinb(asqrt[47] ), .dout(n24434));
  jxor g24177(.dina(n23670), .dinb(n2345), .dout(n24435));
  jand g24178(.dina(n24435), .dinb(asqrt[2] ), .dout(n24436));
  jxor g24179(.dina(n24436), .dinb(n23675), .dout(n24437));
  jnot g24180(.din(n24437), .dout(n24438));
  jand g24181(.dina(n24438), .dinb(n24434), .dout(n24439));
  jor  g24182(.dina(n24439), .dinb(n24433), .dout(n24440));
  jand g24183(.dina(n24440), .dinb(asqrt[48] ), .dout(n24441));
  jor  g24184(.dina(n24440), .dinb(asqrt[48] ), .dout(n24442));
  jxor g24185(.dina(n23677), .dinb(n2108), .dout(n24443));
  jand g24186(.dina(n24443), .dinb(asqrt[2] ), .dout(n24444));
  jxor g24187(.dina(n24444), .dinb(n23682), .dout(n24445));
  jnot g24188(.din(n24445), .dout(n24446));
  jand g24189(.dina(n24446), .dinb(n24442), .dout(n24447));
  jor  g24190(.dina(n24447), .dinb(n24441), .dout(n24448));
  jand g24191(.dina(n24448), .dinb(asqrt[49] ), .dout(n24449));
  jor  g24192(.dina(n24448), .dinb(asqrt[49] ), .dout(n24450));
  jxor g24193(.dina(n23684), .dinb(n1912), .dout(n24451));
  jand g24194(.dina(n24451), .dinb(asqrt[2] ), .dout(n24452));
  jxor g24195(.dina(n24452), .dinb(n23689), .dout(n24453));
  jand g24196(.dina(n24453), .dinb(n24450), .dout(n24454));
  jor  g24197(.dina(n24454), .dinb(n24449), .dout(n24455));
  jand g24198(.dina(n24455), .dinb(asqrt[50] ), .dout(n24456));
  jor  g24199(.dina(n24455), .dinb(asqrt[50] ), .dout(n24457));
  jxor g24200(.dina(n23692), .dinb(n1699), .dout(n24458));
  jand g24201(.dina(n24458), .dinb(asqrt[2] ), .dout(n24459));
  jxor g24202(.dina(n24459), .dinb(n23697), .dout(n24460));
  jnot g24203(.din(n24460), .dout(n24461));
  jand g24204(.dina(n24461), .dinb(n24457), .dout(n24462));
  jor  g24205(.dina(n24462), .dinb(n24456), .dout(n24463));
  jand g24206(.dina(n24463), .dinb(asqrt[51] ), .dout(n24464));
  jor  g24207(.dina(n24463), .dinb(asqrt[51] ), .dout(n24465));
  jxor g24208(.dina(n23699), .dinb(n1516), .dout(n24466));
  jand g24209(.dina(n24466), .dinb(asqrt[2] ), .dout(n24467));
  jxor g24210(.dina(n24467), .dinb(n23704), .dout(n24468));
  jnot g24211(.din(n24468), .dout(n24469));
  jand g24212(.dina(n24469), .dinb(n24465), .dout(n24470));
  jor  g24213(.dina(n24470), .dinb(n24464), .dout(n24471));
  jand g24214(.dina(n24471), .dinb(asqrt[52] ), .dout(n24472));
  jor  g24215(.dina(n24471), .dinb(asqrt[52] ), .dout(n24473));
  jxor g24216(.dina(n23706), .dinb(n1332), .dout(n24474));
  jand g24217(.dina(n24474), .dinb(asqrt[2] ), .dout(n24475));
  jxor g24218(.dina(n24475), .dinb(n23711), .dout(n24476));
  jnot g24219(.din(n24476), .dout(n24477));
  jand g24220(.dina(n24477), .dinb(n24473), .dout(n24478));
  jor  g24221(.dina(n24478), .dinb(n24472), .dout(n24479));
  jand g24222(.dina(n24479), .dinb(asqrt[53] ), .dout(n24480));
  jor  g24223(.dina(n24479), .dinb(asqrt[53] ), .dout(n24481));
  jxor g24224(.dina(n23713), .dinb(n1173), .dout(n24482));
  jand g24225(.dina(n24482), .dinb(asqrt[2] ), .dout(n24483));
  jxor g24226(.dina(n24483), .dinb(n23718), .dout(n24484));
  jnot g24227(.din(n24484), .dout(n24485));
  jand g24228(.dina(n24485), .dinb(n24481), .dout(n24486));
  jor  g24229(.dina(n24486), .dinb(n24480), .dout(n24487));
  jand g24230(.dina(n24487), .dinb(asqrt[54] ), .dout(n24488));
  jor  g24231(.dina(n24487), .dinb(asqrt[54] ), .dout(n24489));
  jxor g24232(.dina(n23720), .dinb(n1008), .dout(n24490));
  jand g24233(.dina(n24490), .dinb(asqrt[2] ), .dout(n24491));
  jxor g24234(.dina(n24491), .dinb(n23725), .dout(n24492));
  jnot g24235(.din(n24492), .dout(n24493));
  jand g24236(.dina(n24493), .dinb(n24489), .dout(n24494));
  jor  g24237(.dina(n24494), .dinb(n24488), .dout(n24495));
  jand g24238(.dina(n24495), .dinb(asqrt[55] ), .dout(n24496));
  jor  g24239(.dina(n24495), .dinb(asqrt[55] ), .dout(n24497));
  jxor g24240(.dina(n23727), .dinb(n884), .dout(n24498));
  jand g24241(.dina(n24498), .dinb(asqrt[2] ), .dout(n24499));
  jxor g24242(.dina(n24499), .dinb(n23732), .dout(n24500));
  jand g24243(.dina(n24500), .dinb(n24497), .dout(n24501));
  jor  g24244(.dina(n24501), .dinb(n24496), .dout(n24502));
  jand g24245(.dina(n24502), .dinb(asqrt[56] ), .dout(n24503));
  jor  g24246(.dina(n24502), .dinb(asqrt[56] ), .dout(n24504));
  jxor g24247(.dina(n23735), .dinb(n743), .dout(n24505));
  jand g24248(.dina(n24505), .dinb(asqrt[2] ), .dout(n24506));
  jxor g24249(.dina(n24506), .dinb(n23740), .dout(n24507));
  jnot g24250(.din(n24507), .dout(n24508));
  jand g24251(.dina(n24508), .dinb(n24504), .dout(n24509));
  jor  g24252(.dina(n24509), .dinb(n24503), .dout(n24510));
  jand g24253(.dina(n24510), .dinb(asqrt[57] ), .dout(n24511));
  jor  g24254(.dina(n24510), .dinb(asqrt[57] ), .dout(n24512));
  jxor g24255(.dina(n23742), .dinb(n635), .dout(n24513));
  jand g24256(.dina(n24513), .dinb(asqrt[2] ), .dout(n24514));
  jxor g24257(.dina(n24514), .dinb(n23747), .dout(n24515));
  jand g24258(.dina(n24515), .dinb(n24512), .dout(n24516));
  jor  g24259(.dina(n24516), .dinb(n24511), .dout(n24517));
  jand g24260(.dina(n24517), .dinb(asqrt[58] ), .dout(n24518));
  jor  g24261(.dina(n24517), .dinb(asqrt[58] ), .dout(n24519));
  jxor g24262(.dina(n23750), .dinb(n515), .dout(n24520));
  jand g24263(.dina(n24520), .dinb(asqrt[2] ), .dout(n24521));
  jxor g24264(.dina(n24521), .dinb(n23755), .dout(n24522));
  jnot g24265(.din(n24522), .dout(n24523));
  jand g24266(.dina(n24523), .dinb(n24519), .dout(n24524));
  jor  g24267(.dina(n24524), .dinb(n24518), .dout(n24525));
  jand g24268(.dina(n24525), .dinb(asqrt[59] ), .dout(n24526));
  jor  g24269(.dina(n24525), .dinb(asqrt[59] ), .dout(n24527));
  jxor g24270(.dina(n23757), .dinb(n443), .dout(n24528));
  jand g24271(.dina(n24528), .dinb(asqrt[2] ), .dout(n24529));
  jxor g24272(.dina(n24529), .dinb(n24080), .dout(n24530));
  jand g24273(.dina(n24530), .dinb(n24527), .dout(n24531));
  jor  g24274(.dina(n24531), .dinb(n24526), .dout(n24532));
  jand g24275(.dina(n24532), .dinb(asqrt[60] ), .dout(n24533));
  jor  g24276(.dina(n24532), .dinb(asqrt[60] ), .dout(n24534));
  jxor g24277(.dina(n23764), .dinb(n352), .dout(n24535));
  jand g24278(.dina(n24535), .dinb(asqrt[2] ), .dout(n24536));
  jxor g24279(.dina(n24536), .dinb(n23769), .dout(n24537));
  jand g24280(.dina(n24537), .dinb(n24534), .dout(n24538));
  jor  g24281(.dina(n24538), .dinb(n24533), .dout(n24539));
  jand g24282(.dina(n24539), .dinb(asqrt[61] ), .dout(n24540));
  jor  g24283(.dina(n24539), .dinb(asqrt[61] ), .dout(n24541));
  jxor g24284(.dina(n23772), .dinb(n294), .dout(n24542));
  jand g24285(.dina(n24542), .dinb(asqrt[2] ), .dout(n24543));
  jxor g24286(.dina(n24543), .dinb(n23777), .dout(n24544));
  jand g24287(.dina(n24544), .dinb(n24541), .dout(n24545));
  jor  g24288(.dina(n24545), .dinb(n24540), .dout(n24546));
  jand g24289(.dina(n24546), .dinb(asqrt[62] ), .dout(n24547));
  jor  g24290(.dina(n24546), .dinb(asqrt[62] ), .dout(n24548));
  jxor g24291(.dina(n23780), .dinb(n239), .dout(n24549));
  jand g24292(.dina(n24549), .dinb(asqrt[2] ), .dout(n24550));
  jxor g24293(.dina(n24550), .dinb(n23785), .dout(n24551));
  jnot g24294(.din(n24551), .dout(n24552));
  jand g24295(.dina(n24552), .dinb(n24548), .dout(n24553));
  jor  g24296(.dina(n24553), .dinb(n24547), .dout(n24554));
  jand g24297(.dina(n23806), .dinb(n24097), .dout(n24555));
  jnot g24298(.din(n24547), .dout(n24556));
  jnot g24299(.din(n24540), .dout(n24557));
  jnot g24300(.din(n24533), .dout(n24558));
  jnot g24301(.din(n24526), .dout(n24559));
  jnot g24302(.din(n24518), .dout(n24560));
  jnot g24303(.din(n24511), .dout(n24561));
  jnot g24304(.din(n24503), .dout(n24562));
  jnot g24305(.din(n24496), .dout(n24563));
  jnot g24306(.din(n24488), .dout(n24564));
  jnot g24307(.din(n24480), .dout(n24565));
  jnot g24308(.din(n24472), .dout(n24566));
  jnot g24309(.din(n24464), .dout(n24567));
  jnot g24310(.din(n24456), .dout(n24568));
  jnot g24311(.din(n24449), .dout(n24569));
  jnot g24312(.din(n24441), .dout(n24570));
  jnot g24313(.din(n24433), .dout(n24571));
  jnot g24314(.din(n24425), .dout(n24572));
  jnot g24315(.din(n24418), .dout(n24573));
  jnot g24316(.din(n24410), .dout(n24574));
  jnot g24317(.din(n24403), .dout(n24575));
  jnot g24318(.din(n24395), .dout(n24576));
  jnot g24319(.din(n24388), .dout(n24577));
  jnot g24320(.din(n24380), .dout(n24578));
  jnot g24321(.din(n24373), .dout(n24579));
  jnot g24322(.din(n24365), .dout(n24580));
  jnot g24323(.din(n24357), .dout(n24581));
  jnot g24324(.din(n24349), .dout(n24582));
  jnot g24325(.din(n24342), .dout(n24583));
  jnot g24326(.din(n24334), .dout(n24584));
  jnot g24327(.din(n24327), .dout(n24585));
  jnot g24328(.din(n24319), .dout(n24586));
  jnot g24329(.din(n24312), .dout(n24587));
  jnot g24330(.din(n24305), .dout(n24588));
  jnot g24331(.din(n24297), .dout(n24589));
  jnot g24332(.din(n24289), .dout(n24590));
  jnot g24333(.din(n24282), .dout(n24591));
  jnot g24334(.din(n24274), .dout(n24592));
  jnot g24335(.din(n24267), .dout(n24593));
  jnot g24336(.din(n24259), .dout(n24594));
  jnot g24337(.din(n24252), .dout(n24595));
  jnot g24338(.din(n24244), .dout(n24596));
  jnot g24339(.din(n24236), .dout(n24597));
  jnot g24340(.din(n24228), .dout(n24598));
  jnot g24341(.din(n24221), .dout(n24599));
  jnot g24342(.din(n24213), .dout(n24600));
  jnot g24343(.din(n24205), .dout(n24601));
  jnot g24344(.din(n24197), .dout(n24602));
  jnot g24345(.din(n24190), .dout(n24603));
  jnot g24346(.din(n24182), .dout(n24604));
  jnot g24347(.din(n24175), .dout(n24605));
  jnot g24348(.din(n24167), .dout(n24606));
  jnot g24349(.din(n24160), .dout(n24607));
  jnot g24350(.din(n24153), .dout(n24608));
  jnot g24351(.din(n24146), .dout(n24609));
  jnot g24352(.din(n24138), .dout(n24610));
  jnot g24353(.din(n24130), .dout(n24611));
  jnot g24354(.din(n24123), .dout(n24612));
  jnot g24355(.din(n24116), .dout(n24613));
  jnot g24356(.din(n24108), .dout(n24614));
  jnot g24357(.din(n23813), .dout(n24615));
  jor  g24358(.dina(n24103), .dinb(n23351), .dout(n24616));
  jnot g24359(.din(n23811), .dout(n24617));
  jand g24360(.dina(n24617), .dinb(n24616), .dout(n24618));
  jand g24361(.dina(n24618), .dinb(n23345), .dout(n24619));
  jor  g24362(.dina(n24103), .dinb(a[4] ), .dout(n24620));
  jand g24363(.dina(n24620), .dinb(a[5] ), .dout(n24621));
  jand g24364(.dina(asqrt[2] ), .dinb(n23353), .dout(n24622));
  jor  g24365(.dina(n24622), .dinb(n24621), .dout(n24623));
  jor  g24366(.dina(n24623), .dinb(n24619), .dout(n24624));
  jand g24367(.dina(n24624), .dinb(n24615), .dout(n24625));
  jand g24368(.dina(n24625), .dinb(n22620), .dout(n24626));
  jor  g24369(.dina(n24112), .dinb(n24626), .dout(n24627));
  jand g24370(.dina(n24627), .dinb(n24614), .dout(n24628));
  jand g24371(.dina(n24628), .dinb(n21887), .dout(n24629));
  jnot g24372(.din(n24120), .dout(n24630));
  jor  g24373(.dina(n24630), .dinb(n24629), .dout(n24631));
  jand g24374(.dina(n24631), .dinb(n24613), .dout(n24632));
  jand g24375(.dina(n24632), .dinb(n21184), .dout(n24633));
  jnot g24376(.din(n24127), .dout(n24634));
  jor  g24377(.dina(n24634), .dinb(n24633), .dout(n24635));
  jand g24378(.dina(n24635), .dinb(n24612), .dout(n24636));
  jand g24379(.dina(n24636), .dinb(n20468), .dout(n24637));
  jor  g24380(.dina(n24134), .dinb(n24637), .dout(n24638));
  jand g24381(.dina(n24638), .dinb(n24611), .dout(n24639));
  jand g24382(.dina(n24639), .dinb(n19791), .dout(n24640));
  jor  g24383(.dina(n24142), .dinb(n24640), .dout(n24641));
  jand g24384(.dina(n24641), .dinb(n24610), .dout(n24642));
  jand g24385(.dina(n24642), .dinb(n19096), .dout(n24643));
  jnot g24386(.din(n24150), .dout(n24644));
  jor  g24387(.dina(n24644), .dinb(n24643), .dout(n24645));
  jand g24388(.dina(n24645), .dinb(n24609), .dout(n24646));
  jand g24389(.dina(n24646), .dinb(n18442), .dout(n24647));
  jnot g24390(.din(n24157), .dout(n24648));
  jor  g24391(.dina(n24648), .dinb(n24647), .dout(n24649));
  jand g24392(.dina(n24649), .dinb(n24608), .dout(n24650));
  jand g24393(.dina(n24650), .dinb(n17769), .dout(n24651));
  jnot g24394(.din(n24164), .dout(n24652));
  jor  g24395(.dina(n24652), .dinb(n24651), .dout(n24653));
  jand g24396(.dina(n24653), .dinb(n24607), .dout(n24654));
  jand g24397(.dina(n24654), .dinb(n17134), .dout(n24655));
  jor  g24398(.dina(n24171), .dinb(n24655), .dout(n24656));
  jand g24399(.dina(n24656), .dinb(n24606), .dout(n24657));
  jand g24400(.dina(n24657), .dinb(n16489), .dout(n24658));
  jnot g24401(.din(n24179), .dout(n24659));
  jor  g24402(.dina(n24659), .dinb(n24658), .dout(n24660));
  jand g24403(.dina(n24660), .dinb(n24605), .dout(n24661));
  jand g24404(.dina(n24661), .dinb(n15878), .dout(n24662));
  jor  g24405(.dina(n24186), .dinb(n24662), .dout(n24663));
  jand g24406(.dina(n24663), .dinb(n24604), .dout(n24664));
  jand g24407(.dina(n24664), .dinb(n15260), .dout(n24665));
  jnot g24408(.din(n24194), .dout(n24666));
  jor  g24409(.dina(n24666), .dinb(n24665), .dout(n24667));
  jand g24410(.dina(n24667), .dinb(n24603), .dout(n24668));
  jand g24411(.dina(n24668), .dinb(n14674), .dout(n24669));
  jor  g24412(.dina(n24201), .dinb(n24669), .dout(n24670));
  jand g24413(.dina(n24670), .dinb(n24602), .dout(n24671));
  jand g24414(.dina(n24671), .dinb(n14078), .dout(n24672));
  jor  g24415(.dina(n24209), .dinb(n24672), .dout(n24673));
  jand g24416(.dina(n24673), .dinb(n24601), .dout(n24674));
  jand g24417(.dina(n24674), .dinb(n13515), .dout(n24675));
  jor  g24418(.dina(n24217), .dinb(n24675), .dout(n24676));
  jand g24419(.dina(n24676), .dinb(n24600), .dout(n24677));
  jand g24420(.dina(n24677), .dinb(n12947), .dout(n24678));
  jnot g24421(.din(n24225), .dout(n24679));
  jor  g24422(.dina(n24679), .dinb(n24678), .dout(n24680));
  jand g24423(.dina(n24680), .dinb(n24599), .dout(n24681));
  jand g24424(.dina(n24681), .dinb(n12410), .dout(n24682));
  jor  g24425(.dina(n24232), .dinb(n24682), .dout(n24683));
  jand g24426(.dina(n24683), .dinb(n24598), .dout(n24684));
  jand g24427(.dina(n24684), .dinb(n11858), .dout(n24685));
  jor  g24428(.dina(n24240), .dinb(n24685), .dout(n24686));
  jand g24429(.dina(n24686), .dinb(n24597), .dout(n24687));
  jand g24430(.dina(n24687), .dinb(n11347), .dout(n24688));
  jor  g24431(.dina(n24248), .dinb(n24688), .dout(n24689));
  jand g24432(.dina(n24689), .dinb(n24596), .dout(n24690));
  jand g24433(.dina(n24690), .dinb(n10824), .dout(n24691));
  jnot g24434(.din(n24256), .dout(n24692));
  jor  g24435(.dina(n24692), .dinb(n24691), .dout(n24693));
  jand g24436(.dina(n24693), .dinb(n24595), .dout(n24694));
  jand g24437(.dina(n24694), .dinb(n10328), .dout(n24695));
  jor  g24438(.dina(n24263), .dinb(n24695), .dout(n24696));
  jand g24439(.dina(n24696), .dinb(n24594), .dout(n24697));
  jand g24440(.dina(n24697), .dinb(n9832), .dout(n24698));
  jnot g24441(.din(n24271), .dout(n24699));
  jor  g24442(.dina(n24699), .dinb(n24698), .dout(n24700));
  jand g24443(.dina(n24700), .dinb(n24593), .dout(n24701));
  jand g24444(.dina(n24701), .dinb(n9369), .dout(n24702));
  jor  g24445(.dina(n24278), .dinb(n24702), .dout(n24703));
  jand g24446(.dina(n24703), .dinb(n24592), .dout(n24704));
  jand g24447(.dina(n24704), .dinb(n8890), .dout(n24705));
  jnot g24448(.din(n24286), .dout(n24706));
  jor  g24449(.dina(n24706), .dinb(n24705), .dout(n24707));
  jand g24450(.dina(n24707), .dinb(n24591), .dout(n24708));
  jand g24451(.dina(n24708), .dinb(n8449), .dout(n24709));
  jor  g24452(.dina(n24293), .dinb(n24709), .dout(n24710));
  jand g24453(.dina(n24710), .dinb(n24590), .dout(n24711));
  jand g24454(.dina(n24711), .dinb(n8003), .dout(n24712));
  jor  g24455(.dina(n24301), .dinb(n24712), .dout(n24713));
  jand g24456(.dina(n24713), .dinb(n24589), .dout(n24714));
  jand g24457(.dina(n24714), .dinb(n7581), .dout(n24715));
  jnot g24458(.din(n24309), .dout(n24716));
  jor  g24459(.dina(n24716), .dinb(n24715), .dout(n24717));
  jand g24460(.dina(n24717), .dinb(n24588), .dout(n24718));
  jand g24461(.dina(n24718), .dinb(n7154), .dout(n24719));
  jnot g24462(.din(n24316), .dout(n24720));
  jor  g24463(.dina(n24720), .dinb(n24719), .dout(n24721));
  jand g24464(.dina(n24721), .dinb(n24587), .dout(n24722));
  jand g24465(.dina(n24722), .dinb(n6758), .dout(n24723));
  jor  g24466(.dina(n24323), .dinb(n24723), .dout(n24724));
  jand g24467(.dina(n24724), .dinb(n24586), .dout(n24725));
  jand g24468(.dina(n24725), .dinb(n6357), .dout(n24726));
  jnot g24469(.din(n24331), .dout(n24727));
  jor  g24470(.dina(n24727), .dinb(n24726), .dout(n24728));
  jand g24471(.dina(n24728), .dinb(n24585), .dout(n24729));
  jand g24472(.dina(n24729), .dinb(n5989), .dout(n24730));
  jor  g24473(.dina(n24338), .dinb(n24730), .dout(n24731));
  jand g24474(.dina(n24731), .dinb(n24584), .dout(n24732));
  jand g24475(.dina(n24732), .dinb(n5606), .dout(n24733));
  jnot g24476(.din(n24346), .dout(n24734));
  jor  g24477(.dina(n24734), .dinb(n24733), .dout(n24735));
  jand g24478(.dina(n24735), .dinb(n24583), .dout(n24736));
  jand g24479(.dina(n24736), .dinb(n5259), .dout(n24737));
  jor  g24480(.dina(n24353), .dinb(n24737), .dout(n24738));
  jand g24481(.dina(n24738), .dinb(n24582), .dout(n24739));
  jand g24482(.dina(n24739), .dinb(n4902), .dout(n24740));
  jor  g24483(.dina(n24361), .dinb(n24740), .dout(n24741));
  jand g24484(.dina(n24741), .dinb(n24581), .dout(n24742));
  jand g24485(.dina(n24742), .dinb(n4582), .dout(n24743));
  jor  g24486(.dina(n24369), .dinb(n24743), .dout(n24744));
  jand g24487(.dina(n24744), .dinb(n24580), .dout(n24745));
  jand g24488(.dina(n24745), .dinb(n4249), .dout(n24746));
  jnot g24489(.din(n24377), .dout(n24747));
  jor  g24490(.dina(n24747), .dinb(n24746), .dout(n24748));
  jand g24491(.dina(n24748), .dinb(n24579), .dout(n24749));
  jand g24492(.dina(n24749), .dinb(n3955), .dout(n24750));
  jor  g24493(.dina(n24384), .dinb(n24750), .dout(n24751));
  jand g24494(.dina(n24751), .dinb(n24578), .dout(n24752));
  jand g24495(.dina(n24752), .dinb(n3642), .dout(n24753));
  jnot g24496(.din(n24392), .dout(n24754));
  jor  g24497(.dina(n24754), .dinb(n24753), .dout(n24755));
  jand g24498(.dina(n24755), .dinb(n24577), .dout(n24756));
  jand g24499(.dina(n24756), .dinb(n3368), .dout(n24757));
  jor  g24500(.dina(n24399), .dinb(n24757), .dout(n24758));
  jand g24501(.dina(n24758), .dinb(n24576), .dout(n24759));
  jand g24502(.dina(n24759), .dinb(n3089), .dout(n24760));
  jnot g24503(.din(n24407), .dout(n24761));
  jor  g24504(.dina(n24761), .dinb(n24760), .dout(n24762));
  jand g24505(.dina(n24762), .dinb(n24575), .dout(n24763));
  jand g24506(.dina(n24763), .dinb(n2833), .dout(n24764));
  jor  g24507(.dina(n24414), .dinb(n24764), .dout(n24765));
  jand g24508(.dina(n24765), .dinb(n24574), .dout(n24766));
  jand g24509(.dina(n24766), .dinb(n2572), .dout(n24767));
  jnot g24510(.din(n24422), .dout(n24768));
  jor  g24511(.dina(n24768), .dinb(n24767), .dout(n24769));
  jand g24512(.dina(n24769), .dinb(n24573), .dout(n24770));
  jand g24513(.dina(n24770), .dinb(n2345), .dout(n24771));
  jor  g24514(.dina(n24429), .dinb(n24771), .dout(n24772));
  jand g24515(.dina(n24772), .dinb(n24572), .dout(n24773));
  jand g24516(.dina(n24773), .dinb(n2108), .dout(n24774));
  jor  g24517(.dina(n24437), .dinb(n24774), .dout(n24775));
  jand g24518(.dina(n24775), .dinb(n24571), .dout(n24776));
  jand g24519(.dina(n24776), .dinb(n1912), .dout(n24777));
  jor  g24520(.dina(n24445), .dinb(n24777), .dout(n24778));
  jand g24521(.dina(n24778), .dinb(n24570), .dout(n24779));
  jand g24522(.dina(n24779), .dinb(n1699), .dout(n24780));
  jnot g24523(.din(n24453), .dout(n24781));
  jor  g24524(.dina(n24781), .dinb(n24780), .dout(n24782));
  jand g24525(.dina(n24782), .dinb(n24569), .dout(n24783));
  jand g24526(.dina(n24783), .dinb(n1516), .dout(n24784));
  jor  g24527(.dina(n24460), .dinb(n24784), .dout(n24785));
  jand g24528(.dina(n24785), .dinb(n24568), .dout(n24786));
  jand g24529(.dina(n24786), .dinb(n1332), .dout(n24787));
  jor  g24530(.dina(n24468), .dinb(n24787), .dout(n24788));
  jand g24531(.dina(n24788), .dinb(n24567), .dout(n24789));
  jand g24532(.dina(n24789), .dinb(n1173), .dout(n24790));
  jor  g24533(.dina(n24476), .dinb(n24790), .dout(n24791));
  jand g24534(.dina(n24791), .dinb(n24566), .dout(n24792));
  jand g24535(.dina(n24792), .dinb(n1008), .dout(n24793));
  jor  g24536(.dina(n24484), .dinb(n24793), .dout(n24794));
  jand g24537(.dina(n24794), .dinb(n24565), .dout(n24795));
  jand g24538(.dina(n24795), .dinb(n884), .dout(n24796));
  jor  g24539(.dina(n24492), .dinb(n24796), .dout(n24797));
  jand g24540(.dina(n24797), .dinb(n24564), .dout(n24798));
  jand g24541(.dina(n24798), .dinb(n743), .dout(n24799));
  jnot g24542(.din(n24500), .dout(n24800));
  jor  g24543(.dina(n24800), .dinb(n24799), .dout(n24801));
  jand g24544(.dina(n24801), .dinb(n24563), .dout(n24802));
  jand g24545(.dina(n24802), .dinb(n635), .dout(n24803));
  jor  g24546(.dina(n24507), .dinb(n24803), .dout(n24804));
  jand g24547(.dina(n24804), .dinb(n24562), .dout(n24805));
  jand g24548(.dina(n24805), .dinb(n515), .dout(n24806));
  jnot g24549(.din(n24515), .dout(n24807));
  jor  g24550(.dina(n24807), .dinb(n24806), .dout(n24808));
  jand g24551(.dina(n24808), .dinb(n24561), .dout(n24809));
  jand g24552(.dina(n24809), .dinb(n443), .dout(n24810));
  jor  g24553(.dina(n24522), .dinb(n24810), .dout(n24811));
  jand g24554(.dina(n24811), .dinb(n24560), .dout(n24812));
  jand g24555(.dina(n24812), .dinb(n352), .dout(n24813));
  jnot g24556(.din(n24530), .dout(n24814));
  jor  g24557(.dina(n24814), .dinb(n24813), .dout(n24815));
  jand g24558(.dina(n24815), .dinb(n24559), .dout(n24816));
  jand g24559(.dina(n24816), .dinb(n294), .dout(n24817));
  jnot g24560(.din(n24537), .dout(n24818));
  jor  g24561(.dina(n24818), .dinb(n24817), .dout(n24819));
  jand g24562(.dina(n24819), .dinb(n24558), .dout(n24820));
  jand g24563(.dina(n24820), .dinb(n239), .dout(n24821));
  jnot g24564(.din(n24544), .dout(n24822));
  jor  g24565(.dina(n24822), .dinb(n24821), .dout(n24823));
  jand g24566(.dina(n24823), .dinb(n24557), .dout(n24824));
  jand g24567(.dina(n24824), .dinb(n221), .dout(n24825));
  jor  g24568(.dina(n24551), .dinb(n24825), .dout(n24826));
  jand g24569(.dina(n24826), .dinb(n24556), .dout(n24827));
  jxor g24570(.dina(n23787), .dinb(n221), .dout(n24828));
  jand g24571(.dina(n24828), .dinb(asqrt[2] ), .dout(n24829));
  jxor g24572(.dina(n24829), .dinb(n23792), .dout(n24830));
  jor  g24573(.dina(n24830), .dinb(n24827), .dout(n24831));
  jor  g24574(.dina(n24831), .dinb(n23795), .dout(n24832));
  jor  g24575(.dina(n24832), .dinb(n24555), .dout(n24833));
  jnot g24576(.din(n24830), .dout(n24834));
  jor  g24577(.dina(n24834), .dinb(n24554), .dout(n24835));
  jand g24578(.dina(n24835), .dinb(n218), .dout(n24836));
  jnot g24579(.din(n24836), .dout(n24837));
  jor  g24580(.dina(n24837), .dinb(n24833), .dout(n24838));
  jand g24581(.dina(n24835), .dinb(asqrt[63] ), .dout(n24839));
  jand g24582(.dina(n24102), .dinb(n23794), .dout(n24840));
  jnot g24583(.din(n24840), .dout(n24841));
  jxor g24584(.dina(n23794), .dinb(n23349), .dout(n24842));
  jand g24585(.dina(n24842), .dinb(n24841), .dout(n24843));
  jnot g24586(.din(n24843), .dout(n24844));
  jand g24587(.dina(n24844), .dinb(n24839), .dout(n24845));
  jnot g24588(.din(n24845), .dout(n24846));
  jand g24589(.dina(n24846), .dinb(n24838), .dout(asqrt[1] ));
  jor  g24590(.dina(asqrt[1] ), .dinb(n24554), .dout(n24848));
  jand g24591(.dina(n24839), .dinb(n24831), .dout(n24849));
  jand g24592(.dina(n24849), .dinb(n24848), .dout(n24850));
  jnot g24593(.din(n24555), .dout(n24851));
  jand g24594(.dina(n24834), .dinb(n24554), .dout(n24852));
  jand g24595(.dina(n24852), .dinb(n23818), .dout(n24853));
  jand g24596(.dina(n24853), .dinb(n24851), .dout(n24854));
  jand g24597(.dina(n24836), .dinb(n24854), .dout(n24855));
  jor  g24598(.dina(n24845), .dinb(n24855), .dout(n24856));
  jxor g24599(.dina(n24539), .dinb(n239), .dout(n24857));
  jor  g24600(.dina(n24857), .dinb(n24856), .dout(n24858));
  jxor g24601(.dina(n24858), .dinb(n24544), .dout(n24859));
  jand g24602(.dina(n24859), .dinb(n221), .dout(n24860));
  jxor g24603(.dina(n24487), .dinb(n884), .dout(n24861));
  jor  g24604(.dina(n24861), .dinb(n24856), .dout(n24862));
  jxor g24605(.dina(n24862), .dinb(n24493), .dout(n24863));
  jor  g24606(.dina(n24863), .dinb(n743), .dout(n24864));
  jxor g24607(.dina(n24479), .dinb(n1008), .dout(n24865));
  jor  g24608(.dina(n24865), .dinb(n24856), .dout(n24866));
  jxor g24609(.dina(n24866), .dinb(n24485), .dout(n24867));
  jand g24610(.dina(n24867), .dinb(n884), .dout(n24868));
  jand g24611(.dina(n24863), .dinb(n743), .dout(n24869));
  jor  g24612(.dina(n24869), .dinb(n24868), .dout(n24870));
  jxor g24613(.dina(n24463), .dinb(n1332), .dout(n24871));
  jor  g24614(.dina(n24871), .dinb(n24856), .dout(n24872));
  jxor g24615(.dina(n24872), .dinb(n24469), .dout(n24873));
  jand g24616(.dina(n24873), .dinb(n1173), .dout(n24874));
  jxor g24617(.dina(n24455), .dinb(n1516), .dout(n24875));
  jor  g24618(.dina(n24875), .dinb(n24856), .dout(n24876));
  jxor g24619(.dina(n24876), .dinb(n24461), .dout(n24877));
  jand g24620(.dina(n24877), .dinb(n1332), .dout(n24878));
  jxor g24621(.dina(n24424), .dinb(n2345), .dout(n24879));
  jor  g24622(.dina(n24879), .dinb(n24856), .dout(n24880));
  jxor g24623(.dina(n24880), .dinb(n24430), .dout(n24881));
  jor  g24624(.dina(n24881), .dinb(n2108), .dout(n24882));
  jxor g24625(.dina(n24417), .dinb(n2572), .dout(n24883));
  jor  g24626(.dina(n24883), .dinb(n24856), .dout(n24884));
  jxor g24627(.dina(n24884), .dinb(n24422), .dout(n24885));
  jand g24628(.dina(n24885), .dinb(n2345), .dout(n24886));
  jxor g24629(.dina(n24394), .dinb(n3368), .dout(n24887));
  jor  g24630(.dina(n24887), .dinb(n24856), .dout(n24888));
  jxor g24631(.dina(n24888), .dinb(n24400), .dout(n24889));
  jand g24632(.dina(n24889), .dinb(n3089), .dout(n24890));
  jxor g24633(.dina(n24364), .dinb(n4582), .dout(n24891));
  jor  g24634(.dina(n24891), .dinb(n24856), .dout(n24892));
  jxor g24635(.dina(n24892), .dinb(n24370), .dout(n24893));
  jor  g24636(.dina(n24893), .dinb(n4249), .dout(n24894));
  jxor g24637(.dina(n24356), .dinb(n4902), .dout(n24895));
  jor  g24638(.dina(n24895), .dinb(n24856), .dout(n24896));
  jxor g24639(.dina(n24896), .dinb(n24362), .dout(n24897));
  jand g24640(.dina(n24897), .dinb(n4582), .dout(n24898));
  jxor g24641(.dina(n24318), .dinb(n6758), .dout(n24899));
  jor  g24642(.dina(n24899), .dinb(n24856), .dout(n24900));
  jxor g24643(.dina(n24900), .dinb(n24324), .dout(n24901));
  jor  g24644(.dina(n24901), .dinb(n6357), .dout(n24902));
  jxor g24645(.dina(n24296), .dinb(n8003), .dout(n24903));
  jor  g24646(.dina(n24903), .dinb(n24856), .dout(n24904));
  jxor g24647(.dina(n24904), .dinb(n24302), .dout(n24905));
  jand g24648(.dina(n24905), .dinb(n7581), .dout(n24906));
  jxor g24649(.dina(n24288), .dinb(n8449), .dout(n24907));
  jor  g24650(.dina(n24907), .dinb(n24856), .dout(n24908));
  jxor g24651(.dina(n24908), .dinb(n24294), .dout(n24909));
  jand g24652(.dina(n24909), .dinb(n8003), .dout(n24910));
  jxor g24653(.dina(n24281), .dinb(n8890), .dout(n24911));
  jor  g24654(.dina(n24911), .dinb(n24856), .dout(n24912));
  jxor g24655(.dina(n24912), .dinb(n24286), .dout(n24913));
  jor  g24656(.dina(n24913), .dinb(n8449), .dout(n24914));
  jxor g24657(.dina(n24251), .dinb(n10824), .dout(n24915));
  jor  g24658(.dina(n24915), .dinb(n24856), .dout(n24916));
  jxor g24659(.dina(n24916), .dinb(n24256), .dout(n24917));
  jand g24660(.dina(n24917), .dinb(n10328), .dout(n24918));
  jxor g24661(.dina(n24243), .dinb(n11347), .dout(n24919));
  jor  g24662(.dina(n24919), .dinb(n24856), .dout(n24920));
  jxor g24663(.dina(n24920), .dinb(n24249), .dout(n24921));
  jand g24664(.dina(n24921), .dinb(n10824), .dout(n24922));
  jxor g24665(.dina(n24227), .dinb(n12410), .dout(n24923));
  jor  g24666(.dina(n24923), .dinb(n24856), .dout(n24924));
  jxor g24667(.dina(n24924), .dinb(n24233), .dout(n24925));
  jor  g24668(.dina(n24925), .dinb(n11858), .dout(n24926));
  jxor g24669(.dina(n24220), .dinb(n12947), .dout(n24927));
  jor  g24670(.dina(n24927), .dinb(n24856), .dout(n24928));
  jxor g24671(.dina(n24928), .dinb(n24225), .dout(n24929));
  jand g24672(.dina(n24929), .dinb(n12410), .dout(n24930));
  jxor g24673(.dina(n24196), .dinb(n14674), .dout(n24931));
  jor  g24674(.dina(n24931), .dinb(n24856), .dout(n24932));
  jxor g24675(.dina(n24932), .dinb(n24202), .dout(n24933));
  jor  g24676(.dina(n24933), .dinb(n14078), .dout(n24934));
  jxor g24677(.dina(n24189), .dinb(n15260), .dout(n24935));
  jor  g24678(.dina(n24935), .dinb(n24856), .dout(n24936));
  jxor g24679(.dina(n24936), .dinb(n24194), .dout(n24937));
  jor  g24680(.dina(n24937), .dinb(n14674), .dout(n24938));
  jxor g24681(.dina(n24174), .dinb(n16489), .dout(n24939));
  jor  g24682(.dina(n24939), .dinb(n24856), .dout(n24940));
  jxor g24683(.dina(n24940), .dinb(n24179), .dout(n24941));
  jor  g24684(.dina(n24941), .dinb(n15878), .dout(n24942));
  jxor g24685(.dina(n24166), .dinb(n17134), .dout(n24943));
  jor  g24686(.dina(n24943), .dinb(n24856), .dout(n24944));
  jxor g24687(.dina(n24944), .dinb(n24172), .dout(n24945));
  jor  g24688(.dina(n24945), .dinb(n16489), .dout(n24946));
  jxor g24689(.dina(n24159), .dinb(n17769), .dout(n24947));
  jor  g24690(.dina(n24947), .dinb(n24856), .dout(n24948));
  jxor g24691(.dina(n24948), .dinb(n24164), .dout(n24949));
  jand g24692(.dina(n24949), .dinb(n17134), .dout(n24950));
  jxor g24693(.dina(n24137), .dinb(n19791), .dout(n24951));
  jor  g24694(.dina(n24951), .dinb(n24856), .dout(n24952));
  jxor g24695(.dina(n24952), .dinb(n24143), .dout(n24953));
  jor  g24696(.dina(n24953), .dinb(n19096), .dout(n24954));
  jand g24697(.dina(n24953), .dinb(n19096), .dout(n24955));
  jxor g24698(.dina(n24129), .dinb(n20468), .dout(n24956));
  jor  g24699(.dina(n24956), .dinb(n24856), .dout(n24957));
  jxor g24700(.dina(n24957), .dinb(n24135), .dout(n24958));
  jor  g24701(.dina(n24958), .dinb(n19791), .dout(n24959));
  jxor g24702(.dina(n24122), .dinb(n21184), .dout(n24960));
  jor  g24703(.dina(n24960), .dinb(n24856), .dout(n24961));
  jxor g24704(.dina(n24961), .dinb(n24127), .dout(n24962));
  jor  g24705(.dina(n24962), .dinb(n20468), .dout(n24963));
  jxor g24706(.dina(n24115), .dinb(n21887), .dout(n24964));
  jor  g24707(.dina(n24964), .dinb(n24856), .dout(n24965));
  jxor g24708(.dina(n24965), .dinb(n24120), .dout(n24966));
  jor  g24709(.dina(n24966), .dinb(n21184), .dout(n24967));
  jand g24710(.dina(asqrt[1] ), .dinb(n23810), .dout(n24968));
  jand g24711(.dina(n24856), .dinb(asqrt[2] ), .dout(n24969));
  jor  g24712(.dina(n24969), .dinb(n24968), .dout(n24970));
  jxor g24713(.dina(n24970), .dinb(a[4] ), .dout(n24971));
  jor  g24714(.dina(n24971), .dinb(n23345), .dout(n24972));
  jnot g24715(.din(a[2] ), .dout(n24973));
  jor  g24716(.dina(a[1] ), .dinb(a[0] ), .dout(n24974));
  jand g24717(.dina(n24974), .dinb(n24973), .dout(n24975));
  jand g24718(.dina(n24856), .dinb(a[2] ), .dout(n24976));
  jor  g24719(.dina(n24976), .dinb(n24975), .dout(n24977));
  jor  g24720(.dina(n24977), .dinb(n24103), .dout(n24978));
  jand g24721(.dina(n24977), .dinb(n24103), .dout(n24979));
  jor  g24722(.dina(n24856), .dinb(a[2] ), .dout(n24980));
  jand g24723(.dina(n24980), .dinb(a[3] ), .dout(n24981));
  jor  g24724(.dina(n24981), .dinb(n24968), .dout(n24982));
  jor  g24725(.dina(n24982), .dinb(n24979), .dout(n24983));
  jand g24726(.dina(n24983), .dinb(n24978), .dout(n24984));
  jand g24727(.dina(n24984), .dinb(n24972), .dout(n24985));
  jxor g24728(.dina(n23812), .dinb(n23345), .dout(n24986));
  jor  g24729(.dina(n24986), .dinb(n24856), .dout(n24987));
  jxor g24730(.dina(n24987), .dinb(n24105), .dout(n24988));
  jand g24731(.dina(n24988), .dinb(n22620), .dout(n24989));
  jand g24732(.dina(n24971), .dinb(n23345), .dout(n24990));
  jor  g24733(.dina(n24990), .dinb(n24989), .dout(n24991));
  jor  g24734(.dina(n24991), .dinb(n24985), .dout(n24992));
  jxor g24735(.dina(n24107), .dinb(n22620), .dout(n24993));
  jor  g24736(.dina(n24993), .dinb(n24856), .dout(n24994));
  jxor g24737(.dina(n24994), .dinb(n24113), .dout(n24995));
  jor  g24738(.dina(n24995), .dinb(n21887), .dout(n24996));
  jor  g24739(.dina(n24988), .dinb(n22620), .dout(n24997));
  jand g24740(.dina(n24997), .dinb(n24996), .dout(n24998));
  jand g24741(.dina(n24998), .dinb(n24992), .dout(n24999));
  jand g24742(.dina(n24966), .dinb(n21184), .dout(n25000));
  jand g24743(.dina(n24995), .dinb(n21887), .dout(n25001));
  jor  g24744(.dina(n25001), .dinb(n25000), .dout(n25002));
  jor  g24745(.dina(n25002), .dinb(n24999), .dout(n25003));
  jand g24746(.dina(n25003), .dinb(n24967), .dout(n25004));
  jand g24747(.dina(n25004), .dinb(n24963), .dout(n25005));
  jand g24748(.dina(n24962), .dinb(n20468), .dout(n25006));
  jand g24749(.dina(n24958), .dinb(n19791), .dout(n25007));
  jor  g24750(.dina(n25007), .dinb(n25006), .dout(n25008));
  jor  g24751(.dina(n25008), .dinb(n25005), .dout(n25009));
  jand g24752(.dina(n25009), .dinb(n24959), .dout(n25010));
  jor  g24753(.dina(n25010), .dinb(n24955), .dout(n25011));
  jxor g24754(.dina(n24145), .dinb(n19096), .dout(n25012));
  jor  g24755(.dina(n25012), .dinb(n24856), .dout(n25013));
  jxor g24756(.dina(n25013), .dinb(n24150), .dout(n25014));
  jor  g24757(.dina(n25014), .dinb(n18442), .dout(n25015));
  jand g24758(.dina(n25015), .dinb(n25011), .dout(n25016));
  jand g24759(.dina(n25016), .dinb(n24954), .dout(n25017));
  jand g24760(.dina(n25014), .dinb(n18442), .dout(n25018));
  jxor g24761(.dina(n24152), .dinb(n18442), .dout(n25019));
  jor  g24762(.dina(n25019), .dinb(n24856), .dout(n25020));
  jxor g24763(.dina(n25020), .dinb(n24157), .dout(n25021));
  jand g24764(.dina(n25021), .dinb(n17769), .dout(n25022));
  jor  g24765(.dina(n25022), .dinb(n25018), .dout(n25023));
  jor  g24766(.dina(n25023), .dinb(n25017), .dout(n25024));
  jor  g24767(.dina(n25021), .dinb(n17769), .dout(n25025));
  jor  g24768(.dina(n24949), .dinb(n17134), .dout(n25026));
  jand g24769(.dina(n25026), .dinb(n25025), .dout(n25027));
  jand g24770(.dina(n25027), .dinb(n25024), .dout(n25028));
  jor  g24771(.dina(n25028), .dinb(n24950), .dout(n25029));
  jand g24772(.dina(n25029), .dinb(n24946), .dout(n25030));
  jand g24773(.dina(n24945), .dinb(n16489), .dout(n25031));
  jand g24774(.dina(n24941), .dinb(n15878), .dout(n25032));
  jor  g24775(.dina(n25032), .dinb(n25031), .dout(n25033));
  jor  g24776(.dina(n25033), .dinb(n25030), .dout(n25034));
  jxor g24777(.dina(n24181), .dinb(n15878), .dout(n25035));
  jor  g24778(.dina(n25035), .dinb(n24856), .dout(n25036));
  jxor g24779(.dina(n25036), .dinb(n24187), .dout(n25037));
  jor  g24780(.dina(n25037), .dinb(n15260), .dout(n25038));
  jand g24781(.dina(n25038), .dinb(n25034), .dout(n25039));
  jand g24782(.dina(n25039), .dinb(n24942), .dout(n25040));
  jand g24783(.dina(n25037), .dinb(n15260), .dout(n25041));
  jand g24784(.dina(n24937), .dinb(n14674), .dout(n25042));
  jor  g24785(.dina(n25042), .dinb(n25041), .dout(n25043));
  jor  g24786(.dina(n25043), .dinb(n25040), .dout(n25044));
  jand g24787(.dina(n25044), .dinb(n24938), .dout(n25045));
  jand g24788(.dina(n24933), .dinb(n14078), .dout(n25046));
  jor  g24789(.dina(n25046), .dinb(n25045), .dout(n25047));
  jxor g24790(.dina(n24204), .dinb(n14078), .dout(n25048));
  jor  g24791(.dina(n25048), .dinb(n24856), .dout(n25049));
  jxor g24792(.dina(n25049), .dinb(n24210), .dout(n25050));
  jor  g24793(.dina(n25050), .dinb(n13515), .dout(n25051));
  jand g24794(.dina(n25051), .dinb(n25047), .dout(n25052));
  jand g24795(.dina(n25052), .dinb(n24934), .dout(n25053));
  jand g24796(.dina(n25050), .dinb(n13515), .dout(n25054));
  jxor g24797(.dina(n24212), .dinb(n13515), .dout(n25055));
  jor  g24798(.dina(n25055), .dinb(n24856), .dout(n25056));
  jxor g24799(.dina(n25056), .dinb(n24218), .dout(n25057));
  jand g24800(.dina(n25057), .dinb(n12947), .dout(n25058));
  jor  g24801(.dina(n25058), .dinb(n25054), .dout(n25059));
  jor  g24802(.dina(n25059), .dinb(n25053), .dout(n25060));
  jor  g24803(.dina(n24929), .dinb(n12410), .dout(n25061));
  jor  g24804(.dina(n25057), .dinb(n12947), .dout(n25062));
  jand g24805(.dina(n25062), .dinb(n25061), .dout(n25063));
  jand g24806(.dina(n25063), .dinb(n25060), .dout(n25064));
  jor  g24807(.dina(n25064), .dinb(n24930), .dout(n25065));
  jand g24808(.dina(n25065), .dinb(n24926), .dout(n25066));
  jand g24809(.dina(n24925), .dinb(n11858), .dout(n25067));
  jxor g24810(.dina(n24235), .dinb(n11858), .dout(n25068));
  jor  g24811(.dina(n25068), .dinb(n24856), .dout(n25069));
  jxor g24812(.dina(n25069), .dinb(n24241), .dout(n25070));
  jand g24813(.dina(n25070), .dinb(n11347), .dout(n25071));
  jor  g24814(.dina(n25071), .dinb(n25067), .dout(n25072));
  jor  g24815(.dina(n25072), .dinb(n25066), .dout(n25073));
  jor  g24816(.dina(n25070), .dinb(n11347), .dout(n25074));
  jor  g24817(.dina(n24921), .dinb(n10824), .dout(n25075));
  jand g24818(.dina(n25075), .dinb(n25074), .dout(n25076));
  jand g24819(.dina(n25076), .dinb(n25073), .dout(n25077));
  jor  g24820(.dina(n25077), .dinb(n24922), .dout(n25078));
  jor  g24821(.dina(n24917), .dinb(n10328), .dout(n25079));
  jand g24822(.dina(n25079), .dinb(n25078), .dout(n25080));
  jxor g24823(.dina(n24258), .dinb(n10328), .dout(n25081));
  jor  g24824(.dina(n25081), .dinb(n24856), .dout(n25082));
  jxor g24825(.dina(n25082), .dinb(n24264), .dout(n25083));
  jand g24826(.dina(n25083), .dinb(n9832), .dout(n25084));
  jor  g24827(.dina(n25084), .dinb(n25080), .dout(n25085));
  jor  g24828(.dina(n25085), .dinb(n24918), .dout(n25086));
  jor  g24829(.dina(n25083), .dinb(n9832), .dout(n25087));
  jxor g24830(.dina(n24266), .dinb(n9832), .dout(n25088));
  jor  g24831(.dina(n25088), .dinb(n24856), .dout(n25089));
  jxor g24832(.dina(n25089), .dinb(n24271), .dout(n25090));
  jor  g24833(.dina(n25090), .dinb(n9369), .dout(n25091));
  jand g24834(.dina(n25091), .dinb(n25087), .dout(n25092));
  jand g24835(.dina(n25092), .dinb(n25086), .dout(n25093));
  jand g24836(.dina(n25090), .dinb(n9369), .dout(n25094));
  jxor g24837(.dina(n24273), .dinb(n9369), .dout(n25095));
  jor  g24838(.dina(n25095), .dinb(n24856), .dout(n25096));
  jxor g24839(.dina(n25096), .dinb(n24279), .dout(n25097));
  jand g24840(.dina(n25097), .dinb(n8890), .dout(n25098));
  jor  g24841(.dina(n25098), .dinb(n25094), .dout(n25099));
  jor  g24842(.dina(n25099), .dinb(n25093), .dout(n25100));
  jor  g24843(.dina(n25097), .dinb(n8890), .dout(n25101));
  jand g24844(.dina(n25101), .dinb(n25100), .dout(n25102));
  jand g24845(.dina(n24913), .dinb(n8449), .dout(n25103));
  jor  g24846(.dina(n25103), .dinb(n25102), .dout(n25104));
  jor  g24847(.dina(n24909), .dinb(n8003), .dout(n25105));
  jand g24848(.dina(n25105), .dinb(n25104), .dout(n25106));
  jand g24849(.dina(n25106), .dinb(n24914), .dout(n25107));
  jor  g24850(.dina(n25107), .dinb(n24910), .dout(n25108));
  jor  g24851(.dina(n24905), .dinb(n7581), .dout(n25109));
  jand g24852(.dina(n25109), .dinb(n25108), .dout(n25110));
  jxor g24853(.dina(n24304), .dinb(n7581), .dout(n25111));
  jor  g24854(.dina(n25111), .dinb(n24856), .dout(n25112));
  jxor g24855(.dina(n25112), .dinb(n24309), .dout(n25113));
  jand g24856(.dina(n25113), .dinb(n7154), .dout(n25114));
  jor  g24857(.dina(n25114), .dinb(n25110), .dout(n25115));
  jor  g24858(.dina(n25115), .dinb(n24906), .dout(n25116));
  jxor g24859(.dina(n24311), .dinb(n7154), .dout(n25117));
  jor  g24860(.dina(n25117), .dinb(n24856), .dout(n25118));
  jxor g24861(.dina(n25118), .dinb(n24316), .dout(n25119));
  jor  g24862(.dina(n25119), .dinb(n6758), .dout(n25120));
  jor  g24863(.dina(n25113), .dinb(n7154), .dout(n25121));
  jand g24864(.dina(n25121), .dinb(n25120), .dout(n25122));
  jand g24865(.dina(n25122), .dinb(n25116), .dout(n25123));
  jand g24866(.dina(n25119), .dinb(n6758), .dout(n25124));
  jand g24867(.dina(n24901), .dinb(n6357), .dout(n25125));
  jor  g24868(.dina(n25125), .dinb(n25124), .dout(n25126));
  jor  g24869(.dina(n25126), .dinb(n25123), .dout(n25127));
  jxor g24870(.dina(n24326), .dinb(n6357), .dout(n25128));
  jor  g24871(.dina(n25128), .dinb(n24856), .dout(n25129));
  jxor g24872(.dina(n25129), .dinb(n24331), .dout(n25130));
  jor  g24873(.dina(n25130), .dinb(n5989), .dout(n25131));
  jand g24874(.dina(n25131), .dinb(n25127), .dout(n25132));
  jand g24875(.dina(n25132), .dinb(n24902), .dout(n25133));
  jand g24876(.dina(n25130), .dinb(n5989), .dout(n25134));
  jxor g24877(.dina(n24333), .dinb(n5989), .dout(n25135));
  jor  g24878(.dina(n25135), .dinb(n24856), .dout(n25136));
  jxor g24879(.dina(n25136), .dinb(n24339), .dout(n25137));
  jand g24880(.dina(n25137), .dinb(n5606), .dout(n25138));
  jor  g24881(.dina(n25138), .dinb(n25134), .dout(n25139));
  jor  g24882(.dina(n25139), .dinb(n25133), .dout(n25140));
  jxor g24883(.dina(n24341), .dinb(n5606), .dout(n25141));
  jor  g24884(.dina(n25141), .dinb(n24856), .dout(n25142));
  jxor g24885(.dina(n25142), .dinb(n24346), .dout(n25143));
  jor  g24886(.dina(n25143), .dinb(n5259), .dout(n25144));
  jor  g24887(.dina(n25137), .dinb(n5606), .dout(n25145));
  jand g24888(.dina(n25145), .dinb(n25144), .dout(n25146));
  jand g24889(.dina(n25146), .dinb(n25140), .dout(n25147));
  jand g24890(.dina(n25143), .dinb(n5259), .dout(n25148));
  jxor g24891(.dina(n24348), .dinb(n5259), .dout(n25149));
  jor  g24892(.dina(n25149), .dinb(n24856), .dout(n25150));
  jxor g24893(.dina(n25150), .dinb(n24354), .dout(n25151));
  jand g24894(.dina(n25151), .dinb(n4902), .dout(n25152));
  jor  g24895(.dina(n25152), .dinb(n25148), .dout(n25153));
  jor  g24896(.dina(n25153), .dinb(n25147), .dout(n25154));
  jor  g24897(.dina(n25151), .dinb(n4902), .dout(n25155));
  jor  g24898(.dina(n24897), .dinb(n4582), .dout(n25156));
  jand g24899(.dina(n25156), .dinb(n25155), .dout(n25157));
  jand g24900(.dina(n25157), .dinb(n25154), .dout(n25158));
  jor  g24901(.dina(n25158), .dinb(n24898), .dout(n25159));
  jand g24902(.dina(n25159), .dinb(n24894), .dout(n25160));
  jand g24903(.dina(n24893), .dinb(n4249), .dout(n25161));
  jxor g24904(.dina(n24372), .dinb(n4249), .dout(n25162));
  jor  g24905(.dina(n25162), .dinb(n24856), .dout(n25163));
  jxor g24906(.dina(n25163), .dinb(n24377), .dout(n25164));
  jand g24907(.dina(n25164), .dinb(n3955), .dout(n25165));
  jor  g24908(.dina(n25165), .dinb(n25161), .dout(n25166));
  jor  g24909(.dina(n25166), .dinb(n25160), .dout(n25167));
  jor  g24910(.dina(n25164), .dinb(n3955), .dout(n25168));
  jxor g24911(.dina(n24379), .dinb(n3955), .dout(n25169));
  jor  g24912(.dina(n25169), .dinb(n24856), .dout(n25170));
  jxor g24913(.dina(n25170), .dinb(n24385), .dout(n25171));
  jor  g24914(.dina(n25171), .dinb(n3642), .dout(n25172));
  jand g24915(.dina(n25172), .dinb(n25168), .dout(n25173));
  jand g24916(.dina(n25173), .dinb(n25167), .dout(n25174));
  jand g24917(.dina(n25171), .dinb(n3642), .dout(n25175));
  jxor g24918(.dina(n24387), .dinb(n3642), .dout(n25176));
  jor  g24919(.dina(n25176), .dinb(n24856), .dout(n25177));
  jxor g24920(.dina(n25177), .dinb(n24392), .dout(n25178));
  jand g24921(.dina(n25178), .dinb(n3368), .dout(n25179));
  jor  g24922(.dina(n25179), .dinb(n25175), .dout(n25180));
  jor  g24923(.dina(n25180), .dinb(n25174), .dout(n25181));
  jor  g24924(.dina(n25178), .dinb(n3368), .dout(n25182));
  jor  g24925(.dina(n24889), .dinb(n3089), .dout(n25183));
  jand g24926(.dina(n25183), .dinb(n25182), .dout(n25184));
  jand g24927(.dina(n25184), .dinb(n25181), .dout(n25185));
  jor  g24928(.dina(n25185), .dinb(n24890), .dout(n25186));
  jxor g24929(.dina(n24402), .dinb(n3089), .dout(n25187));
  jor  g24930(.dina(n25187), .dinb(n24856), .dout(n25188));
  jxor g24931(.dina(n25188), .dinb(n24407), .dout(n25189));
  jor  g24932(.dina(n25189), .dinb(n2833), .dout(n25190));
  jand g24933(.dina(n25190), .dinb(n25186), .dout(n25191));
  jand g24934(.dina(n25189), .dinb(n2833), .dout(n25192));
  jxor g24935(.dina(n24409), .dinb(n2833), .dout(n25193));
  jor  g24936(.dina(n25193), .dinb(n24856), .dout(n25194));
  jxor g24937(.dina(n25194), .dinb(n24415), .dout(n25195));
  jand g24938(.dina(n25195), .dinb(n2572), .dout(n25196));
  jor  g24939(.dina(n25196), .dinb(n25192), .dout(n25197));
  jor  g24940(.dina(n25197), .dinb(n25191), .dout(n25198));
  jor  g24941(.dina(n25195), .dinb(n2572), .dout(n25199));
  jor  g24942(.dina(n24885), .dinb(n2345), .dout(n25200));
  jand g24943(.dina(n25200), .dinb(n25199), .dout(n25201));
  jand g24944(.dina(n25201), .dinb(n25198), .dout(n25202));
  jor  g24945(.dina(n25202), .dinb(n24886), .dout(n25203));
  jand g24946(.dina(n25203), .dinb(n24882), .dout(n25204));
  jand g24947(.dina(n24881), .dinb(n2108), .dout(n25205));
  jxor g24948(.dina(n24432), .dinb(n2108), .dout(n25206));
  jor  g24949(.dina(n25206), .dinb(n24856), .dout(n25207));
  jxor g24950(.dina(n25207), .dinb(n24438), .dout(n25208));
  jand g24951(.dina(n25208), .dinb(n1912), .dout(n25209));
  jor  g24952(.dina(n25209), .dinb(n25205), .dout(n25210));
  jor  g24953(.dina(n25210), .dinb(n25204), .dout(n25211));
  jor  g24954(.dina(n25208), .dinb(n1912), .dout(n25212));
  jxor g24955(.dina(n24440), .dinb(n1912), .dout(n25213));
  jor  g24956(.dina(n25213), .dinb(n24856), .dout(n25214));
  jxor g24957(.dina(n25214), .dinb(n24446), .dout(n25215));
  jor  g24958(.dina(n25215), .dinb(n1699), .dout(n25216));
  jand g24959(.dina(n25216), .dinb(n25212), .dout(n25217));
  jand g24960(.dina(n25217), .dinb(n25211), .dout(n25218));
  jand g24961(.dina(n25215), .dinb(n1699), .dout(n25219));
  jxor g24962(.dina(n24448), .dinb(n1699), .dout(n25220));
  jor  g24963(.dina(n25220), .dinb(n24856), .dout(n25221));
  jxor g24964(.dina(n25221), .dinb(n24453), .dout(n25222));
  jand g24965(.dina(n25222), .dinb(n1516), .dout(n25223));
  jor  g24966(.dina(n25223), .dinb(n25219), .dout(n25224));
  jor  g24967(.dina(n25224), .dinb(n25218), .dout(n25225));
  jor  g24968(.dina(n25222), .dinb(n1516), .dout(n25226));
  jor  g24969(.dina(n24877), .dinb(n1332), .dout(n25227));
  jand g24970(.dina(n25227), .dinb(n25226), .dout(n25228));
  jand g24971(.dina(n25228), .dinb(n25225), .dout(n25229));
  jor  g24972(.dina(n25229), .dinb(n24878), .dout(n25230));
  jor  g24973(.dina(n24873), .dinb(n1173), .dout(n25231));
  jand g24974(.dina(n25231), .dinb(n25230), .dout(n25232));
  jxor g24975(.dina(n24471), .dinb(n1173), .dout(n25233));
  jor  g24976(.dina(n25233), .dinb(n24856), .dout(n25234));
  jxor g24977(.dina(n25234), .dinb(n24477), .dout(n25235));
  jand g24978(.dina(n25235), .dinb(n1008), .dout(n25236));
  jor  g24979(.dina(n25236), .dinb(n25232), .dout(n25237));
  jor  g24980(.dina(n25237), .dinb(n24874), .dout(n25238));
  jor  g24981(.dina(n25235), .dinb(n1008), .dout(n25239));
  jor  g24982(.dina(n24867), .dinb(n884), .dout(n25240));
  jand g24983(.dina(n25240), .dinb(n25239), .dout(n25241));
  jand g24984(.dina(n25241), .dinb(n25238), .dout(n25242));
  jor  g24985(.dina(n25242), .dinb(n24870), .dout(n25243));
  jxor g24986(.dina(n24495), .dinb(n743), .dout(n25244));
  jor  g24987(.dina(n25244), .dinb(n24856), .dout(n25245));
  jxor g24988(.dina(n25245), .dinb(n24500), .dout(n25246));
  jor  g24989(.dina(n25246), .dinb(n635), .dout(n25247));
  jand g24990(.dina(n25247), .dinb(n25243), .dout(n25248));
  jand g24991(.dina(n25248), .dinb(n24864), .dout(n25249));
  jand g24992(.dina(n25246), .dinb(n635), .dout(n25250));
  jxor g24993(.dina(n24502), .dinb(n635), .dout(n25251));
  jor  g24994(.dina(n25251), .dinb(n24856), .dout(n25252));
  jxor g24995(.dina(n25252), .dinb(n24508), .dout(n25253));
  jand g24996(.dina(n25253), .dinb(n515), .dout(n25254));
  jor  g24997(.dina(n25254), .dinb(n25250), .dout(n25255));
  jor  g24998(.dina(n25255), .dinb(n25249), .dout(n25256));
  jor  g24999(.dina(n25253), .dinb(n515), .dout(n25257));
  jxor g25000(.dina(n24510), .dinb(n515), .dout(n25258));
  jor  g25001(.dina(n25258), .dinb(n24856), .dout(n25259));
  jxor g25002(.dina(n25259), .dinb(n24515), .dout(n25260));
  jor  g25003(.dina(n25260), .dinb(n443), .dout(n25261));
  jand g25004(.dina(n25261), .dinb(n25257), .dout(n25262));
  jand g25005(.dina(n25262), .dinb(n25256), .dout(n25263));
  jand g25006(.dina(n25260), .dinb(n443), .dout(n25264));
  jxor g25007(.dina(n24517), .dinb(n443), .dout(n25265));
  jor  g25008(.dina(n25265), .dinb(n24856), .dout(n25266));
  jxor g25009(.dina(n25266), .dinb(n24523), .dout(n25267));
  jand g25010(.dina(n25267), .dinb(n352), .dout(n25268));
  jor  g25011(.dina(n25268), .dinb(n25264), .dout(n25269));
  jor  g25012(.dina(n25269), .dinb(n25263), .dout(n25270));
  jxor g25013(.dina(n24525), .dinb(n352), .dout(n25271));
  jor  g25014(.dina(n25271), .dinb(n24856), .dout(n25272));
  jxor g25015(.dina(n25272), .dinb(n24530), .dout(n25273));
  jor  g25016(.dina(n25273), .dinb(n294), .dout(n25274));
  jor  g25017(.dina(n25267), .dinb(n352), .dout(n25275));
  jand g25018(.dina(n25275), .dinb(n25274), .dout(n25276));
  jand g25019(.dina(n25276), .dinb(n25270), .dout(n25277));
  jand g25020(.dina(n25273), .dinb(n294), .dout(n25278));
  jxor g25021(.dina(n24532), .dinb(n294), .dout(n25279));
  jor  g25022(.dina(n25279), .dinb(n24856), .dout(n25280));
  jxor g25023(.dina(n25280), .dinb(n24537), .dout(n25281));
  jand g25024(.dina(n25281), .dinb(n239), .dout(n25282));
  jor  g25025(.dina(n25282), .dinb(n25278), .dout(n25283));
  jor  g25026(.dina(n25283), .dinb(n25277), .dout(n25284));
  jor  g25027(.dina(n25281), .dinb(n239), .dout(n25285));
  jor  g25028(.dina(n24859), .dinb(n221), .dout(n25286));
  jand g25029(.dina(n25286), .dinb(n25285), .dout(n25287));
  jand g25030(.dina(n25287), .dinb(n25284), .dout(n25288));
  jor  g25031(.dina(n25288), .dinb(n24860), .dout(n25289));
  jxor g25032(.dina(n24546), .dinb(n221), .dout(n25290));
  jor  g25033(.dina(n25290), .dinb(n24856), .dout(n25291));
  jxor g25034(.dina(n25291), .dinb(n24552), .dout(n25292));
  jor  g25035(.dina(n25292), .dinb(n218), .dout(n25293));
  jand g25036(.dina(n25293), .dinb(n25289), .dout(n25294));
  jand g25037(.dina(asqrt[1] ), .dinb(n24852), .dout(n25295));
  jnot g25038(.din(n24835), .dout(n25296));
  jor  g25039(.dina(n25292), .dinb(n25296), .dout(n25297));
  jor  g25040(.dina(n25297), .dinb(n25295), .dout(n25298));
  jand g25041(.dina(n25298), .dinb(n218), .dout(n25299));
  jor  g25042(.dina(n25299), .dinb(n25294), .dout(n25300));
  jor  g25043(.dina(n25300), .dinb(n24850), .dout(asqrt[0] ));
endmodule


