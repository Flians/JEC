/*
rf_c1908:
	jxor: 74
	jspl: 106
	jspl3: 95
	jnot: 41
	jdff: 1045
	jand: 128
	jor: 102

Summary:
	jxor: 74
	jspl: 106
	jspl3: 95
	jnot: 41
	jdff: 1045
	jand: 128
	jor: 102

The maximum logic level gap of any gate:
	rf_c1908: 17
*/

module rf_c1908(gclk, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57);
	input gclk;
	input G101;
	input G104;
	input G107;
	input G110;
	input G113;
	input G116;
	input G119;
	input G122;
	input G125;
	input G128;
	input G131;
	input G134;
	input G137;
	input G140;
	input G143;
	input G146;
	input G210;
	input G214;
	input G217;
	input G221;
	input G224;
	input G227;
	input G234;
	input G237;
	input G469;
	input G472;
	input G475;
	input G478;
	input G898;
	input G900;
	input G902;
	input G952;
	input G953;
	output G3;
	output G6;
	output G9;
	output G12;
	output G30;
	output G45;
	output G48;
	output G15;
	output G18;
	output G21;
	output G24;
	output G27;
	output G33;
	output G36;
	output G39;
	output G42;
	output G75;
	output G51;
	output G54;
	output G60;
	output G63;
	output G66;
	output G69;
	output G72;
	output G57;
	wire n58;
	wire n59;
	wire n60;
	wire n61;
	wire n62;
	wire n63;
	wire n64;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n69;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n188;
	wire n189;
	wire n190;
	wire n192;
	wire n193;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n202;
	wire n204;
	wire n205;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n212;
	wire n213;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n222;
	wire n224;
	wire n225;
	wire n226;
	wire n228;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire [2:0] w_G101_0;
	wire [2:0] w_G104_0;
	wire [2:0] w_G107_0;
	wire [2:0] w_G110_0;
	wire [1:0] w_G110_1;
	wire [1:0] w_G113_0;
	wire [2:0] w_G116_0;
	wire [2:0] w_G119_0;
	wire [2:0] w_G122_0;
	wire [1:0] w_G122_1;
	wire [2:0] w_G125_0;
	wire [2:0] w_G128_0;
	wire [1:0] w_G128_1;
	wire [1:0] w_G131_0;
	wire [2:0] w_G134_0;
	wire [2:0] w_G137_0;
	wire [2:0] w_G140_0;
	wire [2:0] w_G143_0;
	wire [1:0] w_G143_1;
	wire [2:0] w_G146_0;
	wire [2:0] w_G210_0;
	wire [1:0] w_G214_0;
	wire [2:0] w_G217_0;
	wire [1:0] w_G221_0;
	wire [1:0] w_G224_0;
	wire [1:0] w_G227_0;
	wire [2:0] w_G234_0;
	wire [2:0] w_G237_0;
	wire [2:0] w_G469_0;
	wire [1:0] w_G472_0;
	wire [2:0] w_G475_0;
	wire [2:0] w_G478_0;
	wire [2:0] w_G902_0;
	wire [2:0] w_G902_1;
	wire [2:0] w_G902_2;
	wire [2:0] w_G902_3;
	wire [2:0] w_G952_0;
	wire [2:0] w_G953_0;
	wire [2:0] w_G953_1;
	wire [1:0] w_n59_0;
	wire [2:0] w_n60_0;
	wire [2:0] w_n61_0;
	wire [2:0] w_n61_1;
	wire [2:0] w_n61_2;
	wire [2:0] w_n61_3;
	wire [1:0] w_n62_0;
	wire [1:0] w_n67_0;
	wire [1:0] w_n68_0;
	wire [2:0] w_n70_0;
	wire [2:0] w_n70_1;
	wire [2:0] w_n70_2;
	wire [1:0] w_n70_3;
	wire [1:0] w_n71_0;
	wire [1:0] w_n73_0;
	wire [2:0] w_n74_0;
	wire [1:0] w_n74_1;
	wire [1:0] w_n77_0;
	wire [1:0] w_n79_0;
	wire [2:0] w_n81_0;
	wire [1:0] w_n82_0;
	wire [1:0] w_n84_0;
	wire [1:0] w_n86_0;
	wire [2:0] w_n90_0;
	wire [2:0] w_n92_0;
	wire [2:0] w_n92_1;
	wire [2:0] w_n93_0;
	wire [1:0] w_n94_0;
	wire [2:0] w_n95_0;
	wire [2:0] w_n96_0;
	wire [1:0] w_n97_0;
	wire [1:0] w_n101_0;
	wire [1:0] w_n103_0;
	wire [2:0] w_n107_0;
	wire [1:0] w_n108_0;
	wire [1:0] w_n109_0;
	wire [2:0] w_n110_0;
	wire [2:0] w_n112_0;
	wire [1:0] w_n112_1;
	wire [2:0] w_n117_0;
	wire [1:0] w_n118_0;
	wire [1:0] w_n119_0;
	wire [1:0] w_n120_0;
	wire [2:0] w_n121_0;
	wire [1:0] w_n121_1;
	wire [1:0] w_n122_0;
	wire [2:0] w_n130_0;
	wire [1:0] w_n131_0;
	wire [2:0] w_n132_0;
	wire [2:0] w_n141_0;
	wire [1:0] w_n142_0;
	wire [2:0] w_n143_0;
	wire [1:0] w_n143_1;
	wire [2:0] w_n144_0;
	wire [2:0] w_n144_1;
	wire [1:0] w_n145_0;
	wire [1:0] w_n146_0;
	wire [1:0] w_n147_0;
	wire [2:0] w_n151_0;
	wire [1:0] w_n152_0;
	wire [2:0] w_n153_0;
	wire [2:0] w_n154_0;
	wire [1:0] w_n154_1;
	wire [2:0] w_n155_0;
	wire [1:0] w_n156_0;
	wire [2:0] w_n158_0;
	wire [1:0] w_n158_1;
	wire [2:0] w_n159_0;
	wire [1:0] w_n159_1;
	wire [1:0] w_n160_0;
	wire [2:0] w_n161_0;
	wire [1:0] w_n162_0;
	wire [2:0] w_n163_0;
	wire [1:0] w_n164_0;
	wire [2:0] w_n166_0;
	wire [1:0] w_n166_1;
	wire [1:0] w_n167_0;
	wire [2:0] w_n168_0;
	wire [1:0] w_n169_0;
	wire [1:0] w_n172_0;
	wire [2:0] w_n174_0;
	wire [1:0] w_n174_1;
	wire [1:0] w_n175_0;
	wire [1:0] w_n177_0;
	wire [2:0] w_n179_0;
	wire [1:0] w_n180_0;
	wire [2:0] w_n181_0;
	wire [2:0] w_n183_0;
	wire [2:0] w_n184_0;
	wire [1:0] w_n184_1;
	wire [2:0] w_n185_0;
	wire [1:0] w_n186_0;
	wire [2:0] w_n188_0;
	wire [1:0] w_n189_0;
	wire [1:0] w_n190_0;
	wire [2:0] w_n192_0;
	wire [1:0] w_n193_0;
	wire [2:0] w_n196_0;
	wire [2:0] w_n197_0;
	wire [1:0] w_n197_1;
	wire [2:0] w_n198_0;
	wire [1:0] w_n198_1;
	wire [1:0] w_n199_0;
	wire [1:0] w_n200_0;
	wire [1:0] w_n202_0;
	wire [1:0] w_n205_0;
	wire [1:0] w_n207_0;
	wire [1:0] w_n210_0;
	wire [1:0] w_n212_0;
	wire [1:0] w_n213_0;
	wire [2:0] w_n216_0;
	wire [2:0] w_n217_0;
	wire [2:0] w_n218_0;
	wire [1:0] w_n218_1;
	wire [1:0] w_n219_0;
	wire [1:0] w_n220_0;
	wire [1:0] w_n222_0;
	wire [1:0] w_n226_0;
	wire [1:0] w_n228_0;
	wire [2:0] w_n244_0;
	wire [2:0] w_n244_1;
	wire [2:0] w_n244_2;
	wire [1:0] w_n252_0;
	wire [2:0] w_n253_0;
	wire [2:0] w_n254_0;
	wire [1:0] w_n254_1;
	wire [2:0] w_n273_0;
	wire [1:0] w_n274_0;
	wire [1:0] w_n275_0;
	wire [2:0] w_n276_0;
	wire [1:0] w_n276_1;
	wire [1:0] w_n277_0;
	wire [1:0] w_n278_0;
	wire [1:0] w_n280_0;
	wire [2:0] w_n281_0;
	wire [1:0] w_n282_0;
	wire [1:0] w_n286_0;
	wire [2:0] w_n288_0;
	wire [1:0] w_n289_0;
	wire [2:0] w_n290_0;
	wire [1:0] w_n291_0;
	wire [1:0] w_n295_0;
	wire [1:0] w_n308_0;
	wire [1:0] w_n309_0;
	wire [2:0] w_n311_0;
	wire [2:0] w_n314_0;
	wire [1:0] w_n315_0;
	wire [1:0] w_n318_0;
	wire [1:0] w_n325_0;
	wire [1:0] w_n334_0;
	wire [2:0] w_n335_0;
	wire [2:0] w_n335_1;
	wire [1:0] w_n335_2;
	wire [1:0] w_n336_0;
	wire [2:0] w_n340_0;
	wire [2:0] w_n340_1;
	wire [1:0] w_n340_2;
	wire [1:0] w_n346_0;
	wire [1:0] w_n355_0;
	wire [1:0] w_n364_0;
	wire [1:0] w_n372_0;
	wire [1:0] w_n395_0;
	wire w_dff_B_LWkzKn8m7_0;
	wire w_dff_B_Be0JuueW8_0;
	wire w_dff_B_feKD8TAg8_0;
	wire w_dff_B_lkPmwJSH6_0;
	wire w_dff_B_Dus5asfn5_0;
	wire w_dff_B_Mh6gqh832_0;
	wire w_dff_B_Iqg5cNID3_0;
	wire w_dff_B_WhPzckqG5_0;
	wire w_dff_B_Y1HlTLS96_1;
	wire w_dff_B_k74NkQxL3_1;
	wire w_dff_B_3oUgQuJh8_0;
	wire w_dff_B_cnGFPP2K6_0;
	wire w_dff_A_3ue1GCAa6_1;
	wire w_dff_B_pbGQtWSj8_2;
	wire w_dff_B_fXGOIhMh3_2;
	wire w_dff_B_1z3qikvk4_0;
	wire w_dff_B_OjrxPkoz1_0;
	wire w_dff_B_0NusGIpQ1_1;
	wire w_dff_B_hdCoarWM4_1;
	wire w_dff_B_DsJPWdlA2_1;
	wire w_dff_B_u0O1DsPH2_1;
	wire w_dff_B_JakKkpps1_1;
	wire w_dff_B_E6lrRoBW0_1;
	wire w_dff_B_VuZcRjQM4_1;
	wire w_dff_B_q5HVwXmD5_1;
	wire w_dff_B_13uuITfG2_1;
	wire w_dff_B_QL5mamIM6_1;
	wire w_dff_B_LnVkTcjl3_1;
	wire w_dff_B_8v4Z0UIu6_1;
	wire w_dff_B_7u0DeLhZ9_0;
	wire w_dff_B_lYykZK1E7_0;
	wire w_dff_B_fKrfXaD88_0;
	wire w_dff_B_wKbd32w60_0;
	wire w_dff_B_FuQIJ1E44_0;
	wire w_dff_B_H9cCylnh8_0;
	wire w_dff_B_uuXwp87y5_0;
	wire w_dff_B_WQ0cvmw84_0;
	wire w_dff_B_i2Ue4JlN0_0;
	wire w_dff_B_OXR17nlL7_0;
	wire w_dff_B_thlH4yks4_0;
	wire w_dff_B_mimsbmED9_0;
	wire w_dff_B_DzktRynN5_0;
	wire w_dff_B_dr0BwsTl6_0;
	wire w_dff_A_PWhc653A2_0;
	wire w_dff_A_T55N1r1Y9_0;
	wire w_dff_A_KFFnJt7d9_0;
	wire w_dff_A_s8VJWkIA8_0;
	wire w_dff_A_GwVN9RiE3_0;
	wire w_dff_A_jRpf3phO1_0;
	wire w_dff_A_E9kIB8ML0_0;
	wire w_dff_A_6So5Xe162_0;
	wire w_dff_A_vj5pcntQ1_0;
	wire w_dff_A_58eoaMGF4_0;
	wire w_dff_A_z9WPkE0c8_0;
	wire w_dff_A_Tns3PYmN2_0;
	wire w_dff_A_Xs4reAsg9_0;
	wire w_dff_A_yE2KYfAC7_0;
	wire w_dff_A_wK8xo0ih4_0;
	wire w_dff_B_ANQgRK140_1;
	wire w_dff_B_4EnfuEyv7_1;
	wire w_dff_B_Oro06xku4_1;
	wire w_dff_B_XzmnYfwm7_1;
	wire w_dff_B_o5wRrX1u5_1;
	wire w_dff_B_DOqRJtRL1_1;
	wire w_dff_B_RB58VdCH1_1;
	wire w_dff_B_CRDkqrFk2_1;
	wire w_dff_B_8GAmCsxX6_1;
	wire w_dff_B_Rd0PAMwQ7_1;
	wire w_dff_B_jV8dr14K4_1;
	wire w_dff_B_fuB4YbjP6_1;
	wire w_dff_B_74JaBsIo5_0;
	wire w_dff_B_euM955On1_0;
	wire w_dff_B_cQbWAykn8_0;
	wire w_dff_B_luXDGkTp1_0;
	wire w_dff_B_05lhf9A88_0;
	wire w_dff_B_sZFyscMk1_0;
	wire w_dff_B_1vOjhKA85_0;
	wire w_dff_B_E0OyvjAW3_0;
	wire w_dff_B_hPzftarw4_0;
	wire w_dff_B_9TK02zqz0_0;
	wire w_dff_B_zCSJrkjM3_0;
	wire w_dff_B_0eEjCKXP5_0;
	wire w_dff_B_b6LaWH4c2_0;
	wire w_dff_B_Hz6UxcGC4_0;
	wire w_dff_A_WHafdpbG5_0;
	wire w_dff_A_M81hBMB46_0;
	wire w_dff_A_mFIrA8nf3_0;
	wire w_dff_A_SKUTIPTp3_0;
	wire w_dff_A_ZUbskobr6_0;
	wire w_dff_A_FIT1i4QH2_0;
	wire w_dff_A_xWOzoEwx6_0;
	wire w_dff_A_SVMe4flY6_0;
	wire w_dff_A_J79ltrwf6_0;
	wire w_dff_A_mCJiZiea9_0;
	wire w_dff_A_2w90mkWU1_0;
	wire w_dff_A_4SjneQ7j3_0;
	wire w_dff_A_3VrIdUWG7_0;
	wire w_dff_A_TKIxaGy19_0;
	wire w_dff_A_8J7Opxhj7_0;
	wire w_dff_B_SQh2gQdA3_1;
	wire w_dff_B_BJ6Rooop7_1;
	wire w_dff_B_748Igfu64_1;
	wire w_dff_B_DcC6rqkx2_1;
	wire w_dff_B_JVUOG1LR0_1;
	wire w_dff_B_xKDCvSCA8_1;
	wire w_dff_B_6kyTUGvp2_1;
	wire w_dff_B_OAGK93mI9_1;
	wire w_dff_B_hypuAYjm0_1;
	wire w_dff_B_6pDOdZjL4_1;
	wire w_dff_B_7hEdY94K4_1;
	wire w_dff_B_Slxm1lx63_1;
	wire w_dff_B_BBvIKtNP1_0;
	wire w_dff_B_xciTNEE36_0;
	wire w_dff_B_Ro86NhZw8_0;
	wire w_dff_B_jwgBJArJ6_0;
	wire w_dff_B_jGNFm7hT8_0;
	wire w_dff_B_dd85IcJm3_0;
	wire w_dff_B_udz6a51B2_0;
	wire w_dff_B_8R9AMw6g2_0;
	wire w_dff_B_BuFks82O4_0;
	wire w_dff_B_Imz9GHSJ2_0;
	wire w_dff_B_xxDbMDP82_0;
	wire w_dff_B_D7WhIya89_0;
	wire w_dff_B_zyeN6HZ17_0;
	wire w_dff_B_uPAk3PsE8_0;
	wire w_dff_A_dXEIWgDr5_0;
	wire w_dff_A_UblRcr5H7_0;
	wire w_dff_A_GbX3sqRV6_0;
	wire w_dff_A_jNwtQAJy2_0;
	wire w_dff_A_SBVTTQf23_0;
	wire w_dff_A_txZ7Byz38_0;
	wire w_dff_A_8uVVB5dg1_0;
	wire w_dff_A_3CkFEYoY8_0;
	wire w_dff_A_EYRVDabA5_0;
	wire w_dff_A_PsEwy2V65_0;
	wire w_dff_A_3G1Q4sZu6_0;
	wire w_dff_A_fZa86WO57_0;
	wire w_dff_A_DBUrhVvv0_0;
	wire w_dff_A_amj7g5Eo1_0;
	wire w_dff_A_TB6WP7ZL0_0;
	wire w_dff_B_kP0FXXRz4_1;
	wire w_dff_B_v6jcs1Tw1_1;
	wire w_dff_B_7SdlZiU25_1;
	wire w_dff_B_IcRwO1FJ6_1;
	wire w_dff_B_gQBk2m2P4_1;
	wire w_dff_B_iVlEzbxa0_1;
	wire w_dff_B_p0rppZQ87_1;
	wire w_dff_B_2nxCeAFo6_1;
	wire w_dff_B_bzqeEy5W3_1;
	wire w_dff_B_ic9vLmhp3_1;
	wire w_dff_B_233cQcXb5_1;
	wire w_dff_B_LUDNu2k16_1;
	wire w_dff_B_3laqQ3w85_0;
	wire w_dff_B_MRvqB5mu9_0;
	wire w_dff_B_SzAMrhsn1_0;
	wire w_dff_B_tsYHOX1q3_0;
	wire w_dff_B_u7wycnjS7_0;
	wire w_dff_B_rwp3hnEd4_0;
	wire w_dff_B_GKklkikf7_0;
	wire w_dff_B_V3T70aNx7_0;
	wire w_dff_B_Ujlr2ZEg2_0;
	wire w_dff_B_fzpbSU6a7_0;
	wire w_dff_B_rK25yWXp3_0;
	wire w_dff_B_wBy5jWGb1_0;
	wire w_dff_B_VmD68pLY4_0;
	wire w_dff_B_0pIk17TD5_0;
	wire w_dff_A_hJW82m2V4_0;
	wire w_dff_A_qcHMD30S9_0;
	wire w_dff_A_N7O9EOkX8_0;
	wire w_dff_A_j6zj1VIC0_0;
	wire w_dff_A_nhDcfOLW9_0;
	wire w_dff_A_Ckdu4Zry7_0;
	wire w_dff_A_PLKzdo2s9_0;
	wire w_dff_A_25FElTfP6_0;
	wire w_dff_A_tnZHCPXS6_0;
	wire w_dff_A_9I41b1se1_0;
	wire w_dff_A_4Ete7m1f1_0;
	wire w_dff_A_528SSXMD5_0;
	wire w_dff_A_2rWGtBLo2_0;
	wire w_dff_A_5o1TCmD08_0;
	wire w_dff_A_CcABDC6X3_0;
	wire w_dff_B_hhH2xC3T0_1;
	wire w_dff_B_c0dvw7ia2_0;
	wire w_dff_B_DoWwuulz7_0;
	wire w_dff_B_8o2Hng001_0;
	wire w_dff_B_zfNmRqNX3_0;
	wire w_dff_B_boihjMx19_0;
	wire w_dff_B_c1jH6Jpe8_0;
	wire w_dff_B_nhcB0gVo4_0;
	wire w_dff_B_8taZhUz01_0;
	wire w_dff_B_PoYWSBeP3_0;
	wire w_dff_B_rpsa5okZ2_0;
	wire w_dff_B_v1dQ2yPZ9_0;
	wire w_dff_B_NEupvcRc5_0;
	wire w_dff_B_LsTfgIb25_0;
	wire w_dff_B_6ZN0m6354_0;
	wire w_dff_A_mBkQ8FAy0_1;
	wire w_dff_A_YN62kmNa5_1;
	wire w_dff_A_aNi0VYs67_1;
	wire w_dff_A_f5GXX9C38_1;
	wire w_dff_A_DD2Q51WV7_1;
	wire w_dff_A_76QmUyYJ1_1;
	wire w_dff_A_hXQ8m05g6_1;
	wire w_dff_A_zYPqyOQZ3_1;
	wire w_dff_A_iKRB8Wsv9_1;
	wire w_dff_A_MT0lSSNP4_1;
	wire w_dff_A_MfaGeG4A4_1;
	wire w_dff_A_s8bj5XiD9_1;
	wire w_dff_A_7sHtpric0_1;
	wire w_dff_A_XhwenyFf1_1;
	wire w_dff_A_6mnfjbqs5_1;
	wire w_dff_B_6Mcs3N3a4_1;
	wire w_dff_B_IquWU2O29_1;
	wire w_dff_B_TyHydjQp0_1;
	wire w_dff_B_mD54nwjh4_1;
	wire w_dff_B_z8h3506y6_1;
	wire w_dff_B_2GaigCDV5_1;
	wire w_dff_B_lQkRj6Iz3_1;
	wire w_dff_B_LudLZ19a0_1;
	wire w_dff_B_VsWPvjX49_1;
	wire w_dff_B_qbYWJHA10_1;
	wire w_dff_B_O9sw4Yu05_1;
	wire w_dff_B_sSDWAtkI3_1;
	wire w_dff_B_Le9lD93B3_1;
	wire w_dff_B_GnHCDVG52_1;
	wire w_dff_B_PUcHH9zB0_1;
	wire w_dff_B_H800PHkW1_0;
	wire w_dff_B_XO80HZbQ7_0;
	wire w_dff_B_HyClYrg89_0;
	wire w_dff_B_PkibqWmq9_0;
	wire w_dff_B_Hqj4vDCg5_0;
	wire w_dff_B_Hgqy3dFk0_0;
	wire w_dff_B_v8gxKJNi0_0;
	wire w_dff_B_1tux3dAl5_0;
	wire w_dff_B_z6c6gTAI4_0;
	wire w_dff_B_9P16P36S9_0;
	wire w_dff_B_kzZdAeqh0_0;
	wire w_dff_B_nEajhgS89_0;
	wire w_dff_B_vUCbUvtk0_0;
	wire w_dff_B_vItphulR1_0;
	wire w_dff_B_HCeY6Xsg9_0;
	wire w_dff_B_wMfhvqXj8_0;
	wire w_dff_B_V7RppE9K3_0;
	wire w_dff_B_hNunlZQT5_0;
	wire w_dff_B_FabcnBuR2_0;
	wire w_dff_B_EEEa5WqG6_0;
	wire w_dff_B_CBw6WWyj2_0;
	wire w_dff_B_vE20W2EV6_0;
	wire w_dff_B_wJ4gMpo62_0;
	wire w_dff_B_21naDq6z9_0;
	wire w_dff_B_03H9PegJ1_0;
	wire w_dff_B_utAAeGFS6_1;
	wire w_dff_B_vd9YvGa17_1;
	wire w_dff_B_ooi95S6u9_0;
	wire w_dff_B_i5PDVMKi8_0;
	wire w_dff_B_FMRsiVLd6_0;
	wire w_dff_B_6EiM8kwb2_0;
	wire w_dff_B_cyxcypYz0_0;
	wire w_dff_B_N3mjGSh68_0;
	wire w_dff_B_CTe91qRz2_0;
	wire w_dff_B_IgAnoSEi5_0;
	wire w_dff_B_w8VI9R5M8_0;
	wire w_dff_B_fdQnRn6U8_0;
	wire w_dff_B_KCOZqQJA1_0;
	wire w_dff_B_6twX056v2_0;
	wire w_dff_B_oKxb8BLI3_0;
	wire w_dff_B_bNBiZI2c2_1;
	wire w_dff_B_0kZ2z18R8_0;
	wire w_dff_A_A0xHajm72_0;
	wire w_dff_A_2Qa4mDst8_0;
	wire w_dff_A_qkEZTYbq6_2;
	wire w_dff_A_Q9G6vVgF3_2;
	wire w_dff_A_jsAhbsnF8_0;
	wire w_dff_A_AqRVZuO56_2;
	wire w_dff_B_xAj10c8M8_3;
	wire w_dff_B_VWqHtd9m4_0;
	wire w_dff_A_l0EIxeY21_0;
	wire w_dff_A_KXlByAQf7_2;
	wire w_dff_A_jQgXWgqB0_2;
	wire w_dff_A_2MC35eKk5_0;
	wire w_dff_A_bIOKmwFE6_0;
	wire w_dff_A_7hU9kEf18_1;
	wire w_dff_A_HHgnVmET5_1;
	wire w_dff_A_L8M4JS3W9_0;
	wire w_dff_A_e0hOEbT09_2;
	wire w_dff_B_XXYDJJC69_3;
	wire w_dff_A_uOwPDkx45_0;
	wire w_dff_A_ALtmhgTc6_0;
	wire w_dff_A_8RuVw5tC8_1;
	wire w_dff_A_EGYRcwBO5_1;
	wire w_dff_A_9SSMtdeU1_2;
	wire w_dff_A_gtbJ1B1o4_2;
	wire w_dff_A_fOwRUP1N3_2;
	wire w_dff_B_W1OUvgBT0_3;
	wire w_dff_A_Shzbzd048_1;
	wire w_dff_A_W6SoiKOo9_1;
	wire w_dff_A_VFOZdRBQ2_1;
	wire w_dff_A_FvrCfnJD3_1;
	wire w_dff_A_I348fSb59_2;
	wire w_dff_A_Mogc7lRq2_2;
	wire w_dff_A_y4d6FUuI4_2;
	wire w_dff_A_hDLlR9aU9_2;
	wire w_dff_B_fmX5IGTT2_3;
	wire w_dff_B_VihuQQtv3_3;
	wire w_dff_B_iqoVMd6k3_3;
	wire w_dff_B_ylKjk9M09_3;
	wire w_dff_B_ugbwOPxA9_3;
	wire w_dff_B_91GUwpgB9_3;
	wire w_dff_B_PtF5RnJI4_3;
	wire w_dff_B_ews6HzcO6_3;
	wire w_dff_B_x22F5vcs9_3;
	wire w_dff_B_OwRWhq653_3;
	wire w_dff_B_iRIJRMt13_3;
	wire w_dff_B_8eHgVTOX8_3;
	wire w_dff_B_aqMOPiYk9_3;
	wire w_dff_B_AiVg1xue0_3;
	wire w_dff_B_LKvHw9nw2_3;
	wire w_dff_B_XEK9xg8v1_3;
	wire w_dff_B_qrCXNbTi1_1;
	wire w_dff_B_kmet4QdL0_1;
	wire w_dff_B_UIP3Bl9K0_1;
	wire w_dff_B_fC369nER5_1;
	wire w_dff_B_fFhIUMYH7_1;
	wire w_dff_B_MSky3R4C5_1;
	wire w_dff_B_8etoQi9d5_1;
	wire w_dff_B_Z35LIqLt5_1;
	wire w_dff_B_CxMlmehe3_1;
	wire w_dff_B_rM6vO3xV6_1;
	wire w_dff_B_rg16n2yA1_1;
	wire w_dff_B_dn0deQQx3_0;
	wire w_dff_B_rHLRHm304_0;
	wire w_dff_B_dBUl07bo3_0;
	wire w_dff_B_nFgPMPZJ8_0;
	wire w_dff_B_e6POofZE0_0;
	wire w_dff_B_k9as2cgn9_0;
	wire w_dff_B_iJ1Sgwnx8_0;
	wire w_dff_B_MHYNxXFv3_0;
	wire w_dff_B_xh2IlJkJ3_0;
	wire w_dff_B_TpthdZRQ8_0;
	wire w_dff_B_ZItEWuXN2_0;
	wire w_dff_B_VNNNKHBf2_0;
	wire w_dff_B_YYTIRybh0_0;
	wire w_dff_B_dl0Rx4Pp3_0;
	wire w_dff_A_1fyWL2jF4_0;
	wire w_dff_A_73TrNSFc1_0;
	wire w_dff_A_hmd0lHZm7_0;
	wire w_dff_A_oxJmmROU8_0;
	wire w_dff_A_T0lDex9y5_0;
	wire w_dff_A_F0V9QpbM3_0;
	wire w_dff_A_UBbUylUN6_0;
	wire w_dff_A_PVzqeHDp0_0;
	wire w_dff_A_hGkt8E1k4_0;
	wire w_dff_A_mSLNJsGa4_0;
	wire w_dff_A_pMrlqy470_0;
	wire w_dff_A_m6Qx9DAJ2_0;
	wire w_dff_A_LhM1B9Pt1_0;
	wire w_dff_A_fd4PZKEL4_0;
	wire w_dff_A_U46uTslA6_0;
	wire w_dff_B_qRJjuky49_0;
	wire w_dff_B_P1oev6OL7_0;
	wire w_dff_A_O4s2vHtd0_1;
	wire w_dff_A_eRcrnQaJ8_1;
	wire w_dff_B_0F73FT6u8_2;
	wire w_dff_A_CtB0uMGN2_1;
	wire w_dff_A_NtqSXtuH4_1;
	wire w_dff_A_hBG93Yhh6_2;
	wire w_dff_A_7XvFw0v89_2;
	wire w_dff_B_6TFqzJ3w3_3;
	wire w_dff_B_IEPWR7JI3_3;
	wire w_dff_A_DjGGIK7h6_0;
	wire w_dff_A_FKtcFAdn1_1;
	wire w_dff_B_IwweuLLc4_3;
	wire w_dff_A_n1nyfuVj7_1;
	wire w_dff_A_OZ8KK12W0_2;
	wire w_dff_B_xgSN3V3V7_3;
	wire w_dff_A_pbPmsnQ15_0;
	wire w_dff_A_aL9ZvaMz2_0;
	wire w_dff_A_EWqnEigz3_0;
	wire w_dff_A_WrjgMOFJ0_1;
	wire w_dff_A_E73AQ5V10_1;
	wire w_dff_A_CpOdx5Gu0_1;
	wire w_dff_B_wOFWd6LP3_0;
	wire w_dff_B_GAw23NGM7_1;
	wire w_dff_B_nCvU86gK5_0;
	wire w_dff_A_REGWZ8k48_1;
	wire w_dff_A_n2Tcoh2U6_0;
	wire w_dff_B_vBdGNBbj5_3;
	wire w_dff_A_VrzoVLr50_0;
	wire w_dff_A_lnNYhLRA3_0;
	wire w_dff_B_sJq7yOVI7_3;
	wire w_dff_A_IANGZgsD2_0;
	wire w_dff_A_OK5if8aX3_0;
	wire w_dff_A_tmxZjWrt0_2;
	wire w_dff_A_XI8h2cgr0_2;
	wire w_dff_B_E2Ozntam6_2;
	wire w_dff_A_X1itAvbh4_1;
	wire w_dff_A_L4GXIG7G1_1;
	wire w_dff_A_T3WBiKFQ5_2;
	wire w_dff_A_19nn0ZKO9_2;
	wire w_dff_B_RlcOllUj0_1;
	wire w_dff_B_BttTsZuX8_1;
	wire w_dff_B_2NvLaf0d2_1;
	wire w_dff_B_E6KpvIQS1_1;
	wire w_dff_B_tgqTKjST6_1;
	wire w_dff_A_3uMTGr290_0;
	wire w_dff_A_enOvBShm0_0;
	wire w_dff_A_ENUTJ48H9_0;
	wire w_dff_A_8LcSwH8V3_0;
	wire w_dff_A_1W7IgUaM5_0;
	wire w_dff_A_58imru5c5_0;
	wire w_dff_A_TsBU1uMv0_0;
	wire w_dff_A_sPGb23ld7_0;
	wire w_dff_A_k3v7wEYI1_0;
	wire w_dff_A_6AJDCdFE1_0;
	wire w_dff_A_XLhE6Odj0_0;
	wire w_dff_A_sTQzwxcp3_1;
	wire w_dff_B_RiIbFyzW2_3;
	wire w_dff_B_GQ5WKW4Z3_2;
	wire w_dff_A_LPKtXx3w1_1;
	wire w_dff_A_375026EZ7_1;
	wire w_dff_A_4M3NhlzX8_2;
	wire w_dff_A_MM0cDStJ0_2;
	wire w_dff_B_RYP7aEv24_1;
	wire w_dff_B_iB72dv0Z8_1;
	wire w_dff_B_al3r44FB2_1;
	wire w_dff_B_A7iquh0X4_1;
	wire w_dff_B_gkBWQhNm3_1;
	wire w_dff_A_gg5hEwhF8_0;
	wire w_dff_A_WenNg6Ky8_0;
	wire w_dff_A_MwJvXmnu9_0;
	wire w_dff_A_pDQ020eG4_0;
	wire w_dff_A_Q68tyZJT3_0;
	wire w_dff_A_LC3rQaQt4_0;
	wire w_dff_A_ZmC3SGWn1_0;
	wire w_dff_A_Ljyw1Tfj2_0;
	wire w_dff_A_0ya4Ojth2_0;
	wire w_dff_A_gRXzx6lV4_0;
	wire w_dff_A_ehwNMh3i9_0;
	wire w_dff_A_gV3TYRGf2_0;
	wire w_dff_B_wGKmiluw8_1;
	wire w_dff_B_32cs7bWc2_1;
	wire w_dff_A_iMghNJmt4_1;
	wire w_dff_A_r5EtnzcC9_1;
	wire w_dff_A_hAaYs4WB6_1;
	wire w_dff_A_Teu1UDtW7_1;
	wire w_dff_A_Yd45RafL0_1;
	wire w_dff_A_CEab87fn1_1;
	wire w_dff_A_PEcKYvTo2_0;
	wire w_dff_A_09Ithtd01_0;
	wire w_dff_A_0AGzoZu19_0;
	wire w_dff_A_YDij4JRz9_0;
	wire w_dff_A_NYwfiaWO3_0;
	wire w_dff_A_XnX1efKo4_0;
	wire w_dff_A_PYpkFaEB2_0;
	wire w_dff_A_FIvoixvh8_0;
	wire w_dff_A_ULOqf1aM8_0;
	wire w_dff_A_HFst59VX1_0;
	wire w_dff_A_VSiWk4ZR0_0;
	wire w_dff_A_BIDb6lWi9_0;
	wire w_dff_B_Po8Zbi7a6_1;
	wire w_dff_B_Q3GIcbza0_1;
	wire w_dff_B_KYf5x2SV2_1;
	wire w_dff_B_vWcuUjsK6_0;
	wire w_dff_A_uWZcgsMi2_1;
	wire w_dff_A_ScB36H0X3_1;
	wire w_dff_A_4c38AGAK5_1;
	wire w_dff_A_azIz4Y8S7_1;
	wire w_dff_A_xzz8La4D7_1;
	wire w_dff_A_WWtRK1vQ1_1;
	wire w_dff_B_Ecqpcddf1_3;
	wire w_dff_B_3tMQlBob3_3;
	wire w_dff_A_tw9iMYm32_0;
	wire w_dff_A_7f6FhRxn3_0;
	wire w_dff_A_qAr5oImy2_0;
	wire w_dff_A_y39Ir1fy5_1;
	wire w_dff_A_ZNGFzyY63_1;
	wire w_dff_A_SAYeAZFS1_1;
	wire w_dff_B_jF5kPCUT9_1;
	wire w_dff_A_AizOC6QN4_0;
	wire w_dff_A_IZaReYdH1_1;
	wire w_dff_A_GEijYecu8_1;
	wire w_dff_A_5Qhka2Bg4_1;
	wire w_dff_A_E7JR0M4V6_1;
	wire w_dff_A_wSuxgyHR1_1;
	wire w_dff_A_edH96Hus4_1;
	wire w_dff_A_A1IDbqi44_1;
	wire w_dff_A_SI7If7WT8_1;
	wire w_dff_A_m2SUxvgv9_1;
	wire w_dff_A_Wp07xHDd0_1;
	wire w_dff_A_CJMSy18s4_1;
	wire w_dff_A_E0bkq6j93_1;
	wire w_dff_A_o6mUYrvZ4_1;
	wire w_dff_A_6XTcObx51_1;
	wire w_dff_A_nbxBiWfY8_1;
	wire w_dff_A_anU5sl0X7_1;
	wire w_dff_A_AlhORJZi8_1;
	wire w_dff_A_Ji7TlELM7_1;
	wire w_dff_A_zVcPylW94_1;
	wire w_dff_A_FY0A5AWO0_1;
	wire w_dff_A_oQtaNTI90_1;
	wire w_dff_A_7BQyAf1X2_1;
	wire w_dff_A_aCpNVqY13_1;
	wire w_dff_A_LqDRUReX2_1;
	wire w_dff_A_iI3HD5Bp2_1;
	wire w_dff_A_BYruvW6t9_1;
	wire w_dff_A_BsR5A8Rq5_1;
	wire w_dff_B_MxIFyWbc9_3;
	wire w_dff_B_R6cGR84L7_1;
	wire w_dff_A_VuuFiaHe4_2;
	wire w_dff_A_4n5YnmTu4_1;
	wire w_dff_A_IIDNdxzU7_1;
	wire w_dff_A_UNtvUHGa2_2;
	wire w_dff_A_1kIMQEqV3_2;
	wire w_dff_A_yKYSx1j20_1;
	wire w_dff_A_pnq9SN502_1;
	wire w_dff_A_i5PFSqNZ8_1;
	wire w_dff_A_J05vdRn43_1;
	wire w_dff_A_BA8qXEPg4_1;
	wire w_dff_A_J4ywwvin4_1;
	wire w_dff_B_DyUFSELa6_2;
	wire w_dff_B_LVp1aPXk1_2;
	wire w_dff_B_AE97KynP0_2;
	wire w_dff_B_d1Qt6Vw90_2;
	wire w_dff_A_90bTC5ic7_1;
	wire w_dff_A_UVej9Q6S7_1;
	wire w_dff_A_749vA3zO2_2;
	wire w_dff_A_mEDlAG3r4_2;
	wire w_dff_A_cIAEdAzU8_2;
	wire w_dff_A_tPK35H4x3_0;
	wire w_dff_A_UQwIdcxJ2_0;
	wire w_dff_A_xCadTaOD3_0;
	wire w_dff_A_Co9J3NuT7_0;
	wire w_dff_A_dmJ8NtAT6_0;
	wire w_dff_A_5OU4Hzhe9_0;
	wire w_dff_A_ZrJcMgV21_0;
	wire w_dff_A_XOWBeYFi1_0;
	wire w_dff_A_4vKkhNU22_0;
	wire w_dff_A_4opZYrHl7_0;
	wire w_dff_B_aY3Muk5q7_1;
	wire w_dff_B_hdLbOZDB0_1;
	wire w_dff_B_pKaR8eaA2_1;
	wire w_dff_B_Z3x4UZAt1_0;
	wire w_dff_B_qBlcKSpa6_0;
	wire w_dff_B_HZXyvK1o2_0;
	wire w_dff_A_lWle4vzx4_2;
	wire w_dff_A_ND1zml4C2_2;
	wire w_dff_A_zGKtC6DJ0_2;
	wire w_dff_A_qbrnQueL8_2;
	wire w_dff_A_DE4xhmAQ3_0;
	wire w_dff_A_wrXkq0xj6_0;
	wire w_dff_A_F0OlzLAD1_0;
	wire w_dff_A_NYHFwaqr6_0;
	wire w_dff_A_LY3FGZA26_0;
	wire w_dff_A_09DJ5dNl8_0;
	wire w_dff_A_ZsGqYRqj6_0;
	wire w_dff_A_TJWDZQVb4_0;
	wire w_dff_A_dkTleeez0_0;
	wire w_dff_A_KgoQ2qci2_2;
	wire w_dff_A_5C5HgrQm5_2;
	wire w_dff_A_g1cQAKUA6_2;
	wire w_dff_A_iVMlshMV6_2;
	wire w_dff_A_yQejMPDK3_0;
	wire w_dff_B_UXWqgLLL9_3;
	wire w_dff_B_7FRH8gBm4_1;
	wire w_dff_B_wYNYSM4x6_1;
	wire w_dff_B_fMGbrcGh6_1;
	wire w_dff_B_gK9l3Sqx9_1;
	wire w_dff_B_Jx9tTa653_1;
	wire w_dff_A_ID1k2XuY2_0;
	wire w_dff_A_d7FDJCNO2_0;
	wire w_dff_A_XvdFCzrw3_0;
	wire w_dff_A_plQxmdKp7_0;
	wire w_dff_A_vUaupqrr8_0;
	wire w_dff_A_gB9U7PJY9_0;
	wire w_dff_A_cMugvh9q4_0;
	wire w_dff_A_TDbpR4YG0_0;
	wire w_dff_A_2UAMgQJC5_0;
	wire w_dff_A_0FoaCd5f8_0;
	wire w_dff_A_c18q2Jzj9_0;
	wire w_dff_A_O0ethJcU8_0;
	wire w_dff_B_EMzFG6GW9_1;
	wire w_dff_B_2VYMP6Op9_1;
	wire w_dff_B_skuoW42i7_2;
	wire w_dff_A_6D5aWB4x7_0;
	wire w_dff_A_O3vkfvPD5_0;
	wire w_dff_A_xNFSjN763_0;
	wire w_dff_A_euZgJ5on4_0;
	wire w_dff_A_ZlbdMtWu2_0;
	wire w_dff_A_QbEWsmZH7_0;
	wire w_dff_A_TdzEgtCD0_0;
	wire w_dff_A_y8dDQ0a08_0;
	wire w_dff_A_5zEdiTvk8_0;
	wire w_dff_A_RJ5QVG8f1_0;
	wire w_dff_A_wKRISSfC8_0;
	wire w_dff_A_ErJwq7to0_0;
	wire w_dff_A_e3lVX8gh2_2;
	wire w_dff_A_gIN7R3uf1_2;
	wire w_dff_A_mERP0ZkL1_2;
	wire w_dff_A_c70Dbpyw4_2;
	wire w_dff_A_7ZWMuhfi8_2;
	wire w_dff_A_TyI5Y8M08_2;
	wire w_dff_B_WcRU6Qft7_2;
	wire w_dff_B_7quUQe1I0_2;
	wire w_dff_B_pJ0ykcTy3_2;
	wire w_dff_A_aO2f3qcc7_0;
	wire w_dff_A_XNfeC4qt2_0;
	wire w_dff_A_VthqGAlY9_0;
	wire w_dff_A_tqhHZpRV0_0;
	wire w_dff_B_7iPPSUpd2_1;
	wire w_dff_A_5VXt3w777_0;
	wire w_dff_A_7Jpnt4JB2_0;
	wire w_dff_A_PqzGkrR80_0;
	wire w_dff_A_HEbrDUYk4_0;
	wire w_dff_A_xGppPr3k5_1;
	wire w_dff_A_3T0Mu2XP9_2;
	wire w_dff_A_0asksFzo1_1;
	wire w_dff_A_WhLdinJl8_1;
	wire w_dff_A_L7rbIXSV3_1;
	wire w_dff_B_f02cB3R30_1;
	wire w_dff_B_JeWlBlYS1_1;
	wire w_dff_B_hXeRC8QT0_1;
	wire w_dff_A_x1lg016P1_0;
	wire w_dff_A_j272sTqQ3_0;
	wire w_dff_A_gLpiljix5_0;
	wire w_dff_A_9Vav6S578_0;
	wire w_dff_A_vhbPjJiy3_0;
	wire w_dff_A_H88aFHDB1_0;
	wire w_dff_A_DHK4VAkF2_0;
	wire w_dff_A_ft3kdH7l3_0;
	wire w_dff_A_OI8DS2hM9_0;
	wire w_dff_A_oNSKDJch6_0;
	wire w_dff_A_EBXwMR433_0;
	wire w_dff_A_ZhXSyGLz0_0;
	wire w_dff_B_jhzHQqfo5_1;
	wire w_dff_A_hGaPrqic9_0;
	wire w_dff_A_BUEBrPCd2_0;
	wire w_dff_A_hKYDeIqG7_0;
	wire w_dff_A_LK2anFOc8_0;
	wire w_dff_A_GoHPD5xI5_0;
	wire w_dff_A_MP3BtIz50_0;
	wire w_dff_A_2EprVAK18_0;
	wire w_dff_A_e5FFRQJK9_0;
	wire w_dff_A_71AJuITo6_0;
	wire w_dff_A_ABJqDcHw9_0;
	wire w_dff_A_WCLJcx8e0_0;
	wire w_dff_A_wEwstavb2_0;
	wire w_dff_A_guNlDc5m9_1;
	wire w_dff_A_oICwdoW57_1;
	wire w_dff_B_8hXZiefv1_2;
	wire w_dff_A_rfpRIPBm1_0;
	wire w_dff_A_w8A4JYm67_0;
	wire w_dff_A_ADPXycaA9_0;
	wire w_dff_A_FdJbRLZR0_0;
	wire w_dff_A_JAW0FIg22_0;
	wire w_dff_A_LW17otL16_0;
	wire w_dff_A_eFpoyJQ54_0;
	wire w_dff_A_0ztDfp9y9_0;
	wire w_dff_A_7MthCdBr7_0;
	wire w_dff_A_TzaH7j9q2_0;
	wire w_dff_A_yMA7LU7d8_0;
	wire w_dff_A_9wStfIcu0_0;
	wire w_dff_A_Mjp2c5pP9_0;
	wire w_dff_B_FXE00Kze7_1;
	wire w_dff_A_SZ1Nm9Cs6_0;
	wire w_dff_A_b8kOHhoQ6_0;
	wire w_dff_A_3BvIEyqz4_0;
	wire w_dff_A_fl5DajHF6_0;
	wire w_dff_A_f9VF20vk0_0;
	wire w_dff_A_N8KbK16P5_0;
	wire w_dff_A_ZrfOKXBg8_0;
	wire w_dff_A_XTL9CeRp9_0;
	wire w_dff_A_TeErh5ES0_0;
	wire w_dff_A_w9oDyhL51_0;
	wire w_dff_A_DYKoNI6Y5_0;
	wire w_dff_A_w6XTsMsq8_0;
	wire w_dff_A_97FbSwfK4_0;
	wire w_dff_A_GoqsyYIm8_0;
	wire w_dff_A_T4Eaq92Z3_0;
	wire w_dff_A_zElM6zFu1_0;
	wire w_dff_A_DRxUm7kI2_0;
	wire w_dff_A_3yPtjfDy8_0;
	wire w_dff_A_e8loeeor5_0;
	wire w_dff_A_05FENPcz7_0;
	wire w_dff_A_ec6pBWD25_0;
	wire w_dff_A_9IfFmerl9_0;
	wire w_dff_A_W4DPFxFO0_0;
	wire w_dff_A_PB4RuL8e9_0;
	wire w_dff_A_WtxmHIdG9_1;
	wire w_dff_A_ADaMUmKc6_1;
	wire w_dff_A_Xk15ibSQ5_1;
	wire w_dff_A_kOA2vvfP0_1;
	wire w_dff_A_GoWajBuW7_1;
	wire w_dff_A_UdgX3NmM7_1;
	wire w_dff_A_huAXcbKv0_1;
	wire w_dff_A_Jqqv8qbg7_1;
	wire w_dff_A_vATM0Lp49_1;
	wire w_dff_A_RV81MCiQ5_1;
	wire w_dff_A_f7OK7zOE3_1;
	wire w_dff_A_YsiZRDlq9_1;
	wire w_dff_A_lJjo43g72_1;
	wire w_dff_A_d0Eel5RY2_1;
	wire w_dff_A_EyY3UJfQ7_1;
	wire w_dff_A_EeE4pWsK2_2;
	wire w_dff_A_tyLlt4Ug9_1;
	wire w_dff_A_etytuETZ9_1;
	wire w_dff_A_11apbKMy5_1;
	wire w_dff_A_GI9ubTPs6_1;
	wire w_dff_A_1FZCsts23_1;
	wire w_dff_A_S7LbMjC51_1;
	wire w_dff_A_ObpxlGIK4_1;
	wire w_dff_A_0NJh9BDP9_1;
	wire w_dff_A_xzrtJekW4_1;
	wire w_dff_A_wNZ0DuLF0_1;
	wire w_dff_A_95ahYNiN7_1;
	wire w_dff_A_6vbxWAv54_1;
	wire w_dff_A_O4L5RZ7b7_1;
	wire w_dff_A_9G3HKwwo0_1;
	wire w_dff_A_qFoE6ANk9_1;
	wire w_dff_A_fxY1ZImU6_1;
	wire w_dff_A_6FnxbwUU6_1;
	wire w_dff_A_wCCgcxh21_1;
	wire w_dff_A_hjgtmlav3_1;
	wire w_dff_A_ntsyURLv6_1;
	wire w_dff_A_sq6nP6G67_1;
	wire w_dff_A_dSjSA72F1_1;
	wire w_dff_A_hwV4ctbQ9_1;
	wire w_dff_A_RT5C6dx18_1;
	wire w_dff_A_5QxyESWo5_1;
	wire w_dff_A_3twR1F1A9_0;
	wire w_dff_A_lly5St5y0_0;
	wire w_dff_A_E0hdVmTV6_0;
	wire w_dff_A_izuiToZY1_0;
	wire w_dff_A_ASA7AT1X9_0;
	wire w_dff_A_GezeG4B26_1;
	wire w_dff_A_94DAfcxq4_1;
	wire w_dff_A_2Qz32MAY7_1;
	wire w_dff_A_3vajMS4s9_1;
	wire w_dff_A_xnFTH5ZX1_1;
	wire w_dff_A_9v5QviIV3_2;
	wire w_dff_A_tUC0hJ4s2_2;
	wire w_dff_A_uj7b49bG5_2;
	wire w_dff_A_71sARR4R6_2;
	wire w_dff_A_dFpJWWmH4_2;
	wire w_dff_A_eXeabmUB1_2;
	wire w_dff_A_WylMPeS41_2;
	wire w_dff_A_C8ITO4682_1;
	wire w_dff_A_omvqrot23_0;
	wire w_dff_A_z1FKsQwb4_0;
	wire w_dff_A_LVNl98VB2_0;
	wire w_dff_A_YdIrpSVj6_0;
	wire w_dff_A_LJ8Gi4uF8_0;
	wire w_dff_A_DZEGczG83_0;
	wire w_dff_A_KMClJIRV1_0;
	wire w_dff_A_M1oAQNKf2_0;
	wire w_dff_A_cNNtsd1I4_0;
	wire w_dff_A_qtYt3qJj9_0;
	wire w_dff_A_QEH7dcRk1_0;
	wire w_dff_A_wSqvZeYI9_0;
	wire w_dff_A_UaBnAubx0_0;
	wire w_dff_A_c6EKCiTg3_0;
	wire w_dff_A_dAvRHgeN0_0;
	wire w_dff_A_hkaXSMhD4_0;
	wire w_dff_A_ceF5DLAr8_0;
	wire w_dff_A_v9tLWDIF1_0;
	wire w_dff_A_xgo6MV9X2_0;
	wire w_dff_A_CBh5iyhF0_0;
	wire w_dff_A_VLo057qZ4_0;
	wire w_dff_A_TyYdHk1b8_0;
	wire w_dff_A_OnKm0gGs9_0;
	wire w_dff_A_kfRW8fpl9_0;
	wire w_dff_A_1DgrQCxR4_1;
	wire w_dff_A_QPs4KyXP2_1;
	wire w_dff_A_ItqCFU3O9_1;
	wire w_dff_A_uLPdK8m11_1;
	wire w_dff_A_sj9vVAaV6_1;
	wire w_dff_A_c9chWVhq5_1;
	wire w_dff_A_eWvczxoQ7_1;
	wire w_dff_A_NzHc1JiS4_1;
	wire w_dff_A_5CQyyH1w0_1;
	wire w_dff_A_t9EyqNw49_1;
	wire w_dff_A_HKSalTAP3_1;
	wire w_dff_A_CpSt5fEB7_1;
	wire w_dff_A_17b44fcI5_1;
	wire w_dff_A_8BXKGvxZ3_1;
	wire w_dff_A_NfEoZtfz9_1;
	wire w_dff_A_aJrrWy2t9_2;
	wire w_dff_A_aypXjXkt3_2;
	wire w_dff_A_PNIcb18Q8_2;
	wire w_dff_A_OHQTwM1G8_2;
	wire w_dff_A_KHcooSNk5_2;
	wire w_dff_A_4ckL2wm82_2;
	wire w_dff_A_sgmh0wWz7_2;
	wire w_dff_A_NwLwOxON9_2;
	wire w_dff_A_1IFijKqr5_2;
	wire w_dff_A_Dr0R36Qq2_2;
	wire w_dff_A_FAXEgT0e3_2;
	wire w_dff_A_3VXP8UtH9_2;
	wire w_dff_A_PqbbI6gb8_2;
	wire w_dff_A_BnXwzpHc0_2;
	wire w_dff_A_MewQL7980_2;
	wire w_dff_A_jtdazSx98_1;
	wire w_dff_A_32dO2mgZ8_0;
	wire w_dff_A_y6vKYzLK4_0;
	wire w_dff_A_nSLHMqQ46_0;
	wire w_dff_A_q1UogLyh4_0;
	wire w_dff_A_z87XFPGG2_0;
	wire w_dff_A_I9lUJXPJ2_0;
	wire w_dff_A_tkXz10Lf5_0;
	wire w_dff_A_eVRXWvqv9_0;
	wire w_dff_A_YqIhGlMJ0_0;
	wire w_dff_A_7FVeCVei6_0;
	wire w_dff_A_fjjRkyM94_0;
	wire w_dff_A_xokxmThT8_2;
	wire w_dff_B_nhW2gutN0_3;
	wire w_dff_A_zw6Yoo2x9_1;
	wire w_dff_A_QYrbG5kf3_0;
	wire w_dff_A_g1ggyjHE6_0;
	wire w_dff_A_qlAwMW466_0;
	wire w_dff_A_uoLsdpJJ8_0;
	wire w_dff_A_TLRcHvBK0_0;
	wire w_dff_A_G3SHcqRu0_0;
	wire w_dff_A_F5vqeNN54_0;
	wire w_dff_A_4QrWqADd8_0;
	wire w_dff_A_HqrT7uBB3_0;
	wire w_dff_A_uqjWhDGs4_0;
	wire w_dff_A_rEvntC530_0;
	wire w_dff_A_kWji1Z9g6_0;
	wire w_dff_A_ixzV3uN88_0;
	wire w_dff_A_7QMqde7C1_0;
	wire w_dff_A_fTN0M8Nl9_0;
	wire w_dff_A_Xvs9Klv14_0;
	wire w_dff_A_kYAyEiQQ5_0;
	wire w_dff_A_E4mlpWHo2_0;
	wire w_dff_A_hlClqw9d9_0;
	wire w_dff_A_NKLr0QsT4_0;
	wire w_dff_A_9lrOEVyf1_0;
	wire w_dff_A_1jlZLf9J6_0;
	wire w_dff_A_UbfACKGM5_0;
	wire w_dff_A_AQxkgjvZ4_0;
	wire w_dff_A_vFPHv5Kn6_0;
	wire w_dff_A_5uLjVev71_0;
	wire w_dff_A_mhvx7r855_0;
	wire w_dff_A_RNYdsNw95_0;
	wire w_dff_A_LqK2UbH56_0;
	wire w_dff_A_Z7vQxSIJ0_0;
	wire w_dff_A_ge88EaDK2_0;
	wire w_dff_A_MGD9JNrL1_0;
	wire w_dff_A_tNRargS47_0;
	wire w_dff_A_YZHVwf6Q8_0;
	wire w_dff_A_wW6jRfOH3_0;
	wire w_dff_A_uGUkLdGk8_0;
	wire w_dff_B_rrIwJGG22_1;
	wire w_dff_A_QFbJyn4L1_0;
	wire w_dff_A_XUxXPWpj3_0;
	wire w_dff_A_3GdzA8GT8_0;
	wire w_dff_A_qyhQuvCh2_0;
	wire w_dff_A_kP1S94qw3_0;
	wire w_dff_A_np2tc0dK7_0;
	wire w_dff_A_bcKuHTcd4_0;
	wire w_dff_A_ch50iC326_0;
	wire w_dff_A_7pcJFWUh4_0;
	wire w_dff_A_C0Oae3SM7_0;
	wire w_dff_A_nil8ntDj1_0;
	wire w_dff_A_Ooj9orFX9_0;
	wire w_dff_A_iwuOnkwX7_1;
	wire w_dff_A_V2GnYsRI4_1;
	wire w_dff_A_4NJCaWES2_1;
	wire w_dff_A_CZgREzlJ7_1;
	wire w_dff_A_qtqbA7TE2_1;
	wire w_dff_A_xjC3xC1f3_1;
	wire w_dff_A_gjJLpUjO2_1;
	wire w_dff_A_0FBt5On70_1;
	wire w_dff_A_RiPSRki43_1;
	wire w_dff_A_iOJCDytV9_1;
	wire w_dff_A_PtVCZn1s7_1;
	wire w_dff_A_KvChh7Xe5_1;
	wire w_dff_A_tAIPdC814_2;
	wire w_dff_A_uPQtcYLi3_0;
	wire w_dff_A_8dGNuAjS6_1;
	wire w_dff_A_SKEkCR5y1_1;
	wire w_dff_A_bAvRgBrY7_1;
	wire w_dff_A_4a5ZjSeF2_1;
	wire w_dff_A_ML9fB5ek4_1;
	wire w_dff_A_pasSz2kO4_1;
	wire w_dff_A_HJTlownT6_1;
	wire w_dff_A_ZbpgyP838_1;
	wire w_dff_A_f9Epro6U8_1;
	wire w_dff_A_AaxeuSG62_1;
	wire w_dff_A_j6eTlFGV7_1;
	wire w_dff_A_TOF1ISug0_1;
	wire w_dff_A_wOV34ZYg8_1;
	wire w_dff_A_mQkGIWB23_0;
	wire w_dff_A_zXIWKv336_0;
	wire w_dff_A_HiXB6ErV1_0;
	wire w_dff_A_OiKv6x1P3_0;
	wire w_dff_A_MatWtpgi3_0;
	wire w_dff_A_oQ8MpKlk1_0;
	wire w_dff_A_VxZaGK1w3_0;
	wire w_dff_A_9EuIiA1r1_0;
	wire w_dff_A_1MXo40gh8_0;
	wire w_dff_A_UsCn5THH1_0;
	wire w_dff_A_hApYUv2t3_0;
	wire w_dff_A_3crr4E687_0;
	wire w_dff_A_TKgBSNOc3_0;
	wire w_dff_A_GtPlbU3g8_0;
	wire w_dff_A_6wgcFCk43_0;
	wire w_dff_A_p1WLYOiw3_0;
	wire w_dff_A_rEzsa2tP4_0;
	wire w_dff_A_A7GFZBeo0_0;
	wire w_dff_A_hvHGuKJ83_0;
	wire w_dff_A_9nhakWyN2_0;
	wire w_dff_A_WZ3AznBH3_0;
	wire w_dff_A_VkgiVfXZ7_0;
	wire w_dff_A_kaFOH6IU9_0;
	wire w_dff_A_gwoGQgPo3_2;
	wire w_dff_A_0jUAIR0N0_2;
	wire w_dff_B_TYwom6MH1_3;
	wire w_dff_A_Hk3nXfqo8_0;
	wire w_dff_A_BmZUYzin4_0;
	wire w_dff_A_b5eJjfJ28_0;
	wire w_dff_A_CrhC5AA46_0;
	wire w_dff_A_4qiJJOE21_0;
	wire w_dff_A_sSivf5sT5_0;
	wire w_dff_A_Ji5K9ZSn0_0;
	wire w_dff_A_1bPf2LbR7_0;
	wire w_dff_A_j27VBrhb1_0;
	wire w_dff_A_Pr4o3CpU3_0;
	wire w_dff_A_AwtVxnWA7_0;
	wire w_dff_A_etucNoNa4_0;
	wire w_dff_A_tgsGGwUG3_2;
	wire w_dff_A_Jo05WalF4_0;
	wire w_dff_A_lQQ7OrNU9_0;
	wire w_dff_A_Oo8xOv4Z2_0;
	wire w_dff_A_1yTGniJ24_0;
	wire w_dff_A_9CGrs0b87_0;
	wire w_dff_A_irGhth8U4_0;
	wire w_dff_A_1jvHz01S6_2;
	wire w_dff_A_h6B22lMB2_0;
	wire w_dff_A_FLxDXH7i7_0;
	wire w_dff_A_fcLWlC2l7_0;
	wire w_dff_A_3MEcD3C63_0;
	wire w_dff_A_PpPLHoD77_0;
	wire w_dff_A_NWx4ToN48_0;
	wire w_dff_A_B8eR28a40_2;
	wire w_dff_A_yM9yP70s3_0;
	wire w_dff_A_AOZGbwPt8_0;
	wire w_dff_A_3aZ33zEw3_0;
	wire w_dff_A_STmyObGg3_0;
	wire w_dff_A_5zyebfVW4_0;
	wire w_dff_A_y16Uu0qQ7_0;
	wire w_dff_A_0f7i80Nd1_2;
	wire w_dff_A_R4yd7DBk4_0;
	wire w_dff_A_FcBOieOs8_0;
	wire w_dff_A_pLYsoq2Q2_0;
	wire w_dff_A_scRGQsfY4_0;
	wire w_dff_A_SOBVLc7F8_0;
	wire w_dff_A_ZfoTHkX01_0;
	wire w_dff_A_3yefOgGp2_2;
	wire w_dff_A_QjzFVJyZ8_0;
	wire w_dff_A_9cQjYvRQ1_0;
	wire w_dff_A_U4KfyalL5_0;
	wire w_dff_A_AY5bFrSp1_0;
	wire w_dff_A_ASjJGAdI0_0;
	wire w_dff_A_ijmCbDwn1_0;
	wire w_dff_A_ehYWmLY91_2;
	wire w_dff_A_IaTZkgip1_0;
	wire w_dff_A_QLAX8zKf4_0;
	wire w_dff_A_CkySIeNS0_0;
	wire w_dff_A_ukcVafbV1_0;
	wire w_dff_A_u7j7UB2c4_0;
	wire w_dff_A_AYMvHAtF2_0;
	wire w_dff_A_CxV5R3S41_2;
	wire w_dff_A_lByYvY8H8_0;
	wire w_dff_A_D67fBNeB0_0;
	wire w_dff_A_BfppoD9q8_0;
	wire w_dff_A_vt6MVxkA5_0;
	wire w_dff_A_WlEz4kmI8_0;
	wire w_dff_A_pHmFZTGV1_0;
	wire w_dff_A_iA9pP22X1_2;
	wire w_dff_A_IExpIc7W2_0;
	wire w_dff_A_sFpjpHVR7_0;
	wire w_dff_A_Ly8Z3pCD4_0;
	wire w_dff_A_hi7LkfJQ5_0;
	wire w_dff_A_68iq09Iz0_0;
	wire w_dff_A_h4SaEFY61_0;
	wire w_dff_A_OvTispEG5_2;
	wire w_dff_A_x7HgaYxP9_0;
	wire w_dff_A_d0NGJUAT7_0;
	wire w_dff_A_TrxtfwNt8_0;
	wire w_dff_A_Tu2aKiaE8_0;
	wire w_dff_A_8joY4mYZ5_0;
	wire w_dff_A_JJWlIZNC0_0;
	wire w_dff_A_Fko9CuZr6_2;
	wire w_dff_A_2jZUzQMO3_0;
	wire w_dff_A_fFYUbEWo4_0;
	wire w_dff_A_CAVjaFLi4_0;
	wire w_dff_A_Q1qrKJZf1_0;
	wire w_dff_A_xxeOSZzt9_0;
	wire w_dff_A_W8bPgPiJ6_0;
	wire w_dff_A_VxBgzGut5_2;
	wire w_dff_A_UI9HFpeL2_0;
	wire w_dff_A_qJrzVuab9_0;
	wire w_dff_A_4j4wXiaz0_0;
	wire w_dff_A_Aaedy9gb5_0;
	wire w_dff_A_lHlNJP5b7_0;
	wire w_dff_A_edZ4euLr7_0;
	wire w_dff_A_PCaNejM41_2;
	wire w_dff_A_muRMUgys2_0;
	wire w_dff_A_pVO7JxRf3_0;
	wire w_dff_A_cpS9pvUm5_0;
	wire w_dff_A_IhFQEkMO9_0;
	wire w_dff_A_xqSZaXoR3_0;
	wire w_dff_A_mCHTSb2L3_0;
	wire w_dff_A_XeL5ESXH3_2;
	wire w_dff_A_fy9LOIPT8_0;
	wire w_dff_A_xBgBFEHM7_0;
	wire w_dff_A_5gkAEx7I0_0;
	wire w_dff_A_TMpfrc1Q8_0;
	wire w_dff_A_Li6WKKvL4_0;
	wire w_dff_A_o6BgCzU64_0;
	wire w_dff_A_wxTTumbh8_2;
	wire w_dff_A_ilTLLlxC8_0;
	wire w_dff_A_Bz7H5Wjt7_0;
	wire w_dff_A_pI5WLpcv6_0;
	wire w_dff_A_1NG3OYxR8_0;
	wire w_dff_A_jp2Wqpe77_0;
	wire w_dff_A_sZZkANDc0_0;
	wire w_dff_A_5ZGcPxwR6_2;
	wire w_dff_A_BQvTciW99_0;
	wire w_dff_A_0hRpRr789_0;
	wire w_dff_A_DHl6Y7IQ9_0;
	wire w_dff_A_vT75EyGY5_0;
	wire w_dff_A_hm112p493_0;
	wire w_dff_A_teud1nbE4_0;
	wire w_dff_A_5MAg6puK2_2;
	wire w_dff_A_M4OfibrF1_0;
	wire w_dff_A_EzXgRwKQ9_0;
	wire w_dff_A_axJWYsxJ5_0;
	wire w_dff_A_7f5mwdfI9_0;
	wire w_dff_A_8OmdQrkT4_0;
	wire w_dff_A_Y2dIFbtx4_0;
	wire w_dff_A_76IhHjB45_2;
	wire w_dff_A_STzXy76t1_2;
	wire w_dff_A_BblxUM767_2;
	wire w_dff_A_PknvDO025_0;
	jnot g000(.din(w_G146_0[2]),.dout(n58),.clk(gclk));
	jxor g001(.dina(w_G140_0[2]),.dinb(w_G125_0[2]),.dout(n59),.clk(gclk));
	jxor g002(.dina(w_n59_0[1]),.dinb(n58),.dout(n60),.clk(gclk));
	jdff g003(.din(w_G953_1[2]),.dout(n61),.clk(gclk));
	jand g004(.dina(w_n61_3[2]),.dinb(w_G234_0[2]),.dout(n62),.clk(gclk));
	jand g005(.dina(w_n62_0[1]),.dinb(w_G221_0[1]),.dout(n63),.clk(gclk));
	jxor g006(.dina(n63),.dinb(w_G137_0[2]),.dout(n64),.clk(gclk));
	jxor g007(.dina(w_G128_1[1]),.dinb(w_G119_0[2]),.dout(n65),.clk(gclk));
	jor g008(.dina(w_dff_B_HZXyvK1o2_0),.dinb(n64),.dout(n66),.clk(gclk));
	jxor g009(.dina(n66),.dinb(w_G110_1[1]),.dout(n67),.clk(gclk));
	jxor g010(.dina(w_n67_0[1]),.dinb(w_n60_0[2]),.dout(n68),.clk(gclk));
	jor g011(.dina(w_n68_0[1]),.dinb(w_G902_3[2]),.dout(n69),.clk(gclk));
	jnot g012(.din(w_G902_3[1]),.dout(n70),.clk(gclk));
	jand g013(.dina(w_n70_3[1]),.dinb(w_G234_0[1]),.dout(n71),.clk(gclk));
	jnot g014(.din(w_n71_0[1]),.dout(n72),.clk(gclk));
	jand g015(.dina(n72),.dinb(w_G217_0[2]),.dout(n73),.clk(gclk));
	jxor g016(.dina(w_n73_0[1]),.dinb(n69),.dout(n74),.clk(gclk));
	jnot g017(.din(w_G134_0[2]),.dout(n75),.clk(gclk));
	jxor g018(.dina(w_G137_0[1]),.dinb(n75),.dout(n76),.clk(gclk));
	jnot g019(.din(w_G131_0[1]),.dout(n77),.clk(gclk));
	jxor g020(.dina(w_G146_0[1]),.dinb(w_G143_1[1]),.dout(n78),.clk(gclk));
	jxor g021(.dina(n78),.dinb(w_G128_1[0]),.dout(n79),.clk(gclk));
	jxor g022(.dina(w_n79_0[1]),.dinb(w_n77_0[1]),.dout(n80),.clk(gclk));
	jxor g023(.dina(n80),.dinb(w_dff_B_rrIwJGG22_1),.dout(n81),.clk(gclk));
	jnot g024(.din(w_G113_0[1]),.dout(n82),.clk(gclk));
	jxor g025(.dina(w_G119_0[1]),.dinb(w_G116_0[2]),.dout(n83),.clk(gclk));
	jxor g026(.dina(n83),.dinb(w_n82_0[1]),.dout(n84),.clk(gclk));
	jnot g027(.din(w_G210_0[2]),.dout(n85),.clk(gclk));
	jor g028(.dina(w_G953_1[1]),.dinb(w_G237_0[2]),.dout(n86),.clk(gclk));
	jor g029(.dina(w_n86_0[1]),.dinb(n85),.dout(n87),.clk(gclk));
	jxor g030(.dina(n87),.dinb(w_G101_0[2]),.dout(n88),.clk(gclk));
	jxor g031(.dina(n88),.dinb(w_n84_0[1]),.dout(n89),.clk(gclk));
	jxor g032(.dina(n89),.dinb(w_n81_0[2]),.dout(n90),.clk(gclk));
	jand g033(.dina(w_n90_0[2]),.dinb(w_n70_3[0]),.dout(n91),.clk(gclk));
	jxor g034(.dina(n91),.dinb(w_G472_0[1]),.dout(n92),.clk(gclk));
	jand g035(.dina(w_n92_1[2]),.dinb(w_n74_1[1]),.dout(n93),.clk(gclk));
	jor g036(.dina(w_G902_3[0]),.dinb(w_G237_0[1]),.dout(n94),.clk(gclk));
	jand g037(.dina(w_n94_0[1]),.dinb(w_G214_0[1]),.dout(n95),.clk(gclk));
	jnot g038(.din(w_n95_0[2]),.dout(n96),.clk(gclk));
	jand g039(.dina(w_n94_0[0]),.dinb(w_G210_0[1]),.dout(n97),.clk(gclk));
	jnot g040(.din(w_G110_1[0]),.dout(n98),.clk(gclk));
	jxor g041(.dina(w_G122_1[1]),.dinb(n98),.dout(n99),.clk(gclk));
	jxor g042(.dina(w_G107_0[2]),.dinb(w_G104_0[2]),.dout(n100),.clk(gclk));
	jxor g043(.dina(n100),.dinb(w_G101_0[1]),.dout(n101),.clk(gclk));
	jxor g044(.dina(w_n101_0[1]),.dinb(w_n84_0[0]),.dout(n102),.clk(gclk));
	jxor g045(.dina(n102),.dinb(w_dff_B_FXE00Kze7_1),.dout(n103),.clk(gclk));
	jand g046(.dina(w_n61_3[1]),.dinb(w_G224_0[1]),.dout(n104),.clk(gclk));
	jxor g047(.dina(w_n79_0[0]),.dinb(w_G125_0[1]),.dout(n105),.clk(gclk));
	jxor g048(.dina(n105),.dinb(w_dff_B_jhzHQqfo5_1),.dout(n106),.clk(gclk));
	jxor g049(.dina(n106),.dinb(w_n103_0[1]),.dout(n107),.clk(gclk));
	jand g050(.dina(w_n107_0[2]),.dinb(w_n70_2[2]),.dout(n108),.clk(gclk));
	jxor g051(.dina(w_n108_0[1]),.dinb(w_n97_0[1]),.dout(n109),.clk(gclk));
	jand g052(.dina(w_n109_0[1]),.dinb(w_n96_0[2]),.dout(n110),.clk(gclk));
	jnot g053(.din(w_G221_0[0]),.dout(n111),.clk(gclk));
	jor g054(.dina(w_n71_0[0]),.dinb(w_dff_B_7iPPSUpd2_1),.dout(n112),.clk(gclk));
	jxor g055(.dina(w_G140_0[1]),.dinb(w_G110_0[2]),.dout(n113),.clk(gclk));
	jand g056(.dina(w_n61_3[0]),.dinb(w_G227_0[1]),.dout(n114),.clk(gclk));
	jxor g057(.dina(n114),.dinb(w_n101_0[0]),.dout(n115),.clk(gclk));
	jxor g058(.dina(n115),.dinb(w_dff_B_2VYMP6Op9_1),.dout(n116),.clk(gclk));
	jxor g059(.dina(n116),.dinb(w_n81_0[1]),.dout(n117),.clk(gclk));
	jand g060(.dina(w_n117_0[2]),.dinb(w_n70_2[1]),.dout(n118),.clk(gclk));
	jxor g061(.dina(w_n118_0[1]),.dinb(w_G469_0[2]),.dout(n119),.clk(gclk));
	jand g062(.dina(w_n119_0[1]),.dinb(w_n112_1[1]),.dout(n120),.clk(gclk));
	jand g063(.dina(w_n120_0[1]),.dinb(w_n110_0[2]),.dout(n121),.clk(gclk));
	jand g064(.dina(w_n121_1[1]),.dinb(w_n93_0[2]),.dout(n122),.clk(gclk));
	jnot g065(.din(w_G478_0[2]),.dout(n123),.clk(gclk));
	jxor g066(.dina(w_G143_1[0]),.dinb(w_G128_0[2]),.dout(n124),.clk(gclk));
	jand g067(.dina(w_n62_0[0]),.dinb(w_G217_0[1]),.dout(n125),.clk(gclk));
	jxor g068(.dina(w_G122_1[0]),.dinb(w_G116_0[1]),.dout(n126),.clk(gclk));
	jxor g069(.dina(w_G134_0[1]),.dinb(w_G107_0[1]),.dout(n127),.clk(gclk));
	jxor g070(.dina(n127),.dinb(n126),.dout(n128),.clk(gclk));
	jxor g071(.dina(w_dff_B_vWcuUjsK6_0),.dinb(n125),.dout(n129),.clk(gclk));
	jxor g072(.dina(n129),.dinb(w_dff_B_KYf5x2SV2_1),.dout(n130),.clk(gclk));
	jand g073(.dina(w_n130_0[2]),.dinb(w_n70_2[0]),.dout(n131),.clk(gclk));
	jxor g074(.dina(w_n131_0[1]),.dinb(w_dff_B_tgqTKjST6_1),.dout(n132),.clk(gclk));
	jnot g075(.din(w_G475_0[2]),.dout(n133),.clk(gclk));
	jxor g076(.dina(w_G143_0[2]),.dinb(w_n77_0[0]),.dout(n134),.clk(gclk));
	jxor g077(.dina(w_G122_0[2]),.dinb(w_n82_0[0]),.dout(n135),.clk(gclk));
	jxor g078(.dina(n135),.dinb(w_G104_0[1]),.dout(n136),.clk(gclk));
	jnot g079(.din(w_G214_0[0]),.dout(n137),.clk(gclk));
	jor g080(.dina(w_n86_0[0]),.dinb(n137),.dout(n138),.clk(gclk));
	jxor g081(.dina(n138),.dinb(w_n60_0[1]),.dout(n139),.clk(gclk));
	jxor g082(.dina(n139),.dinb(n136),.dout(n140),.clk(gclk));
	jxor g083(.dina(n140),.dinb(w_dff_B_32cs7bWc2_1),.dout(n141),.clk(gclk));
	jand g084(.dina(w_n141_0[2]),.dinb(w_n70_1[2]),.dout(n142),.clk(gclk));
	jxor g085(.dina(w_n142_0[1]),.dinb(w_dff_B_gkBWQhNm3_1),.dout(n143),.clk(gclk));
	jand g086(.dina(w_n143_1[1]),.dinb(w_n132_0[2]),.dout(n144),.clk(gclk));
	jor g087(.dina(w_n61_2[2]),.dinb(w_dff_B_R6cGR84L7_1),.dout(n145),.clk(gclk));
	jand g088(.dina(w_G237_0[0]),.dinb(w_G234_0[0]),.dout(n146),.clk(gclk));
	jor g089(.dina(w_n146_0[1]),.dinb(w_n70_1[1]),.dout(n147),.clk(gclk));
	jor g090(.dina(w_n147_0[1]),.dinb(w_n145_0[1]),.dout(n148),.clk(gclk));
	jnot g091(.din(w_n146_0[0]),.dout(n149),.clk(gclk));
	jand g092(.dina(w_n61_2[1]),.dinb(w_G952_0[2]),.dout(n150),.clk(gclk));
	jand g093(.dina(n150),.dinb(n149),.dout(n151),.clk(gclk));
	jnot g094(.din(w_n151_0[2]),.dout(n152),.clk(gclk));
	jand g095(.dina(w_n152_0[1]),.dinb(w_dff_B_jF5kPCUT9_1),.dout(n153),.clk(gclk));
	jnot g096(.din(w_n153_0[2]),.dout(n154),.clk(gclk));
	jand g097(.dina(w_n154_1[1]),.dinb(w_n144_1[2]),.dout(n155),.clk(gclk));
	jand g098(.dina(w_n155_0[2]),.dinb(w_n122_0[1]),.dout(n156),.clk(gclk));
	jxor g099(.dina(w_n156_0[1]),.dinb(w_G101_0[0]),.dout(w_dff_A_tgsGGwUG3_2),.clk(gclk));
	jnot g100(.din(w_n92_1[1]),.dout(n158),.clk(gclk));
	jand g101(.dina(w_n158_1[1]),.dinb(w_n74_1[0]),.dout(n159),.clk(gclk));
	jand g102(.dina(w_n159_1[1]),.dinb(w_n121_1[0]),.dout(n160),.clk(gclk));
	jxor g103(.dina(w_n142_0[0]),.dinb(w_G475_0[1]),.dout(n161),.clk(gclk));
	jand g104(.dina(w_n161_0[2]),.dinb(w_n132_0[1]),.dout(n162),.clk(gclk));
	jand g105(.dina(w_n162_0[1]),.dinb(w_n154_1[0]),.dout(n163),.clk(gclk));
	jand g106(.dina(w_n163_0[2]),.dinb(w_n160_0[1]),.dout(n164),.clk(gclk));
	jxor g107(.dina(w_n164_0[1]),.dinb(w_G104_0[0]),.dout(w_dff_A_1jvHz01S6_2),.clk(gclk));
	jxor g108(.dina(w_n131_0[0]),.dinb(w_G478_0[1]),.dout(n166),.clk(gclk));
	jand g109(.dina(w_n143_1[0]),.dinb(w_n166_1[1]),.dout(n167),.clk(gclk));
	jand g110(.dina(w_n167_0[1]),.dinb(w_n154_0[2]),.dout(n168),.clk(gclk));
	jand g111(.dina(w_n168_0[2]),.dinb(w_n160_0[0]),.dout(n169),.clk(gclk));
	jxor g112(.dina(w_n169_0[1]),.dinb(w_G107_0[0]),.dout(w_dff_A_B8eR28a40_2),.clk(gclk));
	jnot g113(.din(w_n60_0[0]),.dout(n171),.clk(gclk));
	jxor g114(.dina(w_n67_0[0]),.dinb(w_dff_B_pKaR8eaA2_1),.dout(n172),.clk(gclk));
	jand g115(.dina(w_n172_0[1]),.dinb(w_n70_1[0]),.dout(n173),.clk(gclk));
	jxor g116(.dina(w_n73_0[0]),.dinb(n173),.dout(n174),.clk(gclk));
	jand g117(.dina(w_n158_1[0]),.dinb(w_n174_1[1]),.dout(n175),.clk(gclk));
	jand g118(.dina(w_n175_0[1]),.dinb(w_n155_0[1]),.dout(n176),.clk(gclk));
	jand g119(.dina(n176),.dinb(w_n121_0[2]),.dout(n177),.clk(gclk));
	jxor g120(.dina(w_n177_0[1]),.dinb(w_G110_0[1]),.dout(w_dff_A_0f7i80Nd1_2),.clk(gclk));
	jand g121(.dina(w_n92_1[0]),.dinb(w_n174_1[0]),.dout(n179),.clk(gclk));
	jand g122(.dina(w_n179_0[2]),.dinb(w_n121_0[1]),.dout(n180),.clk(gclk));
	jor g123(.dina(w_n61_2[0]),.dinb(w_dff_B_GAw23NGM7_1),.dout(n181),.clk(gclk));
	jor g124(.dina(w_n181_0[2]),.dinb(w_n147_0[0]),.dout(n182),.clk(gclk));
	jand g125(.dina(w_dff_B_wOFWd6LP3_0),.dinb(w_n152_0[0]),.dout(n183),.clk(gclk));
	jnot g126(.din(w_n183_0[2]),.dout(n184),.clk(gclk));
	jand g127(.dina(w_n184_1[1]),.dinb(w_n167_0[0]),.dout(n185),.clk(gclk));
	jand g128(.dina(w_n185_0[2]),.dinb(w_n180_0[1]),.dout(n186),.clk(gclk));
	jxor g129(.dina(w_n186_0[1]),.dinb(w_G128_0[1]),.dout(w_dff_A_3yefOgGp2_2),.clk(gclk));
	jand g130(.dina(w_n161_0[1]),.dinb(w_n166_1[0]),.dout(n188),.clk(gclk));
	jand g131(.dina(w_n188_0[2]),.dinb(w_n184_1[0]),.dout(n189),.clk(gclk));
	jand g132(.dina(w_n189_0[1]),.dinb(w_n122_0[0]),.dout(n190),.clk(gclk));
	jxor g133(.dina(w_n190_0[1]),.dinb(w_G143_0[1]),.dout(w_dff_A_ehYWmLY91_2),.clk(gclk));
	jand g134(.dina(w_n184_0[2]),.dinb(w_n162_0[0]),.dout(n192),.clk(gclk));
	jand g135(.dina(w_n192_0[2]),.dinb(w_n180_0[0]),.dout(n193),.clk(gclk));
	jxor g136(.dina(w_n193_0[1]),.dinb(w_G146_0[0]),.dout(w_dff_A_CxV5R3S41_2),.clk(gclk));
	jnot g137(.din(w_G469_0[1]),.dout(n195),.clk(gclk));
	jxor g138(.dina(w_n118_0[0]),.dinb(w_dff_B_Jx9tTa653_1),.dout(n196),.clk(gclk));
	jand g139(.dina(w_n196_0[2]),.dinb(w_n112_1[0]),.dout(n197),.clk(gclk));
	jand g140(.dina(w_n197_1[1]),.dinb(w_n110_0[1]),.dout(n198),.clk(gclk));
	jand g141(.dina(w_n198_1[1]),.dinb(w_n93_0[1]),.dout(n199),.clk(gclk));
	jand g142(.dina(w_n199_0[1]),.dinb(w_n163_0[1]),.dout(n200),.clk(gclk));
	jxor g143(.dina(w_n200_0[1]),.dinb(w_G113_0[0]),.dout(w_dff_A_iA9pP22X1_2),.clk(gclk));
	jand g144(.dina(w_n199_0[0]),.dinb(w_n168_0[1]),.dout(n202),.clk(gclk));
	jxor g145(.dina(w_n202_0[1]),.dinb(w_G116_0[0]),.dout(w_dff_A_OvTispEG5_2),.clk(gclk));
	jand g146(.dina(w_n198_1[0]),.dinb(w_n179_0[1]),.dout(n204),.clk(gclk));
	jand g147(.dina(n204),.dinb(w_n155_0[0]),.dout(n205),.clk(gclk));
	jxor g148(.dina(w_n205_0[1]),.dinb(w_G119_0[0]),.dout(w_dff_A_Fko9CuZr6_2),.clk(gclk));
	jand g149(.dina(w_n197_1[0]),.dinb(w_n159_1[0]),.dout(n207),.clk(gclk));
	jand g150(.dina(w_n154_0[1]),.dinb(w_n110_0[0]),.dout(n208),.clk(gclk));
	jand g151(.dina(n208),.dinb(w_n188_0[1]),.dout(n209),.clk(gclk));
	jand g152(.dina(w_dff_B_VWqHtd9m4_0),.dinb(w_n207_0[1]),.dout(n210),.clk(gclk));
	jxor g153(.dina(w_n210_0[1]),.dinb(w_G122_0[1]),.dout(w_dff_A_VxBgzGut5_2),.clk(gclk));
	jand g154(.dina(w_n192_0[1]),.dinb(w_n175_0[0]),.dout(n212),.clk(gclk));
	jand g155(.dina(w_n212_0[1]),.dinb(w_n198_0[2]),.dout(n213),.clk(gclk));
	jxor g156(.dina(w_n213_0[1]),.dinb(w_G125_0[0]),.dout(w_dff_A_PCaNejM41_2),.clk(gclk));
	jnot g157(.din(w_n97_0[0]),.dout(n215),.clk(gclk));
	jxor g158(.dina(w_n108_0[0]),.dinb(w_dff_B_hXeRC8QT0_1),.dout(n216),.clk(gclk));
	jand g159(.dina(w_n216_0[2]),.dinb(w_n96_0[1]),.dout(n217),.clk(gclk));
	jand g160(.dina(w_n217_0[2]),.dinb(w_n120_0[0]),.dout(n218),.clk(gclk));
	jand g161(.dina(w_n218_1[1]),.dinb(w_n93_0[0]),.dout(n219),.clk(gclk));
	jand g162(.dina(w_n219_0[1]),.dinb(w_n192_0[0]),.dout(n220),.clk(gclk));
	jxor g163(.dina(w_n220_0[1]),.dinb(w_G131_0[0]),.dout(w_dff_A_XeL5ESXH3_2),.clk(gclk));
	jand g164(.dina(w_n219_0[0]),.dinb(w_n185_0[1]),.dout(n222),.clk(gclk));
	jxor g165(.dina(w_n222_0[1]),.dinb(w_G134_0[0]),.dout(w_dff_A_wxTTumbh8_2),.clk(gclk));
	jand g166(.dina(w_n184_0[1]),.dinb(w_n144_1[1]),.dout(n224),.clk(gclk));
	jand g167(.dina(w_dff_B_0kZ2z18R8_0),.dinb(w_n179_0[0]),.dout(n225),.clk(gclk));
	jand g168(.dina(n225),.dinb(w_n218_1[0]),.dout(n226),.clk(gclk));
	jxor g169(.dina(w_n226_0[1]),.dinb(w_G137_0[0]),.dout(w_dff_A_5ZGcPxwR6_2),.clk(gclk));
	jand g170(.dina(w_n218_0[2]),.dinb(w_n212_0[0]),.dout(n228),.clk(gclk));
	jxor g171(.dina(w_n228_0[1]),.dinb(w_G140_0[0]),.dout(w_dff_A_5MAg6puK2_2),.clk(gclk));
	jor g172(.dina(w_n177_0[0]),.dinb(w_n169_0[0]),.dout(n230),.clk(gclk));
	jor g173(.dina(w_n202_0[0]),.dinb(w_n164_0[0]),.dout(n231),.clk(gclk));
	jor g174(.dina(n231),.dinb(n230),.dout(n232),.clk(gclk));
	jor g175(.dina(w_n205_0[0]),.dinb(w_n156_0[0]),.dout(n233),.clk(gclk));
	jor g176(.dina(w_n210_0[0]),.dinb(w_n200_0[0]),.dout(n234),.clk(gclk));
	jor g177(.dina(n234),.dinb(n233),.dout(n235),.clk(gclk));
	jor g178(.dina(n235),.dinb(n232),.dout(n236),.clk(gclk));
	jor g179(.dina(w_n220_0[0]),.dinb(w_n193_0[0]),.dout(n237),.clk(gclk));
	jor g180(.dina(w_n222_0[0]),.dinb(w_n186_0[0]),.dout(n238),.clk(gclk));
	jor g181(.dina(n238),.dinb(n237),.dout(n239),.clk(gclk));
	jor g182(.dina(w_n228_0[0]),.dinb(w_n190_0[0]),.dout(n240),.clk(gclk));
	jor g183(.dina(w_n226_0[0]),.dinb(w_n213_0[0]),.dout(n241),.clk(gclk));
	jor g184(.dina(n241),.dinb(n240),.dout(n242),.clk(gclk));
	jor g185(.dina(n242),.dinb(n239),.dout(n243),.clk(gclk));
	jor g186(.dina(n243),.dinb(n236),.dout(n244),.clk(gclk));
	jor g187(.dina(w_n218_0[1]),.dinb(w_n198_0[1]),.dout(n245),.clk(gclk));
	jand g188(.dina(n245),.dinb(w_n144_1[0]),.dout(n246),.clk(gclk));
	jand g189(.dina(w_n217_0[1]),.dinb(w_n197_0[2]),.dout(n247),.clk(gclk));
	jxor g190(.dina(w_n143_0[2]),.dinb(w_n132_0[0]),.dout(n248),.clk(gclk));
	jand g191(.dina(w_dff_B_OjrxPkoz1_0),.dinb(n247),.dout(n249),.clk(gclk));
	jor g192(.dina(w_dff_B_1z3qikvk4_0),.dinb(n246),.dout(n250),.clk(gclk));
	jand g193(.dina(n250),.dinb(w_n159_0[2]),.dout(n251),.clk(gclk));
	jand g194(.dina(w_n217_0[0]),.dinb(w_n144_0[2]),.dout(n252),.clk(gclk));
	jor g195(.dina(w_n92_0[2]),.dinb(w_n174_0[2]),.dout(n253),.clk(gclk));
	jor g196(.dina(w_n158_0[2]),.dinb(w_n74_0[2]),.dout(n254),.clk(gclk));
	jand g197(.dina(w_n197_0[1]),.dinb(w_n254_1[1]),.dout(n255),.clk(gclk));
	jand g198(.dina(n255),.dinb(w_n253_0[2]),.dout(n256),.clk(gclk));
	jand g199(.dina(n256),.dinb(w_n252_0[1]),.dout(n257),.clk(gclk));
	jor g200(.dina(n257),.dinb(n251),.dout(n258),.clk(gclk));
	jand g201(.dina(n258),.dinb(w_n151_0[1]),.dout(n259),.clk(gclk));
	jxor g202(.dina(w_n112_0[2]),.dinb(w_n96_0[0]),.dout(n260),.clk(gclk));
	jand g203(.dina(n260),.dinb(w_n151_0[0]),.dout(n261),.clk(gclk));
	jand g204(.dina(w_dff_B_cnGFPP2K6_0),.dinb(w_n196_0[1]),.dout(n262),.clk(gclk));
	jand g205(.dina(n262),.dinb(w_n216_0[1]),.dout(n263),.clk(gclk));
	jand g206(.dina(w_n159_0[1]),.dinb(w_n144_0[1]),.dout(n264),.clk(gclk));
	jand g207(.dina(n264),.dinb(w_dff_B_k74NkQxL3_1),.dout(n265),.clk(gclk));
	jor g208(.dina(w_dff_B_WhPzckqG5_0),.dinb(n259),.dout(n266),.clk(gclk));
	jor g209(.dina(n266),.dinb(w_n244_2[2]),.dout(n267),.clk(gclk));
	jand g210(.dina(n267),.dinb(w_G952_0[1]),.dout(n268),.clk(gclk));
	jand g211(.dina(w_n252_0[0]),.dinb(w_n207_0[0]),.dout(n269),.clk(gclk));
	jor g212(.dina(n269),.dinb(w_G953_1[0]),.dout(n270),.clk(gclk));
	jor g213(.dina(w_dff_B_Dus5asfn5_0),.dinb(n268),.dout(w_dff_A_76IhHjB45_2),.clk(gclk));
	jnot g214(.din(w_n107_0[1]),.dout(n272),.clk(gclk));
	jor g215(.dina(w_n216_0[0]),.dinb(w_n95_0[1]),.dout(n273),.clk(gclk));
	jnot g216(.din(w_n112_0[1]),.dout(n274),.clk(gclk));
	jor g217(.dina(w_n196_0[0]),.dinb(w_n274_0[1]),.dout(n275),.clk(gclk));
	jor g218(.dina(w_n275_0[1]),.dinb(w_n273_0[2]),.dout(n276),.clk(gclk));
	jor g219(.dina(w_n253_0[1]),.dinb(w_n276_1[1]),.dout(n277),.clk(gclk));
	jnot g220(.din(w_n168_0[0]),.dout(n278),.clk(gclk));
	jor g221(.dina(w_n278_0[1]),.dinb(w_n277_0[1]),.dout(n279),.clk(gclk));
	jor g222(.dina(w_n161_0[0]),.dinb(w_n166_0[2]),.dout(n280),.clk(gclk));
	jor g223(.dina(w_n153_0[1]),.dinb(w_n280_0[1]),.dout(n281),.clk(gclk));
	jor g224(.dina(w_n92_0[1]),.dinb(w_n74_0[1]),.dout(n282),.clk(gclk));
	jor g225(.dina(w_n282_0[1]),.dinb(w_n281_0[2]),.dout(n283),.clk(gclk));
	jor g226(.dina(n283),.dinb(w_n276_1[0]),.dout(n284),.clk(gclk));
	jand g227(.dina(n284),.dinb(n279),.dout(n285),.clk(gclk));
	jnot g228(.din(w_n163_0[0]),.dout(n286),.clk(gclk));
	jor g229(.dina(w_n286_0[1]),.dinb(w_n277_0[0]),.dout(n287),.clk(gclk));
	jor g230(.dina(w_n158_0[1]),.dinb(w_n174_0[1]),.dout(n288),.clk(gclk));
	jor g231(.dina(w_n119_0[0]),.dinb(w_n274_0[0]),.dout(n289),.clk(gclk));
	jor g232(.dina(w_n289_0[1]),.dinb(w_n273_0[1]),.dout(n290),.clk(gclk));
	jor g233(.dina(w_n290_0[2]),.dinb(w_n288_0[2]),.dout(n291),.clk(gclk));
	jor g234(.dina(w_n291_0[1]),.dinb(w_n278_0[0]),.dout(n292),.clk(gclk));
	jand g235(.dina(n292),.dinb(n287),.dout(n293),.clk(gclk));
	jand g236(.dina(n293),.dinb(n285),.dout(n294),.clk(gclk));
	jor g237(.dina(w_n276_0[2]),.dinb(w_n288_0[1]),.dout(n295),.clk(gclk));
	jor g238(.dina(w_n281_0[1]),.dinb(w_n295_0[1]),.dout(n296),.clk(gclk));
	jor g239(.dina(w_n290_0[1]),.dinb(w_n254_1[0]),.dout(n297),.clk(gclk));
	jor g240(.dina(n297),.dinb(w_n281_0[0]),.dout(n298),.clk(gclk));
	jand g241(.dina(n298),.dinb(n296),.dout(n299),.clk(gclk));
	jor g242(.dina(w_n291_0[0]),.dinb(w_n286_0[0]),.dout(n300),.clk(gclk));
	jor g243(.dina(w_n289_0[0]),.dinb(w_n253_0[0]),.dout(n301),.clk(gclk));
	jnot g244(.din(w_n188_0[0]),.dout(n302),.clk(gclk));
	jor g245(.dina(w_n153_0[0]),.dinb(w_n273_0[0]),.dout(n303),.clk(gclk));
	jor g246(.dina(n303),.dinb(n302),.dout(n304),.clk(gclk));
	jor g247(.dina(w_dff_B_nCvU86gK5_0),.dinb(n301),.dout(n305),.clk(gclk));
	jand g248(.dina(n305),.dinb(n300),.dout(n306),.clk(gclk));
	jand g249(.dina(n306),.dinb(n299),.dout(n307),.clk(gclk));
	jand g250(.dina(n307),.dinb(n294),.dout(n308),.clk(gclk));
	jor g251(.dina(w_n254_0[2]),.dinb(w_n276_0[1]),.dout(n309),.clk(gclk));
	jor g252(.dina(w_n143_0[1]),.dinb(w_n166_0[1]),.dout(n310),.clk(gclk));
	jor g253(.dina(w_n183_0[1]),.dinb(n310),.dout(n311),.clk(gclk));
	jor g254(.dina(w_n311_0[2]),.dinb(w_n309_0[1]),.dout(n312),.clk(gclk));
	jor g255(.dina(w_n109_0[0]),.dinb(w_n95_0[0]),.dout(n313),.clk(gclk));
	jor g256(.dina(n313),.dinb(w_n275_0[0]),.dout(n314),.clk(gclk));
	jor g257(.dina(w_n314_0[2]),.dinb(w_n288_0[0]),.dout(n315),.clk(gclk));
	jor g258(.dina(w_n315_0[1]),.dinb(w_n311_0[1]),.dout(n316),.clk(gclk));
	jand g259(.dina(n316),.dinb(n312),.dout(n317),.clk(gclk));
	jnot g260(.din(w_n185_0[0]),.dout(n318),.clk(gclk));
	jor g261(.dina(w_n318_0[1]),.dinb(w_n309_0[0]),.dout(n319),.clk(gclk));
	jor g262(.dina(w_n315_0[0]),.dinb(w_n318_0[0]),.dout(n320),.clk(gclk));
	jand g263(.dina(n320),.dinb(n319),.dout(n321),.clk(gclk));
	jand g264(.dina(n321),.dinb(n317),.dout(n322),.clk(gclk));
	jnot g265(.din(w_n189_0[0]),.dout(n323),.clk(gclk));
	jor g266(.dina(w_dff_B_P1oev6OL7_0),.dinb(w_n295_0[0]),.dout(n324),.clk(gclk));
	jor g267(.dina(w_n311_0[0]),.dinb(w_n282_0[0]),.dout(n325),.clk(gclk));
	jor g268(.dina(w_n314_0[1]),.dinb(w_n325_0[1]),.dout(n326),.clk(gclk));
	jand g269(.dina(n326),.dinb(n324),.dout(n327),.clk(gclk));
	jor g270(.dina(w_n325_0[0]),.dinb(w_n290_0[0]),.dout(n328),.clk(gclk));
	jor g271(.dina(w_n183_0[0]),.dinb(w_n280_0[0]),.dout(n329),.clk(gclk));
	jor g272(.dina(w_dff_B_qRJjuky49_0),.dinb(w_n254_0[1]),.dout(n330),.clk(gclk));
	jor g273(.dina(n330),.dinb(w_n314_0[0]),.dout(n331),.clk(gclk));
	jand g274(.dina(n331),.dinb(n328),.dout(n332),.clk(gclk));
	jand g275(.dina(n332),.dinb(n327),.dout(n333),.clk(gclk));
	jand g276(.dina(n333),.dinb(n322),.dout(n334),.clk(gclk));
	jand g277(.dina(w_n334_0[1]),.dinb(w_n308_0[1]),.dout(n335),.clk(gclk));
	jand g278(.dina(w_G902_2[2]),.dinb(w_G210_0[0]),.dout(n336),.clk(gclk));
	jnot g279(.din(w_n336_0[1]),.dout(n337),.clk(gclk));
	jor g280(.dina(w_dff_B_dr0BwsTl6_0),.dinb(w_n335_2[1]),.dout(n338),.clk(gclk));
	jor g281(.dina(n338),.dinb(w_dff_B_8v4Z0UIu6_1),.dout(n339),.clk(gclk));
	jor g282(.dina(w_n61_1[2]),.dinb(w_G952_0[0]),.dout(n340),.clk(gclk));
	jand g283(.dina(w_n336_0[0]),.dinb(w_n244_2[1]),.dout(n341),.clk(gclk));
	jor g284(.dina(n341),.dinb(w_n107_0[0]),.dout(n342),.clk(gclk));
	jand g285(.dina(n342),.dinb(w_n340_2[1]),.dout(n343),.clk(gclk));
	jand g286(.dina(n343),.dinb(w_dff_B_0NusGIpQ1_1),.dout(G51),.clk(gclk));
	jnot g287(.din(w_n117_0[1]),.dout(n345),.clk(gclk));
	jand g288(.dina(w_G902_2[1]),.dinb(w_G469_0[0]),.dout(n346),.clk(gclk));
	jnot g289(.din(w_n346_0[1]),.dout(n347),.clk(gclk));
	jor g290(.dina(w_dff_B_Hz6UxcGC4_0),.dinb(w_n335_2[0]),.dout(n348),.clk(gclk));
	jor g291(.dina(n348),.dinb(w_dff_B_fuB4YbjP6_1),.dout(n349),.clk(gclk));
	jand g292(.dina(w_n346_0[0]),.dinb(w_n244_2[0]),.dout(n350),.clk(gclk));
	jor g293(.dina(n350),.dinb(w_n117_0[0]),.dout(n351),.clk(gclk));
	jand g294(.dina(n351),.dinb(w_n340_2[0]),.dout(n352),.clk(gclk));
	jand g295(.dina(n352),.dinb(w_dff_B_ANQgRK140_1),.dout(G54),.clk(gclk));
	jnot g296(.din(w_n141_0[1]),.dout(n354),.clk(gclk));
	jand g297(.dina(w_G902_2[0]),.dinb(w_G475_0[0]),.dout(n355),.clk(gclk));
	jnot g298(.din(w_n355_0[1]),.dout(n356),.clk(gclk));
	jor g299(.dina(w_dff_B_uPAk3PsE8_0),.dinb(w_n335_1[2]),.dout(n357),.clk(gclk));
	jor g300(.dina(n357),.dinb(w_dff_B_Slxm1lx63_1),.dout(n358),.clk(gclk));
	jand g301(.dina(w_n355_0[0]),.dinb(w_n244_1[2]),.dout(n359),.clk(gclk));
	jor g302(.dina(n359),.dinb(w_n141_0[0]),.dout(n360),.clk(gclk));
	jand g303(.dina(n360),.dinb(w_n340_1[2]),.dout(n361),.clk(gclk));
	jand g304(.dina(n361),.dinb(w_dff_B_SQh2gQdA3_1),.dout(G60),.clk(gclk));
	jnot g305(.din(w_n130_0[1]),.dout(n363),.clk(gclk));
	jand g306(.dina(w_G902_1[2]),.dinb(w_G478_0[0]),.dout(n364),.clk(gclk));
	jnot g307(.din(w_n364_0[1]),.dout(n365),.clk(gclk));
	jor g308(.dina(w_dff_B_0pIk17TD5_0),.dinb(w_n335_1[1]),.dout(n366),.clk(gclk));
	jor g309(.dina(n366),.dinb(w_dff_B_LUDNu2k16_1),.dout(n367),.clk(gclk));
	jand g310(.dina(w_n364_0[0]),.dinb(w_n244_1[1]),.dout(n368),.clk(gclk));
	jor g311(.dina(n368),.dinb(w_n130_0[0]),.dout(n369),.clk(gclk));
	jand g312(.dina(n369),.dinb(w_n340_1[1]),.dout(n370),.clk(gclk));
	jand g313(.dina(n370),.dinb(w_dff_B_kP0FXXRz4_1),.dout(G63),.clk(gclk));
	jand g314(.dina(w_G902_1[1]),.dinb(w_G217_0[0]),.dout(n372),.clk(gclk));
	jand g315(.dina(w_n372_0[1]),.dinb(w_n244_1[0]),.dout(n373),.clk(gclk));
	jor g316(.dina(n373),.dinb(w_n172_0[0]),.dout(n374),.clk(gclk));
	jnot g317(.din(w_n372_0[0]),.dout(n375),.clk(gclk));
	jor g318(.dina(w_dff_B_6ZN0m6354_0),.dinb(w_n335_1[0]),.dout(n376),.clk(gclk));
	jor g319(.dina(n376),.dinb(w_n68_0[0]),.dout(n377),.clk(gclk));
	jand g320(.dina(n377),.dinb(w_n340_1[0]),.dout(n378),.clk(gclk));
	jand g321(.dina(n378),.dinb(w_dff_B_hhH2xC3T0_1),.dout(G66),.clk(gclk));
	jnot g322(.din(w_n145_0[0]),.dout(n380),.clk(gclk));
	jor g323(.dina(w_n308_0[0]),.dinb(w_G953_0[2]),.dout(n381),.clk(gclk));
	jor g324(.dina(w_n61_1[1]),.dinb(w_G224_0[0]),.dout(n382),.clk(gclk));
	jand g325(.dina(w_dff_B_vItphulR1_0),.dinb(n381),.dout(n383),.clk(gclk));
	jxor g326(.dina(n383),.dinb(w_n103_0[0]),.dout(n384),.clk(gclk));
	jor g327(.dina(n384),.dinb(w_dff_B_PUcHH9zB0_1),.dout(w_dff_A_STzXy76t1_2),.clk(gclk));
	jor g328(.dina(w_n334_0[0]),.dinb(w_G953_0[1]),.dout(n386),.clk(gclk));
	jor g329(.dina(w_n61_1[0]),.dinb(w_G227_0[0]),.dout(n387),.clk(gclk));
	jand g330(.dina(n387),.dinb(w_n181_0[1]),.dout(n388),.clk(gclk));
	jand g331(.dina(w_dff_B_oKxb8BLI3_0),.dinb(n386),.dout(n389),.clk(gclk));
	jnot g332(.din(w_n181_0[0]),.dout(n390),.clk(gclk));
	jxor g333(.dina(w_n81_0[0]),.dinb(w_n59_0[0]),.dout(n391),.clk(gclk));
	jor g334(.dina(n391),.dinb(w_dff_B_vd9YvGa17_1),.dout(n392),.clk(gclk));
	jxor g335(.dina(w_dff_B_03H9PegJ1_0),.dinb(n389),.dout(w_dff_A_BblxUM767_2),.clk(gclk));
	jnot g336(.din(w_n90_0[1]),.dout(n394),.clk(gclk));
	jand g337(.dina(w_G902_1[0]),.dinb(w_G472_0[0]),.dout(n395),.clk(gclk));
	jnot g338(.din(w_n395_0[1]),.dout(n396),.clk(gclk));
	jor g339(.dina(w_dff_B_dl0Rx4Pp3_0),.dinb(w_n335_0[2]),.dout(n397),.clk(gclk));
	jor g340(.dina(n397),.dinb(w_dff_B_rg16n2yA1_1),.dout(n398),.clk(gclk));
	jand g341(.dina(w_n395_0[0]),.dinb(w_n244_0[2]),.dout(n399),.clk(gclk));
	jor g342(.dina(n399),.dinb(w_n90_0[0]),.dout(n400),.clk(gclk));
	jand g343(.dina(n400),.dinb(w_n340_0[2]),.dout(n401),.clk(gclk));
	jand g344(.dina(n401),.dinb(w_dff_B_bNBiZI2c2_1),.dout(G57),.clk(gclk));
	jspl3 jspl3_w_G101_0(.douta(w_dff_A_fjjRkyM94_0),.doutb(w_G101_0[1]),.doutc(w_dff_A_xokxmThT8_2),.din(w_dff_B_nhW2gutN0_3));
	jspl3 jspl3_w_G104_0(.douta(w_dff_A_PB4RuL8e9_0),.doutb(w_dff_A_ADaMUmKc6_1),.doutc(w_G104_0[2]),.din(G104));
	jspl3 jspl3_w_G107_0(.douta(w_dff_A_w6XTsMsq8_0),.doutb(w_G107_0[1]),.doutc(w_G107_0[2]),.din(G107));
	jspl3 jspl3_w_G110_0(.douta(w_G110_0[0]),.doutb(w_dff_A_6FnxbwUU6_1),.doutc(w_G110_0[2]),.din(G110));
	jspl jspl_w_G110_1(.douta(w_G110_1[0]),.doutb(w_dff_A_1FZCsts23_1),.din(w_G110_0[0]));
	jspl jspl_w_G113_0(.douta(w_dff_A_uGUkLdGk8_0),.doutb(w_G113_0[1]),.din(G113));
	jspl3 jspl3_w_G116_0(.douta(w_dff_A_AQxkgjvZ4_0),.doutb(w_G116_0[1]),.doutc(w_G116_0[2]),.din(G116));
	jspl3 jspl3_w_G119_0(.douta(w_dff_A_kWji1Z9g6_0),.doutb(w_G119_0[1]),.doutc(w_G119_0[2]),.din(G119));
	jspl3 jspl3_w_G122_0(.douta(w_G122_0[0]),.doutb(w_dff_A_EyY3UJfQ7_1),.doutc(w_dff_A_EeE4pWsK2_2),.din(G122));
	jspl jspl_w_G122_1(.douta(w_G122_1[0]),.doutb(w_dff_A_Xk15ibSQ5_1),.din(w_G122_0[0]));
	jspl3 jspl3_w_G125_0(.douta(w_dff_A_wEwstavb2_0),.doutb(w_dff_A_oICwdoW57_1),.doutc(w_G125_0[2]),.din(G125));
	jspl3 jspl3_w_G128_0(.douta(w_G128_0[0]),.doutb(w_dff_A_TOF1ISug0_1),.doutc(w_G128_0[2]),.din(G128));
	jspl jspl_w_G128_1(.douta(w_dff_A_uPQtcYLi3_0),.doutb(w_G128_1[1]),.din(w_G128_0[0]));
	jspl jspl_w_G131_0(.douta(w_dff_A_3crr4E687_0),.doutb(w_G131_0[1]),.din(G131));
	jspl3 jspl3_w_G134_0(.douta(w_dff_A_etucNoNa4_0),.doutb(w_G134_0[1]),.doutc(w_G134_0[2]),.din(G134));
	jspl3 jspl3_w_G137_0(.douta(w_dff_A_kaFOH6IU9_0),.doutb(w_G137_0[1]),.doutc(w_dff_A_0jUAIR0N0_2),.din(w_dff_B_TYwom6MH1_3));
	jspl3 jspl3_w_G140_0(.douta(w_dff_A_ErJwq7to0_0),.doutb(w_G140_0[1]),.doutc(w_G140_0[2]),.din(G140));
	jspl3 jspl3_w_G143_0(.douta(w_G143_0[0]),.doutb(w_dff_A_KvChh7Xe5_1),.doutc(w_dff_A_tAIPdC814_2),.din(G143));
	jspl jspl_w_G143_1(.douta(w_G143_1[0]),.doutb(w_G143_1[1]),.din(w_G143_0[0]));
	jspl3 jspl3_w_G146_0(.douta(w_dff_A_Ooj9orFX9_0),.doutb(w_G146_0[1]),.doutc(w_G146_0[2]),.din(G146));
	jspl3 jspl3_w_G210_0(.douta(w_G210_0[0]),.doutb(w_dff_A_jtdazSx98_1),.doutc(w_G210_0[2]),.din(G210));
	jspl jspl_w_G214_0(.douta(w_G214_0[0]),.doutb(w_dff_A_C8ITO4682_1),.din(G214));
	jspl3 jspl3_w_G217_0(.douta(w_G217_0[0]),.doutb(w_dff_A_UVej9Q6S7_1),.doutc(w_dff_A_cIAEdAzU8_2),.din(G217));
	jspl jspl_w_G221_0(.douta(w_G221_0[0]),.doutb(w_dff_A_WhLdinJl8_1),.din(G221));
	jspl jspl_w_G224_0(.douta(w_G224_0[0]),.doutb(w_G224_0[1]),.din(w_dff_B_8hXZiefv1_2));
	jspl jspl_w_G227_0(.douta(w_G227_0[0]),.doutb(w_G227_0[1]),.din(w_dff_B_skuoW42i7_2));
	jspl3 jspl3_w_G234_0(.douta(w_G234_0[0]),.doutb(w_dff_A_xGppPr3k5_1),.doutc(w_dff_A_3T0Mu2XP9_2),.din(G234));
	jspl3 jspl3_w_G237_0(.douta(w_G237_0[0]),.doutb(w_G237_0[1]),.doutc(w_G237_0[2]),.din(G237));
	jspl3 jspl3_w_G469_0(.douta(w_G469_0[0]),.doutb(w_G469_0[1]),.doutc(w_dff_A_TyI5Y8M08_2),.din(G469));
	jspl jspl_w_G472_0(.douta(w_G472_0[0]),.doutb(w_dff_A_J4ywwvin4_1),.din(G472));
	jspl3 jspl3_w_G475_0(.douta(w_G475_0[0]),.doutb(w_dff_A_CEab87fn1_1),.doutc(w_G475_0[2]),.din(G475));
	jspl3 jspl3_w_G478_0(.douta(w_G478_0[0]),.doutb(w_dff_A_WWtRK1vQ1_1),.doutc(w_G478_0[2]),.din(G478));
	jspl3 jspl3_w_G902_0(.douta(w_G902_0[0]),.doutb(w_G902_0[1]),.doutc(w_G902_0[2]),.din(G902));
	jspl3 jspl3_w_G902_1(.douta(w_G902_1[0]),.doutb(w_G902_1[1]),.doutc(w_G902_1[2]),.din(w_G902_0[0]));
	jspl3 jspl3_w_G902_2(.douta(w_G902_2[0]),.doutb(w_G902_2[1]),.doutc(w_G902_2[2]),.din(w_G902_0[1]));
	jspl3 jspl3_w_G902_3(.douta(w_G902_3[0]),.doutb(w_G902_3[1]),.doutc(w_dff_A_WylMPeS41_2),.din(w_G902_0[2]));
	jspl3 jspl3_w_G952_0(.douta(w_G952_0[0]),.doutb(w_dff_A_BsR5A8Rq5_1),.doutc(w_G952_0[2]),.din(w_dff_B_MxIFyWbc9_3));
	jspl3 jspl3_w_G953_0(.douta(w_G953_0[0]),.doutb(w_dff_A_NfEoZtfz9_1),.doutc(w_dff_A_MewQL7980_2),.din(G953));
	jspl3 jspl3_w_G953_1(.douta(w_dff_A_kfRW8fpl9_0),.doutb(w_G953_1[1]),.doutc(w_G953_1[2]),.din(w_G953_0[0]));
	jspl jspl_w_n59_0(.douta(w_dff_A_F0OlzLAD1_0),.doutb(w_n59_0[1]),.din(n59));
	jspl3 jspl3_w_n60_0(.douta(w_n60_0[0]),.doutb(w_n60_0[1]),.doutc(w_dff_A_qbrnQueL8_2),.din(n60));
	jspl3 jspl3_w_n61_0(.douta(w_n61_0[0]),.doutb(w_n61_0[1]),.doutc(w_n61_0[2]),.din(n61));
	jspl3 jspl3_w_n61_1(.douta(w_n61_1[0]),.doutb(w_n61_1[1]),.doutc(w_n61_1[2]),.din(w_n61_0[0]));
	jspl3 jspl3_w_n61_2(.douta(w_n61_2[0]),.doutb(w_n61_2[1]),.doutc(w_n61_2[2]),.din(w_n61_0[1]));
	jspl3 jspl3_w_n61_3(.douta(w_n61_3[0]),.doutb(w_n61_3[1]),.doutc(w_n61_3[2]),.din(w_n61_0[2]));
	jspl jspl_w_n62_0(.douta(w_n62_0[0]),.doutb(w_n62_0[1]),.din(n62));
	jspl jspl_w_n67_0(.douta(w_n67_0[0]),.doutb(w_n67_0[1]),.din(n67));
	jspl jspl_w_n68_0(.douta(w_dff_A_6AJDCdFE1_0),.doutb(w_n68_0[1]),.din(n68));
	jspl3 jspl3_w_n70_0(.douta(w_n70_0[0]),.doutb(w_dff_A_sq6nP6G67_1),.doutc(w_n70_0[2]),.din(n70));
	jspl3 jspl3_w_n70_1(.douta(w_dff_A_dkTleeez0_0),.doutb(w_n70_1[1]),.doutc(w_dff_A_iVMlshMV6_2),.din(w_n70_0[0]));
	jspl3 jspl3_w_n70_2(.douta(w_n70_2[0]),.doutb(w_n70_2[1]),.doutc(w_n70_2[2]),.din(w_n70_0[1]));
	jspl jspl_w_n70_3(.douta(w_dff_A_HEbrDUYk4_0),.doutb(w_n70_3[1]),.din(w_n70_0[2]));
	jspl jspl_w_n71_0(.douta(w_n71_0[0]),.doutb(w_n71_0[1]),.din(n71));
	jspl jspl_w_n73_0(.douta(w_n73_0[0]),.doutb(w_n73_0[1]),.din(w_dff_B_d1Qt6Vw90_2));
	jspl3 jspl3_w_n74_0(.douta(w_n74_0[0]),.doutb(w_n74_0[1]),.doutc(w_n74_0[2]),.din(n74));
	jspl jspl_w_n74_1(.douta(w_n74_1[0]),.doutb(w_n74_1[1]),.din(w_n74_0[0]));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_dff_A_wOV34ZYg8_1),.din(n77));
	jspl jspl_w_n79_0(.douta(w_n79_0[0]),.doutb(w_n79_0[1]),.din(n79));
	jspl3 jspl3_w_n81_0(.douta(w_n81_0[0]),.doutb(w_n81_0[1]),.doutc(w_n81_0[2]),.din(n81));
	jspl jspl_w_n82_0(.douta(w_n82_0[0]),.doutb(w_n82_0[1]),.din(n82));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_dff_A_zw6Yoo2x9_1),.din(n84));
	jspl jspl_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.din(n86));
	jspl3 jspl3_w_n90_0(.douta(w_dff_A_wSqvZeYI9_0),.doutb(w_n90_0[1]),.doutc(w_n90_0[2]),.din(n90));
	jspl3 jspl3_w_n92_0(.douta(w_n92_0[0]),.doutb(w_dff_A_IIDNdxzU7_1),.doutc(w_dff_A_1kIMQEqV3_2),.din(n92));
	jspl3 jspl3_w_n92_1(.douta(w_dff_A_OK5if8aX3_0),.doutb(w_n92_1[1]),.doutc(w_dff_A_XI8h2cgr0_2),.din(w_n92_0[0]));
	jspl3 jspl3_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.doutc(w_n93_0[2]),.din(n93));
	jspl jspl_w_n94_0(.douta(w_n94_0[0]),.doutb(w_n94_0[1]),.din(n94));
	jspl3 jspl3_w_n95_0(.douta(w_dff_A_ASA7AT1X9_0),.doutb(w_dff_A_xnFTH5ZX1_1),.doutc(w_n95_0[2]),.din(n95));
	jspl3 jspl3_w_n96_0(.douta(w_n96_0[0]),.doutb(w_dff_A_FvrCfnJD3_1),.doutc(w_dff_A_hDLlR9aU9_2),.din(n96));
	jspl jspl_w_n97_0(.douta(w_n97_0[0]),.doutb(w_dff_A_5QxyESWo5_1),.din(n97));
	jspl jspl_w_n101_0(.douta(w_n101_0[0]),.doutb(w_n101_0[1]),.din(n101));
	jspl jspl_w_n103_0(.douta(w_dff_A_Mjp2c5pP9_0),.doutb(w_n103_0[1]),.din(n103));
	jspl3 jspl3_w_n107_0(.douta(w_dff_A_ZhXSyGLz0_0),.doutb(w_n107_0[1]),.doutc(w_n107_0[2]),.din(n107));
	jspl jspl_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n109_0(.douta(w_n109_0[0]),.doutb(w_n109_0[1]),.din(n109));
	jspl3 jspl3_w_n110_0(.douta(w_n110_0[0]),.doutb(w_n110_0[1]),.doutc(w_n110_0[2]),.din(n110));
	jspl3 jspl3_w_n112_0(.douta(w_dff_A_tqhHZpRV0_0),.doutb(w_n112_0[1]),.doutc(w_n112_0[2]),.din(n112));
	jspl jspl_w_n112_1(.douta(w_n112_1[0]),.doutb(w_n112_1[1]),.din(w_n112_0[0]));
	jspl3 jspl3_w_n117_0(.douta(w_dff_A_O0ethJcU8_0),.doutb(w_n117_0[1]),.doutc(w_n117_0[2]),.din(n117));
	jspl jspl_w_n118_0(.douta(w_n118_0[0]),.doutb(w_n118_0[1]),.din(n118));
	jspl jspl_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.din(n119));
	jspl jspl_w_n120_0(.douta(w_n120_0[0]),.doutb(w_n120_0[1]),.din(n120));
	jspl3 jspl3_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.doutc(w_dff_A_fOwRUP1N3_2),.din(w_dff_B_W1OUvgBT0_3));
	jspl jspl_w_n121_1(.douta(w_n121_1[0]),.doutb(w_n121_1[1]),.din(w_n121_0[0]));
	jspl jspl_w_n122_0(.douta(w_n122_0[0]),.doutb(w_n122_0[1]),.din(n122));
	jspl3 jspl3_w_n130_0(.douta(w_dff_A_BIDb6lWi9_0),.doutb(w_n130_0[1]),.doutc(w_n130_0[2]),.din(n130));
	jspl jspl_w_n131_0(.douta(w_n131_0[0]),.doutb(w_n131_0[1]),.din(n131));
	jspl3 jspl3_w_n132_0(.douta(w_n132_0[0]),.doutb(w_n132_0[1]),.doutc(w_n132_0[2]),.din(n132));
	jspl3 jspl3_w_n141_0(.douta(w_dff_A_gV3TYRGf2_0),.doutb(w_n141_0[1]),.doutc(w_n141_0[2]),.din(n141));
	jspl jspl_w_n142_0(.douta(w_n142_0[0]),.doutb(w_n142_0[1]),.din(n142));
	jspl3 jspl3_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.doutc(w_n143_0[2]),.din(n143));
	jspl jspl_w_n143_1(.douta(w_n143_1[0]),.doutb(w_n143_1[1]),.din(w_n143_0[0]));
	jspl3 jspl3_w_n144_0(.douta(w_n144_0[0]),.doutb(w_dff_A_EGYRcwBO5_1),.doutc(w_n144_0[2]),.din(n144));
	jspl3 jspl3_w_n144_1(.douta(w_dff_A_ALtmhgTc6_0),.doutb(w_n144_1[1]),.doutc(w_n144_1[2]),.din(w_n144_0[0]));
	jspl jspl_w_n145_0(.douta(w_n145_0[0]),.doutb(w_n145_0[1]),.din(n145));
	jspl jspl_w_n146_0(.douta(w_n146_0[0]),.doutb(w_n146_0[1]),.din(n146));
	jspl jspl_w_n147_0(.douta(w_n147_0[0]),.doutb(w_n147_0[1]),.din(n147));
	jspl3 jspl3_w_n151_0(.douta(w_dff_A_AizOC6QN4_0),.doutb(w_dff_A_CJMSy18s4_1),.doutc(w_n151_0[2]),.din(n151));
	jspl jspl_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.din(n152));
	jspl3 jspl3_w_n153_0(.douta(w_dff_A_qAr5oImy2_0),.doutb(w_dff_A_SAYeAZFS1_1),.doutc(w_n153_0[2]),.din(n153));
	jspl3 jspl3_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.doutc(w_n154_0[2]),.din(w_dff_B_3tMQlBob3_3));
	jspl jspl_w_n154_1(.douta(w_n154_1[0]),.doutb(w_n154_1[1]),.din(w_n154_0[0]));
	jspl3 jspl3_w_n155_0(.douta(w_dff_A_L8M4JS3W9_0),.doutb(w_n155_0[1]),.doutc(w_dff_A_e0hOEbT09_2),.din(w_dff_B_XXYDJJC69_3));
	jspl jspl_w_n156_0(.douta(w_n156_0[0]),.doutb(w_n156_0[1]),.din(n156));
	jspl3 jspl3_w_n158_0(.douta(w_n158_0[0]),.doutb(w_n158_0[1]),.doutc(w_n158_0[2]),.din(w_dff_B_sJq7yOVI7_3));
	jspl jspl_w_n158_1(.douta(w_n158_1[0]),.doutb(w_n158_1[1]),.din(w_n158_0[0]));
	jspl3 jspl3_w_n159_0(.douta(w_n159_0[0]),.doutb(w_n159_0[1]),.doutc(w_dff_A_gtbJ1B1o4_2),.din(n159));
	jspl jspl_w_n159_1(.douta(w_n159_1[0]),.doutb(w_n159_1[1]),.din(w_n159_0[0]));
	jspl jspl_w_n160_0(.douta(w_n160_0[0]),.doutb(w_n160_0[1]),.din(n160));
	jspl3 jspl3_w_n161_0(.douta(w_n161_0[0]),.doutb(w_n161_0[1]),.doutc(w_n161_0[2]),.din(n161));
	jspl jspl_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.din(n162));
	jspl3 jspl3_w_n163_0(.douta(w_n163_0[0]),.doutb(w_dff_A_L4GXIG7G1_1),.doutc(w_dff_A_19nn0ZKO9_2),.din(n163));
	jspl jspl_w_n164_0(.douta(w_n164_0[0]),.doutb(w_n164_0[1]),.din(n164));
	jspl3 jspl3_w_n166_0(.douta(w_n166_0[0]),.doutb(w_n166_0[1]),.doutc(w_n166_0[2]),.din(n166));
	jspl jspl_w_n166_1(.douta(w_n166_1[0]),.doutb(w_n166_1[1]),.din(w_n166_0[0]));
	jspl jspl_w_n167_0(.douta(w_n167_0[0]),.doutb(w_n167_0[1]),.din(n167));
	jspl3 jspl3_w_n168_0(.douta(w_n168_0[0]),.doutb(w_dff_A_375026EZ7_1),.doutc(w_dff_A_MM0cDStJ0_2),.din(n168));
	jspl jspl_w_n169_0(.douta(w_n169_0[0]),.doutb(w_n169_0[1]),.din(n169));
	jspl jspl_w_n172_0(.douta(w_dff_A_4opZYrHl7_0),.doutb(w_n172_0[1]),.din(n172));
	jspl3 jspl3_w_n174_0(.douta(w_n174_0[0]),.doutb(w_n174_0[1]),.doutc(w_n174_0[2]),.din(n174));
	jspl jspl_w_n174_1(.douta(w_n174_1[0]),.doutb(w_n174_1[1]),.din(w_n174_0[0]));
	jspl jspl_w_n175_0(.douta(w_n175_0[0]),.doutb(w_n175_0[1]),.din(n175));
	jspl jspl_w_n177_0(.douta(w_n177_0[0]),.doutb(w_n177_0[1]),.din(n177));
	jspl3 jspl3_w_n179_0(.douta(w_n179_0[0]),.doutb(w_n179_0[1]),.doutc(w_n179_0[2]),.din(n179));
	jspl jspl_w_n180_0(.douta(w_n180_0[0]),.doutb(w_n180_0[1]),.din(n180));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(n181));
	jspl3 jspl3_w_n183_0(.douta(w_dff_A_EWqnEigz3_0),.doutb(w_dff_A_CpOdx5Gu0_1),.doutc(w_n183_0[2]),.din(n183));
	jspl3 jspl3_w_n184_0(.douta(w_n184_0[0]),.doutb(w_n184_0[1]),.doutc(w_n184_0[2]),.din(w_dff_B_IEPWR7JI3_3));
	jspl jspl_w_n184_1(.douta(w_n184_1[0]),.doutb(w_n184_1[1]),.din(w_n184_0[0]));
	jspl3 jspl3_w_n185_0(.douta(w_n185_0[0]),.doutb(w_dff_A_NtqSXtuH4_1),.doutc(w_dff_A_7XvFw0v89_2),.din(n185));
	jspl jspl_w_n186_0(.douta(w_n186_0[0]),.doutb(w_n186_0[1]),.din(n186));
	jspl3 jspl3_w_n188_0(.douta(w_n188_0[0]),.doutb(w_dff_A_REGWZ8k48_1),.doutc(w_n188_0[2]),.din(n188));
	jspl jspl_w_n189_0(.douta(w_n189_0[0]),.doutb(w_dff_A_eRcrnQaJ8_1),.din(n189));
	jspl jspl_w_n190_0(.douta(w_n190_0[0]),.doutb(w_n190_0[1]),.din(n190));
	jspl3 jspl3_w_n192_0(.douta(w_dff_A_jsAhbsnF8_0),.doutb(w_n192_0[1]),.doutc(w_dff_A_AqRVZuO56_2),.din(w_dff_B_xAj10c8M8_3));
	jspl jspl_w_n193_0(.douta(w_n193_0[0]),.doutb(w_n193_0[1]),.din(n193));
	jspl3 jspl3_w_n196_0(.douta(w_n196_0[0]),.doutb(w_n196_0[1]),.doutc(w_n196_0[2]),.din(n196));
	jspl3 jspl3_w_n197_0(.douta(w_n197_0[0]),.doutb(w_dff_A_HHgnVmET5_1),.doutc(w_n197_0[2]),.din(n197));
	jspl jspl_w_n197_1(.douta(w_dff_A_bIOKmwFE6_0),.doutb(w_n197_1[1]),.din(w_n197_0[0]));
	jspl3 jspl3_w_n198_0(.douta(w_dff_A_l0EIxeY21_0),.doutb(w_n198_0[1]),.doutc(w_dff_A_jQgXWgqB0_2),.din(n198));
	jspl jspl_w_n198_1(.douta(w_n198_1[0]),.doutb(w_n198_1[1]),.din(w_n198_0[0]));
	jspl jspl_w_n199_0(.douta(w_n199_0[0]),.doutb(w_n199_0[1]),.din(n199));
	jspl jspl_w_n200_0(.douta(w_n200_0[0]),.doutb(w_n200_0[1]),.din(n200));
	jspl jspl_w_n202_0(.douta(w_n202_0[0]),.doutb(w_n202_0[1]),.din(n202));
	jspl jspl_w_n205_0(.douta(w_n205_0[0]),.doutb(w_n205_0[1]),.din(n205));
	jspl jspl_w_n207_0(.douta(w_n207_0[0]),.doutb(w_n207_0[1]),.din(n207));
	jspl jspl_w_n210_0(.douta(w_n210_0[0]),.doutb(w_n210_0[1]),.din(n210));
	jspl jspl_w_n212_0(.douta(w_n212_0[0]),.doutb(w_n212_0[1]),.din(n212));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_n213_0[1]),.din(n213));
	jspl3 jspl3_w_n216_0(.douta(w_n216_0[0]),.doutb(w_dff_A_L7rbIXSV3_1),.doutc(w_n216_0[2]),.din(n216));
	jspl3 jspl3_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.doutc(w_n217_0[2]),.din(n217));
	jspl3 jspl3_w_n218_0(.douta(w_dff_A_2Qa4mDst8_0),.doutb(w_n218_0[1]),.doutc(w_dff_A_Q9G6vVgF3_2),.din(n218));
	jspl jspl_w_n218_1(.douta(w_dff_A_A0xHajm72_0),.doutb(w_n218_1[1]),.din(w_n218_0[0]));
	jspl jspl_w_n219_0(.douta(w_n219_0[0]),.doutb(w_n219_0[1]),.din(n219));
	jspl jspl_w_n220_0(.douta(w_n220_0[0]),.doutb(w_n220_0[1]),.din(n220));
	jspl jspl_w_n222_0(.douta(w_n222_0[0]),.doutb(w_n222_0[1]),.din(n222));
	jspl jspl_w_n226_0(.douta(w_n226_0[0]),.doutb(w_n226_0[1]),.din(n226));
	jspl jspl_w_n228_0(.douta(w_n228_0[0]),.doutb(w_n228_0[1]),.din(n228));
	jspl3 jspl3_w_n244_0(.douta(w_n244_0[0]),.doutb(w_n244_0[1]),.doutc(w_n244_0[2]),.din(n244));
	jspl3 jspl3_w_n244_1(.douta(w_n244_1[0]),.doutb(w_n244_1[1]),.doutc(w_n244_1[2]),.din(w_n244_0[0]));
	jspl3 jspl3_w_n244_2(.douta(w_n244_2[0]),.doutb(w_n244_2[1]),.doutc(w_n244_2[2]),.din(w_n244_0[1]));
	jspl jspl_w_n252_0(.douta(w_n252_0[0]),.doutb(w_dff_A_3ue1GCAa6_1),.din(w_dff_B_fXGOIhMh3_2));
	jspl3 jspl3_w_n253_0(.douta(w_n253_0[0]),.doutb(w_n253_0[1]),.doutc(w_dff_A_VuuFiaHe4_2),.din(n253));
	jspl3 jspl3_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.doutc(w_n254_0[2]),.din(n254));
	jspl jspl_w_n254_1(.douta(w_n254_1[0]),.doutb(w_n254_1[1]),.din(w_n254_0[0]));
	jspl3 jspl3_w_n273_0(.douta(w_n273_0[0]),.doutb(w_n273_0[1]),.doutc(w_n273_0[2]),.din(n273));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_n274_0[1]),.din(w_dff_B_pJ0ykcTy3_2));
	jspl jspl_w_n275_0(.douta(w_n275_0[0]),.doutb(w_n275_0[1]),.din(n275));
	jspl3 jspl3_w_n276_0(.douta(w_n276_0[0]),.doutb(w_n276_0[1]),.doutc(w_n276_0[2]),.din(w_dff_B_UXWqgLLL9_3));
	jspl jspl_w_n276_1(.douta(w_dff_A_yQejMPDK3_0),.doutb(w_n276_1[1]),.din(w_n276_0[0]));
	jspl jspl_w_n277_0(.douta(w_n277_0[0]),.doutb(w_n277_0[1]),.din(n277));
	jspl jspl_w_n278_0(.douta(w_n278_0[0]),.doutb(w_n278_0[1]),.din(w_dff_B_GQ5WKW4Z3_2));
	jspl jspl_w_n280_0(.douta(w_n280_0[0]),.doutb(w_n280_0[1]),.din(n280));
	jspl3 jspl3_w_n281_0(.douta(w_dff_A_XLhE6Odj0_0),.doutb(w_dff_A_sTQzwxcp3_1),.doutc(w_n281_0[2]),.din(w_dff_B_RiIbFyzW2_3));
	jspl jspl_w_n282_0(.douta(w_n282_0[0]),.doutb(w_n282_0[1]),.din(n282));
	jspl jspl_w_n286_0(.douta(w_n286_0[0]),.doutb(w_n286_0[1]),.din(w_dff_B_E2Ozntam6_2));
	jspl3 jspl3_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.doutc(w_n288_0[2]),.din(n288));
	jspl jspl_w_n289_0(.douta(w_dff_A_lnNYhLRA3_0),.doutb(w_n289_0[1]),.din(n289));
	jspl3 jspl3_w_n290_0(.douta(w_dff_A_n2Tcoh2U6_0),.doutb(w_n290_0[1]),.doutc(w_n290_0[2]),.din(w_dff_B_vBdGNBbj5_3));
	jspl jspl_w_n291_0(.douta(w_n291_0[0]),.doutb(w_n291_0[1]),.din(n291));
	jspl jspl_w_n295_0(.douta(w_n295_0[0]),.doutb(w_n295_0[1]),.din(n295));
	jspl jspl_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.din(n308));
	jspl jspl_w_n309_0(.douta(w_n309_0[0]),.doutb(w_n309_0[1]),.din(n309));
	jspl3 jspl3_w_n311_0(.douta(w_n311_0[0]),.doutb(w_dff_A_n1nyfuVj7_1),.doutc(w_dff_A_OZ8KK12W0_2),.din(w_dff_B_xgSN3V3V7_3));
	jspl3 jspl3_w_n314_0(.douta(w_dff_A_DjGGIK7h6_0),.doutb(w_dff_A_FKtcFAdn1_1),.doutc(w_n314_0[2]),.din(w_dff_B_IwweuLLc4_3));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl jspl_w_n318_0(.douta(w_n318_0[0]),.doutb(w_n318_0[1]),.din(w_dff_B_0F73FT6u8_2));
	jspl jspl_w_n325_0(.douta(w_n325_0[0]),.doutb(w_n325_0[1]),.din(n325));
	jspl jspl_w_n334_0(.douta(w_n334_0[0]),.doutb(w_n334_0[1]),.din(n334));
	jspl3 jspl3_w_n335_0(.douta(w_n335_0[0]),.doutb(w_n335_0[1]),.doutc(w_n335_0[2]),.din(n335));
	jspl3 jspl3_w_n335_1(.douta(w_n335_1[0]),.doutb(w_n335_1[1]),.doutc(w_n335_1[2]),.din(w_n335_0[0]));
	jspl jspl_w_n335_2(.douta(w_n335_2[0]),.doutb(w_n335_2[1]),.din(w_n335_0[1]));
	jspl jspl_w_n336_0(.douta(w_dff_A_wK8xo0ih4_0),.doutb(w_n336_0[1]),.din(n336));
	jspl3 jspl3_w_n340_0(.douta(w_n340_0[0]),.doutb(w_n340_0[1]),.doutc(w_n340_0[2]),.din(w_dff_B_XEK9xg8v1_3));
	jspl3 jspl3_w_n340_1(.douta(w_n340_1[0]),.doutb(w_n340_1[1]),.doutc(w_n340_1[2]),.din(w_n340_0[0]));
	jspl jspl_w_n340_2(.douta(w_n340_2[0]),.doutb(w_n340_2[1]),.din(w_n340_0[1]));
	jspl jspl_w_n346_0(.douta(w_dff_A_8J7Opxhj7_0),.doutb(w_n346_0[1]),.din(n346));
	jspl jspl_w_n355_0(.douta(w_dff_A_TB6WP7ZL0_0),.doutb(w_n355_0[1]),.din(n355));
	jspl jspl_w_n364_0(.douta(w_dff_A_CcABDC6X3_0),.doutb(w_n364_0[1]),.din(n364));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_dff_A_6mnfjbqs5_1),.din(n372));
	jspl jspl_w_n395_0(.douta(w_dff_A_U46uTslA6_0),.doutb(w_n395_0[1]),.din(n395));
	jdff dff_B_LWkzKn8m7_0(.din(n270),.dout(w_dff_B_LWkzKn8m7_0),.clk(gclk));
	jdff dff_B_Be0JuueW8_0(.din(w_dff_B_LWkzKn8m7_0),.dout(w_dff_B_Be0JuueW8_0),.clk(gclk));
	jdff dff_B_feKD8TAg8_0(.din(w_dff_B_Be0JuueW8_0),.dout(w_dff_B_feKD8TAg8_0),.clk(gclk));
	jdff dff_B_lkPmwJSH6_0(.din(w_dff_B_feKD8TAg8_0),.dout(w_dff_B_lkPmwJSH6_0),.clk(gclk));
	jdff dff_B_Dus5asfn5_0(.din(w_dff_B_lkPmwJSH6_0),.dout(w_dff_B_Dus5asfn5_0),.clk(gclk));
	jdff dff_B_Mh6gqh832_0(.din(n265),.dout(w_dff_B_Mh6gqh832_0),.clk(gclk));
	jdff dff_B_Iqg5cNID3_0(.din(w_dff_B_Mh6gqh832_0),.dout(w_dff_B_Iqg5cNID3_0),.clk(gclk));
	jdff dff_B_WhPzckqG5_0(.din(w_dff_B_Iqg5cNID3_0),.dout(w_dff_B_WhPzckqG5_0),.clk(gclk));
	jdff dff_B_Y1HlTLS96_1(.din(n263),.dout(w_dff_B_Y1HlTLS96_1),.clk(gclk));
	jdff dff_B_k74NkQxL3_1(.din(w_dff_B_Y1HlTLS96_1),.dout(w_dff_B_k74NkQxL3_1),.clk(gclk));
	jdff dff_B_3oUgQuJh8_0(.din(n261),.dout(w_dff_B_3oUgQuJh8_0),.clk(gclk));
	jdff dff_B_cnGFPP2K6_0(.din(w_dff_B_3oUgQuJh8_0),.dout(w_dff_B_cnGFPP2K6_0),.clk(gclk));
	jdff dff_A_3ue1GCAa6_1(.dout(w_n252_0[1]),.din(w_dff_A_3ue1GCAa6_1),.clk(gclk));
	jdff dff_B_pbGQtWSj8_2(.din(n252),.dout(w_dff_B_pbGQtWSj8_2),.clk(gclk));
	jdff dff_B_fXGOIhMh3_2(.din(w_dff_B_pbGQtWSj8_2),.dout(w_dff_B_fXGOIhMh3_2),.clk(gclk));
	jdff dff_B_1z3qikvk4_0(.din(n249),.dout(w_dff_B_1z3qikvk4_0),.clk(gclk));
	jdff dff_B_OjrxPkoz1_0(.din(n248),.dout(w_dff_B_OjrxPkoz1_0),.clk(gclk));
	jdff dff_B_0NusGIpQ1_1(.din(n339),.dout(w_dff_B_0NusGIpQ1_1),.clk(gclk));
	jdff dff_B_hdCoarWM4_1(.din(n272),.dout(w_dff_B_hdCoarWM4_1),.clk(gclk));
	jdff dff_B_DsJPWdlA2_1(.din(w_dff_B_hdCoarWM4_1),.dout(w_dff_B_DsJPWdlA2_1),.clk(gclk));
	jdff dff_B_u0O1DsPH2_1(.din(w_dff_B_DsJPWdlA2_1),.dout(w_dff_B_u0O1DsPH2_1),.clk(gclk));
	jdff dff_B_JakKkpps1_1(.din(w_dff_B_u0O1DsPH2_1),.dout(w_dff_B_JakKkpps1_1),.clk(gclk));
	jdff dff_B_E6lrRoBW0_1(.din(w_dff_B_JakKkpps1_1),.dout(w_dff_B_E6lrRoBW0_1),.clk(gclk));
	jdff dff_B_VuZcRjQM4_1(.din(w_dff_B_E6lrRoBW0_1),.dout(w_dff_B_VuZcRjQM4_1),.clk(gclk));
	jdff dff_B_q5HVwXmD5_1(.din(w_dff_B_VuZcRjQM4_1),.dout(w_dff_B_q5HVwXmD5_1),.clk(gclk));
	jdff dff_B_13uuITfG2_1(.din(w_dff_B_q5HVwXmD5_1),.dout(w_dff_B_13uuITfG2_1),.clk(gclk));
	jdff dff_B_QL5mamIM6_1(.din(w_dff_B_13uuITfG2_1),.dout(w_dff_B_QL5mamIM6_1),.clk(gclk));
	jdff dff_B_LnVkTcjl3_1(.din(w_dff_B_QL5mamIM6_1),.dout(w_dff_B_LnVkTcjl3_1),.clk(gclk));
	jdff dff_B_8v4Z0UIu6_1(.din(w_dff_B_LnVkTcjl3_1),.dout(w_dff_B_8v4Z0UIu6_1),.clk(gclk));
	jdff dff_B_7u0DeLhZ9_0(.din(n337),.dout(w_dff_B_7u0DeLhZ9_0),.clk(gclk));
	jdff dff_B_lYykZK1E7_0(.din(w_dff_B_7u0DeLhZ9_0),.dout(w_dff_B_lYykZK1E7_0),.clk(gclk));
	jdff dff_B_fKrfXaD88_0(.din(w_dff_B_lYykZK1E7_0),.dout(w_dff_B_fKrfXaD88_0),.clk(gclk));
	jdff dff_B_wKbd32w60_0(.din(w_dff_B_fKrfXaD88_0),.dout(w_dff_B_wKbd32w60_0),.clk(gclk));
	jdff dff_B_FuQIJ1E44_0(.din(w_dff_B_wKbd32w60_0),.dout(w_dff_B_FuQIJ1E44_0),.clk(gclk));
	jdff dff_B_H9cCylnh8_0(.din(w_dff_B_FuQIJ1E44_0),.dout(w_dff_B_H9cCylnh8_0),.clk(gclk));
	jdff dff_B_uuXwp87y5_0(.din(w_dff_B_H9cCylnh8_0),.dout(w_dff_B_uuXwp87y5_0),.clk(gclk));
	jdff dff_B_WQ0cvmw84_0(.din(w_dff_B_uuXwp87y5_0),.dout(w_dff_B_WQ0cvmw84_0),.clk(gclk));
	jdff dff_B_i2Ue4JlN0_0(.din(w_dff_B_WQ0cvmw84_0),.dout(w_dff_B_i2Ue4JlN0_0),.clk(gclk));
	jdff dff_B_OXR17nlL7_0(.din(w_dff_B_i2Ue4JlN0_0),.dout(w_dff_B_OXR17nlL7_0),.clk(gclk));
	jdff dff_B_thlH4yks4_0(.din(w_dff_B_OXR17nlL7_0),.dout(w_dff_B_thlH4yks4_0),.clk(gclk));
	jdff dff_B_mimsbmED9_0(.din(w_dff_B_thlH4yks4_0),.dout(w_dff_B_mimsbmED9_0),.clk(gclk));
	jdff dff_B_DzktRynN5_0(.din(w_dff_B_mimsbmED9_0),.dout(w_dff_B_DzktRynN5_0),.clk(gclk));
	jdff dff_B_dr0BwsTl6_0(.din(w_dff_B_DzktRynN5_0),.dout(w_dff_B_dr0BwsTl6_0),.clk(gclk));
	jdff dff_A_PWhc653A2_0(.dout(w_n336_0[0]),.din(w_dff_A_PWhc653A2_0),.clk(gclk));
	jdff dff_A_T55N1r1Y9_0(.dout(w_dff_A_PWhc653A2_0),.din(w_dff_A_T55N1r1Y9_0),.clk(gclk));
	jdff dff_A_KFFnJt7d9_0(.dout(w_dff_A_T55N1r1Y9_0),.din(w_dff_A_KFFnJt7d9_0),.clk(gclk));
	jdff dff_A_s8VJWkIA8_0(.dout(w_dff_A_KFFnJt7d9_0),.din(w_dff_A_s8VJWkIA8_0),.clk(gclk));
	jdff dff_A_GwVN9RiE3_0(.dout(w_dff_A_s8VJWkIA8_0),.din(w_dff_A_GwVN9RiE3_0),.clk(gclk));
	jdff dff_A_jRpf3phO1_0(.dout(w_dff_A_GwVN9RiE3_0),.din(w_dff_A_jRpf3phO1_0),.clk(gclk));
	jdff dff_A_E9kIB8ML0_0(.dout(w_dff_A_jRpf3phO1_0),.din(w_dff_A_E9kIB8ML0_0),.clk(gclk));
	jdff dff_A_6So5Xe162_0(.dout(w_dff_A_E9kIB8ML0_0),.din(w_dff_A_6So5Xe162_0),.clk(gclk));
	jdff dff_A_vj5pcntQ1_0(.dout(w_dff_A_6So5Xe162_0),.din(w_dff_A_vj5pcntQ1_0),.clk(gclk));
	jdff dff_A_58eoaMGF4_0(.dout(w_dff_A_vj5pcntQ1_0),.din(w_dff_A_58eoaMGF4_0),.clk(gclk));
	jdff dff_A_z9WPkE0c8_0(.dout(w_dff_A_58eoaMGF4_0),.din(w_dff_A_z9WPkE0c8_0),.clk(gclk));
	jdff dff_A_Tns3PYmN2_0(.dout(w_dff_A_z9WPkE0c8_0),.din(w_dff_A_Tns3PYmN2_0),.clk(gclk));
	jdff dff_A_Xs4reAsg9_0(.dout(w_dff_A_Tns3PYmN2_0),.din(w_dff_A_Xs4reAsg9_0),.clk(gclk));
	jdff dff_A_yE2KYfAC7_0(.dout(w_dff_A_Xs4reAsg9_0),.din(w_dff_A_yE2KYfAC7_0),.clk(gclk));
	jdff dff_A_wK8xo0ih4_0(.dout(w_dff_A_yE2KYfAC7_0),.din(w_dff_A_wK8xo0ih4_0),.clk(gclk));
	jdff dff_B_ANQgRK140_1(.din(n349),.dout(w_dff_B_ANQgRK140_1),.clk(gclk));
	jdff dff_B_4EnfuEyv7_1(.din(n345),.dout(w_dff_B_4EnfuEyv7_1),.clk(gclk));
	jdff dff_B_Oro06xku4_1(.din(w_dff_B_4EnfuEyv7_1),.dout(w_dff_B_Oro06xku4_1),.clk(gclk));
	jdff dff_B_XzmnYfwm7_1(.din(w_dff_B_Oro06xku4_1),.dout(w_dff_B_XzmnYfwm7_1),.clk(gclk));
	jdff dff_B_o5wRrX1u5_1(.din(w_dff_B_XzmnYfwm7_1),.dout(w_dff_B_o5wRrX1u5_1),.clk(gclk));
	jdff dff_B_DOqRJtRL1_1(.din(w_dff_B_o5wRrX1u5_1),.dout(w_dff_B_DOqRJtRL1_1),.clk(gclk));
	jdff dff_B_RB58VdCH1_1(.din(w_dff_B_DOqRJtRL1_1),.dout(w_dff_B_RB58VdCH1_1),.clk(gclk));
	jdff dff_B_CRDkqrFk2_1(.din(w_dff_B_RB58VdCH1_1),.dout(w_dff_B_CRDkqrFk2_1),.clk(gclk));
	jdff dff_B_8GAmCsxX6_1(.din(w_dff_B_CRDkqrFk2_1),.dout(w_dff_B_8GAmCsxX6_1),.clk(gclk));
	jdff dff_B_Rd0PAMwQ7_1(.din(w_dff_B_8GAmCsxX6_1),.dout(w_dff_B_Rd0PAMwQ7_1),.clk(gclk));
	jdff dff_B_jV8dr14K4_1(.din(w_dff_B_Rd0PAMwQ7_1),.dout(w_dff_B_jV8dr14K4_1),.clk(gclk));
	jdff dff_B_fuB4YbjP6_1(.din(w_dff_B_jV8dr14K4_1),.dout(w_dff_B_fuB4YbjP6_1),.clk(gclk));
	jdff dff_B_74JaBsIo5_0(.din(n347),.dout(w_dff_B_74JaBsIo5_0),.clk(gclk));
	jdff dff_B_euM955On1_0(.din(w_dff_B_74JaBsIo5_0),.dout(w_dff_B_euM955On1_0),.clk(gclk));
	jdff dff_B_cQbWAykn8_0(.din(w_dff_B_euM955On1_0),.dout(w_dff_B_cQbWAykn8_0),.clk(gclk));
	jdff dff_B_luXDGkTp1_0(.din(w_dff_B_cQbWAykn8_0),.dout(w_dff_B_luXDGkTp1_0),.clk(gclk));
	jdff dff_B_05lhf9A88_0(.din(w_dff_B_luXDGkTp1_0),.dout(w_dff_B_05lhf9A88_0),.clk(gclk));
	jdff dff_B_sZFyscMk1_0(.din(w_dff_B_05lhf9A88_0),.dout(w_dff_B_sZFyscMk1_0),.clk(gclk));
	jdff dff_B_1vOjhKA85_0(.din(w_dff_B_sZFyscMk1_0),.dout(w_dff_B_1vOjhKA85_0),.clk(gclk));
	jdff dff_B_E0OyvjAW3_0(.din(w_dff_B_1vOjhKA85_0),.dout(w_dff_B_E0OyvjAW3_0),.clk(gclk));
	jdff dff_B_hPzftarw4_0(.din(w_dff_B_E0OyvjAW3_0),.dout(w_dff_B_hPzftarw4_0),.clk(gclk));
	jdff dff_B_9TK02zqz0_0(.din(w_dff_B_hPzftarw4_0),.dout(w_dff_B_9TK02zqz0_0),.clk(gclk));
	jdff dff_B_zCSJrkjM3_0(.din(w_dff_B_9TK02zqz0_0),.dout(w_dff_B_zCSJrkjM3_0),.clk(gclk));
	jdff dff_B_0eEjCKXP5_0(.din(w_dff_B_zCSJrkjM3_0),.dout(w_dff_B_0eEjCKXP5_0),.clk(gclk));
	jdff dff_B_b6LaWH4c2_0(.din(w_dff_B_0eEjCKXP5_0),.dout(w_dff_B_b6LaWH4c2_0),.clk(gclk));
	jdff dff_B_Hz6UxcGC4_0(.din(w_dff_B_b6LaWH4c2_0),.dout(w_dff_B_Hz6UxcGC4_0),.clk(gclk));
	jdff dff_A_WHafdpbG5_0(.dout(w_n346_0[0]),.din(w_dff_A_WHafdpbG5_0),.clk(gclk));
	jdff dff_A_M81hBMB46_0(.dout(w_dff_A_WHafdpbG5_0),.din(w_dff_A_M81hBMB46_0),.clk(gclk));
	jdff dff_A_mFIrA8nf3_0(.dout(w_dff_A_M81hBMB46_0),.din(w_dff_A_mFIrA8nf3_0),.clk(gclk));
	jdff dff_A_SKUTIPTp3_0(.dout(w_dff_A_mFIrA8nf3_0),.din(w_dff_A_SKUTIPTp3_0),.clk(gclk));
	jdff dff_A_ZUbskobr6_0(.dout(w_dff_A_SKUTIPTp3_0),.din(w_dff_A_ZUbskobr6_0),.clk(gclk));
	jdff dff_A_FIT1i4QH2_0(.dout(w_dff_A_ZUbskobr6_0),.din(w_dff_A_FIT1i4QH2_0),.clk(gclk));
	jdff dff_A_xWOzoEwx6_0(.dout(w_dff_A_FIT1i4QH2_0),.din(w_dff_A_xWOzoEwx6_0),.clk(gclk));
	jdff dff_A_SVMe4flY6_0(.dout(w_dff_A_xWOzoEwx6_0),.din(w_dff_A_SVMe4flY6_0),.clk(gclk));
	jdff dff_A_J79ltrwf6_0(.dout(w_dff_A_SVMe4flY6_0),.din(w_dff_A_J79ltrwf6_0),.clk(gclk));
	jdff dff_A_mCJiZiea9_0(.dout(w_dff_A_J79ltrwf6_0),.din(w_dff_A_mCJiZiea9_0),.clk(gclk));
	jdff dff_A_2w90mkWU1_0(.dout(w_dff_A_mCJiZiea9_0),.din(w_dff_A_2w90mkWU1_0),.clk(gclk));
	jdff dff_A_4SjneQ7j3_0(.dout(w_dff_A_2w90mkWU1_0),.din(w_dff_A_4SjneQ7j3_0),.clk(gclk));
	jdff dff_A_3VrIdUWG7_0(.dout(w_dff_A_4SjneQ7j3_0),.din(w_dff_A_3VrIdUWG7_0),.clk(gclk));
	jdff dff_A_TKIxaGy19_0(.dout(w_dff_A_3VrIdUWG7_0),.din(w_dff_A_TKIxaGy19_0),.clk(gclk));
	jdff dff_A_8J7Opxhj7_0(.dout(w_dff_A_TKIxaGy19_0),.din(w_dff_A_8J7Opxhj7_0),.clk(gclk));
	jdff dff_B_SQh2gQdA3_1(.din(n358),.dout(w_dff_B_SQh2gQdA3_1),.clk(gclk));
	jdff dff_B_BJ6Rooop7_1(.din(n354),.dout(w_dff_B_BJ6Rooop7_1),.clk(gclk));
	jdff dff_B_748Igfu64_1(.din(w_dff_B_BJ6Rooop7_1),.dout(w_dff_B_748Igfu64_1),.clk(gclk));
	jdff dff_B_DcC6rqkx2_1(.din(w_dff_B_748Igfu64_1),.dout(w_dff_B_DcC6rqkx2_1),.clk(gclk));
	jdff dff_B_JVUOG1LR0_1(.din(w_dff_B_DcC6rqkx2_1),.dout(w_dff_B_JVUOG1LR0_1),.clk(gclk));
	jdff dff_B_xKDCvSCA8_1(.din(w_dff_B_JVUOG1LR0_1),.dout(w_dff_B_xKDCvSCA8_1),.clk(gclk));
	jdff dff_B_6kyTUGvp2_1(.din(w_dff_B_xKDCvSCA8_1),.dout(w_dff_B_6kyTUGvp2_1),.clk(gclk));
	jdff dff_B_OAGK93mI9_1(.din(w_dff_B_6kyTUGvp2_1),.dout(w_dff_B_OAGK93mI9_1),.clk(gclk));
	jdff dff_B_hypuAYjm0_1(.din(w_dff_B_OAGK93mI9_1),.dout(w_dff_B_hypuAYjm0_1),.clk(gclk));
	jdff dff_B_6pDOdZjL4_1(.din(w_dff_B_hypuAYjm0_1),.dout(w_dff_B_6pDOdZjL4_1),.clk(gclk));
	jdff dff_B_7hEdY94K4_1(.din(w_dff_B_6pDOdZjL4_1),.dout(w_dff_B_7hEdY94K4_1),.clk(gclk));
	jdff dff_B_Slxm1lx63_1(.din(w_dff_B_7hEdY94K4_1),.dout(w_dff_B_Slxm1lx63_1),.clk(gclk));
	jdff dff_B_BBvIKtNP1_0(.din(n356),.dout(w_dff_B_BBvIKtNP1_0),.clk(gclk));
	jdff dff_B_xciTNEE36_0(.din(w_dff_B_BBvIKtNP1_0),.dout(w_dff_B_xciTNEE36_0),.clk(gclk));
	jdff dff_B_Ro86NhZw8_0(.din(w_dff_B_xciTNEE36_0),.dout(w_dff_B_Ro86NhZw8_0),.clk(gclk));
	jdff dff_B_jwgBJArJ6_0(.din(w_dff_B_Ro86NhZw8_0),.dout(w_dff_B_jwgBJArJ6_0),.clk(gclk));
	jdff dff_B_jGNFm7hT8_0(.din(w_dff_B_jwgBJArJ6_0),.dout(w_dff_B_jGNFm7hT8_0),.clk(gclk));
	jdff dff_B_dd85IcJm3_0(.din(w_dff_B_jGNFm7hT8_0),.dout(w_dff_B_dd85IcJm3_0),.clk(gclk));
	jdff dff_B_udz6a51B2_0(.din(w_dff_B_dd85IcJm3_0),.dout(w_dff_B_udz6a51B2_0),.clk(gclk));
	jdff dff_B_8R9AMw6g2_0(.din(w_dff_B_udz6a51B2_0),.dout(w_dff_B_8R9AMw6g2_0),.clk(gclk));
	jdff dff_B_BuFks82O4_0(.din(w_dff_B_8R9AMw6g2_0),.dout(w_dff_B_BuFks82O4_0),.clk(gclk));
	jdff dff_B_Imz9GHSJ2_0(.din(w_dff_B_BuFks82O4_0),.dout(w_dff_B_Imz9GHSJ2_0),.clk(gclk));
	jdff dff_B_xxDbMDP82_0(.din(w_dff_B_Imz9GHSJ2_0),.dout(w_dff_B_xxDbMDP82_0),.clk(gclk));
	jdff dff_B_D7WhIya89_0(.din(w_dff_B_xxDbMDP82_0),.dout(w_dff_B_D7WhIya89_0),.clk(gclk));
	jdff dff_B_zyeN6HZ17_0(.din(w_dff_B_D7WhIya89_0),.dout(w_dff_B_zyeN6HZ17_0),.clk(gclk));
	jdff dff_B_uPAk3PsE8_0(.din(w_dff_B_zyeN6HZ17_0),.dout(w_dff_B_uPAk3PsE8_0),.clk(gclk));
	jdff dff_A_dXEIWgDr5_0(.dout(w_n355_0[0]),.din(w_dff_A_dXEIWgDr5_0),.clk(gclk));
	jdff dff_A_UblRcr5H7_0(.dout(w_dff_A_dXEIWgDr5_0),.din(w_dff_A_UblRcr5H7_0),.clk(gclk));
	jdff dff_A_GbX3sqRV6_0(.dout(w_dff_A_UblRcr5H7_0),.din(w_dff_A_GbX3sqRV6_0),.clk(gclk));
	jdff dff_A_jNwtQAJy2_0(.dout(w_dff_A_GbX3sqRV6_0),.din(w_dff_A_jNwtQAJy2_0),.clk(gclk));
	jdff dff_A_SBVTTQf23_0(.dout(w_dff_A_jNwtQAJy2_0),.din(w_dff_A_SBVTTQf23_0),.clk(gclk));
	jdff dff_A_txZ7Byz38_0(.dout(w_dff_A_SBVTTQf23_0),.din(w_dff_A_txZ7Byz38_0),.clk(gclk));
	jdff dff_A_8uVVB5dg1_0(.dout(w_dff_A_txZ7Byz38_0),.din(w_dff_A_8uVVB5dg1_0),.clk(gclk));
	jdff dff_A_3CkFEYoY8_0(.dout(w_dff_A_8uVVB5dg1_0),.din(w_dff_A_3CkFEYoY8_0),.clk(gclk));
	jdff dff_A_EYRVDabA5_0(.dout(w_dff_A_3CkFEYoY8_0),.din(w_dff_A_EYRVDabA5_0),.clk(gclk));
	jdff dff_A_PsEwy2V65_0(.dout(w_dff_A_EYRVDabA5_0),.din(w_dff_A_PsEwy2V65_0),.clk(gclk));
	jdff dff_A_3G1Q4sZu6_0(.dout(w_dff_A_PsEwy2V65_0),.din(w_dff_A_3G1Q4sZu6_0),.clk(gclk));
	jdff dff_A_fZa86WO57_0(.dout(w_dff_A_3G1Q4sZu6_0),.din(w_dff_A_fZa86WO57_0),.clk(gclk));
	jdff dff_A_DBUrhVvv0_0(.dout(w_dff_A_fZa86WO57_0),.din(w_dff_A_DBUrhVvv0_0),.clk(gclk));
	jdff dff_A_amj7g5Eo1_0(.dout(w_dff_A_DBUrhVvv0_0),.din(w_dff_A_amj7g5Eo1_0),.clk(gclk));
	jdff dff_A_TB6WP7ZL0_0(.dout(w_dff_A_amj7g5Eo1_0),.din(w_dff_A_TB6WP7ZL0_0),.clk(gclk));
	jdff dff_B_kP0FXXRz4_1(.din(n367),.dout(w_dff_B_kP0FXXRz4_1),.clk(gclk));
	jdff dff_B_v6jcs1Tw1_1(.din(n363),.dout(w_dff_B_v6jcs1Tw1_1),.clk(gclk));
	jdff dff_B_7SdlZiU25_1(.din(w_dff_B_v6jcs1Tw1_1),.dout(w_dff_B_7SdlZiU25_1),.clk(gclk));
	jdff dff_B_IcRwO1FJ6_1(.din(w_dff_B_7SdlZiU25_1),.dout(w_dff_B_IcRwO1FJ6_1),.clk(gclk));
	jdff dff_B_gQBk2m2P4_1(.din(w_dff_B_IcRwO1FJ6_1),.dout(w_dff_B_gQBk2m2P4_1),.clk(gclk));
	jdff dff_B_iVlEzbxa0_1(.din(w_dff_B_gQBk2m2P4_1),.dout(w_dff_B_iVlEzbxa0_1),.clk(gclk));
	jdff dff_B_p0rppZQ87_1(.din(w_dff_B_iVlEzbxa0_1),.dout(w_dff_B_p0rppZQ87_1),.clk(gclk));
	jdff dff_B_2nxCeAFo6_1(.din(w_dff_B_p0rppZQ87_1),.dout(w_dff_B_2nxCeAFo6_1),.clk(gclk));
	jdff dff_B_bzqeEy5W3_1(.din(w_dff_B_2nxCeAFo6_1),.dout(w_dff_B_bzqeEy5W3_1),.clk(gclk));
	jdff dff_B_ic9vLmhp3_1(.din(w_dff_B_bzqeEy5W3_1),.dout(w_dff_B_ic9vLmhp3_1),.clk(gclk));
	jdff dff_B_233cQcXb5_1(.din(w_dff_B_ic9vLmhp3_1),.dout(w_dff_B_233cQcXb5_1),.clk(gclk));
	jdff dff_B_LUDNu2k16_1(.din(w_dff_B_233cQcXb5_1),.dout(w_dff_B_LUDNu2k16_1),.clk(gclk));
	jdff dff_B_3laqQ3w85_0(.din(n365),.dout(w_dff_B_3laqQ3w85_0),.clk(gclk));
	jdff dff_B_MRvqB5mu9_0(.din(w_dff_B_3laqQ3w85_0),.dout(w_dff_B_MRvqB5mu9_0),.clk(gclk));
	jdff dff_B_SzAMrhsn1_0(.din(w_dff_B_MRvqB5mu9_0),.dout(w_dff_B_SzAMrhsn1_0),.clk(gclk));
	jdff dff_B_tsYHOX1q3_0(.din(w_dff_B_SzAMrhsn1_0),.dout(w_dff_B_tsYHOX1q3_0),.clk(gclk));
	jdff dff_B_u7wycnjS7_0(.din(w_dff_B_tsYHOX1q3_0),.dout(w_dff_B_u7wycnjS7_0),.clk(gclk));
	jdff dff_B_rwp3hnEd4_0(.din(w_dff_B_u7wycnjS7_0),.dout(w_dff_B_rwp3hnEd4_0),.clk(gclk));
	jdff dff_B_GKklkikf7_0(.din(w_dff_B_rwp3hnEd4_0),.dout(w_dff_B_GKklkikf7_0),.clk(gclk));
	jdff dff_B_V3T70aNx7_0(.din(w_dff_B_GKklkikf7_0),.dout(w_dff_B_V3T70aNx7_0),.clk(gclk));
	jdff dff_B_Ujlr2ZEg2_0(.din(w_dff_B_V3T70aNx7_0),.dout(w_dff_B_Ujlr2ZEg2_0),.clk(gclk));
	jdff dff_B_fzpbSU6a7_0(.din(w_dff_B_Ujlr2ZEg2_0),.dout(w_dff_B_fzpbSU6a7_0),.clk(gclk));
	jdff dff_B_rK25yWXp3_0(.din(w_dff_B_fzpbSU6a7_0),.dout(w_dff_B_rK25yWXp3_0),.clk(gclk));
	jdff dff_B_wBy5jWGb1_0(.din(w_dff_B_rK25yWXp3_0),.dout(w_dff_B_wBy5jWGb1_0),.clk(gclk));
	jdff dff_B_VmD68pLY4_0(.din(w_dff_B_wBy5jWGb1_0),.dout(w_dff_B_VmD68pLY4_0),.clk(gclk));
	jdff dff_B_0pIk17TD5_0(.din(w_dff_B_VmD68pLY4_0),.dout(w_dff_B_0pIk17TD5_0),.clk(gclk));
	jdff dff_A_hJW82m2V4_0(.dout(w_n364_0[0]),.din(w_dff_A_hJW82m2V4_0),.clk(gclk));
	jdff dff_A_qcHMD30S9_0(.dout(w_dff_A_hJW82m2V4_0),.din(w_dff_A_qcHMD30S9_0),.clk(gclk));
	jdff dff_A_N7O9EOkX8_0(.dout(w_dff_A_qcHMD30S9_0),.din(w_dff_A_N7O9EOkX8_0),.clk(gclk));
	jdff dff_A_j6zj1VIC0_0(.dout(w_dff_A_N7O9EOkX8_0),.din(w_dff_A_j6zj1VIC0_0),.clk(gclk));
	jdff dff_A_nhDcfOLW9_0(.dout(w_dff_A_j6zj1VIC0_0),.din(w_dff_A_nhDcfOLW9_0),.clk(gclk));
	jdff dff_A_Ckdu4Zry7_0(.dout(w_dff_A_nhDcfOLW9_0),.din(w_dff_A_Ckdu4Zry7_0),.clk(gclk));
	jdff dff_A_PLKzdo2s9_0(.dout(w_dff_A_Ckdu4Zry7_0),.din(w_dff_A_PLKzdo2s9_0),.clk(gclk));
	jdff dff_A_25FElTfP6_0(.dout(w_dff_A_PLKzdo2s9_0),.din(w_dff_A_25FElTfP6_0),.clk(gclk));
	jdff dff_A_tnZHCPXS6_0(.dout(w_dff_A_25FElTfP6_0),.din(w_dff_A_tnZHCPXS6_0),.clk(gclk));
	jdff dff_A_9I41b1se1_0(.dout(w_dff_A_tnZHCPXS6_0),.din(w_dff_A_9I41b1se1_0),.clk(gclk));
	jdff dff_A_4Ete7m1f1_0(.dout(w_dff_A_9I41b1se1_0),.din(w_dff_A_4Ete7m1f1_0),.clk(gclk));
	jdff dff_A_528SSXMD5_0(.dout(w_dff_A_4Ete7m1f1_0),.din(w_dff_A_528SSXMD5_0),.clk(gclk));
	jdff dff_A_2rWGtBLo2_0(.dout(w_dff_A_528SSXMD5_0),.din(w_dff_A_2rWGtBLo2_0),.clk(gclk));
	jdff dff_A_5o1TCmD08_0(.dout(w_dff_A_2rWGtBLo2_0),.din(w_dff_A_5o1TCmD08_0),.clk(gclk));
	jdff dff_A_CcABDC6X3_0(.dout(w_dff_A_5o1TCmD08_0),.din(w_dff_A_CcABDC6X3_0),.clk(gclk));
	jdff dff_B_hhH2xC3T0_1(.din(n374),.dout(w_dff_B_hhH2xC3T0_1),.clk(gclk));
	jdff dff_B_c0dvw7ia2_0(.din(n375),.dout(w_dff_B_c0dvw7ia2_0),.clk(gclk));
	jdff dff_B_DoWwuulz7_0(.din(w_dff_B_c0dvw7ia2_0),.dout(w_dff_B_DoWwuulz7_0),.clk(gclk));
	jdff dff_B_8o2Hng001_0(.din(w_dff_B_DoWwuulz7_0),.dout(w_dff_B_8o2Hng001_0),.clk(gclk));
	jdff dff_B_zfNmRqNX3_0(.din(w_dff_B_8o2Hng001_0),.dout(w_dff_B_zfNmRqNX3_0),.clk(gclk));
	jdff dff_B_boihjMx19_0(.din(w_dff_B_zfNmRqNX3_0),.dout(w_dff_B_boihjMx19_0),.clk(gclk));
	jdff dff_B_c1jH6Jpe8_0(.din(w_dff_B_boihjMx19_0),.dout(w_dff_B_c1jH6Jpe8_0),.clk(gclk));
	jdff dff_B_nhcB0gVo4_0(.din(w_dff_B_c1jH6Jpe8_0),.dout(w_dff_B_nhcB0gVo4_0),.clk(gclk));
	jdff dff_B_8taZhUz01_0(.din(w_dff_B_nhcB0gVo4_0),.dout(w_dff_B_8taZhUz01_0),.clk(gclk));
	jdff dff_B_PoYWSBeP3_0(.din(w_dff_B_8taZhUz01_0),.dout(w_dff_B_PoYWSBeP3_0),.clk(gclk));
	jdff dff_B_rpsa5okZ2_0(.din(w_dff_B_PoYWSBeP3_0),.dout(w_dff_B_rpsa5okZ2_0),.clk(gclk));
	jdff dff_B_v1dQ2yPZ9_0(.din(w_dff_B_rpsa5okZ2_0),.dout(w_dff_B_v1dQ2yPZ9_0),.clk(gclk));
	jdff dff_B_NEupvcRc5_0(.din(w_dff_B_v1dQ2yPZ9_0),.dout(w_dff_B_NEupvcRc5_0),.clk(gclk));
	jdff dff_B_LsTfgIb25_0(.din(w_dff_B_NEupvcRc5_0),.dout(w_dff_B_LsTfgIb25_0),.clk(gclk));
	jdff dff_B_6ZN0m6354_0(.din(w_dff_B_LsTfgIb25_0),.dout(w_dff_B_6ZN0m6354_0),.clk(gclk));
	jdff dff_A_mBkQ8FAy0_1(.dout(w_n372_0[1]),.din(w_dff_A_mBkQ8FAy0_1),.clk(gclk));
	jdff dff_A_YN62kmNa5_1(.dout(w_dff_A_mBkQ8FAy0_1),.din(w_dff_A_YN62kmNa5_1),.clk(gclk));
	jdff dff_A_aNi0VYs67_1(.dout(w_dff_A_YN62kmNa5_1),.din(w_dff_A_aNi0VYs67_1),.clk(gclk));
	jdff dff_A_f5GXX9C38_1(.dout(w_dff_A_aNi0VYs67_1),.din(w_dff_A_f5GXX9C38_1),.clk(gclk));
	jdff dff_A_DD2Q51WV7_1(.dout(w_dff_A_f5GXX9C38_1),.din(w_dff_A_DD2Q51WV7_1),.clk(gclk));
	jdff dff_A_76QmUyYJ1_1(.dout(w_dff_A_DD2Q51WV7_1),.din(w_dff_A_76QmUyYJ1_1),.clk(gclk));
	jdff dff_A_hXQ8m05g6_1(.dout(w_dff_A_76QmUyYJ1_1),.din(w_dff_A_hXQ8m05g6_1),.clk(gclk));
	jdff dff_A_zYPqyOQZ3_1(.dout(w_dff_A_hXQ8m05g6_1),.din(w_dff_A_zYPqyOQZ3_1),.clk(gclk));
	jdff dff_A_iKRB8Wsv9_1(.dout(w_dff_A_zYPqyOQZ3_1),.din(w_dff_A_iKRB8Wsv9_1),.clk(gclk));
	jdff dff_A_MT0lSSNP4_1(.dout(w_dff_A_iKRB8Wsv9_1),.din(w_dff_A_MT0lSSNP4_1),.clk(gclk));
	jdff dff_A_MfaGeG4A4_1(.dout(w_dff_A_MT0lSSNP4_1),.din(w_dff_A_MfaGeG4A4_1),.clk(gclk));
	jdff dff_A_s8bj5XiD9_1(.dout(w_dff_A_MfaGeG4A4_1),.din(w_dff_A_s8bj5XiD9_1),.clk(gclk));
	jdff dff_A_7sHtpric0_1(.dout(w_dff_A_s8bj5XiD9_1),.din(w_dff_A_7sHtpric0_1),.clk(gclk));
	jdff dff_A_XhwenyFf1_1(.dout(w_dff_A_7sHtpric0_1),.din(w_dff_A_XhwenyFf1_1),.clk(gclk));
	jdff dff_A_6mnfjbqs5_1(.dout(w_dff_A_XhwenyFf1_1),.din(w_dff_A_6mnfjbqs5_1),.clk(gclk));
	jdff dff_B_6Mcs3N3a4_1(.din(n380),.dout(w_dff_B_6Mcs3N3a4_1),.clk(gclk));
	jdff dff_B_IquWU2O29_1(.din(w_dff_B_6Mcs3N3a4_1),.dout(w_dff_B_IquWU2O29_1),.clk(gclk));
	jdff dff_B_TyHydjQp0_1(.din(w_dff_B_IquWU2O29_1),.dout(w_dff_B_TyHydjQp0_1),.clk(gclk));
	jdff dff_B_mD54nwjh4_1(.din(w_dff_B_TyHydjQp0_1),.dout(w_dff_B_mD54nwjh4_1),.clk(gclk));
	jdff dff_B_z8h3506y6_1(.din(w_dff_B_mD54nwjh4_1),.dout(w_dff_B_z8h3506y6_1),.clk(gclk));
	jdff dff_B_2GaigCDV5_1(.din(w_dff_B_z8h3506y6_1),.dout(w_dff_B_2GaigCDV5_1),.clk(gclk));
	jdff dff_B_lQkRj6Iz3_1(.din(w_dff_B_2GaigCDV5_1),.dout(w_dff_B_lQkRj6Iz3_1),.clk(gclk));
	jdff dff_B_LudLZ19a0_1(.din(w_dff_B_lQkRj6Iz3_1),.dout(w_dff_B_LudLZ19a0_1),.clk(gclk));
	jdff dff_B_VsWPvjX49_1(.din(w_dff_B_LudLZ19a0_1),.dout(w_dff_B_VsWPvjX49_1),.clk(gclk));
	jdff dff_B_qbYWJHA10_1(.din(w_dff_B_VsWPvjX49_1),.dout(w_dff_B_qbYWJHA10_1),.clk(gclk));
	jdff dff_B_O9sw4Yu05_1(.din(w_dff_B_qbYWJHA10_1),.dout(w_dff_B_O9sw4Yu05_1),.clk(gclk));
	jdff dff_B_sSDWAtkI3_1(.din(w_dff_B_O9sw4Yu05_1),.dout(w_dff_B_sSDWAtkI3_1),.clk(gclk));
	jdff dff_B_Le9lD93B3_1(.din(w_dff_B_sSDWAtkI3_1),.dout(w_dff_B_Le9lD93B3_1),.clk(gclk));
	jdff dff_B_GnHCDVG52_1(.din(w_dff_B_Le9lD93B3_1),.dout(w_dff_B_GnHCDVG52_1),.clk(gclk));
	jdff dff_B_PUcHH9zB0_1(.din(w_dff_B_GnHCDVG52_1),.dout(w_dff_B_PUcHH9zB0_1),.clk(gclk));
	jdff dff_B_H800PHkW1_0(.din(n382),.dout(w_dff_B_H800PHkW1_0),.clk(gclk));
	jdff dff_B_XO80HZbQ7_0(.din(w_dff_B_H800PHkW1_0),.dout(w_dff_B_XO80HZbQ7_0),.clk(gclk));
	jdff dff_B_HyClYrg89_0(.din(w_dff_B_XO80HZbQ7_0),.dout(w_dff_B_HyClYrg89_0),.clk(gclk));
	jdff dff_B_PkibqWmq9_0(.din(w_dff_B_HyClYrg89_0),.dout(w_dff_B_PkibqWmq9_0),.clk(gclk));
	jdff dff_B_Hqj4vDCg5_0(.din(w_dff_B_PkibqWmq9_0),.dout(w_dff_B_Hqj4vDCg5_0),.clk(gclk));
	jdff dff_B_Hgqy3dFk0_0(.din(w_dff_B_Hqj4vDCg5_0),.dout(w_dff_B_Hgqy3dFk0_0),.clk(gclk));
	jdff dff_B_v8gxKJNi0_0(.din(w_dff_B_Hgqy3dFk0_0),.dout(w_dff_B_v8gxKJNi0_0),.clk(gclk));
	jdff dff_B_1tux3dAl5_0(.din(w_dff_B_v8gxKJNi0_0),.dout(w_dff_B_1tux3dAl5_0),.clk(gclk));
	jdff dff_B_z6c6gTAI4_0(.din(w_dff_B_1tux3dAl5_0),.dout(w_dff_B_z6c6gTAI4_0),.clk(gclk));
	jdff dff_B_9P16P36S9_0(.din(w_dff_B_z6c6gTAI4_0),.dout(w_dff_B_9P16P36S9_0),.clk(gclk));
	jdff dff_B_kzZdAeqh0_0(.din(w_dff_B_9P16P36S9_0),.dout(w_dff_B_kzZdAeqh0_0),.clk(gclk));
	jdff dff_B_nEajhgS89_0(.din(w_dff_B_kzZdAeqh0_0),.dout(w_dff_B_nEajhgS89_0),.clk(gclk));
	jdff dff_B_vUCbUvtk0_0(.din(w_dff_B_nEajhgS89_0),.dout(w_dff_B_vUCbUvtk0_0),.clk(gclk));
	jdff dff_B_vItphulR1_0(.din(w_dff_B_vUCbUvtk0_0),.dout(w_dff_B_vItphulR1_0),.clk(gclk));
	jdff dff_B_HCeY6Xsg9_0(.din(n392),.dout(w_dff_B_HCeY6Xsg9_0),.clk(gclk));
	jdff dff_B_wMfhvqXj8_0(.din(w_dff_B_HCeY6Xsg9_0),.dout(w_dff_B_wMfhvqXj8_0),.clk(gclk));
	jdff dff_B_V7RppE9K3_0(.din(w_dff_B_wMfhvqXj8_0),.dout(w_dff_B_V7RppE9K3_0),.clk(gclk));
	jdff dff_B_hNunlZQT5_0(.din(w_dff_B_V7RppE9K3_0),.dout(w_dff_B_hNunlZQT5_0),.clk(gclk));
	jdff dff_B_FabcnBuR2_0(.din(w_dff_B_hNunlZQT5_0),.dout(w_dff_B_FabcnBuR2_0),.clk(gclk));
	jdff dff_B_EEEa5WqG6_0(.din(w_dff_B_FabcnBuR2_0),.dout(w_dff_B_EEEa5WqG6_0),.clk(gclk));
	jdff dff_B_CBw6WWyj2_0(.din(w_dff_B_EEEa5WqG6_0),.dout(w_dff_B_CBw6WWyj2_0),.clk(gclk));
	jdff dff_B_vE20W2EV6_0(.din(w_dff_B_CBw6WWyj2_0),.dout(w_dff_B_vE20W2EV6_0),.clk(gclk));
	jdff dff_B_wJ4gMpo62_0(.din(w_dff_B_vE20W2EV6_0),.dout(w_dff_B_wJ4gMpo62_0),.clk(gclk));
	jdff dff_B_21naDq6z9_0(.din(w_dff_B_wJ4gMpo62_0),.dout(w_dff_B_21naDq6z9_0),.clk(gclk));
	jdff dff_B_03H9PegJ1_0(.din(w_dff_B_21naDq6z9_0),.dout(w_dff_B_03H9PegJ1_0),.clk(gclk));
	jdff dff_B_utAAeGFS6_1(.din(n390),.dout(w_dff_B_utAAeGFS6_1),.clk(gclk));
	jdff dff_B_vd9YvGa17_1(.din(w_dff_B_utAAeGFS6_1),.dout(w_dff_B_vd9YvGa17_1),.clk(gclk));
	jdff dff_B_ooi95S6u9_0(.din(n388),.dout(w_dff_B_ooi95S6u9_0),.clk(gclk));
	jdff dff_B_i5PDVMKi8_0(.din(w_dff_B_ooi95S6u9_0),.dout(w_dff_B_i5PDVMKi8_0),.clk(gclk));
	jdff dff_B_FMRsiVLd6_0(.din(w_dff_B_i5PDVMKi8_0),.dout(w_dff_B_FMRsiVLd6_0),.clk(gclk));
	jdff dff_B_6EiM8kwb2_0(.din(w_dff_B_FMRsiVLd6_0),.dout(w_dff_B_6EiM8kwb2_0),.clk(gclk));
	jdff dff_B_cyxcypYz0_0(.din(w_dff_B_6EiM8kwb2_0),.dout(w_dff_B_cyxcypYz0_0),.clk(gclk));
	jdff dff_B_N3mjGSh68_0(.din(w_dff_B_cyxcypYz0_0),.dout(w_dff_B_N3mjGSh68_0),.clk(gclk));
	jdff dff_B_CTe91qRz2_0(.din(w_dff_B_N3mjGSh68_0),.dout(w_dff_B_CTe91qRz2_0),.clk(gclk));
	jdff dff_B_IgAnoSEi5_0(.din(w_dff_B_CTe91qRz2_0),.dout(w_dff_B_IgAnoSEi5_0),.clk(gclk));
	jdff dff_B_w8VI9R5M8_0(.din(w_dff_B_IgAnoSEi5_0),.dout(w_dff_B_w8VI9R5M8_0),.clk(gclk));
	jdff dff_B_fdQnRn6U8_0(.din(w_dff_B_w8VI9R5M8_0),.dout(w_dff_B_fdQnRn6U8_0),.clk(gclk));
	jdff dff_B_KCOZqQJA1_0(.din(w_dff_B_fdQnRn6U8_0),.dout(w_dff_B_KCOZqQJA1_0),.clk(gclk));
	jdff dff_B_6twX056v2_0(.din(w_dff_B_KCOZqQJA1_0),.dout(w_dff_B_6twX056v2_0),.clk(gclk));
	jdff dff_B_oKxb8BLI3_0(.din(w_dff_B_6twX056v2_0),.dout(w_dff_B_oKxb8BLI3_0),.clk(gclk));
	jdff dff_B_bNBiZI2c2_1(.din(n398),.dout(w_dff_B_bNBiZI2c2_1),.clk(gclk));
	jdff dff_B_0kZ2z18R8_0(.din(n224),.dout(w_dff_B_0kZ2z18R8_0),.clk(gclk));
	jdff dff_A_A0xHajm72_0(.dout(w_n218_1[0]),.din(w_dff_A_A0xHajm72_0),.clk(gclk));
	jdff dff_A_2Qa4mDst8_0(.dout(w_n218_0[0]),.din(w_dff_A_2Qa4mDst8_0),.clk(gclk));
	jdff dff_A_qkEZTYbq6_2(.dout(w_n218_0[2]),.din(w_dff_A_qkEZTYbq6_2),.clk(gclk));
	jdff dff_A_Q9G6vVgF3_2(.dout(w_dff_A_qkEZTYbq6_2),.din(w_dff_A_Q9G6vVgF3_2),.clk(gclk));
	jdff dff_A_jsAhbsnF8_0(.dout(w_n192_0[0]),.din(w_dff_A_jsAhbsnF8_0),.clk(gclk));
	jdff dff_A_AqRVZuO56_2(.dout(w_n192_0[2]),.din(w_dff_A_AqRVZuO56_2),.clk(gclk));
	jdff dff_B_xAj10c8M8_3(.din(n192),.dout(w_dff_B_xAj10c8M8_3),.clk(gclk));
	jdff dff_B_VWqHtd9m4_0(.din(n209),.dout(w_dff_B_VWqHtd9m4_0),.clk(gclk));
	jdff dff_A_l0EIxeY21_0(.dout(w_n198_0[0]),.din(w_dff_A_l0EIxeY21_0),.clk(gclk));
	jdff dff_A_KXlByAQf7_2(.dout(w_n198_0[2]),.din(w_dff_A_KXlByAQf7_2),.clk(gclk));
	jdff dff_A_jQgXWgqB0_2(.dout(w_dff_A_KXlByAQf7_2),.din(w_dff_A_jQgXWgqB0_2),.clk(gclk));
	jdff dff_A_2MC35eKk5_0(.dout(w_n197_1[0]),.din(w_dff_A_2MC35eKk5_0),.clk(gclk));
	jdff dff_A_bIOKmwFE6_0(.dout(w_dff_A_2MC35eKk5_0),.din(w_dff_A_bIOKmwFE6_0),.clk(gclk));
	jdff dff_A_7hU9kEf18_1(.dout(w_n197_0[1]),.din(w_dff_A_7hU9kEf18_1),.clk(gclk));
	jdff dff_A_HHgnVmET5_1(.dout(w_dff_A_7hU9kEf18_1),.din(w_dff_A_HHgnVmET5_1),.clk(gclk));
	jdff dff_A_L8M4JS3W9_0(.dout(w_n155_0[0]),.din(w_dff_A_L8M4JS3W9_0),.clk(gclk));
	jdff dff_A_e0hOEbT09_2(.dout(w_n155_0[2]),.din(w_dff_A_e0hOEbT09_2),.clk(gclk));
	jdff dff_B_XXYDJJC69_3(.din(n155),.dout(w_dff_B_XXYDJJC69_3),.clk(gclk));
	jdff dff_A_uOwPDkx45_0(.dout(w_n144_1[0]),.din(w_dff_A_uOwPDkx45_0),.clk(gclk));
	jdff dff_A_ALtmhgTc6_0(.dout(w_dff_A_uOwPDkx45_0),.din(w_dff_A_ALtmhgTc6_0),.clk(gclk));
	jdff dff_A_8RuVw5tC8_1(.dout(w_n144_0[1]),.din(w_dff_A_8RuVw5tC8_1),.clk(gclk));
	jdff dff_A_EGYRcwBO5_1(.dout(w_dff_A_8RuVw5tC8_1),.din(w_dff_A_EGYRcwBO5_1),.clk(gclk));
	jdff dff_A_9SSMtdeU1_2(.dout(w_n159_0[2]),.din(w_dff_A_9SSMtdeU1_2),.clk(gclk));
	jdff dff_A_gtbJ1B1o4_2(.dout(w_dff_A_9SSMtdeU1_2),.din(w_dff_A_gtbJ1B1o4_2),.clk(gclk));
	jdff dff_A_fOwRUP1N3_2(.dout(w_n121_0[2]),.din(w_dff_A_fOwRUP1N3_2),.clk(gclk));
	jdff dff_B_W1OUvgBT0_3(.din(n121),.dout(w_dff_B_W1OUvgBT0_3),.clk(gclk));
	jdff dff_A_Shzbzd048_1(.dout(w_n96_0[1]),.din(w_dff_A_Shzbzd048_1),.clk(gclk));
	jdff dff_A_W6SoiKOo9_1(.dout(w_dff_A_Shzbzd048_1),.din(w_dff_A_W6SoiKOo9_1),.clk(gclk));
	jdff dff_A_VFOZdRBQ2_1(.dout(w_dff_A_W6SoiKOo9_1),.din(w_dff_A_VFOZdRBQ2_1),.clk(gclk));
	jdff dff_A_FvrCfnJD3_1(.dout(w_dff_A_VFOZdRBQ2_1),.din(w_dff_A_FvrCfnJD3_1),.clk(gclk));
	jdff dff_A_I348fSb59_2(.dout(w_n96_0[2]),.din(w_dff_A_I348fSb59_2),.clk(gclk));
	jdff dff_A_Mogc7lRq2_2(.dout(w_dff_A_I348fSb59_2),.din(w_dff_A_Mogc7lRq2_2),.clk(gclk));
	jdff dff_A_y4d6FUuI4_2(.dout(w_dff_A_Mogc7lRq2_2),.din(w_dff_A_y4d6FUuI4_2),.clk(gclk));
	jdff dff_A_hDLlR9aU9_2(.dout(w_dff_A_y4d6FUuI4_2),.din(w_dff_A_hDLlR9aU9_2),.clk(gclk));
	jdff dff_B_fmX5IGTT2_3(.din(n340),.dout(w_dff_B_fmX5IGTT2_3),.clk(gclk));
	jdff dff_B_VihuQQtv3_3(.din(w_dff_B_fmX5IGTT2_3),.dout(w_dff_B_VihuQQtv3_3),.clk(gclk));
	jdff dff_B_iqoVMd6k3_3(.din(w_dff_B_VihuQQtv3_3),.dout(w_dff_B_iqoVMd6k3_3),.clk(gclk));
	jdff dff_B_ylKjk9M09_3(.din(w_dff_B_iqoVMd6k3_3),.dout(w_dff_B_ylKjk9M09_3),.clk(gclk));
	jdff dff_B_ugbwOPxA9_3(.din(w_dff_B_ylKjk9M09_3),.dout(w_dff_B_ugbwOPxA9_3),.clk(gclk));
	jdff dff_B_91GUwpgB9_3(.din(w_dff_B_ugbwOPxA9_3),.dout(w_dff_B_91GUwpgB9_3),.clk(gclk));
	jdff dff_B_PtF5RnJI4_3(.din(w_dff_B_91GUwpgB9_3),.dout(w_dff_B_PtF5RnJI4_3),.clk(gclk));
	jdff dff_B_ews6HzcO6_3(.din(w_dff_B_PtF5RnJI4_3),.dout(w_dff_B_ews6HzcO6_3),.clk(gclk));
	jdff dff_B_x22F5vcs9_3(.din(w_dff_B_ews6HzcO6_3),.dout(w_dff_B_x22F5vcs9_3),.clk(gclk));
	jdff dff_B_OwRWhq653_3(.din(w_dff_B_x22F5vcs9_3),.dout(w_dff_B_OwRWhq653_3),.clk(gclk));
	jdff dff_B_iRIJRMt13_3(.din(w_dff_B_OwRWhq653_3),.dout(w_dff_B_iRIJRMt13_3),.clk(gclk));
	jdff dff_B_8eHgVTOX8_3(.din(w_dff_B_iRIJRMt13_3),.dout(w_dff_B_8eHgVTOX8_3),.clk(gclk));
	jdff dff_B_aqMOPiYk9_3(.din(w_dff_B_8eHgVTOX8_3),.dout(w_dff_B_aqMOPiYk9_3),.clk(gclk));
	jdff dff_B_AiVg1xue0_3(.din(w_dff_B_aqMOPiYk9_3),.dout(w_dff_B_AiVg1xue0_3),.clk(gclk));
	jdff dff_B_LKvHw9nw2_3(.din(w_dff_B_AiVg1xue0_3),.dout(w_dff_B_LKvHw9nw2_3),.clk(gclk));
	jdff dff_B_XEK9xg8v1_3(.din(w_dff_B_LKvHw9nw2_3),.dout(w_dff_B_XEK9xg8v1_3),.clk(gclk));
	jdff dff_B_qrCXNbTi1_1(.din(n394),.dout(w_dff_B_qrCXNbTi1_1),.clk(gclk));
	jdff dff_B_kmet4QdL0_1(.din(w_dff_B_qrCXNbTi1_1),.dout(w_dff_B_kmet4QdL0_1),.clk(gclk));
	jdff dff_B_UIP3Bl9K0_1(.din(w_dff_B_kmet4QdL0_1),.dout(w_dff_B_UIP3Bl9K0_1),.clk(gclk));
	jdff dff_B_fC369nER5_1(.din(w_dff_B_UIP3Bl9K0_1),.dout(w_dff_B_fC369nER5_1),.clk(gclk));
	jdff dff_B_fFhIUMYH7_1(.din(w_dff_B_fC369nER5_1),.dout(w_dff_B_fFhIUMYH7_1),.clk(gclk));
	jdff dff_B_MSky3R4C5_1(.din(w_dff_B_fFhIUMYH7_1),.dout(w_dff_B_MSky3R4C5_1),.clk(gclk));
	jdff dff_B_8etoQi9d5_1(.din(w_dff_B_MSky3R4C5_1),.dout(w_dff_B_8etoQi9d5_1),.clk(gclk));
	jdff dff_B_Z35LIqLt5_1(.din(w_dff_B_8etoQi9d5_1),.dout(w_dff_B_Z35LIqLt5_1),.clk(gclk));
	jdff dff_B_CxMlmehe3_1(.din(w_dff_B_Z35LIqLt5_1),.dout(w_dff_B_CxMlmehe3_1),.clk(gclk));
	jdff dff_B_rM6vO3xV6_1(.din(w_dff_B_CxMlmehe3_1),.dout(w_dff_B_rM6vO3xV6_1),.clk(gclk));
	jdff dff_B_rg16n2yA1_1(.din(w_dff_B_rM6vO3xV6_1),.dout(w_dff_B_rg16n2yA1_1),.clk(gclk));
	jdff dff_B_dn0deQQx3_0(.din(n396),.dout(w_dff_B_dn0deQQx3_0),.clk(gclk));
	jdff dff_B_rHLRHm304_0(.din(w_dff_B_dn0deQQx3_0),.dout(w_dff_B_rHLRHm304_0),.clk(gclk));
	jdff dff_B_dBUl07bo3_0(.din(w_dff_B_rHLRHm304_0),.dout(w_dff_B_dBUl07bo3_0),.clk(gclk));
	jdff dff_B_nFgPMPZJ8_0(.din(w_dff_B_dBUl07bo3_0),.dout(w_dff_B_nFgPMPZJ8_0),.clk(gclk));
	jdff dff_B_e6POofZE0_0(.din(w_dff_B_nFgPMPZJ8_0),.dout(w_dff_B_e6POofZE0_0),.clk(gclk));
	jdff dff_B_k9as2cgn9_0(.din(w_dff_B_e6POofZE0_0),.dout(w_dff_B_k9as2cgn9_0),.clk(gclk));
	jdff dff_B_iJ1Sgwnx8_0(.din(w_dff_B_k9as2cgn9_0),.dout(w_dff_B_iJ1Sgwnx8_0),.clk(gclk));
	jdff dff_B_MHYNxXFv3_0(.din(w_dff_B_iJ1Sgwnx8_0),.dout(w_dff_B_MHYNxXFv3_0),.clk(gclk));
	jdff dff_B_xh2IlJkJ3_0(.din(w_dff_B_MHYNxXFv3_0),.dout(w_dff_B_xh2IlJkJ3_0),.clk(gclk));
	jdff dff_B_TpthdZRQ8_0(.din(w_dff_B_xh2IlJkJ3_0),.dout(w_dff_B_TpthdZRQ8_0),.clk(gclk));
	jdff dff_B_ZItEWuXN2_0(.din(w_dff_B_TpthdZRQ8_0),.dout(w_dff_B_ZItEWuXN2_0),.clk(gclk));
	jdff dff_B_VNNNKHBf2_0(.din(w_dff_B_ZItEWuXN2_0),.dout(w_dff_B_VNNNKHBf2_0),.clk(gclk));
	jdff dff_B_YYTIRybh0_0(.din(w_dff_B_VNNNKHBf2_0),.dout(w_dff_B_YYTIRybh0_0),.clk(gclk));
	jdff dff_B_dl0Rx4Pp3_0(.din(w_dff_B_YYTIRybh0_0),.dout(w_dff_B_dl0Rx4Pp3_0),.clk(gclk));
	jdff dff_A_1fyWL2jF4_0(.dout(w_n395_0[0]),.din(w_dff_A_1fyWL2jF4_0),.clk(gclk));
	jdff dff_A_73TrNSFc1_0(.dout(w_dff_A_1fyWL2jF4_0),.din(w_dff_A_73TrNSFc1_0),.clk(gclk));
	jdff dff_A_hmd0lHZm7_0(.dout(w_dff_A_73TrNSFc1_0),.din(w_dff_A_hmd0lHZm7_0),.clk(gclk));
	jdff dff_A_oxJmmROU8_0(.dout(w_dff_A_hmd0lHZm7_0),.din(w_dff_A_oxJmmROU8_0),.clk(gclk));
	jdff dff_A_T0lDex9y5_0(.dout(w_dff_A_oxJmmROU8_0),.din(w_dff_A_T0lDex9y5_0),.clk(gclk));
	jdff dff_A_F0V9QpbM3_0(.dout(w_dff_A_T0lDex9y5_0),.din(w_dff_A_F0V9QpbM3_0),.clk(gclk));
	jdff dff_A_UBbUylUN6_0(.dout(w_dff_A_F0V9QpbM3_0),.din(w_dff_A_UBbUylUN6_0),.clk(gclk));
	jdff dff_A_PVzqeHDp0_0(.dout(w_dff_A_UBbUylUN6_0),.din(w_dff_A_PVzqeHDp0_0),.clk(gclk));
	jdff dff_A_hGkt8E1k4_0(.dout(w_dff_A_PVzqeHDp0_0),.din(w_dff_A_hGkt8E1k4_0),.clk(gclk));
	jdff dff_A_mSLNJsGa4_0(.dout(w_dff_A_hGkt8E1k4_0),.din(w_dff_A_mSLNJsGa4_0),.clk(gclk));
	jdff dff_A_pMrlqy470_0(.dout(w_dff_A_mSLNJsGa4_0),.din(w_dff_A_pMrlqy470_0),.clk(gclk));
	jdff dff_A_m6Qx9DAJ2_0(.dout(w_dff_A_pMrlqy470_0),.din(w_dff_A_m6Qx9DAJ2_0),.clk(gclk));
	jdff dff_A_LhM1B9Pt1_0(.dout(w_dff_A_m6Qx9DAJ2_0),.din(w_dff_A_LhM1B9Pt1_0),.clk(gclk));
	jdff dff_A_fd4PZKEL4_0(.dout(w_dff_A_LhM1B9Pt1_0),.din(w_dff_A_fd4PZKEL4_0),.clk(gclk));
	jdff dff_A_U46uTslA6_0(.dout(w_dff_A_fd4PZKEL4_0),.din(w_dff_A_U46uTslA6_0),.clk(gclk));
	jdff dff_B_qRJjuky49_0(.din(n329),.dout(w_dff_B_qRJjuky49_0),.clk(gclk));
	jdff dff_B_P1oev6OL7_0(.din(n323),.dout(w_dff_B_P1oev6OL7_0),.clk(gclk));
	jdff dff_A_O4s2vHtd0_1(.dout(w_n189_0[1]),.din(w_dff_A_O4s2vHtd0_1),.clk(gclk));
	jdff dff_A_eRcrnQaJ8_1(.dout(w_dff_A_O4s2vHtd0_1),.din(w_dff_A_eRcrnQaJ8_1),.clk(gclk));
	jdff dff_B_0F73FT6u8_2(.din(n318),.dout(w_dff_B_0F73FT6u8_2),.clk(gclk));
	jdff dff_A_CtB0uMGN2_1(.dout(w_n185_0[1]),.din(w_dff_A_CtB0uMGN2_1),.clk(gclk));
	jdff dff_A_NtqSXtuH4_1(.dout(w_dff_A_CtB0uMGN2_1),.din(w_dff_A_NtqSXtuH4_1),.clk(gclk));
	jdff dff_A_hBG93Yhh6_2(.dout(w_n185_0[2]),.din(w_dff_A_hBG93Yhh6_2),.clk(gclk));
	jdff dff_A_7XvFw0v89_2(.dout(w_dff_A_hBG93Yhh6_2),.din(w_dff_A_7XvFw0v89_2),.clk(gclk));
	jdff dff_B_6TFqzJ3w3_3(.din(n184),.dout(w_dff_B_6TFqzJ3w3_3),.clk(gclk));
	jdff dff_B_IEPWR7JI3_3(.din(w_dff_B_6TFqzJ3w3_3),.dout(w_dff_B_IEPWR7JI3_3),.clk(gclk));
	jdff dff_A_DjGGIK7h6_0(.dout(w_n314_0[0]),.din(w_dff_A_DjGGIK7h6_0),.clk(gclk));
	jdff dff_A_FKtcFAdn1_1(.dout(w_n314_0[1]),.din(w_dff_A_FKtcFAdn1_1),.clk(gclk));
	jdff dff_B_IwweuLLc4_3(.din(n314),.dout(w_dff_B_IwweuLLc4_3),.clk(gclk));
	jdff dff_A_n1nyfuVj7_1(.dout(w_n311_0[1]),.din(w_dff_A_n1nyfuVj7_1),.clk(gclk));
	jdff dff_A_OZ8KK12W0_2(.dout(w_n311_0[2]),.din(w_dff_A_OZ8KK12W0_2),.clk(gclk));
	jdff dff_B_xgSN3V3V7_3(.din(n311),.dout(w_dff_B_xgSN3V3V7_3),.clk(gclk));
	jdff dff_A_pbPmsnQ15_0(.dout(w_n183_0[0]),.din(w_dff_A_pbPmsnQ15_0),.clk(gclk));
	jdff dff_A_aL9ZvaMz2_0(.dout(w_dff_A_pbPmsnQ15_0),.din(w_dff_A_aL9ZvaMz2_0),.clk(gclk));
	jdff dff_A_EWqnEigz3_0(.dout(w_dff_A_aL9ZvaMz2_0),.din(w_dff_A_EWqnEigz3_0),.clk(gclk));
	jdff dff_A_WrjgMOFJ0_1(.dout(w_n183_0[1]),.din(w_dff_A_WrjgMOFJ0_1),.clk(gclk));
	jdff dff_A_E73AQ5V10_1(.dout(w_dff_A_WrjgMOFJ0_1),.din(w_dff_A_E73AQ5V10_1),.clk(gclk));
	jdff dff_A_CpOdx5Gu0_1(.dout(w_dff_A_E73AQ5V10_1),.din(w_dff_A_CpOdx5Gu0_1),.clk(gclk));
	jdff dff_B_wOFWd6LP3_0(.din(n182),.dout(w_dff_B_wOFWd6LP3_0),.clk(gclk));
	jdff dff_B_GAw23NGM7_1(.din(G900),.dout(w_dff_B_GAw23NGM7_1),.clk(gclk));
	jdff dff_B_nCvU86gK5_0(.din(n304),.dout(w_dff_B_nCvU86gK5_0),.clk(gclk));
	jdff dff_A_REGWZ8k48_1(.dout(w_n188_0[1]),.din(w_dff_A_REGWZ8k48_1),.clk(gclk));
	jdff dff_A_n2Tcoh2U6_0(.dout(w_n290_0[0]),.din(w_dff_A_n2Tcoh2U6_0),.clk(gclk));
	jdff dff_B_vBdGNBbj5_3(.din(n290),.dout(w_dff_B_vBdGNBbj5_3),.clk(gclk));
	jdff dff_A_VrzoVLr50_0(.dout(w_n289_0[0]),.din(w_dff_A_VrzoVLr50_0),.clk(gclk));
	jdff dff_A_lnNYhLRA3_0(.dout(w_dff_A_VrzoVLr50_0),.din(w_dff_A_lnNYhLRA3_0),.clk(gclk));
	jdff dff_B_sJq7yOVI7_3(.din(n158),.dout(w_dff_B_sJq7yOVI7_3),.clk(gclk));
	jdff dff_A_IANGZgsD2_0(.dout(w_n92_1[0]),.din(w_dff_A_IANGZgsD2_0),.clk(gclk));
	jdff dff_A_OK5if8aX3_0(.dout(w_dff_A_IANGZgsD2_0),.din(w_dff_A_OK5if8aX3_0),.clk(gclk));
	jdff dff_A_tmxZjWrt0_2(.dout(w_n92_1[2]),.din(w_dff_A_tmxZjWrt0_2),.clk(gclk));
	jdff dff_A_XI8h2cgr0_2(.dout(w_dff_A_tmxZjWrt0_2),.din(w_dff_A_XI8h2cgr0_2),.clk(gclk));
	jdff dff_B_E2Ozntam6_2(.din(n286),.dout(w_dff_B_E2Ozntam6_2),.clk(gclk));
	jdff dff_A_X1itAvbh4_1(.dout(w_n163_0[1]),.din(w_dff_A_X1itAvbh4_1),.clk(gclk));
	jdff dff_A_L4GXIG7G1_1(.dout(w_dff_A_X1itAvbh4_1),.din(w_dff_A_L4GXIG7G1_1),.clk(gclk));
	jdff dff_A_T3WBiKFQ5_2(.dout(w_n163_0[2]),.din(w_dff_A_T3WBiKFQ5_2),.clk(gclk));
	jdff dff_A_19nn0ZKO9_2(.dout(w_dff_A_T3WBiKFQ5_2),.din(w_dff_A_19nn0ZKO9_2),.clk(gclk));
	jdff dff_B_RlcOllUj0_1(.din(n123),.dout(w_dff_B_RlcOllUj0_1),.clk(gclk));
	jdff dff_B_BttTsZuX8_1(.din(w_dff_B_RlcOllUj0_1),.dout(w_dff_B_BttTsZuX8_1),.clk(gclk));
	jdff dff_B_2NvLaf0d2_1(.din(w_dff_B_BttTsZuX8_1),.dout(w_dff_B_2NvLaf0d2_1),.clk(gclk));
	jdff dff_B_E6KpvIQS1_1(.din(w_dff_B_2NvLaf0d2_1),.dout(w_dff_B_E6KpvIQS1_1),.clk(gclk));
	jdff dff_B_tgqTKjST6_1(.din(w_dff_B_E6KpvIQS1_1),.dout(w_dff_B_tgqTKjST6_1),.clk(gclk));
	jdff dff_A_3uMTGr290_0(.dout(w_n68_0[0]),.din(w_dff_A_3uMTGr290_0),.clk(gclk));
	jdff dff_A_enOvBShm0_0(.dout(w_dff_A_3uMTGr290_0),.din(w_dff_A_enOvBShm0_0),.clk(gclk));
	jdff dff_A_ENUTJ48H9_0(.dout(w_dff_A_enOvBShm0_0),.din(w_dff_A_ENUTJ48H9_0),.clk(gclk));
	jdff dff_A_8LcSwH8V3_0(.dout(w_dff_A_ENUTJ48H9_0),.din(w_dff_A_8LcSwH8V3_0),.clk(gclk));
	jdff dff_A_1W7IgUaM5_0(.dout(w_dff_A_8LcSwH8V3_0),.din(w_dff_A_1W7IgUaM5_0),.clk(gclk));
	jdff dff_A_58imru5c5_0(.dout(w_dff_A_1W7IgUaM5_0),.din(w_dff_A_58imru5c5_0),.clk(gclk));
	jdff dff_A_TsBU1uMv0_0(.dout(w_dff_A_58imru5c5_0),.din(w_dff_A_TsBU1uMv0_0),.clk(gclk));
	jdff dff_A_sPGb23ld7_0(.dout(w_dff_A_TsBU1uMv0_0),.din(w_dff_A_sPGb23ld7_0),.clk(gclk));
	jdff dff_A_k3v7wEYI1_0(.dout(w_dff_A_sPGb23ld7_0),.din(w_dff_A_k3v7wEYI1_0),.clk(gclk));
	jdff dff_A_6AJDCdFE1_0(.dout(w_dff_A_k3v7wEYI1_0),.din(w_dff_A_6AJDCdFE1_0),.clk(gclk));
	jdff dff_A_XLhE6Odj0_0(.dout(w_n281_0[0]),.din(w_dff_A_XLhE6Odj0_0),.clk(gclk));
	jdff dff_A_sTQzwxcp3_1(.dout(w_n281_0[1]),.din(w_dff_A_sTQzwxcp3_1),.clk(gclk));
	jdff dff_B_RiIbFyzW2_3(.din(n281),.dout(w_dff_B_RiIbFyzW2_3),.clk(gclk));
	jdff dff_B_GQ5WKW4Z3_2(.din(n278),.dout(w_dff_B_GQ5WKW4Z3_2),.clk(gclk));
	jdff dff_A_LPKtXx3w1_1(.dout(w_n168_0[1]),.din(w_dff_A_LPKtXx3w1_1),.clk(gclk));
	jdff dff_A_375026EZ7_1(.dout(w_dff_A_LPKtXx3w1_1),.din(w_dff_A_375026EZ7_1),.clk(gclk));
	jdff dff_A_4M3NhlzX8_2(.dout(w_n168_0[2]),.din(w_dff_A_4M3NhlzX8_2),.clk(gclk));
	jdff dff_A_MM0cDStJ0_2(.dout(w_dff_A_4M3NhlzX8_2),.din(w_dff_A_MM0cDStJ0_2),.clk(gclk));
	jdff dff_B_RYP7aEv24_1(.din(n133),.dout(w_dff_B_RYP7aEv24_1),.clk(gclk));
	jdff dff_B_iB72dv0Z8_1(.din(w_dff_B_RYP7aEv24_1),.dout(w_dff_B_iB72dv0Z8_1),.clk(gclk));
	jdff dff_B_al3r44FB2_1(.din(w_dff_B_iB72dv0Z8_1),.dout(w_dff_B_al3r44FB2_1),.clk(gclk));
	jdff dff_B_A7iquh0X4_1(.din(w_dff_B_al3r44FB2_1),.dout(w_dff_B_A7iquh0X4_1),.clk(gclk));
	jdff dff_B_gkBWQhNm3_1(.din(w_dff_B_A7iquh0X4_1),.dout(w_dff_B_gkBWQhNm3_1),.clk(gclk));
	jdff dff_A_gg5hEwhF8_0(.dout(w_n141_0[0]),.din(w_dff_A_gg5hEwhF8_0),.clk(gclk));
	jdff dff_A_WenNg6Ky8_0(.dout(w_dff_A_gg5hEwhF8_0),.din(w_dff_A_WenNg6Ky8_0),.clk(gclk));
	jdff dff_A_MwJvXmnu9_0(.dout(w_dff_A_WenNg6Ky8_0),.din(w_dff_A_MwJvXmnu9_0),.clk(gclk));
	jdff dff_A_pDQ020eG4_0(.dout(w_dff_A_MwJvXmnu9_0),.din(w_dff_A_pDQ020eG4_0),.clk(gclk));
	jdff dff_A_Q68tyZJT3_0(.dout(w_dff_A_pDQ020eG4_0),.din(w_dff_A_Q68tyZJT3_0),.clk(gclk));
	jdff dff_A_LC3rQaQt4_0(.dout(w_dff_A_Q68tyZJT3_0),.din(w_dff_A_LC3rQaQt4_0),.clk(gclk));
	jdff dff_A_ZmC3SGWn1_0(.dout(w_dff_A_LC3rQaQt4_0),.din(w_dff_A_ZmC3SGWn1_0),.clk(gclk));
	jdff dff_A_Ljyw1Tfj2_0(.dout(w_dff_A_ZmC3SGWn1_0),.din(w_dff_A_Ljyw1Tfj2_0),.clk(gclk));
	jdff dff_A_0ya4Ojth2_0(.dout(w_dff_A_Ljyw1Tfj2_0),.din(w_dff_A_0ya4Ojth2_0),.clk(gclk));
	jdff dff_A_gRXzx6lV4_0(.dout(w_dff_A_0ya4Ojth2_0),.din(w_dff_A_gRXzx6lV4_0),.clk(gclk));
	jdff dff_A_ehwNMh3i9_0(.dout(w_dff_A_gRXzx6lV4_0),.din(w_dff_A_ehwNMh3i9_0),.clk(gclk));
	jdff dff_A_gV3TYRGf2_0(.dout(w_dff_A_ehwNMh3i9_0),.din(w_dff_A_gV3TYRGf2_0),.clk(gclk));
	jdff dff_B_wGKmiluw8_1(.din(n134),.dout(w_dff_B_wGKmiluw8_1),.clk(gclk));
	jdff dff_B_32cs7bWc2_1(.din(w_dff_B_wGKmiluw8_1),.dout(w_dff_B_32cs7bWc2_1),.clk(gclk));
	jdff dff_A_iMghNJmt4_1(.dout(w_G475_0[1]),.din(w_dff_A_iMghNJmt4_1),.clk(gclk));
	jdff dff_A_r5EtnzcC9_1(.dout(w_dff_A_iMghNJmt4_1),.din(w_dff_A_r5EtnzcC9_1),.clk(gclk));
	jdff dff_A_hAaYs4WB6_1(.dout(w_dff_A_r5EtnzcC9_1),.din(w_dff_A_hAaYs4WB6_1),.clk(gclk));
	jdff dff_A_Teu1UDtW7_1(.dout(w_dff_A_hAaYs4WB6_1),.din(w_dff_A_Teu1UDtW7_1),.clk(gclk));
	jdff dff_A_Yd45RafL0_1(.dout(w_dff_A_Teu1UDtW7_1),.din(w_dff_A_Yd45RafL0_1),.clk(gclk));
	jdff dff_A_CEab87fn1_1(.dout(w_dff_A_Yd45RafL0_1),.din(w_dff_A_CEab87fn1_1),.clk(gclk));
	jdff dff_A_PEcKYvTo2_0(.dout(w_n130_0[0]),.din(w_dff_A_PEcKYvTo2_0),.clk(gclk));
	jdff dff_A_09Ithtd01_0(.dout(w_dff_A_PEcKYvTo2_0),.din(w_dff_A_09Ithtd01_0),.clk(gclk));
	jdff dff_A_0AGzoZu19_0(.dout(w_dff_A_09Ithtd01_0),.din(w_dff_A_0AGzoZu19_0),.clk(gclk));
	jdff dff_A_YDij4JRz9_0(.dout(w_dff_A_0AGzoZu19_0),.din(w_dff_A_YDij4JRz9_0),.clk(gclk));
	jdff dff_A_NYwfiaWO3_0(.dout(w_dff_A_YDij4JRz9_0),.din(w_dff_A_NYwfiaWO3_0),.clk(gclk));
	jdff dff_A_XnX1efKo4_0(.dout(w_dff_A_NYwfiaWO3_0),.din(w_dff_A_XnX1efKo4_0),.clk(gclk));
	jdff dff_A_PYpkFaEB2_0(.dout(w_dff_A_XnX1efKo4_0),.din(w_dff_A_PYpkFaEB2_0),.clk(gclk));
	jdff dff_A_FIvoixvh8_0(.dout(w_dff_A_PYpkFaEB2_0),.din(w_dff_A_FIvoixvh8_0),.clk(gclk));
	jdff dff_A_ULOqf1aM8_0(.dout(w_dff_A_FIvoixvh8_0),.din(w_dff_A_ULOqf1aM8_0),.clk(gclk));
	jdff dff_A_HFst59VX1_0(.dout(w_dff_A_ULOqf1aM8_0),.din(w_dff_A_HFst59VX1_0),.clk(gclk));
	jdff dff_A_VSiWk4ZR0_0(.dout(w_dff_A_HFst59VX1_0),.din(w_dff_A_VSiWk4ZR0_0),.clk(gclk));
	jdff dff_A_BIDb6lWi9_0(.dout(w_dff_A_VSiWk4ZR0_0),.din(w_dff_A_BIDb6lWi9_0),.clk(gclk));
	jdff dff_B_Po8Zbi7a6_1(.din(n124),.dout(w_dff_B_Po8Zbi7a6_1),.clk(gclk));
	jdff dff_B_Q3GIcbza0_1(.din(w_dff_B_Po8Zbi7a6_1),.dout(w_dff_B_Q3GIcbza0_1),.clk(gclk));
	jdff dff_B_KYf5x2SV2_1(.din(w_dff_B_Q3GIcbza0_1),.dout(w_dff_B_KYf5x2SV2_1),.clk(gclk));
	jdff dff_B_vWcuUjsK6_0(.din(n128),.dout(w_dff_B_vWcuUjsK6_0),.clk(gclk));
	jdff dff_A_uWZcgsMi2_1(.dout(w_G478_0[1]),.din(w_dff_A_uWZcgsMi2_1),.clk(gclk));
	jdff dff_A_ScB36H0X3_1(.dout(w_dff_A_uWZcgsMi2_1),.din(w_dff_A_ScB36H0X3_1),.clk(gclk));
	jdff dff_A_4c38AGAK5_1(.dout(w_dff_A_ScB36H0X3_1),.din(w_dff_A_4c38AGAK5_1),.clk(gclk));
	jdff dff_A_azIz4Y8S7_1(.dout(w_dff_A_4c38AGAK5_1),.din(w_dff_A_azIz4Y8S7_1),.clk(gclk));
	jdff dff_A_xzz8La4D7_1(.dout(w_dff_A_azIz4Y8S7_1),.din(w_dff_A_xzz8La4D7_1),.clk(gclk));
	jdff dff_A_WWtRK1vQ1_1(.dout(w_dff_A_xzz8La4D7_1),.din(w_dff_A_WWtRK1vQ1_1),.clk(gclk));
	jdff dff_B_Ecqpcddf1_3(.din(n154),.dout(w_dff_B_Ecqpcddf1_3),.clk(gclk));
	jdff dff_B_3tMQlBob3_3(.din(w_dff_B_Ecqpcddf1_3),.dout(w_dff_B_3tMQlBob3_3),.clk(gclk));
	jdff dff_A_tw9iMYm32_0(.dout(w_n153_0[0]),.din(w_dff_A_tw9iMYm32_0),.clk(gclk));
	jdff dff_A_7f6FhRxn3_0(.dout(w_dff_A_tw9iMYm32_0),.din(w_dff_A_7f6FhRxn3_0),.clk(gclk));
	jdff dff_A_qAr5oImy2_0(.dout(w_dff_A_7f6FhRxn3_0),.din(w_dff_A_qAr5oImy2_0),.clk(gclk));
	jdff dff_A_y39Ir1fy5_1(.dout(w_n153_0[1]),.din(w_dff_A_y39Ir1fy5_1),.clk(gclk));
	jdff dff_A_ZNGFzyY63_1(.dout(w_dff_A_y39Ir1fy5_1),.din(w_dff_A_ZNGFzyY63_1),.clk(gclk));
	jdff dff_A_SAYeAZFS1_1(.dout(w_dff_A_ZNGFzyY63_1),.din(w_dff_A_SAYeAZFS1_1),.clk(gclk));
	jdff dff_B_jF5kPCUT9_1(.din(n148),.dout(w_dff_B_jF5kPCUT9_1),.clk(gclk));
	jdff dff_A_AizOC6QN4_0(.dout(w_n151_0[0]),.din(w_dff_A_AizOC6QN4_0),.clk(gclk));
	jdff dff_A_IZaReYdH1_1(.dout(w_n151_0[1]),.din(w_dff_A_IZaReYdH1_1),.clk(gclk));
	jdff dff_A_GEijYecu8_1(.dout(w_dff_A_IZaReYdH1_1),.din(w_dff_A_GEijYecu8_1),.clk(gclk));
	jdff dff_A_5Qhka2Bg4_1(.dout(w_dff_A_GEijYecu8_1),.din(w_dff_A_5Qhka2Bg4_1),.clk(gclk));
	jdff dff_A_E7JR0M4V6_1(.dout(w_dff_A_5Qhka2Bg4_1),.din(w_dff_A_E7JR0M4V6_1),.clk(gclk));
	jdff dff_A_wSuxgyHR1_1(.dout(w_dff_A_E7JR0M4V6_1),.din(w_dff_A_wSuxgyHR1_1),.clk(gclk));
	jdff dff_A_edH96Hus4_1(.dout(w_dff_A_wSuxgyHR1_1),.din(w_dff_A_edH96Hus4_1),.clk(gclk));
	jdff dff_A_A1IDbqi44_1(.dout(w_dff_A_edH96Hus4_1),.din(w_dff_A_A1IDbqi44_1),.clk(gclk));
	jdff dff_A_SI7If7WT8_1(.dout(w_dff_A_A1IDbqi44_1),.din(w_dff_A_SI7If7WT8_1),.clk(gclk));
	jdff dff_A_m2SUxvgv9_1(.dout(w_dff_A_SI7If7WT8_1),.din(w_dff_A_m2SUxvgv9_1),.clk(gclk));
	jdff dff_A_Wp07xHDd0_1(.dout(w_dff_A_m2SUxvgv9_1),.din(w_dff_A_Wp07xHDd0_1),.clk(gclk));
	jdff dff_A_CJMSy18s4_1(.dout(w_dff_A_Wp07xHDd0_1),.din(w_dff_A_CJMSy18s4_1),.clk(gclk));
	jdff dff_A_E0bkq6j93_1(.dout(w_G952_0[1]),.din(w_dff_A_E0bkq6j93_1),.clk(gclk));
	jdff dff_A_o6mUYrvZ4_1(.dout(w_dff_A_E0bkq6j93_1),.din(w_dff_A_o6mUYrvZ4_1),.clk(gclk));
	jdff dff_A_6XTcObx51_1(.dout(w_dff_A_o6mUYrvZ4_1),.din(w_dff_A_6XTcObx51_1),.clk(gclk));
	jdff dff_A_nbxBiWfY8_1(.dout(w_dff_A_6XTcObx51_1),.din(w_dff_A_nbxBiWfY8_1),.clk(gclk));
	jdff dff_A_anU5sl0X7_1(.dout(w_dff_A_nbxBiWfY8_1),.din(w_dff_A_anU5sl0X7_1),.clk(gclk));
	jdff dff_A_AlhORJZi8_1(.dout(w_dff_A_anU5sl0X7_1),.din(w_dff_A_AlhORJZi8_1),.clk(gclk));
	jdff dff_A_Ji7TlELM7_1(.dout(w_dff_A_AlhORJZi8_1),.din(w_dff_A_Ji7TlELM7_1),.clk(gclk));
	jdff dff_A_zVcPylW94_1(.dout(w_dff_A_Ji7TlELM7_1),.din(w_dff_A_zVcPylW94_1),.clk(gclk));
	jdff dff_A_FY0A5AWO0_1(.dout(w_dff_A_zVcPylW94_1),.din(w_dff_A_FY0A5AWO0_1),.clk(gclk));
	jdff dff_A_oQtaNTI90_1(.dout(w_dff_A_FY0A5AWO0_1),.din(w_dff_A_oQtaNTI90_1),.clk(gclk));
	jdff dff_A_7BQyAf1X2_1(.dout(w_dff_A_oQtaNTI90_1),.din(w_dff_A_7BQyAf1X2_1),.clk(gclk));
	jdff dff_A_aCpNVqY13_1(.dout(w_dff_A_7BQyAf1X2_1),.din(w_dff_A_aCpNVqY13_1),.clk(gclk));
	jdff dff_A_LqDRUReX2_1(.dout(w_dff_A_aCpNVqY13_1),.din(w_dff_A_LqDRUReX2_1),.clk(gclk));
	jdff dff_A_iI3HD5Bp2_1(.dout(w_dff_A_LqDRUReX2_1),.din(w_dff_A_iI3HD5Bp2_1),.clk(gclk));
	jdff dff_A_BYruvW6t9_1(.dout(w_dff_A_iI3HD5Bp2_1),.din(w_dff_A_BYruvW6t9_1),.clk(gclk));
	jdff dff_A_BsR5A8Rq5_1(.dout(w_dff_A_BYruvW6t9_1),.din(w_dff_A_BsR5A8Rq5_1),.clk(gclk));
	jdff dff_B_MxIFyWbc9_3(.din(G952),.dout(w_dff_B_MxIFyWbc9_3),.clk(gclk));
	jdff dff_B_R6cGR84L7_1(.din(G898),.dout(w_dff_B_R6cGR84L7_1),.clk(gclk));
	jdff dff_A_VuuFiaHe4_2(.dout(w_n253_0[2]),.din(w_dff_A_VuuFiaHe4_2),.clk(gclk));
	jdff dff_A_4n5YnmTu4_1(.dout(w_n92_0[1]),.din(w_dff_A_4n5YnmTu4_1),.clk(gclk));
	jdff dff_A_IIDNdxzU7_1(.dout(w_dff_A_4n5YnmTu4_1),.din(w_dff_A_IIDNdxzU7_1),.clk(gclk));
	jdff dff_A_UNtvUHGa2_2(.dout(w_n92_0[2]),.din(w_dff_A_UNtvUHGa2_2),.clk(gclk));
	jdff dff_A_1kIMQEqV3_2(.dout(w_dff_A_UNtvUHGa2_2),.din(w_dff_A_1kIMQEqV3_2),.clk(gclk));
	jdff dff_A_yKYSx1j20_1(.dout(w_G472_0[1]),.din(w_dff_A_yKYSx1j20_1),.clk(gclk));
	jdff dff_A_pnq9SN502_1(.dout(w_dff_A_yKYSx1j20_1),.din(w_dff_A_pnq9SN502_1),.clk(gclk));
	jdff dff_A_i5PFSqNZ8_1(.dout(w_dff_A_pnq9SN502_1),.din(w_dff_A_i5PFSqNZ8_1),.clk(gclk));
	jdff dff_A_J05vdRn43_1(.dout(w_dff_A_i5PFSqNZ8_1),.din(w_dff_A_J05vdRn43_1),.clk(gclk));
	jdff dff_A_BA8qXEPg4_1(.dout(w_dff_A_J05vdRn43_1),.din(w_dff_A_BA8qXEPg4_1),.clk(gclk));
	jdff dff_A_J4ywwvin4_1(.dout(w_dff_A_BA8qXEPg4_1),.din(w_dff_A_J4ywwvin4_1),.clk(gclk));
	jdff dff_B_DyUFSELa6_2(.din(n73),.dout(w_dff_B_DyUFSELa6_2),.clk(gclk));
	jdff dff_B_LVp1aPXk1_2(.din(w_dff_B_DyUFSELa6_2),.dout(w_dff_B_LVp1aPXk1_2),.clk(gclk));
	jdff dff_B_AE97KynP0_2(.din(w_dff_B_LVp1aPXk1_2),.dout(w_dff_B_AE97KynP0_2),.clk(gclk));
	jdff dff_B_d1Qt6Vw90_2(.din(w_dff_B_AE97KynP0_2),.dout(w_dff_B_d1Qt6Vw90_2),.clk(gclk));
	jdff dff_A_90bTC5ic7_1(.dout(w_G217_0[1]),.din(w_dff_A_90bTC5ic7_1),.clk(gclk));
	jdff dff_A_UVej9Q6S7_1(.dout(w_dff_A_90bTC5ic7_1),.din(w_dff_A_UVej9Q6S7_1),.clk(gclk));
	jdff dff_A_749vA3zO2_2(.dout(w_G217_0[2]),.din(w_dff_A_749vA3zO2_2),.clk(gclk));
	jdff dff_A_mEDlAG3r4_2(.dout(w_dff_A_749vA3zO2_2),.din(w_dff_A_mEDlAG3r4_2),.clk(gclk));
	jdff dff_A_cIAEdAzU8_2(.dout(w_dff_A_mEDlAG3r4_2),.din(w_dff_A_cIAEdAzU8_2),.clk(gclk));
	jdff dff_A_tPK35H4x3_0(.dout(w_n172_0[0]),.din(w_dff_A_tPK35H4x3_0),.clk(gclk));
	jdff dff_A_UQwIdcxJ2_0(.dout(w_dff_A_tPK35H4x3_0),.din(w_dff_A_UQwIdcxJ2_0),.clk(gclk));
	jdff dff_A_xCadTaOD3_0(.dout(w_dff_A_UQwIdcxJ2_0),.din(w_dff_A_xCadTaOD3_0),.clk(gclk));
	jdff dff_A_Co9J3NuT7_0(.dout(w_dff_A_xCadTaOD3_0),.din(w_dff_A_Co9J3NuT7_0),.clk(gclk));
	jdff dff_A_dmJ8NtAT6_0(.dout(w_dff_A_Co9J3NuT7_0),.din(w_dff_A_dmJ8NtAT6_0),.clk(gclk));
	jdff dff_A_5OU4Hzhe9_0(.dout(w_dff_A_dmJ8NtAT6_0),.din(w_dff_A_5OU4Hzhe9_0),.clk(gclk));
	jdff dff_A_ZrJcMgV21_0(.dout(w_dff_A_5OU4Hzhe9_0),.din(w_dff_A_ZrJcMgV21_0),.clk(gclk));
	jdff dff_A_XOWBeYFi1_0(.dout(w_dff_A_ZrJcMgV21_0),.din(w_dff_A_XOWBeYFi1_0),.clk(gclk));
	jdff dff_A_4vKkhNU22_0(.dout(w_dff_A_XOWBeYFi1_0),.din(w_dff_A_4vKkhNU22_0),.clk(gclk));
	jdff dff_A_4opZYrHl7_0(.dout(w_dff_A_4vKkhNU22_0),.din(w_dff_A_4opZYrHl7_0),.clk(gclk));
	jdff dff_B_aY3Muk5q7_1(.din(n171),.dout(w_dff_B_aY3Muk5q7_1),.clk(gclk));
	jdff dff_B_hdLbOZDB0_1(.din(w_dff_B_aY3Muk5q7_1),.dout(w_dff_B_hdLbOZDB0_1),.clk(gclk));
	jdff dff_B_pKaR8eaA2_1(.din(w_dff_B_hdLbOZDB0_1),.dout(w_dff_B_pKaR8eaA2_1),.clk(gclk));
	jdff dff_B_Z3x4UZAt1_0(.din(n65),.dout(w_dff_B_Z3x4UZAt1_0),.clk(gclk));
	jdff dff_B_qBlcKSpa6_0(.din(w_dff_B_Z3x4UZAt1_0),.dout(w_dff_B_qBlcKSpa6_0),.clk(gclk));
	jdff dff_B_HZXyvK1o2_0(.din(w_dff_B_qBlcKSpa6_0),.dout(w_dff_B_HZXyvK1o2_0),.clk(gclk));
	jdff dff_A_lWle4vzx4_2(.dout(w_n60_0[2]),.din(w_dff_A_lWle4vzx4_2),.clk(gclk));
	jdff dff_A_ND1zml4C2_2(.dout(w_dff_A_lWle4vzx4_2),.din(w_dff_A_ND1zml4C2_2),.clk(gclk));
	jdff dff_A_zGKtC6DJ0_2(.dout(w_dff_A_ND1zml4C2_2),.din(w_dff_A_zGKtC6DJ0_2),.clk(gclk));
	jdff dff_A_qbrnQueL8_2(.dout(w_dff_A_zGKtC6DJ0_2),.din(w_dff_A_qbrnQueL8_2),.clk(gclk));
	jdff dff_A_DE4xhmAQ3_0(.dout(w_n59_0[0]),.din(w_dff_A_DE4xhmAQ3_0),.clk(gclk));
	jdff dff_A_wrXkq0xj6_0(.dout(w_dff_A_DE4xhmAQ3_0),.din(w_dff_A_wrXkq0xj6_0),.clk(gclk));
	jdff dff_A_F0OlzLAD1_0(.dout(w_dff_A_wrXkq0xj6_0),.din(w_dff_A_F0OlzLAD1_0),.clk(gclk));
	jdff dff_A_NYHFwaqr6_0(.dout(w_n70_1[0]),.din(w_dff_A_NYHFwaqr6_0),.clk(gclk));
	jdff dff_A_LY3FGZA26_0(.dout(w_dff_A_NYHFwaqr6_0),.din(w_dff_A_LY3FGZA26_0),.clk(gclk));
	jdff dff_A_09DJ5dNl8_0(.dout(w_dff_A_LY3FGZA26_0),.din(w_dff_A_09DJ5dNl8_0),.clk(gclk));
	jdff dff_A_ZsGqYRqj6_0(.dout(w_dff_A_09DJ5dNl8_0),.din(w_dff_A_ZsGqYRqj6_0),.clk(gclk));
	jdff dff_A_TJWDZQVb4_0(.dout(w_dff_A_ZsGqYRqj6_0),.din(w_dff_A_TJWDZQVb4_0),.clk(gclk));
	jdff dff_A_dkTleeez0_0(.dout(w_dff_A_TJWDZQVb4_0),.din(w_dff_A_dkTleeez0_0),.clk(gclk));
	jdff dff_A_KgoQ2qci2_2(.dout(w_n70_1[2]),.din(w_dff_A_KgoQ2qci2_2),.clk(gclk));
	jdff dff_A_5C5HgrQm5_2(.dout(w_dff_A_KgoQ2qci2_2),.din(w_dff_A_5C5HgrQm5_2),.clk(gclk));
	jdff dff_A_g1cQAKUA6_2(.dout(w_dff_A_5C5HgrQm5_2),.din(w_dff_A_g1cQAKUA6_2),.clk(gclk));
	jdff dff_A_iVMlshMV6_2(.dout(w_dff_A_g1cQAKUA6_2),.din(w_dff_A_iVMlshMV6_2),.clk(gclk));
	jdff dff_A_yQejMPDK3_0(.dout(w_n276_1[0]),.din(w_dff_A_yQejMPDK3_0),.clk(gclk));
	jdff dff_B_UXWqgLLL9_3(.din(n276),.dout(w_dff_B_UXWqgLLL9_3),.clk(gclk));
	jdff dff_B_7FRH8gBm4_1(.din(n195),.dout(w_dff_B_7FRH8gBm4_1),.clk(gclk));
	jdff dff_B_wYNYSM4x6_1(.din(w_dff_B_7FRH8gBm4_1),.dout(w_dff_B_wYNYSM4x6_1),.clk(gclk));
	jdff dff_B_fMGbrcGh6_1(.din(w_dff_B_wYNYSM4x6_1),.dout(w_dff_B_fMGbrcGh6_1),.clk(gclk));
	jdff dff_B_gK9l3Sqx9_1(.din(w_dff_B_fMGbrcGh6_1),.dout(w_dff_B_gK9l3Sqx9_1),.clk(gclk));
	jdff dff_B_Jx9tTa653_1(.din(w_dff_B_gK9l3Sqx9_1),.dout(w_dff_B_Jx9tTa653_1),.clk(gclk));
	jdff dff_A_ID1k2XuY2_0(.dout(w_n117_0[0]),.din(w_dff_A_ID1k2XuY2_0),.clk(gclk));
	jdff dff_A_d7FDJCNO2_0(.dout(w_dff_A_ID1k2XuY2_0),.din(w_dff_A_d7FDJCNO2_0),.clk(gclk));
	jdff dff_A_XvdFCzrw3_0(.dout(w_dff_A_d7FDJCNO2_0),.din(w_dff_A_XvdFCzrw3_0),.clk(gclk));
	jdff dff_A_plQxmdKp7_0(.dout(w_dff_A_XvdFCzrw3_0),.din(w_dff_A_plQxmdKp7_0),.clk(gclk));
	jdff dff_A_vUaupqrr8_0(.dout(w_dff_A_plQxmdKp7_0),.din(w_dff_A_vUaupqrr8_0),.clk(gclk));
	jdff dff_A_gB9U7PJY9_0(.dout(w_dff_A_vUaupqrr8_0),.din(w_dff_A_gB9U7PJY9_0),.clk(gclk));
	jdff dff_A_cMugvh9q4_0(.dout(w_dff_A_gB9U7PJY9_0),.din(w_dff_A_cMugvh9q4_0),.clk(gclk));
	jdff dff_A_TDbpR4YG0_0(.dout(w_dff_A_cMugvh9q4_0),.din(w_dff_A_TDbpR4YG0_0),.clk(gclk));
	jdff dff_A_2UAMgQJC5_0(.dout(w_dff_A_TDbpR4YG0_0),.din(w_dff_A_2UAMgQJC5_0),.clk(gclk));
	jdff dff_A_0FoaCd5f8_0(.dout(w_dff_A_2UAMgQJC5_0),.din(w_dff_A_0FoaCd5f8_0),.clk(gclk));
	jdff dff_A_c18q2Jzj9_0(.dout(w_dff_A_0FoaCd5f8_0),.din(w_dff_A_c18q2Jzj9_0),.clk(gclk));
	jdff dff_A_O0ethJcU8_0(.dout(w_dff_A_c18q2Jzj9_0),.din(w_dff_A_O0ethJcU8_0),.clk(gclk));
	jdff dff_B_EMzFG6GW9_1(.din(n113),.dout(w_dff_B_EMzFG6GW9_1),.clk(gclk));
	jdff dff_B_2VYMP6Op9_1(.din(w_dff_B_EMzFG6GW9_1),.dout(w_dff_B_2VYMP6Op9_1),.clk(gclk));
	jdff dff_B_skuoW42i7_2(.din(G227),.dout(w_dff_B_skuoW42i7_2),.clk(gclk));
	jdff dff_A_6D5aWB4x7_0(.dout(w_G140_0[0]),.din(w_dff_A_6D5aWB4x7_0),.clk(gclk));
	jdff dff_A_O3vkfvPD5_0(.dout(w_dff_A_6D5aWB4x7_0),.din(w_dff_A_O3vkfvPD5_0),.clk(gclk));
	jdff dff_A_xNFSjN763_0(.dout(w_dff_A_O3vkfvPD5_0),.din(w_dff_A_xNFSjN763_0),.clk(gclk));
	jdff dff_A_euZgJ5on4_0(.dout(w_dff_A_xNFSjN763_0),.din(w_dff_A_euZgJ5on4_0),.clk(gclk));
	jdff dff_A_ZlbdMtWu2_0(.dout(w_dff_A_euZgJ5on4_0),.din(w_dff_A_ZlbdMtWu2_0),.clk(gclk));
	jdff dff_A_QbEWsmZH7_0(.dout(w_dff_A_ZlbdMtWu2_0),.din(w_dff_A_QbEWsmZH7_0),.clk(gclk));
	jdff dff_A_TdzEgtCD0_0(.dout(w_dff_A_QbEWsmZH7_0),.din(w_dff_A_TdzEgtCD0_0),.clk(gclk));
	jdff dff_A_y8dDQ0a08_0(.dout(w_dff_A_TdzEgtCD0_0),.din(w_dff_A_y8dDQ0a08_0),.clk(gclk));
	jdff dff_A_5zEdiTvk8_0(.dout(w_dff_A_y8dDQ0a08_0),.din(w_dff_A_5zEdiTvk8_0),.clk(gclk));
	jdff dff_A_RJ5QVG8f1_0(.dout(w_dff_A_5zEdiTvk8_0),.din(w_dff_A_RJ5QVG8f1_0),.clk(gclk));
	jdff dff_A_wKRISSfC8_0(.dout(w_dff_A_RJ5QVG8f1_0),.din(w_dff_A_wKRISSfC8_0),.clk(gclk));
	jdff dff_A_ErJwq7to0_0(.dout(w_dff_A_wKRISSfC8_0),.din(w_dff_A_ErJwq7to0_0),.clk(gclk));
	jdff dff_A_e3lVX8gh2_2(.dout(w_G469_0[2]),.din(w_dff_A_e3lVX8gh2_2),.clk(gclk));
	jdff dff_A_gIN7R3uf1_2(.dout(w_dff_A_e3lVX8gh2_2),.din(w_dff_A_gIN7R3uf1_2),.clk(gclk));
	jdff dff_A_mERP0ZkL1_2(.dout(w_dff_A_gIN7R3uf1_2),.din(w_dff_A_mERP0ZkL1_2),.clk(gclk));
	jdff dff_A_c70Dbpyw4_2(.dout(w_dff_A_mERP0ZkL1_2),.din(w_dff_A_c70Dbpyw4_2),.clk(gclk));
	jdff dff_A_7ZWMuhfi8_2(.dout(w_dff_A_c70Dbpyw4_2),.din(w_dff_A_7ZWMuhfi8_2),.clk(gclk));
	jdff dff_A_TyI5Y8M08_2(.dout(w_dff_A_7ZWMuhfi8_2),.din(w_dff_A_TyI5Y8M08_2),.clk(gclk));
	jdff dff_B_WcRU6Qft7_2(.din(n274),.dout(w_dff_B_WcRU6Qft7_2),.clk(gclk));
	jdff dff_B_7quUQe1I0_2(.din(w_dff_B_WcRU6Qft7_2),.dout(w_dff_B_7quUQe1I0_2),.clk(gclk));
	jdff dff_B_pJ0ykcTy3_2(.din(w_dff_B_7quUQe1I0_2),.dout(w_dff_B_pJ0ykcTy3_2),.clk(gclk));
	jdff dff_A_aO2f3qcc7_0(.dout(w_n112_0[0]),.din(w_dff_A_aO2f3qcc7_0),.clk(gclk));
	jdff dff_A_XNfeC4qt2_0(.dout(w_dff_A_aO2f3qcc7_0),.din(w_dff_A_XNfeC4qt2_0),.clk(gclk));
	jdff dff_A_VthqGAlY9_0(.dout(w_dff_A_XNfeC4qt2_0),.din(w_dff_A_VthqGAlY9_0),.clk(gclk));
	jdff dff_A_tqhHZpRV0_0(.dout(w_dff_A_VthqGAlY9_0),.din(w_dff_A_tqhHZpRV0_0),.clk(gclk));
	jdff dff_B_7iPPSUpd2_1(.din(n111),.dout(w_dff_B_7iPPSUpd2_1),.clk(gclk));
	jdff dff_A_5VXt3w777_0(.dout(w_n70_3[0]),.din(w_dff_A_5VXt3w777_0),.clk(gclk));
	jdff dff_A_7Jpnt4JB2_0(.dout(w_dff_A_5VXt3w777_0),.din(w_dff_A_7Jpnt4JB2_0),.clk(gclk));
	jdff dff_A_PqzGkrR80_0(.dout(w_dff_A_7Jpnt4JB2_0),.din(w_dff_A_PqzGkrR80_0),.clk(gclk));
	jdff dff_A_HEbrDUYk4_0(.dout(w_dff_A_PqzGkrR80_0),.din(w_dff_A_HEbrDUYk4_0),.clk(gclk));
	jdff dff_A_xGppPr3k5_1(.dout(w_G234_0[1]),.din(w_dff_A_xGppPr3k5_1),.clk(gclk));
	jdff dff_A_3T0Mu2XP9_2(.dout(w_G234_0[2]),.din(w_dff_A_3T0Mu2XP9_2),.clk(gclk));
	jdff dff_A_0asksFzo1_1(.dout(w_G221_0[1]),.din(w_dff_A_0asksFzo1_1),.clk(gclk));
	jdff dff_A_WhLdinJl8_1(.dout(w_dff_A_0asksFzo1_1),.din(w_dff_A_WhLdinJl8_1),.clk(gclk));
	jdff dff_A_L7rbIXSV3_1(.dout(w_n216_0[1]),.din(w_dff_A_L7rbIXSV3_1),.clk(gclk));
	jdff dff_B_f02cB3R30_1(.din(n215),.dout(w_dff_B_f02cB3R30_1),.clk(gclk));
	jdff dff_B_JeWlBlYS1_1(.din(w_dff_B_f02cB3R30_1),.dout(w_dff_B_JeWlBlYS1_1),.clk(gclk));
	jdff dff_B_hXeRC8QT0_1(.din(w_dff_B_JeWlBlYS1_1),.dout(w_dff_B_hXeRC8QT0_1),.clk(gclk));
	jdff dff_A_x1lg016P1_0(.dout(w_n107_0[0]),.din(w_dff_A_x1lg016P1_0),.clk(gclk));
	jdff dff_A_j272sTqQ3_0(.dout(w_dff_A_x1lg016P1_0),.din(w_dff_A_j272sTqQ3_0),.clk(gclk));
	jdff dff_A_gLpiljix5_0(.dout(w_dff_A_j272sTqQ3_0),.din(w_dff_A_gLpiljix5_0),.clk(gclk));
	jdff dff_A_9Vav6S578_0(.dout(w_dff_A_gLpiljix5_0),.din(w_dff_A_9Vav6S578_0),.clk(gclk));
	jdff dff_A_vhbPjJiy3_0(.dout(w_dff_A_9Vav6S578_0),.din(w_dff_A_vhbPjJiy3_0),.clk(gclk));
	jdff dff_A_H88aFHDB1_0(.dout(w_dff_A_vhbPjJiy3_0),.din(w_dff_A_H88aFHDB1_0),.clk(gclk));
	jdff dff_A_DHK4VAkF2_0(.dout(w_dff_A_H88aFHDB1_0),.din(w_dff_A_DHK4VAkF2_0),.clk(gclk));
	jdff dff_A_ft3kdH7l3_0(.dout(w_dff_A_DHK4VAkF2_0),.din(w_dff_A_ft3kdH7l3_0),.clk(gclk));
	jdff dff_A_OI8DS2hM9_0(.dout(w_dff_A_ft3kdH7l3_0),.din(w_dff_A_OI8DS2hM9_0),.clk(gclk));
	jdff dff_A_oNSKDJch6_0(.dout(w_dff_A_OI8DS2hM9_0),.din(w_dff_A_oNSKDJch6_0),.clk(gclk));
	jdff dff_A_EBXwMR433_0(.dout(w_dff_A_oNSKDJch6_0),.din(w_dff_A_EBXwMR433_0),.clk(gclk));
	jdff dff_A_ZhXSyGLz0_0(.dout(w_dff_A_EBXwMR433_0),.din(w_dff_A_ZhXSyGLz0_0),.clk(gclk));
	jdff dff_B_jhzHQqfo5_1(.din(n104),.dout(w_dff_B_jhzHQqfo5_1),.clk(gclk));
	jdff dff_A_hGaPrqic9_0(.dout(w_G125_0[0]),.din(w_dff_A_hGaPrqic9_0),.clk(gclk));
	jdff dff_A_BUEBrPCd2_0(.dout(w_dff_A_hGaPrqic9_0),.din(w_dff_A_BUEBrPCd2_0),.clk(gclk));
	jdff dff_A_hKYDeIqG7_0(.dout(w_dff_A_BUEBrPCd2_0),.din(w_dff_A_hKYDeIqG7_0),.clk(gclk));
	jdff dff_A_LK2anFOc8_0(.dout(w_dff_A_hKYDeIqG7_0),.din(w_dff_A_LK2anFOc8_0),.clk(gclk));
	jdff dff_A_GoHPD5xI5_0(.dout(w_dff_A_LK2anFOc8_0),.din(w_dff_A_GoHPD5xI5_0),.clk(gclk));
	jdff dff_A_MP3BtIz50_0(.dout(w_dff_A_GoHPD5xI5_0),.din(w_dff_A_MP3BtIz50_0),.clk(gclk));
	jdff dff_A_2EprVAK18_0(.dout(w_dff_A_MP3BtIz50_0),.din(w_dff_A_2EprVAK18_0),.clk(gclk));
	jdff dff_A_e5FFRQJK9_0(.dout(w_dff_A_2EprVAK18_0),.din(w_dff_A_e5FFRQJK9_0),.clk(gclk));
	jdff dff_A_71AJuITo6_0(.dout(w_dff_A_e5FFRQJK9_0),.din(w_dff_A_71AJuITo6_0),.clk(gclk));
	jdff dff_A_ABJqDcHw9_0(.dout(w_dff_A_71AJuITo6_0),.din(w_dff_A_ABJqDcHw9_0),.clk(gclk));
	jdff dff_A_WCLJcx8e0_0(.dout(w_dff_A_ABJqDcHw9_0),.din(w_dff_A_WCLJcx8e0_0),.clk(gclk));
	jdff dff_A_wEwstavb2_0(.dout(w_dff_A_WCLJcx8e0_0),.din(w_dff_A_wEwstavb2_0),.clk(gclk));
	jdff dff_A_guNlDc5m9_1(.dout(w_G125_0[1]),.din(w_dff_A_guNlDc5m9_1),.clk(gclk));
	jdff dff_A_oICwdoW57_1(.dout(w_dff_A_guNlDc5m9_1),.din(w_dff_A_oICwdoW57_1),.clk(gclk));
	jdff dff_B_8hXZiefv1_2(.din(G224),.dout(w_dff_B_8hXZiefv1_2),.clk(gclk));
	jdff dff_A_rfpRIPBm1_0(.dout(w_n103_0[0]),.din(w_dff_A_rfpRIPBm1_0),.clk(gclk));
	jdff dff_A_w8A4JYm67_0(.dout(w_dff_A_rfpRIPBm1_0),.din(w_dff_A_w8A4JYm67_0),.clk(gclk));
	jdff dff_A_ADPXycaA9_0(.dout(w_dff_A_w8A4JYm67_0),.din(w_dff_A_ADPXycaA9_0),.clk(gclk));
	jdff dff_A_FdJbRLZR0_0(.dout(w_dff_A_ADPXycaA9_0),.din(w_dff_A_FdJbRLZR0_0),.clk(gclk));
	jdff dff_A_JAW0FIg22_0(.dout(w_dff_A_FdJbRLZR0_0),.din(w_dff_A_JAW0FIg22_0),.clk(gclk));
	jdff dff_A_LW17otL16_0(.dout(w_dff_A_JAW0FIg22_0),.din(w_dff_A_LW17otL16_0),.clk(gclk));
	jdff dff_A_eFpoyJQ54_0(.dout(w_dff_A_LW17otL16_0),.din(w_dff_A_eFpoyJQ54_0),.clk(gclk));
	jdff dff_A_0ztDfp9y9_0(.dout(w_dff_A_eFpoyJQ54_0),.din(w_dff_A_0ztDfp9y9_0),.clk(gclk));
	jdff dff_A_7MthCdBr7_0(.dout(w_dff_A_0ztDfp9y9_0),.din(w_dff_A_7MthCdBr7_0),.clk(gclk));
	jdff dff_A_TzaH7j9q2_0(.dout(w_dff_A_7MthCdBr7_0),.din(w_dff_A_TzaH7j9q2_0),.clk(gclk));
	jdff dff_A_yMA7LU7d8_0(.dout(w_dff_A_TzaH7j9q2_0),.din(w_dff_A_yMA7LU7d8_0),.clk(gclk));
	jdff dff_A_9wStfIcu0_0(.dout(w_dff_A_yMA7LU7d8_0),.din(w_dff_A_9wStfIcu0_0),.clk(gclk));
	jdff dff_A_Mjp2c5pP9_0(.dout(w_dff_A_9wStfIcu0_0),.din(w_dff_A_Mjp2c5pP9_0),.clk(gclk));
	jdff dff_B_FXE00Kze7_1(.din(n99),.dout(w_dff_B_FXE00Kze7_1),.clk(gclk));
	jdff dff_A_SZ1Nm9Cs6_0(.dout(w_G107_0[0]),.din(w_dff_A_SZ1Nm9Cs6_0),.clk(gclk));
	jdff dff_A_b8kOHhoQ6_0(.dout(w_dff_A_SZ1Nm9Cs6_0),.din(w_dff_A_b8kOHhoQ6_0),.clk(gclk));
	jdff dff_A_3BvIEyqz4_0(.dout(w_dff_A_b8kOHhoQ6_0),.din(w_dff_A_3BvIEyqz4_0),.clk(gclk));
	jdff dff_A_fl5DajHF6_0(.dout(w_dff_A_3BvIEyqz4_0),.din(w_dff_A_fl5DajHF6_0),.clk(gclk));
	jdff dff_A_f9VF20vk0_0(.dout(w_dff_A_fl5DajHF6_0),.din(w_dff_A_f9VF20vk0_0),.clk(gclk));
	jdff dff_A_N8KbK16P5_0(.dout(w_dff_A_f9VF20vk0_0),.din(w_dff_A_N8KbK16P5_0),.clk(gclk));
	jdff dff_A_ZrfOKXBg8_0(.dout(w_dff_A_N8KbK16P5_0),.din(w_dff_A_ZrfOKXBg8_0),.clk(gclk));
	jdff dff_A_XTL9CeRp9_0(.dout(w_dff_A_ZrfOKXBg8_0),.din(w_dff_A_XTL9CeRp9_0),.clk(gclk));
	jdff dff_A_TeErh5ES0_0(.dout(w_dff_A_XTL9CeRp9_0),.din(w_dff_A_TeErh5ES0_0),.clk(gclk));
	jdff dff_A_w9oDyhL51_0(.dout(w_dff_A_TeErh5ES0_0),.din(w_dff_A_w9oDyhL51_0),.clk(gclk));
	jdff dff_A_DYKoNI6Y5_0(.dout(w_dff_A_w9oDyhL51_0),.din(w_dff_A_DYKoNI6Y5_0),.clk(gclk));
	jdff dff_A_w6XTsMsq8_0(.dout(w_dff_A_DYKoNI6Y5_0),.din(w_dff_A_w6XTsMsq8_0),.clk(gclk));
	jdff dff_A_97FbSwfK4_0(.dout(w_G104_0[0]),.din(w_dff_A_97FbSwfK4_0),.clk(gclk));
	jdff dff_A_GoqsyYIm8_0(.dout(w_dff_A_97FbSwfK4_0),.din(w_dff_A_GoqsyYIm8_0),.clk(gclk));
	jdff dff_A_T4Eaq92Z3_0(.dout(w_dff_A_GoqsyYIm8_0),.din(w_dff_A_T4Eaq92Z3_0),.clk(gclk));
	jdff dff_A_zElM6zFu1_0(.dout(w_dff_A_T4Eaq92Z3_0),.din(w_dff_A_zElM6zFu1_0),.clk(gclk));
	jdff dff_A_DRxUm7kI2_0(.dout(w_dff_A_zElM6zFu1_0),.din(w_dff_A_DRxUm7kI2_0),.clk(gclk));
	jdff dff_A_3yPtjfDy8_0(.dout(w_dff_A_DRxUm7kI2_0),.din(w_dff_A_3yPtjfDy8_0),.clk(gclk));
	jdff dff_A_e8loeeor5_0(.dout(w_dff_A_3yPtjfDy8_0),.din(w_dff_A_e8loeeor5_0),.clk(gclk));
	jdff dff_A_05FENPcz7_0(.dout(w_dff_A_e8loeeor5_0),.din(w_dff_A_05FENPcz7_0),.clk(gclk));
	jdff dff_A_ec6pBWD25_0(.dout(w_dff_A_05FENPcz7_0),.din(w_dff_A_ec6pBWD25_0),.clk(gclk));
	jdff dff_A_9IfFmerl9_0(.dout(w_dff_A_ec6pBWD25_0),.din(w_dff_A_9IfFmerl9_0),.clk(gclk));
	jdff dff_A_W4DPFxFO0_0(.dout(w_dff_A_9IfFmerl9_0),.din(w_dff_A_W4DPFxFO0_0),.clk(gclk));
	jdff dff_A_PB4RuL8e9_0(.dout(w_dff_A_W4DPFxFO0_0),.din(w_dff_A_PB4RuL8e9_0),.clk(gclk));
	jdff dff_A_WtxmHIdG9_1(.dout(w_G104_0[1]),.din(w_dff_A_WtxmHIdG9_1),.clk(gclk));
	jdff dff_A_ADaMUmKc6_1(.dout(w_dff_A_WtxmHIdG9_1),.din(w_dff_A_ADaMUmKc6_1),.clk(gclk));
	jdff dff_A_Xk15ibSQ5_1(.dout(w_G122_1[1]),.din(w_dff_A_Xk15ibSQ5_1),.clk(gclk));
	jdff dff_A_kOA2vvfP0_1(.dout(w_G122_0[1]),.din(w_dff_A_kOA2vvfP0_1),.clk(gclk));
	jdff dff_A_GoWajBuW7_1(.dout(w_dff_A_kOA2vvfP0_1),.din(w_dff_A_GoWajBuW7_1),.clk(gclk));
	jdff dff_A_UdgX3NmM7_1(.dout(w_dff_A_GoWajBuW7_1),.din(w_dff_A_UdgX3NmM7_1),.clk(gclk));
	jdff dff_A_huAXcbKv0_1(.dout(w_dff_A_UdgX3NmM7_1),.din(w_dff_A_huAXcbKv0_1),.clk(gclk));
	jdff dff_A_Jqqv8qbg7_1(.dout(w_dff_A_huAXcbKv0_1),.din(w_dff_A_Jqqv8qbg7_1),.clk(gclk));
	jdff dff_A_vATM0Lp49_1(.dout(w_dff_A_Jqqv8qbg7_1),.din(w_dff_A_vATM0Lp49_1),.clk(gclk));
	jdff dff_A_RV81MCiQ5_1(.dout(w_dff_A_vATM0Lp49_1),.din(w_dff_A_RV81MCiQ5_1),.clk(gclk));
	jdff dff_A_f7OK7zOE3_1(.dout(w_dff_A_RV81MCiQ5_1),.din(w_dff_A_f7OK7zOE3_1),.clk(gclk));
	jdff dff_A_YsiZRDlq9_1(.dout(w_dff_A_f7OK7zOE3_1),.din(w_dff_A_YsiZRDlq9_1),.clk(gclk));
	jdff dff_A_lJjo43g72_1(.dout(w_dff_A_YsiZRDlq9_1),.din(w_dff_A_lJjo43g72_1),.clk(gclk));
	jdff dff_A_d0Eel5RY2_1(.dout(w_dff_A_lJjo43g72_1),.din(w_dff_A_d0Eel5RY2_1),.clk(gclk));
	jdff dff_A_EyY3UJfQ7_1(.dout(w_dff_A_d0Eel5RY2_1),.din(w_dff_A_EyY3UJfQ7_1),.clk(gclk));
	jdff dff_A_EeE4pWsK2_2(.dout(w_G122_0[2]),.din(w_dff_A_EeE4pWsK2_2),.clk(gclk));
	jdff dff_A_tyLlt4Ug9_1(.dout(w_G110_1[1]),.din(w_dff_A_tyLlt4Ug9_1),.clk(gclk));
	jdff dff_A_etytuETZ9_1(.dout(w_dff_A_tyLlt4Ug9_1),.din(w_dff_A_etytuETZ9_1),.clk(gclk));
	jdff dff_A_11apbKMy5_1(.dout(w_dff_A_etytuETZ9_1),.din(w_dff_A_11apbKMy5_1),.clk(gclk));
	jdff dff_A_GI9ubTPs6_1(.dout(w_dff_A_11apbKMy5_1),.din(w_dff_A_GI9ubTPs6_1),.clk(gclk));
	jdff dff_A_1FZCsts23_1(.dout(w_dff_A_GI9ubTPs6_1),.din(w_dff_A_1FZCsts23_1),.clk(gclk));
	jdff dff_A_S7LbMjC51_1(.dout(w_G110_0[1]),.din(w_dff_A_S7LbMjC51_1),.clk(gclk));
	jdff dff_A_ObpxlGIK4_1(.dout(w_dff_A_S7LbMjC51_1),.din(w_dff_A_ObpxlGIK4_1),.clk(gclk));
	jdff dff_A_0NJh9BDP9_1(.dout(w_dff_A_ObpxlGIK4_1),.din(w_dff_A_0NJh9BDP9_1),.clk(gclk));
	jdff dff_A_xzrtJekW4_1(.dout(w_dff_A_0NJh9BDP9_1),.din(w_dff_A_xzrtJekW4_1),.clk(gclk));
	jdff dff_A_wNZ0DuLF0_1(.dout(w_dff_A_xzrtJekW4_1),.din(w_dff_A_wNZ0DuLF0_1),.clk(gclk));
	jdff dff_A_95ahYNiN7_1(.dout(w_dff_A_wNZ0DuLF0_1),.din(w_dff_A_95ahYNiN7_1),.clk(gclk));
	jdff dff_A_6vbxWAv54_1(.dout(w_dff_A_95ahYNiN7_1),.din(w_dff_A_6vbxWAv54_1),.clk(gclk));
	jdff dff_A_O4L5RZ7b7_1(.dout(w_dff_A_6vbxWAv54_1),.din(w_dff_A_O4L5RZ7b7_1),.clk(gclk));
	jdff dff_A_9G3HKwwo0_1(.dout(w_dff_A_O4L5RZ7b7_1),.din(w_dff_A_9G3HKwwo0_1),.clk(gclk));
	jdff dff_A_qFoE6ANk9_1(.dout(w_dff_A_9G3HKwwo0_1),.din(w_dff_A_qFoE6ANk9_1),.clk(gclk));
	jdff dff_A_fxY1ZImU6_1(.dout(w_dff_A_qFoE6ANk9_1),.din(w_dff_A_fxY1ZImU6_1),.clk(gclk));
	jdff dff_A_6FnxbwUU6_1(.dout(w_dff_A_fxY1ZImU6_1),.din(w_dff_A_6FnxbwUU6_1),.clk(gclk));
	jdff dff_A_wCCgcxh21_1(.dout(w_n70_0[1]),.din(w_dff_A_wCCgcxh21_1),.clk(gclk));
	jdff dff_A_hjgtmlav3_1(.dout(w_dff_A_wCCgcxh21_1),.din(w_dff_A_hjgtmlav3_1),.clk(gclk));
	jdff dff_A_ntsyURLv6_1(.dout(w_dff_A_hjgtmlav3_1),.din(w_dff_A_ntsyURLv6_1),.clk(gclk));
	jdff dff_A_sq6nP6G67_1(.dout(w_dff_A_ntsyURLv6_1),.din(w_dff_A_sq6nP6G67_1),.clk(gclk));
	jdff dff_A_dSjSA72F1_1(.dout(w_n97_0[1]),.din(w_dff_A_dSjSA72F1_1),.clk(gclk));
	jdff dff_A_hwV4ctbQ9_1(.dout(w_dff_A_dSjSA72F1_1),.din(w_dff_A_hwV4ctbQ9_1),.clk(gclk));
	jdff dff_A_RT5C6dx18_1(.dout(w_dff_A_hwV4ctbQ9_1),.din(w_dff_A_RT5C6dx18_1),.clk(gclk));
	jdff dff_A_5QxyESWo5_1(.dout(w_dff_A_RT5C6dx18_1),.din(w_dff_A_5QxyESWo5_1),.clk(gclk));
	jdff dff_A_3twR1F1A9_0(.dout(w_n95_0[0]),.din(w_dff_A_3twR1F1A9_0),.clk(gclk));
	jdff dff_A_lly5St5y0_0(.dout(w_dff_A_3twR1F1A9_0),.din(w_dff_A_lly5St5y0_0),.clk(gclk));
	jdff dff_A_E0hdVmTV6_0(.dout(w_dff_A_lly5St5y0_0),.din(w_dff_A_E0hdVmTV6_0),.clk(gclk));
	jdff dff_A_izuiToZY1_0(.dout(w_dff_A_E0hdVmTV6_0),.din(w_dff_A_izuiToZY1_0),.clk(gclk));
	jdff dff_A_ASA7AT1X9_0(.dout(w_dff_A_izuiToZY1_0),.din(w_dff_A_ASA7AT1X9_0),.clk(gclk));
	jdff dff_A_GezeG4B26_1(.dout(w_n95_0[1]),.din(w_dff_A_GezeG4B26_1),.clk(gclk));
	jdff dff_A_94DAfcxq4_1(.dout(w_dff_A_GezeG4B26_1),.din(w_dff_A_94DAfcxq4_1),.clk(gclk));
	jdff dff_A_2Qz32MAY7_1(.dout(w_dff_A_94DAfcxq4_1),.din(w_dff_A_2Qz32MAY7_1),.clk(gclk));
	jdff dff_A_3vajMS4s9_1(.dout(w_dff_A_2Qz32MAY7_1),.din(w_dff_A_3vajMS4s9_1),.clk(gclk));
	jdff dff_A_xnFTH5ZX1_1(.dout(w_dff_A_3vajMS4s9_1),.din(w_dff_A_xnFTH5ZX1_1),.clk(gclk));
	jdff dff_A_9v5QviIV3_2(.dout(w_G902_3[2]),.din(w_dff_A_9v5QviIV3_2),.clk(gclk));
	jdff dff_A_tUC0hJ4s2_2(.dout(w_dff_A_9v5QviIV3_2),.din(w_dff_A_tUC0hJ4s2_2),.clk(gclk));
	jdff dff_A_uj7b49bG5_2(.dout(w_dff_A_tUC0hJ4s2_2),.din(w_dff_A_uj7b49bG5_2),.clk(gclk));
	jdff dff_A_71sARR4R6_2(.dout(w_dff_A_uj7b49bG5_2),.din(w_dff_A_71sARR4R6_2),.clk(gclk));
	jdff dff_A_dFpJWWmH4_2(.dout(w_dff_A_71sARR4R6_2),.din(w_dff_A_dFpJWWmH4_2),.clk(gclk));
	jdff dff_A_eXeabmUB1_2(.dout(w_dff_A_dFpJWWmH4_2),.din(w_dff_A_eXeabmUB1_2),.clk(gclk));
	jdff dff_A_WylMPeS41_2(.dout(w_dff_A_eXeabmUB1_2),.din(w_dff_A_WylMPeS41_2),.clk(gclk));
	jdff dff_A_C8ITO4682_1(.dout(w_G214_0[1]),.din(w_dff_A_C8ITO4682_1),.clk(gclk));
	jdff dff_A_omvqrot23_0(.dout(w_n90_0[0]),.din(w_dff_A_omvqrot23_0),.clk(gclk));
	jdff dff_A_z1FKsQwb4_0(.dout(w_dff_A_omvqrot23_0),.din(w_dff_A_z1FKsQwb4_0),.clk(gclk));
	jdff dff_A_LVNl98VB2_0(.dout(w_dff_A_z1FKsQwb4_0),.din(w_dff_A_LVNl98VB2_0),.clk(gclk));
	jdff dff_A_YdIrpSVj6_0(.dout(w_dff_A_LVNl98VB2_0),.din(w_dff_A_YdIrpSVj6_0),.clk(gclk));
	jdff dff_A_LJ8Gi4uF8_0(.dout(w_dff_A_YdIrpSVj6_0),.din(w_dff_A_LJ8Gi4uF8_0),.clk(gclk));
	jdff dff_A_DZEGczG83_0(.dout(w_dff_A_LJ8Gi4uF8_0),.din(w_dff_A_DZEGczG83_0),.clk(gclk));
	jdff dff_A_KMClJIRV1_0(.dout(w_dff_A_DZEGczG83_0),.din(w_dff_A_KMClJIRV1_0),.clk(gclk));
	jdff dff_A_M1oAQNKf2_0(.dout(w_dff_A_KMClJIRV1_0),.din(w_dff_A_M1oAQNKf2_0),.clk(gclk));
	jdff dff_A_cNNtsd1I4_0(.dout(w_dff_A_M1oAQNKf2_0),.din(w_dff_A_cNNtsd1I4_0),.clk(gclk));
	jdff dff_A_qtYt3qJj9_0(.dout(w_dff_A_cNNtsd1I4_0),.din(w_dff_A_qtYt3qJj9_0),.clk(gclk));
	jdff dff_A_QEH7dcRk1_0(.dout(w_dff_A_qtYt3qJj9_0),.din(w_dff_A_QEH7dcRk1_0),.clk(gclk));
	jdff dff_A_wSqvZeYI9_0(.dout(w_dff_A_QEH7dcRk1_0),.din(w_dff_A_wSqvZeYI9_0),.clk(gclk));
	jdff dff_A_UaBnAubx0_0(.dout(w_G953_1[0]),.din(w_dff_A_UaBnAubx0_0),.clk(gclk));
	jdff dff_A_c6EKCiTg3_0(.dout(w_dff_A_UaBnAubx0_0),.din(w_dff_A_c6EKCiTg3_0),.clk(gclk));
	jdff dff_A_dAvRHgeN0_0(.dout(w_dff_A_c6EKCiTg3_0),.din(w_dff_A_dAvRHgeN0_0),.clk(gclk));
	jdff dff_A_hkaXSMhD4_0(.dout(w_dff_A_dAvRHgeN0_0),.din(w_dff_A_hkaXSMhD4_0),.clk(gclk));
	jdff dff_A_ceF5DLAr8_0(.dout(w_dff_A_hkaXSMhD4_0),.din(w_dff_A_ceF5DLAr8_0),.clk(gclk));
	jdff dff_A_v9tLWDIF1_0(.dout(w_dff_A_ceF5DLAr8_0),.din(w_dff_A_v9tLWDIF1_0),.clk(gclk));
	jdff dff_A_xgo6MV9X2_0(.dout(w_dff_A_v9tLWDIF1_0),.din(w_dff_A_xgo6MV9X2_0),.clk(gclk));
	jdff dff_A_CBh5iyhF0_0(.dout(w_dff_A_xgo6MV9X2_0),.din(w_dff_A_CBh5iyhF0_0),.clk(gclk));
	jdff dff_A_VLo057qZ4_0(.dout(w_dff_A_CBh5iyhF0_0),.din(w_dff_A_VLo057qZ4_0),.clk(gclk));
	jdff dff_A_TyYdHk1b8_0(.dout(w_dff_A_VLo057qZ4_0),.din(w_dff_A_TyYdHk1b8_0),.clk(gclk));
	jdff dff_A_OnKm0gGs9_0(.dout(w_dff_A_TyYdHk1b8_0),.din(w_dff_A_OnKm0gGs9_0),.clk(gclk));
	jdff dff_A_kfRW8fpl9_0(.dout(w_dff_A_OnKm0gGs9_0),.din(w_dff_A_kfRW8fpl9_0),.clk(gclk));
	jdff dff_A_1DgrQCxR4_1(.dout(w_G953_0[1]),.din(w_dff_A_1DgrQCxR4_1),.clk(gclk));
	jdff dff_A_QPs4KyXP2_1(.dout(w_dff_A_1DgrQCxR4_1),.din(w_dff_A_QPs4KyXP2_1),.clk(gclk));
	jdff dff_A_ItqCFU3O9_1(.dout(w_dff_A_QPs4KyXP2_1),.din(w_dff_A_ItqCFU3O9_1),.clk(gclk));
	jdff dff_A_uLPdK8m11_1(.dout(w_dff_A_ItqCFU3O9_1),.din(w_dff_A_uLPdK8m11_1),.clk(gclk));
	jdff dff_A_sj9vVAaV6_1(.dout(w_dff_A_uLPdK8m11_1),.din(w_dff_A_sj9vVAaV6_1),.clk(gclk));
	jdff dff_A_c9chWVhq5_1(.dout(w_dff_A_sj9vVAaV6_1),.din(w_dff_A_c9chWVhq5_1),.clk(gclk));
	jdff dff_A_eWvczxoQ7_1(.dout(w_dff_A_c9chWVhq5_1),.din(w_dff_A_eWvczxoQ7_1),.clk(gclk));
	jdff dff_A_NzHc1JiS4_1(.dout(w_dff_A_eWvczxoQ7_1),.din(w_dff_A_NzHc1JiS4_1),.clk(gclk));
	jdff dff_A_5CQyyH1w0_1(.dout(w_dff_A_NzHc1JiS4_1),.din(w_dff_A_5CQyyH1w0_1),.clk(gclk));
	jdff dff_A_t9EyqNw49_1(.dout(w_dff_A_5CQyyH1w0_1),.din(w_dff_A_t9EyqNw49_1),.clk(gclk));
	jdff dff_A_HKSalTAP3_1(.dout(w_dff_A_t9EyqNw49_1),.din(w_dff_A_HKSalTAP3_1),.clk(gclk));
	jdff dff_A_CpSt5fEB7_1(.dout(w_dff_A_HKSalTAP3_1),.din(w_dff_A_CpSt5fEB7_1),.clk(gclk));
	jdff dff_A_17b44fcI5_1(.dout(w_dff_A_CpSt5fEB7_1),.din(w_dff_A_17b44fcI5_1),.clk(gclk));
	jdff dff_A_8BXKGvxZ3_1(.dout(w_dff_A_17b44fcI5_1),.din(w_dff_A_8BXKGvxZ3_1),.clk(gclk));
	jdff dff_A_NfEoZtfz9_1(.dout(w_dff_A_8BXKGvxZ3_1),.din(w_dff_A_NfEoZtfz9_1),.clk(gclk));
	jdff dff_A_aJrrWy2t9_2(.dout(w_G953_0[2]),.din(w_dff_A_aJrrWy2t9_2),.clk(gclk));
	jdff dff_A_aypXjXkt3_2(.dout(w_dff_A_aJrrWy2t9_2),.din(w_dff_A_aypXjXkt3_2),.clk(gclk));
	jdff dff_A_PNIcb18Q8_2(.dout(w_dff_A_aypXjXkt3_2),.din(w_dff_A_PNIcb18Q8_2),.clk(gclk));
	jdff dff_A_OHQTwM1G8_2(.dout(w_dff_A_PNIcb18Q8_2),.din(w_dff_A_OHQTwM1G8_2),.clk(gclk));
	jdff dff_A_KHcooSNk5_2(.dout(w_dff_A_OHQTwM1G8_2),.din(w_dff_A_KHcooSNk5_2),.clk(gclk));
	jdff dff_A_4ckL2wm82_2(.dout(w_dff_A_KHcooSNk5_2),.din(w_dff_A_4ckL2wm82_2),.clk(gclk));
	jdff dff_A_sgmh0wWz7_2(.dout(w_dff_A_4ckL2wm82_2),.din(w_dff_A_sgmh0wWz7_2),.clk(gclk));
	jdff dff_A_NwLwOxON9_2(.dout(w_dff_A_sgmh0wWz7_2),.din(w_dff_A_NwLwOxON9_2),.clk(gclk));
	jdff dff_A_1IFijKqr5_2(.dout(w_dff_A_NwLwOxON9_2),.din(w_dff_A_1IFijKqr5_2),.clk(gclk));
	jdff dff_A_Dr0R36Qq2_2(.dout(w_dff_A_1IFijKqr5_2),.din(w_dff_A_Dr0R36Qq2_2),.clk(gclk));
	jdff dff_A_FAXEgT0e3_2(.dout(w_dff_A_Dr0R36Qq2_2),.din(w_dff_A_FAXEgT0e3_2),.clk(gclk));
	jdff dff_A_3VXP8UtH9_2(.dout(w_dff_A_FAXEgT0e3_2),.din(w_dff_A_3VXP8UtH9_2),.clk(gclk));
	jdff dff_A_PqbbI6gb8_2(.dout(w_dff_A_3VXP8UtH9_2),.din(w_dff_A_PqbbI6gb8_2),.clk(gclk));
	jdff dff_A_BnXwzpHc0_2(.dout(w_dff_A_PqbbI6gb8_2),.din(w_dff_A_BnXwzpHc0_2),.clk(gclk));
	jdff dff_A_MewQL7980_2(.dout(w_dff_A_BnXwzpHc0_2),.din(w_dff_A_MewQL7980_2),.clk(gclk));
	jdff dff_A_jtdazSx98_1(.dout(w_G210_0[1]),.din(w_dff_A_jtdazSx98_1),.clk(gclk));
	jdff dff_A_32dO2mgZ8_0(.dout(w_G101_0[0]),.din(w_dff_A_32dO2mgZ8_0),.clk(gclk));
	jdff dff_A_y6vKYzLK4_0(.dout(w_dff_A_32dO2mgZ8_0),.din(w_dff_A_y6vKYzLK4_0),.clk(gclk));
	jdff dff_A_nSLHMqQ46_0(.dout(w_dff_A_y6vKYzLK4_0),.din(w_dff_A_nSLHMqQ46_0),.clk(gclk));
	jdff dff_A_q1UogLyh4_0(.dout(w_dff_A_nSLHMqQ46_0),.din(w_dff_A_q1UogLyh4_0),.clk(gclk));
	jdff dff_A_z87XFPGG2_0(.dout(w_dff_A_q1UogLyh4_0),.din(w_dff_A_z87XFPGG2_0),.clk(gclk));
	jdff dff_A_I9lUJXPJ2_0(.dout(w_dff_A_z87XFPGG2_0),.din(w_dff_A_I9lUJXPJ2_0),.clk(gclk));
	jdff dff_A_tkXz10Lf5_0(.dout(w_dff_A_I9lUJXPJ2_0),.din(w_dff_A_tkXz10Lf5_0),.clk(gclk));
	jdff dff_A_eVRXWvqv9_0(.dout(w_dff_A_tkXz10Lf5_0),.din(w_dff_A_eVRXWvqv9_0),.clk(gclk));
	jdff dff_A_YqIhGlMJ0_0(.dout(w_dff_A_eVRXWvqv9_0),.din(w_dff_A_YqIhGlMJ0_0),.clk(gclk));
	jdff dff_A_7FVeCVei6_0(.dout(w_dff_A_YqIhGlMJ0_0),.din(w_dff_A_7FVeCVei6_0),.clk(gclk));
	jdff dff_A_fjjRkyM94_0(.dout(w_dff_A_7FVeCVei6_0),.din(w_dff_A_fjjRkyM94_0),.clk(gclk));
	jdff dff_A_xokxmThT8_2(.dout(w_G101_0[2]),.din(w_dff_A_xokxmThT8_2),.clk(gclk));
	jdff dff_B_nhW2gutN0_3(.din(G101),.dout(w_dff_B_nhW2gutN0_3),.clk(gclk));
	jdff dff_A_zw6Yoo2x9_1(.dout(w_n84_0[1]),.din(w_dff_A_zw6Yoo2x9_1),.clk(gclk));
	jdff dff_A_QYrbG5kf3_0(.dout(w_G119_0[0]),.din(w_dff_A_QYrbG5kf3_0),.clk(gclk));
	jdff dff_A_g1ggyjHE6_0(.dout(w_dff_A_QYrbG5kf3_0),.din(w_dff_A_g1ggyjHE6_0),.clk(gclk));
	jdff dff_A_qlAwMW466_0(.dout(w_dff_A_g1ggyjHE6_0),.din(w_dff_A_qlAwMW466_0),.clk(gclk));
	jdff dff_A_uoLsdpJJ8_0(.dout(w_dff_A_qlAwMW466_0),.din(w_dff_A_uoLsdpJJ8_0),.clk(gclk));
	jdff dff_A_TLRcHvBK0_0(.dout(w_dff_A_uoLsdpJJ8_0),.din(w_dff_A_TLRcHvBK0_0),.clk(gclk));
	jdff dff_A_G3SHcqRu0_0(.dout(w_dff_A_TLRcHvBK0_0),.din(w_dff_A_G3SHcqRu0_0),.clk(gclk));
	jdff dff_A_F5vqeNN54_0(.dout(w_dff_A_G3SHcqRu0_0),.din(w_dff_A_F5vqeNN54_0),.clk(gclk));
	jdff dff_A_4QrWqADd8_0(.dout(w_dff_A_F5vqeNN54_0),.din(w_dff_A_4QrWqADd8_0),.clk(gclk));
	jdff dff_A_HqrT7uBB3_0(.dout(w_dff_A_4QrWqADd8_0),.din(w_dff_A_HqrT7uBB3_0),.clk(gclk));
	jdff dff_A_uqjWhDGs4_0(.dout(w_dff_A_HqrT7uBB3_0),.din(w_dff_A_uqjWhDGs4_0),.clk(gclk));
	jdff dff_A_rEvntC530_0(.dout(w_dff_A_uqjWhDGs4_0),.din(w_dff_A_rEvntC530_0),.clk(gclk));
	jdff dff_A_kWji1Z9g6_0(.dout(w_dff_A_rEvntC530_0),.din(w_dff_A_kWji1Z9g6_0),.clk(gclk));
	jdff dff_A_ixzV3uN88_0(.dout(w_G116_0[0]),.din(w_dff_A_ixzV3uN88_0),.clk(gclk));
	jdff dff_A_7QMqde7C1_0(.dout(w_dff_A_ixzV3uN88_0),.din(w_dff_A_7QMqde7C1_0),.clk(gclk));
	jdff dff_A_fTN0M8Nl9_0(.dout(w_dff_A_7QMqde7C1_0),.din(w_dff_A_fTN0M8Nl9_0),.clk(gclk));
	jdff dff_A_Xvs9Klv14_0(.dout(w_dff_A_fTN0M8Nl9_0),.din(w_dff_A_Xvs9Klv14_0),.clk(gclk));
	jdff dff_A_kYAyEiQQ5_0(.dout(w_dff_A_Xvs9Klv14_0),.din(w_dff_A_kYAyEiQQ5_0),.clk(gclk));
	jdff dff_A_E4mlpWHo2_0(.dout(w_dff_A_kYAyEiQQ5_0),.din(w_dff_A_E4mlpWHo2_0),.clk(gclk));
	jdff dff_A_hlClqw9d9_0(.dout(w_dff_A_E4mlpWHo2_0),.din(w_dff_A_hlClqw9d9_0),.clk(gclk));
	jdff dff_A_NKLr0QsT4_0(.dout(w_dff_A_hlClqw9d9_0),.din(w_dff_A_NKLr0QsT4_0),.clk(gclk));
	jdff dff_A_9lrOEVyf1_0(.dout(w_dff_A_NKLr0QsT4_0),.din(w_dff_A_9lrOEVyf1_0),.clk(gclk));
	jdff dff_A_1jlZLf9J6_0(.dout(w_dff_A_9lrOEVyf1_0),.din(w_dff_A_1jlZLf9J6_0),.clk(gclk));
	jdff dff_A_UbfACKGM5_0(.dout(w_dff_A_1jlZLf9J6_0),.din(w_dff_A_UbfACKGM5_0),.clk(gclk));
	jdff dff_A_AQxkgjvZ4_0(.dout(w_dff_A_UbfACKGM5_0),.din(w_dff_A_AQxkgjvZ4_0),.clk(gclk));
	jdff dff_A_vFPHv5Kn6_0(.dout(w_G113_0[0]),.din(w_dff_A_vFPHv5Kn6_0),.clk(gclk));
	jdff dff_A_5uLjVev71_0(.dout(w_dff_A_vFPHv5Kn6_0),.din(w_dff_A_5uLjVev71_0),.clk(gclk));
	jdff dff_A_mhvx7r855_0(.dout(w_dff_A_5uLjVev71_0),.din(w_dff_A_mhvx7r855_0),.clk(gclk));
	jdff dff_A_RNYdsNw95_0(.dout(w_dff_A_mhvx7r855_0),.din(w_dff_A_RNYdsNw95_0),.clk(gclk));
	jdff dff_A_LqK2UbH56_0(.dout(w_dff_A_RNYdsNw95_0),.din(w_dff_A_LqK2UbH56_0),.clk(gclk));
	jdff dff_A_Z7vQxSIJ0_0(.dout(w_dff_A_LqK2UbH56_0),.din(w_dff_A_Z7vQxSIJ0_0),.clk(gclk));
	jdff dff_A_ge88EaDK2_0(.dout(w_dff_A_Z7vQxSIJ0_0),.din(w_dff_A_ge88EaDK2_0),.clk(gclk));
	jdff dff_A_MGD9JNrL1_0(.dout(w_dff_A_ge88EaDK2_0),.din(w_dff_A_MGD9JNrL1_0),.clk(gclk));
	jdff dff_A_tNRargS47_0(.dout(w_dff_A_MGD9JNrL1_0),.din(w_dff_A_tNRargS47_0),.clk(gclk));
	jdff dff_A_YZHVwf6Q8_0(.dout(w_dff_A_tNRargS47_0),.din(w_dff_A_YZHVwf6Q8_0),.clk(gclk));
	jdff dff_A_wW6jRfOH3_0(.dout(w_dff_A_YZHVwf6Q8_0),.din(w_dff_A_wW6jRfOH3_0),.clk(gclk));
	jdff dff_A_uGUkLdGk8_0(.dout(w_dff_A_wW6jRfOH3_0),.din(w_dff_A_uGUkLdGk8_0),.clk(gclk));
	jdff dff_B_rrIwJGG22_1(.din(n76),.dout(w_dff_B_rrIwJGG22_1),.clk(gclk));
	jdff dff_A_QFbJyn4L1_0(.dout(w_G146_0[0]),.din(w_dff_A_QFbJyn4L1_0),.clk(gclk));
	jdff dff_A_XUxXPWpj3_0(.dout(w_dff_A_QFbJyn4L1_0),.din(w_dff_A_XUxXPWpj3_0),.clk(gclk));
	jdff dff_A_3GdzA8GT8_0(.dout(w_dff_A_XUxXPWpj3_0),.din(w_dff_A_3GdzA8GT8_0),.clk(gclk));
	jdff dff_A_qyhQuvCh2_0(.dout(w_dff_A_3GdzA8GT8_0),.din(w_dff_A_qyhQuvCh2_0),.clk(gclk));
	jdff dff_A_kP1S94qw3_0(.dout(w_dff_A_qyhQuvCh2_0),.din(w_dff_A_kP1S94qw3_0),.clk(gclk));
	jdff dff_A_np2tc0dK7_0(.dout(w_dff_A_kP1S94qw3_0),.din(w_dff_A_np2tc0dK7_0),.clk(gclk));
	jdff dff_A_bcKuHTcd4_0(.dout(w_dff_A_np2tc0dK7_0),.din(w_dff_A_bcKuHTcd4_0),.clk(gclk));
	jdff dff_A_ch50iC326_0(.dout(w_dff_A_bcKuHTcd4_0),.din(w_dff_A_ch50iC326_0),.clk(gclk));
	jdff dff_A_7pcJFWUh4_0(.dout(w_dff_A_ch50iC326_0),.din(w_dff_A_7pcJFWUh4_0),.clk(gclk));
	jdff dff_A_C0Oae3SM7_0(.dout(w_dff_A_7pcJFWUh4_0),.din(w_dff_A_C0Oae3SM7_0),.clk(gclk));
	jdff dff_A_nil8ntDj1_0(.dout(w_dff_A_C0Oae3SM7_0),.din(w_dff_A_nil8ntDj1_0),.clk(gclk));
	jdff dff_A_Ooj9orFX9_0(.dout(w_dff_A_nil8ntDj1_0),.din(w_dff_A_Ooj9orFX9_0),.clk(gclk));
	jdff dff_A_iwuOnkwX7_1(.dout(w_G143_0[1]),.din(w_dff_A_iwuOnkwX7_1),.clk(gclk));
	jdff dff_A_V2GnYsRI4_1(.dout(w_dff_A_iwuOnkwX7_1),.din(w_dff_A_V2GnYsRI4_1),.clk(gclk));
	jdff dff_A_4NJCaWES2_1(.dout(w_dff_A_V2GnYsRI4_1),.din(w_dff_A_4NJCaWES2_1),.clk(gclk));
	jdff dff_A_CZgREzlJ7_1(.dout(w_dff_A_4NJCaWES2_1),.din(w_dff_A_CZgREzlJ7_1),.clk(gclk));
	jdff dff_A_qtqbA7TE2_1(.dout(w_dff_A_CZgREzlJ7_1),.din(w_dff_A_qtqbA7TE2_1),.clk(gclk));
	jdff dff_A_xjC3xC1f3_1(.dout(w_dff_A_qtqbA7TE2_1),.din(w_dff_A_xjC3xC1f3_1),.clk(gclk));
	jdff dff_A_gjJLpUjO2_1(.dout(w_dff_A_xjC3xC1f3_1),.din(w_dff_A_gjJLpUjO2_1),.clk(gclk));
	jdff dff_A_0FBt5On70_1(.dout(w_dff_A_gjJLpUjO2_1),.din(w_dff_A_0FBt5On70_1),.clk(gclk));
	jdff dff_A_RiPSRki43_1(.dout(w_dff_A_0FBt5On70_1),.din(w_dff_A_RiPSRki43_1),.clk(gclk));
	jdff dff_A_iOJCDytV9_1(.dout(w_dff_A_RiPSRki43_1),.din(w_dff_A_iOJCDytV9_1),.clk(gclk));
	jdff dff_A_PtVCZn1s7_1(.dout(w_dff_A_iOJCDytV9_1),.din(w_dff_A_PtVCZn1s7_1),.clk(gclk));
	jdff dff_A_KvChh7Xe5_1(.dout(w_dff_A_PtVCZn1s7_1),.din(w_dff_A_KvChh7Xe5_1),.clk(gclk));
	jdff dff_A_tAIPdC814_2(.dout(w_G143_0[2]),.din(w_dff_A_tAIPdC814_2),.clk(gclk));
	jdff dff_A_uPQtcYLi3_0(.dout(w_G128_1[0]),.din(w_dff_A_uPQtcYLi3_0),.clk(gclk));
	jdff dff_A_8dGNuAjS6_1(.dout(w_G128_0[1]),.din(w_dff_A_8dGNuAjS6_1),.clk(gclk));
	jdff dff_A_SKEkCR5y1_1(.dout(w_dff_A_8dGNuAjS6_1),.din(w_dff_A_SKEkCR5y1_1),.clk(gclk));
	jdff dff_A_bAvRgBrY7_1(.dout(w_dff_A_SKEkCR5y1_1),.din(w_dff_A_bAvRgBrY7_1),.clk(gclk));
	jdff dff_A_4a5ZjSeF2_1(.dout(w_dff_A_bAvRgBrY7_1),.din(w_dff_A_4a5ZjSeF2_1),.clk(gclk));
	jdff dff_A_ML9fB5ek4_1(.dout(w_dff_A_4a5ZjSeF2_1),.din(w_dff_A_ML9fB5ek4_1),.clk(gclk));
	jdff dff_A_pasSz2kO4_1(.dout(w_dff_A_ML9fB5ek4_1),.din(w_dff_A_pasSz2kO4_1),.clk(gclk));
	jdff dff_A_HJTlownT6_1(.dout(w_dff_A_pasSz2kO4_1),.din(w_dff_A_HJTlownT6_1),.clk(gclk));
	jdff dff_A_ZbpgyP838_1(.dout(w_dff_A_HJTlownT6_1),.din(w_dff_A_ZbpgyP838_1),.clk(gclk));
	jdff dff_A_f9Epro6U8_1(.dout(w_dff_A_ZbpgyP838_1),.din(w_dff_A_f9Epro6U8_1),.clk(gclk));
	jdff dff_A_AaxeuSG62_1(.dout(w_dff_A_f9Epro6U8_1),.din(w_dff_A_AaxeuSG62_1),.clk(gclk));
	jdff dff_A_j6eTlFGV7_1(.dout(w_dff_A_AaxeuSG62_1),.din(w_dff_A_j6eTlFGV7_1),.clk(gclk));
	jdff dff_A_TOF1ISug0_1(.dout(w_dff_A_j6eTlFGV7_1),.din(w_dff_A_TOF1ISug0_1),.clk(gclk));
	jdff dff_A_wOV34ZYg8_1(.dout(w_n77_0[1]),.din(w_dff_A_wOV34ZYg8_1),.clk(gclk));
	jdff dff_A_mQkGIWB23_0(.dout(w_G131_0[0]),.din(w_dff_A_mQkGIWB23_0),.clk(gclk));
	jdff dff_A_zXIWKv336_0(.dout(w_dff_A_mQkGIWB23_0),.din(w_dff_A_zXIWKv336_0),.clk(gclk));
	jdff dff_A_HiXB6ErV1_0(.dout(w_dff_A_zXIWKv336_0),.din(w_dff_A_HiXB6ErV1_0),.clk(gclk));
	jdff dff_A_OiKv6x1P3_0(.dout(w_dff_A_HiXB6ErV1_0),.din(w_dff_A_OiKv6x1P3_0),.clk(gclk));
	jdff dff_A_MatWtpgi3_0(.dout(w_dff_A_OiKv6x1P3_0),.din(w_dff_A_MatWtpgi3_0),.clk(gclk));
	jdff dff_A_oQ8MpKlk1_0(.dout(w_dff_A_MatWtpgi3_0),.din(w_dff_A_oQ8MpKlk1_0),.clk(gclk));
	jdff dff_A_VxZaGK1w3_0(.dout(w_dff_A_oQ8MpKlk1_0),.din(w_dff_A_VxZaGK1w3_0),.clk(gclk));
	jdff dff_A_9EuIiA1r1_0(.dout(w_dff_A_VxZaGK1w3_0),.din(w_dff_A_9EuIiA1r1_0),.clk(gclk));
	jdff dff_A_1MXo40gh8_0(.dout(w_dff_A_9EuIiA1r1_0),.din(w_dff_A_1MXo40gh8_0),.clk(gclk));
	jdff dff_A_UsCn5THH1_0(.dout(w_dff_A_1MXo40gh8_0),.din(w_dff_A_UsCn5THH1_0),.clk(gclk));
	jdff dff_A_hApYUv2t3_0(.dout(w_dff_A_UsCn5THH1_0),.din(w_dff_A_hApYUv2t3_0),.clk(gclk));
	jdff dff_A_3crr4E687_0(.dout(w_dff_A_hApYUv2t3_0),.din(w_dff_A_3crr4E687_0),.clk(gclk));
	jdff dff_A_TKgBSNOc3_0(.dout(w_G137_0[0]),.din(w_dff_A_TKgBSNOc3_0),.clk(gclk));
	jdff dff_A_GtPlbU3g8_0(.dout(w_dff_A_TKgBSNOc3_0),.din(w_dff_A_GtPlbU3g8_0),.clk(gclk));
	jdff dff_A_6wgcFCk43_0(.dout(w_dff_A_GtPlbU3g8_0),.din(w_dff_A_6wgcFCk43_0),.clk(gclk));
	jdff dff_A_p1WLYOiw3_0(.dout(w_dff_A_6wgcFCk43_0),.din(w_dff_A_p1WLYOiw3_0),.clk(gclk));
	jdff dff_A_rEzsa2tP4_0(.dout(w_dff_A_p1WLYOiw3_0),.din(w_dff_A_rEzsa2tP4_0),.clk(gclk));
	jdff dff_A_A7GFZBeo0_0(.dout(w_dff_A_rEzsa2tP4_0),.din(w_dff_A_A7GFZBeo0_0),.clk(gclk));
	jdff dff_A_hvHGuKJ83_0(.dout(w_dff_A_A7GFZBeo0_0),.din(w_dff_A_hvHGuKJ83_0),.clk(gclk));
	jdff dff_A_9nhakWyN2_0(.dout(w_dff_A_hvHGuKJ83_0),.din(w_dff_A_9nhakWyN2_0),.clk(gclk));
	jdff dff_A_WZ3AznBH3_0(.dout(w_dff_A_9nhakWyN2_0),.din(w_dff_A_WZ3AznBH3_0),.clk(gclk));
	jdff dff_A_VkgiVfXZ7_0(.dout(w_dff_A_WZ3AznBH3_0),.din(w_dff_A_VkgiVfXZ7_0),.clk(gclk));
	jdff dff_A_kaFOH6IU9_0(.dout(w_dff_A_VkgiVfXZ7_0),.din(w_dff_A_kaFOH6IU9_0),.clk(gclk));
	jdff dff_A_gwoGQgPo3_2(.dout(w_G137_0[2]),.din(w_dff_A_gwoGQgPo3_2),.clk(gclk));
	jdff dff_A_0jUAIR0N0_2(.dout(w_dff_A_gwoGQgPo3_2),.din(w_dff_A_0jUAIR0N0_2),.clk(gclk));
	jdff dff_B_TYwom6MH1_3(.din(G137),.dout(w_dff_B_TYwom6MH1_3),.clk(gclk));
	jdff dff_A_Hk3nXfqo8_0(.dout(w_G134_0[0]),.din(w_dff_A_Hk3nXfqo8_0),.clk(gclk));
	jdff dff_A_BmZUYzin4_0(.dout(w_dff_A_Hk3nXfqo8_0),.din(w_dff_A_BmZUYzin4_0),.clk(gclk));
	jdff dff_A_b5eJjfJ28_0(.dout(w_dff_A_BmZUYzin4_0),.din(w_dff_A_b5eJjfJ28_0),.clk(gclk));
	jdff dff_A_CrhC5AA46_0(.dout(w_dff_A_b5eJjfJ28_0),.din(w_dff_A_CrhC5AA46_0),.clk(gclk));
	jdff dff_A_4qiJJOE21_0(.dout(w_dff_A_CrhC5AA46_0),.din(w_dff_A_4qiJJOE21_0),.clk(gclk));
	jdff dff_A_sSivf5sT5_0(.dout(w_dff_A_4qiJJOE21_0),.din(w_dff_A_sSivf5sT5_0),.clk(gclk));
	jdff dff_A_Ji5K9ZSn0_0(.dout(w_dff_A_sSivf5sT5_0),.din(w_dff_A_Ji5K9ZSn0_0),.clk(gclk));
	jdff dff_A_1bPf2LbR7_0(.dout(w_dff_A_Ji5K9ZSn0_0),.din(w_dff_A_1bPf2LbR7_0),.clk(gclk));
	jdff dff_A_j27VBrhb1_0(.dout(w_dff_A_1bPf2LbR7_0),.din(w_dff_A_j27VBrhb1_0),.clk(gclk));
	jdff dff_A_Pr4o3CpU3_0(.dout(w_dff_A_j27VBrhb1_0),.din(w_dff_A_Pr4o3CpU3_0),.clk(gclk));
	jdff dff_A_AwtVxnWA7_0(.dout(w_dff_A_Pr4o3CpU3_0),.din(w_dff_A_AwtVxnWA7_0),.clk(gclk));
	jdff dff_A_etucNoNa4_0(.dout(w_dff_A_AwtVxnWA7_0),.din(w_dff_A_etucNoNa4_0),.clk(gclk));
	jdff dff_A_tgsGGwUG3_2(.dout(w_dff_A_Jo05WalF4_0),.din(w_dff_A_tgsGGwUG3_2),.clk(gclk));
	jdff dff_A_Jo05WalF4_0(.dout(w_dff_A_lQQ7OrNU9_0),.din(w_dff_A_Jo05WalF4_0),.clk(gclk));
	jdff dff_A_lQQ7OrNU9_0(.dout(w_dff_A_Oo8xOv4Z2_0),.din(w_dff_A_lQQ7OrNU9_0),.clk(gclk));
	jdff dff_A_Oo8xOv4Z2_0(.dout(w_dff_A_1yTGniJ24_0),.din(w_dff_A_Oo8xOv4Z2_0),.clk(gclk));
	jdff dff_A_1yTGniJ24_0(.dout(w_dff_A_9CGrs0b87_0),.din(w_dff_A_1yTGniJ24_0),.clk(gclk));
	jdff dff_A_9CGrs0b87_0(.dout(w_dff_A_irGhth8U4_0),.din(w_dff_A_9CGrs0b87_0),.clk(gclk));
	jdff dff_A_irGhth8U4_0(.dout(G3),.din(w_dff_A_irGhth8U4_0),.clk(gclk));
	jdff dff_A_1jvHz01S6_2(.dout(w_dff_A_h6B22lMB2_0),.din(w_dff_A_1jvHz01S6_2),.clk(gclk));
	jdff dff_A_h6B22lMB2_0(.dout(w_dff_A_FLxDXH7i7_0),.din(w_dff_A_h6B22lMB2_0),.clk(gclk));
	jdff dff_A_FLxDXH7i7_0(.dout(w_dff_A_fcLWlC2l7_0),.din(w_dff_A_FLxDXH7i7_0),.clk(gclk));
	jdff dff_A_fcLWlC2l7_0(.dout(w_dff_A_3MEcD3C63_0),.din(w_dff_A_fcLWlC2l7_0),.clk(gclk));
	jdff dff_A_3MEcD3C63_0(.dout(w_dff_A_PpPLHoD77_0),.din(w_dff_A_3MEcD3C63_0),.clk(gclk));
	jdff dff_A_PpPLHoD77_0(.dout(w_dff_A_NWx4ToN48_0),.din(w_dff_A_PpPLHoD77_0),.clk(gclk));
	jdff dff_A_NWx4ToN48_0(.dout(G6),.din(w_dff_A_NWx4ToN48_0),.clk(gclk));
	jdff dff_A_B8eR28a40_2(.dout(w_dff_A_yM9yP70s3_0),.din(w_dff_A_B8eR28a40_2),.clk(gclk));
	jdff dff_A_yM9yP70s3_0(.dout(w_dff_A_AOZGbwPt8_0),.din(w_dff_A_yM9yP70s3_0),.clk(gclk));
	jdff dff_A_AOZGbwPt8_0(.dout(w_dff_A_3aZ33zEw3_0),.din(w_dff_A_AOZGbwPt8_0),.clk(gclk));
	jdff dff_A_3aZ33zEw3_0(.dout(w_dff_A_STmyObGg3_0),.din(w_dff_A_3aZ33zEw3_0),.clk(gclk));
	jdff dff_A_STmyObGg3_0(.dout(w_dff_A_5zyebfVW4_0),.din(w_dff_A_STmyObGg3_0),.clk(gclk));
	jdff dff_A_5zyebfVW4_0(.dout(w_dff_A_y16Uu0qQ7_0),.din(w_dff_A_5zyebfVW4_0),.clk(gclk));
	jdff dff_A_y16Uu0qQ7_0(.dout(G9),.din(w_dff_A_y16Uu0qQ7_0),.clk(gclk));
	jdff dff_A_0f7i80Nd1_2(.dout(w_dff_A_R4yd7DBk4_0),.din(w_dff_A_0f7i80Nd1_2),.clk(gclk));
	jdff dff_A_R4yd7DBk4_0(.dout(w_dff_A_FcBOieOs8_0),.din(w_dff_A_R4yd7DBk4_0),.clk(gclk));
	jdff dff_A_FcBOieOs8_0(.dout(w_dff_A_pLYsoq2Q2_0),.din(w_dff_A_FcBOieOs8_0),.clk(gclk));
	jdff dff_A_pLYsoq2Q2_0(.dout(w_dff_A_scRGQsfY4_0),.din(w_dff_A_pLYsoq2Q2_0),.clk(gclk));
	jdff dff_A_scRGQsfY4_0(.dout(w_dff_A_SOBVLc7F8_0),.din(w_dff_A_scRGQsfY4_0),.clk(gclk));
	jdff dff_A_SOBVLc7F8_0(.dout(w_dff_A_ZfoTHkX01_0),.din(w_dff_A_SOBVLc7F8_0),.clk(gclk));
	jdff dff_A_ZfoTHkX01_0(.dout(G12),.din(w_dff_A_ZfoTHkX01_0),.clk(gclk));
	jdff dff_A_3yefOgGp2_2(.dout(w_dff_A_QjzFVJyZ8_0),.din(w_dff_A_3yefOgGp2_2),.clk(gclk));
	jdff dff_A_QjzFVJyZ8_0(.dout(w_dff_A_9cQjYvRQ1_0),.din(w_dff_A_QjzFVJyZ8_0),.clk(gclk));
	jdff dff_A_9cQjYvRQ1_0(.dout(w_dff_A_U4KfyalL5_0),.din(w_dff_A_9cQjYvRQ1_0),.clk(gclk));
	jdff dff_A_U4KfyalL5_0(.dout(w_dff_A_AY5bFrSp1_0),.din(w_dff_A_U4KfyalL5_0),.clk(gclk));
	jdff dff_A_AY5bFrSp1_0(.dout(w_dff_A_ASjJGAdI0_0),.din(w_dff_A_AY5bFrSp1_0),.clk(gclk));
	jdff dff_A_ASjJGAdI0_0(.dout(w_dff_A_ijmCbDwn1_0),.din(w_dff_A_ASjJGAdI0_0),.clk(gclk));
	jdff dff_A_ijmCbDwn1_0(.dout(G30),.din(w_dff_A_ijmCbDwn1_0),.clk(gclk));
	jdff dff_A_ehYWmLY91_2(.dout(w_dff_A_IaTZkgip1_0),.din(w_dff_A_ehYWmLY91_2),.clk(gclk));
	jdff dff_A_IaTZkgip1_0(.dout(w_dff_A_QLAX8zKf4_0),.din(w_dff_A_IaTZkgip1_0),.clk(gclk));
	jdff dff_A_QLAX8zKf4_0(.dout(w_dff_A_CkySIeNS0_0),.din(w_dff_A_QLAX8zKf4_0),.clk(gclk));
	jdff dff_A_CkySIeNS0_0(.dout(w_dff_A_ukcVafbV1_0),.din(w_dff_A_CkySIeNS0_0),.clk(gclk));
	jdff dff_A_ukcVafbV1_0(.dout(w_dff_A_u7j7UB2c4_0),.din(w_dff_A_ukcVafbV1_0),.clk(gclk));
	jdff dff_A_u7j7UB2c4_0(.dout(w_dff_A_AYMvHAtF2_0),.din(w_dff_A_u7j7UB2c4_0),.clk(gclk));
	jdff dff_A_AYMvHAtF2_0(.dout(G45),.din(w_dff_A_AYMvHAtF2_0),.clk(gclk));
	jdff dff_A_CxV5R3S41_2(.dout(w_dff_A_lByYvY8H8_0),.din(w_dff_A_CxV5R3S41_2),.clk(gclk));
	jdff dff_A_lByYvY8H8_0(.dout(w_dff_A_D67fBNeB0_0),.din(w_dff_A_lByYvY8H8_0),.clk(gclk));
	jdff dff_A_D67fBNeB0_0(.dout(w_dff_A_BfppoD9q8_0),.din(w_dff_A_D67fBNeB0_0),.clk(gclk));
	jdff dff_A_BfppoD9q8_0(.dout(w_dff_A_vt6MVxkA5_0),.din(w_dff_A_BfppoD9q8_0),.clk(gclk));
	jdff dff_A_vt6MVxkA5_0(.dout(w_dff_A_WlEz4kmI8_0),.din(w_dff_A_vt6MVxkA5_0),.clk(gclk));
	jdff dff_A_WlEz4kmI8_0(.dout(w_dff_A_pHmFZTGV1_0),.din(w_dff_A_WlEz4kmI8_0),.clk(gclk));
	jdff dff_A_pHmFZTGV1_0(.dout(G48),.din(w_dff_A_pHmFZTGV1_0),.clk(gclk));
	jdff dff_A_iA9pP22X1_2(.dout(w_dff_A_IExpIc7W2_0),.din(w_dff_A_iA9pP22X1_2),.clk(gclk));
	jdff dff_A_IExpIc7W2_0(.dout(w_dff_A_sFpjpHVR7_0),.din(w_dff_A_IExpIc7W2_0),.clk(gclk));
	jdff dff_A_sFpjpHVR7_0(.dout(w_dff_A_Ly8Z3pCD4_0),.din(w_dff_A_sFpjpHVR7_0),.clk(gclk));
	jdff dff_A_Ly8Z3pCD4_0(.dout(w_dff_A_hi7LkfJQ5_0),.din(w_dff_A_Ly8Z3pCD4_0),.clk(gclk));
	jdff dff_A_hi7LkfJQ5_0(.dout(w_dff_A_68iq09Iz0_0),.din(w_dff_A_hi7LkfJQ5_0),.clk(gclk));
	jdff dff_A_68iq09Iz0_0(.dout(w_dff_A_h4SaEFY61_0),.din(w_dff_A_68iq09Iz0_0),.clk(gclk));
	jdff dff_A_h4SaEFY61_0(.dout(G15),.din(w_dff_A_h4SaEFY61_0),.clk(gclk));
	jdff dff_A_OvTispEG5_2(.dout(w_dff_A_x7HgaYxP9_0),.din(w_dff_A_OvTispEG5_2),.clk(gclk));
	jdff dff_A_x7HgaYxP9_0(.dout(w_dff_A_d0NGJUAT7_0),.din(w_dff_A_x7HgaYxP9_0),.clk(gclk));
	jdff dff_A_d0NGJUAT7_0(.dout(w_dff_A_TrxtfwNt8_0),.din(w_dff_A_d0NGJUAT7_0),.clk(gclk));
	jdff dff_A_TrxtfwNt8_0(.dout(w_dff_A_Tu2aKiaE8_0),.din(w_dff_A_TrxtfwNt8_0),.clk(gclk));
	jdff dff_A_Tu2aKiaE8_0(.dout(w_dff_A_8joY4mYZ5_0),.din(w_dff_A_Tu2aKiaE8_0),.clk(gclk));
	jdff dff_A_8joY4mYZ5_0(.dout(w_dff_A_JJWlIZNC0_0),.din(w_dff_A_8joY4mYZ5_0),.clk(gclk));
	jdff dff_A_JJWlIZNC0_0(.dout(G18),.din(w_dff_A_JJWlIZNC0_0),.clk(gclk));
	jdff dff_A_Fko9CuZr6_2(.dout(w_dff_A_2jZUzQMO3_0),.din(w_dff_A_Fko9CuZr6_2),.clk(gclk));
	jdff dff_A_2jZUzQMO3_0(.dout(w_dff_A_fFYUbEWo4_0),.din(w_dff_A_2jZUzQMO3_0),.clk(gclk));
	jdff dff_A_fFYUbEWo4_0(.dout(w_dff_A_CAVjaFLi4_0),.din(w_dff_A_fFYUbEWo4_0),.clk(gclk));
	jdff dff_A_CAVjaFLi4_0(.dout(w_dff_A_Q1qrKJZf1_0),.din(w_dff_A_CAVjaFLi4_0),.clk(gclk));
	jdff dff_A_Q1qrKJZf1_0(.dout(w_dff_A_xxeOSZzt9_0),.din(w_dff_A_Q1qrKJZf1_0),.clk(gclk));
	jdff dff_A_xxeOSZzt9_0(.dout(w_dff_A_W8bPgPiJ6_0),.din(w_dff_A_xxeOSZzt9_0),.clk(gclk));
	jdff dff_A_W8bPgPiJ6_0(.dout(G21),.din(w_dff_A_W8bPgPiJ6_0),.clk(gclk));
	jdff dff_A_VxBgzGut5_2(.dout(w_dff_A_UI9HFpeL2_0),.din(w_dff_A_VxBgzGut5_2),.clk(gclk));
	jdff dff_A_UI9HFpeL2_0(.dout(w_dff_A_qJrzVuab9_0),.din(w_dff_A_UI9HFpeL2_0),.clk(gclk));
	jdff dff_A_qJrzVuab9_0(.dout(w_dff_A_4j4wXiaz0_0),.din(w_dff_A_qJrzVuab9_0),.clk(gclk));
	jdff dff_A_4j4wXiaz0_0(.dout(w_dff_A_Aaedy9gb5_0),.din(w_dff_A_4j4wXiaz0_0),.clk(gclk));
	jdff dff_A_Aaedy9gb5_0(.dout(w_dff_A_lHlNJP5b7_0),.din(w_dff_A_Aaedy9gb5_0),.clk(gclk));
	jdff dff_A_lHlNJP5b7_0(.dout(w_dff_A_edZ4euLr7_0),.din(w_dff_A_lHlNJP5b7_0),.clk(gclk));
	jdff dff_A_edZ4euLr7_0(.dout(G24),.din(w_dff_A_edZ4euLr7_0),.clk(gclk));
	jdff dff_A_PCaNejM41_2(.dout(w_dff_A_muRMUgys2_0),.din(w_dff_A_PCaNejM41_2),.clk(gclk));
	jdff dff_A_muRMUgys2_0(.dout(w_dff_A_pVO7JxRf3_0),.din(w_dff_A_muRMUgys2_0),.clk(gclk));
	jdff dff_A_pVO7JxRf3_0(.dout(w_dff_A_cpS9pvUm5_0),.din(w_dff_A_pVO7JxRf3_0),.clk(gclk));
	jdff dff_A_cpS9pvUm5_0(.dout(w_dff_A_IhFQEkMO9_0),.din(w_dff_A_cpS9pvUm5_0),.clk(gclk));
	jdff dff_A_IhFQEkMO9_0(.dout(w_dff_A_xqSZaXoR3_0),.din(w_dff_A_IhFQEkMO9_0),.clk(gclk));
	jdff dff_A_xqSZaXoR3_0(.dout(w_dff_A_mCHTSb2L3_0),.din(w_dff_A_xqSZaXoR3_0),.clk(gclk));
	jdff dff_A_mCHTSb2L3_0(.dout(G27),.din(w_dff_A_mCHTSb2L3_0),.clk(gclk));
	jdff dff_A_XeL5ESXH3_2(.dout(w_dff_A_fy9LOIPT8_0),.din(w_dff_A_XeL5ESXH3_2),.clk(gclk));
	jdff dff_A_fy9LOIPT8_0(.dout(w_dff_A_xBgBFEHM7_0),.din(w_dff_A_fy9LOIPT8_0),.clk(gclk));
	jdff dff_A_xBgBFEHM7_0(.dout(w_dff_A_5gkAEx7I0_0),.din(w_dff_A_xBgBFEHM7_0),.clk(gclk));
	jdff dff_A_5gkAEx7I0_0(.dout(w_dff_A_TMpfrc1Q8_0),.din(w_dff_A_5gkAEx7I0_0),.clk(gclk));
	jdff dff_A_TMpfrc1Q8_0(.dout(w_dff_A_Li6WKKvL4_0),.din(w_dff_A_TMpfrc1Q8_0),.clk(gclk));
	jdff dff_A_Li6WKKvL4_0(.dout(w_dff_A_o6BgCzU64_0),.din(w_dff_A_Li6WKKvL4_0),.clk(gclk));
	jdff dff_A_o6BgCzU64_0(.dout(G33),.din(w_dff_A_o6BgCzU64_0),.clk(gclk));
	jdff dff_A_wxTTumbh8_2(.dout(w_dff_A_ilTLLlxC8_0),.din(w_dff_A_wxTTumbh8_2),.clk(gclk));
	jdff dff_A_ilTLLlxC8_0(.dout(w_dff_A_Bz7H5Wjt7_0),.din(w_dff_A_ilTLLlxC8_0),.clk(gclk));
	jdff dff_A_Bz7H5Wjt7_0(.dout(w_dff_A_pI5WLpcv6_0),.din(w_dff_A_Bz7H5Wjt7_0),.clk(gclk));
	jdff dff_A_pI5WLpcv6_0(.dout(w_dff_A_1NG3OYxR8_0),.din(w_dff_A_pI5WLpcv6_0),.clk(gclk));
	jdff dff_A_1NG3OYxR8_0(.dout(w_dff_A_jp2Wqpe77_0),.din(w_dff_A_1NG3OYxR8_0),.clk(gclk));
	jdff dff_A_jp2Wqpe77_0(.dout(w_dff_A_sZZkANDc0_0),.din(w_dff_A_jp2Wqpe77_0),.clk(gclk));
	jdff dff_A_sZZkANDc0_0(.dout(G36),.din(w_dff_A_sZZkANDc0_0),.clk(gclk));
	jdff dff_A_5ZGcPxwR6_2(.dout(w_dff_A_BQvTciW99_0),.din(w_dff_A_5ZGcPxwR6_2),.clk(gclk));
	jdff dff_A_BQvTciW99_0(.dout(w_dff_A_0hRpRr789_0),.din(w_dff_A_BQvTciW99_0),.clk(gclk));
	jdff dff_A_0hRpRr789_0(.dout(w_dff_A_DHl6Y7IQ9_0),.din(w_dff_A_0hRpRr789_0),.clk(gclk));
	jdff dff_A_DHl6Y7IQ9_0(.dout(w_dff_A_vT75EyGY5_0),.din(w_dff_A_DHl6Y7IQ9_0),.clk(gclk));
	jdff dff_A_vT75EyGY5_0(.dout(w_dff_A_hm112p493_0),.din(w_dff_A_vT75EyGY5_0),.clk(gclk));
	jdff dff_A_hm112p493_0(.dout(w_dff_A_teud1nbE4_0),.din(w_dff_A_hm112p493_0),.clk(gclk));
	jdff dff_A_teud1nbE4_0(.dout(G39),.din(w_dff_A_teud1nbE4_0),.clk(gclk));
	jdff dff_A_5MAg6puK2_2(.dout(w_dff_A_M4OfibrF1_0),.din(w_dff_A_5MAg6puK2_2),.clk(gclk));
	jdff dff_A_M4OfibrF1_0(.dout(w_dff_A_EzXgRwKQ9_0),.din(w_dff_A_M4OfibrF1_0),.clk(gclk));
	jdff dff_A_EzXgRwKQ9_0(.dout(w_dff_A_axJWYsxJ5_0),.din(w_dff_A_EzXgRwKQ9_0),.clk(gclk));
	jdff dff_A_axJWYsxJ5_0(.dout(w_dff_A_7f5mwdfI9_0),.din(w_dff_A_axJWYsxJ5_0),.clk(gclk));
	jdff dff_A_7f5mwdfI9_0(.dout(w_dff_A_8OmdQrkT4_0),.din(w_dff_A_7f5mwdfI9_0),.clk(gclk));
	jdff dff_A_8OmdQrkT4_0(.dout(w_dff_A_Y2dIFbtx4_0),.din(w_dff_A_8OmdQrkT4_0),.clk(gclk));
	jdff dff_A_Y2dIFbtx4_0(.dout(G42),.din(w_dff_A_Y2dIFbtx4_0),.clk(gclk));
	jdff dff_A_76IhHjB45_2(.dout(G75),.din(w_dff_A_76IhHjB45_2),.clk(gclk));
	jdff dff_A_STzXy76t1_2(.dout(G69),.din(w_dff_A_STzXy76t1_2),.clk(gclk));
	jdff dff_A_BblxUM767_2(.dout(w_dff_A_PknvDO025_0),.din(w_dff_A_BblxUM767_2),.clk(gclk));
	jdff dff_A_PknvDO025_0(.dout(G72),.din(w_dff_A_PknvDO025_0),.clk(gclk));
endmodule

