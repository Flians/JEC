/*

c7552:
	jxor: 242
	jspl: 295
	jspl3: 359
	jnot: 215
	jdff: 6368
	jor: 391
	jand: 479

Summary:
	jxor: 242
	jspl: 295
	jspl3: 359
	jnot: 215
	jdff: 6368
	jor: 391
	jand: 479
*/

module c7552(gclk, G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41, G44, G47, G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106, G109, G110, G111, G112, G113, G114, G115, G118, G121, G124, G127, G130, G133, G134, G135, G138, G141, G144, G147, G150, G151, G152, G153, G154, G155, G156, G157, G158, G159, G160, G161, G162, G163, G164, G165, G166, G167, G168, G169, G170, G171, G172, G173, G174, G175, G176, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G187, G188, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G216, G217, G218, G219, G220, G221, G222, G223, G224, G225, G226, G227, G228, G229, G230, G231, G232, G233, G234, G235, G236, G237, G238, G239, G240, G339, G1197, G1455, G1459, G1462, G1469, G1480, G1486, G1492, G1496, G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239, G2247, G2253, G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729, G3737, G3743, G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420, G4427, G4432, G4437, G4526, G4528, G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490, G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550, G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524, G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284, G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270, G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249, G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336, G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359, G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399);
	input gclk;
	input G1;
	input G5;
	input G9;
	input G12;
	input G15;
	input G18;
	input G23;
	input G26;
	input G29;
	input G32;
	input G35;
	input G38;
	input G41;
	input G44;
	input G47;
	input G50;
	input G53;
	input G54;
	input G55;
	input G56;
	input G57;
	input G58;
	input G59;
	input G60;
	input G61;
	input G62;
	input G63;
	input G64;
	input G65;
	input G66;
	input G69;
	input G70;
	input G73;
	input G74;
	input G75;
	input G76;
	input G77;
	input G78;
	input G79;
	input G80;
	input G81;
	input G82;
	input G83;
	input G84;
	input G85;
	input G86;
	input G87;
	input G88;
	input G89;
	input G94;
	input G97;
	input G100;
	input G103;
	input G106;
	input G109;
	input G110;
	input G111;
	input G112;
	input G113;
	input G114;
	input G115;
	input G118;
	input G121;
	input G124;
	input G127;
	input G130;
	input G133;
	input G134;
	input G135;
	input G138;
	input G141;
	input G144;
	input G147;
	input G150;
	input G151;
	input G152;
	input G153;
	input G154;
	input G155;
	input G156;
	input G157;
	input G158;
	input G159;
	input G160;
	input G161;
	input G162;
	input G163;
	input G164;
	input G165;
	input G166;
	input G167;
	input G168;
	input G169;
	input G170;
	input G171;
	input G172;
	input G173;
	input G174;
	input G175;
	input G176;
	input G177;
	input G178;
	input G179;
	input G180;
	input G181;
	input G182;
	input G183;
	input G184;
	input G185;
	input G186;
	input G187;
	input G188;
	input G189;
	input G190;
	input G191;
	input G192;
	input G193;
	input G194;
	input G195;
	input G196;
	input G197;
	input G198;
	input G199;
	input G200;
	input G201;
	input G202;
	input G203;
	input G204;
	input G205;
	input G206;
	input G207;
	input G208;
	input G209;
	input G210;
	input G211;
	input G212;
	input G213;
	input G214;
	input G215;
	input G216;
	input G217;
	input G218;
	input G219;
	input G220;
	input G221;
	input G222;
	input G223;
	input G224;
	input G225;
	input G226;
	input G227;
	input G228;
	input G229;
	input G230;
	input G231;
	input G232;
	input G233;
	input G234;
	input G235;
	input G236;
	input G237;
	input G238;
	input G239;
	input G240;
	input G339;
	input G1197;
	input G1455;
	input G1459;
	input G1462;
	input G1469;
	input G1480;
	input G1486;
	input G1492;
	input G1496;
	input G2204;
	input G2208;
	input G2211;
	input G2218;
	input G2224;
	input G2230;
	input G2236;
	input G2239;
	input G2247;
	input G2253;
	input G2256;
	input G3698;
	input G3701;
	input G3705;
	input G3711;
	input G3717;
	input G3723;
	input G3729;
	input G3737;
	input G3743;
	input G3749;
	input G4393;
	input G4394;
	input G4400;
	input G4405;
	input G4410;
	input G4415;
	input G4420;
	input G4427;
	input G4432;
	input G4437;
	input G4526;
	input G4528;
	output G2;
	output G3;
	output G450;
	output G448;
	output G444;
	output G442;
	output G440;
	output G438;
	output G496;
	output G494;
	output G492;
	output G490;
	output G488;
	output G486;
	output G484;
	output G482;
	output G480;
	output G560;
	output G542;
	output G558;
	output G556;
	output G554;
	output G552;
	output G550;
	output G548;
	output G546;
	output G544;
	output G540;
	output G538;
	output G536;
	output G534;
	output G532;
	output G530;
	output G528;
	output G526;
	output G524;
	output G279;
	output G436;
	output G478;
	output G522;
	output G402;
	output G404;
	output G406;
	output G408;
	output G410;
	output G432;
	output G446;
	output G284;
	output G286;
	output G289;
	output G292;
	output G341;
	output G281;
	output G453;
	output G278;
	output G373;
	output G246;
	output G258;
	output G264;
	output G270;
	output G388;
	output G391;
	output G394;
	output G397;
	output G376;
	output G379;
	output G382;
	output G385;
	output G412;
	output G414;
	output G416;
	output G249;
	output G295;
	output G324;
	output G252;
	output G276;
	output G310;
	output G313;
	output G316;
	output G319;
	output G327;
	output G330;
	output G333;
	output G336;
	output G418;
	output G273;
	output G298;
	output G301;
	output G304;
	output G307;
	output G344;
	output G422;
	output G469;
	output G419;
	output G471;
	output G359;
	output G362;
	output G365;
	output G368;
	output G347;
	output G350;
	output G353;
	output G356;
	output G321;
	output G338;
	output G370;
	output G399;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n345;
	wire n347;
	wire n348;
	wire n349;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1082;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1102;
	wire n1103;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1356;
	wire n1357;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1384;
	wire n1385;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1399;
	wire n1400;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1413;
	wire n1414;
	wire n1416;
	wire n1417;
	wire n1419;
	wire n1421;
	wire n1423;
	wire n1424;
	wire n1426;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire[2:0] w_G1_0;
	wire[2:0] w_G1_1;
	wire[2:0] w_G5_0;
	wire[1:0] w_G5_1;
	wire[2:0] w_G15_0;
	wire[2:0] w_G18_0;
	wire[2:0] w_G18_1;
	wire[2:0] w_G18_2;
	wire[2:0] w_G18_3;
	wire[2:0] w_G18_4;
	wire[2:0] w_G18_5;
	wire[2:0] w_G18_6;
	wire[2:0] w_G18_7;
	wire[2:0] w_G18_8;
	wire[2:0] w_G18_9;
	wire[2:0] w_G18_10;
	wire[2:0] w_G18_11;
	wire[2:0] w_G18_12;
	wire[2:0] w_G18_13;
	wire[2:0] w_G18_14;
	wire[2:0] w_G18_15;
	wire[2:0] w_G18_16;
	wire[2:0] w_G18_17;
	wire[2:0] w_G18_18;
	wire[2:0] w_G18_19;
	wire[2:0] w_G18_20;
	wire[2:0] w_G18_21;
	wire[2:0] w_G18_22;
	wire[2:0] w_G18_23;
	wire[2:0] w_G18_24;
	wire[2:0] w_G18_25;
	wire[2:0] w_G18_26;
	wire[2:0] w_G18_27;
	wire[2:0] w_G18_28;
	wire[2:0] w_G18_29;
	wire[2:0] w_G18_30;
	wire[2:0] w_G18_31;
	wire[2:0] w_G18_32;
	wire[2:0] w_G18_33;
	wire[2:0] w_G18_34;
	wire[2:0] w_G18_35;
	wire[2:0] w_G18_36;
	wire[2:0] w_G18_37;
	wire[2:0] w_G18_38;
	wire[2:0] w_G18_39;
	wire[2:0] w_G18_40;
	wire[2:0] w_G18_41;
	wire[2:0] w_G18_42;
	wire[2:0] w_G18_43;
	wire[2:0] w_G18_44;
	wire[2:0] w_G18_45;
	wire[2:0] w_G18_46;
	wire[2:0] w_G18_47;
	wire[2:0] w_G18_48;
	wire[2:0] w_G18_49;
	wire[1:0] w_G29_0;
	wire[2:0] w_G38_0;
	wire[2:0] w_G38_1;
	wire[2:0] w_G38_2;
	wire[1:0] w_G41_0;
	wire[1:0] w_G70_0;
	wire[1:0] w_G89_0;
	wire[2:0] w_G106_0;
	wire[1:0] w_G106_1;
	wire[1:0] w_G209_0;
	wire[1:0] w_G238_0;
	wire[2:0] w_G1455_0;
	wire[1:0] w_G1459_0;
	wire[1:0] w_G1462_0;
	wire[1:0] w_G1469_0;
	wire[2:0] w_G1480_0;
	wire[1:0] w_G1486_0;
	wire[2:0] w_G1492_0;
	wire[1:0] w_G1492_1;
	wire[2:0] w_G1496_0;
	wire[1:0] w_G1496_1;
	wire[2:0] w_G2204_0;
	wire[1:0] w_G2208_0;
	wire[2:0] w_G2211_0;
	wire[2:0] w_G2218_0;
	wire[2:0] w_G2224_0;
	wire[1:0] w_G2224_1;
	wire[2:0] w_G2230_0;
	wire[2:0] w_G2236_0;
	wire[2:0] w_G2239_0;
	wire[1:0] w_G2239_1;
	wire[2:0] w_G2247_0;
	wire[2:0] w_G2253_0;
	wire[1:0] w_G2256_0;
	wire[1:0] w_G3698_0;
	wire[2:0] w_G3701_0;
	wire[1:0] w_G3701_1;
	wire[2:0] w_G3705_0;
	wire[2:0] w_G3705_1;
	wire[1:0] w_G3711_0;
	wire[2:0] w_G3717_0;
	wire[2:0] w_G3723_0;
	wire[2:0] w_G3729_0;
	wire[1:0] w_G3729_1;
	wire[2:0] w_G3737_0;
	wire[2:0] w_G3743_0;
	wire[2:0] w_G3749_0;
	wire[1:0] w_G4393_0;
	wire[2:0] w_G4394_0;
	wire[1:0] w_G4394_1;
	wire[2:0] w_G4400_0;
	wire[1:0] w_G4400_1;
	wire[2:0] w_G4405_0;
	wire[1:0] w_G4405_1;
	wire[2:0] w_G4410_0;
	wire[2:0] w_G4415_0;
	wire[1:0] w_G4415_1;
	wire[2:0] w_G4420_0;
	wire[1:0] w_G4420_1;
	wire[2:0] w_G4427_0;
	wire[2:0] w_G4432_0;
	wire[2:0] w_G4437_0;
	wire[2:0] w_G4526_0;
	wire[2:0] w_G4526_1;
	wire[2:0] w_G4526_2;
	wire[2:0] w_G4528_0;
	wire w_G404_0;
	wire G404_fa_;
	wire w_G406_0;
	wire G406_fa_;
	wire w_G408_0;
	wire G408_fa_;
	wire w_G410_0;
	wire G410_fa_;
	wire w_G412_0;
	wire G412_fa_;
	wire w_G414_0;
	wire G414_fa_;
	wire w_G416_0;
	wire G416_fa_;
	wire w_G252_0;
	wire G252_fa_;
	wire[1:0] w_n345_0;
	wire[1:0] w_n347_0;
	wire[1:0] w_n349_0;
	wire[1:0] w_n353_0;
	wire[2:0] w_n354_0;
	wire[2:0] w_n355_0;
	wire[2:0] w_n355_1;
	wire[2:0] w_n355_2;
	wire[2:0] w_n355_3;
	wire[2:0] w_n355_4;
	wire[2:0] w_n355_5;
	wire[2:0] w_n355_6;
	wire[2:0] w_n355_7;
	wire[2:0] w_n355_8;
	wire[2:0] w_n355_9;
	wire[2:0] w_n355_10;
	wire[2:0] w_n355_11;
	wire[2:0] w_n355_12;
	wire[2:0] w_n355_13;
	wire[2:0] w_n355_14;
	wire[2:0] w_n355_15;
	wire[2:0] w_n355_16;
	wire[2:0] w_n355_17;
	wire[2:0] w_n355_18;
	wire[2:0] w_n355_19;
	wire[2:0] w_n355_20;
	wire[2:0] w_n355_21;
	wire[2:0] w_n355_22;
	wire[2:0] w_n355_23;
	wire[2:0] w_n355_24;
	wire[2:0] w_n355_25;
	wire[2:0] w_n355_26;
	wire[2:0] w_n355_27;
	wire[2:0] w_n355_28;
	wire[2:0] w_n355_29;
	wire[2:0] w_n355_30;
	wire[2:0] w_n355_31;
	wire[2:0] w_n355_32;
	wire[2:0] w_n355_33;
	wire[2:0] w_n355_34;
	wire[2:0] w_n355_35;
	wire[1:0] w_n357_0;
	wire[1:0] w_n358_0;
	wire[2:0] w_n359_0;
	wire[1:0] w_n359_1;
	wire[2:0] w_n361_0;
	wire[2:0] w_n362_0;
	wire[2:0] w_n363_0;
	wire[2:0] w_n364_0;
	wire[2:0] w_n366_0;
	wire[1:0] w_n367_0;
	wire[1:0] w_n368_0;
	wire[1:0] w_n369_0;
	wire[2:0] w_n370_0;
	wire[2:0] w_n371_0;
	wire[1:0] w_n372_0;
	wire[2:0] w_n373_0;
	wire[2:0] w_n373_1;
	wire[2:0] w_n373_2;
	wire[2:0] w_n373_3;
	wire[2:0] w_n373_4;
	wire[2:0] w_n373_5;
	wire[2:0] w_n373_6;
	wire[2:0] w_n373_7;
	wire[2:0] w_n373_8;
	wire[2:0] w_n373_9;
	wire[1:0] w_n374_0;
	wire[2:0] w_n375_0;
	wire[2:0] w_n377_0;
	wire[2:0] w_n377_1;
	wire[1:0] w_n378_0;
	wire[2:0] w_n379_0;
	wire[1:0] w_n380_0;
	wire[2:0] w_n383_0;
	wire[1:0] w_n385_0;
	wire[1:0] w_n386_0;
	wire[2:0] w_n387_0;
	wire[1:0] w_n387_1;
	wire[2:0] w_n388_0;
	wire[2:0] w_n388_1;
	wire[2:0] w_n389_0;
	wire[1:0] w_n389_1;
	wire[2:0] w_n391_0;
	wire[2:0] w_n392_0;
	wire[2:0] w_n393_0;
	wire[1:0] w_n393_1;
	wire[1:0] w_n394_0;
	wire[2:0] w_n395_0;
	wire[1:0] w_n395_1;
	wire[2:0] w_n396_0;
	wire[2:0] w_n396_1;
	wire[1:0] w_n397_0;
	wire[2:0] w_n405_0;
	wire[1:0] w_n407_0;
	wire[2:0] w_n409_0;
	wire[1:0] w_n409_1;
	wire[2:0] w_n411_0;
	wire[1:0] w_n411_1;
	wire[2:0] w_n413_0;
	wire[1:0] w_n413_1;
	wire[2:0] w_n414_0;
	wire[1:0] w_n414_1;
	wire[1:0] w_n415_0;
	wire[2:0] w_n416_0;
	wire[1:0] w_n418_0;
	wire[1:0] w_n419_0;
	wire[1:0] w_n420_0;
	wire[2:0] w_n421_0;
	wire[1:0] w_n422_0;
	wire[2:0] w_n423_0;
	wire[1:0] w_n424_0;
	wire[2:0] w_n425_0;
	wire[1:0] w_n425_1;
	wire[2:0] w_n426_0;
	wire[1:0] w_n427_0;
	wire[2:0] w_n428_0;
	wire[2:0] w_n429_0;
	wire[1:0] w_n430_0;
	wire[1:0] w_n431_0;
	wire[2:0] w_n432_0;
	wire[2:0] w_n433_0;
	wire[2:0] w_n433_1;
	wire[1:0] w_n434_0;
	wire[1:0] w_n435_0;
	wire[2:0] w_n436_0;
	wire[2:0] w_n437_0;
	wire[1:0] w_n438_0;
	wire[1:0] w_n440_0;
	wire[2:0] w_n444_0;
	wire[2:0] w_n445_0;
	wire[2:0] w_n447_0;
	wire[2:0] w_n449_0;
	wire[1:0] w_n449_1;
	wire[2:0] w_n450_0;
	wire[2:0] w_n451_0;
	wire[2:0] w_n453_0;
	wire[1:0] w_n453_1;
	wire[2:0] w_n456_0;
	wire[1:0] w_n457_0;
	wire[2:0] w_n459_0;
	wire[2:0] w_n460_0;
	wire[2:0] w_n460_1;
	wire[2:0] w_n462_0;
	wire[2:0] w_n463_0;
	wire[1:0] w_n463_1;
	wire[2:0] w_n464_0;
	wire[1:0] w_n465_0;
	wire[1:0] w_n466_0;
	wire[1:0] w_n467_0;
	wire[2:0] w_n469_0;
	wire[1:0] w_n469_1;
	wire[2:0] w_n470_0;
	wire[2:0] w_n471_0;
	wire[1:0] w_n472_0;
	wire[2:0] w_n474_0;
	wire[2:0] w_n475_0;
	wire[2:0] w_n476_0;
	wire[1:0] w_n477_0;
	wire[2:0] w_n479_0;
	wire[1:0] w_n479_1;
	wire[2:0] w_n480_0;
	wire[1:0] w_n480_1;
	wire[1:0] w_n481_0;
	wire[1:0] w_n485_0;
	wire[1:0] w_n486_0;
	wire[2:0] w_n487_0;
	wire[2:0] w_n489_0;
	wire[2:0] w_n491_0;
	wire[1:0] w_n491_1;
	wire[2:0] w_n495_0;
	wire[1:0] w_n495_1;
	wire[2:0] w_n496_0;
	wire[2:0] w_n497_0;
	wire[1:0] w_n497_1;
	wire[1:0] w_n499_0;
	wire[1:0] w_n500_0;
	wire[2:0] w_n501_0;
	wire[1:0] w_n503_0;
	wire[2:0] w_n504_0;
	wire[1:0] w_n504_1;
	wire[1:0] w_n505_0;
	wire[1:0] w_n507_0;
	wire[2:0] w_n509_0;
	wire[1:0] w_n511_0;
	wire[2:0] w_n512_0;
	wire[2:0] w_n513_0;
	wire[1:0] w_n513_1;
	wire[1:0] w_n514_0;
	wire[1:0] w_n516_0;
	wire[2:0] w_n517_0;
	wire[1:0] w_n517_1;
	wire[2:0] w_n518_0;
	wire[2:0] w_n518_1;
	wire[1:0] w_n520_0;
	wire[1:0] w_n522_0;
	wire[2:0] w_n523_0;
	wire[2:0] w_n524_0;
	wire[2:0] w_n524_1;
	wire[2:0] w_n526_0;
	wire[1:0] w_n528_0;
	wire[1:0] w_n530_0;
	wire[2:0] w_n531_0;
	wire[1:0] w_n531_1;
	wire[2:0] w_n536_0;
	wire[1:0] w_n538_0;
	wire[2:0] w_n539_0;
	wire[1:0] w_n539_1;
	wire[1:0] w_n544_0;
	wire[1:0] w_n546_0;
	wire[2:0] w_n547_0;
	wire[1:0] w_n547_1;
	wire[1:0] w_n548_0;
	wire[1:0] w_n550_0;
	wire[1:0] w_n552_0;
	wire[1:0] w_n554_0;
	wire[2:0] w_n555_0;
	wire[1:0] w_n555_1;
	wire[2:0] w_n556_0;
	wire[1:0] w_n558_0;
	wire[1:0] w_n560_0;
	wire[1:0] w_n562_0;
	wire[2:0] w_n563_0;
	wire[1:0] w_n563_1;
	wire[2:0] w_n564_0;
	wire[1:0] w_n565_0;
	wire[2:0] w_n566_0;
	wire[2:0] w_n568_0;
	wire[2:0] w_n570_0;
	wire[2:0] w_n570_1;
	wire[2:0] w_n572_0;
	wire[1:0] w_n572_1;
	wire[2:0] w_n573_0;
	wire[1:0] w_n573_1;
	wire[2:0] w_n574_0;
	wire[2:0] w_n575_0;
	wire[1:0] w_n575_1;
	wire[2:0] w_n576_0;
	wire[1:0] w_n577_0;
	wire[2:0] w_n578_0;
	wire[2:0] w_n580_0;
	wire[2:0] w_n581_0;
	wire[2:0] w_n582_0;
	wire[1:0] w_n584_0;
	wire[2:0] w_n585_0;
	wire[1:0] w_n585_1;
	wire[2:0] w_n586_0;
	wire[1:0] w_n588_0;
	wire[2:0] w_n590_0;
	wire[1:0] w_n592_0;
	wire[2:0] w_n593_0;
	wire[1:0] w_n593_1;
	wire[2:0] w_n594_0;
	wire[2:0] w_n595_0;
	wire[1:0] w_n597_0;
	wire[2:0] w_n598_0;
	wire[1:0] w_n598_1;
	wire[2:0] w_n599_0;
	wire[1:0] w_n600_0;
	wire[1:0] w_n602_0;
	wire[2:0] w_n603_0;
	wire[1:0] w_n603_1;
	wire[1:0] w_n604_0;
	wire[2:0] w_n605_0;
	wire[1:0] w_n609_0;
	wire[1:0] w_n610_0;
	wire[1:0] w_n612_0;
	wire[2:0] w_n613_0;
	wire[2:0] w_n615_0;
	wire[1:0] w_n616_0;
	wire[2:0] w_n618_0;
	wire[2:0] w_n619_0;
	wire[2:0] w_n622_0;
	wire[1:0] w_n624_0;
	wire[2:0] w_n625_0;
	wire[1:0] w_n625_1;
	wire[2:0] w_n626_0;
	wire[1:0] w_n626_1;
	wire[2:0] w_n627_0;
	wire[1:0] w_n629_0;
	wire[2:0] w_n630_0;
	wire[2:0] w_n631_0;
	wire[2:0] w_n632_0;
	wire[1:0] w_n632_1;
	wire[1:0] w_n634_0;
	wire[2:0] w_n635_0;
	wire[1:0] w_n635_1;
	wire[2:0] w_n636_0;
	wire[2:0] w_n641_0;
	wire[2:0] w_n642_0;
	wire[1:0] w_n644_0;
	wire[1:0] w_n645_0;
	wire[1:0] w_n646_0;
	wire[1:0] w_n647_0;
	wire[1:0] w_n649_0;
	wire[1:0] w_n651_0;
	wire[1:0] w_n652_0;
	wire[1:0] w_n653_0;
	wire[2:0] w_n654_0;
	wire[1:0] w_n655_0;
	wire[1:0] w_n656_0;
	wire[2:0] w_n657_0;
	wire[1:0] w_n659_0;
	wire[2:0] w_n660_0;
	wire[2:0] w_n661_0;
	wire[1:0] w_n662_0;
	wire[2:0] w_n663_0;
	wire[1:0] w_n663_1;
	wire[1:0] w_n664_0;
	wire[1:0] w_n666_0;
	wire[1:0] w_n669_0;
	wire[1:0] w_n671_0;
	wire[2:0] w_n673_0;
	wire[1:0] w_n674_0;
	wire[2:0] w_n676_0;
	wire[1:0] w_n678_0;
	wire[2:0] w_n680_0;
	wire[2:0] w_n680_1;
	wire[2:0] w_n680_2;
	wire[1:0] w_n682_0;
	wire[1:0] w_n683_0;
	wire[1:0] w_n687_0;
	wire[1:0] w_n689_0;
	wire[1:0] w_n690_0;
	wire[1:0] w_n693_0;
	wire[1:0] w_n694_0;
	wire[1:0] w_n695_0;
	wire[1:0] w_n696_0;
	wire[1:0] w_n698_0;
	wire[2:0] w_n700_0;
	wire[1:0] w_n700_1;
	wire[2:0] w_n703_0;
	wire[2:0] w_n703_1;
	wire[1:0] w_n705_0;
	wire[2:0] w_n707_0;
	wire[2:0] w_n707_1;
	wire[2:0] w_n709_0;
	wire[1:0] w_n709_1;
	wire[2:0] w_n711_0;
	wire[1:0] w_n711_1;
	wire[2:0] w_n712_0;
	wire[1:0] w_n713_0;
	wire[2:0] w_n715_0;
	wire[1:0] w_n715_1;
	wire[2:0] w_n718_0;
	wire[1:0] w_n719_0;
	wire[2:0] w_n720_0;
	wire[2:0] w_n723_0;
	wire[1:0] w_n724_0;
	wire[1:0] w_n725_0;
	wire[2:0] w_n726_0;
	wire[1:0] w_n726_1;
	wire[2:0] w_n729_0;
	wire[1:0] w_n729_1;
	wire[2:0] w_n734_0;
	wire[1:0] w_n736_0;
	wire[2:0] w_n737_0;
	wire[1:0] w_n737_1;
	wire[2:0] w_n741_0;
	wire[1:0] w_n741_1;
	wire[1:0] w_n743_0;
	wire[2:0] w_n744_0;
	wire[2:0] w_n747_0;
	wire[1:0] w_n749_0;
	wire[1:0] w_n754_0;
	wire[2:0] w_n755_0;
	wire[1:0] w_n755_1;
	wire[2:0] w_n758_0;
	wire[1:0] w_n758_1;
	wire[1:0] w_n760_0;
	wire[2:0] w_n761_0;
	wire[2:0] w_n764_0;
	wire[1:0] w_n766_0;
	wire[1:0] w_n767_0;
	wire[2:0] w_n768_0;
	wire[2:0] w_n772_0;
	wire[1:0] w_n773_0;
	wire[1:0] w_n774_0;
	wire[1:0] w_n775_0;
	wire[2:0] w_n776_0;
	wire[2:0] w_n780_0;
	wire[1:0] w_n781_0;
	wire[2:0] w_n796_0;
	wire[1:0] w_n796_1;
	wire[2:0] w_n800_0;
	wire[1:0] w_n800_1;
	wire[2:0] w_n803_0;
	wire[2:0] w_n806_0;
	wire[1:0] w_n808_0;
	wire[2:0] w_n810_0;
	wire[1:0] w_n810_1;
	wire[2:0] w_n814_0;
	wire[1:0] w_n814_1;
	wire[2:0] w_n817_0;
	wire[2:0] w_n820_0;
	wire[1:0] w_n822_0;
	wire[2:0] w_n824_0;
	wire[2:0] w_n827_0;
	wire[2:0] w_n845_0;
	wire[1:0] w_n845_1;
	wire[2:0] w_n848_0;
	wire[1:0] w_n848_1;
	wire[2:0] w_n851_0;
	wire[2:0] w_n854_0;
	wire[1:0] w_n856_0;
	wire[2:0] w_n858_0;
	wire[2:0] w_n862_0;
	wire[1:0] w_n863_0;
	wire[1:0] w_n864_0;
	wire[2:0] w_n866_0;
	wire[2:0] w_n870_0;
	wire[1:0] w_n871_0;
	wire[2:0] w_n885_0;
	wire[2:0] w_n888_0;
	wire[2:0] w_n891_0;
	wire[2:0] w_n894_0;
	wire[1:0] w_n895_0;
	wire[2:0] w_n900_0;
	wire[2:0] w_n903_0;
	wire[1:0] w_n905_0;
	wire[2:0] w_n916_0;
	wire[2:0] w_n919_0;
	wire[2:0] w_n926_0;
	wire[2:0] w_n930_0;
	wire[2:0] w_n935_0;
	wire[2:0] w_n938_0;
	wire[2:0] w_n944_0;
	wire[2:0] w_n947_0;
	wire[2:0] w_n950_0;
	wire[1:0] w_n950_1;
	wire[2:0] w_n953_0;
	wire[1:0] w_n953_1;
	wire[2:0] w_n966_0;
	wire[2:0] w_n970_0;
	wire[2:0] w_n973_0;
	wire[1:0] w_n973_1;
	wire[2:0] w_n977_0;
	wire[1:0] w_n977_1;
	wire[2:0] w_n980_0;
	wire[2:0] w_n983_0;
	wire[1:0] w_n985_0;
	wire[2:0] w_n987_0;
	wire[2:0] w_n991_0;
	wire[1:0] w_n992_0;
	wire[2:0] w_n995_0;
	wire[2:0] w_n999_0;
	wire[1:0] w_n1000_0;
	wire[1:0] w_n1003_0;
	wire[1:0] w_n1007_0;
	wire[1:0] w_n1008_0;
	wire[1:0] w_n1042_0;
	wire[2:0] w_n1059_0;
	wire[2:0] w_n1067_0;
	wire[2:0] w_n1069_0;
	wire[1:0] w_n1070_0;
	wire[1:0] w_n1073_0;
	wire[1:0] w_n1078_0;
	wire[2:0] w_n1084_0;
	wire[1:0] w_n1086_0;
	wire[1:0] w_n1090_0;
	wire[2:0] w_n1092_0;
	wire[2:0] w_n1094_0;
	wire[1:0] w_n1096_0;
	wire[1:0] w_n1099_0;
	wire[1:0] w_n1105_0;
	wire[1:0] w_n1106_0;
	wire[1:0] w_n1108_0;
	wire[1:0] w_n1113_0;
	wire[1:0] w_n1118_0;
	wire[1:0] w_n1127_0;
	wire[1:0] w_n1137_0;
	wire[1:0] w_n1150_0;
	wire[1:0] w_n1172_0;
	wire[1:0] w_n1307_0;
	wire[1:0] w_n1308_0;
	wire[1:0] w_n1309_0;
	wire[1:0] w_n1310_0;
	wire[2:0] w_n1312_0;
	wire[1:0] w_n1312_1;
	wire[1:0] w_n1316_0;
	wire[1:0] w_n1317_0;
	wire[2:0] w_n1321_0;
	wire[1:0] w_n1321_1;
	wire[1:0] w_n1323_0;
	wire[1:0] w_n1333_0;
	wire[2:0] w_n1337_0;
	wire[1:0] w_n1337_1;
	wire[2:0] w_n1340_0;
	wire[1:0] w_n1343_0;
	wire[1:0] w_n1344_0;
	wire[1:0] w_n1359_0;
	wire[1:0] w_n1364_0;
	wire[1:0] w_n1369_0;
	wire[1:0] w_n1370_0;
	wire[1:0] w_n1372_0;
	wire[1:0] w_n1387_0;
	wire[1:0] w_n1388_0;
	wire[1:0] w_n1396_0;
	wire[1:0] w_n1402_0;
	wire[1:0] w_n1408_0;
	wire[1:0] w_n1419_0;
	wire[1:0] w_n1426_0;
	wire[1:0] w_n1431_0;
	wire[1:0] w_n1433_0;
	wire[1:0] w_n1440_0;
	wire[2:0] w_n1452_0;
	wire[1:0] w_n1458_0;
	wire[1:0] w_n1486_0;
	wire[1:0] w_n1492_0;
	wire[1:0] w_n1506_0;
	wire[1:0] w_n1511_0;
	wire[1:0] w_n1518_0;
	wire[1:0] w_n1529_0;
	wire[1:0] w_n1531_0;
	wire[1:0] w_n1534_0;
	wire[1:0] w_n1536_0;
	wire[1:0] w_n1543_0;
	wire[1:0] w_n1554_0;
	wire[2:0] w_n1562_0;
	wire[1:0] w_n1587_0;
	wire[1:0] w_n1597_0;
	wire[1:0] w_n1605_0;
	wire[1:0] w_n1607_0;
	wire[1:0] w_n1610_0;
	wire[1:0] w_n1620_0;
	wire[1:0] w_n1624_0;
	wire w_dff_A_T5tMKu6E2_0;
	wire w_dff_A_oNTQhwtA1_1;
	wire w_dff_A_1a3BOk4N7_2;
	wire w_dff_B_zOw0FkEF5_2;
	wire w_dff_B_6U6LXPHR6_0;
	wire w_dff_B_TjLqO1u54_1;
	wire w_dff_B_97wWmE6h6_1;
	wire w_dff_B_4VCGVyj24_1;
	wire w_dff_B_ufsFaH6f3_1;
	wire w_dff_B_CyEW83ti4_1;
	wire w_dff_B_1jFsO2pC0_1;
	wire w_dff_B_2hcssRmX0_1;
	wire w_dff_B_Fh2yl14E5_1;
	wire w_dff_B_RRky67T19_1;
	wire w_dff_B_qIlkOmM51_1;
	wire w_dff_B_3HpaRzXJ5_1;
	wire w_dff_B_kaDHWLyL4_1;
	wire w_dff_B_rPJsex3M4_1;
	wire w_dff_B_JcuS8AgU8_1;
	wire w_dff_B_0kzfT6xZ6_1;
	wire w_dff_B_SROuIGVL6_1;
	wire w_dff_B_Tw8HPB605_1;
	wire w_dff_B_QEsPxDpC0_1;
	wire w_dff_B_QtIF5Vso0_0;
	wire w_dff_B_QMWRNQhZ5_0;
	wire w_dff_B_li2eQKuw8_0;
	wire w_dff_B_HpNPKjcS6_0;
	wire w_dff_B_RFd3dZtY3_0;
	wire w_dff_B_if3aMaBK6_0;
	wire w_dff_B_4nECUVdc6_0;
	wire w_dff_B_Vc1PWlxZ1_0;
	wire w_dff_B_KWdKesqb8_0;
	wire w_dff_B_qOsK37uE5_0;
	wire w_dff_B_n2qIGD8l4_0;
	wire w_dff_B_3OPqg3A28_0;
	wire w_dff_B_o4x9k8Hm3_0;
	wire w_dff_B_dDhKryAR8_0;
	wire w_dff_B_lLGJXY3r1_0;
	wire w_dff_B_mjsGBemm5_0;
	wire w_dff_B_junc3TOI5_1;
	wire w_dff_B_2yB9OqOV3_1;
	wire w_dff_B_Et9qnbCU0_1;
	wire w_dff_B_ANo0zDnp6_1;
	wire w_dff_B_qkNvFZIn9_1;
	wire w_dff_B_Mmpnp9mB6_1;
	wire w_dff_B_07ZkajnW5_1;
	wire w_dff_B_Mu0xTX3i7_1;
	wire w_dff_B_gHZo3aqe3_1;
	wire w_dff_B_imUXYW195_0;
	wire w_dff_B_JO3UKFHT7_0;
	wire w_dff_B_v38kqikO1_0;
	wire w_dff_B_kcXzZ2IU4_0;
	wire w_dff_B_Bm2F6y6y6_0;
	wire w_dff_B_H57zb1K81_0;
	wire w_dff_B_Xa7VGz1K9_0;
	wire w_dff_B_6E66sqbu1_0;
	wire w_dff_B_73ua5IHw6_0;
	wire w_dff_B_2ocE5viI8_0;
	wire w_dff_B_uGZGQZJL0_0;
	wire w_dff_B_GScmS10K5_0;
	wire w_dff_B_VJyiFUPr6_0;
	wire w_dff_B_v7D954u79_0;
	wire w_dff_B_0sRoyxnh1_0;
	wire w_dff_B_c7MJRDtg1_0;
	wire w_dff_B_ZR0Rcscs5_0;
	wire w_dff_B_kJItpt9r0_1;
	wire w_dff_B_4WtbBNc87_1;
	wire w_dff_A_CphRJuGg1_0;
	wire w_dff_B_55reXz6K6_1;
	wire w_dff_B_AQ3bK5jI6_1;
	wire w_dff_B_9ccSpmjd7_1;
	wire w_dff_B_QBQeBDuX0_1;
	wire w_dff_B_ikunosyf0_1;
	wire w_dff_B_2xlYf5BN1_1;
	wire w_dff_B_KJhSDUHe8_1;
	wire w_dff_B_AtHwi2QQ7_1;
	wire w_dff_B_UggBC4N44_1;
	wire w_dff_B_lwHLunpJ9_1;
	wire w_dff_B_2rjIlNi35_1;
	wire w_dff_B_Gkd9alQJ7_1;
	wire w_dff_B_Xp10PR8c9_1;
	wire w_dff_B_3C0Jcu5e6_1;
	wire w_dff_B_XhyAd35E2_1;
	wire w_dff_B_iUyAeNp71_1;
	wire w_dff_B_LYCb3kK50_1;
	wire w_dff_B_BEKYu4Ds1_1;
	wire w_dff_B_n5fF0UMc1_1;
	wire w_dff_B_0hEaJtkG7_1;
	wire w_dff_B_ABL8kD7e8_1;
	wire w_dff_B_6oJjkDGb9_1;
	wire w_dff_B_BpEyDqFM3_1;
	wire w_dff_B_TTQ6jrHG5_1;
	wire w_dff_B_kD2uZm3u0_1;
	wire w_dff_B_PLBi3gOJ4_1;
	wire w_dff_B_PkwjJBL94_1;
	wire w_dff_B_eeLuYLuh1_1;
	wire w_dff_B_AN1m9qJC1_1;
	wire w_dff_B_2GmbTt8p1_1;
	wire w_dff_B_tnrcfJL44_0;
	wire w_dff_B_YTrADmT94_0;
	wire w_dff_B_JUkwTrJG5_0;
	wire w_dff_B_87pkms7O0_0;
	wire w_dff_B_V7NRqf8f6_0;
	wire w_dff_B_uwiXtHGO0_0;
	wire w_dff_B_xsDK7qTa1_0;
	wire w_dff_B_2xUTUYxk9_0;
	wire w_dff_B_DalyDTKL9_0;
	wire w_dff_B_hrGNiiTO6_0;
	wire w_dff_B_B3aBrb1W9_0;
	wire w_dff_B_hc5zIjFW5_0;
	wire w_dff_B_NzmYv2Ju3_0;
	wire w_dff_B_JFomYLpH8_0;
	wire w_dff_B_VNYPqclP3_0;
	wire w_dff_B_ZwTl6rAk0_0;
	wire w_dff_B_mwrMtZeR5_1;
	wire w_dff_B_QCwqzs4K5_1;
	wire w_dff_B_KrCqQOpC8_1;
	wire w_dff_B_VYSGL44K4_1;
	wire w_dff_B_y0iAhE1x1_1;
	wire w_dff_B_gaAUvedO2_1;
	wire w_dff_B_DDaQ0Nhf4_1;
	wire w_dff_B_Awj8k4IR0_1;
	wire w_dff_B_djD8XoOW9_1;
	wire w_dff_B_l9p2k1Q35_1;
	wire w_dff_B_CXoIoVTw8_1;
	wire w_dff_B_4QyVYSAf5_1;
	wire w_dff_B_H3Db3hF04_1;
	wire w_dff_B_H15ONvw94_1;
	wire w_dff_B_5Te35amx6_1;
	wire w_dff_B_d2014slu1_1;
	wire w_dff_B_Fv9Tf1Do3_1;
	wire w_dff_B_IeXeeWmW2_1;
	wire w_dff_B_BbmWtOQG4_1;
	wire w_dff_B_h8N6Mso09_1;
	wire w_dff_B_Esn3nXfG9_1;
	wire w_dff_B_3XYmJmJV0_1;
	wire w_dff_B_c8bI1Gsq5_1;
	wire w_dff_B_VFnSsohA1_1;
	wire w_dff_B_9EZCnDqB9_0;
	wire w_dff_B_krIL2Sla4_0;
	wire w_dff_B_vIDtoBo01_0;
	wire w_dff_B_WfQNlUCq7_0;
	wire w_dff_B_oI7Ro3ve0_0;
	wire w_dff_B_RZ1doWGM3_0;
	wire w_dff_B_bTzE2Vb16_0;
	wire w_dff_B_UKak35Q27_0;
	wire w_dff_B_47WPA4wK6_0;
	wire w_dff_B_sy7JW3no2_0;
	wire w_dff_B_SEsKKMeJ7_0;
	wire w_dff_B_clx5t3Ka4_0;
	wire w_dff_B_hr7f8krV9_0;
	wire w_dff_B_AdyRxg5x1_0;
	wire w_dff_B_AL4TOg2N8_0;
	wire w_dff_B_zMHrUpc90_0;
	wire w_dff_B_yE5DwyML5_1;
	wire w_dff_B_FWBTaxcO4_1;
	wire w_dff_B_9aw3Afxr6_0;
	wire w_dff_A_Eg7cyhMt0_1;
	wire w_dff_A_KeH7Nrrb3_1;
	wire w_dff_B_Ddj01x9g8_0;
	wire w_dff_B_O1JLdrLw2_1;
	wire w_dff_A_enWUTCuu1_1;
	wire w_dff_B_E8nBb3DH5_2;
	wire w_dff_B_XAAgdeGg2_1;
	wire w_dff_B_I5FCwES43_1;
	wire w_dff_B_MlLdonTk2_1;
	wire w_dff_B_sGNYDTMf1_1;
	wire w_dff_B_2G7vtFay6_1;
	wire w_dff_B_Dt6dA6I30_1;
	wire w_dff_A_JsJXQnTB5_1;
	wire w_dff_A_RZ0RSApD5_1;
	wire w_dff_A_oi0Er4UG6_1;
	wire w_dff_A_M57ltLga8_1;
	wire w_dff_B_wkAoRgPc7_3;
	wire w_dff_B_PmmN9UCR7_3;
	wire w_dff_B_AhAyDMWW2_3;
	wire w_dff_B_5lKdJiw20_3;
	wire w_dff_B_Fx4k30Tr9_3;
	wire w_dff_B_dF9Rz8HV0_3;
	wire w_dff_B_QlWGqAmt3_3;
	wire w_dff_B_QH6vNJpY5_3;
	wire w_dff_B_5cdujKON1_3;
	wire w_dff_B_QrESFXZm3_3;
	wire w_dff_B_wUXpcn6J7_3;
	wire w_dff_B_wBxjDCTh1_3;
	wire w_dff_B_AuPEkyDQ4_3;
	wire w_dff_B_9XVIZCmG7_3;
	wire w_dff_B_pplEk7n83_3;
	wire w_dff_B_WO7SOUzB9_3;
	wire w_dff_B_RgiMDdgi4_3;
	wire w_dff_B_3CbOvO5n8_3;
	wire w_dff_B_4R7OiaOD7_3;
	wire w_dff_B_rj9Ym2rU0_3;
	wire w_dff_B_fV29Gfar9_3;
	wire w_dff_B_HSiGjv8v6_3;
	wire w_dff_B_3zJjK5z10_3;
	wire w_dff_B_KT5fBCnk8_3;
	wire w_dff_B_HX5r9EjC7_0;
	wire w_dff_B_ppAVmaDk9_1;
	wire w_dff_B_jGtEyOsT0_1;
	wire w_dff_B_APeBZFjU6_1;
	wire w_dff_B_jzw1SDOq0_1;
	wire w_dff_B_NUTPwWig2_1;
	wire w_dff_B_aFKDUAAb1_1;
	wire w_dff_B_pYbMP1xr9_1;
	wire w_dff_B_WWZoYfmp3_1;
	wire w_dff_B_BqJSAS7T3_1;
	wire w_dff_B_7XmpVo0t3_1;
	wire w_dff_B_5QrLIniJ8_1;
	wire w_dff_B_ANLS58eZ7_1;
	wire w_dff_B_VZtkMsey5_1;
	wire w_dff_B_ZdGQvklp9_1;
	wire w_dff_B_T1FzLBe52_1;
	wire w_dff_B_g0FDj0mJ9_1;
	wire w_dff_B_ZsfmaTUk9_1;
	wire w_dff_B_yhjINwvk2_1;
	wire w_dff_B_D2oOjfBR4_1;
	wire w_dff_B_le0XpBTs7_1;
	wire w_dff_B_A7AGMUKI9_1;
	wire w_dff_B_fnd0kqBg8_1;
	wire w_dff_B_2nEbmhW49_1;
	wire w_dff_B_WRoDaIlx8_1;
	wire w_dff_B_c96qlGPT9_1;
	wire w_dff_B_DIMC7OCW0_1;
	wire w_dff_B_0xnUJhc19_1;
	wire w_dff_B_CEqWA62t8_1;
	wire w_dff_B_ahWALvHo2_1;
	wire w_dff_B_oOPoAVln8_1;
	wire w_dff_B_1JamPVks3_1;
	wire w_dff_B_bwgk3luk8_1;
	wire w_dff_B_1NeJ41o38_1;
	wire w_dff_B_Zh41odSJ6_1;
	wire w_dff_B_ROdLkkHL3_1;
	wire w_dff_B_lsmqHwtk6_1;
	wire w_dff_B_LXeHp9zA5_1;
	wire w_dff_B_xkwPng879_1;
	wire w_dff_B_YUPn6mdh1_1;
	wire w_dff_B_SnQXJfha5_1;
	wire w_dff_B_Y4vEEvQ13_1;
	wire w_dff_B_3PRK96Yo5_0;
	wire w_dff_B_CexrjSCz3_0;
	wire w_dff_B_n1cRIjSk2_0;
	wire w_dff_B_U8Mv3Hj79_0;
	wire w_dff_B_ZSzFuQvI4_0;
	wire w_dff_B_oaJJPAP00_0;
	wire w_dff_B_SphKZ9Px2_0;
	wire w_dff_B_w7bN5dAK4_0;
	wire w_dff_B_0Tk8qq6q4_0;
	wire w_dff_B_0r9O8Azb5_0;
	wire w_dff_B_qT45hAnc6_0;
	wire w_dff_B_jnT5tqD47_0;
	wire w_dff_B_AduYHKX63_1;
	wire w_dff_B_77aJXqCp8_1;
	wire w_dff_B_9VJ5u3Ms8_1;
	wire w_dff_B_lDVCWs0x5_1;
	wire w_dff_B_woLyC5fT9_0;
	wire w_dff_B_A6CLlKNI3_0;
	wire w_dff_B_T6Uv8ky34_1;
	wire w_dff_B_rCzq5duE1_0;
	wire w_dff_B_H3R4MueT7_0;
	wire w_dff_B_XuQVTKfc1_0;
	wire w_dff_B_qNMshn2w7_1;
	wire w_dff_B_xTcMbHgz3_1;
	wire w_dff_B_ZYclXlcM2_1;
	wire w_dff_B_RQkOQna85_1;
	wire w_dff_B_BkNagHHh6_1;
	wire w_dff_B_iPp6XAEi3_0;
	wire w_dff_B_duw1jA3D8_0;
	wire w_dff_B_TLv5oiTp8_0;
	wire w_dff_A_nWFur3Lc4_0;
	wire w_dff_A_zKfZMW4N9_0;
	wire w_dff_A_o6NPZiL11_0;
	wire w_dff_A_XqgRxEJy4_0;
	wire w_dff_B_3gV6bLg16_1;
	wire w_dff_A_c6ksV2It6_0;
	wire w_dff_A_Tss7Uoax4_1;
	wire w_dff_A_lzsf9YNj2_1;
	wire w_dff_B_Xus4ekrH4_2;
	wire w_dff_B_mvlVMQb49_0;
	wire w_dff_B_pZ8lh82s2_0;
	wire w_dff_B_CT3fc92M1_0;
	wire w_dff_B_xd3cfJjR0_0;
	wire w_dff_B_EmzoD31v6_0;
	wire w_dff_B_nwKB96Tv8_0;
	wire w_dff_B_HKXq822L7_1;
	wire w_dff_B_Lhoo9HH01_0;
	wire w_dff_B_F8nFENal5_0;
	wire w_dff_B_uu1JPCKy3_0;
	wire w_dff_B_1qaZhbnY0_0;
	wire w_dff_B_Z1wa6H460_0;
	wire w_dff_B_JueNAneB1_0;
	wire w_dff_B_nd8RMhdZ1_0;
	wire w_dff_B_7kP8I6Nv7_0;
	wire w_dff_B_HtoLOBwu0_0;
	wire w_dff_B_p4w6oiXH2_0;
	wire w_dff_B_EAGu5l770_0;
	wire w_dff_B_funZwnL82_0;
	wire w_dff_B_tSORCQTA6_0;
	wire w_dff_B_vpZpWSVG6_0;
	wire w_dff_B_D3MvhOYV3_0;
	wire w_dff_B_DRHH5VbM8_0;
	wire w_dff_B_Y2y7A30A9_0;
	wire w_dff_B_vgFcF65u4_0;
	wire w_dff_B_oCrv8doN3_1;
	wire w_dff_B_RmpkDI601_1;
	wire w_dff_B_DUUq7Zzj9_1;
	wire w_dff_B_jXWBPfOv2_0;
	wire w_dff_B_Z1KLiv0J5_0;
	wire w_dff_B_wzfHBs9Y7_0;
	wire w_dff_B_BlvzTLvr5_0;
	wire w_dff_A_VkhTzqs80_0;
	wire w_dff_A_RAnhR2Ke5_0;
	wire w_dff_B_gEZBHIQa1_0;
	wire w_dff_B_XLgbErkX1_1;
	wire w_dff_A_G2KgPMH80_1;
	wire w_dff_A_AEaRPL7B0_1;
	wire w_dff_B_TlGkzb2R8_1;
	wire w_dff_B_Q8Ztu0Pv0_1;
	wire w_dff_B_ASG2Rf5Z3_1;
	wire w_dff_B_ebtfvnBV1_1;
	wire w_dff_B_O7vbFofv9_1;
	wire w_dff_B_xilKJ2bD4_1;
	wire w_dff_B_wzUqhPo52_1;
	wire w_dff_B_uJ1Livi89_1;
	wire w_dff_B_3b6CDBYm8_1;
	wire w_dff_B_3lPQYY2G2_1;
	wire w_dff_B_ec7G6yed2_1;
	wire w_dff_B_eolntUTj5_1;
	wire w_dff_B_M9uQLkgk0_1;
	wire w_dff_B_jgexdI7w1_1;
	wire w_dff_B_9JvjqUzm1_1;
	wire w_dff_B_vvv6rMzV4_1;
	wire w_dff_B_Y04GqOKy9_1;
	wire w_dff_B_Z6wYFNCf8_1;
	wire w_dff_B_mzBNgqCu9_1;
	wire w_dff_B_ki0A4K324_1;
	wire w_dff_B_fjpEQ3Jo4_1;
	wire w_dff_B_qcZSPAcg4_1;
	wire w_dff_B_NzjvkRve8_1;
	wire w_dff_B_9m8w8OCT8_1;
	wire w_dff_B_N7BvwqaP7_1;
	wire w_dff_B_L4ss8y1M3_1;
	wire w_dff_B_EPO0p1Pn7_1;
	wire w_dff_B_D8ohgkie5_1;
	wire w_dff_B_aoyY9Iwj9_1;
	wire w_dff_B_DVk0kigS7_1;
	wire w_dff_B_ZozvfSql1_1;
	wire w_dff_B_iwN74MFK9_1;
	wire w_dff_B_CTYAs7z95_1;
	wire w_dff_B_vw8GA2Eg7_1;
	wire w_dff_B_OKTHmd9v8_1;
	wire w_dff_B_lzn87cmm9_1;
	wire w_dff_B_zxTxP1KQ0_1;
	wire w_dff_B_MzmrHBrI1_1;
	wire w_dff_B_z8PSb0fK2_1;
	wire w_dff_B_dvejynQC0_1;
	wire w_dff_B_pUvmZt6c4_1;
	wire w_dff_B_rwaob1yQ1_1;
	wire w_dff_B_S3HLASqu6_1;
	wire w_dff_B_pgbUEQQb9_1;
	wire w_dff_B_O5C0QGcS7_1;
	wire w_dff_B_MqArCBY05_1;
	wire w_dff_B_MqfVkYW82_1;
	wire w_dff_B_iJvWAqwt9_1;
	wire w_dff_B_scPDfLPg7_1;
	wire w_dff_B_OT03VlAw2_1;
	wire w_dff_B_zSoaRWf89_1;
	wire w_dff_B_Ii4PdT4b5_1;
	wire w_dff_B_TBzUmDJr7_1;
	wire w_dff_B_EXIhrkNU4_1;
	wire w_dff_B_ThSv8kmx6_1;
	wire w_dff_B_8pYQJq272_2;
	wire w_dff_B_YMbh9Iu96_2;
	wire w_dff_B_45it95Sr4_2;
	wire w_dff_B_yYsuVKir5_2;
	wire w_dff_B_VaF2Ke1S9_2;
	wire w_dff_B_Pikv11Vr8_2;
	wire w_dff_B_eAeKRf8c3_2;
	wire w_dff_B_VvI9QdN05_2;
	wire w_dff_B_J8I8Ps9A3_2;
	wire w_dff_B_8gcKVKG65_2;
	wire w_dff_B_yIEjn4Pn5_2;
	wire w_dff_B_jcZbdmaF2_2;
	wire w_dff_B_skB34im25_2;
	wire w_dff_B_KbuqKSM01_2;
	wire w_dff_B_JNirCrmu0_2;
	wire w_dff_B_ylluQ5Kf2_2;
	wire w_dff_B_5e84sic98_2;
	wire w_dff_B_IjfXU1yO3_2;
	wire w_dff_B_mhnhOjzv2_2;
	wire w_dff_B_5Oakuo148_2;
	wire w_dff_B_CCM2iDWJ7_2;
	wire w_dff_B_7XyHSN1D7_2;
	wire w_dff_B_MDSQJJpu9_2;
	wire w_dff_B_KuG2qXsX3_2;
	wire w_dff_B_pbgTkE6x3_2;
	wire w_dff_B_rTO6oFH15_2;
	wire w_dff_B_U29MVMUq1_2;
	wire w_dff_B_0BnnNxp55_2;
	wire w_dff_B_Q4fjijCy2_2;
	wire w_dff_B_1mZL0dUv3_2;
	wire w_dff_B_DgRzcWjQ8_2;
	wire w_dff_B_8Hf5oHJP8_2;
	wire w_dff_B_7jsBZXdH1_2;
	wire w_dff_B_vKV2T5HU2_2;
	wire w_dff_B_P7c0iDiS3_2;
	wire w_dff_B_rfCKVihw4_2;
	wire w_dff_B_Nl5YtmKF3_2;
	wire w_dff_B_m6VlBMTA1_2;
	wire w_dff_B_yT0YB5Gr3_2;
	wire w_dff_B_TpIjfnur2_2;
	wire w_dff_B_oVRGp3Sp6_2;
	wire w_dff_B_H3Kw4QSz6_2;
	wire w_dff_B_vbgj8Y442_2;
	wire w_dff_B_zoCGWlAW4_2;
	wire w_dff_B_OBL6shLY8_2;
	wire w_dff_B_QidyfkZl2_2;
	wire w_dff_B_Deppp6vs2_2;
	wire w_dff_B_jhV68JHR4_2;
	wire w_dff_B_39WsdQ8F9_2;
	wire w_dff_B_b4yFNX0X3_2;
	wire w_dff_B_pLRVB3053_2;
	wire w_dff_B_qgVOwGVd2_2;
	wire w_dff_B_zHXr17j86_2;
	wire w_dff_B_i2F67teG0_2;
	wire w_dff_B_O0tNs1sG8_2;
	wire w_dff_B_WRdAaSLj6_2;
	wire w_dff_B_uth7opkF7_2;
	wire w_dff_B_HxE8CPM29_2;
	wire w_dff_B_CRNLJUNR4_2;
	wire w_dff_B_EqhbmTAQ8_2;
	wire w_dff_B_uElOBBtR3_1;
	wire w_dff_B_tS23SFrS2_1;
	wire w_dff_B_yxjpoCoZ8_1;
	wire w_dff_B_Hf9LsCV74_1;
	wire w_dff_B_CRQGqpHS3_1;
	wire w_dff_B_yW36kaxx7_1;
	wire w_dff_B_UqoebJiW5_1;
	wire w_dff_B_BNnp8BfI5_1;
	wire w_dff_B_pquUCSvW2_1;
	wire w_dff_B_3IVVGFyI8_1;
	wire w_dff_B_c1ijh12B7_0;
	wire w_dff_B_9MZ870eG6_0;
	wire w_dff_B_cOu8ZMnh0_0;
	wire w_dff_B_HOFjcere8_0;
	wire w_dff_B_2K5IGgkt5_0;
	wire w_dff_B_OR3YWzNO8_0;
	wire w_dff_B_cmBMnGhB7_0;
	wire w_dff_B_I71mcKFI5_0;
	wire w_dff_B_1RmXZwGf4_0;
	wire w_dff_B_5zLcyl1i2_0;
	wire w_dff_B_OSNyLonq1_1;
	wire w_dff_B_3qIHyXp94_0;
	wire w_dff_B_faRuQwHF6_1;
	wire w_dff_B_Rfv0VYib5_1;
	wire w_dff_B_OcEbHR1J6_1;
	wire w_dff_B_XmbktWK82_1;
	wire w_dff_B_FzkDygg79_1;
	wire w_dff_B_L7PyJuBi0_0;
	wire w_dff_B_OBgwpE531_0;
	wire w_dff_B_hnkeOZ9E8_0;
	wire w_dff_B_WoLNCHGJ7_0;
	wire w_dff_B_0tWcuBVx4_1;
	wire w_dff_B_B1RoABjt7_0;
	wire w_dff_B_d49urWCg8_1;
	wire w_dff_B_GoIcQ4gX1_1;
	wire w_dff_B_jlJHHk7H2_1;
	wire w_dff_B_GzZMZkHb1_1;
	wire w_dff_B_eAJK5NMH4_0;
	wire w_dff_B_0aYxZ4TB8_0;
	wire w_dff_B_LOeSXeM65_0;
	wire w_dff_B_0hoj0HAF7_0;
	wire w_dff_B_4vA8AQV10_1;
	wire w_dff_B_cfkoG1Vt8_1;
	wire w_dff_B_VN3Zm8r59_0;
	wire w_dff_B_rrXjb51L9_0;
	wire w_dff_B_RJRmwaaI4_0;
	wire w_dff_B_QrpMF2wn8_0;
	wire w_dff_B_yAVd0J5N4_0;
	wire w_dff_B_dzW4rya13_0;
	wire w_dff_B_m3XKlcFu2_0;
	wire w_dff_B_79UrQMsw7_0;
	wire w_dff_B_DMptHjD75_0;
	wire w_dff_B_zHUjpYCt9_0;
	wire w_dff_A_qESbXHkL9_0;
	wire w_dff_B_xys7zFVf2_0;
	wire w_dff_B_VXgU1qD85_1;
	wire w_dff_B_vQInOfKG2_1;
	wire w_dff_B_27Kqg1wR5_1;
	wire w_dff_B_t2sPzaDQ7_1;
	wire w_dff_B_Jjg7lsSH3_1;
	wire w_dff_A_7g4YtcYM3_0;
	wire w_dff_A_IBrD16ts4_0;
	wire w_dff_B_DIYmvKh25_0;
	wire w_dff_A_ntrVif4o4_0;
	wire w_dff_A_3E42TCUS7_0;
	wire w_dff_B_hwMRptnW4_0;
	wire w_dff_B_w0VPXIFy1_0;
	wire w_dff_A_KqBYPGeX1_2;
	wire w_dff_B_9Rdq1LAr7_0;
	wire w_dff_B_D0eYQcHv3_1;
	wire w_dff_B_xjXDcDOB3_1;
	wire w_dff_B_LU0uSKLW4_0;
	wire w_dff_A_zDNHOQQv8_1;
	wire w_dff_B_XImWSt9X0_0;
	wire w_dff_B_s4LIctIT6_0;
	wire w_dff_B_NahVCNbJ8_0;
	wire w_dff_B_DKVgnHfT6_0;
	wire w_dff_B_ms9OW3LG2_0;
	wire w_dff_B_yv5Uv9zV8_0;
	wire w_dff_B_MikmA2wz1_0;
	wire w_dff_B_JsIfzC3e0_0;
	wire w_dff_B_V5tqYNKC5_0;
	wire w_dff_B_tSwZ6JNW4_0;
	wire w_dff_B_fgoR0sKj5_0;
	wire w_dff_B_v55vyGEp0_0;
	wire w_dff_B_ljr0nkmZ3_0;
	wire w_dff_B_qaOf45IT1_0;
	wire w_dff_B_eOJ5LWf19_0;
	wire w_dff_B_y2n6IbNe1_0;
	wire w_dff_B_7M8GAmf22_0;
	wire w_dff_B_7T05TSdV1_0;
	wire w_dff_B_aXUeyR8z8_0;
	wire w_dff_B_emtolqjk2_0;
	wire w_dff_B_YnrrQu3O9_0;
	wire w_dff_B_XkSaNPgG2_0;
	wire w_dff_A_DLyspXo41_0;
	wire w_dff_B_uZxkjb4b3_0;
	wire w_dff_A_1UvK5pWl9_0;
	wire w_dff_B_mW1xUD1e1_1;
	wire w_dff_B_OCSbmqRp2_1;
	wire w_dff_B_IVfu9r9O7_0;
	wire w_dff_B_LRbrNLwJ6_0;
	wire w_dff_B_b4hPWs5V6_0;
	wire w_dff_B_6ARVs7Pz3_0;
	wire w_dff_B_DPX5VXjw8_0;
	wire w_dff_B_aRJmjQrm7_0;
	wire w_dff_B_b9rs7CCj0_0;
	wire w_dff_A_izC37lvh5_0;
	wire w_dff_A_m8kotUJU7_2;
	wire w_dff_A_frr3oQK92_2;
	wire w_dff_B_7CQ1qRfY7_1;
	wire w_dff_B_1nQ57FpA3_1;
	wire w_dff_B_W4jNgWOn8_0;
	wire w_dff_A_UYOAdUYd4_0;
	wire w_dff_B_xDZu6nOM6_0;
	wire w_dff_B_wC0aYQQN6_1;
	wire w_dff_A_QYDi2JN64_1;
	wire w_dff_B_XtbsRcWL8_0;
	wire w_dff_B_p0CF3ola8_0;
	wire w_dff_B_V6haeHWd2_0;
	wire w_dff_B_nLQv1jO69_0;
	wire w_dff_B_USso0eYK3_0;
	wire w_dff_B_bOdZZeZW2_0;
	wire w_dff_B_E6bjujDE2_0;
	wire w_dff_B_LNa1SlTM1_1;
	wire w_dff_A_6CCpYkzY5_0;
	wire w_dff_B_89Ljj37K2_0;
	wire w_dff_B_XrjS3DjW1_0;
	wire w_dff_A_WiualOEz8_0;
	wire w_dff_B_ECjMh99R0_0;
	wire w_dff_B_KjMdpMqY3_0;
	wire w_dff_B_RMyClBpC5_0;
	wire w_dff_B_rVfVfTqS2_0;
	wire w_dff_B_0KB6iv9g0_0;
	wire w_dff_B_n52irTqO9_0;
	wire w_dff_B_aZGGt5d13_0;
	wire w_dff_B_xix0vYG33_0;
	wire w_dff_B_7UccTtN25_0;
	wire w_dff_B_BLQwtI809_0;
	wire w_dff_B_jP0SD0ms6_0;
	wire w_dff_B_6C2O4IGp8_0;
	wire w_dff_B_cJHpgVha7_0;
	wire w_dff_B_9QxBzGL67_0;
	wire w_dff_B_NiDkIno62_0;
	wire w_dff_B_Ol64LYX28_0;
	wire w_dff_B_pJwGi2Fx0_0;
	wire w_dff_A_8zHwxbIv2_0;
	wire w_dff_B_IEzZQimm6_0;
	wire w_dff_B_Gu6ly2qK5_0;
	wire w_dff_B_mqK82V5A0_3;
	wire w_dff_B_wtxMmLdS3_3;
	wire w_dff_B_glwqR3mg8_3;
	wire w_dff_B_gDlJkdk08_3;
	wire w_dff_B_w2khVVI92_3;
	wire w_dff_B_wjdCyHom4_3;
	wire w_dff_B_fQo03E7Z0_3;
	wire w_dff_B_3TTKgxND6_3;
	wire w_dff_B_NZMT5rI36_3;
	wire w_dff_B_gfChancj5_3;
	wire w_dff_B_9Vcbey5X0_3;
	wire w_dff_B_ZaKJrtyT2_3;
	wire w_dff_B_Ms6c9Mpd4_3;
	wire w_dff_B_RjQ30wm96_3;
	wire w_dff_B_J1XDUVKt9_3;
	wire w_dff_B_JehOWxDS7_3;
	wire w_dff_B_ZOzfa1qW7_3;
	wire w_dff_B_VtjMCQ885_3;
	wire w_dff_B_gQ0MuVuL1_3;
	wire w_dff_B_V9cJFCcC3_3;
	wire w_dff_B_1Fi2TARt0_3;
	wire w_dff_B_GckgrVIi4_3;
	wire w_dff_B_EHKo0wt72_3;
	wire w_dff_B_ek1NjZSI8_3;
	wire w_dff_B_kHfJAVQO1_3;
	wire w_dff_B_NZfRnSj54_3;
	wire w_dff_B_n6fv7dQd7_3;
	wire w_dff_B_mtwyelTu3_3;
	wire w_dff_B_zDoaU84N9_3;
	wire w_dff_B_SBGlCL4L1_3;
	wire w_dff_B_ZasoEgxn9_3;
	wire w_dff_B_d5C4eOE93_3;
	wire w_dff_B_CCdq6dpQ9_3;
	wire w_dff_B_szjUyLJN5_3;
	wire w_dff_B_dHTH04tO0_0;
	wire w_dff_B_DmaoDgws5_1;
	wire w_dff_B_30yG8BV70_1;
	wire w_dff_B_3XibVL1S4_1;
	wire w_dff_B_OGgz2ypa1_1;
	wire w_dff_B_1VIWuLj67_1;
	wire w_dff_B_OlBKJfqu5_1;
	wire w_dff_B_5Pq49O0v9_1;
	wire w_dff_B_uTJXqnZl7_1;
	wire w_dff_B_Yi9paHfp6_1;
	wire w_dff_B_V9DTpW9O1_1;
	wire w_dff_B_p00NvwVE7_1;
	wire w_dff_B_uLZz6l8T7_1;
	wire w_dff_B_DHuRrOr86_1;
	wire w_dff_B_TO8jfICl5_1;
	wire w_dff_B_LnQ2JwSt4_1;
	wire w_dff_B_nyPLHBkH6_1;
	wire w_dff_B_WTuTZ1VK3_1;
	wire w_dff_B_tykZTdNa8_1;
	wire w_dff_B_jv7ZM1Es7_1;
	wire w_dff_B_ZqqTC3111_1;
	wire w_dff_B_bZ6p0Aom4_1;
	wire w_dff_B_KwgvnGu60_1;
	wire w_dff_B_3rsUJrOM6_1;
	wire w_dff_B_D5qV4Rt37_1;
	wire w_dff_B_2NXbjwEV1_1;
	wire w_dff_B_f42ZBbJr1_1;
	wire w_dff_B_9zhpym730_1;
	wire w_dff_B_blCWD16m3_1;
	wire w_dff_B_lvyyLC6r9_1;
	wire w_dff_B_1nnbtCHl1_1;
	wire w_dff_B_0ZOCEZBN8_1;
	wire w_dff_B_gxOD9HZV4_1;
	wire w_dff_B_iQfw0NuI9_1;
	wire w_dff_B_CBDC1UjX4_1;
	wire w_dff_A_q2N10pwF2_0;
	wire w_dff_A_7dQjV6FX7_0;
	wire w_dff_A_9tvWxzFK6_0;
	wire w_dff_A_3UfxVOXQ3_0;
	wire w_dff_A_H3nBd0GW2_0;
	wire w_dff_A_s1PhLqMt0_0;
	wire w_dff_A_F8FekCd93_0;
	wire w_dff_A_egLKs2CI2_0;
	wire w_dff_A_qM3wT2Px9_0;
	wire w_dff_A_QfczoNKq7_0;
	wire w_dff_A_2FtDRXID7_0;
	wire w_dff_A_7BRGPNsc5_0;
	wire w_dff_A_G0qAYfci7_0;
	wire w_dff_A_PFfIZ3qv7_0;
	wire w_dff_A_g9dEiv1b4_0;
	wire w_dff_A_eP3SQm9B0_0;
	wire w_dff_A_TbXDGri54_0;
	wire w_dff_A_muDG5zJw4_0;
	wire w_dff_A_XvIzNUqa4_0;
	wire w_dff_A_D6QNu48D3_0;
	wire w_dff_A_O5DWwDki5_0;
	wire w_dff_A_j6ndADna4_0;
	wire w_dff_A_VMpfbThm6_0;
	wire w_dff_A_teUtjFgE9_0;
	wire w_dff_A_6jwelbXS9_0;
	wire w_dff_A_5kExzYhZ0_0;
	wire w_dff_A_dG7aaPpF8_0;
	wire w_dff_A_R1RA9pMz7_0;
	wire w_dff_A_lcqFBfw92_0;
	wire w_dff_A_jqKepCQL4_0;
	wire w_dff_A_xp6NkX0r8_0;
	wire w_dff_A_d1LKsnvV4_0;
	wire w_dff_A_Nq8HOIKa7_0;
	wire w_dff_A_bTX9z9f33_0;
	wire w_dff_A_8FTKaedz4_1;
	wire w_dff_A_9ehyRf9E8_0;
	wire w_dff_A_pwqs1dkK6_0;
	wire w_dff_A_njhFUcHG4_1;
	wire w_dff_A_mIsh5nKZ1_1;
	wire w_dff_B_ZU6tV9hk4_3;
	wire w_dff_B_b2tLbgnK7_3;
	wire w_dff_B_HLQVfAld4_3;
	wire w_dff_B_HHiri41I1_3;
	wire w_dff_B_Oh6wSpcm7_3;
	wire w_dff_B_2cH0qWM34_3;
	wire w_dff_B_lDJ72o1Y7_3;
	wire w_dff_B_nSDZTnrN0_3;
	wire w_dff_B_pQZv2jl38_3;
	wire w_dff_B_EFnZsD9u6_3;
	wire w_dff_B_kOYPSxsu0_3;
	wire w_dff_B_1KbbxszE4_3;
	wire w_dff_B_24ZEiQPO2_3;
	wire w_dff_B_mfW44h273_3;
	wire w_dff_B_G63aBnyk4_3;
	wire w_dff_B_0ieYwiaR6_3;
	wire w_dff_B_U6KM1CAw4_3;
	wire w_dff_B_A2IaMNhV9_3;
	wire w_dff_B_7h0BXQlo3_3;
	wire w_dff_B_ezhxHhaj2_3;
	wire w_dff_B_LFVQ22Rs9_3;
	wire w_dff_B_A71FCdqi3_3;
	wire w_dff_B_igpqo0ga5_3;
	wire w_dff_B_VlldJtQx4_3;
	wire w_dff_B_2zhIbBKE7_3;
	wire w_dff_B_L0VxVvAx3_3;
	wire w_dff_B_x0f5if7o1_3;
	wire w_dff_B_tzYvNAlR7_3;
	wire w_dff_B_I55Vq5pF0_3;
	wire w_dff_B_1vIWxpLO5_3;
	wire w_dff_B_JdA71qNN2_3;
	wire w_dff_B_CQ4A5VLN4_3;
	wire w_dff_B_XV3MfLLv5_1;
	wire w_dff_A_IK4xxIxf6_2;
	wire w_dff_B_xYNrf7is3_3;
	wire w_dff_B_BXBFnrXY1_3;
	wire w_dff_B_9Rqn8m6M7_3;
	wire w_dff_B_JENYrdUh5_3;
	wire w_dff_B_w9mgrB452_3;
	wire w_dff_B_OWfkJWGJ0_3;
	wire w_dff_B_7ti0uLSR2_3;
	wire w_dff_B_4iREe2qE0_3;
	wire w_dff_B_VwsYQFrQ9_3;
	wire w_dff_B_SjaM4DmG8_3;
	wire w_dff_B_lsV7hKWi3_3;
	wire w_dff_B_Ks4Iu0u74_3;
	wire w_dff_B_IQakFRgW9_3;
	wire w_dff_B_8JLSYnvn7_3;
	wire w_dff_B_kMDuHP7i0_3;
	wire w_dff_B_hty7O9MI2_3;
	wire w_dff_B_PnJUayvo0_3;
	wire w_dff_B_QhQzerc22_3;
	wire w_dff_B_Tks1g2cz1_3;
	wire w_dff_B_mxagUY3t3_3;
	wire w_dff_B_fCeMwCYK0_3;
	wire w_dff_B_2goDnZLM2_3;
	wire w_dff_B_7ogavWEc8_3;
	wire w_dff_B_WgSmYDol3_3;
	wire w_dff_B_2w72tr4c5_3;
	wire w_dff_B_rZoPdTTN8_3;
	wire w_dff_B_kRYUO83D3_3;
	wire w_dff_B_pscKGlGo7_3;
	wire w_dff_B_AwBuAuDI2_3;
	wire w_dff_B_wi1ZHICE9_3;
	wire w_dff_B_hbKJ8em88_3;
	wire w_dff_B_qfDuvjXL3_3;
	wire w_dff_B_i0IAEUFQ6_3;
	wire w_dff_B_cbk2BWzk1_3;
	wire w_dff_B_iwCZEiy92_1;
	wire w_dff_B_lwAhtTXJ6_1;
	wire w_dff_B_mvZEa8Yb1_1;
	wire w_dff_B_rNLNxwjw9_1;
	wire w_dff_B_0RPQMNlp9_1;
	wire w_dff_B_ItB9DSYK4_1;
	wire w_dff_B_nY6fBif09_1;
	wire w_dff_B_CzZm3sKM5_0;
	wire w_dff_B_IJqXK7xy4_0;
	wire w_dff_B_CQOPHmxj9_0;
	wire w_dff_B_U6uUJYMY4_0;
	wire w_dff_B_CjtaEvzf9_0;
	wire w_dff_B_YU0fqcTE2_0;
	wire w_dff_B_ITbNaMFb3_0;
	wire w_dff_B_CmeW8RsZ9_0;
	wire w_dff_B_n5Wlgp9y2_0;
	wire w_dff_B_maMs4OPL4_0;
	wire w_dff_B_wWZT8jzU8_0;
	wire w_dff_B_AulaXLNa1_0;
	wire w_dff_B_ksX8i8EM9_0;
	wire w_dff_B_5QgMdvmu0_0;
	wire w_dff_B_Kl87ZlXS5_0;
	wire w_dff_B_njTeZRjP2_0;
	wire w_dff_B_heeQ53XN0_0;
	wire w_dff_B_2uSCymEX3_0;
	wire w_dff_B_Dlngj57s1_0;
	wire w_dff_B_jplcTCD69_0;
	wire w_dff_B_JHL2yQWh1_0;
	wire w_dff_B_WStrZEZs9_0;
	wire w_dff_B_gYFDldi45_0;
	wire w_dff_B_0WgCKNXn7_0;
	wire w_dff_B_rTWBlQkd3_0;
	wire w_dff_B_rJHql58A8_0;
	wire w_dff_B_jzMC9Zpr9_0;
	wire w_dff_B_NQhUAtfH7_0;
	wire w_dff_B_jEpyes7S5_0;
	wire w_dff_B_xtUd53kq0_0;
	wire w_dff_B_QKsJMYwe8_0;
	wire w_dff_B_mN2iOQhY1_0;
	wire w_dff_B_ZIMfv6Ft0_0;
	wire w_dff_B_mQHKKZk18_0;
	wire w_dff_B_KQMtYEJ24_0;
	wire w_dff_B_voiF3B4n6_0;
	wire w_dff_B_GZw9fVJM1_0;
	wire w_dff_B_oBeFwSQN7_0;
	wire w_dff_B_3Bok2QBk2_0;
	wire w_dff_B_GwYFLE550_0;
	wire w_dff_B_YcQLb1wr8_0;
	wire w_dff_B_4e0S8qxo6_0;
	wire w_dff_B_entIfyXW2_0;
	wire w_dff_B_8XGtxMwR9_0;
	wire w_dff_B_a0nVU4kh9_0;
	wire w_dff_B_QxABoxwe4_0;
	wire w_dff_B_Ldyh76fx6_0;
	wire w_dff_B_F4gtk9VZ6_0;
	wire w_dff_B_Jr8WZMTC0_0;
	wire w_dff_B_hmSVbWko1_0;
	wire w_dff_B_5kx1C4oU1_0;
	wire w_dff_B_ib85P0Do7_0;
	wire w_dff_B_4iHWD0pp4_0;
	wire w_dff_B_HRGL5uT05_0;
	wire w_dff_B_4jen2nQk7_0;
	wire w_dff_B_dtd8IRAi8_0;
	wire w_dff_B_9mp0lpax4_0;
	wire w_dff_B_BhWBXVsX9_0;
	wire w_dff_B_eN8HR6yF0_0;
	wire w_dff_B_4aYXOa487_0;
	wire w_dff_B_6OTOHNuf9_0;
	wire w_dff_B_fg5nQDsy0_0;
	wire w_dff_B_adcEbKvM5_0;
	wire w_dff_B_jhGPRTPu7_0;
	wire w_dff_B_cVQd0kbu9_0;
	wire w_dff_B_4junVqrn3_0;
	wire w_dff_B_HQvhTqdr8_0;
	wire w_dff_B_RDVU7uQd1_0;
	wire w_dff_B_rUyNkDps8_0;
	wire w_dff_B_ifkGSxQ64_0;
	wire w_dff_B_06H5CUu42_0;
	wire w_dff_B_KBTEMHY11_0;
	wire w_dff_B_JQAzfofo1_1;
	wire w_dff_B_MzXGszdx7_0;
	wire w_dff_B_pZjI0ZAQ9_0;
	wire w_dff_B_m0O3PEqb1_0;
	wire w_dff_B_wnS3s8PN9_0;
	wire w_dff_B_zVPfz9jM0_1;
	wire w_dff_B_LIpDOmxh0_1;
	wire w_dff_B_yNI3N9J80_0;
	wire w_dff_B_pBgev0qp1_0;
	wire w_dff_B_DBz0h19I2_0;
	wire w_dff_B_ykHznQu92_0;
	wire w_dff_A_OPGzQBy28_0;
	wire w_dff_A_sdWPMgqU9_0;
	wire w_dff_A_ZAU6hFYu9_0;
	wire w_dff_A_877u7CnR6_0;
	wire w_dff_A_Kx8IwE3u5_2;
	wire w_dff_A_Y4qbgTZr0_2;
	wire w_dff_A_WGaGkLAH1_2;
	wire w_dff_A_AKv7wvjL7_1;
	wire w_dff_A_CzCbI9Ji8_2;
	wire w_dff_A_qD5rT4n13_2;
	wire w_dff_A_D8tpZV5o0_2;
	wire w_dff_A_3KaTgZGL4_2;
	wire w_dff_A_RAPm4VBC9_2;
	wire w_dff_A_yBzZvtQJ0_2;
	wire w_dff_A_wGwfwR1B1_2;
	wire w_dff_A_LuJYgc4V1_2;
	wire w_dff_A_X7GV8CaJ3_2;
	wire w_dff_A_G3RKkQxr8_2;
	wire w_dff_A_3niIIym51_2;
	wire w_dff_A_Xsw30ZU44_2;
	wire w_dff_A_X3eG48iL9_2;
	wire w_dff_A_sVAdGYO23_2;
	wire w_dff_A_dapvPtw94_2;
	wire w_dff_A_5PYuZQCK5_2;
	wire w_dff_A_zGzwXonD2_2;
	wire w_dff_A_5JlJnPZS8_2;
	wire w_dff_A_jZ4S0nXB2_2;
	wire w_dff_A_ZzzLr51u8_2;
	wire w_dff_A_uDXqbVQo7_2;
	wire w_dff_B_5FSA70jg8_3;
	wire w_dff_B_QY12PvqX4_3;
	wire w_dff_B_h8YYfvGs6_3;
	wire w_dff_B_HCiw0wR69_0;
	wire w_dff_B_v9P2Ef6F8_0;
	wire w_dff_B_tDajx7HY7_0;
	wire w_dff_B_SdnNc85e9_0;
	wire w_dff_B_ZnjrzCG81_0;
	wire w_dff_B_JGBqApfD5_0;
	wire w_dff_B_hl2s3UDQ1_0;
	wire w_dff_B_poRSKr6K7_0;
	wire w_dff_B_wlYSBYug4_0;
	wire w_dff_B_Y8LRYdsQ7_0;
	wire w_dff_B_YYdb0WtZ2_0;
	wire w_dff_B_AfLOuRbE6_0;
	wire w_dff_B_Guu9W5lT3_0;
	wire w_dff_B_Hh445aZ72_0;
	wire w_dff_B_MNXvU4Yq5_0;
	wire w_dff_B_GCFSsGMy4_0;
	wire w_dff_B_Oqzd83765_0;
	wire w_dff_B_YcZj1Ee59_0;
	wire w_dff_B_CYuVarN33_0;
	wire w_dff_B_19gLca623_1;
	wire w_dff_B_oVKeCFhR0_0;
	wire w_dff_B_p3iDl0LL3_0;
	wire w_dff_B_pA3M7hlw5_0;
	wire w_dff_B_nXw0z1C79_0;
	wire w_dff_B_RmEVGv169_0;
	wire w_dff_B_Q2TMaCkN0_0;
	wire w_dff_B_ioWVW5cq5_0;
	wire w_dff_B_zUMtOvXg5_0;
	wire w_dff_B_dTYmxbU09_0;
	wire w_dff_B_m2bOGnqx5_0;
	wire w_dff_B_vYd0JbmH8_0;
	wire w_dff_B_Exw3ZbQ40_0;
	wire w_dff_B_bbqsGEX53_0;
	wire w_dff_B_dgleFurm4_0;
	wire w_dff_B_HSpi26eR3_0;
	wire w_dff_B_WPVgTrKh4_0;
	wire w_dff_B_SliFyK364_0;
	wire w_dff_B_DDPPv2SI4_0;
	wire w_dff_B_a64E0SVz4_0;
	wire w_dff_B_eBmcZyFn2_0;
	wire w_dff_B_XqyKNomX4_0;
	wire w_dff_B_vnvmDqhx9_0;
	wire w_dff_B_JOn9JoTf0_0;
	wire w_dff_B_OWbI6Hs37_1;
	wire w_dff_A_zDaaqjFq9_1;
	wire w_dff_A_bIs27t4o1_1;
	wire w_dff_A_jSGZbhrz3_1;
	wire w_dff_A_igY0Jrt43_1;
	wire w_dff_A_HZ0CV9l05_1;
	wire w_dff_A_UQWJPadr1_1;
	wire w_dff_A_Y6r6FIxN5_1;
	wire w_dff_A_px2Qhygn8_1;
	wire w_dff_A_ikDAEHbm8_1;
	wire w_dff_A_HuNo3HCd3_1;
	wire w_dff_A_deX5kzSy0_1;
	wire w_dff_A_xgkS52bQ8_1;
	wire w_dff_A_sefBpE1U3_1;
	wire w_dff_A_cC0Afoxr2_1;
	wire w_dff_A_fJZpjdl66_1;
	wire w_dff_A_Vm4uW51n2_1;
	wire w_dff_A_Gr6F1muv4_1;
	wire w_dff_A_YlEPGzQx4_1;
	wire w_dff_A_9s3g67sC1_1;
	wire w_dff_A_zxHTcwwh6_1;
	wire w_dff_A_KjWqLPWo4_1;
	wire w_dff_A_rwnUHiRA0_1;
	wire w_dff_A_OdH2NJne7_1;
	wire w_dff_A_8iBegAz22_1;
	wire w_dff_A_3hTYa1n72_1;
	wire w_dff_A_IBQBu9xf7_0;
	wire w_dff_A_1wkanVuV3_0;
	wire w_dff_B_yp0UUsgy3_2;
	wire w_dff_B_HhkjUhcZ3_2;
	wire w_dff_B_REaPs5VA1_2;
	wire w_dff_B_bJorngyd9_2;
	wire w_dff_B_M4dntbBX2_0;
	wire w_dff_B_Uh9VKXdS1_0;
	wire w_dff_B_LscSTxLd5_0;
	wire w_dff_B_gkVVzPnk3_0;
	wire w_dff_B_vtGtHBCI9_0;
	wire w_dff_B_8BqA5M6p5_0;
	wire w_dff_B_js9pqa8p6_0;
	wire w_dff_B_F4FwegUn5_0;
	wire w_dff_B_pYsChYHg4_0;
	wire w_dff_B_FpcoZgm93_0;
	wire w_dff_B_5UE2RiJF5_0;
	wire w_dff_B_Rwj7kJJZ2_0;
	wire w_dff_B_hYHRqDqo2_0;
	wire w_dff_B_wVCtVCBj2_0;
	wire w_dff_B_kKCJNrL00_0;
	wire w_dff_B_1pfcmRyW4_0;
	wire w_dff_B_zCPKfWUA2_0;
	wire w_dff_B_PBm2BaFD9_0;
	wire w_dff_B_uU2xQCE56_0;
	wire w_dff_A_5gGzOLJl8_1;
	wire w_dff_A_YmHdbC4Z9_1;
	wire w_dff_A_b2PEHwBn9_1;
	wire w_dff_A_4MNvW2gx6_1;
	wire w_dff_A_14FdSpXK1_1;
	wire w_dff_A_4s24rNNu7_1;
	wire w_dff_A_XIhn4XGv7_1;
	wire w_dff_A_zb1yipxd6_1;
	wire w_dff_A_LfnEtyXp6_1;
	wire w_dff_A_VHqQA4S40_1;
	wire w_dff_A_2r4QNp145_1;
	wire w_dff_A_Z0u7eusa9_1;
	wire w_dff_A_wBacaGYp0_1;
	wire w_dff_A_sqLm0VZW5_1;
	wire w_dff_A_GCDSgynG5_1;
	wire w_dff_A_QjUPw4BJ8_1;
	wire w_dff_A_kvK8H9oF0_1;
	wire w_dff_A_Ip0fJTsx9_1;
	wire w_dff_A_4EbeUOuD3_1;
	wire w_dff_A_HhEuQ8gq0_1;
	wire w_dff_A_8rcwYPhX6_1;
	wire w_dff_A_EfqEAZC60_0;
	wire w_dff_A_vPrYrtUM3_0;
	wire w_dff_A_kFKHFjBJ0_0;
	wire w_dff_A_MgolSiJF5_0;
	wire w_dff_A_z3DODmv08_0;
	wire w_dff_A_Bu2R6wKw1_0;
	wire w_dff_A_jHGQd42d4_0;
	wire w_dff_A_IOekg5D68_0;
	wire w_dff_A_vnP7HZqA6_0;
	wire w_dff_A_RnAshcBa2_0;
	wire w_dff_A_I9Yk1Ke74_0;
	wire w_dff_A_vsYzurLH9_0;
	wire w_dff_A_iXw4laOV6_0;
	wire w_dff_A_gwCZCdB63_0;
	wire w_dff_A_zF9GTniw8_0;
	wire w_dff_A_veFTmxyv3_0;
	wire w_dff_A_m1cyPN2n6_0;
	wire w_dff_A_dUxSFAs18_0;
	wire w_dff_A_FCcBznTD9_0;
	wire w_dff_A_OEP0ppCs1_0;
	wire w_dff_A_MnDcgg263_0;
	wire w_dff_B_rg8UwGAd5_1;
	wire w_dff_B_iQSqXYyW4_1;
	wire w_dff_B_ynPXtwQx8_1;
	wire w_dff_B_V1qUrEA61_1;
	wire w_dff_B_CZwh5s0v2_1;
	wire w_dff_B_v7OCEp2r2_1;
	wire w_dff_B_OTYgK7iz0_1;
	wire w_dff_A_D1dZChUW1_1;
	wire w_dff_A_Sz70AeEL0_1;
	wire w_dff_A_YpLn6Q9P6_1;
	wire w_dff_A_NoKSTi4d3_1;
	wire w_dff_A_zMO4Xgwz1_1;
	wire w_dff_A_KHAYfGor3_1;
	wire w_dff_B_IkFwriAd7_0;
	wire w_dff_B_9usL6MWy7_0;
	wire w_dff_B_HHDruGVr0_0;
	wire w_dff_B_WLMEmKxs3_0;
	wire w_dff_B_XsDpzbJf8_0;
	wire w_dff_B_xi4K8tC28_0;
	wire w_dff_B_sY5i52Hl1_0;
	wire w_dff_B_joWPS9LO5_0;
	wire w_dff_B_hY2aYXSu0_0;
	wire w_dff_B_uqJpKo9i4_0;
	wire w_dff_B_NNmZswSL9_0;
	wire w_dff_B_7OObS6FG5_0;
	wire w_dff_B_hBJ7awXS7_0;
	wire w_dff_B_2INUkVPi7_0;
	wire w_dff_B_BhkEQldm1_0;
	wire w_dff_B_aOla3Zsa1_0;
	wire w_dff_B_ttYZu3Rs4_0;
	wire w_dff_B_To1HMDCp2_0;
	wire w_dff_B_IiTdSLe73_1;
	wire w_dff_B_LAE2XKGt9_0;
	wire w_dff_B_uytsovJ87_0;
	wire w_dff_B_ejmQ3Efr8_0;
	wire w_dff_B_qP1Nuk7T4_0;
	wire w_dff_B_GdGqE3hQ0_0;
	wire w_dff_B_7sNWLq7L1_0;
	wire w_dff_B_PdBQmugf1_0;
	wire w_dff_B_qLIsIgXK4_0;
	wire w_dff_B_p90kH7vl4_0;
	wire w_dff_A_YDtMt7ws4_2;
	wire w_dff_A_T1F6XDXd7_0;
	wire w_dff_A_5Nhhcxai6_0;
	wire w_dff_A_y9fJLhst5_0;
	wire w_dff_A_ZAY3sdbH0_1;
	wire w_dff_A_stjFbjlk7_0;
	wire w_dff_B_6cDj0TJ59_2;
	wire w_dff_B_DdHJJIrb7_2;
	wire w_dff_B_2lLYqGG66_2;
	wire w_dff_B_6DXf3yZk1_2;
	wire w_dff_B_8QKTm6sM2_2;
	wire w_dff_B_FWWtzdEu6_2;
	wire w_dff_B_TW6PJP5p4_2;
	wire w_dff_B_zsXdLKoc7_2;
	wire w_dff_B_Eio5xOfu0_1;
	wire w_dff_A_TS9rw5RI0_0;
	wire w_dff_A_5c0RCyZl8_0;
	wire w_dff_A_1BRvXLhZ3_2;
	wire w_dff_A_dHJt4ITd3_2;
	wire w_dff_A_J3NkEjqI6_2;
	wire w_dff_A_mN4Y5ULW5_0;
	wire w_dff_A_ryf5ao1F6_2;
	wire w_dff_A_tK7K9Fkw6_2;
	wire w_dff_A_OMEH5hXN6_2;
	wire w_dff_A_LQdGDyaf3_0;
	wire w_dff_A_fc7Tr0NP2_2;
	wire w_dff_B_rRADiHUb3_1;
	wire w_dff_B_TgN42e2d3_1;
	wire w_dff_B_yU4SBeVL3_1;
	wire w_dff_B_Dor57Wdg2_1;
	wire w_dff_B_sSf5Vc6P5_1;
	wire w_dff_B_65cDIrOJ4_1;
	wire w_dff_B_rnc7HdhT9_1;
	wire w_dff_B_JlSU60wd0_1;
	wire w_dff_A_vv1u85RS6_0;
	wire w_dff_A_I1sQzuSs6_0;
	wire w_dff_A_ShlfCCAp3_0;
	wire w_dff_A_au2HequK3_0;
	wire w_dff_A_XYNYSsfo3_0;
	wire w_dff_A_lCo0J2P36_0;
	wire w_dff_A_3VcDMBVU6_0;
	wire w_dff_A_YkEiM8el4_0;
	wire w_dff_A_zFoCX1fE6_0;
	wire w_dff_A_lGEjnJqf7_0;
	wire w_dff_A_B4Uvi9wh0_0;
	wire w_dff_A_WIvLSdsG7_0;
	wire w_dff_A_86Hw0UjG9_0;
	wire w_dff_A_wCl0FIRY7_0;
	wire w_dff_A_1HXuwVzF8_0;
	wire w_dff_A_7w42ZpaP5_0;
	wire w_dff_A_XnA6JFnX3_0;
	wire w_dff_A_Ofx3yYQi7_0;
	wire w_dff_A_XV5Ix2l99_0;
	wire w_dff_A_o4RdDaLv8_0;
	wire w_dff_A_FqsXpHRE5_0;
	wire w_dff_A_4SfiI0QB4_0;
	wire w_dff_A_g8uNbSA76_0;
	wire w_dff_A_tt9k7NbA3_0;
	wire w_dff_A_sXSo4oBX0_0;
	wire w_dff_A_rFX5MMDq0_0;
	wire w_dff_A_O4x9BQG24_0;
	wire w_dff_A_Bazhx6cq3_0;
	wire w_dff_A_W95FR43n2_0;
	wire w_dff_A_f4rNf0jd1_0;
	wire w_dff_A_uH96gR3q6_2;
	wire w_dff_A_BqSshFE30_2;
	wire w_dff_A_73TXpqed6_2;
	wire w_dff_A_GpE9zX9c1_2;
	wire w_dff_A_Cek6xykY5_2;
	wire w_dff_B_KbplI2i71_1;
	wire w_dff_B_8DgCpoAW7_1;
	wire w_dff_B_zR2UjtQK0_1;
	wire w_dff_B_oHTIevSM9_1;
	wire w_dff_B_mcCwunEQ9_1;
	wire w_dff_B_9OZxQn1N4_1;
	wire w_dff_B_AK0tmjSl2_1;
	wire w_dff_B_MHuP8Hc85_1;
	wire w_dff_B_SGl2lSaj0_1;
	wire w_dff_B_6E6gNwgW2_1;
	wire w_dff_B_3psTi4QW0_1;
	wire w_dff_B_RIBcg9Vm5_1;
	wire w_dff_B_pvs0lKTW6_1;
	wire w_dff_B_kMzW6HNz0_1;
	wire w_dff_B_vvt3UTDS2_1;
	wire w_dff_B_8K8sOztk2_1;
	wire w_dff_B_lqwY6KzP5_1;
	wire w_dff_B_LMwXuSfa5_1;
	wire w_dff_B_9wMV4Wy31_1;
	wire w_dff_B_zAJOaNse4_1;
	wire w_dff_B_TOfUppsf6_1;
	wire w_dff_B_0NfPig3K9_1;
	wire w_dff_B_G1p4miaA2_1;
	wire w_dff_B_arAO3LTb2_1;
	wire w_dff_B_h2ZseJna0_1;
	wire w_dff_B_6Xsr2TIy5_1;
	wire w_dff_B_Ubk3OkEW4_1;
	wire w_dff_B_VNQEIJ2B7_1;
	wire w_dff_B_CCgQi8H14_1;
	wire w_dff_B_Oav8gulg4_1;
	wire w_dff_B_RQNtAc8l7_1;
	wire w_dff_B_ZIFG6nf48_0;
	wire w_dff_B_VPTJctPF0_0;
	wire w_dff_B_filD7DCD1_0;
	wire w_dff_B_oFAVvcJc8_0;
	wire w_dff_B_OwzwZ3Pz2_0;
	wire w_dff_B_ZfF76pED0_0;
	wire w_dff_B_zsKa5CVc3_0;
	wire w_dff_B_Jf18p4N64_0;
	wire w_dff_B_v77hwnGl8_0;
	wire w_dff_B_PiQIMHru8_0;
	wire w_dff_B_few3mHEU3_0;
	wire w_dff_B_CGo767pF6_0;
	wire w_dff_B_KQYFpcZO3_0;
	wire w_dff_B_yJ0NXdhk6_0;
	wire w_dff_B_HHrZ6Q6R0_0;
	wire w_dff_B_1uPdd0nj8_0;
	wire w_dff_B_EttT5PON4_0;
	wire w_dff_B_nDchxqvr3_0;
	wire w_dff_B_EO5KVPZn6_0;
	wire w_dff_B_kwGuXUXQ2_0;
	wire w_dff_B_y6jLaFWv5_1;
	wire w_dff_B_fY56sq2l1_1;
	wire w_dff_B_BiUg6YDy3_0;
	wire w_dff_B_u2tlrm4O5_0;
	wire w_dff_B_W66BIxzs5_0;
	wire w_dff_B_e1JuA95y3_0;
	wire w_dff_B_INzzAuzd4_0;
	wire w_dff_A_FajkBpHE7_1;
	wire w_dff_A_UBZNhFsc9_1;
	wire w_dff_A_sSjpLx367_1;
	wire w_dff_A_l0oPRfmY3_1;
	wire w_dff_A_BmyqDzfJ2_1;
	wire w_dff_A_8eK0kAel7_1;
	wire w_dff_A_wcfNUdRJ4_1;
	wire w_dff_A_7pTc6CZs1_1;
	wire w_dff_A_TqpQzs9O1_1;
	wire w_dff_A_IOVYzYAs3_1;
	wire w_dff_A_Oc2YygRX0_1;
	wire w_dff_A_S6VsueXs1_1;
	wire w_dff_A_Z5MDXOdj9_1;
	wire w_dff_A_l8Z1Tr2Y5_1;
	wire w_dff_A_1KjP9csF4_1;
	wire w_dff_A_3U1leG9n6_1;
	wire w_dff_A_V2tacE9T4_1;
	wire w_dff_A_XroujTcU7_1;
	wire w_dff_A_XiW6w5JV9_1;
	wire w_dff_A_OCUELDqV1_1;
	wire w_dff_A_xIq35Qv42_1;
	wire w_dff_A_o6T7RTMj2_1;
	wire w_dff_A_hTFS2Vpd0_1;
	wire w_dff_A_QtcHqgc40_1;
	wire w_dff_A_WB2CvrJW5_1;
	wire w_dff_B_JiERR1Iq0_0;
	wire w_dff_B_2ARvBBtH9_0;
	wire w_dff_B_qzHqw6h73_0;
	wire w_dff_B_xnTx0TVi2_1;
	wire w_dff_B_lP1eYBD99_1;
	wire w_dff_B_y1FHGEko7_1;
	wire w_dff_B_57MVZArM1_1;
	wire w_dff_B_azEqYxyT5_1;
	wire w_dff_A_f8cSmmCn9_1;
	wire w_dff_A_35OU87DK2_1;
	wire w_dff_A_RgOlcgrK5_1;
	wire w_dff_A_wHuEb2lj3_1;
	wire w_dff_A_KFaKO4vd4_1;
	wire w_dff_A_XQnY0Vo61_1;
	wire w_dff_A_nZPq9cQh5_1;
	wire w_dff_A_hXUpu4BD6_1;
	wire w_dff_A_6bLof3eb8_1;
	wire w_dff_A_gBSzMHpX3_1;
	wire w_dff_A_JhXtz3Ss1_1;
	wire w_dff_A_3SwhL6qs9_1;
	wire w_dff_A_SuPxILcn6_1;
	wire w_dff_A_QeM17DCO2_1;
	wire w_dff_A_UZfkibCq1_1;
	wire w_dff_A_wG4CRCBj7_1;
	wire w_dff_A_HQZuX8Zv8_1;
	wire w_dff_A_3LeyG6A52_1;
	wire w_dff_A_W3yrwK1G2_1;
	wire w_dff_A_cTh2FNYV6_1;
	wire w_dff_A_UJXvJUo44_1;
	wire w_dff_A_TWZkus282_1;
	wire w_dff_B_a3SJFK7E1_2;
	wire w_dff_A_9CY54BSs3_0;
	wire w_dff_A_XHzGi9Jr4_0;
	wire w_dff_A_22JjTXqe3_0;
	wire w_dff_A_cr1hPzEY8_0;
	wire w_dff_A_1E9O2vqX7_0;
	wire w_dff_B_FyQNE8XS5_1;
	wire w_dff_B_hMyXcZCq6_1;
	wire w_dff_B_mYAMaaH61_1;
	wire w_dff_B_KfqJFjZz0_1;
	wire w_dff_B_2XDJCDok9_1;
	wire w_dff_B_ocGeuNd14_1;
	wire w_dff_B_tQ5mKweV1_1;
	wire w_dff_B_vSOESnuB6_1;
	wire w_dff_B_4vwUtX5y7_1;
	wire w_dff_B_vonLHBY13_1;
	wire w_dff_B_83Vkj7219_1;
	wire w_dff_B_7yZszsJV6_1;
	wire w_dff_B_NxWmUapD7_1;
	wire w_dff_B_KH17Yc3t7_1;
	wire w_dff_B_JVgoryDw9_1;
	wire w_dff_B_jYNCGmAX8_1;
	wire w_dff_B_L0Q5T17N2_1;
	wire w_dff_B_1CLltA5J4_1;
	wire w_dff_B_Gx05KMYm4_1;
	wire w_dff_B_q8x3KuWt4_1;
	wire w_dff_B_9SzYDlrH2_1;
	wire w_dff_B_Kfiz4VTJ4_1;
	wire w_dff_B_dckUumh78_1;
	wire w_dff_B_k78dmU431_1;
	wire w_dff_B_hGk3aXMW6_1;
	wire w_dff_B_XOV5dNNa5_1;
	wire w_dff_B_2KWgNVkv5_1;
	wire w_dff_B_KmzGxk4w4_1;
	wire w_dff_B_UuxtBApE6_1;
	wire w_dff_B_kgdgUzU63_1;
	wire w_dff_B_mjnOfVEj5_1;
	wire w_dff_B_jjJdIxsd7_1;
	wire w_dff_B_lspRqeE73_1;
	wire w_dff_B_gwTe6ssh4_1;
	wire w_dff_B_Md7ixU3w3_1;
	wire w_dff_B_wuHD7whs2_1;
	wire w_dff_B_0UrAc8Nk5_1;
	wire w_dff_B_6aehAtxn9_1;
	wire w_dff_B_kLm88onJ5_1;
	wire w_dff_B_XbUdJMHW0_1;
	wire w_dff_B_Jgu0j0xR7_1;
	wire w_dff_B_FZiKhB0O5_1;
	wire w_dff_B_WfgI7hsW9_1;
	wire w_dff_B_sP7NPzcD3_1;
	wire w_dff_B_LFetKh0N2_1;
	wire w_dff_B_s1j3VRCI0_1;
	wire w_dff_B_JQFZhxoG3_1;
	wire w_dff_B_KCDDsFAB6_1;
	wire w_dff_B_wkaufNKd8_1;
	wire w_dff_B_6ityTnxH3_1;
	wire w_dff_B_nc4DORdT0_1;
	wire w_dff_B_t5VmvgvV9_1;
	wire w_dff_B_Wxi7Li0q3_1;
	wire w_dff_B_iItRIaRy7_1;
	wire w_dff_B_6gFcWADp7_1;
	wire w_dff_B_NFuqLFRS5_1;
	wire w_dff_B_e1Nbm4jB5_1;
	wire w_dff_B_BE6TCiES2_1;
	wire w_dff_B_rEz2ctfc6_1;
	wire w_dff_B_v5nlcT5a1_1;
	wire w_dff_B_gSYitMou4_1;
	wire w_dff_B_uUUtTRDO4_1;
	wire w_dff_B_i8HOPdLC2_1;
	wire w_dff_B_k7zfV01k8_1;
	wire w_dff_B_YUnwslQ83_1;
	wire w_dff_B_GX9SKCAI0_1;
	wire w_dff_B_RbCXqxy93_1;
	wire w_dff_B_xweBRsBM1_1;
	wire w_dff_B_7dwATRM32_1;
	wire w_dff_B_exD9w7Jj8_1;
	wire w_dff_B_X8LozdNv4_1;
	wire w_dff_B_wFA1FKeK2_1;
	wire w_dff_B_tKBrGSFa3_1;
	wire w_dff_B_LwvcJn2Y5_1;
	wire w_dff_B_1mrE3lYF9_1;
	wire w_dff_B_qtVtrj7r8_1;
	wire w_dff_B_ZsmpZskx1_1;
	wire w_dff_B_Le4P70Ot2_1;
	wire w_dff_B_jB6DICeT0_1;
	wire w_dff_B_ycODkcrf4_1;
	wire w_dff_B_IYIgiYo72_1;
	wire w_dff_B_hJRc0dPJ1_1;
	wire w_dff_B_iV4lKNpO6_1;
	wire w_dff_B_JtWnfbAq1_1;
	wire w_dff_B_yDGNHflk5_1;
	wire w_dff_B_A6e4ZRcf8_1;
	wire w_dff_B_xJrEr7jx1_1;
	wire w_dff_B_OdY8VVL85_1;
	wire w_dff_B_2D0Xl9bl6_1;
	wire w_dff_B_hxBAdlmy9_1;
	wire w_dff_B_Hyo3IW770_1;
	wire w_dff_B_HyuUShvg7_1;
	wire w_dff_B_618PvWUD2_1;
	wire w_dff_B_mGx99hM97_1;
	wire w_dff_B_oARdvx0O9_1;
	wire w_dff_B_jUTm8CVk7_1;
	wire w_dff_B_QDCFzGIp4_1;
	wire w_dff_B_HLGIwBVv4_1;
	wire w_dff_B_aU46LyhX4_1;
	wire w_dff_B_b3E2JgJ75_1;
	wire w_dff_B_nzMu3MQf1_1;
	wire w_dff_B_Na4DGaBP4_1;
	wire w_dff_B_0DGm8ZVX2_1;
	wire w_dff_B_wjyj0WKK4_1;
	wire w_dff_B_8MXny79A3_1;
	wire w_dff_B_rXONjn159_1;
	wire w_dff_B_kFcP249J9_1;
	wire w_dff_B_sjs9PK3f1_1;
	wire w_dff_B_mQgQ7USW3_1;
	wire w_dff_B_pBpIIhvz7_1;
	wire w_dff_B_67vwr24W4_1;
	wire w_dff_B_Ccl6R05j0_1;
	wire w_dff_B_YiFqbGVX2_1;
	wire w_dff_B_SMa0Ue6V0_1;
	wire w_dff_B_m25LymCS0_1;
	wire w_dff_B_1FZOIzhJ1_1;
	wire w_dff_B_LoQlbB2L8_1;
	wire w_dff_B_VmyuVrLh6_1;
	wire w_dff_B_nO889iOG1_1;
	wire w_dff_B_Ywhl824d5_1;
	wire w_dff_B_mDKbaS6F0_1;
	wire w_dff_B_xwiRNtQZ0_1;
	wire w_dff_B_vkejMAam6_1;
	wire w_dff_B_5A6KfDUS4_1;
	wire w_dff_B_MRxhsvNs4_1;
	wire w_dff_B_5YEcKngC6_1;
	wire w_dff_B_iNFNxHr21_1;
	wire w_dff_B_AbJ7Z0fu5_1;
	wire w_dff_B_KAjw9nXX1_1;
	wire w_dff_B_UXF6fFBc8_1;
	wire w_dff_B_omzyU4fI5_1;
	wire w_dff_B_k1nw84Sn9_1;
	wire w_dff_B_PDI63GOE2_1;
	wire w_dff_B_vobuiUjm5_1;
	wire w_dff_B_c6slsYjW3_1;
	wire w_dff_B_CjjnwJBo7_1;
	wire w_dff_B_BQ9Dt4NL1_1;
	wire w_dff_B_DyYlIAEO6_1;
	wire w_dff_B_FIIhOPuE1_1;
	wire w_dff_B_ia5UFewF2_1;
	wire w_dff_B_aIuIpuQN4_1;
	wire w_dff_B_RzXcr7NG3_1;
	wire w_dff_B_5dSlsuGz1_1;
	wire w_dff_B_wTcfhqba2_1;
	wire w_dff_B_S7MtSNHF6_1;
	wire w_dff_B_x4A1eFdW1_1;
	wire w_dff_B_iue93fgv9_1;
	wire w_dff_B_MFWxDZjZ4_1;
	wire w_dff_B_AIGBwvCy8_1;
	wire w_dff_B_tHIbB0nD0_1;
	wire w_dff_B_kCkRmjlp8_1;
	wire w_dff_B_u2NDm4Ji8_1;
	wire w_dff_B_QscYYWEd6_1;
	wire w_dff_B_yIrNcaTs8_1;
	wire w_dff_B_2Clwai8F5_1;
	wire w_dff_B_TnMGmJki1_1;
	wire w_dff_B_uvmzdZ8J0_1;
	wire w_dff_B_NhtVaw2U4_1;
	wire w_dff_B_yX9Qr8n53_1;
	wire w_dff_B_xOVJDA0A4_1;
	wire w_dff_B_CF214jRL6_1;
	wire w_dff_B_xNzka8Gs5_1;
	wire w_dff_B_U0u26TLn6_1;
	wire w_dff_B_pUClwu2V7_1;
	wire w_dff_B_CazNRacx3_1;
	wire w_dff_B_bxQZ3oYx8_1;
	wire w_dff_B_nTwStTD28_1;
	wire w_dff_B_zsWtJ7c32_1;
	wire w_dff_B_Lf3YjB8x2_1;
	wire w_dff_B_o5iXYbXe4_1;
	wire w_dff_B_uMs40pPp2_1;
	wire w_dff_A_5PzhnG0g9_0;
	wire w_dff_B_G2sRD8PB5_2;
	wire w_dff_B_4pyoJNWl4_2;
	wire w_dff_B_qjv0Lg5Z6_2;
	wire w_dff_B_3MkCsW2U8_2;
	wire w_dff_B_kQ10nz9p1_2;
	wire w_dff_B_1TB3yJBA4_2;
	wire w_dff_B_0cVblnQ83_2;
	wire w_dff_B_mqZiUbpZ1_2;
	wire w_dff_B_zfdWl9Zc2_2;
	wire w_dff_B_a08hvitt5_2;
	wire w_dff_B_YKOnaPrb3_2;
	wire w_dff_B_vnqouHvk9_2;
	wire w_dff_B_FHxVOqjL8_2;
	wire w_dff_B_JAcY4Fv07_2;
	wire w_dff_B_PK82reXo3_2;
	wire w_dff_B_NM65Ng3H3_2;
	wire w_dff_B_BVVFdk8K6_2;
	wire w_dff_B_YG7X9TBI8_2;
	wire w_dff_B_GtGNpjkY6_0;
	wire w_dff_B_MksgHUwL4_0;
	wire w_dff_B_prF0gspV3_0;
	wire w_dff_B_hYk4TRTn1_0;
	wire w_dff_B_aBFwM9Tn0_0;
	wire w_dff_B_Le84nWLh8_0;
	wire w_dff_B_zRQ6A17J5_0;
	wire w_dff_B_3apr6BjE8_0;
	wire w_dff_B_tZ7XdPbV2_0;
	wire w_dff_B_wyiDseBh1_0;
	wire w_dff_B_94EGorVZ2_0;
	wire w_dff_B_7RpELD2L9_0;
	wire w_dff_B_g4GfoDlH0_0;
	wire w_dff_B_tUEC23Bw2_0;
	wire w_dff_B_LWWXeHGo1_0;
	wire w_dff_B_fdGn16v56_0;
	wire w_dff_B_vE0mNmXg8_0;
	wire w_dff_B_QVuiiY506_0;
	wire w_dff_B_SWav6wUL2_0;
	wire w_dff_B_2jcijqAw9_0;
	wire w_dff_B_icxVN9Xl1_0;
	wire w_dff_B_rEnROenV5_0;
	wire w_dff_B_g9ZzwNWj2_0;
	wire w_dff_B_U9Uof8Zi7_0;
	wire w_dff_B_aJjHLNgA8_0;
	wire w_dff_B_NbkvPVtR2_0;
	wire w_dff_A_95i5VaAd0_1;
	wire w_dff_A_2vsiFvqM0_1;
	wire w_dff_A_2x4lTKbJ3_1;
	wire w_dff_A_lxuxghtD1_1;
	wire w_dff_A_c5R14jvO5_1;
	wire w_dff_A_6E9jmO564_1;
	wire w_dff_A_6kuqJZYv6_1;
	wire w_dff_A_drh3cEUA6_1;
	wire w_dff_B_ekGaqtbt1_1;
	wire w_dff_B_em3F549f2_1;
	wire w_dff_A_OOfnODKZ7_1;
	wire w_dff_A_PbHA0OyO1_1;
	wire w_dff_A_ii7swT7v9_1;
	wire w_dff_A_ojVSGgJo3_1;
	wire w_dff_A_KuaHP4KI2_1;
	wire w_dff_A_EKFCEww64_1;
	wire w_dff_A_n05DZqeF9_1;
	wire w_dff_A_1mhXccgt4_1;
	wire w_dff_A_sb2m2DnT4_1;
	wire w_dff_A_gEWU635e2_1;
	wire w_dff_A_FMnkG7ba4_1;
	wire w_dff_A_yYzzaMCv0_1;
	wire w_dff_A_o5MYQtDW6_1;
	wire w_dff_A_eO6sFnFc8_1;
	wire w_dff_A_JcHFkQZf7_1;
	wire w_dff_A_FFasYZI84_1;
	wire w_dff_A_8QdHh2Jl3_1;
	wire w_dff_A_RA75SVgC6_1;
	wire w_dff_A_eLsNsyci3_1;
	wire w_dff_A_ZAfiIHrD6_1;
	wire w_dff_A_mU4icPyt6_1;
	wire w_dff_A_Hk5LcA3I3_1;
	wire w_dff_A_OLArNwdu6_1;
	wire w_dff_A_450TeNIi1_1;
	wire w_dff_A_448yc5vn0_1;
	wire w_dff_A_WzubKg2U0_1;
	wire w_dff_A_2DXACgZw7_1;
	wire w_dff_A_BCmgUvh55_1;
	wire w_dff_B_6BwQGnYJ8_2;
	wire w_dff_B_5rJKp6IJ3_2;
	wire w_dff_A_26WJXEW48_2;
	wire w_dff_A_8lV63m5T9_2;
	wire w_dff_A_Kk9NeGaH9_2;
	wire w_dff_A_Qq3bdX2w1_2;
	wire w_dff_A_xYp5hSQi3_2;
	wire w_dff_A_3GavLteP2_2;
	wire w_dff_A_soFWozYs9_2;
	wire w_dff_A_PKlY2QPT2_2;
	wire w_dff_A_Eeg1FAdI2_2;
	wire w_dff_A_ehGKBBX01_2;
	wire w_dff_A_WYxLSF3l4_2;
	wire w_dff_A_qGSlH1az1_2;
	wire w_dff_A_BwZ8dWmo5_2;
	wire w_dff_A_gc5Xm6gJ7_2;
	wire w_dff_A_GZw4V4NJ9_2;
	wire w_dff_A_11tYlTAR9_2;
	wire w_dff_A_ntvZ2byh4_2;
	wire w_dff_A_PBxKXlHt8_2;
	wire w_dff_A_VxsJxqaG4_2;
	wire w_dff_A_HYr82aQo3_2;
	wire w_dff_A_nMrlwQhx4_2;
	wire w_dff_A_S6hBsDT89_2;
	wire w_dff_A_Fb0cOCXF9_2;
	wire w_dff_B_D0gJOx8J1_1;
	wire w_dff_B_JOGLfg5g2_1;
	wire w_dff_B_QDr4lZed4_1;
	wire w_dff_B_V0Nq0Ly36_1;
	wire w_dff_B_EgzQaDCc9_1;
	wire w_dff_B_NLcblhT63_1;
	wire w_dff_B_B0usU2pS8_1;
	wire w_dff_B_eSJ1HwC54_1;
	wire w_dff_B_K0MX5dgt9_1;
	wire w_dff_A_Auvk7I1V0_2;
	wire w_dff_A_fUBhY7kh0_2;
	wire w_dff_A_Utp2DALW4_2;
	wire w_dff_A_LSik3jui9_2;
	wire w_dff_A_X1zzGqSG2_2;
	wire w_dff_A_GFpTUtin8_2;
	wire w_dff_A_AlyYxMXm2_2;
	wire w_dff_A_GbjKeSl74_2;
	wire w_dff_A_gyv9OaHD0_2;
	wire w_dff_A_1wuB2zG22_2;
	wire w_dff_A_Qtp3fshZ6_2;
	wire w_dff_A_sYSJHyLy6_2;
	wire w_dff_A_XNjKxdey5_2;
	wire w_dff_A_wpMgTIkY9_2;
	wire w_dff_A_20HUvQGN2_2;
	wire w_dff_A_OKMVvEvr9_2;
	wire w_dff_A_rgZNpjYs0_2;
	wire w_dff_A_7wVfDs5L1_2;
	wire w_dff_A_wSxouZwt2_2;
	wire w_dff_A_YoTaRUFu5_2;
	wire w_dff_A_Xph7QObS9_2;
	wire w_dff_A_Dvp3fPxA5_2;
	wire w_dff_A_hkYNGdsl8_2;
	wire w_dff_A_qBUx1Ono8_2;
	wire w_dff_A_DhCr42MS9_2;
	wire w_dff_B_2gdIxIEi6_1;
	wire w_dff_A_TIdTR1mS2_0;
	wire w_dff_A_w8WYQ7RD0_1;
	wire w_dff_A_y3yCDxrG6_1;
	wire w_dff_A_RerjHRQO9_1;
	wire w_dff_A_KXCRNkLg3_1;
	wire w_dff_A_jBhf4Lxe5_1;
	wire w_dff_A_OhkghTEl0_1;
	wire w_dff_A_x97otNYY5_1;
	wire w_dff_A_zUzEgu3P4_1;
	wire w_dff_A_N4XDKADg7_1;
	wire w_dff_A_sdnuuLMM9_1;
	wire w_dff_A_f3gOcPDY1_1;
	wire w_dff_A_NKn7JzbY6_1;
	wire w_dff_A_onvQ0Hb92_1;
	wire w_dff_A_eK6BNmJJ1_1;
	wire w_dff_A_OED5NbrK0_1;
	wire w_dff_A_Y7X0RcEi9_1;
	wire w_dff_A_CWUemXRA2_1;
	wire w_dff_A_4AWYKe2d6_1;
	wire w_dff_A_bfFZYIRT3_1;
	wire w_dff_A_PlTYs98K0_1;
	wire w_dff_A_LRCSOgBY0_1;
	wire w_dff_A_USyveyuP5_1;
	wire w_dff_A_rjpMRCjg1_1;
	wire w_dff_A_fvwy0dSg3_1;
	wire w_dff_A_HqRy27oo6_1;
	wire w_dff_A_ukSRDnTv1_1;
	wire w_dff_A_cDnUIF5z5_1;
	wire w_dff_A_WADLSwTz5_1;
	wire w_dff_A_RpciiL6M2_1;
	wire w_dff_A_j8rANZNm7_1;
	wire w_dff_A_jYbaV7PM9_1;
	wire w_dff_A_SX3eBsGe0_1;
	wire w_dff_B_6lWvEOl36_0;
	wire w_dff_A_N6RBtDlV2_0;
	wire w_dff_A_0ZPv1UgA1_0;
	wire w_dff_A_h0z2qC435_1;
	wire w_dff_A_zqEgeehC9_1;
	wire w_dff_A_sOUMJ5Uv7_0;
	wire w_dff_A_W7zyNWZK3_0;
	wire w_dff_A_76V8GQ9D3_0;
	wire w_dff_A_j9cYzXVv8_0;
	wire w_dff_A_Hs3YZ0n28_0;
	wire w_dff_B_CaE08qKQ8_2;
	wire w_dff_A_HCOW2wxX5_0;
	wire w_dff_A_sDvOWC695_0;
	wire w_dff_A_Mk3Y9kGR3_1;
	wire w_dff_A_8hA8yP7X7_1;
	wire w_dff_A_d1f47uPV5_0;
	wire w_dff_A_esoiYOnO9_2;
	wire w_dff_A_GkomEHwd6_0;
	wire w_dff_A_unS6yNBJ5_0;
	wire w_dff_A_K6p4i9Ny4_2;
	wire w_dff_A_NJOsFSPx2_2;
	wire w_dff_A_bWBHz9yJ3_2;
	wire w_dff_A_xElJ8NFB3_2;
	wire w_dff_A_ZQmCDssD9_2;
	wire w_dff_A_SR6dHKWw2_2;
	wire w_dff_A_GJFWv1ec1_2;
	wire w_dff_A_FYbWQtoV8_0;
	wire w_dff_A_MM8c0lGK3_0;
	wire w_dff_B_xc9uFfJ31_0;
	wire w_dff_A_w7Q4eY0z2_1;
	wire w_dff_A_SuyAG6dD7_1;
	wire w_dff_A_OAyUsTmf6_2;
	wire w_dff_A_Zkr9sd264_2;
	wire w_dff_B_wQ2PMfI50_1;
	wire w_dff_B_rfSBHnSX5_1;
	wire w_dff_B_aCJDbkf27_1;
	wire w_dff_B_15NAMZfR8_1;
	wire w_dff_B_ySkQdOIf1_1;
	wire w_dff_B_Lz3C0pVl2_1;
	wire w_dff_B_iKfYZPQF9_1;
	wire w_dff_B_ln7zhQeV7_1;
	wire w_dff_B_wm5BKaSa1_1;
	wire w_dff_B_1zNhJcEm4_1;
	wire w_dff_B_dJbhAIgp7_1;
	wire w_dff_B_sdnlnBax3_1;
	wire w_dff_B_wQ1lNVpq3_1;
	wire w_dff_B_lvLgAINt7_1;
	wire w_dff_B_fmePZ4cR4_1;
	wire w_dff_B_SmiIqvJS0_1;
	wire w_dff_B_60ORWjGP0_1;
	wire w_dff_B_RWneN9S12_1;
	wire w_dff_B_WWYGcvMe7_1;
	wire w_dff_B_hmkJm5fk9_0;
	wire w_dff_B_LLCjecBY0_0;
	wire w_dff_B_m4UXWIJG9_0;
	wire w_dff_B_60MmKkKi2_0;
	wire w_dff_B_HPyX5hiM0_0;
	wire w_dff_B_DiZlY0Yg3_0;
	wire w_dff_B_GEykmAI96_0;
	wire w_dff_B_Xy1yLjEo5_0;
	wire w_dff_B_yVh2irt11_0;
	wire w_dff_B_Hul66GOv5_0;
	wire w_dff_B_rbbKn9bM4_0;
	wire w_dff_B_TtJHkCmy5_0;
	wire w_dff_B_EnLLDslU7_0;
	wire w_dff_B_eaqtGupW1_0;
	wire w_dff_A_53r8eIzj3_0;
	wire w_dff_A_h6UuGasn2_0;
	wire w_dff_A_NEgK3E738_0;
	wire w_dff_A_X1ENr5nY4_0;
	wire w_dff_A_BDQPPL190_0;
	wire w_dff_A_ejiq0jjN4_0;
	wire w_dff_A_UW2SCsm97_0;
	wire w_dff_A_74tjy7kl5_0;
	wire w_dff_A_B6lVHn3M9_0;
	wire w_dff_A_aDpe2EhD5_0;
	wire w_dff_A_FmcT6jx85_0;
	wire w_dff_A_kO7549DR1_0;
	wire w_dff_A_tsQ1su0p6_0;
	wire w_dff_A_a3tr2dka2_0;
	wire w_dff_A_iQeXEwhg6_0;
	wire w_dff_B_HYJttRAU5_1;
	wire w_dff_B_kDrfp6vL7_1;
	wire w_dff_B_gokY1vEq5_1;
	wire w_dff_B_BKExFhTI0_1;
	wire w_dff_B_a29utAwe0_1;
	wire w_dff_B_rGygypLd3_1;
	wire w_dff_B_CdlzwAyf0_1;
	wire w_dff_B_J0VlKb5g2_1;
	wire w_dff_B_9bmPxkie9_1;
	wire w_dff_B_FraTEUNL8_1;
	wire w_dff_B_MJ4rqQGV0_1;
	wire w_dff_B_UsLOLSfz0_1;
	wire w_dff_B_0FtXJN2A7_1;
	wire w_dff_B_oQpbIVWX8_1;
	wire w_dff_B_K601PMIT9_1;
	wire w_dff_B_XxnRDXtu6_1;
	wire w_dff_B_LOLKaIid3_1;
	wire w_dff_B_Uz1Zm8eK4_1;
	wire w_dff_B_CtHFdiwh9_1;
	wire w_dff_B_mmI1cXgL2_1;
	wire w_dff_B_BLjKThjL5_1;
	wire w_dff_B_gVy1CQY12_1;
	wire w_dff_B_ORUcWxsl2_1;
	wire w_dff_B_aFFUNSsZ1_1;
	wire w_dff_B_Ii41U4s57_1;
	wire w_dff_B_iDlq5Qbu8_1;
	wire w_dff_B_jnmVzGmV2_1;
	wire w_dff_B_wug3JZzv1_1;
	wire w_dff_B_pVU240ri1_1;
	wire w_dff_B_PJ3UrIzK9_1;
	wire w_dff_B_WC41jezt4_1;
	wire w_dff_B_QMvArpxz2_1;
	wire w_dff_B_DYUbNjOo5_1;
	wire w_dff_B_W33OGnFZ9_1;
	wire w_dff_A_amAYhCsa7_1;
	wire w_dff_A_GpTyvR8n3_1;
	wire w_dff_A_tIBXdVDf5_1;
	wire w_dff_A_UUAEIRxE0_1;
	wire w_dff_A_EqCf6LOY1_1;
	wire w_dff_A_tBMhYuYz7_1;
	wire w_dff_A_EbzSqyfX0_1;
	wire w_dff_A_o4hKN4Nk7_1;
	wire w_dff_A_NcVEOXhi5_1;
	wire w_dff_A_SjxkgvLG3_1;
	wire w_dff_A_LaQBvpyP2_1;
	wire w_dff_A_ouPtDqXW0_1;
	wire w_dff_A_UgnEGHoV7_1;
	wire w_dff_A_RfMCjFwd9_1;
	wire w_dff_A_OkbB5HG98_1;
	wire w_dff_A_jBLPjwIz9_1;
	wire w_dff_A_jhMpSaWM5_1;
	wire w_dff_A_SsTPKTdV9_1;
	wire w_dff_A_cC4jDxwZ0_1;
	wire w_dff_A_wrJvwDwI0_0;
	wire w_dff_A_MOh5qngo9_0;
	wire w_dff_A_W5BhSzPy5_0;
	wire w_dff_A_IADBaKt47_0;
	wire w_dff_A_Klcoe3uJ0_0;
	wire w_dff_A_PL2uC0MR5_0;
	wire w_dff_A_edNij6l28_0;
	wire w_dff_A_Xr05sfnV4_0;
	wire w_dff_A_bABSf4G24_0;
	wire w_dff_A_X09YGMTN7_0;
	wire w_dff_A_k30zt85Z7_0;
	wire w_dff_A_5t6lLZ050_0;
	wire w_dff_A_Bcu7KTF06_0;
	wire w_dff_A_DbDF4rQJ7_0;
	wire w_dff_A_xSbZG5Ba2_0;
	wire w_dff_A_hdv4s7Pz1_0;
	wire w_dff_A_XiWMazXS0_0;
	wire w_dff_A_FNKjGO625_0;
	wire w_dff_A_T6Ux1lWC6_0;
	wire w_dff_A_aJryGNPj1_0;
	wire w_dff_A_gNaQHZmM1_1;
	wire w_dff_A_xuIBbaxg9_1;
	wire w_dff_A_kxZRG5zq2_1;
	wire w_dff_A_QdAeCn2i2_1;
	wire w_dff_A_BcsaBom17_1;
	wire w_dff_A_gODWlgmR5_1;
	wire w_dff_A_3JcRLIeR3_1;
	wire w_dff_A_faKNPZ6T9_1;
	wire w_dff_A_ANRzoikc5_1;
	wire w_dff_A_Kh3lZXq61_1;
	wire w_dff_A_3c3ITUf51_1;
	wire w_dff_A_GaVM0qnd6_1;
	wire w_dff_A_lNJnqCOM6_1;
	wire w_dff_A_JRCDhjtx9_1;
	wire w_dff_A_cDo7qvmm0_1;
	wire w_dff_A_ZAEKEhuG8_1;
	wire w_dff_A_WMbwGSev8_1;
	wire w_dff_A_PrlsKesa0_1;
	wire w_dff_A_h6i8hGZv5_1;
	wire w_dff_A_RGcGofez3_1;
	wire w_dff_A_BopCeC6t1_1;
	wire w_dff_A_xavBH0ie1_1;
	wire w_dff_A_aB5MWU2t6_1;
	wire w_dff_A_NoNtTVNC3_1;
	wire w_dff_A_tcdEHWon4_1;
	wire w_dff_A_lSrIxcek8_1;
	wire w_dff_A_Ih3zeL8h5_1;
	wire w_dff_A_oJjRbQZT4_1;
	wire w_dff_A_MnWO2fIl3_1;
	wire w_dff_A_TO7YJ9K24_1;
	wire w_dff_A_CxsKsmNL5_1;
	wire w_dff_A_p53AzdjF4_1;
	wire w_dff_A_JCFtJ09t4_1;
	wire w_dff_A_tIeBY7ZP5_1;
	wire w_dff_A_Y1AugM6I4_1;
	wire w_dff_A_Rus3fZtn4_1;
	wire w_dff_A_38b6xME91_1;
	wire w_dff_A_3boJ5GZc9_1;
	wire w_dff_A_bOSuo1ok3_1;
	wire w_dff_A_DKf7sUZJ4_1;
	wire w_dff_A_w2kgbuby9_1;
	wire w_dff_A_cy97yl1b8_1;
	wire w_dff_A_TKdoqjWU0_1;
	wire w_dff_A_CuFBcBUB5_1;
	wire w_dff_A_m61EdLbR0_1;
	wire w_dff_A_uxma2TSc2_1;
	wire w_dff_A_YvnfCmG75_1;
	wire w_dff_A_n1su2Csh1_1;
	wire w_dff_A_p0RGQNFY8_1;
	wire w_dff_A_xt7GjEEB2_1;
	wire w_dff_A_tAXEGNpo0_1;
	wire w_dff_A_9Jayynfx4_1;
	wire w_dff_A_RhW9o69O3_1;
	wire w_dff_A_1RskFi178_1;
	wire w_dff_A_N7mi49Vo4_1;
	wire w_dff_A_VbIRRRyl1_1;
	wire w_dff_A_msWSaFgt3_1;
	wire w_dff_A_Aak0B7AL6_0;
	wire w_dff_A_P05SiyRm0_0;
	wire w_dff_A_R0djuMDo8_0;
	wire w_dff_A_ZK73vVpY6_0;
	wire w_dff_A_Kw7ugb9f3_0;
	wire w_dff_A_HeY7sfu61_0;
	wire w_dff_A_m2ZkOJmp7_0;
	wire w_dff_A_cCxWXWnh5_0;
	wire w_dff_A_lVYM9zJJ2_0;
	wire w_dff_A_kq8E1F326_0;
	wire w_dff_A_9te5rlwh6_0;
	wire w_dff_A_wOFbS5LS0_0;
	wire w_dff_A_EBLLEKGN7_0;
	wire w_dff_A_T1FhP12T4_0;
	wire w_dff_A_rBfVoVXJ8_0;
	wire w_dff_A_QcH6RXIT7_0;
	wire w_dff_A_h3i2shtr9_0;
	wire w_dff_A_BvmYfvAB1_0;
	wire w_dff_A_VJ2PfoYk9_0;
	wire w_dff_B_WyeZXHbr1_1;
	wire w_dff_B_4X3kPJrL4_1;
	wire w_dff_B_g08RlGq63_1;
	wire w_dff_A_jMcenfR22_0;
	wire w_dff_A_fbyIUOcx5_0;
	wire w_dff_A_4cOLjCDA2_0;
	wire w_dff_A_CNbKM23z5_0;
	wire w_dff_A_vrYdFfq63_0;
	wire w_dff_A_AhgtTm8d6_0;
	wire w_dff_A_Vm7Bi5zH8_0;
	wire w_dff_A_HxeLPVrN7_0;
	wire w_dff_A_v4MGICBa5_0;
	wire w_dff_A_1thZgHSK8_0;
	wire w_dff_A_sX3ENFkg6_0;
	wire w_dff_A_s6oeVN8V5_0;
	wire w_dff_A_6jXzVsJW9_0;
	wire w_dff_A_bktw3wX13_0;
	wire w_dff_A_gb6Wb1IB8_0;
	wire w_dff_A_zp2ffKLE6_0;
	wire w_dff_A_bXSlSjE39_0;
	wire w_dff_A_hLKCT2WW2_0;
	wire w_dff_A_i8ufmyLE3_0;
	wire w_dff_B_JtsGdVzx3_1;
	wire w_dff_B_2dzCEDNR0_1;
	wire w_dff_A_deUKMUkG8_0;
	wire w_dff_A_morsh9Fq2_0;
	wire w_dff_A_LLfcPI5v9_0;
	wire w_dff_A_wG0ZifpE8_2;
	wire w_dff_A_VKErXlhW5_2;
	wire w_dff_A_Td4dErbD5_1;
	wire w_dff_A_RJv3wE9p0_1;
	wire w_dff_A_sXwtEneV7_1;
	wire w_dff_A_LqLvx6vs9_1;
	wire w_dff_A_Y9Y3BmyK7_1;
	wire w_dff_A_euV10qq49_1;
	wire w_dff_A_zxgVdpJs7_1;
	wire w_dff_A_fA7HAnm02_1;
	wire w_dff_A_VfDpkJqr1_1;
	wire w_dff_A_nlt2YmsH7_1;
	wire w_dff_A_DPtj4cdg5_1;
	wire w_dff_A_af5DXFEl3_1;
	wire w_dff_A_6giP8EKq3_1;
	wire w_dff_A_Dw9AWMnf6_1;
	wire w_dff_A_F0DtYoY39_1;
	wire w_dff_A_ctsS75dJ9_1;
	wire w_dff_A_dtPwwUCt7_1;
	wire w_dff_A_H8CTkzRh7_1;
	wire w_dff_A_HOC6O1zJ7_1;
	wire w_dff_A_CVe3MJHb0_1;
	wire w_dff_A_uttDgsHk0_1;
	wire w_dff_A_ywD6YQRO6_1;
	wire w_dff_A_l3fDYImI1_1;
	wire w_dff_A_AdtOCzBY1_1;
	wire w_dff_A_ixqYGm1o7_0;
	wire w_dff_A_Wv6rvCIi5_0;
	wire w_dff_A_YgJCA40H7_0;
	wire w_dff_A_FoBgatEC9_0;
	wire w_dff_A_SLK28GeL0_0;
	wire w_dff_A_fw7sQ5W87_0;
	wire w_dff_A_bjHvmDvY6_0;
	wire w_dff_A_TqdS7yiw2_0;
	wire w_dff_A_jeJvfZqg1_0;
	wire w_dff_A_EJyWmnr29_0;
	wire w_dff_A_ljWnEnYu4_0;
	wire w_dff_A_LxUaOaY84_0;
	wire w_dff_A_OJIukkaT8_0;
	wire w_dff_A_cq1EfrJU1_0;
	wire w_dff_A_Jsq2I9WM1_0;
	wire w_dff_A_dqOX5aeL9_0;
	wire w_dff_A_jgP0GqKZ1_0;
	wire w_dff_A_vVf75h6x2_0;
	wire w_dff_A_nB36qrht8_0;
	wire w_dff_A_wDM6Fowa2_0;
	wire w_dff_A_zEyFOwDZ0_0;
	wire w_dff_A_PjQxVjRq2_0;
	wire w_dff_A_7dEHGSlS3_2;
	wire w_dff_A_Unfq8XEe0_2;
	wire w_dff_A_XBArIg9C2_2;
	wire w_dff_A_93PiUjLl4_2;
	wire w_dff_A_5f2KQPVj1_2;
	wire w_dff_A_dqu1Ec3R5_2;
	wire w_dff_A_dxGJRV5L1_2;
	wire w_dff_A_kMabNZBW6_2;
	wire w_dff_A_du08SVZh0_2;
	wire w_dff_A_9PwJ1itP8_2;
	wire w_dff_A_s2YSep9r3_2;
	wire w_dff_A_4mgP7Jwu0_2;
	wire w_dff_A_V2A7bli74_2;
	wire w_dff_A_eZTe3fYw8_2;
	wire w_dff_A_IkjMENBR8_2;
	wire w_dff_A_pe96QAlF8_2;
	wire w_dff_A_c4aHzUs29_2;
	wire w_dff_A_z62fQYdD3_2;
	wire w_dff_A_4SEeGFhv8_2;
	wire w_dff_A_KOHVLl2s2_2;
	wire w_dff_A_UYgUFvLc4_2;
	wire w_dff_A_W2yMJyFv7_2;
	wire w_dff_A_qzEOAB5K5_2;
	wire w_dff_B_YBVMhFrw4_0;
	wire w_dff_B_sPQTSDO91_0;
	wire w_dff_A_rbide4Po5_1;
	wire w_dff_A_nz0WVmC46_1;
	wire w_dff_A_pR8aIAKi6_2;
	wire w_dff_A_1SPzV9KS9_2;
	wire w_dff_A_sGQoS01B7_1;
	wire w_dff_A_qrDWNDAB0_1;
	wire w_dff_A_MnOJFYCr0_1;
	wire w_dff_A_4jd6T85v2_1;
	wire w_dff_A_6rNoCX3n4_1;
	wire w_dff_A_NotIBoFg4_1;
	wire w_dff_A_CblEHEA98_1;
	wire w_dff_A_o9EmDkHT5_1;
	wire w_dff_A_c25rgt6U1_1;
	wire w_dff_A_iP8JrcrQ8_1;
	wire w_dff_A_5uCsJvHT3_1;
	wire w_dff_A_Ar5yrfF34_1;
	wire w_dff_A_8K2was2a9_1;
	wire w_dff_A_KE3zLGnF9_1;
	wire w_dff_A_60TIwxxS2_1;
	wire w_dff_A_8QjpGOze1_1;
	wire w_dff_A_3ICgD0yx3_1;
	wire w_dff_A_zQHypauh2_1;
	wire w_dff_A_Y2HCjpeZ3_1;
	wire w_dff_A_QrAtwv8C7_1;
	wire w_dff_A_Pf1AyaWd1_1;
	wire w_dff_A_WN2omO4Y4_1;
	wire w_dff_A_BKSl8FZe3_1;
	wire w_dff_A_NgHy1mTr1_1;
	wire w_dff_A_pqVDuJwH0_1;
	wire w_dff_A_ioEIHelg3_1;
	wire w_dff_A_CheGRkuj5_1;
	wire w_dff_A_p3LiCpr75_1;
	wire w_dff_A_iNqFcuDB5_1;
	wire w_dff_B_ahLzISW37_0;
	wire w_dff_B_F3PASO123_0;
	wire w_dff_A_sqRzoyHI0_1;
	wire w_dff_A_AEUcQ3Nn0_1;
	wire w_dff_A_tCymbE621_2;
	wire w_dff_A_CoRA3fFb5_2;
	wire w_dff_A_tavuTiH99_1;
	wire w_dff_A_WktiMIxJ5_1;
	wire w_dff_A_DQVx4nYE2_1;
	wire w_dff_A_ejDtG6IA4_1;
	wire w_dff_A_PZWFXNLs9_1;
	wire w_dff_A_R86NxYsJ6_1;
	wire w_dff_A_C5vvK6m33_1;
	wire w_dff_A_kOnaPuB27_1;
	wire w_dff_A_3sMKEa3p7_1;
	wire w_dff_A_JhgKSz0k8_1;
	wire w_dff_A_nvpwnhzr6_1;
	wire w_dff_A_XTQAwFBM3_1;
	wire w_dff_A_043I4qEv6_1;
	wire w_dff_A_1tZbmfKg6_1;
	wire w_dff_A_YjaYXnGM2_1;
	wire w_dff_A_52dVQub69_1;
	wire w_dff_A_JNAGShZX7_1;
	wire w_dff_A_hLm5jJZp3_1;
	wire w_dff_A_lNNwIN8B6_1;
	wire w_dff_A_OewrYHc16_1;
	wire w_dff_A_v2heRr9F6_1;
	wire w_dff_A_dWEs66E19_1;
	wire w_dff_A_BhADi4hU3_1;
	wire w_dff_A_all0LASw7_1;
	wire w_dff_A_ZOi4iXss8_1;
	wire w_dff_A_D2x2x57p3_1;
	wire w_dff_A_VuCtGG891_1;
	wire w_dff_A_nDvXNVFL7_1;
	wire w_dff_A_T7jq9jDO9_1;
	wire w_dff_A_bhpvO7y81_2;
	wire w_dff_A_2iW2PPZY8_1;
	wire w_dff_B_KFM86BYY5_0;
	wire w_dff_B_L0FO5yLy8_0;
	wire w_dff_B_7VdUCKjH3_2;
	wire w_dff_B_faLwkV1V1_2;
	wire w_dff_A_caASnzbL5_0;
	wire w_dff_A_VoAJ2kes2_0;
	wire w_dff_A_v13rWSEn4_0;
	wire w_dff_A_l1y0aVPn7_0;
	wire w_dff_A_AEtra7w43_1;
	wire w_dff_B_l2wkP1F76_2;
	wire w_dff_B_4kkUNG699_2;
	wire w_dff_B_Q6mApC7R4_2;
	wire w_dff_B_8NkWGC5a1_2;
	wire w_dff_A_pOGrQRJ74_1;
	wire w_dff_A_4cFrbtet4_1;
	wire w_dff_A_ttM2uUXo0_1;
	wire w_dff_A_G6gEQHXt7_1;
	wire w_dff_A_TvL30THj2_1;
	wire w_dff_A_5cxykv8L1_1;
	wire w_dff_A_zCXWJnRx8_1;
	wire w_dff_A_13AGVodk3_1;
	wire w_dff_A_X2WrYvLe1_1;
	wire w_dff_A_oMdgqgGd7_1;
	wire w_dff_A_2OckOhek1_1;
	wire w_dff_A_o4723JXm7_1;
	wire w_dff_A_GpWcJurk9_1;
	wire w_dff_A_qY5T57XT4_1;
	wire w_dff_A_k2u2chqi7_1;
	wire w_dff_A_GTWvrOJQ6_1;
	wire w_dff_A_TF61Uxpp9_1;
	wire w_dff_A_41JQzHdh9_1;
	wire w_dff_A_pDyqnRQE7_1;
	wire w_dff_A_lhbev20A3_1;
	wire w_dff_A_4O90wrX25_1;
	wire w_dff_A_yQmnoKOA2_1;
	wire w_dff_A_r1MOO3YE6_1;
	wire w_dff_A_wJUIGS9O9_1;
	wire w_dff_A_LN73Blkg7_1;
	wire w_dff_A_k81yAa526_1;
	wire w_dff_A_UaCQODc75_0;
	wire w_dff_A_UjtKMMZn4_0;
	wire w_dff_A_ptbWX0HT0_0;
	wire w_dff_A_K3ootG9A8_0;
	wire w_dff_A_UpRHNI212_0;
	wire w_dff_A_Go9qbMMu2_0;
	wire w_dff_A_yC46ZHJd7_0;
	wire w_dff_A_8k6Kz5o43_0;
	wire w_dff_A_2qiBYBpj5_0;
	wire w_dff_A_WPKsUuVp2_0;
	wire w_dff_A_s4JpMiZd2_0;
	wire w_dff_A_WQ8eqC0R4_0;
	wire w_dff_A_jQedEa9h7_0;
	wire w_dff_A_mimc7q7d7_0;
	wire w_dff_A_meMNJLVk2_0;
	wire w_dff_A_5flPCkGW2_0;
	wire w_dff_A_whrHmqgw8_0;
	wire w_dff_A_5S1UkWTf8_0;
	wire w_dff_A_SHWbbS468_0;
	wire w_dff_A_rEpJmsOW1_0;
	wire w_dff_A_Oaej3STT6_0;
	wire w_dff_A_dNXNp3CK8_0;
	wire w_dff_A_J2DPbQwi1_0;
	wire w_dff_A_pcoKWbB46_0;
	wire w_dff_A_gldFSnIi1_0;
	wire w_dff_A_j2LrPGVh2_0;
	wire w_dff_A_bYv9v9ah0_0;
	wire w_dff_A_mm9xl4ny1_0;
	wire w_dff_A_G1k9tSbX4_1;
	wire w_dff_A_3dcrqoOw5_1;
	wire w_dff_A_OOnyHpnr0_1;
	wire w_dff_A_HOEtFrdf6_2;
	wire w_dff_A_mggUfphE7_2;
	wire w_dff_A_GiEsqJZu5_2;
	wire w_dff_A_23iTfWE05_2;
	wire w_dff_A_Rf91Ri1L3_1;
	wire w_dff_A_hpJFL3sK0_1;
	wire w_dff_A_Z26zVEXv0_1;
	wire w_dff_A_vjieTZMz6_1;
	wire w_dff_A_cdWFS5cL6_1;
	wire w_dff_A_ky4Amsyu1_1;
	wire w_dff_A_hgSBaEk42_1;
	wire w_dff_A_OlHMVJ4s3_1;
	wire w_dff_A_t7KsHmnV8_1;
	wire w_dff_A_pN6C2wDF7_1;
	wire w_dff_A_SDN5vM8n2_1;
	wire w_dff_A_nfEqkOvf0_1;
	wire w_dff_A_uyfU2R556_1;
	wire w_dff_A_P376HyIw7_1;
	wire w_dff_A_NFZRabpp8_1;
	wire w_dff_A_X7Ynu4Cz3_1;
	wire w_dff_A_QipKPhqW4_1;
	wire w_dff_A_NcPLJRFM8_1;
	wire w_dff_A_vJhYnvck0_1;
	wire w_dff_A_qc4czDye1_1;
	wire w_dff_A_KeAGqp0V3_1;
	wire w_dff_A_L9VoewlE4_2;
	wire w_dff_A_qzCVUCyk7_2;
	wire w_dff_A_bPgGgxjM5_2;
	wire w_dff_A_gKC5si9E3_2;
	wire w_dff_A_9UTW68s00_2;
	wire w_dff_B_awopLnNH5_1;
	wire w_dff_A_k54MonoF7_0;
	wire w_dff_A_XFZsADoa1_0;
	wire w_dff_A_6Fzfy2Kw6_0;
	wire w_dff_A_WOMwj1407_0;
	wire w_dff_A_lTbCl6VD0_0;
	wire w_dff_A_Jaufee2s4_0;
	wire w_dff_A_3K3HuQsC1_0;
	wire w_dff_A_I8bYwQpi8_0;
	wire w_dff_A_tr4JXemg5_0;
	wire w_dff_A_uVdBUZgR5_0;
	wire w_dff_A_lJRI20IG7_0;
	wire w_dff_A_OggVfmVL6_0;
	wire w_dff_A_fbyLv0JS6_0;
	wire w_dff_A_JLadxANj4_0;
	wire w_dff_A_TaoVFQzy5_0;
	wire w_dff_A_CUw2PL7y8_0;
	wire w_dff_A_3Ykac4vI4_0;
	wire w_dff_A_2HLiQELv2_0;
	wire w_dff_A_gEPW8tZJ0_0;
	wire w_dff_A_tPxeaxz58_0;
	wire w_dff_A_XZ6FJpzZ7_0;
	wire w_dff_A_mXitxHfX8_0;
	wire w_dff_A_MM3YtLNQ1_0;
	wire w_dff_A_D83NkRkf2_0;
	wire w_dff_A_Prlrm1Jf5_0;
	wire w_dff_A_zpjBqJBo4_0;
	wire w_dff_A_PAbldBJs3_0;
	wire w_dff_A_mzPJmmpA5_0;
	wire w_dff_A_D6r6m7ZR6_1;
	wire w_dff_A_Cd2kLbxp1_1;
	wire w_dff_A_i6aS6Uzj7_1;
	wire w_dff_A_HZaM7yQs6_1;
	wire w_dff_A_p4hK0S748_1;
	wire w_dff_A_cs9eMcnY5_1;
	wire w_dff_A_OVY1ZdqL7_1;
	wire w_dff_A_QI2cO9NY5_1;
	wire w_dff_A_q5JZpPPZ4_1;
	wire w_dff_A_9ojgAUoF7_1;
	wire w_dff_A_uNPmcJ450_1;
	wire w_dff_A_Gu8katj50_1;
	wire w_dff_A_BFuNihQf4_1;
	wire w_dff_A_0jMCvRlY8_1;
	wire w_dff_A_y8KDwPwL0_1;
	wire w_dff_A_gD5kEaY65_1;
	wire w_dff_A_gLfuqoBq6_1;
	wire w_dff_A_BKMi7xRg3_1;
	wire w_dff_A_9CRIjJAW2_1;
	wire w_dff_A_l1Pl7gFq8_1;
	wire w_dff_A_R2MjCZWp0_1;
	wire w_dff_A_rlbrlT4k6_1;
	wire w_dff_A_ATBdNKld5_1;
	wire w_dff_A_boWxus9s7_1;
	wire w_dff_A_1m3cni3m7_1;
	wire w_dff_A_g6KYlXOQ2_1;
	wire w_dff_A_N4yhrShC2_1;
	wire w_dff_A_g1jzQxd28_1;
	wire w_dff_A_rYATWfRs2_1;
	wire w_dff_A_6p8k5DXg7_1;
	wire w_dff_A_VTlxaBkL6_1;
	wire w_dff_A_fIiVjdhg4_1;
	wire w_dff_A_oMDMfYxR4_1;
	wire w_dff_A_wc1m5kDg1_2;
	wire w_dff_A_NoJhKZFu6_2;
	wire w_dff_A_lJjdzwwr6_2;
	wire w_dff_A_nXayk9as8_2;
	wire w_dff_A_JsuecAtg8_2;
	wire w_dff_A_OJNo70x40_2;
	wire w_dff_A_qlnCXpzK1_2;
	wire w_dff_B_OMw2dKd80_0;
	wire w_dff_B_ysREwqJz0_0;
	wire w_dff_A_MTwDKs0H0_1;
	wire w_dff_A_GH49b0Su4_1;
	wire w_dff_A_wc2lkZX18_2;
	wire w_dff_A_ma0gtraA9_2;
	wire w_dff_A_R1Gxr56t4_1;
	wire w_dff_A_MfAaBqbI0_1;
	wire w_dff_A_G8sCmpI01_1;
	wire w_dff_A_Goj5lNI45_1;
	wire w_dff_A_awJpdhdt3_1;
	wire w_dff_B_EvTmIQ8u7_0;
	wire w_dff_B_MgTpLvgR6_3;
	wire w_dff_B_bNAyFE7f2_3;
	wire w_dff_A_3S1neNv82_2;
	wire w_dff_A_ykxDAA0P3_2;
	wire w_dff_A_tFbW4tOx3_2;
	wire w_dff_A_tvye38Pp7_2;
	wire w_dff_A_enhqDaiv4_2;
	wire w_dff_A_eItKloPp7_2;
	wire w_dff_A_0d6vNpb52_2;
	wire w_dff_A_yf62CRGq7_2;
	wire w_dff_A_LsuuyCNT7_2;
	wire w_dff_A_KA1S5kW75_2;
	wire w_dff_A_mMLIqVbr8_2;
	wire w_dff_A_qRfaVIaL4_2;
	wire w_dff_A_KYEyjIBc4_2;
	wire w_dff_A_jtDziYMX8_2;
	wire w_dff_A_JwZ5fufX0_2;
	wire w_dff_A_JO1coacm2_2;
	wire w_dff_A_Y0CwjJpz5_2;
	wire w_dff_A_nM01yALH0_2;
	wire w_dff_A_h2uaSdnx1_2;
	wire w_dff_A_DKY0ehu74_2;
	wire w_dff_A_5knmi0wC6_2;
	wire w_dff_A_DNUoJNJS9_2;
	wire w_dff_B_OMd4cECq2_1;
	wire w_dff_B_jcpkSiok6_1;
	wire w_dff_A_Do1sJfAz5_0;
	wire w_dff_A_NouzY9c38_0;
	wire w_dff_A_2CwuWeYS2_0;
	wire w_dff_A_rczZvGLY6_0;
	wire w_dff_A_3czVK9Hi5_0;
	wire w_dff_A_UPXzAwwS1_0;
	wire w_dff_A_Z7s8AnT55_0;
	wire w_dff_A_OCEYguF52_0;
	wire w_dff_A_cyVtxLIv9_0;
	wire w_dff_A_D8iRD0d30_0;
	wire w_dff_A_c88lOILW2_0;
	wire w_dff_A_rC09rrzG1_0;
	wire w_dff_A_T9WLxHLB0_0;
	wire w_dff_A_4rOCjNwl0_0;
	wire w_dff_A_oPhxW1jV8_0;
	wire w_dff_A_bPiOyOgD4_0;
	wire w_dff_A_Wv6O4urJ2_0;
	wire w_dff_A_S34mABln7_0;
	wire w_dff_A_4gEplQKp0_0;
	wire w_dff_A_B17cHXGn9_0;
	wire w_dff_A_zcWYUNbH5_0;
	wire w_dff_A_DJvvuMLZ3_0;
	wire w_dff_B_92yrD0BR6_1;
	wire w_dff_B_p7xMscoi9_1;
	wire w_dff_B_Ou96JSKD7_1;
	wire w_dff_A_lSOvDucG9_1;
	wire w_dff_A_0og9mOzJ2_1;
	wire w_dff_A_g8jwiIRc6_1;
	wire w_dff_A_562oG0IR3_1;
	wire w_dff_A_ooJOZcO43_1;
	wire w_dff_A_bQ5XIrnC0_1;
	wire w_dff_A_y6vuZmFO8_1;
	wire w_dff_A_77w7c0Vu9_1;
	wire w_dff_A_jT8ITcZl9_1;
	wire w_dff_A_u9H8DKzF4_1;
	wire w_dff_A_XUMC7h4P2_1;
	wire w_dff_A_MxfbuE8l9_1;
	wire w_dff_A_R0ntPxkG1_1;
	wire w_dff_A_D3ZAsYJc5_1;
	wire w_dff_A_1HMHWy0a3_1;
	wire w_dff_A_ql5cb95U8_1;
	wire w_dff_A_llMvCMUc7_1;
	wire w_dff_A_7myUnSTh2_1;
	wire w_dff_A_zp1yClKZ0_1;
	wire w_dff_A_3JW7lJiX4_1;
	wire w_dff_A_yZhDyhzO9_1;
	wire w_dff_A_moLcn9wU0_1;
	wire w_dff_A_56ri7JEp4_1;
	wire w_dff_A_GpfJrIyz1_1;
	wire w_dff_A_RFn9ktMs9_1;
	wire w_dff_A_VUVo3DE22_1;
	wire w_dff_A_5PZGs2378_1;
	wire w_dff_A_WsaBE3856_1;
	wire w_dff_A_TkcaGzHM1_1;
	wire w_dff_A_j2HZZJ2b8_1;
	wire w_dff_A_g3jquSgD0_1;
	wire w_dff_A_OZRE09i87_1;
	wire w_dff_A_etf9XN9x5_1;
	wire w_dff_A_0t2k46q24_1;
	wire w_dff_A_AJeRGgbJ2_1;
	wire w_dff_A_LYO3CrNn0_1;
	wire w_dff_A_SruZ1Knl4_1;
	wire w_dff_A_39mH9nLB8_1;
	wire w_dff_A_dh5nasNr4_1;
	wire w_dff_A_7mirB95L5_1;
	wire w_dff_A_OwyZFgff2_1;
	wire w_dff_A_2XPP5Prc7_1;
	wire w_dff_A_twyROc2w9_1;
	wire w_dff_A_L9IcrBII0_1;
	wire w_dff_A_Awvm9W7S9_1;
	wire w_dff_A_HhO3Cjdg8_1;
	wire w_dff_A_3z9xDdNO9_1;
	wire w_dff_A_yFnz547Q7_1;
	wire w_dff_A_6Fi2hSCE6_1;
	wire w_dff_A_S05y18lQ3_1;
	wire w_dff_A_OaUA8Du73_1;
	wire w_dff_A_uO1vhw4H7_1;
	wire w_dff_A_a66fwNCD5_1;
	wire w_dff_A_CO40dOUl0_2;
	wire w_dff_A_k6HhHNvI3_0;
	wire w_dff_A_CH0mOYP28_0;
	wire w_dff_A_IbM43Zvt2_0;
	wire w_dff_A_fLryOFyT8_0;
	wire w_dff_A_RIoNaBDg0_0;
	wire w_dff_A_vvyyG51H5_0;
	wire w_dff_A_Njb6Iykp2_0;
	wire w_dff_A_puOeH4213_0;
	wire w_dff_A_ZdalX3Tx6_0;
	wire w_dff_A_2YY4HiPW9_0;
	wire w_dff_A_o2mStPB95_0;
	wire w_dff_A_Zj86wMtU0_0;
	wire w_dff_A_F6N1Egpz5_0;
	wire w_dff_A_4stGaW3o8_0;
	wire w_dff_A_JX6KbI918_0;
	wire w_dff_A_PMK8qwEG7_0;
	wire w_dff_A_THvPmz6x0_0;
	wire w_dff_A_vsMZr1rU0_0;
	wire w_dff_A_K85VhOl68_0;
	wire w_dff_A_dEaryAQz7_0;
	wire w_dff_A_pgfyR0812_0;
	wire w_dff_A_FM1OgzgO3_0;
	wire w_dff_A_jWP61y9L6_0;
	wire w_dff_A_rMjcHjkf5_0;
	wire w_dff_A_ZCXL6AFb6_0;
	wire w_dff_A_NuFAHOKH5_1;
	wire w_dff_A_ugyEEQqb4_1;
	wire w_dff_A_B3uSnQhe1_1;
	wire w_dff_A_82knghJg4_1;
	wire w_dff_A_HVGFICnp9_1;
	wire w_dff_A_dueqnUqy6_1;
	wire w_dff_A_WAfWcaXV9_1;
	wire w_dff_A_Iv52h5mp0_1;
	wire w_dff_A_w8Fw9Eu57_1;
	wire w_dff_A_Uq9F3kxL2_1;
	wire w_dff_A_OfCpVxKO8_1;
	wire w_dff_A_zMsGmvg76_1;
	wire w_dff_A_Iq2PYwmo5_1;
	wire w_dff_A_lfKF9niy6_1;
	wire w_dff_A_pmBDn31b6_1;
	wire w_dff_A_W8PxzLLF1_1;
	wire w_dff_A_xjJsVOJO5_1;
	wire w_dff_A_fNhn1uZ19_1;
	wire w_dff_A_ugVYufGk2_1;
	wire w_dff_A_1xdISX657_1;
	wire w_dff_A_W9ZblWwJ6_1;
	wire w_dff_A_o4UjdsTI3_1;
	wire w_dff_A_6iqiNvZX1_1;
	wire w_dff_A_Y3GMXjN15_1;
	wire w_dff_A_sZMFraKx5_1;
	wire w_dff_A_tq65jwS84_1;
	wire w_dff_A_7jupj86t9_0;
	wire w_dff_A_9dsEoGvg6_0;
	wire w_dff_B_izHlvbbm7_0;
	wire w_dff_B_tyt6915Y6_2;
	wire w_dff_B_pwi9h59w5_2;
	wire w_dff_A_zLwudB9B5_2;
	wire w_dff_A_h8kQPKRa5_2;
	wire w_dff_A_FZhp2flj2_2;
	wire w_dff_A_qd8jTaPx2_2;
	wire w_dff_A_AlzcVAKM9_0;
	wire w_dff_A_v8n0XNNu5_0;
	wire w_dff_A_Jo1ugJtU2_0;
	wire w_dff_A_HuFmlrno0_0;
	wire w_dff_A_W8Uej57R9_0;
	wire w_dff_A_kUCYf8kN2_0;
	wire w_dff_A_q113nbdl4_0;
	wire w_dff_A_uQdRHUcm2_0;
	wire w_dff_A_dn66hNLH8_0;
	wire w_dff_A_al6QU0vJ8_0;
	wire w_dff_A_SgCnDcuy9_0;
	wire w_dff_A_GmdPsuQo1_0;
	wire w_dff_A_cLtwMcub9_0;
	wire w_dff_A_KaPls0NG1_0;
	wire w_dff_A_AX3bxqO52_0;
	wire w_dff_A_ycP2fRZk4_0;
	wire w_dff_A_e8tZFNsW7_0;
	wire w_dff_A_D74tUqf23_0;
	wire w_dff_A_wEIpCUQT9_0;
	wire w_dff_A_Bo2UcP7W5_0;
	wire w_dff_A_5tmLieRe6_0;
	wire w_dff_A_iFw9RA5e3_0;
	wire w_dff_A_qpvyfEgP9_0;
	wire w_dff_A_VOzBRYgO8_0;
	wire w_dff_A_vbI13Ixl4_0;
	wire w_dff_A_gzmndNtt5_0;
	wire w_dff_A_rYllZkbH4_0;
	wire w_dff_A_30iM3TXy2_0;
	wire w_dff_A_I0MZ7KOz8_2;
	wire w_dff_A_cN3hT0l91_2;
	wire w_dff_A_mQ10DAUR1_2;
	wire w_dff_A_HEOQgHfq2_2;
	wire w_dff_A_nyssFGsN8_0;
	wire w_dff_A_xlQYpSbL7_0;
	wire w_dff_B_pPgfFLMk6_0;
	wire w_dff_B_crLlfJIw9_2;
	wire w_dff_B_yLX4YxfI0_2;
	wire w_dff_A_89EwIiis5_1;
	wire w_dff_A_4QrBMBET5_1;
	wire w_dff_A_6K5JmWpr5_1;
	wire w_dff_A_eWcErX501_1;
	wire w_dff_A_tv0ZjUZ57_1;
	wire w_dff_A_oVUZjhSq8_1;
	wire w_dff_A_3g6Hn5Wv6_1;
	wire w_dff_A_lD5UgCw14_1;
	wire w_dff_A_djG3bFr94_1;
	wire w_dff_A_fh94tmfL3_1;
	wire w_dff_A_AIwIqTYA4_1;
	wire w_dff_A_IEwPQ85E2_1;
	wire w_dff_A_OrKqRh162_1;
	wire w_dff_A_okEJVrfg6_1;
	wire w_dff_A_nw04RoSO9_1;
	wire w_dff_A_WmPSiICV0_1;
	wire w_dff_A_m7AHlMkS4_1;
	wire w_dff_A_VKcbacxA9_1;
	wire w_dff_A_ehaYp7VW2_1;
	wire w_dff_A_UBHMCOdy3_1;
	wire w_dff_A_jesx9sLH6_1;
	wire w_dff_A_PCNN4v9u3_1;
	wire w_dff_A_tSFY5sVH4_1;
	wire w_dff_A_hVxrw2tu1_1;
	wire w_dff_A_Mr3Sy99q2_1;
	wire w_dff_A_jD4VLyHv4_1;
	wire w_dff_A_ap7CsYDg3_1;
	wire w_dff_A_9jLdaajW3_1;
	wire w_dff_A_3hHbEkJw4_2;
	wire w_dff_A_8axD2BKd8_0;
	wire w_dff_A_LH9Vwqk78_0;
	wire w_dff_B_pvlpNQrM0_0;
	wire w_dff_A_4rk7qgCu2_1;
	wire w_dff_A_pev09nyh0_1;
	wire w_dff_A_guDKXsto8_2;
	wire w_dff_A_jXiXJTM48_2;
	wire w_dff_A_9yVFVzBQ3_1;
	wire w_dff_A_F7C2nutF1_1;
	wire w_dff_A_uDvPeQvH9_1;
	wire w_dff_A_frfO4gwx4_1;
	wire w_dff_A_WDOYyWZJ6_1;
	wire w_dff_A_snsW2rGW9_1;
	wire w_dff_A_UoATPuIy5_1;
	wire w_dff_A_cQUnQXGj7_1;
	wire w_dff_A_JZORpoAV6_1;
	wire w_dff_A_08ZtQnWK9_1;
	wire w_dff_A_zeoIeoUY5_1;
	wire w_dff_A_Y6WMetcc5_1;
	wire w_dff_A_FcIjmJT88_1;
	wire w_dff_A_2eb6slmX3_1;
	wire w_dff_A_0YdkfY6u0_1;
	wire w_dff_A_gGaIcq9W3_1;
	wire w_dff_A_kBnKYt0K2_1;
	wire w_dff_A_YcTFhvGB5_1;
	wire w_dff_A_kpUOp8HU8_1;
	wire w_dff_A_DepCaV7C1_1;
	wire w_dff_A_4TZPQH0r0_1;
	wire w_dff_A_3DskEiN37_1;
	wire w_dff_A_34dwUmOG1_1;
	wire w_dff_A_sRtAdeT96_1;
	wire w_dff_A_MNoAWPjX9_1;
	wire w_dff_A_8rxtEIsp6_1;
	wire w_dff_A_nmnVDEYr4_1;
	wire w_dff_A_hAWpOiWd7_1;
	wire w_dff_A_v8tUjL8T1_1;
	wire w_dff_A_05tgbhy02_1;
	wire w_dff_A_4MiPJ3LA3_1;
	wire w_dff_A_YgznzAnD1_1;
	wire w_dff_A_nfmxpdLb1_2;
	wire w_dff_A_ViNW4HgW0_2;
	wire w_dff_A_uUmampzn9_2;
	wire w_dff_A_FlRIwn5i0_2;
	wire w_dff_A_zbBR5lUA8_2;
	wire w_dff_A_U9vXyqPk9_2;
	wire w_dff_A_9jIVbu968_2;
	wire w_dff_A_sPaykXaM7_2;
	wire w_dff_A_BrJWuiaC8_2;
	wire w_dff_A_pBcZMKd46_2;
	wire w_dff_A_cbDPx23U4_2;
	wire w_dff_A_IM4vO9031_2;
	wire w_dff_A_7aLLXZtZ3_2;
	wire w_dff_A_thblUgG17_2;
	wire w_dff_A_v28JbT4a6_2;
	wire w_dff_A_3cqgQiJx0_2;
	wire w_dff_A_GKzDMjvo6_2;
	wire w_dff_A_ICIwWuyt6_2;
	wire w_dff_A_OeNZrCCi6_2;
	wire w_dff_A_kOs2V4Nv4_2;
	wire w_dff_A_ilpsLJRE7_2;
	wire w_dff_A_Br6KRhQR9_2;
	wire w_dff_A_FJAcj8Gr8_2;
	wire w_dff_A_loqtJTl15_2;
	wire w_dff_A_FOEQd2I65_2;
	wire w_dff_A_wbREUSQ84_2;
	wire w_dff_A_f32nalKt1_2;
	wire w_dff_A_Inqk3ZfN9_2;
	wire w_dff_A_QFFXqi4l6_1;
	wire w_dff_A_O5vJ67dP6_1;
	wire w_dff_A_EordcHI36_1;
	wire w_dff_A_KlMKcVk09_1;
	wire w_dff_A_NiwAgNE42_1;
	wire w_dff_A_i48I0sIY1_1;
	wire w_dff_A_zmM9YdNU5_1;
	wire w_dff_A_20t1uaI64_1;
	wire w_dff_A_Q55RE2jL8_1;
	wire w_dff_A_BQ9zBtmF0_1;
	wire w_dff_A_8yxk20K62_1;
	wire w_dff_A_zuVLIfE58_1;
	wire w_dff_A_hSSvffpZ8_1;
	wire w_dff_A_wPLjj0o73_1;
	wire w_dff_A_a3104nWL0_1;
	wire w_dff_A_WaqrZ3HL7_1;
	wire w_dff_A_Gvx5zwgd8_1;
	wire w_dff_A_4TlbubFC3_1;
	wire w_dff_A_N13YSZie3_1;
	wire w_dff_A_PnztjSvN8_1;
	wire w_dff_A_bFibu95c6_1;
	wire w_dff_A_2JN3ySKm1_1;
	wire w_dff_A_mgyvRonx9_1;
	wire w_dff_A_y2pkpJJP4_1;
	wire w_dff_A_VWfB6z6I2_1;
	wire w_dff_A_pyjGeP4F9_1;
	wire w_dff_A_2ltKX4H53_1;
	wire w_dff_A_DHeldumB4_1;
	wire w_dff_A_CSmNRdhO9_1;
	wire w_dff_A_NlcaFYkA4_0;
	wire w_dff_A_LlyypmAA3_0;
	wire w_dff_B_zfCEdJOT5_0;
	wire w_dff_A_BhsS0mFn0_1;
	wire w_dff_A_AczDAVgJ8_1;
	wire w_dff_A_7rlPCFmP0_2;
	wire w_dff_A_0BKpP0JF3_2;
	wire w_dff_A_iyFxE0WN7_1;
	wire w_dff_A_0p0bLv4h5_1;
	wire w_dff_A_rTrW1eUT5_1;
	wire w_dff_A_4GrWIc1s1_1;
	wire w_dff_A_NTQ1reO15_1;
	wire w_dff_A_IiPd0a298_1;
	wire w_dff_A_u0Xv4gTN7_1;
	wire w_dff_A_7nLFGb9G2_1;
	wire w_dff_A_PXQxivjl1_1;
	wire w_dff_A_NNCNc2w56_1;
	wire w_dff_A_jcUFpHuc8_1;
	wire w_dff_A_WDfCFM9k1_1;
	wire w_dff_A_v1AG3zii7_1;
	wire w_dff_A_EoMrbiIW1_1;
	wire w_dff_A_IkXlJV928_1;
	wire w_dff_A_TdtnEfxh9_1;
	wire w_dff_A_jHgTChG39_1;
	wire w_dff_A_5NzEaXDh7_1;
	wire w_dff_A_nEagDW6k0_1;
	wire w_dff_A_AjcqR7Yg2_1;
	wire w_dff_A_JDaC1WEL3_1;
	wire w_dff_A_Q1QpMwcF1_1;
	wire w_dff_A_ClCaIhFk2_1;
	wire w_dff_A_1yihF3513_1;
	wire w_dff_A_xn5aMBvj8_1;
	wire w_dff_A_6esJE98D4_1;
	wire w_dff_A_O2Q6WSYo9_1;
	wire w_dff_A_5LsLCVbA5_1;
	wire w_dff_A_ZZDoLTrp5_1;
	wire w_dff_A_f4VrnYDr7_1;
	wire w_dff_A_ton5okTs8_1;
	wire w_dff_A_alS2OU0O7_1;
	wire w_dff_A_NIIPZnVf3_0;
	wire w_dff_A_e43K4zLq2_0;
	wire w_dff_B_l5zNm9Gi9_0;
	wire w_dff_A_Ifa0eeTd3_1;
	wire w_dff_A_Dr6I3zdZ5_1;
	wire w_dff_A_NewWcorh8_2;
	wire w_dff_A_6dGCM4iH7_2;
	wire w_dff_A_DY1kktFA4_2;
	wire w_dff_A_Mwxo8oJu9_2;
	wire w_dff_A_QK14DYwA1_2;
	wire w_dff_A_rB8GOIbM9_2;
	wire w_dff_B_A4tUEeHk1_0;
	wire w_dff_B_DmC11cly1_2;
	wire w_dff_B_RleEmAtv9_2;
	wire w_dff_A_hpoEgCU05_0;
	wire w_dff_A_7eMha8en1_0;
	wire w_dff_A_RvVpfsPN9_0;
	wire w_dff_A_hwt4BvMM2_0;
	wire w_dff_B_103VmZWn5_1;
	wire w_dff_B_agReMxmj6_1;
	wire w_dff_B_93yrlnIL7_1;
	wire w_dff_B_plq1XYuG0_1;
	wire w_dff_B_zgrmvCJ14_1;
	wire w_dff_B_aAFM1OFQ8_1;
	wire w_dff_B_FbAYhA0K9_1;
	wire w_dff_B_rmoIH8jC0_1;
	wire w_dff_B_sPOB1pyl2_1;
	wire w_dff_B_6uk0RQrf1_1;
	wire w_dff_B_Kvf6QrTG2_1;
	wire w_dff_B_NUAUviSo4_1;
	wire w_dff_B_3oV9plvU5_1;
	wire w_dff_B_mDdB53xk4_1;
	wire w_dff_B_UjeyhpaG1_1;
	wire w_dff_B_IwQzJvZb6_0;
	wire w_dff_B_aT7TYaF82_0;
	wire w_dff_B_yjpXPO2h6_0;
	wire w_dff_B_uPo0wcI66_0;
	wire w_dff_B_z66APjTh5_0;
	wire w_dff_B_C8X1P6Dm0_0;
	wire w_dff_B_jYtn8H0s7_0;
	wire w_dff_B_mJfFUkk79_0;
	wire w_dff_B_fXaCUOCl5_0;
	wire w_dff_B_moMo4PEw5_0;
	wire w_dff_B_CCxRpgky9_0;
	wire w_dff_B_vAnRDzCG8_1;
	wire w_dff_B_tHfsW3vq4_1;
	wire w_dff_B_YY2AIPKe1_0;
	wire w_dff_B_X6ducswn4_0;
	wire w_dff_B_kTVk2DZi1_0;
	wire w_dff_B_TDlfsMvs7_0;
	wire w_dff_B_4oBtaw2G0_0;
	wire w_dff_B_IlZDseQj4_0;
	wire w_dff_B_fc44wMvx8_0;
	wire w_dff_A_TT291i8o6_0;
	wire w_dff_A_VhyWcYjA2_0;
	wire w_dff_A_sziBKZFJ9_0;
	wire w_dff_A_zUERrm125_0;
	wire w_dff_A_b1SzQC9W3_0;
	wire w_dff_A_732wFWfy2_0;
	wire w_dff_A_y1uIFPlM4_0;
	wire w_dff_A_GgwafJLG3_1;
	wire w_dff_A_NXy2NtW05_1;
	wire w_dff_A_FD2nd6Wv3_1;
	wire w_dff_A_8TwFusgJ7_1;
	wire w_dff_A_KCyGJCE62_1;
	wire w_dff_A_kaQ6s8Sg9_1;
	wire w_dff_A_7W0PCMHr4_1;
	wire w_dff_B_m84ttWlY6_0;
	wire w_dff_B_bt5CqlH54_0;
	wire w_dff_B_anNSMSO76_0;
	wire w_dff_B_uz5JdEPA2_0;
	wire w_dff_A_G5VoCGkp6_1;
	wire w_dff_A_J7u78SKN9_1;
	wire w_dff_A_UyfMFkSm2_1;
	wire w_dff_A_HgLKnW4C8_1;
	wire w_dff_A_oAA3E9by7_1;
	wire w_dff_A_lfbYJuDe3_1;
	wire w_dff_A_TKUk1gsn4_1;
	wire w_dff_B_8KIOEasC4_1;
	wire w_dff_B_waw4KLp83_1;
	wire w_dff_B_hDLAAMvA5_1;
	wire w_dff_B_KVrrMNTG3_1;
	wire w_dff_B_in5wwlVu7_1;
	wire w_dff_B_YuPztimZ1_1;
	wire w_dff_B_QRt6WBdp0_0;
	wire w_dff_B_One0Agdz9_0;
	wire w_dff_B_cX7DX5Th0_0;
	wire w_dff_A_ecD2UVhc6_1;
	wire w_dff_A_cOHiFweG9_1;
	wire w_dff_A_FekR1ssV9_1;
	wire w_dff_A_Q9SO47pB3_1;
	wire w_dff_A_aIS6u4cB4_1;
	wire w_dff_A_OvrM5F6E5_1;
	wire w_dff_A_02qyTdDV4_1;
	wire w_dff_A_EWnY6QVI2_1;
	wire w_dff_A_Wi9IFu6e2_1;
	wire w_dff_A_x9ng5r8N3_1;
	wire w_dff_A_JTN3oEue1_1;
	wire w_dff_A_rS5PolOt7_1;
	wire w_dff_A_agESjHom7_1;
	wire w_dff_A_Lbuzz2I51_1;
	wire w_dff_A_GpqMXNZU8_1;
	wire w_dff_B_pTgNxzNA1_0;
	wire w_dff_B_JwPkVB3w4_0;
	wire w_dff_B_FYsF2bfK2_1;
	wire w_dff_B_gCAW2DAF2_1;
	wire w_dff_B_CFxhFbna6_1;
	wire w_dff_B_58RorVq24_1;
	wire w_dff_B_cIwl27WB0_1;
	wire w_dff_B_hLttKi5x0_1;
	wire w_dff_B_iO8JwX4U0_1;
	wire w_dff_B_1kx18BGy0_1;
	wire w_dff_B_odRQHQ3C6_1;
	wire w_dff_B_LXOtIWEn4_1;
	wire w_dff_B_UiFwSTNy9_1;
	wire w_dff_B_nRC0Yr099_1;
	wire w_dff_B_TmRP1p7q3_0;
	wire w_dff_A_nIsRN38t6_1;
	wire w_dff_B_d2XB5cjq2_2;
	wire w_dff_B_B4ZEY8c77_2;
	wire w_dff_B_LTthsse71_0;
	wire w_dff_B_WdonE3CV6_0;
	wire w_dff_B_KphS10fo0_0;
	wire w_dff_B_kAHKnmBg9_0;
	wire w_dff_B_jn8IgKiS4_0;
	wire w_dff_B_Xh53Gc1B2_1;
	wire w_dff_B_4MLFFKzK1_1;
	wire w_dff_B_vpfiJFkd0_1;
	wire w_dff_A_iAdNOIPv3_0;
	wire w_dff_A_JoU9a7Oq1_0;
	wire w_dff_A_9uE2buWy8_0;
	wire w_dff_A_z6sf7Fkn6_0;
	wire w_dff_A_EAxVI1FH9_1;
	wire w_dff_A_eGotZmrQ3_1;
	wire w_dff_A_NNu9KYcg2_1;
	wire w_dff_A_D1LYb21k7_1;
	wire w_dff_A_pSgudIjE3_1;
	wire w_dff_A_1wY814jb9_1;
	wire w_dff_A_ZryUnmGD4_1;
	wire w_dff_A_36IVZN5a9_1;
	wire w_dff_A_yPI8eKWu7_1;
	wire w_dff_A_63KGx8rG5_1;
	wire w_dff_A_8SRdCOxw0_1;
	wire w_dff_A_q3UANLk35_1;
	wire w_dff_A_hEif0nC70_1;
	wire w_dff_A_AmjgDKJK9_1;
	wire w_dff_A_OLJlUU8w0_1;
	wire w_dff_A_ZZCWqlCV2_1;
	wire w_dff_B_FCmJPHfS7_0;
	wire w_dff_B_td1CobWD0_0;
	wire w_dff_B_x6SATIH07_0;
	wire w_dff_B_ryPHwt8F6_0;
	wire w_dff_B_d2U7s5oQ6_0;
	wire w_dff_B_oaIbomvf7_0;
	wire w_dff_B_aaz4RO4F3_0;
	wire w_dff_A_Wi6E2LJo4_1;
	wire w_dff_A_9nftVOMq4_1;
	wire w_dff_A_cyHA4Zav3_1;
	wire w_dff_A_Qg8qfCDN1_1;
	wire w_dff_A_pLDhhI3T2_1;
	wire w_dff_A_g2n6lwlj0_1;
	wire w_dff_A_fPjZS4nm8_1;
	wire w_dff_A_3utLmtf54_1;
	wire w_dff_A_WPovrqbZ6_1;
	wire w_dff_A_5CgJH34Z8_1;
	wire w_dff_A_px9vcTcr0_1;
	wire w_dff_A_OEHqpfUh9_1;
	wire w_dff_A_v1SmNGQr8_1;
	wire w_dff_A_IgszziJX7_1;
	wire w_dff_A_3vVToo9h8_1;
	wire w_dff_A_67SlbUFS4_1;
	wire w_dff_A_GSGGZwE50_1;
	wire w_dff_A_mN7i3Yrl0_1;
	wire w_dff_A_DFF7w8UG3_1;
	wire w_dff_A_9ELLg1NZ1_1;
	wire w_dff_B_XYDuZhvK7_2;
	wire w_dff_A_9g2qfnBI4_2;
	wire w_dff_B_OjPSi83b8_1;
	wire w_dff_B_hevlZQKt0_0;
	wire w_dff_A_AZjeSlZO9_0;
	wire w_dff_A_jggx32xI4_0;
	wire w_dff_A_Tuk0jMnd9_2;
	wire w_dff_A_2cU5pr8u4_2;
	wire w_dff_A_7yLK3So26_1;
	wire w_dff_A_akYgauwP8_1;
	wire w_dff_A_1s9AXgTT6_1;
	wire w_dff_A_4CLa4k1Y8_1;
	wire w_dff_A_0KLLPL4s9_1;
	wire w_dff_A_pvdZHmJR1_1;
	wire w_dff_A_8YpAQu4S6_1;
	wire w_dff_A_S3pMlIGa0_1;
	wire w_dff_A_EXrf9peh3_1;
	wire w_dff_A_NILS2dXM9_1;
	wire w_dff_A_rMlBMTFf2_1;
	wire w_dff_A_NCqt1J6M7_1;
	wire w_dff_A_7c2tpUQI9_1;
	wire w_dff_A_p8haoUJq4_1;
	wire w_dff_A_lmL2Uuze4_1;
	wire w_dff_A_PDstxXkQ3_1;
	wire w_dff_A_gUul2mw15_1;
	wire w_dff_A_voPurD9a3_1;
	wire w_dff_A_Rdj7FWHn1_1;
	wire w_dff_A_zlS3VSDO0_1;
	wire w_dff_A_powAz74V9_0;
	wire w_dff_A_PbcLaPLQ3_1;
	wire w_dff_A_RExE2HPu3_1;
	wire w_dff_A_prtf9rx73_1;
	wire w_dff_A_YMpjr2zA1_1;
	wire w_dff_A_pytR5S3c5_1;
	wire w_dff_A_gj1an2Kd8_1;
	wire w_dff_A_NDBWt4Gi7_1;
	wire w_dff_A_x0vXnbmk4_1;
	wire w_dff_A_gjE7Cwl60_1;
	wire w_dff_A_EWvrhSlB1_1;
	wire w_dff_A_d3yFPxrF5_1;
	wire w_dff_A_gk5TTWpK9_1;
	wire w_dff_A_alYCBDb98_1;
	wire w_dff_A_zcKipE6K2_1;
	wire w_dff_A_6ToQmENd2_1;
	wire w_dff_B_mkdFzHJL4_0;
	wire w_dff_A_xgd73YNd1_0;
	wire w_dff_A_EwimlYRb6_0;
	wire w_dff_A_IojLoow58_0;
	wire w_dff_A_KWRn9VrQ3_0;
	wire w_dff_A_Bg8ECj7Q6_0;
	wire w_dff_A_J61Cz9ao4_0;
	wire w_dff_A_pDZnYLP57_0;
	wire w_dff_A_QjDMdVsT3_0;
	wire w_dff_A_MqXFakvJ1_0;
	wire w_dff_A_9JHRMoDA2_0;
	wire w_dff_A_SybwssI75_0;
	wire w_dff_A_8KsBEpC97_0;
	wire w_dff_A_bPfJXG0X2_0;
	wire w_dff_A_euClOofw5_0;
	wire w_dff_A_xOFp0yv78_0;
	wire w_dff_A_35YdLmI60_0;
	wire w_dff_A_s4tbPafp6_0;
	wire w_dff_A_q5tRPNSs9_0;
	wire w_dff_B_zif2k5jg5_1;
	wire w_dff_A_Dj3DA7wv9_2;
	wire w_dff_A_7Tau7gTA6_2;
	wire w_dff_A_gicobGyc3_2;
	wire w_dff_A_w1ybD9kK7_2;
	wire w_dff_A_ds8IdZiz7_2;
	wire w_dff_A_0cnjByHZ7_2;
	wire w_dff_A_zOr7Kzy26_2;
	wire w_dff_A_rZ8T6MVo3_2;
	wire w_dff_A_fwufgFKK9_2;
	wire w_dff_A_8eEiDzOi0_2;
	wire w_dff_A_eveQR6kS6_2;
	wire w_dff_A_q3PuDnq04_2;
	wire w_dff_A_u52IRCK89_2;
	wire w_dff_A_9eJ9HbSg4_2;
	wire w_dff_A_vSC06nqv4_2;
	wire w_dff_A_hafLcM778_2;
	wire w_dff_A_E8kYfVRo1_2;
	wire w_dff_A_ijuTNTL78_0;
	wire w_dff_A_6Z1d3v7H1_0;
	wire w_dff_A_BXjGEBES7_0;
	wire w_dff_A_fdpv6NKn2_0;
	wire w_dff_A_HRaddUvR5_0;
	wire w_dff_A_sENznjUR7_0;
	wire w_dff_A_6ITc35Vn3_0;
	wire w_dff_A_jvKDct7U9_0;
	wire w_dff_A_66c7i4qM5_0;
	wire w_dff_A_P7wMnUqo9_0;
	wire w_dff_A_JbXlZfCK4_0;
	wire w_dff_A_RLwTPzdA1_0;
	wire w_dff_A_BouNLdYb9_0;
	wire w_dff_A_9M46Ac4o7_0;
	wire w_dff_A_B8cVVLXC0_0;
	wire w_dff_A_rITaSCkS6_0;
	wire w_dff_A_ndPhYgKa6_0;
	wire w_dff_A_5oso5I1j9_0;
	wire w_dff_B_kgtB5zK48_1;
	wire w_dff_B_6Hnef3P70_0;
	wire w_dff_B_qEqpUElT1_2;
	wire w_dff_B_V2dp9oao7_2;
	wire w_dff_A_O38cRWwB9_0;
	wire w_dff_A_bqzeMAZm9_0;
	wire w_dff_A_b5cgMnwu5_0;
	wire w_dff_A_HBJIOJCi0_0;
	wire w_dff_B_1uxc9meZ2_1;
	wire w_dff_B_FI8IhTCi2_0;
	wire w_dff_B_Ku9p1LZk8_2;
	wire w_dff_B_9w2r0qCf1_2;
	wire w_dff_A_cBpxTyuL7_1;
	wire w_dff_B_stDaMQtR2_2;
	wire w_dff_A_JOmmXEPd3_2;
	wire w_dff_A_lvSU19PP7_2;
	wire w_dff_A_Z9nIQoCp2_2;
	wire w_dff_A_H8YYUOsO4_2;
	wire w_dff_A_mEQNs6C42_2;
	wire w_dff_B_eprve7413_1;
	wire w_dff_B_kh9eKsd88_0;
	wire w_dff_A_5S4Af8175_1;
	wire w_dff_A_iDCFiOTb3_1;
	wire w_dff_A_KCLPAnYJ7_2;
	wire w_dff_A_eBZdL6T88_2;
	wire w_dff_A_nRpXKqVf5_1;
	wire w_dff_A_etaTxasj8_1;
	wire w_dff_A_6hNQKIf72_1;
	wire w_dff_A_7nXfocmh8_1;
	wire w_dff_A_tTzWUmWD5_1;
	wire w_dff_A_JQtcVcW30_1;
	wire w_dff_A_GUwOCB6M5_1;
	wire w_dff_A_HnVWsxJd4_1;
	wire w_dff_A_ckG5mk5n5_1;
	wire w_dff_A_cBVGppdq7_1;
	wire w_dff_A_b5O9x9WL1_1;
	wire w_dff_A_ChrPDoUt9_1;
	wire w_dff_A_kxNOyO7N4_1;
	wire w_dff_B_Ik4vbIEX3_1;
	wire w_dff_B_QQ6alOl00_1;
	wire w_dff_B_X2FDpMm36_1;
	wire w_dff_B_MHByK6Eq9_1;
	wire w_dff_B_iYETiQbB5_1;
	wire w_dff_B_Venm6auk9_1;
	wire w_dff_B_qb6YZBQ74_1;
	wire w_dff_B_NzvuBmVy4_1;
	wire w_dff_B_BEuDBo4u4_1;
	wire w_dff_B_0kqVoX2y3_1;
	wire w_dff_B_vNMvTpCU8_1;
	wire w_dff_B_Nlt59Phy8_1;
	wire w_dff_B_RyXZpfk67_1;
	wire w_dff_B_4PI7nKJX5_1;
	wire w_dff_B_DkdIHtIg6_1;
	wire w_dff_A_PMlK8EoZ3_1;
	wire w_dff_A_NNm5HebY3_1;
	wire w_dff_A_vFPzkZcD1_1;
	wire w_dff_A_IRf6ExwL3_1;
	wire w_dff_A_rNK7SLuU1_1;
	wire w_dff_A_CE8TZrZ11_1;
	wire w_dff_A_vtLg4Pz35_1;
	wire w_dff_B_YrCqxNbT4_1;
	wire w_dff_B_SB8hL7Ki5_1;
	wire w_dff_B_gUpevgBD3_1;
	wire w_dff_B_HE2ZpfZg5_1;
	wire w_dff_B_UcisGcxM6_1;
	wire w_dff_B_N4pNtpjI3_1;
	wire w_dff_B_iu005BEr3_1;
	wire w_dff_B_RA7GSw6j4_1;
	wire w_dff_B_gopcol739_1;
	wire w_dff_B_wxZYj8iP6_1;
	wire w_dff_B_FeOV8fMy1_1;
	wire w_dff_B_QAni6bGw5_1;
	wire w_dff_B_M54LwU609_1;
	wire w_dff_A_vJugByyt6_0;
	wire w_dff_A_BaT3VEvH7_0;
	wire w_dff_A_0ZUkzLIF1_0;
	wire w_dff_A_blumDytY3_0;
	wire w_dff_A_Kd3z0hum8_0;
	wire w_dff_A_V6ue6u8k0_0;
	wire w_dff_A_ebunmQqZ3_0;
	wire w_dff_A_LjYP9uA77_0;
	wire w_dff_A_SzYy73Gq8_0;
	wire w_dff_A_vXJCbXxc0_0;
	wire w_dff_A_SFSrMxs73_0;
	wire w_dff_A_N94m8ke02_1;
	wire w_dff_A_8SPwT7SL5_1;
	wire w_dff_A_AlL3C5b40_1;
	wire w_dff_A_G5mp3rok0_1;
	wire w_dff_A_DxZAQzaO9_1;
	wire w_dff_A_YMitZxPN7_1;
	wire w_dff_A_tc6v9mLJ2_1;
	wire w_dff_A_D7MDysKd6_1;
	wire w_dff_A_4a1uEYYr2_1;
	wire w_dff_A_3oJZCltt9_1;
	wire w_dff_A_LQDSPVtc1_1;
	wire w_dff_A_iGsFYc2f1_1;
	wire w_dff_A_8ygS51Vp9_1;
	wire w_dff_A_tZIMvvsQ3_1;
	wire w_dff_A_9eFk9Aht4_1;
	wire w_dff_A_bvENYMJC6_2;
	wire w_dff_A_8HZhCT4c0_2;
	wire w_dff_A_QLaHShLO6_0;
	wire w_dff_A_wYCagy7e1_1;
	wire w_dff_A_BA1F0Zgy1_2;
	wire w_dff_A_EzDBjIMm5_2;
	wire w_dff_A_JTbuxVf88_2;
	wire w_dff_A_dPBMJ54I4_0;
	wire w_dff_A_6RKzcdbo6_0;
	wire w_dff_A_3cuPesp66_0;
	wire w_dff_A_Z193WOGo5_0;
	wire w_dff_A_KhFQ59lS2_0;
	wire w_dff_A_C08UO7vJ2_1;
	wire w_dff_A_p8TbQbTy4_1;
	wire w_dff_A_4S11vnnI9_1;
	wire w_dff_A_TZznZrcF6_1;
	wire w_dff_A_VK935xeR7_1;
	wire w_dff_A_Lsy9KzB41_1;
	wire w_dff_A_7hPF4fB09_1;
	wire w_dff_B_KJ16u6mD3_2;
	wire w_dff_B_CVqjWA7C4_2;
	wire w_dff_B_7Y9ChrHQ0_2;
	wire w_dff_B_aHyXyoDH8_2;
	wire w_dff_B_iZ6gBjLr1_2;
	wire w_dff_B_E97Us8X46_2;
	wire w_dff_B_K5x5SohI6_2;
	wire w_dff_B_cMRHQBCL1_2;
	wire w_dff_A_ysMVdwFZ3_0;
	wire w_dff_A_gPzslvf37_0;
	wire w_dff_A_vuvPEHOq4_0;
	wire w_dff_A_6AioAxSI3_0;
	wire w_dff_A_PWTQCgE72_0;
	wire w_dff_A_vCz0QbXB2_0;
	wire w_dff_A_kU1oxVam1_0;
	wire w_dff_A_71DzBzYo3_2;
	wire w_dff_A_3sBOF4St6_2;
	wire w_dff_A_dB2iJaPX3_2;
	wire w_dff_A_p9pMCzO73_2;
	wire w_dff_A_p3KhwOOd0_2;
	wire w_dff_A_W2jkEVHY0_2;
	wire w_dff_A_oTKXff7P4_2;
	wire w_dff_A_miJ4WaIk0_2;
	wire w_dff_A_IZiN2qeO5_2;
	wire w_dff_A_GY5bjR3s4_2;
	wire w_dff_A_GXXDDDUQ5_2;
	wire w_dff_A_2Cawg4TM3_0;
	wire w_dff_A_xgz65GIG9_0;
	wire w_dff_A_Wfs2Q56b3_0;
	wire w_dff_A_t67qWl7n1_0;
	wire w_dff_A_kCaYLmSo8_0;
	wire w_dff_A_CugJAFDh4_0;
	wire w_dff_A_l2nWqKwK2_0;
	wire w_dff_A_IAVF5e637_1;
	wire w_dff_A_pkWrhgyj1_1;
	wire w_dff_A_azkasoZy5_1;
	wire w_dff_A_6d1kYrZC2_1;
	wire w_dff_A_BvaK4DRU8_1;
	wire w_dff_A_M2QEomtA6_1;
	wire w_dff_A_CZEXJRqe6_1;
	wire w_dff_A_4esIxRVH1_1;
	wire w_dff_A_5xWiSkwM3_1;
	wire w_dff_A_L9qQU0RR2_1;
	wire w_dff_A_k2kAb4RG9_1;
	wire w_dff_A_mon5JnRv2_1;
	wire w_dff_A_lqffWO2G4_0;
	wire w_dff_A_acD5kKi72_1;
	wire w_dff_A_B8ZxuV172_1;
	wire w_dff_A_Au93wacp1_1;
	wire w_dff_A_3gxpf3SG0_1;
	wire w_dff_A_CUgKotio2_1;
	wire w_dff_A_JmJgEfVy3_1;
	wire w_dff_A_9j9WAkp86_1;
	wire w_dff_A_UhJAmNbx4_1;
	wire w_dff_A_W0e2XS114_1;
	wire w_dff_A_SJvgTQ1q5_1;
	wire w_dff_A_kOxryNfs6_1;
	wire w_dff_A_OpJIBC5E1_1;
	wire w_dff_A_zYOezuNr4_1;
	wire w_dff_A_tXO1PP5z8_1;
	wire w_dff_A_yeAsge4y4_1;
	wire w_dff_A_0TdKwvQd0_1;
	wire w_dff_B_qIPZoZRM4_1;
	wire w_dff_B_Riboc5A53_0;
	wire w_dff_B_XccfJ9tn6_2;
	wire w_dff_B_ihvAxHVv3_2;
	wire w_dff_A_xgTb31pd1_0;
	wire w_dff_A_v88eWpYU9_0;
	wire w_dff_A_1WAWknsy7_0;
	wire w_dff_A_lTrelQPG1_0;
	wire w_dff_B_dQ2S0xJ08_1;
	wire w_dff_B_p60qXJgH6_0;
	wire w_dff_A_f9O9ovBw2_1;
	wire w_dff_A_dLMjmZVF5_1;
	wire w_dff_A_1px5iE7k2_2;
	wire w_dff_A_TgcstwJn7_2;
	wire w_dff_A_jCIFrJNW2_1;
	wire w_dff_A_7Htipfr83_1;
	wire w_dff_A_XpHdLBPY4_1;
	wire w_dff_A_9wSeb58Q6_1;
	wire w_dff_A_N3WShLZG1_0;
	wire w_dff_A_DvtYQeO81_0;
	wire w_dff_A_4FiJ6Abm9_0;
	wire w_dff_A_kabXAEER0_0;
	wire w_dff_A_PPGF0MwR1_0;
	wire w_dff_A_PNH8FUOz4_0;
	wire w_dff_A_sNYJcCNi8_0;
	wire w_dff_A_kB8hMKWp6_0;
	wire w_dff_A_u3019IJd7_0;
	wire w_dff_A_wcaFuKEE8_0;
	wire w_dff_A_bGViTR6f4_0;
	wire w_dff_A_a9XS4HMB7_0;
	wire w_dff_A_hz18Lgjr9_0;
	wire w_dff_A_NvpZ0mFy4_0;
	wire w_dff_A_WVd6taLi7_0;
	wire w_dff_A_UHRhb0km1_0;
	wire w_dff_A_8o1EvQQ89_0;
	wire w_dff_A_DPHt0NE36_0;
	wire w_dff_A_amYwbKsM0_0;
	wire w_dff_A_Wq2N3hnR2_0;
	wire w_dff_A_V1PNa2iC3_0;
	wire w_dff_A_IkU1o7ym0_0;
	wire w_dff_A_fwOiAooC4_0;
	wire w_dff_A_OvfXvPDW2_0;
	wire w_dff_A_D2ClmSTB0_0;
	wire w_dff_A_BEQMLTWM3_0;
	wire w_dff_A_8x3bmntu0_0;
	wire w_dff_A_p4US44f95_2;
	wire w_dff_A_u22XtAVW7_2;
	wire w_dff_A_736VvCll4_2;
	wire w_dff_A_nlQeMzFL1_2;
	wire w_dff_A_pundBuOL3_2;
	wire w_dff_A_rSR9TcK67_2;
	wire w_dff_A_uweABs4V3_2;
	wire w_dff_A_Jnt2VpNM3_2;
	wire w_dff_A_hUGxjfsN8_2;
	wire w_dff_A_2HpiObd17_2;
	wire w_dff_A_xAiIsYas7_2;
	wire w_dff_A_atlK1W1j0_2;
	wire w_dff_A_YRz67tca0_2;
	wire w_dff_A_7r7a95wO4_2;
	wire w_dff_B_5J78YsqT1_1;
	wire w_dff_B_3iz5PsYf1_0;
	wire w_dff_B_VwWmTBK90_2;
	wire w_dff_B_7TqLiHyu6_2;
	wire w_dff_A_Pkfnl6f13_2;
	wire w_dff_A_iuaibS5Y5_2;
	wire w_dff_A_yzUKPOdA1_2;
	wire w_dff_A_IutNNJpv4_2;
	wire w_dff_A_OC50sEMX8_1;
	wire w_dff_A_jAzB48uU8_1;
	wire w_dff_A_Av1rnJiU2_1;
	wire w_dff_A_RaQj24hW2_1;
	wire w_dff_A_bW3y7cdp8_1;
	wire w_dff_A_e4WQQvfR9_1;
	wire w_dff_A_MVe4SJEJ1_1;
	wire w_dff_A_B2WhMACO0_1;
	wire w_dff_A_SZ5m0Uam4_1;
	wire w_dff_A_sOGc9nEV3_1;
	wire w_dff_A_S9zR2MoY0_1;
	wire w_dff_A_DxrbamLN8_1;
	wire w_dff_A_ddPo7jrP3_1;
	wire w_dff_A_fVl5iCD92_1;
	wire w_dff_A_b6AGPVkI5_1;
	wire w_dff_A_ygwklOHH0_1;
	wire w_dff_B_38xGnxtj6_1;
	wire w_dff_B_7tTp421h9_0;
	wire w_dff_B_PVbhmyMo4_2;
	wire w_dff_B_BCtcMeMM9_2;
	wire w_dff_A_xmQWixmU5_0;
	wire w_dff_A_jNF1ql180_0;
	wire w_dff_A_Og3rJbXB4_0;
	wire w_dff_A_sFIkmB0G0_0;
	wire w_dff_A_7fuK7RtU0_0;
	wire w_dff_A_6izLRkuO9_0;
	wire w_dff_A_rXlwLnIN3_0;
	wire w_dff_A_T1k0BBKT5_0;
	wire w_dff_A_E6ImUlFE7_0;
	wire w_dff_A_yPefPCJk6_0;
	wire w_dff_A_tz40ulXB7_0;
	wire w_dff_A_42BOIvwl5_0;
	wire w_dff_A_fuCPdAOi6_0;
	wire w_dff_A_kEQhtFmE3_0;
	wire w_dff_A_Glr05qO79_0;
	wire w_dff_A_C08EW8Rb1_0;
	wire w_dff_A_qittnX8T7_0;
	wire w_dff_A_LvjM02uI6_0;
	wire w_dff_A_hLOoceXz1_1;
	wire w_dff_A_oYqyl08q4_1;
	wire w_dff_A_MNSi9QRU8_1;
	wire w_dff_A_mvKoU86b7_2;
	wire w_dff_A_tuR61V1o1_2;
	wire w_dff_B_9C4K4mYd5_3;
	wire w_dff_B_8mpWh9QD7_3;
	wire w_dff_B_t9qFBe8s0_1;
	wire w_dff_B_kRuWr5Ze3_0;
	wire w_dff_B_N7qyj0SS7_2;
	wire w_dff_B_O4P7ekHV9_2;
	wire w_dff_A_0KBxwsSj2_0;
	wire w_dff_A_aLmk8uKN5_0;
	wire w_dff_A_jyj8FSGN1_0;
	wire w_dff_A_lnZFptbP4_0;
	wire w_dff_B_1MnPFWTn6_1;
	wire w_dff_B_CzRc0bBz7_1;
	wire w_dff_B_e2BLbAhW4_1;
	wire w_dff_B_UDhXF6iJ1_1;
	wire w_dff_B_BEhZtLA78_1;
	wire w_dff_B_BoOkr2Ex8_1;
	wire w_dff_B_kc1tfybA7_1;
	wire w_dff_B_O1q6X0h10_1;
	wire w_dff_B_jdSfgv1h5_1;
	wire w_dff_B_88xv0lQT3_1;
	wire w_dff_B_ldq4NBgL5_1;
	wire w_dff_B_xycWIFKM6_1;
	wire w_dff_B_WyXqx9GF2_1;
	wire w_dff_B_Sf0ECSPo6_1;
	wire w_dff_B_eVzLRdWj1_1;
	wire w_dff_B_1qfAXtC86_1;
	wire w_dff_B_nguaJ4fU0_1;
	wire w_dff_B_Ok5coIGX5_1;
	wire w_dff_A_FBA4pPba7_0;
	wire w_dff_A_SMOczHxq3_0;
	wire w_dff_A_BzVI7Hmc4_0;
	wire w_dff_A_otTBf6UK0_1;
	wire w_dff_A_t8eUGYfF0_1;
	wire w_dff_A_mFwHVCmR1_1;
	wire w_dff_A_B4YaPbWH1_1;
	wire w_dff_A_EaGWucWr5_1;
	wire w_dff_A_1g1knSvq5_1;
	wire w_dff_A_KEpOUmLI6_1;
	wire w_dff_A_Z9KREoSp5_0;
	wire w_dff_A_cQ64OiLb2_0;
	wire w_dff_A_jwrJUxZu5_0;
	wire w_dff_A_YAzPImYi1_0;
	wire w_dff_A_0D7DRRfH4_0;
	wire w_dff_A_qSCmXCoz6_0;
	wire w_dff_A_9ieRz2IT8_0;
	wire w_dff_A_ulwkfI8V2_0;
	wire w_dff_A_I9cviMoA4_0;
	wire w_dff_A_rE0JRAc74_0;
	wire w_dff_A_RjDBOhul3_0;
	wire w_dff_A_KNCJspG11_1;
	wire w_dff_A_Rb3tevW70_1;
	wire w_dff_A_YLKPixlB3_1;
	wire w_dff_A_2EbvKKd93_1;
	wire w_dff_A_hxTGiEPx4_1;
	wire w_dff_A_GiUdOuoH4_1;
	wire w_dff_A_ZO06GEhO5_1;
	wire w_dff_A_OJGNnBwV2_1;
	wire w_dff_A_7qzebuRD8_1;
	wire w_dff_A_vsLeinxy3_1;
	wire w_dff_A_FUS7ZetH6_1;
	wire w_dff_A_wcIRTCIK3_1;
	wire w_dff_A_2tPgZb2z2_1;
	wire w_dff_A_McxqYnwG5_2;
	wire w_dff_A_eXL2fdfm5_2;
	wire w_dff_A_WDwcHOGF9_2;
	wire w_dff_A_Oc5dMlRx2_2;
	wire w_dff_A_aKAJ4X310_2;
	wire w_dff_A_hU48JwK29_2;
	wire w_dff_A_Cn0Vxd4t7_2;
	wire w_dff_A_t8LjUqfe9_2;
	wire w_dff_A_RqBsZQBk7_2;
	wire w_dff_A_i9EFuq3a5_2;
	wire w_dff_A_45OF1Ef03_2;
	wire w_dff_A_CYddlKxF6_2;
	wire w_dff_A_WKfWzS9X7_2;
	wire w_dff_B_a7EzQSxI7_0;
	wire w_dff_B_T3gQHh6T4_0;
	wire w_dff_B_CfL1mf701_0;
	wire w_dff_B_96jNs8Ki9_0;
	wire w_dff_B_BJI2hD937_0;
	wire w_dff_B_6qVgfeOH7_0;
	wire w_dff_B_8AUtE38n6_0;
	wire w_dff_B_mNlrzDub2_0;
	wire w_dff_B_CuGglQsX9_0;
	wire w_dff_B_yktIWuvJ8_0;
	wire w_dff_B_3p4fg0Jy6_0;
	wire w_dff_B_HUTbIaS43_1;
	wire w_dff_B_ngg18DwO4_1;
	wire w_dff_B_rJyFWDR91_1;
	wire w_dff_A_KF6NnfZB2_0;
	wire w_dff_A_tNhpBkgq5_0;
	wire w_dff_B_zRmf5Vmx7_0;
	wire w_dff_B_0ZuZZlVW5_0;
	wire w_dff_B_kradYcl35_1;
	wire w_dff_B_R2AitHJL1_1;
	wire w_dff_B_Ak1eFJ806_1;
	wire w_dff_B_uud4iB130_0;
	wire w_dff_B_XkQg6ELH9_0;
	wire w_dff_B_oGy0A1gd7_0;
	wire w_dff_B_DeW867u91_0;
	wire w_dff_B_YhKwkhYb7_0;
	wire w_dff_A_4kWqaBCf0_0;
	wire w_dff_A_zAzTDnyc4_0;
	wire w_dff_A_WUvdjBcC0_0;
	wire w_dff_B_2Jgxhcxe8_0;
	wire w_dff_A_bDMyFFig2_0;
	wire w_dff_A_feYm9Cay4_0;
	wire w_dff_A_6n6nbIef7_0;
	wire w_dff_A_TuTJ2ZQJ1_0;
	wire w_dff_A_qHTQzuGI7_0;
	wire w_dff_B_oHa9ooEO4_0;
	wire w_dff_B_AkmfGLxS3_1;
	wire w_dff_A_bu5l24mo1_1;
	wire w_dff_B_2qDZexht2_2;
	wire w_dff_B_wFidWInp6_0;
	wire w_dff_B_2hPWlplO9_0;
	wire w_dff_B_BZvg9vHT9_0;
	wire w_dff_B_kzPwRbqB8_0;
	wire w_dff_B_veFixvxm7_0;
	wire w_dff_A_xbYiXmtF2_1;
	wire w_dff_A_TjyU1OXs3_1;
	wire w_dff_A_oB7sxDnQ9_1;
	wire w_dff_A_8sBd1jj22_1;
	wire w_dff_A_ZXN5ixdo4_1;
	wire w_dff_A_BWNUhscW4_1;
	wire w_dff_A_LXIdQTAd3_1;
	wire w_dff_A_DhEd4Yhf6_1;
	wire w_dff_A_YPCb7Y197_1;
	wire w_dff_A_7QPIrrcj9_1;
	wire w_dff_A_i5KSLdrG3_1;
	wire w_dff_A_sSgBY74Z6_1;
	wire w_dff_A_hoDPsrQ82_1;
	wire w_dff_A_tp6F6lUs4_1;
	wire w_dff_A_nT099fAz5_1;
	wire w_dff_B_eZX0uqCU7_1;
	wire w_dff_B_ZbK3sXt04_1;
	wire w_dff_A_XiAuJxIm0_0;
	wire w_dff_A_y5kFTxXt5_0;
	wire w_dff_A_FxK24AHN5_0;
	wire w_dff_A_6EreClJn7_0;
	wire w_dff_A_Kz2uNPy41_0;
	wire w_dff_B_0UPOrKaP0_1;
	wire w_dff_B_hy0ml6fJ9_1;
	wire w_dff_A_eBmxvIUd3_0;
	wire w_dff_A_VLtttGbJ4_0;
	wire w_dff_A_mzrBUT0E4_1;
	wire w_dff_A_9XOtSCNm2_1;
	wire w_dff_A_njp2cFh33_1;
	wire w_dff_A_0PcztyWg5_1;
	wire w_dff_A_AX8YAVEV9_1;
	wire w_dff_A_QO3Ew3Hl7_1;
	wire w_dff_A_qsGsNXAh3_1;
	wire w_dff_A_n6YmIM1H6_1;
	wire w_dff_A_lUsHpICq5_1;
	wire w_dff_A_C2x1klrX5_0;
	wire w_dff_A_rMM9sWQL4_0;
	wire w_dff_A_3b07Xonv3_0;
	wire w_dff_A_MqzgzvAT4_0;
	wire w_dff_A_WYCJ9KX06_0;
	wire w_dff_A_GzP3BLua7_0;
	wire w_dff_A_tKkvh8lj4_0;
	wire w_dff_A_v394gfxm8_0;
	wire w_dff_A_EusGPNz78_0;
	wire w_dff_A_fpwKEp9r3_0;
	wire w_dff_A_MqdtD7bv8_1;
	wire w_dff_A_HL4xyrhO9_1;
	wire w_dff_A_am7P2UTf1_1;
	wire w_dff_A_3ZRPYQxP9_1;
	wire w_dff_A_2l3z9mCJ6_1;
	wire w_dff_A_zcN8Ytqm3_1;
	wire w_dff_A_ZeXlIfVU6_1;
	wire w_dff_A_IYz19oPn3_1;
	wire w_dff_A_OCLlUMon3_1;
	wire w_dff_A_OziQOkLQ4_1;
	wire w_dff_A_Xv9SHgSe6_1;
	wire w_dff_A_hJkd0q0H7_1;
	wire w_dff_A_uLJhR1De9_2;
	wire w_dff_B_bFXeCJWI1_1;
	wire w_dff_B_P2NvOeP18_1;
	wire w_dff_B_SPEF7vWy2_1;
	wire w_dff_B_C1GdZ4kY1_1;
	wire w_dff_A_Bwd6QaoA3_0;
	wire w_dff_A_S7RxhA6h0_0;
	wire w_dff_A_k4tZXlm27_0;
	wire w_dff_B_okLIaUll6_2;
	wire w_dff_A_g3iSUOi77_1;
	wire w_dff_A_g47FT1Sz5_1;
	wire w_dff_A_R2bpxslN8_1;
	wire w_dff_A_fUruxAvU7_1;
	wire w_dff_A_lqYBdj6U0_2;
	wire w_dff_B_QnNTBcV28_1;
	wire w_dff_A_eMdK6NeO2_1;
	wire w_dff_A_T6DH3wwq8_1;
	wire w_dff_A_KrLgufYI9_2;
	wire w_dff_A_mb2OTymV4_2;
	wire w_dff_A_SLcNwMxy7_0;
	wire w_dff_A_lC4qb3jX0_0;
	wire w_dff_A_lZXB9Ylo4_0;
	wire w_dff_B_9jMRwUAO9_2;
	wire w_dff_B_kPkQ15z64_2;
	wire w_dff_B_kKtfS4rA8_2;
	wire w_dff_A_jX290eNI2_0;
	wire w_dff_A_s8xnPzOq5_1;
	wire w_dff_A_SxvGIu5g6_1;
	wire w_dff_B_W9vLfPdA9_3;
	wire w_dff_B_uwGCQ1Gp5_3;
	wire w_dff_B_RgcyJSHo2_3;
	wire w_dff_B_bzl0gWHi7_3;
	wire w_dff_B_yRq3ZuRu6_3;
	wire w_dff_B_zJt5tn4C4_3;
	wire w_dff_B_baY7IJcr3_3;
	wire w_dff_B_GA7pTdUZ8_3;
	wire w_dff_B_T8FdJU7K8_3;
	wire w_dff_B_5RF7sKrM0_3;
	wire w_dff_B_ldnKndYB2_3;
	wire w_dff_A_F0MUBJYi3_0;
	wire w_dff_A_WzpvETxh7_0;
	wire w_dff_A_NvDLcwJC7_0;
	wire w_dff_A_6afAvTiA1_0;
	wire w_dff_A_AWdn3BLB4_0;
	wire w_dff_A_Avu9ZOkc3_0;
	wire w_dff_A_0begA1fN1_0;
	wire w_dff_A_ffGYkaM04_0;
	wire w_dff_A_R7Bcrq286_0;
	wire w_dff_A_QsS64q9h6_0;
	wire w_dff_A_N02OklIP5_0;
	wire w_dff_A_zFcb95415_0;
	wire w_dff_A_D0l4WvQv4_0;
	wire w_dff_A_ehAwgVB08_0;
	wire w_dff_A_yBL0tugy4_2;
	wire w_dff_A_gm1J99Qc7_2;
	wire w_dff_A_HXkUXqia7_2;
	wire w_dff_A_rFBNmaJz8_2;
	wire w_dff_A_M7wVrncw9_2;
	wire w_dff_A_G0fSlt6T2_1;
	wire w_dff_A_bXAyjwwu1_1;
	wire w_dff_A_Fw08xDqB0_1;
	wire w_dff_A_ehkbIuDh9_1;
	wire w_dff_A_pSxPcOGY3_1;
	wire w_dff_A_XCpN15Zn1_2;
	wire w_dff_A_3jDpRkMg1_2;
	wire w_dff_A_MmY3BLUr3_2;
	wire w_dff_A_uHvhsYT62_2;
	wire w_dff_A_geXDWWpj9_2;
	wire w_dff_A_2cAierZb3_2;
	wire w_dff_A_Jg55DGE26_2;
	wire w_dff_A_lQlJXt8t3_2;
	wire w_dff_A_RiQyqCRg9_2;
	wire w_dff_A_hphdq8121_2;
	wire w_dff_A_qtSG9lwf5_2;
	wire w_dff_A_XLa1vGuz1_2;
	wire w_dff_A_1RvgfV2T7_2;
	wire w_dff_B_cI4nzNZ88_0;
	wire w_dff_B_L2qPwmGX6_0;
	wire w_dff_B_9P2eLogb0_1;
	wire w_dff_B_GtBINyod8_1;
	wire w_dff_B_FekjwbPH0_0;
	wire w_dff_A_yC57tngl3_0;
	wire w_dff_A_oEs2wZ5J3_0;
	wire w_dff_A_zXTFClyW9_1;
	wire w_dff_A_ekkaAfHZ3_1;
	wire w_dff_A_MNZ06QkH1_2;
	wire w_dff_A_LqdujMuD7_2;
	wire w_dff_A_qWObL3q60_1;
	wire w_dff_A_EC2x0mWa3_1;
	wire w_dff_A_xWPT1tlm4_1;
	wire w_dff_A_WmoD18nh9_1;
	wire w_dff_A_UpOGuhrs6_1;
	wire w_dff_A_OtXKASWw2_1;
	wire w_dff_A_0OPGAQxC3_1;
	wire w_dff_A_Ym2u3F2I1_1;
	wire w_dff_A_QJDwRvtH6_1;
	wire w_dff_B_txm5M3Xs0_2;
	wire w_dff_B_TNGCVpEa1_2;
	wire w_dff_A_wLnESNMi5_1;
	wire w_dff_A_f82UZDuO2_1;
	wire w_dff_B_0P5kGAq49_2;
	wire w_dff_B_n6OpHj769_2;
	wire w_dff_B_wfvo8goK1_1;
	wire w_dff_B_s7RfLXDr5_0;
	wire w_dff_A_SUobC3IH6_1;
	wire w_dff_A_DlWciL399_1;
	wire w_dff_A_v7RoWmpE5_1;
	wire w_dff_A_h7Gae4JC6_1;
	wire w_dff_A_T2l5DZtf0_1;
	wire w_dff_A_ZWMNnxvV5_2;
	wire w_dff_A_vKGARMXT5_2;
	wire w_dff_A_51wQeFao0_2;
	wire w_dff_A_erKoI9zu3_2;
	wire w_dff_A_27MsNwcw0_2;
	wire w_dff_A_8FAGhlia4_2;
	wire w_dff_A_9C1hqSRx7_2;
	wire w_dff_A_GbsbaBAM0_2;
	wire w_dff_A_6BvlZLHM4_2;
	wire w_dff_A_3WkyXO8q5_2;
	wire w_dff_A_D6zaqLRz9_2;
	wire w_dff_A_9nPoXgzs7_2;
	wire w_dff_B_8cvNMGpq8_1;
	wire w_dff_B_M6rCd2HD1_0;
	wire w_dff_A_mz1xwCoR0_0;
	wire w_dff_A_Tr8DNePw2_0;
	wire w_dff_A_W2sQknpv5_2;
	wire w_dff_A_fwUXfxUZ0_2;
	wire w_dff_A_DJ3DCg119_1;
	wire w_dff_A_10wQNGWj8_1;
	wire w_dff_A_q9efD5AW6_1;
	wire w_dff_A_grsjDkSy3_1;
	wire w_dff_A_CpakcBnU6_1;
	wire w_dff_A_4WvY5A2k1_1;
	wire w_dff_A_2PIS5woK2_1;
	wire w_dff_A_vwftn3eC3_1;
	wire w_dff_A_3dPNGlx54_1;
	wire w_dff_A_z9Is80aF2_1;
	wire w_dff_A_vMJgKACb1_1;
	wire w_dff_A_cQUJLcfI9_1;
	wire w_dff_A_dju4lfQv3_1;
	wire w_dff_B_a2pNsB9Y1_1;
	wire w_dff_B_7QV1unCt1_0;
	wire w_dff_A_bNwzzcrN2_2;
	wire w_dff_A_C8AfzeSp8_2;
	wire w_dff_A_kepke5qS6_2;
	wire w_dff_A_d6USlwJ36_2;
	wire w_dff_A_DB2Wrj6J1_1;
	wire w_dff_A_Olvsr9NF6_1;
	wire w_dff_A_RWSabYOR2_1;
	wire w_dff_A_0St775YA1_1;
	wire w_dff_A_IM7OfCDf7_1;
	wire w_dff_A_AaWoBz0U8_1;
	wire w_dff_A_eRNhunRI9_1;
	wire w_dff_A_4qWlNzCh6_1;
	wire w_dff_A_qjV563ti3_1;
	wire w_dff_A_0FiDF4Wn0_1;
	wire w_dff_B_50ilp20S7_2;
	wire w_dff_B_xjUMoG9V3_1;
	wire w_dff_B_fE0qDrAB4_0;
	wire w_dff_A_lQ3831J44_1;
	wire w_dff_A_JBmjHym93_1;
	wire w_dff_A_97Q6vCgf6_2;
	wire w_dff_A_lw13vdjv0_2;
	wire w_dff_A_m6ftOYds0_1;
	wire w_dff_A_FTlmgWLO4_1;
	wire w_dff_A_udDzy56d3_1;
	wire w_dff_A_5JKO9HUY8_1;
	wire w_dff_B_L7ehRztw8_1;
	wire w_dff_B_P7u6YAzT2_1;
	wire w_dff_B_NtNfFnlQ6_1;
	wire w_dff_B_FWwsQ1OX3_1;
	wire w_dff_B_7GV5nmRp3_1;
	wire w_dff_B_APXEe3xc8_1;
	wire w_dff_B_bb6ohPrX4_1;
	wire w_dff_B_0ty9xCX39_1;
	wire w_dff_B_C1fNn5vN1_1;
	wire w_dff_B_PyqZRoxv3_1;
	wire w_dff_B_8ReLGgYj4_1;
	wire w_dff_B_Dn49nIRW9_1;
	wire w_dff_B_sYlCGmio9_1;
	wire w_dff_A_tVHP3ub39_1;
	wire w_dff_A_We4CQKko3_1;
	wire w_dff_A_OLYZPrwD4_1;
	wire w_dff_A_2MoRzi234_1;
	wire w_dff_A_pjFj03hC5_1;
	wire w_dff_A_i2BNmNkV7_1;
	wire w_dff_A_rkCiUCNi9_1;
	wire w_dff_A_jmIQUttQ0_1;
	wire w_dff_A_VAADDw1t6_1;
	wire w_dff_A_4ffNxxmu7_1;
	wire w_dff_A_o6MVf1uf5_1;
	wire w_dff_A_uPsZQYsd5_1;
	wire w_dff_A_wxbAMaeY6_2;
	wire w_dff_A_u55ca3qf7_2;
	wire w_dff_A_4V5MLa2f1_2;
	wire w_dff_A_RzDvUsnI8_2;
	wire w_dff_A_wFuCSSMj3_0;
	wire w_dff_A_1fbhWlmc2_0;
	wire w_dff_A_HIs4Qe9V0_0;
	wire w_dff_A_QcjPCR3s1_0;
	wire w_dff_A_eytVzZhE5_0;
	wire w_dff_A_TnK07E4D0_0;
	wire w_dff_A_Dnw5UdAG5_0;
	wire w_dff_A_l9F1dX233_0;
	wire w_dff_A_CQBBE4km1_0;
	wire w_dff_A_aUNklMmy4_1;
	wire w_dff_A_mnGL5ekG2_1;
	wire w_dff_A_a31CDdwQ9_1;
	wire w_dff_A_tYeMHNTp3_1;
	wire w_dff_A_wdpgfduw9_1;
	wire w_dff_A_dijHIl8Y2_1;
	wire w_dff_A_u7CR8iOw3_1;
	wire w_dff_A_HwbULfST9_0;
	wire w_dff_B_rBPl433c7_2;
	wire w_dff_B_IL6LlgCz6_2;
	wire w_dff_A_QSMjHyq86_1;
	wire w_dff_A_R5PM2Q5y9_1;
	wire w_dff_A_G23F854o3_1;
	wire w_dff_A_2MAJkVPS5_1;
	wire w_dff_A_rNwQE5Az1_1;
	wire w_dff_B_iivay0ji0_3;
	wire w_dff_A_TcgSIRFV1_0;
	wire w_dff_A_8kUJOeFo4_0;
	wire w_dff_A_EVwhCroP0_0;
	wire w_dff_A_0ekPl5pE5_0;
	wire w_dff_A_pk4VvjxV7_2;
	wire w_dff_A_8VRlv9Ky3_2;
	wire w_dff_A_JJz8ZuTB3_2;
	wire w_dff_A_lEOyIBCx6_2;
	wire w_dff_A_JeMr8D3h9_2;
	wire w_dff_A_BtE9KoFR5_2;
	wire w_dff_A_GIscOO4y1_0;
	wire w_dff_A_AA1GIeGo7_0;
	wire w_dff_A_6OPMGmh60_0;
	wire w_dff_B_oEDRfFsY6_3;
	wire w_dff_A_lQtzHlbT7_0;
	wire w_dff_A_8gH7ZCXd4_1;
	wire w_dff_A_abmFYAEM6_0;
	wire w_dff_A_OUvp96IM3_1;
	wire w_dff_A_hfbqRdsU0_1;
	wire w_dff_A_4yJLPBI18_1;
	wire w_dff_A_fMw4awqK4_1;
	wire w_dff_A_G5JbCDNA5_2;
	wire w_dff_A_qhiPFY6g6_2;
	wire w_dff_B_1i2SLdk65_1;
	wire w_dff_B_ELLLUtH34_0;
	wire w_dff_A_jCHUc5Ti2_1;
	wire w_dff_A_k5oACphD2_0;
	wire w_dff_A_xecZ0YzB1_0;
	wire w_dff_A_FIyIO9se7_2;
	wire w_dff_A_XWBOdunm4_2;
	wire w_dff_A_uabqrrnq4_1;
	wire w_dff_A_nAghyw0R2_1;
	wire w_dff_A_v1DPICNN5_1;
	wire w_dff_A_EBj3uFbd5_1;
	wire w_dff_A_726Qwzzu5_1;
	wire w_dff_A_4jEPWjE13_1;
	wire w_dff_A_WZmF5jrl7_1;
	wire w_dff_A_ZCmzAjkn2_2;
	wire w_dff_A_1wCTM7hN2_2;
	wire w_dff_A_LKOjZSAq4_2;
	wire w_dff_B_pxBIfhne4_1;
	wire w_dff_B_q1q8bvml7_0;
	wire w_dff_A_byP7oCMA1_1;
	wire w_dff_A_3QSoSmmK1_1;
	wire w_dff_A_VAhCKBDb7_2;
	wire w_dff_A_MQZwyx2v6_2;
	wire w_dff_A_rw8FVwEy8_1;
	wire w_dff_A_AhzntgmX8_1;
	wire w_dff_A_HOmbI2og8_1;
	wire w_dff_A_ky1Zb9sY5_1;
	wire w_dff_A_Ifwq6ZIh7_0;
	wire w_dff_A_NutrcOz82_0;
	wire w_dff_A_eVsK6hWb2_0;
	wire w_dff_A_XDICiVpS9_0;
	wire w_dff_A_RoLXqBJa7_0;
	wire w_dff_A_ZnXxb8QY4_0;
	wire w_dff_A_kpVQThfN9_0;
	wire w_dff_A_r2JoQ3I74_0;
	wire w_dff_A_lEWmyDbc0_0;
	wire w_dff_A_pumRDhR26_1;
	wire w_dff_A_KfabqNKi2_1;
	wire w_dff_A_sWU4GC0H7_1;
	wire w_dff_A_ZNiXlFuF1_1;
	wire w_dff_B_9E1ofxPW9_1;
	wire w_dff_B_xFCehTzh4_0;
	wire w_dff_A_9oWdtRfv0_2;
	wire w_dff_A_ghbSHbT54_1;
	wire w_dff_A_6JY6j7Qz2_1;
	wire w_dff_A_nFnDtmKI9_2;
	wire w_dff_A_f2nqb3SF5_2;
	wire w_dff_A_cxdFok9Y7_1;
	wire w_dff_A_K1Y39WDO9_1;
	wire w_dff_A_1mrJC09w4_1;
	wire w_dff_A_EXeMCmjT5_1;
	wire w_dff_A_22M6stkl3_1;
	wire w_dff_A_S4BFoTEg6_0;
	wire w_dff_A_cUjB2sxD9_0;
	wire w_dff_A_2FGcljJN8_0;
	wire w_dff_A_Q0WvdquK7_0;
	wire w_dff_A_WgqfywFy7_0;
	wire w_dff_A_ooOM0ng85_0;
	wire w_dff_A_iG3EWeGa5_0;
	wire w_dff_A_jshj2HiV8_0;
	wire w_dff_A_tW6X4tx01_0;
	wire w_dff_A_J9C4wcfI8_0;
	wire w_dff_A_qysSZoJr1_0;
	wire w_dff_A_yU5Vka497_0;
	wire w_dff_A_Ph4Tfi194_0;
	wire w_dff_A_5QfYp62S4_0;
	wire w_dff_A_l4sKdUgq2_0;
	wire w_dff_A_9kWW4kCv6_0;
	wire w_dff_A_8ALYuyfL6_0;
	wire w_dff_A_FAb7LJJY5_0;
	wire w_dff_A_Fv2hj1QM1_0;
	wire w_dff_A_XKd3H5AC1_0;
	wire w_dff_A_o5d3wDgu8_0;
	wire w_dff_A_zeVGAt1I0_0;
	wire w_dff_A_eXbbmxP21_0;
	wire w_dff_A_RmA6BJyc6_0;
	wire w_dff_A_hMn7lFQn0_0;
	wire w_dff_A_oaFdoqsV7_0;
	wire w_dff_A_LUm5Lnf42_0;
	wire w_dff_A_hXiG1aqj1_0;
	wire w_dff_A_amNfyYye3_0;
	wire w_dff_A_dySuGVcc0_0;
	wire w_dff_A_ESk33UDh2_0;
	wire w_dff_A_HBJBjulU5_0;
	wire w_dff_A_wKp5vQlJ0_0;
	wire w_dff_A_TYsgP5zn3_0;
	wire w_dff_A_J41lkMAy3_0;
	wire w_dff_A_PgBZ7IZV6_0;
	wire w_dff_A_aowgxbNX0_0;
	wire w_dff_A_HVDuQ0YC1_0;
	wire w_dff_A_FXX2zFPh3_1;
	wire w_dff_A_kb1Jqb6t5_0;
	wire w_dff_A_ESnj91XR7_0;
	wire w_dff_A_uP4QCxyX4_0;
	wire w_dff_A_96M8kcMJ0_0;
	wire w_dff_A_GVrsSbyC8_0;
	wire w_dff_A_Yvn67Gvx1_0;
	wire w_dff_A_WAnU2WVe6_0;
	wire w_dff_A_Ak3wK5Nx7_0;
	wire w_dff_A_wdjaViia8_0;
	wire w_dff_A_YdebARPe6_0;
	wire w_dff_A_Ca4iiYRE3_0;
	wire w_dff_A_2bRzvp8s6_0;
	wire w_dff_A_tDHIY1q45_0;
	wire w_dff_A_Tki5cdCZ2_0;
	wire w_dff_A_8wxorWK81_0;
	wire w_dff_A_BkjYdNYj3_0;
	wire w_dff_A_8VhYLVrL6_0;
	wire w_dff_A_pYU1CmHc1_0;
	wire w_dff_A_GWI359iE7_0;
	wire w_dff_A_1x7sEI0E9_0;
	wire w_dff_A_FuxWOYa01_0;
	wire w_dff_A_bRszjOR23_0;
	wire w_dff_A_bRuHXpf80_0;
	wire w_dff_A_KpBloNhI2_0;
	wire w_dff_A_7PtS6bqi0_0;
	wire w_dff_A_7t5sQ2k68_0;
	wire w_dff_A_ErKWJn080_0;
	wire w_dff_A_WgoReFDp1_0;
	wire w_dff_A_qS46TXoT6_0;
	wire w_dff_A_gdDr2Rt98_0;
	wire w_dff_A_Z8a0uKeH2_0;
	wire w_dff_A_dKOU73DZ5_0;
	wire w_dff_A_S0bU80Qj9_0;
	wire w_dff_A_0ouWjXHq3_0;
	wire w_dff_A_2asVuN543_0;
	wire w_dff_A_VzLzMeMV6_0;
	wire w_dff_A_pN6dqDnS3_0;
	wire w_dff_A_2rLl3HX90_0;
	wire w_dff_A_APRPgR7j9_1;
	wire w_dff_A_joyYYdNZ9_0;
	wire w_dff_A_Jf93922w9_0;
	wire w_dff_A_Gr38YLUF1_0;
	wire w_dff_A_7f7gfzmx5_0;
	wire w_dff_A_9e0u9XDq2_0;
	wire w_dff_A_jxaGMBcM1_0;
	wire w_dff_A_A4CM5ywT6_0;
	wire w_dff_A_PeUX5KYj9_0;
	wire w_dff_A_1SIO7G3m7_0;
	wire w_dff_A_vseIl3hp2_0;
	wire w_dff_A_cJ6w0haZ7_0;
	wire w_dff_A_NJQndC2a4_0;
	wire w_dff_A_TGfx6qn55_0;
	wire w_dff_A_lhQJjV5B4_0;
	wire w_dff_A_t1E4pHzx1_0;
	wire w_dff_A_GCmU1yjW9_0;
	wire w_dff_A_4ePGndEy2_0;
	wire w_dff_A_deH99ELa8_0;
	wire w_dff_A_EhrpGzo54_0;
	wire w_dff_A_Pb2Rtkhx1_0;
	wire w_dff_A_hikMJNge3_0;
	wire w_dff_A_ReDCaeiz6_0;
	wire w_dff_A_rPRVe1h62_0;
	wire w_dff_A_4zA1Yrov6_0;
	wire w_dff_A_7SFxjS3U8_0;
	wire w_dff_A_atmgDZ0b6_0;
	wire w_dff_A_E5BsM33q3_0;
	wire w_dff_A_jEDbpPey0_0;
	wire w_dff_A_LHPxXMxu9_0;
	wire w_dff_A_HFeGHG6V1_0;
	wire w_dff_A_9ymznQRo8_0;
	wire w_dff_A_VOfRLEwm1_0;
	wire w_dff_A_FsAWgeSX1_0;
	wire w_dff_A_ruaAMZbA3_0;
	wire w_dff_A_yy8WFVP23_0;
	wire w_dff_A_GLO2zFsA6_0;
	wire w_dff_A_2DVGfjUz6_0;
	wire w_dff_A_Kpoxo9Ac0_0;
	wire w_dff_A_NJEEXzqd5_1;
	wire w_dff_A_pLDhAxMW8_0;
	wire w_dff_A_HrgcHspM1_0;
	wire w_dff_A_vItZSYUu0_0;
	wire w_dff_A_C2s8FxDV2_0;
	wire w_dff_A_50huoxlO8_0;
	wire w_dff_A_ymn8d7Ed9_0;
	wire w_dff_A_N2s6VMqI2_0;
	wire w_dff_A_4x2ySOQx5_0;
	wire w_dff_A_rJQDC5Ul8_0;
	wire w_dff_A_lzE6P0r60_0;
	wire w_dff_A_Kvpt5Jz93_0;
	wire w_dff_A_rR3p43uK6_0;
	wire w_dff_A_qvSXeoiA3_0;
	wire w_dff_A_EpUsK3Ox6_0;
	wire w_dff_A_qIxks7bg9_0;
	wire w_dff_A_hw0WMDrl4_0;
	wire w_dff_A_JMjM0Poi2_0;
	wire w_dff_A_1oOQQzJq1_0;
	wire w_dff_A_YYIfwsKE6_0;
	wire w_dff_A_7cCxsnQj9_0;
	wire w_dff_A_V0sMGLOD2_0;
	wire w_dff_A_JZ9MfmNk1_0;
	wire w_dff_A_bLjutzPT2_0;
	wire w_dff_A_19OpLNiN2_0;
	wire w_dff_A_ozZ9DEEF6_0;
	wire w_dff_A_Nrvh4t3X0_0;
	wire w_dff_A_psu5GN3F5_0;
	wire w_dff_A_BMjsK2cp1_0;
	wire w_dff_A_hFHxa1pX2_0;
	wire w_dff_A_swjjkuwg7_0;
	wire w_dff_A_DPx1y6bV7_0;
	wire w_dff_A_2gyv21uI6_0;
	wire w_dff_A_TK11w9Mu1_0;
	wire w_dff_A_UsPHTIis6_0;
	wire w_dff_A_ePDkRL1W0_0;
	wire w_dff_A_mM7rX9mh2_0;
	wire w_dff_A_lMMfu7Xz6_0;
	wire w_dff_A_iLl64GnQ8_0;
	wire w_dff_A_pjeMTmIZ9_1;
	wire w_dff_A_5VHOhAeF2_0;
	wire w_dff_A_U9QzQQ9X1_0;
	wire w_dff_A_VQFCUgMN2_0;
	wire w_dff_A_zIT6kIx26_0;
	wire w_dff_A_XMBCQbZP8_0;
	wire w_dff_A_cr8nApi83_0;
	wire w_dff_A_HUnZAv1t8_0;
	wire w_dff_A_DS8rsTnH4_0;
	wire w_dff_A_RUxLkkNd4_0;
	wire w_dff_A_De5hgCDX4_0;
	wire w_dff_A_VPO65Toq8_0;
	wire w_dff_A_KpwmRhmd8_0;
	wire w_dff_A_HZKXD9XM7_0;
	wire w_dff_A_UpxB5qYb2_0;
	wire w_dff_A_hbYWN6iI1_0;
	wire w_dff_A_sulSAXgm5_0;
	wire w_dff_A_TFdCJt3D0_0;
	wire w_dff_A_aD0Xtqq53_0;
	wire w_dff_A_qXy8SuO81_0;
	wire w_dff_A_N3PHSIqS1_0;
	wire w_dff_A_sqfIr7R24_0;
	wire w_dff_A_0fVAjGjA0_0;
	wire w_dff_A_GE8rLY793_0;
	wire w_dff_A_NtiNDVCG5_0;
	wire w_dff_A_7xeFGeCz4_0;
	wire w_dff_A_eGcgMxIJ4_0;
	wire w_dff_A_C5PEqtWi0_0;
	wire w_dff_A_rxe9sFe13_0;
	wire w_dff_A_XNvkBDgL3_0;
	wire w_dff_A_IJNGve9L7_0;
	wire w_dff_A_Nsd9QtNA2_0;
	wire w_dff_A_YaqgMtqt4_0;
	wire w_dff_A_ieI7m9dX1_0;
	wire w_dff_A_YHyu4QRf7_0;
	wire w_dff_A_Rp9Mh0v21_0;
	wire w_dff_A_tc341b1e3_0;
	wire w_dff_A_H0i7A5Jk0_0;
	wire w_dff_A_R6NsU4lJ8_0;
	wire w_dff_A_wpKXgQFK7_1;
	wire w_dff_A_NRfkR5Rg5_0;
	wire w_dff_A_aSrchFsx3_0;
	wire w_dff_A_1uZ6WErQ9_0;
	wire w_dff_A_T7iW3xuc1_0;
	wire w_dff_A_MooRyZOh2_0;
	wire w_dff_A_w5D30tJ44_0;
	wire w_dff_A_YJxLTvYM8_0;
	wire w_dff_A_rSipwpsY5_0;
	wire w_dff_A_ZBXtti1C9_0;
	wire w_dff_A_MVqZHUEl9_0;
	wire w_dff_A_yI3eLD4U0_0;
	wire w_dff_A_S25IkXfV5_0;
	wire w_dff_A_r3ahwtRx7_0;
	wire w_dff_A_VsEkdvk80_0;
	wire w_dff_A_BRkNOJsf7_0;
	wire w_dff_A_iiKzEKlV2_0;
	wire w_dff_A_k9Irk9G35_0;
	wire w_dff_A_jOe8RLtg7_0;
	wire w_dff_A_V3hm9Lmh5_0;
	wire w_dff_A_X8aFoeJu3_0;
	wire w_dff_A_X9wJXq9V7_0;
	wire w_dff_A_9oMvkVNg9_0;
	wire w_dff_A_2weA3CNg6_0;
	wire w_dff_A_9vnvz8Io1_0;
	wire w_dff_A_oCtwRTgz3_0;
	wire w_dff_A_jG079AtQ9_0;
	wire w_dff_A_LGRfUNvg7_0;
	wire w_dff_A_S2o33HEF5_0;
	wire w_dff_A_0vdKzqsL4_0;
	wire w_dff_A_UtkowifO0_0;
	wire w_dff_A_8QSAcOa86_0;
	wire w_dff_A_YMEXzMq00_0;
	wire w_dff_A_uHVHlb2t0_0;
	wire w_dff_A_dxfDkiid8_0;
	wire w_dff_A_WRg3cFNA0_0;
	wire w_dff_A_mv9TeVLQ0_0;
	wire w_dff_A_N4kyoXmk4_0;
	wire w_dff_A_T5ewH2rZ8_0;
	wire w_dff_A_anzn7UR03_1;
	wire w_dff_A_v6uTtzOE0_0;
	wire w_dff_A_2eVirea68_0;
	wire w_dff_A_OlmaOuYn5_0;
	wire w_dff_A_adIBZ9nD8_0;
	wire w_dff_A_a8gVUd2g9_0;
	wire w_dff_A_39vzzhvZ8_0;
	wire w_dff_A_EQM940HP3_0;
	wire w_dff_A_FlIdlKtr1_0;
	wire w_dff_A_Ecx36kOV9_0;
	wire w_dff_A_2ENfJecH1_0;
	wire w_dff_A_l6Op9T8j6_0;
	wire w_dff_A_gZOGycUB6_0;
	wire w_dff_A_wClD1ypr4_0;
	wire w_dff_A_FxuEfVco8_0;
	wire w_dff_A_oJZOEiA06_0;
	wire w_dff_A_HBxp9Q4m2_0;
	wire w_dff_A_FKBI3KL28_0;
	wire w_dff_A_uYj6YSfL4_0;
	wire w_dff_A_QfirL6wC1_0;
	wire w_dff_A_pibm4Z2y9_0;
	wire w_dff_A_DLSmdPvn1_0;
	wire w_dff_A_0BWT3AG56_0;
	wire w_dff_A_gd1pvYuj4_0;
	wire w_dff_A_UDJaqCAE2_0;
	wire w_dff_A_tW2S6lpC2_0;
	wire w_dff_A_bGAxGVPH0_0;
	wire w_dff_A_3MM7oVWi2_0;
	wire w_dff_A_fF2TI0ro4_0;
	wire w_dff_A_1kksXPnv6_0;
	wire w_dff_A_2N90lZmI6_0;
	wire w_dff_A_6CPn6VuH5_0;
	wire w_dff_A_oKpCBGvs8_0;
	wire w_dff_A_prIP4twm0_0;
	wire w_dff_A_hXNc79B47_0;
	wire w_dff_A_mMTCwnvF9_0;
	wire w_dff_A_zRJ58SpW8_0;
	wire w_dff_A_emxznUEz5_0;
	wire w_dff_A_w4IbDKxW6_0;
	wire w_dff_A_SmHHSwBU9_1;
	wire w_dff_A_IllnQw2i3_0;
	wire w_dff_A_MoIg7aE97_0;
	wire w_dff_A_RTuxeuop9_0;
	wire w_dff_A_cs9yoYxh6_0;
	wire w_dff_A_9vD9Msxf3_0;
	wire w_dff_A_YE8pMHkq1_0;
	wire w_dff_A_vmCRhtlb3_0;
	wire w_dff_A_bksCjaE00_0;
	wire w_dff_A_8XGRIX9H7_0;
	wire w_dff_A_aDQZd3382_0;
	wire w_dff_A_8Y9VSXqN9_0;
	wire w_dff_A_fO4se0o44_0;
	wire w_dff_A_tR5P0jYG9_0;
	wire w_dff_A_B1PheY4K2_0;
	wire w_dff_A_O1scLa9C1_0;
	wire w_dff_A_I7VUaWfu0_0;
	wire w_dff_A_X8IZP3vW9_0;
	wire w_dff_A_pmSQrNhR3_0;
	wire w_dff_A_zTi8jiHI0_0;
	wire w_dff_A_GnmzxZgJ0_0;
	wire w_dff_A_Wfdp2Woa9_0;
	wire w_dff_A_NiBiFuvV6_0;
	wire w_dff_A_GBKZmWoa2_0;
	wire w_dff_A_9RgFqwdU7_0;
	wire w_dff_A_kMmQEkZV6_0;
	wire w_dff_A_IfwIk9Mo6_0;
	wire w_dff_A_qFwxWb6H9_0;
	wire w_dff_A_9T4GLeUL7_0;
	wire w_dff_A_pnPsdKjh3_0;
	wire w_dff_A_7IIicVW07_0;
	wire w_dff_A_KQoFEcxO5_0;
	wire w_dff_A_vx3J51w74_0;
	wire w_dff_A_XJDpRknC7_0;
	wire w_dff_A_AdZ9fheF7_0;
	wire w_dff_A_5KNDTQtG6_0;
	wire w_dff_A_id4zQhtR6_0;
	wire w_dff_A_0YQTmjmN1_0;
	wire w_dff_A_OSb0Z9x99_0;
	wire w_dff_A_80xgeO6u2_1;
	wire w_dff_A_ezgQ9NYB2_0;
	wire w_dff_A_biwJmZpO0_0;
	wire w_dff_A_JkUfybyo6_0;
	wire w_dff_A_v58gaw6T7_0;
	wire w_dff_A_bzeXVAKH7_0;
	wire w_dff_A_z3P9eGGF9_0;
	wire w_dff_A_APjyFnb33_0;
	wire w_dff_A_YWuP8LU71_0;
	wire w_dff_A_5dRQYwzG2_0;
	wire w_dff_A_0llwhG3y7_0;
	wire w_dff_A_FYuuIKS63_0;
	wire w_dff_A_6dW1B7MK5_0;
	wire w_dff_A_nOmjzmaC0_0;
	wire w_dff_A_8plihuOL8_0;
	wire w_dff_A_LNIor2Xf0_0;
	wire w_dff_A_CEBDPqtw5_0;
	wire w_dff_A_16OuaOQH2_0;
	wire w_dff_A_AVimHYPv4_0;
	wire w_dff_A_vvESrzoA1_0;
	wire w_dff_A_yATOE5Va9_0;
	wire w_dff_A_EcludsJw6_0;
	wire w_dff_A_pY3RRJxD2_0;
	wire w_dff_A_WFNoR3kn7_0;
	wire w_dff_A_MHpEk0p79_0;
	wire w_dff_A_WOmtw4fb2_0;
	wire w_dff_A_ZmMtlInh1_0;
	wire w_dff_A_RHUMRomJ5_0;
	wire w_dff_A_dJNh6HjZ3_0;
	wire w_dff_A_RbrVPB010_0;
	wire w_dff_A_g0nl9VDs2_0;
	wire w_dff_A_9IjAxkMp3_0;
	wire w_dff_A_SuYkeoy75_0;
	wire w_dff_A_pxcwxjmd6_0;
	wire w_dff_A_ec3ctuvZ9_0;
	wire w_dff_A_Tf1nq2nt0_0;
	wire w_dff_A_cRrTHZtY5_0;
	wire w_dff_A_mxSh4hRX4_0;
	wire w_dff_A_8yyeYsUc3_0;
	wire w_dff_A_YVg7X2Az1_1;
	wire w_dff_A_MXaWD79m3_0;
	wire w_dff_A_jLdr1f5V8_0;
	wire w_dff_A_UFyh85405_0;
	wire w_dff_A_p1eiRlI63_0;
	wire w_dff_A_FNKxDVsY5_0;
	wire w_dff_A_GpjnpPWB6_0;
	wire w_dff_A_WRkQc04j3_0;
	wire w_dff_A_t4dCEtDO0_0;
	wire w_dff_A_GbRewRmk2_0;
	wire w_dff_A_AO0R8pZt7_0;
	wire w_dff_A_Sd5Okzlu6_0;
	wire w_dff_A_utuPAZp03_0;
	wire w_dff_A_i314Kx4Z4_0;
	wire w_dff_A_8cMlb01G5_0;
	wire w_dff_A_aeMYdjSe5_0;
	wire w_dff_A_VYRWkyGi3_0;
	wire w_dff_A_CiJDJtQR6_0;
	wire w_dff_A_KW1APJHx1_0;
	wire w_dff_A_8FTIaBrG0_0;
	wire w_dff_A_cEPE2HEn9_0;
	wire w_dff_A_fGni8lWD1_0;
	wire w_dff_A_UXajtxwi9_0;
	wire w_dff_A_AOieRl762_0;
	wire w_dff_A_e9d9JLwp0_0;
	wire w_dff_A_gQNRETQP8_0;
	wire w_dff_A_1IKU9MDR5_0;
	wire w_dff_A_YtYnKT9c6_0;
	wire w_dff_A_lhyrcOQn2_0;
	wire w_dff_A_xUhD7t390_0;
	wire w_dff_A_nkJ6LJve5_0;
	wire w_dff_A_xznqdVAg2_0;
	wire w_dff_A_SCLFNjAf3_0;
	wire w_dff_A_lmcW9Wyn7_0;
	wire w_dff_A_vlXgyy7X4_0;
	wire w_dff_A_lKgm11G57_0;
	wire w_dff_A_4uC7qwO28_0;
	wire w_dff_A_JYBOTeNq5_0;
	wire w_dff_A_cRtgBYsu5_0;
	wire w_dff_A_mpaoxbKU2_1;
	wire w_dff_A_cYZ2IKGn7_0;
	wire w_dff_A_cycveu3Z7_0;
	wire w_dff_A_CIoCGSL70_0;
	wire w_dff_A_J2ionYCO1_0;
	wire w_dff_A_K2yjXhet7_0;
	wire w_dff_A_anAyCNaC6_0;
	wire w_dff_A_zJlDiPSJ3_0;
	wire w_dff_A_g9kp4wvI9_0;
	wire w_dff_A_omvzH8zG3_0;
	wire w_dff_A_ccqN55Ia5_0;
	wire w_dff_A_6gbjhOCs0_0;
	wire w_dff_A_4MBoiJ1d1_0;
	wire w_dff_A_O8VjdEiG0_0;
	wire w_dff_A_xioW0aD39_0;
	wire w_dff_A_1CvV8QTk9_0;
	wire w_dff_A_tR8aNwGo7_0;
	wire w_dff_A_nBYRpbld3_0;
	wire w_dff_A_kvRiJ8q16_0;
	wire w_dff_A_qWhhbW5h1_0;
	wire w_dff_A_dfq6BZrT7_0;
	wire w_dff_A_VyTe9x7Q3_0;
	wire w_dff_A_vJ6wse6q6_0;
	wire w_dff_A_XbiUDmNj9_0;
	wire w_dff_A_r2vlyFyq6_0;
	wire w_dff_A_uPjsHCum6_0;
	wire w_dff_A_KJTLbru53_0;
	wire w_dff_A_bfFVPh7U2_0;
	wire w_dff_A_g2brIlxC0_0;
	wire w_dff_A_nCLp73rZ4_0;
	wire w_dff_A_5XSOq4r64_0;
	wire w_dff_A_j5H86hvk2_0;
	wire w_dff_A_m4SKr0up3_0;
	wire w_dff_A_4Eq57y9q2_0;
	wire w_dff_A_TNHctidh2_0;
	wire w_dff_A_YOpylAWh6_0;
	wire w_dff_A_X8mRE8At2_0;
	wire w_dff_A_TFZIlna89_0;
	wire w_dff_A_NG80fwJf3_0;
	wire w_dff_A_gICE3Ix18_1;
	wire w_dff_A_hAy73yhW6_0;
	wire w_dff_A_mIioMXJ75_0;
	wire w_dff_A_OkALlnOw5_0;
	wire w_dff_A_UhZFbW2Y2_0;
	wire w_dff_A_JS6anSuB8_0;
	wire w_dff_A_bhDUjaVG7_0;
	wire w_dff_A_qk8ezBHH1_0;
	wire w_dff_A_jftG65BW3_0;
	wire w_dff_A_W60Ja46K7_0;
	wire w_dff_A_aRka5JIz5_0;
	wire w_dff_A_jlLkGC4H5_0;
	wire w_dff_A_RkGwdNfh5_0;
	wire w_dff_A_XvFD3BqM1_0;
	wire w_dff_A_NgdQUWgm4_0;
	wire w_dff_A_gMMartza4_0;
	wire w_dff_A_3NpBXOue6_0;
	wire w_dff_A_yBAykUBv1_0;
	wire w_dff_A_rStL3uCh5_0;
	wire w_dff_A_pY3iuBvZ6_0;
	wire w_dff_A_2v8gQzCh1_0;
	wire w_dff_A_7iOw09Wk2_0;
	wire w_dff_A_3EDjtkm78_0;
	wire w_dff_A_LpddJ1ql4_0;
	wire w_dff_A_AERKqKoX2_0;
	wire w_dff_A_Q0Nw8LDx6_0;
	wire w_dff_A_NxLKSlcU2_0;
	wire w_dff_A_rJYzxeyq1_0;
	wire w_dff_A_qWbwLqEz2_0;
	wire w_dff_A_Ck2igJu86_0;
	wire w_dff_A_ASAKMGb29_0;
	wire w_dff_A_APh0v85o0_0;
	wire w_dff_A_cfYMOmt40_0;
	wire w_dff_A_lDPvVcJx8_0;
	wire w_dff_A_0gcyLViY4_0;
	wire w_dff_A_7sM2PFdl2_0;
	wire w_dff_A_Gkt4wVHe7_0;
	wire w_dff_A_wZMYVtAT5_0;
	wire w_dff_A_dR862AWT0_0;
	wire w_dff_A_m3c6GcYD1_1;
	wire w_dff_A_neS8Pgns2_0;
	wire w_dff_A_rdz9Xd5D5_0;
	wire w_dff_A_ztTt08Oi4_0;
	wire w_dff_A_943GbJWl9_0;
	wire w_dff_A_xTFEDmBO1_0;
	wire w_dff_A_nPOe1cdb0_0;
	wire w_dff_A_rXh3dXAu9_0;
	wire w_dff_A_9PXEMyFt7_0;
	wire w_dff_A_UwqongY06_0;
	wire w_dff_A_w0K9tAnF1_0;
	wire w_dff_A_Fb82YPe71_0;
	wire w_dff_A_mstaH5dM2_0;
	wire w_dff_A_S8OODCLB7_0;
	wire w_dff_A_js3HKh461_0;
	wire w_dff_A_oKqEzSjx9_0;
	wire w_dff_A_QJVmFa2Y6_0;
	wire w_dff_A_f87hGuYl5_0;
	wire w_dff_A_XG7333ai6_0;
	wire w_dff_A_cxYubjPU6_0;
	wire w_dff_A_j34uCqX86_0;
	wire w_dff_A_luFbhypQ6_0;
	wire w_dff_A_sM0bIXdM6_0;
	wire w_dff_A_HwhAxqBb0_0;
	wire w_dff_A_vNnowdhk0_0;
	wire w_dff_A_MWNV53vX6_0;
	wire w_dff_A_oLMKUFjx2_0;
	wire w_dff_A_8kp5LDLQ8_0;
	wire w_dff_A_qfQRVDYx2_0;
	wire w_dff_A_m1mERx9q2_0;
	wire w_dff_A_N7UUOuJD4_0;
	wire w_dff_A_Tng41wUW5_0;
	wire w_dff_A_lhCvl2OA6_0;
	wire w_dff_A_2N58DUVH5_0;
	wire w_dff_A_49fNHbAV5_0;
	wire w_dff_A_tvUAzi222_0;
	wire w_dff_A_JnVh7jBS1_0;
	wire w_dff_A_23cXEvfi6_0;
	wire w_dff_A_veXBQrut6_0;
	wire w_dff_A_DbjIJw5y8_1;
	wire w_dff_A_QYSelc0D7_0;
	wire w_dff_A_Tq1uZKXt2_0;
	wire w_dff_A_97EzWTwg3_0;
	wire w_dff_A_FWtycdES8_0;
	wire w_dff_A_R0yC1cZQ9_0;
	wire w_dff_A_Rhv9BR7e1_0;
	wire w_dff_A_dhGNVNjb8_0;
	wire w_dff_A_cmhEXjT05_0;
	wire w_dff_A_UtPqRUnd7_0;
	wire w_dff_A_TRUcJJt18_0;
	wire w_dff_A_64Xz9RBk9_0;
	wire w_dff_A_0l3uT3AI1_0;
	wire w_dff_A_2Ty6CJTh4_0;
	wire w_dff_A_RZ7SBawl7_0;
	wire w_dff_A_Y3wCbXW99_0;
	wire w_dff_A_aqLYkpf27_0;
	wire w_dff_A_Ydp6s5eV0_0;
	wire w_dff_A_vV0R2ADP3_0;
	wire w_dff_A_xz0c9TPD2_0;
	wire w_dff_A_kVaBKblE5_0;
	wire w_dff_A_JzBG10k53_0;
	wire w_dff_A_0QyNtdmT3_0;
	wire w_dff_A_PnpAtMP68_0;
	wire w_dff_A_3zeNyRdK4_0;
	wire w_dff_A_PfcutuxV2_0;
	wire w_dff_A_q7AOk8wm3_0;
	wire w_dff_A_313SaAKf7_0;
	wire w_dff_A_5ST6FeWs7_0;
	wire w_dff_A_VcOPj1xB5_0;
	wire w_dff_A_XrKAWLTg1_0;
	wire w_dff_A_fS3KHqaN9_0;
	wire w_dff_A_dXsAKbSW6_0;
	wire w_dff_A_GcSKwiS31_0;
	wire w_dff_A_hOyQfFMB6_0;
	wire w_dff_A_DFrt3KYs7_0;
	wire w_dff_A_5X3ERRQL3_0;
	wire w_dff_A_4rFzbcav9_0;
	wire w_dff_A_P2HSYyjk1_0;
	wire w_dff_A_b76irSqt9_1;
	wire w_dff_A_reT6XF4V4_0;
	wire w_dff_A_kXX141018_0;
	wire w_dff_A_S3KLaESd4_0;
	wire w_dff_A_P7ViR7n67_0;
	wire w_dff_A_yQLnTgxJ9_0;
	wire w_dff_A_NZ7CLybj4_0;
	wire w_dff_A_cpmCXHgA6_0;
	wire w_dff_A_ILKfShA53_0;
	wire w_dff_A_kzQ9x1E33_0;
	wire w_dff_A_T3Fq2j7j1_0;
	wire w_dff_A_oUahWUZq1_0;
	wire w_dff_A_h4gozfmx1_0;
	wire w_dff_A_Wt2eAbIB6_0;
	wire w_dff_A_bYX0Rqqi9_0;
	wire w_dff_A_a3awiYBU0_0;
	wire w_dff_A_DFBPr1fE6_0;
	wire w_dff_A_lYij1PQv5_0;
	wire w_dff_A_Nz1EZmFF7_0;
	wire w_dff_A_8WRbKEq50_0;
	wire w_dff_A_cvG73VD89_0;
	wire w_dff_A_OUkmg86w7_0;
	wire w_dff_A_CNqfQS2a6_0;
	wire w_dff_A_BdPQEPs52_0;
	wire w_dff_A_EOBdxKmj9_0;
	wire w_dff_A_VwxVqiaW2_0;
	wire w_dff_A_vkFrLgkq8_0;
	wire w_dff_A_DK06YMd55_0;
	wire w_dff_A_bZTLqbwK9_0;
	wire w_dff_A_0FG6J8lp3_0;
	wire w_dff_A_qVey2nH26_0;
	wire w_dff_A_o7YYdPZb8_0;
	wire w_dff_A_8e3NSgGz4_0;
	wire w_dff_A_ZdajZTpo7_0;
	wire w_dff_A_G7pNbg3o5_0;
	wire w_dff_A_t15XqLDb6_0;
	wire w_dff_A_i0uMMR9k8_0;
	wire w_dff_A_RNq0drEK1_0;
	wire w_dff_A_hp9W9RQd6_0;
	wire w_dff_A_TsLfMgku7_1;
	wire w_dff_A_f1O61jzJ1_0;
	wire w_dff_A_Lg3biNeC0_0;
	wire w_dff_A_PCzP35HW3_0;
	wire w_dff_A_X7bcaziw6_0;
	wire w_dff_A_Ew4NW7Qv0_0;
	wire w_dff_A_HR0ph5xB1_0;
	wire w_dff_A_hvp87gTd3_0;
	wire w_dff_A_SnrefMJk4_0;
	wire w_dff_A_3j0jRYW06_0;
	wire w_dff_A_6uMRXNgg4_0;
	wire w_dff_A_6ZoRoiwh3_0;
	wire w_dff_A_YPFnoJnQ3_0;
	wire w_dff_A_fHfI0eZM9_0;
	wire w_dff_A_gRuPA4TU2_0;
	wire w_dff_A_XOH9Vxbi6_0;
	wire w_dff_A_cxzg8MLS7_0;
	wire w_dff_A_IIkQb37F3_0;
	wire w_dff_A_3SrfgKcy4_0;
	wire w_dff_A_H0zE0MqB5_0;
	wire w_dff_A_jEJsBPDI2_0;
	wire w_dff_A_lwdGFB0M9_0;
	wire w_dff_A_E43OOoqb7_0;
	wire w_dff_A_ExYbjIgL7_0;
	wire w_dff_A_N99zULwH4_0;
	wire w_dff_A_Q7DsiNFS6_0;
	wire w_dff_A_Bp9PA9I03_0;
	wire w_dff_A_WHA63cDu3_0;
	wire w_dff_A_88bYetJ04_0;
	wire w_dff_A_aYKkb3F38_0;
	wire w_dff_A_yvuYe1cI1_0;
	wire w_dff_A_ecqAn2cX8_0;
	wire w_dff_A_Qx3u5Vze8_0;
	wire w_dff_A_yLz1uhqc8_0;
	wire w_dff_A_Ec1mXMq14_0;
	wire w_dff_A_Tw0LEMIy5_0;
	wire w_dff_A_eZMBy8LW3_0;
	wire w_dff_A_1VKNnZiP6_0;
	wire w_dff_A_53yowiEy8_0;
	wire w_dff_A_2530MqCy4_1;
	wire w_dff_A_u3ZY1c3w1_0;
	wire w_dff_A_FKw4GYPd0_0;
	wire w_dff_A_2dWXPccF2_0;
	wire w_dff_A_Mxelbxml5_0;
	wire w_dff_A_2HIeRP1a8_0;
	wire w_dff_A_YSnFNhfn7_0;
	wire w_dff_A_dGIOdedb0_0;
	wire w_dff_A_5G15qr067_0;
	wire w_dff_A_m6Kg4wvX6_0;
	wire w_dff_A_9xIV4Aai7_0;
	wire w_dff_A_hP868HXy7_0;
	wire w_dff_A_PmkPx5z52_0;
	wire w_dff_A_7pZIGqW44_0;
	wire w_dff_A_8IEzc5wK7_0;
	wire w_dff_A_SUYVqbea4_0;
	wire w_dff_A_yf7d9Imp7_0;
	wire w_dff_A_sRS5qING4_0;
	wire w_dff_A_T6eia1x64_0;
	wire w_dff_A_rofsiZJc8_0;
	wire w_dff_A_ACNn2aBM3_0;
	wire w_dff_A_uMhffgGd6_0;
	wire w_dff_A_AhsZBdRY8_0;
	wire w_dff_A_iv2h2Ekl5_0;
	wire w_dff_A_lchCOYYE6_0;
	wire w_dff_A_QyxtzM7w5_0;
	wire w_dff_A_pgBbFTUJ7_0;
	wire w_dff_A_VE8bT0ec1_0;
	wire w_dff_A_ULACfosk9_0;
	wire w_dff_A_W8pp6NW67_0;
	wire w_dff_A_5ojiMLSw4_0;
	wire w_dff_A_7kMqU2V71_0;
	wire w_dff_A_bazroMft3_0;
	wire w_dff_A_hI6L4BFx2_0;
	wire w_dff_A_S71oothp2_0;
	wire w_dff_A_1au17JYi4_0;
	wire w_dff_A_ge44J7sP0_0;
	wire w_dff_A_7uUriDOv6_0;
	wire w_dff_A_8sQcEexO1_0;
	wire w_dff_A_LItvViFw0_1;
	wire w_dff_A_hEONwuQo9_0;
	wire w_dff_A_Sup9vN4O5_0;
	wire w_dff_A_owix1sHB2_0;
	wire w_dff_A_RzDwBfp12_0;
	wire w_dff_A_m5KEiS5a3_0;
	wire w_dff_A_T6Tluu1o6_0;
	wire w_dff_A_82rB9WJf6_0;
	wire w_dff_A_JfPR4Bnq9_0;
	wire w_dff_A_KrnNDBXj2_0;
	wire w_dff_A_HKzJ4Kr05_0;
	wire w_dff_A_2z7kxOfK8_0;
	wire w_dff_A_tXpRaclm5_0;
	wire w_dff_A_56rCdv0G7_0;
	wire w_dff_A_idQtLsYp5_0;
	wire w_dff_A_PTbWvBUr4_0;
	wire w_dff_A_oiwUN3C77_0;
	wire w_dff_A_EKyhdG104_0;
	wire w_dff_A_HteDVVk90_0;
	wire w_dff_A_PjyJv4ia5_0;
	wire w_dff_A_qsz4TLkT1_0;
	wire w_dff_A_TBilviF56_0;
	wire w_dff_A_5Hc8v8rE9_0;
	wire w_dff_A_ew6xvEHu8_0;
	wire w_dff_A_NxL9531h2_0;
	wire w_dff_A_W2Baw9qX6_0;
	wire w_dff_A_hV6JXWaV1_0;
	wire w_dff_A_SFVzwpxV7_0;
	wire w_dff_A_fioC63og8_0;
	wire w_dff_A_2D4uhXIu5_0;
	wire w_dff_A_SeTkpVWa2_0;
	wire w_dff_A_gTkDgGKf8_0;
	wire w_dff_A_6Zc7PEBQ8_0;
	wire w_dff_A_XsDY4orp4_0;
	wire w_dff_A_edTETl5E2_0;
	wire w_dff_A_RbL5fwkj5_0;
	wire w_dff_A_U06ymaAX7_0;
	wire w_dff_A_pnwIKx1Y2_0;
	wire w_dff_A_YjjJQKyr1_0;
	wire w_dff_A_vnhaT5SN9_1;
	wire w_dff_A_G9tMNoQa9_0;
	wire w_dff_A_omjDHzPE6_0;
	wire w_dff_A_eLKOlVg81_0;
	wire w_dff_A_oNeJbNLr0_0;
	wire w_dff_A_w8jiqpA43_0;
	wire w_dff_A_L9fEAcTQ1_0;
	wire w_dff_A_Wuql2Nan2_0;
	wire w_dff_A_c5Cq1KLm0_0;
	wire w_dff_A_FtI0Pbei6_0;
	wire w_dff_A_PmH1NPZn3_0;
	wire w_dff_A_qBjKAfGX9_0;
	wire w_dff_A_Wad7dzZ72_0;
	wire w_dff_A_LEBHHY8y6_0;
	wire w_dff_A_7VEdD81l7_0;
	wire w_dff_A_Hes6odD83_0;
	wire w_dff_A_ewM9UXo09_0;
	wire w_dff_A_6EZDpP983_0;
	wire w_dff_A_lPteOT4K6_0;
	wire w_dff_A_G0J0sIXi6_0;
	wire w_dff_A_M4Q3ZGpu8_0;
	wire w_dff_A_68M00IZ28_0;
	wire w_dff_A_1QHzNTzL8_0;
	wire w_dff_A_ZMmhDyv55_0;
	wire w_dff_A_pi1Tr7P82_0;
	wire w_dff_A_ip5Ey8nq0_0;
	wire w_dff_A_j5kHKfiM9_0;
	wire w_dff_A_eLn2iFOw5_0;
	wire w_dff_A_LSff1cIb9_0;
	wire w_dff_A_XCbC5SHI0_0;
	wire w_dff_A_z3hAff878_0;
	wire w_dff_A_QGjGK16B2_0;
	wire w_dff_A_brRFeKfR2_0;
	wire w_dff_A_KkmY2knc5_0;
	wire w_dff_A_BaWrWveG5_0;
	wire w_dff_A_NZQMJ2Hb8_0;
	wire w_dff_A_BAMtfML29_0;
	wire w_dff_A_7MQyo9mS8_0;
	wire w_dff_A_IKXSTLAS2_0;
	wire w_dff_A_LUDcVW948_1;
	wire w_dff_A_X9YYyhJt4_0;
	wire w_dff_A_dfLPMELM5_0;
	wire w_dff_A_WBm55wzQ7_0;
	wire w_dff_A_qund6fSy6_0;
	wire w_dff_A_kbMK0lRx7_0;
	wire w_dff_A_jfdW6br75_0;
	wire w_dff_A_bTQNog3I2_0;
	wire w_dff_A_8pSMHK1a6_0;
	wire w_dff_A_xgzBJHGm1_0;
	wire w_dff_A_hU2l9HEg1_0;
	wire w_dff_A_D3qznDfe4_0;
	wire w_dff_A_JTWzKiJT7_0;
	wire w_dff_A_sRxDq0wE5_0;
	wire w_dff_A_xu2u7iYx8_0;
	wire w_dff_A_HX08QI1R4_0;
	wire w_dff_A_W7tll8Kn7_0;
	wire w_dff_A_w6Uqyi141_0;
	wire w_dff_A_UxCJXwjV5_0;
	wire w_dff_A_znO0lCOk1_0;
	wire w_dff_A_05UaASIe7_0;
	wire w_dff_A_Yb3OQUze3_0;
	wire w_dff_A_MLoAZUGu2_0;
	wire w_dff_A_HGdACXJw5_0;
	wire w_dff_A_wAlFokZx2_0;
	wire w_dff_A_84w4AuBQ4_0;
	wire w_dff_A_v8wXJQ4y2_0;
	wire w_dff_A_F5wxTxZB3_0;
	wire w_dff_A_wk8UXeRf8_0;
	wire w_dff_A_HS9Bc7a39_0;
	wire w_dff_A_2TsYyfjP2_0;
	wire w_dff_A_a4Pl5pdD8_0;
	wire w_dff_A_rJrvrkpQ6_0;
	wire w_dff_A_7hE47G178_0;
	wire w_dff_A_Dzu1FWcg0_0;
	wire w_dff_A_WKTmC0dz8_0;
	wire w_dff_A_GS4gIo068_0;
	wire w_dff_A_klrKteQO1_0;
	wire w_dff_A_i2I4SPfK6_0;
	wire w_dff_A_YgGp9OAD8_1;
	wire w_dff_A_0QlK25Ds0_0;
	wire w_dff_A_zIPE5OUr0_0;
	wire w_dff_A_uaGCy09q6_0;
	wire w_dff_A_GwBIRKze0_0;
	wire w_dff_A_EE7qzUBt2_0;
	wire w_dff_A_3Sn0e4Ym4_0;
	wire w_dff_A_i515ZKvw2_0;
	wire w_dff_A_Bf7dUFB88_0;
	wire w_dff_A_LQzbzHAh7_0;
	wire w_dff_A_3kC3B4rI8_0;
	wire w_dff_A_NQmCufV21_0;
	wire w_dff_A_iT40sNiM0_0;
	wire w_dff_A_gkCiHrCh7_0;
	wire w_dff_A_BKY44R154_0;
	wire w_dff_A_zb4o4c8M6_0;
	wire w_dff_A_SJtMSAf81_0;
	wire w_dff_A_KflnuDOR8_0;
	wire w_dff_A_i8eqpaAh1_0;
	wire w_dff_A_UXEqZ9wj2_0;
	wire w_dff_A_ySpLjSze5_0;
	wire w_dff_A_05agX0Ev1_0;
	wire w_dff_A_F5elunu49_0;
	wire w_dff_A_XtB4WoBz8_0;
	wire w_dff_A_S6EMwAXX9_0;
	wire w_dff_A_nGSzjTJM9_0;
	wire w_dff_A_emgDBOkS0_0;
	wire w_dff_A_ecjFM3G38_0;
	wire w_dff_A_nhhOIW3N3_0;
	wire w_dff_A_Ag1zIeCj0_0;
	wire w_dff_A_1VwfO0Fo5_0;
	wire w_dff_A_45jw5LT38_0;
	wire w_dff_A_FmChxGpk6_0;
	wire w_dff_A_JCxyAt8p3_0;
	wire w_dff_A_4SCFmmLB0_0;
	wire w_dff_A_eMK9UIsO4_0;
	wire w_dff_A_6UmeON7q0_0;
	wire w_dff_A_0nYxeyv95_0;
	wire w_dff_A_GY6VqlmW0_0;
	wire w_dff_A_0NogE0yY4_1;
	wire w_dff_A_Nvdx9tAO0_0;
	wire w_dff_A_Ott9JlcE6_0;
	wire w_dff_A_kzTENg772_0;
	wire w_dff_A_LCANN16k2_0;
	wire w_dff_A_Lkyqgqbx3_0;
	wire w_dff_A_zu0QWtS43_0;
	wire w_dff_A_OGLDDCL70_0;
	wire w_dff_A_z6yUUIVR2_0;
	wire w_dff_A_GBbJVQwi5_0;
	wire w_dff_A_8DZfy4kQ5_0;
	wire w_dff_A_RjhtBDwM8_0;
	wire w_dff_A_CdEYTqNb2_0;
	wire w_dff_A_evSR5vPu2_0;
	wire w_dff_A_0gEGOtzx8_0;
	wire w_dff_A_bFOhM57K2_0;
	wire w_dff_A_IwRwMLat5_0;
	wire w_dff_A_FafZDnee1_0;
	wire w_dff_A_Hzm2QZ7G8_0;
	wire w_dff_A_VKymOSal2_0;
	wire w_dff_A_PorutfbF3_0;
	wire w_dff_A_qJeIaSCR4_0;
	wire w_dff_A_234ifCIy2_0;
	wire w_dff_A_3zfAX6XL4_0;
	wire w_dff_A_9a46uQbX8_0;
	wire w_dff_A_fgPiidmh7_0;
	wire w_dff_A_knJEV6iV6_0;
	wire w_dff_A_ZDYYDH1t9_0;
	wire w_dff_A_PeQX62QY1_0;
	wire w_dff_A_16dSxHqO9_0;
	wire w_dff_A_xOsVZGl18_0;
	wire w_dff_A_0BcjZkzi9_0;
	wire w_dff_A_gFbqdkQx3_0;
	wire w_dff_A_bRh5qoeL9_0;
	wire w_dff_A_nhbAUFk49_0;
	wire w_dff_A_WZGRpOHd1_0;
	wire w_dff_A_P9H4QUlG4_0;
	wire w_dff_A_zkyjy38M1_0;
	wire w_dff_A_yETswr8r4_0;
	wire w_dff_A_B1CtAN1E0_1;
	wire w_dff_A_x0z06xRE3_0;
	wire w_dff_A_RFDGyIYF6_0;
	wire w_dff_A_QEehQPA88_0;
	wire w_dff_A_qrPugM7A5_0;
	wire w_dff_A_UAMn1Up06_0;
	wire w_dff_A_gMuqVDUc9_0;
	wire w_dff_A_aUGvikyU2_0;
	wire w_dff_A_FiS1OJIh8_0;
	wire w_dff_A_Zl9N27pS1_0;
	wire w_dff_A_6a4R9skz6_0;
	wire w_dff_A_ysZsao199_0;
	wire w_dff_A_C2rjcaTl9_0;
	wire w_dff_A_jeNX7dG11_0;
	wire w_dff_A_7xhBNyUp1_0;
	wire w_dff_A_190ctC065_0;
	wire w_dff_A_eTZUHcvB5_0;
	wire w_dff_A_5mB3WdhG2_0;
	wire w_dff_A_geMJTZzl9_0;
	wire w_dff_A_s3bH4qku5_0;
	wire w_dff_A_1ce1HdOi2_0;
	wire w_dff_A_ADOZWDe22_0;
	wire w_dff_A_WvcocX5X9_0;
	wire w_dff_A_SbKRXqAB1_0;
	wire w_dff_A_wLr2L8Pe8_0;
	wire w_dff_A_aVeR2SgY8_0;
	wire w_dff_A_qN2rgI7h4_0;
	wire w_dff_A_d2Leqkyp2_0;
	wire w_dff_A_bGGfmgPl6_0;
	wire w_dff_A_go56ikbc7_0;
	wire w_dff_A_f3CHvaWl7_0;
	wire w_dff_A_jqQC6r8m8_0;
	wire w_dff_A_aBGzrkyQ3_0;
	wire w_dff_A_Za1zlMD60_0;
	wire w_dff_A_qzfSJFPC9_0;
	wire w_dff_A_rT8MbJeM2_0;
	wire w_dff_A_gJXzCv1j1_0;
	wire w_dff_A_Vi5XxNHS2_0;
	wire w_dff_A_L53p63RB4_0;
	wire w_dff_A_OfvxdAZI9_1;
	wire w_dff_A_u6w11RdQ8_0;
	wire w_dff_A_gVfvJfFu9_0;
	wire w_dff_A_6qP8pnkO8_0;
	wire w_dff_A_0evuJGdV0_0;
	wire w_dff_A_gQNLP9a55_0;
	wire w_dff_A_WguEMg0S5_0;
	wire w_dff_A_3kZrnrwH9_0;
	wire w_dff_A_72MKYkRT3_0;
	wire w_dff_A_oQxkLytR8_0;
	wire w_dff_A_OnQOin4c2_0;
	wire w_dff_A_mAzHswCT5_0;
	wire w_dff_A_O64vvKgi2_0;
	wire w_dff_A_r6ffcCki1_0;
	wire w_dff_A_UMKyvzuM8_0;
	wire w_dff_A_AyJ4YQeu2_0;
	wire w_dff_A_0RHyS6RY9_0;
	wire w_dff_A_lN8WtdiX8_0;
	wire w_dff_A_09I1zbWa9_0;
	wire w_dff_A_zX5IKqPQ7_0;
	wire w_dff_A_lhmmAC7S3_0;
	wire w_dff_A_4auHpJRm7_0;
	wire w_dff_A_2i9WPWth9_0;
	wire w_dff_A_aPEbTLQu3_0;
	wire w_dff_A_K4uzrSny2_0;
	wire w_dff_A_Y16NZxXz7_0;
	wire w_dff_A_Kz7a0dJK3_0;
	wire w_dff_A_Qxtx3XIQ0_0;
	wire w_dff_A_F6jp2qLA6_0;
	wire w_dff_A_h61LNy6v1_0;
	wire w_dff_A_n7aRZqte7_0;
	wire w_dff_A_1wnQql9o7_0;
	wire w_dff_A_Geec7v7P3_0;
	wire w_dff_A_BSKXJ16d3_0;
	wire w_dff_A_3nrr3Pyi6_0;
	wire w_dff_A_c6DmA7c72_0;
	wire w_dff_A_seyxrpUW8_0;
	wire w_dff_A_KVv70fzu6_0;
	wire w_dff_A_cWBRYjaq1_0;
	wire w_dff_A_raA4ZSOf6_1;
	wire w_dff_A_JsonzD2n9_0;
	wire w_dff_A_1FEFb6k40_0;
	wire w_dff_A_27xWi6MH1_0;
	wire w_dff_A_RRigINkF0_0;
	wire w_dff_A_dNvhmzVZ6_0;
	wire w_dff_A_YifYED4m2_0;
	wire w_dff_A_YwG0u98N9_0;
	wire w_dff_A_agu1s1IU2_0;
	wire w_dff_A_H8w1aGhe8_0;
	wire w_dff_A_b20fpsaN7_0;
	wire w_dff_A_6o3FVUH64_0;
	wire w_dff_A_6YCWbd2H3_0;
	wire w_dff_A_JXZK6Gig5_0;
	wire w_dff_A_u4giKg3J1_0;
	wire w_dff_A_tnzplJ4T0_0;
	wire w_dff_A_CIdePGpv1_0;
	wire w_dff_A_xYfrSgnN8_0;
	wire w_dff_A_8c83QNxC2_0;
	wire w_dff_A_JTDxKvRv8_0;
	wire w_dff_A_UnKXg5GR2_0;
	wire w_dff_A_aZvQrLwx4_0;
	wire w_dff_A_3LWuqz2S5_0;
	wire w_dff_A_5NwHhuGE2_0;
	wire w_dff_A_NKpto9AQ6_0;
	wire w_dff_A_PhVbRa9F6_0;
	wire w_dff_A_vJ3Libtc0_0;
	wire w_dff_A_jJSL0Y978_0;
	wire w_dff_A_fPdXwmPX5_0;
	wire w_dff_A_rQPHKf2f9_0;
	wire w_dff_A_2uHhfrbJ5_0;
	wire w_dff_A_H7igYsBG8_0;
	wire w_dff_A_PCJQs6Ti8_0;
	wire w_dff_A_ZLxdT2nR1_0;
	wire w_dff_A_1WBCEbt64_0;
	wire w_dff_A_qEqrCszF4_0;
	wire w_dff_A_D1bRoyE32_0;
	wire w_dff_A_zl51YVJi4_0;
	wire w_dff_A_AYvTdkIM1_0;
	wire w_dff_A_cdzx6Owo0_1;
	wire w_dff_A_Q2vYo6iT3_0;
	wire w_dff_A_I2nAqOy29_0;
	wire w_dff_A_hEW80LHj8_0;
	wire w_dff_A_5AqO0yc54_0;
	wire w_dff_A_sFVRGxik1_0;
	wire w_dff_A_fBSuky5A1_0;
	wire w_dff_A_78wQVgxb4_0;
	wire w_dff_A_uRcIAe7U4_0;
	wire w_dff_A_XopxEOvI9_0;
	wire w_dff_A_DQ2lfse11_0;
	wire w_dff_A_rlQG7AFW3_0;
	wire w_dff_A_FmaAT13e0_0;
	wire w_dff_A_lYEkRAoq4_0;
	wire w_dff_A_3K9slGGc9_0;
	wire w_dff_A_8Lc4IL521_0;
	wire w_dff_A_10MirRNo9_0;
	wire w_dff_A_4ZLUGN9Y2_0;
	wire w_dff_A_CIYjPe135_0;
	wire w_dff_A_lRt2hjzH2_0;
	wire w_dff_A_HYYqvbGz5_0;
	wire w_dff_A_fNzDb7rS7_0;
	wire w_dff_A_h4oIc3Mn2_0;
	wire w_dff_A_tX8PkE9y2_0;
	wire w_dff_A_BOgF5B9s8_0;
	wire w_dff_A_uV0C22BX2_0;
	wire w_dff_A_GZxWhTm66_0;
	wire w_dff_A_azJgPFh68_0;
	wire w_dff_A_Gf4MZAsF8_0;
	wire w_dff_A_AfH548px0_0;
	wire w_dff_A_12qmTvYC5_0;
	wire w_dff_A_zOE9RhDo4_0;
	wire w_dff_A_nT8oR8Zy9_0;
	wire w_dff_A_wdPlmwse4_0;
	wire w_dff_A_0iLuSKBQ0_0;
	wire w_dff_A_c4LIxd3n2_0;
	wire w_dff_A_QgJWroce0_0;
	wire w_dff_A_nbgJAfPH5_0;
	wire w_dff_A_RHmuEuxu0_0;
	wire w_dff_A_34A5K7yA7_1;
	wire w_dff_A_YYy4sqko7_0;
	wire w_dff_A_O6WxUSNV2_0;
	wire w_dff_A_Hww3Vx2F3_0;
	wire w_dff_A_nZ8o2BWI4_0;
	wire w_dff_A_wn9mJYof6_0;
	wire w_dff_A_pjOWfvd54_0;
	wire w_dff_A_Kr9kCJOH5_0;
	wire w_dff_A_wg2BCycD8_0;
	wire w_dff_A_MYe3cHNE2_0;
	wire w_dff_A_w9IBA8XL6_0;
	wire w_dff_A_2nDwcplW4_0;
	wire w_dff_A_h535TGIq5_0;
	wire w_dff_A_rOou0g5I4_0;
	wire w_dff_A_cgo5ybVO1_0;
	wire w_dff_A_AI6EbtoA9_0;
	wire w_dff_A_YDJNwgpP5_0;
	wire w_dff_A_QPrX51YL7_0;
	wire w_dff_A_Es8ZUgLv8_0;
	wire w_dff_A_0GRQwzjl4_0;
	wire w_dff_A_mLHrelrP7_0;
	wire w_dff_A_8cuvPt7V1_0;
	wire w_dff_A_NwBWVVcX1_0;
	wire w_dff_A_Dx9qxdNX2_0;
	wire w_dff_A_F4ma6W6j2_0;
	wire w_dff_A_rEMHaQ3A4_0;
	wire w_dff_A_6Fu8ZWVr2_0;
	wire w_dff_A_NAg3yQwV2_0;
	wire w_dff_A_bWPxweDt0_0;
	wire w_dff_A_FZEVdlcS9_0;
	wire w_dff_A_JxgndWWk8_0;
	wire w_dff_A_0cIJTg6E1_0;
	wire w_dff_A_2DR5c3VK1_0;
	wire w_dff_A_YJoPn7qq5_0;
	wire w_dff_A_Ixrh25oI7_0;
	wire w_dff_A_XvcRrPbp4_0;
	wire w_dff_A_2AAweAFa4_0;
	wire w_dff_A_KKwDUADl4_0;
	wire w_dff_A_tCT5eKfd3_0;
	wire w_dff_A_kb3quiGP8_1;
	wire w_dff_A_sws1mcak6_0;
	wire w_dff_A_eHVzY1QB8_0;
	wire w_dff_A_7T5N5bgl5_0;
	wire w_dff_A_YN3Svbd34_0;
	wire w_dff_A_tWWm99yc8_0;
	wire w_dff_A_t2wWbrph2_0;
	wire w_dff_A_4Z18cAcd1_0;
	wire w_dff_A_YRGoSWNz9_0;
	wire w_dff_A_jGCQWyix8_0;
	wire w_dff_A_jgC289Hi2_0;
	wire w_dff_A_dno8tfrB2_0;
	wire w_dff_A_4i6coCeV3_0;
	wire w_dff_A_jzC4GcB65_0;
	wire w_dff_A_XACZ4ObN1_0;
	wire w_dff_A_8unOYwrm5_0;
	wire w_dff_A_JZ8Zvg5O6_0;
	wire w_dff_A_qZ7Ldncm9_0;
	wire w_dff_A_LbQ70CBp4_0;
	wire w_dff_A_815YWJ2x8_0;
	wire w_dff_A_vH264ND87_0;
	wire w_dff_A_flJHiBxc1_0;
	wire w_dff_A_G0wH6e5i3_0;
	wire w_dff_A_DltdmxHx7_0;
	wire w_dff_A_ByPB2ARu6_0;
	wire w_dff_A_Olq6KVgr2_0;
	wire w_dff_A_vs1JXJ5y8_0;
	wire w_dff_A_Xfkpeue67_0;
	wire w_dff_A_aR3Sna410_0;
	wire w_dff_A_6VorzEux4_0;
	wire w_dff_A_ELM2bTzb3_0;
	wire w_dff_A_YJuaxuA56_0;
	wire w_dff_A_7PtTTNbd7_0;
	wire w_dff_A_blD2RiJn5_0;
	wire w_dff_A_nVDlxkkq5_0;
	wire w_dff_A_yGDEcFTE9_0;
	wire w_dff_A_lx6OzEzQ5_0;
	wire w_dff_A_mbyBwvos9_0;
	wire w_dff_A_Vj1kNBeA7_0;
	wire w_dff_A_5GiWzOQF0_1;
	wire w_dff_A_aEpl5dPU0_0;
	wire w_dff_A_5oSoT8jO1_0;
	wire w_dff_A_rwVjqHsJ6_0;
	wire w_dff_A_dp23amMn5_0;
	wire w_dff_A_WJcD30dT3_0;
	wire w_dff_A_scoYqcGf7_0;
	wire w_dff_A_jBFjaZrK3_0;
	wire w_dff_A_hZNQNLVY3_0;
	wire w_dff_A_1ahuj7sp4_0;
	wire w_dff_A_eC30xmAe9_0;
	wire w_dff_A_aEG3ns3P3_0;
	wire w_dff_A_EWZHG3wT8_0;
	wire w_dff_A_WXYRMgKc2_0;
	wire w_dff_A_WqG2lU4F2_0;
	wire w_dff_A_n2XbPuEm2_0;
	wire w_dff_A_dodAIOqs3_0;
	wire w_dff_A_5eikFxYu7_0;
	wire w_dff_A_aFKANECi0_0;
	wire w_dff_A_MeBg5q7G5_0;
	wire w_dff_A_sMTyoztj8_0;
	wire w_dff_A_MZSXbWH45_0;
	wire w_dff_A_749LB0Xs8_0;
	wire w_dff_A_pudogwcz5_0;
	wire w_dff_A_Tj3pnvvU6_0;
	wire w_dff_A_Aioi3WAO4_0;
	wire w_dff_A_00lnqNId7_0;
	wire w_dff_A_yNqaZA5K5_0;
	wire w_dff_A_Jt4d8DcT6_0;
	wire w_dff_A_Ag6yEwyO8_0;
	wire w_dff_A_GgSRjkx82_0;
	wire w_dff_A_ghQsRmtn1_0;
	wire w_dff_A_SvIOz8Nl1_0;
	wire w_dff_A_ZItLgTyd3_0;
	wire w_dff_A_8rHoO3FM4_0;
	wire w_dff_A_kld8f9Z77_0;
	wire w_dff_A_Kj5KJFDM7_0;
	wire w_dff_A_2KX31jHY6_0;
	wire w_dff_A_0nfS8F1I7_0;
	wire w_dff_A_vkEKZ9tY8_1;
	wire w_dff_A_3Hga92oZ0_0;
	wire w_dff_A_khtVPgM78_0;
	wire w_dff_A_11Wyybou4_0;
	wire w_dff_A_WoMGRrGq8_0;
	wire w_dff_A_M3jD6m6m0_0;
	wire w_dff_A_dp2iTbNE4_0;
	wire w_dff_A_2zauRqPv3_0;
	wire w_dff_A_Iv07XKB11_0;
	wire w_dff_A_AYcvrKBm4_0;
	wire w_dff_A_USkBZdhj3_0;
	wire w_dff_A_Hl6BNh9y6_0;
	wire w_dff_A_gq3eAXEG8_0;
	wire w_dff_A_qNoK2uQk1_0;
	wire w_dff_A_1SmrEwel9_0;
	wire w_dff_A_YydFjzVM7_0;
	wire w_dff_A_W2mIK5yg7_0;
	wire w_dff_A_03IhAZp77_0;
	wire w_dff_A_aB6KPaFm9_0;
	wire w_dff_A_skQ4Dmx88_0;
	wire w_dff_A_YWqL8S1h1_0;
	wire w_dff_A_AKbjk9nv2_0;
	wire w_dff_A_F8RXZ21P3_0;
	wire w_dff_A_T8jB2xNd3_0;
	wire w_dff_A_dJsbkDX95_0;
	wire w_dff_A_axCQjWg46_0;
	wire w_dff_A_FjIr2JJr1_0;
	wire w_dff_A_zInnHBRp3_0;
	wire w_dff_A_yBWDkHuo3_0;
	wire w_dff_A_xuEmGywE2_0;
	wire w_dff_A_5OVNLf8I4_0;
	wire w_dff_A_oHn3GFpu5_0;
	wire w_dff_A_zEXVDgTy4_0;
	wire w_dff_A_0fTmNK6w1_0;
	wire w_dff_A_PW9dBE841_0;
	wire w_dff_A_h5mQSizS4_0;
	wire w_dff_A_cROyc4D50_0;
	wire w_dff_A_ZInPEIfL0_0;
	wire w_dff_A_5DMb0lvz5_0;
	wire w_dff_A_Y0XsnTNc9_1;
	wire w_dff_A_T7a8vy667_0;
	wire w_dff_A_QjisMclL7_0;
	wire w_dff_A_V1nFNSGM9_0;
	wire w_dff_A_l7ShLEp08_0;
	wire w_dff_A_ogvvfXQc4_0;
	wire w_dff_A_daaCWMT53_0;
	wire w_dff_A_cbH8fffg2_0;
	wire w_dff_A_YKAcz1qg2_0;
	wire w_dff_A_YYzpSPer0_0;
	wire w_dff_A_WbSzd5fG5_0;
	wire w_dff_A_Vxafupq79_0;
	wire w_dff_A_obNLe7ck8_0;
	wire w_dff_A_RRVBhwzk0_0;
	wire w_dff_A_sZ87DjIv2_0;
	wire w_dff_A_7vDfyxsn6_0;
	wire w_dff_A_puks27fJ6_0;
	wire w_dff_A_TCDd4YRd4_0;
	wire w_dff_A_gopMhbKD8_0;
	wire w_dff_A_ZX7d4pxK9_0;
	wire w_dff_A_fPIXqN9E5_0;
	wire w_dff_A_LSPT52hn1_0;
	wire w_dff_A_GqLBgOHo7_0;
	wire w_dff_A_j42bWZsS5_0;
	wire w_dff_A_M8vHD1Ac8_0;
	wire w_dff_A_O4HCTYPZ1_0;
	wire w_dff_A_pd5eUize2_0;
	wire w_dff_A_y6qSF2Ev1_0;
	wire w_dff_A_w3E732Vl5_0;
	wire w_dff_A_D5suDTaQ3_0;
	wire w_dff_A_bu96vTmr7_0;
	wire w_dff_A_5rZ717lo4_0;
	wire w_dff_A_2toj0yy12_0;
	wire w_dff_A_vcT4gfum4_0;
	wire w_dff_A_xovUDJzy7_0;
	wire w_dff_A_2Pbeh5Cg0_0;
	wire w_dff_A_aPMfGfWe8_0;
	wire w_dff_A_P0SWuub67_0;
	wire w_dff_A_yVsYAMKi6_0;
	wire w_dff_A_o22oslEs2_1;
	wire w_dff_A_SWudl3fH6_0;
	wire w_dff_A_kFYwmWPx8_0;
	wire w_dff_A_GjjemOjO5_0;
	wire w_dff_A_Wd24Repo5_0;
	wire w_dff_A_mcIabQoo0_0;
	wire w_dff_A_vNWVtsxY0_0;
	wire w_dff_A_LbyYWF4Z8_0;
	wire w_dff_A_SNaNUHVy7_0;
	wire w_dff_A_iLDs1PeX6_0;
	wire w_dff_A_icN3eGbN8_0;
	wire w_dff_A_3qNU8Oj16_0;
	wire w_dff_A_iGRTyvPk4_0;
	wire w_dff_A_lrSiQmtD4_0;
	wire w_dff_A_yN2i2zPk7_0;
	wire w_dff_A_Lt70lOct4_0;
	wire w_dff_A_UE6mAHTh1_0;
	wire w_dff_A_MvkKaeaj4_0;
	wire w_dff_A_tgX9iR9T3_0;
	wire w_dff_A_OmA1Ya523_0;
	wire w_dff_A_aw5W9kgK5_0;
	wire w_dff_A_QxQyy5JU8_0;
	wire w_dff_A_mVzhrwoW5_0;
	wire w_dff_A_fBcNLUnm6_0;
	wire w_dff_A_v2B4HLeQ0_0;
	wire w_dff_A_4IbIkKsT0_0;
	wire w_dff_A_Hg0LsFs22_0;
	wire w_dff_A_jxZF3BAR8_0;
	wire w_dff_A_PSWajxFq8_0;
	wire w_dff_A_3cptEHxw6_0;
	wire w_dff_A_DNGDY2Ph1_0;
	wire w_dff_A_FCCMkWCz6_0;
	wire w_dff_A_suDbfMfF5_0;
	wire w_dff_A_BIMIoinK2_0;
	wire w_dff_A_Qmvh1YgZ5_0;
	wire w_dff_A_ma8oUp8w2_0;
	wire w_dff_A_ODou38dY2_0;
	wire w_dff_A_krEJdneQ4_0;
	wire w_dff_A_Hf7d0RiV9_0;
	wire w_dff_A_HR72Rhmh8_1;
	wire w_dff_A_L4mAU5u48_0;
	wire w_dff_A_Up0ZXbfK1_0;
	wire w_dff_A_aCiQFfaL4_0;
	wire w_dff_A_NOXl3xAN5_0;
	wire w_dff_A_JXLM4iq89_0;
	wire w_dff_A_UaeNUpip8_0;
	wire w_dff_A_HjgzRhnt0_0;
	wire w_dff_A_6lXovPbp7_0;
	wire w_dff_A_O9BjyBi62_0;
	wire w_dff_A_ltnuCPoY6_0;
	wire w_dff_A_1dPmnWAJ4_0;
	wire w_dff_A_mljuEguS8_0;
	wire w_dff_A_T7uqPioX1_0;
	wire w_dff_A_lsku68HW7_0;
	wire w_dff_A_p1O28qaI2_0;
	wire w_dff_A_YVGVUQl08_0;
	wire w_dff_A_xGPAdEvR3_0;
	wire w_dff_A_gH1sdyky3_0;
	wire w_dff_A_JSSzHHmi4_0;
	wire w_dff_A_o9yy6nCv3_0;
	wire w_dff_A_LNP5akWZ2_0;
	wire w_dff_A_q0fcwMf04_0;
	wire w_dff_A_bfcZ9Axs7_0;
	wire w_dff_A_kwuIIMe07_0;
	wire w_dff_A_2tNBqF4j3_0;
	wire w_dff_A_ifLkofgn5_0;
	wire w_dff_A_17OsI95U8_0;
	wire w_dff_A_Bhm3YoXP9_0;
	wire w_dff_A_UD468PUo7_0;
	wire w_dff_A_uWKsv6AY7_0;
	wire w_dff_A_fJGcvVX29_0;
	wire w_dff_A_UlHOXTTj5_0;
	wire w_dff_A_0qOKb5Iz9_0;
	wire w_dff_A_HSPwinYF8_0;
	wire w_dff_A_vnHQNcEU3_0;
	wire w_dff_A_I4409HAU4_0;
	wire w_dff_A_CWbfRxkb1_0;
	wire w_dff_A_Lh4jv2Bj5_0;
	wire w_dff_A_p7sM1NwD4_1;
	wire w_dff_A_ZwzT2qxk8_0;
	wire w_dff_A_60tzlkKa4_0;
	wire w_dff_A_M8i6pD6M0_0;
	wire w_dff_A_DJpZwrAq2_0;
	wire w_dff_A_BV8BsgHy2_0;
	wire w_dff_A_XOhjJSgs0_0;
	wire w_dff_A_3nNodtXk4_0;
	wire w_dff_A_CdQnmaiK3_0;
	wire w_dff_A_34PWiVlI1_0;
	wire w_dff_A_5Be4p3Dh1_0;
	wire w_dff_A_36NETdFm6_0;
	wire w_dff_A_Q8eqRP257_0;
	wire w_dff_A_iWGNhWis4_0;
	wire w_dff_A_qsE37HYN4_0;
	wire w_dff_A_PsNvbgbS2_0;
	wire w_dff_A_A8yPce9r5_0;
	wire w_dff_A_DSKIPWAX9_0;
	wire w_dff_A_5I0lhWkl6_0;
	wire w_dff_A_hHgjl12u8_0;
	wire w_dff_A_tS3kruGW0_0;
	wire w_dff_A_G6YL1vPH1_0;
	wire w_dff_A_DEhrCFrZ9_0;
	wire w_dff_A_dXGZVzsO6_0;
	wire w_dff_A_rSHqQfRY7_0;
	wire w_dff_A_ZOlQ0VHj1_0;
	wire w_dff_A_k866hyE98_0;
	wire w_dff_A_woUojX6s0_0;
	wire w_dff_A_LKGX8AmU1_0;
	wire w_dff_A_dgIvbyZM9_0;
	wire w_dff_A_mhqGb4EO9_0;
	wire w_dff_A_CijkUDh53_0;
	wire w_dff_A_vAxk4ePj9_0;
	wire w_dff_A_VyuPYwbb9_0;
	wire w_dff_A_hWwlbegk8_0;
	wire w_dff_A_JByeqisy2_0;
	wire w_dff_A_a1bUKP9I2_0;
	wire w_dff_A_4hl7L4aQ1_0;
	wire w_dff_A_eHE9IdWZ8_0;
	wire w_dff_A_vAZbA4Z74_1;
	wire w_dff_A_2MMp62kH6_0;
	wire w_dff_A_Uezq7o1B3_0;
	wire w_dff_A_BhLPUd8a5_0;
	wire w_dff_A_DjgBeDDH9_0;
	wire w_dff_A_PGkMPdFJ2_0;
	wire w_dff_A_yEbciAXi2_0;
	wire w_dff_A_dbq3GH680_0;
	wire w_dff_A_xEQ4c4kd0_0;
	wire w_dff_A_4M4XRUCz6_0;
	wire w_dff_A_SgUjyxAP9_0;
	wire w_dff_A_vrW4C4ix7_0;
	wire w_dff_A_m7BdAZj59_0;
	wire w_dff_A_3kbH9r0a1_0;
	wire w_dff_A_0AAUV0yJ2_0;
	wire w_dff_A_pjfqcciz7_0;
	wire w_dff_A_8wtueMno8_0;
	wire w_dff_A_WB0DWFEg4_0;
	wire w_dff_A_gjvpN5Wr2_0;
	wire w_dff_A_QbzNtfmz9_0;
	wire w_dff_A_Pugu3RvD2_0;
	wire w_dff_A_dw9GOxEv1_0;
	wire w_dff_A_AR1CtIRJ8_0;
	wire w_dff_A_lh3xLDUg4_0;
	wire w_dff_A_CwQlRBn45_0;
	wire w_dff_A_UUSNmJRB2_0;
	wire w_dff_A_RxD0gh791_0;
	wire w_dff_A_GU26L0L16_0;
	wire w_dff_A_Q8SU1OhR9_0;
	wire w_dff_A_7YbTRTcE1_0;
	wire w_dff_A_UKvk0YiI1_0;
	wire w_dff_A_kpItN9ID0_0;
	wire w_dff_A_KwL4tTzp8_0;
	wire w_dff_A_zxTDcH0z3_0;
	wire w_dff_A_70CmHYck2_0;
	wire w_dff_A_fJ82zzi54_0;
	wire w_dff_A_zAl7ihCX2_0;
	wire w_dff_A_HZt1AhWg5_0;
	wire w_dff_A_sFNRtXSA0_0;
	wire w_dff_A_mt2rqSeK3_1;
	wire w_dff_A_xbmFH1iK5_0;
	wire w_dff_A_xbiJKr2Z6_0;
	wire w_dff_A_ofcDf6b19_0;
	wire w_dff_A_qpW2n5U76_0;
	wire w_dff_A_LFeS4H0z5_0;
	wire w_dff_A_qGOcPXK40_0;
	wire w_dff_A_C734e5R69_0;
	wire w_dff_A_ZaUUDSYa3_0;
	wire w_dff_A_l3d6zRP65_0;
	wire w_dff_A_YbJHumxK4_0;
	wire w_dff_A_sFKswxqH0_0;
	wire w_dff_A_xv7CYBWv2_0;
	wire w_dff_A_79wXGOJO1_0;
	wire w_dff_A_fMCP0aMa3_0;
	wire w_dff_A_VSwDGCem0_0;
	wire w_dff_A_1pvS7Uzg9_0;
	wire w_dff_A_Tl4ODZsD9_0;
	wire w_dff_A_typFEyuf4_0;
	wire w_dff_A_2tOivj167_0;
	wire w_dff_A_lToGJ2b27_0;
	wire w_dff_A_0o5o424W3_0;
	wire w_dff_A_YOz7mk6i7_0;
	wire w_dff_A_rORy3Q6Z9_0;
	wire w_dff_A_S9ryIOuu0_0;
	wire w_dff_A_YPgn7Exi0_0;
	wire w_dff_A_dsE7BO5X6_0;
	wire w_dff_A_rfFe7aCU5_0;
	wire w_dff_A_a6mlJYpW4_0;
	wire w_dff_A_MbLrLki79_0;
	wire w_dff_A_7XMwCsdi2_0;
	wire w_dff_A_KCKSzwGq7_0;
	wire w_dff_A_zshp0VFt3_0;
	wire w_dff_A_DMiGRzAQ7_0;
	wire w_dff_A_mtQZz3yC9_0;
	wire w_dff_A_ov4lPmoW6_0;
	wire w_dff_A_KyCXR99V6_0;
	wire w_dff_A_VvZqcXFo5_0;
	wire w_dff_A_PHcpn06L7_0;
	wire w_dff_A_TSybH3fu9_1;
	wire w_dff_A_wUfJfbab4_0;
	wire w_dff_A_dxnGsKwm7_0;
	wire w_dff_A_111G5MnE0_0;
	wire w_dff_A_ruUpCu2q4_0;
	wire w_dff_A_iviRMjc33_0;
	wire w_dff_A_YM5RG50y9_0;
	wire w_dff_A_ueBud0cC9_0;
	wire w_dff_A_k6wISBbL2_0;
	wire w_dff_A_0IzXZe2J3_0;
	wire w_dff_A_dGVSNvSl7_0;
	wire w_dff_A_O5oDpgQH9_0;
	wire w_dff_A_0b6JbqDN7_0;
	wire w_dff_A_vgVSCNHd1_0;
	wire w_dff_A_Pv71OZNk7_0;
	wire w_dff_A_NhKCvbut6_0;
	wire w_dff_A_C3Qvz7a30_0;
	wire w_dff_A_LC7wDpGe7_0;
	wire w_dff_A_6BkqTbXD3_0;
	wire w_dff_A_NFdnTzuk7_0;
	wire w_dff_A_p78Ohcai2_0;
	wire w_dff_A_zvbxpQgT1_0;
	wire w_dff_A_voC7HsMn0_0;
	wire w_dff_A_7BzzUeIZ2_0;
	wire w_dff_A_qz6BamNr6_0;
	wire w_dff_A_4uXHtAva8_0;
	wire w_dff_A_DMAjX8Vy8_0;
	wire w_dff_A_K06MPBqo0_0;
	wire w_dff_A_cpZusPVZ8_0;
	wire w_dff_A_hX9yW4Hs7_0;
	wire w_dff_A_17jpNigM5_0;
	wire w_dff_A_PABwR32d7_0;
	wire w_dff_A_EHAb92WK2_0;
	wire w_dff_A_nsGyaO1J4_0;
	wire w_dff_A_yiwkFo8X6_0;
	wire w_dff_A_Ii6OrUsK4_0;
	wire w_dff_A_iuSd4yFD0_0;
	wire w_dff_A_F8U0IhfW5_0;
	wire w_dff_A_l1LtiW1L5_1;
	wire w_dff_A_n2eZmFw13_0;
	wire w_dff_A_VD6nyx6i9_0;
	wire w_dff_A_0ZU42tqb6_0;
	wire w_dff_A_oHR3riFy7_0;
	wire w_dff_A_fyxfenTr9_0;
	wire w_dff_A_c8uAtUer9_0;
	wire w_dff_A_hItoQ4gS7_0;
	wire w_dff_A_sWW8MIeX3_0;
	wire w_dff_A_z7J0neZo6_0;
	wire w_dff_A_aSMoqDED7_0;
	wire w_dff_A_zCw2bg9x2_0;
	wire w_dff_A_oJswhKXS1_0;
	wire w_dff_A_lnHBadhK4_0;
	wire w_dff_A_eK7qKMgm7_0;
	wire w_dff_A_ON5FvVXy1_0;
	wire w_dff_A_gRqDjITU4_0;
	wire w_dff_A_9rkra2Mh0_0;
	wire w_dff_A_hwZxyIz79_0;
	wire w_dff_A_jE3CuK5s3_0;
	wire w_dff_A_r74hzztW8_0;
	wire w_dff_A_6Kr9jzom6_0;
	wire w_dff_A_Z4OIoiN49_0;
	wire w_dff_A_6ntirba20_0;
	wire w_dff_A_gAa2w9kM6_0;
	wire w_dff_A_awoxwtPU7_0;
	wire w_dff_A_GceHtWRX7_0;
	wire w_dff_A_q2X91lZv2_0;
	wire w_dff_A_9W89dofE4_0;
	wire w_dff_A_SzKoG7Nf0_0;
	wire w_dff_A_Vqyhnwny2_0;
	wire w_dff_A_x5mplucE6_0;
	wire w_dff_A_t6Eg007H0_0;
	wire w_dff_A_npW94Dfe7_0;
	wire w_dff_A_e8DteCl24_0;
	wire w_dff_A_nXOA6hWi9_0;
	wire w_dff_A_t2C4BIya5_0;
	wire w_dff_A_yd6bdb4p1_0;
	wire w_dff_A_5XalOgPE1_0;
	wire w_dff_A_gDU3XBye5_1;
	wire w_dff_A_XaqKY3Uv8_0;
	wire w_dff_A_HT7RyJrq9_0;
	wire w_dff_A_uKdcXXce1_0;
	wire w_dff_A_S55DiAsQ2_0;
	wire w_dff_A_14iiDsQQ6_0;
	wire w_dff_A_2ERLpZRJ8_0;
	wire w_dff_A_ZOuhXUfD9_0;
	wire w_dff_A_VPTkTMMH5_0;
	wire w_dff_A_bUiwIDly7_0;
	wire w_dff_A_KLJ1kaQ70_0;
	wire w_dff_A_ycUmO0n55_0;
	wire w_dff_A_c5ukUARk7_0;
	wire w_dff_A_p1RpYnfq1_0;
	wire w_dff_A_T0MSFy8n7_0;
	wire w_dff_A_5OZjwaVm4_0;
	wire w_dff_A_iQbagzNJ7_0;
	wire w_dff_A_Om19IT620_0;
	wire w_dff_A_GqV94TZb7_0;
	wire w_dff_A_C8BBNJca9_0;
	wire w_dff_A_DQPdZpQ47_0;
	wire w_dff_A_36kNi4lH9_0;
	wire w_dff_A_nrs4xXtW1_0;
	wire w_dff_A_RoCASpEY7_0;
	wire w_dff_A_N94buLv33_0;
	wire w_dff_A_iHESPorf3_0;
	wire w_dff_A_uwyn9o5o1_0;
	wire w_dff_A_BjG5g2wx7_0;
	wire w_dff_A_0UFCBU9A4_0;
	wire w_dff_A_dIPEFoYA6_0;
	wire w_dff_A_In1Y5C103_0;
	wire w_dff_A_sl6JrQzi9_0;
	wire w_dff_A_RKaIDixn2_0;
	wire w_dff_A_oi7ybY5V9_0;
	wire w_dff_A_Stah2Cq73_0;
	wire w_dff_A_1oAPG64a6_0;
	wire w_dff_A_GGRN8gwU6_0;
	wire w_dff_A_ocRhdTu39_0;
	wire w_dff_A_j5NQvppo7_0;
	wire w_dff_A_A1UvnyQh2_1;
	wire w_dff_A_juuvXi4i5_0;
	wire w_dff_A_r73q4xdv6_0;
	wire w_dff_A_aAZO6Nog0_0;
	wire w_dff_A_ER8IkTw92_0;
	wire w_dff_A_o4IQMRov5_0;
	wire w_dff_A_r3uHDbat4_0;
	wire w_dff_A_kRzEGgJu7_0;
	wire w_dff_A_qf4wB7cb9_0;
	wire w_dff_A_Y8vkjRUW5_0;
	wire w_dff_A_cXCYdfaI5_0;
	wire w_dff_A_i97WNmP72_0;
	wire w_dff_A_NC1IORo18_0;
	wire w_dff_A_8K3toON05_0;
	wire w_dff_A_VlbAE4hi5_0;
	wire w_dff_A_1ZcrHtIr3_0;
	wire w_dff_A_1C1ZgeCE3_0;
	wire w_dff_A_cPO6wbOn0_0;
	wire w_dff_A_wQdq0cQ51_0;
	wire w_dff_A_HecgiphY4_0;
	wire w_dff_A_F0iMQwZu7_0;
	wire w_dff_A_QKYiXZuG4_0;
	wire w_dff_A_kbNUKgLM4_0;
	wire w_dff_A_jQFjtW4i1_0;
	wire w_dff_A_tvsClI7Q6_0;
	wire w_dff_A_wG3InMlT3_0;
	wire w_dff_A_8jX9fUtF4_0;
	wire w_dff_A_tgINGoiR5_0;
	wire w_dff_A_aglNXVMK6_0;
	wire w_dff_A_YqUCq5HW9_0;
	wire w_dff_A_asljbY750_0;
	wire w_dff_A_m4NMEdVN7_0;
	wire w_dff_A_rQfQiJ3b0_0;
	wire w_dff_A_oxLrrY4h2_0;
	wire w_dff_A_2fnleoYj8_0;
	wire w_dff_A_QKaa79P86_0;
	wire w_dff_A_y6VYdPWv5_0;
	wire w_dff_A_F6Zd8z8H0_0;
	wire w_dff_A_7xpMx7Hg3_0;
	wire w_dff_A_ytKocOgQ9_2;
	wire w_dff_A_u5xFHdfj4_0;
	wire w_dff_A_WjhAFeTN3_0;
	wire w_dff_A_i0Qe0xZI2_0;
	wire w_dff_A_uu0dqjlh6_0;
	wire w_dff_A_MUSNqhkS9_0;
	wire w_dff_A_CdTwKHOO1_0;
	wire w_dff_A_zDHfvWjw4_0;
	wire w_dff_A_REomNbKK3_0;
	wire w_dff_A_1PiOxjdb9_0;
	wire w_dff_A_lVT4Lv2J2_0;
	wire w_dff_A_17kDSziH4_0;
	wire w_dff_A_PseaJE7S1_0;
	wire w_dff_A_kt8TGQsx6_0;
	wire w_dff_A_9VH95EMP3_0;
	wire w_dff_A_m7SZCh5R7_0;
	wire w_dff_A_HLy6FROn2_0;
	wire w_dff_A_vVOcTRRB1_0;
	wire w_dff_A_qxxy23fn0_0;
	wire w_dff_A_LUMijow94_0;
	wire w_dff_A_QcqMtWdv5_0;
	wire w_dff_A_BU6FsyXU0_0;
	wire w_dff_A_iYOqQ03s6_0;
	wire w_dff_A_F17JKdJi0_0;
	wire w_dff_A_zcTBT6Mo7_0;
	wire w_dff_A_aCEpFAws8_0;
	wire w_dff_A_hYJjWxaU4_0;
	wire w_dff_A_edeUIN8j2_0;
	wire w_dff_A_oRNrh9pK4_0;
	wire w_dff_A_ADmdLgf23_0;
	wire w_dff_A_SmSVMTgY7_0;
	wire w_dff_A_sgXfAoIJ8_0;
	wire w_dff_A_IfOjwXXJ5_0;
	wire w_dff_A_MZSXz5CL7_0;
	wire w_dff_A_nwL4j4is7_0;
	wire w_dff_A_NOAIjAV92_0;
	wire w_dff_A_i8ISFjqi3_0;
	wire w_dff_A_lap6QBdo1_0;
	wire w_dff_A_J1N7OnNX3_1;
	wire w_dff_A_cZlyu6Op5_0;
	wire w_dff_A_2iWyQBWE1_0;
	wire w_dff_A_WQuOi4cU9_0;
	wire w_dff_A_GYvyVxEJ1_0;
	wire w_dff_A_z4eYSgZB9_0;
	wire w_dff_A_G22fjfJg1_0;
	wire w_dff_A_0BtYIAYk7_0;
	wire w_dff_A_c0Qgxy8h0_0;
	wire w_dff_A_ZlbS6m6V5_0;
	wire w_dff_A_3fKf1FqW7_0;
	wire w_dff_A_m6vayyXN6_0;
	wire w_dff_A_zHOyvh6I5_0;
	wire w_dff_A_3xsB2VpR0_0;
	wire w_dff_A_F6GOwVeM8_0;
	wire w_dff_A_qFyn40Y37_0;
	wire w_dff_A_KheC66zi1_0;
	wire w_dff_A_FThAYanL2_0;
	wire w_dff_A_FxhLIXlx9_0;
	wire w_dff_A_kMh4pZ8s4_0;
	wire w_dff_A_xER7NfyN8_0;
	wire w_dff_A_6CAWJEE01_0;
	wire w_dff_A_1TxotZe58_0;
	wire w_dff_A_0vSiCIxz0_0;
	wire w_dff_A_ONIgy8xa7_0;
	wire w_dff_A_sAWWlxPQ1_0;
	wire w_dff_A_K6eae1RU0_0;
	wire w_dff_A_39OMQxVR5_0;
	wire w_dff_A_ryC3YZ0i3_0;
	wire w_dff_A_RcZpSoEr1_0;
	wire w_dff_A_Qj9Fo3y39_0;
	wire w_dff_A_I02JL7wp8_0;
	wire w_dff_A_XnvXlk3W7_0;
	wire w_dff_A_SBLRncLt0_0;
	wire w_dff_A_kGAyADmM3_0;
	wire w_dff_A_4JNmywKz3_0;
	wire w_dff_A_vKZYkuMo0_1;
	wire w_dff_A_y1wWVzf25_0;
	wire w_dff_A_xJ6PQyQB2_0;
	wire w_dff_A_9fONwAQG3_0;
	wire w_dff_A_NVCuZiQI8_0;
	wire w_dff_A_k0TrAN6J8_0;
	wire w_dff_A_BNaTlAM82_0;
	wire w_dff_A_L0AVxZpo7_0;
	wire w_dff_A_iqtFYjiF8_0;
	wire w_dff_A_gnHKDHsb3_0;
	wire w_dff_A_IjITfvdX3_0;
	wire w_dff_A_9zsa2Fmy4_0;
	wire w_dff_A_qLyNy7Xk7_0;
	wire w_dff_A_ADjBySD68_0;
	wire w_dff_A_P0c72Ign7_0;
	wire w_dff_A_y0rhxQyx4_0;
	wire w_dff_A_N1tgLf6D6_0;
	wire w_dff_A_D96EK0Sb7_0;
	wire w_dff_A_Jm0BlKwW1_0;
	wire w_dff_A_p335ytl93_0;
	wire w_dff_A_sOloWGCk6_0;
	wire w_dff_A_mIMorqH67_0;
	wire w_dff_A_HS6lVqRg9_0;
	wire w_dff_A_BHAdBjoz8_0;
	wire w_dff_A_w7EP3kX83_0;
	wire w_dff_A_efElcyDT8_0;
	wire w_dff_A_nBnFMORK2_0;
	wire w_dff_A_vAcffl565_0;
	wire w_dff_A_MnEcJrgw4_0;
	wire w_dff_A_iRZ7G1i57_0;
	wire w_dff_A_9JtKrjYg0_0;
	wire w_dff_A_4VhiGOsD6_0;
	wire w_dff_A_RkOevjGX8_0;
	wire w_dff_A_bX2iq0xp7_0;
	wire w_dff_A_Mm3jRJD58_0;
	wire w_dff_A_UO7Ui96n4_0;
	wire w_dff_A_pWywJuT40_1;
	wire w_dff_A_OmcSt8XA9_0;
	wire w_dff_A_G3whShqi9_0;
	wire w_dff_A_CZWnj7yt0_0;
	wire w_dff_A_WKcQ9D6q1_0;
	wire w_dff_A_SuqlomHn0_0;
	wire w_dff_A_52SSafLD6_0;
	wire w_dff_A_rhyFH44k0_0;
	wire w_dff_A_Jvz11xS98_0;
	wire w_dff_A_ohBE1dOx0_0;
	wire w_dff_A_YcrqZh111_0;
	wire w_dff_A_z2qtqzGQ5_0;
	wire w_dff_A_BYl4qxk40_0;
	wire w_dff_A_pNKDWu4z1_0;
	wire w_dff_A_J3a95Kom8_0;
	wire w_dff_A_EsWQiaez5_0;
	wire w_dff_A_fGLI1hom9_0;
	wire w_dff_A_lqZ1YNqm0_0;
	wire w_dff_A_aES1XdRl7_0;
	wire w_dff_A_XezniCnN2_0;
	wire w_dff_A_G1qFyNAM7_0;
	wire w_dff_A_77v2BGaR4_0;
	wire w_dff_A_imZMvE2Z6_0;
	wire w_dff_A_90aUtIOG5_0;
	wire w_dff_A_0v7KErAQ1_0;
	wire w_dff_A_nx3FjhIU3_0;
	wire w_dff_A_s9cDMHhc8_0;
	wire w_dff_A_hE3LesJc5_0;
	wire w_dff_A_VqfrfqeV1_0;
	wire w_dff_A_L7xPMk6m2_0;
	wire w_dff_A_oxMLrf1v5_0;
	wire w_dff_A_BNGkmhFq8_0;
	wire w_dff_A_LIqfwZBR1_0;
	wire w_dff_A_4Vgnq3KN2_0;
	wire w_dff_A_B2VwcZ5K1_0;
	wire w_dff_A_tswiLVgG9_0;
	wire w_dff_A_4rlRYtVI6_1;
	wire w_dff_A_lVJCs9ZF4_0;
	wire w_dff_A_BzvzbFi90_0;
	wire w_dff_A_8ApUZZPu5_0;
	wire w_dff_A_5p3tVPcr1_0;
	wire w_dff_A_9nnseZvV1_0;
	wire w_dff_A_J3LHzdNO5_0;
	wire w_dff_A_xUbCm4fK5_0;
	wire w_dff_A_FGV63dXO2_0;
	wire w_dff_A_3dJgQMh64_0;
	wire w_dff_A_V0NOh91S7_0;
	wire w_dff_A_9ujKsLdH3_0;
	wire w_dff_A_czrNmvtQ8_0;
	wire w_dff_A_kYBm0jpd5_0;
	wire w_dff_A_NNGpHLtA3_0;
	wire w_dff_A_NK0zeahi0_0;
	wire w_dff_A_vrxORiO87_0;
	wire w_dff_A_iRnrcSFN8_0;
	wire w_dff_A_vRfM4m8o0_0;
	wire w_dff_A_wWnhpshe5_0;
	wire w_dff_A_JzeHmLeB7_0;
	wire w_dff_A_6UzM0ipI4_0;
	wire w_dff_A_Z4IxsRvl0_0;
	wire w_dff_A_hemLPamn5_0;
	wire w_dff_A_K8mVxuH75_0;
	wire w_dff_A_RPtz7jam2_0;
	wire w_dff_A_hgm0GLFr8_0;
	wire w_dff_A_cEMixir65_0;
	wire w_dff_A_lHSRB4If0_0;
	wire w_dff_A_7DiyNd2U7_0;
	wire w_dff_A_NEKHCgtP6_0;
	wire w_dff_A_fJ9wCbnK3_0;
	wire w_dff_A_PBtBLRCE7_0;
	wire w_dff_A_2sK6pDFq1_0;
	wire w_dff_A_zKLxZxQ44_0;
	wire w_dff_A_jA7dYkxF0_0;
	wire w_dff_A_Vu8cR4Jp7_1;
	wire w_dff_A_5i8cpLHb5_0;
	wire w_dff_A_DMpA8Top1_0;
	wire w_dff_A_qwTR4BgR4_0;
	wire w_dff_A_dmW5sze64_0;
	wire w_dff_A_nyK44cbR3_0;
	wire w_dff_A_wStYp6HT4_0;
	wire w_dff_A_VaIU62lX1_0;
	wire w_dff_A_s3ZZiT9V0_0;
	wire w_dff_A_fcSOBhbo1_0;
	wire w_dff_A_64DurM4V4_0;
	wire w_dff_A_ZHpPe69W6_0;
	wire w_dff_A_jKtpQYMP9_0;
	wire w_dff_A_gPhuUl9e5_0;
	wire w_dff_A_rdnhWoVd3_0;
	wire w_dff_A_kaewQR4S1_0;
	wire w_dff_A_K3hv1RBr7_0;
	wire w_dff_A_VVggvK314_0;
	wire w_dff_A_TYQzpptT9_0;
	wire w_dff_A_5nTvMQDm1_0;
	wire w_dff_A_Rd1xvNJk0_0;
	wire w_dff_A_lpTnLFOU4_0;
	wire w_dff_A_Kdortbxs2_0;
	wire w_dff_A_jF6WUCVy7_0;
	wire w_dff_A_fknDQMDx4_0;
	wire w_dff_A_tmDtVvh60_0;
	wire w_dff_A_AP9pPwuU0_0;
	wire w_dff_A_qEDjwCFU2_0;
	wire w_dff_A_ZxQnCWNX0_0;
	wire w_dff_A_N3niM0mL6_0;
	wire w_dff_A_MESrp0w46_0;
	wire w_dff_A_VydHrt5f2_0;
	wire w_dff_A_KwPWcltU3_0;
	wire w_dff_A_O6iDQXGb4_0;
	wire w_dff_A_pK8l7x282_0;
	wire w_dff_A_oZ17SNP94_0;
	wire w_dff_A_3k3A0XI34_0;
	wire w_dff_A_B6U3A0sW5_0;
	wire w_dff_A_cUs6tElO5_0;
	wire w_dff_A_5vq1NzK46_1;
	wire w_dff_A_RWhZPeyn5_0;
	wire w_dff_A_69t1KPyU5_0;
	wire w_dff_A_oRLo3DGd9_0;
	wire w_dff_A_bG0dqtIO2_0;
	wire w_dff_A_4d62k3gL4_0;
	wire w_dff_A_AqzIaTTa0_0;
	wire w_dff_A_LrVSuCY69_0;
	wire w_dff_A_ZTk8f71O4_0;
	wire w_dff_A_DzSrgD5D8_0;
	wire w_dff_A_J5bLCuQa5_0;
	wire w_dff_A_HKjWBDn83_0;
	wire w_dff_A_kyJOby1d8_0;
	wire w_dff_A_EtL645nO0_0;
	wire w_dff_A_R05f0I603_0;
	wire w_dff_A_lNBHcHsV8_0;
	wire w_dff_A_nfPGEAUK3_0;
	wire w_dff_A_PNtiR7ui6_0;
	wire w_dff_A_4w1V4leJ9_0;
	wire w_dff_A_xTQhv5cJ1_0;
	wire w_dff_A_d9pzY2252_0;
	wire w_dff_A_ZXUZEbvX1_0;
	wire w_dff_A_tFuMzwrz1_0;
	wire w_dff_A_fnFz8lJJ6_0;
	wire w_dff_A_YX0uaIbB1_0;
	wire w_dff_A_cE95QgSE5_0;
	wire w_dff_A_ATLcBc094_0;
	wire w_dff_A_OyHI66Sc8_0;
	wire w_dff_A_v9n2gnZu9_0;
	wire w_dff_A_3HL1oRR98_0;
	wire w_dff_A_RBvs5vBl3_0;
	wire w_dff_A_9UTDv1vd6_0;
	wire w_dff_A_BWBcdv017_0;
	wire w_dff_A_eyrzJ9co8_0;
	wire w_dff_A_HUPnCAvo6_0;
	wire w_dff_A_Q1owd4z01_0;
	wire w_dff_A_N90zrYVj4_0;
	wire w_dff_A_xgtMHEqH5_0;
	wire w_dff_A_7DFVRbGw8_0;
	wire w_dff_A_wmykSRR86_2;
	wire w_dff_A_Z51GU5HB7_0;
	wire w_dff_A_zGrKeZqZ5_0;
	wire w_dff_A_PXuxDnnM5_0;
	wire w_dff_A_ol68DJzv4_0;
	wire w_dff_A_AOORy8nP5_0;
	wire w_dff_A_XCwxvokX3_0;
	wire w_dff_A_F6HjEGE46_0;
	wire w_dff_A_5lelyWJW0_0;
	wire w_dff_A_YIzQye5Q8_0;
	wire w_dff_A_imD8Z55Y9_0;
	wire w_dff_A_OHJsVG1g2_0;
	wire w_dff_A_GHJmHHPj3_0;
	wire w_dff_A_WpU0gC1M2_0;
	wire w_dff_A_C3w5BKHM3_0;
	wire w_dff_A_WhEpmYTP2_0;
	wire w_dff_A_T97Vuu3R3_0;
	wire w_dff_A_GRGcX3AD1_0;
	wire w_dff_A_8A0qKjGt6_0;
	wire w_dff_A_Vkh5GnhK1_0;
	wire w_dff_A_5B6xlWj57_0;
	wire w_dff_A_Dx3Vfwf22_0;
	wire w_dff_A_MZjFnhSg8_0;
	wire w_dff_A_gtXoUYHa9_0;
	wire w_dff_A_fS6QIagt1_0;
	wire w_dff_A_VjFsIsaQ0_0;
	wire w_dff_A_uRNgKGz43_0;
	wire w_dff_A_lggBUf2K4_0;
	wire w_dff_A_eGhgYgQh1_0;
	wire w_dff_A_Ffwg5ycn5_0;
	wire w_dff_A_3F30JImT4_0;
	wire w_dff_A_VUe7KyNH7_0;
	wire w_dff_A_7TtxzLVg4_0;
	wire w_dff_A_cus4gAfG4_0;
	wire w_dff_A_WQRpURD65_0;
	wire w_dff_A_lyW3cX1Q4_0;
	wire w_dff_A_Kr8Zppao6_0;
	wire w_dff_A_LK3Lj7IW8_1;
	wire w_dff_A_vv713Bvq1_0;
	wire w_dff_A_zEbL5uDi0_0;
	wire w_dff_A_SQp6LKnd4_0;
	wire w_dff_A_PQYNnWu59_0;
	wire w_dff_A_ZyBpAdI46_0;
	wire w_dff_A_YTqWs3Sx5_0;
	wire w_dff_A_Nyh6K99J5_0;
	wire w_dff_A_vbwYQ40B2_0;
	wire w_dff_A_fm3Ygbhl8_0;
	wire w_dff_A_nGFsQlsp1_0;
	wire w_dff_A_0EKOTzA42_0;
	wire w_dff_A_D2xOMZRz9_0;
	wire w_dff_A_KgnTolMr3_0;
	wire w_dff_A_lJp42sc29_0;
	wire w_dff_A_ghXbvJ1f8_0;
	wire w_dff_A_uy9TUzlO2_0;
	wire w_dff_A_2hZ8ETyn4_0;
	wire w_dff_A_7jQfeHko0_0;
	wire w_dff_A_A8HAJWnj9_0;
	wire w_dff_A_HVcHDPwV4_0;
	wire w_dff_A_SMhDs7gf6_0;
	wire w_dff_A_af1a85sD4_0;
	wire w_dff_A_fqstAJLj5_0;
	wire w_dff_A_bJdLdHTK8_0;
	wire w_dff_A_3tPXQOIt0_0;
	wire w_dff_A_UJc8fYiZ0_0;
	wire w_dff_A_TERPNisl1_0;
	wire w_dff_A_8RV9zaeB0_0;
	wire w_dff_A_Fq8lh1uI3_0;
	wire w_dff_A_PLbobi7e6_0;
	wire w_dff_A_gAWdG71D4_0;
	wire w_dff_A_YQMTkIYH3_0;
	wire w_dff_A_x8BFfMcg6_0;
	wire w_dff_A_c0YvDkVh3_0;
	wire w_dff_A_bZSNPdQs8_0;
	wire w_dff_A_xcQwQ9SM8_0;
	wire w_dff_A_m9WXrRFw4_0;
	wire w_dff_A_Zda8mllT3_2;
	wire w_dff_A_ANWSoPVe0_0;
	wire w_dff_A_ENPSlR9V8_0;
	wire w_dff_A_tr6UedhH1_0;
	wire w_dff_A_o2mxWgGN3_0;
	wire w_dff_A_fPCIrz2y1_0;
	wire w_dff_A_DZkV7ReE7_0;
	wire w_dff_A_S5GL391M7_0;
	wire w_dff_A_wlig9YlB9_0;
	wire w_dff_A_c84YCPeC5_0;
	wire w_dff_A_kT4Seda37_0;
	wire w_dff_A_feMNgSdp0_0;
	wire w_dff_A_I0Tdke2j5_0;
	wire w_dff_A_CT9V92q39_0;
	wire w_dff_A_rWJd1lxd0_0;
	wire w_dff_A_xmgpYhAA6_0;
	wire w_dff_A_ysMsFMnY4_0;
	wire w_dff_A_CxL67Ksl0_0;
	wire w_dff_A_GXVuplTV8_0;
	wire w_dff_A_rlfxZZjm3_0;
	wire w_dff_A_HR6Im4lF0_0;
	wire w_dff_A_GTRhtGmT5_0;
	wire w_dff_A_9sztd85p7_0;
	wire w_dff_A_bDzlcFXt1_0;
	wire w_dff_A_mpb3HOcT8_0;
	wire w_dff_A_B7fRJPiM1_0;
	wire w_dff_A_olsAFkr41_0;
	wire w_dff_A_u7o8P4pA6_0;
	wire w_dff_A_LEKUdH8H6_0;
	wire w_dff_A_VjIfLl0q2_0;
	wire w_dff_A_AtfvshBG0_0;
	wire w_dff_A_yVvlo2nG3_0;
	wire w_dff_A_amVJRz0l2_0;
	wire w_dff_A_kgUi1bYH3_0;
	wire w_dff_A_VkzLy2zk9_0;
	wire w_dff_A_1Q23ub1H0_0;
	wire w_dff_A_9KmSwSEi9_0;
	wire w_dff_A_D8xH8Oi22_2;
	wire w_dff_A_QeaqzpoA3_0;
	wire w_dff_A_UlKbVGnf9_0;
	wire w_dff_A_RUH0X1aq1_0;
	wire w_dff_A_LTjQI9qp2_0;
	wire w_dff_A_EFgoXyTb1_0;
	wire w_dff_A_TQYILxmN6_0;
	wire w_dff_A_EV6b3my62_0;
	wire w_dff_A_c4hGrQpA7_0;
	wire w_dff_A_wrxJuxDE4_0;
	wire w_dff_A_16Mm9h3l1_0;
	wire w_dff_A_I8wEl9ob2_0;
	wire w_dff_A_1wzQhIEN6_0;
	wire w_dff_A_Xqd6tnkC1_0;
	wire w_dff_A_RLLruLqB2_0;
	wire w_dff_A_nJtGxlW45_0;
	wire w_dff_A_J17VpB8y7_0;
	wire w_dff_A_3KaJR61b6_0;
	wire w_dff_A_ImVMVU8X4_0;
	wire w_dff_A_UvYnuncs2_0;
	wire w_dff_A_FmvigApb9_0;
	wire w_dff_A_JoVMRdbh2_0;
	wire w_dff_A_NsS6ZsxL4_0;
	wire w_dff_A_GQLbrFlD0_0;
	wire w_dff_A_tFinVVOt8_0;
	wire w_dff_A_qsDEeN3N2_0;
	wire w_dff_A_7tya0M0h9_0;
	wire w_dff_A_hwszIDsf6_0;
	wire w_dff_A_NKkSuLOP3_0;
	wire w_dff_A_lKQqMRGc9_0;
	wire w_dff_A_1yF2FMkm4_0;
	wire w_dff_A_UEzsUctU8_0;
	wire w_dff_A_fgRZTT0e8_0;
	wire w_dff_A_hvkTvSRV7_0;
	wire w_dff_A_guDGb1dG0_0;
	wire w_dff_A_2lOuxi4F3_0;
	wire w_dff_A_GbPQfCGT0_1;
	wire w_dff_A_irDydLFs4_0;
	wire w_dff_A_cDmpTu5Y2_0;
	wire w_dff_A_kNrv0VxV9_0;
	wire w_dff_A_tWLpSJRW1_0;
	wire w_dff_A_u55keSlm9_0;
	wire w_dff_A_Q8wsBj6h9_0;
	wire w_dff_A_tplCoRQI2_0;
	wire w_dff_A_I7o8meEr5_0;
	wire w_dff_A_TLkILGK99_0;
	wire w_dff_A_J2LBPLHi3_0;
	wire w_dff_A_Rf6o4KNF3_0;
	wire w_dff_A_LV1LWeau9_0;
	wire w_dff_A_bamJNO4J8_0;
	wire w_dff_A_Dk3ozH7T4_0;
	wire w_dff_A_gbygC4fj8_0;
	wire w_dff_A_qtCeMX6g6_0;
	wire w_dff_A_3lANmBzG1_0;
	wire w_dff_A_Hp2aH8Te5_0;
	wire w_dff_A_5EEAs0TA0_0;
	wire w_dff_A_vQZG6WeP3_0;
	wire w_dff_A_53xjXXvi9_0;
	wire w_dff_A_DTKax7gg9_0;
	wire w_dff_A_1bQCAe5l2_0;
	wire w_dff_A_ad9ZMT4Z0_0;
	wire w_dff_A_H6MSNFsM6_0;
	wire w_dff_A_SdmCZUZD1_0;
	wire w_dff_A_1N1Kpv939_0;
	wire w_dff_A_qUdhMDYJ4_0;
	wire w_dff_A_HCAzTAlZ3_0;
	wire w_dff_A_lsPXM3Wn5_0;
	wire w_dff_A_e0E61vYZ3_0;
	wire w_dff_A_ApsbvxKn4_0;
	wire w_dff_A_pnoAOqv47_0;
	wire w_dff_A_QMTuUWtV1_0;
	wire w_dff_A_SnxHDgde9_0;
	wire w_dff_A_c9brB2b12_0;
	wire w_dff_A_f2PAfZVx0_0;
	wire w_dff_A_9eF0pr3b7_2;
	wire w_dff_A_U5aihzHX7_0;
	wire w_dff_A_Ebt2Dh5G4_0;
	wire w_dff_A_UOIeNXiL8_0;
	wire w_dff_A_igtWn4hb3_0;
	wire w_dff_A_U5APrh1d1_0;
	wire w_dff_A_vP9pbXTf6_0;
	wire w_dff_A_dHhyIdd24_0;
	wire w_dff_A_57JAJ3C18_0;
	wire w_dff_A_WK4SPcEo0_0;
	wire w_dff_A_fMxxyZX77_0;
	wire w_dff_A_YqKXUNoP6_0;
	wire w_dff_A_alhtDkAp7_0;
	wire w_dff_A_F3hDwAHE7_0;
	wire w_dff_A_AhqxXLdX3_0;
	wire w_dff_A_m9g9MC1d9_0;
	wire w_dff_A_pj3aacqR7_0;
	wire w_dff_A_aghY5Z0G6_0;
	wire w_dff_A_ylHZq5le6_0;
	wire w_dff_A_Jl4jzpA91_0;
	wire w_dff_A_K7RRo5073_0;
	wire w_dff_A_ETH7nLvz9_0;
	wire w_dff_A_yWt2LeYO8_0;
	wire w_dff_A_HBWfBKkJ9_0;
	wire w_dff_A_Y2KUgy323_0;
	wire w_dff_A_y9BS71jB9_0;
	wire w_dff_A_KJ5YL3Fu2_0;
	wire w_dff_A_esaUVrAh2_0;
	wire w_dff_A_ozpON0Wj9_0;
	wire w_dff_A_H5pdPkaq8_0;
	wire w_dff_A_s8gxRBU05_0;
	wire w_dff_A_0XLYwrdL8_0;
	wire w_dff_A_CF594JrW0_0;
	wire w_dff_A_Z2hBtZLw1_0;
	wire w_dff_A_IWgvaZ752_0;
	wire w_dff_A_4HyqLyIS7_0;
	wire w_dff_A_VajKcQKi2_1;
	wire w_dff_A_iGg4Nv891_0;
	wire w_dff_A_25goQeuA9_0;
	wire w_dff_A_HatPLPWP1_0;
	wire w_dff_A_qzThAfp04_0;
	wire w_dff_A_AhGh7UAO2_0;
	wire w_dff_A_ibjJ9Hns4_0;
	wire w_dff_A_BCoYnTiM9_0;
	wire w_dff_A_26Aud73p7_0;
	wire w_dff_A_TfnDFASo2_0;
	wire w_dff_A_v2o9LzU17_0;
	wire w_dff_A_N9P4dUAr8_0;
	wire w_dff_A_tGlkqVm22_0;
	wire w_dff_A_VjHpNReM8_0;
	wire w_dff_A_2j0VGHDN6_0;
	wire w_dff_A_IzYZAoVZ8_0;
	wire w_dff_A_0nnwbXVY7_0;
	wire w_dff_A_KEowFla87_0;
	wire w_dff_A_Tpchak8d5_0;
	wire w_dff_A_av91L8Q51_0;
	wire w_dff_A_SZXiAgwB9_0;
	wire w_dff_A_eucxQIuR4_0;
	wire w_dff_A_uMrkjlE98_0;
	wire w_dff_A_PZEL2WM43_0;
	wire w_dff_A_eko1wODP7_0;
	wire w_dff_A_KAN9EA0y5_0;
	wire w_dff_A_Bv3P9Ohy5_0;
	wire w_dff_A_7viZ92165_0;
	wire w_dff_A_vXMDM2cu8_0;
	wire w_dff_A_ij20ieMK5_0;
	wire w_dff_A_QygmYoyv5_0;
	wire w_dff_A_bL4S26bH5_0;
	wire w_dff_A_Cg2zNbpT6_0;
	wire w_dff_A_FGeTxGOj4_0;
	wire w_dff_A_OPflZcUf0_0;
	wire w_dff_A_pCjmLV2F7_0;
	wire w_dff_A_RYBntYTO7_0;
	wire w_dff_A_3y7xPflI7_0;
	wire w_dff_A_iliYjplN9_0;
	wire w_dff_A_yJxiPeRD1_2;
	wire w_dff_A_iHVGdYtC5_0;
	wire w_dff_A_Z8YN3F5L8_0;
	wire w_dff_A_rGU61j2x4_0;
	wire w_dff_A_EUtMwiv20_0;
	wire w_dff_A_JK7lKOAd9_0;
	wire w_dff_A_u0WiDjz06_0;
	wire w_dff_A_fGrgpTCd4_0;
	wire w_dff_A_cMg4yR6h7_0;
	wire w_dff_A_VcRvXCnt1_0;
	wire w_dff_A_ppGeXKRj7_0;
	wire w_dff_A_uUrkPgJd2_0;
	wire w_dff_A_gwWwRlz55_0;
	wire w_dff_A_8885U0Yd4_0;
	wire w_dff_A_z6AFslYN4_0;
	wire w_dff_A_HAPUPDnJ5_0;
	wire w_dff_A_ifnRkYcn9_0;
	wire w_dff_A_PUCYaq8L6_0;
	wire w_dff_A_q5YU6Sbn5_0;
	wire w_dff_A_bojcxAPn8_0;
	wire w_dff_A_fnS28SFh7_0;
	wire w_dff_A_fK8fBM9u7_0;
	wire w_dff_A_xW1zuY2b6_0;
	wire w_dff_A_4oh8RdhF9_0;
	wire w_dff_A_E2dOlFAB5_0;
	wire w_dff_A_5eKDupkb3_0;
	wire w_dff_A_L0tboVp27_0;
	wire w_dff_A_0aDugl4U4_0;
	wire w_dff_A_qlUrri2u5_0;
	wire w_dff_A_ZrAVO2IU7_0;
	wire w_dff_A_4LD1nPrA5_0;
	wire w_dff_A_MlgP1iY98_0;
	wire w_dff_A_fvKcz1on6_0;
	wire w_dff_A_9iFHD7mZ9_0;
	wire w_dff_A_W9gYILl37_0;
	wire w_dff_A_kviH5ehM8_0;
	wire w_dff_A_kp2e2jZt0_0;
	wire w_dff_A_MC5uGbXK2_0;
	wire w_dff_A_62FaZpmK6_2;
	wire w_dff_A_g69OA2CD8_0;
	wire w_dff_A_QuiRtBwq1_0;
	wire w_dff_A_TlIzQDNG4_0;
	wire w_dff_A_Z7FljO0j8_0;
	wire w_dff_A_1jhYuCaq9_0;
	wire w_dff_A_a04esJpm8_0;
	wire w_dff_A_wf0HrOHu5_0;
	wire w_dff_A_p28Vpuyy9_0;
	wire w_dff_A_aRu70x720_0;
	wire w_dff_A_Y0bK5UJ64_0;
	wire w_dff_A_LFn6pe3n6_0;
	wire w_dff_A_sutW7no98_0;
	wire w_dff_A_lmvuzq220_0;
	wire w_dff_A_KCalkvOR0_0;
	wire w_dff_A_Tmn7GQBH2_0;
	wire w_dff_A_BvtVsQ6g7_0;
	wire w_dff_A_hWK0YZrx1_0;
	wire w_dff_A_xOLgtix93_0;
	wire w_dff_A_EkoUja323_0;
	wire w_dff_A_hZjZiFLp0_0;
	wire w_dff_A_rccexe282_0;
	wire w_dff_A_tSTR4kib9_0;
	wire w_dff_A_taBGw0sO5_0;
	wire w_dff_A_LFuVQOqR2_0;
	wire w_dff_A_99dDVmuY5_0;
	wire w_dff_A_cUEa9D5Z8_0;
	wire w_dff_A_46SttGKm0_0;
	wire w_dff_A_38FWKvTq4_0;
	wire w_dff_A_XYDVWFAH6_0;
	wire w_dff_A_scyCPkrx4_0;
	wire w_dff_A_Wiugym454_0;
	wire w_dff_A_fDL61mJj8_0;
	wire w_dff_A_ajNjXzv73_2;
	wire w_dff_A_TT4aLrxh8_0;
	wire w_dff_A_b0mGOHEG0_0;
	wire w_dff_A_OnzrlcE83_0;
	wire w_dff_A_Ni1LBTDx6_0;
	wire w_dff_A_51H5h98E4_0;
	wire w_dff_A_IQtwMLvQ3_0;
	wire w_dff_A_AT6yNBzT9_0;
	wire w_dff_A_YHG8H1Bh1_0;
	wire w_dff_A_3hIjCyoX8_0;
	wire w_dff_A_AVEnn40H0_0;
	wire w_dff_A_Q0KcgJhF3_2;
	wire w_dff_A_KOl0W78C0_0;
	wire w_dff_A_Z3KaIGIt9_0;
	wire w_dff_A_kh0fWH8s9_0;
	wire w_dff_A_RIu0V3s05_0;
	wire w_dff_A_L2FBgBar5_0;
	wire w_dff_A_os08S9Zl1_0;
	wire w_dff_A_s9YsBpMv2_0;
	wire w_dff_A_nrhjltUI8_0;
	wire w_dff_A_ZpScyhoT6_0;
	wire w_dff_A_Mdo2LnXM0_0;
	wire w_dff_A_x51Q2GgN5_2;
	wire w_dff_A_QXfTuB9g2_0;
	wire w_dff_A_8AmfZoAq5_0;
	wire w_dff_A_IbzWtfJ57_0;
	wire w_dff_A_nQDqItJ52_0;
	wire w_dff_A_1A2juYv22_0;
	wire w_dff_A_7kVhfNGW5_0;
	wire w_dff_A_4FGNoSC30_0;
	wire w_dff_A_XsqEqve71_0;
	wire w_dff_A_6XKQXWdV0_0;
	wire w_dff_A_axiQnByq7_0;
	wire w_dff_A_1zmDcDJv6_0;
	wire w_dff_A_2JzmCsOe5_0;
	wire w_dff_A_m5nnqRn43_0;
	wire w_dff_A_bZxY0xT66_0;
	wire w_dff_A_HtTAx8rO5_0;
	wire w_dff_A_PobgbFdN5_0;
	wire w_dff_A_1D3r5Csv8_0;
	wire w_dff_A_zP4AdlFR4_0;
	wire w_dff_A_R5K8hbGX9_0;
	wire w_dff_A_YzPpywWF1_0;
	wire w_dff_A_IqpCznLV2_0;
	wire w_dff_A_74miDqLV3_0;
	wire w_dff_A_cnOsFqtO4_0;
	wire w_dff_A_w1xkvhtt2_0;
	wire w_dff_A_tgXJYLwI4_2;
	wire w_dff_A_e8n7Ar3U3_0;
	wire w_dff_A_wv5xUv0L1_0;
	wire w_dff_A_shkJdoO66_0;
	wire w_dff_A_lDZ4pdgI4_0;
	wire w_dff_A_e8Lf7LST4_0;
	wire w_dff_A_TTlPoZiz7_0;
	wire w_dff_A_8DBmWNwx2_0;
	wire w_dff_A_QYoWCk942_0;
	wire w_dff_A_qwXBWzUf1_0;
	wire w_dff_A_J92Njuev3_0;
	wire w_dff_A_lF18xUBi2_0;
	wire w_dff_A_PbYKugJO5_0;
	wire w_dff_A_MFIzeAoe9_0;
	wire w_dff_A_zTlAwahR5_0;
	wire w_dff_A_Cjn9rNU64_0;
	wire w_dff_A_WR4UX0mG1_0;
	wire w_dff_A_SjN8FEkV4_0;
	wire w_dff_A_nVanINLU6_0;
	wire w_dff_A_KdBdRfhE9_0;
	wire w_dff_A_64vzetlD5_0;
	wire w_dff_A_KB6jdD1o0_0;
	wire w_dff_A_gyCzG5ON0_0;
	wire w_dff_A_Vn7EchJy1_0;
	wire w_dff_A_AZGuGxhX2_0;
	wire w_dff_A_4NLTdJkF2_0;
	wire w_dff_A_zOyK1N2d6_0;
	wire w_dff_A_hkO5sPZ89_2;
	wire w_dff_A_hDf1sSif9_0;
	wire w_dff_A_FKu6O3aV5_0;
	wire w_dff_A_rcWQz1U65_0;
	wire w_dff_A_uFpE2Po36_0;
	wire w_dff_A_keeOhkK75_0;
	wire w_dff_A_MsShcQ7S4_0;
	wire w_dff_A_oNjxtp9A8_0;
	wire w_dff_A_rC0muEOt1_0;
	wire w_dff_A_erigIFGs7_0;
	wire w_dff_A_8NSbKSdI9_0;
	wire w_dff_A_IR4XtSOk8_0;
	wire w_dff_A_y9o18sIB9_0;
	wire w_dff_A_TEolZjW42_0;
	wire w_dff_A_DqLLjM5I8_0;
	wire w_dff_A_EIhcovon5_0;
	wire w_dff_A_XqDFxfmS0_0;
	wire w_dff_A_fxpMamxY8_0;
	wire w_dff_A_2lMCaGUg2_0;
	wire w_dff_A_B7BVzTId6_0;
	wire w_dff_A_9Hiq8nFQ8_0;
	wire w_dff_A_M2FgQ2rq9_0;
	wire w_dff_A_dEMzwWWl4_0;
	wire w_dff_A_G2oBSjtg8_0;
	wire w_dff_A_8LK18O1Z3_0;
	wire w_dff_A_LQJK2jlo1_0;
	wire w_dff_A_MA2zVwB88_0;
	wire w_dff_A_4vkxo6Gj6_0;
	wire w_dff_A_8RB6P5rK6_0;
	wire w_dff_A_aT2yF8k26_0;
	wire w_dff_A_pvUyVpXg5_2;
	wire w_dff_A_aQnNbj4A1_0;
	wire w_dff_A_GM2XjGwi6_0;
	wire w_dff_A_afYCStxr6_0;
	wire w_dff_A_ArzSCmgO4_0;
	wire w_dff_A_ANBeOubi5_0;
	wire w_dff_A_PirPFoVG9_0;
	wire w_dff_A_6Km1af7F4_0;
	wire w_dff_A_1AOz8bgR5_0;
	wire w_dff_A_TQyB4yGi6_0;
	wire w_dff_A_JPi4u3Gg9_0;
	wire w_dff_A_XgAjAylE0_0;
	wire w_dff_A_R8HW4Iw66_0;
	wire w_dff_A_AMDfN9IF8_0;
	wire w_dff_A_bG1X534F1_0;
	wire w_dff_A_Olh0tCaK3_0;
	wire w_dff_A_ICOjzVrE7_0;
	wire w_dff_A_V4d4Pfi78_0;
	wire w_dff_A_U9Mlowu36_0;
	wire w_dff_A_o7ACEmcQ1_0;
	wire w_dff_A_ByUSFJiO5_0;
	wire w_dff_A_cEuF0Rzi9_0;
	wire w_dff_A_9957mxCD8_0;
	wire w_dff_A_HFWFTiPj0_0;
	wire w_dff_A_HlwiP6gc5_0;
	wire w_dff_A_5oN3giQS6_0;
	wire w_dff_A_K0kl6G7I1_0;
	wire w_dff_A_Y37qaQCu8_0;
	wire w_dff_A_GWYdknZy7_0;
	wire w_dff_A_CoNVsJtZ1_0;
	wire w_dff_A_663F91Cz0_0;
	wire w_dff_A_GuechTS56_2;
	wire w_dff_A_DreT6W6u5_0;
	wire w_dff_A_YOm0inDL0_0;
	wire w_dff_A_e4jPZs2m6_0;
	wire w_dff_A_Vr572Rtv1_0;
	wire w_dff_A_DOUAVlbY7_0;
	wire w_dff_A_FcKAJZuq1_0;
	wire w_dff_A_fJ3zIYMN2_0;
	wire w_dff_A_6S90kLS13_0;
	wire w_dff_A_kdPz2qcZ8_0;
	wire w_dff_A_Vm79z5F93_0;
	wire w_dff_A_AWdaB3Ec6_0;
	wire w_dff_A_zaIDG96W8_0;
	wire w_dff_A_gZJ7ln329_0;
	wire w_dff_A_KUkinsFk0_0;
	wire w_dff_A_Ype3lJny5_0;
	wire w_dff_A_C3XdZN2U6_0;
	wire w_dff_A_Z9f3GqZY4_0;
	wire w_dff_A_VhDx769O3_0;
	wire w_dff_A_l23cfTzy2_0;
	wire w_dff_A_ZvFxzFFl6_2;
	wire w_dff_A_yl4c68K17_0;
	wire w_dff_A_BWACLAwZ7_0;
	wire w_dff_A_pYW6OGzw3_0;
	wire w_dff_A_HByCGAtg4_0;
	wire w_dff_A_7yPhfK087_0;
	wire w_dff_A_nzCs7fQd0_0;
	wire w_dff_A_mM4BEOBM8_0;
	wire w_dff_A_vW1ke1cG7_0;
	wire w_dff_A_rGreo9cd6_0;
	wire w_dff_A_eJJTBJwz2_0;
	wire w_dff_A_6YfKyfQg2_0;
	wire w_dff_A_eMGdGFOn4_0;
	wire w_dff_A_x134uNko5_0;
	wire w_dff_A_nU6I5wxd2_0;
	wire w_dff_A_l6yd9qmU7_0;
	wire w_dff_A_EcGTPUBE1_0;
	wire w_dff_A_1kgivv1n3_0;
	wire w_dff_A_H0wMBfXf4_0;
	wire w_dff_A_dEMtNCfJ5_0;
	wire w_dff_A_zKLkmPlr7_0;
	wire w_dff_A_YqoFysBa9_0;
	wire w_dff_A_5w4VshfQ8_2;
	wire w_dff_A_q7n93WK18_0;
	wire w_dff_A_lvbsOgSD4_0;
	wire w_dff_A_wFHhGfu92_0;
	wire w_dff_A_Tu5a0fAV7_0;
	wire w_dff_A_3St9h9bx2_0;
	wire w_dff_A_NyrB6F5Q5_0;
	wire w_dff_A_0f8N24lP9_0;
	wire w_dff_A_b621w5zO5_0;
	wire w_dff_A_XRs9b6JG2_0;
	wire w_dff_A_TjQF7fUR9_0;
	wire w_dff_A_mY6ane3F4_0;
	wire w_dff_A_fxNW82Go9_0;
	wire w_dff_A_DFuXy87B4_0;
	wire w_dff_A_O5b2Z5p05_0;
	wire w_dff_A_VrUYWFm31_0;
	wire w_dff_A_imV7IoPg4_0;
	wire w_dff_A_Wb9TkMDO0_0;
	wire w_dff_A_6Lsfjqr59_0;
	wire w_dff_A_8wj6Wm7R1_0;
	wire w_dff_A_vdQfoMTJ6_0;
	wire w_dff_A_kL0ot33z2_0;
	wire w_dff_A_DUPrbXiE4_2;
	wire w_dff_A_2ivTuG0o4_0;
	wire w_dff_A_Quh7QA6X1_0;
	wire w_dff_A_4yJtbFSK1_0;
	wire w_dff_A_N5r2sCJW6_0;
	wire w_dff_A_41HNgVQJ9_0;
	wire w_dff_A_ZiYWAXPU8_0;
	wire w_dff_A_khwVr4Ex7_0;
	wire w_dff_A_B0hqfcLv2_0;
	wire w_dff_A_oNali3mg7_0;
	wire w_dff_A_DgZ3Dx7Y1_0;
	wire w_dff_A_7KBxL5iM3_0;
	wire w_dff_A_wm5El60a6_0;
	wire w_dff_A_EfTPYhTn4_0;
	wire w_dff_A_zxSMasvo1_0;
	wire w_dff_A_hZVaN7bZ1_0;
	wire w_dff_A_ulTVmNjv0_0;
	wire w_dff_A_ZhR5ERnX7_0;
	wire w_dff_A_UiJ7KuGz5_0;
	wire w_dff_A_1LaUYo8R6_0;
	wire w_dff_A_I61dxXyN6_0;
	wire w_dff_A_mtaQzUXW4_0;
	wire w_dff_A_lLR2aZWF8_0;
	wire w_dff_A_uEdtUAss8_0;
	wire w_dff_A_CNbvXIlX4_1;
	wire w_dff_A_8LJshTeN7_0;
	wire w_dff_A_cmvwVrDb7_0;
	wire w_dff_A_7D5mA9my9_0;
	wire w_dff_A_C5C6CeiH3_0;
	wire w_dff_A_vmR9uS2j2_0;
	wire w_dff_A_NRrrW3Nn8_0;
	wire w_dff_A_Gixi2GFr1_0;
	wire w_dff_A_BLTyQRrj2_0;
	wire w_dff_A_L4MvBRI58_0;
	wire w_dff_A_NoZQupbt3_0;
	wire w_dff_A_WfXEtKLE8_0;
	wire w_dff_A_rClWGEqo3_0;
	wire w_dff_A_ZjEpd6U45_0;
	wire w_dff_A_voZF0aPA0_0;
	wire w_dff_A_MJm2m4Ol4_0;
	wire w_dff_A_IXPfjlOj1_0;
	wire w_dff_A_bJTur37y6_0;
	wire w_dff_A_Gv9xqr5e8_0;
	wire w_dff_A_T6kEokzt6_0;
	wire w_dff_A_Sj8e0U7L1_0;
	wire w_dff_A_bFkTP5Xb4_0;
	wire w_dff_A_EOVDFatY7_0;
	wire w_dff_A_lMf3jntd4_0;
	wire w_dff_A_JTfPbw8A4_0;
	wire w_dff_A_w0Bp0l8X8_0;
	wire w_dff_A_ZhHw2eDs6_0;
	wire w_dff_A_CbgiTCht4_0;
	wire w_dff_A_UmDLHC9r2_1;
	wire w_dff_A_fpzQTFJ88_0;
	wire w_dff_A_apvPFEcu1_0;
	wire w_dff_A_NKZ9uYqh1_0;
	wire w_dff_A_tb2fT9FA9_0;
	wire w_dff_A_cS7YiuoZ3_0;
	wire w_dff_A_2djp1TUH2_0;
	wire w_dff_A_54QTNkBY3_0;
	wire w_dff_A_PHxgHErl7_0;
	wire w_dff_A_TTVQ65Tf8_0;
	wire w_dff_A_6Tm1qKK22_0;
	wire w_dff_A_gRYMJjOw4_0;
	wire w_dff_A_JhLcErlz3_0;
	wire w_dff_A_S8VLBB1r3_0;
	wire w_dff_A_1MEE1oU61_0;
	wire w_dff_A_Xq4Wyqyy4_0;
	wire w_dff_A_yue0ZhoI1_0;
	wire w_dff_A_eNDQTfor1_0;
	wire w_dff_A_jACVARD91_0;
	wire w_dff_A_ZEp5Uszh1_0;
	wire w_dff_A_SseCrQIB5_0;
	wire w_dff_A_9lLQRbp46_0;
	wire w_dff_A_L5Jy556h1_0;
	wire w_dff_A_3nug4nro5_0;
	wire w_dff_A_yRGTWnt00_0;
	wire w_dff_A_lSvp8Sbu1_0;
	wire w_dff_A_udFZ3Dq62_0;
	wire w_dff_A_BsUIBrL06_0;
	wire w_dff_A_XdoZMduP1_0;
	wire w_dff_A_x2zyQsxn2_0;
	wire w_dff_A_R88Dkp5e7_1;
	wire w_dff_A_PgfZ5iMz1_0;
	wire w_dff_A_5ar995Zr9_0;
	wire w_dff_A_bvX4qXK23_0;
	wire w_dff_A_ygLL3ad08_0;
	wire w_dff_A_jKnj2jlE8_0;
	wire w_dff_A_RtyD8z916_0;
	wire w_dff_A_fRKrrvAt0_0;
	wire w_dff_A_Z9UaPxn51_0;
	wire w_dff_A_nSMqXAOa3_0;
	wire w_dff_A_iYlIXvBp6_0;
	wire w_dff_A_OPtxso7F4_0;
	wire w_dff_A_donPucLe5_0;
	wire w_dff_A_S39SYTDx8_0;
	wire w_dff_A_KTChpuad1_0;
	wire w_dff_A_ElT9XbFR7_0;
	wire w_dff_A_5D3gpbdx6_0;
	wire w_dff_A_SUhHr1jl9_0;
	wire w_dff_A_rViJZvoT5_0;
	wire w_dff_A_cSgCoskL8_0;
	wire w_dff_A_V478lIvK7_0;
	wire w_dff_A_s8s7KUzL3_0;
	wire w_dff_A_imoyar1A6_0;
	wire w_dff_A_scCGR20z6_0;
	wire w_dff_A_VshQyyec1_0;
	wire w_dff_A_ZrAtgBOy7_0;
	wire w_dff_A_iwnZEO5h9_0;
	wire w_dff_A_VdZczkdE1_0;
	wire w_dff_A_eEEDelEM6_0;
	wire w_dff_A_5fdEYc6z9_2;
	wire w_dff_A_EORhwlQA5_0;
	wire w_dff_A_BCtXgJXy4_0;
	wire w_dff_A_HpSA6GNa2_0;
	wire w_dff_A_Z6W0c00I9_0;
	wire w_dff_A_iHS23Xyr0_0;
	wire w_dff_A_JTPkDerP5_0;
	wire w_dff_A_vVBTWctA0_0;
	wire w_dff_A_CIEdHvQv7_0;
	wire w_dff_A_7tpVCytZ9_0;
	wire w_dff_A_hO2CJKlI2_0;
	wire w_dff_A_3zfTOB0e0_2;
	wire w_dff_A_lSxQCspR5_0;
	wire w_dff_A_X4Ne4JLj5_0;
	wire w_dff_A_1OHz36ns6_0;
	wire w_dff_A_WYSgW46M0_0;
	wire w_dff_A_z71eXQPj8_0;
	wire w_dff_A_6RbivZWz4_0;
	wire w_dff_A_4LaOOQ7W1_0;
	wire w_dff_A_FovQvqSJ1_0;
	wire w_dff_A_fS9GxS7v6_0;
	wire w_dff_A_k5zg3SHu2_0;
	wire w_dff_A_fKN3Ov279_2;
	wire w_dff_A_kLygOFrb5_0;
	wire w_dff_A_A8k1YTxs7_0;
	wire w_dff_A_fWYw82rE4_0;
	wire w_dff_A_0iaYpmVK7_1;
	wire w_dff_A_nd7AJyg36_0;
	wire w_dff_A_f2JQRMEI9_0;
	wire w_dff_A_9moGAJdc7_0;
	wire w_dff_A_074rv2Fs0_0;
	wire w_dff_A_AfXj7ETA8_0;
	wire w_dff_A_YekKFm1z6_0;
	wire w_dff_A_kU9ikpeo2_0;
	wire w_dff_A_zLDth2L44_0;
	wire w_dff_A_CrMRH2oI7_0;
	wire w_dff_A_lE2sFZxr7_0;
	wire w_dff_A_4b11MPkO2_0;
	wire w_dff_A_AqDBN58x7_0;
	wire w_dff_A_055wRPif3_0;
	wire w_dff_A_RevDtGVB1_0;
	wire w_dff_A_4L3ylKuf4_0;
	wire w_dff_A_mQpxvKvk7_0;
	wire w_dff_A_Na6gBKa89_0;
	wire w_dff_A_xZ5XmhYy0_0;
	wire w_dff_A_N22YiHxz7_0;
	wire w_dff_A_8x1oYZfP3_0;
	wire w_dff_A_BYw8wZjg9_2;
	wire w_dff_A_V6aVPXsc1_0;
	wire w_dff_A_Bd28jUTQ4_0;
	wire w_dff_A_QMYkzvZA8_0;
	wire w_dff_A_VLQlYb5f8_0;
	wire w_dff_A_xPeoULhC5_0;
	wire w_dff_A_3tjmx9Te0_2;
	wire w_dff_A_EtOCEjPl6_0;
	wire w_dff_A_Bd5eKFnI8_0;
	wire w_dff_A_3N0DEjoK4_0;
	wire w_dff_A_hygaRTBY6_0;
	wire w_dff_A_gZ1v9epB1_2;
	wire w_dff_A_D7ucvZLP8_0;
	wire w_dff_A_5bO1MY4L3_0;
	wire w_dff_A_dvDrvt444_0;
	wire w_dff_A_2FUZ899C1_0;
	wire w_dff_A_XUGEsEnh5_0;
	wire w_dff_A_DNmFV2Mc1_0;
	wire w_dff_A_wP1tavFb2_0;
	wire w_dff_A_Tp7fuB0T8_0;
	wire w_dff_A_F2Gv4zZ05_2;
	wire w_dff_A_gy11JA5I7_0;
	wire w_dff_A_s76ba72r2_0;
	wire w_dff_A_ldh5CQJd0_0;
	wire w_dff_A_jwyxDsZy2_0;
	wire w_dff_A_7rEevuaQ2_0;
	wire w_dff_A_ffhrifTG8_0;
	wire w_dff_A_iu1Ysb078_0;
	wire w_dff_A_YhiS2eGY6_0;
	wire w_dff_A_7obnZiGZ1_2;
	wire w_dff_A_FE5QoXE37_0;
	wire w_dff_A_UdtblJ0F2_2;
	wire w_dff_A_6NY2N59Y3_0;
	wire w_dff_A_PsLnarY76_2;
	wire w_dff_A_xYPcZIYe7_0;
	wire w_dff_A_YlBNGGZi2_2;
	wire w_dff_A_8nPXRQOf6_0;
	wire w_dff_A_exSyuo865_0;
	wire w_dff_A_jtwMi6hO8_0;
	wire w_dff_A_QR7dOgq43_0;
	wire w_dff_A_Kk5KURfM1_0;
	wire w_dff_A_crNFTGrv7_0;
	wire w_dff_A_1BREmXEr6_0;
	wire w_dff_A_qJ50bqhN4_0;
	wire w_dff_A_BjosxPRc4_0;
	wire w_dff_A_4Ad49jj66_0;
	wire w_dff_A_8z8uGJbX4_0;
	wire w_dff_A_1Glriinb3_0;
	wire w_dff_A_LC1YCvD15_0;
	wire w_dff_A_gmEY2Ycu3_0;
	wire w_dff_A_wI6qLgtO3_0;
	wire w_dff_A_p0wxxp632_0;
	wire w_dff_A_9nSFi8Nl6_0;
	wire w_dff_A_CD2gKyok9_0;
	wire w_dff_A_mzpcjNh41_0;
	wire w_dff_A_MXOMLNmN4_0;
	wire w_dff_A_tXdazhKJ0_0;
	wire w_dff_A_gkBkkFd59_0;
	wire w_dff_A_wdOZv0zc9_0;
	wire w_dff_A_XcZolYWe6_0;
	wire w_dff_A_PSGSlOxf2_2;
	wire w_dff_A_yyOA2ltG6_0;
	wire w_dff_A_tgoJ9R3q8_0;
	wire w_dff_A_nRmN2kCU9_0;
	wire w_dff_A_kZHY9oCh1_0;
	wire w_dff_A_hZVgUNuc6_0;
	wire w_dff_A_FicGj5tX6_2;
	wire w_dff_A_VbWxeYIa1_0;
	wire w_dff_A_2btqfOnt3_0;
	wire w_dff_A_pY1t3G7j6_0;
	wire w_dff_A_4TrwIiOk1_0;
	wire w_dff_A_I9bGlMmw8_0;
	wire w_dff_A_IHdVYUXP2_2;
	wire w_dff_A_n66B77iq3_0;
	wire w_dff_A_h3tYHDBo0_0;
	wire w_dff_A_uCdvdXR31_0;
	wire w_dff_A_ThQPVUZP2_0;
	wire w_dff_A_LPZCpK0T7_0;
	wire w_dff_A_aKlzg0Oe8_2;
	wire w_dff_A_XKCHa7yq9_0;
	wire w_dff_A_9lGyOzaR7_0;
	wire w_dff_A_hbCd1HdE8_0;
	wire w_dff_A_yh5GrPfm0_0;
	wire w_dff_A_2uPZWpXo8_0;
	wire w_dff_A_LKzkoi9k2_0;
	wire w_dff_A_DgiL5ows8_0;
	wire w_dff_A_6BxXv4053_2;
	wire w_dff_A_T7FLFExf7_0;
	wire w_dff_A_gxXrxuWL9_0;
	wire w_dff_A_CUaJcXwy6_0;
	wire w_dff_A_rj3gX9H63_0;
	wire w_dff_A_LR5uCdEj9_0;
	wire w_dff_A_stHxCVM24_0;
	wire w_dff_A_KtULCR773_0;
	wire w_dff_A_4IIErU4q7_0;
	wire w_dff_A_h8jLWbDh0_0;
	wire w_dff_A_bFHILsoQ2_0;
	wire w_dff_A_uJlXdGCo4_0;
	wire w_dff_A_OA4O4XbX5_0;
	wire w_dff_A_mV9ksafz0_0;
	wire w_dff_A_EPDQAWEU0_0;
	wire w_dff_A_LQYxvjbz1_0;
	wire w_dff_A_O7a0owzQ8_0;
	wire w_dff_A_zp7is1dU1_0;
	wire w_dff_A_evLEjbNM1_0;
	wire w_dff_A_V10yD3eU5_0;
	wire w_dff_A_3gY2Zx692_2;
	wire w_dff_A_YEfry8FO8_0;
	wire w_dff_A_aRxRy8Qx1_2;
	wire w_dff_A_M26jmssu0_0;
	wire w_dff_A_pGz0TzDp7_2;
	wire w_dff_A_1Ze2UWsQ7_0;
	wire w_dff_A_tRBRv4QH4_0;
	wire w_dff_A_ArwEOjAo5_0;
	wire w_dff_A_K1LKraZY5_0;
	wire w_dff_A_FnHRRYsr4_0;
	wire w_dff_A_mGv8qgAs6_0;
	wire w_dff_A_1iNBjEtb2_0;
	wire w_dff_A_TZUlzPwn3_0;
	wire w_dff_A_0bS4kFjy0_0;
	wire w_dff_A_n88kCQf22_0;
	wire w_dff_A_rvnlIuCq0_0;
	wire w_dff_A_cbZfSeR66_0;
	wire w_dff_A_4RSug8h85_0;
	wire w_dff_A_Cuc6i5YH6_0;
	wire w_dff_A_bC7cKcKa8_0;
	wire w_dff_A_jXnLANAr8_0;
	wire w_dff_A_f6XPnz5h0_0;
	wire w_dff_A_39LSarcR8_2;
	wire w_dff_A_Or38g4ww3_0;
	wire w_dff_A_frBTXjWn8_0;
	wire w_dff_A_wCld7PdR6_0;
	wire w_dff_A_Dk1DG5NK1_0;
	wire w_dff_A_NDIquvQZ6_0;
	wire w_dff_A_lpfcRF452_0;
	wire w_dff_A_hTgLSKpD6_0;
	wire w_dff_A_eshq81ff7_0;
	wire w_dff_A_oeDvoZ4n8_0;
	wire w_dff_A_KXMEQTyr6_0;
	wire w_dff_A_XPTkbgQm6_0;
	wire w_dff_A_IJAOBrqm7_0;
	wire w_dff_A_E1DccclB9_0;
	wire w_dff_A_R2ygSeKK7_0;
	wire w_dff_A_aQ9HZ5sN7_0;
	wire w_dff_A_uzccgCpY4_0;
	wire w_dff_A_WEZgCqLO8_0;
	wire w_dff_A_Ok6uAbWN4_2;
	wire w_dff_A_0ayCAdl21_0;
	wire w_dff_A_Hai4Bxo74_0;
	wire w_dff_A_fUvfw16W8_0;
	wire w_dff_A_cWyOtGep6_0;
	wire w_dff_A_IHHwLxq40_0;
	wire w_dff_A_hrMgtwa86_0;
	wire w_dff_A_F4nXchMr5_0;
	wire w_dff_A_kZcCp9ng2_0;
	wire w_dff_A_l4l0kOFP9_0;
	wire w_dff_A_9vqlPN4g2_0;
	wire w_dff_A_GLPquVQM1_0;
	wire w_dff_A_e8yGQNQJ4_0;
	wire w_dff_A_RqlPRQDE2_0;
	wire w_dff_A_VBz0642q7_0;
	wire w_dff_A_1tUKpQca0_0;
	wire w_dff_A_QUQ54itN9_0;
	wire w_dff_A_Bmbl6rZ65_0;
	wire w_dff_A_N1mAsmmi2_2;
	wire w_dff_A_e86IiVHH3_0;
	wire w_dff_A_M36832ah7_0;
	wire w_dff_A_e0Orb4lA6_0;
	wire w_dff_A_5eBgw1Tk2_0;
	wire w_dff_A_JcuY7N3g4_0;
	wire w_dff_A_zPNojqUB6_0;
	wire w_dff_A_BrEpKekj3_0;
	wire w_dff_A_encOh2s40_0;
	wire w_dff_A_9cJOMgqh0_0;
	wire w_dff_A_fRd1r4RP4_0;
	wire w_dff_A_CZbadehM3_0;
	wire w_dff_A_lswNp0EP2_0;
	wire w_dff_A_qlGniEvj2_0;
	wire w_dff_A_N007mEEt9_0;
	wire w_dff_A_DS3zjS1V5_0;
	wire w_dff_A_b5ZoaKfv0_0;
	wire w_dff_A_Z8oRwTuK9_0;
	wire w_dff_A_HerJdIIO9_2;
	wire w_dff_A_Zw4k2O9c9_0;
	wire w_dff_A_ORQZ0sdf8_0;
	wire w_dff_A_T46XX8Qa8_0;
	wire w_dff_A_erjosBMk0_0;
	wire w_dff_A_fuPWfSGP0_0;
	wire w_dff_A_YvaQSWAJ8_0;
	wire w_dff_A_7bjsJIrq2_0;
	wire w_dff_A_D9Te1xWZ6_0;
	wire w_dff_A_PhUca8Jx0_0;
	wire w_dff_A_aWMShC4i6_0;
	wire w_dff_A_WbEsNmol1_0;
	wire w_dff_A_szg5BwvA8_0;
	wire w_dff_A_cmrFAdAy7_2;
	wire w_dff_A_JJeTwaYA8_0;
	wire w_dff_A_dii8jI0N8_0;
	wire w_dff_A_ubCvPUdn0_0;
	wire w_dff_A_3LMAsPgj4_0;
	wire w_dff_A_6j41Zqs12_0;
	wire w_dff_A_73sxFhUA2_0;
	wire w_dff_A_9b2rEQ9O6_0;
	wire w_dff_A_opntaJuZ7_0;
	wire w_dff_A_ftHqaEUe4_0;
	wire w_dff_A_JTd57Y9V7_0;
	wire w_dff_A_fZnjr7TN2_0;
	wire w_dff_A_8MpDjeCt8_0;
	wire w_dff_A_7kOYqbgg5_0;
	wire w_dff_A_zYA4qFmc0_2;
	wire w_dff_A_xCaeHS7k4_0;
	wire w_dff_A_91RMdsVf8_0;
	wire w_dff_A_buf0kbXX3_0;
	wire w_dff_A_kfjrNXJh5_0;
	wire w_dff_A_BLuQR1Qx7_0;
	wire w_dff_A_HYhVbmDM8_0;
	wire w_dff_A_FkCRMnaE6_0;
	wire w_dff_A_uRo3uB4I6_0;
	wire w_dff_A_rdB7BPKt8_0;
	wire w_dff_A_UbmbXZi94_0;
	wire w_dff_A_3Wdne82Z6_0;
	wire w_dff_A_4roMcrxw9_0;
	wire w_dff_A_8fCtJaLk4_0;
	wire w_dff_A_KNA2aBHr1_0;
	wire w_dff_A_FNRnCz2S2_0;
	wire w_dff_A_IpwnXTLg0_2;
	wire w_dff_A_1KQy76900_0;
	wire w_dff_A_NNJdX76P6_0;
	wire w_dff_A_LtTshqNf1_0;
	wire w_dff_A_2YNl0r4s9_0;
	wire w_dff_A_HDpytnws8_0;
	wire w_dff_A_LEfRcKZu6_0;
	wire w_dff_A_kQQnB38u1_0;
	wire w_dff_A_EfBYDn0W6_0;
	wire w_dff_A_5rgiUtMz3_0;
	wire w_dff_A_bDmVCKah5_0;
	wire w_dff_A_4UV6Aa7P7_0;
	wire w_dff_A_Kh6KxNtQ8_0;
	wire w_dff_A_HhDMNim98_0;
	wire w_dff_A_UZQTJyrc7_0;
	wire w_dff_A_KGm3qQhT2_0;
	wire w_dff_A_CJf3sWow9_0;
	wire w_dff_A_wIhJ1ELX0_0;
	wire w_dff_A_DxbKqrBV1_2;
	wire w_dff_A_BsORI0N07_0;
	wire w_dff_A_RdRs7Zcf0_0;
	wire w_dff_A_74jZjFLF0_0;
	wire w_dff_A_ZVxD6Kul4_0;
	wire w_dff_A_ihJQiTas3_0;
	wire w_dff_A_SofaJqix2_2;
	wire w_dff_A_jT5X6nYq2_2;
	wire w_dff_A_T7aJU2ej9_0;
	wire w_dff_A_TfS78Cxh5_0;
	wire w_dff_A_52IkDmef8_0;
	wire w_dff_A_AHIN5y2A5_0;
	wire w_dff_A_87HskYOj1_0;
	wire w_dff_A_koxF0wgk2_0;
	wire w_dff_A_JuP36eVp6_0;
	wire w_dff_A_pe6aqDYz1_0;
	wire w_dff_A_dQ9g9yfS3_0;
	wire w_dff_A_1jKm0Lkr1_0;
	wire w_dff_A_l9tCs6TB9_0;
	wire w_dff_A_q059EdLg0_0;
	wire w_dff_A_3lC6Xhkx8_0;
	wire w_dff_A_d6aRNQxc8_0;
	wire w_dff_A_xxupOa4X3_0;
	wire w_dff_A_U4owkrqr3_0;
	wire w_dff_A_3UnuSp1X4_2;
	wire w_dff_A_K8LeKm9Q2_0;
	wire w_dff_A_GC3ghFZB9_0;
	wire w_dff_A_ESuSZBGM1_0;
	wire w_dff_A_uTtzCnn51_0;
	wire w_dff_A_yEjBOBBS7_0;
	wire w_dff_A_nbJmh1Ss8_0;
	wire w_dff_A_ynywxUvS5_0;
	wire w_dff_A_NKEk5aAE6_0;
	wire w_dff_A_TNlNeo4I2_0;
	wire w_dff_A_cZ4FOvJs2_0;
	wire w_dff_A_IiVWy0E29_0;
	wire w_dff_A_3m5eUpMJ9_0;
	wire w_dff_A_8HyNi9Vr8_0;
	wire w_dff_A_QzauXjnj9_0;
	wire w_dff_A_QHuSf2Ia6_0;
	wire w_dff_A_zS6HEnMW4_0;
	wire w_dff_A_wyp349xj3_0;
	wire w_dff_A_OSd91su29_0;
	wire w_dff_A_yCUoTRVp8_0;
	wire w_dff_A_iKhB3adl6_0;
	jnot g0000(.din(w_G15_0[2]),.dout(w_dff_A_TSybH3fu9_1),.clk(gclk));
	jor g0001(.dina(G57),.dinb(w_G5_1[1]),.dout(w_dff_A_ytKocOgQ9_2),.clk(gclk));
	jnot g0002(.din(G184),.dout(n317),.clk(gclk));
	jnot g0003(.din(G228),.dout(n318),.clk(gclk));
	jor g0004(.dina(n318),.dinb(n317),.dout(n319),.clk(gclk));
	jnot g0005(.din(G150),.dout(n320),.clk(gclk));
	jnot g0006(.din(G240),.dout(n321),.clk(gclk));
	jor g0007(.dina(n321),.dinb(n320),.dout(n322),.clk(gclk));
	jor g0008(.dina(n322),.dinb(n319),.dout(G404_fa_),.clk(gclk));
	jnot g0009(.din(G210),.dout(n324),.clk(gclk));
	jnot g0010(.din(G218),.dout(n325),.clk(gclk));
	jor g0011(.dina(n325),.dinb(n324),.dout(n326),.clk(gclk));
	jnot g0012(.din(G152),.dout(n327),.clk(gclk));
	jnot g0013(.din(G230),.dout(n328),.clk(gclk));
	jor g0014(.dina(n328),.dinb(n327),.dout(n329),.clk(gclk));
	jor g0015(.dina(n329),.dinb(n326),.dout(G406_fa_),.clk(gclk));
	jnot g0016(.din(G183),.dout(n331),.clk(gclk));
	jnot g0017(.din(G185),.dout(n332),.clk(gclk));
	jor g0018(.dina(n332),.dinb(n331),.dout(n333),.clk(gclk));
	jnot g0019(.din(G182),.dout(n334),.clk(gclk));
	jnot g0020(.din(G186),.dout(n335),.clk(gclk));
	jor g0021(.dina(n335),.dinb(n334),.dout(n336),.clk(gclk));
	jor g0022(.dina(n336),.dinb(n333),.dout(G408_fa_),.clk(gclk));
	jnot g0023(.din(G172),.dout(n338),.clk(gclk));
	jnot g0024(.din(G188),.dout(n339),.clk(gclk));
	jor g0025(.dina(n339),.dinb(n338),.dout(n340),.clk(gclk));
	jnot g0026(.din(G162),.dout(n341),.clk(gclk));
	jnot g0027(.din(G199),.dout(n342),.clk(gclk));
	jor g0028(.dina(n342),.dinb(n341),.dout(n343),.clk(gclk));
	jor g0029(.dina(n343),.dinb(n340),.dout(G410_fa_),.clk(gclk));
	jnot g0030(.din(G1197),.dout(n345),.clk(gclk));
	jor g0031(.dina(w_n345_0[1]),.dinb(w_G5_1[0]),.dout(w_dff_A_wmykSRR86_2),.clk(gclk));
	jnot g0032(.din(G134),.dout(n347),.clk(gclk));
	jnot g0033(.din(G133),.dout(n348),.clk(gclk));
	jor g0034(.dina(n348),.dinb(w_G5_0[2]),.dout(n349),.clk(gclk));
	jor g0035(.dina(w_n349_0[1]),.dinb(w_n347_0[1]),.dout(w_dff_A_D8xH8Oi22_2),.clk(gclk));
	jand g0036(.dina(G163),.dinb(w_G1_1[2]),.dout(w_dff_A_yJxiPeRD1_2),.clk(gclk));
	jnot g0037(.din(w_G41_0[1]),.dout(n352),.clk(gclk));
	jor g0038(.dina(n352),.dinb(w_G18_49[2]),.dout(n353),.clk(gclk));
	jor g0039(.dina(w_n353_0[1]),.dinb(w_G3701_1[1]),.dout(n354),.clk(gclk));
	jnot g0040(.din(w_G18_49[1]),.dout(n355),.clk(gclk));
	jand g0041(.dina(w_G3701_1[0]),.dinb(w_n355_35[2]),.dout(n356),.clk(gclk));
	jand g0042(.dina(n356),.dinb(w_n353_0[0]),.dout(n357),.clk(gclk));
	jnot g0043(.din(w_n357_0[1]),.dout(n358),.clk(gclk));
	jand g0044(.dina(w_n358_0[1]),.dinb(w_n354_0[2]),.dout(n359),.clk(gclk));
	jxor g0045(.dina(w_n359_1[1]),.dinb(w_G4526_2[2]),.dout(w_dff_A_62FaZpmK6_2),.clk(gclk));
	jnot g0046(.din(w_G38_2[2]),.dout(n361),.clk(gclk));
	jand g0047(.dina(w_G4528_0[2]),.dinb(w_G1492_1[1]),.dout(n362),.clk(gclk));
	jxor g0048(.dina(w_n362_0[2]),.dinb(w_n361_0[2]),.dout(n363),.clk(gclk));
	jand g0049(.dina(w_G4528_0[1]),.dinb(w_G1496_1[1]),.dout(n364),.clk(gclk));
	jor g0050(.dina(w_n364_0[2]),.dinb(w_n361_0[1]),.dout(n365),.clk(gclk));
	jnot g0051(.din(w_G1496_1[0]),.dout(n366),.clk(gclk));
	jnot g0052(.din(w_G4528_0[0]),.dout(n367),.clk(gclk));
	jor g0053(.dina(w_n367_0[1]),.dinb(w_G38_2[1]),.dout(n368),.clk(gclk));
	jor g0054(.dina(w_n368_0[1]),.dinb(w_n366_0[2]),.dout(n369),.clk(gclk));
	jand g0055(.dina(w_n369_0[1]),.dinb(w_dff_B_XV3MfLLv5_1),.dout(n370),.clk(gclk));
	jnot g0056(.din(w_G1486_0[1]),.dout(n371),.clk(gclk));
	jand g0057(.dina(G12),.dinb(G9),.dout(n372),.clk(gclk));
	jnot g0058(.din(w_n372_0[1]),.dout(n373),.clk(gclk));
	jor g0059(.dina(w_dff_B_xc9uFfJ31_0),.dinb(w_n355_35[1]),.dout(n374),.clk(gclk));
	jand g0060(.dina(w_n374_0[1]),.dinb(w_n373_9[2]),.dout(n375),.clk(gclk));
	jand g0061(.dina(w_n375_0[2]),.dinb(w_n371_0[2]),.dout(n376),.clk(gclk));
	jxor g0062(.dina(w_n375_0[1]),.dinb(w_n371_0[1]),.dout(n377),.clk(gclk));
	jor g0063(.dina(w_dff_B_l5zNm9Gi9_0),.dinb(w_n355_35[0]),.dout(n378),.clk(gclk));
	jand g0064(.dina(w_n378_0[1]),.dinb(w_n373_9[1]),.dout(n379),.clk(gclk));
	jnot g0065(.din(w_n379_0[2]),.dout(n380),.clk(gclk));
	jand g0066(.dina(w_n380_0[1]),.dinb(w_G1480_0[2]),.dout(n381),.clk(gclk));
	jnot g0067(.din(n381),.dout(n382),.clk(gclk));
	jnot g0068(.din(w_G1480_0[1]),.dout(n383),.clk(gclk));
	jand g0069(.dina(w_n379_0[1]),.dinb(w_n383_0[2]),.dout(n384),.clk(gclk));
	jnot g0070(.din(w_G106_1[1]),.dout(n385),.clk(gclk));
	jor g0071(.dina(w_dff_B_A4tUEeHk1_0),.dinb(w_n355_34[2]),.dout(n386),.clk(gclk));
	jand g0072(.dina(w_n386_0[1]),.dinb(w_n373_9[0]),.dout(n387),.clk(gclk));
	jxor g0073(.dina(w_n387_1[1]),.dinb(w_n385_0[1]),.dout(n388),.clk(gclk));
	jnot g0074(.din(w_G1462_0[1]),.dout(n389),.clk(gclk));
	jor g0075(.dina(w_G209_0[1]),.dinb(w_n355_34[1]),.dout(n390),.clk(gclk));
	jand g0076(.dina(n390),.dinb(w_n373_8[2]),.dout(n391),.clk(gclk));
	jand g0077(.dina(w_n391_0[2]),.dinb(w_n389_1[1]),.dout(n392),.clk(gclk));
	jnot g0078(.din(w_G1469_0[1]),.dout(n393),.clk(gclk));
	jor g0079(.dina(w_dff_B_6lWvEOl36_0),.dinb(w_n355_34[0]),.dout(n394),.clk(gclk));
	jand g0080(.dina(w_n394_0[1]),.dinb(w_n373_8[1]),.dout(n395),.clk(gclk));
	jxor g0081(.dina(w_n395_1[1]),.dinb(w_n393_1[1]),.dout(n396),.clk(gclk));
	jand g0082(.dina(w_n396_1[2]),.dinb(w_n392_0[2]),.dout(n397),.clk(gclk));
	jand g0083(.dina(w_n397_0[1]),.dinb(w_n388_1[2]),.dout(n398),.clk(gclk));
	jnot g0084(.din(n398),.dout(n399),.clk(gclk));
	jand g0085(.dina(w_n387_1[0]),.dinb(w_n385_0[0]),.dout(n400),.clk(gclk));
	jnot g0086(.din(n400),.dout(n401),.clk(gclk));
	jnot g0087(.din(w_n387_0[2]),.dout(n402),.clk(gclk));
	jand g0088(.dina(n402),.dinb(w_G106_1[0]),.dout(n403),.clk(gclk));
	jand g0089(.dina(w_n395_1[0]),.dinb(w_n393_1[0]),.dout(n404),.clk(gclk));
	jnot g0090(.din(n404),.dout(n405),.clk(gclk));
	jor g0091(.dina(w_n405_0[2]),.dinb(n403),.dout(n406),.clk(gclk));
	jand g0092(.dina(n406),.dinb(w_dff_B_2gdIxIEi6_1),.dout(n407),.clk(gclk));
	jand g0093(.dina(w_n407_0[1]),.dinb(n399),.dout(n408),.clk(gclk));
	jnot g0094(.din(n408),.dout(n409),.clk(gclk));
	jor g0095(.dina(w_n409_1[1]),.dinb(w_dff_B_K0MX5dgt9_1),.dout(n410),.clk(gclk));
	jand g0096(.dina(n410),.dinb(w_dff_B_V0Nq0Ly36_1),.dout(n411),.clk(gclk));
	jand g0097(.dina(w_n411_1[1]),.dinb(w_n377_1[2]),.dout(n412),.clk(gclk));
	jor g0098(.dina(n412),.dinb(w_dff_B_JlSU60wd0_1),.dout(n413),.clk(gclk));
	jxor g0099(.dina(w_n391_0[1]),.dinb(w_n389_1[0]),.dout(n414),.clk(gclk));
	jand g0100(.dina(w_n414_1[1]),.dinb(w_n396_1[1]),.dout(n415),.clk(gclk));
	jxor g0101(.dina(w_n379_0[0]),.dinb(w_n383_0[1]),.dout(n416),.clk(gclk));
	jand g0102(.dina(w_n416_0[2]),.dinb(w_n388_1[1]),.dout(n417),.clk(gclk));
	jand g0103(.dina(n417),.dinb(w_n415_0[1]),.dout(n418),.clk(gclk));
	jand g0104(.dina(w_n418_0[1]),.dinb(w_n377_1[1]),.dout(n419),.clk(gclk));
	jor g0105(.dina(w_n419_0[1]),.dinb(w_n413_1[1]),.dout(n420),.clk(gclk));
	jnot g0106(.din(w_G2256_0[1]),.dout(n421),.clk(gclk));
	jor g0107(.dina(w_dff_B_zfCEdJOT5_0),.dinb(w_n355_33[2]),.dout(n422),.clk(gclk));
	jand g0108(.dina(w_n422_0[1]),.dinb(w_n373_8[0]),.dout(n423),.clk(gclk));
	jand g0109(.dina(w_n423_0[2]),.dinb(w_n421_0[2]),.dout(n424),.clk(gclk));
	jxor g0110(.dina(w_n423_0[1]),.dinb(w_n421_0[1]),.dout(n425),.clk(gclk));
	jnot g0111(.din(w_G2253_0[2]),.dout(n426),.clk(gclk));
	jor g0112(.dina(w_dff_B_pvlpNQrM0_0),.dinb(w_n355_33[1]),.dout(n427),.clk(gclk));
	jand g0113(.dina(w_n427_0[1]),.dinb(w_n373_7[2]),.dout(n428),.clk(gclk));
	jxor g0114(.dina(w_n428_0[2]),.dinb(w_n426_0[2]),.dout(n429),.clk(gclk));
	jnot g0115(.din(w_G2247_0[2]),.dout(n430),.clk(gclk));
	jor g0116(.dina(w_dff_B_pPgfFLMk6_0),.dinb(w_n355_33[0]),.dout(n431),.clk(gclk));
	jand g0117(.dina(w_n431_0[1]),.dinb(w_n373_7[1]),.dout(n432),.clk(gclk));
	jxor g0118(.dina(w_n432_0[2]),.dinb(w_n430_0[1]),.dout(n433),.clk(gclk));
	jnot g0119(.din(w_G2239_1[1]),.dout(n434),.clk(gclk));
	jor g0120(.dina(w_dff_B_izHlvbbm7_0),.dinb(w_n355_32[2]),.dout(n435),.clk(gclk));
	jand g0121(.dina(w_n435_0[1]),.dinb(w_n373_7[0]),.dout(n436),.clk(gclk));
	jxor g0122(.dina(w_n436_0[2]),.dinb(w_n434_0[1]),.dout(n437),.clk(gclk));
	jand g0123(.dina(w_n437_0[2]),.dinb(w_n433_1[2]),.dout(n438),.clk(gclk));
	jand g0124(.dina(w_n438_0[1]),.dinb(w_n429_0[2]),.dout(n439),.clk(gclk));
	jnot g0125(.din(w_n428_0[1]),.dout(n440),.clk(gclk));
	jand g0126(.dina(w_n440_0[1]),.dinb(w_G2253_0[1]),.dout(n441),.clk(gclk));
	jnot g0127(.din(n441),.dout(n442),.clk(gclk));
	jand g0128(.dina(w_n428_0[0]),.dinb(w_n426_0[1]),.dout(n443),.clk(gclk));
	jand g0129(.dina(w_n432_0[1]),.dinb(w_n430_0[0]),.dout(n444),.clk(gclk));
	jand g0130(.dina(w_n436_0[1]),.dinb(w_n434_0[0]),.dout(n445),.clk(gclk));
	jand g0131(.dina(w_n445_0[2]),.dinb(w_n433_1[1]),.dout(n446),.clk(gclk));
	jor g0132(.dina(n446),.dinb(w_n444_0[2]),.dout(n447),.clk(gclk));
	jor g0133(.dina(w_n447_0[2]),.dinb(w_dff_B_Ou96JSKD7_1),.dout(n448),.clk(gclk));
	jand g0134(.dina(n448),.dinb(w_dff_B_92yrD0BR6_1),.dout(n449),.clk(gclk));
	jor g0135(.dina(w_n449_1[1]),.dinb(w_dff_B_jcpkSiok6_1),.dout(n450),.clk(gclk));
	jnot g0136(.din(w_G2236_0[2]),.dout(n451),.clk(gclk));
	jor g0137(.dina(w_dff_B_EvTmIQ8u7_0),.dinb(w_n355_32[1]),.dout(n452),.clk(gclk));
	jand g0138(.dina(n452),.dinb(w_n373_6[2]),.dout(n453),.clk(gclk));
	jand g0139(.dina(w_n453_1[1]),.dinb(w_n451_0[2]),.dout(n454),.clk(gclk));
	jor g0140(.dina(w_n453_1[0]),.dinb(w_n451_0[1]),.dout(n455),.clk(gclk));
	jnot g0141(.din(w_G2230_0[2]),.dout(n456),.clk(gclk));
	jand g0142(.dina(w_dff_B_ysREwqJz0_0),.dinb(w_n355_32[0]),.dout(n457),.clk(gclk));
	jand g0143(.dina(G158),.dinb(w_G18_49[0]),.dout(n458),.clk(gclk));
	jor g0144(.dina(w_dff_B_OMw2dKd80_0),.dinb(w_n457_0[1]),.dout(n459),.clk(gclk));
	jand g0145(.dina(w_n459_0[2]),.dinb(w_n456_0[2]),.dout(n460),.clk(gclk));
	jand g0146(.dina(w_n460_1[2]),.dinb(n455),.dout(n461),.clk(gclk));
	jor g0147(.dina(n461),.dinb(w_dff_B_awopLnNH5_1),.dout(n462),.clk(gclk));
	jxor g0148(.dina(w_n453_0[2]),.dinb(w_n451_0[0]),.dout(n463),.clk(gclk));
	jxor g0149(.dina(w_n459_0[1]),.dinb(w_n456_0[1]),.dout(n464),.clk(gclk));
	jand g0150(.dina(w_n464_0[2]),.dinb(w_n463_1[1]),.dout(n465),.clk(gclk));
	jnot g0151(.din(w_G2224_1[1]),.dout(n466),.clk(gclk));
	jand g0152(.dina(w_dff_B_L0FO5yLy8_0),.dinb(w_n355_31[2]),.dout(n467),.clk(gclk));
	jand g0153(.dina(G159),.dinb(w_G18_48[2]),.dout(n468),.clk(gclk));
	jor g0154(.dina(w_dff_B_KFM86BYY5_0),.dinb(w_n467_0[1]),.dout(n469),.clk(gclk));
	jxor g0155(.dina(w_n469_1[1]),.dinb(w_n466_0[1]),.dout(n470),.clk(gclk));
	jnot g0156(.din(w_G2218_0[2]),.dout(n471),.clk(gclk));
	jand g0157(.dina(w_dff_B_F3PASO123_0),.dinb(w_n355_31[1]),.dout(n472),.clk(gclk));
	jand g0158(.dina(G160),.dinb(w_G18_48[1]),.dout(n473),.clk(gclk));
	jor g0159(.dina(w_dff_B_ahLzISW37_0),.dinb(w_n472_0[1]),.dout(n474),.clk(gclk));
	jxor g0160(.dina(w_n474_0[2]),.dinb(w_n471_0[2]),.dout(n475),.clk(gclk));
	jnot g0161(.din(w_G2211_0[2]),.dout(n476),.clk(gclk));
	jand g0162(.dina(w_dff_B_sPQTSDO91_0),.dinb(w_n355_31[0]),.dout(n477),.clk(gclk));
	jand g0163(.dina(G151),.dinb(w_G18_48[0]),.dout(n478),.clk(gclk));
	jor g0164(.dina(w_dff_B_YBVMhFrw4_0),.dinb(w_n477_0[1]),.dout(n479),.clk(gclk));
	jxor g0165(.dina(w_n479_1[1]),.dinb(w_n476_0[2]),.dout(n480),.clk(gclk));
	jand g0166(.dina(w_n480_1[1]),.dinb(w_n475_0[2]),.dout(n481),.clk(gclk));
	jand g0167(.dina(w_n481_0[1]),.dinb(w_n470_0[2]),.dout(n482),.clk(gclk));
	jnot g0168(.din(w_n469_1[0]),.dout(n483),.clk(gclk));
	jand g0169(.dina(n483),.dinb(w_G2224_1[0]),.dout(n484),.clk(gclk));
	jnot g0170(.din(w_n474_0[1]),.dout(n485),.clk(gclk));
	jand g0171(.dina(w_n485_0[1]),.dinb(w_G2218_0[1]),.dout(n486),.clk(gclk));
	jand g0172(.dina(w_n479_1[0]),.dinb(w_n476_0[1]),.dout(n487),.clk(gclk));
	jnot g0173(.din(w_n487_0[2]),.dout(n488),.clk(gclk));
	jor g0174(.dina(n488),.dinb(w_n486_0[1]),.dout(n489),.clk(gclk));
	jand g0175(.dina(w_n469_0[2]),.dinb(w_n466_0[0]),.dout(n490),.clk(gclk));
	jand g0176(.dina(w_n474_0[0]),.dinb(w_n471_0[1]),.dout(n491),.clk(gclk));
	jor g0177(.dina(w_n491_1[1]),.dinb(n490),.dout(n492),.clk(gclk));
	jnot g0178(.din(n492),.dout(n493),.clk(gclk));
	jand g0179(.dina(n493),.dinb(w_n489_0[2]),.dout(n494),.clk(gclk));
	jor g0180(.dina(n494),.dinb(w_dff_B_2dzCEDNR0_1),.dout(n495),.clk(gclk));
	jnot g0181(.din(w_n495_1[1]),.dout(n496),.clk(gclk));
	jor g0182(.dina(w_n496_0[2]),.dinb(w_dff_B_g08RlGq63_1),.dout(n497),.clk(gclk));
	jand g0183(.dina(w_n497_1[1]),.dinb(w_n465_0[1]),.dout(n498),.clk(gclk));
	jor g0184(.dina(n498),.dinb(w_n462_0[2]),.dout(n499),.clk(gclk));
	jand g0185(.dina(w_n496_0[1]),.dinb(w_n465_0[0]),.dout(n500),.clk(gclk));
	jnot g0186(.din(w_G4437_0[2]),.dout(n501),.clk(gclk));
	jand g0187(.dina(G219),.dinb(w_G18_47[2]),.dout(n502),.clk(gclk));
	jand g0188(.dina(w_dff_B_hevlZQKt0_0),.dinb(w_n355_30[2]),.dout(n503),.clk(gclk));
	jor g0189(.dina(w_n503_0[1]),.dinb(w_dff_B_OjPSi83b8_1),.dout(n504),.clk(gclk));
	jand g0190(.dina(w_n504_1[1]),.dinb(w_n501_0[2]),.dout(n505),.clk(gclk));
	jnot g0191(.din(w_n504_1[0]),.dout(n506),.clk(gclk));
	jand g0192(.dina(n506),.dinb(w_G4437_0[1]),.dout(n507),.clk(gclk));
	jnot g0193(.din(w_n507_0[1]),.dout(n508),.clk(gclk));
	jnot g0194(.din(w_G4432_0[2]),.dout(n509),.clk(gclk));
	jand g0195(.dina(G220),.dinb(w_G18_47[1]),.dout(n510),.clk(gclk));
	jand g0196(.dina(w_dff_B_kh9eKsd88_0),.dinb(w_n355_30[1]),.dout(n511),.clk(gclk));
	jor g0197(.dina(w_n511_0[1]),.dinb(w_dff_B_eprve7413_1),.dout(n512),.clk(gclk));
	jxor g0198(.dina(w_n512_0[2]),.dinb(w_n509_0[2]),.dout(n513),.clk(gclk));
	jnot g0199(.din(w_G4420_1[1]),.dout(n514),.clk(gclk));
	jand g0200(.dina(G222),.dinb(w_G18_47[0]),.dout(n515),.clk(gclk));
	jand g0201(.dina(w_dff_B_6Hnef3P70_0),.dinb(w_n355_30[0]),.dout(n516),.clk(gclk));
	jor g0202(.dina(w_n516_0[1]),.dinb(w_dff_B_kgtB5zK48_1),.dout(n517),.clk(gclk));
	jand g0203(.dina(w_n517_1[1]),.dinb(w_n514_0[1]),.dout(n518),.clk(gclk));
	jnot g0204(.din(w_n518_1[2]),.dout(n519),.clk(gclk));
	jnot g0205(.din(w_G4427_0[2]),.dout(n520),.clk(gclk));
	jand g0206(.dina(G221),.dinb(w_G18_46[2]),.dout(n521),.clk(gclk));
	jand g0207(.dina(w_dff_B_FI8IhTCi2_0),.dinb(w_n355_29[2]),.dout(n522),.clk(gclk));
	jor g0208(.dina(w_n522_0[1]),.dinb(w_dff_B_1uxc9meZ2_1),.dout(n523),.clk(gclk));
	jxor g0209(.dina(w_n523_0[2]),.dinb(w_n520_0[1]),.dout(n524),.clk(gclk));
	jnot g0210(.din(w_n517_1[0]),.dout(n525),.clk(gclk));
	jand g0211(.dina(n525),.dinb(w_G4420_1[0]),.dout(n526),.clk(gclk));
	jnot g0212(.din(w_n526_0[2]),.dout(n527),.clk(gclk));
	jnot g0213(.din(w_G4415_1[1]),.dout(n528),.clk(gclk));
	jand g0214(.dina(G223),.dinb(w_G18_46[1]),.dout(n529),.clk(gclk));
	jand g0215(.dina(w_dff_B_kRuWr5Ze3_0),.dinb(w_n355_29[1]),.dout(n530),.clk(gclk));
	jor g0216(.dina(w_n530_0[1]),.dinb(w_dff_B_t9qFBe8s0_1),.dout(n531),.clk(gclk));
	jand g0217(.dina(w_n531_1[1]),.dinb(w_n528_0[1]),.dout(n532),.clk(gclk));
	jnot g0218(.din(w_n531_1[0]),.dout(n533),.clk(gclk));
	jand g0219(.dina(n533),.dinb(w_G4415_1[0]),.dout(n534),.clk(gclk));
	jnot g0220(.din(n534),.dout(n535),.clk(gclk));
	jnot g0221(.din(w_G4410_0[2]),.dout(n536),.clk(gclk));
	jand g0222(.dina(G224),.dinb(w_G18_46[0]),.dout(n537),.clk(gclk));
	jand g0223(.dina(w_dff_B_p60qXJgH6_0),.dinb(w_n355_29[0]),.dout(n538),.clk(gclk));
	jor g0224(.dina(w_n538_0[1]),.dinb(w_dff_B_dQ2S0xJ08_1),.dout(n539),.clk(gclk));
	jand g0225(.dina(w_n539_1[1]),.dinb(w_n536_0[2]),.dout(n540),.clk(gclk));
	jnot g0226(.din(w_n539_1[0]),.dout(n541),.clk(gclk));
	jand g0227(.dina(n541),.dinb(w_G4410_0[1]),.dout(n542),.clk(gclk));
	jnot g0228(.din(n542),.dout(n543),.clk(gclk));
	jnot g0229(.din(w_G4405_1[1]),.dout(n544),.clk(gclk));
	jand g0230(.dina(G225),.dinb(w_G18_45[2]),.dout(n545),.clk(gclk));
	jand g0231(.dina(w_dff_B_Riboc5A53_0),.dinb(w_n355_28[2]),.dout(n546),.clk(gclk));
	jor g0232(.dina(w_n546_0[1]),.dinb(w_dff_B_qIPZoZRM4_1),.dout(n547),.clk(gclk));
	jand g0233(.dina(w_n547_1[1]),.dinb(w_n544_0[1]),.dout(n548),.clk(gclk));
	jnot g0234(.din(w_n547_1[0]),.dout(n549),.clk(gclk));
	jand g0235(.dina(n549),.dinb(w_G4405_1[0]),.dout(n550),.clk(gclk));
	jnot g0236(.din(w_n550_0[1]),.dout(n551),.clk(gclk));
	jnot g0237(.din(w_G4400_1[1]),.dout(n552),.clk(gclk));
	jand g0238(.dina(G226),.dinb(w_G18_45[1]),.dout(n553),.clk(gclk));
	jand g0239(.dina(w_dff_B_7tTp421h9_0),.dinb(w_n355_28[1]),.dout(n554),.clk(gclk));
	jor g0240(.dina(w_n554_0[1]),.dinb(w_dff_B_38xGnxtj6_1),.dout(n555),.clk(gclk));
	jand g0241(.dina(w_n555_1[1]),.dinb(w_n552_0[1]),.dout(n556),.clk(gclk));
	jnot g0242(.din(w_n555_1[0]),.dout(n557),.clk(gclk));
	jand g0243(.dina(n557),.dinb(w_G4400_1[0]),.dout(n558),.clk(gclk));
	jnot g0244(.din(w_n558_0[1]),.dout(n559),.clk(gclk));
	jnot g0245(.din(w_G4394_1[1]),.dout(n560),.clk(gclk));
	jand g0246(.dina(G217),.dinb(w_G18_45[0]),.dout(n561),.clk(gclk));
	jand g0247(.dina(w_dff_B_3iz5PsYf1_0),.dinb(w_n355_28[0]),.dout(n562),.clk(gclk));
	jor g0248(.dina(w_n562_0[1]),.dinb(w_dff_B_5J78YsqT1_1),.dout(n563),.clk(gclk));
	jand g0249(.dina(w_n563_1[1]),.dinb(w_n560_0[1]),.dout(n564),.clk(gclk));
	jand g0250(.dina(w_n564_0[2]),.dinb(n559),.dout(n565),.clk(gclk));
	jor g0251(.dina(w_n565_0[1]),.dinb(w_n556_0[2]),.dout(n566),.clk(gclk));
	jand g0252(.dina(w_n566_0[2]),.dinb(w_dff_B_M54LwU609_1),.dout(n567),.clk(gclk));
	jor g0253(.dina(n567),.dinb(w_n548_0[1]),.dout(n568),.clk(gclk));
	jand g0254(.dina(w_n568_0[2]),.dinb(w_dff_B_FeOV8fMy1_1),.dout(n569),.clk(gclk));
	jor g0255(.dina(n569),.dinb(w_dff_B_iu005BEr3_1),.dout(n570),.clk(gclk));
	jand g0256(.dina(w_n570_1[2]),.dinb(w_dff_B_DkdIHtIg6_1),.dout(n571),.clk(gclk));
	jor g0257(.dina(n571),.dinb(w_dff_B_BEuDBo4u4_1),.dout(n572),.clk(gclk));
	jxor g0258(.dina(w_n531_0[2]),.dinb(w_n528_0[0]),.dout(n573),.clk(gclk));
	jxor g0259(.dina(w_n555_0[2]),.dinb(w_n552_0[0]),.dout(n574),.clk(gclk));
	jxor g0260(.dina(w_n563_1[0]),.dinb(w_n560_0[0]),.dout(n575),.clk(gclk));
	jand g0261(.dina(w_n575_1[1]),.dinb(w_n574_0[2]),.dout(n576),.clk(gclk));
	jxor g0262(.dina(w_n539_0[2]),.dinb(w_n536_0[1]),.dout(n577),.clk(gclk));
	jxor g0263(.dina(w_n547_0[2]),.dinb(w_n544_0[0]),.dout(n578),.clk(gclk));
	jand g0264(.dina(w_n578_0[2]),.dinb(w_n577_0[1]),.dout(n579),.clk(gclk));
	jand g0265(.dina(n579),.dinb(w_n576_0[2]),.dout(n580),.clk(gclk));
	jand g0266(.dina(w_n580_0[2]),.dinb(w_n573_1[1]),.dout(n581),.clk(gclk));
	jnot g0267(.din(w_G3749_0[2]),.dout(n582),.clk(gclk));
	jand g0268(.dina(G231),.dinb(w_G18_44[2]),.dout(n583),.clk(gclk));
	jand g0269(.dina(w_dff_B_M6rCd2HD1_0),.dinb(w_n355_27[2]),.dout(n584),.clk(gclk));
	jor g0270(.dina(w_n584_0[1]),.dinb(w_dff_B_8cvNMGpq8_1),.dout(n585),.clk(gclk));
	jand g0271(.dina(w_n585_1[1]),.dinb(w_n582_0[2]),.dout(n586),.clk(gclk));
	jnot g0272(.din(w_n585_1[0]),.dout(n587),.clk(gclk));
	jand g0273(.dina(n587),.dinb(w_G3749_0[1]),.dout(n588),.clk(gclk));
	jnot g0274(.din(w_n588_0[1]),.dout(n589),.clk(gclk));
	jnot g0275(.din(w_G3743_0[2]),.dout(n590),.clk(gclk));
	jand g0276(.dina(G232),.dinb(w_G18_44[1]),.dout(n591),.clk(gclk));
	jand g0277(.dina(w_dff_B_s7RfLXDr5_0),.dinb(w_n355_27[1]),.dout(n592),.clk(gclk));
	jor g0278(.dina(w_n592_0[1]),.dinb(w_dff_B_wfvo8goK1_1),.dout(n593),.clk(gclk));
	jxor g0279(.dina(w_n593_1[1]),.dinb(w_n590_0[2]),.dout(n594),.clk(gclk));
	jnot g0280(.din(w_G3737_0[2]),.dout(n595),.clk(gclk));
	jand g0281(.dina(G233),.dinb(w_G18_44[0]),.dout(n596),.clk(gclk));
	jand g0282(.dina(w_dff_B_fE0qDrAB4_0),.dinb(w_n355_27[0]),.dout(n597),.clk(gclk));
	jor g0283(.dina(w_n597_0[1]),.dinb(w_dff_B_xjUMoG9V3_1),.dout(n598),.clk(gclk));
	jxor g0284(.dina(w_n598_1[1]),.dinb(w_n595_0[2]),.dout(n599),.clk(gclk));
	jnot g0285(.din(w_G3729_1[1]),.dout(n600),.clk(gclk));
	jand g0286(.dina(G234),.dinb(w_G18_43[2]),.dout(n601),.clk(gclk));
	jand g0287(.dina(w_dff_B_7QV1unCt1_0),.dinb(w_n355_26[2]),.dout(n602),.clk(gclk));
	jor g0288(.dina(w_n602_0[1]),.dinb(w_dff_B_a2pNsB9Y1_1),.dout(n603),.clk(gclk));
	jxor g0289(.dina(w_n603_1[1]),.dinb(w_n600_0[1]),.dout(n604),.clk(gclk));
	jand g0290(.dina(w_n604_0[1]),.dinb(w_n599_0[2]),.dout(n605),.clk(gclk));
	jand g0291(.dina(w_n605_0[2]),.dinb(w_n594_0[2]),.dout(n606),.clk(gclk));
	jnot g0292(.din(n606),.dout(n607),.clk(gclk));
	jnot g0293(.din(w_n593_1[0]),.dout(n608),.clk(gclk));
	jand g0294(.dina(n608),.dinb(w_G3743_0[1]),.dout(n609),.clk(gclk));
	jand g0295(.dina(w_n593_0[2]),.dinb(w_n590_0[1]),.dout(n610),.clk(gclk));
	jnot g0296(.din(w_n610_0[1]),.dout(n611),.clk(gclk));
	jand g0297(.dina(w_n598_1[0]),.dinb(w_n595_0[1]),.dout(n612),.clk(gclk));
	jand g0298(.dina(w_n603_1[0]),.dinb(w_n600_0[0]),.dout(n613),.clk(gclk));
	jand g0299(.dina(w_n613_0[2]),.dinb(w_n599_0[1]),.dout(n614),.clk(gclk));
	jor g0300(.dina(n614),.dinb(w_n612_0[1]),.dout(n615),.clk(gclk));
	jnot g0301(.din(w_n615_0[2]),.dout(n616),.clk(gclk));
	jand g0302(.dina(w_n616_0[1]),.dinb(w_dff_B_hy0ml6fJ9_1),.dout(n617),.clk(gclk));
	jor g0303(.dina(n617),.dinb(w_n609_0[1]),.dout(n618),.clk(gclk));
	jand g0304(.dina(w_n618_0[2]),.dinb(w_dff_B_ZbK3sXt04_1),.dout(n619),.clk(gclk));
	jnot g0305(.din(w_n619_0[2]),.dout(n620),.clk(gclk));
	jnot g0306(.din(w_n618_0[1]),.dout(n621),.clk(gclk));
	jnot g0307(.din(w_G3723_0[2]),.dout(n622),.clk(gclk));
	jand g0308(.dina(G235),.dinb(w_G18_43[1]),.dout(n623),.clk(gclk));
	jand g0309(.dina(w_dff_B_xFCehTzh4_0),.dinb(w_n355_26[1]),.dout(n624),.clk(gclk));
	jor g0310(.dina(w_n624_0[1]),.dinb(w_dff_B_9E1ofxPW9_1),.dout(n625),.clk(gclk));
	jxor g0311(.dina(w_n625_1[1]),.dinb(w_n622_0[2]),.dout(n626),.clk(gclk));
	jnot g0312(.din(w_G3717_0[2]),.dout(n627),.clk(gclk));
	jand g0313(.dina(G236),.dinb(w_G18_43[0]),.dout(n628),.clk(gclk));
	jand g0314(.dina(w_dff_B_q1q8bvml7_0),.dinb(w_n355_26[0]),.dout(n629),.clk(gclk));
	jor g0315(.dina(w_n629_0[1]),.dinb(w_dff_B_pxBIfhne4_1),.dout(n630),.clk(gclk));
	jxor g0316(.dina(w_n630_0[2]),.dinb(w_n627_0[2]),.dout(n631),.clk(gclk));
	jnot g0317(.din(w_G3711_0[1]),.dout(n632),.clk(gclk));
	jand g0318(.dina(G237),.dinb(w_G18_42[2]),.dout(n633),.clk(gclk));
	jand g0319(.dina(w_dff_B_ELLLUtH34_0),.dinb(w_n355_25[2]),.dout(n634),.clk(gclk));
	jor g0320(.dina(w_n634_0[1]),.dinb(w_dff_B_1i2SLdk65_1),.dout(n635),.clk(gclk));
	jxor g0321(.dina(w_n635_1[1]),.dinb(w_n632_1[1]),.dout(n636),.clk(gclk));
	jnot g0322(.din(w_G238_0[1]),.dout(n637),.clk(gclk));
	jor g0323(.dina(n637),.dinb(w_n355_25[1]),.dout(n638),.clk(gclk));
	jnot g0324(.din(w_G29_0[1]),.dout(n639),.clk(gclk));
	jor g0325(.dina(n639),.dinb(w_G18_42[1]),.dout(n640),.clk(gclk));
	jand g0326(.dina(n640),.dinb(n638),.dout(n641),.clk(gclk));
	jxor g0327(.dina(w_n641_0[2]),.dinb(w_G3705_1[2]),.dout(n642),.clk(gclk));
	jand g0328(.dina(w_n642_0[2]),.dinb(w_n359_1[0]),.dout(n643),.clk(gclk));
	jand g0329(.dina(n643),.dinb(w_n636_0[2]),.dout(n644),.clk(gclk));
	jand g0330(.dina(w_n644_0[1]),.dinb(w_n631_0[2]),.dout(n645),.clk(gclk));
	jand g0331(.dina(w_n645_0[1]),.dinb(w_n626_1[1]),.dout(n646),.clk(gclk));
	jand g0332(.dina(w_n625_1[0]),.dinb(w_n622_0[1]),.dout(n647),.clk(gclk));
	jnot g0333(.din(w_n625_0[2]),.dout(n648),.clk(gclk));
	jand g0334(.dina(n648),.dinb(w_G3723_0[1]),.dout(n649),.clk(gclk));
	jnot g0335(.din(w_n649_0[1]),.dout(n650),.clk(gclk));
	jnot g0336(.din(w_n630_0[1]),.dout(n651),.clk(gclk));
	jand g0337(.dina(w_n651_0[1]),.dinb(w_G3717_0[1]),.dout(n652),.clk(gclk));
	jnot g0338(.din(w_n652_0[1]),.dout(n653),.clk(gclk));
	jand g0339(.dina(w_n630_0[0]),.dinb(w_n627_0[1]),.dout(n654),.clk(gclk));
	jand g0340(.dina(w_n635_1[0]),.dinb(w_n632_1[0]),.dout(n655),.clk(gclk));
	jor g0341(.dina(w_n635_0[2]),.dinb(w_n632_0[2]),.dout(n656),.clk(gclk));
	jnot g0342(.din(w_G3705_1[1]),.dout(n657),.clk(gclk));
	jand g0343(.dina(w_G238_0[0]),.dinb(w_G18_42[0]),.dout(n658),.clk(gclk));
	jand g0344(.dina(w_G29_0[0]),.dinb(w_n355_25[0]),.dout(n659),.clk(gclk));
	jor g0345(.dina(w_n659_0[1]),.dinb(w_dff_B_QnNTBcV28_1),.dout(n660),.clk(gclk));
	jor g0346(.dina(w_n660_0[2]),.dinb(w_n657_0[2]),.dout(n661),.clk(gclk));
	jnot g0347(.din(w_G3701_0[2]),.dout(n662),.clk(gclk));
	jand g0348(.dina(w_G41_0[0]),.dinb(w_n355_24[2]),.dout(n663),.clk(gclk));
	jand g0349(.dina(w_n663_1[1]),.dinb(w_n662_0[1]),.dout(n664),.clk(gclk));
	jand g0350(.dina(w_n660_0[1]),.dinb(w_n657_0[1]),.dout(n665),.clk(gclk));
	jor g0351(.dina(n665),.dinb(w_n664_0[1]),.dout(n666),.clk(gclk));
	jand g0352(.dina(w_n666_0[1]),.dinb(w_n661_0[2]),.dout(n667),.clk(gclk));
	jand g0353(.dina(n667),.dinb(w_n656_0[1]),.dout(n668),.clk(gclk));
	jor g0354(.dina(n668),.dinb(w_n655_0[1]),.dout(n669),.clk(gclk));
	jor g0355(.dina(w_n669_0[1]),.dinb(w_n654_0[2]),.dout(n670),.clk(gclk));
	jand g0356(.dina(n670),.dinb(w_n653_0[1]),.dout(n671),.clk(gclk));
	jand g0357(.dina(w_n671_0[1]),.dinb(w_dff_B_C1GdZ4kY1_1),.dout(n672),.clk(gclk));
	jor g0358(.dina(n672),.dinb(w_n647_0[1]),.dout(n673),.clk(gclk));
	jor g0359(.dina(w_n673_0[2]),.dinb(w_n646_0[1]),.dout(n674),.clk(gclk));
	jor g0360(.dina(w_n673_0[1]),.dinb(w_G4526_2[1]),.dout(n675),.clk(gclk));
	jand g0361(.dina(n675),.dinb(w_n674_0[1]),.dout(n676),.clk(gclk));
	jor g0362(.dina(w_n676_0[2]),.dinb(w_dff_B_Ok5coIGX5_1),.dout(n677),.clk(gclk));
	jand g0363(.dina(n677),.dinb(w_dff_B_Sf0ECSPo6_1),.dout(n678),.clk(gclk));
	jand g0364(.dina(w_n678_0[1]),.dinb(w_dff_B_88xv0lQT3_1),.dout(n679),.clk(gclk));
	jor g0365(.dina(n679),.dinb(w_n586_0[2]),.dout(n680),.clk(gclk));
	jand g0366(.dina(w_n680_2[2]),.dinb(w_n581_0[2]),.dout(n681),.clk(gclk));
	jor g0367(.dina(n681),.dinb(w_n572_1[1]),.dout(n682),.clk(gclk));
	jand g0368(.dina(w_n682_0[1]),.dinb(w_dff_B_W33OGnFZ9_1),.dout(n683),.clk(gclk));
	jand g0369(.dina(w_n683_0[1]),.dinb(w_n524_1[2]),.dout(n684),.clk(gclk));
	jand g0370(.dina(n684),.dinb(w_dff_B_mmI1cXgL2_1),.dout(n685),.clk(gclk));
	jand g0371(.dina(n685),.dinb(w_n513_1[1]),.dout(n686),.clk(gclk));
	jand g0372(.dina(w_n512_0[1]),.dinb(w_n509_0[1]),.dout(n687),.clk(gclk));
	jnot g0373(.din(w_n687_0[1]),.dout(n688),.clk(gclk));
	jnot g0374(.din(w_n512_0[0]),.dout(n689),.clk(gclk));
	jand g0375(.dina(w_n689_0[1]),.dinb(w_G4432_0[1]),.dout(n690),.clk(gclk));
	jand g0376(.dina(w_n523_0[1]),.dinb(w_n520_0[0]),.dout(n691),.clk(gclk));
	jand g0377(.dina(w_n524_1[1]),.dinb(w_n518_1[1]),.dout(n692),.clk(gclk));
	jor g0378(.dina(n692),.dinb(w_dff_B_zif2k5jg5_1),.dout(n693),.clk(gclk));
	jnot g0379(.din(w_n693_0[1]),.dout(n694),.clk(gclk));
	jor g0380(.dina(w_n694_0[1]),.dinb(w_n690_0[1]),.dout(n695),.clk(gclk));
	jand g0381(.dina(w_n695_0[1]),.dinb(w_dff_B_gokY1vEq5_1),.dout(n696),.clk(gclk));
	jnot g0382(.din(w_n696_0[1]),.dout(n697),.clk(gclk));
	jor g0383(.dina(w_dff_B_eaqtGupW1_0),.dinb(n686),.dout(n698),.clk(gclk));
	jand g0384(.dina(w_n698_0[1]),.dinb(w_dff_B_WWYGcvMe7_1),.dout(n699),.clk(gclk));
	jor g0385(.dina(n699),.dinb(w_n505_0[1]),.dout(n700),.clk(gclk));
	jor g0386(.dina(w_n700_1[1]),.dinb(w_n462_0[1]),.dout(n701),.clk(gclk));
	jor g0387(.dina(n701),.dinb(w_n500_0[1]),.dout(n702),.clk(gclk));
	jand g0388(.dina(n702),.dinb(w_n499_0[1]),.dout(n703),.clk(gclk));
	jor g0389(.dina(w_n703_1[2]),.dinb(w_n449_1[0]),.dout(n704),.clk(gclk));
	jand g0390(.dina(n704),.dinb(w_n450_0[2]),.dout(n705),.clk(gclk));
	jand g0391(.dina(w_n705_0[1]),.dinb(w_n425_1[1]),.dout(n706),.clk(gclk));
	jor g0392(.dina(n706),.dinb(w_n424_0[1]),.dout(n707),.clk(gclk));
	jor g0393(.dina(w_n707_1[2]),.dinb(w_n413_1[0]),.dout(n708),.clk(gclk));
	jand g0394(.dina(n708),.dinb(w_n420_0[1]),.dout(n709),.clk(gclk));
	jand g0395(.dina(w_n709_1[1]),.dinb(w_n370_0[2]),.dout(n710),.clk(gclk));
	jand g0396(.dina(n710),.dinb(w_n363_0[2]),.dout(n711),.clk(gclk));
	jnot g0397(.din(w_n362_0[1]),.dout(n712),.clk(gclk));
	jand g0398(.dina(w_n712_0[2]),.dinb(w_G38_2[0]),.dout(n713),.clk(gclk));
	jand g0399(.dina(w_n366_0[1]),.dinb(w_G38_1[2]),.dout(n714),.clk(gclk));
	jor g0400(.dina(w_dff_B_dHTH04tO0_0),.dinb(w_n713_0[1]),.dout(n715),.clk(gclk));
	jor g0401(.dina(w_n715_1[1]),.dinb(w_n711_1[1]),.dout(G246),.clk(gclk));
	jand g0402(.dina(w_G2204_0[2]),.dinb(w_G1455_0[2]),.dout(n717),.clk(gclk));
	jor g0403(.dina(w_dff_B_HX5r9EjC7_0),.dinb(w_n368_0[0]),.dout(n718),.clk(gclk));
	jor g0404(.dina(w_dff_B_hwMRptnW4_0),.dinb(w_n355_24[1]),.dout(n719),.clk(gclk));
	jand g0405(.dina(w_n719_0[1]),.dinb(w_n373_6[1]),.dout(n720),.clk(gclk));
	jor g0406(.dina(w_n371_0[0]),.dinb(w_n355_24[0]),.dout(n721),.clk(gclk));
	jor g0407(.dina(G88),.dinb(w_G18_41[2]),.dout(n722),.clk(gclk));
	jand g0408(.dina(w_dff_B_b9rs7CCj0_0),.dinb(n721),.dout(n723),.clk(gclk));
	jxor g0409(.dina(w_n723_0[2]),.dinb(w_n720_0[2]),.dout(n724),.clk(gclk));
	jor g0410(.dina(w_dff_B_DIYmvKh25_0),.dinb(w_n355_23[2]),.dout(n725),.clk(gclk));
	jand g0411(.dina(w_n725_0[1]),.dinb(w_n373_6[0]),.dout(n726),.clk(gclk));
	jor g0412(.dina(w_n383_0[0]),.dinb(w_n355_23[1]),.dout(n727),.clk(gclk));
	jor g0413(.dina(G112),.dinb(w_G18_41[1]),.dout(n728),.clk(gclk));
	jand g0414(.dina(w_dff_B_aRJmjQrm7_0),.dinb(n727),.dout(n729),.clk(gclk));
	jor g0415(.dina(w_n729_1[1]),.dinb(w_n726_1[1]),.dout(n730),.clk(gclk));
	jand g0416(.dina(w_n729_1[0]),.dinb(w_n726_1[0]),.dout(n731),.clk(gclk));
	jor g0417(.dina(w_n389_0[2]),.dinb(w_n355_23[0]),.dout(n732),.clk(gclk));
	jor g0418(.dina(G113),.dinb(w_G18_41[0]),.dout(n733),.clk(gclk));
	jand g0419(.dina(w_dff_B_b4hPWs5V6_0),.dinb(n732),.dout(n734),.clk(gclk));
	jand g0420(.dina(w_n734_0[2]),.dinb(w_n373_5[2]),.dout(n735),.clk(gclk));
	jor g0421(.dina(w_dff_B_9Rdq1LAr7_0),.dinb(w_n355_22[2]),.dout(n736),.clk(gclk));
	jand g0422(.dina(w_n736_0[1]),.dinb(w_n373_5[1]),.dout(n737),.clk(gclk));
	jand g0423(.dina(w_G106_0[2]),.dinb(w_G18_40[2]),.dout(n738),.clk(gclk));
	jnot g0424(.din(n738),.dout(n739),.clk(gclk));
	jor g0425(.dina(G87),.dinb(w_G18_40[1]),.dout(n740),.clk(gclk));
	jand g0426(.dina(w_dff_B_DPX5VXjw8_0),.dinb(n739),.dout(n741),.clk(gclk));
	jxor g0427(.dina(w_n741_1[1]),.dinb(w_n737_1[1]),.dout(n742),.clk(gclk));
	jor g0428(.dina(w_dff_B_w0VPXIFy1_0),.dinb(w_n355_22[1]),.dout(n743),.clk(gclk));
	jand g0429(.dina(w_n743_0[1]),.dinb(w_n373_5[0]),.dout(n744),.clk(gclk));
	jor g0430(.dina(w_n393_0[2]),.dinb(w_n355_22[0]),.dout(n745),.clk(gclk));
	jor g0431(.dina(G111),.dinb(w_G18_40[0]),.dout(n746),.clk(gclk));
	jand g0432(.dina(w_dff_B_6ARVs7Pz3_0),.dinb(n745),.dout(n747),.clk(gclk));
	jxor g0433(.dina(w_n747_0[2]),.dinb(w_n744_0[2]),.dout(n748),.clk(gclk));
	jand g0434(.dina(n748),.dinb(n742),.dout(n749),.clk(gclk));
	jand g0435(.dina(w_n749_0[1]),.dinb(w_dff_B_Dt6dA6I30_1),.dout(n750),.clk(gclk));
	jor g0436(.dina(n750),.dinb(w_dff_B_2G7vtFay6_1),.dout(n751),.clk(gclk));
	jand g0437(.dina(n751),.dinb(w_dff_B_MlLdonTk2_1),.dout(n752),.clk(gclk));
	jand g0438(.dina(n752),.dinb(w_n724_0[1]),.dout(n753),.clk(gclk));
	jor g0439(.dina(w_dff_B_dzW4rya13_0),.dinb(w_n355_21[2]),.dout(n754),.clk(gclk));
	jand g0440(.dina(w_n754_0[1]),.dinb(w_n373_4[2]),.dout(n755),.clk(gclk));
	jor g0441(.dina(w_n421_0[0]),.dinb(w_n355_21[1]),.dout(n756),.clk(gclk));
	jor g0442(.dina(G110),.dinb(w_G18_39[2]),.dout(n757),.clk(gclk));
	jand g0443(.dina(w_dff_B_BLQwtI809_0),.dinb(n756),.dout(n758),.clk(gclk));
	jxor g0444(.dina(w_n758_1[1]),.dinb(w_n755_1[1]),.dout(n759),.clk(gclk));
	jor g0445(.dina(w_dff_B_yAVd0J5N4_0),.dinb(w_n355_21[0]),.dout(n760),.clk(gclk));
	jand g0446(.dina(w_n760_0[1]),.dinb(w_n373_4[1]),.dout(n761),.clk(gclk));
	jor g0447(.dina(w_n426_0[0]),.dinb(w_n355_20[2]),.dout(n762),.clk(gclk));
	jor g0448(.dina(G109),.dinb(w_G18_39[1]),.dout(n763),.clk(gclk));
	jand g0449(.dina(w_dff_B_7UccTtN25_0),.dinb(n762),.dout(n764),.clk(gclk));
	jxor g0450(.dina(w_n764_0[2]),.dinb(w_n761_0[2]),.dout(n765),.clk(gclk));
	jand g0451(.dina(n765),.dinb(n759),.dout(n766),.clk(gclk));
	jor g0452(.dina(w_dff_B_79UrQMsw7_0),.dinb(w_n355_20[1]),.dout(n767),.clk(gclk));
	jand g0453(.dina(w_n767_0[1]),.dinb(w_n373_4[0]),.dout(n768),.clk(gclk));
	jand g0454(.dina(w_G2247_0[1]),.dinb(w_G18_39[0]),.dout(n769),.clk(gclk));
	jnot g0455(.din(n769),.dout(n770),.clk(gclk));
	jor g0456(.dina(G86),.dinb(w_G18_38[2]),.dout(n771),.clk(gclk));
	jand g0457(.dina(w_dff_B_Gu6ly2qK5_0),.dinb(n770),.dout(n772),.clk(gclk));
	jand g0458(.dina(w_n772_0[2]),.dinb(w_n768_0[2]),.dout(n773),.clk(gclk));
	jor g0459(.dina(w_n772_0[1]),.dinb(w_n768_0[1]),.dout(n774),.clk(gclk));
	jor g0460(.dina(w_dff_B_m3XKlcFu2_0),.dinb(w_n355_20[0]),.dout(n775),.clk(gclk));
	jand g0461(.dina(w_n775_0[1]),.dinb(w_n373_3[2]),.dout(n776),.clk(gclk));
	jand g0462(.dina(w_G2239_1[0]),.dinb(w_G18_38[1]),.dout(n777),.clk(gclk));
	jnot g0463(.din(n777),.dout(n778),.clk(gclk));
	jor g0464(.dina(G63),.dinb(w_G18_38[0]),.dout(n779),.clk(gclk));
	jand g0465(.dina(w_dff_B_IEzZQimm6_0),.dinb(n778),.dout(n780),.clk(gclk));
	jand g0466(.dina(w_n780_0[2]),.dinb(w_n776_0[2]),.dout(n781),.clk(gclk));
	jand g0467(.dina(w_n781_0[1]),.dinb(w_n774_0[1]),.dout(n782),.clk(gclk));
	jor g0468(.dina(n782),.dinb(w_n773_0[1]),.dout(n783),.clk(gclk));
	jand g0469(.dina(n783),.dinb(w_n766_0[1]),.dout(n784),.clk(gclk));
	jand g0470(.dina(w_n758_1[0]),.dinb(w_n755_1[0]),.dout(n785),.clk(gclk));
	jor g0471(.dina(w_n758_0[2]),.dinb(w_n755_0[2]),.dout(n786),.clk(gclk));
	jand g0472(.dina(w_n764_0[1]),.dinb(w_n761_0[1]),.dout(n787),.clk(gclk));
	jand g0473(.dina(n787),.dinb(n786),.dout(n788),.clk(gclk));
	jor g0474(.dina(n788),.dinb(w_dff_B_O1JLdrLw2_1),.dout(n789),.clk(gclk));
	jor g0475(.dina(w_dff_B_Ddj01x9g8_0),.dinb(n784),.dout(n790),.clk(gclk));
	jnot g0476(.din(w_n773_0[0]),.dout(n791),.clk(gclk));
	jnot g0477(.din(w_n781_0[0]),.dout(n792),.clk(gclk));
	jand g0478(.dina(n792),.dinb(n791),.dout(n793),.clk(gclk));
	jand g0479(.dina(n793),.dinb(w_n766_0[0]),.dout(n794),.clk(gclk));
	jor g0480(.dina(w_dff_B_zHUjpYCt9_0),.dinb(w_n355_19[2]),.dout(n795),.clk(gclk));
	jand g0481(.dina(n795),.dinb(w_n373_3[1]),.dout(n796),.clk(gclk));
	jand g0482(.dina(w_G2236_0[1]),.dinb(w_G18_37[2]),.dout(n797),.clk(gclk));
	jnot g0483(.din(n797),.dout(n798),.clk(gclk));
	jor g0484(.dina(G64),.dinb(w_G18_37[1]),.dout(n799),.clk(gclk));
	jand g0485(.dina(w_dff_B_9QxBzGL67_0),.dinb(n798),.dout(n800),.clk(gclk));
	jxor g0486(.dina(w_n800_1[1]),.dinb(w_n796_1[1]),.dout(n801),.clk(gclk));
	jand g0487(.dina(G178),.dinb(w_G18_37[0]),.dout(n802),.clk(gclk));
	jor g0488(.dina(w_dff_B_DMptHjD75_0),.dinb(w_n457_0[0]),.dout(n803),.clk(gclk));
	jor g0489(.dina(w_n456_0[0]),.dinb(w_n355_19[1]),.dout(n804),.clk(gclk));
	jor g0490(.dina(G85),.dinb(w_G18_36[2]),.dout(n805),.clk(gclk));
	jand g0491(.dina(w_dff_B_cJHpgVha7_0),.dinb(n804),.dout(n806),.clk(gclk));
	jxor g0492(.dina(w_n806_0[2]),.dinb(w_n803_0[2]),.dout(n807),.clk(gclk));
	jand g0493(.dina(n807),.dinb(n801),.dout(n808),.clk(gclk));
	jand g0494(.dina(G179),.dinb(w_G18_36[1]),.dout(n809),.clk(gclk));
	jor g0495(.dina(w_dff_B_QrpMF2wn8_0),.dinb(w_n467_0[0]),.dout(n810),.clk(gclk));
	jand g0496(.dina(w_G2224_0[2]),.dinb(w_G18_36[0]),.dout(n811),.clk(gclk));
	jnot g0497(.din(n811),.dout(n812),.clk(gclk));
	jor g0498(.dina(G84),.dinb(w_G18_35[2]),.dout(n813),.clk(gclk));
	jand g0499(.dina(w_dff_B_6C2O4IGp8_0),.dinb(n812),.dout(n814),.clk(gclk));
	jxor g0500(.dina(w_n814_1[1]),.dinb(w_n810_1[1]),.dout(n815),.clk(gclk));
	jand g0501(.dina(G180),.dinb(w_G18_35[1]),.dout(n816),.clk(gclk));
	jor g0502(.dina(w_dff_B_RJRmwaaI4_0),.dinb(w_n472_0[0]),.dout(n817),.clk(gclk));
	jor g0503(.dina(w_n471_0[0]),.dinb(w_n355_19[0]),.dout(n818),.clk(gclk));
	jor g0504(.dina(G83),.dinb(w_G18_35[0]),.dout(n819),.clk(gclk));
	jand g0505(.dina(w_dff_B_jP0SD0ms6_0),.dinb(n818),.dout(n820),.clk(gclk));
	jxor g0506(.dina(w_n820_0[2]),.dinb(w_n817_0[2]),.dout(n821),.clk(gclk));
	jand g0507(.dina(n821),.dinb(n815),.dout(n822),.clk(gclk));
	jand g0508(.dina(G171),.dinb(w_G18_34[2]),.dout(n823),.clk(gclk));
	jor g0509(.dina(w_dff_B_xys7zFVf2_0),.dinb(w_n477_0[0]),.dout(n824),.clk(gclk));
	jor g0510(.dina(w_n476_0[0]),.dinb(w_n355_18[2]),.dout(n825),.clk(gclk));
	jor g0511(.dina(G65),.dinb(w_G18_34[1]),.dout(n826),.clk(gclk));
	jand g0512(.dina(w_dff_B_pJwGi2Fx0_0),.dinb(n825),.dout(n827),.clk(gclk));
	jand g0513(.dina(w_n827_0[2]),.dinb(w_n824_0[2]),.dout(n828),.clk(gclk));
	jand g0514(.dina(w_dff_B_9aw3Afxr6_0),.dinb(w_n822_0[1]),.dout(n829),.clk(gclk));
	jand g0515(.dina(w_n814_1[0]),.dinb(w_n810_1[0]),.dout(n830),.clk(gclk));
	jor g0516(.dina(w_n814_0[2]),.dinb(w_n810_0[2]),.dout(n831),.clk(gclk));
	jand g0517(.dina(w_n820_0[1]),.dinb(w_n817_0[1]),.dout(n832),.clk(gclk));
	jand g0518(.dina(n832),.dinb(n831),.dout(n833),.clk(gclk));
	jor g0519(.dina(n833),.dinb(w_dff_B_FWBTaxcO4_1),.dout(n834),.clk(gclk));
	jor g0520(.dina(n834),.dinb(n829),.dout(n835),.clk(gclk));
	jand g0521(.dina(n835),.dinb(w_n808_0[1]),.dout(n836),.clk(gclk));
	jand g0522(.dina(w_n800_1[0]),.dinb(w_n796_1[0]),.dout(n837),.clk(gclk));
	jor g0523(.dina(w_n800_0[2]),.dinb(w_n796_0[2]),.dout(n838),.clk(gclk));
	jand g0524(.dina(w_n806_0[1]),.dinb(w_n803_0[1]),.dout(n839),.clk(gclk));
	jand g0525(.dina(n839),.dinb(n838),.dout(n840),.clk(gclk));
	jor g0526(.dina(n840),.dinb(w_dff_B_yE5DwyML5_1),.dout(n841),.clk(gclk));
	jor g0527(.dina(w_dff_B_zMHrUpc90_0),.dinb(n836),.dout(n842),.clk(gclk));
	jand g0528(.dina(w_n822_0[0]),.dinb(w_n808_0[0]),.dout(n843),.clk(gclk));
	jand g0529(.dina(G189),.dinb(w_G18_34[0]),.dout(n844),.clk(gclk));
	jor g0530(.dina(w_dff_B_XImWSt9X0_0),.dinb(w_n503_0[0]),.dout(n845),.clk(gclk));
	jor g0531(.dina(w_n501_0[1]),.dinb(w_n355_18[1]),.dout(n846),.clk(gclk));
	jor g0532(.dina(G62),.dinb(w_G18_33[2]),.dout(n847),.clk(gclk));
	jand g0533(.dina(w_dff_B_E6bjujDE2_0),.dinb(n846),.dout(n848),.clk(gclk));
	jxor g0534(.dina(w_n848_1[1]),.dinb(w_n845_1[1]),.dout(n849),.clk(gclk));
	jand g0535(.dina(G190),.dinb(w_G18_33[1]),.dout(n850),.clk(gclk));
	jor g0536(.dina(w_dff_B_LU0uSKLW4_0),.dinb(w_n511_0[0]),.dout(n851),.clk(gclk));
	jor g0537(.dina(w_n509_0[0]),.dinb(w_n355_18[0]),.dout(n852),.clk(gclk));
	jor g0538(.dina(G61),.dinb(w_G18_33[0]),.dout(n853),.clk(gclk));
	jand g0539(.dina(w_dff_B_bOdZZeZW2_0),.dinb(n852),.dout(n854),.clk(gclk));
	jxor g0540(.dina(w_n854_0[2]),.dinb(w_n851_0[2]),.dout(n855),.clk(gclk));
	jand g0541(.dina(n855),.dinb(n849),.dout(n856),.clk(gclk));
	jand g0542(.dina(G191),.dinb(w_G18_32[2]),.dout(n857),.clk(gclk));
	jor g0543(.dina(w_dff_B_tSwZ6JNW4_0),.dinb(w_n522_0[0]),.dout(n858),.clk(gclk));
	jand g0544(.dina(w_G4427_0[1]),.dinb(w_G18_32[1]),.dout(n859),.clk(gclk));
	jnot g0545(.din(n859),.dout(n860),.clk(gclk));
	jor g0546(.dina(G60),.dinb(w_G18_32[0]),.dout(n861),.clk(gclk));
	jand g0547(.dina(w_dff_B_USso0eYK3_0),.dinb(n860),.dout(n862),.clk(gclk));
	jand g0548(.dina(w_n862_0[2]),.dinb(w_n858_0[2]),.dout(n863),.clk(gclk));
	jor g0549(.dina(w_n862_0[1]),.dinb(w_n858_0[1]),.dout(n864),.clk(gclk));
	jand g0550(.dina(G192),.dinb(w_G18_31[2]),.dout(n865),.clk(gclk));
	jor g0551(.dina(w_dff_B_V5tqYNKC5_0),.dinb(w_n516_0[0]),.dout(n866),.clk(gclk));
	jand g0552(.dina(w_G4420_0[2]),.dinb(w_G18_31[1]),.dout(n867),.clk(gclk));
	jnot g0553(.din(n867),.dout(n868),.clk(gclk));
	jor g0554(.dina(G79),.dinb(w_G18_31[0]),.dout(n869),.clk(gclk));
	jand g0555(.dina(w_dff_B_nLQv1jO69_0),.dinb(n868),.dout(n870),.clk(gclk));
	jand g0556(.dina(w_n870_0[2]),.dinb(w_n866_0[2]),.dout(n871),.clk(gclk));
	jand g0557(.dina(w_n871_0[1]),.dinb(w_n864_0[1]),.dout(n872),.clk(gclk));
	jor g0558(.dina(n872),.dinb(w_n863_0[1]),.dout(n873),.clk(gclk));
	jand g0559(.dina(n873),.dinb(w_n856_0[1]),.dout(n874),.clk(gclk));
	jand g0560(.dina(w_n848_1[0]),.dinb(w_n845_1[0]),.dout(n875),.clk(gclk));
	jor g0561(.dina(w_n848_0[2]),.dinb(w_n845_0[2]),.dout(n876),.clk(gclk));
	jand g0562(.dina(w_n854_0[1]),.dinb(w_n851_0[1]),.dout(n877),.clk(gclk));
	jand g0563(.dina(n877),.dinb(n876),.dout(n878),.clk(gclk));
	jor g0564(.dina(n878),.dinb(w_dff_B_XLgbErkX1_1),.dout(n879),.clk(gclk));
	jor g0565(.dina(w_dff_B_gEZBHIQa1_0),.dinb(n874),.dout(n880),.clk(gclk));
	jor g0566(.dina(w_n870_0[1]),.dinb(w_n866_0[1]),.dout(n881),.clk(gclk));
	jand g0567(.dina(n881),.dinb(w_n864_0[0]),.dout(n882),.clk(gclk));
	jand g0568(.dina(n882),.dinb(w_n856_0[0]),.dout(n883),.clk(gclk));
	jand g0569(.dina(G205),.dinb(w_G18_30[2]),.dout(n884),.clk(gclk));
	jor g0570(.dina(w_dff_B_eOJ5LWf19_0),.dinb(w_n629_0[0]),.dout(n885),.clk(gclk));
	jor g0571(.dina(w_n627_0[0]),.dinb(w_n355_17[2]),.dout(n886),.clk(gclk));
	jor g0572(.dina(G75),.dinb(w_G18_30[1]),.dout(n887),.clk(gclk));
	jand g0573(.dina(w_dff_B_RMyClBpC5_0),.dinb(n886),.dout(n888),.clk(gclk));
	jor g0574(.dina(w_n888_0[2]),.dinb(w_n885_0[2]),.dout(n889),.clk(gclk));
	jand g0575(.dina(G206),.dinb(w_G18_30[0]),.dout(n890),.clk(gclk));
	jor g0576(.dina(w_dff_B_ljr0nkmZ3_0),.dinb(w_n634_0[0]),.dout(n891),.clk(gclk));
	jor g0577(.dina(w_n632_0[1]),.dinb(w_n355_17[1]),.dout(n892),.clk(gclk));
	jor g0578(.dina(G76),.dinb(w_G18_29[2]),.dout(n893),.clk(gclk));
	jand g0579(.dina(w_dff_B_0KB6iv9g0_0),.dinb(n892),.dout(n894),.clk(gclk));
	jand g0580(.dina(w_n894_0[2]),.dinb(w_n891_0[2]),.dout(n895),.clk(gclk));
	jor g0581(.dina(w_G89_0[1]),.dinb(w_G70_0[1]),.dout(n896),.clk(gclk));
	jand g0582(.dina(w_dff_B_BlvzTLvr5_0),.dinb(w_n663_1[0]),.dout(n897),.clk(gclk));
	jor g0583(.dina(w_dff_B_wzfHBs9Y7_0),.dinb(w_n895_0[1]),.dout(n898),.clk(gclk));
	jand g0584(.dina(G207),.dinb(w_G18_29[1]),.dout(n899),.clk(gclk));
	jor g0585(.dina(w_dff_B_v55vyGEp0_0),.dinb(w_n659_0[0]),.dout(n900),.clk(gclk));
	jor g0586(.dina(w_n657_0[0]),.dinb(w_n355_17[0]),.dout(n901),.clk(gclk));
	jor g0587(.dina(G74),.dinb(w_G18_29[0]),.dout(n902),.clk(gclk));
	jand g0588(.dina(w_dff_B_rVfVfTqS2_0),.dinb(n901),.dout(n903),.clk(gclk));
	jand g0589(.dina(w_n903_0[2]),.dinb(w_n900_0[2]),.dout(n904),.clk(gclk));
	jor g0590(.dina(w_G70_0[0]),.dinb(w_G18_28[2]),.dout(n905),.clk(gclk));
	jand g0591(.dina(w_n905_0[1]),.dinb(w_G89_0[0]),.dout(n906),.clk(gclk));
	jor g0592(.dina(w_dff_B_Z1KLiv0J5_0),.dinb(n904),.dout(n907),.clk(gclk));
	jor g0593(.dina(n907),.dinb(n898),.dout(n908),.clk(gclk));
	jor g0594(.dina(w_n903_0[1]),.dinb(w_n900_0[1]),.dout(n909),.clk(gclk));
	jor g0595(.dina(w_n894_0[1]),.dinb(w_n891_0[1]),.dout(n910),.clk(gclk));
	jand g0596(.dina(n910),.dinb(n909),.dout(n911),.clk(gclk));
	jor g0597(.dina(n911),.dinb(w_n895_0[0]),.dout(n912),.clk(gclk));
	jand g0598(.dina(n912),.dinb(n908),.dout(n913),.clk(gclk));
	jand g0599(.dina(n913),.dinb(w_dff_B_DUUq7Zzj9_1),.dout(n914),.clk(gclk));
	jand g0600(.dina(G204),.dinb(w_G18_28[1]),.dout(n915),.clk(gclk));
	jor g0601(.dina(w_dff_B_qaOf45IT1_0),.dinb(w_n624_0[0]),.dout(n916),.clk(gclk));
	jor g0602(.dina(w_n622_0[0]),.dinb(w_n355_16[2]),.dout(n917),.clk(gclk));
	jor g0603(.dina(G73),.dinb(w_G18_28[0]),.dout(n918),.clk(gclk));
	jand g0604(.dina(w_dff_B_ECjMh99R0_0),.dinb(n917),.dout(n919),.clk(gclk));
	jand g0605(.dina(w_n919_0[2]),.dinb(w_n916_0[2]),.dout(n920),.clk(gclk));
	jand g0606(.dina(w_n888_0[1]),.dinb(w_n885_0[1]),.dout(n921),.clk(gclk));
	jor g0607(.dina(n921),.dinb(n920),.dout(n922),.clk(gclk));
	jor g0608(.dina(w_dff_B_vgFcF65u4_0),.dinb(n914),.dout(n923),.clk(gclk));
	jor g0609(.dina(w_n919_0[1]),.dinb(w_n916_0[1]),.dout(n924),.clk(gclk));
	jand g0610(.dina(G203),.dinb(w_G18_27[2]),.dout(n925),.clk(gclk));
	jor g0611(.dina(w_dff_B_uZxkjb4b3_0),.dinb(w_n602_0[0]),.dout(n926),.clk(gclk));
	jand g0612(.dina(w_G3729_1[0]),.dinb(w_G18_27[1]),.dout(n927),.clk(gclk));
	jnot g0613(.din(n927),.dout(n928),.clk(gclk));
	jor g0614(.dina(G53),.dinb(w_G18_27[0]),.dout(n929),.clk(gclk));
	jand g0615(.dina(w_dff_B_XrjS3DjW1_0),.dinb(n928),.dout(n930),.clk(gclk));
	jor g0616(.dina(w_n930_0[2]),.dinb(w_n926_0[2]),.dout(n931),.clk(gclk));
	jand g0617(.dina(n931),.dinb(n924),.dout(n932),.clk(gclk));
	jand g0618(.dina(w_dff_B_D3MvhOYV3_0),.dinb(n923),.dout(n933),.clk(gclk));
	jand g0619(.dina(G202),.dinb(w_G18_26[2]),.dout(n934),.clk(gclk));
	jor g0620(.dina(w_dff_B_XkSaNPgG2_0),.dinb(w_n597_0[0]),.dout(n935),.clk(gclk));
	jor g0621(.dina(w_n595_0[0]),.dinb(w_n355_16[1]),.dout(n936),.clk(gclk));
	jor g0622(.dina(G54),.dinb(w_G18_26[1]),.dout(n937),.clk(gclk));
	jand g0623(.dina(w_dff_B_89Ljj37K2_0),.dinb(n936),.dout(n938),.clk(gclk));
	jand g0624(.dina(w_n938_0[2]),.dinb(w_n935_0[2]),.dout(n939),.clk(gclk));
	jand g0625(.dina(w_n930_0[1]),.dinb(w_n926_0[1]),.dout(n940),.clk(gclk));
	jor g0626(.dina(n940),.dinb(n939),.dout(n941),.clk(gclk));
	jor g0627(.dina(w_dff_B_EAGu5l770_0),.dinb(n933),.dout(n942),.clk(gclk));
	jand g0628(.dina(G201),.dinb(w_G18_26[0]),.dout(n943),.clk(gclk));
	jor g0629(.dina(w_dff_B_YnrrQu3O9_0),.dinb(w_n592_0[0]),.dout(n944),.clk(gclk));
	jor g0630(.dina(w_n590_0[0]),.dinb(w_n355_16[0]),.dout(n945),.clk(gclk));
	jor g0631(.dina(G55),.dinb(w_G18_25[2]),.dout(n946),.clk(gclk));
	jand g0632(.dina(w_dff_B_aZGGt5d13_0),.dinb(n945),.dout(n947),.clk(gclk));
	jxor g0633(.dina(w_n947_0[2]),.dinb(w_n944_0[2]),.dout(n948),.clk(gclk));
	jand g0634(.dina(G200),.dinb(w_G18_25[1]),.dout(n949),.clk(gclk));
	jor g0635(.dina(w_dff_B_emtolqjk2_0),.dinb(w_n584_0[0]),.dout(n950),.clk(gclk));
	jor g0636(.dina(w_n582_0[1]),.dinb(w_n355_15[2]),.dout(n951),.clk(gclk));
	jor g0637(.dina(G56),.dinb(w_G18_25[0]),.dout(n952),.clk(gclk));
	jand g0638(.dina(w_dff_B_n52irTqO9_0),.dinb(n951),.dout(n953),.clk(gclk));
	jxor g0639(.dina(w_n953_1[1]),.dinb(w_n950_1[1]),.dout(n954),.clk(gclk));
	jand g0640(.dina(n954),.dinb(n948),.dout(n955),.clk(gclk));
	jor g0641(.dina(w_n938_0[1]),.dinb(w_n935_0[1]),.dout(n956),.clk(gclk));
	jand g0642(.dina(w_dff_B_JueNAneB1_0),.dinb(n955),.dout(n957),.clk(gclk));
	jand g0643(.dina(w_dff_B_Z1wa6H460_0),.dinb(n942),.dout(n958),.clk(gclk));
	jand g0644(.dina(w_n953_1[0]),.dinb(w_n950_1[0]),.dout(n959),.clk(gclk));
	jand g0645(.dina(w_n947_0[1]),.dinb(w_n944_0[1]),.dout(n960),.clk(gclk));
	jor g0646(.dina(w_n953_0[2]),.dinb(w_n950_0[2]),.dout(n961),.clk(gclk));
	jand g0647(.dina(n961),.dinb(n960),.dout(n962),.clk(gclk));
	jor g0648(.dina(n962),.dinb(w_dff_B_HKXq822L7_1),.dout(n963),.clk(gclk));
	jor g0649(.dina(w_dff_B_nwKB96Tv8_0),.dinb(n958),.dout(n964),.clk(gclk));
	jand g0650(.dina(G187),.dinb(w_G18_24[2]),.dout(n965),.clk(gclk));
	jor g0651(.dina(w_dff_B_DKVgnHfT6_0),.dinb(w_n562_0[0]),.dout(n966),.clk(gclk));
	jand g0652(.dina(w_G4394_1[0]),.dinb(w_G18_24[1]),.dout(n967),.clk(gclk));
	jnot g0653(.din(n967),.dout(n968),.clk(gclk));
	jor g0654(.dina(G77),.dinb(w_G18_24[0]),.dout(n969),.clk(gclk));
	jand g0655(.dina(w_dff_B_XtbsRcWL8_0),.dinb(n968),.dout(n970),.clk(gclk));
	jor g0656(.dina(w_n970_0[2]),.dinb(w_n966_0[2]),.dout(n971),.clk(gclk));
	jand g0657(.dina(G193),.dinb(w_G18_23[2]),.dout(n972),.clk(gclk));
	jor g0658(.dina(w_dff_B_yv5Uv9zV8_0),.dinb(w_n530_0[0]),.dout(n973),.clk(gclk));
	jand g0659(.dina(w_G4415_0[2]),.dinb(w_G18_23[1]),.dout(n974),.clk(gclk));
	jnot g0660(.din(n974),.dout(n975),.clk(gclk));
	jor g0661(.dina(G80),.dinb(w_G18_23[0]),.dout(n976),.clk(gclk));
	jand g0662(.dina(w_dff_B_V6haeHWd2_0),.dinb(n975),.dout(n977),.clk(gclk));
	jxor g0663(.dina(w_n977_1[1]),.dinb(w_n973_1[1]),.dout(n978),.clk(gclk));
	jand g0664(.dina(G194),.dinb(w_G18_22[2]),.dout(n979),.clk(gclk));
	jor g0665(.dina(w_dff_B_ms9OW3LG2_0),.dinb(w_n538_0[0]),.dout(n980),.clk(gclk));
	jor g0666(.dina(w_n536_0[0]),.dinb(w_n355_15[1]),.dout(n981),.clk(gclk));
	jor g0667(.dina(G81),.dinb(w_G18_22[1]),.dout(n982),.clk(gclk));
	jand g0668(.dina(w_dff_B_p0CF3ola8_0),.dinb(n981),.dout(n983),.clk(gclk));
	jxor g0669(.dina(w_n983_0[2]),.dinb(w_n980_0[2]),.dout(n984),.clk(gclk));
	jand g0670(.dina(n984),.dinb(n978),.dout(n985),.clk(gclk));
	jand g0671(.dina(G196),.dinb(w_G18_22[0]),.dout(n986),.clk(gclk));
	jor g0672(.dina(w_dff_B_JsIfzC3e0_0),.dinb(w_n554_0[0]),.dout(n987),.clk(gclk));
	jand g0673(.dina(w_G4400_0[2]),.dinb(w_G18_21[2]),.dout(n988),.clk(gclk));
	jnot g0674(.din(n988),.dout(n989),.clk(gclk));
	jor g0675(.dina(G78),.dinb(w_G18_21[1]),.dout(n990),.clk(gclk));
	jand g0676(.dina(w_dff_B_xDZu6nOM6_0),.dinb(n989),.dout(n991),.clk(gclk));
	jand g0677(.dina(w_n991_0[2]),.dinb(w_n987_0[2]),.dout(n992),.clk(gclk));
	jnot g0678(.din(w_n992_0[1]),.dout(n993),.clk(gclk));
	jand g0679(.dina(G195),.dinb(w_G18_21[0]),.dout(n994),.clk(gclk));
	jor g0680(.dina(w_dff_B_MikmA2wz1_0),.dinb(w_n546_0[0]),.dout(n995),.clk(gclk));
	jand g0681(.dina(w_G4405_0[2]),.dinb(w_G18_20[2]),.dout(n996),.clk(gclk));
	jnot g0682(.din(n996),.dout(n997),.clk(gclk));
	jor g0683(.dina(G59),.dinb(w_G18_20[1]),.dout(n998),.clk(gclk));
	jand g0684(.dina(w_dff_B_W4jNgWOn8_0),.dinb(n997),.dout(n999),.clk(gclk));
	jor g0685(.dina(w_n999_0[2]),.dinb(w_n995_0[2]),.dout(n1000),.clk(gclk));
	jand g0686(.dina(w_n1000_0[1]),.dinb(n993),.dout(n1001),.clk(gclk));
	jor g0687(.dina(w_n991_0[1]),.dinb(w_n987_0[1]),.dout(n1002),.clk(gclk));
	jand g0688(.dina(w_n999_0[1]),.dinb(w_n995_0[1]),.dout(n1003),.clk(gclk));
	jnot g0689(.din(w_n1003_0[1]),.dout(n1004),.clk(gclk));
	jand g0690(.dina(n1004),.dinb(w_dff_B_3gV6bLg16_1),.dout(n1005),.clk(gclk));
	jand g0691(.dina(n1005),.dinb(n1001),.dout(n1006),.clk(gclk));
	jand g0692(.dina(n1006),.dinb(w_n985_0[1]),.dout(n1007),.clk(gclk));
	jand g0693(.dina(w_n970_0[1]),.dinb(w_n966_0[1]),.dout(n1008),.clk(gclk));
	jnot g0694(.din(w_n1008_0[1]),.dout(n1009),.clk(gclk));
	jand g0695(.dina(w_dff_B_TLv5oiTp8_0),.dinb(w_n1007_0[1]),.dout(n1010),.clk(gclk));
	jand g0696(.dina(n1010),.dinb(w_dff_B_BkNagHHh6_1),.dout(n1011),.clk(gclk));
	jand g0697(.dina(w_dff_B_XuQVTKfc1_0),.dinb(n964),.dout(n1012),.clk(gclk));
	jand g0698(.dina(w_n977_1[0]),.dinb(w_n973_1[0]),.dout(n1013),.clk(gclk));
	jor g0699(.dina(w_n977_0[2]),.dinb(w_n973_0[2]),.dout(n1014),.clk(gclk));
	jand g0700(.dina(w_n983_0[1]),.dinb(w_n980_0[1]),.dout(n1015),.clk(gclk));
	jand g0701(.dina(n1015),.dinb(n1014),.dout(n1016),.clk(gclk));
	jor g0702(.dina(n1016),.dinb(w_dff_B_T6Uv8ky34_1),.dout(n1017),.clk(gclk));
	jand g0703(.dina(w_n1008_0[0]),.dinb(w_n1007_0[0]),.dout(n1018),.clk(gclk));
	jand g0704(.dina(w_n1000_0[0]),.dinb(w_n992_0[0]),.dout(n1019),.clk(gclk));
	jor g0705(.dina(n1019),.dinb(w_n1003_0[0]),.dout(n1020),.clk(gclk));
	jand g0706(.dina(n1020),.dinb(w_n985_0[0]),.dout(n1021),.clk(gclk));
	jor g0707(.dina(w_dff_B_A6CLlKNI3_0),.dinb(n1018),.dout(n1022),.clk(gclk));
	jor g0708(.dina(n1022),.dinb(w_dff_B_lDVCWs0x5_1),.dout(n1023),.clk(gclk));
	jor g0709(.dina(w_dff_B_jnT5tqD47_0),.dinb(n1012),.dout(n1024),.clk(gclk));
	jnot g0710(.din(w_n863_0[0]),.dout(n1025),.clk(gclk));
	jnot g0711(.din(w_n871_0[0]),.dout(n1026),.clk(gclk));
	jand g0712(.dina(n1026),.dinb(n1025),.dout(n1027),.clk(gclk));
	jand g0713(.dina(w_dff_B_0Tk8qq6q4_0),.dinb(n1024),.dout(n1028),.clk(gclk));
	jand g0714(.dina(n1028),.dinb(w_dff_B_Y4vEEvQ13_1),.dout(n1029),.clk(gclk));
	jor g0715(.dina(n1029),.dinb(w_dff_B_1JamPVks3_1),.dout(G252_fa_),.clk(gclk));
	jxor g0716(.dina(w_n827_0[1]),.dinb(w_n824_0[1]),.dout(n1031),.clk(gclk));
	jand g0717(.dina(w_dff_B_AdyRxg5x1_0),.dinb(w_G252_0),.dout(n1032),.clk(gclk));
	jand g0718(.dina(n1032),.dinb(w_dff_B_VFnSsohA1_1),.dout(n1033),.clk(gclk));
	jor g0719(.dina(n1033),.dinb(w_dff_B_CXoIoVTw8_1),.dout(n1034),.clk(gclk));
	jor g0720(.dina(w_n780_0[1]),.dinb(w_n776_0[1]),.dout(n1035),.clk(gclk));
	jand g0721(.dina(n1035),.dinb(w_n774_0[0]),.dout(n1036),.clk(gclk));
	jand g0722(.dina(w_dff_B_ZwTl6rAk0_0),.dinb(n1034),.dout(n1037),.clk(gclk));
	jand g0723(.dina(n1037),.dinb(w_dff_B_2GmbTt8p1_1),.dout(n1038),.clk(gclk));
	jor g0724(.dina(n1038),.dinb(w_dff_B_XhyAd35E2_1),.dout(n1039),.clk(gclk));
	jxor g0725(.dina(w_n734_0[1]),.dinb(w_n373_3[0]),.dout(n1040),.clk(gclk));
	jxor g0726(.dina(w_n729_0[2]),.dinb(w_n726_0[2]),.dout(n1041),.clk(gclk));
	jand g0727(.dina(n1041),.dinb(w_n724_0[0]),.dout(n1042),.clk(gclk));
	jand g0728(.dina(w_n1042_0[1]),.dinb(w_n749_0[0]),.dout(n1043),.clk(gclk));
	jand g0729(.dina(n1043),.dinb(w_dff_B_4WtbBNc87_1),.dout(n1044),.clk(gclk));
	jand g0730(.dina(w_dff_B_ZR0Rcscs5_0),.dinb(n1039),.dout(n1045),.clk(gclk));
	jor g0731(.dina(w_G2204_0[1]),.dinb(w_G1455_0[1]),.dout(n1046),.clk(gclk));
	jor g0732(.dina(n1046),.dinb(w_n367_0[0]),.dout(n1047),.clk(gclk));
	jand g0733(.dina(n1047),.dinb(w_G38_1[1]),.dout(n1048),.clk(gclk));
	jand g0734(.dina(w_n723_0[1]),.dinb(w_n720_0[1]),.dout(n1049),.clk(gclk));
	jand g0735(.dina(w_n741_1[0]),.dinb(w_n737_1[0]),.dout(n1050),.clk(gclk));
	jor g0736(.dina(w_n741_0[2]),.dinb(w_n737_0[2]),.dout(n1051),.clk(gclk));
	jand g0737(.dina(w_n747_0[1]),.dinb(w_n744_0[1]),.dout(n1052),.clk(gclk));
	jand g0738(.dina(n1052),.dinb(n1051),.dout(n1053),.clk(gclk));
	jor g0739(.dina(n1053),.dinb(w_dff_B_gHZo3aqe3_1),.dout(n1054),.clk(gclk));
	jand g0740(.dina(n1054),.dinb(w_n1042_0[0]),.dout(n1055),.clk(gclk));
	jor g0741(.dina(n1055),.dinb(w_dff_B_Mu0xTX3i7_1),.dout(n1056),.clk(gclk));
	jor g0742(.dina(n1056),.dinb(w_dff_B_qkNvFZIn9_1),.dout(n1057),.clk(gclk));
	jor g0743(.dina(w_dff_B_mjsGBemm5_0),.dinb(n1045),.dout(n1058),.clk(gclk));
	jor g0744(.dina(n1058),.dinb(w_dff_B_QEsPxDpC0_1),.dout(n1059),.clk(gclk));
	jand g0745(.dina(w_n1059_0[2]),.dinb(w_n718_0[2]),.dout(w_dff_A_ajNjXzv73_2),.clk(gclk));
	jnot g0746(.din(w_n644_0[0]),.dout(n1061),.clk(gclk));
	jnot g0747(.din(w_n655_0[0]),.dout(n1062),.clk(gclk));
	jnot g0748(.din(w_n656_0[0]),.dout(n1063),.clk(gclk));
	jand g0749(.dina(w_n641_0[1]),.dinb(w_G3705_1[0]),.dout(n1064),.clk(gclk));
	jor g0750(.dina(w_n641_0[0]),.dinb(w_G3705_0[2]),.dout(n1065),.clk(gclk));
	jand g0751(.dina(n1065),.dinb(w_n354_0[1]),.dout(n1066),.clk(gclk));
	jor g0752(.dina(n1066),.dinb(w_dff_B_sYlCGmio9_1),.dout(n1067),.clk(gclk));
	jor g0753(.dina(w_n1067_0[2]),.dinb(w_dff_B_Dn49nIRW9_1),.dout(n1068),.clk(gclk));
	jand g0754(.dina(n1068),.dinb(w_dff_B_8ReLGgYj4_1),.dout(n1069),.clk(gclk));
	jand g0755(.dina(w_n1069_0[2]),.dinb(n1061),.dout(n1070),.clk(gclk));
	jnot g0756(.din(w_n1070_0[1]),.dout(n1071),.clk(gclk));
	jor g0757(.dina(w_n669_0[0]),.dinb(w_G4526_2[0]),.dout(n1072),.clk(gclk));
	jand g0758(.dina(w_dff_B_6U6LXPHR6_0),.dinb(n1071),.dout(n1073),.clk(gclk));
	jor g0759(.dina(w_n1073_0[1]),.dinb(w_n654_0[1]),.dout(n1074),.clk(gclk));
	jand g0760(.dina(n1074),.dinb(w_n653_0[0]),.dout(n1075),.clk(gclk));
	jxor g0761(.dina(n1075),.dinb(w_n626_1[0]),.dout(w_dff_A_x51Q2GgN5_2),.clk(gclk));
	jxor g0762(.dina(w_n1073_0[0]),.dinb(w_n631_0[1]),.dout(w_dff_A_tgXJYLwI4_2),.clk(gclk));
	jand g0763(.dina(w_n359_0[2]),.dinb(w_G4526_1[2]),.dout(n1078),.clk(gclk));
	jor g0764(.dina(w_n666_0[0]),.dinb(w_n1078_0[1]),.dout(n1079),.clk(gclk));
	jand g0765(.dina(n1079),.dinb(w_n661_0[1]),.dout(n1080),.clk(gclk));
	jxor g0766(.dina(n1080),.dinb(w_n636_0[1]),.dout(w_dff_A_hkO5sPZ89_2),.clk(gclk));
	jor g0767(.dina(w_n1078_0[0]),.dinb(w_n664_0[0]),.dout(n1082),.clk(gclk));
	jxor g0768(.dina(n1082),.dinb(w_n642_0[1]),.dout(w_dff_A_pvUyVpXg5_2),.clk(gclk));
	jxor g0769(.dina(w_n585_0[2]),.dinb(w_n582_0[0]),.dout(n1084),.clk(gclk));
	jor g0770(.dina(w_n1084_0[2]),.dinb(w_n678_0[0]),.dout(n1085),.clk(gclk));
	jnot g0771(.din(w_n646_0[0]),.dout(n1086),.clk(gclk));
	jnot g0772(.din(w_n647_0[0]),.dout(n1087),.clk(gclk));
	jnot g0773(.din(w_n654_0[0]),.dout(n1088),.clk(gclk));
	jand g0774(.dina(w_n1069_0[1]),.dinb(w_dff_B_C1fNn5vN1_1),.dout(n1089),.clk(gclk));
	jor g0775(.dina(n1089),.dinb(w_n652_0[0]),.dout(n1090),.clk(gclk));
	jor g0776(.dina(w_n1090_0[1]),.dinb(w_n649_0[0]),.dout(n1091),.clk(gclk));
	jand g0777(.dina(n1091),.dinb(w_dff_B_APXEe3xc8_1),.dout(n1092),.clk(gclk));
	jand g0778(.dina(w_n1092_0[2]),.dinb(w_n1086_0[1]),.dout(n1093),.clk(gclk));
	jnot g0779(.din(w_G4526_1[1]),.dout(n1094),.clk(gclk));
	jand g0780(.dina(w_n1092_0[1]),.dinb(w_n1094_0[2]),.dout(n1095),.clk(gclk));
	jor g0781(.dina(n1095),.dinb(n1093),.dout(n1096),.clk(gclk));
	jand g0782(.dina(w_n1096_0[1]),.dinb(w_n618_0[0]),.dout(n1097),.clk(gclk));
	jor g0783(.dina(n1097),.dinb(w_n619_0[1]),.dout(n1098),.clk(gclk));
	jor g0784(.dina(n1098),.dinb(w_n588_0[0]),.dout(n1099),.clk(gclk));
	jor g0785(.dina(w_n1099_0[1]),.dinb(w_n586_0[1]),.dout(n1100),.clk(gclk));
	jand g0786(.dina(n1100),.dinb(w_dff_B_TjLqO1u54_1),.dout(w_dff_A_GuechTS56_2),.clk(gclk));
	jand g0787(.dina(w_n676_0[1]),.dinb(w_n605_0[1]),.dout(n1102),.clk(gclk));
	jor g0788(.dina(n1102),.dinb(w_n615_0[1]),.dout(n1103),.clk(gclk));
	jxor g0789(.dina(n1103),.dinb(w_n594_0[1]),.dout(w_dff_A_ZvFxzFFl6_2),.clk(gclk));
	jnot g0790(.din(w_n599_0[0]),.dout(n1105),.clk(gclk));
	jnot g0791(.din(w_n613_0[1]),.dout(n1106),.clk(gclk));
	jnot g0792(.din(w_n603_0[2]),.dout(n1107),.clk(gclk));
	jand g0793(.dina(n1107),.dinb(w_G3729_0[2]),.dout(n1108),.clk(gclk));
	jor g0794(.dina(w_n1096_0[0]),.dinb(w_n1108_0[1]),.dout(n1109),.clk(gclk));
	jand g0795(.dina(n1109),.dinb(w_n1106_0[1]),.dout(n1110),.clk(gclk));
	jxor g0796(.dina(n1110),.dinb(w_n1105_0[1]),.dout(w_dff_A_5w4VshfQ8_2),.clk(gclk));
	jxor g0797(.dina(w_n676_0[0]),.dinb(w_n604_0[0]),.dout(w_dff_A_DUPrbXiE4_2),.clk(gclk));
	jnot g0798(.din(w_n436_0[0]),.dout(n1113),.clk(gclk));
	jor g0799(.dina(w_n1113_0[1]),.dinb(w_n431_0[0]),.dout(n1114),.clk(gclk));
	jnot g0800(.din(w_n432_0[0]),.dout(n1115),.clk(gclk));
	jor g0801(.dina(w_n435_0[0]),.dinb(n1115),.dout(n1116),.clk(gclk));
	jand g0802(.dina(n1116),.dinb(n1114),.dout(n1117),.clk(gclk));
	jnot g0803(.din(w_n459_0[0]),.dout(n1118),.clk(gclk));
	jxor g0804(.dina(w_n1118_0[1]),.dinb(w_n453_0[1]),.dout(n1119),.clk(gclk));
	jxor g0805(.dina(w_dff_B_LOeSXeM65_0),.dinb(n1117),.dout(n1120),.clk(gclk));
	jxor g0806(.dina(w_n485_0[0]),.dinb(w_n469_0[1]),.dout(n1121),.clk(gclk));
	jor g0807(.dina(w_n440_0[0]),.dinb(w_n422_0[0]),.dout(n1122),.clk(gclk));
	jnot g0808(.din(w_n423_0[0]),.dout(n1123),.clk(gclk));
	jor g0809(.dina(w_n427_0[0]),.dinb(n1123),.dout(n1124),.clk(gclk));
	jand g0810(.dina(n1124),.dinb(n1122),.dout(n1125),.clk(gclk));
	jnot g0811(.din(G141),.dout(n1126),.clk(gclk));
	jor g0812(.dina(n1126),.dinb(w_G18_20[0]),.dout(n1127),.clk(gclk));
	jnot g0813(.din(G161),.dout(n1128),.clk(gclk));
	jor g0814(.dina(n1128),.dinb(w_n355_15[0]),.dout(n1129),.clk(gclk));
	jand g0815(.dina(n1129),.dinb(w_n1127_0[1]),.dout(n1130),.clk(gclk));
	jxor g0816(.dina(n1130),.dinb(w_n479_0[2]),.dout(n1131),.clk(gclk));
	jxor g0817(.dina(w_dff_B_0aYxZ4TB8_0),.dinb(n1125),.dout(n1132),.clk(gclk));
	jxor g0818(.dina(n1132),.dinb(w_dff_B_GzZMZkHb1_1),.dout(n1133),.clk(gclk));
	jxor g0819(.dina(n1133),.dinb(w_dff_B_GoIcQ4gX1_1),.dout(n1134),.clk(gclk));
	jxor g0820(.dina(w_n603_0[1]),.dinb(w_n598_0[2]),.dout(n1135),.clk(gclk));
	jand g0821(.dina(G239),.dinb(w_G18_19[2]),.dout(n1136),.clk(gclk));
	jand g0822(.dina(w_dff_B_7T05TSdV1_0),.dinb(w_n355_14[2]),.dout(n1137),.clk(gclk));
	jor g0823(.dina(w_n1137_0[1]),.dinb(w_dff_B_d49urWCg8_1),.dout(n1138),.clk(gclk));
	jxor g0824(.dina(w_dff_B_B1RoABjt7_0),.dinb(w_n651_0[0]),.dout(n1139),.clk(gclk));
	jxor g0825(.dina(n1139),.dinb(w_dff_B_0tWcuBVx4_1),.dout(n1140),.clk(gclk));
	jand g0826(.dina(G229),.dinb(w_G18_19[1]),.dout(n1141),.clk(gclk));
	jor g0827(.dina(w_dff_B_WoLNCHGJ7_0),.dinb(w_n663_0[2]),.dout(n1142),.clk(gclk));
	jxor g0828(.dina(n1142),.dinb(w_n660_0[0]),.dout(n1143),.clk(gclk));
	jxor g0829(.dina(w_n635_0[1]),.dinb(w_n625_0[1]),.dout(n1144),.clk(gclk));
	jxor g0830(.dina(n1144),.dinb(n1143),.dout(n1145),.clk(gclk));
	jxor g0831(.dina(w_n593_0[1]),.dinb(w_n585_0[1]),.dout(n1146),.clk(gclk));
	jxor g0832(.dina(w_dff_B_hnkeOZ9E8_0),.dinb(n1145),.dout(n1147),.clk(gclk));
	jxor g0833(.dina(n1147),.dinb(n1140),.dout(n1148),.clk(gclk));
	jor g0834(.dina(w_dff_B_OBgwpE531_0),.dinb(n1134),.dout(n1149),.clk(gclk));
	jor g0835(.dina(w_n372_0[0]),.dinb(w_n355_14[1]),.dout(n1150),.clk(gclk));
	jxor g0836(.dina(G212),.dinb(G211),.dout(n1151),.clk(gclk));
	jxor g0837(.dina(n1151),.dinb(w_G209_0[0]),.dout(n1152),.clk(gclk));
	jor g0838(.dina(n1152),.dinb(w_n1150_0[1]),.dout(n1153),.clk(gclk));
	jnot g0839(.din(w_n386_0[0]),.dout(n1154),.clk(gclk));
	jand g0840(.dina(w_n395_0[2]),.dinb(n1154),.dout(n1155),.clk(gclk));
	jnot g0841(.din(w_n394_0[0]),.dout(n1156),.clk(gclk));
	jand g0842(.dina(n1156),.dinb(w_n387_0[1]),.dout(n1157),.clk(gclk));
	jor g0843(.dina(n1157),.dinb(n1155),.dout(n1158),.clk(gclk));
	jor g0844(.dina(w_n380_0[0]),.dinb(w_n374_0[0]),.dout(n1159),.clk(gclk));
	jnot g0845(.din(w_n375_0[0]),.dout(n1160),.clk(gclk));
	jor g0846(.dina(w_n378_0[0]),.dinb(n1160),.dout(n1161),.clk(gclk));
	jand g0847(.dina(n1161),.dinb(n1159),.dout(n1162),.clk(gclk));
	jxor g0848(.dina(n1162),.dinb(w_dff_B_FzkDygg79_1),.dout(n1163),.clk(gclk));
	jxor g0849(.dina(n1163),.dinb(w_dff_B_XmbktWK82_1),.dout(n1164),.clk(gclk));
	jxor g0850(.dina(w_n689_0[0]),.dinb(w_n504_0[2]),.dout(n1165),.clk(gclk));
	jxor g0851(.dina(w_n523_0[0]),.dinb(w_n517_0[2]),.dout(n1166),.clk(gclk));
	jxor g0852(.dina(w_dff_B_3qIHyXp94_0),.dinb(n1165),.dout(n1167),.clk(gclk));
	jxor g0853(.dina(w_n555_0[1]),.dinb(w_n539_0[1]),.dout(n1168),.clk(gclk));
	jxor g0854(.dina(w_n547_0[1]),.dinb(w_n531_0[1]),.dout(n1169),.clk(gclk));
	jxor g0855(.dina(n1169),.dinb(n1168),.dout(n1170),.clk(gclk));
	jand g0856(.dina(G227),.dinb(w_G18_19[0]),.dout(n1171),.clk(gclk));
	jand g0857(.dina(w_dff_B_NahVCNbJ8_0),.dinb(w_n355_14[0]),.dout(n1172),.clk(gclk));
	jor g0858(.dina(w_n1172_0[1]),.dinb(w_dff_B_OSNyLonq1_1),.dout(n1173),.clk(gclk));
	jxor g0859(.dina(n1173),.dinb(w_n563_0[2]),.dout(n1174),.clk(gclk));
	jxor g0860(.dina(w_dff_B_5zLcyl1i2_0),.dinb(n1170),.dout(n1175),.clk(gclk));
	jxor g0861(.dina(n1175),.dinb(n1167),.dout(n1176),.clk(gclk));
	jor g0862(.dina(w_dff_B_1RmXZwGf4_0),.dinb(n1164),.dout(n1177),.clk(gclk));
	jor g0863(.dina(w_dff_B_I71mcKFI5_0),.dinb(n1149),.dout(G412_fa_),.clk(gclk));
	jnot g0864(.din(w_n772_0[0]),.dout(n1179),.clk(gclk));
	jxor g0865(.dina(w_n780_0[0]),.dinb(n1179),.dout(n1180),.clk(gclk));
	jnot g0866(.din(w_G2208_0[1]),.dout(n1181),.clk(gclk));
	jor g0867(.dina(n1181),.dinb(w_n355_13[2]),.dout(n1182),.clk(gclk));
	jor g0868(.dina(G82),.dinb(w_G18_18[2]),.dout(n1183),.clk(gclk));
	jand g0869(.dina(w_dff_B_Ol64LYX28_0),.dinb(n1182),.dout(n1184),.clk(gclk));
	jxor g0870(.dina(n1184),.dinb(w_n827_0[0]),.dout(n1185),.clk(gclk));
	jxor g0871(.dina(w_dff_B_NiDkIno62_0),.dinb(n1180),.dout(n1186),.clk(gclk));
	jxor g0872(.dina(w_n806_0[0]),.dinb(w_n800_0[1]),.dout(n1187),.clk(gclk));
	jxor g0873(.dina(w_n820_0[0]),.dinb(w_n814_0[1]),.dout(n1188),.clk(gclk));
	jxor g0874(.dina(n1188),.dinb(n1187),.dout(n1189),.clk(gclk));
	jxor g0875(.dina(w_n764_0[0]),.dinb(w_n758_0[1]),.dout(n1190),.clk(gclk));
	jxor g0876(.dina(w_dff_B_xix0vYG33_0),.dinb(n1189),.dout(n1191),.clk(gclk));
	jxor g0877(.dina(n1191),.dinb(n1186),.dout(n1192),.clk(gclk));
	jxor g0878(.dina(w_n953_0[1]),.dinb(w_n947_0[0]),.dout(n1193),.clk(gclk));
	jxor g0879(.dina(w_n903_0[0]),.dinb(w_n894_0[0]),.dout(n1194),.clk(gclk));
	jxor g0880(.dina(n1194),.dinb(n1193),.dout(n1195),.clk(gclk));
	jnot g0881(.din(w_G3698_0[1]),.dout(n1196),.clk(gclk));
	jor g0882(.dina(n1196),.dinb(w_n355_13[1]),.dout(n1197),.clk(gclk));
	jor g0883(.dina(G69),.dinb(w_G18_18[1]),.dout(n1198),.clk(gclk));
	jand g0884(.dina(w_dff_B_KjMdpMqY3_0),.dinb(n1197),.dout(n1199),.clk(gclk));
	jxor g0885(.dina(n1199),.dinb(w_n888_0[0]),.dout(n1200),.clk(gclk));
	jor g0886(.dina(w_n662_0[0]),.dinb(w_n355_13[0]),.dout(n1201),.clk(gclk));
	jand g0887(.dina(n1201),.dinb(w_n905_0[0]),.dout(n1202),.clk(gclk));
	jxor g0888(.dina(n1202),.dinb(w_n919_0[0]),.dout(n1203),.clk(gclk));
	jxor g0889(.dina(n1203),.dinb(n1200),.dout(n1204),.clk(gclk));
	jnot g0890(.din(w_n930_0[0]),.dout(n1205),.clk(gclk));
	jxor g0891(.dina(w_n938_0[0]),.dinb(n1205),.dout(n1206),.clk(gclk));
	jxor g0892(.dina(n1206),.dinb(n1204),.dout(n1207),.clk(gclk));
	jxor g0893(.dina(n1207),.dinb(w_dff_B_LNa1SlTM1_1),.dout(n1208),.clk(gclk));
	jor g0894(.dina(n1208),.dinb(n1192),.dout(n1209),.clk(gclk));
	jxor g0895(.dina(w_n854_0[0]),.dinb(w_n848_0[1]),.dout(n1210),.clk(gclk));
	jxor g0896(.dina(w_n870_0[0]),.dinb(w_n862_0[0]),.dout(n1211),.clk(gclk));
	jxor g0897(.dina(n1211),.dinb(n1210),.dout(n1212),.clk(gclk));
	jxor g0898(.dina(w_n983_0[0]),.dinb(w_n977_0[1]),.dout(n1213),.clk(gclk));
	jand g0899(.dina(w_G4393_0[1]),.dinb(w_G18_18[0]),.dout(n1214),.clk(gclk));
	jnot g0900(.din(G58),.dout(n1215),.clk(gclk));
	jand g0901(.dina(n1215),.dinb(w_n355_12[2]),.dout(n1216),.clk(gclk));
	jor g0902(.dina(n1216),.dinb(w_dff_B_wC0aYQQN6_1),.dout(n1217),.clk(gclk));
	jxor g0903(.dina(n1217),.dinb(w_n970_0[0]),.dout(n1218),.clk(gclk));
	jxor g0904(.dina(w_n999_0[0]),.dinb(w_n991_0[0]),.dout(n1219),.clk(gclk));
	jxor g0905(.dina(n1219),.dinb(n1218),.dout(n1220),.clk(gclk));
	jxor g0906(.dina(n1220),.dinb(w_dff_B_1nQ57FpA3_1),.dout(n1221),.clk(gclk));
	jxor g0907(.dina(n1221),.dinb(w_dff_B_7CQ1qRfY7_1),.dout(n1222),.clk(gclk));
	jxor g0908(.dina(w_n366_0[0]),.dinb(w_G1492_1[0]),.dout(n1223),.clk(gclk));
	jor g0909(.dina(n1223),.dinb(w_n355_12[1]),.dout(n1224),.clk(gclk));
	jnot g0910(.din(w_G1455_0[0]),.dout(n1225),.clk(gclk));
	jxor g0911(.dina(w_G2204_0[0]),.dinb(n1225),.dout(n1226),.clk(gclk));
	jor g0912(.dina(n1226),.dinb(w_G18_17[2]),.dout(n1227),.clk(gclk));
	jand g0913(.dina(n1227),.dinb(n1224),.dout(n1228),.clk(gclk));
	jxor g0914(.dina(w_n729_0[1]),.dinb(w_n723_0[0]),.dout(n1229),.clk(gclk));
	jxor g0915(.dina(w_n747_0[0]),.dinb(w_n741_0[1]),.dout(n1230),.clk(gclk));
	jxor g0916(.dina(n1230),.dinb(n1229),.dout(n1231),.clk(gclk));
	jnot g0917(.din(w_G1459_0[1]),.dout(n1232),.clk(gclk));
	jor g0918(.dina(n1232),.dinb(w_n355_12[0]),.dout(n1233),.clk(gclk));
	jor g0919(.dina(G114),.dinb(w_G18_17[1]),.dout(n1234),.clk(gclk));
	jand g0920(.dina(w_dff_B_LRbrNLwJ6_0),.dinb(n1233),.dout(n1235),.clk(gclk));
	jxor g0921(.dina(n1235),.dinb(w_n734_0[0]),.dout(n1236),.clk(gclk));
	jxor g0922(.dina(w_dff_B_IVfu9r9O7_0),.dinb(n1231),.dout(n1237),.clk(gclk));
	jxor g0923(.dina(n1237),.dinb(w_dff_B_OCSbmqRp2_1),.dout(n1238),.clk(gclk));
	jor g0924(.dina(n1238),.dinb(n1222),.dout(n1239),.clk(gclk));
	jor g0925(.dina(n1239),.dinb(n1209),.dout(G414_fa_),.clk(gclk));
	jnot g0926(.din(w_n935_0[0]),.dout(n1241),.clk(gclk));
	jxor g0927(.dina(n1241),.dinb(w_n926_0[0]),.dout(n1242),.clk(gclk));
	jxor g0928(.dina(w_n950_0[1]),.dinb(w_n944_0[0]),.dout(n1243),.clk(gclk));
	jxor g0929(.dina(w_dff_B_aXUeyR8z8_0),.dinb(n1242),.dout(n1244),.clk(gclk));
	jand g0930(.dina(G208),.dinb(w_G18_17[0]),.dout(n1245),.clk(gclk));
	jor g0931(.dina(w_dff_B_7M8GAmf22_0),.dinb(w_n1137_0[0]),.dout(n1246),.clk(gclk));
	jand g0932(.dina(G198),.dinb(w_G18_16[2]),.dout(n1247),.clk(gclk));
	jor g0933(.dina(w_dff_B_y2n6IbNe1_0),.dinb(w_n663_0[1]),.dout(n1248),.clk(gclk));
	jxor g0934(.dina(n1248),.dinb(n1246),.dout(n1249),.clk(gclk));
	jxor g0935(.dina(w_n916_0[0]),.dinb(w_n885_0[0]),.dout(n1250),.clk(gclk));
	jxor g0936(.dina(n1250),.dinb(n1249),.dout(n1251),.clk(gclk));
	jxor g0937(.dina(w_n900_0[0]),.dinb(w_n891_0[0]),.dout(n1252),.clk(gclk));
	jxor g0938(.dina(w_dff_B_fgoR0sKj5_0),.dinb(n1251),.dout(n1253),.clk(gclk));
	jxor g0939(.dina(n1253),.dinb(n1244),.dout(n1254),.clk(gclk));
	jxor g0940(.dina(w_n866_0[0]),.dinb(w_n858_0[0]),.dout(n1255),.clk(gclk));
	jxor g0941(.dina(w_n995_0[0]),.dinb(w_n987_0[0]),.dout(n1256),.clk(gclk));
	jxor g0942(.dina(n1256),.dinb(n1255),.dout(n1257),.clk(gclk));
	jxor g0943(.dina(w_n980_0[0]),.dinb(w_n973_0[1]),.dout(n1258),.clk(gclk));
	jand g0944(.dina(G197),.dinb(w_G18_16[1]),.dout(n1259),.clk(gclk));
	jor g0945(.dina(w_dff_B_s4LIctIT6_0),.dinb(w_n1172_0[0]),.dout(n1260),.clk(gclk));
	jxor g0946(.dina(n1260),.dinb(w_n966_0[0]),.dout(n1261),.clk(gclk));
	jxor g0947(.dina(n1261),.dinb(n1258),.dout(n1262),.clk(gclk));
	jnot g0948(.din(w_n851_0[0]),.dout(n1263),.clk(gclk));
	jxor g0949(.dina(n1263),.dinb(w_n845_0[1]),.dout(n1264),.clk(gclk));
	jxor g0950(.dina(n1264),.dinb(n1262),.dout(n1265),.clk(gclk));
	jxor g0951(.dina(n1265),.dinb(w_dff_B_xjXDcDOB3_1),.dout(n1266),.clk(gclk));
	jor g0952(.dina(n1266),.dinb(n1254),.dout(n1267),.clk(gclk));
	jxor g0953(.dina(G165),.dinb(G164),.dout(n1268),.clk(gclk));
	jxor g0954(.dina(n1268),.dinb(w_dff_B_D0eYQcHv3_1),.dout(n1269),.clk(gclk));
	jor g0955(.dina(n1269),.dinb(w_n1150_0[0]),.dout(n1270),.clk(gclk));
	jnot g0956(.din(w_n736_0[0]),.dout(n1271),.clk(gclk));
	jand g0957(.dina(w_n744_0[0]),.dinb(n1271),.dout(n1272),.clk(gclk));
	jnot g0958(.din(w_n743_0[0]),.dout(n1273),.clk(gclk));
	jand g0959(.dina(n1273),.dinb(w_n737_0[1]),.dout(n1274),.clk(gclk));
	jor g0960(.dina(n1274),.dinb(n1272),.dout(n1275),.clk(gclk));
	jnot g0961(.din(w_n726_0[1]),.dout(n1276),.clk(gclk));
	jor g0962(.dina(n1276),.dinb(w_n719_0[0]),.dout(n1277),.clk(gclk));
	jnot g0963(.din(w_n720_0[0]),.dout(n1278),.clk(gclk));
	jor g0964(.dina(w_n725_0[0]),.dinb(n1278),.dout(n1279),.clk(gclk));
	jand g0965(.dina(n1279),.dinb(n1277),.dout(n1280),.clk(gclk));
	jxor g0966(.dina(n1280),.dinb(w_dff_B_Jjg7lsSH3_1),.dout(n1281),.clk(gclk));
	jxor g0967(.dina(n1281),.dinb(w_dff_B_t2sPzaDQ7_1),.dout(n1282),.clk(gclk));
	jor g0968(.dina(n1282),.dinb(n1267),.dout(n1283),.clk(gclk));
	jnot g0969(.din(G181),.dout(n1284),.clk(gclk));
	jor g0970(.dina(n1284),.dinb(w_n355_11[2]),.dout(n1285),.clk(gclk));
	jand g0971(.dina(n1285),.dinb(w_n1127_0[0]),.dout(n1286),.clk(gclk));
	jxor g0972(.dina(n1286),.dinb(w_n824_0[0]),.dout(n1287),.clk(gclk));
	jxor g0973(.dina(w_n803_0[0]),.dinb(w_n796_0[1]),.dout(n1288),.clk(gclk));
	jxor g0974(.dina(n1288),.dinb(n1287),.dout(n1289),.clk(gclk));
	jnot g0975(.din(w_n767_0[0]),.dout(n1290),.clk(gclk));
	jand g0976(.dina(w_n776_0[0]),.dinb(n1290),.dout(n1291),.clk(gclk));
	jnot g0977(.din(w_n775_0[0]),.dout(n1292),.clk(gclk));
	jand g0978(.dina(n1292),.dinb(w_n768_0[0]),.dout(n1293),.clk(gclk));
	jor g0979(.dina(n1293),.dinb(n1291),.dout(n1294),.clk(gclk));
	jnot g0980(.din(w_n754_0[0]),.dout(n1295),.clk(gclk));
	jand g0981(.dina(w_n761_0[0]),.dinb(n1295),.dout(n1296),.clk(gclk));
	jnot g0982(.din(w_n760_0[0]),.dout(n1297),.clk(gclk));
	jand g0983(.dina(n1297),.dinb(w_n755_0[1]),.dout(n1298),.clk(gclk));
	jor g0984(.dina(n1298),.dinb(n1296),.dout(n1299),.clk(gclk));
	jxor g0985(.dina(n1299),.dinb(n1294),.dout(n1300),.clk(gclk));
	jxor g0986(.dina(w_n817_0[0]),.dinb(w_n810_0[1]),.dout(n1301),.clk(gclk));
	jxor g0987(.dina(w_dff_B_rrXjb51L9_0),.dinb(n1300),.dout(n1302),.clk(gclk));
	jxor g0988(.dina(n1302),.dinb(w_dff_B_cfkoG1Vt8_1),.dout(n1303),.clk(gclk));
	jor g0989(.dina(w_dff_B_0hoj0HAF7_0),.dinb(n1283),.dout(G416_fa_),.clk(gclk));
	jnot g0990(.din(w_n480_1[0]),.dout(n1305),.clk(gclk));
	jnot g0991(.din(w_n505_0[0]),.dout(n1306),.clk(gclk));
	jnot g0992(.din(w_n513_1[0]),.dout(n1307),.clk(gclk));
	jnot g0993(.din(w_n524_1[0]),.dout(n1308),.clk(gclk));
	jnot g0994(.din(w_n572_1[0]),.dout(n1309),.clk(gclk));
	jnot g0995(.din(w_n581_0[1]),.dout(n1310),.clk(gclk));
	jnot g0996(.din(w_n586_0[0]),.dout(n1311),.clk(gclk));
	jand g0997(.dina(w_n1099_0[0]),.dinb(w_dff_B_nRC0Yr099_1),.dout(n1312),.clk(gclk));
	jor g0998(.dina(w_n1312_1[1]),.dinb(w_n1310_0[1]),.dout(n1313),.clk(gclk));
	jand g0999(.dina(n1313),.dinb(w_n1309_0[1]),.dout(n1314),.clk(gclk));
	jor g1000(.dina(n1314),.dinb(w_n526_0[1]),.dout(n1315),.clk(gclk));
	jor g1001(.dina(n1315),.dinb(w_n1308_0[1]),.dout(n1316),.clk(gclk));
	jor g1002(.dina(w_n1316_0[1]),.dinb(w_n518_1[0]),.dout(n1317),.clk(gclk));
	jor g1003(.dina(w_n1317_0[1]),.dinb(w_n1307_0[1]),.dout(n1318),.clk(gclk));
	jand g1004(.dina(w_n696_0[0]),.dinb(n1318),.dout(n1319),.clk(gclk));
	jor g1005(.dina(n1319),.dinb(w_n507_0[0]),.dout(n1320),.clk(gclk));
	jand g1006(.dina(n1320),.dinb(w_dff_B_uMs40pPp2_1),.dout(n1321),.clk(gclk));
	jxor g1007(.dina(w_n1321_1[1]),.dinb(w_dff_B_fnd0kqBg8_1),.dout(w_dff_A_3zfTOB0e0_2),.clk(gclk));
	jnot g1008(.din(w_n414_1[0]),.dout(n1323),.clk(gclk));
	jnot g1009(.din(w_n424_0[0]),.dout(n1324),.clk(gclk));
	jnot g1010(.din(w_n425_1[0]),.dout(n1325),.clk(gclk));
	jnot g1011(.din(w_n450_0[1]),.dout(n1326),.clk(gclk));
	jnot g1012(.din(w_n449_0[2]),.dout(n1327),.clk(gclk));
	jnot g1013(.din(w_n499_0[0]),.dout(n1328),.clk(gclk));
	jnot g1014(.din(w_n500_0[0]),.dout(n1329),.clk(gclk));
	jnot g1015(.din(w_n462_0[0]),.dout(n1330),.clk(gclk));
	jand g1016(.dina(w_n1321_1[0]),.dinb(w_dff_B_tHIbB0nD0_1),.dout(n1331),.clk(gclk));
	jand g1017(.dina(n1331),.dinb(w_dff_B_UXF6fFBc8_1),.dout(n1332),.clk(gclk));
	jor g1018(.dina(n1332),.dinb(w_dff_B_YiFqbGVX2_1),.dout(n1333),.clk(gclk));
	jand g1019(.dina(w_n1333_0[1]),.dinb(w_dff_B_QDCFzGIp4_1),.dout(n1334),.clk(gclk));
	jor g1020(.dina(n1334),.dinb(w_dff_B_qtVtrj7r8_1),.dout(n1335),.clk(gclk));
	jor g1021(.dina(n1335),.dinb(w_dff_B_6gFcWADp7_1),.dout(n1336),.clk(gclk));
	jand g1022(.dina(n1336),.dinb(w_dff_B_KmzGxk4w4_1),.dout(n1337),.clk(gclk));
	jxor g1023(.dina(w_n1337_1[1]),.dinb(w_n1323_0[1]),.dout(w_dff_A_fKN3Ov279_2),.clk(gclk));
	jand g1024(.dina(w_n1118_0[0]),.dinb(w_G2230_0[1]),.dout(n1339),.clk(gclk));
	jnot g1025(.din(n1339),.dout(n1340),.clk(gclk));
	jand g1026(.dina(w_n1321_0[2]),.dinb(w_n495_1[0]),.dout(n1341),.clk(gclk));
	jnot g1027(.din(n1341),.dout(n1342),.clk(gclk));
	jand g1028(.dina(n1342),.dinb(w_n497_1[0]),.dout(n1343),.clk(gclk));
	jand g1029(.dina(w_n1343_0[1]),.dinb(w_n1340_0[2]),.dout(n1344),.clk(gclk));
	jor g1030(.dina(w_n1344_0[1]),.dinb(w_n460_1[1]),.dout(n1345),.clk(gclk));
	jxor g1031(.dina(n1345),.dinb(w_n463_1[0]),.dout(w_dff_A_BYw8wZjg9_2),.clk(gclk));
	jor g1032(.dina(w_n1343_0[0]),.dinb(w_n464_0[1]),.dout(n1347),.clk(gclk));
	jnot g1033(.din(w_n1344_0[0]),.dout(n1348),.clk(gclk));
	jor g1034(.dina(n1348),.dinb(w_n460_1[0]),.dout(n1349),.clk(gclk));
	jand g1035(.dina(n1349),.dinb(w_dff_B_Q8Ztu0Pv0_1),.dout(w_dff_A_3tjmx9Te0_2),.clk(gclk));
	jnot g1036(.din(w_n489_0[1]),.dout(n1351),.clk(gclk));
	jor g1037(.dina(n1351),.dinb(w_n491_1[0]),.dout(n1352),.clk(gclk));
	jand g1038(.dina(w_n700_1[0]),.dinb(w_n481_0[0]),.dout(n1353),.clk(gclk));
	jor g1039(.dina(n1353),.dinb(w_dff_B_qcZSPAcg4_1),.dout(n1354),.clk(gclk));
	jxor g1040(.dina(n1354),.dinb(w_n470_0[1]),.dout(w_dff_A_gZ1v9epB1_2),.clk(gclk));
	jand g1041(.dina(w_n700_0[2]),.dinb(w_n480_0[2]),.dout(n1356),.clk(gclk));
	jor g1042(.dina(n1356),.dinb(w_n487_0[1]),.dout(n1357),.clk(gclk));
	jxor g1043(.dina(n1357),.dinb(w_n475_0[1]),.dout(w_dff_A_F2Gv4zZ05_2),.clk(gclk));
	jor g1044(.dina(w_n418_0[0]),.dinb(w_n411_1[0]),.dout(n1359),.clk(gclk));
	jor g1045(.dina(w_n707_1[1]),.dinb(w_n411_0[2]),.dout(n1360),.clk(gclk));
	jand g1046(.dina(n1360),.dinb(w_n1359_0[1]),.dout(n1361),.clk(gclk));
	jxor g1047(.dina(n1361),.dinb(w_n377_1[0]),.dout(w_dff_A_7obnZiGZ1_2),.clk(gclk));
	jand g1048(.dina(w_n415_0[0]),.dinb(w_n388_1[0]),.dout(n1363),.clk(gclk));
	jor g1049(.dina(w_dff_B_qzHqw6h73_0),.dinb(w_n409_1[0]),.dout(n1364),.clk(gclk));
	jor g1050(.dina(w_n707_1[0]),.dinb(w_n409_0[2]),.dout(n1365),.clk(gclk));
	jand g1051(.dina(n1365),.dinb(w_n1364_0[1]),.dout(n1366),.clk(gclk));
	jxor g1052(.dina(n1366),.dinb(w_n416_0[1]),.dout(w_dff_A_UdtblJ0F2_2),.clk(gclk));
	jnot g1053(.din(w_n388_0[2]),.dout(n1368),.clk(gclk));
	jnot g1054(.din(w_n396_1[0]),.dout(n1369),.clk(gclk));
	jnot g1055(.din(w_n392_0[1]),.dout(n1370),.clk(gclk));
	jor g1056(.dina(w_n1337_1[0]),.dinb(w_n1323_0[0]),.dout(n1371),.clk(gclk));
	jand g1057(.dina(n1371),.dinb(w_n1370_0[1]),.dout(n1372),.clk(gclk));
	jor g1058(.dina(w_n1372_0[1]),.dinb(w_n1369_0[1]),.dout(n1373),.clk(gclk));
	jand g1059(.dina(n1373),.dinb(w_n405_0[1]),.dout(n1374),.clk(gclk));
	jxor g1060(.dina(n1374),.dinb(w_dff_B_ThSv8kmx6_1),.dout(G333),.clk(gclk));
	jxor g1061(.dina(w_n1372_0[0]),.dinb(w_n1369_0[0]),.dout(w_dff_A_PsLnarY76_2),.clk(gclk));
	jor g1062(.dina(w_G416_0),.dinb(w_G414_0),.dout(n1377),.clk(gclk));
	jor g1063(.dina(w_G408_0),.dinb(w_G404_0),.dout(n1378),.clk(gclk));
	jor g1064(.dina(w_G410_0),.dinb(w_G406_0),.dout(n1379),.clk(gclk));
	jor g1065(.dina(w_dff_B_cmBMnGhB7_0),.dinb(w_G412_0),.dout(n1380),.clk(gclk));
	jor g1066(.dina(n1380),.dinb(w_dff_B_3IVVGFyI8_1),.dout(n1381),.clk(gclk));
	jor g1067(.dina(n1381),.dinb(w_dff_B_tS23SFrS2_1),.dout(w_dff_A_YlBNGGZi2_2),.clk(gclk));
	jxor g1068(.dina(w_n705_0[0]),.dinb(w_n425_0[2]),.dout(w_dff_A_PSGSlOxf2_2),.clk(gclk));
	jand g1069(.dina(w_n703_1[1]),.dinb(w_n438_0[0]),.dout(n1384),.clk(gclk));
	jor g1070(.dina(n1384),.dinb(w_n447_0[1]),.dout(n1385),.clk(gclk));
	jxor g1071(.dina(n1385),.dinb(w_n429_0[1]),.dout(w_dff_A_FicGj5tX6_2),.clk(gclk));
	jand g1072(.dina(w_n1113_0[0]),.dinb(w_G2239_0[2]),.dout(n1387),.clk(gclk));
	jnot g1073(.din(w_n1387_0[1]),.dout(n1388),.clk(gclk));
	jor g1074(.dina(w_n703_1[0]),.dinb(w_n445_0[1]),.dout(n1389),.clk(gclk));
	jand g1075(.dina(n1389),.dinb(w_n1388_0[1]),.dout(n1390),.clk(gclk));
	jxor g1076(.dina(n1390),.dinb(w_n433_1[0]),.dout(w_dff_A_IHdVYUXP2_2),.clk(gclk));
	jxor g1077(.dina(w_n703_0[2]),.dinb(w_n437_0[1]),.dout(w_dff_A_aKlzg0Oe8_2),.clk(gclk));
	jxor g1078(.dina(w_n680_2[1]),.dinb(w_n575_1[0]),.dout(w_dff_A_6BxXv4053_2),.clk(gclk));
	jor g1079(.dina(w_n712_0[1]),.dinb(w_G38_1[0]),.dout(n1394),.clk(gclk));
	jor g1080(.dina(w_n713_0[0]),.dinb(w_n709_1[0]),.dout(n1395),.clk(gclk));
	jand g1081(.dina(n1395),.dinb(w_dff_B_CBDC1UjX4_1),.dout(n1396),.clk(gclk));
	jxor g1082(.dina(w_n1396_0[1]),.dinb(w_n370_0[1]),.dout(G422),.clk(gclk));
	jxor g1083(.dina(w_n709_0[2]),.dinb(w_n363_0[1]),.dout(w_dff_A_3gY2Zx692_2),.clk(gclk));
	jand g1084(.dina(w_n680_2[0]),.dinb(w_n580_0[1]),.dout(n1399),.clk(gclk));
	jor g1085(.dina(n1399),.dinb(w_n570_1[1]),.dout(n1400),.clk(gclk));
	jxor g1086(.dina(n1400),.dinb(w_n573_1[0]),.dout(w_dff_A_pGz0TzDp7_2),.clk(gclk));
	jnot g1087(.din(w_n577_0[0]),.dout(n1402),.clk(gclk));
	jnot g1088(.din(w_n548_0[0]),.dout(n1403),.clk(gclk));
	jnot g1089(.din(w_n566_0[1]),.dout(n1404),.clk(gclk));
	jnot g1090(.din(w_n576_0[1]),.dout(n1405),.clk(gclk));
	jand g1091(.dina(w_dff_B_cX7DX5Th0_0),.dinb(n1404),.dout(n1406),.clk(gclk));
	jor g1092(.dina(n1406),.dinb(w_n550_0[0]),.dout(n1407),.clk(gclk));
	jand g1093(.dina(n1407),.dinb(w_dff_B_YuPztimZ1_1),.dout(n1408),.clk(gclk));
	jnot g1094(.din(w_n568_0[1]),.dout(n1409),.clk(gclk));
	jand g1095(.dina(w_n1312_1[0]),.dinb(w_dff_B_nY6fBif09_1),.dout(n1410),.clk(gclk));
	jor g1096(.dina(n1410),.dinb(w_n1408_0[1]),.dout(n1411),.clk(gclk));
	jxor g1097(.dina(n1411),.dinb(w_n1402_0[1]),.dout(w_dff_A_39LSarcR8_2),.clk(gclk));
	jand g1098(.dina(w_n680_1[2]),.dinb(w_n576_0[0]),.dout(n1413),.clk(gclk));
	jor g1099(.dina(n1413),.dinb(w_n566_0[0]),.dout(n1414),.clk(gclk));
	jxor g1100(.dina(n1414),.dinb(w_n578_0[1]),.dout(w_dff_A_Ok6uAbWN4_2),.clk(gclk));
	jand g1101(.dina(w_n680_1[1]),.dinb(w_n575_0[2]),.dout(n1416),.clk(gclk));
	jor g1102(.dina(n1416),.dinb(w_n564_0[1]),.dout(n1417),.clk(gclk));
	jxor g1103(.dina(n1417),.dinb(w_n574_0[1]),.dout(w_dff_A_N1mAsmmi2_2),.clk(gclk));
	jxor g1104(.dina(w_n504_0[1]),.dinb(w_n501_0[0]),.dout(n1419),.clk(gclk));
	jxor g1105(.dina(w_n1419_0[1]),.dinb(w_n698_0[0]),.dout(w_dff_A_HerJdIIO9_2),.clk(gclk));
	jand g1106(.dina(w_n694_0[0]),.dinb(w_n1317_0[0]),.dout(n1421),.clk(gclk));
	jxor g1107(.dina(n1421),.dinb(w_n1307_0[0]),.dout(w_dff_A_cmrFAdAy7_2),.clk(gclk));
	jxor g1108(.dina(w_n524_0[2]),.dinb(w_n518_0[2]),.dout(n1423),.clk(gclk));
	jor g1109(.dina(w_dff_B_njTeZRjP2_0),.dinb(w_n683_0[0]),.dout(n1424),.clk(gclk));
	jand g1110(.dina(n1424),.dinb(w_n1316_0[0]),.dout(w_dff_A_zYA4qFmc0_2),.clk(gclk));
	jxor g1111(.dina(w_n517_0[1]),.dinb(w_n514_0[0]),.dout(n1426),.clk(gclk));
	jxor g1112(.dina(w_n1426_0[1]),.dinb(w_n682_0[0]),.dout(w_dff_A_IpwnXTLg0_2),.clk(gclk));
	jxor g1113(.dina(w_n429_0[0]),.dinb(w_n425_0[1]),.dout(n1431),.clk(gclk));
	jor g1114(.dina(w_n1388_0[0]),.dinb(w_n444_0[1]),.dout(n1432),.clk(gclk));
	jnot g1115(.din(w_n447_0[0]),.dout(n1433),.clk(gclk));
	jor g1116(.dina(w_n1433_0[1]),.dinb(w_n1387_0[0]),.dout(n1434),.clk(gclk));
	jand g1117(.dina(n1434),.dinb(w_dff_B_OWbI6Hs37_1),.dout(n1435),.clk(gclk));
	jxor g1118(.dina(n1435),.dinb(w_n1431_0[1]),.dout(n1436),.clk(gclk));
	jxor g1119(.dina(w_n449_0[1]),.dinb(w_n433_0[2]),.dout(n1437),.clk(gclk));
	jxor g1120(.dina(w_dff_B_JOn9JoTf0_0),.dinb(n1436),.dout(n1438),.clk(gclk));
	jand g1121(.dina(w_dff_B_vnvmDqhx9_0),.dinb(w_n1333_0[0]),.dout(n1439),.clk(gclk));
	jxor g1122(.dina(w_n445_0[0]),.dinb(w_n433_0[1]),.dout(n1440),.clk(gclk));
	jnot g1123(.din(w_n1440_0[1]),.dout(n1441),.clk(gclk));
	jand g1124(.dina(w_dff_B_pA3M7hlw5_0),.dinb(w_n1433_0[0]),.dout(n1442),.clk(gclk));
	jor g1125(.dina(w_n437_0[0]),.dinb(w_n444_0[0]),.dout(n1443),.clk(gclk));
	jand g1126(.dina(n1443),.dinb(w_n1440_0[0]),.dout(n1444),.clk(gclk));
	jor g1127(.dina(w_dff_B_p3iDl0LL3_0),.dinb(n1442),.dout(n1445),.clk(gclk));
	jxor g1128(.dina(w_n1431_0[0]),.dinb(w_n450_0[0]),.dout(n1446),.clk(gclk));
	jxor g1129(.dina(n1446),.dinb(w_dff_B_19gLca623_1),.dout(n1447),.clk(gclk));
	jand g1130(.dina(w_dff_B_CYuVarN33_0),.dinb(w_n703_0[1]),.dout(n1448),.clk(gclk));
	jor g1131(.dina(n1448),.dinb(n1439),.dout(n1449),.clk(gclk));
	jand g1132(.dina(w_n497_0[2]),.dinb(w_n1340_0[1]),.dout(n1450),.clk(gclk));
	jor g1133(.dina(n1450),.dinb(w_n460_0[2]),.dout(n1451),.clk(gclk));
	jxor g1134(.dina(w_n480_0[1]),.dinb(w_n475_0[0]),.dout(n1452),.clk(gclk));
	jand g1135(.dina(w_n1452_0[2]),.dinb(w_n495_0[2]),.dout(n1453),.clk(gclk));
	jnot g1136(.din(w_n1452_0[1]),.dout(n1454),.clk(gclk));
	jand g1137(.dina(w_dff_B_ykHznQu92_0),.dinb(w_n497_0[1]),.dout(n1455),.clk(gclk));
	jor g1138(.dina(n1455),.dinb(w_dff_B_LIpDOmxh0_1),.dout(n1456),.clk(gclk));
	jnot g1139(.din(w_n479_0[1]),.dout(n1457),.clk(gclk));
	jand g1140(.dina(n1457),.dinb(w_G2211_0[1]),.dout(n1458),.clk(gclk));
	jnot g1141(.din(w_n1458_0[1]),.dout(n1459),.clk(gclk));
	jor g1142(.dina(n1459),.dinb(w_n491_0[2]),.dout(n1460),.clk(gclk));
	jor g1143(.dina(w_n1458_0[0]),.dinb(w_n486_0[0]),.dout(n1461),.clk(gclk));
	jand g1144(.dina(w_dff_B_wnS3s8PN9_0),.dinb(n1460),.dout(n1462),.clk(gclk));
	jxor g1145(.dina(n1462),.dinb(w_n463_0[2]),.dout(n1463),.clk(gclk));
	jxor g1146(.dina(w_dff_B_m0O3PEqb1_0),.dinb(n1456),.dout(n1464),.clk(gclk));
	jxor g1147(.dina(n1464),.dinb(w_dff_B_JQAzfofo1_1),.dout(n1465),.clk(gclk));
	jand g1148(.dina(w_dff_B_KBTEMHY11_0),.dinb(w_n700_0[1]),.dout(n1466),.clk(gclk));
	jand g1149(.dina(w_n496_0[0]),.dinb(w_n1340_0[0]),.dout(n1467),.clk(gclk));
	jor g1150(.dina(n1467),.dinb(w_n460_0[1]),.dout(n1468),.clk(gclk));
	jor g1151(.dina(w_n487_0[0]),.dinb(w_n491_0[1]),.dout(n1469),.clk(gclk));
	jand g1152(.dina(w_dff_B_eN8HR6yF0_0),.dinb(w_n489_0[0]),.dout(n1470),.clk(gclk));
	jxor g1153(.dina(n1470),.dinb(w_n463_0[1]),.dout(n1471),.clk(gclk));
	jxor g1154(.dina(n1471),.dinb(w_n495_0[1]),.dout(n1472),.clk(gclk));
	jxor g1155(.dina(n1472),.dinb(w_n1452_0[0]),.dout(n1473),.clk(gclk));
	jxor g1156(.dina(w_dff_B_BhWBXVsX9_0),.dinb(n1468),.dout(n1474),.clk(gclk));
	jand g1157(.dina(w_dff_B_9mp0lpax4_0),.dinb(w_n1321_0[1]),.dout(n1475),.clk(gclk));
	jor g1158(.dina(n1475),.dinb(n1466),.dout(n1476),.clk(gclk));
	jxor g1159(.dina(w_n470_0[0]),.dinb(w_n464_0[0]),.dout(n1477),.clk(gclk));
	jxor g1160(.dina(w_dff_B_4e0S8qxo6_0),.dinb(n1476),.dout(n1478),.clk(gclk));
	jxor g1161(.dina(w_dff_B_2uSCymEX3_0),.dinb(n1449),.dout(w_dff_A_DxbKqrBV1_2),.clk(gclk));
	jxor g1162(.dina(w_n416_0[0]),.dinb(w_n388_0[1]),.dout(n1480),.clk(gclk));
	jxor g1163(.dina(w_n411_0[1]),.dinb(w_n377_0[2]),.dout(n1481),.clk(gclk));
	jand g1164(.dina(w_n407_0[0]),.dinb(w_n1370_0[0]),.dout(n1482),.clk(gclk));
	jand g1165(.dina(w_n409_0[1]),.dinb(w_n392_0[0]),.dout(n1483),.clk(gclk));
	jor g1166(.dina(n1483),.dinb(w_dff_B_em3F549f2_1),.dout(n1484),.clk(gclk));
	jnot g1167(.din(w_n397_0[0]),.dout(n1485),.clk(gclk));
	jand g1168(.dina(n1485),.dinb(w_n405_0[0]),.dout(n1486),.clk(gclk));
	jxor g1169(.dina(w_n414_0[2]),.dinb(w_n396_0[2]),.dout(n1487),.clk(gclk));
	jxor g1170(.dina(w_dff_B_NbkvPVtR2_0),.dinb(w_n1486_0[1]),.dout(n1488),.clk(gclk));
	jxor g1171(.dina(w_dff_B_U9Uof8Zi7_0),.dinb(n1484),.dout(n1489),.clk(gclk));
	jxor g1172(.dina(n1489),.dinb(n1481),.dout(n1490),.clk(gclk));
	jor g1173(.dina(w_dff_B_icxVN9Xl1_0),.dinb(w_n707_0[2]),.dout(n1491),.clk(gclk));
	jor g1174(.dina(w_n391_0[0]),.dinb(w_n389_0[1]),.dout(n1492),.clk(gclk));
	jor g1175(.dina(w_n395_0[1]),.dinb(w_n393_0[1]),.dout(n1493),.clk(gclk));
	jand g1176(.dina(n1493),.dinb(w_n1492_0[1]),.dout(n1494),.clk(gclk));
	jnot g1177(.din(w_n1492_0[0]),.dout(n1495),.clk(gclk));
	jand g1178(.dina(w_n1486_0[0]),.dinb(w_dff_B_azEqYxyT5_1),.dout(n1496),.clk(gclk));
	jor g1179(.dina(n1496),.dinb(w_dff_B_y1FHGEko7_1),.dout(n1497),.clk(gclk));
	jxor g1180(.dina(w_n396_0[1]),.dinb(w_n377_0[1]),.dout(n1498),.clk(gclk));
	jxor g1181(.dina(w_dff_B_INzzAuzd4_0),.dinb(w_n1364_0[0]),.dout(n1499),.clk(gclk));
	jxor g1182(.dina(n1499),.dinb(w_dff_B_fY56sq2l1_1),.dout(n1500),.clk(gclk));
	jxor g1183(.dina(n1500),.dinb(w_n414_0[1]),.dout(n1501),.clk(gclk));
	jxor g1184(.dina(n1501),.dinb(w_n1359_0[0]),.dout(n1502),.clk(gclk));
	jor g1185(.dina(w_dff_B_kwGuXUXQ2_0),.dinb(w_n1337_0[2]),.dout(n1503),.clk(gclk));
	jand g1186(.dina(n1503),.dinb(n1491),.dout(n1504),.clk(gclk));
	jxor g1187(.dina(n1504),.dinb(w_dff_B_RQNtAc8l7_1),.dout(n1505),.clk(gclk));
	jand g1188(.dina(w_n362_0[0]),.dinb(w_G38_0[2]),.dout(n1506),.clk(gclk));
	jnot g1189(.din(w_n364_0[1]),.dout(n1507),.clk(gclk));
	jor g1190(.dina(n1507),.dinb(w_n1506_0[1]),.dout(n1508),.clk(gclk));
	jnot g1191(.din(w_n1506_0[0]),.dout(n1509),.clk(gclk));
	jor g1192(.dina(n1509),.dinb(w_G1496_0[2]),.dout(n1510),.clk(gclk));
	jand g1193(.dina(n1510),.dinb(w_dff_B_Eio5xOfu0_1),.dout(n1511),.clk(gclk));
	jand g1194(.dina(w_n1511_0[1]),.dinb(w_n413_0[2]),.dout(n1512),.clk(gclk));
	jnot g1195(.din(w_n413_0[1]),.dout(n1513),.clk(gclk));
	jand g1196(.dina(w_n712_0[0]),.dinb(w_n361_0[0]),.dout(n1514),.clk(gclk));
	jor g1197(.dina(w_n364_0[0]),.dinb(n1514),.dout(n1515),.clk(gclk));
	jor g1198(.dina(w_n369_0[0]),.dinb(w_G1492_0[2]),.dout(n1516),.clk(gclk));
	jand g1199(.dina(n1516),.dinb(n1515),.dout(n1517),.clk(gclk));
	jand g1200(.dina(w_dff_B_p90kH7vl4_0),.dinb(n1513),.dout(n1518),.clk(gclk));
	jor g1201(.dina(w_n1518_0[1]),.dinb(w_dff_B_IiTdSLe73_1),.dout(n1519),.clk(gclk));
	jor g1202(.dina(w_dff_B_To1HMDCp2_0),.dinb(w_n707_0[1]),.dout(n1520),.clk(gclk));
	jnot g1203(.din(w_n419_0[0]),.dout(n1521),.clk(gclk));
	jand g1204(.dina(w_n1518_0[0]),.dinb(w_dff_B_OTYgK7iz0_1),.dout(n1522),.clk(gclk));
	jand g1205(.dina(w_n1511_0[0]),.dinb(w_n420_0[0]),.dout(n1523),.clk(gclk));
	jor g1206(.dina(w_dff_B_uU2xQCE56_0),.dinb(n1522),.dout(n1524),.clk(gclk));
	jor g1207(.dina(w_dff_B_PBm2BaFD9_0),.dinb(w_n1337_0[1]),.dout(n1525),.clk(gclk));
	jand g1208(.dina(n1525),.dinb(n1520),.dout(n1526),.clk(gclk));
	jxor g1209(.dina(w_dff_B_M4dntbBX2_0),.dinb(n1505),.dout(w_dff_A_SofaJqix2_2),.clk(gclk));
	jor g1210(.dina(w_n693_0[0]),.dinb(w_n687_0[0]),.dout(n1528),.clk(gclk));
	jand g1211(.dina(w_dff_B_mkdFzHJL4_0),.dinb(w_n695_0[0]),.dout(n1529),.clk(gclk));
	jor g1212(.dina(w_n1529_0[1]),.dinb(w_n513_0[2]),.dout(n1530),.clk(gclk));
	jxor g1213(.dina(w_n1419_0[0]),.dinb(w_n1308_0[0]),.dout(n1531),.clk(gclk));
	jxor g1214(.dina(w_n1531_0[1]),.dinb(w_n526_0[0]),.dout(n1532),.clk(gclk));
	jxor g1215(.dina(w_dff_B_aaz4RO4F3_0),.dinb(n1530),.dout(n1533),.clk(gclk));
	jand g1216(.dina(w_dff_B_ryPHwt8F6_0),.dinb(w_n1309_0[0]),.dout(n1534),.clk(gclk));
	jand g1217(.dina(w_n1534_0[1]),.dinb(w_n1310_0[0]),.dout(n1535),.clk(gclk));
	jand g1218(.dina(w_n1426_0[0]),.dinb(w_n524_0[1]),.dout(n1536),.clk(gclk));
	jnot g1219(.din(w_n1536_0[1]),.dout(n1537),.clk(gclk));
	jor g1220(.dina(n1537),.dinb(w_n690_0[0]),.dout(n1538),.clk(gclk));
	jor g1221(.dina(w_n1536_0[0]),.dinb(w_n1529_0[0]),.dout(n1539),.clk(gclk));
	jand g1222(.dina(n1539),.dinb(w_dff_B_vpfiJFkd0_1),.dout(n1540),.clk(gclk));
	jxor g1223(.dina(w_n518_0[1]),.dinb(w_n513_0[1]),.dout(n1541),.clk(gclk));
	jxor g1224(.dina(w_dff_B_jn8IgKiS4_0),.dinb(w_n1531_0[0]),.dout(n1542),.clk(gclk));
	jxor g1225(.dina(w_dff_B_kAHKnmBg9_0),.dinb(n1540),.dout(n1543),.clk(gclk));
	jor g1226(.dina(w_n581_0[0]),.dinb(w_n572_0[2]),.dout(n1544),.clk(gclk));
	jand g1227(.dina(n1544),.dinb(w_n1543_0[1]),.dout(n1545),.clk(gclk));
	jor g1228(.dina(w_dff_B_TmRP1p7q3_0),.dinb(n1535),.dout(n1546),.clk(gclk));
	jand g1229(.dina(n1546),.dinb(w_n680_1[0]),.dout(n1547),.clk(gclk));
	jand g1230(.dina(w_n1543_0[0]),.dinb(w_n572_0[1]),.dout(n1548),.clk(gclk));
	jor g1231(.dina(w_dff_B_JwPkVB3w4_0),.dinb(w_n1534_0[0]),.dout(n1549),.clk(gclk));
	jand g1232(.dina(w_dff_B_pTgNxzNA1_0),.dinb(w_n1312_0[2]),.dout(n1550),.clk(gclk));
	jor g1233(.dina(n1550),.dinb(n1547),.dout(n1551),.clk(gclk));
	jxor g1234(.dina(w_n578_0[0]),.dinb(w_n1402_0[0]),.dout(n1552),.clk(gclk));
	jnot g1235(.din(w_n563_0[1]),.dout(n1553),.clk(gclk));
	jand g1236(.dina(n1553),.dinb(w_G4394_0[2]),.dout(n1554),.clk(gclk));
	jnot g1237(.din(w_n1554_0[1]),.dout(n1555),.clk(gclk));
	jand g1238(.dina(n1555),.dinb(w_n558_0[0]),.dout(n1556),.clk(gclk));
	jand g1239(.dina(w_n1554_0[0]),.dinb(w_n556_0[1]),.dout(n1557),.clk(gclk));
	jor g1240(.dina(w_dff_B_uz5JdEPA2_0),.dinb(n1556),.dout(n1558),.clk(gclk));
	jxor g1241(.dina(n1558),.dinb(w_n573_0[2]),.dout(n1559),.clk(gclk));
	jxor g1242(.dina(w_dff_B_anNSMSO76_0),.dinb(w_n1408_0[0]),.dout(n1560),.clk(gclk));
	jnot g1243(.din(w_n570_1[0]),.dout(n1561),.clk(gclk));
	jxor g1244(.dina(w_n575_0[1]),.dinb(w_n574_0[0]),.dout(n1562),.clk(gclk));
	jnot g1245(.din(w_n1562_0[2]),.dout(n1563),.clk(gclk));
	jor g1246(.dina(w_dff_B_fc44wMvx8_0),.dinb(n1561),.dout(n1564),.clk(gclk));
	jor g1247(.dina(w_n1562_0[1]),.dinb(w_n570_0[2]),.dout(n1565),.clk(gclk));
	jor g1248(.dina(n1565),.dinb(w_n580_0[0]),.dout(n1566),.clk(gclk));
	jand g1249(.dina(n1566),.dinb(n1564),.dout(n1567),.clk(gclk));
	jxor g1250(.dina(n1567),.dinb(w_dff_B_tHfsW3vq4_1),.dout(n1568),.clk(gclk));
	jor g1251(.dina(w_dff_B_CCxRpgky9_0),.dinb(w_n1312_0[1]),.dout(n1569),.clk(gclk));
	jxor g1252(.dina(w_n1562_0[0]),.dinb(w_n570_0[1]),.dout(n1570),.clk(gclk));
	jnot g1253(.din(w_n565_0[0]),.dout(n1571),.clk(gclk));
	jor g1254(.dina(w_n564_0[0]),.dinb(w_n556_0[0]),.dout(n1572),.clk(gclk));
	jand g1255(.dina(w_dff_B_fXaCUOCl5_0),.dinb(n1571),.dout(n1573),.clk(gclk));
	jxor g1256(.dina(n1573),.dinb(w_n573_0[1]),.dout(n1574),.clk(gclk));
	jxor g1257(.dina(n1574),.dinb(w_n568_0[0]),.dout(n1575),.clk(gclk));
	jxor g1258(.dina(w_dff_B_C8X1P6Dm0_0),.dinb(n1570),.dout(n1576),.clk(gclk));
	jor g1259(.dina(w_dff_B_uPo0wcI66_0),.dinb(w_n680_0[2]),.dout(n1577),.clk(gclk));
	jand g1260(.dina(n1577),.dinb(n1569),.dout(n1578),.clk(gclk));
	jxor g1261(.dina(n1578),.dinb(w_dff_B_UjeyhpaG1_1),.dout(n1579),.clk(gclk));
	jxor g1262(.dina(n1579),.dinb(w_dff_B_103VmZWn5_1),.dout(w_dff_A_jT5X6nYq2_2),.clk(gclk));
	jxor g1263(.dina(w_n1084_0[1]),.dinb(w_n1108_0[0]),.dout(n1581),.clk(gclk));
	jxor g1264(.dina(n1581),.dinb(w_n1105_0[0]),.dout(n1582),.clk(gclk));
	jand g1265(.dina(w_n616_0[0]),.dinb(w_n609_0[0]),.dout(n1583),.clk(gclk));
	jand g1266(.dina(w_n615_0[0]),.dinb(w_n610_0[0]),.dout(n1584),.clk(gclk));
	jor g1267(.dina(w_dff_B_FekjwbPH0_0),.dinb(n1583),.dout(n1585),.clk(gclk));
	jxor g1268(.dina(n1585),.dinb(w_dff_B_GtBINyod8_1),.dout(n1586),.clk(gclk));
	jand g1269(.dina(w_dff_B_L2qPwmGX6_0),.dinb(w_n1092_0[0]),.dout(n1587),.clk(gclk));
	jand g1270(.dina(w_n1587_0[1]),.dinb(w_n1086_0[0]),.dout(n1588),.clk(gclk));
	jnot g1271(.din(w_n598_0[1]),.dout(n1589),.clk(gclk));
	jand g1272(.dina(n1589),.dinb(w_G3737_0[1]),.dout(n1590),.clk(gclk));
	jand g1273(.dina(w_n1106_0[0]),.dinb(n1590),.dout(n1591),.clk(gclk));
	jand g1274(.dina(w_n613_0[0]),.dinb(w_n612_0[0]),.dout(n1592),.clk(gclk));
	jor g1275(.dina(w_dff_B_veFixvxm7_0),.dinb(n1591),.dout(n1593),.clk(gclk));
	jor g1276(.dina(n1593),.dinb(w_n605_0[0]),.dout(n1594),.clk(gclk));
	jxor g1277(.dina(w_n1084_0[0]),.dinb(w_n594_0[0]),.dout(n1595),.clk(gclk));
	jxor g1278(.dina(w_dff_B_kzPwRbqB8_0),.dinb(n1594),.dout(n1596),.clk(gclk));
	jxor g1279(.dina(w_dff_B_wFidWInp6_0),.dinb(w_n619_0[0]),.dout(n1597),.clk(gclk));
	jand g1280(.dina(w_n1597_0[1]),.dinb(w_n674_0[0]),.dout(n1598),.clk(gclk));
	jor g1281(.dina(n1598),.dinb(w_n1094_0[1]),.dout(n1599),.clk(gclk));
	jor g1282(.dina(n1599),.dinb(w_dff_B_AkmfGLxS3_1),.dout(n1600),.clk(gclk));
	jand g1283(.dina(w_n1597_0[0]),.dinb(w_n673_0[0]),.dout(n1601),.clk(gclk));
	jor g1284(.dina(n1601),.dinb(w_n1587_0[0]),.dout(n1602),.clk(gclk));
	jor g1285(.dina(n1602),.dinb(w_G4526_1[0]),.dout(n1603),.clk(gclk));
	jand g1286(.dina(w_dff_B_oHa9ooEO4_0),.dinb(n1600),.dout(n1604),.clk(gclk));
	jxor g1287(.dina(w_n642_0[0]),.dinb(w_n359_0[1]),.dout(n1605),.clk(gclk));
	jxor g1288(.dina(w_n1605_0[1]),.dinb(w_n1067_0[1]),.dout(n1606),.clk(gclk));
	jxor g1289(.dina(w_dff_B_2Jgxhcxe8_0),.dinb(w_n1069_0[0]),.dout(n1607),.clk(gclk));
	jnot g1290(.din(w_n1607_0[1]),.dout(n1608),.clk(gclk));
	jxor g1291(.dina(w_n626_0[2]),.dinb(w_n354_0[0]),.dout(n1609),.clk(gclk));
	jxor g1292(.dina(w_dff_B_YhKwkhYb7_0),.dinb(w_n671_0[0]),.dout(n1610),.clk(gclk));
	jor g1293(.dina(w_n1610_0[1]),.dinb(w_dff_B_Ak1eFJ806_1),.dout(n1611),.clk(gclk));
	jnot g1294(.din(w_n1610_0[0]),.dout(n1612),.clk(gclk));
	jor g1295(.dina(n1612),.dinb(w_n1607_0[0]),.dout(n1613),.clk(gclk));
	jand g1296(.dina(n1613),.dinb(w_n1094_0[0]),.dout(n1614),.clk(gclk));
	jand g1297(.dina(n1614),.dinb(w_dff_B_R2AitHJL1_1),.dout(n1615),.clk(gclk));
	jand g1298(.dina(w_n1067_0[0]),.dinb(w_n357_0[0]),.dout(n1616),.clk(gclk));
	jand g1299(.dina(w_n661_0[0]),.dinb(w_n358_0[0]),.dout(n1617),.clk(gclk));
	jor g1300(.dina(w_dff_B_0ZuZZlVW5_0),.dinb(n1616),.dout(n1618),.clk(gclk));
	jxor g1301(.dina(n1618),.dinb(w_n626_0[1]),.dout(n1619),.clk(gclk));
	jxor g1302(.dina(n1619),.dinb(w_n1070_0[0]),.dout(n1620),.clk(gclk));
	jnot g1303(.din(w_n1620_0[1]),.dout(n1621),.clk(gclk));
	jnot g1304(.din(w_n645_0[0]),.dout(n1622),.clk(gclk));
	jand g1305(.dina(w_n1090_0[0]),.dinb(w_dff_B_rJyFWDR91_1),.dout(n1623),.clk(gclk));
	jxor g1306(.dina(n1623),.dinb(w_n1605_0[0]),.dout(n1624),.clk(gclk));
	jnot g1307(.din(w_n1624_0[1]),.dout(n1625),.clk(gclk));
	jor g1308(.dina(n1625),.dinb(w_dff_B_ngg18DwO4_1),.dout(n1626),.clk(gclk));
	jor g1309(.dina(w_n1624_0[0]),.dinb(w_n1620_0[0]),.dout(n1627),.clk(gclk));
	jand g1310(.dina(n1627),.dinb(w_G4526_0[2]),.dout(n1628),.clk(gclk));
	jand g1311(.dina(n1628),.dinb(n1626),.dout(n1629),.clk(gclk));
	jor g1312(.dina(n1629),.dinb(n1615),.dout(n1630),.clk(gclk));
	jxor g1313(.dina(w_n636_0[0]),.dinb(w_n631_0[0]),.dout(n1631),.clk(gclk));
	jxor g1314(.dina(w_dff_B_3p4fg0Jy6_0),.dinb(n1630),.dout(n1632),.clk(gclk));
	jxor g1315(.dina(n1632),.dinb(n1604),.dout(w_dff_A_3UnuSp1X4_2),.clk(gclk));
	buf g1316(.din(w_G1_1[1]),.dout(w_dff_A_22M6stkl3_1));
	buf g1317(.din(w_G1_1[0]),.dout(w_dff_A_FXX2zFPh3_1));
	buf g1318(.din(w_G1459_0[0]),.dout(w_dff_A_APRPgR7j9_1));
	buf g1319(.din(w_G1469_0[0]),.dout(w_dff_A_NJEEXzqd5_1));
	buf g1320(.din(w_G1480_0[0]),.dout(w_dff_A_pjeMTmIZ9_1));
	buf g1321(.din(w_G1486_0[0]),.dout(w_dff_A_wpKXgQFK7_1));
	buf g1322(.din(w_G1492_0[1]),.dout(w_dff_A_anzn7UR03_1));
	buf g1323(.din(w_G1496_0[1]),.dout(w_dff_A_SmHHSwBU9_1));
	buf g1324(.din(w_G2208_0[0]),.dout(w_dff_A_80xgeO6u2_1));
	buf g1325(.din(w_G2218_0[0]),.dout(w_dff_A_YVg7X2Az1_1));
	buf g1326(.din(w_G2224_0[1]),.dout(w_dff_A_mpaoxbKU2_1));
	buf g1327(.din(w_G2230_0[0]),.dout(w_dff_A_gICE3Ix18_1));
	buf g1328(.din(w_G2236_0[0]),.dout(w_dff_A_m3c6GcYD1_1));
	buf g1329(.din(w_G2239_0[1]),.dout(w_dff_A_DbjIJw5y8_1));
	buf g1330(.din(w_G2247_0[0]),.dout(w_dff_A_b76irSqt9_1));
	buf g1331(.din(w_G2253_0[0]),.dout(w_dff_A_TsLfMgku7_1));
	buf g1332(.din(w_G2256_0[0]),.dout(w_dff_A_2530MqCy4_1));
	buf g1333(.din(w_G3698_0[0]),.dout(w_dff_A_LItvViFw0_1));
	buf g1334(.din(w_G3701_0[1]),.dout(w_dff_A_vnhaT5SN9_1));
	buf g1335(.din(w_G3705_0[1]),.dout(w_dff_A_LUDcVW948_1));
	buf g1336(.din(w_G3711_0[0]),.dout(w_dff_A_YgGp9OAD8_1));
	buf g1337(.din(w_G3717_0[0]),.dout(w_dff_A_0NogE0yY4_1));
	buf g1338(.din(w_G3723_0[0]),.dout(w_dff_A_B1CtAN1E0_1));
	buf g1339(.din(w_G3729_0[1]),.dout(w_dff_A_OfvxdAZI9_1));
	buf g1340(.din(w_G3737_0[0]),.dout(w_dff_A_raA4ZSOf6_1));
	buf g1341(.din(w_G3743_0[0]),.dout(w_dff_A_cdzx6Owo0_1));
	buf g1342(.din(w_G3749_0[0]),.dout(w_dff_A_34A5K7yA7_1));
	buf g1343(.din(w_G4393_0[0]),.dout(w_dff_A_kb3quiGP8_1));
	buf g1344(.din(w_G4400_0[1]),.dout(w_dff_A_5GiWzOQF0_1));
	buf g1345(.din(w_G4405_0[1]),.dout(w_dff_A_vkEKZ9tY8_1));
	buf g1346(.din(w_G4410_0[0]),.dout(w_dff_A_Y0XsnTNc9_1));
	buf g1347(.din(w_G4415_0[1]),.dout(w_dff_A_o22oslEs2_1));
	buf g1348(.din(w_G4420_0[1]),.dout(w_dff_A_HR72Rhmh8_1));
	buf g1349(.din(w_G4427_0[0]),.dout(w_dff_A_p7sM1NwD4_1));
	buf g1350(.din(w_G4432_0[0]),.dout(w_dff_A_vAZbA4Z74_1));
	buf g1351(.din(w_G4437_0[0]),.dout(w_dff_A_mt2rqSeK3_1));
	buf g1352(.din(w_G1462_0[0]),.dout(w_dff_A_l1LtiW1L5_1));
	buf g1353(.din(w_G2211_0[0]),.dout(w_dff_A_gDU3XBye5_1));
	buf g1354(.din(w_G4394_0[1]),.dout(w_dff_A_A1UvnyQh2_1));
	buf g1355(.din(w_G1_0[2]),.dout(w_dff_A_Vu8cR4Jp7_1));
	buf g1356(.din(w_G106_0[1]),.dout(w_dff_A_5vq1NzK46_1));
	jnot g1357(.din(w_G15_0[1]),.dout(w_dff_A_LK3Lj7IW8_1),.clk(gclk));
	jor g1358(.dina(w_n345_0[0]),.dinb(w_G5_0[1]),.dout(w_dff_A_Zda8mllT3_2),.clk(gclk));
	jnot g1359(.din(w_G15_0[0]),.dout(w_dff_A_GbPQfCGT0_1),.clk(gclk));
	jor g1360(.dina(w_n349_0[0]),.dinb(w_n347_0[0]),.dout(w_dff_A_9eF0pr3b7_2),.clk(gclk));
	buf g1361(.din(w_G1_0[1]),.dout(w_dff_A_VajKcQKi2_1));
	jand g1362(.dina(w_n1059_0[1]),.dinb(w_n718_0[1]),.dout(w_dff_A_Q0KcgJhF3_2),.clk(gclk));
	jor g1363(.dina(w_n715_1[0]),.dinb(w_n711_1[0]),.dout(G270),.clk(gclk));
	jand g1364(.dina(w_n1059_0[0]),.dinb(w_n718_0[0]),.dout(w_dff_A_5fdEYc6z9_2),.clk(gclk));
	jor g1365(.dina(w_n715_0[2]),.dinb(w_n711_0[2]),.dout(G276),.clk(gclk));
	jor g1366(.dina(w_n715_0[1]),.dinb(w_n711_0[1]),.dout(G273),.clk(gclk));
	jxor g1367(.dina(w_n1396_0[0]),.dinb(w_n370_0[0]),.dout(G469),.clk(gclk));
	jxor g1368(.dina(w_n709_0[1]),.dinb(w_n363_0[0]),.dout(w_dff_A_aRxRy8Qx1_2),.clk(gclk));
	jspl3 jspl3_w_G1_0(.douta(w_G1_0[0]),.doutb(w_G1_0[1]),.doutc(w_G1_0[2]),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_G1_1[0]),.doutb(w_G1_1[1]),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl3 jspl3_w_G5_0(.douta(w_G5_0[0]),.doutb(w_dff_A_oNTQhwtA1_1),.doutc(w_dff_A_1a3BOk4N7_2),.din(G5));
	jspl jspl_w_G5_1(.douta(w_dff_A_T5tMKu6E2_0),.doutb(w_G5_1[1]),.din(w_G5_0[0]));
	jspl3 jspl3_w_G15_0(.douta(w_G15_0[0]),.doutb(w_G15_0[1]),.doutc(w_G15_0[2]),.din(G15));
	jspl3 jspl3_w_G18_0(.douta(w_G18_0[0]),.doutb(w_G18_0[1]),.doutc(w_G18_0[2]),.din(G18));
	jspl3 jspl3_w_G18_1(.douta(w_G18_1[0]),.doutb(w_G18_1[1]),.doutc(w_G18_1[2]),.din(w_G18_0[0]));
	jspl3 jspl3_w_G18_2(.douta(w_G18_2[0]),.doutb(w_G18_2[1]),.doutc(w_G18_2[2]),.din(w_G18_0[1]));
	jspl3 jspl3_w_G18_3(.douta(w_G18_3[0]),.doutb(w_G18_3[1]),.doutc(w_G18_3[2]),.din(w_G18_0[2]));
	jspl3 jspl3_w_G18_4(.douta(w_G18_4[0]),.doutb(w_G18_4[1]),.doutc(w_G18_4[2]),.din(w_G18_1[0]));
	jspl3 jspl3_w_G18_5(.douta(w_G18_5[0]),.doutb(w_G18_5[1]),.doutc(w_G18_5[2]),.din(w_G18_1[1]));
	jspl3 jspl3_w_G18_6(.douta(w_G18_6[0]),.doutb(w_G18_6[1]),.doutc(w_G18_6[2]),.din(w_G18_1[2]));
	jspl3 jspl3_w_G18_7(.douta(w_G18_7[0]),.doutb(w_G18_7[1]),.doutc(w_G18_7[2]),.din(w_G18_2[0]));
	jspl3 jspl3_w_G18_8(.douta(w_G18_8[0]),.doutb(w_G18_8[1]),.doutc(w_G18_8[2]),.din(w_G18_2[1]));
	jspl3 jspl3_w_G18_9(.douta(w_G18_9[0]),.doutb(w_G18_9[1]),.doutc(w_G18_9[2]),.din(w_G18_2[2]));
	jspl3 jspl3_w_G18_10(.douta(w_G18_10[0]),.doutb(w_G18_10[1]),.doutc(w_G18_10[2]),.din(w_G18_3[0]));
	jspl3 jspl3_w_G18_11(.douta(w_G18_11[0]),.doutb(w_G18_11[1]),.doutc(w_G18_11[2]),.din(w_G18_3[1]));
	jspl3 jspl3_w_G18_12(.douta(w_G18_12[0]),.doutb(w_G18_12[1]),.doutc(w_G18_12[2]),.din(w_G18_3[2]));
	jspl3 jspl3_w_G18_13(.douta(w_G18_13[0]),.doutb(w_G18_13[1]),.doutc(w_G18_13[2]),.din(w_G18_4[0]));
	jspl3 jspl3_w_G18_14(.douta(w_G18_14[0]),.doutb(w_G18_14[1]),.doutc(w_G18_14[2]),.din(w_G18_4[1]));
	jspl3 jspl3_w_G18_15(.douta(w_G18_15[0]),.doutb(w_G18_15[1]),.doutc(w_G18_15[2]),.din(w_G18_4[2]));
	jspl3 jspl3_w_G18_16(.douta(w_G18_16[0]),.doutb(w_G18_16[1]),.doutc(w_G18_16[2]),.din(w_G18_5[0]));
	jspl3 jspl3_w_G18_17(.douta(w_G18_17[0]),.doutb(w_G18_17[1]),.doutc(w_dff_A_frr3oQK92_2),.din(w_G18_5[1]));
	jspl3 jspl3_w_G18_18(.douta(w_G18_18[0]),.doutb(w_G18_18[1]),.doutc(w_G18_18[2]),.din(w_G18_5[2]));
	jspl3 jspl3_w_G18_19(.douta(w_G18_19[0]),.doutb(w_G18_19[1]),.doutc(w_G18_19[2]),.din(w_G18_6[0]));
	jspl3 jspl3_w_G18_20(.douta(w_dff_A_UYOAdUYd4_0),.doutb(w_G18_20[1]),.doutc(w_G18_20[2]),.din(w_G18_6[1]));
	jspl3 jspl3_w_G18_21(.douta(w_G18_21[0]),.doutb(w_G18_21[1]),.doutc(w_G18_21[2]),.din(w_G18_6[2]));
	jspl3 jspl3_w_G18_22(.douta(w_G18_22[0]),.doutb(w_G18_22[1]),.doutc(w_G18_22[2]),.din(w_G18_7[0]));
	jspl3 jspl3_w_G18_23(.douta(w_G18_23[0]),.doutb(w_G18_23[1]),.doutc(w_G18_23[2]),.din(w_G18_7[1]));
	jspl3 jspl3_w_G18_24(.douta(w_G18_24[0]),.doutb(w_G18_24[1]),.doutc(w_G18_24[2]),.din(w_G18_7[2]));
	jspl3 jspl3_w_G18_25(.douta(w_G18_25[0]),.doutb(w_G18_25[1]),.doutc(w_G18_25[2]),.din(w_G18_8[0]));
	jspl3 jspl3_w_G18_26(.douta(w_G18_26[0]),.doutb(w_G18_26[1]),.doutc(w_G18_26[2]),.din(w_G18_8[1]));
	jspl3 jspl3_w_G18_27(.douta(w_G18_27[0]),.doutb(w_G18_27[1]),.doutc(w_G18_27[2]),.din(w_G18_8[2]));
	jspl3 jspl3_w_G18_28(.douta(w_G18_28[0]),.doutb(w_G18_28[1]),.doutc(w_G18_28[2]),.din(w_G18_9[0]));
	jspl3 jspl3_w_G18_29(.douta(w_G18_29[0]),.doutb(w_G18_29[1]),.doutc(w_G18_29[2]),.din(w_G18_9[1]));
	jspl3 jspl3_w_G18_30(.douta(w_G18_30[0]),.doutb(w_G18_30[1]),.doutc(w_G18_30[2]),.din(w_G18_9[2]));
	jspl3 jspl3_w_G18_31(.douta(w_G18_31[0]),.doutb(w_G18_31[1]),.doutc(w_G18_31[2]),.din(w_G18_10[0]));
	jspl3 jspl3_w_G18_32(.douta(w_G18_32[0]),.doutb(w_G18_32[1]),.doutc(w_G18_32[2]),.din(w_G18_10[1]));
	jspl3 jspl3_w_G18_33(.douta(w_G18_33[0]),.doutb(w_G18_33[1]),.doutc(w_G18_33[2]),.din(w_G18_10[2]));
	jspl3 jspl3_w_G18_34(.douta(w_G18_34[0]),.doutb(w_G18_34[1]),.doutc(w_G18_34[2]),.din(w_G18_11[0]));
	jspl3 jspl3_w_G18_35(.douta(w_G18_35[0]),.doutb(w_G18_35[1]),.doutc(w_G18_35[2]),.din(w_G18_11[1]));
	jspl3 jspl3_w_G18_36(.douta(w_G18_36[0]),.doutb(w_G18_36[1]),.doutc(w_G18_36[2]),.din(w_G18_11[2]));
	jspl3 jspl3_w_G18_37(.douta(w_G18_37[0]),.doutb(w_G18_37[1]),.doutc(w_G18_37[2]),.din(w_G18_12[0]));
	jspl3 jspl3_w_G18_38(.douta(w_G18_38[0]),.doutb(w_G18_38[1]),.doutc(w_G18_38[2]),.din(w_G18_12[1]));
	jspl3 jspl3_w_G18_39(.douta(w_G18_39[0]),.doutb(w_G18_39[1]),.doutc(w_G18_39[2]),.din(w_G18_12[2]));
	jspl3 jspl3_w_G18_40(.douta(w_G18_40[0]),.doutb(w_G18_40[1]),.doutc(w_G18_40[2]),.din(w_G18_13[0]));
	jspl3 jspl3_w_G18_41(.douta(w_G18_41[0]),.doutb(w_G18_41[1]),.doutc(w_G18_41[2]),.din(w_G18_13[1]));
	jspl3 jspl3_w_G18_42(.douta(w_G18_42[0]),.doutb(w_dff_A_jCHUc5Ti2_1),.doutc(w_G18_42[2]),.din(w_G18_13[2]));
	jspl3 jspl3_w_G18_43(.douta(w_G18_43[0]),.doutb(w_G18_43[1]),.doutc(w_G18_43[2]),.din(w_G18_14[0]));
	jspl3 jspl3_w_G18_44(.douta(w_G18_44[0]),.doutb(w_G18_44[1]),.doutc(w_G18_44[2]),.din(w_G18_14[1]));
	jspl3 jspl3_w_G18_45(.douta(w_G18_45[0]),.doutb(w_G18_45[1]),.doutc(w_G18_45[2]),.din(w_G18_14[2]));
	jspl3 jspl3_w_G18_46(.douta(w_G18_46[0]),.doutb(w_G18_46[1]),.doutc(w_G18_46[2]),.din(w_G18_15[0]));
	jspl3 jspl3_w_G18_47(.douta(w_G18_47[0]),.doutb(w_G18_47[1]),.doutc(w_G18_47[2]),.din(w_G18_15[1]));
	jspl3 jspl3_w_G18_48(.douta(w_G18_48[0]),.doutb(w_G18_48[1]),.doutc(w_G18_48[2]),.din(w_G18_15[2]));
	jspl3 jspl3_w_G18_49(.douta(w_G18_49[0]),.doutb(w_G18_49[1]),.doutc(w_dff_A_9oWdtRfv0_2),.din(w_G18_16[0]));
	jspl jspl_w_G29_0(.douta(w_dff_A_TcgSIRFV1_0),.doutb(w_G29_0[1]),.din(G29));
	jspl3 jspl3_w_G38_0(.douta(w_dff_A_LQdGDyaf3_0),.doutb(w_G38_0[1]),.doutc(w_dff_A_fc7Tr0NP2_2),.din(G38));
	jspl3 jspl3_w_G38_1(.douta(w_dff_A_bTX9z9f33_0),.doutb(w_dff_A_8FTKaedz4_1),.doutc(w_G38_1[2]),.din(w_G38_0[0]));
	jspl3 jspl3_w_G38_2(.douta(w_dff_A_y9fJLhst5_0),.doutb(w_dff_A_ZAY3sdbH0_1),.doutc(w_G38_2[2]),.din(w_G38_0[1]));
	jspl jspl_w_G41_0(.douta(w_dff_A_lQtzHlbT7_0),.doutb(w_G41_0[1]),.din(G41));
	jspl jspl_w_G70_0(.douta(w_G70_0[0]),.doutb(w_G70_0[1]),.din(G70));
	jspl jspl_w_G89_0(.douta(w_dff_A_VkhTzqs80_0),.doutb(w_G89_0[1]),.din(G89));
	jspl3 jspl3_w_G106_0(.douta(w_G106_0[0]),.doutb(w_G106_0[1]),.doutc(w_G106_0[2]),.din(G106));
	jspl jspl_w_G106_1(.douta(w_dff_A_hwt4BvMM2_0),.doutb(w_G106_1[1]),.din(w_G106_0[0]));
	jspl jspl_w_G209_0(.douta(w_G209_0[0]),.doutb(w_G209_0[1]),.din(w_dff_B_CaE08qKQ8_2));
	jspl jspl_w_G238_0(.douta(w_G238_0[0]),.doutb(w_G238_0[1]),.din(G238));
	jspl3 jspl3_w_G1455_0(.douta(w_G1455_0[0]),.doutb(w_G1455_0[1]),.doutc(w_G1455_0[2]),.din(G1455));
	jspl jspl_w_G1459_0(.douta(w_G1459_0[0]),.doutb(w_G1459_0[1]),.din(G1459));
	jspl jspl_w_G1462_0(.douta(w_G1462_0[0]),.doutb(w_G1462_0[1]),.din(G1462));
	jspl jspl_w_G1469_0(.douta(w_G1469_0[0]),.doutb(w_G1469_0[1]),.din(G1469));
	jspl3 jspl3_w_G1480_0(.douta(w_G1480_0[0]),.doutb(w_G1480_0[1]),.doutc(w_dff_A_rB8GOIbM9_2),.din(G1480));
	jspl jspl_w_G1486_0(.douta(w_G1486_0[0]),.doutb(w_G1486_0[1]),.din(G1486));
	jspl3 jspl3_w_G1492_0(.douta(w_G1492_0[0]),.doutb(w_G1492_0[1]),.doutc(w_dff_A_OMEH5hXN6_2),.din(G1492));
	jspl jspl_w_G1492_1(.douta(w_dff_A_mN4Y5ULW5_0),.doutb(w_G1492_1[1]),.din(w_G1492_0[0]));
	jspl3 jspl3_w_G1496_0(.douta(w_G1496_0[0]),.doutb(w_G1496_0[1]),.doutc(w_dff_A_J3NkEjqI6_2),.din(G1496));
	jspl jspl_w_G1496_1(.douta(w_G1496_1[0]),.doutb(w_G1496_1[1]),.din(w_G1496_0[0]));
	jspl3 jspl3_w_G2204_0(.douta(w_dff_A_izC37lvh5_0),.doutb(w_G2204_0[1]),.doutc(w_G2204_0[2]),.din(G2204));
	jspl jspl_w_G2208_0(.douta(w_G2208_0[0]),.doutb(w_G2208_0[1]),.din(G2208));
	jspl3 jspl3_w_G2211_0(.douta(w_G2211_0[0]),.doutb(w_dff_A_4jd6T85v2_1),.doutc(w_G2211_0[2]),.din(G2211));
	jspl3 jspl3_w_G2218_0(.douta(w_G2218_0[0]),.doutb(w_dff_A_ejDtG6IA4_1),.doutc(w_G2218_0[2]),.din(G2218));
	jspl3 jspl3_w_G2224_0(.douta(w_G2224_0[0]),.doutb(w_G2224_0[1]),.doutc(w_G2224_0[2]),.din(G2224));
	jspl jspl_w_G2224_1(.douta(w_dff_A_l1y0aVPn7_0),.doutb(w_G2224_1[1]),.din(w_G2224_0[0]));
	jspl3 jspl3_w_G2230_0(.douta(w_G2230_0[0]),.doutb(w_dff_A_Goj5lNI45_1),.doutc(w_G2230_0[2]),.din(G2230));
	jspl3 jspl3_w_G2236_0(.douta(w_G2236_0[0]),.doutb(w_G2236_0[1]),.doutc(w_G2236_0[2]),.din(G2236));
	jspl3 jspl3_w_G2239_0(.douta(w_G2239_0[0]),.doutb(w_G2239_0[1]),.doutc(w_dff_A_qd8jTaPx2_2),.din(G2239));
	jspl jspl_w_G2239_1(.douta(w_G2239_1[0]),.doutb(w_G2239_1[1]),.din(w_G2239_0[0]));
	jspl3 jspl3_w_G2247_0(.douta(w_G2247_0[0]),.doutb(w_G2247_0[1]),.doutc(w_G2247_0[2]),.din(G2247));
	jspl3 jspl3_w_G2253_0(.douta(w_G2253_0[0]),.doutb(w_dff_A_frfO4gwx4_1),.doutc(w_G2253_0[2]),.din(G2253));
	jspl jspl_w_G2256_0(.douta(w_G2256_0[0]),.doutb(w_G2256_0[1]),.din(G2256));
	jspl jspl_w_G3698_0(.douta(w_G3698_0[0]),.doutb(w_G3698_0[1]),.din(G3698));
	jspl3 jspl3_w_G3701_0(.douta(w_dff_A_abmFYAEM6_0),.doutb(w_G3701_0[1]),.doutc(w_G3701_0[2]),.din(G3701));
	jspl jspl_w_G3701_1(.douta(w_G3701_1[0]),.doutb(w_dff_A_8gH7ZCXd4_1),.din(w_G3701_0[0]));
	jspl3 jspl3_w_G3705_0(.douta(w_G3705_0[0]),.doutb(w_G3705_0[1]),.doutc(w_dff_A_BtE9KoFR5_2),.din(G3705));
	jspl3 jspl3_w_G3705_1(.douta(w_dff_A_0ekPl5pE5_0),.doutb(w_G3705_1[1]),.doutc(w_dff_A_JJz8ZuTB3_2),.din(w_G3705_0[0]));
	jspl jspl_w_G3711_0(.douta(w_G3711_0[0]),.doutb(w_G3711_0[1]),.din(G3711));
	jspl3 jspl3_w_G3717_0(.douta(w_G3717_0[0]),.doutb(w_dff_A_ky1Zb9sY5_1),.doutc(w_G3717_0[2]),.din(G3717));
	jspl3 jspl3_w_G3723_0(.douta(w_G3723_0[0]),.doutb(w_dff_A_EXeMCmjT5_1),.doutc(w_G3723_0[2]),.din(G3723));
	jspl3 jspl3_w_G3729_0(.douta(w_G3729_0[0]),.doutb(w_G3729_0[1]),.doutc(w_dff_A_d6USlwJ36_2),.din(G3729));
	jspl jspl_w_G3729_1(.douta(w_G3729_1[0]),.doutb(w_G3729_1[1]),.din(w_G3729_0[0]));
	jspl3 jspl3_w_G3737_0(.douta(w_G3737_0[0]),.doutb(w_dff_A_5JKO9HUY8_1),.doutc(w_G3737_0[2]),.din(G3737));
	jspl3 jspl3_w_G3743_0(.douta(w_G3743_0[0]),.doutb(w_dff_A_h7Gae4JC6_1),.doutc(w_G3743_0[2]),.din(G3743));
	jspl3 jspl3_w_G3749_0(.douta(w_G3749_0[0]),.doutb(w_dff_A_grsjDkSy3_1),.doutc(w_G3749_0[2]),.din(G3749));
	jspl jspl_w_G4393_0(.douta(w_G4393_0[0]),.doutb(w_G4393_0[1]),.din(G4393));
	jspl3 jspl3_w_G4394_0(.douta(w_G4394_0[0]),.doutb(w_G4394_0[1]),.doutc(w_dff_A_IutNNJpv4_2),.din(G4394));
	jspl jspl_w_G4394_1(.douta(w_G4394_1[0]),.doutb(w_G4394_1[1]),.din(w_G4394_0[0]));
	jspl3 jspl3_w_G4400_0(.douta(w_G4400_0[0]),.doutb(w_G4400_0[1]),.doutc(w_G4400_0[2]),.din(G4400));
	jspl jspl_w_G4400_1(.douta(w_dff_A_sFIkmB0G0_0),.doutb(w_G4400_1[1]),.din(w_G4400_0[0]));
	jspl3 jspl3_w_G4405_0(.douta(w_G4405_0[0]),.doutb(w_G4405_0[1]),.doutc(w_G4405_0[2]),.din(G4405));
	jspl jspl_w_G4405_1(.douta(w_dff_A_lTrelQPG1_0),.doutb(w_G4405_1[1]),.din(w_G4405_0[0]));
	jspl3 jspl3_w_G4410_0(.douta(w_G4410_0[0]),.doutb(w_dff_A_9wSeb58Q6_1),.doutc(w_G4410_0[2]),.din(G4410));
	jspl3 jspl3_w_G4415_0(.douta(w_G4415_0[0]),.doutb(w_G4415_0[1]),.doutc(w_G4415_0[2]),.din(G4415));
	jspl jspl_w_G4415_1(.douta(w_dff_A_lnZFptbP4_0),.doutb(w_G4415_1[1]),.din(w_G4415_0[0]));
	jspl3 jspl3_w_G4420_0(.douta(w_G4420_0[0]),.doutb(w_G4420_0[1]),.doutc(w_G4420_0[2]),.din(G4420));
	jspl jspl_w_G4420_1(.douta(w_dff_A_HBJIOJCi0_0),.doutb(w_G4420_1[1]),.din(w_G4420_0[0]));
	jspl3 jspl3_w_G4427_0(.douta(w_G4427_0[0]),.doutb(w_G4427_0[1]),.doutc(w_G4427_0[2]),.din(G4427));
	jspl3 jspl3_w_G4432_0(.douta(w_G4432_0[0]),.doutb(w_dff_A_7nXfocmh8_1),.doutc(w_G4432_0[2]),.din(G4432));
	jspl3 jspl3_w_G4437_0(.douta(w_G4437_0[0]),.doutb(w_dff_A_4CLa4k1Y8_1),.doutc(w_G4437_0[2]),.din(G4437));
	jspl3 jspl3_w_G4526_0(.douta(w_G4526_0[0]),.doutb(w_dff_A_pSxPcOGY3_1),.doutc(w_dff_A_1RvgfV2T7_2),.din(G4526));
	jspl3 jspl3_w_G4526_1(.douta(w_dff_A_ehAwgVB08_0),.doutb(w_G4526_1[1]),.doutc(w_dff_A_M7wVrncw9_2),.din(w_G4526_0[0]));
	jspl3 jspl3_w_G4526_2(.douta(w_dff_A_BzVI7Hmc4_0),.doutb(w_dff_A_KEpOUmLI6_1),.doutc(w_G4526_2[2]),.din(w_G4526_0[1]));
	jspl3 jspl3_w_G4528_0(.douta(w_G4528_0[0]),.doutb(w_G4528_0[1]),.doutc(w_G4528_0[2]),.din(G4528));
	jspl jspl_w_G404_0(.douta(w_G404_0),.doutb(w_dff_A_J1N7OnNX3_1),.din(G404_fa_));
	jspl jspl_w_G406_0(.douta(w_G406_0),.doutb(w_dff_A_vKZYkuMo0_1),.din(G406_fa_));
	jspl jspl_w_G408_0(.douta(w_G408_0),.doutb(w_dff_A_pWywJuT40_1),.din(G408_fa_));
	jspl jspl_w_G410_0(.douta(w_G410_0),.doutb(w_dff_A_4rlRYtVI6_1),.din(G410_fa_));
	jspl jspl_w_G412_0(.douta(w_G412_0),.doutb(w_dff_A_CNbvXIlX4_1),.din(G412_fa_));
	jspl jspl_w_G414_0(.douta(w_dff_A_1UvK5pWl9_0),.doutb(w_dff_A_UmDLHC9r2_1),.din(G414_fa_));
	jspl jspl_w_G416_0(.douta(w_G416_0),.doutb(w_dff_A_R88Dkp5e7_1),.din(G416_fa_));
	jspl jspl_w_G252_0(.douta(w_G252_0),.doutb(w_dff_A_0iaYpmVK7_1),.din(G252_fa_));
	jspl jspl_w_n345_0(.douta(w_n345_0[0]),.doutb(w_n345_0[1]),.din(n345));
	jspl jspl_w_n347_0(.douta(w_n347_0[0]),.doutb(w_n347_0[1]),.din(w_dff_B_zOw0FkEF5_2));
	jspl jspl_w_n349_0(.douta(w_n349_0[0]),.doutb(w_n349_0[1]),.din(n349));
	jspl jspl_w_n353_0(.douta(w_n353_0[0]),.doutb(w_n353_0[1]),.din(n353));
	jspl3 jspl3_w_n354_0(.douta(w_n354_0[0]),.doutb(w_n354_0[1]),.doutc(w_n354_0[2]),.din(w_dff_B_oEDRfFsY6_3));
	jspl3 jspl3_w_n355_0(.douta(w_n355_0[0]),.doutb(w_n355_0[1]),.doutc(w_n355_0[2]),.din(n355));
	jspl3 jspl3_w_n355_1(.douta(w_n355_1[0]),.doutb(w_n355_1[1]),.doutc(w_n355_1[2]),.din(w_n355_0[0]));
	jspl3 jspl3_w_n355_2(.douta(w_n355_2[0]),.doutb(w_n355_2[1]),.doutc(w_n355_2[2]),.din(w_n355_0[1]));
	jspl3 jspl3_w_n355_3(.douta(w_n355_3[0]),.doutb(w_n355_3[1]),.doutc(w_n355_3[2]),.din(w_n355_0[2]));
	jspl3 jspl3_w_n355_4(.douta(w_n355_4[0]),.doutb(w_n355_4[1]),.doutc(w_n355_4[2]),.din(w_n355_1[0]));
	jspl3 jspl3_w_n355_5(.douta(w_n355_5[0]),.doutb(w_n355_5[1]),.doutc(w_n355_5[2]),.din(w_n355_1[1]));
	jspl3 jspl3_w_n355_6(.douta(w_n355_6[0]),.doutb(w_n355_6[1]),.doutc(w_n355_6[2]),.din(w_n355_1[2]));
	jspl3 jspl3_w_n355_7(.douta(w_n355_7[0]),.doutb(w_n355_7[1]),.doutc(w_n355_7[2]),.din(w_n355_2[0]));
	jspl3 jspl3_w_n355_8(.douta(w_n355_8[0]),.doutb(w_n355_8[1]),.doutc(w_n355_8[2]),.din(w_n355_2[1]));
	jspl3 jspl3_w_n355_9(.douta(w_n355_9[0]),.doutb(w_n355_9[1]),.doutc(w_n355_9[2]),.din(w_n355_2[2]));
	jspl3 jspl3_w_n355_10(.douta(w_n355_10[0]),.doutb(w_n355_10[1]),.doutc(w_n355_10[2]),.din(w_n355_3[0]));
	jspl3 jspl3_w_n355_11(.douta(w_n355_11[0]),.doutb(w_n355_11[1]),.doutc(w_n355_11[2]),.din(w_n355_3[1]));
	jspl3 jspl3_w_n355_12(.douta(w_n355_12[0]),.doutb(w_dff_A_QYDi2JN64_1),.doutc(w_n355_12[2]),.din(w_n355_3[2]));
	jspl3 jspl3_w_n355_13(.douta(w_n355_13[0]),.doutb(w_n355_13[1]),.doutc(w_n355_13[2]),.din(w_n355_4[0]));
	jspl3 jspl3_w_n355_14(.douta(w_n355_14[0]),.doutb(w_n355_14[1]),.doutc(w_n355_14[2]),.din(w_n355_4[1]));
	jspl3 jspl3_w_n355_15(.douta(w_n355_15[0]),.doutb(w_n355_15[1]),.doutc(w_n355_15[2]),.din(w_n355_4[2]));
	jspl3 jspl3_w_n355_16(.douta(w_n355_16[0]),.doutb(w_n355_16[1]),.doutc(w_n355_16[2]),.din(w_n355_5[0]));
	jspl3 jspl3_w_n355_17(.douta(w_n355_17[0]),.doutb(w_n355_17[1]),.doutc(w_n355_17[2]),.din(w_n355_5[1]));
	jspl3 jspl3_w_n355_18(.douta(w_n355_18[0]),.doutb(w_n355_18[1]),.doutc(w_n355_18[2]),.din(w_n355_5[2]));
	jspl3 jspl3_w_n355_19(.douta(w_n355_19[0]),.doutb(w_n355_19[1]),.doutc(w_n355_19[2]),.din(w_n355_6[0]));
	jspl3 jspl3_w_n355_20(.douta(w_n355_20[0]),.doutb(w_n355_20[1]),.doutc(w_n355_20[2]),.din(w_n355_6[1]));
	jspl3 jspl3_w_n355_21(.douta(w_n355_21[0]),.doutb(w_n355_21[1]),.doutc(w_n355_21[2]),.din(w_n355_6[2]));
	jspl3 jspl3_w_n355_22(.douta(w_n355_22[0]),.doutb(w_n355_22[1]),.doutc(w_n355_22[2]),.din(w_n355_7[0]));
	jspl3 jspl3_w_n355_23(.douta(w_n355_23[0]),.doutb(w_n355_23[1]),.doutc(w_n355_23[2]),.din(w_n355_7[1]));
	jspl3 jspl3_w_n355_24(.douta(w_n355_24[0]),.doutb(w_n355_24[1]),.doutc(w_n355_24[2]),.din(w_n355_7[2]));
	jspl3 jspl3_w_n355_25(.douta(w_n355_25[0]),.doutb(w_n355_25[1]),.doutc(w_n355_25[2]),.din(w_n355_8[0]));
	jspl3 jspl3_w_n355_26(.douta(w_n355_26[0]),.doutb(w_n355_26[1]),.doutc(w_n355_26[2]),.din(w_n355_8[1]));
	jspl3 jspl3_w_n355_27(.douta(w_n355_27[0]),.doutb(w_n355_27[1]),.doutc(w_n355_27[2]),.din(w_n355_8[2]));
	jspl3 jspl3_w_n355_28(.douta(w_n355_28[0]),.doutb(w_n355_28[1]),.doutc(w_n355_28[2]),.din(w_n355_9[0]));
	jspl3 jspl3_w_n355_29(.douta(w_n355_29[0]),.doutb(w_n355_29[1]),.doutc(w_n355_29[2]),.din(w_n355_9[1]));
	jspl3 jspl3_w_n355_30(.douta(w_n355_30[0]),.doutb(w_n355_30[1]),.doutc(w_n355_30[2]),.din(w_n355_9[2]));
	jspl3 jspl3_w_n355_31(.douta(w_n355_31[0]),.doutb(w_n355_31[1]),.doutc(w_n355_31[2]),.din(w_n355_10[0]));
	jspl3 jspl3_w_n355_32(.douta(w_n355_32[0]),.doutb(w_n355_32[1]),.doutc(w_n355_32[2]),.din(w_n355_10[1]));
	jspl3 jspl3_w_n355_33(.douta(w_n355_33[0]),.doutb(w_n355_33[1]),.doutc(w_n355_33[2]),.din(w_n355_10[2]));
	jspl3 jspl3_w_n355_34(.douta(w_n355_34[0]),.doutb(w_n355_34[1]),.doutc(w_n355_34[2]),.din(w_n355_11[0]));
	jspl3 jspl3_w_n355_35(.douta(w_n355_35[0]),.doutb(w_n355_35[1]),.doutc(w_n355_35[2]),.din(w_n355_11[1]));
	jspl jspl_w_n357_0(.douta(w_dff_A_6OPMGmh60_0),.doutb(w_n357_0[1]),.din(n357));
	jspl jspl_w_n358_0(.douta(w_n358_0[0]),.doutb(w_n358_0[1]),.din(n358));
	jspl3 jspl3_w_n359_0(.douta(w_n359_0[0]),.doutb(w_n359_0[1]),.doutc(w_n359_0[2]),.din(n359));
	jspl jspl_w_n359_1(.douta(w_n359_1[0]),.doutb(w_n359_1[1]),.din(w_n359_0[0]));
	jspl3 jspl3_w_n361_0(.douta(w_dff_A_T1F6XDXd7_0),.doutb(w_n361_0[1]),.doutc(w_n361_0[2]),.din(n361));
	jspl3 jspl3_w_n362_0(.douta(w_n362_0[0]),.doutb(w_n362_0[1]),.doutc(w_n362_0[2]),.din(n362));
	jspl3 jspl3_w_n363_0(.douta(w_n363_0[0]),.doutb(w_n363_0[1]),.doutc(w_dff_A_IK4xxIxf6_2),.din(w_dff_B_cbk2BWzk1_3));
	jspl3 jspl3_w_n364_0(.douta(w_dff_A_5c0RCyZl8_0),.doutb(w_n364_0[1]),.doutc(w_n364_0[2]),.din(n364));
	jspl3 jspl3_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.doutc(w_dff_A_YDtMt7ws4_2),.din(n366));
	jspl jspl_w_n367_0(.douta(w_n367_0[0]),.doutb(w_n367_0[1]),.din(n367));
	jspl jspl_w_n368_0(.douta(w_n368_0[0]),.doutb(w_n368_0[1]),.din(n368));
	jspl jspl_w_n369_0(.douta(w_n369_0[0]),.doutb(w_n369_0[1]),.din(n369));
	jspl3 jspl3_w_n370_0(.douta(w_dff_A_pwqs1dkK6_0),.doutb(w_dff_A_mIsh5nKZ1_1),.doutc(w_n370_0[2]),.din(w_dff_B_CQ4A5VLN4_3));
	jspl3 jspl3_w_n371_0(.douta(w_n371_0[0]),.doutb(w_dff_A_SuyAG6dD7_1),.doutc(w_dff_A_Zkr9sd264_2),.din(n371));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.din(n372));
	jspl3 jspl3_w_n373_0(.douta(w_n373_0[0]),.doutb(w_n373_0[1]),.doutc(w_n373_0[2]),.din(n373));
	jspl3 jspl3_w_n373_1(.douta(w_n373_1[0]),.doutb(w_n373_1[1]),.doutc(w_n373_1[2]),.din(w_n373_0[0]));
	jspl3 jspl3_w_n373_2(.douta(w_n373_2[0]),.doutb(w_n373_2[1]),.doutc(w_n373_2[2]),.din(w_n373_0[1]));
	jspl3 jspl3_w_n373_3(.douta(w_dff_A_qESbXHkL9_0),.doutb(w_n373_3[1]),.doutc(w_n373_3[2]),.din(w_n373_0[2]));
	jspl3 jspl3_w_n373_4(.douta(w_n373_4[0]),.doutb(w_n373_4[1]),.doutc(w_n373_4[2]),.din(w_n373_1[0]));
	jspl3 jspl3_w_n373_5(.douta(w_n373_5[0]),.doutb(w_n373_5[1]),.doutc(w_dff_A_KqBYPGeX1_2),.din(w_n373_1[1]));
	jspl3 jspl3_w_n373_6(.douta(w_n373_6[0]),.doutb(w_n373_6[1]),.doutc(w_n373_6[2]),.din(w_n373_1[2]));
	jspl3 jspl3_w_n373_7(.douta(w_n373_7[0]),.doutb(w_n373_7[1]),.doutc(w_n373_7[2]),.din(w_n373_2[0]));
	jspl3 jspl3_w_n373_8(.douta(w_n373_8[0]),.doutb(w_n373_8[1]),.doutc(w_n373_8[2]),.din(w_n373_2[1]));
	jspl3 jspl3_w_n373_9(.douta(w_n373_9[0]),.doutb(w_n373_9[1]),.doutc(w_n373_9[2]),.din(w_n373_2[2]));
	jspl jspl_w_n374_0(.douta(w_dff_A_MM8c0lGK3_0),.doutb(w_n374_0[1]),.din(n374));
	jspl3 jspl3_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.doutc(w_n375_0[2]),.din(n375));
	jspl3 jspl3_w_n377_0(.douta(w_dff_A_unS6yNBJ5_0),.doutb(w_n377_0[1]),.doutc(w_dff_A_GJFWv1ec1_2),.din(n377));
	jspl3 jspl3_w_n377_1(.douta(w_dff_A_f4rNf0jd1_0),.doutb(w_n377_1[1]),.doutc(w_dff_A_Cek6xykY5_2),.din(w_n377_0[0]));
	jspl jspl_w_n378_0(.douta(w_dff_A_e43K4zLq2_0),.doutb(w_n378_0[1]),.din(n378));
	jspl3 jspl3_w_n379_0(.douta(w_n379_0[0]),.doutb(w_n379_0[1]),.doutc(w_n379_0[2]),.din(n379));
	jspl jspl_w_n380_0(.douta(w_n380_0[0]),.doutb(w_n380_0[1]),.din(n380));
	jspl3 jspl3_w_n383_0(.douta(w_n383_0[0]),.doutb(w_dff_A_Dr6I3zdZ5_1),.doutc(w_dff_A_6dGCM4iH7_2),.din(n383));
	jspl jspl_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.din(w_dff_B_RleEmAtv9_2));
	jspl jspl_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.din(n386));
	jspl3 jspl3_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.doutc(w_n387_0[2]),.din(n387));
	jspl jspl_w_n387_1(.douta(w_n387_1[0]),.doutb(w_n387_1[1]),.din(w_n387_0[0]));
	jspl3 jspl3_w_n388_0(.douta(w_n388_0[0]),.doutb(w_n388_0[1]),.doutc(w_n388_0[2]),.din(n388));
	jspl3 jspl3_w_n388_1(.douta(w_dff_A_d1f47uPV5_0),.doutb(w_n388_1[1]),.doutc(w_dff_A_esoiYOnO9_2),.din(w_n388_0[0]));
	jspl3 jspl3_w_n389_0(.douta(w_dff_A_sDvOWC695_0),.doutb(w_dff_A_8hA8yP7X7_1),.doutc(w_n389_0[2]),.din(n389));
	jspl jspl_w_n389_1(.douta(w_n389_1[0]),.doutb(w_n389_1[1]),.din(w_n389_0[0]));
	jspl3 jspl3_w_n391_0(.douta(w_n391_0[0]),.doutb(w_n391_0[1]),.doutc(w_n391_0[2]),.din(n391));
	jspl3 jspl3_w_n392_0(.douta(w_dff_A_Hs3YZ0n28_0),.doutb(w_n392_0[1]),.doutc(w_n392_0[2]),.din(n392));
	jspl3 jspl3_w_n393_0(.douta(w_dff_A_0ZPv1UgA1_0),.doutb(w_dff_A_zqEgeehC9_1),.doutc(w_n393_0[2]),.din(n393));
	jspl jspl_w_n393_1(.douta(w_n393_1[0]),.doutb(w_n393_1[1]),.din(w_n393_0[0]));
	jspl jspl_w_n394_0(.douta(w_n394_0[0]),.doutb(w_n394_0[1]),.din(n394));
	jspl3 jspl3_w_n395_0(.douta(w_n395_0[0]),.doutb(w_n395_0[1]),.doutc(w_n395_0[2]),.din(n395));
	jspl jspl_w_n395_1(.douta(w_n395_1[0]),.doutb(w_n395_1[1]),.din(w_n395_0[0]));
	jspl3 jspl3_w_n396_0(.douta(w_n396_0[0]),.doutb(w_n396_0[1]),.doutc(w_n396_0[2]),.din(n396));
	jspl3 jspl3_w_n396_1(.douta(w_n396_1[0]),.doutb(w_n396_1[1]),.doutc(w_n396_1[2]),.din(w_n396_0[0]));
	jspl jspl_w_n397_0(.douta(w_n397_0[0]),.doutb(w_n397_0[1]),.din(n397));
	jspl3 jspl3_w_n405_0(.douta(w_dff_A_TIdTR1mS2_0),.doutb(w_dff_A_SX3eBsGe0_1),.doutc(w_n405_0[2]),.din(n405));
	jspl jspl_w_n407_0(.douta(w_n407_0[0]),.doutb(w_n407_0[1]),.din(n407));
	jspl3 jspl3_w_n409_0(.douta(w_n409_0[0]),.doutb(w_n409_0[1]),.doutc(w_dff_A_DhCr42MS9_2),.din(n409));
	jspl jspl_w_n409_1(.douta(w_n409_1[0]),.doutb(w_n409_1[1]),.din(w_n409_0[0]));
	jspl3 jspl3_w_n411_0(.douta(w_n411_0[0]),.doutb(w_n411_0[1]),.doutc(w_dff_A_Fb0cOCXF9_2),.din(n411));
	jspl jspl_w_n411_1(.douta(w_n411_1[0]),.doutb(w_n411_1[1]),.din(w_n411_0[0]));
	jspl3 jspl3_w_n413_0(.douta(w_n413_0[0]),.doutb(w_n413_0[1]),.doutc(w_n413_0[2]),.din(n413));
	jspl jspl_w_n413_1(.douta(w_dff_A_MnDcgg263_0),.doutb(w_n413_1[1]),.din(w_n413_0[0]));
	jspl3 jspl3_w_n414_0(.douta(w_n414_0[0]),.doutb(w_dff_A_drh3cEUA6_1),.doutc(w_n414_0[2]),.din(n414));
	jspl jspl_w_n414_1(.douta(w_n414_1[0]),.doutb(w_n414_1[1]),.din(w_n414_0[0]));
	jspl jspl_w_n415_0(.douta(w_n415_0[0]),.doutb(w_n415_0[1]),.din(n415));
	jspl3 jspl3_w_n416_0(.douta(w_n416_0[0]),.doutb(w_dff_A_alS2OU0O7_1),.doutc(w_n416_0[2]),.din(n416));
	jspl jspl_w_n418_0(.douta(w_dff_A_1E9O2vqX7_0),.doutb(w_n418_0[1]),.din(n418));
	jspl jspl_w_n419_0(.douta(w_n419_0[0]),.doutb(w_dff_A_KHAYfGor3_1),.din(n419));
	jspl jspl_w_n420_0(.douta(w_n420_0[0]),.doutb(w_dff_A_8rcwYPhX6_1),.din(n420));
	jspl3 jspl3_w_n421_0(.douta(w_n421_0[0]),.doutb(w_dff_A_AczDAVgJ8_1),.doutc(w_dff_A_0BKpP0JF3_2),.din(n421));
	jspl jspl_w_n422_0(.douta(w_dff_A_LlyypmAA3_0),.doutb(w_n422_0[1]),.din(n422));
	jspl3 jspl3_w_n423_0(.douta(w_n423_0[0]),.doutb(w_n423_0[1]),.doutc(w_n423_0[2]),.din(n423));
	jspl jspl_w_n424_0(.douta(w_n424_0[0]),.doutb(w_dff_A_CSmNRdhO9_1),.din(n424));
	jspl3 jspl3_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.doutc(w_dff_A_Inqk3ZfN9_2),.din(n425));
	jspl jspl_w_n425_1(.douta(w_n425_1[0]),.doutb(w_dff_A_YgznzAnD1_1),.din(w_n425_0[0]));
	jspl3 jspl3_w_n426_0(.douta(w_n426_0[0]),.doutb(w_dff_A_pev09nyh0_1),.doutc(w_dff_A_jXiXJTM48_2),.din(n426));
	jspl jspl_w_n427_0(.douta(w_dff_A_LH9Vwqk78_0),.doutb(w_n427_0[1]),.din(n427));
	jspl3 jspl3_w_n428_0(.douta(w_n428_0[0]),.doutb(w_n428_0[1]),.doutc(w_n428_0[2]),.din(n428));
	jspl3 jspl3_w_n429_0(.douta(w_n429_0[0]),.doutb(w_dff_A_9jLdaajW3_1),.doutc(w_dff_A_3hHbEkJw4_2),.din(n429));
	jspl jspl_w_n430_0(.douta(w_n430_0[0]),.doutb(w_n430_0[1]),.din(w_dff_B_yLX4YxfI0_2));
	jspl jspl_w_n431_0(.douta(w_dff_A_xlQYpSbL7_0),.doutb(w_n431_0[1]),.din(n431));
	jspl3 jspl3_w_n432_0(.douta(w_n432_0[0]),.doutb(w_n432_0[1]),.doutc(w_n432_0[2]),.din(n432));
	jspl3 jspl3_w_n433_0(.douta(w_n433_0[0]),.doutb(w_n433_0[1]),.doutc(w_dff_A_HEOQgHfq2_2),.din(n433));
	jspl3 jspl3_w_n433_1(.douta(w_dff_A_30iM3TXy2_0),.doutb(w_n433_1[1]),.doutc(w_n433_1[2]),.din(w_n433_0[0]));
	jspl jspl_w_n434_0(.douta(w_n434_0[0]),.doutb(w_n434_0[1]),.din(w_dff_B_pwi9h59w5_2));
	jspl jspl_w_n435_0(.douta(w_dff_A_9dsEoGvg6_0),.doutb(w_n435_0[1]),.din(n435));
	jspl3 jspl3_w_n436_0(.douta(w_n436_0[0]),.doutb(w_n436_0[1]),.doutc(w_n436_0[2]),.din(n436));
	jspl3 jspl3_w_n437_0(.douta(w_n437_0[0]),.doutb(w_dff_A_tq65jwS84_1),.doutc(w_n437_0[2]),.din(n437));
	jspl jspl_w_n438_0(.douta(w_dff_A_ZCXL6AFb6_0),.doutb(w_n438_0[1]),.din(n438));
	jspl jspl_w_n440_0(.douta(w_n440_0[0]),.doutb(w_n440_0[1]),.din(n440));
	jspl3 jspl3_w_n444_0(.douta(w_n444_0[0]),.doutb(w_dff_A_a66fwNCD5_1),.doutc(w_dff_A_CO40dOUl0_2),.din(n444));
	jspl3 jspl3_w_n445_0(.douta(w_n445_0[0]),.doutb(w_dff_A_OaUA8Du73_1),.doutc(w_n445_0[2]),.din(n445));
	jspl3 jspl3_w_n447_0(.douta(w_n447_0[0]),.doutb(w_dff_A_RFn9ktMs9_1),.doutc(w_n447_0[2]),.din(n447));
	jspl3 jspl3_w_n449_0(.douta(w_n449_0[0]),.doutb(w_n449_0[1]),.doutc(w_n449_0[2]),.din(n449));
	jspl jspl_w_n449_1(.douta(w_dff_A_DJvvuMLZ3_0),.doutb(w_n449_1[1]),.din(w_n449_0[0]));
	jspl3 jspl3_w_n450_0(.douta(w_n450_0[0]),.doutb(w_n450_0[1]),.doutc(w_dff_A_DNUoJNJS9_2),.din(n450));
	jspl3 jspl3_w_n451_0(.douta(w_n451_0[0]),.doutb(w_n451_0[1]),.doutc(w_n451_0[2]),.din(w_dff_B_bNAyFE7f2_3));
	jspl3 jspl3_w_n453_0(.douta(w_n453_0[0]),.doutb(w_dff_A_awJpdhdt3_1),.doutc(w_n453_0[2]),.din(n453));
	jspl jspl_w_n453_1(.douta(w_n453_1[0]),.doutb(w_n453_1[1]),.din(w_n453_0[0]));
	jspl3 jspl3_w_n456_0(.douta(w_n456_0[0]),.doutb(w_dff_A_GH49b0Su4_1),.doutc(w_dff_A_ma0gtraA9_2),.din(n456));
	jspl jspl_w_n457_0(.douta(w_n457_0[0]),.doutb(w_n457_0[1]),.din(n457));
	jspl3 jspl3_w_n459_0(.douta(w_n459_0[0]),.doutb(w_n459_0[1]),.doutc(w_n459_0[2]),.din(n459));
	jspl3 jspl3_w_n460_0(.douta(w_n460_0[0]),.doutb(w_dff_A_oMDMfYxR4_1),.doutc(w_dff_A_qlnCXpzK1_2),.din(n460));
	jspl3 jspl3_w_n460_1(.douta(w_dff_A_mzPJmmpA5_0),.doutb(w_dff_A_N4yhrShC2_1),.doutc(w_n460_1[2]),.din(w_n460_0[0]));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_dff_A_KeAGqp0V3_1),.doutc(w_dff_A_9UTW68s00_2),.din(n462));
	jspl3 jspl3_w_n463_0(.douta(w_n463_0[0]),.doutb(w_dff_A_OOnyHpnr0_1),.doutc(w_dff_A_23iTfWE05_2),.din(n463));
	jspl jspl_w_n463_1(.douta(w_dff_A_mm9xl4ny1_0),.doutb(w_n463_1[1]),.din(w_n463_0[0]));
	jspl3 jspl3_w_n464_0(.douta(w_n464_0[0]),.doutb(w_dff_A_k81yAa526_1),.doutc(w_n464_0[2]),.din(n464));
	jspl jspl_w_n465_0(.douta(w_n465_0[0]),.doutb(w_dff_A_AEtra7w43_1),.din(w_dff_B_8NkWGC5a1_2));
	jspl jspl_w_n466_0(.douta(w_n466_0[0]),.doutb(w_n466_0[1]),.din(w_dff_B_faLwkV1V1_2));
	jspl jspl_w_n467_0(.douta(w_n467_0[0]),.doutb(w_n467_0[1]),.din(n467));
	jspl3 jspl3_w_n469_0(.douta(w_n469_0[0]),.doutb(w_dff_A_2iW2PPZY8_1),.doutc(w_n469_0[2]),.din(n469));
	jspl jspl_w_n469_1(.douta(w_n469_1[0]),.doutb(w_n469_1[1]),.din(w_n469_0[0]));
	jspl3 jspl3_w_n470_0(.douta(w_n470_0[0]),.doutb(w_dff_A_T7jq9jDO9_1),.doutc(w_dff_A_bhpvO7y81_2),.din(n470));
	jspl3 jspl3_w_n471_0(.douta(w_n471_0[0]),.doutb(w_dff_A_AEUcQ3Nn0_1),.doutc(w_dff_A_CoRA3fFb5_2),.din(n471));
	jspl jspl_w_n472_0(.douta(w_n472_0[0]),.doutb(w_n472_0[1]),.din(n472));
	jspl3 jspl3_w_n474_0(.douta(w_n474_0[0]),.doutb(w_n474_0[1]),.doutc(w_n474_0[2]),.din(n474));
	jspl3 jspl3_w_n475_0(.douta(w_n475_0[0]),.doutb(w_dff_A_iNqFcuDB5_1),.doutc(w_n475_0[2]),.din(n475));
	jspl3 jspl3_w_n476_0(.douta(w_n476_0[0]),.doutb(w_dff_A_nz0WVmC46_1),.doutc(w_dff_A_1SPzV9KS9_2),.din(n476));
	jspl jspl_w_n477_0(.douta(w_n477_0[0]),.doutb(w_n477_0[1]),.din(n477));
	jspl3 jspl3_w_n479_0(.douta(w_n479_0[0]),.doutb(w_n479_0[1]),.doutc(w_n479_0[2]),.din(n479));
	jspl jspl_w_n479_1(.douta(w_n479_1[0]),.doutb(w_n479_1[1]),.din(w_n479_0[0]));
	jspl3 jspl3_w_n480_0(.douta(w_n480_0[0]),.doutb(w_n480_0[1]),.doutc(w_dff_A_qzEOAB5K5_2),.din(n480));
	jspl jspl_w_n480_1(.douta(w_n480_1[0]),.doutb(w_n480_1[1]),.din(w_n480_0[0]));
	jspl jspl_w_n481_0(.douta(w_dff_A_PjQxVjRq2_0),.doutb(w_n481_0[1]),.din(n481));
	jspl jspl_w_n485_0(.douta(w_n485_0[0]),.doutb(w_n485_0[1]),.din(n485));
	jspl jspl_w_n486_0(.douta(w_n486_0[0]),.doutb(w_n486_0[1]),.din(n486));
	jspl3 jspl3_w_n487_0(.douta(w_n487_0[0]),.doutb(w_dff_A_AdtOCzBY1_1),.doutc(w_n487_0[2]),.din(n487));
	jspl3 jspl3_w_n489_0(.douta(w_n489_0[0]),.doutb(w_n489_0[1]),.doutc(w_n489_0[2]),.din(n489));
	jspl3 jspl3_w_n491_0(.douta(w_n491_0[0]),.doutb(w_n491_0[1]),.doutc(w_dff_A_VKErXlhW5_2),.din(n491));
	jspl jspl_w_n491_1(.douta(w_dff_A_LLfcPI5v9_0),.doutb(w_n491_1[1]),.din(w_n491_0[0]));
	jspl3 jspl3_w_n495_0(.douta(w_n495_0[0]),.doutb(w_n495_0[1]),.doutc(w_n495_0[2]),.din(n495));
	jspl jspl_w_n495_1(.douta(w_dff_A_i8ufmyLE3_0),.doutb(w_n495_1[1]),.din(w_n495_0[0]));
	jspl3 jspl3_w_n496_0(.douta(w_n496_0[0]),.doutb(w_n496_0[1]),.doutc(w_n496_0[2]),.din(n496));
	jspl3 jspl3_w_n497_0(.douta(w_n497_0[0]),.doutb(w_n497_0[1]),.doutc(w_n497_0[2]),.din(n497));
	jspl jspl_w_n497_1(.douta(w_dff_A_VJ2PfoYk9_0),.doutb(w_n497_1[1]),.din(w_n497_0[0]));
	jspl jspl_w_n499_0(.douta(w_n499_0[0]),.doutb(w_dff_A_msWSaFgt3_1),.din(n499));
	jspl jspl_w_n500_0(.douta(w_n500_0[0]),.doutb(w_dff_A_DKf7sUZJ4_1),.din(n500));
	jspl3 jspl3_w_n501_0(.douta(w_dff_A_jggx32xI4_0),.doutb(w_n501_0[1]),.doutc(w_dff_A_2cU5pr8u4_2),.din(n501));
	jspl jspl_w_n503_0(.douta(w_n503_0[0]),.doutb(w_n503_0[1]),.din(n503));
	jspl3 jspl3_w_n504_0(.douta(w_n504_0[0]),.doutb(w_n504_0[1]),.doutc(w_dff_A_9g2qfnBI4_2),.din(n504));
	jspl jspl_w_n504_1(.douta(w_n504_1[0]),.doutb(w_n504_1[1]),.din(w_n504_0[0]));
	jspl jspl_w_n505_0(.douta(w_n505_0[0]),.doutb(w_dff_A_xavBH0ie1_1),.din(n505));
	jspl jspl_w_n507_0(.douta(w_dff_A_aJryGNPj1_0),.doutb(w_n507_0[1]),.din(n507));
	jspl3 jspl3_w_n509_0(.douta(w_n509_0[0]),.doutb(w_dff_A_iDCFiOTb3_1),.doutc(w_dff_A_eBZdL6T88_2),.din(n509));
	jspl jspl_w_n511_0(.douta(w_n511_0[0]),.doutb(w_n511_0[1]),.din(n511));
	jspl3 jspl3_w_n512_0(.douta(w_n512_0[0]),.doutb(w_n512_0[1]),.doutc(w_n512_0[2]),.din(n512));
	jspl3 jspl3_w_n513_0(.douta(w_n513_0[0]),.doutb(w_n513_0[1]),.doutc(w_dff_A_mEQNs6C42_2),.din(n513));
	jspl jspl_w_n513_1(.douta(w_n513_1[0]),.doutb(w_dff_A_cC4jDxwZ0_1),.din(w_n513_0[0]));
	jspl jspl_w_n514_0(.douta(w_n514_0[0]),.doutb(w_n514_0[1]),.din(w_dff_B_V2dp9oao7_2));
	jspl jspl_w_n516_0(.douta(w_n516_0[0]),.doutb(w_n516_0[1]),.din(n516));
	jspl3 jspl3_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.doutc(w_n517_0[2]),.din(n517));
	jspl jspl_w_n517_1(.douta(w_n517_1[0]),.doutb(w_n517_1[1]),.din(w_n517_0[0]));
	jspl3 jspl3_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.doutc(w_n518_0[2]),.din(n518));
	jspl3 jspl3_w_n518_1(.douta(w_dff_A_5oso5I1j9_0),.doutb(w_n518_1[1]),.doutc(w_n518_1[2]),.din(w_n518_0[0]));
	jspl jspl_w_n520_0(.douta(w_n520_0[0]),.doutb(w_n520_0[1]),.din(w_dff_B_9w2r0qCf1_2));
	jspl jspl_w_n522_0(.douta(w_n522_0[0]),.doutb(w_n522_0[1]),.din(n522));
	jspl3 jspl3_w_n523_0(.douta(w_n523_0[0]),.doutb(w_n523_0[1]),.doutc(w_n523_0[2]),.din(n523));
	jspl3 jspl3_w_n524_0(.douta(w_n524_0[0]),.doutb(w_n524_0[1]),.doutc(w_n524_0[2]),.din(n524));
	jspl3 jspl3_w_n524_1(.douta(w_n524_1[0]),.doutb(w_n524_1[1]),.doutc(w_dff_A_E8kYfVRo1_2),.din(w_n524_0[0]));
	jspl3 jspl3_w_n526_0(.douta(w_dff_A_powAz74V9_0),.doutb(w_dff_A_6ToQmENd2_1),.doutc(w_n526_0[2]),.din(n526));
	jspl jspl_w_n528_0(.douta(w_n528_0[0]),.doutb(w_n528_0[1]),.din(w_dff_B_O4P7ekHV9_2));
	jspl jspl_w_n530_0(.douta(w_n530_0[0]),.doutb(w_n530_0[1]),.din(n530));
	jspl3 jspl3_w_n531_0(.douta(w_n531_0[0]),.doutb(w_n531_0[1]),.doutc(w_n531_0[2]),.din(n531));
	jspl jspl_w_n531_1(.douta(w_n531_1[0]),.doutb(w_n531_1[1]),.din(w_n531_0[0]));
	jspl3 jspl3_w_n536_0(.douta(w_n536_0[0]),.doutb(w_dff_A_dLMjmZVF5_1),.doutc(w_dff_A_TgcstwJn7_2),.din(n536));
	jspl jspl_w_n538_0(.douta(w_n538_0[0]),.doutb(w_n538_0[1]),.din(n538));
	jspl3 jspl3_w_n539_0(.douta(w_n539_0[0]),.doutb(w_n539_0[1]),.doutc(w_n539_0[2]),.din(n539));
	jspl jspl_w_n539_1(.douta(w_n539_1[0]),.doutb(w_n539_1[1]),.din(w_n539_0[0]));
	jspl jspl_w_n544_0(.douta(w_n544_0[0]),.doutb(w_n544_0[1]),.din(w_dff_B_ihvAxHVv3_2));
	jspl jspl_w_n546_0(.douta(w_n546_0[0]),.doutb(w_n546_0[1]),.din(n546));
	jspl3 jspl3_w_n547_0(.douta(w_n547_0[0]),.doutb(w_n547_0[1]),.doutc(w_n547_0[2]),.din(n547));
	jspl jspl_w_n547_1(.douta(w_n547_1[0]),.doutb(w_n547_1[1]),.din(w_n547_0[0]));
	jspl jspl_w_n548_0(.douta(w_n548_0[0]),.doutb(w_dff_A_VK935xeR7_1),.din(n548));
	jspl jspl_w_n550_0(.douta(w_dff_A_KhFQ59lS2_0),.doutb(w_n550_0[1]),.din(n550));
	jspl jspl_w_n552_0(.douta(w_n552_0[0]),.doutb(w_n552_0[1]),.din(w_dff_B_BCtcMeMM9_2));
	jspl jspl_w_n554_0(.douta(w_n554_0[0]),.doutb(w_n554_0[1]),.din(n554));
	jspl3 jspl3_w_n555_0(.douta(w_n555_0[0]),.doutb(w_n555_0[1]),.doutc(w_n555_0[2]),.din(n555));
	jspl jspl_w_n555_1(.douta(w_n555_1[0]),.doutb(w_n555_1[1]),.din(w_n555_0[0]));
	jspl3 jspl3_w_n556_0(.douta(w_n556_0[0]),.doutb(w_dff_A_wYCagy7e1_1),.doutc(w_dff_A_JTbuxVf88_2),.din(n556));
	jspl jspl_w_n558_0(.douta(w_dff_A_QLaHShLO6_0),.doutb(w_n558_0[1]),.din(n558));
	jspl jspl_w_n560_0(.douta(w_n560_0[0]),.doutb(w_n560_0[1]),.din(w_dff_B_7TqLiHyu6_2));
	jspl jspl_w_n562_0(.douta(w_n562_0[0]),.doutb(w_n562_0[1]),.din(n562));
	jspl3 jspl3_w_n563_0(.douta(w_n563_0[0]),.doutb(w_n563_0[1]),.doutc(w_n563_0[2]),.din(n563));
	jspl jspl_w_n563_1(.douta(w_n563_1[0]),.doutb(w_n563_1[1]),.din(w_n563_0[0]));
	jspl3 jspl3_w_n564_0(.douta(w_n564_0[0]),.doutb(w_dff_A_9eFk9Aht4_1),.doutc(w_dff_A_8HZhCT4c0_2),.din(n564));
	jspl jspl_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.din(n565));
	jspl3 jspl3_w_n566_0(.douta(w_dff_A_SFSrMxs73_0),.doutb(w_n566_0[1]),.doutc(w_n566_0[2]),.din(n566));
	jspl3 jspl3_w_n568_0(.douta(w_n568_0[0]),.doutb(w_n568_0[1]),.doutc(w_n568_0[2]),.din(n568));
	jspl3 jspl3_w_n570_0(.douta(w_n570_0[0]),.doutb(w_n570_0[1]),.doutc(w_n570_0[2]),.din(n570));
	jspl3 jspl3_w_n570_1(.douta(w_n570_1[0]),.doutb(w_dff_A_vtLg4Pz35_1),.doutc(w_n570_1[2]),.din(w_n570_0[0]));
	jspl3 jspl3_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.doutc(w_n572_0[2]),.din(n572));
	jspl jspl_w_n572_1(.douta(w_n572_1[0]),.doutb(w_dff_A_kxNOyO7N4_1),.din(w_n572_0[0]));
	jspl3 jspl3_w_n573_0(.douta(w_n573_0[0]),.doutb(w_dff_A_MNSi9QRU8_1),.doutc(w_dff_A_tuR61V1o1_2),.din(w_dff_B_8mpWh9QD7_3));
	jspl jspl_w_n573_1(.douta(w_dff_A_LvjM02uI6_0),.doutb(w_n573_1[1]),.din(w_n573_0[0]));
	jspl3 jspl3_w_n574_0(.douta(w_n574_0[0]),.doutb(w_dff_A_ygwklOHH0_1),.doutc(w_n574_0[2]),.din(n574));
	jspl3 jspl3_w_n575_0(.douta(w_n575_0[0]),.doutb(w_n575_0[1]),.doutc(w_dff_A_7r7a95wO4_2),.din(n575));
	jspl jspl_w_n575_1(.douta(w_dff_A_8x3bmntu0_0),.doutb(w_n575_1[1]),.din(w_n575_0[0]));
	jspl3 jspl3_w_n576_0(.douta(w_dff_A_hz18Lgjr9_0),.doutb(w_n576_0[1]),.doutc(w_n576_0[2]),.din(n576));
	jspl jspl_w_n577_0(.douta(w_n577_0[0]),.doutb(w_n577_0[1]),.din(n577));
	jspl3 jspl3_w_n578_0(.douta(w_dff_A_lqffWO2G4_0),.doutb(w_dff_A_0TdKwvQd0_1),.doutc(w_n578_0[2]),.din(n578));
	jspl3 jspl3_w_n580_0(.douta(w_dff_A_l2nWqKwK2_0),.doutb(w_dff_A_mon5JnRv2_1),.doutc(w_n580_0[2]),.din(n580));
	jspl3 jspl3_w_n581_0(.douta(w_dff_A_kU1oxVam1_0),.doutb(w_n581_0[1]),.doutc(w_dff_A_GXXDDDUQ5_2),.din(n581));
	jspl3 jspl3_w_n582_0(.douta(w_dff_A_Tr8DNePw2_0),.doutb(w_n582_0[1]),.doutc(w_dff_A_fwUXfxUZ0_2),.din(n582));
	jspl jspl_w_n584_0(.douta(w_n584_0[0]),.doutb(w_n584_0[1]),.din(n584));
	jspl3 jspl3_w_n585_0(.douta(w_n585_0[0]),.doutb(w_n585_0[1]),.doutc(w_n585_0[2]),.din(n585));
	jspl jspl_w_n585_1(.douta(w_n585_1[0]),.doutb(w_n585_1[1]),.din(w_n585_0[0]));
	jspl3 jspl3_w_n586_0(.douta(w_n586_0[0]),.doutb(w_dff_A_2tPgZb2z2_1),.doutc(w_dff_A_WKfWzS9X7_2),.din(n586));
	jspl jspl_w_n588_0(.douta(w_dff_A_RjDBOhul3_0),.doutb(w_n588_0[1]),.din(n588));
	jspl3 jspl3_w_n590_0(.douta(w_n590_0[0]),.doutb(w_dff_A_ekkaAfHZ3_1),.doutc(w_dff_A_LqdujMuD7_2),.din(n590));
	jspl jspl_w_n592_0(.douta(w_n592_0[0]),.doutb(w_n592_0[1]),.din(n592));
	jspl3 jspl3_w_n593_0(.douta(w_n593_0[0]),.doutb(w_n593_0[1]),.doutc(w_n593_0[2]),.din(n593));
	jspl jspl_w_n593_1(.douta(w_n593_1[0]),.doutb(w_n593_1[1]),.din(w_n593_0[0]));
	jspl3 jspl3_w_n594_0(.douta(w_n594_0[0]),.doutb(w_dff_A_hJkd0q0H7_1),.doutc(w_dff_A_uLJhR1De9_2),.din(n594));
	jspl3 jspl3_w_n595_0(.douta(w_n595_0[0]),.doutb(w_dff_A_JBmjHym93_1),.doutc(w_dff_A_lw13vdjv0_2),.din(n595));
	jspl jspl_w_n597_0(.douta(w_n597_0[0]),.doutb(w_n597_0[1]),.din(n597));
	jspl3 jspl3_w_n598_0(.douta(w_n598_0[0]),.doutb(w_n598_0[1]),.doutc(w_n598_0[2]),.din(n598));
	jspl jspl_w_n598_1(.douta(w_n598_1[0]),.doutb(w_n598_1[1]),.din(w_n598_0[0]));
	jspl3 jspl3_w_n599_0(.douta(w_n599_0[0]),.doutb(w_n599_0[1]),.doutc(w_n599_0[2]),.din(n599));
	jspl jspl_w_n600_0(.douta(w_n600_0[0]),.doutb(w_n600_0[1]),.din(w_dff_B_TNGCVpEa1_2));
	jspl jspl_w_n602_0(.douta(w_n602_0[0]),.doutb(w_n602_0[1]),.din(n602));
	jspl3 jspl3_w_n603_0(.douta(w_n603_0[0]),.doutb(w_n603_0[1]),.doutc(w_n603_0[2]),.din(n603));
	jspl jspl_w_n603_1(.douta(w_n603_1[0]),.doutb(w_n603_1[1]),.din(w_n603_0[0]));
	jspl jspl_w_n604_0(.douta(w_dff_A_fpwKEp9r3_0),.doutb(w_n604_0[1]),.din(n604));
	jspl3 jspl3_w_n605_0(.douta(w_dff_A_VLtttGbJ4_0),.doutb(w_dff_A_lUsHpICq5_1),.doutc(w_n605_0[2]),.din(n605));
	jspl jspl_w_n609_0(.douta(w_n609_0[0]),.doutb(w_dff_A_f82UZDuO2_1),.din(w_dff_B_n6OpHj769_2));
	jspl jspl_w_n610_0(.douta(w_dff_A_oEs2wZ5J3_0),.doutb(w_n610_0[1]),.din(n610));
	jspl jspl_w_n612_0(.douta(w_n612_0[0]),.doutb(w_dff_A_wLnESNMi5_1),.din(n612));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.doutc(w_n613_0[2]),.din(n613));
	jspl3 jspl3_w_n615_0(.douta(w_n615_0[0]),.doutb(w_dff_A_QJDwRvtH6_1),.doutc(w_n615_0[2]),.din(n615));
	jspl jspl_w_n616_0(.douta(w_n616_0[0]),.doutb(w_n616_0[1]),.din(n616));
	jspl3 jspl3_w_n618_0(.douta(w_dff_A_Kz2uNPy41_0),.doutb(w_n618_0[1]),.doutc(w_n618_0[2]),.din(n618));
	jspl3 jspl3_w_n619_0(.douta(w_n619_0[0]),.doutb(w_dff_A_nT099fAz5_1),.doutc(w_n619_0[2]),.din(n619));
	jspl3 jspl3_w_n622_0(.douta(w_n622_0[0]),.doutb(w_dff_A_6JY6j7Qz2_1),.doutc(w_dff_A_f2nqb3SF5_2),.din(n622));
	jspl jspl_w_n624_0(.douta(w_n624_0[0]),.doutb(w_n624_0[1]),.din(n624));
	jspl3 jspl3_w_n625_0(.douta(w_n625_0[0]),.doutb(w_n625_0[1]),.doutc(w_n625_0[2]),.din(n625));
	jspl jspl_w_n625_1(.douta(w_n625_1[0]),.doutb(w_n625_1[1]),.din(w_n625_0[0]));
	jspl3 jspl3_w_n626_0(.douta(w_dff_A_lEWmyDbc0_0),.doutb(w_dff_A_ZNiXlFuF1_1),.doutc(w_n626_0[2]),.din(n626));
	jspl jspl_w_n626_1(.douta(w_dff_A_RoLXqBJa7_0),.doutb(w_n626_1[1]),.din(w_n626_0[0]));
	jspl3 jspl3_w_n627_0(.douta(w_n627_0[0]),.doutb(w_dff_A_3QSoSmmK1_1),.doutc(w_dff_A_MQZwyx2v6_2),.din(n627));
	jspl jspl_w_n629_0(.douta(w_n629_0[0]),.doutb(w_n629_0[1]),.din(n629));
	jspl3 jspl3_w_n630_0(.douta(w_n630_0[0]),.doutb(w_n630_0[1]),.doutc(w_n630_0[2]),.din(n630));
	jspl3 jspl3_w_n631_0(.douta(w_n631_0[0]),.doutb(w_dff_A_WZmF5jrl7_1),.doutc(w_dff_A_LKOjZSAq4_2),.din(n631));
	jspl3 jspl3_w_n632_0(.douta(w_dff_A_xecZ0YzB1_0),.doutb(w_n632_0[1]),.doutc(w_dff_A_XWBOdunm4_2),.din(n632));
	jspl jspl_w_n632_1(.douta(w_n632_1[0]),.doutb(w_n632_1[1]),.din(w_n632_0[0]));
	jspl jspl_w_n634_0(.douta(w_n634_0[0]),.doutb(w_n634_0[1]),.din(n634));
	jspl3 jspl3_w_n635_0(.douta(w_n635_0[0]),.doutb(w_n635_0[1]),.doutc(w_n635_0[2]),.din(n635));
	jspl jspl_w_n635_1(.douta(w_n635_1[0]),.doutb(w_n635_1[1]),.din(w_n635_0[0]));
	jspl3 jspl3_w_n636_0(.douta(w_n636_0[0]),.doutb(w_dff_A_fMw4awqK4_1),.doutc(w_dff_A_qhiPFY6g6_2),.din(n636));
	jspl3 jspl3_w_n641_0(.douta(w_n641_0[0]),.doutb(w_n641_0[1]),.doutc(w_n641_0[2]),.din(n641));
	jspl3 jspl3_w_n642_0(.douta(w_n642_0[0]),.doutb(w_dff_A_rNwQE5Az1_1),.doutc(w_n642_0[2]),.din(w_dff_B_iivay0ji0_3));
	jspl jspl_w_n644_0(.douta(w_n644_0[0]),.doutb(w_n644_0[1]),.din(n644));
	jspl jspl_w_n645_0(.douta(w_n645_0[0]),.doutb(w_n645_0[1]),.din(n645));
	jspl jspl_w_n646_0(.douta(w_n646_0[0]),.doutb(w_dff_A_G23F854o3_1),.din(n646));
	jspl jspl_w_n647_0(.douta(w_n647_0[0]),.doutb(w_dff_A_u7CR8iOw3_1),.din(n647));
	jspl jspl_w_n649_0(.douta(w_dff_A_CQBBE4km1_0),.doutb(w_n649_0[1]),.din(n649));
	jspl jspl_w_n651_0(.douta(w_n651_0[0]),.doutb(w_n651_0[1]),.din(n651));
	jspl jspl_w_n652_0(.douta(w_dff_A_QcjPCR3s1_0),.doutb(w_n652_0[1]),.din(n652));
	jspl jspl_w_n653_0(.douta(w_dff_A_lZXB9Ylo4_0),.doutb(w_n653_0[1]),.din(w_dff_B_kKtfS4rA8_2));
	jspl3 jspl3_w_n654_0(.douta(w_n654_0[0]),.doutb(w_dff_A_uPsZQYsd5_1),.doutc(w_dff_A_RzDvUsnI8_2),.din(n654));
	jspl jspl_w_n655_0(.douta(w_n655_0[0]),.doutb(w_dff_A_pjFj03hC5_1),.din(n655));
	jspl jspl_w_n656_0(.douta(w_n656_0[0]),.doutb(w_dff_A_We4CQKko3_1),.din(n656));
	jspl3 jspl3_w_n657_0(.douta(w_n657_0[0]),.doutb(w_dff_A_T6DH3wwq8_1),.doutc(w_dff_A_mb2OTymV4_2),.din(n657));
	jspl jspl_w_n659_0(.douta(w_n659_0[0]),.doutb(w_n659_0[1]),.din(n659));
	jspl3 jspl3_w_n660_0(.douta(w_n660_0[0]),.doutb(w_n660_0[1]),.doutc(w_n660_0[2]),.din(n660));
	jspl3 jspl3_w_n661_0(.douta(w_n661_0[0]),.doutb(w_dff_A_fUruxAvU7_1),.doutc(w_dff_A_lqYBdj6U0_2),.din(n661));
	jspl jspl_w_n662_0(.douta(w_n662_0[0]),.doutb(w_dff_A_g3iSUOi77_1),.din(n662));
	jspl3 jspl3_w_n663_0(.douta(w_n663_0[0]),.doutb(w_n663_0[1]),.doutc(w_n663_0[2]),.din(n663));
	jspl jspl_w_n663_1(.douta(w_n663_1[0]),.doutb(w_n663_1[1]),.din(w_n663_0[0]));
	jspl jspl_w_n664_0(.douta(w_dff_A_k4tZXlm27_0),.doutb(w_n664_0[1]),.din(w_dff_B_okLIaUll6_2));
	jspl jspl_w_n666_0(.douta(w_dff_A_Bwd6QaoA3_0),.doutb(w_n666_0[1]),.din(n666));
	jspl jspl_w_n669_0(.douta(w_n669_0[0]),.doutb(w_n669_0[1]),.din(n669));
	jspl jspl_w_n671_0(.douta(w_n671_0[0]),.doutb(w_n671_0[1]),.din(n671));
	jspl3 jspl3_w_n673_0(.douta(w_n673_0[0]),.doutb(w_n673_0[1]),.doutc(w_n673_0[2]),.din(n673));
	jspl jspl_w_n674_0(.douta(w_n674_0[0]),.doutb(w_n674_0[1]),.din(n674));
	jspl3 jspl3_w_n676_0(.douta(w_n676_0[0]),.doutb(w_n676_0[1]),.doutc(w_n676_0[2]),.din(n676));
	jspl jspl_w_n678_0(.douta(w_n678_0[0]),.doutb(w_n678_0[1]),.din(n678));
	jspl3 jspl3_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.doutc(w_n680_0[2]),.din(n680));
	jspl3 jspl3_w_n680_1(.douta(w_n680_1[0]),.doutb(w_n680_1[1]),.doutc(w_n680_1[2]),.din(w_n680_0[0]));
	jspl3 jspl3_w_n680_2(.douta(w_n680_2[0]),.doutb(w_n680_2[1]),.doutc(w_n680_2[2]),.din(w_n680_0[1]));
	jspl jspl_w_n682_0(.douta(w_n682_0[0]),.doutb(w_n682_0[1]),.din(n682));
	jspl jspl_w_n683_0(.douta(w_n683_0[0]),.doutb(w_n683_0[1]),.din(n683));
	jspl jspl_w_n687_0(.douta(w_dff_A_EwimlYRb6_0),.doutb(w_n687_0[1]),.din(n687));
	jspl jspl_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.din(n689));
	jspl jspl_w_n690_0(.douta(w_n690_0[0]),.doutb(w_dff_A_cBpxTyuL7_1),.din(w_dff_B_stDaMQtR2_2));
	jspl jspl_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.din(n693));
	jspl jspl_w_n694_0(.douta(w_dff_A_q5tRPNSs9_0),.doutb(w_n694_0[1]),.din(n694));
	jspl jspl_w_n695_0(.douta(w_n695_0[0]),.doutb(w_n695_0[1]),.din(n695));
	jspl jspl_w_n696_0(.douta(w_dff_A_iQeXEwhg6_0),.doutb(w_n696_0[1]),.din(n696));
	jspl jspl_w_n698_0(.douta(w_n698_0[0]),.doutb(w_n698_0[1]),.din(n698));
	jspl3 jspl3_w_n700_0(.douta(w_n700_0[0]),.doutb(w_n700_0[1]),.doutc(w_n700_0[2]),.din(n700));
	jspl jspl_w_n700_1(.douta(w_n700_1[0]),.doutb(w_n700_1[1]),.din(w_n700_0[0]));
	jspl3 jspl3_w_n703_0(.douta(w_n703_0[0]),.doutb(w_n703_0[1]),.doutc(w_n703_0[2]),.din(n703));
	jspl3 jspl3_w_n703_1(.douta(w_n703_1[0]),.doutb(w_n703_1[1]),.doutc(w_n703_1[2]),.din(w_n703_0[0]));
	jspl jspl_w_n705_0(.douta(w_n705_0[0]),.doutb(w_n705_0[1]),.din(n705));
	jspl3 jspl3_w_n707_0(.douta(w_n707_0[0]),.doutb(w_n707_0[1]),.doutc(w_n707_0[2]),.din(n707));
	jspl3 jspl3_w_n707_1(.douta(w_n707_1[0]),.doutb(w_n707_1[1]),.doutc(w_n707_1[2]),.din(w_n707_0[0]));
	jspl3 jspl3_w_n709_0(.douta(w_n709_0[0]),.doutb(w_n709_0[1]),.doutc(w_n709_0[2]),.din(n709));
	jspl jspl_w_n709_1(.douta(w_n709_1[0]),.doutb(w_n709_1[1]),.din(w_n709_0[0]));
	jspl3 jspl3_w_n711_0(.douta(w_n711_0[0]),.doutb(w_n711_0[1]),.doutc(w_n711_0[2]),.din(n711));
	jspl jspl_w_n711_1(.douta(w_n711_1[0]),.doutb(w_n711_1[1]),.din(w_n711_0[0]));
	jspl3 jspl3_w_n712_0(.douta(w_n712_0[0]),.doutb(w_n712_0[1]),.doutc(w_n712_0[2]),.din(n712));
	jspl jspl_w_n713_0(.douta(w_dff_A_Nq8HOIKa7_0),.doutb(w_n713_0[1]),.din(n713));
	jspl3 jspl3_w_n715_0(.douta(w_n715_0[0]),.doutb(w_n715_0[1]),.doutc(w_n715_0[2]),.din(w_dff_B_szjUyLJN5_3));
	jspl jspl_w_n715_1(.douta(w_n715_1[0]),.doutb(w_n715_1[1]),.din(w_n715_0[0]));
	jspl3 jspl3_w_n718_0(.douta(w_n718_0[0]),.doutb(w_n718_0[1]),.doutc(w_n718_0[2]),.din(w_dff_B_KT5fBCnk8_3));
	jspl jspl_w_n719_0(.douta(w_dff_A_3E42TCUS7_0),.doutb(w_n719_0[1]),.din(n719));
	jspl3 jspl3_w_n720_0(.douta(w_n720_0[0]),.doutb(w_n720_0[1]),.doutc(w_n720_0[2]),.din(n720));
	jspl3 jspl3_w_n723_0(.douta(w_n723_0[0]),.doutb(w_n723_0[1]),.doutc(w_n723_0[2]),.din(n723));
	jspl jspl_w_n724_0(.douta(w_n724_0[0]),.doutb(w_dff_A_M57ltLga8_1),.din(n724));
	jspl jspl_w_n725_0(.douta(w_dff_A_IBrD16ts4_0),.doutb(w_n725_0[1]),.din(n725));
	jspl3 jspl3_w_n726_0(.douta(w_n726_0[0]),.doutb(w_n726_0[1]),.doutc(w_n726_0[2]),.din(n726));
	jspl jspl_w_n726_1(.douta(w_n726_1[0]),.doutb(w_n726_1[1]),.din(w_n726_0[0]));
	jspl3 jspl3_w_n729_0(.douta(w_n729_0[0]),.doutb(w_n729_0[1]),.doutc(w_n729_0[2]),.din(n729));
	jspl jspl_w_n729_1(.douta(w_n729_1[0]),.doutb(w_n729_1[1]),.din(w_n729_0[0]));
	jspl3 jspl3_w_n734_0(.douta(w_n734_0[0]),.doutb(w_n734_0[1]),.doutc(w_n734_0[2]),.din(n734));
	jspl jspl_w_n736_0(.douta(w_n736_0[0]),.doutb(w_n736_0[1]),.din(n736));
	jspl3 jspl3_w_n737_0(.douta(w_n737_0[0]),.doutb(w_n737_0[1]),.doutc(w_n737_0[2]),.din(n737));
	jspl jspl_w_n737_1(.douta(w_n737_1[0]),.doutb(w_n737_1[1]),.din(w_n737_0[0]));
	jspl3 jspl3_w_n741_0(.douta(w_n741_0[0]),.doutb(w_n741_0[1]),.doutc(w_n741_0[2]),.din(n741));
	jspl jspl_w_n741_1(.douta(w_n741_1[0]),.doutb(w_n741_1[1]),.din(w_n741_0[0]));
	jspl jspl_w_n743_0(.douta(w_n743_0[0]),.doutb(w_n743_0[1]),.din(n743));
	jspl3 jspl3_w_n744_0(.douta(w_n744_0[0]),.doutb(w_n744_0[1]),.doutc(w_n744_0[2]),.din(n744));
	jspl3 jspl3_w_n747_0(.douta(w_n747_0[0]),.doutb(w_n747_0[1]),.doutc(w_n747_0[2]),.din(n747));
	jspl jspl_w_n749_0(.douta(w_n749_0[0]),.doutb(w_n749_0[1]),.din(n749));
	jspl jspl_w_n754_0(.douta(w_n754_0[0]),.doutb(w_n754_0[1]),.din(n754));
	jspl3 jspl3_w_n755_0(.douta(w_n755_0[0]),.doutb(w_n755_0[1]),.doutc(w_n755_0[2]),.din(n755));
	jspl jspl_w_n755_1(.douta(w_n755_1[0]),.doutb(w_n755_1[1]),.din(w_n755_0[0]));
	jspl3 jspl3_w_n758_0(.douta(w_n758_0[0]),.doutb(w_n758_0[1]),.doutc(w_n758_0[2]),.din(n758));
	jspl jspl_w_n758_1(.douta(w_n758_1[0]),.doutb(w_n758_1[1]),.din(w_n758_0[0]));
	jspl jspl_w_n760_0(.douta(w_n760_0[0]),.doutb(w_n760_0[1]),.din(n760));
	jspl3 jspl3_w_n761_0(.douta(w_n761_0[0]),.doutb(w_n761_0[1]),.doutc(w_n761_0[2]),.din(n761));
	jspl3 jspl3_w_n764_0(.douta(w_n764_0[0]),.doutb(w_n764_0[1]),.doutc(w_n764_0[2]),.din(n764));
	jspl jspl_w_n766_0(.douta(w_n766_0[0]),.doutb(w_n766_0[1]),.din(w_dff_B_E8nBb3DH5_2));
	jspl jspl_w_n767_0(.douta(w_n767_0[0]),.doutb(w_n767_0[1]),.din(n767));
	jspl3 jspl3_w_n768_0(.douta(w_n768_0[0]),.doutb(w_n768_0[1]),.doutc(w_n768_0[2]),.din(n768));
	jspl3 jspl3_w_n772_0(.douta(w_n772_0[0]),.doutb(w_n772_0[1]),.doutc(w_n772_0[2]),.din(n772));
	jspl jspl_w_n773_0(.douta(w_n773_0[0]),.doutb(w_dff_A_enWUTCuu1_1),.din(n773));
	jspl jspl_w_n774_0(.douta(w_n774_0[0]),.doutb(w_n774_0[1]),.din(n774));
	jspl jspl_w_n775_0(.douta(w_n775_0[0]),.doutb(w_n775_0[1]),.din(n775));
	jspl3 jspl3_w_n776_0(.douta(w_n776_0[0]),.doutb(w_n776_0[1]),.doutc(w_n776_0[2]),.din(n776));
	jspl3 jspl3_w_n780_0(.douta(w_dff_A_8zHwxbIv2_0),.doutb(w_n780_0[1]),.doutc(w_n780_0[2]),.din(n780));
	jspl jspl_w_n781_0(.douta(w_n781_0[0]),.doutb(w_n781_0[1]),.din(n781));
	jspl3 jspl3_w_n796_0(.douta(w_n796_0[0]),.doutb(w_n796_0[1]),.doutc(w_n796_0[2]),.din(n796));
	jspl jspl_w_n796_1(.douta(w_n796_1[0]),.doutb(w_n796_1[1]),.din(w_n796_0[0]));
	jspl3 jspl3_w_n800_0(.douta(w_n800_0[0]),.doutb(w_n800_0[1]),.doutc(w_n800_0[2]),.din(n800));
	jspl jspl_w_n800_1(.douta(w_n800_1[0]),.doutb(w_n800_1[1]),.din(w_n800_0[0]));
	jspl3 jspl3_w_n803_0(.douta(w_n803_0[0]),.doutb(w_n803_0[1]),.doutc(w_n803_0[2]),.din(n803));
	jspl3 jspl3_w_n806_0(.douta(w_n806_0[0]),.doutb(w_n806_0[1]),.doutc(w_n806_0[2]),.din(n806));
	jspl jspl_w_n808_0(.douta(w_n808_0[0]),.doutb(w_dff_A_KeH7Nrrb3_1),.din(n808));
	jspl3 jspl3_w_n810_0(.douta(w_n810_0[0]),.doutb(w_n810_0[1]),.doutc(w_n810_0[2]),.din(n810));
	jspl jspl_w_n810_1(.douta(w_n810_1[0]),.doutb(w_n810_1[1]),.din(w_n810_0[0]));
	jspl3 jspl3_w_n814_0(.douta(w_n814_0[0]),.doutb(w_n814_0[1]),.doutc(w_n814_0[2]),.din(n814));
	jspl jspl_w_n814_1(.douta(w_n814_1[0]),.doutb(w_n814_1[1]),.din(w_n814_0[0]));
	jspl3 jspl3_w_n817_0(.douta(w_n817_0[0]),.doutb(w_n817_0[1]),.doutc(w_n817_0[2]),.din(n817));
	jspl3 jspl3_w_n820_0(.douta(w_n820_0[0]),.doutb(w_n820_0[1]),.doutc(w_n820_0[2]),.din(n820));
	jspl jspl_w_n822_0(.douta(w_n822_0[0]),.doutb(w_n822_0[1]),.din(n822));
	jspl3 jspl3_w_n824_0(.douta(w_n824_0[0]),.doutb(w_n824_0[1]),.doutc(w_n824_0[2]),.din(n824));
	jspl3 jspl3_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.doutc(w_n827_0[2]),.din(n827));
	jspl3 jspl3_w_n845_0(.douta(w_n845_0[0]),.doutb(w_dff_A_zDNHOQQv8_1),.doutc(w_n845_0[2]),.din(n845));
	jspl jspl_w_n845_1(.douta(w_n845_1[0]),.doutb(w_n845_1[1]),.din(w_n845_0[0]));
	jspl3 jspl3_w_n848_0(.douta(w_n848_0[0]),.doutb(w_n848_0[1]),.doutc(w_n848_0[2]),.din(n848));
	jspl jspl_w_n848_1(.douta(w_n848_1[0]),.doutb(w_n848_1[1]),.din(w_n848_0[0]));
	jspl3 jspl3_w_n851_0(.douta(w_n851_0[0]),.doutb(w_n851_0[1]),.doutc(w_n851_0[2]),.din(n851));
	jspl3 jspl3_w_n854_0(.douta(w_n854_0[0]),.doutb(w_n854_0[1]),.doutc(w_n854_0[2]),.din(n854));
	jspl jspl_w_n856_0(.douta(w_n856_0[0]),.doutb(w_dff_A_AEaRPL7B0_1),.din(n856));
	jspl3 jspl3_w_n858_0(.douta(w_n858_0[0]),.doutb(w_n858_0[1]),.doutc(w_n858_0[2]),.din(n858));
	jspl3 jspl3_w_n862_0(.douta(w_n862_0[0]),.doutb(w_n862_0[1]),.doutc(w_n862_0[2]),.din(n862));
	jspl jspl_w_n863_0(.douta(w_n863_0[0]),.doutb(w_dff_A_G2KgPMH80_1),.din(n863));
	jspl jspl_w_n864_0(.douta(w_n864_0[0]),.doutb(w_n864_0[1]),.din(n864));
	jspl3 jspl3_w_n866_0(.douta(w_n866_0[0]),.doutb(w_n866_0[1]),.doutc(w_n866_0[2]),.din(n866));
	jspl3 jspl3_w_n870_0(.douta(w_n870_0[0]),.doutb(w_n870_0[1]),.doutc(w_n870_0[2]),.din(n870));
	jspl jspl_w_n871_0(.douta(w_n871_0[0]),.doutb(w_n871_0[1]),.din(n871));
	jspl3 jspl3_w_n885_0(.douta(w_n885_0[0]),.doutb(w_n885_0[1]),.doutc(w_n885_0[2]),.din(n885));
	jspl3 jspl3_w_n888_0(.douta(w_n888_0[0]),.doutb(w_n888_0[1]),.doutc(w_n888_0[2]),.din(n888));
	jspl3 jspl3_w_n891_0(.douta(w_n891_0[0]),.doutb(w_n891_0[1]),.doutc(w_n891_0[2]),.din(n891));
	jspl3 jspl3_w_n894_0(.douta(w_n894_0[0]),.doutb(w_n894_0[1]),.doutc(w_n894_0[2]),.din(n894));
	jspl jspl_w_n895_0(.douta(w_dff_A_RAnhR2Ke5_0),.doutb(w_n895_0[1]),.din(n895));
	jspl3 jspl3_w_n900_0(.douta(w_n900_0[0]),.doutb(w_n900_0[1]),.doutc(w_n900_0[2]),.din(n900));
	jspl3 jspl3_w_n903_0(.douta(w_n903_0[0]),.doutb(w_n903_0[1]),.doutc(w_n903_0[2]),.din(n903));
	jspl jspl_w_n905_0(.douta(w_dff_A_WiualOEz8_0),.doutb(w_n905_0[1]),.din(n905));
	jspl3 jspl3_w_n916_0(.douta(w_n916_0[0]),.doutb(w_n916_0[1]),.doutc(w_n916_0[2]),.din(n916));
	jspl3 jspl3_w_n919_0(.douta(w_n919_0[0]),.doutb(w_n919_0[1]),.doutc(w_n919_0[2]),.din(n919));
	jspl3 jspl3_w_n926_0(.douta(w_dff_A_DLyspXo41_0),.doutb(w_n926_0[1]),.doutc(w_n926_0[2]),.din(n926));
	jspl3 jspl3_w_n930_0(.douta(w_n930_0[0]),.doutb(w_n930_0[1]),.doutc(w_n930_0[2]),.din(n930));
	jspl3 jspl3_w_n935_0(.douta(w_n935_0[0]),.doutb(w_n935_0[1]),.doutc(w_n935_0[2]),.din(n935));
	jspl3 jspl3_w_n938_0(.douta(w_dff_A_6CCpYkzY5_0),.doutb(w_n938_0[1]),.doutc(w_n938_0[2]),.din(n938));
	jspl3 jspl3_w_n944_0(.douta(w_n944_0[0]),.doutb(w_n944_0[1]),.doutc(w_n944_0[2]),.din(n944));
	jspl3 jspl3_w_n947_0(.douta(w_n947_0[0]),.doutb(w_n947_0[1]),.doutc(w_n947_0[2]),.din(n947));
	jspl3 jspl3_w_n950_0(.douta(w_n950_0[0]),.doutb(w_n950_0[1]),.doutc(w_n950_0[2]),.din(n950));
	jspl jspl_w_n950_1(.douta(w_n950_1[0]),.doutb(w_n950_1[1]),.din(w_n950_0[0]));
	jspl3 jspl3_w_n953_0(.douta(w_n953_0[0]),.doutb(w_n953_0[1]),.doutc(w_n953_0[2]),.din(n953));
	jspl jspl_w_n953_1(.douta(w_n953_1[0]),.doutb(w_n953_1[1]),.din(w_n953_0[0]));
	jspl3 jspl3_w_n966_0(.douta(w_n966_0[0]),.doutb(w_n966_0[1]),.doutc(w_n966_0[2]),.din(n966));
	jspl3 jspl3_w_n970_0(.douta(w_n970_0[0]),.doutb(w_n970_0[1]),.doutc(w_n970_0[2]),.din(n970));
	jspl3 jspl3_w_n973_0(.douta(w_n973_0[0]),.doutb(w_n973_0[1]),.doutc(w_n973_0[2]),.din(n973));
	jspl jspl_w_n973_1(.douta(w_n973_1[0]),.doutb(w_n973_1[1]),.din(w_n973_0[0]));
	jspl3 jspl3_w_n977_0(.douta(w_n977_0[0]),.doutb(w_n977_0[1]),.doutc(w_n977_0[2]),.din(n977));
	jspl jspl_w_n977_1(.douta(w_n977_1[0]),.doutb(w_n977_1[1]),.din(w_n977_0[0]));
	jspl3 jspl3_w_n980_0(.douta(w_n980_0[0]),.doutb(w_n980_0[1]),.doutc(w_n980_0[2]),.din(n980));
	jspl3 jspl3_w_n983_0(.douta(w_n983_0[0]),.doutb(w_n983_0[1]),.doutc(w_n983_0[2]),.din(n983));
	jspl jspl_w_n985_0(.douta(w_n985_0[0]),.doutb(w_dff_A_lzsf9YNj2_1),.din(w_dff_B_Xus4ekrH4_2));
	jspl3 jspl3_w_n987_0(.douta(w_n987_0[0]),.doutb(w_n987_0[1]),.doutc(w_n987_0[2]),.din(n987));
	jspl3 jspl3_w_n991_0(.douta(w_n991_0[0]),.doutb(w_n991_0[1]),.doutc(w_n991_0[2]),.din(n991));
	jspl jspl_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.din(n992));
	jspl3 jspl3_w_n995_0(.douta(w_n995_0[0]),.doutb(w_n995_0[1]),.doutc(w_n995_0[2]),.din(n995));
	jspl3 jspl3_w_n999_0(.douta(w_n999_0[0]),.doutb(w_n999_0[1]),.doutc(w_n999_0[2]),.din(n999));
	jspl jspl_w_n1000_0(.douta(w_n1000_0[0]),.doutb(w_dff_A_Tss7Uoax4_1),.din(n1000));
	jspl jspl_w_n1003_0(.douta(w_dff_A_c6ksV2It6_0),.doutb(w_n1003_0[1]),.din(n1003));
	jspl jspl_w_n1007_0(.douta(w_n1007_0[0]),.doutb(w_n1007_0[1]),.din(n1007));
	jspl jspl_w_n1008_0(.douta(w_dff_A_XqgRxEJy4_0),.doutb(w_n1008_0[1]),.din(n1008));
	jspl jspl_w_n1042_0(.douta(w_dff_A_CphRJuGg1_0),.doutb(w_n1042_0[1]),.din(n1042));
	jspl3 jspl3_w_n1059_0(.douta(w_n1059_0[0]),.doutb(w_n1059_0[1]),.doutc(w_n1059_0[2]),.din(n1059));
	jspl3 jspl3_w_n1067_0(.douta(w_n1067_0[0]),.doutb(w_n1067_0[1]),.doutc(w_n1067_0[2]),.din(n1067));
	jspl3 jspl3_w_n1069_0(.douta(w_n1069_0[0]),.doutb(w_n1069_0[1]),.doutc(w_n1069_0[2]),.din(n1069));
	jspl jspl_w_n1070_0(.douta(w_n1070_0[0]),.doutb(w_n1070_0[1]),.din(n1070));
	jspl jspl_w_n1073_0(.douta(w_n1073_0[0]),.doutb(w_n1073_0[1]),.din(n1073));
	jspl jspl_w_n1078_0(.douta(w_n1078_0[0]),.doutb(w_n1078_0[1]),.din(n1078));
	jspl3 jspl3_w_n1084_0(.douta(w_n1084_0[0]),.doutb(w_dff_A_T2l5DZtf0_1),.doutc(w_dff_A_9nPoXgzs7_2),.din(n1084));
	jspl jspl_w_n1086_0(.douta(w_dff_A_HwbULfST9_0),.doutb(w_n1086_0[1]),.din(w_dff_B_IL6LlgCz6_2));
	jspl jspl_w_n1090_0(.douta(w_n1090_0[0]),.doutb(w_n1090_0[1]),.din(n1090));
	jspl3 jspl3_w_n1092_0(.douta(w_n1092_0[0]),.doutb(w_n1092_0[1]),.doutc(w_n1092_0[2]),.din(n1092));
	jspl3 jspl3_w_n1094_0(.douta(w_dff_A_jX290eNI2_0),.doutb(w_dff_A_SxvGIu5g6_1),.doutc(w_n1094_0[2]),.din(w_dff_B_ldnKndYB2_3));
	jspl jspl_w_n1096_0(.douta(w_n1096_0[0]),.doutb(w_n1096_0[1]),.din(n1096));
	jspl jspl_w_n1099_0(.douta(w_n1099_0[0]),.doutb(w_n1099_0[1]),.din(n1099));
	jspl jspl_w_n1105_0(.douta(w_n1105_0[0]),.doutb(w_dff_A_0FiDF4Wn0_1),.din(w_dff_B_50ilp20S7_2));
	jspl jspl_w_n1106_0(.douta(w_n1106_0[0]),.doutb(w_dff_A_7QPIrrcj9_1),.din(n1106));
	jspl jspl_w_n1108_0(.douta(w_n1108_0[0]),.doutb(w_dff_A_dju4lfQv3_1),.din(n1108));
	jspl jspl_w_n1113_0(.douta(w_n1113_0[0]),.doutb(w_n1113_0[1]),.din(n1113));
	jspl jspl_w_n1118_0(.douta(w_n1118_0[0]),.doutb(w_n1118_0[1]),.din(n1118));
	jspl jspl_w_n1127_0(.douta(w_n1127_0[0]),.doutb(w_n1127_0[1]),.din(n1127));
	jspl jspl_w_n1137_0(.douta(w_n1137_0[0]),.doutb(w_n1137_0[1]),.din(n1137));
	jspl jspl_w_n1150_0(.douta(w_n1150_0[0]),.doutb(w_n1150_0[1]),.din(n1150));
	jspl jspl_w_n1172_0(.douta(w_n1172_0[0]),.doutb(w_n1172_0[1]),.din(n1172));
	jspl jspl_w_n1307_0(.douta(w_dff_A_5PzhnG0g9_0),.doutb(w_n1307_0[1]),.din(w_dff_B_YG7X9TBI8_2));
	jspl jspl_w_n1308_0(.douta(w_n1308_0[0]),.doutb(w_dff_A_zlS3VSDO0_1),.din(n1308));
	jspl jspl_w_n1309_0(.douta(w_n1309_0[0]),.doutb(w_dff_A_HnVWsxJd4_1),.din(n1309));
	jspl jspl_w_n1310_0(.douta(w_n1310_0[0]),.doutb(w_dff_A_7hPF4fB09_1),.din(w_dff_B_cMRHQBCL1_2));
	jspl3 jspl3_w_n1312_0(.douta(w_n1312_0[0]),.doutb(w_n1312_0[1]),.doutc(w_n1312_0[2]),.din(n1312));
	jspl jspl_w_n1312_1(.douta(w_n1312_1[0]),.doutb(w_n1312_1[1]),.din(w_n1312_0[0]));
	jspl jspl_w_n1316_0(.douta(w_n1316_0[0]),.doutb(w_n1316_0[1]),.din(n1316));
	jspl jspl_w_n1317_0(.douta(w_n1317_0[0]),.doutb(w_n1317_0[1]),.din(n1317));
	jspl3 jspl3_w_n1321_0(.douta(w_n1321_0[0]),.doutb(w_n1321_0[1]),.doutc(w_n1321_0[2]),.din(n1321));
	jspl jspl_w_n1321_1(.douta(w_n1321_1[0]),.doutb(w_n1321_1[1]),.din(w_n1321_0[0]));
	jspl jspl_w_n1323_0(.douta(w_n1323_0[0]),.doutb(w_n1323_0[1]),.din(w_dff_B_Q4fjijCy2_2));
	jspl jspl_w_n1333_0(.douta(w_n1333_0[0]),.doutb(w_n1333_0[1]),.din(n1333));
	jspl3 jspl3_w_n1337_0(.douta(w_n1337_0[0]),.doutb(w_n1337_0[1]),.doutc(w_n1337_0[2]),.din(n1337));
	jspl jspl_w_n1337_1(.douta(w_n1337_1[0]),.doutb(w_n1337_1[1]),.din(w_n1337_0[0]));
	jspl3 jspl3_w_n1340_0(.douta(w_n1340_0[0]),.doutb(w_dff_A_AKv7wvjL7_1),.doutc(w_dff_A_uDXqbVQo7_2),.din(w_dff_B_h8YYfvGs6_3));
	jspl jspl_w_n1343_0(.douta(w_n1343_0[0]),.doutb(w_n1343_0[1]),.din(n1343));
	jspl jspl_w_n1344_0(.douta(w_n1344_0[0]),.doutb(w_n1344_0[1]),.din(n1344));
	jspl jspl_w_n1359_0(.douta(w_n1359_0[0]),.doutb(w_dff_A_TWZkus282_1),.din(w_dff_B_a3SJFK7E1_2));
	jspl jspl_w_n1364_0(.douta(w_n1364_0[0]),.doutb(w_dff_A_WB2CvrJW5_1),.din(n1364));
	jspl jspl_w_n1369_0(.douta(w_n1369_0[0]),.doutb(w_n1369_0[1]),.din(w_dff_B_EqhbmTAQ8_2));
	jspl jspl_w_n1370_0(.douta(w_n1370_0[0]),.doutb(w_dff_A_BCmgUvh55_1),.din(w_dff_B_5rJKp6IJ3_2));
	jspl jspl_w_n1372_0(.douta(w_n1372_0[0]),.doutb(w_n1372_0[1]),.din(n1372));
	jspl jspl_w_n1387_0(.douta(w_dff_A_1wkanVuV3_0),.doutb(w_n1387_0[1]),.din(n1387));
	jspl jspl_w_n1388_0(.douta(w_n1388_0[0]),.doutb(w_dff_A_3hTYa1n72_1),.din(n1388));
	jspl jspl_w_n1396_0(.douta(w_n1396_0[0]),.doutb(w_n1396_0[1]),.din(n1396));
	jspl jspl_w_n1402_0(.douta(w_n1402_0[0]),.doutb(w_dff_A_GpqMXNZU8_1),.din(n1402));
	jspl jspl_w_n1408_0(.douta(w_n1408_0[0]),.doutb(w_dff_A_TKUk1gsn4_1),.din(n1408));
	jspl jspl_w_n1419_0(.douta(w_n1419_0[0]),.doutb(w_dff_A_9ELLg1NZ1_1),.din(w_dff_B_XYDuZhvK7_2));
	jspl jspl_w_n1426_0(.douta(w_n1426_0[0]),.doutb(w_dff_A_ZZCWqlCV2_1),.din(n1426));
	jspl jspl_w_n1431_0(.douta(w_n1431_0[0]),.doutb(w_n1431_0[1]),.din(w_dff_B_bJorngyd9_2));
	jspl jspl_w_n1433_0(.douta(w_n1433_0[0]),.doutb(w_n1433_0[1]),.din(n1433));
	jspl jspl_w_n1440_0(.douta(w_n1440_0[0]),.doutb(w_n1440_0[1]),.din(n1440));
	jspl3 jspl3_w_n1452_0(.douta(w_dff_A_877u7CnR6_0),.doutb(w_n1452_0[1]),.doutc(w_dff_A_WGaGkLAH1_2),.din(n1452));
	jspl jspl_w_n1458_0(.douta(w_n1458_0[0]),.doutb(w_n1458_0[1]),.din(n1458));
	jspl jspl_w_n1486_0(.douta(w_n1486_0[0]),.doutb(w_n1486_0[1]),.din(n1486));
	jspl jspl_w_n1492_0(.douta(w_n1492_0[0]),.doutb(w_n1492_0[1]),.din(n1492));
	jspl jspl_w_n1506_0(.douta(w_n1506_0[0]),.doutb(w_n1506_0[1]),.din(n1506));
	jspl jspl_w_n1511_0(.douta(w_dff_A_stjFbjlk7_0),.doutb(w_n1511_0[1]),.din(w_dff_B_zsXdLKoc7_2));
	jspl jspl_w_n1518_0(.douta(w_n1518_0[0]),.doutb(w_n1518_0[1]),.din(n1518));
	jspl jspl_w_n1529_0(.douta(w_n1529_0[0]),.doutb(w_n1529_0[1]),.din(n1529));
	jspl jspl_w_n1531_0(.douta(w_n1531_0[0]),.doutb(w_n1531_0[1]),.din(n1531));
	jspl jspl_w_n1534_0(.douta(w_n1534_0[0]),.doutb(w_n1534_0[1]),.din(n1534));
	jspl jspl_w_n1536_0(.douta(w_dff_A_z6sf7Fkn6_0),.doutb(w_n1536_0[1]),.din(n1536));
	jspl jspl_w_n1543_0(.douta(w_n1543_0[0]),.doutb(w_dff_A_nIsRN38t6_1),.din(w_dff_B_B4ZEY8c77_2));
	jspl jspl_w_n1554_0(.douta(w_n1554_0[0]),.doutb(w_n1554_0[1]),.din(n1554));
	jspl3 jspl3_w_n1562_0(.douta(w_dff_A_y1uIFPlM4_0),.doutb(w_dff_A_7W0PCMHr4_1),.doutc(w_n1562_0[2]),.din(n1562));
	jspl jspl_w_n1587_0(.douta(w_n1587_0[0]),.doutb(w_n1587_0[1]),.din(n1587));
	jspl jspl_w_n1597_0(.douta(w_n1597_0[0]),.doutb(w_dff_A_bu5l24mo1_1),.din(w_dff_B_2qDZexht2_2));
	jspl jspl_w_n1605_0(.douta(w_dff_A_qHTQzuGI7_0),.doutb(w_n1605_0[1]),.din(n1605));
	jspl jspl_w_n1607_0(.douta(w_dff_A_WUvdjBcC0_0),.doutb(w_n1607_0[1]),.din(n1607));
	jspl jspl_w_n1610_0(.douta(w_n1610_0[0]),.doutb(w_n1610_0[1]),.din(n1610));
	jspl jspl_w_n1620_0(.douta(w_dff_A_tNhpBkgq5_0),.doutb(w_n1620_0[1]),.din(n1620));
	jspl jspl_w_n1624_0(.douta(w_n1624_0[0]),.doutb(w_n1624_0[1]),.din(n1624));
	jdff dff_A_T5tMKu6E2_0(.dout(w_G5_1[0]),.din(w_dff_A_T5tMKu6E2_0),.clk(gclk));
	jdff dff_A_oNTQhwtA1_1(.dout(w_G5_0[1]),.din(w_dff_A_oNTQhwtA1_1),.clk(gclk));
	jdff dff_A_1a3BOk4N7_2(.dout(w_G5_0[2]),.din(w_dff_A_1a3BOk4N7_2),.clk(gclk));
	jdff dff_B_zOw0FkEF5_2(.din(n347),.dout(w_dff_B_zOw0FkEF5_2),.clk(gclk));
	jdff dff_B_6U6LXPHR6_0(.din(n1072),.dout(w_dff_B_6U6LXPHR6_0),.clk(gclk));
	jdff dff_B_TjLqO1u54_1(.din(n1085),.dout(w_dff_B_TjLqO1u54_1),.clk(gclk));
	jdff dff_B_97wWmE6h6_1(.din(n753),.dout(w_dff_B_97wWmE6h6_1),.clk(gclk));
	jdff dff_B_4VCGVyj24_1(.din(w_dff_B_97wWmE6h6_1),.dout(w_dff_B_4VCGVyj24_1),.clk(gclk));
	jdff dff_B_ufsFaH6f3_1(.din(w_dff_B_4VCGVyj24_1),.dout(w_dff_B_ufsFaH6f3_1),.clk(gclk));
	jdff dff_B_CyEW83ti4_1(.din(w_dff_B_ufsFaH6f3_1),.dout(w_dff_B_CyEW83ti4_1),.clk(gclk));
	jdff dff_B_1jFsO2pC0_1(.din(w_dff_B_CyEW83ti4_1),.dout(w_dff_B_1jFsO2pC0_1),.clk(gclk));
	jdff dff_B_2hcssRmX0_1(.din(w_dff_B_1jFsO2pC0_1),.dout(w_dff_B_2hcssRmX0_1),.clk(gclk));
	jdff dff_B_Fh2yl14E5_1(.din(w_dff_B_2hcssRmX0_1),.dout(w_dff_B_Fh2yl14E5_1),.clk(gclk));
	jdff dff_B_RRky67T19_1(.din(w_dff_B_Fh2yl14E5_1),.dout(w_dff_B_RRky67T19_1),.clk(gclk));
	jdff dff_B_qIlkOmM51_1(.din(w_dff_B_RRky67T19_1),.dout(w_dff_B_qIlkOmM51_1),.clk(gclk));
	jdff dff_B_3HpaRzXJ5_1(.din(w_dff_B_qIlkOmM51_1),.dout(w_dff_B_3HpaRzXJ5_1),.clk(gclk));
	jdff dff_B_kaDHWLyL4_1(.din(w_dff_B_3HpaRzXJ5_1),.dout(w_dff_B_kaDHWLyL4_1),.clk(gclk));
	jdff dff_B_rPJsex3M4_1(.din(w_dff_B_kaDHWLyL4_1),.dout(w_dff_B_rPJsex3M4_1),.clk(gclk));
	jdff dff_B_JcuS8AgU8_1(.din(w_dff_B_rPJsex3M4_1),.dout(w_dff_B_JcuS8AgU8_1),.clk(gclk));
	jdff dff_B_0kzfT6xZ6_1(.din(w_dff_B_JcuS8AgU8_1),.dout(w_dff_B_0kzfT6xZ6_1),.clk(gclk));
	jdff dff_B_SROuIGVL6_1(.din(w_dff_B_0kzfT6xZ6_1),.dout(w_dff_B_SROuIGVL6_1),.clk(gclk));
	jdff dff_B_Tw8HPB605_1(.din(w_dff_B_SROuIGVL6_1),.dout(w_dff_B_Tw8HPB605_1),.clk(gclk));
	jdff dff_B_QEsPxDpC0_1(.din(w_dff_B_Tw8HPB605_1),.dout(w_dff_B_QEsPxDpC0_1),.clk(gclk));
	jdff dff_B_QtIF5Vso0_0(.din(n1057),.dout(w_dff_B_QtIF5Vso0_0),.clk(gclk));
	jdff dff_B_QMWRNQhZ5_0(.din(w_dff_B_QtIF5Vso0_0),.dout(w_dff_B_QMWRNQhZ5_0),.clk(gclk));
	jdff dff_B_li2eQKuw8_0(.din(w_dff_B_QMWRNQhZ5_0),.dout(w_dff_B_li2eQKuw8_0),.clk(gclk));
	jdff dff_B_HpNPKjcS6_0(.din(w_dff_B_li2eQKuw8_0),.dout(w_dff_B_HpNPKjcS6_0),.clk(gclk));
	jdff dff_B_RFd3dZtY3_0(.din(w_dff_B_HpNPKjcS6_0),.dout(w_dff_B_RFd3dZtY3_0),.clk(gclk));
	jdff dff_B_if3aMaBK6_0(.din(w_dff_B_RFd3dZtY3_0),.dout(w_dff_B_if3aMaBK6_0),.clk(gclk));
	jdff dff_B_4nECUVdc6_0(.din(w_dff_B_if3aMaBK6_0),.dout(w_dff_B_4nECUVdc6_0),.clk(gclk));
	jdff dff_B_Vc1PWlxZ1_0(.din(w_dff_B_4nECUVdc6_0),.dout(w_dff_B_Vc1PWlxZ1_0),.clk(gclk));
	jdff dff_B_KWdKesqb8_0(.din(w_dff_B_Vc1PWlxZ1_0),.dout(w_dff_B_KWdKesqb8_0),.clk(gclk));
	jdff dff_B_qOsK37uE5_0(.din(w_dff_B_KWdKesqb8_0),.dout(w_dff_B_qOsK37uE5_0),.clk(gclk));
	jdff dff_B_n2qIGD8l4_0(.din(w_dff_B_qOsK37uE5_0),.dout(w_dff_B_n2qIGD8l4_0),.clk(gclk));
	jdff dff_B_3OPqg3A28_0(.din(w_dff_B_n2qIGD8l4_0),.dout(w_dff_B_3OPqg3A28_0),.clk(gclk));
	jdff dff_B_o4x9k8Hm3_0(.din(w_dff_B_3OPqg3A28_0),.dout(w_dff_B_o4x9k8Hm3_0),.clk(gclk));
	jdff dff_B_dDhKryAR8_0(.din(w_dff_B_o4x9k8Hm3_0),.dout(w_dff_B_dDhKryAR8_0),.clk(gclk));
	jdff dff_B_lLGJXY3r1_0(.din(w_dff_B_dDhKryAR8_0),.dout(w_dff_B_lLGJXY3r1_0),.clk(gclk));
	jdff dff_B_mjsGBemm5_0(.din(w_dff_B_lLGJXY3r1_0),.dout(w_dff_B_mjsGBemm5_0),.clk(gclk));
	jdff dff_B_junc3TOI5_1(.din(n1048),.dout(w_dff_B_junc3TOI5_1),.clk(gclk));
	jdff dff_B_2yB9OqOV3_1(.din(w_dff_B_junc3TOI5_1),.dout(w_dff_B_2yB9OqOV3_1),.clk(gclk));
	jdff dff_B_Et9qnbCU0_1(.din(w_dff_B_2yB9OqOV3_1),.dout(w_dff_B_Et9qnbCU0_1),.clk(gclk));
	jdff dff_B_ANo0zDnp6_1(.din(w_dff_B_Et9qnbCU0_1),.dout(w_dff_B_ANo0zDnp6_1),.clk(gclk));
	jdff dff_B_qkNvFZIn9_1(.din(w_dff_B_ANo0zDnp6_1),.dout(w_dff_B_qkNvFZIn9_1),.clk(gclk));
	jdff dff_B_Mmpnp9mB6_1(.din(n1049),.dout(w_dff_B_Mmpnp9mB6_1),.clk(gclk));
	jdff dff_B_07ZkajnW5_1(.din(w_dff_B_Mmpnp9mB6_1),.dout(w_dff_B_07ZkajnW5_1),.clk(gclk));
	jdff dff_B_Mu0xTX3i7_1(.din(w_dff_B_07ZkajnW5_1),.dout(w_dff_B_Mu0xTX3i7_1),.clk(gclk));
	jdff dff_B_gHZo3aqe3_1(.din(n1050),.dout(w_dff_B_gHZo3aqe3_1),.clk(gclk));
	jdff dff_B_imUXYW195_0(.din(n1044),.dout(w_dff_B_imUXYW195_0),.clk(gclk));
	jdff dff_B_JO3UKFHT7_0(.din(w_dff_B_imUXYW195_0),.dout(w_dff_B_JO3UKFHT7_0),.clk(gclk));
	jdff dff_B_v38kqikO1_0(.din(w_dff_B_JO3UKFHT7_0),.dout(w_dff_B_v38kqikO1_0),.clk(gclk));
	jdff dff_B_kcXzZ2IU4_0(.din(w_dff_B_v38kqikO1_0),.dout(w_dff_B_kcXzZ2IU4_0),.clk(gclk));
	jdff dff_B_Bm2F6y6y6_0(.din(w_dff_B_kcXzZ2IU4_0),.dout(w_dff_B_Bm2F6y6y6_0),.clk(gclk));
	jdff dff_B_H57zb1K81_0(.din(w_dff_B_Bm2F6y6y6_0),.dout(w_dff_B_H57zb1K81_0),.clk(gclk));
	jdff dff_B_Xa7VGz1K9_0(.din(w_dff_B_H57zb1K81_0),.dout(w_dff_B_Xa7VGz1K9_0),.clk(gclk));
	jdff dff_B_6E66sqbu1_0(.din(w_dff_B_Xa7VGz1K9_0),.dout(w_dff_B_6E66sqbu1_0),.clk(gclk));
	jdff dff_B_73ua5IHw6_0(.din(w_dff_B_6E66sqbu1_0),.dout(w_dff_B_73ua5IHw6_0),.clk(gclk));
	jdff dff_B_2ocE5viI8_0(.din(w_dff_B_73ua5IHw6_0),.dout(w_dff_B_2ocE5viI8_0),.clk(gclk));
	jdff dff_B_uGZGQZJL0_0(.din(w_dff_B_2ocE5viI8_0),.dout(w_dff_B_uGZGQZJL0_0),.clk(gclk));
	jdff dff_B_GScmS10K5_0(.din(w_dff_B_uGZGQZJL0_0),.dout(w_dff_B_GScmS10K5_0),.clk(gclk));
	jdff dff_B_VJyiFUPr6_0(.din(w_dff_B_GScmS10K5_0),.dout(w_dff_B_VJyiFUPr6_0),.clk(gclk));
	jdff dff_B_v7D954u79_0(.din(w_dff_B_VJyiFUPr6_0),.dout(w_dff_B_v7D954u79_0),.clk(gclk));
	jdff dff_B_0sRoyxnh1_0(.din(w_dff_B_v7D954u79_0),.dout(w_dff_B_0sRoyxnh1_0),.clk(gclk));
	jdff dff_B_c7MJRDtg1_0(.din(w_dff_B_0sRoyxnh1_0),.dout(w_dff_B_c7MJRDtg1_0),.clk(gclk));
	jdff dff_B_ZR0Rcscs5_0(.din(w_dff_B_c7MJRDtg1_0),.dout(w_dff_B_ZR0Rcscs5_0),.clk(gclk));
	jdff dff_B_kJItpt9r0_1(.din(n1040),.dout(w_dff_B_kJItpt9r0_1),.clk(gclk));
	jdff dff_B_4WtbBNc87_1(.din(w_dff_B_kJItpt9r0_1),.dout(w_dff_B_4WtbBNc87_1),.clk(gclk));
	jdff dff_A_CphRJuGg1_0(.dout(w_n1042_0[0]),.din(w_dff_A_CphRJuGg1_0),.clk(gclk));
	jdff dff_B_55reXz6K6_1(.din(n790),.dout(w_dff_B_55reXz6K6_1),.clk(gclk));
	jdff dff_B_AQ3bK5jI6_1(.din(w_dff_B_55reXz6K6_1),.dout(w_dff_B_AQ3bK5jI6_1),.clk(gclk));
	jdff dff_B_9ccSpmjd7_1(.din(w_dff_B_AQ3bK5jI6_1),.dout(w_dff_B_9ccSpmjd7_1),.clk(gclk));
	jdff dff_B_QBQeBDuX0_1(.din(w_dff_B_9ccSpmjd7_1),.dout(w_dff_B_QBQeBDuX0_1),.clk(gclk));
	jdff dff_B_ikunosyf0_1(.din(w_dff_B_QBQeBDuX0_1),.dout(w_dff_B_ikunosyf0_1),.clk(gclk));
	jdff dff_B_2xlYf5BN1_1(.din(w_dff_B_ikunosyf0_1),.dout(w_dff_B_2xlYf5BN1_1),.clk(gclk));
	jdff dff_B_KJhSDUHe8_1(.din(w_dff_B_2xlYf5BN1_1),.dout(w_dff_B_KJhSDUHe8_1),.clk(gclk));
	jdff dff_B_AtHwi2QQ7_1(.din(w_dff_B_KJhSDUHe8_1),.dout(w_dff_B_AtHwi2QQ7_1),.clk(gclk));
	jdff dff_B_UggBC4N44_1(.din(w_dff_B_AtHwi2QQ7_1),.dout(w_dff_B_UggBC4N44_1),.clk(gclk));
	jdff dff_B_lwHLunpJ9_1(.din(w_dff_B_UggBC4N44_1),.dout(w_dff_B_lwHLunpJ9_1),.clk(gclk));
	jdff dff_B_2rjIlNi35_1(.din(w_dff_B_lwHLunpJ9_1),.dout(w_dff_B_2rjIlNi35_1),.clk(gclk));
	jdff dff_B_Gkd9alQJ7_1(.din(w_dff_B_2rjIlNi35_1),.dout(w_dff_B_Gkd9alQJ7_1),.clk(gclk));
	jdff dff_B_Xp10PR8c9_1(.din(w_dff_B_Gkd9alQJ7_1),.dout(w_dff_B_Xp10PR8c9_1),.clk(gclk));
	jdff dff_B_3C0Jcu5e6_1(.din(w_dff_B_Xp10PR8c9_1),.dout(w_dff_B_3C0Jcu5e6_1),.clk(gclk));
	jdff dff_B_XhyAd35E2_1(.din(w_dff_B_3C0Jcu5e6_1),.dout(w_dff_B_XhyAd35E2_1),.clk(gclk));
	jdff dff_B_iUyAeNp71_1(.din(n794),.dout(w_dff_B_iUyAeNp71_1),.clk(gclk));
	jdff dff_B_LYCb3kK50_1(.din(w_dff_B_iUyAeNp71_1),.dout(w_dff_B_LYCb3kK50_1),.clk(gclk));
	jdff dff_B_BEKYu4Ds1_1(.din(w_dff_B_LYCb3kK50_1),.dout(w_dff_B_BEKYu4Ds1_1),.clk(gclk));
	jdff dff_B_n5fF0UMc1_1(.din(w_dff_B_BEKYu4Ds1_1),.dout(w_dff_B_n5fF0UMc1_1),.clk(gclk));
	jdff dff_B_0hEaJtkG7_1(.din(w_dff_B_n5fF0UMc1_1),.dout(w_dff_B_0hEaJtkG7_1),.clk(gclk));
	jdff dff_B_ABL8kD7e8_1(.din(w_dff_B_0hEaJtkG7_1),.dout(w_dff_B_ABL8kD7e8_1),.clk(gclk));
	jdff dff_B_6oJjkDGb9_1(.din(w_dff_B_ABL8kD7e8_1),.dout(w_dff_B_6oJjkDGb9_1),.clk(gclk));
	jdff dff_B_BpEyDqFM3_1(.din(w_dff_B_6oJjkDGb9_1),.dout(w_dff_B_BpEyDqFM3_1),.clk(gclk));
	jdff dff_B_TTQ6jrHG5_1(.din(w_dff_B_BpEyDqFM3_1),.dout(w_dff_B_TTQ6jrHG5_1),.clk(gclk));
	jdff dff_B_kD2uZm3u0_1(.din(w_dff_B_TTQ6jrHG5_1),.dout(w_dff_B_kD2uZm3u0_1),.clk(gclk));
	jdff dff_B_PLBi3gOJ4_1(.din(w_dff_B_kD2uZm3u0_1),.dout(w_dff_B_PLBi3gOJ4_1),.clk(gclk));
	jdff dff_B_PkwjJBL94_1(.din(w_dff_B_PLBi3gOJ4_1),.dout(w_dff_B_PkwjJBL94_1),.clk(gclk));
	jdff dff_B_eeLuYLuh1_1(.din(w_dff_B_PkwjJBL94_1),.dout(w_dff_B_eeLuYLuh1_1),.clk(gclk));
	jdff dff_B_AN1m9qJC1_1(.din(w_dff_B_eeLuYLuh1_1),.dout(w_dff_B_AN1m9qJC1_1),.clk(gclk));
	jdff dff_B_2GmbTt8p1_1(.din(w_dff_B_AN1m9qJC1_1),.dout(w_dff_B_2GmbTt8p1_1),.clk(gclk));
	jdff dff_B_tnrcfJL44_0(.din(n1036),.dout(w_dff_B_tnrcfJL44_0),.clk(gclk));
	jdff dff_B_YTrADmT94_0(.din(w_dff_B_tnrcfJL44_0),.dout(w_dff_B_YTrADmT94_0),.clk(gclk));
	jdff dff_B_JUkwTrJG5_0(.din(w_dff_B_YTrADmT94_0),.dout(w_dff_B_JUkwTrJG5_0),.clk(gclk));
	jdff dff_B_87pkms7O0_0(.din(w_dff_B_JUkwTrJG5_0),.dout(w_dff_B_87pkms7O0_0),.clk(gclk));
	jdff dff_B_V7NRqf8f6_0(.din(w_dff_B_87pkms7O0_0),.dout(w_dff_B_V7NRqf8f6_0),.clk(gclk));
	jdff dff_B_uwiXtHGO0_0(.din(w_dff_B_V7NRqf8f6_0),.dout(w_dff_B_uwiXtHGO0_0),.clk(gclk));
	jdff dff_B_xsDK7qTa1_0(.din(w_dff_B_uwiXtHGO0_0),.dout(w_dff_B_xsDK7qTa1_0),.clk(gclk));
	jdff dff_B_2xUTUYxk9_0(.din(w_dff_B_xsDK7qTa1_0),.dout(w_dff_B_2xUTUYxk9_0),.clk(gclk));
	jdff dff_B_DalyDTKL9_0(.din(w_dff_B_2xUTUYxk9_0),.dout(w_dff_B_DalyDTKL9_0),.clk(gclk));
	jdff dff_B_hrGNiiTO6_0(.din(w_dff_B_DalyDTKL9_0),.dout(w_dff_B_hrGNiiTO6_0),.clk(gclk));
	jdff dff_B_B3aBrb1W9_0(.din(w_dff_B_hrGNiiTO6_0),.dout(w_dff_B_B3aBrb1W9_0),.clk(gclk));
	jdff dff_B_hc5zIjFW5_0(.din(w_dff_B_B3aBrb1W9_0),.dout(w_dff_B_hc5zIjFW5_0),.clk(gclk));
	jdff dff_B_NzmYv2Ju3_0(.din(w_dff_B_hc5zIjFW5_0),.dout(w_dff_B_NzmYv2Ju3_0),.clk(gclk));
	jdff dff_B_JFomYLpH8_0(.din(w_dff_B_NzmYv2Ju3_0),.dout(w_dff_B_JFomYLpH8_0),.clk(gclk));
	jdff dff_B_VNYPqclP3_0(.din(w_dff_B_JFomYLpH8_0),.dout(w_dff_B_VNYPqclP3_0),.clk(gclk));
	jdff dff_B_ZwTl6rAk0_0(.din(w_dff_B_VNYPqclP3_0),.dout(w_dff_B_ZwTl6rAk0_0),.clk(gclk));
	jdff dff_B_mwrMtZeR5_1(.din(n842),.dout(w_dff_B_mwrMtZeR5_1),.clk(gclk));
	jdff dff_B_QCwqzs4K5_1(.din(w_dff_B_mwrMtZeR5_1),.dout(w_dff_B_QCwqzs4K5_1),.clk(gclk));
	jdff dff_B_KrCqQOpC8_1(.din(w_dff_B_QCwqzs4K5_1),.dout(w_dff_B_KrCqQOpC8_1),.clk(gclk));
	jdff dff_B_VYSGL44K4_1(.din(w_dff_B_KrCqQOpC8_1),.dout(w_dff_B_VYSGL44K4_1),.clk(gclk));
	jdff dff_B_y0iAhE1x1_1(.din(w_dff_B_VYSGL44K4_1),.dout(w_dff_B_y0iAhE1x1_1),.clk(gclk));
	jdff dff_B_gaAUvedO2_1(.din(w_dff_B_y0iAhE1x1_1),.dout(w_dff_B_gaAUvedO2_1),.clk(gclk));
	jdff dff_B_DDaQ0Nhf4_1(.din(w_dff_B_gaAUvedO2_1),.dout(w_dff_B_DDaQ0Nhf4_1),.clk(gclk));
	jdff dff_B_Awj8k4IR0_1(.din(w_dff_B_DDaQ0Nhf4_1),.dout(w_dff_B_Awj8k4IR0_1),.clk(gclk));
	jdff dff_B_djD8XoOW9_1(.din(w_dff_B_Awj8k4IR0_1),.dout(w_dff_B_djD8XoOW9_1),.clk(gclk));
	jdff dff_B_l9p2k1Q35_1(.din(w_dff_B_djD8XoOW9_1),.dout(w_dff_B_l9p2k1Q35_1),.clk(gclk));
	jdff dff_B_CXoIoVTw8_1(.din(w_dff_B_l9p2k1Q35_1),.dout(w_dff_B_CXoIoVTw8_1),.clk(gclk));
	jdff dff_B_4QyVYSAf5_1(.din(n843),.dout(w_dff_B_4QyVYSAf5_1),.clk(gclk));
	jdff dff_B_H3Db3hF04_1(.din(w_dff_B_4QyVYSAf5_1),.dout(w_dff_B_H3Db3hF04_1),.clk(gclk));
	jdff dff_B_H15ONvw94_1(.din(w_dff_B_H3Db3hF04_1),.dout(w_dff_B_H15ONvw94_1),.clk(gclk));
	jdff dff_B_5Te35amx6_1(.din(w_dff_B_H15ONvw94_1),.dout(w_dff_B_5Te35amx6_1),.clk(gclk));
	jdff dff_B_d2014slu1_1(.din(w_dff_B_5Te35amx6_1),.dout(w_dff_B_d2014slu1_1),.clk(gclk));
	jdff dff_B_Fv9Tf1Do3_1(.din(w_dff_B_d2014slu1_1),.dout(w_dff_B_Fv9Tf1Do3_1),.clk(gclk));
	jdff dff_B_IeXeeWmW2_1(.din(w_dff_B_Fv9Tf1Do3_1),.dout(w_dff_B_IeXeeWmW2_1),.clk(gclk));
	jdff dff_B_BbmWtOQG4_1(.din(w_dff_B_IeXeeWmW2_1),.dout(w_dff_B_BbmWtOQG4_1),.clk(gclk));
	jdff dff_B_h8N6Mso09_1(.din(w_dff_B_BbmWtOQG4_1),.dout(w_dff_B_h8N6Mso09_1),.clk(gclk));
	jdff dff_B_Esn3nXfG9_1(.din(w_dff_B_h8N6Mso09_1),.dout(w_dff_B_Esn3nXfG9_1),.clk(gclk));
	jdff dff_B_3XYmJmJV0_1(.din(w_dff_B_Esn3nXfG9_1),.dout(w_dff_B_3XYmJmJV0_1),.clk(gclk));
	jdff dff_B_c8bI1Gsq5_1(.din(w_dff_B_3XYmJmJV0_1),.dout(w_dff_B_c8bI1Gsq5_1),.clk(gclk));
	jdff dff_B_VFnSsohA1_1(.din(w_dff_B_c8bI1Gsq5_1),.dout(w_dff_B_VFnSsohA1_1),.clk(gclk));
	jdff dff_B_9EZCnDqB9_0(.din(n1031),.dout(w_dff_B_9EZCnDqB9_0),.clk(gclk));
	jdff dff_B_krIL2Sla4_0(.din(w_dff_B_9EZCnDqB9_0),.dout(w_dff_B_krIL2Sla4_0),.clk(gclk));
	jdff dff_B_vIDtoBo01_0(.din(w_dff_B_krIL2Sla4_0),.dout(w_dff_B_vIDtoBo01_0),.clk(gclk));
	jdff dff_B_WfQNlUCq7_0(.din(w_dff_B_vIDtoBo01_0),.dout(w_dff_B_WfQNlUCq7_0),.clk(gclk));
	jdff dff_B_oI7Ro3ve0_0(.din(w_dff_B_WfQNlUCq7_0),.dout(w_dff_B_oI7Ro3ve0_0),.clk(gclk));
	jdff dff_B_RZ1doWGM3_0(.din(w_dff_B_oI7Ro3ve0_0),.dout(w_dff_B_RZ1doWGM3_0),.clk(gclk));
	jdff dff_B_bTzE2Vb16_0(.din(w_dff_B_RZ1doWGM3_0),.dout(w_dff_B_bTzE2Vb16_0),.clk(gclk));
	jdff dff_B_UKak35Q27_0(.din(w_dff_B_bTzE2Vb16_0),.dout(w_dff_B_UKak35Q27_0),.clk(gclk));
	jdff dff_B_47WPA4wK6_0(.din(w_dff_B_UKak35Q27_0),.dout(w_dff_B_47WPA4wK6_0),.clk(gclk));
	jdff dff_B_sy7JW3no2_0(.din(w_dff_B_47WPA4wK6_0),.dout(w_dff_B_sy7JW3no2_0),.clk(gclk));
	jdff dff_B_SEsKKMeJ7_0(.din(w_dff_B_sy7JW3no2_0),.dout(w_dff_B_SEsKKMeJ7_0),.clk(gclk));
	jdff dff_B_clx5t3Ka4_0(.din(w_dff_B_SEsKKMeJ7_0),.dout(w_dff_B_clx5t3Ka4_0),.clk(gclk));
	jdff dff_B_hr7f8krV9_0(.din(w_dff_B_clx5t3Ka4_0),.dout(w_dff_B_hr7f8krV9_0),.clk(gclk));
	jdff dff_B_AdyRxg5x1_0(.din(w_dff_B_hr7f8krV9_0),.dout(w_dff_B_AdyRxg5x1_0),.clk(gclk));
	jdff dff_B_AL4TOg2N8_0(.din(n841),.dout(w_dff_B_AL4TOg2N8_0),.clk(gclk));
	jdff dff_B_zMHrUpc90_0(.din(w_dff_B_AL4TOg2N8_0),.dout(w_dff_B_zMHrUpc90_0),.clk(gclk));
	jdff dff_B_yE5DwyML5_1(.din(n837),.dout(w_dff_B_yE5DwyML5_1),.clk(gclk));
	jdff dff_B_FWBTaxcO4_1(.din(n830),.dout(w_dff_B_FWBTaxcO4_1),.clk(gclk));
	jdff dff_B_9aw3Afxr6_0(.din(n828),.dout(w_dff_B_9aw3Afxr6_0),.clk(gclk));
	jdff dff_A_Eg7cyhMt0_1(.dout(w_n808_0[1]),.din(w_dff_A_Eg7cyhMt0_1),.clk(gclk));
	jdff dff_A_KeH7Nrrb3_1(.dout(w_dff_A_Eg7cyhMt0_1),.din(w_dff_A_KeH7Nrrb3_1),.clk(gclk));
	jdff dff_B_Ddj01x9g8_0(.din(n789),.dout(w_dff_B_Ddj01x9g8_0),.clk(gclk));
	jdff dff_B_O1JLdrLw2_1(.din(n785),.dout(w_dff_B_O1JLdrLw2_1),.clk(gclk));
	jdff dff_A_enWUTCuu1_1(.dout(w_n773_0[1]),.din(w_dff_A_enWUTCuu1_1),.clk(gclk));
	jdff dff_B_E8nBb3DH5_2(.din(n766),.dout(w_dff_B_E8nBb3DH5_2),.clk(gclk));
	jdff dff_B_XAAgdeGg2_1(.din(n730),.dout(w_dff_B_XAAgdeGg2_1),.clk(gclk));
	jdff dff_B_I5FCwES43_1(.din(w_dff_B_XAAgdeGg2_1),.dout(w_dff_B_I5FCwES43_1),.clk(gclk));
	jdff dff_B_MlLdonTk2_1(.din(w_dff_B_I5FCwES43_1),.dout(w_dff_B_MlLdonTk2_1),.clk(gclk));
	jdff dff_B_sGNYDTMf1_1(.din(n731),.dout(w_dff_B_sGNYDTMf1_1),.clk(gclk));
	jdff dff_B_2G7vtFay6_1(.din(w_dff_B_sGNYDTMf1_1),.dout(w_dff_B_2G7vtFay6_1),.clk(gclk));
	jdff dff_B_Dt6dA6I30_1(.din(n735),.dout(w_dff_B_Dt6dA6I30_1),.clk(gclk));
	jdff dff_A_JsJXQnTB5_1(.dout(w_n724_0[1]),.din(w_dff_A_JsJXQnTB5_1),.clk(gclk));
	jdff dff_A_RZ0RSApD5_1(.dout(w_dff_A_JsJXQnTB5_1),.din(w_dff_A_RZ0RSApD5_1),.clk(gclk));
	jdff dff_A_oi0Er4UG6_1(.dout(w_dff_A_RZ0RSApD5_1),.din(w_dff_A_oi0Er4UG6_1),.clk(gclk));
	jdff dff_A_M57ltLga8_1(.dout(w_dff_A_oi0Er4UG6_1),.din(w_dff_A_M57ltLga8_1),.clk(gclk));
	jdff dff_B_wkAoRgPc7_3(.din(n718),.dout(w_dff_B_wkAoRgPc7_3),.clk(gclk));
	jdff dff_B_PmmN9UCR7_3(.din(w_dff_B_wkAoRgPc7_3),.dout(w_dff_B_PmmN9UCR7_3),.clk(gclk));
	jdff dff_B_AhAyDMWW2_3(.din(w_dff_B_PmmN9UCR7_3),.dout(w_dff_B_AhAyDMWW2_3),.clk(gclk));
	jdff dff_B_5lKdJiw20_3(.din(w_dff_B_AhAyDMWW2_3),.dout(w_dff_B_5lKdJiw20_3),.clk(gclk));
	jdff dff_B_Fx4k30Tr9_3(.din(w_dff_B_5lKdJiw20_3),.dout(w_dff_B_Fx4k30Tr9_3),.clk(gclk));
	jdff dff_B_dF9Rz8HV0_3(.din(w_dff_B_Fx4k30Tr9_3),.dout(w_dff_B_dF9Rz8HV0_3),.clk(gclk));
	jdff dff_B_QlWGqAmt3_3(.din(w_dff_B_dF9Rz8HV0_3),.dout(w_dff_B_QlWGqAmt3_3),.clk(gclk));
	jdff dff_B_QH6vNJpY5_3(.din(w_dff_B_QlWGqAmt3_3),.dout(w_dff_B_QH6vNJpY5_3),.clk(gclk));
	jdff dff_B_5cdujKON1_3(.din(w_dff_B_QH6vNJpY5_3),.dout(w_dff_B_5cdujKON1_3),.clk(gclk));
	jdff dff_B_QrESFXZm3_3(.din(w_dff_B_5cdujKON1_3),.dout(w_dff_B_QrESFXZm3_3),.clk(gclk));
	jdff dff_B_wUXpcn6J7_3(.din(w_dff_B_QrESFXZm3_3),.dout(w_dff_B_wUXpcn6J7_3),.clk(gclk));
	jdff dff_B_wBxjDCTh1_3(.din(w_dff_B_wUXpcn6J7_3),.dout(w_dff_B_wBxjDCTh1_3),.clk(gclk));
	jdff dff_B_AuPEkyDQ4_3(.din(w_dff_B_wBxjDCTh1_3),.dout(w_dff_B_AuPEkyDQ4_3),.clk(gclk));
	jdff dff_B_9XVIZCmG7_3(.din(w_dff_B_AuPEkyDQ4_3),.dout(w_dff_B_9XVIZCmG7_3),.clk(gclk));
	jdff dff_B_pplEk7n83_3(.din(w_dff_B_9XVIZCmG7_3),.dout(w_dff_B_pplEk7n83_3),.clk(gclk));
	jdff dff_B_WO7SOUzB9_3(.din(w_dff_B_pplEk7n83_3),.dout(w_dff_B_WO7SOUzB9_3),.clk(gclk));
	jdff dff_B_RgiMDdgi4_3(.din(w_dff_B_WO7SOUzB9_3),.dout(w_dff_B_RgiMDdgi4_3),.clk(gclk));
	jdff dff_B_3CbOvO5n8_3(.din(w_dff_B_RgiMDdgi4_3),.dout(w_dff_B_3CbOvO5n8_3),.clk(gclk));
	jdff dff_B_4R7OiaOD7_3(.din(w_dff_B_3CbOvO5n8_3),.dout(w_dff_B_4R7OiaOD7_3),.clk(gclk));
	jdff dff_B_rj9Ym2rU0_3(.din(w_dff_B_4R7OiaOD7_3),.dout(w_dff_B_rj9Ym2rU0_3),.clk(gclk));
	jdff dff_B_fV29Gfar9_3(.din(w_dff_B_rj9Ym2rU0_3),.dout(w_dff_B_fV29Gfar9_3),.clk(gclk));
	jdff dff_B_HSiGjv8v6_3(.din(w_dff_B_fV29Gfar9_3),.dout(w_dff_B_HSiGjv8v6_3),.clk(gclk));
	jdff dff_B_3zJjK5z10_3(.din(w_dff_B_HSiGjv8v6_3),.dout(w_dff_B_3zJjK5z10_3),.clk(gclk));
	jdff dff_B_KT5fBCnk8_3(.din(w_dff_B_3zJjK5z10_3),.dout(w_dff_B_KT5fBCnk8_3),.clk(gclk));
	jdff dff_B_HX5r9EjC7_0(.din(n717),.dout(w_dff_B_HX5r9EjC7_0),.clk(gclk));
	jdff dff_B_ppAVmaDk9_1(.din(n1305),.dout(w_dff_B_ppAVmaDk9_1),.clk(gclk));
	jdff dff_B_jGtEyOsT0_1(.din(w_dff_B_ppAVmaDk9_1),.dout(w_dff_B_jGtEyOsT0_1),.clk(gclk));
	jdff dff_B_APeBZFjU6_1(.din(w_dff_B_jGtEyOsT0_1),.dout(w_dff_B_APeBZFjU6_1),.clk(gclk));
	jdff dff_B_jzw1SDOq0_1(.din(w_dff_B_APeBZFjU6_1),.dout(w_dff_B_jzw1SDOq0_1),.clk(gclk));
	jdff dff_B_NUTPwWig2_1(.din(w_dff_B_jzw1SDOq0_1),.dout(w_dff_B_NUTPwWig2_1),.clk(gclk));
	jdff dff_B_aFKDUAAb1_1(.din(w_dff_B_NUTPwWig2_1),.dout(w_dff_B_aFKDUAAb1_1),.clk(gclk));
	jdff dff_B_pYbMP1xr9_1(.din(w_dff_B_aFKDUAAb1_1),.dout(w_dff_B_pYbMP1xr9_1),.clk(gclk));
	jdff dff_B_WWZoYfmp3_1(.din(w_dff_B_pYbMP1xr9_1),.dout(w_dff_B_WWZoYfmp3_1),.clk(gclk));
	jdff dff_B_BqJSAS7T3_1(.din(w_dff_B_WWZoYfmp3_1),.dout(w_dff_B_BqJSAS7T3_1),.clk(gclk));
	jdff dff_B_7XmpVo0t3_1(.din(w_dff_B_BqJSAS7T3_1),.dout(w_dff_B_7XmpVo0t3_1),.clk(gclk));
	jdff dff_B_5QrLIniJ8_1(.din(w_dff_B_7XmpVo0t3_1),.dout(w_dff_B_5QrLIniJ8_1),.clk(gclk));
	jdff dff_B_ANLS58eZ7_1(.din(w_dff_B_5QrLIniJ8_1),.dout(w_dff_B_ANLS58eZ7_1),.clk(gclk));
	jdff dff_B_VZtkMsey5_1(.din(w_dff_B_ANLS58eZ7_1),.dout(w_dff_B_VZtkMsey5_1),.clk(gclk));
	jdff dff_B_ZdGQvklp9_1(.din(w_dff_B_VZtkMsey5_1),.dout(w_dff_B_ZdGQvklp9_1),.clk(gclk));
	jdff dff_B_T1FzLBe52_1(.din(w_dff_B_ZdGQvklp9_1),.dout(w_dff_B_T1FzLBe52_1),.clk(gclk));
	jdff dff_B_g0FDj0mJ9_1(.din(w_dff_B_T1FzLBe52_1),.dout(w_dff_B_g0FDj0mJ9_1),.clk(gclk));
	jdff dff_B_ZsfmaTUk9_1(.din(w_dff_B_g0FDj0mJ9_1),.dout(w_dff_B_ZsfmaTUk9_1),.clk(gclk));
	jdff dff_B_yhjINwvk2_1(.din(w_dff_B_ZsfmaTUk9_1),.dout(w_dff_B_yhjINwvk2_1),.clk(gclk));
	jdff dff_B_D2oOjfBR4_1(.din(w_dff_B_yhjINwvk2_1),.dout(w_dff_B_D2oOjfBR4_1),.clk(gclk));
	jdff dff_B_le0XpBTs7_1(.din(w_dff_B_D2oOjfBR4_1),.dout(w_dff_B_le0XpBTs7_1),.clk(gclk));
	jdff dff_B_A7AGMUKI9_1(.din(w_dff_B_le0XpBTs7_1),.dout(w_dff_B_A7AGMUKI9_1),.clk(gclk));
	jdff dff_B_fnd0kqBg8_1(.din(w_dff_B_A7AGMUKI9_1),.dout(w_dff_B_fnd0kqBg8_1),.clk(gclk));
	jdff dff_B_2nEbmhW49_1(.din(n880),.dout(w_dff_B_2nEbmhW49_1),.clk(gclk));
	jdff dff_B_WRoDaIlx8_1(.din(w_dff_B_2nEbmhW49_1),.dout(w_dff_B_WRoDaIlx8_1),.clk(gclk));
	jdff dff_B_c96qlGPT9_1(.din(w_dff_B_WRoDaIlx8_1),.dout(w_dff_B_c96qlGPT9_1),.clk(gclk));
	jdff dff_B_DIMC7OCW0_1(.din(w_dff_B_c96qlGPT9_1),.dout(w_dff_B_DIMC7OCW0_1),.clk(gclk));
	jdff dff_B_0xnUJhc19_1(.din(w_dff_B_DIMC7OCW0_1),.dout(w_dff_B_0xnUJhc19_1),.clk(gclk));
	jdff dff_B_CEqWA62t8_1(.din(w_dff_B_0xnUJhc19_1),.dout(w_dff_B_CEqWA62t8_1),.clk(gclk));
	jdff dff_B_ahWALvHo2_1(.din(w_dff_B_CEqWA62t8_1),.dout(w_dff_B_ahWALvHo2_1),.clk(gclk));
	jdff dff_B_oOPoAVln8_1(.din(w_dff_B_ahWALvHo2_1),.dout(w_dff_B_oOPoAVln8_1),.clk(gclk));
	jdff dff_B_1JamPVks3_1(.din(w_dff_B_oOPoAVln8_1),.dout(w_dff_B_1JamPVks3_1),.clk(gclk));
	jdff dff_B_bwgk3luk8_1(.din(n883),.dout(w_dff_B_bwgk3luk8_1),.clk(gclk));
	jdff dff_B_1NeJ41o38_1(.din(w_dff_B_bwgk3luk8_1),.dout(w_dff_B_1NeJ41o38_1),.clk(gclk));
	jdff dff_B_Zh41odSJ6_1(.din(w_dff_B_1NeJ41o38_1),.dout(w_dff_B_Zh41odSJ6_1),.clk(gclk));
	jdff dff_B_ROdLkkHL3_1(.din(w_dff_B_Zh41odSJ6_1),.dout(w_dff_B_ROdLkkHL3_1),.clk(gclk));
	jdff dff_B_lsmqHwtk6_1(.din(w_dff_B_ROdLkkHL3_1),.dout(w_dff_B_lsmqHwtk6_1),.clk(gclk));
	jdff dff_B_LXeHp9zA5_1(.din(w_dff_B_lsmqHwtk6_1),.dout(w_dff_B_LXeHp9zA5_1),.clk(gclk));
	jdff dff_B_xkwPng879_1(.din(w_dff_B_LXeHp9zA5_1),.dout(w_dff_B_xkwPng879_1),.clk(gclk));
	jdff dff_B_YUPn6mdh1_1(.din(w_dff_B_xkwPng879_1),.dout(w_dff_B_YUPn6mdh1_1),.clk(gclk));
	jdff dff_B_SnQXJfha5_1(.din(w_dff_B_YUPn6mdh1_1),.dout(w_dff_B_SnQXJfha5_1),.clk(gclk));
	jdff dff_B_Y4vEEvQ13_1(.din(w_dff_B_SnQXJfha5_1),.dout(w_dff_B_Y4vEEvQ13_1),.clk(gclk));
	jdff dff_B_3PRK96Yo5_0(.din(n1027),.dout(w_dff_B_3PRK96Yo5_0),.clk(gclk));
	jdff dff_B_CexrjSCz3_0(.din(w_dff_B_3PRK96Yo5_0),.dout(w_dff_B_CexrjSCz3_0),.clk(gclk));
	jdff dff_B_n1cRIjSk2_0(.din(w_dff_B_CexrjSCz3_0),.dout(w_dff_B_n1cRIjSk2_0),.clk(gclk));
	jdff dff_B_U8Mv3Hj79_0(.din(w_dff_B_n1cRIjSk2_0),.dout(w_dff_B_U8Mv3Hj79_0),.clk(gclk));
	jdff dff_B_ZSzFuQvI4_0(.din(w_dff_B_U8Mv3Hj79_0),.dout(w_dff_B_ZSzFuQvI4_0),.clk(gclk));
	jdff dff_B_oaJJPAP00_0(.din(w_dff_B_ZSzFuQvI4_0),.dout(w_dff_B_oaJJPAP00_0),.clk(gclk));
	jdff dff_B_SphKZ9Px2_0(.din(w_dff_B_oaJJPAP00_0),.dout(w_dff_B_SphKZ9Px2_0),.clk(gclk));
	jdff dff_B_w7bN5dAK4_0(.din(w_dff_B_SphKZ9Px2_0),.dout(w_dff_B_w7bN5dAK4_0),.clk(gclk));
	jdff dff_B_0Tk8qq6q4_0(.din(w_dff_B_w7bN5dAK4_0),.dout(w_dff_B_0Tk8qq6q4_0),.clk(gclk));
	jdff dff_B_0r9O8Azb5_0(.din(n1023),.dout(w_dff_B_0r9O8Azb5_0),.clk(gclk));
	jdff dff_B_qT45hAnc6_0(.din(w_dff_B_0r9O8Azb5_0),.dout(w_dff_B_qT45hAnc6_0),.clk(gclk));
	jdff dff_B_jnT5tqD47_0(.din(w_dff_B_qT45hAnc6_0),.dout(w_dff_B_jnT5tqD47_0),.clk(gclk));
	jdff dff_B_AduYHKX63_1(.din(n1017),.dout(w_dff_B_AduYHKX63_1),.clk(gclk));
	jdff dff_B_77aJXqCp8_1(.din(w_dff_B_AduYHKX63_1),.dout(w_dff_B_77aJXqCp8_1),.clk(gclk));
	jdff dff_B_9VJ5u3Ms8_1(.din(w_dff_B_77aJXqCp8_1),.dout(w_dff_B_9VJ5u3Ms8_1),.clk(gclk));
	jdff dff_B_lDVCWs0x5_1(.din(w_dff_B_9VJ5u3Ms8_1),.dout(w_dff_B_lDVCWs0x5_1),.clk(gclk));
	jdff dff_B_woLyC5fT9_0(.din(n1021),.dout(w_dff_B_woLyC5fT9_0),.clk(gclk));
	jdff dff_B_A6CLlKNI3_0(.din(w_dff_B_woLyC5fT9_0),.dout(w_dff_B_A6CLlKNI3_0),.clk(gclk));
	jdff dff_B_T6Uv8ky34_1(.din(n1013),.dout(w_dff_B_T6Uv8ky34_1),.clk(gclk));
	jdff dff_B_rCzq5duE1_0(.din(n1011),.dout(w_dff_B_rCzq5duE1_0),.clk(gclk));
	jdff dff_B_H3R4MueT7_0(.din(w_dff_B_rCzq5duE1_0),.dout(w_dff_B_H3R4MueT7_0),.clk(gclk));
	jdff dff_B_XuQVTKfc1_0(.din(w_dff_B_H3R4MueT7_0),.dout(w_dff_B_XuQVTKfc1_0),.clk(gclk));
	jdff dff_B_qNMshn2w7_1(.din(n971),.dout(w_dff_B_qNMshn2w7_1),.clk(gclk));
	jdff dff_B_xTcMbHgz3_1(.din(w_dff_B_qNMshn2w7_1),.dout(w_dff_B_xTcMbHgz3_1),.clk(gclk));
	jdff dff_B_ZYclXlcM2_1(.din(w_dff_B_xTcMbHgz3_1),.dout(w_dff_B_ZYclXlcM2_1),.clk(gclk));
	jdff dff_B_RQkOQna85_1(.din(w_dff_B_ZYclXlcM2_1),.dout(w_dff_B_RQkOQna85_1),.clk(gclk));
	jdff dff_B_BkNagHHh6_1(.din(w_dff_B_RQkOQna85_1),.dout(w_dff_B_BkNagHHh6_1),.clk(gclk));
	jdff dff_B_iPp6XAEi3_0(.din(n1009),.dout(w_dff_B_iPp6XAEi3_0),.clk(gclk));
	jdff dff_B_duw1jA3D8_0(.din(w_dff_B_iPp6XAEi3_0),.dout(w_dff_B_duw1jA3D8_0),.clk(gclk));
	jdff dff_B_TLv5oiTp8_0(.din(w_dff_B_duw1jA3D8_0),.dout(w_dff_B_TLv5oiTp8_0),.clk(gclk));
	jdff dff_A_nWFur3Lc4_0(.dout(w_n1008_0[0]),.din(w_dff_A_nWFur3Lc4_0),.clk(gclk));
	jdff dff_A_zKfZMW4N9_0(.dout(w_dff_A_nWFur3Lc4_0),.din(w_dff_A_zKfZMW4N9_0),.clk(gclk));
	jdff dff_A_o6NPZiL11_0(.dout(w_dff_A_zKfZMW4N9_0),.din(w_dff_A_o6NPZiL11_0),.clk(gclk));
	jdff dff_A_XqgRxEJy4_0(.dout(w_dff_A_o6NPZiL11_0),.din(w_dff_A_XqgRxEJy4_0),.clk(gclk));
	jdff dff_B_3gV6bLg16_1(.din(n1002),.dout(w_dff_B_3gV6bLg16_1),.clk(gclk));
	jdff dff_A_c6ksV2It6_0(.dout(w_n1003_0[0]),.din(w_dff_A_c6ksV2It6_0),.clk(gclk));
	jdff dff_A_Tss7Uoax4_1(.dout(w_n1000_0[1]),.din(w_dff_A_Tss7Uoax4_1),.clk(gclk));
	jdff dff_A_lzsf9YNj2_1(.dout(w_n985_0[1]),.din(w_dff_A_lzsf9YNj2_1),.clk(gclk));
	jdff dff_B_Xus4ekrH4_2(.din(n985),.dout(w_dff_B_Xus4ekrH4_2),.clk(gclk));
	jdff dff_B_mvlVMQb49_0(.din(n963),.dout(w_dff_B_mvlVMQb49_0),.clk(gclk));
	jdff dff_B_pZ8lh82s2_0(.din(w_dff_B_mvlVMQb49_0),.dout(w_dff_B_pZ8lh82s2_0),.clk(gclk));
	jdff dff_B_CT3fc92M1_0(.din(w_dff_B_pZ8lh82s2_0),.dout(w_dff_B_CT3fc92M1_0),.clk(gclk));
	jdff dff_B_xd3cfJjR0_0(.din(w_dff_B_CT3fc92M1_0),.dout(w_dff_B_xd3cfJjR0_0),.clk(gclk));
	jdff dff_B_EmzoD31v6_0(.din(w_dff_B_xd3cfJjR0_0),.dout(w_dff_B_EmzoD31v6_0),.clk(gclk));
	jdff dff_B_nwKB96Tv8_0(.din(w_dff_B_EmzoD31v6_0),.dout(w_dff_B_nwKB96Tv8_0),.clk(gclk));
	jdff dff_B_HKXq822L7_1(.din(n959),.dout(w_dff_B_HKXq822L7_1),.clk(gclk));
	jdff dff_B_Lhoo9HH01_0(.din(n957),.dout(w_dff_B_Lhoo9HH01_0),.clk(gclk));
	jdff dff_B_F8nFENal5_0(.din(w_dff_B_Lhoo9HH01_0),.dout(w_dff_B_F8nFENal5_0),.clk(gclk));
	jdff dff_B_uu1JPCKy3_0(.din(w_dff_B_F8nFENal5_0),.dout(w_dff_B_uu1JPCKy3_0),.clk(gclk));
	jdff dff_B_1qaZhbnY0_0(.din(w_dff_B_uu1JPCKy3_0),.dout(w_dff_B_1qaZhbnY0_0),.clk(gclk));
	jdff dff_B_Z1wa6H460_0(.din(w_dff_B_1qaZhbnY0_0),.dout(w_dff_B_Z1wa6H460_0),.clk(gclk));
	jdff dff_B_JueNAneB1_0(.din(n956),.dout(w_dff_B_JueNAneB1_0),.clk(gclk));
	jdff dff_B_nd8RMhdZ1_0(.din(n941),.dout(w_dff_B_nd8RMhdZ1_0),.clk(gclk));
	jdff dff_B_7kP8I6Nv7_0(.din(w_dff_B_nd8RMhdZ1_0),.dout(w_dff_B_7kP8I6Nv7_0),.clk(gclk));
	jdff dff_B_HtoLOBwu0_0(.din(w_dff_B_7kP8I6Nv7_0),.dout(w_dff_B_HtoLOBwu0_0),.clk(gclk));
	jdff dff_B_p4w6oiXH2_0(.din(w_dff_B_HtoLOBwu0_0),.dout(w_dff_B_p4w6oiXH2_0),.clk(gclk));
	jdff dff_B_EAGu5l770_0(.din(w_dff_B_p4w6oiXH2_0),.dout(w_dff_B_EAGu5l770_0),.clk(gclk));
	jdff dff_B_funZwnL82_0(.din(n932),.dout(w_dff_B_funZwnL82_0),.clk(gclk));
	jdff dff_B_tSORCQTA6_0(.din(w_dff_B_funZwnL82_0),.dout(w_dff_B_tSORCQTA6_0),.clk(gclk));
	jdff dff_B_vpZpWSVG6_0(.din(w_dff_B_tSORCQTA6_0),.dout(w_dff_B_vpZpWSVG6_0),.clk(gclk));
	jdff dff_B_D3MvhOYV3_0(.din(w_dff_B_vpZpWSVG6_0),.dout(w_dff_B_D3MvhOYV3_0),.clk(gclk));
	jdff dff_B_DRHH5VbM8_0(.din(n922),.dout(w_dff_B_DRHH5VbM8_0),.clk(gclk));
	jdff dff_B_Y2y7A30A9_0(.din(w_dff_B_DRHH5VbM8_0),.dout(w_dff_B_Y2y7A30A9_0),.clk(gclk));
	jdff dff_B_vgFcF65u4_0(.din(w_dff_B_Y2y7A30A9_0),.dout(w_dff_B_vgFcF65u4_0),.clk(gclk));
	jdff dff_B_oCrv8doN3_1(.din(n889),.dout(w_dff_B_oCrv8doN3_1),.clk(gclk));
	jdff dff_B_RmpkDI601_1(.din(w_dff_B_oCrv8doN3_1),.dout(w_dff_B_RmpkDI601_1),.clk(gclk));
	jdff dff_B_DUUq7Zzj9_1(.din(w_dff_B_RmpkDI601_1),.dout(w_dff_B_DUUq7Zzj9_1),.clk(gclk));
	jdff dff_B_jXWBPfOv2_0(.din(n906),.dout(w_dff_B_jXWBPfOv2_0),.clk(gclk));
	jdff dff_B_Z1KLiv0J5_0(.din(w_dff_B_jXWBPfOv2_0),.dout(w_dff_B_Z1KLiv0J5_0),.clk(gclk));
	jdff dff_B_wzfHBs9Y7_0(.din(n897),.dout(w_dff_B_wzfHBs9Y7_0),.clk(gclk));
	jdff dff_B_BlvzTLvr5_0(.din(n896),.dout(w_dff_B_BlvzTLvr5_0),.clk(gclk));
	jdff dff_A_VkhTzqs80_0(.dout(w_G89_0[0]),.din(w_dff_A_VkhTzqs80_0),.clk(gclk));
	jdff dff_A_RAnhR2Ke5_0(.dout(w_n895_0[0]),.din(w_dff_A_RAnhR2Ke5_0),.clk(gclk));
	jdff dff_B_gEZBHIQa1_0(.din(n879),.dout(w_dff_B_gEZBHIQa1_0),.clk(gclk));
	jdff dff_B_XLgbErkX1_1(.din(n875),.dout(w_dff_B_XLgbErkX1_1),.clk(gclk));
	jdff dff_A_G2KgPMH80_1(.dout(w_n863_0[1]),.din(w_dff_A_G2KgPMH80_1),.clk(gclk));
	jdff dff_A_AEaRPL7B0_1(.dout(w_n856_0[1]),.din(w_dff_A_AEaRPL7B0_1),.clk(gclk));
	jdff dff_B_TlGkzb2R8_1(.din(n1347),.dout(w_dff_B_TlGkzb2R8_1),.clk(gclk));
	jdff dff_B_Q8Ztu0Pv0_1(.din(w_dff_B_TlGkzb2R8_1),.dout(w_dff_B_Q8Ztu0Pv0_1),.clk(gclk));
	jdff dff_B_ASG2Rf5Z3_1(.din(n1352),.dout(w_dff_B_ASG2Rf5Z3_1),.clk(gclk));
	jdff dff_B_ebtfvnBV1_1(.din(w_dff_B_ASG2Rf5Z3_1),.dout(w_dff_B_ebtfvnBV1_1),.clk(gclk));
	jdff dff_B_O7vbFofv9_1(.din(w_dff_B_ebtfvnBV1_1),.dout(w_dff_B_O7vbFofv9_1),.clk(gclk));
	jdff dff_B_xilKJ2bD4_1(.din(w_dff_B_O7vbFofv9_1),.dout(w_dff_B_xilKJ2bD4_1),.clk(gclk));
	jdff dff_B_wzUqhPo52_1(.din(w_dff_B_xilKJ2bD4_1),.dout(w_dff_B_wzUqhPo52_1),.clk(gclk));
	jdff dff_B_uJ1Livi89_1(.din(w_dff_B_wzUqhPo52_1),.dout(w_dff_B_uJ1Livi89_1),.clk(gclk));
	jdff dff_B_3b6CDBYm8_1(.din(w_dff_B_uJ1Livi89_1),.dout(w_dff_B_3b6CDBYm8_1),.clk(gclk));
	jdff dff_B_3lPQYY2G2_1(.din(w_dff_B_3b6CDBYm8_1),.dout(w_dff_B_3lPQYY2G2_1),.clk(gclk));
	jdff dff_B_ec7G6yed2_1(.din(w_dff_B_3lPQYY2G2_1),.dout(w_dff_B_ec7G6yed2_1),.clk(gclk));
	jdff dff_B_eolntUTj5_1(.din(w_dff_B_ec7G6yed2_1),.dout(w_dff_B_eolntUTj5_1),.clk(gclk));
	jdff dff_B_M9uQLkgk0_1(.din(w_dff_B_eolntUTj5_1),.dout(w_dff_B_M9uQLkgk0_1),.clk(gclk));
	jdff dff_B_jgexdI7w1_1(.din(w_dff_B_M9uQLkgk0_1),.dout(w_dff_B_jgexdI7w1_1),.clk(gclk));
	jdff dff_B_9JvjqUzm1_1(.din(w_dff_B_jgexdI7w1_1),.dout(w_dff_B_9JvjqUzm1_1),.clk(gclk));
	jdff dff_B_vvv6rMzV4_1(.din(w_dff_B_9JvjqUzm1_1),.dout(w_dff_B_vvv6rMzV4_1),.clk(gclk));
	jdff dff_B_Y04GqOKy9_1(.din(w_dff_B_vvv6rMzV4_1),.dout(w_dff_B_Y04GqOKy9_1),.clk(gclk));
	jdff dff_B_Z6wYFNCf8_1(.din(w_dff_B_Y04GqOKy9_1),.dout(w_dff_B_Z6wYFNCf8_1),.clk(gclk));
	jdff dff_B_mzBNgqCu9_1(.din(w_dff_B_Z6wYFNCf8_1),.dout(w_dff_B_mzBNgqCu9_1),.clk(gclk));
	jdff dff_B_ki0A4K324_1(.din(w_dff_B_mzBNgqCu9_1),.dout(w_dff_B_ki0A4K324_1),.clk(gclk));
	jdff dff_B_fjpEQ3Jo4_1(.din(w_dff_B_ki0A4K324_1),.dout(w_dff_B_fjpEQ3Jo4_1),.clk(gclk));
	jdff dff_B_qcZSPAcg4_1(.din(w_dff_B_fjpEQ3Jo4_1),.dout(w_dff_B_qcZSPAcg4_1),.clk(gclk));
	jdff dff_B_NzjvkRve8_1(.din(n1368),.dout(w_dff_B_NzjvkRve8_1),.clk(gclk));
	jdff dff_B_9m8w8OCT8_1(.din(w_dff_B_NzjvkRve8_1),.dout(w_dff_B_9m8w8OCT8_1),.clk(gclk));
	jdff dff_B_N7BvwqaP7_1(.din(w_dff_B_9m8w8OCT8_1),.dout(w_dff_B_N7BvwqaP7_1),.clk(gclk));
	jdff dff_B_L4ss8y1M3_1(.din(w_dff_B_N7BvwqaP7_1),.dout(w_dff_B_L4ss8y1M3_1),.clk(gclk));
	jdff dff_B_EPO0p1Pn7_1(.din(w_dff_B_L4ss8y1M3_1),.dout(w_dff_B_EPO0p1Pn7_1),.clk(gclk));
	jdff dff_B_D8ohgkie5_1(.din(w_dff_B_EPO0p1Pn7_1),.dout(w_dff_B_D8ohgkie5_1),.clk(gclk));
	jdff dff_B_aoyY9Iwj9_1(.din(w_dff_B_D8ohgkie5_1),.dout(w_dff_B_aoyY9Iwj9_1),.clk(gclk));
	jdff dff_B_DVk0kigS7_1(.din(w_dff_B_aoyY9Iwj9_1),.dout(w_dff_B_DVk0kigS7_1),.clk(gclk));
	jdff dff_B_ZozvfSql1_1(.din(w_dff_B_DVk0kigS7_1),.dout(w_dff_B_ZozvfSql1_1),.clk(gclk));
	jdff dff_B_iwN74MFK9_1(.din(w_dff_B_ZozvfSql1_1),.dout(w_dff_B_iwN74MFK9_1),.clk(gclk));
	jdff dff_B_CTYAs7z95_1(.din(w_dff_B_iwN74MFK9_1),.dout(w_dff_B_CTYAs7z95_1),.clk(gclk));
	jdff dff_B_vw8GA2Eg7_1(.din(w_dff_B_CTYAs7z95_1),.dout(w_dff_B_vw8GA2Eg7_1),.clk(gclk));
	jdff dff_B_OKTHmd9v8_1(.din(w_dff_B_vw8GA2Eg7_1),.dout(w_dff_B_OKTHmd9v8_1),.clk(gclk));
	jdff dff_B_lzn87cmm9_1(.din(w_dff_B_OKTHmd9v8_1),.dout(w_dff_B_lzn87cmm9_1),.clk(gclk));
	jdff dff_B_zxTxP1KQ0_1(.din(w_dff_B_lzn87cmm9_1),.dout(w_dff_B_zxTxP1KQ0_1),.clk(gclk));
	jdff dff_B_MzmrHBrI1_1(.din(w_dff_B_zxTxP1KQ0_1),.dout(w_dff_B_MzmrHBrI1_1),.clk(gclk));
	jdff dff_B_z8PSb0fK2_1(.din(w_dff_B_MzmrHBrI1_1),.dout(w_dff_B_z8PSb0fK2_1),.clk(gclk));
	jdff dff_B_dvejynQC0_1(.din(w_dff_B_z8PSb0fK2_1),.dout(w_dff_B_dvejynQC0_1),.clk(gclk));
	jdff dff_B_pUvmZt6c4_1(.din(w_dff_B_dvejynQC0_1),.dout(w_dff_B_pUvmZt6c4_1),.clk(gclk));
	jdff dff_B_rwaob1yQ1_1(.din(w_dff_B_pUvmZt6c4_1),.dout(w_dff_B_rwaob1yQ1_1),.clk(gclk));
	jdff dff_B_S3HLASqu6_1(.din(w_dff_B_rwaob1yQ1_1),.dout(w_dff_B_S3HLASqu6_1),.clk(gclk));
	jdff dff_B_pgbUEQQb9_1(.din(w_dff_B_S3HLASqu6_1),.dout(w_dff_B_pgbUEQQb9_1),.clk(gclk));
	jdff dff_B_O5C0QGcS7_1(.din(w_dff_B_pgbUEQQb9_1),.dout(w_dff_B_O5C0QGcS7_1),.clk(gclk));
	jdff dff_B_MqArCBY05_1(.din(w_dff_B_O5C0QGcS7_1),.dout(w_dff_B_MqArCBY05_1),.clk(gclk));
	jdff dff_B_MqfVkYW82_1(.din(w_dff_B_MqArCBY05_1),.dout(w_dff_B_MqfVkYW82_1),.clk(gclk));
	jdff dff_B_iJvWAqwt9_1(.din(w_dff_B_MqfVkYW82_1),.dout(w_dff_B_iJvWAqwt9_1),.clk(gclk));
	jdff dff_B_scPDfLPg7_1(.din(w_dff_B_iJvWAqwt9_1),.dout(w_dff_B_scPDfLPg7_1),.clk(gclk));
	jdff dff_B_OT03VlAw2_1(.din(w_dff_B_scPDfLPg7_1),.dout(w_dff_B_OT03VlAw2_1),.clk(gclk));
	jdff dff_B_zSoaRWf89_1(.din(w_dff_B_OT03VlAw2_1),.dout(w_dff_B_zSoaRWf89_1),.clk(gclk));
	jdff dff_B_Ii4PdT4b5_1(.din(w_dff_B_zSoaRWf89_1),.dout(w_dff_B_Ii4PdT4b5_1),.clk(gclk));
	jdff dff_B_TBzUmDJr7_1(.din(w_dff_B_Ii4PdT4b5_1),.dout(w_dff_B_TBzUmDJr7_1),.clk(gclk));
	jdff dff_B_EXIhrkNU4_1(.din(w_dff_B_TBzUmDJr7_1),.dout(w_dff_B_EXIhrkNU4_1),.clk(gclk));
	jdff dff_B_ThSv8kmx6_1(.din(w_dff_B_EXIhrkNU4_1),.dout(w_dff_B_ThSv8kmx6_1),.clk(gclk));
	jdff dff_B_8pYQJq272_2(.din(n1323),.dout(w_dff_B_8pYQJq272_2),.clk(gclk));
	jdff dff_B_YMbh9Iu96_2(.din(w_dff_B_8pYQJq272_2),.dout(w_dff_B_YMbh9Iu96_2),.clk(gclk));
	jdff dff_B_45it95Sr4_2(.din(w_dff_B_YMbh9Iu96_2),.dout(w_dff_B_45it95Sr4_2),.clk(gclk));
	jdff dff_B_yYsuVKir5_2(.din(w_dff_B_45it95Sr4_2),.dout(w_dff_B_yYsuVKir5_2),.clk(gclk));
	jdff dff_B_VaF2Ke1S9_2(.din(w_dff_B_yYsuVKir5_2),.dout(w_dff_B_VaF2Ke1S9_2),.clk(gclk));
	jdff dff_B_Pikv11Vr8_2(.din(w_dff_B_VaF2Ke1S9_2),.dout(w_dff_B_Pikv11Vr8_2),.clk(gclk));
	jdff dff_B_eAeKRf8c3_2(.din(w_dff_B_Pikv11Vr8_2),.dout(w_dff_B_eAeKRf8c3_2),.clk(gclk));
	jdff dff_B_VvI9QdN05_2(.din(w_dff_B_eAeKRf8c3_2),.dout(w_dff_B_VvI9QdN05_2),.clk(gclk));
	jdff dff_B_J8I8Ps9A3_2(.din(w_dff_B_VvI9QdN05_2),.dout(w_dff_B_J8I8Ps9A3_2),.clk(gclk));
	jdff dff_B_8gcKVKG65_2(.din(w_dff_B_J8I8Ps9A3_2),.dout(w_dff_B_8gcKVKG65_2),.clk(gclk));
	jdff dff_B_yIEjn4Pn5_2(.din(w_dff_B_8gcKVKG65_2),.dout(w_dff_B_yIEjn4Pn5_2),.clk(gclk));
	jdff dff_B_jcZbdmaF2_2(.din(w_dff_B_yIEjn4Pn5_2),.dout(w_dff_B_jcZbdmaF2_2),.clk(gclk));
	jdff dff_B_skB34im25_2(.din(w_dff_B_jcZbdmaF2_2),.dout(w_dff_B_skB34im25_2),.clk(gclk));
	jdff dff_B_KbuqKSM01_2(.din(w_dff_B_skB34im25_2),.dout(w_dff_B_KbuqKSM01_2),.clk(gclk));
	jdff dff_B_JNirCrmu0_2(.din(w_dff_B_KbuqKSM01_2),.dout(w_dff_B_JNirCrmu0_2),.clk(gclk));
	jdff dff_B_ylluQ5Kf2_2(.din(w_dff_B_JNirCrmu0_2),.dout(w_dff_B_ylluQ5Kf2_2),.clk(gclk));
	jdff dff_B_5e84sic98_2(.din(w_dff_B_ylluQ5Kf2_2),.dout(w_dff_B_5e84sic98_2),.clk(gclk));
	jdff dff_B_IjfXU1yO3_2(.din(w_dff_B_5e84sic98_2),.dout(w_dff_B_IjfXU1yO3_2),.clk(gclk));
	jdff dff_B_mhnhOjzv2_2(.din(w_dff_B_IjfXU1yO3_2),.dout(w_dff_B_mhnhOjzv2_2),.clk(gclk));
	jdff dff_B_5Oakuo148_2(.din(w_dff_B_mhnhOjzv2_2),.dout(w_dff_B_5Oakuo148_2),.clk(gclk));
	jdff dff_B_CCM2iDWJ7_2(.din(w_dff_B_5Oakuo148_2),.dout(w_dff_B_CCM2iDWJ7_2),.clk(gclk));
	jdff dff_B_7XyHSN1D7_2(.din(w_dff_B_CCM2iDWJ7_2),.dout(w_dff_B_7XyHSN1D7_2),.clk(gclk));
	jdff dff_B_MDSQJJpu9_2(.din(w_dff_B_7XyHSN1D7_2),.dout(w_dff_B_MDSQJJpu9_2),.clk(gclk));
	jdff dff_B_KuG2qXsX3_2(.din(w_dff_B_MDSQJJpu9_2),.dout(w_dff_B_KuG2qXsX3_2),.clk(gclk));
	jdff dff_B_pbgTkE6x3_2(.din(w_dff_B_KuG2qXsX3_2),.dout(w_dff_B_pbgTkE6x3_2),.clk(gclk));
	jdff dff_B_rTO6oFH15_2(.din(w_dff_B_pbgTkE6x3_2),.dout(w_dff_B_rTO6oFH15_2),.clk(gclk));
	jdff dff_B_U29MVMUq1_2(.din(w_dff_B_rTO6oFH15_2),.dout(w_dff_B_U29MVMUq1_2),.clk(gclk));
	jdff dff_B_0BnnNxp55_2(.din(w_dff_B_U29MVMUq1_2),.dout(w_dff_B_0BnnNxp55_2),.clk(gclk));
	jdff dff_B_Q4fjijCy2_2(.din(w_dff_B_0BnnNxp55_2),.dout(w_dff_B_Q4fjijCy2_2),.clk(gclk));
	jdff dff_B_1mZL0dUv3_2(.din(n1369),.dout(w_dff_B_1mZL0dUv3_2),.clk(gclk));
	jdff dff_B_DgRzcWjQ8_2(.din(w_dff_B_1mZL0dUv3_2),.dout(w_dff_B_DgRzcWjQ8_2),.clk(gclk));
	jdff dff_B_8Hf5oHJP8_2(.din(w_dff_B_DgRzcWjQ8_2),.dout(w_dff_B_8Hf5oHJP8_2),.clk(gclk));
	jdff dff_B_7jsBZXdH1_2(.din(w_dff_B_8Hf5oHJP8_2),.dout(w_dff_B_7jsBZXdH1_2),.clk(gclk));
	jdff dff_B_vKV2T5HU2_2(.din(w_dff_B_7jsBZXdH1_2),.dout(w_dff_B_vKV2T5HU2_2),.clk(gclk));
	jdff dff_B_P7c0iDiS3_2(.din(w_dff_B_vKV2T5HU2_2),.dout(w_dff_B_P7c0iDiS3_2),.clk(gclk));
	jdff dff_B_rfCKVihw4_2(.din(w_dff_B_P7c0iDiS3_2),.dout(w_dff_B_rfCKVihw4_2),.clk(gclk));
	jdff dff_B_Nl5YtmKF3_2(.din(w_dff_B_rfCKVihw4_2),.dout(w_dff_B_Nl5YtmKF3_2),.clk(gclk));
	jdff dff_B_m6VlBMTA1_2(.din(w_dff_B_Nl5YtmKF3_2),.dout(w_dff_B_m6VlBMTA1_2),.clk(gclk));
	jdff dff_B_yT0YB5Gr3_2(.din(w_dff_B_m6VlBMTA1_2),.dout(w_dff_B_yT0YB5Gr3_2),.clk(gclk));
	jdff dff_B_TpIjfnur2_2(.din(w_dff_B_yT0YB5Gr3_2),.dout(w_dff_B_TpIjfnur2_2),.clk(gclk));
	jdff dff_B_oVRGp3Sp6_2(.din(w_dff_B_TpIjfnur2_2),.dout(w_dff_B_oVRGp3Sp6_2),.clk(gclk));
	jdff dff_B_H3Kw4QSz6_2(.din(w_dff_B_oVRGp3Sp6_2),.dout(w_dff_B_H3Kw4QSz6_2),.clk(gclk));
	jdff dff_B_vbgj8Y442_2(.din(w_dff_B_H3Kw4QSz6_2),.dout(w_dff_B_vbgj8Y442_2),.clk(gclk));
	jdff dff_B_zoCGWlAW4_2(.din(w_dff_B_vbgj8Y442_2),.dout(w_dff_B_zoCGWlAW4_2),.clk(gclk));
	jdff dff_B_OBL6shLY8_2(.din(w_dff_B_zoCGWlAW4_2),.dout(w_dff_B_OBL6shLY8_2),.clk(gclk));
	jdff dff_B_QidyfkZl2_2(.din(w_dff_B_OBL6shLY8_2),.dout(w_dff_B_QidyfkZl2_2),.clk(gclk));
	jdff dff_B_Deppp6vs2_2(.din(w_dff_B_QidyfkZl2_2),.dout(w_dff_B_Deppp6vs2_2),.clk(gclk));
	jdff dff_B_jhV68JHR4_2(.din(w_dff_B_Deppp6vs2_2),.dout(w_dff_B_jhV68JHR4_2),.clk(gclk));
	jdff dff_B_39WsdQ8F9_2(.din(w_dff_B_jhV68JHR4_2),.dout(w_dff_B_39WsdQ8F9_2),.clk(gclk));
	jdff dff_B_b4yFNX0X3_2(.din(w_dff_B_39WsdQ8F9_2),.dout(w_dff_B_b4yFNX0X3_2),.clk(gclk));
	jdff dff_B_pLRVB3053_2(.din(w_dff_B_b4yFNX0X3_2),.dout(w_dff_B_pLRVB3053_2),.clk(gclk));
	jdff dff_B_qgVOwGVd2_2(.din(w_dff_B_pLRVB3053_2),.dout(w_dff_B_qgVOwGVd2_2),.clk(gclk));
	jdff dff_B_zHXr17j86_2(.din(w_dff_B_qgVOwGVd2_2),.dout(w_dff_B_zHXr17j86_2),.clk(gclk));
	jdff dff_B_i2F67teG0_2(.din(w_dff_B_zHXr17j86_2),.dout(w_dff_B_i2F67teG0_2),.clk(gclk));
	jdff dff_B_O0tNs1sG8_2(.din(w_dff_B_i2F67teG0_2),.dout(w_dff_B_O0tNs1sG8_2),.clk(gclk));
	jdff dff_B_WRdAaSLj6_2(.din(w_dff_B_O0tNs1sG8_2),.dout(w_dff_B_WRdAaSLj6_2),.clk(gclk));
	jdff dff_B_uth7opkF7_2(.din(w_dff_B_WRdAaSLj6_2),.dout(w_dff_B_uth7opkF7_2),.clk(gclk));
	jdff dff_B_HxE8CPM29_2(.din(w_dff_B_uth7opkF7_2),.dout(w_dff_B_HxE8CPM29_2),.clk(gclk));
	jdff dff_B_CRNLJUNR4_2(.din(w_dff_B_HxE8CPM29_2),.dout(w_dff_B_CRNLJUNR4_2),.clk(gclk));
	jdff dff_B_EqhbmTAQ8_2(.din(w_dff_B_CRNLJUNR4_2),.dout(w_dff_B_EqhbmTAQ8_2),.clk(gclk));
	jdff dff_B_uElOBBtR3_1(.din(n1377),.dout(w_dff_B_uElOBBtR3_1),.clk(gclk));
	jdff dff_B_tS23SFrS2_1(.din(w_dff_B_uElOBBtR3_1),.dout(w_dff_B_tS23SFrS2_1),.clk(gclk));
	jdff dff_B_yxjpoCoZ8_1(.din(n1378),.dout(w_dff_B_yxjpoCoZ8_1),.clk(gclk));
	jdff dff_B_Hf9LsCV74_1(.din(w_dff_B_yxjpoCoZ8_1),.dout(w_dff_B_Hf9LsCV74_1),.clk(gclk));
	jdff dff_B_CRQGqpHS3_1(.din(w_dff_B_Hf9LsCV74_1),.dout(w_dff_B_CRQGqpHS3_1),.clk(gclk));
	jdff dff_B_yW36kaxx7_1(.din(w_dff_B_CRQGqpHS3_1),.dout(w_dff_B_yW36kaxx7_1),.clk(gclk));
	jdff dff_B_UqoebJiW5_1(.din(w_dff_B_yW36kaxx7_1),.dout(w_dff_B_UqoebJiW5_1),.clk(gclk));
	jdff dff_B_BNnp8BfI5_1(.din(w_dff_B_UqoebJiW5_1),.dout(w_dff_B_BNnp8BfI5_1),.clk(gclk));
	jdff dff_B_pquUCSvW2_1(.din(w_dff_B_BNnp8BfI5_1),.dout(w_dff_B_pquUCSvW2_1),.clk(gclk));
	jdff dff_B_3IVVGFyI8_1(.din(w_dff_B_pquUCSvW2_1),.dout(w_dff_B_3IVVGFyI8_1),.clk(gclk));
	jdff dff_B_c1ijh12B7_0(.din(n1379),.dout(w_dff_B_c1ijh12B7_0),.clk(gclk));
	jdff dff_B_9MZ870eG6_0(.din(w_dff_B_c1ijh12B7_0),.dout(w_dff_B_9MZ870eG6_0),.clk(gclk));
	jdff dff_B_cOu8ZMnh0_0(.din(w_dff_B_9MZ870eG6_0),.dout(w_dff_B_cOu8ZMnh0_0),.clk(gclk));
	jdff dff_B_HOFjcere8_0(.din(w_dff_B_cOu8ZMnh0_0),.dout(w_dff_B_HOFjcere8_0),.clk(gclk));
	jdff dff_B_2K5IGgkt5_0(.din(w_dff_B_HOFjcere8_0),.dout(w_dff_B_2K5IGgkt5_0),.clk(gclk));
	jdff dff_B_OR3YWzNO8_0(.din(w_dff_B_2K5IGgkt5_0),.dout(w_dff_B_OR3YWzNO8_0),.clk(gclk));
	jdff dff_B_cmBMnGhB7_0(.din(w_dff_B_OR3YWzNO8_0),.dout(w_dff_B_cmBMnGhB7_0),.clk(gclk));
	jdff dff_B_I71mcKFI5_0(.din(n1177),.dout(w_dff_B_I71mcKFI5_0),.clk(gclk));
	jdff dff_B_1RmXZwGf4_0(.din(n1176),.dout(w_dff_B_1RmXZwGf4_0),.clk(gclk));
	jdff dff_B_5zLcyl1i2_0(.din(n1174),.dout(w_dff_B_5zLcyl1i2_0),.clk(gclk));
	jdff dff_B_OSNyLonq1_1(.din(n1171),.dout(w_dff_B_OSNyLonq1_1),.clk(gclk));
	jdff dff_B_3qIHyXp94_0(.din(n1166),.dout(w_dff_B_3qIHyXp94_0),.clk(gclk));
	jdff dff_B_faRuQwHF6_1(.din(n1153),.dout(w_dff_B_faRuQwHF6_1),.clk(gclk));
	jdff dff_B_Rfv0VYib5_1(.din(w_dff_B_faRuQwHF6_1),.dout(w_dff_B_Rfv0VYib5_1),.clk(gclk));
	jdff dff_B_OcEbHR1J6_1(.din(w_dff_B_Rfv0VYib5_1),.dout(w_dff_B_OcEbHR1J6_1),.clk(gclk));
	jdff dff_B_XmbktWK82_1(.din(w_dff_B_OcEbHR1J6_1),.dout(w_dff_B_XmbktWK82_1),.clk(gclk));
	jdff dff_B_FzkDygg79_1(.din(n1158),.dout(w_dff_B_FzkDygg79_1),.clk(gclk));
	jdff dff_B_L7PyJuBi0_0(.din(n1148),.dout(w_dff_B_L7PyJuBi0_0),.clk(gclk));
	jdff dff_B_OBgwpE531_0(.din(w_dff_B_L7PyJuBi0_0),.dout(w_dff_B_OBgwpE531_0),.clk(gclk));
	jdff dff_B_hnkeOZ9E8_0(.din(n1146),.dout(w_dff_B_hnkeOZ9E8_0),.clk(gclk));
	jdff dff_B_WoLNCHGJ7_0(.din(n1141),.dout(w_dff_B_WoLNCHGJ7_0),.clk(gclk));
	jdff dff_B_0tWcuBVx4_1(.din(n1135),.dout(w_dff_B_0tWcuBVx4_1),.clk(gclk));
	jdff dff_B_B1RoABjt7_0(.din(n1138),.dout(w_dff_B_B1RoABjt7_0),.clk(gclk));
	jdff dff_B_d49urWCg8_1(.din(n1136),.dout(w_dff_B_d49urWCg8_1),.clk(gclk));
	jdff dff_B_GoIcQ4gX1_1(.din(n1120),.dout(w_dff_B_GoIcQ4gX1_1),.clk(gclk));
	jdff dff_B_jlJHHk7H2_1(.din(n1121),.dout(w_dff_B_jlJHHk7H2_1),.clk(gclk));
	jdff dff_B_GzZMZkHb1_1(.din(w_dff_B_jlJHHk7H2_1),.dout(w_dff_B_GzZMZkHb1_1),.clk(gclk));
	jdff dff_B_eAJK5NMH4_0(.din(n1131),.dout(w_dff_B_eAJK5NMH4_0),.clk(gclk));
	jdff dff_B_0aYxZ4TB8_0(.din(w_dff_B_eAJK5NMH4_0),.dout(w_dff_B_0aYxZ4TB8_0),.clk(gclk));
	jdff dff_B_LOeSXeM65_0(.din(n1119),.dout(w_dff_B_LOeSXeM65_0),.clk(gclk));
	jdff dff_B_0hoj0HAF7_0(.din(n1303),.dout(w_dff_B_0hoj0HAF7_0),.clk(gclk));
	jdff dff_B_4vA8AQV10_1(.din(n1289),.dout(w_dff_B_4vA8AQV10_1),.clk(gclk));
	jdff dff_B_cfkoG1Vt8_1(.din(w_dff_B_4vA8AQV10_1),.dout(w_dff_B_cfkoG1Vt8_1),.clk(gclk));
	jdff dff_B_VN3Zm8r59_0(.din(n1301),.dout(w_dff_B_VN3Zm8r59_0),.clk(gclk));
	jdff dff_B_rrXjb51L9_0(.din(w_dff_B_VN3Zm8r59_0),.dout(w_dff_B_rrXjb51L9_0),.clk(gclk));
	jdff dff_B_RJRmwaaI4_0(.din(n816),.dout(w_dff_B_RJRmwaaI4_0),.clk(gclk));
	jdff dff_B_QrpMF2wn8_0(.din(n809),.dout(w_dff_B_QrpMF2wn8_0),.clk(gclk));
	jdff dff_B_yAVd0J5N4_0(.din(G174),.dout(w_dff_B_yAVd0J5N4_0),.clk(gclk));
	jdff dff_B_dzW4rya13_0(.din(G173),.dout(w_dff_B_dzW4rya13_0),.clk(gclk));
	jdff dff_B_m3XKlcFu2_0(.din(G176),.dout(w_dff_B_m3XKlcFu2_0),.clk(gclk));
	jdff dff_B_79UrQMsw7_0(.din(G175),.dout(w_dff_B_79UrQMsw7_0),.clk(gclk));
	jdff dff_B_DMptHjD75_0(.din(n802),.dout(w_dff_B_DMptHjD75_0),.clk(gclk));
	jdff dff_B_zHUjpYCt9_0(.din(G177),.dout(w_dff_B_zHUjpYCt9_0),.clk(gclk));
	jdff dff_A_qESbXHkL9_0(.dout(w_n373_3[0]),.din(w_dff_A_qESbXHkL9_0),.clk(gclk));
	jdff dff_B_xys7zFVf2_0(.din(n823),.dout(w_dff_B_xys7zFVf2_0),.clk(gclk));
	jdff dff_B_VXgU1qD85_1(.din(n1270),.dout(w_dff_B_VXgU1qD85_1),.clk(gclk));
	jdff dff_B_vQInOfKG2_1(.din(w_dff_B_VXgU1qD85_1),.dout(w_dff_B_vQInOfKG2_1),.clk(gclk));
	jdff dff_B_27Kqg1wR5_1(.din(w_dff_B_vQInOfKG2_1),.dout(w_dff_B_27Kqg1wR5_1),.clk(gclk));
	jdff dff_B_t2sPzaDQ7_1(.din(w_dff_B_27Kqg1wR5_1),.dout(w_dff_B_t2sPzaDQ7_1),.clk(gclk));
	jdff dff_B_Jjg7lsSH3_1(.din(n1275),.dout(w_dff_B_Jjg7lsSH3_1),.clk(gclk));
	jdff dff_A_7g4YtcYM3_0(.dout(w_n725_0[0]),.din(w_dff_A_7g4YtcYM3_0),.clk(gclk));
	jdff dff_A_IBrD16ts4_0(.dout(w_dff_A_7g4YtcYM3_0),.din(w_dff_A_IBrD16ts4_0),.clk(gclk));
	jdff dff_B_DIYmvKh25_0(.din(G167),.dout(w_dff_B_DIYmvKh25_0),.clk(gclk));
	jdff dff_A_ntrVif4o4_0(.dout(w_n719_0[0]),.din(w_dff_A_ntrVif4o4_0),.clk(gclk));
	jdff dff_A_3E42TCUS7_0(.dout(w_dff_A_ntrVif4o4_0),.din(w_dff_A_3E42TCUS7_0),.clk(gclk));
	jdff dff_B_hwMRptnW4_0(.din(G166),.dout(w_dff_B_hwMRptnW4_0),.clk(gclk));
	jdff dff_B_w0VPXIFy1_0(.din(G169),.dout(w_dff_B_w0VPXIFy1_0),.clk(gclk));
	jdff dff_A_KqBYPGeX1_2(.dout(w_n373_5[2]),.din(w_dff_A_KqBYPGeX1_2),.clk(gclk));
	jdff dff_B_9Rdq1LAr7_0(.din(G168),.dout(w_dff_B_9Rdq1LAr7_0),.clk(gclk));
	jdff dff_B_D0eYQcHv3_1(.din(G170),.dout(w_dff_B_D0eYQcHv3_1),.clk(gclk));
	jdff dff_B_xjXDcDOB3_1(.din(n1257),.dout(w_dff_B_xjXDcDOB3_1),.clk(gclk));
	jdff dff_B_LU0uSKLW4_0(.din(n850),.dout(w_dff_B_LU0uSKLW4_0),.clk(gclk));
	jdff dff_A_zDNHOQQv8_1(.dout(w_n845_0[1]),.din(w_dff_A_zDNHOQQv8_1),.clk(gclk));
	jdff dff_B_XImWSt9X0_0(.din(n844),.dout(w_dff_B_XImWSt9X0_0),.clk(gclk));
	jdff dff_B_s4LIctIT6_0(.din(n1259),.dout(w_dff_B_s4LIctIT6_0),.clk(gclk));
	jdff dff_B_NahVCNbJ8_0(.din(G115),.dout(w_dff_B_NahVCNbJ8_0),.clk(gclk));
	jdff dff_B_DKVgnHfT6_0(.din(n965),.dout(w_dff_B_DKVgnHfT6_0),.clk(gclk));
	jdff dff_B_ms9OW3LG2_0(.din(n979),.dout(w_dff_B_ms9OW3LG2_0),.clk(gclk));
	jdff dff_B_yv5Uv9zV8_0(.din(n972),.dout(w_dff_B_yv5Uv9zV8_0),.clk(gclk));
	jdff dff_B_MikmA2wz1_0(.din(n994),.dout(w_dff_B_MikmA2wz1_0),.clk(gclk));
	jdff dff_B_JsIfzC3e0_0(.din(n986),.dout(w_dff_B_JsIfzC3e0_0),.clk(gclk));
	jdff dff_B_V5tqYNKC5_0(.din(n865),.dout(w_dff_B_V5tqYNKC5_0),.clk(gclk));
	jdff dff_B_tSwZ6JNW4_0(.din(n857),.dout(w_dff_B_tSwZ6JNW4_0),.clk(gclk));
	jdff dff_B_fgoR0sKj5_0(.din(n1252),.dout(w_dff_B_fgoR0sKj5_0),.clk(gclk));
	jdff dff_B_v55vyGEp0_0(.din(n899),.dout(w_dff_B_v55vyGEp0_0),.clk(gclk));
	jdff dff_B_ljr0nkmZ3_0(.din(n890),.dout(w_dff_B_ljr0nkmZ3_0),.clk(gclk));
	jdff dff_B_qaOf45IT1_0(.din(n915),.dout(w_dff_B_qaOf45IT1_0),.clk(gclk));
	jdff dff_B_eOJ5LWf19_0(.din(n884),.dout(w_dff_B_eOJ5LWf19_0),.clk(gclk));
	jdff dff_B_y2n6IbNe1_0(.din(n1247),.dout(w_dff_B_y2n6IbNe1_0),.clk(gclk));
	jdff dff_B_7M8GAmf22_0(.din(n1245),.dout(w_dff_B_7M8GAmf22_0),.clk(gclk));
	jdff dff_B_7T05TSdV1_0(.din(G44),.dout(w_dff_B_7T05TSdV1_0),.clk(gclk));
	jdff dff_B_aXUeyR8z8_0(.din(n1243),.dout(w_dff_B_aXUeyR8z8_0),.clk(gclk));
	jdff dff_B_emtolqjk2_0(.din(n949),.dout(w_dff_B_emtolqjk2_0),.clk(gclk));
	jdff dff_B_YnrrQu3O9_0(.din(n943),.dout(w_dff_B_YnrrQu3O9_0),.clk(gclk));
	jdff dff_B_XkSaNPgG2_0(.din(n934),.dout(w_dff_B_XkSaNPgG2_0),.clk(gclk));
	jdff dff_A_DLyspXo41_0(.dout(w_n926_0[0]),.din(w_dff_A_DLyspXo41_0),.clk(gclk));
	jdff dff_B_uZxkjb4b3_0(.din(n925),.dout(w_dff_B_uZxkjb4b3_0),.clk(gclk));
	jdff dff_A_1UvK5pWl9_0(.dout(w_G414_0),.din(w_dff_A_1UvK5pWl9_0),.clk(gclk));
	jdff dff_B_mW1xUD1e1_1(.din(n1228),.dout(w_dff_B_mW1xUD1e1_1),.clk(gclk));
	jdff dff_B_OCSbmqRp2_1(.din(w_dff_B_mW1xUD1e1_1),.dout(w_dff_B_OCSbmqRp2_1),.clk(gclk));
	jdff dff_B_IVfu9r9O7_0(.din(n1236),.dout(w_dff_B_IVfu9r9O7_0),.clk(gclk));
	jdff dff_B_LRbrNLwJ6_0(.din(n1234),.dout(w_dff_B_LRbrNLwJ6_0),.clk(gclk));
	jdff dff_B_b4hPWs5V6_0(.din(n733),.dout(w_dff_B_b4hPWs5V6_0),.clk(gclk));
	jdff dff_B_6ARVs7Pz3_0(.din(n746),.dout(w_dff_B_6ARVs7Pz3_0),.clk(gclk));
	jdff dff_B_DPX5VXjw8_0(.din(n740),.dout(w_dff_B_DPX5VXjw8_0),.clk(gclk));
	jdff dff_B_aRJmjQrm7_0(.din(n728),.dout(w_dff_B_aRJmjQrm7_0),.clk(gclk));
	jdff dff_B_b9rs7CCj0_0(.din(n722),.dout(w_dff_B_b9rs7CCj0_0),.clk(gclk));
	jdff dff_A_izC37lvh5_0(.dout(w_G2204_0[0]),.din(w_dff_A_izC37lvh5_0),.clk(gclk));
	jdff dff_A_m8kotUJU7_2(.dout(w_G18_17[2]),.din(w_dff_A_m8kotUJU7_2),.clk(gclk));
	jdff dff_A_frr3oQK92_2(.dout(w_dff_A_m8kotUJU7_2),.din(w_dff_A_frr3oQK92_2),.clk(gclk));
	jdff dff_B_7CQ1qRfY7_1(.din(n1212),.dout(w_dff_B_7CQ1qRfY7_1),.clk(gclk));
	jdff dff_B_1nQ57FpA3_1(.din(n1213),.dout(w_dff_B_1nQ57FpA3_1),.clk(gclk));
	jdff dff_B_W4jNgWOn8_0(.din(n998),.dout(w_dff_B_W4jNgWOn8_0),.clk(gclk));
	jdff dff_A_UYOAdUYd4_0(.dout(w_G18_20[0]),.din(w_dff_A_UYOAdUYd4_0),.clk(gclk));
	jdff dff_B_xDZu6nOM6_0(.din(n990),.dout(w_dff_B_xDZu6nOM6_0),.clk(gclk));
	jdff dff_B_wC0aYQQN6_1(.din(n1214),.dout(w_dff_B_wC0aYQQN6_1),.clk(gclk));
	jdff dff_A_QYDi2JN64_1(.dout(w_n355_12[1]),.din(w_dff_A_QYDi2JN64_1),.clk(gclk));
	jdff dff_B_XtbsRcWL8_0(.din(n969),.dout(w_dff_B_XtbsRcWL8_0),.clk(gclk));
	jdff dff_B_p0CF3ola8_0(.din(n982),.dout(w_dff_B_p0CF3ola8_0),.clk(gclk));
	jdff dff_B_V6haeHWd2_0(.din(n976),.dout(w_dff_B_V6haeHWd2_0),.clk(gclk));
	jdff dff_B_nLQv1jO69_0(.din(n869),.dout(w_dff_B_nLQv1jO69_0),.clk(gclk));
	jdff dff_B_USso0eYK3_0(.din(n861),.dout(w_dff_B_USso0eYK3_0),.clk(gclk));
	jdff dff_B_bOdZZeZW2_0(.din(n853),.dout(w_dff_B_bOdZZeZW2_0),.clk(gclk));
	jdff dff_B_E6bjujDE2_0(.din(n847),.dout(w_dff_B_E6bjujDE2_0),.clk(gclk));
	jdff dff_B_LNa1SlTM1_1(.din(n1195),.dout(w_dff_B_LNa1SlTM1_1),.clk(gclk));
	jdff dff_A_6CCpYkzY5_0(.dout(w_n938_0[0]),.din(w_dff_A_6CCpYkzY5_0),.clk(gclk));
	jdff dff_B_89Ljj37K2_0(.din(n937),.dout(w_dff_B_89Ljj37K2_0),.clk(gclk));
	jdff dff_B_XrjS3DjW1_0(.din(n929),.dout(w_dff_B_XrjS3DjW1_0),.clk(gclk));
	jdff dff_A_WiualOEz8_0(.dout(w_n905_0[0]),.din(w_dff_A_WiualOEz8_0),.clk(gclk));
	jdff dff_B_ECjMh99R0_0(.din(n918),.dout(w_dff_B_ECjMh99R0_0),.clk(gclk));
	jdff dff_B_KjMdpMqY3_0(.din(n1198),.dout(w_dff_B_KjMdpMqY3_0),.clk(gclk));
	jdff dff_B_RMyClBpC5_0(.din(n887),.dout(w_dff_B_RMyClBpC5_0),.clk(gclk));
	jdff dff_B_rVfVfTqS2_0(.din(n902),.dout(w_dff_B_rVfVfTqS2_0),.clk(gclk));
	jdff dff_B_0KB6iv9g0_0(.din(n893),.dout(w_dff_B_0KB6iv9g0_0),.clk(gclk));
	jdff dff_B_n52irTqO9_0(.din(n952),.dout(w_dff_B_n52irTqO9_0),.clk(gclk));
	jdff dff_B_aZGGt5d13_0(.din(n946),.dout(w_dff_B_aZGGt5d13_0),.clk(gclk));
	jdff dff_B_xix0vYG33_0(.din(n1190),.dout(w_dff_B_xix0vYG33_0),.clk(gclk));
	jdff dff_B_7UccTtN25_0(.din(n763),.dout(w_dff_B_7UccTtN25_0),.clk(gclk));
	jdff dff_B_BLQwtI809_0(.din(n757),.dout(w_dff_B_BLQwtI809_0),.clk(gclk));
	jdff dff_B_jP0SD0ms6_0(.din(n819),.dout(w_dff_B_jP0SD0ms6_0),.clk(gclk));
	jdff dff_B_6C2O4IGp8_0(.din(n813),.dout(w_dff_B_6C2O4IGp8_0),.clk(gclk));
	jdff dff_B_cJHpgVha7_0(.din(n805),.dout(w_dff_B_cJHpgVha7_0),.clk(gclk));
	jdff dff_B_9QxBzGL67_0(.din(n799),.dout(w_dff_B_9QxBzGL67_0),.clk(gclk));
	jdff dff_B_NiDkIno62_0(.din(n1185),.dout(w_dff_B_NiDkIno62_0),.clk(gclk));
	jdff dff_B_Ol64LYX28_0(.din(n1183),.dout(w_dff_B_Ol64LYX28_0),.clk(gclk));
	jdff dff_B_pJwGi2Fx0_0(.din(n826),.dout(w_dff_B_pJwGi2Fx0_0),.clk(gclk));
	jdff dff_A_8zHwxbIv2_0(.dout(w_n780_0[0]),.din(w_dff_A_8zHwxbIv2_0),.clk(gclk));
	jdff dff_B_IEzZQimm6_0(.din(n779),.dout(w_dff_B_IEzZQimm6_0),.clk(gclk));
	jdff dff_B_Gu6ly2qK5_0(.din(n771),.dout(w_dff_B_Gu6ly2qK5_0),.clk(gclk));
	jdff dff_B_mqK82V5A0_3(.din(n715),.dout(w_dff_B_mqK82V5A0_3),.clk(gclk));
	jdff dff_B_wtxMmLdS3_3(.din(w_dff_B_mqK82V5A0_3),.dout(w_dff_B_wtxMmLdS3_3),.clk(gclk));
	jdff dff_B_glwqR3mg8_3(.din(w_dff_B_wtxMmLdS3_3),.dout(w_dff_B_glwqR3mg8_3),.clk(gclk));
	jdff dff_B_gDlJkdk08_3(.din(w_dff_B_glwqR3mg8_3),.dout(w_dff_B_gDlJkdk08_3),.clk(gclk));
	jdff dff_B_w2khVVI92_3(.din(w_dff_B_gDlJkdk08_3),.dout(w_dff_B_w2khVVI92_3),.clk(gclk));
	jdff dff_B_wjdCyHom4_3(.din(w_dff_B_w2khVVI92_3),.dout(w_dff_B_wjdCyHom4_3),.clk(gclk));
	jdff dff_B_fQo03E7Z0_3(.din(w_dff_B_wjdCyHom4_3),.dout(w_dff_B_fQo03E7Z0_3),.clk(gclk));
	jdff dff_B_3TTKgxND6_3(.din(w_dff_B_fQo03E7Z0_3),.dout(w_dff_B_3TTKgxND6_3),.clk(gclk));
	jdff dff_B_NZMT5rI36_3(.din(w_dff_B_3TTKgxND6_3),.dout(w_dff_B_NZMT5rI36_3),.clk(gclk));
	jdff dff_B_gfChancj5_3(.din(w_dff_B_NZMT5rI36_3),.dout(w_dff_B_gfChancj5_3),.clk(gclk));
	jdff dff_B_9Vcbey5X0_3(.din(w_dff_B_gfChancj5_3),.dout(w_dff_B_9Vcbey5X0_3),.clk(gclk));
	jdff dff_B_ZaKJrtyT2_3(.din(w_dff_B_9Vcbey5X0_3),.dout(w_dff_B_ZaKJrtyT2_3),.clk(gclk));
	jdff dff_B_Ms6c9Mpd4_3(.din(w_dff_B_ZaKJrtyT2_3),.dout(w_dff_B_Ms6c9Mpd4_3),.clk(gclk));
	jdff dff_B_RjQ30wm96_3(.din(w_dff_B_Ms6c9Mpd4_3),.dout(w_dff_B_RjQ30wm96_3),.clk(gclk));
	jdff dff_B_J1XDUVKt9_3(.din(w_dff_B_RjQ30wm96_3),.dout(w_dff_B_J1XDUVKt9_3),.clk(gclk));
	jdff dff_B_JehOWxDS7_3(.din(w_dff_B_J1XDUVKt9_3),.dout(w_dff_B_JehOWxDS7_3),.clk(gclk));
	jdff dff_B_ZOzfa1qW7_3(.din(w_dff_B_JehOWxDS7_3),.dout(w_dff_B_ZOzfa1qW7_3),.clk(gclk));
	jdff dff_B_VtjMCQ885_3(.din(w_dff_B_ZOzfa1qW7_3),.dout(w_dff_B_VtjMCQ885_3),.clk(gclk));
	jdff dff_B_gQ0MuVuL1_3(.din(w_dff_B_VtjMCQ885_3),.dout(w_dff_B_gQ0MuVuL1_3),.clk(gclk));
	jdff dff_B_V9cJFCcC3_3(.din(w_dff_B_gQ0MuVuL1_3),.dout(w_dff_B_V9cJFCcC3_3),.clk(gclk));
	jdff dff_B_1Fi2TARt0_3(.din(w_dff_B_V9cJFCcC3_3),.dout(w_dff_B_1Fi2TARt0_3),.clk(gclk));
	jdff dff_B_GckgrVIi4_3(.din(w_dff_B_1Fi2TARt0_3),.dout(w_dff_B_GckgrVIi4_3),.clk(gclk));
	jdff dff_B_EHKo0wt72_3(.din(w_dff_B_GckgrVIi4_3),.dout(w_dff_B_EHKo0wt72_3),.clk(gclk));
	jdff dff_B_ek1NjZSI8_3(.din(w_dff_B_EHKo0wt72_3),.dout(w_dff_B_ek1NjZSI8_3),.clk(gclk));
	jdff dff_B_kHfJAVQO1_3(.din(w_dff_B_ek1NjZSI8_3),.dout(w_dff_B_kHfJAVQO1_3),.clk(gclk));
	jdff dff_B_NZfRnSj54_3(.din(w_dff_B_kHfJAVQO1_3),.dout(w_dff_B_NZfRnSj54_3),.clk(gclk));
	jdff dff_B_n6fv7dQd7_3(.din(w_dff_B_NZfRnSj54_3),.dout(w_dff_B_n6fv7dQd7_3),.clk(gclk));
	jdff dff_B_mtwyelTu3_3(.din(w_dff_B_n6fv7dQd7_3),.dout(w_dff_B_mtwyelTu3_3),.clk(gclk));
	jdff dff_B_zDoaU84N9_3(.din(w_dff_B_mtwyelTu3_3),.dout(w_dff_B_zDoaU84N9_3),.clk(gclk));
	jdff dff_B_SBGlCL4L1_3(.din(w_dff_B_zDoaU84N9_3),.dout(w_dff_B_SBGlCL4L1_3),.clk(gclk));
	jdff dff_B_ZasoEgxn9_3(.din(w_dff_B_SBGlCL4L1_3),.dout(w_dff_B_ZasoEgxn9_3),.clk(gclk));
	jdff dff_B_d5C4eOE93_3(.din(w_dff_B_ZasoEgxn9_3),.dout(w_dff_B_d5C4eOE93_3),.clk(gclk));
	jdff dff_B_CCdq6dpQ9_3(.din(w_dff_B_d5C4eOE93_3),.dout(w_dff_B_CCdq6dpQ9_3),.clk(gclk));
	jdff dff_B_szjUyLJN5_3(.din(w_dff_B_CCdq6dpQ9_3),.dout(w_dff_B_szjUyLJN5_3),.clk(gclk));
	jdff dff_B_dHTH04tO0_0(.din(n714),.dout(w_dff_B_dHTH04tO0_0),.clk(gclk));
	jdff dff_B_DmaoDgws5_1(.din(n1394),.dout(w_dff_B_DmaoDgws5_1),.clk(gclk));
	jdff dff_B_30yG8BV70_1(.din(w_dff_B_DmaoDgws5_1),.dout(w_dff_B_30yG8BV70_1),.clk(gclk));
	jdff dff_B_3XibVL1S4_1(.din(w_dff_B_30yG8BV70_1),.dout(w_dff_B_3XibVL1S4_1),.clk(gclk));
	jdff dff_B_OGgz2ypa1_1(.din(w_dff_B_3XibVL1S4_1),.dout(w_dff_B_OGgz2ypa1_1),.clk(gclk));
	jdff dff_B_1VIWuLj67_1(.din(w_dff_B_OGgz2ypa1_1),.dout(w_dff_B_1VIWuLj67_1),.clk(gclk));
	jdff dff_B_OlBKJfqu5_1(.din(w_dff_B_1VIWuLj67_1),.dout(w_dff_B_OlBKJfqu5_1),.clk(gclk));
	jdff dff_B_5Pq49O0v9_1(.din(w_dff_B_OlBKJfqu5_1),.dout(w_dff_B_5Pq49O0v9_1),.clk(gclk));
	jdff dff_B_uTJXqnZl7_1(.din(w_dff_B_5Pq49O0v9_1),.dout(w_dff_B_uTJXqnZl7_1),.clk(gclk));
	jdff dff_B_Yi9paHfp6_1(.din(w_dff_B_uTJXqnZl7_1),.dout(w_dff_B_Yi9paHfp6_1),.clk(gclk));
	jdff dff_B_V9DTpW9O1_1(.din(w_dff_B_Yi9paHfp6_1),.dout(w_dff_B_V9DTpW9O1_1),.clk(gclk));
	jdff dff_B_p00NvwVE7_1(.din(w_dff_B_V9DTpW9O1_1),.dout(w_dff_B_p00NvwVE7_1),.clk(gclk));
	jdff dff_B_uLZz6l8T7_1(.din(w_dff_B_p00NvwVE7_1),.dout(w_dff_B_uLZz6l8T7_1),.clk(gclk));
	jdff dff_B_DHuRrOr86_1(.din(w_dff_B_uLZz6l8T7_1),.dout(w_dff_B_DHuRrOr86_1),.clk(gclk));
	jdff dff_B_TO8jfICl5_1(.din(w_dff_B_DHuRrOr86_1),.dout(w_dff_B_TO8jfICl5_1),.clk(gclk));
	jdff dff_B_LnQ2JwSt4_1(.din(w_dff_B_TO8jfICl5_1),.dout(w_dff_B_LnQ2JwSt4_1),.clk(gclk));
	jdff dff_B_nyPLHBkH6_1(.din(w_dff_B_LnQ2JwSt4_1),.dout(w_dff_B_nyPLHBkH6_1),.clk(gclk));
	jdff dff_B_WTuTZ1VK3_1(.din(w_dff_B_nyPLHBkH6_1),.dout(w_dff_B_WTuTZ1VK3_1),.clk(gclk));
	jdff dff_B_tykZTdNa8_1(.din(w_dff_B_WTuTZ1VK3_1),.dout(w_dff_B_tykZTdNa8_1),.clk(gclk));
	jdff dff_B_jv7ZM1Es7_1(.din(w_dff_B_tykZTdNa8_1),.dout(w_dff_B_jv7ZM1Es7_1),.clk(gclk));
	jdff dff_B_ZqqTC3111_1(.din(w_dff_B_jv7ZM1Es7_1),.dout(w_dff_B_ZqqTC3111_1),.clk(gclk));
	jdff dff_B_bZ6p0Aom4_1(.din(w_dff_B_ZqqTC3111_1),.dout(w_dff_B_bZ6p0Aom4_1),.clk(gclk));
	jdff dff_B_KwgvnGu60_1(.din(w_dff_B_bZ6p0Aom4_1),.dout(w_dff_B_KwgvnGu60_1),.clk(gclk));
	jdff dff_B_3rsUJrOM6_1(.din(w_dff_B_KwgvnGu60_1),.dout(w_dff_B_3rsUJrOM6_1),.clk(gclk));
	jdff dff_B_D5qV4Rt37_1(.din(w_dff_B_3rsUJrOM6_1),.dout(w_dff_B_D5qV4Rt37_1),.clk(gclk));
	jdff dff_B_2NXbjwEV1_1(.din(w_dff_B_D5qV4Rt37_1),.dout(w_dff_B_2NXbjwEV1_1),.clk(gclk));
	jdff dff_B_f42ZBbJr1_1(.din(w_dff_B_2NXbjwEV1_1),.dout(w_dff_B_f42ZBbJr1_1),.clk(gclk));
	jdff dff_B_9zhpym730_1(.din(w_dff_B_f42ZBbJr1_1),.dout(w_dff_B_9zhpym730_1),.clk(gclk));
	jdff dff_B_blCWD16m3_1(.din(w_dff_B_9zhpym730_1),.dout(w_dff_B_blCWD16m3_1),.clk(gclk));
	jdff dff_B_lvyyLC6r9_1(.din(w_dff_B_blCWD16m3_1),.dout(w_dff_B_lvyyLC6r9_1),.clk(gclk));
	jdff dff_B_1nnbtCHl1_1(.din(w_dff_B_lvyyLC6r9_1),.dout(w_dff_B_1nnbtCHl1_1),.clk(gclk));
	jdff dff_B_0ZOCEZBN8_1(.din(w_dff_B_1nnbtCHl1_1),.dout(w_dff_B_0ZOCEZBN8_1),.clk(gclk));
	jdff dff_B_gxOD9HZV4_1(.din(w_dff_B_0ZOCEZBN8_1),.dout(w_dff_B_gxOD9HZV4_1),.clk(gclk));
	jdff dff_B_iQfw0NuI9_1(.din(w_dff_B_gxOD9HZV4_1),.dout(w_dff_B_iQfw0NuI9_1),.clk(gclk));
	jdff dff_B_CBDC1UjX4_1(.din(w_dff_B_iQfw0NuI9_1),.dout(w_dff_B_CBDC1UjX4_1),.clk(gclk));
	jdff dff_A_q2N10pwF2_0(.dout(w_n713_0[0]),.din(w_dff_A_q2N10pwF2_0),.clk(gclk));
	jdff dff_A_7dQjV6FX7_0(.dout(w_dff_A_q2N10pwF2_0),.din(w_dff_A_7dQjV6FX7_0),.clk(gclk));
	jdff dff_A_9tvWxzFK6_0(.dout(w_dff_A_7dQjV6FX7_0),.din(w_dff_A_9tvWxzFK6_0),.clk(gclk));
	jdff dff_A_3UfxVOXQ3_0(.dout(w_dff_A_9tvWxzFK6_0),.din(w_dff_A_3UfxVOXQ3_0),.clk(gclk));
	jdff dff_A_H3nBd0GW2_0(.dout(w_dff_A_3UfxVOXQ3_0),.din(w_dff_A_H3nBd0GW2_0),.clk(gclk));
	jdff dff_A_s1PhLqMt0_0(.dout(w_dff_A_H3nBd0GW2_0),.din(w_dff_A_s1PhLqMt0_0),.clk(gclk));
	jdff dff_A_F8FekCd93_0(.dout(w_dff_A_s1PhLqMt0_0),.din(w_dff_A_F8FekCd93_0),.clk(gclk));
	jdff dff_A_egLKs2CI2_0(.dout(w_dff_A_F8FekCd93_0),.din(w_dff_A_egLKs2CI2_0),.clk(gclk));
	jdff dff_A_qM3wT2Px9_0(.dout(w_dff_A_egLKs2CI2_0),.din(w_dff_A_qM3wT2Px9_0),.clk(gclk));
	jdff dff_A_QfczoNKq7_0(.dout(w_dff_A_qM3wT2Px9_0),.din(w_dff_A_QfczoNKq7_0),.clk(gclk));
	jdff dff_A_2FtDRXID7_0(.dout(w_dff_A_QfczoNKq7_0),.din(w_dff_A_2FtDRXID7_0),.clk(gclk));
	jdff dff_A_7BRGPNsc5_0(.dout(w_dff_A_2FtDRXID7_0),.din(w_dff_A_7BRGPNsc5_0),.clk(gclk));
	jdff dff_A_G0qAYfci7_0(.dout(w_dff_A_7BRGPNsc5_0),.din(w_dff_A_G0qAYfci7_0),.clk(gclk));
	jdff dff_A_PFfIZ3qv7_0(.dout(w_dff_A_G0qAYfci7_0),.din(w_dff_A_PFfIZ3qv7_0),.clk(gclk));
	jdff dff_A_g9dEiv1b4_0(.dout(w_dff_A_PFfIZ3qv7_0),.din(w_dff_A_g9dEiv1b4_0),.clk(gclk));
	jdff dff_A_eP3SQm9B0_0(.dout(w_dff_A_g9dEiv1b4_0),.din(w_dff_A_eP3SQm9B0_0),.clk(gclk));
	jdff dff_A_TbXDGri54_0(.dout(w_dff_A_eP3SQm9B0_0),.din(w_dff_A_TbXDGri54_0),.clk(gclk));
	jdff dff_A_muDG5zJw4_0(.dout(w_dff_A_TbXDGri54_0),.din(w_dff_A_muDG5zJw4_0),.clk(gclk));
	jdff dff_A_XvIzNUqa4_0(.dout(w_dff_A_muDG5zJw4_0),.din(w_dff_A_XvIzNUqa4_0),.clk(gclk));
	jdff dff_A_D6QNu48D3_0(.dout(w_dff_A_XvIzNUqa4_0),.din(w_dff_A_D6QNu48D3_0),.clk(gclk));
	jdff dff_A_O5DWwDki5_0(.dout(w_dff_A_D6QNu48D3_0),.din(w_dff_A_O5DWwDki5_0),.clk(gclk));
	jdff dff_A_j6ndADna4_0(.dout(w_dff_A_O5DWwDki5_0),.din(w_dff_A_j6ndADna4_0),.clk(gclk));
	jdff dff_A_VMpfbThm6_0(.dout(w_dff_A_j6ndADna4_0),.din(w_dff_A_VMpfbThm6_0),.clk(gclk));
	jdff dff_A_teUtjFgE9_0(.dout(w_dff_A_VMpfbThm6_0),.din(w_dff_A_teUtjFgE9_0),.clk(gclk));
	jdff dff_A_6jwelbXS9_0(.dout(w_dff_A_teUtjFgE9_0),.din(w_dff_A_6jwelbXS9_0),.clk(gclk));
	jdff dff_A_5kExzYhZ0_0(.dout(w_dff_A_6jwelbXS9_0),.din(w_dff_A_5kExzYhZ0_0),.clk(gclk));
	jdff dff_A_dG7aaPpF8_0(.dout(w_dff_A_5kExzYhZ0_0),.din(w_dff_A_dG7aaPpF8_0),.clk(gclk));
	jdff dff_A_R1RA9pMz7_0(.dout(w_dff_A_dG7aaPpF8_0),.din(w_dff_A_R1RA9pMz7_0),.clk(gclk));
	jdff dff_A_lcqFBfw92_0(.dout(w_dff_A_R1RA9pMz7_0),.din(w_dff_A_lcqFBfw92_0),.clk(gclk));
	jdff dff_A_jqKepCQL4_0(.dout(w_dff_A_lcqFBfw92_0),.din(w_dff_A_jqKepCQL4_0),.clk(gclk));
	jdff dff_A_xp6NkX0r8_0(.dout(w_dff_A_jqKepCQL4_0),.din(w_dff_A_xp6NkX0r8_0),.clk(gclk));
	jdff dff_A_d1LKsnvV4_0(.dout(w_dff_A_xp6NkX0r8_0),.din(w_dff_A_d1LKsnvV4_0),.clk(gclk));
	jdff dff_A_Nq8HOIKa7_0(.dout(w_dff_A_d1LKsnvV4_0),.din(w_dff_A_Nq8HOIKa7_0),.clk(gclk));
	jdff dff_A_bTX9z9f33_0(.dout(w_G38_1[0]),.din(w_dff_A_bTX9z9f33_0),.clk(gclk));
	jdff dff_A_8FTKaedz4_1(.dout(w_G38_1[1]),.din(w_dff_A_8FTKaedz4_1),.clk(gclk));
	jdff dff_A_9ehyRf9E8_0(.dout(w_n370_0[0]),.din(w_dff_A_9ehyRf9E8_0),.clk(gclk));
	jdff dff_A_pwqs1dkK6_0(.dout(w_dff_A_9ehyRf9E8_0),.din(w_dff_A_pwqs1dkK6_0),.clk(gclk));
	jdff dff_A_njhFUcHG4_1(.dout(w_n370_0[1]),.din(w_dff_A_njhFUcHG4_1),.clk(gclk));
	jdff dff_A_mIsh5nKZ1_1(.dout(w_dff_A_njhFUcHG4_1),.din(w_dff_A_mIsh5nKZ1_1),.clk(gclk));
	jdff dff_B_ZU6tV9hk4_3(.din(n370),.dout(w_dff_B_ZU6tV9hk4_3),.clk(gclk));
	jdff dff_B_b2tLbgnK7_3(.din(w_dff_B_ZU6tV9hk4_3),.dout(w_dff_B_b2tLbgnK7_3),.clk(gclk));
	jdff dff_B_HLQVfAld4_3(.din(w_dff_B_b2tLbgnK7_3),.dout(w_dff_B_HLQVfAld4_3),.clk(gclk));
	jdff dff_B_HHiri41I1_3(.din(w_dff_B_HLQVfAld4_3),.dout(w_dff_B_HHiri41I1_3),.clk(gclk));
	jdff dff_B_Oh6wSpcm7_3(.din(w_dff_B_HHiri41I1_3),.dout(w_dff_B_Oh6wSpcm7_3),.clk(gclk));
	jdff dff_B_2cH0qWM34_3(.din(w_dff_B_Oh6wSpcm7_3),.dout(w_dff_B_2cH0qWM34_3),.clk(gclk));
	jdff dff_B_lDJ72o1Y7_3(.din(w_dff_B_2cH0qWM34_3),.dout(w_dff_B_lDJ72o1Y7_3),.clk(gclk));
	jdff dff_B_nSDZTnrN0_3(.din(w_dff_B_lDJ72o1Y7_3),.dout(w_dff_B_nSDZTnrN0_3),.clk(gclk));
	jdff dff_B_pQZv2jl38_3(.din(w_dff_B_nSDZTnrN0_3),.dout(w_dff_B_pQZv2jl38_3),.clk(gclk));
	jdff dff_B_EFnZsD9u6_3(.din(w_dff_B_pQZv2jl38_3),.dout(w_dff_B_EFnZsD9u6_3),.clk(gclk));
	jdff dff_B_kOYPSxsu0_3(.din(w_dff_B_EFnZsD9u6_3),.dout(w_dff_B_kOYPSxsu0_3),.clk(gclk));
	jdff dff_B_1KbbxszE4_3(.din(w_dff_B_kOYPSxsu0_3),.dout(w_dff_B_1KbbxszE4_3),.clk(gclk));
	jdff dff_B_24ZEiQPO2_3(.din(w_dff_B_1KbbxszE4_3),.dout(w_dff_B_24ZEiQPO2_3),.clk(gclk));
	jdff dff_B_mfW44h273_3(.din(w_dff_B_24ZEiQPO2_3),.dout(w_dff_B_mfW44h273_3),.clk(gclk));
	jdff dff_B_G63aBnyk4_3(.din(w_dff_B_mfW44h273_3),.dout(w_dff_B_G63aBnyk4_3),.clk(gclk));
	jdff dff_B_0ieYwiaR6_3(.din(w_dff_B_G63aBnyk4_3),.dout(w_dff_B_0ieYwiaR6_3),.clk(gclk));
	jdff dff_B_U6KM1CAw4_3(.din(w_dff_B_0ieYwiaR6_3),.dout(w_dff_B_U6KM1CAw4_3),.clk(gclk));
	jdff dff_B_A2IaMNhV9_3(.din(w_dff_B_U6KM1CAw4_3),.dout(w_dff_B_A2IaMNhV9_3),.clk(gclk));
	jdff dff_B_7h0BXQlo3_3(.din(w_dff_B_A2IaMNhV9_3),.dout(w_dff_B_7h0BXQlo3_3),.clk(gclk));
	jdff dff_B_ezhxHhaj2_3(.din(w_dff_B_7h0BXQlo3_3),.dout(w_dff_B_ezhxHhaj2_3),.clk(gclk));
	jdff dff_B_LFVQ22Rs9_3(.din(w_dff_B_ezhxHhaj2_3),.dout(w_dff_B_LFVQ22Rs9_3),.clk(gclk));
	jdff dff_B_A71FCdqi3_3(.din(w_dff_B_LFVQ22Rs9_3),.dout(w_dff_B_A71FCdqi3_3),.clk(gclk));
	jdff dff_B_igpqo0ga5_3(.din(w_dff_B_A71FCdqi3_3),.dout(w_dff_B_igpqo0ga5_3),.clk(gclk));
	jdff dff_B_VlldJtQx4_3(.din(w_dff_B_igpqo0ga5_3),.dout(w_dff_B_VlldJtQx4_3),.clk(gclk));
	jdff dff_B_2zhIbBKE7_3(.din(w_dff_B_VlldJtQx4_3),.dout(w_dff_B_2zhIbBKE7_3),.clk(gclk));
	jdff dff_B_L0VxVvAx3_3(.din(w_dff_B_2zhIbBKE7_3),.dout(w_dff_B_L0VxVvAx3_3),.clk(gclk));
	jdff dff_B_x0f5if7o1_3(.din(w_dff_B_L0VxVvAx3_3),.dout(w_dff_B_x0f5if7o1_3),.clk(gclk));
	jdff dff_B_tzYvNAlR7_3(.din(w_dff_B_x0f5if7o1_3),.dout(w_dff_B_tzYvNAlR7_3),.clk(gclk));
	jdff dff_B_I55Vq5pF0_3(.din(w_dff_B_tzYvNAlR7_3),.dout(w_dff_B_I55Vq5pF0_3),.clk(gclk));
	jdff dff_B_1vIWxpLO5_3(.din(w_dff_B_I55Vq5pF0_3),.dout(w_dff_B_1vIWxpLO5_3),.clk(gclk));
	jdff dff_B_JdA71qNN2_3(.din(w_dff_B_1vIWxpLO5_3),.dout(w_dff_B_JdA71qNN2_3),.clk(gclk));
	jdff dff_B_CQ4A5VLN4_3(.din(w_dff_B_JdA71qNN2_3),.dout(w_dff_B_CQ4A5VLN4_3),.clk(gclk));
	jdff dff_B_XV3MfLLv5_1(.din(n365),.dout(w_dff_B_XV3MfLLv5_1),.clk(gclk));
	jdff dff_A_IK4xxIxf6_2(.dout(w_n363_0[2]),.din(w_dff_A_IK4xxIxf6_2),.clk(gclk));
	jdff dff_B_xYNrf7is3_3(.din(n363),.dout(w_dff_B_xYNrf7is3_3),.clk(gclk));
	jdff dff_B_BXBFnrXY1_3(.din(w_dff_B_xYNrf7is3_3),.dout(w_dff_B_BXBFnrXY1_3),.clk(gclk));
	jdff dff_B_9Rqn8m6M7_3(.din(w_dff_B_BXBFnrXY1_3),.dout(w_dff_B_9Rqn8m6M7_3),.clk(gclk));
	jdff dff_B_JENYrdUh5_3(.din(w_dff_B_9Rqn8m6M7_3),.dout(w_dff_B_JENYrdUh5_3),.clk(gclk));
	jdff dff_B_w9mgrB452_3(.din(w_dff_B_JENYrdUh5_3),.dout(w_dff_B_w9mgrB452_3),.clk(gclk));
	jdff dff_B_OWfkJWGJ0_3(.din(w_dff_B_w9mgrB452_3),.dout(w_dff_B_OWfkJWGJ0_3),.clk(gclk));
	jdff dff_B_7ti0uLSR2_3(.din(w_dff_B_OWfkJWGJ0_3),.dout(w_dff_B_7ti0uLSR2_3),.clk(gclk));
	jdff dff_B_4iREe2qE0_3(.din(w_dff_B_7ti0uLSR2_3),.dout(w_dff_B_4iREe2qE0_3),.clk(gclk));
	jdff dff_B_VwsYQFrQ9_3(.din(w_dff_B_4iREe2qE0_3),.dout(w_dff_B_VwsYQFrQ9_3),.clk(gclk));
	jdff dff_B_SjaM4DmG8_3(.din(w_dff_B_VwsYQFrQ9_3),.dout(w_dff_B_SjaM4DmG8_3),.clk(gclk));
	jdff dff_B_lsV7hKWi3_3(.din(w_dff_B_SjaM4DmG8_3),.dout(w_dff_B_lsV7hKWi3_3),.clk(gclk));
	jdff dff_B_Ks4Iu0u74_3(.din(w_dff_B_lsV7hKWi3_3),.dout(w_dff_B_Ks4Iu0u74_3),.clk(gclk));
	jdff dff_B_IQakFRgW9_3(.din(w_dff_B_Ks4Iu0u74_3),.dout(w_dff_B_IQakFRgW9_3),.clk(gclk));
	jdff dff_B_8JLSYnvn7_3(.din(w_dff_B_IQakFRgW9_3),.dout(w_dff_B_8JLSYnvn7_3),.clk(gclk));
	jdff dff_B_kMDuHP7i0_3(.din(w_dff_B_8JLSYnvn7_3),.dout(w_dff_B_kMDuHP7i0_3),.clk(gclk));
	jdff dff_B_hty7O9MI2_3(.din(w_dff_B_kMDuHP7i0_3),.dout(w_dff_B_hty7O9MI2_3),.clk(gclk));
	jdff dff_B_PnJUayvo0_3(.din(w_dff_B_hty7O9MI2_3),.dout(w_dff_B_PnJUayvo0_3),.clk(gclk));
	jdff dff_B_QhQzerc22_3(.din(w_dff_B_PnJUayvo0_3),.dout(w_dff_B_QhQzerc22_3),.clk(gclk));
	jdff dff_B_Tks1g2cz1_3(.din(w_dff_B_QhQzerc22_3),.dout(w_dff_B_Tks1g2cz1_3),.clk(gclk));
	jdff dff_B_mxagUY3t3_3(.din(w_dff_B_Tks1g2cz1_3),.dout(w_dff_B_mxagUY3t3_3),.clk(gclk));
	jdff dff_B_fCeMwCYK0_3(.din(w_dff_B_mxagUY3t3_3),.dout(w_dff_B_fCeMwCYK0_3),.clk(gclk));
	jdff dff_B_2goDnZLM2_3(.din(w_dff_B_fCeMwCYK0_3),.dout(w_dff_B_2goDnZLM2_3),.clk(gclk));
	jdff dff_B_7ogavWEc8_3(.din(w_dff_B_2goDnZLM2_3),.dout(w_dff_B_7ogavWEc8_3),.clk(gclk));
	jdff dff_B_WgSmYDol3_3(.din(w_dff_B_7ogavWEc8_3),.dout(w_dff_B_WgSmYDol3_3),.clk(gclk));
	jdff dff_B_2w72tr4c5_3(.din(w_dff_B_WgSmYDol3_3),.dout(w_dff_B_2w72tr4c5_3),.clk(gclk));
	jdff dff_B_rZoPdTTN8_3(.din(w_dff_B_2w72tr4c5_3),.dout(w_dff_B_rZoPdTTN8_3),.clk(gclk));
	jdff dff_B_kRYUO83D3_3(.din(w_dff_B_rZoPdTTN8_3),.dout(w_dff_B_kRYUO83D3_3),.clk(gclk));
	jdff dff_B_pscKGlGo7_3(.din(w_dff_B_kRYUO83D3_3),.dout(w_dff_B_pscKGlGo7_3),.clk(gclk));
	jdff dff_B_AwBuAuDI2_3(.din(w_dff_B_pscKGlGo7_3),.dout(w_dff_B_AwBuAuDI2_3),.clk(gclk));
	jdff dff_B_wi1ZHICE9_3(.din(w_dff_B_AwBuAuDI2_3),.dout(w_dff_B_wi1ZHICE9_3),.clk(gclk));
	jdff dff_B_hbKJ8em88_3(.din(w_dff_B_wi1ZHICE9_3),.dout(w_dff_B_hbKJ8em88_3),.clk(gclk));
	jdff dff_B_qfDuvjXL3_3(.din(w_dff_B_hbKJ8em88_3),.dout(w_dff_B_qfDuvjXL3_3),.clk(gclk));
	jdff dff_B_i0IAEUFQ6_3(.din(w_dff_B_qfDuvjXL3_3),.dout(w_dff_B_i0IAEUFQ6_3),.clk(gclk));
	jdff dff_B_cbk2BWzk1_3(.din(w_dff_B_i0IAEUFQ6_3),.dout(w_dff_B_cbk2BWzk1_3),.clk(gclk));
	jdff dff_B_iwCZEiy92_1(.din(n1409),.dout(w_dff_B_iwCZEiy92_1),.clk(gclk));
	jdff dff_B_lwAhtTXJ6_1(.din(w_dff_B_iwCZEiy92_1),.dout(w_dff_B_lwAhtTXJ6_1),.clk(gclk));
	jdff dff_B_mvZEa8Yb1_1(.din(w_dff_B_lwAhtTXJ6_1),.dout(w_dff_B_mvZEa8Yb1_1),.clk(gclk));
	jdff dff_B_rNLNxwjw9_1(.din(w_dff_B_mvZEa8Yb1_1),.dout(w_dff_B_rNLNxwjw9_1),.clk(gclk));
	jdff dff_B_0RPQMNlp9_1(.din(w_dff_B_rNLNxwjw9_1),.dout(w_dff_B_0RPQMNlp9_1),.clk(gclk));
	jdff dff_B_ItB9DSYK4_1(.din(w_dff_B_0RPQMNlp9_1),.dout(w_dff_B_ItB9DSYK4_1),.clk(gclk));
	jdff dff_B_nY6fBif09_1(.din(w_dff_B_ItB9DSYK4_1),.dout(w_dff_B_nY6fBif09_1),.clk(gclk));
	jdff dff_B_CzZm3sKM5_0(.din(n1423),.dout(w_dff_B_CzZm3sKM5_0),.clk(gclk));
	jdff dff_B_IJqXK7xy4_0(.din(w_dff_B_CzZm3sKM5_0),.dout(w_dff_B_IJqXK7xy4_0),.clk(gclk));
	jdff dff_B_CQOPHmxj9_0(.din(w_dff_B_IJqXK7xy4_0),.dout(w_dff_B_CQOPHmxj9_0),.clk(gclk));
	jdff dff_B_U6uUJYMY4_0(.din(w_dff_B_CQOPHmxj9_0),.dout(w_dff_B_U6uUJYMY4_0),.clk(gclk));
	jdff dff_B_CjtaEvzf9_0(.din(w_dff_B_U6uUJYMY4_0),.dout(w_dff_B_CjtaEvzf9_0),.clk(gclk));
	jdff dff_B_YU0fqcTE2_0(.din(w_dff_B_CjtaEvzf9_0),.dout(w_dff_B_YU0fqcTE2_0),.clk(gclk));
	jdff dff_B_ITbNaMFb3_0(.din(w_dff_B_YU0fqcTE2_0),.dout(w_dff_B_ITbNaMFb3_0),.clk(gclk));
	jdff dff_B_CmeW8RsZ9_0(.din(w_dff_B_ITbNaMFb3_0),.dout(w_dff_B_CmeW8RsZ9_0),.clk(gclk));
	jdff dff_B_n5Wlgp9y2_0(.din(w_dff_B_CmeW8RsZ9_0),.dout(w_dff_B_n5Wlgp9y2_0),.clk(gclk));
	jdff dff_B_maMs4OPL4_0(.din(w_dff_B_n5Wlgp9y2_0),.dout(w_dff_B_maMs4OPL4_0),.clk(gclk));
	jdff dff_B_wWZT8jzU8_0(.din(w_dff_B_maMs4OPL4_0),.dout(w_dff_B_wWZT8jzU8_0),.clk(gclk));
	jdff dff_B_AulaXLNa1_0(.din(w_dff_B_wWZT8jzU8_0),.dout(w_dff_B_AulaXLNa1_0),.clk(gclk));
	jdff dff_B_ksX8i8EM9_0(.din(w_dff_B_AulaXLNa1_0),.dout(w_dff_B_ksX8i8EM9_0),.clk(gclk));
	jdff dff_B_5QgMdvmu0_0(.din(w_dff_B_ksX8i8EM9_0),.dout(w_dff_B_5QgMdvmu0_0),.clk(gclk));
	jdff dff_B_Kl87ZlXS5_0(.din(w_dff_B_5QgMdvmu0_0),.dout(w_dff_B_Kl87ZlXS5_0),.clk(gclk));
	jdff dff_B_njTeZRjP2_0(.din(w_dff_B_Kl87ZlXS5_0),.dout(w_dff_B_njTeZRjP2_0),.clk(gclk));
	jdff dff_B_heeQ53XN0_0(.din(n1478),.dout(w_dff_B_heeQ53XN0_0),.clk(gclk));
	jdff dff_B_2uSCymEX3_0(.din(w_dff_B_heeQ53XN0_0),.dout(w_dff_B_2uSCymEX3_0),.clk(gclk));
	jdff dff_B_Dlngj57s1_0(.din(n1477),.dout(w_dff_B_Dlngj57s1_0),.clk(gclk));
	jdff dff_B_jplcTCD69_0(.din(w_dff_B_Dlngj57s1_0),.dout(w_dff_B_jplcTCD69_0),.clk(gclk));
	jdff dff_B_JHL2yQWh1_0(.din(w_dff_B_jplcTCD69_0),.dout(w_dff_B_JHL2yQWh1_0),.clk(gclk));
	jdff dff_B_WStrZEZs9_0(.din(w_dff_B_JHL2yQWh1_0),.dout(w_dff_B_WStrZEZs9_0),.clk(gclk));
	jdff dff_B_gYFDldi45_0(.din(w_dff_B_WStrZEZs9_0),.dout(w_dff_B_gYFDldi45_0),.clk(gclk));
	jdff dff_B_0WgCKNXn7_0(.din(w_dff_B_gYFDldi45_0),.dout(w_dff_B_0WgCKNXn7_0),.clk(gclk));
	jdff dff_B_rTWBlQkd3_0(.din(w_dff_B_0WgCKNXn7_0),.dout(w_dff_B_rTWBlQkd3_0),.clk(gclk));
	jdff dff_B_rJHql58A8_0(.din(w_dff_B_rTWBlQkd3_0),.dout(w_dff_B_rJHql58A8_0),.clk(gclk));
	jdff dff_B_jzMC9Zpr9_0(.din(w_dff_B_rJHql58A8_0),.dout(w_dff_B_jzMC9Zpr9_0),.clk(gclk));
	jdff dff_B_NQhUAtfH7_0(.din(w_dff_B_jzMC9Zpr9_0),.dout(w_dff_B_NQhUAtfH7_0),.clk(gclk));
	jdff dff_B_jEpyes7S5_0(.din(w_dff_B_NQhUAtfH7_0),.dout(w_dff_B_jEpyes7S5_0),.clk(gclk));
	jdff dff_B_xtUd53kq0_0(.din(w_dff_B_jEpyes7S5_0),.dout(w_dff_B_xtUd53kq0_0),.clk(gclk));
	jdff dff_B_QKsJMYwe8_0(.din(w_dff_B_xtUd53kq0_0),.dout(w_dff_B_QKsJMYwe8_0),.clk(gclk));
	jdff dff_B_mN2iOQhY1_0(.din(w_dff_B_QKsJMYwe8_0),.dout(w_dff_B_mN2iOQhY1_0),.clk(gclk));
	jdff dff_B_ZIMfv6Ft0_0(.din(w_dff_B_mN2iOQhY1_0),.dout(w_dff_B_ZIMfv6Ft0_0),.clk(gclk));
	jdff dff_B_mQHKKZk18_0(.din(w_dff_B_ZIMfv6Ft0_0),.dout(w_dff_B_mQHKKZk18_0),.clk(gclk));
	jdff dff_B_KQMtYEJ24_0(.din(w_dff_B_mQHKKZk18_0),.dout(w_dff_B_KQMtYEJ24_0),.clk(gclk));
	jdff dff_B_voiF3B4n6_0(.din(w_dff_B_KQMtYEJ24_0),.dout(w_dff_B_voiF3B4n6_0),.clk(gclk));
	jdff dff_B_GZw9fVJM1_0(.din(w_dff_B_voiF3B4n6_0),.dout(w_dff_B_GZw9fVJM1_0),.clk(gclk));
	jdff dff_B_oBeFwSQN7_0(.din(w_dff_B_GZw9fVJM1_0),.dout(w_dff_B_oBeFwSQN7_0),.clk(gclk));
	jdff dff_B_3Bok2QBk2_0(.din(w_dff_B_oBeFwSQN7_0),.dout(w_dff_B_3Bok2QBk2_0),.clk(gclk));
	jdff dff_B_GwYFLE550_0(.din(w_dff_B_3Bok2QBk2_0),.dout(w_dff_B_GwYFLE550_0),.clk(gclk));
	jdff dff_B_YcQLb1wr8_0(.din(w_dff_B_GwYFLE550_0),.dout(w_dff_B_YcQLb1wr8_0),.clk(gclk));
	jdff dff_B_4e0S8qxo6_0(.din(w_dff_B_YcQLb1wr8_0),.dout(w_dff_B_4e0S8qxo6_0),.clk(gclk));
	jdff dff_B_entIfyXW2_0(.din(n1474),.dout(w_dff_B_entIfyXW2_0),.clk(gclk));
	jdff dff_B_8XGtxMwR9_0(.din(w_dff_B_entIfyXW2_0),.dout(w_dff_B_8XGtxMwR9_0),.clk(gclk));
	jdff dff_B_a0nVU4kh9_0(.din(w_dff_B_8XGtxMwR9_0),.dout(w_dff_B_a0nVU4kh9_0),.clk(gclk));
	jdff dff_B_QxABoxwe4_0(.din(w_dff_B_a0nVU4kh9_0),.dout(w_dff_B_QxABoxwe4_0),.clk(gclk));
	jdff dff_B_Ldyh76fx6_0(.din(w_dff_B_QxABoxwe4_0),.dout(w_dff_B_Ldyh76fx6_0),.clk(gclk));
	jdff dff_B_F4gtk9VZ6_0(.din(w_dff_B_Ldyh76fx6_0),.dout(w_dff_B_F4gtk9VZ6_0),.clk(gclk));
	jdff dff_B_Jr8WZMTC0_0(.din(w_dff_B_F4gtk9VZ6_0),.dout(w_dff_B_Jr8WZMTC0_0),.clk(gclk));
	jdff dff_B_hmSVbWko1_0(.din(w_dff_B_Jr8WZMTC0_0),.dout(w_dff_B_hmSVbWko1_0),.clk(gclk));
	jdff dff_B_5kx1C4oU1_0(.din(w_dff_B_hmSVbWko1_0),.dout(w_dff_B_5kx1C4oU1_0),.clk(gclk));
	jdff dff_B_ib85P0Do7_0(.din(w_dff_B_5kx1C4oU1_0),.dout(w_dff_B_ib85P0Do7_0),.clk(gclk));
	jdff dff_B_4iHWD0pp4_0(.din(w_dff_B_ib85P0Do7_0),.dout(w_dff_B_4iHWD0pp4_0),.clk(gclk));
	jdff dff_B_HRGL5uT05_0(.din(w_dff_B_4iHWD0pp4_0),.dout(w_dff_B_HRGL5uT05_0),.clk(gclk));
	jdff dff_B_4jen2nQk7_0(.din(w_dff_B_HRGL5uT05_0),.dout(w_dff_B_4jen2nQk7_0),.clk(gclk));
	jdff dff_B_dtd8IRAi8_0(.din(w_dff_B_4jen2nQk7_0),.dout(w_dff_B_dtd8IRAi8_0),.clk(gclk));
	jdff dff_B_9mp0lpax4_0(.din(w_dff_B_dtd8IRAi8_0),.dout(w_dff_B_9mp0lpax4_0),.clk(gclk));
	jdff dff_B_BhWBXVsX9_0(.din(n1473),.dout(w_dff_B_BhWBXVsX9_0),.clk(gclk));
	jdff dff_B_eN8HR6yF0_0(.din(n1469),.dout(w_dff_B_eN8HR6yF0_0),.clk(gclk));
	jdff dff_B_4aYXOa487_0(.din(n1465),.dout(w_dff_B_4aYXOa487_0),.clk(gclk));
	jdff dff_B_6OTOHNuf9_0(.din(w_dff_B_4aYXOa487_0),.dout(w_dff_B_6OTOHNuf9_0),.clk(gclk));
	jdff dff_B_fg5nQDsy0_0(.din(w_dff_B_6OTOHNuf9_0),.dout(w_dff_B_fg5nQDsy0_0),.clk(gclk));
	jdff dff_B_adcEbKvM5_0(.din(w_dff_B_fg5nQDsy0_0),.dout(w_dff_B_adcEbKvM5_0),.clk(gclk));
	jdff dff_B_jhGPRTPu7_0(.din(w_dff_B_adcEbKvM5_0),.dout(w_dff_B_jhGPRTPu7_0),.clk(gclk));
	jdff dff_B_cVQd0kbu9_0(.din(w_dff_B_jhGPRTPu7_0),.dout(w_dff_B_cVQd0kbu9_0),.clk(gclk));
	jdff dff_B_4junVqrn3_0(.din(w_dff_B_cVQd0kbu9_0),.dout(w_dff_B_4junVqrn3_0),.clk(gclk));
	jdff dff_B_HQvhTqdr8_0(.din(w_dff_B_4junVqrn3_0),.dout(w_dff_B_HQvhTqdr8_0),.clk(gclk));
	jdff dff_B_RDVU7uQd1_0(.din(w_dff_B_HQvhTqdr8_0),.dout(w_dff_B_RDVU7uQd1_0),.clk(gclk));
	jdff dff_B_rUyNkDps8_0(.din(w_dff_B_RDVU7uQd1_0),.dout(w_dff_B_rUyNkDps8_0),.clk(gclk));
	jdff dff_B_ifkGSxQ64_0(.din(w_dff_B_rUyNkDps8_0),.dout(w_dff_B_ifkGSxQ64_0),.clk(gclk));
	jdff dff_B_06H5CUu42_0(.din(w_dff_B_ifkGSxQ64_0),.dout(w_dff_B_06H5CUu42_0),.clk(gclk));
	jdff dff_B_KBTEMHY11_0(.din(w_dff_B_06H5CUu42_0),.dout(w_dff_B_KBTEMHY11_0),.clk(gclk));
	jdff dff_B_JQAzfofo1_1(.din(n1451),.dout(w_dff_B_JQAzfofo1_1),.clk(gclk));
	jdff dff_B_MzXGszdx7_0(.din(n1463),.dout(w_dff_B_MzXGszdx7_0),.clk(gclk));
	jdff dff_B_pZjI0ZAQ9_0(.din(w_dff_B_MzXGszdx7_0),.dout(w_dff_B_pZjI0ZAQ9_0),.clk(gclk));
	jdff dff_B_m0O3PEqb1_0(.din(w_dff_B_pZjI0ZAQ9_0),.dout(w_dff_B_m0O3PEqb1_0),.clk(gclk));
	jdff dff_B_wnS3s8PN9_0(.din(n1461),.dout(w_dff_B_wnS3s8PN9_0),.clk(gclk));
	jdff dff_B_zVPfz9jM0_1(.din(n1453),.dout(w_dff_B_zVPfz9jM0_1),.clk(gclk));
	jdff dff_B_LIpDOmxh0_1(.din(w_dff_B_zVPfz9jM0_1),.dout(w_dff_B_LIpDOmxh0_1),.clk(gclk));
	jdff dff_B_yNI3N9J80_0(.din(n1454),.dout(w_dff_B_yNI3N9J80_0),.clk(gclk));
	jdff dff_B_pBgev0qp1_0(.din(w_dff_B_yNI3N9J80_0),.dout(w_dff_B_pBgev0qp1_0),.clk(gclk));
	jdff dff_B_DBz0h19I2_0(.din(w_dff_B_pBgev0qp1_0),.dout(w_dff_B_DBz0h19I2_0),.clk(gclk));
	jdff dff_B_ykHznQu92_0(.din(w_dff_B_DBz0h19I2_0),.dout(w_dff_B_ykHznQu92_0),.clk(gclk));
	jdff dff_A_OPGzQBy28_0(.dout(w_n1452_0[0]),.din(w_dff_A_OPGzQBy28_0),.clk(gclk));
	jdff dff_A_sdWPMgqU9_0(.dout(w_dff_A_OPGzQBy28_0),.din(w_dff_A_sdWPMgqU9_0),.clk(gclk));
	jdff dff_A_ZAU6hFYu9_0(.dout(w_dff_A_sdWPMgqU9_0),.din(w_dff_A_ZAU6hFYu9_0),.clk(gclk));
	jdff dff_A_877u7CnR6_0(.dout(w_dff_A_ZAU6hFYu9_0),.din(w_dff_A_877u7CnR6_0),.clk(gclk));
	jdff dff_A_Kx8IwE3u5_2(.dout(w_n1452_0[2]),.din(w_dff_A_Kx8IwE3u5_2),.clk(gclk));
	jdff dff_A_Y4qbgTZr0_2(.dout(w_dff_A_Kx8IwE3u5_2),.din(w_dff_A_Y4qbgTZr0_2),.clk(gclk));
	jdff dff_A_WGaGkLAH1_2(.dout(w_dff_A_Y4qbgTZr0_2),.din(w_dff_A_WGaGkLAH1_2),.clk(gclk));
	jdff dff_A_AKv7wvjL7_1(.dout(w_n1340_0[1]),.din(w_dff_A_AKv7wvjL7_1),.clk(gclk));
	jdff dff_A_CzCbI9Ji8_2(.dout(w_n1340_0[2]),.din(w_dff_A_CzCbI9Ji8_2),.clk(gclk));
	jdff dff_A_qD5rT4n13_2(.dout(w_dff_A_CzCbI9Ji8_2),.din(w_dff_A_qD5rT4n13_2),.clk(gclk));
	jdff dff_A_D8tpZV5o0_2(.dout(w_dff_A_qD5rT4n13_2),.din(w_dff_A_D8tpZV5o0_2),.clk(gclk));
	jdff dff_A_3KaTgZGL4_2(.dout(w_dff_A_D8tpZV5o0_2),.din(w_dff_A_3KaTgZGL4_2),.clk(gclk));
	jdff dff_A_RAPm4VBC9_2(.dout(w_dff_A_3KaTgZGL4_2),.din(w_dff_A_RAPm4VBC9_2),.clk(gclk));
	jdff dff_A_yBzZvtQJ0_2(.dout(w_dff_A_RAPm4VBC9_2),.din(w_dff_A_yBzZvtQJ0_2),.clk(gclk));
	jdff dff_A_wGwfwR1B1_2(.dout(w_dff_A_yBzZvtQJ0_2),.din(w_dff_A_wGwfwR1B1_2),.clk(gclk));
	jdff dff_A_LuJYgc4V1_2(.dout(w_dff_A_wGwfwR1B1_2),.din(w_dff_A_LuJYgc4V1_2),.clk(gclk));
	jdff dff_A_X7GV8CaJ3_2(.dout(w_dff_A_LuJYgc4V1_2),.din(w_dff_A_X7GV8CaJ3_2),.clk(gclk));
	jdff dff_A_G3RKkQxr8_2(.dout(w_dff_A_X7GV8CaJ3_2),.din(w_dff_A_G3RKkQxr8_2),.clk(gclk));
	jdff dff_A_3niIIym51_2(.dout(w_dff_A_G3RKkQxr8_2),.din(w_dff_A_3niIIym51_2),.clk(gclk));
	jdff dff_A_Xsw30ZU44_2(.dout(w_dff_A_3niIIym51_2),.din(w_dff_A_Xsw30ZU44_2),.clk(gclk));
	jdff dff_A_X3eG48iL9_2(.dout(w_dff_A_Xsw30ZU44_2),.din(w_dff_A_X3eG48iL9_2),.clk(gclk));
	jdff dff_A_sVAdGYO23_2(.dout(w_dff_A_X3eG48iL9_2),.din(w_dff_A_sVAdGYO23_2),.clk(gclk));
	jdff dff_A_dapvPtw94_2(.dout(w_dff_A_sVAdGYO23_2),.din(w_dff_A_dapvPtw94_2),.clk(gclk));
	jdff dff_A_5PYuZQCK5_2(.dout(w_dff_A_dapvPtw94_2),.din(w_dff_A_5PYuZQCK5_2),.clk(gclk));
	jdff dff_A_zGzwXonD2_2(.dout(w_dff_A_5PYuZQCK5_2),.din(w_dff_A_zGzwXonD2_2),.clk(gclk));
	jdff dff_A_5JlJnPZS8_2(.dout(w_dff_A_zGzwXonD2_2),.din(w_dff_A_5JlJnPZS8_2),.clk(gclk));
	jdff dff_A_jZ4S0nXB2_2(.dout(w_dff_A_5JlJnPZS8_2),.din(w_dff_A_jZ4S0nXB2_2),.clk(gclk));
	jdff dff_A_ZzzLr51u8_2(.dout(w_dff_A_jZ4S0nXB2_2),.din(w_dff_A_ZzzLr51u8_2),.clk(gclk));
	jdff dff_A_uDXqbVQo7_2(.dout(w_dff_A_ZzzLr51u8_2),.din(w_dff_A_uDXqbVQo7_2),.clk(gclk));
	jdff dff_B_5FSA70jg8_3(.din(n1340),.dout(w_dff_B_5FSA70jg8_3),.clk(gclk));
	jdff dff_B_QY12PvqX4_3(.din(w_dff_B_5FSA70jg8_3),.dout(w_dff_B_QY12PvqX4_3),.clk(gclk));
	jdff dff_B_h8YYfvGs6_3(.din(w_dff_B_QY12PvqX4_3),.dout(w_dff_B_h8YYfvGs6_3),.clk(gclk));
	jdff dff_B_HCiw0wR69_0(.din(n1447),.dout(w_dff_B_HCiw0wR69_0),.clk(gclk));
	jdff dff_B_v9P2Ef6F8_0(.din(w_dff_B_HCiw0wR69_0),.dout(w_dff_B_v9P2Ef6F8_0),.clk(gclk));
	jdff dff_B_tDajx7HY7_0(.din(w_dff_B_v9P2Ef6F8_0),.dout(w_dff_B_tDajx7HY7_0),.clk(gclk));
	jdff dff_B_SdnNc85e9_0(.din(w_dff_B_tDajx7HY7_0),.dout(w_dff_B_SdnNc85e9_0),.clk(gclk));
	jdff dff_B_ZnjrzCG81_0(.din(w_dff_B_SdnNc85e9_0),.dout(w_dff_B_ZnjrzCG81_0),.clk(gclk));
	jdff dff_B_JGBqApfD5_0(.din(w_dff_B_ZnjrzCG81_0),.dout(w_dff_B_JGBqApfD5_0),.clk(gclk));
	jdff dff_B_hl2s3UDQ1_0(.din(w_dff_B_JGBqApfD5_0),.dout(w_dff_B_hl2s3UDQ1_0),.clk(gclk));
	jdff dff_B_poRSKr6K7_0(.din(w_dff_B_hl2s3UDQ1_0),.dout(w_dff_B_poRSKr6K7_0),.clk(gclk));
	jdff dff_B_wlYSBYug4_0(.din(w_dff_B_poRSKr6K7_0),.dout(w_dff_B_wlYSBYug4_0),.clk(gclk));
	jdff dff_B_Y8LRYdsQ7_0(.din(w_dff_B_wlYSBYug4_0),.dout(w_dff_B_Y8LRYdsQ7_0),.clk(gclk));
	jdff dff_B_YYdb0WtZ2_0(.din(w_dff_B_Y8LRYdsQ7_0),.dout(w_dff_B_YYdb0WtZ2_0),.clk(gclk));
	jdff dff_B_AfLOuRbE6_0(.din(w_dff_B_YYdb0WtZ2_0),.dout(w_dff_B_AfLOuRbE6_0),.clk(gclk));
	jdff dff_B_Guu9W5lT3_0(.din(w_dff_B_AfLOuRbE6_0),.dout(w_dff_B_Guu9W5lT3_0),.clk(gclk));
	jdff dff_B_Hh445aZ72_0(.din(w_dff_B_Guu9W5lT3_0),.dout(w_dff_B_Hh445aZ72_0),.clk(gclk));
	jdff dff_B_MNXvU4Yq5_0(.din(w_dff_B_Hh445aZ72_0),.dout(w_dff_B_MNXvU4Yq5_0),.clk(gclk));
	jdff dff_B_GCFSsGMy4_0(.din(w_dff_B_MNXvU4Yq5_0),.dout(w_dff_B_GCFSsGMy4_0),.clk(gclk));
	jdff dff_B_Oqzd83765_0(.din(w_dff_B_GCFSsGMy4_0),.dout(w_dff_B_Oqzd83765_0),.clk(gclk));
	jdff dff_B_YcZj1Ee59_0(.din(w_dff_B_Oqzd83765_0),.dout(w_dff_B_YcZj1Ee59_0),.clk(gclk));
	jdff dff_B_CYuVarN33_0(.din(w_dff_B_YcZj1Ee59_0),.dout(w_dff_B_CYuVarN33_0),.clk(gclk));
	jdff dff_B_19gLca623_1(.din(n1445),.dout(w_dff_B_19gLca623_1),.clk(gclk));
	jdff dff_B_oVKeCFhR0_0(.din(n1444),.dout(w_dff_B_oVKeCFhR0_0),.clk(gclk));
	jdff dff_B_p3iDl0LL3_0(.din(w_dff_B_oVKeCFhR0_0),.dout(w_dff_B_p3iDl0LL3_0),.clk(gclk));
	jdff dff_B_pA3M7hlw5_0(.din(n1441),.dout(w_dff_B_pA3M7hlw5_0),.clk(gclk));
	jdff dff_B_nXw0z1C79_0(.din(n1438),.dout(w_dff_B_nXw0z1C79_0),.clk(gclk));
	jdff dff_B_RmEVGv169_0(.din(w_dff_B_nXw0z1C79_0),.dout(w_dff_B_RmEVGv169_0),.clk(gclk));
	jdff dff_B_Q2TMaCkN0_0(.din(w_dff_B_RmEVGv169_0),.dout(w_dff_B_Q2TMaCkN0_0),.clk(gclk));
	jdff dff_B_ioWVW5cq5_0(.din(w_dff_B_Q2TMaCkN0_0),.dout(w_dff_B_ioWVW5cq5_0),.clk(gclk));
	jdff dff_B_zUMtOvXg5_0(.din(w_dff_B_ioWVW5cq5_0),.dout(w_dff_B_zUMtOvXg5_0),.clk(gclk));
	jdff dff_B_dTYmxbU09_0(.din(w_dff_B_zUMtOvXg5_0),.dout(w_dff_B_dTYmxbU09_0),.clk(gclk));
	jdff dff_B_m2bOGnqx5_0(.din(w_dff_B_dTYmxbU09_0),.dout(w_dff_B_m2bOGnqx5_0),.clk(gclk));
	jdff dff_B_vYd0JbmH8_0(.din(w_dff_B_m2bOGnqx5_0),.dout(w_dff_B_vYd0JbmH8_0),.clk(gclk));
	jdff dff_B_Exw3ZbQ40_0(.din(w_dff_B_vYd0JbmH8_0),.dout(w_dff_B_Exw3ZbQ40_0),.clk(gclk));
	jdff dff_B_bbqsGEX53_0(.din(w_dff_B_Exw3ZbQ40_0),.dout(w_dff_B_bbqsGEX53_0),.clk(gclk));
	jdff dff_B_dgleFurm4_0(.din(w_dff_B_bbqsGEX53_0),.dout(w_dff_B_dgleFurm4_0),.clk(gclk));
	jdff dff_B_HSpi26eR3_0(.din(w_dff_B_dgleFurm4_0),.dout(w_dff_B_HSpi26eR3_0),.clk(gclk));
	jdff dff_B_WPVgTrKh4_0(.din(w_dff_B_HSpi26eR3_0),.dout(w_dff_B_WPVgTrKh4_0),.clk(gclk));
	jdff dff_B_SliFyK364_0(.din(w_dff_B_WPVgTrKh4_0),.dout(w_dff_B_SliFyK364_0),.clk(gclk));
	jdff dff_B_DDPPv2SI4_0(.din(w_dff_B_SliFyK364_0),.dout(w_dff_B_DDPPv2SI4_0),.clk(gclk));
	jdff dff_B_a64E0SVz4_0(.din(w_dff_B_DDPPv2SI4_0),.dout(w_dff_B_a64E0SVz4_0),.clk(gclk));
	jdff dff_B_eBmcZyFn2_0(.din(w_dff_B_a64E0SVz4_0),.dout(w_dff_B_eBmcZyFn2_0),.clk(gclk));
	jdff dff_B_XqyKNomX4_0(.din(w_dff_B_eBmcZyFn2_0),.dout(w_dff_B_XqyKNomX4_0),.clk(gclk));
	jdff dff_B_vnvmDqhx9_0(.din(w_dff_B_XqyKNomX4_0),.dout(w_dff_B_vnvmDqhx9_0),.clk(gclk));
	jdff dff_B_JOn9JoTf0_0(.din(n1437),.dout(w_dff_B_JOn9JoTf0_0),.clk(gclk));
	jdff dff_B_OWbI6Hs37_1(.din(n1432),.dout(w_dff_B_OWbI6Hs37_1),.clk(gclk));
	jdff dff_A_zDaaqjFq9_1(.dout(w_n1388_0[1]),.din(w_dff_A_zDaaqjFq9_1),.clk(gclk));
	jdff dff_A_bIs27t4o1_1(.dout(w_dff_A_zDaaqjFq9_1),.din(w_dff_A_bIs27t4o1_1),.clk(gclk));
	jdff dff_A_jSGZbhrz3_1(.dout(w_dff_A_bIs27t4o1_1),.din(w_dff_A_jSGZbhrz3_1),.clk(gclk));
	jdff dff_A_igY0Jrt43_1(.dout(w_dff_A_jSGZbhrz3_1),.din(w_dff_A_igY0Jrt43_1),.clk(gclk));
	jdff dff_A_HZ0CV9l05_1(.dout(w_dff_A_igY0Jrt43_1),.din(w_dff_A_HZ0CV9l05_1),.clk(gclk));
	jdff dff_A_UQWJPadr1_1(.dout(w_dff_A_HZ0CV9l05_1),.din(w_dff_A_UQWJPadr1_1),.clk(gclk));
	jdff dff_A_Y6r6FIxN5_1(.dout(w_dff_A_UQWJPadr1_1),.din(w_dff_A_Y6r6FIxN5_1),.clk(gclk));
	jdff dff_A_px2Qhygn8_1(.dout(w_dff_A_Y6r6FIxN5_1),.din(w_dff_A_px2Qhygn8_1),.clk(gclk));
	jdff dff_A_ikDAEHbm8_1(.dout(w_dff_A_px2Qhygn8_1),.din(w_dff_A_ikDAEHbm8_1),.clk(gclk));
	jdff dff_A_HuNo3HCd3_1(.dout(w_dff_A_ikDAEHbm8_1),.din(w_dff_A_HuNo3HCd3_1),.clk(gclk));
	jdff dff_A_deX5kzSy0_1(.dout(w_dff_A_HuNo3HCd3_1),.din(w_dff_A_deX5kzSy0_1),.clk(gclk));
	jdff dff_A_xgkS52bQ8_1(.dout(w_dff_A_deX5kzSy0_1),.din(w_dff_A_xgkS52bQ8_1),.clk(gclk));
	jdff dff_A_sefBpE1U3_1(.dout(w_dff_A_xgkS52bQ8_1),.din(w_dff_A_sefBpE1U3_1),.clk(gclk));
	jdff dff_A_cC0Afoxr2_1(.dout(w_dff_A_sefBpE1U3_1),.din(w_dff_A_cC0Afoxr2_1),.clk(gclk));
	jdff dff_A_fJZpjdl66_1(.dout(w_dff_A_cC0Afoxr2_1),.din(w_dff_A_fJZpjdl66_1),.clk(gclk));
	jdff dff_A_Vm4uW51n2_1(.dout(w_dff_A_fJZpjdl66_1),.din(w_dff_A_Vm4uW51n2_1),.clk(gclk));
	jdff dff_A_Gr6F1muv4_1(.dout(w_dff_A_Vm4uW51n2_1),.din(w_dff_A_Gr6F1muv4_1),.clk(gclk));
	jdff dff_A_YlEPGzQx4_1(.dout(w_dff_A_Gr6F1muv4_1),.din(w_dff_A_YlEPGzQx4_1),.clk(gclk));
	jdff dff_A_9s3g67sC1_1(.dout(w_dff_A_YlEPGzQx4_1),.din(w_dff_A_9s3g67sC1_1),.clk(gclk));
	jdff dff_A_zxHTcwwh6_1(.dout(w_dff_A_9s3g67sC1_1),.din(w_dff_A_zxHTcwwh6_1),.clk(gclk));
	jdff dff_A_KjWqLPWo4_1(.dout(w_dff_A_zxHTcwwh6_1),.din(w_dff_A_KjWqLPWo4_1),.clk(gclk));
	jdff dff_A_rwnUHiRA0_1(.dout(w_dff_A_KjWqLPWo4_1),.din(w_dff_A_rwnUHiRA0_1),.clk(gclk));
	jdff dff_A_OdH2NJne7_1(.dout(w_dff_A_rwnUHiRA0_1),.din(w_dff_A_OdH2NJne7_1),.clk(gclk));
	jdff dff_A_8iBegAz22_1(.dout(w_dff_A_OdH2NJne7_1),.din(w_dff_A_8iBegAz22_1),.clk(gclk));
	jdff dff_A_3hTYa1n72_1(.dout(w_dff_A_8iBegAz22_1),.din(w_dff_A_3hTYa1n72_1),.clk(gclk));
	jdff dff_A_IBQBu9xf7_0(.dout(w_n1387_0[0]),.din(w_dff_A_IBQBu9xf7_0),.clk(gclk));
	jdff dff_A_1wkanVuV3_0(.dout(w_dff_A_IBQBu9xf7_0),.din(w_dff_A_1wkanVuV3_0),.clk(gclk));
	jdff dff_B_yp0UUsgy3_2(.din(n1431),.dout(w_dff_B_yp0UUsgy3_2),.clk(gclk));
	jdff dff_B_HhkjUhcZ3_2(.din(w_dff_B_yp0UUsgy3_2),.dout(w_dff_B_HhkjUhcZ3_2),.clk(gclk));
	jdff dff_B_REaPs5VA1_2(.din(w_dff_B_HhkjUhcZ3_2),.dout(w_dff_B_REaPs5VA1_2),.clk(gclk));
	jdff dff_B_bJorngyd9_2(.din(w_dff_B_REaPs5VA1_2),.dout(w_dff_B_bJorngyd9_2),.clk(gclk));
	jdff dff_B_M4dntbBX2_0(.din(n1526),.dout(w_dff_B_M4dntbBX2_0),.clk(gclk));
	jdff dff_B_Uh9VKXdS1_0(.din(n1524),.dout(w_dff_B_Uh9VKXdS1_0),.clk(gclk));
	jdff dff_B_LscSTxLd5_0(.din(w_dff_B_Uh9VKXdS1_0),.dout(w_dff_B_LscSTxLd5_0),.clk(gclk));
	jdff dff_B_gkVVzPnk3_0(.din(w_dff_B_LscSTxLd5_0),.dout(w_dff_B_gkVVzPnk3_0),.clk(gclk));
	jdff dff_B_vtGtHBCI9_0(.din(w_dff_B_gkVVzPnk3_0),.dout(w_dff_B_vtGtHBCI9_0),.clk(gclk));
	jdff dff_B_8BqA5M6p5_0(.din(w_dff_B_vtGtHBCI9_0),.dout(w_dff_B_8BqA5M6p5_0),.clk(gclk));
	jdff dff_B_js9pqa8p6_0(.din(w_dff_B_8BqA5M6p5_0),.dout(w_dff_B_js9pqa8p6_0),.clk(gclk));
	jdff dff_B_F4FwegUn5_0(.din(w_dff_B_js9pqa8p6_0),.dout(w_dff_B_F4FwegUn5_0),.clk(gclk));
	jdff dff_B_pYsChYHg4_0(.din(w_dff_B_F4FwegUn5_0),.dout(w_dff_B_pYsChYHg4_0),.clk(gclk));
	jdff dff_B_FpcoZgm93_0(.din(w_dff_B_pYsChYHg4_0),.dout(w_dff_B_FpcoZgm93_0),.clk(gclk));
	jdff dff_B_5UE2RiJF5_0(.din(w_dff_B_FpcoZgm93_0),.dout(w_dff_B_5UE2RiJF5_0),.clk(gclk));
	jdff dff_B_Rwj7kJJZ2_0(.din(w_dff_B_5UE2RiJF5_0),.dout(w_dff_B_Rwj7kJJZ2_0),.clk(gclk));
	jdff dff_B_hYHRqDqo2_0(.din(w_dff_B_Rwj7kJJZ2_0),.dout(w_dff_B_hYHRqDqo2_0),.clk(gclk));
	jdff dff_B_wVCtVCBj2_0(.din(w_dff_B_hYHRqDqo2_0),.dout(w_dff_B_wVCtVCBj2_0),.clk(gclk));
	jdff dff_B_kKCJNrL00_0(.din(w_dff_B_wVCtVCBj2_0),.dout(w_dff_B_kKCJNrL00_0),.clk(gclk));
	jdff dff_B_1pfcmRyW4_0(.din(w_dff_B_kKCJNrL00_0),.dout(w_dff_B_1pfcmRyW4_0),.clk(gclk));
	jdff dff_B_zCPKfWUA2_0(.din(w_dff_B_1pfcmRyW4_0),.dout(w_dff_B_zCPKfWUA2_0),.clk(gclk));
	jdff dff_B_PBm2BaFD9_0(.din(w_dff_B_zCPKfWUA2_0),.dout(w_dff_B_PBm2BaFD9_0),.clk(gclk));
	jdff dff_B_uU2xQCE56_0(.din(n1523),.dout(w_dff_B_uU2xQCE56_0),.clk(gclk));
	jdff dff_A_5gGzOLJl8_1(.dout(w_n420_0[1]),.din(w_dff_A_5gGzOLJl8_1),.clk(gclk));
	jdff dff_A_YmHdbC4Z9_1(.dout(w_dff_A_5gGzOLJl8_1),.din(w_dff_A_YmHdbC4Z9_1),.clk(gclk));
	jdff dff_A_b2PEHwBn9_1(.dout(w_dff_A_YmHdbC4Z9_1),.din(w_dff_A_b2PEHwBn9_1),.clk(gclk));
	jdff dff_A_4MNvW2gx6_1(.dout(w_dff_A_b2PEHwBn9_1),.din(w_dff_A_4MNvW2gx6_1),.clk(gclk));
	jdff dff_A_14FdSpXK1_1(.dout(w_dff_A_4MNvW2gx6_1),.din(w_dff_A_14FdSpXK1_1),.clk(gclk));
	jdff dff_A_4s24rNNu7_1(.dout(w_dff_A_14FdSpXK1_1),.din(w_dff_A_4s24rNNu7_1),.clk(gclk));
	jdff dff_A_XIhn4XGv7_1(.dout(w_dff_A_4s24rNNu7_1),.din(w_dff_A_XIhn4XGv7_1),.clk(gclk));
	jdff dff_A_zb1yipxd6_1(.dout(w_dff_A_XIhn4XGv7_1),.din(w_dff_A_zb1yipxd6_1),.clk(gclk));
	jdff dff_A_LfnEtyXp6_1(.dout(w_dff_A_zb1yipxd6_1),.din(w_dff_A_LfnEtyXp6_1),.clk(gclk));
	jdff dff_A_VHqQA4S40_1(.dout(w_dff_A_LfnEtyXp6_1),.din(w_dff_A_VHqQA4S40_1),.clk(gclk));
	jdff dff_A_2r4QNp145_1(.dout(w_dff_A_VHqQA4S40_1),.din(w_dff_A_2r4QNp145_1),.clk(gclk));
	jdff dff_A_Z0u7eusa9_1(.dout(w_dff_A_2r4QNp145_1),.din(w_dff_A_Z0u7eusa9_1),.clk(gclk));
	jdff dff_A_wBacaGYp0_1(.dout(w_dff_A_Z0u7eusa9_1),.din(w_dff_A_wBacaGYp0_1),.clk(gclk));
	jdff dff_A_sqLm0VZW5_1(.dout(w_dff_A_wBacaGYp0_1),.din(w_dff_A_sqLm0VZW5_1),.clk(gclk));
	jdff dff_A_GCDSgynG5_1(.dout(w_dff_A_sqLm0VZW5_1),.din(w_dff_A_GCDSgynG5_1),.clk(gclk));
	jdff dff_A_QjUPw4BJ8_1(.dout(w_dff_A_GCDSgynG5_1),.din(w_dff_A_QjUPw4BJ8_1),.clk(gclk));
	jdff dff_A_kvK8H9oF0_1(.dout(w_dff_A_QjUPw4BJ8_1),.din(w_dff_A_kvK8H9oF0_1),.clk(gclk));
	jdff dff_A_Ip0fJTsx9_1(.dout(w_dff_A_kvK8H9oF0_1),.din(w_dff_A_Ip0fJTsx9_1),.clk(gclk));
	jdff dff_A_4EbeUOuD3_1(.dout(w_dff_A_Ip0fJTsx9_1),.din(w_dff_A_4EbeUOuD3_1),.clk(gclk));
	jdff dff_A_HhEuQ8gq0_1(.dout(w_dff_A_4EbeUOuD3_1),.din(w_dff_A_HhEuQ8gq0_1),.clk(gclk));
	jdff dff_A_8rcwYPhX6_1(.dout(w_dff_A_HhEuQ8gq0_1),.din(w_dff_A_8rcwYPhX6_1),.clk(gclk));
	jdff dff_A_EfqEAZC60_0(.dout(w_n413_1[0]),.din(w_dff_A_EfqEAZC60_0),.clk(gclk));
	jdff dff_A_vPrYrtUM3_0(.dout(w_dff_A_EfqEAZC60_0),.din(w_dff_A_vPrYrtUM3_0),.clk(gclk));
	jdff dff_A_kFKHFjBJ0_0(.dout(w_dff_A_vPrYrtUM3_0),.din(w_dff_A_kFKHFjBJ0_0),.clk(gclk));
	jdff dff_A_MgolSiJF5_0(.dout(w_dff_A_kFKHFjBJ0_0),.din(w_dff_A_MgolSiJF5_0),.clk(gclk));
	jdff dff_A_z3DODmv08_0(.dout(w_dff_A_MgolSiJF5_0),.din(w_dff_A_z3DODmv08_0),.clk(gclk));
	jdff dff_A_Bu2R6wKw1_0(.dout(w_dff_A_z3DODmv08_0),.din(w_dff_A_Bu2R6wKw1_0),.clk(gclk));
	jdff dff_A_jHGQd42d4_0(.dout(w_dff_A_Bu2R6wKw1_0),.din(w_dff_A_jHGQd42d4_0),.clk(gclk));
	jdff dff_A_IOekg5D68_0(.dout(w_dff_A_jHGQd42d4_0),.din(w_dff_A_IOekg5D68_0),.clk(gclk));
	jdff dff_A_vnP7HZqA6_0(.dout(w_dff_A_IOekg5D68_0),.din(w_dff_A_vnP7HZqA6_0),.clk(gclk));
	jdff dff_A_RnAshcBa2_0(.dout(w_dff_A_vnP7HZqA6_0),.din(w_dff_A_RnAshcBa2_0),.clk(gclk));
	jdff dff_A_I9Yk1Ke74_0(.dout(w_dff_A_RnAshcBa2_0),.din(w_dff_A_I9Yk1Ke74_0),.clk(gclk));
	jdff dff_A_vsYzurLH9_0(.dout(w_dff_A_I9Yk1Ke74_0),.din(w_dff_A_vsYzurLH9_0),.clk(gclk));
	jdff dff_A_iXw4laOV6_0(.dout(w_dff_A_vsYzurLH9_0),.din(w_dff_A_iXw4laOV6_0),.clk(gclk));
	jdff dff_A_gwCZCdB63_0(.dout(w_dff_A_iXw4laOV6_0),.din(w_dff_A_gwCZCdB63_0),.clk(gclk));
	jdff dff_A_zF9GTniw8_0(.dout(w_dff_A_gwCZCdB63_0),.din(w_dff_A_zF9GTniw8_0),.clk(gclk));
	jdff dff_A_veFTmxyv3_0(.dout(w_dff_A_zF9GTniw8_0),.din(w_dff_A_veFTmxyv3_0),.clk(gclk));
	jdff dff_A_m1cyPN2n6_0(.dout(w_dff_A_veFTmxyv3_0),.din(w_dff_A_m1cyPN2n6_0),.clk(gclk));
	jdff dff_A_dUxSFAs18_0(.dout(w_dff_A_m1cyPN2n6_0),.din(w_dff_A_dUxSFAs18_0),.clk(gclk));
	jdff dff_A_FCcBznTD9_0(.dout(w_dff_A_dUxSFAs18_0),.din(w_dff_A_FCcBznTD9_0),.clk(gclk));
	jdff dff_A_OEP0ppCs1_0(.dout(w_dff_A_FCcBznTD9_0),.din(w_dff_A_OEP0ppCs1_0),.clk(gclk));
	jdff dff_A_MnDcgg263_0(.dout(w_dff_A_OEP0ppCs1_0),.din(w_dff_A_MnDcgg263_0),.clk(gclk));
	jdff dff_B_rg8UwGAd5_1(.din(n1521),.dout(w_dff_B_rg8UwGAd5_1),.clk(gclk));
	jdff dff_B_iQSqXYyW4_1(.din(w_dff_B_rg8UwGAd5_1),.dout(w_dff_B_iQSqXYyW4_1),.clk(gclk));
	jdff dff_B_ynPXtwQx8_1(.din(w_dff_B_iQSqXYyW4_1),.dout(w_dff_B_ynPXtwQx8_1),.clk(gclk));
	jdff dff_B_V1qUrEA61_1(.din(w_dff_B_ynPXtwQx8_1),.dout(w_dff_B_V1qUrEA61_1),.clk(gclk));
	jdff dff_B_CZwh5s0v2_1(.din(w_dff_B_V1qUrEA61_1),.dout(w_dff_B_CZwh5s0v2_1),.clk(gclk));
	jdff dff_B_v7OCEp2r2_1(.din(w_dff_B_CZwh5s0v2_1),.dout(w_dff_B_v7OCEp2r2_1),.clk(gclk));
	jdff dff_B_OTYgK7iz0_1(.din(w_dff_B_v7OCEp2r2_1),.dout(w_dff_B_OTYgK7iz0_1),.clk(gclk));
	jdff dff_A_D1dZChUW1_1(.dout(w_n419_0[1]),.din(w_dff_A_D1dZChUW1_1),.clk(gclk));
	jdff dff_A_Sz70AeEL0_1(.dout(w_dff_A_D1dZChUW1_1),.din(w_dff_A_Sz70AeEL0_1),.clk(gclk));
	jdff dff_A_YpLn6Q9P6_1(.dout(w_dff_A_Sz70AeEL0_1),.din(w_dff_A_YpLn6Q9P6_1),.clk(gclk));
	jdff dff_A_NoKSTi4d3_1(.dout(w_dff_A_YpLn6Q9P6_1),.din(w_dff_A_NoKSTi4d3_1),.clk(gclk));
	jdff dff_A_zMO4Xgwz1_1(.dout(w_dff_A_NoKSTi4d3_1),.din(w_dff_A_zMO4Xgwz1_1),.clk(gclk));
	jdff dff_A_KHAYfGor3_1(.dout(w_dff_A_zMO4Xgwz1_1),.din(w_dff_A_KHAYfGor3_1),.clk(gclk));
	jdff dff_B_IkFwriAd7_0(.din(n1519),.dout(w_dff_B_IkFwriAd7_0),.clk(gclk));
	jdff dff_B_9usL6MWy7_0(.din(w_dff_B_IkFwriAd7_0),.dout(w_dff_B_9usL6MWy7_0),.clk(gclk));
	jdff dff_B_HHDruGVr0_0(.din(w_dff_B_9usL6MWy7_0),.dout(w_dff_B_HHDruGVr0_0),.clk(gclk));
	jdff dff_B_WLMEmKxs3_0(.din(w_dff_B_HHDruGVr0_0),.dout(w_dff_B_WLMEmKxs3_0),.clk(gclk));
	jdff dff_B_XsDpzbJf8_0(.din(w_dff_B_WLMEmKxs3_0),.dout(w_dff_B_XsDpzbJf8_0),.clk(gclk));
	jdff dff_B_xi4K8tC28_0(.din(w_dff_B_XsDpzbJf8_0),.dout(w_dff_B_xi4K8tC28_0),.clk(gclk));
	jdff dff_B_sY5i52Hl1_0(.din(w_dff_B_xi4K8tC28_0),.dout(w_dff_B_sY5i52Hl1_0),.clk(gclk));
	jdff dff_B_joWPS9LO5_0(.din(w_dff_B_sY5i52Hl1_0),.dout(w_dff_B_joWPS9LO5_0),.clk(gclk));
	jdff dff_B_hY2aYXSu0_0(.din(w_dff_B_joWPS9LO5_0),.dout(w_dff_B_hY2aYXSu0_0),.clk(gclk));
	jdff dff_B_uqJpKo9i4_0(.din(w_dff_B_hY2aYXSu0_0),.dout(w_dff_B_uqJpKo9i4_0),.clk(gclk));
	jdff dff_B_NNmZswSL9_0(.din(w_dff_B_uqJpKo9i4_0),.dout(w_dff_B_NNmZswSL9_0),.clk(gclk));
	jdff dff_B_7OObS6FG5_0(.din(w_dff_B_NNmZswSL9_0),.dout(w_dff_B_7OObS6FG5_0),.clk(gclk));
	jdff dff_B_hBJ7awXS7_0(.din(w_dff_B_7OObS6FG5_0),.dout(w_dff_B_hBJ7awXS7_0),.clk(gclk));
	jdff dff_B_2INUkVPi7_0(.din(w_dff_B_hBJ7awXS7_0),.dout(w_dff_B_2INUkVPi7_0),.clk(gclk));
	jdff dff_B_BhkEQldm1_0(.din(w_dff_B_2INUkVPi7_0),.dout(w_dff_B_BhkEQldm1_0),.clk(gclk));
	jdff dff_B_aOla3Zsa1_0(.din(w_dff_B_BhkEQldm1_0),.dout(w_dff_B_aOla3Zsa1_0),.clk(gclk));
	jdff dff_B_ttYZu3Rs4_0(.din(w_dff_B_aOla3Zsa1_0),.dout(w_dff_B_ttYZu3Rs4_0),.clk(gclk));
	jdff dff_B_To1HMDCp2_0(.din(w_dff_B_ttYZu3Rs4_0),.dout(w_dff_B_To1HMDCp2_0),.clk(gclk));
	jdff dff_B_IiTdSLe73_1(.din(n1512),.dout(w_dff_B_IiTdSLe73_1),.clk(gclk));
	jdff dff_B_LAE2XKGt9_0(.din(n1517),.dout(w_dff_B_LAE2XKGt9_0),.clk(gclk));
	jdff dff_B_uytsovJ87_0(.din(w_dff_B_LAE2XKGt9_0),.dout(w_dff_B_uytsovJ87_0),.clk(gclk));
	jdff dff_B_ejmQ3Efr8_0(.din(w_dff_B_uytsovJ87_0),.dout(w_dff_B_ejmQ3Efr8_0),.clk(gclk));
	jdff dff_B_qP1Nuk7T4_0(.din(w_dff_B_ejmQ3Efr8_0),.dout(w_dff_B_qP1Nuk7T4_0),.clk(gclk));
	jdff dff_B_GdGqE3hQ0_0(.din(w_dff_B_qP1Nuk7T4_0),.dout(w_dff_B_GdGqE3hQ0_0),.clk(gclk));
	jdff dff_B_7sNWLq7L1_0(.din(w_dff_B_GdGqE3hQ0_0),.dout(w_dff_B_7sNWLq7L1_0),.clk(gclk));
	jdff dff_B_PdBQmugf1_0(.din(w_dff_B_7sNWLq7L1_0),.dout(w_dff_B_PdBQmugf1_0),.clk(gclk));
	jdff dff_B_qLIsIgXK4_0(.din(w_dff_B_PdBQmugf1_0),.dout(w_dff_B_qLIsIgXK4_0),.clk(gclk));
	jdff dff_B_p90kH7vl4_0(.din(w_dff_B_qLIsIgXK4_0),.dout(w_dff_B_p90kH7vl4_0),.clk(gclk));
	jdff dff_A_YDtMt7ws4_2(.dout(w_n366_0[2]),.din(w_dff_A_YDtMt7ws4_2),.clk(gclk));
	jdff dff_A_T1F6XDXd7_0(.dout(w_n361_0[0]),.din(w_dff_A_T1F6XDXd7_0),.clk(gclk));
	jdff dff_A_5Nhhcxai6_0(.dout(w_G38_2[0]),.din(w_dff_A_5Nhhcxai6_0),.clk(gclk));
	jdff dff_A_y9fJLhst5_0(.dout(w_dff_A_5Nhhcxai6_0),.din(w_dff_A_y9fJLhst5_0),.clk(gclk));
	jdff dff_A_ZAY3sdbH0_1(.dout(w_G38_2[1]),.din(w_dff_A_ZAY3sdbH0_1),.clk(gclk));
	jdff dff_A_stjFbjlk7_0(.dout(w_n1511_0[0]),.din(w_dff_A_stjFbjlk7_0),.clk(gclk));
	jdff dff_B_6cDj0TJ59_2(.din(n1511),.dout(w_dff_B_6cDj0TJ59_2),.clk(gclk));
	jdff dff_B_DdHJJIrb7_2(.din(w_dff_B_6cDj0TJ59_2),.dout(w_dff_B_DdHJJIrb7_2),.clk(gclk));
	jdff dff_B_2lLYqGG66_2(.din(w_dff_B_DdHJJIrb7_2),.dout(w_dff_B_2lLYqGG66_2),.clk(gclk));
	jdff dff_B_6DXf3yZk1_2(.din(w_dff_B_2lLYqGG66_2),.dout(w_dff_B_6DXf3yZk1_2),.clk(gclk));
	jdff dff_B_8QKTm6sM2_2(.din(w_dff_B_6DXf3yZk1_2),.dout(w_dff_B_8QKTm6sM2_2),.clk(gclk));
	jdff dff_B_FWWtzdEu6_2(.din(w_dff_B_8QKTm6sM2_2),.dout(w_dff_B_FWWtzdEu6_2),.clk(gclk));
	jdff dff_B_TW6PJP5p4_2(.din(w_dff_B_FWWtzdEu6_2),.dout(w_dff_B_TW6PJP5p4_2),.clk(gclk));
	jdff dff_B_zsXdLKoc7_2(.din(w_dff_B_TW6PJP5p4_2),.dout(w_dff_B_zsXdLKoc7_2),.clk(gclk));
	jdff dff_B_Eio5xOfu0_1(.din(n1508),.dout(w_dff_B_Eio5xOfu0_1),.clk(gclk));
	jdff dff_A_TS9rw5RI0_0(.dout(w_n364_0[0]),.din(w_dff_A_TS9rw5RI0_0),.clk(gclk));
	jdff dff_A_5c0RCyZl8_0(.dout(w_dff_A_TS9rw5RI0_0),.din(w_dff_A_5c0RCyZl8_0),.clk(gclk));
	jdff dff_A_1BRvXLhZ3_2(.dout(w_G1496_0[2]),.din(w_dff_A_1BRvXLhZ3_2),.clk(gclk));
	jdff dff_A_dHJt4ITd3_2(.dout(w_dff_A_1BRvXLhZ3_2),.din(w_dff_A_dHJt4ITd3_2),.clk(gclk));
	jdff dff_A_J3NkEjqI6_2(.dout(w_dff_A_dHJt4ITd3_2),.din(w_dff_A_J3NkEjqI6_2),.clk(gclk));
	jdff dff_A_mN4Y5ULW5_0(.dout(w_G1492_1[0]),.din(w_dff_A_mN4Y5ULW5_0),.clk(gclk));
	jdff dff_A_ryf5ao1F6_2(.dout(w_G1492_0[2]),.din(w_dff_A_ryf5ao1F6_2),.clk(gclk));
	jdff dff_A_tK7K9Fkw6_2(.dout(w_dff_A_ryf5ao1F6_2),.din(w_dff_A_tK7K9Fkw6_2),.clk(gclk));
	jdff dff_A_OMEH5hXN6_2(.dout(w_dff_A_tK7K9Fkw6_2),.din(w_dff_A_OMEH5hXN6_2),.clk(gclk));
	jdff dff_A_LQdGDyaf3_0(.dout(w_G38_0[0]),.din(w_dff_A_LQdGDyaf3_0),.clk(gclk));
	jdff dff_A_fc7Tr0NP2_2(.dout(w_G38_0[2]),.din(w_dff_A_fc7Tr0NP2_2),.clk(gclk));
	jdff dff_B_rRADiHUb3_1(.din(n376),.dout(w_dff_B_rRADiHUb3_1),.clk(gclk));
	jdff dff_B_TgN42e2d3_1(.din(w_dff_B_rRADiHUb3_1),.dout(w_dff_B_TgN42e2d3_1),.clk(gclk));
	jdff dff_B_yU4SBeVL3_1(.din(w_dff_B_TgN42e2d3_1),.dout(w_dff_B_yU4SBeVL3_1),.clk(gclk));
	jdff dff_B_Dor57Wdg2_1(.din(w_dff_B_yU4SBeVL3_1),.dout(w_dff_B_Dor57Wdg2_1),.clk(gclk));
	jdff dff_B_sSf5Vc6P5_1(.din(w_dff_B_Dor57Wdg2_1),.dout(w_dff_B_sSf5Vc6P5_1),.clk(gclk));
	jdff dff_B_65cDIrOJ4_1(.din(w_dff_B_sSf5Vc6P5_1),.dout(w_dff_B_65cDIrOJ4_1),.clk(gclk));
	jdff dff_B_rnc7HdhT9_1(.din(w_dff_B_65cDIrOJ4_1),.dout(w_dff_B_rnc7HdhT9_1),.clk(gclk));
	jdff dff_B_JlSU60wd0_1(.din(w_dff_B_rnc7HdhT9_1),.dout(w_dff_B_JlSU60wd0_1),.clk(gclk));
	jdff dff_A_vv1u85RS6_0(.dout(w_n377_1[0]),.din(w_dff_A_vv1u85RS6_0),.clk(gclk));
	jdff dff_A_I1sQzuSs6_0(.dout(w_dff_A_vv1u85RS6_0),.din(w_dff_A_I1sQzuSs6_0),.clk(gclk));
	jdff dff_A_ShlfCCAp3_0(.dout(w_dff_A_I1sQzuSs6_0),.din(w_dff_A_ShlfCCAp3_0),.clk(gclk));
	jdff dff_A_au2HequK3_0(.dout(w_dff_A_ShlfCCAp3_0),.din(w_dff_A_au2HequK3_0),.clk(gclk));
	jdff dff_A_XYNYSsfo3_0(.dout(w_dff_A_au2HequK3_0),.din(w_dff_A_XYNYSsfo3_0),.clk(gclk));
	jdff dff_A_lCo0J2P36_0(.dout(w_dff_A_XYNYSsfo3_0),.din(w_dff_A_lCo0J2P36_0),.clk(gclk));
	jdff dff_A_3VcDMBVU6_0(.dout(w_dff_A_lCo0J2P36_0),.din(w_dff_A_3VcDMBVU6_0),.clk(gclk));
	jdff dff_A_YkEiM8el4_0(.dout(w_dff_A_3VcDMBVU6_0),.din(w_dff_A_YkEiM8el4_0),.clk(gclk));
	jdff dff_A_zFoCX1fE6_0(.dout(w_dff_A_YkEiM8el4_0),.din(w_dff_A_zFoCX1fE6_0),.clk(gclk));
	jdff dff_A_lGEjnJqf7_0(.dout(w_dff_A_zFoCX1fE6_0),.din(w_dff_A_lGEjnJqf7_0),.clk(gclk));
	jdff dff_A_B4Uvi9wh0_0(.dout(w_dff_A_lGEjnJqf7_0),.din(w_dff_A_B4Uvi9wh0_0),.clk(gclk));
	jdff dff_A_WIvLSdsG7_0(.dout(w_dff_A_B4Uvi9wh0_0),.din(w_dff_A_WIvLSdsG7_0),.clk(gclk));
	jdff dff_A_86Hw0UjG9_0(.dout(w_dff_A_WIvLSdsG7_0),.din(w_dff_A_86Hw0UjG9_0),.clk(gclk));
	jdff dff_A_wCl0FIRY7_0(.dout(w_dff_A_86Hw0UjG9_0),.din(w_dff_A_wCl0FIRY7_0),.clk(gclk));
	jdff dff_A_1HXuwVzF8_0(.dout(w_dff_A_wCl0FIRY7_0),.din(w_dff_A_1HXuwVzF8_0),.clk(gclk));
	jdff dff_A_7w42ZpaP5_0(.dout(w_dff_A_1HXuwVzF8_0),.din(w_dff_A_7w42ZpaP5_0),.clk(gclk));
	jdff dff_A_XnA6JFnX3_0(.dout(w_dff_A_7w42ZpaP5_0),.din(w_dff_A_XnA6JFnX3_0),.clk(gclk));
	jdff dff_A_Ofx3yYQi7_0(.dout(w_dff_A_XnA6JFnX3_0),.din(w_dff_A_Ofx3yYQi7_0),.clk(gclk));
	jdff dff_A_XV5Ix2l99_0(.dout(w_dff_A_Ofx3yYQi7_0),.din(w_dff_A_XV5Ix2l99_0),.clk(gclk));
	jdff dff_A_o4RdDaLv8_0(.dout(w_dff_A_XV5Ix2l99_0),.din(w_dff_A_o4RdDaLv8_0),.clk(gclk));
	jdff dff_A_FqsXpHRE5_0(.dout(w_dff_A_o4RdDaLv8_0),.din(w_dff_A_FqsXpHRE5_0),.clk(gclk));
	jdff dff_A_4SfiI0QB4_0(.dout(w_dff_A_FqsXpHRE5_0),.din(w_dff_A_4SfiI0QB4_0),.clk(gclk));
	jdff dff_A_g8uNbSA76_0(.dout(w_dff_A_4SfiI0QB4_0),.din(w_dff_A_g8uNbSA76_0),.clk(gclk));
	jdff dff_A_tt9k7NbA3_0(.dout(w_dff_A_g8uNbSA76_0),.din(w_dff_A_tt9k7NbA3_0),.clk(gclk));
	jdff dff_A_sXSo4oBX0_0(.dout(w_dff_A_tt9k7NbA3_0),.din(w_dff_A_sXSo4oBX0_0),.clk(gclk));
	jdff dff_A_rFX5MMDq0_0(.dout(w_dff_A_sXSo4oBX0_0),.din(w_dff_A_rFX5MMDq0_0),.clk(gclk));
	jdff dff_A_O4x9BQG24_0(.dout(w_dff_A_rFX5MMDq0_0),.din(w_dff_A_O4x9BQG24_0),.clk(gclk));
	jdff dff_A_Bazhx6cq3_0(.dout(w_dff_A_O4x9BQG24_0),.din(w_dff_A_Bazhx6cq3_0),.clk(gclk));
	jdff dff_A_W95FR43n2_0(.dout(w_dff_A_Bazhx6cq3_0),.din(w_dff_A_W95FR43n2_0),.clk(gclk));
	jdff dff_A_f4rNf0jd1_0(.dout(w_dff_A_W95FR43n2_0),.din(w_dff_A_f4rNf0jd1_0),.clk(gclk));
	jdff dff_A_uH96gR3q6_2(.dout(w_n377_1[2]),.din(w_dff_A_uH96gR3q6_2),.clk(gclk));
	jdff dff_A_BqSshFE30_2(.dout(w_dff_A_uH96gR3q6_2),.din(w_dff_A_BqSshFE30_2),.clk(gclk));
	jdff dff_A_73TXpqed6_2(.dout(w_dff_A_BqSshFE30_2),.din(w_dff_A_73TXpqed6_2),.clk(gclk));
	jdff dff_A_GpE9zX9c1_2(.dout(w_dff_A_73TXpqed6_2),.din(w_dff_A_GpE9zX9c1_2),.clk(gclk));
	jdff dff_A_Cek6xykY5_2(.dout(w_dff_A_GpE9zX9c1_2),.din(w_dff_A_Cek6xykY5_2),.clk(gclk));
	jdff dff_B_KbplI2i71_1(.din(n1480),.dout(w_dff_B_KbplI2i71_1),.clk(gclk));
	jdff dff_B_8DgCpoAW7_1(.din(w_dff_B_KbplI2i71_1),.dout(w_dff_B_8DgCpoAW7_1),.clk(gclk));
	jdff dff_B_zR2UjtQK0_1(.din(w_dff_B_8DgCpoAW7_1),.dout(w_dff_B_zR2UjtQK0_1),.clk(gclk));
	jdff dff_B_oHTIevSM9_1(.din(w_dff_B_zR2UjtQK0_1),.dout(w_dff_B_oHTIevSM9_1),.clk(gclk));
	jdff dff_B_mcCwunEQ9_1(.din(w_dff_B_oHTIevSM9_1),.dout(w_dff_B_mcCwunEQ9_1),.clk(gclk));
	jdff dff_B_9OZxQn1N4_1(.din(w_dff_B_mcCwunEQ9_1),.dout(w_dff_B_9OZxQn1N4_1),.clk(gclk));
	jdff dff_B_AK0tmjSl2_1(.din(w_dff_B_9OZxQn1N4_1),.dout(w_dff_B_AK0tmjSl2_1),.clk(gclk));
	jdff dff_B_MHuP8Hc85_1(.din(w_dff_B_AK0tmjSl2_1),.dout(w_dff_B_MHuP8Hc85_1),.clk(gclk));
	jdff dff_B_SGl2lSaj0_1(.din(w_dff_B_MHuP8Hc85_1),.dout(w_dff_B_SGl2lSaj0_1),.clk(gclk));
	jdff dff_B_6E6gNwgW2_1(.din(w_dff_B_SGl2lSaj0_1),.dout(w_dff_B_6E6gNwgW2_1),.clk(gclk));
	jdff dff_B_3psTi4QW0_1(.din(w_dff_B_6E6gNwgW2_1),.dout(w_dff_B_3psTi4QW0_1),.clk(gclk));
	jdff dff_B_RIBcg9Vm5_1(.din(w_dff_B_3psTi4QW0_1),.dout(w_dff_B_RIBcg9Vm5_1),.clk(gclk));
	jdff dff_B_pvs0lKTW6_1(.din(w_dff_B_RIBcg9Vm5_1),.dout(w_dff_B_pvs0lKTW6_1),.clk(gclk));
	jdff dff_B_kMzW6HNz0_1(.din(w_dff_B_pvs0lKTW6_1),.dout(w_dff_B_kMzW6HNz0_1),.clk(gclk));
	jdff dff_B_vvt3UTDS2_1(.din(w_dff_B_kMzW6HNz0_1),.dout(w_dff_B_vvt3UTDS2_1),.clk(gclk));
	jdff dff_B_8K8sOztk2_1(.din(w_dff_B_vvt3UTDS2_1),.dout(w_dff_B_8K8sOztk2_1),.clk(gclk));
	jdff dff_B_lqwY6KzP5_1(.din(w_dff_B_8K8sOztk2_1),.dout(w_dff_B_lqwY6KzP5_1),.clk(gclk));
	jdff dff_B_LMwXuSfa5_1(.din(w_dff_B_lqwY6KzP5_1),.dout(w_dff_B_LMwXuSfa5_1),.clk(gclk));
	jdff dff_B_9wMV4Wy31_1(.din(w_dff_B_LMwXuSfa5_1),.dout(w_dff_B_9wMV4Wy31_1),.clk(gclk));
	jdff dff_B_zAJOaNse4_1(.din(w_dff_B_9wMV4Wy31_1),.dout(w_dff_B_zAJOaNse4_1),.clk(gclk));
	jdff dff_B_TOfUppsf6_1(.din(w_dff_B_zAJOaNse4_1),.dout(w_dff_B_TOfUppsf6_1),.clk(gclk));
	jdff dff_B_0NfPig3K9_1(.din(w_dff_B_TOfUppsf6_1),.dout(w_dff_B_0NfPig3K9_1),.clk(gclk));
	jdff dff_B_G1p4miaA2_1(.din(w_dff_B_0NfPig3K9_1),.dout(w_dff_B_G1p4miaA2_1),.clk(gclk));
	jdff dff_B_arAO3LTb2_1(.din(w_dff_B_G1p4miaA2_1),.dout(w_dff_B_arAO3LTb2_1),.clk(gclk));
	jdff dff_B_h2ZseJna0_1(.din(w_dff_B_arAO3LTb2_1),.dout(w_dff_B_h2ZseJna0_1),.clk(gclk));
	jdff dff_B_6Xsr2TIy5_1(.din(w_dff_B_h2ZseJna0_1),.dout(w_dff_B_6Xsr2TIy5_1),.clk(gclk));
	jdff dff_B_Ubk3OkEW4_1(.din(w_dff_B_6Xsr2TIy5_1),.dout(w_dff_B_Ubk3OkEW4_1),.clk(gclk));
	jdff dff_B_VNQEIJ2B7_1(.din(w_dff_B_Ubk3OkEW4_1),.dout(w_dff_B_VNQEIJ2B7_1),.clk(gclk));
	jdff dff_B_CCgQi8H14_1(.din(w_dff_B_VNQEIJ2B7_1),.dout(w_dff_B_CCgQi8H14_1),.clk(gclk));
	jdff dff_B_Oav8gulg4_1(.din(w_dff_B_CCgQi8H14_1),.dout(w_dff_B_Oav8gulg4_1),.clk(gclk));
	jdff dff_B_RQNtAc8l7_1(.din(w_dff_B_Oav8gulg4_1),.dout(w_dff_B_RQNtAc8l7_1),.clk(gclk));
	jdff dff_B_ZIFG6nf48_0(.din(n1502),.dout(w_dff_B_ZIFG6nf48_0),.clk(gclk));
	jdff dff_B_VPTJctPF0_0(.din(w_dff_B_ZIFG6nf48_0),.dout(w_dff_B_VPTJctPF0_0),.clk(gclk));
	jdff dff_B_filD7DCD1_0(.din(w_dff_B_VPTJctPF0_0),.dout(w_dff_B_filD7DCD1_0),.clk(gclk));
	jdff dff_B_oFAVvcJc8_0(.din(w_dff_B_filD7DCD1_0),.dout(w_dff_B_oFAVvcJc8_0),.clk(gclk));
	jdff dff_B_OwzwZ3Pz2_0(.din(w_dff_B_oFAVvcJc8_0),.dout(w_dff_B_OwzwZ3Pz2_0),.clk(gclk));
	jdff dff_B_ZfF76pED0_0(.din(w_dff_B_OwzwZ3Pz2_0),.dout(w_dff_B_ZfF76pED0_0),.clk(gclk));
	jdff dff_B_zsKa5CVc3_0(.din(w_dff_B_ZfF76pED0_0),.dout(w_dff_B_zsKa5CVc3_0),.clk(gclk));
	jdff dff_B_Jf18p4N64_0(.din(w_dff_B_zsKa5CVc3_0),.dout(w_dff_B_Jf18p4N64_0),.clk(gclk));
	jdff dff_B_v77hwnGl8_0(.din(w_dff_B_Jf18p4N64_0),.dout(w_dff_B_v77hwnGl8_0),.clk(gclk));
	jdff dff_B_PiQIMHru8_0(.din(w_dff_B_v77hwnGl8_0),.dout(w_dff_B_PiQIMHru8_0),.clk(gclk));
	jdff dff_B_few3mHEU3_0(.din(w_dff_B_PiQIMHru8_0),.dout(w_dff_B_few3mHEU3_0),.clk(gclk));
	jdff dff_B_CGo767pF6_0(.din(w_dff_B_few3mHEU3_0),.dout(w_dff_B_CGo767pF6_0),.clk(gclk));
	jdff dff_B_KQYFpcZO3_0(.din(w_dff_B_CGo767pF6_0),.dout(w_dff_B_KQYFpcZO3_0),.clk(gclk));
	jdff dff_B_yJ0NXdhk6_0(.din(w_dff_B_KQYFpcZO3_0),.dout(w_dff_B_yJ0NXdhk6_0),.clk(gclk));
	jdff dff_B_HHrZ6Q6R0_0(.din(w_dff_B_yJ0NXdhk6_0),.dout(w_dff_B_HHrZ6Q6R0_0),.clk(gclk));
	jdff dff_B_1uPdd0nj8_0(.din(w_dff_B_HHrZ6Q6R0_0),.dout(w_dff_B_1uPdd0nj8_0),.clk(gclk));
	jdff dff_B_EttT5PON4_0(.din(w_dff_B_1uPdd0nj8_0),.dout(w_dff_B_EttT5PON4_0),.clk(gclk));
	jdff dff_B_nDchxqvr3_0(.din(w_dff_B_EttT5PON4_0),.dout(w_dff_B_nDchxqvr3_0),.clk(gclk));
	jdff dff_B_EO5KVPZn6_0(.din(w_dff_B_nDchxqvr3_0),.dout(w_dff_B_EO5KVPZn6_0),.clk(gclk));
	jdff dff_B_kwGuXUXQ2_0(.din(w_dff_B_EO5KVPZn6_0),.dout(w_dff_B_kwGuXUXQ2_0),.clk(gclk));
	jdff dff_B_y6jLaFWv5_1(.din(n1497),.dout(w_dff_B_y6jLaFWv5_1),.clk(gclk));
	jdff dff_B_fY56sq2l1_1(.din(w_dff_B_y6jLaFWv5_1),.dout(w_dff_B_fY56sq2l1_1),.clk(gclk));
	jdff dff_B_BiUg6YDy3_0(.din(n1498),.dout(w_dff_B_BiUg6YDy3_0),.clk(gclk));
	jdff dff_B_u2tlrm4O5_0(.din(w_dff_B_BiUg6YDy3_0),.dout(w_dff_B_u2tlrm4O5_0),.clk(gclk));
	jdff dff_B_W66BIxzs5_0(.din(w_dff_B_u2tlrm4O5_0),.dout(w_dff_B_W66BIxzs5_0),.clk(gclk));
	jdff dff_B_e1JuA95y3_0(.din(w_dff_B_W66BIxzs5_0),.dout(w_dff_B_e1JuA95y3_0),.clk(gclk));
	jdff dff_B_INzzAuzd4_0(.din(w_dff_B_e1JuA95y3_0),.dout(w_dff_B_INzzAuzd4_0),.clk(gclk));
	jdff dff_A_FajkBpHE7_1(.dout(w_n1364_0[1]),.din(w_dff_A_FajkBpHE7_1),.clk(gclk));
	jdff dff_A_UBZNhFsc9_1(.dout(w_dff_A_FajkBpHE7_1),.din(w_dff_A_UBZNhFsc9_1),.clk(gclk));
	jdff dff_A_sSjpLx367_1(.dout(w_dff_A_UBZNhFsc9_1),.din(w_dff_A_sSjpLx367_1),.clk(gclk));
	jdff dff_A_l0oPRfmY3_1(.dout(w_dff_A_sSjpLx367_1),.din(w_dff_A_l0oPRfmY3_1),.clk(gclk));
	jdff dff_A_BmyqDzfJ2_1(.dout(w_dff_A_l0oPRfmY3_1),.din(w_dff_A_BmyqDzfJ2_1),.clk(gclk));
	jdff dff_A_8eK0kAel7_1(.dout(w_dff_A_BmyqDzfJ2_1),.din(w_dff_A_8eK0kAel7_1),.clk(gclk));
	jdff dff_A_wcfNUdRJ4_1(.dout(w_dff_A_8eK0kAel7_1),.din(w_dff_A_wcfNUdRJ4_1),.clk(gclk));
	jdff dff_A_7pTc6CZs1_1(.dout(w_dff_A_wcfNUdRJ4_1),.din(w_dff_A_7pTc6CZs1_1),.clk(gclk));
	jdff dff_A_TqpQzs9O1_1(.dout(w_dff_A_7pTc6CZs1_1),.din(w_dff_A_TqpQzs9O1_1),.clk(gclk));
	jdff dff_A_IOVYzYAs3_1(.dout(w_dff_A_TqpQzs9O1_1),.din(w_dff_A_IOVYzYAs3_1),.clk(gclk));
	jdff dff_A_Oc2YygRX0_1(.dout(w_dff_A_IOVYzYAs3_1),.din(w_dff_A_Oc2YygRX0_1),.clk(gclk));
	jdff dff_A_S6VsueXs1_1(.dout(w_dff_A_Oc2YygRX0_1),.din(w_dff_A_S6VsueXs1_1),.clk(gclk));
	jdff dff_A_Z5MDXOdj9_1(.dout(w_dff_A_S6VsueXs1_1),.din(w_dff_A_Z5MDXOdj9_1),.clk(gclk));
	jdff dff_A_l8Z1Tr2Y5_1(.dout(w_dff_A_Z5MDXOdj9_1),.din(w_dff_A_l8Z1Tr2Y5_1),.clk(gclk));
	jdff dff_A_1KjP9csF4_1(.dout(w_dff_A_l8Z1Tr2Y5_1),.din(w_dff_A_1KjP9csF4_1),.clk(gclk));
	jdff dff_A_3U1leG9n6_1(.dout(w_dff_A_1KjP9csF4_1),.din(w_dff_A_3U1leG9n6_1),.clk(gclk));
	jdff dff_A_V2tacE9T4_1(.dout(w_dff_A_3U1leG9n6_1),.din(w_dff_A_V2tacE9T4_1),.clk(gclk));
	jdff dff_A_XroujTcU7_1(.dout(w_dff_A_V2tacE9T4_1),.din(w_dff_A_XroujTcU7_1),.clk(gclk));
	jdff dff_A_XiW6w5JV9_1(.dout(w_dff_A_XroujTcU7_1),.din(w_dff_A_XiW6w5JV9_1),.clk(gclk));
	jdff dff_A_OCUELDqV1_1(.dout(w_dff_A_XiW6w5JV9_1),.din(w_dff_A_OCUELDqV1_1),.clk(gclk));
	jdff dff_A_xIq35Qv42_1(.dout(w_dff_A_OCUELDqV1_1),.din(w_dff_A_xIq35Qv42_1),.clk(gclk));
	jdff dff_A_o6T7RTMj2_1(.dout(w_dff_A_xIq35Qv42_1),.din(w_dff_A_o6T7RTMj2_1),.clk(gclk));
	jdff dff_A_hTFS2Vpd0_1(.dout(w_dff_A_o6T7RTMj2_1),.din(w_dff_A_hTFS2Vpd0_1),.clk(gclk));
	jdff dff_A_QtcHqgc40_1(.dout(w_dff_A_hTFS2Vpd0_1),.din(w_dff_A_QtcHqgc40_1),.clk(gclk));
	jdff dff_A_WB2CvrJW5_1(.dout(w_dff_A_QtcHqgc40_1),.din(w_dff_A_WB2CvrJW5_1),.clk(gclk));
	jdff dff_B_JiERR1Iq0_0(.din(n1363),.dout(w_dff_B_JiERR1Iq0_0),.clk(gclk));
	jdff dff_B_2ARvBBtH9_0(.din(w_dff_B_JiERR1Iq0_0),.dout(w_dff_B_2ARvBBtH9_0),.clk(gclk));
	jdff dff_B_qzHqw6h73_0(.din(w_dff_B_2ARvBBtH9_0),.dout(w_dff_B_qzHqw6h73_0),.clk(gclk));
	jdff dff_B_xnTx0TVi2_1(.din(n1494),.dout(w_dff_B_xnTx0TVi2_1),.clk(gclk));
	jdff dff_B_lP1eYBD99_1(.din(w_dff_B_xnTx0TVi2_1),.dout(w_dff_B_lP1eYBD99_1),.clk(gclk));
	jdff dff_B_y1FHGEko7_1(.din(w_dff_B_lP1eYBD99_1),.dout(w_dff_B_y1FHGEko7_1),.clk(gclk));
	jdff dff_B_57MVZArM1_1(.din(n1495),.dout(w_dff_B_57MVZArM1_1),.clk(gclk));
	jdff dff_B_azEqYxyT5_1(.din(w_dff_B_57MVZArM1_1),.dout(w_dff_B_azEqYxyT5_1),.clk(gclk));
	jdff dff_A_f8cSmmCn9_1(.dout(w_n1359_0[1]),.din(w_dff_A_f8cSmmCn9_1),.clk(gclk));
	jdff dff_A_35OU87DK2_1(.dout(w_dff_A_f8cSmmCn9_1),.din(w_dff_A_35OU87DK2_1),.clk(gclk));
	jdff dff_A_RgOlcgrK5_1(.dout(w_dff_A_35OU87DK2_1),.din(w_dff_A_RgOlcgrK5_1),.clk(gclk));
	jdff dff_A_wHuEb2lj3_1(.dout(w_dff_A_RgOlcgrK5_1),.din(w_dff_A_wHuEb2lj3_1),.clk(gclk));
	jdff dff_A_KFaKO4vd4_1(.dout(w_dff_A_wHuEb2lj3_1),.din(w_dff_A_KFaKO4vd4_1),.clk(gclk));
	jdff dff_A_XQnY0Vo61_1(.dout(w_dff_A_KFaKO4vd4_1),.din(w_dff_A_XQnY0Vo61_1),.clk(gclk));
	jdff dff_A_nZPq9cQh5_1(.dout(w_dff_A_XQnY0Vo61_1),.din(w_dff_A_nZPq9cQh5_1),.clk(gclk));
	jdff dff_A_hXUpu4BD6_1(.dout(w_dff_A_nZPq9cQh5_1),.din(w_dff_A_hXUpu4BD6_1),.clk(gclk));
	jdff dff_A_6bLof3eb8_1(.dout(w_dff_A_hXUpu4BD6_1),.din(w_dff_A_6bLof3eb8_1),.clk(gclk));
	jdff dff_A_gBSzMHpX3_1(.dout(w_dff_A_6bLof3eb8_1),.din(w_dff_A_gBSzMHpX3_1),.clk(gclk));
	jdff dff_A_JhXtz3Ss1_1(.dout(w_dff_A_gBSzMHpX3_1),.din(w_dff_A_JhXtz3Ss1_1),.clk(gclk));
	jdff dff_A_3SwhL6qs9_1(.dout(w_dff_A_JhXtz3Ss1_1),.din(w_dff_A_3SwhL6qs9_1),.clk(gclk));
	jdff dff_A_SuPxILcn6_1(.dout(w_dff_A_3SwhL6qs9_1),.din(w_dff_A_SuPxILcn6_1),.clk(gclk));
	jdff dff_A_QeM17DCO2_1(.dout(w_dff_A_SuPxILcn6_1),.din(w_dff_A_QeM17DCO2_1),.clk(gclk));
	jdff dff_A_UZfkibCq1_1(.dout(w_dff_A_QeM17DCO2_1),.din(w_dff_A_UZfkibCq1_1),.clk(gclk));
	jdff dff_A_wG4CRCBj7_1(.dout(w_dff_A_UZfkibCq1_1),.din(w_dff_A_wG4CRCBj7_1),.clk(gclk));
	jdff dff_A_HQZuX8Zv8_1(.dout(w_dff_A_wG4CRCBj7_1),.din(w_dff_A_HQZuX8Zv8_1),.clk(gclk));
	jdff dff_A_3LeyG6A52_1(.dout(w_dff_A_HQZuX8Zv8_1),.din(w_dff_A_3LeyG6A52_1),.clk(gclk));
	jdff dff_A_W3yrwK1G2_1(.dout(w_dff_A_3LeyG6A52_1),.din(w_dff_A_W3yrwK1G2_1),.clk(gclk));
	jdff dff_A_cTh2FNYV6_1(.dout(w_dff_A_W3yrwK1G2_1),.din(w_dff_A_cTh2FNYV6_1),.clk(gclk));
	jdff dff_A_UJXvJUo44_1(.dout(w_dff_A_cTh2FNYV6_1),.din(w_dff_A_UJXvJUo44_1),.clk(gclk));
	jdff dff_A_TWZkus282_1(.dout(w_dff_A_UJXvJUo44_1),.din(w_dff_A_TWZkus282_1),.clk(gclk));
	jdff dff_B_a3SJFK7E1_2(.din(n1359),.dout(w_dff_B_a3SJFK7E1_2),.clk(gclk));
	jdff dff_A_9CY54BSs3_0(.dout(w_n418_0[0]),.din(w_dff_A_9CY54BSs3_0),.clk(gclk));
	jdff dff_A_XHzGi9Jr4_0(.dout(w_dff_A_9CY54BSs3_0),.din(w_dff_A_XHzGi9Jr4_0),.clk(gclk));
	jdff dff_A_22JjTXqe3_0(.dout(w_dff_A_XHzGi9Jr4_0),.din(w_dff_A_22JjTXqe3_0),.clk(gclk));
	jdff dff_A_cr1hPzEY8_0(.dout(w_dff_A_22JjTXqe3_0),.din(w_dff_A_cr1hPzEY8_0),.clk(gclk));
	jdff dff_A_1E9O2vqX7_0(.dout(w_dff_A_cr1hPzEY8_0),.din(w_dff_A_1E9O2vqX7_0),.clk(gclk));
	jdff dff_B_FyQNE8XS5_1(.din(n1324),.dout(w_dff_B_FyQNE8XS5_1),.clk(gclk));
	jdff dff_B_hMyXcZCq6_1(.din(w_dff_B_FyQNE8XS5_1),.dout(w_dff_B_hMyXcZCq6_1),.clk(gclk));
	jdff dff_B_mYAMaaH61_1(.din(w_dff_B_hMyXcZCq6_1),.dout(w_dff_B_mYAMaaH61_1),.clk(gclk));
	jdff dff_B_KfqJFjZz0_1(.din(w_dff_B_mYAMaaH61_1),.dout(w_dff_B_KfqJFjZz0_1),.clk(gclk));
	jdff dff_B_2XDJCDok9_1(.din(w_dff_B_KfqJFjZz0_1),.dout(w_dff_B_2XDJCDok9_1),.clk(gclk));
	jdff dff_B_ocGeuNd14_1(.din(w_dff_B_2XDJCDok9_1),.dout(w_dff_B_ocGeuNd14_1),.clk(gclk));
	jdff dff_B_tQ5mKweV1_1(.din(w_dff_B_ocGeuNd14_1),.dout(w_dff_B_tQ5mKweV1_1),.clk(gclk));
	jdff dff_B_vSOESnuB6_1(.din(w_dff_B_tQ5mKweV1_1),.dout(w_dff_B_vSOESnuB6_1),.clk(gclk));
	jdff dff_B_4vwUtX5y7_1(.din(w_dff_B_vSOESnuB6_1),.dout(w_dff_B_4vwUtX5y7_1),.clk(gclk));
	jdff dff_B_vonLHBY13_1(.din(w_dff_B_4vwUtX5y7_1),.dout(w_dff_B_vonLHBY13_1),.clk(gclk));
	jdff dff_B_83Vkj7219_1(.din(w_dff_B_vonLHBY13_1),.dout(w_dff_B_83Vkj7219_1),.clk(gclk));
	jdff dff_B_7yZszsJV6_1(.din(w_dff_B_83Vkj7219_1),.dout(w_dff_B_7yZszsJV6_1),.clk(gclk));
	jdff dff_B_NxWmUapD7_1(.din(w_dff_B_7yZszsJV6_1),.dout(w_dff_B_NxWmUapD7_1),.clk(gclk));
	jdff dff_B_KH17Yc3t7_1(.din(w_dff_B_NxWmUapD7_1),.dout(w_dff_B_KH17Yc3t7_1),.clk(gclk));
	jdff dff_B_JVgoryDw9_1(.din(w_dff_B_KH17Yc3t7_1),.dout(w_dff_B_JVgoryDw9_1),.clk(gclk));
	jdff dff_B_jYNCGmAX8_1(.din(w_dff_B_JVgoryDw9_1),.dout(w_dff_B_jYNCGmAX8_1),.clk(gclk));
	jdff dff_B_L0Q5T17N2_1(.din(w_dff_B_jYNCGmAX8_1),.dout(w_dff_B_L0Q5T17N2_1),.clk(gclk));
	jdff dff_B_1CLltA5J4_1(.din(w_dff_B_L0Q5T17N2_1),.dout(w_dff_B_1CLltA5J4_1),.clk(gclk));
	jdff dff_B_Gx05KMYm4_1(.din(w_dff_B_1CLltA5J4_1),.dout(w_dff_B_Gx05KMYm4_1),.clk(gclk));
	jdff dff_B_q8x3KuWt4_1(.din(w_dff_B_Gx05KMYm4_1),.dout(w_dff_B_q8x3KuWt4_1),.clk(gclk));
	jdff dff_B_9SzYDlrH2_1(.din(w_dff_B_q8x3KuWt4_1),.dout(w_dff_B_9SzYDlrH2_1),.clk(gclk));
	jdff dff_B_Kfiz4VTJ4_1(.din(w_dff_B_9SzYDlrH2_1),.dout(w_dff_B_Kfiz4VTJ4_1),.clk(gclk));
	jdff dff_B_dckUumh78_1(.din(w_dff_B_Kfiz4VTJ4_1),.dout(w_dff_B_dckUumh78_1),.clk(gclk));
	jdff dff_B_k78dmU431_1(.din(w_dff_B_dckUumh78_1),.dout(w_dff_B_k78dmU431_1),.clk(gclk));
	jdff dff_B_hGk3aXMW6_1(.din(w_dff_B_k78dmU431_1),.dout(w_dff_B_hGk3aXMW6_1),.clk(gclk));
	jdff dff_B_XOV5dNNa5_1(.din(w_dff_B_hGk3aXMW6_1),.dout(w_dff_B_XOV5dNNa5_1),.clk(gclk));
	jdff dff_B_2KWgNVkv5_1(.din(w_dff_B_XOV5dNNa5_1),.dout(w_dff_B_2KWgNVkv5_1),.clk(gclk));
	jdff dff_B_KmzGxk4w4_1(.din(w_dff_B_2KWgNVkv5_1),.dout(w_dff_B_KmzGxk4w4_1),.clk(gclk));
	jdff dff_B_UuxtBApE6_1(.din(n1325),.dout(w_dff_B_UuxtBApE6_1),.clk(gclk));
	jdff dff_B_kgdgUzU63_1(.din(w_dff_B_UuxtBApE6_1),.dout(w_dff_B_kgdgUzU63_1),.clk(gclk));
	jdff dff_B_mjnOfVEj5_1(.din(w_dff_B_kgdgUzU63_1),.dout(w_dff_B_mjnOfVEj5_1),.clk(gclk));
	jdff dff_B_jjJdIxsd7_1(.din(w_dff_B_mjnOfVEj5_1),.dout(w_dff_B_jjJdIxsd7_1),.clk(gclk));
	jdff dff_B_lspRqeE73_1(.din(w_dff_B_jjJdIxsd7_1),.dout(w_dff_B_lspRqeE73_1),.clk(gclk));
	jdff dff_B_gwTe6ssh4_1(.din(w_dff_B_lspRqeE73_1),.dout(w_dff_B_gwTe6ssh4_1),.clk(gclk));
	jdff dff_B_Md7ixU3w3_1(.din(w_dff_B_gwTe6ssh4_1),.dout(w_dff_B_Md7ixU3w3_1),.clk(gclk));
	jdff dff_B_wuHD7whs2_1(.din(w_dff_B_Md7ixU3w3_1),.dout(w_dff_B_wuHD7whs2_1),.clk(gclk));
	jdff dff_B_0UrAc8Nk5_1(.din(w_dff_B_wuHD7whs2_1),.dout(w_dff_B_0UrAc8Nk5_1),.clk(gclk));
	jdff dff_B_6aehAtxn9_1(.din(w_dff_B_0UrAc8Nk5_1),.dout(w_dff_B_6aehAtxn9_1),.clk(gclk));
	jdff dff_B_kLm88onJ5_1(.din(w_dff_B_6aehAtxn9_1),.dout(w_dff_B_kLm88onJ5_1),.clk(gclk));
	jdff dff_B_XbUdJMHW0_1(.din(w_dff_B_kLm88onJ5_1),.dout(w_dff_B_XbUdJMHW0_1),.clk(gclk));
	jdff dff_B_Jgu0j0xR7_1(.din(w_dff_B_XbUdJMHW0_1),.dout(w_dff_B_Jgu0j0xR7_1),.clk(gclk));
	jdff dff_B_FZiKhB0O5_1(.din(w_dff_B_Jgu0j0xR7_1),.dout(w_dff_B_FZiKhB0O5_1),.clk(gclk));
	jdff dff_B_WfgI7hsW9_1(.din(w_dff_B_FZiKhB0O5_1),.dout(w_dff_B_WfgI7hsW9_1),.clk(gclk));
	jdff dff_B_sP7NPzcD3_1(.din(w_dff_B_WfgI7hsW9_1),.dout(w_dff_B_sP7NPzcD3_1),.clk(gclk));
	jdff dff_B_LFetKh0N2_1(.din(w_dff_B_sP7NPzcD3_1),.dout(w_dff_B_LFetKh0N2_1),.clk(gclk));
	jdff dff_B_s1j3VRCI0_1(.din(w_dff_B_LFetKh0N2_1),.dout(w_dff_B_s1j3VRCI0_1),.clk(gclk));
	jdff dff_B_JQFZhxoG3_1(.din(w_dff_B_s1j3VRCI0_1),.dout(w_dff_B_JQFZhxoG3_1),.clk(gclk));
	jdff dff_B_KCDDsFAB6_1(.din(w_dff_B_JQFZhxoG3_1),.dout(w_dff_B_KCDDsFAB6_1),.clk(gclk));
	jdff dff_B_wkaufNKd8_1(.din(w_dff_B_KCDDsFAB6_1),.dout(w_dff_B_wkaufNKd8_1),.clk(gclk));
	jdff dff_B_6ityTnxH3_1(.din(w_dff_B_wkaufNKd8_1),.dout(w_dff_B_6ityTnxH3_1),.clk(gclk));
	jdff dff_B_nc4DORdT0_1(.din(w_dff_B_6ityTnxH3_1),.dout(w_dff_B_nc4DORdT0_1),.clk(gclk));
	jdff dff_B_t5VmvgvV9_1(.din(w_dff_B_nc4DORdT0_1),.dout(w_dff_B_t5VmvgvV9_1),.clk(gclk));
	jdff dff_B_Wxi7Li0q3_1(.din(w_dff_B_t5VmvgvV9_1),.dout(w_dff_B_Wxi7Li0q3_1),.clk(gclk));
	jdff dff_B_iItRIaRy7_1(.din(w_dff_B_Wxi7Li0q3_1),.dout(w_dff_B_iItRIaRy7_1),.clk(gclk));
	jdff dff_B_6gFcWADp7_1(.din(w_dff_B_iItRIaRy7_1),.dout(w_dff_B_6gFcWADp7_1),.clk(gclk));
	jdff dff_B_NFuqLFRS5_1(.din(n1326),.dout(w_dff_B_NFuqLFRS5_1),.clk(gclk));
	jdff dff_B_e1Nbm4jB5_1(.din(w_dff_B_NFuqLFRS5_1),.dout(w_dff_B_e1Nbm4jB5_1),.clk(gclk));
	jdff dff_B_BE6TCiES2_1(.din(w_dff_B_e1Nbm4jB5_1),.dout(w_dff_B_BE6TCiES2_1),.clk(gclk));
	jdff dff_B_rEz2ctfc6_1(.din(w_dff_B_BE6TCiES2_1),.dout(w_dff_B_rEz2ctfc6_1),.clk(gclk));
	jdff dff_B_v5nlcT5a1_1(.din(w_dff_B_rEz2ctfc6_1),.dout(w_dff_B_v5nlcT5a1_1),.clk(gclk));
	jdff dff_B_gSYitMou4_1(.din(w_dff_B_v5nlcT5a1_1),.dout(w_dff_B_gSYitMou4_1),.clk(gclk));
	jdff dff_B_uUUtTRDO4_1(.din(w_dff_B_gSYitMou4_1),.dout(w_dff_B_uUUtTRDO4_1),.clk(gclk));
	jdff dff_B_i8HOPdLC2_1(.din(w_dff_B_uUUtTRDO4_1),.dout(w_dff_B_i8HOPdLC2_1),.clk(gclk));
	jdff dff_B_k7zfV01k8_1(.din(w_dff_B_i8HOPdLC2_1),.dout(w_dff_B_k7zfV01k8_1),.clk(gclk));
	jdff dff_B_YUnwslQ83_1(.din(w_dff_B_k7zfV01k8_1),.dout(w_dff_B_YUnwslQ83_1),.clk(gclk));
	jdff dff_B_GX9SKCAI0_1(.din(w_dff_B_YUnwslQ83_1),.dout(w_dff_B_GX9SKCAI0_1),.clk(gclk));
	jdff dff_B_RbCXqxy93_1(.din(w_dff_B_GX9SKCAI0_1),.dout(w_dff_B_RbCXqxy93_1),.clk(gclk));
	jdff dff_B_xweBRsBM1_1(.din(w_dff_B_RbCXqxy93_1),.dout(w_dff_B_xweBRsBM1_1),.clk(gclk));
	jdff dff_B_7dwATRM32_1(.din(w_dff_B_xweBRsBM1_1),.dout(w_dff_B_7dwATRM32_1),.clk(gclk));
	jdff dff_B_exD9w7Jj8_1(.din(w_dff_B_7dwATRM32_1),.dout(w_dff_B_exD9w7Jj8_1),.clk(gclk));
	jdff dff_B_X8LozdNv4_1(.din(w_dff_B_exD9w7Jj8_1),.dout(w_dff_B_X8LozdNv4_1),.clk(gclk));
	jdff dff_B_wFA1FKeK2_1(.din(w_dff_B_X8LozdNv4_1),.dout(w_dff_B_wFA1FKeK2_1),.clk(gclk));
	jdff dff_B_tKBrGSFa3_1(.din(w_dff_B_wFA1FKeK2_1),.dout(w_dff_B_tKBrGSFa3_1),.clk(gclk));
	jdff dff_B_LwvcJn2Y5_1(.din(w_dff_B_tKBrGSFa3_1),.dout(w_dff_B_LwvcJn2Y5_1),.clk(gclk));
	jdff dff_B_1mrE3lYF9_1(.din(w_dff_B_LwvcJn2Y5_1),.dout(w_dff_B_1mrE3lYF9_1),.clk(gclk));
	jdff dff_B_qtVtrj7r8_1(.din(w_dff_B_1mrE3lYF9_1),.dout(w_dff_B_qtVtrj7r8_1),.clk(gclk));
	jdff dff_B_ZsmpZskx1_1(.din(n1327),.dout(w_dff_B_ZsmpZskx1_1),.clk(gclk));
	jdff dff_B_Le4P70Ot2_1(.din(w_dff_B_ZsmpZskx1_1),.dout(w_dff_B_Le4P70Ot2_1),.clk(gclk));
	jdff dff_B_jB6DICeT0_1(.din(w_dff_B_Le4P70Ot2_1),.dout(w_dff_B_jB6DICeT0_1),.clk(gclk));
	jdff dff_B_ycODkcrf4_1(.din(w_dff_B_jB6DICeT0_1),.dout(w_dff_B_ycODkcrf4_1),.clk(gclk));
	jdff dff_B_IYIgiYo72_1(.din(w_dff_B_ycODkcrf4_1),.dout(w_dff_B_IYIgiYo72_1),.clk(gclk));
	jdff dff_B_hJRc0dPJ1_1(.din(w_dff_B_IYIgiYo72_1),.dout(w_dff_B_hJRc0dPJ1_1),.clk(gclk));
	jdff dff_B_iV4lKNpO6_1(.din(w_dff_B_hJRc0dPJ1_1),.dout(w_dff_B_iV4lKNpO6_1),.clk(gclk));
	jdff dff_B_JtWnfbAq1_1(.din(w_dff_B_iV4lKNpO6_1),.dout(w_dff_B_JtWnfbAq1_1),.clk(gclk));
	jdff dff_B_yDGNHflk5_1(.din(w_dff_B_JtWnfbAq1_1),.dout(w_dff_B_yDGNHflk5_1),.clk(gclk));
	jdff dff_B_A6e4ZRcf8_1(.din(w_dff_B_yDGNHflk5_1),.dout(w_dff_B_A6e4ZRcf8_1),.clk(gclk));
	jdff dff_B_xJrEr7jx1_1(.din(w_dff_B_A6e4ZRcf8_1),.dout(w_dff_B_xJrEr7jx1_1),.clk(gclk));
	jdff dff_B_OdY8VVL85_1(.din(w_dff_B_xJrEr7jx1_1),.dout(w_dff_B_OdY8VVL85_1),.clk(gclk));
	jdff dff_B_2D0Xl9bl6_1(.din(w_dff_B_OdY8VVL85_1),.dout(w_dff_B_2D0Xl9bl6_1),.clk(gclk));
	jdff dff_B_hxBAdlmy9_1(.din(w_dff_B_2D0Xl9bl6_1),.dout(w_dff_B_hxBAdlmy9_1),.clk(gclk));
	jdff dff_B_Hyo3IW770_1(.din(w_dff_B_hxBAdlmy9_1),.dout(w_dff_B_Hyo3IW770_1),.clk(gclk));
	jdff dff_B_HyuUShvg7_1(.din(w_dff_B_Hyo3IW770_1),.dout(w_dff_B_HyuUShvg7_1),.clk(gclk));
	jdff dff_B_618PvWUD2_1(.din(w_dff_B_HyuUShvg7_1),.dout(w_dff_B_618PvWUD2_1),.clk(gclk));
	jdff dff_B_mGx99hM97_1(.din(w_dff_B_618PvWUD2_1),.dout(w_dff_B_mGx99hM97_1),.clk(gclk));
	jdff dff_B_oARdvx0O9_1(.din(w_dff_B_mGx99hM97_1),.dout(w_dff_B_oARdvx0O9_1),.clk(gclk));
	jdff dff_B_jUTm8CVk7_1(.din(w_dff_B_oARdvx0O9_1),.dout(w_dff_B_jUTm8CVk7_1),.clk(gclk));
	jdff dff_B_QDCFzGIp4_1(.din(w_dff_B_jUTm8CVk7_1),.dout(w_dff_B_QDCFzGIp4_1),.clk(gclk));
	jdff dff_B_HLGIwBVv4_1(.din(n1328),.dout(w_dff_B_HLGIwBVv4_1),.clk(gclk));
	jdff dff_B_aU46LyhX4_1(.din(w_dff_B_HLGIwBVv4_1),.dout(w_dff_B_aU46LyhX4_1),.clk(gclk));
	jdff dff_B_b3E2JgJ75_1(.din(w_dff_B_aU46LyhX4_1),.dout(w_dff_B_b3E2JgJ75_1),.clk(gclk));
	jdff dff_B_nzMu3MQf1_1(.din(w_dff_B_b3E2JgJ75_1),.dout(w_dff_B_nzMu3MQf1_1),.clk(gclk));
	jdff dff_B_Na4DGaBP4_1(.din(w_dff_B_nzMu3MQf1_1),.dout(w_dff_B_Na4DGaBP4_1),.clk(gclk));
	jdff dff_B_0DGm8ZVX2_1(.din(w_dff_B_Na4DGaBP4_1),.dout(w_dff_B_0DGm8ZVX2_1),.clk(gclk));
	jdff dff_B_wjyj0WKK4_1(.din(w_dff_B_0DGm8ZVX2_1),.dout(w_dff_B_wjyj0WKK4_1),.clk(gclk));
	jdff dff_B_8MXny79A3_1(.din(w_dff_B_wjyj0WKK4_1),.dout(w_dff_B_8MXny79A3_1),.clk(gclk));
	jdff dff_B_rXONjn159_1(.din(w_dff_B_8MXny79A3_1),.dout(w_dff_B_rXONjn159_1),.clk(gclk));
	jdff dff_B_kFcP249J9_1(.din(w_dff_B_rXONjn159_1),.dout(w_dff_B_kFcP249J9_1),.clk(gclk));
	jdff dff_B_sjs9PK3f1_1(.din(w_dff_B_kFcP249J9_1),.dout(w_dff_B_sjs9PK3f1_1),.clk(gclk));
	jdff dff_B_mQgQ7USW3_1(.din(w_dff_B_sjs9PK3f1_1),.dout(w_dff_B_mQgQ7USW3_1),.clk(gclk));
	jdff dff_B_pBpIIhvz7_1(.din(w_dff_B_mQgQ7USW3_1),.dout(w_dff_B_pBpIIhvz7_1),.clk(gclk));
	jdff dff_B_67vwr24W4_1(.din(w_dff_B_pBpIIhvz7_1),.dout(w_dff_B_67vwr24W4_1),.clk(gclk));
	jdff dff_B_Ccl6R05j0_1(.din(w_dff_B_67vwr24W4_1),.dout(w_dff_B_Ccl6R05j0_1),.clk(gclk));
	jdff dff_B_YiFqbGVX2_1(.din(w_dff_B_Ccl6R05j0_1),.dout(w_dff_B_YiFqbGVX2_1),.clk(gclk));
	jdff dff_B_SMa0Ue6V0_1(.din(n1329),.dout(w_dff_B_SMa0Ue6V0_1),.clk(gclk));
	jdff dff_B_m25LymCS0_1(.din(w_dff_B_SMa0Ue6V0_1),.dout(w_dff_B_m25LymCS0_1),.clk(gclk));
	jdff dff_B_1FZOIzhJ1_1(.din(w_dff_B_m25LymCS0_1),.dout(w_dff_B_1FZOIzhJ1_1),.clk(gclk));
	jdff dff_B_LoQlbB2L8_1(.din(w_dff_B_1FZOIzhJ1_1),.dout(w_dff_B_LoQlbB2L8_1),.clk(gclk));
	jdff dff_B_VmyuVrLh6_1(.din(w_dff_B_LoQlbB2L8_1),.dout(w_dff_B_VmyuVrLh6_1),.clk(gclk));
	jdff dff_B_nO889iOG1_1(.din(w_dff_B_VmyuVrLh6_1),.dout(w_dff_B_nO889iOG1_1),.clk(gclk));
	jdff dff_B_Ywhl824d5_1(.din(w_dff_B_nO889iOG1_1),.dout(w_dff_B_Ywhl824d5_1),.clk(gclk));
	jdff dff_B_mDKbaS6F0_1(.din(w_dff_B_Ywhl824d5_1),.dout(w_dff_B_mDKbaS6F0_1),.clk(gclk));
	jdff dff_B_xwiRNtQZ0_1(.din(w_dff_B_mDKbaS6F0_1),.dout(w_dff_B_xwiRNtQZ0_1),.clk(gclk));
	jdff dff_B_vkejMAam6_1(.din(w_dff_B_xwiRNtQZ0_1),.dout(w_dff_B_vkejMAam6_1),.clk(gclk));
	jdff dff_B_5A6KfDUS4_1(.din(w_dff_B_vkejMAam6_1),.dout(w_dff_B_5A6KfDUS4_1),.clk(gclk));
	jdff dff_B_MRxhsvNs4_1(.din(w_dff_B_5A6KfDUS4_1),.dout(w_dff_B_MRxhsvNs4_1),.clk(gclk));
	jdff dff_B_5YEcKngC6_1(.din(w_dff_B_MRxhsvNs4_1),.dout(w_dff_B_5YEcKngC6_1),.clk(gclk));
	jdff dff_B_iNFNxHr21_1(.din(w_dff_B_5YEcKngC6_1),.dout(w_dff_B_iNFNxHr21_1),.clk(gclk));
	jdff dff_B_AbJ7Z0fu5_1(.din(w_dff_B_iNFNxHr21_1),.dout(w_dff_B_AbJ7Z0fu5_1),.clk(gclk));
	jdff dff_B_KAjw9nXX1_1(.din(w_dff_B_AbJ7Z0fu5_1),.dout(w_dff_B_KAjw9nXX1_1),.clk(gclk));
	jdff dff_B_UXF6fFBc8_1(.din(w_dff_B_KAjw9nXX1_1),.dout(w_dff_B_UXF6fFBc8_1),.clk(gclk));
	jdff dff_B_omzyU4fI5_1(.din(n1330),.dout(w_dff_B_omzyU4fI5_1),.clk(gclk));
	jdff dff_B_k1nw84Sn9_1(.din(w_dff_B_omzyU4fI5_1),.dout(w_dff_B_k1nw84Sn9_1),.clk(gclk));
	jdff dff_B_PDI63GOE2_1(.din(w_dff_B_k1nw84Sn9_1),.dout(w_dff_B_PDI63GOE2_1),.clk(gclk));
	jdff dff_B_vobuiUjm5_1(.din(w_dff_B_PDI63GOE2_1),.dout(w_dff_B_vobuiUjm5_1),.clk(gclk));
	jdff dff_B_c6slsYjW3_1(.din(w_dff_B_vobuiUjm5_1),.dout(w_dff_B_c6slsYjW3_1),.clk(gclk));
	jdff dff_B_CjjnwJBo7_1(.din(w_dff_B_c6slsYjW3_1),.dout(w_dff_B_CjjnwJBo7_1),.clk(gclk));
	jdff dff_B_BQ9Dt4NL1_1(.din(w_dff_B_CjjnwJBo7_1),.dout(w_dff_B_BQ9Dt4NL1_1),.clk(gclk));
	jdff dff_B_DyYlIAEO6_1(.din(w_dff_B_BQ9Dt4NL1_1),.dout(w_dff_B_DyYlIAEO6_1),.clk(gclk));
	jdff dff_B_FIIhOPuE1_1(.din(w_dff_B_DyYlIAEO6_1),.dout(w_dff_B_FIIhOPuE1_1),.clk(gclk));
	jdff dff_B_ia5UFewF2_1(.din(w_dff_B_FIIhOPuE1_1),.dout(w_dff_B_ia5UFewF2_1),.clk(gclk));
	jdff dff_B_aIuIpuQN4_1(.din(w_dff_B_ia5UFewF2_1),.dout(w_dff_B_aIuIpuQN4_1),.clk(gclk));
	jdff dff_B_RzXcr7NG3_1(.din(w_dff_B_aIuIpuQN4_1),.dout(w_dff_B_RzXcr7NG3_1),.clk(gclk));
	jdff dff_B_5dSlsuGz1_1(.din(w_dff_B_RzXcr7NG3_1),.dout(w_dff_B_5dSlsuGz1_1),.clk(gclk));
	jdff dff_B_wTcfhqba2_1(.din(w_dff_B_5dSlsuGz1_1),.dout(w_dff_B_wTcfhqba2_1),.clk(gclk));
	jdff dff_B_S7MtSNHF6_1(.din(w_dff_B_wTcfhqba2_1),.dout(w_dff_B_S7MtSNHF6_1),.clk(gclk));
	jdff dff_B_x4A1eFdW1_1(.din(w_dff_B_S7MtSNHF6_1),.dout(w_dff_B_x4A1eFdW1_1),.clk(gclk));
	jdff dff_B_iue93fgv9_1(.din(w_dff_B_x4A1eFdW1_1),.dout(w_dff_B_iue93fgv9_1),.clk(gclk));
	jdff dff_B_MFWxDZjZ4_1(.din(w_dff_B_iue93fgv9_1),.dout(w_dff_B_MFWxDZjZ4_1),.clk(gclk));
	jdff dff_B_AIGBwvCy8_1(.din(w_dff_B_MFWxDZjZ4_1),.dout(w_dff_B_AIGBwvCy8_1),.clk(gclk));
	jdff dff_B_tHIbB0nD0_1(.din(w_dff_B_AIGBwvCy8_1),.dout(w_dff_B_tHIbB0nD0_1),.clk(gclk));
	jdff dff_B_kCkRmjlp8_1(.din(n1306),.dout(w_dff_B_kCkRmjlp8_1),.clk(gclk));
	jdff dff_B_u2NDm4Ji8_1(.din(w_dff_B_kCkRmjlp8_1),.dout(w_dff_B_u2NDm4Ji8_1),.clk(gclk));
	jdff dff_B_QscYYWEd6_1(.din(w_dff_B_u2NDm4Ji8_1),.dout(w_dff_B_QscYYWEd6_1),.clk(gclk));
	jdff dff_B_yIrNcaTs8_1(.din(w_dff_B_QscYYWEd6_1),.dout(w_dff_B_yIrNcaTs8_1),.clk(gclk));
	jdff dff_B_2Clwai8F5_1(.din(w_dff_B_yIrNcaTs8_1),.dout(w_dff_B_2Clwai8F5_1),.clk(gclk));
	jdff dff_B_TnMGmJki1_1(.din(w_dff_B_2Clwai8F5_1),.dout(w_dff_B_TnMGmJki1_1),.clk(gclk));
	jdff dff_B_uvmzdZ8J0_1(.din(w_dff_B_TnMGmJki1_1),.dout(w_dff_B_uvmzdZ8J0_1),.clk(gclk));
	jdff dff_B_NhtVaw2U4_1(.din(w_dff_B_uvmzdZ8J0_1),.dout(w_dff_B_NhtVaw2U4_1),.clk(gclk));
	jdff dff_B_yX9Qr8n53_1(.din(w_dff_B_NhtVaw2U4_1),.dout(w_dff_B_yX9Qr8n53_1),.clk(gclk));
	jdff dff_B_xOVJDA0A4_1(.din(w_dff_B_yX9Qr8n53_1),.dout(w_dff_B_xOVJDA0A4_1),.clk(gclk));
	jdff dff_B_CF214jRL6_1(.din(w_dff_B_xOVJDA0A4_1),.dout(w_dff_B_CF214jRL6_1),.clk(gclk));
	jdff dff_B_xNzka8Gs5_1(.din(w_dff_B_CF214jRL6_1),.dout(w_dff_B_xNzka8Gs5_1),.clk(gclk));
	jdff dff_B_U0u26TLn6_1(.din(w_dff_B_xNzka8Gs5_1),.dout(w_dff_B_U0u26TLn6_1),.clk(gclk));
	jdff dff_B_pUClwu2V7_1(.din(w_dff_B_U0u26TLn6_1),.dout(w_dff_B_pUClwu2V7_1),.clk(gclk));
	jdff dff_B_CazNRacx3_1(.din(w_dff_B_pUClwu2V7_1),.dout(w_dff_B_CazNRacx3_1),.clk(gclk));
	jdff dff_B_bxQZ3oYx8_1(.din(w_dff_B_CazNRacx3_1),.dout(w_dff_B_bxQZ3oYx8_1),.clk(gclk));
	jdff dff_B_nTwStTD28_1(.din(w_dff_B_bxQZ3oYx8_1),.dout(w_dff_B_nTwStTD28_1),.clk(gclk));
	jdff dff_B_zsWtJ7c32_1(.din(w_dff_B_nTwStTD28_1),.dout(w_dff_B_zsWtJ7c32_1),.clk(gclk));
	jdff dff_B_Lf3YjB8x2_1(.din(w_dff_B_zsWtJ7c32_1),.dout(w_dff_B_Lf3YjB8x2_1),.clk(gclk));
	jdff dff_B_o5iXYbXe4_1(.din(w_dff_B_Lf3YjB8x2_1),.dout(w_dff_B_o5iXYbXe4_1),.clk(gclk));
	jdff dff_B_uMs40pPp2_1(.din(w_dff_B_o5iXYbXe4_1),.dout(w_dff_B_uMs40pPp2_1),.clk(gclk));
	jdff dff_A_5PzhnG0g9_0(.dout(w_n1307_0[0]),.din(w_dff_A_5PzhnG0g9_0),.clk(gclk));
	jdff dff_B_G2sRD8PB5_2(.din(n1307),.dout(w_dff_B_G2sRD8PB5_2),.clk(gclk));
	jdff dff_B_4pyoJNWl4_2(.din(w_dff_B_G2sRD8PB5_2),.dout(w_dff_B_4pyoJNWl4_2),.clk(gclk));
	jdff dff_B_qjv0Lg5Z6_2(.din(w_dff_B_4pyoJNWl4_2),.dout(w_dff_B_qjv0Lg5Z6_2),.clk(gclk));
	jdff dff_B_3MkCsW2U8_2(.din(w_dff_B_qjv0Lg5Z6_2),.dout(w_dff_B_3MkCsW2U8_2),.clk(gclk));
	jdff dff_B_kQ10nz9p1_2(.din(w_dff_B_3MkCsW2U8_2),.dout(w_dff_B_kQ10nz9p1_2),.clk(gclk));
	jdff dff_B_1TB3yJBA4_2(.din(w_dff_B_kQ10nz9p1_2),.dout(w_dff_B_1TB3yJBA4_2),.clk(gclk));
	jdff dff_B_0cVblnQ83_2(.din(w_dff_B_1TB3yJBA4_2),.dout(w_dff_B_0cVblnQ83_2),.clk(gclk));
	jdff dff_B_mqZiUbpZ1_2(.din(w_dff_B_0cVblnQ83_2),.dout(w_dff_B_mqZiUbpZ1_2),.clk(gclk));
	jdff dff_B_zfdWl9Zc2_2(.din(w_dff_B_mqZiUbpZ1_2),.dout(w_dff_B_zfdWl9Zc2_2),.clk(gclk));
	jdff dff_B_a08hvitt5_2(.din(w_dff_B_zfdWl9Zc2_2),.dout(w_dff_B_a08hvitt5_2),.clk(gclk));
	jdff dff_B_YKOnaPrb3_2(.din(w_dff_B_a08hvitt5_2),.dout(w_dff_B_YKOnaPrb3_2),.clk(gclk));
	jdff dff_B_vnqouHvk9_2(.din(w_dff_B_YKOnaPrb3_2),.dout(w_dff_B_vnqouHvk9_2),.clk(gclk));
	jdff dff_B_FHxVOqjL8_2(.din(w_dff_B_vnqouHvk9_2),.dout(w_dff_B_FHxVOqjL8_2),.clk(gclk));
	jdff dff_B_JAcY4Fv07_2(.din(w_dff_B_FHxVOqjL8_2),.dout(w_dff_B_JAcY4Fv07_2),.clk(gclk));
	jdff dff_B_PK82reXo3_2(.din(w_dff_B_JAcY4Fv07_2),.dout(w_dff_B_PK82reXo3_2),.clk(gclk));
	jdff dff_B_NM65Ng3H3_2(.din(w_dff_B_PK82reXo3_2),.dout(w_dff_B_NM65Ng3H3_2),.clk(gclk));
	jdff dff_B_BVVFdk8K6_2(.din(w_dff_B_NM65Ng3H3_2),.dout(w_dff_B_BVVFdk8K6_2),.clk(gclk));
	jdff dff_B_YG7X9TBI8_2(.din(w_dff_B_BVVFdk8K6_2),.dout(w_dff_B_YG7X9TBI8_2),.clk(gclk));
	jdff dff_B_GtGNpjkY6_0(.din(n1490),.dout(w_dff_B_GtGNpjkY6_0),.clk(gclk));
	jdff dff_B_MksgHUwL4_0(.din(w_dff_B_GtGNpjkY6_0),.dout(w_dff_B_MksgHUwL4_0),.clk(gclk));
	jdff dff_B_prF0gspV3_0(.din(w_dff_B_MksgHUwL4_0),.dout(w_dff_B_prF0gspV3_0),.clk(gclk));
	jdff dff_B_hYk4TRTn1_0(.din(w_dff_B_prF0gspV3_0),.dout(w_dff_B_hYk4TRTn1_0),.clk(gclk));
	jdff dff_B_aBFwM9Tn0_0(.din(w_dff_B_hYk4TRTn1_0),.dout(w_dff_B_aBFwM9Tn0_0),.clk(gclk));
	jdff dff_B_Le84nWLh8_0(.din(w_dff_B_aBFwM9Tn0_0),.dout(w_dff_B_Le84nWLh8_0),.clk(gclk));
	jdff dff_B_zRQ6A17J5_0(.din(w_dff_B_Le84nWLh8_0),.dout(w_dff_B_zRQ6A17J5_0),.clk(gclk));
	jdff dff_B_3apr6BjE8_0(.din(w_dff_B_zRQ6A17J5_0),.dout(w_dff_B_3apr6BjE8_0),.clk(gclk));
	jdff dff_B_tZ7XdPbV2_0(.din(w_dff_B_3apr6BjE8_0),.dout(w_dff_B_tZ7XdPbV2_0),.clk(gclk));
	jdff dff_B_wyiDseBh1_0(.din(w_dff_B_tZ7XdPbV2_0),.dout(w_dff_B_wyiDseBh1_0),.clk(gclk));
	jdff dff_B_94EGorVZ2_0(.din(w_dff_B_wyiDseBh1_0),.dout(w_dff_B_94EGorVZ2_0),.clk(gclk));
	jdff dff_B_7RpELD2L9_0(.din(w_dff_B_94EGorVZ2_0),.dout(w_dff_B_7RpELD2L9_0),.clk(gclk));
	jdff dff_B_g4GfoDlH0_0(.din(w_dff_B_7RpELD2L9_0),.dout(w_dff_B_g4GfoDlH0_0),.clk(gclk));
	jdff dff_B_tUEC23Bw2_0(.din(w_dff_B_g4GfoDlH0_0),.dout(w_dff_B_tUEC23Bw2_0),.clk(gclk));
	jdff dff_B_LWWXeHGo1_0(.din(w_dff_B_tUEC23Bw2_0),.dout(w_dff_B_LWWXeHGo1_0),.clk(gclk));
	jdff dff_B_fdGn16v56_0(.din(w_dff_B_LWWXeHGo1_0),.dout(w_dff_B_fdGn16v56_0),.clk(gclk));
	jdff dff_B_vE0mNmXg8_0(.din(w_dff_B_fdGn16v56_0),.dout(w_dff_B_vE0mNmXg8_0),.clk(gclk));
	jdff dff_B_QVuiiY506_0(.din(w_dff_B_vE0mNmXg8_0),.dout(w_dff_B_QVuiiY506_0),.clk(gclk));
	jdff dff_B_SWav6wUL2_0(.din(w_dff_B_QVuiiY506_0),.dout(w_dff_B_SWav6wUL2_0),.clk(gclk));
	jdff dff_B_2jcijqAw9_0(.din(w_dff_B_SWav6wUL2_0),.dout(w_dff_B_2jcijqAw9_0),.clk(gclk));
	jdff dff_B_icxVN9Xl1_0(.din(w_dff_B_2jcijqAw9_0),.dout(w_dff_B_icxVN9Xl1_0),.clk(gclk));
	jdff dff_B_rEnROenV5_0(.din(n1488),.dout(w_dff_B_rEnROenV5_0),.clk(gclk));
	jdff dff_B_g9ZzwNWj2_0(.din(w_dff_B_rEnROenV5_0),.dout(w_dff_B_g9ZzwNWj2_0),.clk(gclk));
	jdff dff_B_U9Uof8Zi7_0(.din(w_dff_B_g9ZzwNWj2_0),.dout(w_dff_B_U9Uof8Zi7_0),.clk(gclk));
	jdff dff_B_aJjHLNgA8_0(.din(n1487),.dout(w_dff_B_aJjHLNgA8_0),.clk(gclk));
	jdff dff_B_NbkvPVtR2_0(.din(w_dff_B_aJjHLNgA8_0),.dout(w_dff_B_NbkvPVtR2_0),.clk(gclk));
	jdff dff_A_95i5VaAd0_1(.dout(w_n414_0[1]),.din(w_dff_A_95i5VaAd0_1),.clk(gclk));
	jdff dff_A_2vsiFvqM0_1(.dout(w_dff_A_95i5VaAd0_1),.din(w_dff_A_2vsiFvqM0_1),.clk(gclk));
	jdff dff_A_2x4lTKbJ3_1(.dout(w_dff_A_2vsiFvqM0_1),.din(w_dff_A_2x4lTKbJ3_1),.clk(gclk));
	jdff dff_A_lxuxghtD1_1(.dout(w_dff_A_2x4lTKbJ3_1),.din(w_dff_A_lxuxghtD1_1),.clk(gclk));
	jdff dff_A_c5R14jvO5_1(.dout(w_dff_A_lxuxghtD1_1),.din(w_dff_A_c5R14jvO5_1),.clk(gclk));
	jdff dff_A_6E9jmO564_1(.dout(w_dff_A_c5R14jvO5_1),.din(w_dff_A_6E9jmO564_1),.clk(gclk));
	jdff dff_A_6kuqJZYv6_1(.dout(w_dff_A_6E9jmO564_1),.din(w_dff_A_6kuqJZYv6_1),.clk(gclk));
	jdff dff_A_drh3cEUA6_1(.dout(w_dff_A_6kuqJZYv6_1),.din(w_dff_A_drh3cEUA6_1),.clk(gclk));
	jdff dff_B_ekGaqtbt1_1(.din(n1482),.dout(w_dff_B_ekGaqtbt1_1),.clk(gclk));
	jdff dff_B_em3F549f2_1(.din(w_dff_B_ekGaqtbt1_1),.dout(w_dff_B_em3F549f2_1),.clk(gclk));
	jdff dff_A_OOfnODKZ7_1(.dout(w_n1370_0[1]),.din(w_dff_A_OOfnODKZ7_1),.clk(gclk));
	jdff dff_A_PbHA0OyO1_1(.dout(w_dff_A_OOfnODKZ7_1),.din(w_dff_A_PbHA0OyO1_1),.clk(gclk));
	jdff dff_A_ii7swT7v9_1(.dout(w_dff_A_PbHA0OyO1_1),.din(w_dff_A_ii7swT7v9_1),.clk(gclk));
	jdff dff_A_ojVSGgJo3_1(.dout(w_dff_A_ii7swT7v9_1),.din(w_dff_A_ojVSGgJo3_1),.clk(gclk));
	jdff dff_A_KuaHP4KI2_1(.dout(w_dff_A_ojVSGgJo3_1),.din(w_dff_A_KuaHP4KI2_1),.clk(gclk));
	jdff dff_A_EKFCEww64_1(.dout(w_dff_A_KuaHP4KI2_1),.din(w_dff_A_EKFCEww64_1),.clk(gclk));
	jdff dff_A_n05DZqeF9_1(.dout(w_dff_A_EKFCEww64_1),.din(w_dff_A_n05DZqeF9_1),.clk(gclk));
	jdff dff_A_1mhXccgt4_1(.dout(w_dff_A_n05DZqeF9_1),.din(w_dff_A_1mhXccgt4_1),.clk(gclk));
	jdff dff_A_sb2m2DnT4_1(.dout(w_dff_A_1mhXccgt4_1),.din(w_dff_A_sb2m2DnT4_1),.clk(gclk));
	jdff dff_A_gEWU635e2_1(.dout(w_dff_A_sb2m2DnT4_1),.din(w_dff_A_gEWU635e2_1),.clk(gclk));
	jdff dff_A_FMnkG7ba4_1(.dout(w_dff_A_gEWU635e2_1),.din(w_dff_A_FMnkG7ba4_1),.clk(gclk));
	jdff dff_A_yYzzaMCv0_1(.dout(w_dff_A_FMnkG7ba4_1),.din(w_dff_A_yYzzaMCv0_1),.clk(gclk));
	jdff dff_A_o5MYQtDW6_1(.dout(w_dff_A_yYzzaMCv0_1),.din(w_dff_A_o5MYQtDW6_1),.clk(gclk));
	jdff dff_A_eO6sFnFc8_1(.dout(w_dff_A_o5MYQtDW6_1),.din(w_dff_A_eO6sFnFc8_1),.clk(gclk));
	jdff dff_A_JcHFkQZf7_1(.dout(w_dff_A_eO6sFnFc8_1),.din(w_dff_A_JcHFkQZf7_1),.clk(gclk));
	jdff dff_A_FFasYZI84_1(.dout(w_dff_A_JcHFkQZf7_1),.din(w_dff_A_FFasYZI84_1),.clk(gclk));
	jdff dff_A_8QdHh2Jl3_1(.dout(w_dff_A_FFasYZI84_1),.din(w_dff_A_8QdHh2Jl3_1),.clk(gclk));
	jdff dff_A_RA75SVgC6_1(.dout(w_dff_A_8QdHh2Jl3_1),.din(w_dff_A_RA75SVgC6_1),.clk(gclk));
	jdff dff_A_eLsNsyci3_1(.dout(w_dff_A_RA75SVgC6_1),.din(w_dff_A_eLsNsyci3_1),.clk(gclk));
	jdff dff_A_ZAfiIHrD6_1(.dout(w_dff_A_eLsNsyci3_1),.din(w_dff_A_ZAfiIHrD6_1),.clk(gclk));
	jdff dff_A_mU4icPyt6_1(.dout(w_dff_A_ZAfiIHrD6_1),.din(w_dff_A_mU4icPyt6_1),.clk(gclk));
	jdff dff_A_Hk5LcA3I3_1(.dout(w_dff_A_mU4icPyt6_1),.din(w_dff_A_Hk5LcA3I3_1),.clk(gclk));
	jdff dff_A_OLArNwdu6_1(.dout(w_dff_A_Hk5LcA3I3_1),.din(w_dff_A_OLArNwdu6_1),.clk(gclk));
	jdff dff_A_450TeNIi1_1(.dout(w_dff_A_OLArNwdu6_1),.din(w_dff_A_450TeNIi1_1),.clk(gclk));
	jdff dff_A_448yc5vn0_1(.dout(w_dff_A_450TeNIi1_1),.din(w_dff_A_448yc5vn0_1),.clk(gclk));
	jdff dff_A_WzubKg2U0_1(.dout(w_dff_A_448yc5vn0_1),.din(w_dff_A_WzubKg2U0_1),.clk(gclk));
	jdff dff_A_2DXACgZw7_1(.dout(w_dff_A_WzubKg2U0_1),.din(w_dff_A_2DXACgZw7_1),.clk(gclk));
	jdff dff_A_BCmgUvh55_1(.dout(w_dff_A_2DXACgZw7_1),.din(w_dff_A_BCmgUvh55_1),.clk(gclk));
	jdff dff_B_6BwQGnYJ8_2(.din(n1370),.dout(w_dff_B_6BwQGnYJ8_2),.clk(gclk));
	jdff dff_B_5rJKp6IJ3_2(.din(w_dff_B_6BwQGnYJ8_2),.dout(w_dff_B_5rJKp6IJ3_2),.clk(gclk));
	jdff dff_A_26WJXEW48_2(.dout(w_n411_0[2]),.din(w_dff_A_26WJXEW48_2),.clk(gclk));
	jdff dff_A_8lV63m5T9_2(.dout(w_dff_A_26WJXEW48_2),.din(w_dff_A_8lV63m5T9_2),.clk(gclk));
	jdff dff_A_Kk9NeGaH9_2(.dout(w_dff_A_8lV63m5T9_2),.din(w_dff_A_Kk9NeGaH9_2),.clk(gclk));
	jdff dff_A_Qq3bdX2w1_2(.dout(w_dff_A_Kk9NeGaH9_2),.din(w_dff_A_Qq3bdX2w1_2),.clk(gclk));
	jdff dff_A_xYp5hSQi3_2(.dout(w_dff_A_Qq3bdX2w1_2),.din(w_dff_A_xYp5hSQi3_2),.clk(gclk));
	jdff dff_A_3GavLteP2_2(.dout(w_dff_A_xYp5hSQi3_2),.din(w_dff_A_3GavLteP2_2),.clk(gclk));
	jdff dff_A_soFWozYs9_2(.dout(w_dff_A_3GavLteP2_2),.din(w_dff_A_soFWozYs9_2),.clk(gclk));
	jdff dff_A_PKlY2QPT2_2(.dout(w_dff_A_soFWozYs9_2),.din(w_dff_A_PKlY2QPT2_2),.clk(gclk));
	jdff dff_A_Eeg1FAdI2_2(.dout(w_dff_A_PKlY2QPT2_2),.din(w_dff_A_Eeg1FAdI2_2),.clk(gclk));
	jdff dff_A_ehGKBBX01_2(.dout(w_dff_A_Eeg1FAdI2_2),.din(w_dff_A_ehGKBBX01_2),.clk(gclk));
	jdff dff_A_WYxLSF3l4_2(.dout(w_dff_A_ehGKBBX01_2),.din(w_dff_A_WYxLSF3l4_2),.clk(gclk));
	jdff dff_A_qGSlH1az1_2(.dout(w_dff_A_WYxLSF3l4_2),.din(w_dff_A_qGSlH1az1_2),.clk(gclk));
	jdff dff_A_BwZ8dWmo5_2(.dout(w_dff_A_qGSlH1az1_2),.din(w_dff_A_BwZ8dWmo5_2),.clk(gclk));
	jdff dff_A_gc5Xm6gJ7_2(.dout(w_dff_A_BwZ8dWmo5_2),.din(w_dff_A_gc5Xm6gJ7_2),.clk(gclk));
	jdff dff_A_GZw4V4NJ9_2(.dout(w_dff_A_gc5Xm6gJ7_2),.din(w_dff_A_GZw4V4NJ9_2),.clk(gclk));
	jdff dff_A_11tYlTAR9_2(.dout(w_dff_A_GZw4V4NJ9_2),.din(w_dff_A_11tYlTAR9_2),.clk(gclk));
	jdff dff_A_ntvZ2byh4_2(.dout(w_dff_A_11tYlTAR9_2),.din(w_dff_A_ntvZ2byh4_2),.clk(gclk));
	jdff dff_A_PBxKXlHt8_2(.dout(w_dff_A_ntvZ2byh4_2),.din(w_dff_A_PBxKXlHt8_2),.clk(gclk));
	jdff dff_A_VxsJxqaG4_2(.dout(w_dff_A_PBxKXlHt8_2),.din(w_dff_A_VxsJxqaG4_2),.clk(gclk));
	jdff dff_A_HYr82aQo3_2(.dout(w_dff_A_VxsJxqaG4_2),.din(w_dff_A_HYr82aQo3_2),.clk(gclk));
	jdff dff_A_nMrlwQhx4_2(.dout(w_dff_A_HYr82aQo3_2),.din(w_dff_A_nMrlwQhx4_2),.clk(gclk));
	jdff dff_A_S6hBsDT89_2(.dout(w_dff_A_nMrlwQhx4_2),.din(w_dff_A_S6hBsDT89_2),.clk(gclk));
	jdff dff_A_Fb0cOCXF9_2(.dout(w_dff_A_S6hBsDT89_2),.din(w_dff_A_Fb0cOCXF9_2),.clk(gclk));
	jdff dff_B_D0gJOx8J1_1(.din(n382),.dout(w_dff_B_D0gJOx8J1_1),.clk(gclk));
	jdff dff_B_JOGLfg5g2_1(.din(w_dff_B_D0gJOx8J1_1),.dout(w_dff_B_JOGLfg5g2_1),.clk(gclk));
	jdff dff_B_QDr4lZed4_1(.din(w_dff_B_JOGLfg5g2_1),.dout(w_dff_B_QDr4lZed4_1),.clk(gclk));
	jdff dff_B_V0Nq0Ly36_1(.din(w_dff_B_QDr4lZed4_1),.dout(w_dff_B_V0Nq0Ly36_1),.clk(gclk));
	jdff dff_B_EgzQaDCc9_1(.din(n384),.dout(w_dff_B_EgzQaDCc9_1),.clk(gclk));
	jdff dff_B_NLcblhT63_1(.din(w_dff_B_EgzQaDCc9_1),.dout(w_dff_B_NLcblhT63_1),.clk(gclk));
	jdff dff_B_B0usU2pS8_1(.din(w_dff_B_NLcblhT63_1),.dout(w_dff_B_B0usU2pS8_1),.clk(gclk));
	jdff dff_B_eSJ1HwC54_1(.din(w_dff_B_B0usU2pS8_1),.dout(w_dff_B_eSJ1HwC54_1),.clk(gclk));
	jdff dff_B_K0MX5dgt9_1(.din(w_dff_B_eSJ1HwC54_1),.dout(w_dff_B_K0MX5dgt9_1),.clk(gclk));
	jdff dff_A_Auvk7I1V0_2(.dout(w_n409_0[2]),.din(w_dff_A_Auvk7I1V0_2),.clk(gclk));
	jdff dff_A_fUBhY7kh0_2(.dout(w_dff_A_Auvk7I1V0_2),.din(w_dff_A_fUBhY7kh0_2),.clk(gclk));
	jdff dff_A_Utp2DALW4_2(.dout(w_dff_A_fUBhY7kh0_2),.din(w_dff_A_Utp2DALW4_2),.clk(gclk));
	jdff dff_A_LSik3jui9_2(.dout(w_dff_A_Utp2DALW4_2),.din(w_dff_A_LSik3jui9_2),.clk(gclk));
	jdff dff_A_X1zzGqSG2_2(.dout(w_dff_A_LSik3jui9_2),.din(w_dff_A_X1zzGqSG2_2),.clk(gclk));
	jdff dff_A_GFpTUtin8_2(.dout(w_dff_A_X1zzGqSG2_2),.din(w_dff_A_GFpTUtin8_2),.clk(gclk));
	jdff dff_A_AlyYxMXm2_2(.dout(w_dff_A_GFpTUtin8_2),.din(w_dff_A_AlyYxMXm2_2),.clk(gclk));
	jdff dff_A_GbjKeSl74_2(.dout(w_dff_A_AlyYxMXm2_2),.din(w_dff_A_GbjKeSl74_2),.clk(gclk));
	jdff dff_A_gyv9OaHD0_2(.dout(w_dff_A_GbjKeSl74_2),.din(w_dff_A_gyv9OaHD0_2),.clk(gclk));
	jdff dff_A_1wuB2zG22_2(.dout(w_dff_A_gyv9OaHD0_2),.din(w_dff_A_1wuB2zG22_2),.clk(gclk));
	jdff dff_A_Qtp3fshZ6_2(.dout(w_dff_A_1wuB2zG22_2),.din(w_dff_A_Qtp3fshZ6_2),.clk(gclk));
	jdff dff_A_sYSJHyLy6_2(.dout(w_dff_A_Qtp3fshZ6_2),.din(w_dff_A_sYSJHyLy6_2),.clk(gclk));
	jdff dff_A_XNjKxdey5_2(.dout(w_dff_A_sYSJHyLy6_2),.din(w_dff_A_XNjKxdey5_2),.clk(gclk));
	jdff dff_A_wpMgTIkY9_2(.dout(w_dff_A_XNjKxdey5_2),.din(w_dff_A_wpMgTIkY9_2),.clk(gclk));
	jdff dff_A_20HUvQGN2_2(.dout(w_dff_A_wpMgTIkY9_2),.din(w_dff_A_20HUvQGN2_2),.clk(gclk));
	jdff dff_A_OKMVvEvr9_2(.dout(w_dff_A_20HUvQGN2_2),.din(w_dff_A_OKMVvEvr9_2),.clk(gclk));
	jdff dff_A_rgZNpjYs0_2(.dout(w_dff_A_OKMVvEvr9_2),.din(w_dff_A_rgZNpjYs0_2),.clk(gclk));
	jdff dff_A_7wVfDs5L1_2(.dout(w_dff_A_rgZNpjYs0_2),.din(w_dff_A_7wVfDs5L1_2),.clk(gclk));
	jdff dff_A_wSxouZwt2_2(.dout(w_dff_A_7wVfDs5L1_2),.din(w_dff_A_wSxouZwt2_2),.clk(gclk));
	jdff dff_A_YoTaRUFu5_2(.dout(w_dff_A_wSxouZwt2_2),.din(w_dff_A_YoTaRUFu5_2),.clk(gclk));
	jdff dff_A_Xph7QObS9_2(.dout(w_dff_A_YoTaRUFu5_2),.din(w_dff_A_Xph7QObS9_2),.clk(gclk));
	jdff dff_A_Dvp3fPxA5_2(.dout(w_dff_A_Xph7QObS9_2),.din(w_dff_A_Dvp3fPxA5_2),.clk(gclk));
	jdff dff_A_hkYNGdsl8_2(.dout(w_dff_A_Dvp3fPxA5_2),.din(w_dff_A_hkYNGdsl8_2),.clk(gclk));
	jdff dff_A_qBUx1Ono8_2(.dout(w_dff_A_hkYNGdsl8_2),.din(w_dff_A_qBUx1Ono8_2),.clk(gclk));
	jdff dff_A_DhCr42MS9_2(.dout(w_dff_A_qBUx1Ono8_2),.din(w_dff_A_DhCr42MS9_2),.clk(gclk));
	jdff dff_B_2gdIxIEi6_1(.din(n401),.dout(w_dff_B_2gdIxIEi6_1),.clk(gclk));
	jdff dff_A_TIdTR1mS2_0(.dout(w_n405_0[0]),.din(w_dff_A_TIdTR1mS2_0),.clk(gclk));
	jdff dff_A_w8WYQ7RD0_1(.dout(w_n405_0[1]),.din(w_dff_A_w8WYQ7RD0_1),.clk(gclk));
	jdff dff_A_y3yCDxrG6_1(.dout(w_dff_A_w8WYQ7RD0_1),.din(w_dff_A_y3yCDxrG6_1),.clk(gclk));
	jdff dff_A_RerjHRQO9_1(.dout(w_dff_A_y3yCDxrG6_1),.din(w_dff_A_RerjHRQO9_1),.clk(gclk));
	jdff dff_A_KXCRNkLg3_1(.dout(w_dff_A_RerjHRQO9_1),.din(w_dff_A_KXCRNkLg3_1),.clk(gclk));
	jdff dff_A_jBhf4Lxe5_1(.dout(w_dff_A_KXCRNkLg3_1),.din(w_dff_A_jBhf4Lxe5_1),.clk(gclk));
	jdff dff_A_OhkghTEl0_1(.dout(w_dff_A_jBhf4Lxe5_1),.din(w_dff_A_OhkghTEl0_1),.clk(gclk));
	jdff dff_A_x97otNYY5_1(.dout(w_dff_A_OhkghTEl0_1),.din(w_dff_A_x97otNYY5_1),.clk(gclk));
	jdff dff_A_zUzEgu3P4_1(.dout(w_dff_A_x97otNYY5_1),.din(w_dff_A_zUzEgu3P4_1),.clk(gclk));
	jdff dff_A_N4XDKADg7_1(.dout(w_dff_A_zUzEgu3P4_1),.din(w_dff_A_N4XDKADg7_1),.clk(gclk));
	jdff dff_A_sdnuuLMM9_1(.dout(w_dff_A_N4XDKADg7_1),.din(w_dff_A_sdnuuLMM9_1),.clk(gclk));
	jdff dff_A_f3gOcPDY1_1(.dout(w_dff_A_sdnuuLMM9_1),.din(w_dff_A_f3gOcPDY1_1),.clk(gclk));
	jdff dff_A_NKn7JzbY6_1(.dout(w_dff_A_f3gOcPDY1_1),.din(w_dff_A_NKn7JzbY6_1),.clk(gclk));
	jdff dff_A_onvQ0Hb92_1(.dout(w_dff_A_NKn7JzbY6_1),.din(w_dff_A_onvQ0Hb92_1),.clk(gclk));
	jdff dff_A_eK6BNmJJ1_1(.dout(w_dff_A_onvQ0Hb92_1),.din(w_dff_A_eK6BNmJJ1_1),.clk(gclk));
	jdff dff_A_OED5NbrK0_1(.dout(w_dff_A_eK6BNmJJ1_1),.din(w_dff_A_OED5NbrK0_1),.clk(gclk));
	jdff dff_A_Y7X0RcEi9_1(.dout(w_dff_A_OED5NbrK0_1),.din(w_dff_A_Y7X0RcEi9_1),.clk(gclk));
	jdff dff_A_CWUemXRA2_1(.dout(w_dff_A_Y7X0RcEi9_1),.din(w_dff_A_CWUemXRA2_1),.clk(gclk));
	jdff dff_A_4AWYKe2d6_1(.dout(w_dff_A_CWUemXRA2_1),.din(w_dff_A_4AWYKe2d6_1),.clk(gclk));
	jdff dff_A_bfFZYIRT3_1(.dout(w_dff_A_4AWYKe2d6_1),.din(w_dff_A_bfFZYIRT3_1),.clk(gclk));
	jdff dff_A_PlTYs98K0_1(.dout(w_dff_A_bfFZYIRT3_1),.din(w_dff_A_PlTYs98K0_1),.clk(gclk));
	jdff dff_A_LRCSOgBY0_1(.dout(w_dff_A_PlTYs98K0_1),.din(w_dff_A_LRCSOgBY0_1),.clk(gclk));
	jdff dff_A_USyveyuP5_1(.dout(w_dff_A_LRCSOgBY0_1),.din(w_dff_A_USyveyuP5_1),.clk(gclk));
	jdff dff_A_rjpMRCjg1_1(.dout(w_dff_A_USyveyuP5_1),.din(w_dff_A_rjpMRCjg1_1),.clk(gclk));
	jdff dff_A_fvwy0dSg3_1(.dout(w_dff_A_rjpMRCjg1_1),.din(w_dff_A_fvwy0dSg3_1),.clk(gclk));
	jdff dff_A_HqRy27oo6_1(.dout(w_dff_A_fvwy0dSg3_1),.din(w_dff_A_HqRy27oo6_1),.clk(gclk));
	jdff dff_A_ukSRDnTv1_1(.dout(w_dff_A_HqRy27oo6_1),.din(w_dff_A_ukSRDnTv1_1),.clk(gclk));
	jdff dff_A_cDnUIF5z5_1(.dout(w_dff_A_ukSRDnTv1_1),.din(w_dff_A_cDnUIF5z5_1),.clk(gclk));
	jdff dff_A_WADLSwTz5_1(.dout(w_dff_A_cDnUIF5z5_1),.din(w_dff_A_WADLSwTz5_1),.clk(gclk));
	jdff dff_A_RpciiL6M2_1(.dout(w_dff_A_WADLSwTz5_1),.din(w_dff_A_RpciiL6M2_1),.clk(gclk));
	jdff dff_A_j8rANZNm7_1(.dout(w_dff_A_RpciiL6M2_1),.din(w_dff_A_j8rANZNm7_1),.clk(gclk));
	jdff dff_A_jYbaV7PM9_1(.dout(w_dff_A_j8rANZNm7_1),.din(w_dff_A_jYbaV7PM9_1),.clk(gclk));
	jdff dff_A_SX3eBsGe0_1(.dout(w_dff_A_jYbaV7PM9_1),.din(w_dff_A_SX3eBsGe0_1),.clk(gclk));
	jdff dff_B_6lWvEOl36_0(.din(G216),.dout(w_dff_B_6lWvEOl36_0),.clk(gclk));
	jdff dff_A_N6RBtDlV2_0(.dout(w_n393_0[0]),.din(w_dff_A_N6RBtDlV2_0),.clk(gclk));
	jdff dff_A_0ZPv1UgA1_0(.dout(w_dff_A_N6RBtDlV2_0),.din(w_dff_A_0ZPv1UgA1_0),.clk(gclk));
	jdff dff_A_h0z2qC435_1(.dout(w_n393_0[1]),.din(w_dff_A_h0z2qC435_1),.clk(gclk));
	jdff dff_A_zqEgeehC9_1(.dout(w_dff_A_h0z2qC435_1),.din(w_dff_A_zqEgeehC9_1),.clk(gclk));
	jdff dff_A_sOUMJ5Uv7_0(.dout(w_n392_0[0]),.din(w_dff_A_sOUMJ5Uv7_0),.clk(gclk));
	jdff dff_A_W7zyNWZK3_0(.dout(w_dff_A_sOUMJ5Uv7_0),.din(w_dff_A_W7zyNWZK3_0),.clk(gclk));
	jdff dff_A_76V8GQ9D3_0(.dout(w_dff_A_W7zyNWZK3_0),.din(w_dff_A_76V8GQ9D3_0),.clk(gclk));
	jdff dff_A_j9cYzXVv8_0(.dout(w_dff_A_76V8GQ9D3_0),.din(w_dff_A_j9cYzXVv8_0),.clk(gclk));
	jdff dff_A_Hs3YZ0n28_0(.dout(w_dff_A_j9cYzXVv8_0),.din(w_dff_A_Hs3YZ0n28_0),.clk(gclk));
	jdff dff_B_CaE08qKQ8_2(.din(G209),.dout(w_dff_B_CaE08qKQ8_2),.clk(gclk));
	jdff dff_A_HCOW2wxX5_0(.dout(w_n389_0[0]),.din(w_dff_A_HCOW2wxX5_0),.clk(gclk));
	jdff dff_A_sDvOWC695_0(.dout(w_dff_A_HCOW2wxX5_0),.din(w_dff_A_sDvOWC695_0),.clk(gclk));
	jdff dff_A_Mk3Y9kGR3_1(.dout(w_n389_0[1]),.din(w_dff_A_Mk3Y9kGR3_1),.clk(gclk));
	jdff dff_A_8hA8yP7X7_1(.dout(w_dff_A_Mk3Y9kGR3_1),.din(w_dff_A_8hA8yP7X7_1),.clk(gclk));
	jdff dff_A_d1f47uPV5_0(.dout(w_n388_1[0]),.din(w_dff_A_d1f47uPV5_0),.clk(gclk));
	jdff dff_A_esoiYOnO9_2(.dout(w_n388_1[2]),.din(w_dff_A_esoiYOnO9_2),.clk(gclk));
	jdff dff_A_GkomEHwd6_0(.dout(w_n377_0[0]),.din(w_dff_A_GkomEHwd6_0),.clk(gclk));
	jdff dff_A_unS6yNBJ5_0(.dout(w_dff_A_GkomEHwd6_0),.din(w_dff_A_unS6yNBJ5_0),.clk(gclk));
	jdff dff_A_K6p4i9Ny4_2(.dout(w_n377_0[2]),.din(w_dff_A_K6p4i9Ny4_2),.clk(gclk));
	jdff dff_A_NJOsFSPx2_2(.dout(w_dff_A_K6p4i9Ny4_2),.din(w_dff_A_NJOsFSPx2_2),.clk(gclk));
	jdff dff_A_bWBHz9yJ3_2(.dout(w_dff_A_NJOsFSPx2_2),.din(w_dff_A_bWBHz9yJ3_2),.clk(gclk));
	jdff dff_A_xElJ8NFB3_2(.dout(w_dff_A_bWBHz9yJ3_2),.din(w_dff_A_xElJ8NFB3_2),.clk(gclk));
	jdff dff_A_ZQmCDssD9_2(.dout(w_dff_A_xElJ8NFB3_2),.din(w_dff_A_ZQmCDssD9_2),.clk(gclk));
	jdff dff_A_SR6dHKWw2_2(.dout(w_dff_A_ZQmCDssD9_2),.din(w_dff_A_SR6dHKWw2_2),.clk(gclk));
	jdff dff_A_GJFWv1ec1_2(.dout(w_dff_A_SR6dHKWw2_2),.din(w_dff_A_GJFWv1ec1_2),.clk(gclk));
	jdff dff_A_FYbWQtoV8_0(.dout(w_n374_0[0]),.din(w_dff_A_FYbWQtoV8_0),.clk(gclk));
	jdff dff_A_MM8c0lGK3_0(.dout(w_dff_A_FYbWQtoV8_0),.din(w_dff_A_MM8c0lGK3_0),.clk(gclk));
	jdff dff_B_xc9uFfJ31_0(.din(G213),.dout(w_dff_B_xc9uFfJ31_0),.clk(gclk));
	jdff dff_A_w7Q4eY0z2_1(.dout(w_n371_0[1]),.din(w_dff_A_w7Q4eY0z2_1),.clk(gclk));
	jdff dff_A_SuyAG6dD7_1(.dout(w_dff_A_w7Q4eY0z2_1),.din(w_dff_A_SuyAG6dD7_1),.clk(gclk));
	jdff dff_A_OAyUsTmf6_2(.dout(w_n371_0[2]),.din(w_dff_A_OAyUsTmf6_2),.clk(gclk));
	jdff dff_A_Zkr9sd264_2(.dout(w_dff_A_OAyUsTmf6_2),.din(w_dff_A_Zkr9sd264_2),.clk(gclk));
	jdff dff_B_wQ2PMfI50_1(.din(n508),.dout(w_dff_B_wQ2PMfI50_1),.clk(gclk));
	jdff dff_B_rfSBHnSX5_1(.din(w_dff_B_wQ2PMfI50_1),.dout(w_dff_B_rfSBHnSX5_1),.clk(gclk));
	jdff dff_B_aCJDbkf27_1(.din(w_dff_B_rfSBHnSX5_1),.dout(w_dff_B_aCJDbkf27_1),.clk(gclk));
	jdff dff_B_15NAMZfR8_1(.din(w_dff_B_aCJDbkf27_1),.dout(w_dff_B_15NAMZfR8_1),.clk(gclk));
	jdff dff_B_ySkQdOIf1_1(.din(w_dff_B_15NAMZfR8_1),.dout(w_dff_B_ySkQdOIf1_1),.clk(gclk));
	jdff dff_B_Lz3C0pVl2_1(.din(w_dff_B_ySkQdOIf1_1),.dout(w_dff_B_Lz3C0pVl2_1),.clk(gclk));
	jdff dff_B_iKfYZPQF9_1(.din(w_dff_B_Lz3C0pVl2_1),.dout(w_dff_B_iKfYZPQF9_1),.clk(gclk));
	jdff dff_B_ln7zhQeV7_1(.din(w_dff_B_iKfYZPQF9_1),.dout(w_dff_B_ln7zhQeV7_1),.clk(gclk));
	jdff dff_B_wm5BKaSa1_1(.din(w_dff_B_ln7zhQeV7_1),.dout(w_dff_B_wm5BKaSa1_1),.clk(gclk));
	jdff dff_B_1zNhJcEm4_1(.din(w_dff_B_wm5BKaSa1_1),.dout(w_dff_B_1zNhJcEm4_1),.clk(gclk));
	jdff dff_B_dJbhAIgp7_1(.din(w_dff_B_1zNhJcEm4_1),.dout(w_dff_B_dJbhAIgp7_1),.clk(gclk));
	jdff dff_B_sdnlnBax3_1(.din(w_dff_B_dJbhAIgp7_1),.dout(w_dff_B_sdnlnBax3_1),.clk(gclk));
	jdff dff_B_wQ1lNVpq3_1(.din(w_dff_B_sdnlnBax3_1),.dout(w_dff_B_wQ1lNVpq3_1),.clk(gclk));
	jdff dff_B_lvLgAINt7_1(.din(w_dff_B_wQ1lNVpq3_1),.dout(w_dff_B_lvLgAINt7_1),.clk(gclk));
	jdff dff_B_fmePZ4cR4_1(.din(w_dff_B_lvLgAINt7_1),.dout(w_dff_B_fmePZ4cR4_1),.clk(gclk));
	jdff dff_B_SmiIqvJS0_1(.din(w_dff_B_fmePZ4cR4_1),.dout(w_dff_B_SmiIqvJS0_1),.clk(gclk));
	jdff dff_B_60ORWjGP0_1(.din(w_dff_B_SmiIqvJS0_1),.dout(w_dff_B_60ORWjGP0_1),.clk(gclk));
	jdff dff_B_RWneN9S12_1(.din(w_dff_B_60ORWjGP0_1),.dout(w_dff_B_RWneN9S12_1),.clk(gclk));
	jdff dff_B_WWYGcvMe7_1(.din(w_dff_B_RWneN9S12_1),.dout(w_dff_B_WWYGcvMe7_1),.clk(gclk));
	jdff dff_B_hmkJm5fk9_0(.din(n697),.dout(w_dff_B_hmkJm5fk9_0),.clk(gclk));
	jdff dff_B_LLCjecBY0_0(.din(w_dff_B_hmkJm5fk9_0),.dout(w_dff_B_LLCjecBY0_0),.clk(gclk));
	jdff dff_B_m4UXWIJG9_0(.din(w_dff_B_LLCjecBY0_0),.dout(w_dff_B_m4UXWIJG9_0),.clk(gclk));
	jdff dff_B_60MmKkKi2_0(.din(w_dff_B_m4UXWIJG9_0),.dout(w_dff_B_60MmKkKi2_0),.clk(gclk));
	jdff dff_B_HPyX5hiM0_0(.din(w_dff_B_60MmKkKi2_0),.dout(w_dff_B_HPyX5hiM0_0),.clk(gclk));
	jdff dff_B_DiZlY0Yg3_0(.din(w_dff_B_HPyX5hiM0_0),.dout(w_dff_B_DiZlY0Yg3_0),.clk(gclk));
	jdff dff_B_GEykmAI96_0(.din(w_dff_B_DiZlY0Yg3_0),.dout(w_dff_B_GEykmAI96_0),.clk(gclk));
	jdff dff_B_Xy1yLjEo5_0(.din(w_dff_B_GEykmAI96_0),.dout(w_dff_B_Xy1yLjEo5_0),.clk(gclk));
	jdff dff_B_yVh2irt11_0(.din(w_dff_B_Xy1yLjEo5_0),.dout(w_dff_B_yVh2irt11_0),.clk(gclk));
	jdff dff_B_Hul66GOv5_0(.din(w_dff_B_yVh2irt11_0),.dout(w_dff_B_Hul66GOv5_0),.clk(gclk));
	jdff dff_B_rbbKn9bM4_0(.din(w_dff_B_Hul66GOv5_0),.dout(w_dff_B_rbbKn9bM4_0),.clk(gclk));
	jdff dff_B_TtJHkCmy5_0(.din(w_dff_B_rbbKn9bM4_0),.dout(w_dff_B_TtJHkCmy5_0),.clk(gclk));
	jdff dff_B_EnLLDslU7_0(.din(w_dff_B_TtJHkCmy5_0),.dout(w_dff_B_EnLLDslU7_0),.clk(gclk));
	jdff dff_B_eaqtGupW1_0(.din(w_dff_B_EnLLDslU7_0),.dout(w_dff_B_eaqtGupW1_0),.clk(gclk));
	jdff dff_A_53r8eIzj3_0(.dout(w_n696_0[0]),.din(w_dff_A_53r8eIzj3_0),.clk(gclk));
	jdff dff_A_h6UuGasn2_0(.dout(w_dff_A_53r8eIzj3_0),.din(w_dff_A_h6UuGasn2_0),.clk(gclk));
	jdff dff_A_NEgK3E738_0(.dout(w_dff_A_h6UuGasn2_0),.din(w_dff_A_NEgK3E738_0),.clk(gclk));
	jdff dff_A_X1ENr5nY4_0(.dout(w_dff_A_NEgK3E738_0),.din(w_dff_A_X1ENr5nY4_0),.clk(gclk));
	jdff dff_A_BDQPPL190_0(.dout(w_dff_A_X1ENr5nY4_0),.din(w_dff_A_BDQPPL190_0),.clk(gclk));
	jdff dff_A_ejiq0jjN4_0(.dout(w_dff_A_BDQPPL190_0),.din(w_dff_A_ejiq0jjN4_0),.clk(gclk));
	jdff dff_A_UW2SCsm97_0(.dout(w_dff_A_ejiq0jjN4_0),.din(w_dff_A_UW2SCsm97_0),.clk(gclk));
	jdff dff_A_74tjy7kl5_0(.dout(w_dff_A_UW2SCsm97_0),.din(w_dff_A_74tjy7kl5_0),.clk(gclk));
	jdff dff_A_B6lVHn3M9_0(.dout(w_dff_A_74tjy7kl5_0),.din(w_dff_A_B6lVHn3M9_0),.clk(gclk));
	jdff dff_A_aDpe2EhD5_0(.dout(w_dff_A_B6lVHn3M9_0),.din(w_dff_A_aDpe2EhD5_0),.clk(gclk));
	jdff dff_A_FmcT6jx85_0(.dout(w_dff_A_aDpe2EhD5_0),.din(w_dff_A_FmcT6jx85_0),.clk(gclk));
	jdff dff_A_kO7549DR1_0(.dout(w_dff_A_FmcT6jx85_0),.din(w_dff_A_kO7549DR1_0),.clk(gclk));
	jdff dff_A_tsQ1su0p6_0(.dout(w_dff_A_kO7549DR1_0),.din(w_dff_A_tsQ1su0p6_0),.clk(gclk));
	jdff dff_A_a3tr2dka2_0(.dout(w_dff_A_tsQ1su0p6_0),.din(w_dff_A_a3tr2dka2_0),.clk(gclk));
	jdff dff_A_iQeXEwhg6_0(.dout(w_dff_A_a3tr2dka2_0),.din(w_dff_A_iQeXEwhg6_0),.clk(gclk));
	jdff dff_B_HYJttRAU5_1(.din(n688),.dout(w_dff_B_HYJttRAU5_1),.clk(gclk));
	jdff dff_B_kDrfp6vL7_1(.din(w_dff_B_HYJttRAU5_1),.dout(w_dff_B_kDrfp6vL7_1),.clk(gclk));
	jdff dff_B_gokY1vEq5_1(.din(w_dff_B_kDrfp6vL7_1),.dout(w_dff_B_gokY1vEq5_1),.clk(gclk));
	jdff dff_B_BKExFhTI0_1(.din(n519),.dout(w_dff_B_BKExFhTI0_1),.clk(gclk));
	jdff dff_B_a29utAwe0_1(.din(w_dff_B_BKExFhTI0_1),.dout(w_dff_B_a29utAwe0_1),.clk(gclk));
	jdff dff_B_rGygypLd3_1(.din(w_dff_B_a29utAwe0_1),.dout(w_dff_B_rGygypLd3_1),.clk(gclk));
	jdff dff_B_CdlzwAyf0_1(.din(w_dff_B_rGygypLd3_1),.dout(w_dff_B_CdlzwAyf0_1),.clk(gclk));
	jdff dff_B_J0VlKb5g2_1(.din(w_dff_B_CdlzwAyf0_1),.dout(w_dff_B_J0VlKb5g2_1),.clk(gclk));
	jdff dff_B_9bmPxkie9_1(.din(w_dff_B_J0VlKb5g2_1),.dout(w_dff_B_9bmPxkie9_1),.clk(gclk));
	jdff dff_B_FraTEUNL8_1(.din(w_dff_B_9bmPxkie9_1),.dout(w_dff_B_FraTEUNL8_1),.clk(gclk));
	jdff dff_B_MJ4rqQGV0_1(.din(w_dff_B_FraTEUNL8_1),.dout(w_dff_B_MJ4rqQGV0_1),.clk(gclk));
	jdff dff_B_UsLOLSfz0_1(.din(w_dff_B_MJ4rqQGV0_1),.dout(w_dff_B_UsLOLSfz0_1),.clk(gclk));
	jdff dff_B_0FtXJN2A7_1(.din(w_dff_B_UsLOLSfz0_1),.dout(w_dff_B_0FtXJN2A7_1),.clk(gclk));
	jdff dff_B_oQpbIVWX8_1(.din(w_dff_B_0FtXJN2A7_1),.dout(w_dff_B_oQpbIVWX8_1),.clk(gclk));
	jdff dff_B_K601PMIT9_1(.din(w_dff_B_oQpbIVWX8_1),.dout(w_dff_B_K601PMIT9_1),.clk(gclk));
	jdff dff_B_XxnRDXtu6_1(.din(w_dff_B_K601PMIT9_1),.dout(w_dff_B_XxnRDXtu6_1),.clk(gclk));
	jdff dff_B_LOLKaIid3_1(.din(w_dff_B_XxnRDXtu6_1),.dout(w_dff_B_LOLKaIid3_1),.clk(gclk));
	jdff dff_B_Uz1Zm8eK4_1(.din(w_dff_B_LOLKaIid3_1),.dout(w_dff_B_Uz1Zm8eK4_1),.clk(gclk));
	jdff dff_B_CtHFdiwh9_1(.din(w_dff_B_Uz1Zm8eK4_1),.dout(w_dff_B_CtHFdiwh9_1),.clk(gclk));
	jdff dff_B_mmI1cXgL2_1(.din(w_dff_B_CtHFdiwh9_1),.dout(w_dff_B_mmI1cXgL2_1),.clk(gclk));
	jdff dff_B_BLjKThjL5_1(.din(n527),.dout(w_dff_B_BLjKThjL5_1),.clk(gclk));
	jdff dff_B_gVy1CQY12_1(.din(w_dff_B_BLjKThjL5_1),.dout(w_dff_B_gVy1CQY12_1),.clk(gclk));
	jdff dff_B_ORUcWxsl2_1(.din(w_dff_B_gVy1CQY12_1),.dout(w_dff_B_ORUcWxsl2_1),.clk(gclk));
	jdff dff_B_aFFUNSsZ1_1(.din(w_dff_B_ORUcWxsl2_1),.dout(w_dff_B_aFFUNSsZ1_1),.clk(gclk));
	jdff dff_B_Ii41U4s57_1(.din(w_dff_B_aFFUNSsZ1_1),.dout(w_dff_B_Ii41U4s57_1),.clk(gclk));
	jdff dff_B_iDlq5Qbu8_1(.din(w_dff_B_Ii41U4s57_1),.dout(w_dff_B_iDlq5Qbu8_1),.clk(gclk));
	jdff dff_B_jnmVzGmV2_1(.din(w_dff_B_iDlq5Qbu8_1),.dout(w_dff_B_jnmVzGmV2_1),.clk(gclk));
	jdff dff_B_wug3JZzv1_1(.din(w_dff_B_jnmVzGmV2_1),.dout(w_dff_B_wug3JZzv1_1),.clk(gclk));
	jdff dff_B_pVU240ri1_1(.din(w_dff_B_wug3JZzv1_1),.dout(w_dff_B_pVU240ri1_1),.clk(gclk));
	jdff dff_B_PJ3UrIzK9_1(.din(w_dff_B_pVU240ri1_1),.dout(w_dff_B_PJ3UrIzK9_1),.clk(gclk));
	jdff dff_B_WC41jezt4_1(.din(w_dff_B_PJ3UrIzK9_1),.dout(w_dff_B_WC41jezt4_1),.clk(gclk));
	jdff dff_B_QMvArpxz2_1(.din(w_dff_B_WC41jezt4_1),.dout(w_dff_B_QMvArpxz2_1),.clk(gclk));
	jdff dff_B_DYUbNjOo5_1(.din(w_dff_B_QMvArpxz2_1),.dout(w_dff_B_DYUbNjOo5_1),.clk(gclk));
	jdff dff_B_W33OGnFZ9_1(.din(w_dff_B_DYUbNjOo5_1),.dout(w_dff_B_W33OGnFZ9_1),.clk(gclk));
	jdff dff_A_amAYhCsa7_1(.dout(w_n513_1[1]),.din(w_dff_A_amAYhCsa7_1),.clk(gclk));
	jdff dff_A_GpTyvR8n3_1(.dout(w_dff_A_amAYhCsa7_1),.din(w_dff_A_GpTyvR8n3_1),.clk(gclk));
	jdff dff_A_tIBXdVDf5_1(.dout(w_dff_A_GpTyvR8n3_1),.din(w_dff_A_tIBXdVDf5_1),.clk(gclk));
	jdff dff_A_UUAEIRxE0_1(.dout(w_dff_A_tIBXdVDf5_1),.din(w_dff_A_UUAEIRxE0_1),.clk(gclk));
	jdff dff_A_EqCf6LOY1_1(.dout(w_dff_A_UUAEIRxE0_1),.din(w_dff_A_EqCf6LOY1_1),.clk(gclk));
	jdff dff_A_tBMhYuYz7_1(.dout(w_dff_A_EqCf6LOY1_1),.din(w_dff_A_tBMhYuYz7_1),.clk(gclk));
	jdff dff_A_EbzSqyfX0_1(.dout(w_dff_A_tBMhYuYz7_1),.din(w_dff_A_EbzSqyfX0_1),.clk(gclk));
	jdff dff_A_o4hKN4Nk7_1(.dout(w_dff_A_EbzSqyfX0_1),.din(w_dff_A_o4hKN4Nk7_1),.clk(gclk));
	jdff dff_A_NcVEOXhi5_1(.dout(w_dff_A_o4hKN4Nk7_1),.din(w_dff_A_NcVEOXhi5_1),.clk(gclk));
	jdff dff_A_SjxkgvLG3_1(.dout(w_dff_A_NcVEOXhi5_1),.din(w_dff_A_SjxkgvLG3_1),.clk(gclk));
	jdff dff_A_LaQBvpyP2_1(.dout(w_dff_A_SjxkgvLG3_1),.din(w_dff_A_LaQBvpyP2_1),.clk(gclk));
	jdff dff_A_ouPtDqXW0_1(.dout(w_dff_A_LaQBvpyP2_1),.din(w_dff_A_ouPtDqXW0_1),.clk(gclk));
	jdff dff_A_UgnEGHoV7_1(.dout(w_dff_A_ouPtDqXW0_1),.din(w_dff_A_UgnEGHoV7_1),.clk(gclk));
	jdff dff_A_RfMCjFwd9_1(.dout(w_dff_A_UgnEGHoV7_1),.din(w_dff_A_RfMCjFwd9_1),.clk(gclk));
	jdff dff_A_OkbB5HG98_1(.dout(w_dff_A_RfMCjFwd9_1),.din(w_dff_A_OkbB5HG98_1),.clk(gclk));
	jdff dff_A_jBLPjwIz9_1(.dout(w_dff_A_OkbB5HG98_1),.din(w_dff_A_jBLPjwIz9_1),.clk(gclk));
	jdff dff_A_jhMpSaWM5_1(.dout(w_dff_A_jBLPjwIz9_1),.din(w_dff_A_jhMpSaWM5_1),.clk(gclk));
	jdff dff_A_SsTPKTdV9_1(.dout(w_dff_A_jhMpSaWM5_1),.din(w_dff_A_SsTPKTdV9_1),.clk(gclk));
	jdff dff_A_cC4jDxwZ0_1(.dout(w_dff_A_SsTPKTdV9_1),.din(w_dff_A_cC4jDxwZ0_1),.clk(gclk));
	jdff dff_A_wrJvwDwI0_0(.dout(w_n507_0[0]),.din(w_dff_A_wrJvwDwI0_0),.clk(gclk));
	jdff dff_A_MOh5qngo9_0(.dout(w_dff_A_wrJvwDwI0_0),.din(w_dff_A_MOh5qngo9_0),.clk(gclk));
	jdff dff_A_W5BhSzPy5_0(.dout(w_dff_A_MOh5qngo9_0),.din(w_dff_A_W5BhSzPy5_0),.clk(gclk));
	jdff dff_A_IADBaKt47_0(.dout(w_dff_A_W5BhSzPy5_0),.din(w_dff_A_IADBaKt47_0),.clk(gclk));
	jdff dff_A_Klcoe3uJ0_0(.dout(w_dff_A_IADBaKt47_0),.din(w_dff_A_Klcoe3uJ0_0),.clk(gclk));
	jdff dff_A_PL2uC0MR5_0(.dout(w_dff_A_Klcoe3uJ0_0),.din(w_dff_A_PL2uC0MR5_0),.clk(gclk));
	jdff dff_A_edNij6l28_0(.dout(w_dff_A_PL2uC0MR5_0),.din(w_dff_A_edNij6l28_0),.clk(gclk));
	jdff dff_A_Xr05sfnV4_0(.dout(w_dff_A_edNij6l28_0),.din(w_dff_A_Xr05sfnV4_0),.clk(gclk));
	jdff dff_A_bABSf4G24_0(.dout(w_dff_A_Xr05sfnV4_0),.din(w_dff_A_bABSf4G24_0),.clk(gclk));
	jdff dff_A_X09YGMTN7_0(.dout(w_dff_A_bABSf4G24_0),.din(w_dff_A_X09YGMTN7_0),.clk(gclk));
	jdff dff_A_k30zt85Z7_0(.dout(w_dff_A_X09YGMTN7_0),.din(w_dff_A_k30zt85Z7_0),.clk(gclk));
	jdff dff_A_5t6lLZ050_0(.dout(w_dff_A_k30zt85Z7_0),.din(w_dff_A_5t6lLZ050_0),.clk(gclk));
	jdff dff_A_Bcu7KTF06_0(.dout(w_dff_A_5t6lLZ050_0),.din(w_dff_A_Bcu7KTF06_0),.clk(gclk));
	jdff dff_A_DbDF4rQJ7_0(.dout(w_dff_A_Bcu7KTF06_0),.din(w_dff_A_DbDF4rQJ7_0),.clk(gclk));
	jdff dff_A_xSbZG5Ba2_0(.dout(w_dff_A_DbDF4rQJ7_0),.din(w_dff_A_xSbZG5Ba2_0),.clk(gclk));
	jdff dff_A_hdv4s7Pz1_0(.dout(w_dff_A_xSbZG5Ba2_0),.din(w_dff_A_hdv4s7Pz1_0),.clk(gclk));
	jdff dff_A_XiWMazXS0_0(.dout(w_dff_A_hdv4s7Pz1_0),.din(w_dff_A_XiWMazXS0_0),.clk(gclk));
	jdff dff_A_FNKjGO625_0(.dout(w_dff_A_XiWMazXS0_0),.din(w_dff_A_FNKjGO625_0),.clk(gclk));
	jdff dff_A_T6Ux1lWC6_0(.dout(w_dff_A_FNKjGO625_0),.din(w_dff_A_T6Ux1lWC6_0),.clk(gclk));
	jdff dff_A_aJryGNPj1_0(.dout(w_dff_A_T6Ux1lWC6_0),.din(w_dff_A_aJryGNPj1_0),.clk(gclk));
	jdff dff_A_gNaQHZmM1_1(.dout(w_n505_0[1]),.din(w_dff_A_gNaQHZmM1_1),.clk(gclk));
	jdff dff_A_xuIBbaxg9_1(.dout(w_dff_A_gNaQHZmM1_1),.din(w_dff_A_xuIBbaxg9_1),.clk(gclk));
	jdff dff_A_kxZRG5zq2_1(.dout(w_dff_A_xuIBbaxg9_1),.din(w_dff_A_kxZRG5zq2_1),.clk(gclk));
	jdff dff_A_QdAeCn2i2_1(.dout(w_dff_A_kxZRG5zq2_1),.din(w_dff_A_QdAeCn2i2_1),.clk(gclk));
	jdff dff_A_BcsaBom17_1(.dout(w_dff_A_QdAeCn2i2_1),.din(w_dff_A_BcsaBom17_1),.clk(gclk));
	jdff dff_A_gODWlgmR5_1(.dout(w_dff_A_BcsaBom17_1),.din(w_dff_A_gODWlgmR5_1),.clk(gclk));
	jdff dff_A_3JcRLIeR3_1(.dout(w_dff_A_gODWlgmR5_1),.din(w_dff_A_3JcRLIeR3_1),.clk(gclk));
	jdff dff_A_faKNPZ6T9_1(.dout(w_dff_A_3JcRLIeR3_1),.din(w_dff_A_faKNPZ6T9_1),.clk(gclk));
	jdff dff_A_ANRzoikc5_1(.dout(w_dff_A_faKNPZ6T9_1),.din(w_dff_A_ANRzoikc5_1),.clk(gclk));
	jdff dff_A_Kh3lZXq61_1(.dout(w_dff_A_ANRzoikc5_1),.din(w_dff_A_Kh3lZXq61_1),.clk(gclk));
	jdff dff_A_3c3ITUf51_1(.dout(w_dff_A_Kh3lZXq61_1),.din(w_dff_A_3c3ITUf51_1),.clk(gclk));
	jdff dff_A_GaVM0qnd6_1(.dout(w_dff_A_3c3ITUf51_1),.din(w_dff_A_GaVM0qnd6_1),.clk(gclk));
	jdff dff_A_lNJnqCOM6_1(.dout(w_dff_A_GaVM0qnd6_1),.din(w_dff_A_lNJnqCOM6_1),.clk(gclk));
	jdff dff_A_JRCDhjtx9_1(.dout(w_dff_A_lNJnqCOM6_1),.din(w_dff_A_JRCDhjtx9_1),.clk(gclk));
	jdff dff_A_cDo7qvmm0_1(.dout(w_dff_A_JRCDhjtx9_1),.din(w_dff_A_cDo7qvmm0_1),.clk(gclk));
	jdff dff_A_ZAEKEhuG8_1(.dout(w_dff_A_cDo7qvmm0_1),.din(w_dff_A_ZAEKEhuG8_1),.clk(gclk));
	jdff dff_A_WMbwGSev8_1(.dout(w_dff_A_ZAEKEhuG8_1),.din(w_dff_A_WMbwGSev8_1),.clk(gclk));
	jdff dff_A_PrlsKesa0_1(.dout(w_dff_A_WMbwGSev8_1),.din(w_dff_A_PrlsKesa0_1),.clk(gclk));
	jdff dff_A_h6i8hGZv5_1(.dout(w_dff_A_PrlsKesa0_1),.din(w_dff_A_h6i8hGZv5_1),.clk(gclk));
	jdff dff_A_RGcGofez3_1(.dout(w_dff_A_h6i8hGZv5_1),.din(w_dff_A_RGcGofez3_1),.clk(gclk));
	jdff dff_A_BopCeC6t1_1(.dout(w_dff_A_RGcGofez3_1),.din(w_dff_A_BopCeC6t1_1),.clk(gclk));
	jdff dff_A_xavBH0ie1_1(.dout(w_dff_A_BopCeC6t1_1),.din(w_dff_A_xavBH0ie1_1),.clk(gclk));
	jdff dff_A_aB5MWU2t6_1(.dout(w_n500_0[1]),.din(w_dff_A_aB5MWU2t6_1),.clk(gclk));
	jdff dff_A_NoNtTVNC3_1(.dout(w_dff_A_aB5MWU2t6_1),.din(w_dff_A_NoNtTVNC3_1),.clk(gclk));
	jdff dff_A_tcdEHWon4_1(.dout(w_dff_A_NoNtTVNC3_1),.din(w_dff_A_tcdEHWon4_1),.clk(gclk));
	jdff dff_A_lSrIxcek8_1(.dout(w_dff_A_tcdEHWon4_1),.din(w_dff_A_lSrIxcek8_1),.clk(gclk));
	jdff dff_A_Ih3zeL8h5_1(.dout(w_dff_A_lSrIxcek8_1),.din(w_dff_A_Ih3zeL8h5_1),.clk(gclk));
	jdff dff_A_oJjRbQZT4_1(.dout(w_dff_A_Ih3zeL8h5_1),.din(w_dff_A_oJjRbQZT4_1),.clk(gclk));
	jdff dff_A_MnWO2fIl3_1(.dout(w_dff_A_oJjRbQZT4_1),.din(w_dff_A_MnWO2fIl3_1),.clk(gclk));
	jdff dff_A_TO7YJ9K24_1(.dout(w_dff_A_MnWO2fIl3_1),.din(w_dff_A_TO7YJ9K24_1),.clk(gclk));
	jdff dff_A_CxsKsmNL5_1(.dout(w_dff_A_TO7YJ9K24_1),.din(w_dff_A_CxsKsmNL5_1),.clk(gclk));
	jdff dff_A_p53AzdjF4_1(.dout(w_dff_A_CxsKsmNL5_1),.din(w_dff_A_p53AzdjF4_1),.clk(gclk));
	jdff dff_A_JCFtJ09t4_1(.dout(w_dff_A_p53AzdjF4_1),.din(w_dff_A_JCFtJ09t4_1),.clk(gclk));
	jdff dff_A_tIeBY7ZP5_1(.dout(w_dff_A_JCFtJ09t4_1),.din(w_dff_A_tIeBY7ZP5_1),.clk(gclk));
	jdff dff_A_Y1AugM6I4_1(.dout(w_dff_A_tIeBY7ZP5_1),.din(w_dff_A_Y1AugM6I4_1),.clk(gclk));
	jdff dff_A_Rus3fZtn4_1(.dout(w_dff_A_Y1AugM6I4_1),.din(w_dff_A_Rus3fZtn4_1),.clk(gclk));
	jdff dff_A_38b6xME91_1(.dout(w_dff_A_Rus3fZtn4_1),.din(w_dff_A_38b6xME91_1),.clk(gclk));
	jdff dff_A_3boJ5GZc9_1(.dout(w_dff_A_38b6xME91_1),.din(w_dff_A_3boJ5GZc9_1),.clk(gclk));
	jdff dff_A_bOSuo1ok3_1(.dout(w_dff_A_3boJ5GZc9_1),.din(w_dff_A_bOSuo1ok3_1),.clk(gclk));
	jdff dff_A_DKf7sUZJ4_1(.dout(w_dff_A_bOSuo1ok3_1),.din(w_dff_A_DKf7sUZJ4_1),.clk(gclk));
	jdff dff_A_w2kgbuby9_1(.dout(w_n499_0[1]),.din(w_dff_A_w2kgbuby9_1),.clk(gclk));
	jdff dff_A_cy97yl1b8_1(.dout(w_dff_A_w2kgbuby9_1),.din(w_dff_A_cy97yl1b8_1),.clk(gclk));
	jdff dff_A_TKdoqjWU0_1(.dout(w_dff_A_cy97yl1b8_1),.din(w_dff_A_TKdoqjWU0_1),.clk(gclk));
	jdff dff_A_CuFBcBUB5_1(.dout(w_dff_A_TKdoqjWU0_1),.din(w_dff_A_CuFBcBUB5_1),.clk(gclk));
	jdff dff_A_m61EdLbR0_1(.dout(w_dff_A_CuFBcBUB5_1),.din(w_dff_A_m61EdLbR0_1),.clk(gclk));
	jdff dff_A_uxma2TSc2_1(.dout(w_dff_A_m61EdLbR0_1),.din(w_dff_A_uxma2TSc2_1),.clk(gclk));
	jdff dff_A_YvnfCmG75_1(.dout(w_dff_A_uxma2TSc2_1),.din(w_dff_A_YvnfCmG75_1),.clk(gclk));
	jdff dff_A_n1su2Csh1_1(.dout(w_dff_A_YvnfCmG75_1),.din(w_dff_A_n1su2Csh1_1),.clk(gclk));
	jdff dff_A_p0RGQNFY8_1(.dout(w_dff_A_n1su2Csh1_1),.din(w_dff_A_p0RGQNFY8_1),.clk(gclk));
	jdff dff_A_xt7GjEEB2_1(.dout(w_dff_A_p0RGQNFY8_1),.din(w_dff_A_xt7GjEEB2_1),.clk(gclk));
	jdff dff_A_tAXEGNpo0_1(.dout(w_dff_A_xt7GjEEB2_1),.din(w_dff_A_tAXEGNpo0_1),.clk(gclk));
	jdff dff_A_9Jayynfx4_1(.dout(w_dff_A_tAXEGNpo0_1),.din(w_dff_A_9Jayynfx4_1),.clk(gclk));
	jdff dff_A_RhW9o69O3_1(.dout(w_dff_A_9Jayynfx4_1),.din(w_dff_A_RhW9o69O3_1),.clk(gclk));
	jdff dff_A_1RskFi178_1(.dout(w_dff_A_RhW9o69O3_1),.din(w_dff_A_1RskFi178_1),.clk(gclk));
	jdff dff_A_N7mi49Vo4_1(.dout(w_dff_A_1RskFi178_1),.din(w_dff_A_N7mi49Vo4_1),.clk(gclk));
	jdff dff_A_VbIRRRyl1_1(.dout(w_dff_A_N7mi49Vo4_1),.din(w_dff_A_VbIRRRyl1_1),.clk(gclk));
	jdff dff_A_msWSaFgt3_1(.dout(w_dff_A_VbIRRRyl1_1),.din(w_dff_A_msWSaFgt3_1),.clk(gclk));
	jdff dff_A_Aak0B7AL6_0(.dout(w_n497_1[0]),.din(w_dff_A_Aak0B7AL6_0),.clk(gclk));
	jdff dff_A_P05SiyRm0_0(.dout(w_dff_A_Aak0B7AL6_0),.din(w_dff_A_P05SiyRm0_0),.clk(gclk));
	jdff dff_A_R0djuMDo8_0(.dout(w_dff_A_P05SiyRm0_0),.din(w_dff_A_R0djuMDo8_0),.clk(gclk));
	jdff dff_A_ZK73vVpY6_0(.dout(w_dff_A_R0djuMDo8_0),.din(w_dff_A_ZK73vVpY6_0),.clk(gclk));
	jdff dff_A_Kw7ugb9f3_0(.dout(w_dff_A_ZK73vVpY6_0),.din(w_dff_A_Kw7ugb9f3_0),.clk(gclk));
	jdff dff_A_HeY7sfu61_0(.dout(w_dff_A_Kw7ugb9f3_0),.din(w_dff_A_HeY7sfu61_0),.clk(gclk));
	jdff dff_A_m2ZkOJmp7_0(.dout(w_dff_A_HeY7sfu61_0),.din(w_dff_A_m2ZkOJmp7_0),.clk(gclk));
	jdff dff_A_cCxWXWnh5_0(.dout(w_dff_A_m2ZkOJmp7_0),.din(w_dff_A_cCxWXWnh5_0),.clk(gclk));
	jdff dff_A_lVYM9zJJ2_0(.dout(w_dff_A_cCxWXWnh5_0),.din(w_dff_A_lVYM9zJJ2_0),.clk(gclk));
	jdff dff_A_kq8E1F326_0(.dout(w_dff_A_lVYM9zJJ2_0),.din(w_dff_A_kq8E1F326_0),.clk(gclk));
	jdff dff_A_9te5rlwh6_0(.dout(w_dff_A_kq8E1F326_0),.din(w_dff_A_9te5rlwh6_0),.clk(gclk));
	jdff dff_A_wOFbS5LS0_0(.dout(w_dff_A_9te5rlwh6_0),.din(w_dff_A_wOFbS5LS0_0),.clk(gclk));
	jdff dff_A_EBLLEKGN7_0(.dout(w_dff_A_wOFbS5LS0_0),.din(w_dff_A_EBLLEKGN7_0),.clk(gclk));
	jdff dff_A_T1FhP12T4_0(.dout(w_dff_A_EBLLEKGN7_0),.din(w_dff_A_T1FhP12T4_0),.clk(gclk));
	jdff dff_A_rBfVoVXJ8_0(.dout(w_dff_A_T1FhP12T4_0),.din(w_dff_A_rBfVoVXJ8_0),.clk(gclk));
	jdff dff_A_QcH6RXIT7_0(.dout(w_dff_A_rBfVoVXJ8_0),.din(w_dff_A_QcH6RXIT7_0),.clk(gclk));
	jdff dff_A_h3i2shtr9_0(.dout(w_dff_A_QcH6RXIT7_0),.din(w_dff_A_h3i2shtr9_0),.clk(gclk));
	jdff dff_A_BvmYfvAB1_0(.dout(w_dff_A_h3i2shtr9_0),.din(w_dff_A_BvmYfvAB1_0),.clk(gclk));
	jdff dff_A_VJ2PfoYk9_0(.dout(w_dff_A_BvmYfvAB1_0),.din(w_dff_A_VJ2PfoYk9_0),.clk(gclk));
	jdff dff_B_WyeZXHbr1_1(.din(n482),.dout(w_dff_B_WyeZXHbr1_1),.clk(gclk));
	jdff dff_B_4X3kPJrL4_1(.din(w_dff_B_WyeZXHbr1_1),.dout(w_dff_B_4X3kPJrL4_1),.clk(gclk));
	jdff dff_B_g08RlGq63_1(.din(w_dff_B_4X3kPJrL4_1),.dout(w_dff_B_g08RlGq63_1),.clk(gclk));
	jdff dff_A_jMcenfR22_0(.dout(w_n495_1[0]),.din(w_dff_A_jMcenfR22_0),.clk(gclk));
	jdff dff_A_fbyIUOcx5_0(.dout(w_dff_A_jMcenfR22_0),.din(w_dff_A_fbyIUOcx5_0),.clk(gclk));
	jdff dff_A_4cOLjCDA2_0(.dout(w_dff_A_fbyIUOcx5_0),.din(w_dff_A_4cOLjCDA2_0),.clk(gclk));
	jdff dff_A_CNbKM23z5_0(.dout(w_dff_A_4cOLjCDA2_0),.din(w_dff_A_CNbKM23z5_0),.clk(gclk));
	jdff dff_A_vrYdFfq63_0(.dout(w_dff_A_CNbKM23z5_0),.din(w_dff_A_vrYdFfq63_0),.clk(gclk));
	jdff dff_A_AhgtTm8d6_0(.dout(w_dff_A_vrYdFfq63_0),.din(w_dff_A_AhgtTm8d6_0),.clk(gclk));
	jdff dff_A_Vm7Bi5zH8_0(.dout(w_dff_A_AhgtTm8d6_0),.din(w_dff_A_Vm7Bi5zH8_0),.clk(gclk));
	jdff dff_A_HxeLPVrN7_0(.dout(w_dff_A_Vm7Bi5zH8_0),.din(w_dff_A_HxeLPVrN7_0),.clk(gclk));
	jdff dff_A_v4MGICBa5_0(.dout(w_dff_A_HxeLPVrN7_0),.din(w_dff_A_v4MGICBa5_0),.clk(gclk));
	jdff dff_A_1thZgHSK8_0(.dout(w_dff_A_v4MGICBa5_0),.din(w_dff_A_1thZgHSK8_0),.clk(gclk));
	jdff dff_A_sX3ENFkg6_0(.dout(w_dff_A_1thZgHSK8_0),.din(w_dff_A_sX3ENFkg6_0),.clk(gclk));
	jdff dff_A_s6oeVN8V5_0(.dout(w_dff_A_sX3ENFkg6_0),.din(w_dff_A_s6oeVN8V5_0),.clk(gclk));
	jdff dff_A_6jXzVsJW9_0(.dout(w_dff_A_s6oeVN8V5_0),.din(w_dff_A_6jXzVsJW9_0),.clk(gclk));
	jdff dff_A_bktw3wX13_0(.dout(w_dff_A_6jXzVsJW9_0),.din(w_dff_A_bktw3wX13_0),.clk(gclk));
	jdff dff_A_gb6Wb1IB8_0(.dout(w_dff_A_bktw3wX13_0),.din(w_dff_A_gb6Wb1IB8_0),.clk(gclk));
	jdff dff_A_zp2ffKLE6_0(.dout(w_dff_A_gb6Wb1IB8_0),.din(w_dff_A_zp2ffKLE6_0),.clk(gclk));
	jdff dff_A_bXSlSjE39_0(.dout(w_dff_A_zp2ffKLE6_0),.din(w_dff_A_bXSlSjE39_0),.clk(gclk));
	jdff dff_A_hLKCT2WW2_0(.dout(w_dff_A_bXSlSjE39_0),.din(w_dff_A_hLKCT2WW2_0),.clk(gclk));
	jdff dff_A_i8ufmyLE3_0(.dout(w_dff_A_hLKCT2WW2_0),.din(w_dff_A_i8ufmyLE3_0),.clk(gclk));
	jdff dff_B_JtsGdVzx3_1(.din(n484),.dout(w_dff_B_JtsGdVzx3_1),.clk(gclk));
	jdff dff_B_2dzCEDNR0_1(.din(w_dff_B_JtsGdVzx3_1),.dout(w_dff_B_2dzCEDNR0_1),.clk(gclk));
	jdff dff_A_deUKMUkG8_0(.dout(w_n491_1[0]),.din(w_dff_A_deUKMUkG8_0),.clk(gclk));
	jdff dff_A_morsh9Fq2_0(.dout(w_dff_A_deUKMUkG8_0),.din(w_dff_A_morsh9Fq2_0),.clk(gclk));
	jdff dff_A_LLfcPI5v9_0(.dout(w_dff_A_morsh9Fq2_0),.din(w_dff_A_LLfcPI5v9_0),.clk(gclk));
	jdff dff_A_wG0ZifpE8_2(.dout(w_n491_0[2]),.din(w_dff_A_wG0ZifpE8_2),.clk(gclk));
	jdff dff_A_VKErXlhW5_2(.dout(w_dff_A_wG0ZifpE8_2),.din(w_dff_A_VKErXlhW5_2),.clk(gclk));
	jdff dff_A_Td4dErbD5_1(.dout(w_n487_0[1]),.din(w_dff_A_Td4dErbD5_1),.clk(gclk));
	jdff dff_A_RJv3wE9p0_1(.dout(w_dff_A_Td4dErbD5_1),.din(w_dff_A_RJv3wE9p0_1),.clk(gclk));
	jdff dff_A_sXwtEneV7_1(.dout(w_dff_A_RJv3wE9p0_1),.din(w_dff_A_sXwtEneV7_1),.clk(gclk));
	jdff dff_A_LqLvx6vs9_1(.dout(w_dff_A_sXwtEneV7_1),.din(w_dff_A_LqLvx6vs9_1),.clk(gclk));
	jdff dff_A_Y9Y3BmyK7_1(.dout(w_dff_A_LqLvx6vs9_1),.din(w_dff_A_Y9Y3BmyK7_1),.clk(gclk));
	jdff dff_A_euV10qq49_1(.dout(w_dff_A_Y9Y3BmyK7_1),.din(w_dff_A_euV10qq49_1),.clk(gclk));
	jdff dff_A_zxgVdpJs7_1(.dout(w_dff_A_euV10qq49_1),.din(w_dff_A_zxgVdpJs7_1),.clk(gclk));
	jdff dff_A_fA7HAnm02_1(.dout(w_dff_A_zxgVdpJs7_1),.din(w_dff_A_fA7HAnm02_1),.clk(gclk));
	jdff dff_A_VfDpkJqr1_1(.dout(w_dff_A_fA7HAnm02_1),.din(w_dff_A_VfDpkJqr1_1),.clk(gclk));
	jdff dff_A_nlt2YmsH7_1(.dout(w_dff_A_VfDpkJqr1_1),.din(w_dff_A_nlt2YmsH7_1),.clk(gclk));
	jdff dff_A_DPtj4cdg5_1(.dout(w_dff_A_nlt2YmsH7_1),.din(w_dff_A_DPtj4cdg5_1),.clk(gclk));
	jdff dff_A_af5DXFEl3_1(.dout(w_dff_A_DPtj4cdg5_1),.din(w_dff_A_af5DXFEl3_1),.clk(gclk));
	jdff dff_A_6giP8EKq3_1(.dout(w_dff_A_af5DXFEl3_1),.din(w_dff_A_6giP8EKq3_1),.clk(gclk));
	jdff dff_A_Dw9AWMnf6_1(.dout(w_dff_A_6giP8EKq3_1),.din(w_dff_A_Dw9AWMnf6_1),.clk(gclk));
	jdff dff_A_F0DtYoY39_1(.dout(w_dff_A_Dw9AWMnf6_1),.din(w_dff_A_F0DtYoY39_1),.clk(gclk));
	jdff dff_A_ctsS75dJ9_1(.dout(w_dff_A_F0DtYoY39_1),.din(w_dff_A_ctsS75dJ9_1),.clk(gclk));
	jdff dff_A_dtPwwUCt7_1(.dout(w_dff_A_ctsS75dJ9_1),.din(w_dff_A_dtPwwUCt7_1),.clk(gclk));
	jdff dff_A_H8CTkzRh7_1(.dout(w_dff_A_dtPwwUCt7_1),.din(w_dff_A_H8CTkzRh7_1),.clk(gclk));
	jdff dff_A_HOC6O1zJ7_1(.dout(w_dff_A_H8CTkzRh7_1),.din(w_dff_A_HOC6O1zJ7_1),.clk(gclk));
	jdff dff_A_CVe3MJHb0_1(.dout(w_dff_A_HOC6O1zJ7_1),.din(w_dff_A_CVe3MJHb0_1),.clk(gclk));
	jdff dff_A_uttDgsHk0_1(.dout(w_dff_A_CVe3MJHb0_1),.din(w_dff_A_uttDgsHk0_1),.clk(gclk));
	jdff dff_A_ywD6YQRO6_1(.dout(w_dff_A_uttDgsHk0_1),.din(w_dff_A_ywD6YQRO6_1),.clk(gclk));
	jdff dff_A_l3fDYImI1_1(.dout(w_dff_A_ywD6YQRO6_1),.din(w_dff_A_l3fDYImI1_1),.clk(gclk));
	jdff dff_A_AdtOCzBY1_1(.dout(w_dff_A_l3fDYImI1_1),.din(w_dff_A_AdtOCzBY1_1),.clk(gclk));
	jdff dff_A_ixqYGm1o7_0(.dout(w_n481_0[0]),.din(w_dff_A_ixqYGm1o7_0),.clk(gclk));
	jdff dff_A_Wv6rvCIi5_0(.dout(w_dff_A_ixqYGm1o7_0),.din(w_dff_A_Wv6rvCIi5_0),.clk(gclk));
	jdff dff_A_YgJCA40H7_0(.dout(w_dff_A_Wv6rvCIi5_0),.din(w_dff_A_YgJCA40H7_0),.clk(gclk));
	jdff dff_A_FoBgatEC9_0(.dout(w_dff_A_YgJCA40H7_0),.din(w_dff_A_FoBgatEC9_0),.clk(gclk));
	jdff dff_A_SLK28GeL0_0(.dout(w_dff_A_FoBgatEC9_0),.din(w_dff_A_SLK28GeL0_0),.clk(gclk));
	jdff dff_A_fw7sQ5W87_0(.dout(w_dff_A_SLK28GeL0_0),.din(w_dff_A_fw7sQ5W87_0),.clk(gclk));
	jdff dff_A_bjHvmDvY6_0(.dout(w_dff_A_fw7sQ5W87_0),.din(w_dff_A_bjHvmDvY6_0),.clk(gclk));
	jdff dff_A_TqdS7yiw2_0(.dout(w_dff_A_bjHvmDvY6_0),.din(w_dff_A_TqdS7yiw2_0),.clk(gclk));
	jdff dff_A_jeJvfZqg1_0(.dout(w_dff_A_TqdS7yiw2_0),.din(w_dff_A_jeJvfZqg1_0),.clk(gclk));
	jdff dff_A_EJyWmnr29_0(.dout(w_dff_A_jeJvfZqg1_0),.din(w_dff_A_EJyWmnr29_0),.clk(gclk));
	jdff dff_A_ljWnEnYu4_0(.dout(w_dff_A_EJyWmnr29_0),.din(w_dff_A_ljWnEnYu4_0),.clk(gclk));
	jdff dff_A_LxUaOaY84_0(.dout(w_dff_A_ljWnEnYu4_0),.din(w_dff_A_LxUaOaY84_0),.clk(gclk));
	jdff dff_A_OJIukkaT8_0(.dout(w_dff_A_LxUaOaY84_0),.din(w_dff_A_OJIukkaT8_0),.clk(gclk));
	jdff dff_A_cq1EfrJU1_0(.dout(w_dff_A_OJIukkaT8_0),.din(w_dff_A_cq1EfrJU1_0),.clk(gclk));
	jdff dff_A_Jsq2I9WM1_0(.dout(w_dff_A_cq1EfrJU1_0),.din(w_dff_A_Jsq2I9WM1_0),.clk(gclk));
	jdff dff_A_dqOX5aeL9_0(.dout(w_dff_A_Jsq2I9WM1_0),.din(w_dff_A_dqOX5aeL9_0),.clk(gclk));
	jdff dff_A_jgP0GqKZ1_0(.dout(w_dff_A_dqOX5aeL9_0),.din(w_dff_A_jgP0GqKZ1_0),.clk(gclk));
	jdff dff_A_vVf75h6x2_0(.dout(w_dff_A_jgP0GqKZ1_0),.din(w_dff_A_vVf75h6x2_0),.clk(gclk));
	jdff dff_A_nB36qrht8_0(.dout(w_dff_A_vVf75h6x2_0),.din(w_dff_A_nB36qrht8_0),.clk(gclk));
	jdff dff_A_wDM6Fowa2_0(.dout(w_dff_A_nB36qrht8_0),.din(w_dff_A_wDM6Fowa2_0),.clk(gclk));
	jdff dff_A_zEyFOwDZ0_0(.dout(w_dff_A_wDM6Fowa2_0),.din(w_dff_A_zEyFOwDZ0_0),.clk(gclk));
	jdff dff_A_PjQxVjRq2_0(.dout(w_dff_A_zEyFOwDZ0_0),.din(w_dff_A_PjQxVjRq2_0),.clk(gclk));
	jdff dff_A_7dEHGSlS3_2(.dout(w_n480_0[2]),.din(w_dff_A_7dEHGSlS3_2),.clk(gclk));
	jdff dff_A_Unfq8XEe0_2(.dout(w_dff_A_7dEHGSlS3_2),.din(w_dff_A_Unfq8XEe0_2),.clk(gclk));
	jdff dff_A_XBArIg9C2_2(.dout(w_dff_A_Unfq8XEe0_2),.din(w_dff_A_XBArIg9C2_2),.clk(gclk));
	jdff dff_A_93PiUjLl4_2(.dout(w_dff_A_XBArIg9C2_2),.din(w_dff_A_93PiUjLl4_2),.clk(gclk));
	jdff dff_A_5f2KQPVj1_2(.dout(w_dff_A_93PiUjLl4_2),.din(w_dff_A_5f2KQPVj1_2),.clk(gclk));
	jdff dff_A_dqu1Ec3R5_2(.dout(w_dff_A_5f2KQPVj1_2),.din(w_dff_A_dqu1Ec3R5_2),.clk(gclk));
	jdff dff_A_dxGJRV5L1_2(.dout(w_dff_A_dqu1Ec3R5_2),.din(w_dff_A_dxGJRV5L1_2),.clk(gclk));
	jdff dff_A_kMabNZBW6_2(.dout(w_dff_A_dxGJRV5L1_2),.din(w_dff_A_kMabNZBW6_2),.clk(gclk));
	jdff dff_A_du08SVZh0_2(.dout(w_dff_A_kMabNZBW6_2),.din(w_dff_A_du08SVZh0_2),.clk(gclk));
	jdff dff_A_9PwJ1itP8_2(.dout(w_dff_A_du08SVZh0_2),.din(w_dff_A_9PwJ1itP8_2),.clk(gclk));
	jdff dff_A_s2YSep9r3_2(.dout(w_dff_A_9PwJ1itP8_2),.din(w_dff_A_s2YSep9r3_2),.clk(gclk));
	jdff dff_A_4mgP7Jwu0_2(.dout(w_dff_A_s2YSep9r3_2),.din(w_dff_A_4mgP7Jwu0_2),.clk(gclk));
	jdff dff_A_V2A7bli74_2(.dout(w_dff_A_4mgP7Jwu0_2),.din(w_dff_A_V2A7bli74_2),.clk(gclk));
	jdff dff_A_eZTe3fYw8_2(.dout(w_dff_A_V2A7bli74_2),.din(w_dff_A_eZTe3fYw8_2),.clk(gclk));
	jdff dff_A_IkjMENBR8_2(.dout(w_dff_A_eZTe3fYw8_2),.din(w_dff_A_IkjMENBR8_2),.clk(gclk));
	jdff dff_A_pe96QAlF8_2(.dout(w_dff_A_IkjMENBR8_2),.din(w_dff_A_pe96QAlF8_2),.clk(gclk));
	jdff dff_A_c4aHzUs29_2(.dout(w_dff_A_pe96QAlF8_2),.din(w_dff_A_c4aHzUs29_2),.clk(gclk));
	jdff dff_A_z62fQYdD3_2(.dout(w_dff_A_c4aHzUs29_2),.din(w_dff_A_z62fQYdD3_2),.clk(gclk));
	jdff dff_A_4SEeGFhv8_2(.dout(w_dff_A_z62fQYdD3_2),.din(w_dff_A_4SEeGFhv8_2),.clk(gclk));
	jdff dff_A_KOHVLl2s2_2(.dout(w_dff_A_4SEeGFhv8_2),.din(w_dff_A_KOHVLl2s2_2),.clk(gclk));
	jdff dff_A_UYgUFvLc4_2(.dout(w_dff_A_KOHVLl2s2_2),.din(w_dff_A_UYgUFvLc4_2),.clk(gclk));
	jdff dff_A_W2yMJyFv7_2(.dout(w_dff_A_UYgUFvLc4_2),.din(w_dff_A_W2yMJyFv7_2),.clk(gclk));
	jdff dff_A_qzEOAB5K5_2(.dout(w_dff_A_W2yMJyFv7_2),.din(w_dff_A_qzEOAB5K5_2),.clk(gclk));
	jdff dff_B_YBVMhFrw4_0(.din(n478),.dout(w_dff_B_YBVMhFrw4_0),.clk(gclk));
	jdff dff_B_sPQTSDO91_0(.din(G147),.dout(w_dff_B_sPQTSDO91_0),.clk(gclk));
	jdff dff_A_rbide4Po5_1(.dout(w_n476_0[1]),.din(w_dff_A_rbide4Po5_1),.clk(gclk));
	jdff dff_A_nz0WVmC46_1(.dout(w_dff_A_rbide4Po5_1),.din(w_dff_A_nz0WVmC46_1),.clk(gclk));
	jdff dff_A_pR8aIAKi6_2(.dout(w_n476_0[2]),.din(w_dff_A_pR8aIAKi6_2),.clk(gclk));
	jdff dff_A_1SPzV9KS9_2(.dout(w_dff_A_pR8aIAKi6_2),.din(w_dff_A_1SPzV9KS9_2),.clk(gclk));
	jdff dff_A_sGQoS01B7_1(.dout(w_G2211_0[1]),.din(w_dff_A_sGQoS01B7_1),.clk(gclk));
	jdff dff_A_qrDWNDAB0_1(.dout(w_dff_A_sGQoS01B7_1),.din(w_dff_A_qrDWNDAB0_1),.clk(gclk));
	jdff dff_A_MnOJFYCr0_1(.dout(w_dff_A_qrDWNDAB0_1),.din(w_dff_A_MnOJFYCr0_1),.clk(gclk));
	jdff dff_A_4jd6T85v2_1(.dout(w_dff_A_MnOJFYCr0_1),.din(w_dff_A_4jd6T85v2_1),.clk(gclk));
	jdff dff_A_6rNoCX3n4_1(.dout(w_n475_0[1]),.din(w_dff_A_6rNoCX3n4_1),.clk(gclk));
	jdff dff_A_NotIBoFg4_1(.dout(w_dff_A_6rNoCX3n4_1),.din(w_dff_A_NotIBoFg4_1),.clk(gclk));
	jdff dff_A_CblEHEA98_1(.dout(w_dff_A_NotIBoFg4_1),.din(w_dff_A_CblEHEA98_1),.clk(gclk));
	jdff dff_A_o9EmDkHT5_1(.dout(w_dff_A_CblEHEA98_1),.din(w_dff_A_o9EmDkHT5_1),.clk(gclk));
	jdff dff_A_c25rgt6U1_1(.dout(w_dff_A_o9EmDkHT5_1),.din(w_dff_A_c25rgt6U1_1),.clk(gclk));
	jdff dff_A_iP8JrcrQ8_1(.dout(w_dff_A_c25rgt6U1_1),.din(w_dff_A_iP8JrcrQ8_1),.clk(gclk));
	jdff dff_A_5uCsJvHT3_1(.dout(w_dff_A_iP8JrcrQ8_1),.din(w_dff_A_5uCsJvHT3_1),.clk(gclk));
	jdff dff_A_Ar5yrfF34_1(.dout(w_dff_A_5uCsJvHT3_1),.din(w_dff_A_Ar5yrfF34_1),.clk(gclk));
	jdff dff_A_8K2was2a9_1(.dout(w_dff_A_Ar5yrfF34_1),.din(w_dff_A_8K2was2a9_1),.clk(gclk));
	jdff dff_A_KE3zLGnF9_1(.dout(w_dff_A_8K2was2a9_1),.din(w_dff_A_KE3zLGnF9_1),.clk(gclk));
	jdff dff_A_60TIwxxS2_1(.dout(w_dff_A_KE3zLGnF9_1),.din(w_dff_A_60TIwxxS2_1),.clk(gclk));
	jdff dff_A_8QjpGOze1_1(.dout(w_dff_A_60TIwxxS2_1),.din(w_dff_A_8QjpGOze1_1),.clk(gclk));
	jdff dff_A_3ICgD0yx3_1(.dout(w_dff_A_8QjpGOze1_1),.din(w_dff_A_3ICgD0yx3_1),.clk(gclk));
	jdff dff_A_zQHypauh2_1(.dout(w_dff_A_3ICgD0yx3_1),.din(w_dff_A_zQHypauh2_1),.clk(gclk));
	jdff dff_A_Y2HCjpeZ3_1(.dout(w_dff_A_zQHypauh2_1),.din(w_dff_A_Y2HCjpeZ3_1),.clk(gclk));
	jdff dff_A_QrAtwv8C7_1(.dout(w_dff_A_Y2HCjpeZ3_1),.din(w_dff_A_QrAtwv8C7_1),.clk(gclk));
	jdff dff_A_Pf1AyaWd1_1(.dout(w_dff_A_QrAtwv8C7_1),.din(w_dff_A_Pf1AyaWd1_1),.clk(gclk));
	jdff dff_A_WN2omO4Y4_1(.dout(w_dff_A_Pf1AyaWd1_1),.din(w_dff_A_WN2omO4Y4_1),.clk(gclk));
	jdff dff_A_BKSl8FZe3_1(.dout(w_dff_A_WN2omO4Y4_1),.din(w_dff_A_BKSl8FZe3_1),.clk(gclk));
	jdff dff_A_NgHy1mTr1_1(.dout(w_dff_A_BKSl8FZe3_1),.din(w_dff_A_NgHy1mTr1_1),.clk(gclk));
	jdff dff_A_pqVDuJwH0_1(.dout(w_dff_A_NgHy1mTr1_1),.din(w_dff_A_pqVDuJwH0_1),.clk(gclk));
	jdff dff_A_ioEIHelg3_1(.dout(w_dff_A_pqVDuJwH0_1),.din(w_dff_A_ioEIHelg3_1),.clk(gclk));
	jdff dff_A_CheGRkuj5_1(.dout(w_dff_A_ioEIHelg3_1),.din(w_dff_A_CheGRkuj5_1),.clk(gclk));
	jdff dff_A_p3LiCpr75_1(.dout(w_dff_A_CheGRkuj5_1),.din(w_dff_A_p3LiCpr75_1),.clk(gclk));
	jdff dff_A_iNqFcuDB5_1(.dout(w_dff_A_p3LiCpr75_1),.din(w_dff_A_iNqFcuDB5_1),.clk(gclk));
	jdff dff_B_ahLzISW37_0(.din(n473),.dout(w_dff_B_ahLzISW37_0),.clk(gclk));
	jdff dff_B_F3PASO123_0(.din(G138),.dout(w_dff_B_F3PASO123_0),.clk(gclk));
	jdff dff_A_sqRzoyHI0_1(.dout(w_n471_0[1]),.din(w_dff_A_sqRzoyHI0_1),.clk(gclk));
	jdff dff_A_AEUcQ3Nn0_1(.dout(w_dff_A_sqRzoyHI0_1),.din(w_dff_A_AEUcQ3Nn0_1),.clk(gclk));
	jdff dff_A_tCymbE621_2(.dout(w_n471_0[2]),.din(w_dff_A_tCymbE621_2),.clk(gclk));
	jdff dff_A_CoRA3fFb5_2(.dout(w_dff_A_tCymbE621_2),.din(w_dff_A_CoRA3fFb5_2),.clk(gclk));
	jdff dff_A_tavuTiH99_1(.dout(w_G2218_0[1]),.din(w_dff_A_tavuTiH99_1),.clk(gclk));
	jdff dff_A_WktiMIxJ5_1(.dout(w_dff_A_tavuTiH99_1),.din(w_dff_A_WktiMIxJ5_1),.clk(gclk));
	jdff dff_A_DQVx4nYE2_1(.dout(w_dff_A_WktiMIxJ5_1),.din(w_dff_A_DQVx4nYE2_1),.clk(gclk));
	jdff dff_A_ejDtG6IA4_1(.dout(w_dff_A_DQVx4nYE2_1),.din(w_dff_A_ejDtG6IA4_1),.clk(gclk));
	jdff dff_A_PZWFXNLs9_1(.dout(w_n470_0[1]),.din(w_dff_A_PZWFXNLs9_1),.clk(gclk));
	jdff dff_A_R86NxYsJ6_1(.dout(w_dff_A_PZWFXNLs9_1),.din(w_dff_A_R86NxYsJ6_1),.clk(gclk));
	jdff dff_A_C5vvK6m33_1(.dout(w_dff_A_R86NxYsJ6_1),.din(w_dff_A_C5vvK6m33_1),.clk(gclk));
	jdff dff_A_kOnaPuB27_1(.dout(w_dff_A_C5vvK6m33_1),.din(w_dff_A_kOnaPuB27_1),.clk(gclk));
	jdff dff_A_3sMKEa3p7_1(.dout(w_dff_A_kOnaPuB27_1),.din(w_dff_A_3sMKEa3p7_1),.clk(gclk));
	jdff dff_A_JhgKSz0k8_1(.dout(w_dff_A_3sMKEa3p7_1),.din(w_dff_A_JhgKSz0k8_1),.clk(gclk));
	jdff dff_A_nvpwnhzr6_1(.dout(w_dff_A_JhgKSz0k8_1),.din(w_dff_A_nvpwnhzr6_1),.clk(gclk));
	jdff dff_A_XTQAwFBM3_1(.dout(w_dff_A_nvpwnhzr6_1),.din(w_dff_A_XTQAwFBM3_1),.clk(gclk));
	jdff dff_A_043I4qEv6_1(.dout(w_dff_A_XTQAwFBM3_1),.din(w_dff_A_043I4qEv6_1),.clk(gclk));
	jdff dff_A_1tZbmfKg6_1(.dout(w_dff_A_043I4qEv6_1),.din(w_dff_A_1tZbmfKg6_1),.clk(gclk));
	jdff dff_A_YjaYXnGM2_1(.dout(w_dff_A_1tZbmfKg6_1),.din(w_dff_A_YjaYXnGM2_1),.clk(gclk));
	jdff dff_A_52dVQub69_1(.dout(w_dff_A_YjaYXnGM2_1),.din(w_dff_A_52dVQub69_1),.clk(gclk));
	jdff dff_A_JNAGShZX7_1(.dout(w_dff_A_52dVQub69_1),.din(w_dff_A_JNAGShZX7_1),.clk(gclk));
	jdff dff_A_hLm5jJZp3_1(.dout(w_dff_A_JNAGShZX7_1),.din(w_dff_A_hLm5jJZp3_1),.clk(gclk));
	jdff dff_A_lNNwIN8B6_1(.dout(w_dff_A_hLm5jJZp3_1),.din(w_dff_A_lNNwIN8B6_1),.clk(gclk));
	jdff dff_A_OewrYHc16_1(.dout(w_dff_A_lNNwIN8B6_1),.din(w_dff_A_OewrYHc16_1),.clk(gclk));
	jdff dff_A_v2heRr9F6_1(.dout(w_dff_A_OewrYHc16_1),.din(w_dff_A_v2heRr9F6_1),.clk(gclk));
	jdff dff_A_dWEs66E19_1(.dout(w_dff_A_v2heRr9F6_1),.din(w_dff_A_dWEs66E19_1),.clk(gclk));
	jdff dff_A_BhADi4hU3_1(.dout(w_dff_A_dWEs66E19_1),.din(w_dff_A_BhADi4hU3_1),.clk(gclk));
	jdff dff_A_all0LASw7_1(.dout(w_dff_A_BhADi4hU3_1),.din(w_dff_A_all0LASw7_1),.clk(gclk));
	jdff dff_A_ZOi4iXss8_1(.dout(w_dff_A_all0LASw7_1),.din(w_dff_A_ZOi4iXss8_1),.clk(gclk));
	jdff dff_A_D2x2x57p3_1(.dout(w_dff_A_ZOi4iXss8_1),.din(w_dff_A_D2x2x57p3_1),.clk(gclk));
	jdff dff_A_VuCtGG891_1(.dout(w_dff_A_D2x2x57p3_1),.din(w_dff_A_VuCtGG891_1),.clk(gclk));
	jdff dff_A_nDvXNVFL7_1(.dout(w_dff_A_VuCtGG891_1),.din(w_dff_A_nDvXNVFL7_1),.clk(gclk));
	jdff dff_A_T7jq9jDO9_1(.dout(w_dff_A_nDvXNVFL7_1),.din(w_dff_A_T7jq9jDO9_1),.clk(gclk));
	jdff dff_A_bhpvO7y81_2(.dout(w_n470_0[2]),.din(w_dff_A_bhpvO7y81_2),.clk(gclk));
	jdff dff_A_2iW2PPZY8_1(.dout(w_n469_0[1]),.din(w_dff_A_2iW2PPZY8_1),.clk(gclk));
	jdff dff_B_KFM86BYY5_0(.din(n468),.dout(w_dff_B_KFM86BYY5_0),.clk(gclk));
	jdff dff_B_L0FO5yLy8_0(.din(G144),.dout(w_dff_B_L0FO5yLy8_0),.clk(gclk));
	jdff dff_B_7VdUCKjH3_2(.din(n466),.dout(w_dff_B_7VdUCKjH3_2),.clk(gclk));
	jdff dff_B_faLwkV1V1_2(.din(w_dff_B_7VdUCKjH3_2),.dout(w_dff_B_faLwkV1V1_2),.clk(gclk));
	jdff dff_A_caASnzbL5_0(.dout(w_G2224_1[0]),.din(w_dff_A_caASnzbL5_0),.clk(gclk));
	jdff dff_A_VoAJ2kes2_0(.dout(w_dff_A_caASnzbL5_0),.din(w_dff_A_VoAJ2kes2_0),.clk(gclk));
	jdff dff_A_v13rWSEn4_0(.dout(w_dff_A_VoAJ2kes2_0),.din(w_dff_A_v13rWSEn4_0),.clk(gclk));
	jdff dff_A_l1y0aVPn7_0(.dout(w_dff_A_v13rWSEn4_0),.din(w_dff_A_l1y0aVPn7_0),.clk(gclk));
	jdff dff_A_AEtra7w43_1(.dout(w_n465_0[1]),.din(w_dff_A_AEtra7w43_1),.clk(gclk));
	jdff dff_B_l2wkP1F76_2(.din(n465),.dout(w_dff_B_l2wkP1F76_2),.clk(gclk));
	jdff dff_B_4kkUNG699_2(.din(w_dff_B_l2wkP1F76_2),.dout(w_dff_B_4kkUNG699_2),.clk(gclk));
	jdff dff_B_Q6mApC7R4_2(.din(w_dff_B_4kkUNG699_2),.dout(w_dff_B_Q6mApC7R4_2),.clk(gclk));
	jdff dff_B_8NkWGC5a1_2(.din(w_dff_B_Q6mApC7R4_2),.dout(w_dff_B_8NkWGC5a1_2),.clk(gclk));
	jdff dff_A_pOGrQRJ74_1(.dout(w_n464_0[1]),.din(w_dff_A_pOGrQRJ74_1),.clk(gclk));
	jdff dff_A_4cFrbtet4_1(.dout(w_dff_A_pOGrQRJ74_1),.din(w_dff_A_4cFrbtet4_1),.clk(gclk));
	jdff dff_A_ttM2uUXo0_1(.dout(w_dff_A_4cFrbtet4_1),.din(w_dff_A_ttM2uUXo0_1),.clk(gclk));
	jdff dff_A_G6gEQHXt7_1(.dout(w_dff_A_ttM2uUXo0_1),.din(w_dff_A_G6gEQHXt7_1),.clk(gclk));
	jdff dff_A_TvL30THj2_1(.dout(w_dff_A_G6gEQHXt7_1),.din(w_dff_A_TvL30THj2_1),.clk(gclk));
	jdff dff_A_5cxykv8L1_1(.dout(w_dff_A_TvL30THj2_1),.din(w_dff_A_5cxykv8L1_1),.clk(gclk));
	jdff dff_A_zCXWJnRx8_1(.dout(w_dff_A_5cxykv8L1_1),.din(w_dff_A_zCXWJnRx8_1),.clk(gclk));
	jdff dff_A_13AGVodk3_1(.dout(w_dff_A_zCXWJnRx8_1),.din(w_dff_A_13AGVodk3_1),.clk(gclk));
	jdff dff_A_X2WrYvLe1_1(.dout(w_dff_A_13AGVodk3_1),.din(w_dff_A_X2WrYvLe1_1),.clk(gclk));
	jdff dff_A_oMdgqgGd7_1(.dout(w_dff_A_X2WrYvLe1_1),.din(w_dff_A_oMdgqgGd7_1),.clk(gclk));
	jdff dff_A_2OckOhek1_1(.dout(w_dff_A_oMdgqgGd7_1),.din(w_dff_A_2OckOhek1_1),.clk(gclk));
	jdff dff_A_o4723JXm7_1(.dout(w_dff_A_2OckOhek1_1),.din(w_dff_A_o4723JXm7_1),.clk(gclk));
	jdff dff_A_GpWcJurk9_1(.dout(w_dff_A_o4723JXm7_1),.din(w_dff_A_GpWcJurk9_1),.clk(gclk));
	jdff dff_A_qY5T57XT4_1(.dout(w_dff_A_GpWcJurk9_1),.din(w_dff_A_qY5T57XT4_1),.clk(gclk));
	jdff dff_A_k2u2chqi7_1(.dout(w_dff_A_qY5T57XT4_1),.din(w_dff_A_k2u2chqi7_1),.clk(gclk));
	jdff dff_A_GTWvrOJQ6_1(.dout(w_dff_A_k2u2chqi7_1),.din(w_dff_A_GTWvrOJQ6_1),.clk(gclk));
	jdff dff_A_TF61Uxpp9_1(.dout(w_dff_A_GTWvrOJQ6_1),.din(w_dff_A_TF61Uxpp9_1),.clk(gclk));
	jdff dff_A_41JQzHdh9_1(.dout(w_dff_A_TF61Uxpp9_1),.din(w_dff_A_41JQzHdh9_1),.clk(gclk));
	jdff dff_A_pDyqnRQE7_1(.dout(w_dff_A_41JQzHdh9_1),.din(w_dff_A_pDyqnRQE7_1),.clk(gclk));
	jdff dff_A_lhbev20A3_1(.dout(w_dff_A_pDyqnRQE7_1),.din(w_dff_A_lhbev20A3_1),.clk(gclk));
	jdff dff_A_4O90wrX25_1(.dout(w_dff_A_lhbev20A3_1),.din(w_dff_A_4O90wrX25_1),.clk(gclk));
	jdff dff_A_yQmnoKOA2_1(.dout(w_dff_A_4O90wrX25_1),.din(w_dff_A_yQmnoKOA2_1),.clk(gclk));
	jdff dff_A_r1MOO3YE6_1(.dout(w_dff_A_yQmnoKOA2_1),.din(w_dff_A_r1MOO3YE6_1),.clk(gclk));
	jdff dff_A_wJUIGS9O9_1(.dout(w_dff_A_r1MOO3YE6_1),.din(w_dff_A_wJUIGS9O9_1),.clk(gclk));
	jdff dff_A_LN73Blkg7_1(.dout(w_dff_A_wJUIGS9O9_1),.din(w_dff_A_LN73Blkg7_1),.clk(gclk));
	jdff dff_A_k81yAa526_1(.dout(w_dff_A_LN73Blkg7_1),.din(w_dff_A_k81yAa526_1),.clk(gclk));
	jdff dff_A_UaCQODc75_0(.dout(w_n463_1[0]),.din(w_dff_A_UaCQODc75_0),.clk(gclk));
	jdff dff_A_UjtKMMZn4_0(.dout(w_dff_A_UaCQODc75_0),.din(w_dff_A_UjtKMMZn4_0),.clk(gclk));
	jdff dff_A_ptbWX0HT0_0(.dout(w_dff_A_UjtKMMZn4_0),.din(w_dff_A_ptbWX0HT0_0),.clk(gclk));
	jdff dff_A_K3ootG9A8_0(.dout(w_dff_A_ptbWX0HT0_0),.din(w_dff_A_K3ootG9A8_0),.clk(gclk));
	jdff dff_A_UpRHNI212_0(.dout(w_dff_A_K3ootG9A8_0),.din(w_dff_A_UpRHNI212_0),.clk(gclk));
	jdff dff_A_Go9qbMMu2_0(.dout(w_dff_A_UpRHNI212_0),.din(w_dff_A_Go9qbMMu2_0),.clk(gclk));
	jdff dff_A_yC46ZHJd7_0(.dout(w_dff_A_Go9qbMMu2_0),.din(w_dff_A_yC46ZHJd7_0),.clk(gclk));
	jdff dff_A_8k6Kz5o43_0(.dout(w_dff_A_yC46ZHJd7_0),.din(w_dff_A_8k6Kz5o43_0),.clk(gclk));
	jdff dff_A_2qiBYBpj5_0(.dout(w_dff_A_8k6Kz5o43_0),.din(w_dff_A_2qiBYBpj5_0),.clk(gclk));
	jdff dff_A_WPKsUuVp2_0(.dout(w_dff_A_2qiBYBpj5_0),.din(w_dff_A_WPKsUuVp2_0),.clk(gclk));
	jdff dff_A_s4JpMiZd2_0(.dout(w_dff_A_WPKsUuVp2_0),.din(w_dff_A_s4JpMiZd2_0),.clk(gclk));
	jdff dff_A_WQ8eqC0R4_0(.dout(w_dff_A_s4JpMiZd2_0),.din(w_dff_A_WQ8eqC0R4_0),.clk(gclk));
	jdff dff_A_jQedEa9h7_0(.dout(w_dff_A_WQ8eqC0R4_0),.din(w_dff_A_jQedEa9h7_0),.clk(gclk));
	jdff dff_A_mimc7q7d7_0(.dout(w_dff_A_jQedEa9h7_0),.din(w_dff_A_mimc7q7d7_0),.clk(gclk));
	jdff dff_A_meMNJLVk2_0(.dout(w_dff_A_mimc7q7d7_0),.din(w_dff_A_meMNJLVk2_0),.clk(gclk));
	jdff dff_A_5flPCkGW2_0(.dout(w_dff_A_meMNJLVk2_0),.din(w_dff_A_5flPCkGW2_0),.clk(gclk));
	jdff dff_A_whrHmqgw8_0(.dout(w_dff_A_5flPCkGW2_0),.din(w_dff_A_whrHmqgw8_0),.clk(gclk));
	jdff dff_A_5S1UkWTf8_0(.dout(w_dff_A_whrHmqgw8_0),.din(w_dff_A_5S1UkWTf8_0),.clk(gclk));
	jdff dff_A_SHWbbS468_0(.dout(w_dff_A_5S1UkWTf8_0),.din(w_dff_A_SHWbbS468_0),.clk(gclk));
	jdff dff_A_rEpJmsOW1_0(.dout(w_dff_A_SHWbbS468_0),.din(w_dff_A_rEpJmsOW1_0),.clk(gclk));
	jdff dff_A_Oaej3STT6_0(.dout(w_dff_A_rEpJmsOW1_0),.din(w_dff_A_Oaej3STT6_0),.clk(gclk));
	jdff dff_A_dNXNp3CK8_0(.dout(w_dff_A_Oaej3STT6_0),.din(w_dff_A_dNXNp3CK8_0),.clk(gclk));
	jdff dff_A_J2DPbQwi1_0(.dout(w_dff_A_dNXNp3CK8_0),.din(w_dff_A_J2DPbQwi1_0),.clk(gclk));
	jdff dff_A_pcoKWbB46_0(.dout(w_dff_A_J2DPbQwi1_0),.din(w_dff_A_pcoKWbB46_0),.clk(gclk));
	jdff dff_A_gldFSnIi1_0(.dout(w_dff_A_pcoKWbB46_0),.din(w_dff_A_gldFSnIi1_0),.clk(gclk));
	jdff dff_A_j2LrPGVh2_0(.dout(w_dff_A_gldFSnIi1_0),.din(w_dff_A_j2LrPGVh2_0),.clk(gclk));
	jdff dff_A_bYv9v9ah0_0(.dout(w_dff_A_j2LrPGVh2_0),.din(w_dff_A_bYv9v9ah0_0),.clk(gclk));
	jdff dff_A_mm9xl4ny1_0(.dout(w_dff_A_bYv9v9ah0_0),.din(w_dff_A_mm9xl4ny1_0),.clk(gclk));
	jdff dff_A_G1k9tSbX4_1(.dout(w_n463_0[1]),.din(w_dff_A_G1k9tSbX4_1),.clk(gclk));
	jdff dff_A_3dcrqoOw5_1(.dout(w_dff_A_G1k9tSbX4_1),.din(w_dff_A_3dcrqoOw5_1),.clk(gclk));
	jdff dff_A_OOnyHpnr0_1(.dout(w_dff_A_3dcrqoOw5_1),.din(w_dff_A_OOnyHpnr0_1),.clk(gclk));
	jdff dff_A_HOEtFrdf6_2(.dout(w_n463_0[2]),.din(w_dff_A_HOEtFrdf6_2),.clk(gclk));
	jdff dff_A_mggUfphE7_2(.dout(w_dff_A_HOEtFrdf6_2),.din(w_dff_A_mggUfphE7_2),.clk(gclk));
	jdff dff_A_GiEsqJZu5_2(.dout(w_dff_A_mggUfphE7_2),.din(w_dff_A_GiEsqJZu5_2),.clk(gclk));
	jdff dff_A_23iTfWE05_2(.dout(w_dff_A_GiEsqJZu5_2),.din(w_dff_A_23iTfWE05_2),.clk(gclk));
	jdff dff_A_Rf91Ri1L3_1(.dout(w_n462_0[1]),.din(w_dff_A_Rf91Ri1L3_1),.clk(gclk));
	jdff dff_A_hpJFL3sK0_1(.dout(w_dff_A_Rf91Ri1L3_1),.din(w_dff_A_hpJFL3sK0_1),.clk(gclk));
	jdff dff_A_Z26zVEXv0_1(.dout(w_dff_A_hpJFL3sK0_1),.din(w_dff_A_Z26zVEXv0_1),.clk(gclk));
	jdff dff_A_vjieTZMz6_1(.dout(w_dff_A_Z26zVEXv0_1),.din(w_dff_A_vjieTZMz6_1),.clk(gclk));
	jdff dff_A_cdWFS5cL6_1(.dout(w_dff_A_vjieTZMz6_1),.din(w_dff_A_cdWFS5cL6_1),.clk(gclk));
	jdff dff_A_ky4Amsyu1_1(.dout(w_dff_A_cdWFS5cL6_1),.din(w_dff_A_ky4Amsyu1_1),.clk(gclk));
	jdff dff_A_hgSBaEk42_1(.dout(w_dff_A_ky4Amsyu1_1),.din(w_dff_A_hgSBaEk42_1),.clk(gclk));
	jdff dff_A_OlHMVJ4s3_1(.dout(w_dff_A_hgSBaEk42_1),.din(w_dff_A_OlHMVJ4s3_1),.clk(gclk));
	jdff dff_A_t7KsHmnV8_1(.dout(w_dff_A_OlHMVJ4s3_1),.din(w_dff_A_t7KsHmnV8_1),.clk(gclk));
	jdff dff_A_pN6C2wDF7_1(.dout(w_dff_A_t7KsHmnV8_1),.din(w_dff_A_pN6C2wDF7_1),.clk(gclk));
	jdff dff_A_SDN5vM8n2_1(.dout(w_dff_A_pN6C2wDF7_1),.din(w_dff_A_SDN5vM8n2_1),.clk(gclk));
	jdff dff_A_nfEqkOvf0_1(.dout(w_dff_A_SDN5vM8n2_1),.din(w_dff_A_nfEqkOvf0_1),.clk(gclk));
	jdff dff_A_uyfU2R556_1(.dout(w_dff_A_nfEqkOvf0_1),.din(w_dff_A_uyfU2R556_1),.clk(gclk));
	jdff dff_A_P376HyIw7_1(.dout(w_dff_A_uyfU2R556_1),.din(w_dff_A_P376HyIw7_1),.clk(gclk));
	jdff dff_A_NFZRabpp8_1(.dout(w_dff_A_P376HyIw7_1),.din(w_dff_A_NFZRabpp8_1),.clk(gclk));
	jdff dff_A_X7Ynu4Cz3_1(.dout(w_dff_A_NFZRabpp8_1),.din(w_dff_A_X7Ynu4Cz3_1),.clk(gclk));
	jdff dff_A_QipKPhqW4_1(.dout(w_dff_A_X7Ynu4Cz3_1),.din(w_dff_A_QipKPhqW4_1),.clk(gclk));
	jdff dff_A_NcPLJRFM8_1(.dout(w_dff_A_QipKPhqW4_1),.din(w_dff_A_NcPLJRFM8_1),.clk(gclk));
	jdff dff_A_vJhYnvck0_1(.dout(w_dff_A_NcPLJRFM8_1),.din(w_dff_A_vJhYnvck0_1),.clk(gclk));
	jdff dff_A_qc4czDye1_1(.dout(w_dff_A_vJhYnvck0_1),.din(w_dff_A_qc4czDye1_1),.clk(gclk));
	jdff dff_A_KeAGqp0V3_1(.dout(w_dff_A_qc4czDye1_1),.din(w_dff_A_KeAGqp0V3_1),.clk(gclk));
	jdff dff_A_L9VoewlE4_2(.dout(w_n462_0[2]),.din(w_dff_A_L9VoewlE4_2),.clk(gclk));
	jdff dff_A_qzCVUCyk7_2(.dout(w_dff_A_L9VoewlE4_2),.din(w_dff_A_qzCVUCyk7_2),.clk(gclk));
	jdff dff_A_bPgGgxjM5_2(.dout(w_dff_A_qzCVUCyk7_2),.din(w_dff_A_bPgGgxjM5_2),.clk(gclk));
	jdff dff_A_gKC5si9E3_2(.dout(w_dff_A_bPgGgxjM5_2),.din(w_dff_A_gKC5si9E3_2),.clk(gclk));
	jdff dff_A_9UTW68s00_2(.dout(w_dff_A_gKC5si9E3_2),.din(w_dff_A_9UTW68s00_2),.clk(gclk));
	jdff dff_B_awopLnNH5_1(.din(n454),.dout(w_dff_B_awopLnNH5_1),.clk(gclk));
	jdff dff_A_k54MonoF7_0(.dout(w_n460_1[0]),.din(w_dff_A_k54MonoF7_0),.clk(gclk));
	jdff dff_A_XFZsADoa1_0(.dout(w_dff_A_k54MonoF7_0),.din(w_dff_A_XFZsADoa1_0),.clk(gclk));
	jdff dff_A_6Fzfy2Kw6_0(.dout(w_dff_A_XFZsADoa1_0),.din(w_dff_A_6Fzfy2Kw6_0),.clk(gclk));
	jdff dff_A_WOMwj1407_0(.dout(w_dff_A_6Fzfy2Kw6_0),.din(w_dff_A_WOMwj1407_0),.clk(gclk));
	jdff dff_A_lTbCl6VD0_0(.dout(w_dff_A_WOMwj1407_0),.din(w_dff_A_lTbCl6VD0_0),.clk(gclk));
	jdff dff_A_Jaufee2s4_0(.dout(w_dff_A_lTbCl6VD0_0),.din(w_dff_A_Jaufee2s4_0),.clk(gclk));
	jdff dff_A_3K3HuQsC1_0(.dout(w_dff_A_Jaufee2s4_0),.din(w_dff_A_3K3HuQsC1_0),.clk(gclk));
	jdff dff_A_I8bYwQpi8_0(.dout(w_dff_A_3K3HuQsC1_0),.din(w_dff_A_I8bYwQpi8_0),.clk(gclk));
	jdff dff_A_tr4JXemg5_0(.dout(w_dff_A_I8bYwQpi8_0),.din(w_dff_A_tr4JXemg5_0),.clk(gclk));
	jdff dff_A_uVdBUZgR5_0(.dout(w_dff_A_tr4JXemg5_0),.din(w_dff_A_uVdBUZgR5_0),.clk(gclk));
	jdff dff_A_lJRI20IG7_0(.dout(w_dff_A_uVdBUZgR5_0),.din(w_dff_A_lJRI20IG7_0),.clk(gclk));
	jdff dff_A_OggVfmVL6_0(.dout(w_dff_A_lJRI20IG7_0),.din(w_dff_A_OggVfmVL6_0),.clk(gclk));
	jdff dff_A_fbyLv0JS6_0(.dout(w_dff_A_OggVfmVL6_0),.din(w_dff_A_fbyLv0JS6_0),.clk(gclk));
	jdff dff_A_JLadxANj4_0(.dout(w_dff_A_fbyLv0JS6_0),.din(w_dff_A_JLadxANj4_0),.clk(gclk));
	jdff dff_A_TaoVFQzy5_0(.dout(w_dff_A_JLadxANj4_0),.din(w_dff_A_TaoVFQzy5_0),.clk(gclk));
	jdff dff_A_CUw2PL7y8_0(.dout(w_dff_A_TaoVFQzy5_0),.din(w_dff_A_CUw2PL7y8_0),.clk(gclk));
	jdff dff_A_3Ykac4vI4_0(.dout(w_dff_A_CUw2PL7y8_0),.din(w_dff_A_3Ykac4vI4_0),.clk(gclk));
	jdff dff_A_2HLiQELv2_0(.dout(w_dff_A_3Ykac4vI4_0),.din(w_dff_A_2HLiQELv2_0),.clk(gclk));
	jdff dff_A_gEPW8tZJ0_0(.dout(w_dff_A_2HLiQELv2_0),.din(w_dff_A_gEPW8tZJ0_0),.clk(gclk));
	jdff dff_A_tPxeaxz58_0(.dout(w_dff_A_gEPW8tZJ0_0),.din(w_dff_A_tPxeaxz58_0),.clk(gclk));
	jdff dff_A_XZ6FJpzZ7_0(.dout(w_dff_A_tPxeaxz58_0),.din(w_dff_A_XZ6FJpzZ7_0),.clk(gclk));
	jdff dff_A_mXitxHfX8_0(.dout(w_dff_A_XZ6FJpzZ7_0),.din(w_dff_A_mXitxHfX8_0),.clk(gclk));
	jdff dff_A_MM3YtLNQ1_0(.dout(w_dff_A_mXitxHfX8_0),.din(w_dff_A_MM3YtLNQ1_0),.clk(gclk));
	jdff dff_A_D83NkRkf2_0(.dout(w_dff_A_MM3YtLNQ1_0),.din(w_dff_A_D83NkRkf2_0),.clk(gclk));
	jdff dff_A_Prlrm1Jf5_0(.dout(w_dff_A_D83NkRkf2_0),.din(w_dff_A_Prlrm1Jf5_0),.clk(gclk));
	jdff dff_A_zpjBqJBo4_0(.dout(w_dff_A_Prlrm1Jf5_0),.din(w_dff_A_zpjBqJBo4_0),.clk(gclk));
	jdff dff_A_PAbldBJs3_0(.dout(w_dff_A_zpjBqJBo4_0),.din(w_dff_A_PAbldBJs3_0),.clk(gclk));
	jdff dff_A_mzPJmmpA5_0(.dout(w_dff_A_PAbldBJs3_0),.din(w_dff_A_mzPJmmpA5_0),.clk(gclk));
	jdff dff_A_D6r6m7ZR6_1(.dout(w_n460_1[1]),.din(w_dff_A_D6r6m7ZR6_1),.clk(gclk));
	jdff dff_A_Cd2kLbxp1_1(.dout(w_dff_A_D6r6m7ZR6_1),.din(w_dff_A_Cd2kLbxp1_1),.clk(gclk));
	jdff dff_A_i6aS6Uzj7_1(.dout(w_dff_A_Cd2kLbxp1_1),.din(w_dff_A_i6aS6Uzj7_1),.clk(gclk));
	jdff dff_A_HZaM7yQs6_1(.dout(w_dff_A_i6aS6Uzj7_1),.din(w_dff_A_HZaM7yQs6_1),.clk(gclk));
	jdff dff_A_p4hK0S748_1(.dout(w_dff_A_HZaM7yQs6_1),.din(w_dff_A_p4hK0S748_1),.clk(gclk));
	jdff dff_A_cs9eMcnY5_1(.dout(w_dff_A_p4hK0S748_1),.din(w_dff_A_cs9eMcnY5_1),.clk(gclk));
	jdff dff_A_OVY1ZdqL7_1(.dout(w_dff_A_cs9eMcnY5_1),.din(w_dff_A_OVY1ZdqL7_1),.clk(gclk));
	jdff dff_A_QI2cO9NY5_1(.dout(w_dff_A_OVY1ZdqL7_1),.din(w_dff_A_QI2cO9NY5_1),.clk(gclk));
	jdff dff_A_q5JZpPPZ4_1(.dout(w_dff_A_QI2cO9NY5_1),.din(w_dff_A_q5JZpPPZ4_1),.clk(gclk));
	jdff dff_A_9ojgAUoF7_1(.dout(w_dff_A_q5JZpPPZ4_1),.din(w_dff_A_9ojgAUoF7_1),.clk(gclk));
	jdff dff_A_uNPmcJ450_1(.dout(w_dff_A_9ojgAUoF7_1),.din(w_dff_A_uNPmcJ450_1),.clk(gclk));
	jdff dff_A_Gu8katj50_1(.dout(w_dff_A_uNPmcJ450_1),.din(w_dff_A_Gu8katj50_1),.clk(gclk));
	jdff dff_A_BFuNihQf4_1(.dout(w_dff_A_Gu8katj50_1),.din(w_dff_A_BFuNihQf4_1),.clk(gclk));
	jdff dff_A_0jMCvRlY8_1(.dout(w_dff_A_BFuNihQf4_1),.din(w_dff_A_0jMCvRlY8_1),.clk(gclk));
	jdff dff_A_y8KDwPwL0_1(.dout(w_dff_A_0jMCvRlY8_1),.din(w_dff_A_y8KDwPwL0_1),.clk(gclk));
	jdff dff_A_gD5kEaY65_1(.dout(w_dff_A_y8KDwPwL0_1),.din(w_dff_A_gD5kEaY65_1),.clk(gclk));
	jdff dff_A_gLfuqoBq6_1(.dout(w_dff_A_gD5kEaY65_1),.din(w_dff_A_gLfuqoBq6_1),.clk(gclk));
	jdff dff_A_BKMi7xRg3_1(.dout(w_dff_A_gLfuqoBq6_1),.din(w_dff_A_BKMi7xRg3_1),.clk(gclk));
	jdff dff_A_9CRIjJAW2_1(.dout(w_dff_A_BKMi7xRg3_1),.din(w_dff_A_9CRIjJAW2_1),.clk(gclk));
	jdff dff_A_l1Pl7gFq8_1(.dout(w_dff_A_9CRIjJAW2_1),.din(w_dff_A_l1Pl7gFq8_1),.clk(gclk));
	jdff dff_A_R2MjCZWp0_1(.dout(w_dff_A_l1Pl7gFq8_1),.din(w_dff_A_R2MjCZWp0_1),.clk(gclk));
	jdff dff_A_rlbrlT4k6_1(.dout(w_dff_A_R2MjCZWp0_1),.din(w_dff_A_rlbrlT4k6_1),.clk(gclk));
	jdff dff_A_ATBdNKld5_1(.dout(w_dff_A_rlbrlT4k6_1),.din(w_dff_A_ATBdNKld5_1),.clk(gclk));
	jdff dff_A_boWxus9s7_1(.dout(w_dff_A_ATBdNKld5_1),.din(w_dff_A_boWxus9s7_1),.clk(gclk));
	jdff dff_A_1m3cni3m7_1(.dout(w_dff_A_boWxus9s7_1),.din(w_dff_A_1m3cni3m7_1),.clk(gclk));
	jdff dff_A_g6KYlXOQ2_1(.dout(w_dff_A_1m3cni3m7_1),.din(w_dff_A_g6KYlXOQ2_1),.clk(gclk));
	jdff dff_A_N4yhrShC2_1(.dout(w_dff_A_g6KYlXOQ2_1),.din(w_dff_A_N4yhrShC2_1),.clk(gclk));
	jdff dff_A_g1jzQxd28_1(.dout(w_n460_0[1]),.din(w_dff_A_g1jzQxd28_1),.clk(gclk));
	jdff dff_A_rYATWfRs2_1(.dout(w_dff_A_g1jzQxd28_1),.din(w_dff_A_rYATWfRs2_1),.clk(gclk));
	jdff dff_A_6p8k5DXg7_1(.dout(w_dff_A_rYATWfRs2_1),.din(w_dff_A_6p8k5DXg7_1),.clk(gclk));
	jdff dff_A_VTlxaBkL6_1(.dout(w_dff_A_6p8k5DXg7_1),.din(w_dff_A_VTlxaBkL6_1),.clk(gclk));
	jdff dff_A_fIiVjdhg4_1(.dout(w_dff_A_VTlxaBkL6_1),.din(w_dff_A_fIiVjdhg4_1),.clk(gclk));
	jdff dff_A_oMDMfYxR4_1(.dout(w_dff_A_fIiVjdhg4_1),.din(w_dff_A_oMDMfYxR4_1),.clk(gclk));
	jdff dff_A_wc1m5kDg1_2(.dout(w_n460_0[2]),.din(w_dff_A_wc1m5kDg1_2),.clk(gclk));
	jdff dff_A_NoJhKZFu6_2(.dout(w_dff_A_wc1m5kDg1_2),.din(w_dff_A_NoJhKZFu6_2),.clk(gclk));
	jdff dff_A_lJjdzwwr6_2(.dout(w_dff_A_NoJhKZFu6_2),.din(w_dff_A_lJjdzwwr6_2),.clk(gclk));
	jdff dff_A_nXayk9as8_2(.dout(w_dff_A_lJjdzwwr6_2),.din(w_dff_A_nXayk9as8_2),.clk(gclk));
	jdff dff_A_JsuecAtg8_2(.dout(w_dff_A_nXayk9as8_2),.din(w_dff_A_JsuecAtg8_2),.clk(gclk));
	jdff dff_A_OJNo70x40_2(.dout(w_dff_A_JsuecAtg8_2),.din(w_dff_A_OJNo70x40_2),.clk(gclk));
	jdff dff_A_qlnCXpzK1_2(.dout(w_dff_A_OJNo70x40_2),.din(w_dff_A_qlnCXpzK1_2),.clk(gclk));
	jdff dff_B_OMw2dKd80_0(.din(n458),.dout(w_dff_B_OMw2dKd80_0),.clk(gclk));
	jdff dff_B_ysREwqJz0_0(.din(G135),.dout(w_dff_B_ysREwqJz0_0),.clk(gclk));
	jdff dff_A_MTwDKs0H0_1(.dout(w_n456_0[1]),.din(w_dff_A_MTwDKs0H0_1),.clk(gclk));
	jdff dff_A_GH49b0Su4_1(.dout(w_dff_A_MTwDKs0H0_1),.din(w_dff_A_GH49b0Su4_1),.clk(gclk));
	jdff dff_A_wc2lkZX18_2(.dout(w_n456_0[2]),.din(w_dff_A_wc2lkZX18_2),.clk(gclk));
	jdff dff_A_ma0gtraA9_2(.dout(w_dff_A_wc2lkZX18_2),.din(w_dff_A_ma0gtraA9_2),.clk(gclk));
	jdff dff_A_R1Gxr56t4_1(.dout(w_G2230_0[1]),.din(w_dff_A_R1Gxr56t4_1),.clk(gclk));
	jdff dff_A_MfAaBqbI0_1(.dout(w_dff_A_R1Gxr56t4_1),.din(w_dff_A_MfAaBqbI0_1),.clk(gclk));
	jdff dff_A_G8sCmpI01_1(.dout(w_dff_A_MfAaBqbI0_1),.din(w_dff_A_G8sCmpI01_1),.clk(gclk));
	jdff dff_A_Goj5lNI45_1(.dout(w_dff_A_G8sCmpI01_1),.din(w_dff_A_Goj5lNI45_1),.clk(gclk));
	jdff dff_A_awJpdhdt3_1(.dout(w_n453_0[1]),.din(w_dff_A_awJpdhdt3_1),.clk(gclk));
	jdff dff_B_EvTmIQ8u7_0(.din(G157),.dout(w_dff_B_EvTmIQ8u7_0),.clk(gclk));
	jdff dff_B_MgTpLvgR6_3(.din(n451),.dout(w_dff_B_MgTpLvgR6_3),.clk(gclk));
	jdff dff_B_bNAyFE7f2_3(.din(w_dff_B_MgTpLvgR6_3),.dout(w_dff_B_bNAyFE7f2_3),.clk(gclk));
	jdff dff_A_3S1neNv82_2(.dout(w_n450_0[2]),.din(w_dff_A_3S1neNv82_2),.clk(gclk));
	jdff dff_A_ykxDAA0P3_2(.dout(w_dff_A_3S1neNv82_2),.din(w_dff_A_ykxDAA0P3_2),.clk(gclk));
	jdff dff_A_tFbW4tOx3_2(.dout(w_dff_A_ykxDAA0P3_2),.din(w_dff_A_tFbW4tOx3_2),.clk(gclk));
	jdff dff_A_tvye38Pp7_2(.dout(w_dff_A_tFbW4tOx3_2),.din(w_dff_A_tvye38Pp7_2),.clk(gclk));
	jdff dff_A_enhqDaiv4_2(.dout(w_dff_A_tvye38Pp7_2),.din(w_dff_A_enhqDaiv4_2),.clk(gclk));
	jdff dff_A_eItKloPp7_2(.dout(w_dff_A_enhqDaiv4_2),.din(w_dff_A_eItKloPp7_2),.clk(gclk));
	jdff dff_A_0d6vNpb52_2(.dout(w_dff_A_eItKloPp7_2),.din(w_dff_A_0d6vNpb52_2),.clk(gclk));
	jdff dff_A_yf62CRGq7_2(.dout(w_dff_A_0d6vNpb52_2),.din(w_dff_A_yf62CRGq7_2),.clk(gclk));
	jdff dff_A_LsuuyCNT7_2(.dout(w_dff_A_yf62CRGq7_2),.din(w_dff_A_LsuuyCNT7_2),.clk(gclk));
	jdff dff_A_KA1S5kW75_2(.dout(w_dff_A_LsuuyCNT7_2),.din(w_dff_A_KA1S5kW75_2),.clk(gclk));
	jdff dff_A_mMLIqVbr8_2(.dout(w_dff_A_KA1S5kW75_2),.din(w_dff_A_mMLIqVbr8_2),.clk(gclk));
	jdff dff_A_qRfaVIaL4_2(.dout(w_dff_A_mMLIqVbr8_2),.din(w_dff_A_qRfaVIaL4_2),.clk(gclk));
	jdff dff_A_KYEyjIBc4_2(.dout(w_dff_A_qRfaVIaL4_2),.din(w_dff_A_KYEyjIBc4_2),.clk(gclk));
	jdff dff_A_jtDziYMX8_2(.dout(w_dff_A_KYEyjIBc4_2),.din(w_dff_A_jtDziYMX8_2),.clk(gclk));
	jdff dff_A_JwZ5fufX0_2(.dout(w_dff_A_jtDziYMX8_2),.din(w_dff_A_JwZ5fufX0_2),.clk(gclk));
	jdff dff_A_JO1coacm2_2(.dout(w_dff_A_JwZ5fufX0_2),.din(w_dff_A_JO1coacm2_2),.clk(gclk));
	jdff dff_A_Y0CwjJpz5_2(.dout(w_dff_A_JO1coacm2_2),.din(w_dff_A_Y0CwjJpz5_2),.clk(gclk));
	jdff dff_A_nM01yALH0_2(.dout(w_dff_A_Y0CwjJpz5_2),.din(w_dff_A_nM01yALH0_2),.clk(gclk));
	jdff dff_A_h2uaSdnx1_2(.dout(w_dff_A_nM01yALH0_2),.din(w_dff_A_h2uaSdnx1_2),.clk(gclk));
	jdff dff_A_DKY0ehu74_2(.dout(w_dff_A_h2uaSdnx1_2),.din(w_dff_A_DKY0ehu74_2),.clk(gclk));
	jdff dff_A_5knmi0wC6_2(.dout(w_dff_A_DKY0ehu74_2),.din(w_dff_A_5knmi0wC6_2),.clk(gclk));
	jdff dff_A_DNUoJNJS9_2(.dout(w_dff_A_5knmi0wC6_2),.din(w_dff_A_DNUoJNJS9_2),.clk(gclk));
	jdff dff_B_OMd4cECq2_1(.din(n439),.dout(w_dff_B_OMd4cECq2_1),.clk(gclk));
	jdff dff_B_jcpkSiok6_1(.din(w_dff_B_OMd4cECq2_1),.dout(w_dff_B_jcpkSiok6_1),.clk(gclk));
	jdff dff_A_Do1sJfAz5_0(.dout(w_n449_1[0]),.din(w_dff_A_Do1sJfAz5_0),.clk(gclk));
	jdff dff_A_NouzY9c38_0(.dout(w_dff_A_Do1sJfAz5_0),.din(w_dff_A_NouzY9c38_0),.clk(gclk));
	jdff dff_A_2CwuWeYS2_0(.dout(w_dff_A_NouzY9c38_0),.din(w_dff_A_2CwuWeYS2_0),.clk(gclk));
	jdff dff_A_rczZvGLY6_0(.dout(w_dff_A_2CwuWeYS2_0),.din(w_dff_A_rczZvGLY6_0),.clk(gclk));
	jdff dff_A_3czVK9Hi5_0(.dout(w_dff_A_rczZvGLY6_0),.din(w_dff_A_3czVK9Hi5_0),.clk(gclk));
	jdff dff_A_UPXzAwwS1_0(.dout(w_dff_A_3czVK9Hi5_0),.din(w_dff_A_UPXzAwwS1_0),.clk(gclk));
	jdff dff_A_Z7s8AnT55_0(.dout(w_dff_A_UPXzAwwS1_0),.din(w_dff_A_Z7s8AnT55_0),.clk(gclk));
	jdff dff_A_OCEYguF52_0(.dout(w_dff_A_Z7s8AnT55_0),.din(w_dff_A_OCEYguF52_0),.clk(gclk));
	jdff dff_A_cyVtxLIv9_0(.dout(w_dff_A_OCEYguF52_0),.din(w_dff_A_cyVtxLIv9_0),.clk(gclk));
	jdff dff_A_D8iRD0d30_0(.dout(w_dff_A_cyVtxLIv9_0),.din(w_dff_A_D8iRD0d30_0),.clk(gclk));
	jdff dff_A_c88lOILW2_0(.dout(w_dff_A_D8iRD0d30_0),.din(w_dff_A_c88lOILW2_0),.clk(gclk));
	jdff dff_A_rC09rrzG1_0(.dout(w_dff_A_c88lOILW2_0),.din(w_dff_A_rC09rrzG1_0),.clk(gclk));
	jdff dff_A_T9WLxHLB0_0(.dout(w_dff_A_rC09rrzG1_0),.din(w_dff_A_T9WLxHLB0_0),.clk(gclk));
	jdff dff_A_4rOCjNwl0_0(.dout(w_dff_A_T9WLxHLB0_0),.din(w_dff_A_4rOCjNwl0_0),.clk(gclk));
	jdff dff_A_oPhxW1jV8_0(.dout(w_dff_A_4rOCjNwl0_0),.din(w_dff_A_oPhxW1jV8_0),.clk(gclk));
	jdff dff_A_bPiOyOgD4_0(.dout(w_dff_A_oPhxW1jV8_0),.din(w_dff_A_bPiOyOgD4_0),.clk(gclk));
	jdff dff_A_Wv6O4urJ2_0(.dout(w_dff_A_bPiOyOgD4_0),.din(w_dff_A_Wv6O4urJ2_0),.clk(gclk));
	jdff dff_A_S34mABln7_0(.dout(w_dff_A_Wv6O4urJ2_0),.din(w_dff_A_S34mABln7_0),.clk(gclk));
	jdff dff_A_4gEplQKp0_0(.dout(w_dff_A_S34mABln7_0),.din(w_dff_A_4gEplQKp0_0),.clk(gclk));
	jdff dff_A_B17cHXGn9_0(.dout(w_dff_A_4gEplQKp0_0),.din(w_dff_A_B17cHXGn9_0),.clk(gclk));
	jdff dff_A_zcWYUNbH5_0(.dout(w_dff_A_B17cHXGn9_0),.din(w_dff_A_zcWYUNbH5_0),.clk(gclk));
	jdff dff_A_DJvvuMLZ3_0(.dout(w_dff_A_zcWYUNbH5_0),.din(w_dff_A_DJvvuMLZ3_0),.clk(gclk));
	jdff dff_B_92yrD0BR6_1(.din(n442),.dout(w_dff_B_92yrD0BR6_1),.clk(gclk));
	jdff dff_B_p7xMscoi9_1(.din(n443),.dout(w_dff_B_p7xMscoi9_1),.clk(gclk));
	jdff dff_B_Ou96JSKD7_1(.din(w_dff_B_p7xMscoi9_1),.dout(w_dff_B_Ou96JSKD7_1),.clk(gclk));
	jdff dff_A_lSOvDucG9_1(.dout(w_n447_0[1]),.din(w_dff_A_lSOvDucG9_1),.clk(gclk));
	jdff dff_A_0og9mOzJ2_1(.dout(w_dff_A_lSOvDucG9_1),.din(w_dff_A_0og9mOzJ2_1),.clk(gclk));
	jdff dff_A_g8jwiIRc6_1(.dout(w_dff_A_0og9mOzJ2_1),.din(w_dff_A_g8jwiIRc6_1),.clk(gclk));
	jdff dff_A_562oG0IR3_1(.dout(w_dff_A_g8jwiIRc6_1),.din(w_dff_A_562oG0IR3_1),.clk(gclk));
	jdff dff_A_ooJOZcO43_1(.dout(w_dff_A_562oG0IR3_1),.din(w_dff_A_ooJOZcO43_1),.clk(gclk));
	jdff dff_A_bQ5XIrnC0_1(.dout(w_dff_A_ooJOZcO43_1),.din(w_dff_A_bQ5XIrnC0_1),.clk(gclk));
	jdff dff_A_y6vuZmFO8_1(.dout(w_dff_A_bQ5XIrnC0_1),.din(w_dff_A_y6vuZmFO8_1),.clk(gclk));
	jdff dff_A_77w7c0Vu9_1(.dout(w_dff_A_y6vuZmFO8_1),.din(w_dff_A_77w7c0Vu9_1),.clk(gclk));
	jdff dff_A_jT8ITcZl9_1(.dout(w_dff_A_77w7c0Vu9_1),.din(w_dff_A_jT8ITcZl9_1),.clk(gclk));
	jdff dff_A_u9H8DKzF4_1(.dout(w_dff_A_jT8ITcZl9_1),.din(w_dff_A_u9H8DKzF4_1),.clk(gclk));
	jdff dff_A_XUMC7h4P2_1(.dout(w_dff_A_u9H8DKzF4_1),.din(w_dff_A_XUMC7h4P2_1),.clk(gclk));
	jdff dff_A_MxfbuE8l9_1(.dout(w_dff_A_XUMC7h4P2_1),.din(w_dff_A_MxfbuE8l9_1),.clk(gclk));
	jdff dff_A_R0ntPxkG1_1(.dout(w_dff_A_MxfbuE8l9_1),.din(w_dff_A_R0ntPxkG1_1),.clk(gclk));
	jdff dff_A_D3ZAsYJc5_1(.dout(w_dff_A_R0ntPxkG1_1),.din(w_dff_A_D3ZAsYJc5_1),.clk(gclk));
	jdff dff_A_1HMHWy0a3_1(.dout(w_dff_A_D3ZAsYJc5_1),.din(w_dff_A_1HMHWy0a3_1),.clk(gclk));
	jdff dff_A_ql5cb95U8_1(.dout(w_dff_A_1HMHWy0a3_1),.din(w_dff_A_ql5cb95U8_1),.clk(gclk));
	jdff dff_A_llMvCMUc7_1(.dout(w_dff_A_ql5cb95U8_1),.din(w_dff_A_llMvCMUc7_1),.clk(gclk));
	jdff dff_A_7myUnSTh2_1(.dout(w_dff_A_llMvCMUc7_1),.din(w_dff_A_7myUnSTh2_1),.clk(gclk));
	jdff dff_A_zp1yClKZ0_1(.dout(w_dff_A_7myUnSTh2_1),.din(w_dff_A_zp1yClKZ0_1),.clk(gclk));
	jdff dff_A_3JW7lJiX4_1(.dout(w_dff_A_zp1yClKZ0_1),.din(w_dff_A_3JW7lJiX4_1),.clk(gclk));
	jdff dff_A_yZhDyhzO9_1(.dout(w_dff_A_3JW7lJiX4_1),.din(w_dff_A_yZhDyhzO9_1),.clk(gclk));
	jdff dff_A_moLcn9wU0_1(.dout(w_dff_A_yZhDyhzO9_1),.din(w_dff_A_moLcn9wU0_1),.clk(gclk));
	jdff dff_A_56ri7JEp4_1(.dout(w_dff_A_moLcn9wU0_1),.din(w_dff_A_56ri7JEp4_1),.clk(gclk));
	jdff dff_A_GpfJrIyz1_1(.dout(w_dff_A_56ri7JEp4_1),.din(w_dff_A_GpfJrIyz1_1),.clk(gclk));
	jdff dff_A_RFn9ktMs9_1(.dout(w_dff_A_GpfJrIyz1_1),.din(w_dff_A_RFn9ktMs9_1),.clk(gclk));
	jdff dff_A_VUVo3DE22_1(.dout(w_n445_0[1]),.din(w_dff_A_VUVo3DE22_1),.clk(gclk));
	jdff dff_A_5PZGs2378_1(.dout(w_dff_A_VUVo3DE22_1),.din(w_dff_A_5PZGs2378_1),.clk(gclk));
	jdff dff_A_WsaBE3856_1(.dout(w_dff_A_5PZGs2378_1),.din(w_dff_A_WsaBE3856_1),.clk(gclk));
	jdff dff_A_TkcaGzHM1_1(.dout(w_dff_A_WsaBE3856_1),.din(w_dff_A_TkcaGzHM1_1),.clk(gclk));
	jdff dff_A_j2HZZJ2b8_1(.dout(w_dff_A_TkcaGzHM1_1),.din(w_dff_A_j2HZZJ2b8_1),.clk(gclk));
	jdff dff_A_g3jquSgD0_1(.dout(w_dff_A_j2HZZJ2b8_1),.din(w_dff_A_g3jquSgD0_1),.clk(gclk));
	jdff dff_A_OZRE09i87_1(.dout(w_dff_A_g3jquSgD0_1),.din(w_dff_A_OZRE09i87_1),.clk(gclk));
	jdff dff_A_etf9XN9x5_1(.dout(w_dff_A_OZRE09i87_1),.din(w_dff_A_etf9XN9x5_1),.clk(gclk));
	jdff dff_A_0t2k46q24_1(.dout(w_dff_A_etf9XN9x5_1),.din(w_dff_A_0t2k46q24_1),.clk(gclk));
	jdff dff_A_AJeRGgbJ2_1(.dout(w_dff_A_0t2k46q24_1),.din(w_dff_A_AJeRGgbJ2_1),.clk(gclk));
	jdff dff_A_LYO3CrNn0_1(.dout(w_dff_A_AJeRGgbJ2_1),.din(w_dff_A_LYO3CrNn0_1),.clk(gclk));
	jdff dff_A_SruZ1Knl4_1(.dout(w_dff_A_LYO3CrNn0_1),.din(w_dff_A_SruZ1Knl4_1),.clk(gclk));
	jdff dff_A_39mH9nLB8_1(.dout(w_dff_A_SruZ1Knl4_1),.din(w_dff_A_39mH9nLB8_1),.clk(gclk));
	jdff dff_A_dh5nasNr4_1(.dout(w_dff_A_39mH9nLB8_1),.din(w_dff_A_dh5nasNr4_1),.clk(gclk));
	jdff dff_A_7mirB95L5_1(.dout(w_dff_A_dh5nasNr4_1),.din(w_dff_A_7mirB95L5_1),.clk(gclk));
	jdff dff_A_OwyZFgff2_1(.dout(w_dff_A_7mirB95L5_1),.din(w_dff_A_OwyZFgff2_1),.clk(gclk));
	jdff dff_A_2XPP5Prc7_1(.dout(w_dff_A_OwyZFgff2_1),.din(w_dff_A_2XPP5Prc7_1),.clk(gclk));
	jdff dff_A_twyROc2w9_1(.dout(w_dff_A_2XPP5Prc7_1),.din(w_dff_A_twyROc2w9_1),.clk(gclk));
	jdff dff_A_L9IcrBII0_1(.dout(w_dff_A_twyROc2w9_1),.din(w_dff_A_L9IcrBII0_1),.clk(gclk));
	jdff dff_A_Awvm9W7S9_1(.dout(w_dff_A_L9IcrBII0_1),.din(w_dff_A_Awvm9W7S9_1),.clk(gclk));
	jdff dff_A_HhO3Cjdg8_1(.dout(w_dff_A_Awvm9W7S9_1),.din(w_dff_A_HhO3Cjdg8_1),.clk(gclk));
	jdff dff_A_3z9xDdNO9_1(.dout(w_dff_A_HhO3Cjdg8_1),.din(w_dff_A_3z9xDdNO9_1),.clk(gclk));
	jdff dff_A_yFnz547Q7_1(.dout(w_dff_A_3z9xDdNO9_1),.din(w_dff_A_yFnz547Q7_1),.clk(gclk));
	jdff dff_A_6Fi2hSCE6_1(.dout(w_dff_A_yFnz547Q7_1),.din(w_dff_A_6Fi2hSCE6_1),.clk(gclk));
	jdff dff_A_S05y18lQ3_1(.dout(w_dff_A_6Fi2hSCE6_1),.din(w_dff_A_S05y18lQ3_1),.clk(gclk));
	jdff dff_A_OaUA8Du73_1(.dout(w_dff_A_S05y18lQ3_1),.din(w_dff_A_OaUA8Du73_1),.clk(gclk));
	jdff dff_A_uO1vhw4H7_1(.dout(w_n444_0[1]),.din(w_dff_A_uO1vhw4H7_1),.clk(gclk));
	jdff dff_A_a66fwNCD5_1(.dout(w_dff_A_uO1vhw4H7_1),.din(w_dff_A_a66fwNCD5_1),.clk(gclk));
	jdff dff_A_CO40dOUl0_2(.dout(w_n444_0[2]),.din(w_dff_A_CO40dOUl0_2),.clk(gclk));
	jdff dff_A_k6HhHNvI3_0(.dout(w_n438_0[0]),.din(w_dff_A_k6HhHNvI3_0),.clk(gclk));
	jdff dff_A_CH0mOYP28_0(.dout(w_dff_A_k6HhHNvI3_0),.din(w_dff_A_CH0mOYP28_0),.clk(gclk));
	jdff dff_A_IbM43Zvt2_0(.dout(w_dff_A_CH0mOYP28_0),.din(w_dff_A_IbM43Zvt2_0),.clk(gclk));
	jdff dff_A_fLryOFyT8_0(.dout(w_dff_A_IbM43Zvt2_0),.din(w_dff_A_fLryOFyT8_0),.clk(gclk));
	jdff dff_A_RIoNaBDg0_0(.dout(w_dff_A_fLryOFyT8_0),.din(w_dff_A_RIoNaBDg0_0),.clk(gclk));
	jdff dff_A_vvyyG51H5_0(.dout(w_dff_A_RIoNaBDg0_0),.din(w_dff_A_vvyyG51H5_0),.clk(gclk));
	jdff dff_A_Njb6Iykp2_0(.dout(w_dff_A_vvyyG51H5_0),.din(w_dff_A_Njb6Iykp2_0),.clk(gclk));
	jdff dff_A_puOeH4213_0(.dout(w_dff_A_Njb6Iykp2_0),.din(w_dff_A_puOeH4213_0),.clk(gclk));
	jdff dff_A_ZdalX3Tx6_0(.dout(w_dff_A_puOeH4213_0),.din(w_dff_A_ZdalX3Tx6_0),.clk(gclk));
	jdff dff_A_2YY4HiPW9_0(.dout(w_dff_A_ZdalX3Tx6_0),.din(w_dff_A_2YY4HiPW9_0),.clk(gclk));
	jdff dff_A_o2mStPB95_0(.dout(w_dff_A_2YY4HiPW9_0),.din(w_dff_A_o2mStPB95_0),.clk(gclk));
	jdff dff_A_Zj86wMtU0_0(.dout(w_dff_A_o2mStPB95_0),.din(w_dff_A_Zj86wMtU0_0),.clk(gclk));
	jdff dff_A_F6N1Egpz5_0(.dout(w_dff_A_Zj86wMtU0_0),.din(w_dff_A_F6N1Egpz5_0),.clk(gclk));
	jdff dff_A_4stGaW3o8_0(.dout(w_dff_A_F6N1Egpz5_0),.din(w_dff_A_4stGaW3o8_0),.clk(gclk));
	jdff dff_A_JX6KbI918_0(.dout(w_dff_A_4stGaW3o8_0),.din(w_dff_A_JX6KbI918_0),.clk(gclk));
	jdff dff_A_PMK8qwEG7_0(.dout(w_dff_A_JX6KbI918_0),.din(w_dff_A_PMK8qwEG7_0),.clk(gclk));
	jdff dff_A_THvPmz6x0_0(.dout(w_dff_A_PMK8qwEG7_0),.din(w_dff_A_THvPmz6x0_0),.clk(gclk));
	jdff dff_A_vsMZr1rU0_0(.dout(w_dff_A_THvPmz6x0_0),.din(w_dff_A_vsMZr1rU0_0),.clk(gclk));
	jdff dff_A_K85VhOl68_0(.dout(w_dff_A_vsMZr1rU0_0),.din(w_dff_A_K85VhOl68_0),.clk(gclk));
	jdff dff_A_dEaryAQz7_0(.dout(w_dff_A_K85VhOl68_0),.din(w_dff_A_dEaryAQz7_0),.clk(gclk));
	jdff dff_A_pgfyR0812_0(.dout(w_dff_A_dEaryAQz7_0),.din(w_dff_A_pgfyR0812_0),.clk(gclk));
	jdff dff_A_FM1OgzgO3_0(.dout(w_dff_A_pgfyR0812_0),.din(w_dff_A_FM1OgzgO3_0),.clk(gclk));
	jdff dff_A_jWP61y9L6_0(.dout(w_dff_A_FM1OgzgO3_0),.din(w_dff_A_jWP61y9L6_0),.clk(gclk));
	jdff dff_A_rMjcHjkf5_0(.dout(w_dff_A_jWP61y9L6_0),.din(w_dff_A_rMjcHjkf5_0),.clk(gclk));
	jdff dff_A_ZCXL6AFb6_0(.dout(w_dff_A_rMjcHjkf5_0),.din(w_dff_A_ZCXL6AFb6_0),.clk(gclk));
	jdff dff_A_NuFAHOKH5_1(.dout(w_n437_0[1]),.din(w_dff_A_NuFAHOKH5_1),.clk(gclk));
	jdff dff_A_ugyEEQqb4_1(.dout(w_dff_A_NuFAHOKH5_1),.din(w_dff_A_ugyEEQqb4_1),.clk(gclk));
	jdff dff_A_B3uSnQhe1_1(.dout(w_dff_A_ugyEEQqb4_1),.din(w_dff_A_B3uSnQhe1_1),.clk(gclk));
	jdff dff_A_82knghJg4_1(.dout(w_dff_A_B3uSnQhe1_1),.din(w_dff_A_82knghJg4_1),.clk(gclk));
	jdff dff_A_HVGFICnp9_1(.dout(w_dff_A_82knghJg4_1),.din(w_dff_A_HVGFICnp9_1),.clk(gclk));
	jdff dff_A_dueqnUqy6_1(.dout(w_dff_A_HVGFICnp9_1),.din(w_dff_A_dueqnUqy6_1),.clk(gclk));
	jdff dff_A_WAfWcaXV9_1(.dout(w_dff_A_dueqnUqy6_1),.din(w_dff_A_WAfWcaXV9_1),.clk(gclk));
	jdff dff_A_Iv52h5mp0_1(.dout(w_dff_A_WAfWcaXV9_1),.din(w_dff_A_Iv52h5mp0_1),.clk(gclk));
	jdff dff_A_w8Fw9Eu57_1(.dout(w_dff_A_Iv52h5mp0_1),.din(w_dff_A_w8Fw9Eu57_1),.clk(gclk));
	jdff dff_A_Uq9F3kxL2_1(.dout(w_dff_A_w8Fw9Eu57_1),.din(w_dff_A_Uq9F3kxL2_1),.clk(gclk));
	jdff dff_A_OfCpVxKO8_1(.dout(w_dff_A_Uq9F3kxL2_1),.din(w_dff_A_OfCpVxKO8_1),.clk(gclk));
	jdff dff_A_zMsGmvg76_1(.dout(w_dff_A_OfCpVxKO8_1),.din(w_dff_A_zMsGmvg76_1),.clk(gclk));
	jdff dff_A_Iq2PYwmo5_1(.dout(w_dff_A_zMsGmvg76_1),.din(w_dff_A_Iq2PYwmo5_1),.clk(gclk));
	jdff dff_A_lfKF9niy6_1(.dout(w_dff_A_Iq2PYwmo5_1),.din(w_dff_A_lfKF9niy6_1),.clk(gclk));
	jdff dff_A_pmBDn31b6_1(.dout(w_dff_A_lfKF9niy6_1),.din(w_dff_A_pmBDn31b6_1),.clk(gclk));
	jdff dff_A_W8PxzLLF1_1(.dout(w_dff_A_pmBDn31b6_1),.din(w_dff_A_W8PxzLLF1_1),.clk(gclk));
	jdff dff_A_xjJsVOJO5_1(.dout(w_dff_A_W8PxzLLF1_1),.din(w_dff_A_xjJsVOJO5_1),.clk(gclk));
	jdff dff_A_fNhn1uZ19_1(.dout(w_dff_A_xjJsVOJO5_1),.din(w_dff_A_fNhn1uZ19_1),.clk(gclk));
	jdff dff_A_ugVYufGk2_1(.dout(w_dff_A_fNhn1uZ19_1),.din(w_dff_A_ugVYufGk2_1),.clk(gclk));
	jdff dff_A_1xdISX657_1(.dout(w_dff_A_ugVYufGk2_1),.din(w_dff_A_1xdISX657_1),.clk(gclk));
	jdff dff_A_W9ZblWwJ6_1(.dout(w_dff_A_1xdISX657_1),.din(w_dff_A_W9ZblWwJ6_1),.clk(gclk));
	jdff dff_A_o4UjdsTI3_1(.dout(w_dff_A_W9ZblWwJ6_1),.din(w_dff_A_o4UjdsTI3_1),.clk(gclk));
	jdff dff_A_6iqiNvZX1_1(.dout(w_dff_A_o4UjdsTI3_1),.din(w_dff_A_6iqiNvZX1_1),.clk(gclk));
	jdff dff_A_Y3GMXjN15_1(.dout(w_dff_A_6iqiNvZX1_1),.din(w_dff_A_Y3GMXjN15_1),.clk(gclk));
	jdff dff_A_sZMFraKx5_1(.dout(w_dff_A_Y3GMXjN15_1),.din(w_dff_A_sZMFraKx5_1),.clk(gclk));
	jdff dff_A_tq65jwS84_1(.dout(w_dff_A_sZMFraKx5_1),.din(w_dff_A_tq65jwS84_1),.clk(gclk));
	jdff dff_A_7jupj86t9_0(.dout(w_n435_0[0]),.din(w_dff_A_7jupj86t9_0),.clk(gclk));
	jdff dff_A_9dsEoGvg6_0(.dout(w_dff_A_7jupj86t9_0),.din(w_dff_A_9dsEoGvg6_0),.clk(gclk));
	jdff dff_B_izHlvbbm7_0(.din(G156),.dout(w_dff_B_izHlvbbm7_0),.clk(gclk));
	jdff dff_B_tyt6915Y6_2(.din(n434),.dout(w_dff_B_tyt6915Y6_2),.clk(gclk));
	jdff dff_B_pwi9h59w5_2(.din(w_dff_B_tyt6915Y6_2),.dout(w_dff_B_pwi9h59w5_2),.clk(gclk));
	jdff dff_A_zLwudB9B5_2(.dout(w_G2239_0[2]),.din(w_dff_A_zLwudB9B5_2),.clk(gclk));
	jdff dff_A_h8kQPKRa5_2(.dout(w_dff_A_zLwudB9B5_2),.din(w_dff_A_h8kQPKRa5_2),.clk(gclk));
	jdff dff_A_FZhp2flj2_2(.dout(w_dff_A_h8kQPKRa5_2),.din(w_dff_A_FZhp2flj2_2),.clk(gclk));
	jdff dff_A_qd8jTaPx2_2(.dout(w_dff_A_FZhp2flj2_2),.din(w_dff_A_qd8jTaPx2_2),.clk(gclk));
	jdff dff_A_AlzcVAKM9_0(.dout(w_n433_1[0]),.din(w_dff_A_AlzcVAKM9_0),.clk(gclk));
	jdff dff_A_v8n0XNNu5_0(.dout(w_dff_A_AlzcVAKM9_0),.din(w_dff_A_v8n0XNNu5_0),.clk(gclk));
	jdff dff_A_Jo1ugJtU2_0(.dout(w_dff_A_v8n0XNNu5_0),.din(w_dff_A_Jo1ugJtU2_0),.clk(gclk));
	jdff dff_A_HuFmlrno0_0(.dout(w_dff_A_Jo1ugJtU2_0),.din(w_dff_A_HuFmlrno0_0),.clk(gclk));
	jdff dff_A_W8Uej57R9_0(.dout(w_dff_A_HuFmlrno0_0),.din(w_dff_A_W8Uej57R9_0),.clk(gclk));
	jdff dff_A_kUCYf8kN2_0(.dout(w_dff_A_W8Uej57R9_0),.din(w_dff_A_kUCYf8kN2_0),.clk(gclk));
	jdff dff_A_q113nbdl4_0(.dout(w_dff_A_kUCYf8kN2_0),.din(w_dff_A_q113nbdl4_0),.clk(gclk));
	jdff dff_A_uQdRHUcm2_0(.dout(w_dff_A_q113nbdl4_0),.din(w_dff_A_uQdRHUcm2_0),.clk(gclk));
	jdff dff_A_dn66hNLH8_0(.dout(w_dff_A_uQdRHUcm2_0),.din(w_dff_A_dn66hNLH8_0),.clk(gclk));
	jdff dff_A_al6QU0vJ8_0(.dout(w_dff_A_dn66hNLH8_0),.din(w_dff_A_al6QU0vJ8_0),.clk(gclk));
	jdff dff_A_SgCnDcuy9_0(.dout(w_dff_A_al6QU0vJ8_0),.din(w_dff_A_SgCnDcuy9_0),.clk(gclk));
	jdff dff_A_GmdPsuQo1_0(.dout(w_dff_A_SgCnDcuy9_0),.din(w_dff_A_GmdPsuQo1_0),.clk(gclk));
	jdff dff_A_cLtwMcub9_0(.dout(w_dff_A_GmdPsuQo1_0),.din(w_dff_A_cLtwMcub9_0),.clk(gclk));
	jdff dff_A_KaPls0NG1_0(.dout(w_dff_A_cLtwMcub9_0),.din(w_dff_A_KaPls0NG1_0),.clk(gclk));
	jdff dff_A_AX3bxqO52_0(.dout(w_dff_A_KaPls0NG1_0),.din(w_dff_A_AX3bxqO52_0),.clk(gclk));
	jdff dff_A_ycP2fRZk4_0(.dout(w_dff_A_AX3bxqO52_0),.din(w_dff_A_ycP2fRZk4_0),.clk(gclk));
	jdff dff_A_e8tZFNsW7_0(.dout(w_dff_A_ycP2fRZk4_0),.din(w_dff_A_e8tZFNsW7_0),.clk(gclk));
	jdff dff_A_D74tUqf23_0(.dout(w_dff_A_e8tZFNsW7_0),.din(w_dff_A_D74tUqf23_0),.clk(gclk));
	jdff dff_A_wEIpCUQT9_0(.dout(w_dff_A_D74tUqf23_0),.din(w_dff_A_wEIpCUQT9_0),.clk(gclk));
	jdff dff_A_Bo2UcP7W5_0(.dout(w_dff_A_wEIpCUQT9_0),.din(w_dff_A_Bo2UcP7W5_0),.clk(gclk));
	jdff dff_A_5tmLieRe6_0(.dout(w_dff_A_Bo2UcP7W5_0),.din(w_dff_A_5tmLieRe6_0),.clk(gclk));
	jdff dff_A_iFw9RA5e3_0(.dout(w_dff_A_5tmLieRe6_0),.din(w_dff_A_iFw9RA5e3_0),.clk(gclk));
	jdff dff_A_qpvyfEgP9_0(.dout(w_dff_A_iFw9RA5e3_0),.din(w_dff_A_qpvyfEgP9_0),.clk(gclk));
	jdff dff_A_VOzBRYgO8_0(.dout(w_dff_A_qpvyfEgP9_0),.din(w_dff_A_VOzBRYgO8_0),.clk(gclk));
	jdff dff_A_vbI13Ixl4_0(.dout(w_dff_A_VOzBRYgO8_0),.din(w_dff_A_vbI13Ixl4_0),.clk(gclk));
	jdff dff_A_gzmndNtt5_0(.dout(w_dff_A_vbI13Ixl4_0),.din(w_dff_A_gzmndNtt5_0),.clk(gclk));
	jdff dff_A_rYllZkbH4_0(.dout(w_dff_A_gzmndNtt5_0),.din(w_dff_A_rYllZkbH4_0),.clk(gclk));
	jdff dff_A_30iM3TXy2_0(.dout(w_dff_A_rYllZkbH4_0),.din(w_dff_A_30iM3TXy2_0),.clk(gclk));
	jdff dff_A_I0MZ7KOz8_2(.dout(w_n433_0[2]),.din(w_dff_A_I0MZ7KOz8_2),.clk(gclk));
	jdff dff_A_cN3hT0l91_2(.dout(w_dff_A_I0MZ7KOz8_2),.din(w_dff_A_cN3hT0l91_2),.clk(gclk));
	jdff dff_A_mQ10DAUR1_2(.dout(w_dff_A_cN3hT0l91_2),.din(w_dff_A_mQ10DAUR1_2),.clk(gclk));
	jdff dff_A_HEOQgHfq2_2(.dout(w_dff_A_mQ10DAUR1_2),.din(w_dff_A_HEOQgHfq2_2),.clk(gclk));
	jdff dff_A_nyssFGsN8_0(.dout(w_n431_0[0]),.din(w_dff_A_nyssFGsN8_0),.clk(gclk));
	jdff dff_A_xlQYpSbL7_0(.dout(w_dff_A_nyssFGsN8_0),.din(w_dff_A_xlQYpSbL7_0),.clk(gclk));
	jdff dff_B_pPgfFLMk6_0(.din(G155),.dout(w_dff_B_pPgfFLMk6_0),.clk(gclk));
	jdff dff_B_crLlfJIw9_2(.din(n430),.dout(w_dff_B_crLlfJIw9_2),.clk(gclk));
	jdff dff_B_yLX4YxfI0_2(.din(w_dff_B_crLlfJIw9_2),.dout(w_dff_B_yLX4YxfI0_2),.clk(gclk));
	jdff dff_A_89EwIiis5_1(.dout(w_n429_0[1]),.din(w_dff_A_89EwIiis5_1),.clk(gclk));
	jdff dff_A_4QrBMBET5_1(.dout(w_dff_A_89EwIiis5_1),.din(w_dff_A_4QrBMBET5_1),.clk(gclk));
	jdff dff_A_6K5JmWpr5_1(.dout(w_dff_A_4QrBMBET5_1),.din(w_dff_A_6K5JmWpr5_1),.clk(gclk));
	jdff dff_A_eWcErX501_1(.dout(w_dff_A_6K5JmWpr5_1),.din(w_dff_A_eWcErX501_1),.clk(gclk));
	jdff dff_A_tv0ZjUZ57_1(.dout(w_dff_A_eWcErX501_1),.din(w_dff_A_tv0ZjUZ57_1),.clk(gclk));
	jdff dff_A_oVUZjhSq8_1(.dout(w_dff_A_tv0ZjUZ57_1),.din(w_dff_A_oVUZjhSq8_1),.clk(gclk));
	jdff dff_A_3g6Hn5Wv6_1(.dout(w_dff_A_oVUZjhSq8_1),.din(w_dff_A_3g6Hn5Wv6_1),.clk(gclk));
	jdff dff_A_lD5UgCw14_1(.dout(w_dff_A_3g6Hn5Wv6_1),.din(w_dff_A_lD5UgCw14_1),.clk(gclk));
	jdff dff_A_djG3bFr94_1(.dout(w_dff_A_lD5UgCw14_1),.din(w_dff_A_djG3bFr94_1),.clk(gclk));
	jdff dff_A_fh94tmfL3_1(.dout(w_dff_A_djG3bFr94_1),.din(w_dff_A_fh94tmfL3_1),.clk(gclk));
	jdff dff_A_AIwIqTYA4_1(.dout(w_dff_A_fh94tmfL3_1),.din(w_dff_A_AIwIqTYA4_1),.clk(gclk));
	jdff dff_A_IEwPQ85E2_1(.dout(w_dff_A_AIwIqTYA4_1),.din(w_dff_A_IEwPQ85E2_1),.clk(gclk));
	jdff dff_A_OrKqRh162_1(.dout(w_dff_A_IEwPQ85E2_1),.din(w_dff_A_OrKqRh162_1),.clk(gclk));
	jdff dff_A_okEJVrfg6_1(.dout(w_dff_A_OrKqRh162_1),.din(w_dff_A_okEJVrfg6_1),.clk(gclk));
	jdff dff_A_nw04RoSO9_1(.dout(w_dff_A_okEJVrfg6_1),.din(w_dff_A_nw04RoSO9_1),.clk(gclk));
	jdff dff_A_WmPSiICV0_1(.dout(w_dff_A_nw04RoSO9_1),.din(w_dff_A_WmPSiICV0_1),.clk(gclk));
	jdff dff_A_m7AHlMkS4_1(.dout(w_dff_A_WmPSiICV0_1),.din(w_dff_A_m7AHlMkS4_1),.clk(gclk));
	jdff dff_A_VKcbacxA9_1(.dout(w_dff_A_m7AHlMkS4_1),.din(w_dff_A_VKcbacxA9_1),.clk(gclk));
	jdff dff_A_ehaYp7VW2_1(.dout(w_dff_A_VKcbacxA9_1),.din(w_dff_A_ehaYp7VW2_1),.clk(gclk));
	jdff dff_A_UBHMCOdy3_1(.dout(w_dff_A_ehaYp7VW2_1),.din(w_dff_A_UBHMCOdy3_1),.clk(gclk));
	jdff dff_A_jesx9sLH6_1(.dout(w_dff_A_UBHMCOdy3_1),.din(w_dff_A_jesx9sLH6_1),.clk(gclk));
	jdff dff_A_PCNN4v9u3_1(.dout(w_dff_A_jesx9sLH6_1),.din(w_dff_A_PCNN4v9u3_1),.clk(gclk));
	jdff dff_A_tSFY5sVH4_1(.dout(w_dff_A_PCNN4v9u3_1),.din(w_dff_A_tSFY5sVH4_1),.clk(gclk));
	jdff dff_A_hVxrw2tu1_1(.dout(w_dff_A_tSFY5sVH4_1),.din(w_dff_A_hVxrw2tu1_1),.clk(gclk));
	jdff dff_A_Mr3Sy99q2_1(.dout(w_dff_A_hVxrw2tu1_1),.din(w_dff_A_Mr3Sy99q2_1),.clk(gclk));
	jdff dff_A_jD4VLyHv4_1(.dout(w_dff_A_Mr3Sy99q2_1),.din(w_dff_A_jD4VLyHv4_1),.clk(gclk));
	jdff dff_A_ap7CsYDg3_1(.dout(w_dff_A_jD4VLyHv4_1),.din(w_dff_A_ap7CsYDg3_1),.clk(gclk));
	jdff dff_A_9jLdaajW3_1(.dout(w_dff_A_ap7CsYDg3_1),.din(w_dff_A_9jLdaajW3_1),.clk(gclk));
	jdff dff_A_3hHbEkJw4_2(.dout(w_n429_0[2]),.din(w_dff_A_3hHbEkJw4_2),.clk(gclk));
	jdff dff_A_8axD2BKd8_0(.dout(w_n427_0[0]),.din(w_dff_A_8axD2BKd8_0),.clk(gclk));
	jdff dff_A_LH9Vwqk78_0(.dout(w_dff_A_8axD2BKd8_0),.din(w_dff_A_LH9Vwqk78_0),.clk(gclk));
	jdff dff_B_pvlpNQrM0_0(.din(G154),.dout(w_dff_B_pvlpNQrM0_0),.clk(gclk));
	jdff dff_A_4rk7qgCu2_1(.dout(w_n426_0[1]),.din(w_dff_A_4rk7qgCu2_1),.clk(gclk));
	jdff dff_A_pev09nyh0_1(.dout(w_dff_A_4rk7qgCu2_1),.din(w_dff_A_pev09nyh0_1),.clk(gclk));
	jdff dff_A_guDKXsto8_2(.dout(w_n426_0[2]),.din(w_dff_A_guDKXsto8_2),.clk(gclk));
	jdff dff_A_jXiXJTM48_2(.dout(w_dff_A_guDKXsto8_2),.din(w_dff_A_jXiXJTM48_2),.clk(gclk));
	jdff dff_A_9yVFVzBQ3_1(.dout(w_G2253_0[1]),.din(w_dff_A_9yVFVzBQ3_1),.clk(gclk));
	jdff dff_A_F7C2nutF1_1(.dout(w_dff_A_9yVFVzBQ3_1),.din(w_dff_A_F7C2nutF1_1),.clk(gclk));
	jdff dff_A_uDvPeQvH9_1(.dout(w_dff_A_F7C2nutF1_1),.din(w_dff_A_uDvPeQvH9_1),.clk(gclk));
	jdff dff_A_frfO4gwx4_1(.dout(w_dff_A_uDvPeQvH9_1),.din(w_dff_A_frfO4gwx4_1),.clk(gclk));
	jdff dff_A_WDOYyWZJ6_1(.dout(w_n425_1[1]),.din(w_dff_A_WDOYyWZJ6_1),.clk(gclk));
	jdff dff_A_snsW2rGW9_1(.dout(w_dff_A_WDOYyWZJ6_1),.din(w_dff_A_snsW2rGW9_1),.clk(gclk));
	jdff dff_A_UoATPuIy5_1(.dout(w_dff_A_snsW2rGW9_1),.din(w_dff_A_UoATPuIy5_1),.clk(gclk));
	jdff dff_A_cQUnQXGj7_1(.dout(w_dff_A_UoATPuIy5_1),.din(w_dff_A_cQUnQXGj7_1),.clk(gclk));
	jdff dff_A_JZORpoAV6_1(.dout(w_dff_A_cQUnQXGj7_1),.din(w_dff_A_JZORpoAV6_1),.clk(gclk));
	jdff dff_A_08ZtQnWK9_1(.dout(w_dff_A_JZORpoAV6_1),.din(w_dff_A_08ZtQnWK9_1),.clk(gclk));
	jdff dff_A_zeoIeoUY5_1(.dout(w_dff_A_08ZtQnWK9_1),.din(w_dff_A_zeoIeoUY5_1),.clk(gclk));
	jdff dff_A_Y6WMetcc5_1(.dout(w_dff_A_zeoIeoUY5_1),.din(w_dff_A_Y6WMetcc5_1),.clk(gclk));
	jdff dff_A_FcIjmJT88_1(.dout(w_dff_A_Y6WMetcc5_1),.din(w_dff_A_FcIjmJT88_1),.clk(gclk));
	jdff dff_A_2eb6slmX3_1(.dout(w_dff_A_FcIjmJT88_1),.din(w_dff_A_2eb6slmX3_1),.clk(gclk));
	jdff dff_A_0YdkfY6u0_1(.dout(w_dff_A_2eb6slmX3_1),.din(w_dff_A_0YdkfY6u0_1),.clk(gclk));
	jdff dff_A_gGaIcq9W3_1(.dout(w_dff_A_0YdkfY6u0_1),.din(w_dff_A_gGaIcq9W3_1),.clk(gclk));
	jdff dff_A_kBnKYt0K2_1(.dout(w_dff_A_gGaIcq9W3_1),.din(w_dff_A_kBnKYt0K2_1),.clk(gclk));
	jdff dff_A_YcTFhvGB5_1(.dout(w_dff_A_kBnKYt0K2_1),.din(w_dff_A_YcTFhvGB5_1),.clk(gclk));
	jdff dff_A_kpUOp8HU8_1(.dout(w_dff_A_YcTFhvGB5_1),.din(w_dff_A_kpUOp8HU8_1),.clk(gclk));
	jdff dff_A_DepCaV7C1_1(.dout(w_dff_A_kpUOp8HU8_1),.din(w_dff_A_DepCaV7C1_1),.clk(gclk));
	jdff dff_A_4TZPQH0r0_1(.dout(w_dff_A_DepCaV7C1_1),.din(w_dff_A_4TZPQH0r0_1),.clk(gclk));
	jdff dff_A_3DskEiN37_1(.dout(w_dff_A_4TZPQH0r0_1),.din(w_dff_A_3DskEiN37_1),.clk(gclk));
	jdff dff_A_34dwUmOG1_1(.dout(w_dff_A_3DskEiN37_1),.din(w_dff_A_34dwUmOG1_1),.clk(gclk));
	jdff dff_A_sRtAdeT96_1(.dout(w_dff_A_34dwUmOG1_1),.din(w_dff_A_sRtAdeT96_1),.clk(gclk));
	jdff dff_A_MNoAWPjX9_1(.dout(w_dff_A_sRtAdeT96_1),.din(w_dff_A_MNoAWPjX9_1),.clk(gclk));
	jdff dff_A_8rxtEIsp6_1(.dout(w_dff_A_MNoAWPjX9_1),.din(w_dff_A_8rxtEIsp6_1),.clk(gclk));
	jdff dff_A_nmnVDEYr4_1(.dout(w_dff_A_8rxtEIsp6_1),.din(w_dff_A_nmnVDEYr4_1),.clk(gclk));
	jdff dff_A_hAWpOiWd7_1(.dout(w_dff_A_nmnVDEYr4_1),.din(w_dff_A_hAWpOiWd7_1),.clk(gclk));
	jdff dff_A_v8tUjL8T1_1(.dout(w_dff_A_hAWpOiWd7_1),.din(w_dff_A_v8tUjL8T1_1),.clk(gclk));
	jdff dff_A_05tgbhy02_1(.dout(w_dff_A_v8tUjL8T1_1),.din(w_dff_A_05tgbhy02_1),.clk(gclk));
	jdff dff_A_4MiPJ3LA3_1(.dout(w_dff_A_05tgbhy02_1),.din(w_dff_A_4MiPJ3LA3_1),.clk(gclk));
	jdff dff_A_YgznzAnD1_1(.dout(w_dff_A_4MiPJ3LA3_1),.din(w_dff_A_YgznzAnD1_1),.clk(gclk));
	jdff dff_A_nfmxpdLb1_2(.dout(w_n425_0[2]),.din(w_dff_A_nfmxpdLb1_2),.clk(gclk));
	jdff dff_A_ViNW4HgW0_2(.dout(w_dff_A_nfmxpdLb1_2),.din(w_dff_A_ViNW4HgW0_2),.clk(gclk));
	jdff dff_A_uUmampzn9_2(.dout(w_dff_A_ViNW4HgW0_2),.din(w_dff_A_uUmampzn9_2),.clk(gclk));
	jdff dff_A_FlRIwn5i0_2(.dout(w_dff_A_uUmampzn9_2),.din(w_dff_A_FlRIwn5i0_2),.clk(gclk));
	jdff dff_A_zbBR5lUA8_2(.dout(w_dff_A_FlRIwn5i0_2),.din(w_dff_A_zbBR5lUA8_2),.clk(gclk));
	jdff dff_A_U9vXyqPk9_2(.dout(w_dff_A_zbBR5lUA8_2),.din(w_dff_A_U9vXyqPk9_2),.clk(gclk));
	jdff dff_A_9jIVbu968_2(.dout(w_dff_A_U9vXyqPk9_2),.din(w_dff_A_9jIVbu968_2),.clk(gclk));
	jdff dff_A_sPaykXaM7_2(.dout(w_dff_A_9jIVbu968_2),.din(w_dff_A_sPaykXaM7_2),.clk(gclk));
	jdff dff_A_BrJWuiaC8_2(.dout(w_dff_A_sPaykXaM7_2),.din(w_dff_A_BrJWuiaC8_2),.clk(gclk));
	jdff dff_A_pBcZMKd46_2(.dout(w_dff_A_BrJWuiaC8_2),.din(w_dff_A_pBcZMKd46_2),.clk(gclk));
	jdff dff_A_cbDPx23U4_2(.dout(w_dff_A_pBcZMKd46_2),.din(w_dff_A_cbDPx23U4_2),.clk(gclk));
	jdff dff_A_IM4vO9031_2(.dout(w_dff_A_cbDPx23U4_2),.din(w_dff_A_IM4vO9031_2),.clk(gclk));
	jdff dff_A_7aLLXZtZ3_2(.dout(w_dff_A_IM4vO9031_2),.din(w_dff_A_7aLLXZtZ3_2),.clk(gclk));
	jdff dff_A_thblUgG17_2(.dout(w_dff_A_7aLLXZtZ3_2),.din(w_dff_A_thblUgG17_2),.clk(gclk));
	jdff dff_A_v28JbT4a6_2(.dout(w_dff_A_thblUgG17_2),.din(w_dff_A_v28JbT4a6_2),.clk(gclk));
	jdff dff_A_3cqgQiJx0_2(.dout(w_dff_A_v28JbT4a6_2),.din(w_dff_A_3cqgQiJx0_2),.clk(gclk));
	jdff dff_A_GKzDMjvo6_2(.dout(w_dff_A_3cqgQiJx0_2),.din(w_dff_A_GKzDMjvo6_2),.clk(gclk));
	jdff dff_A_ICIwWuyt6_2(.dout(w_dff_A_GKzDMjvo6_2),.din(w_dff_A_ICIwWuyt6_2),.clk(gclk));
	jdff dff_A_OeNZrCCi6_2(.dout(w_dff_A_ICIwWuyt6_2),.din(w_dff_A_OeNZrCCi6_2),.clk(gclk));
	jdff dff_A_kOs2V4Nv4_2(.dout(w_dff_A_OeNZrCCi6_2),.din(w_dff_A_kOs2V4Nv4_2),.clk(gclk));
	jdff dff_A_ilpsLJRE7_2(.dout(w_dff_A_kOs2V4Nv4_2),.din(w_dff_A_ilpsLJRE7_2),.clk(gclk));
	jdff dff_A_Br6KRhQR9_2(.dout(w_dff_A_ilpsLJRE7_2),.din(w_dff_A_Br6KRhQR9_2),.clk(gclk));
	jdff dff_A_FJAcj8Gr8_2(.dout(w_dff_A_Br6KRhQR9_2),.din(w_dff_A_FJAcj8Gr8_2),.clk(gclk));
	jdff dff_A_loqtJTl15_2(.dout(w_dff_A_FJAcj8Gr8_2),.din(w_dff_A_loqtJTl15_2),.clk(gclk));
	jdff dff_A_FOEQd2I65_2(.dout(w_dff_A_loqtJTl15_2),.din(w_dff_A_FOEQd2I65_2),.clk(gclk));
	jdff dff_A_wbREUSQ84_2(.dout(w_dff_A_FOEQd2I65_2),.din(w_dff_A_wbREUSQ84_2),.clk(gclk));
	jdff dff_A_f32nalKt1_2(.dout(w_dff_A_wbREUSQ84_2),.din(w_dff_A_f32nalKt1_2),.clk(gclk));
	jdff dff_A_Inqk3ZfN9_2(.dout(w_dff_A_f32nalKt1_2),.din(w_dff_A_Inqk3ZfN9_2),.clk(gclk));
	jdff dff_A_QFFXqi4l6_1(.dout(w_n424_0[1]),.din(w_dff_A_QFFXqi4l6_1),.clk(gclk));
	jdff dff_A_O5vJ67dP6_1(.dout(w_dff_A_QFFXqi4l6_1),.din(w_dff_A_O5vJ67dP6_1),.clk(gclk));
	jdff dff_A_EordcHI36_1(.dout(w_dff_A_O5vJ67dP6_1),.din(w_dff_A_EordcHI36_1),.clk(gclk));
	jdff dff_A_KlMKcVk09_1(.dout(w_dff_A_EordcHI36_1),.din(w_dff_A_KlMKcVk09_1),.clk(gclk));
	jdff dff_A_NiwAgNE42_1(.dout(w_dff_A_KlMKcVk09_1),.din(w_dff_A_NiwAgNE42_1),.clk(gclk));
	jdff dff_A_i48I0sIY1_1(.dout(w_dff_A_NiwAgNE42_1),.din(w_dff_A_i48I0sIY1_1),.clk(gclk));
	jdff dff_A_zmM9YdNU5_1(.dout(w_dff_A_i48I0sIY1_1),.din(w_dff_A_zmM9YdNU5_1),.clk(gclk));
	jdff dff_A_20t1uaI64_1(.dout(w_dff_A_zmM9YdNU5_1),.din(w_dff_A_20t1uaI64_1),.clk(gclk));
	jdff dff_A_Q55RE2jL8_1(.dout(w_dff_A_20t1uaI64_1),.din(w_dff_A_Q55RE2jL8_1),.clk(gclk));
	jdff dff_A_BQ9zBtmF0_1(.dout(w_dff_A_Q55RE2jL8_1),.din(w_dff_A_BQ9zBtmF0_1),.clk(gclk));
	jdff dff_A_8yxk20K62_1(.dout(w_dff_A_BQ9zBtmF0_1),.din(w_dff_A_8yxk20K62_1),.clk(gclk));
	jdff dff_A_zuVLIfE58_1(.dout(w_dff_A_8yxk20K62_1),.din(w_dff_A_zuVLIfE58_1),.clk(gclk));
	jdff dff_A_hSSvffpZ8_1(.dout(w_dff_A_zuVLIfE58_1),.din(w_dff_A_hSSvffpZ8_1),.clk(gclk));
	jdff dff_A_wPLjj0o73_1(.dout(w_dff_A_hSSvffpZ8_1),.din(w_dff_A_wPLjj0o73_1),.clk(gclk));
	jdff dff_A_a3104nWL0_1(.dout(w_dff_A_wPLjj0o73_1),.din(w_dff_A_a3104nWL0_1),.clk(gclk));
	jdff dff_A_WaqrZ3HL7_1(.dout(w_dff_A_a3104nWL0_1),.din(w_dff_A_WaqrZ3HL7_1),.clk(gclk));
	jdff dff_A_Gvx5zwgd8_1(.dout(w_dff_A_WaqrZ3HL7_1),.din(w_dff_A_Gvx5zwgd8_1),.clk(gclk));
	jdff dff_A_4TlbubFC3_1(.dout(w_dff_A_Gvx5zwgd8_1),.din(w_dff_A_4TlbubFC3_1),.clk(gclk));
	jdff dff_A_N13YSZie3_1(.dout(w_dff_A_4TlbubFC3_1),.din(w_dff_A_N13YSZie3_1),.clk(gclk));
	jdff dff_A_PnztjSvN8_1(.dout(w_dff_A_N13YSZie3_1),.din(w_dff_A_PnztjSvN8_1),.clk(gclk));
	jdff dff_A_bFibu95c6_1(.dout(w_dff_A_PnztjSvN8_1),.din(w_dff_A_bFibu95c6_1),.clk(gclk));
	jdff dff_A_2JN3ySKm1_1(.dout(w_dff_A_bFibu95c6_1),.din(w_dff_A_2JN3ySKm1_1),.clk(gclk));
	jdff dff_A_mgyvRonx9_1(.dout(w_dff_A_2JN3ySKm1_1),.din(w_dff_A_mgyvRonx9_1),.clk(gclk));
	jdff dff_A_y2pkpJJP4_1(.dout(w_dff_A_mgyvRonx9_1),.din(w_dff_A_y2pkpJJP4_1),.clk(gclk));
	jdff dff_A_VWfB6z6I2_1(.dout(w_dff_A_y2pkpJJP4_1),.din(w_dff_A_VWfB6z6I2_1),.clk(gclk));
	jdff dff_A_pyjGeP4F9_1(.dout(w_dff_A_VWfB6z6I2_1),.din(w_dff_A_pyjGeP4F9_1),.clk(gclk));
	jdff dff_A_2ltKX4H53_1(.dout(w_dff_A_pyjGeP4F9_1),.din(w_dff_A_2ltKX4H53_1),.clk(gclk));
	jdff dff_A_DHeldumB4_1(.dout(w_dff_A_2ltKX4H53_1),.din(w_dff_A_DHeldumB4_1),.clk(gclk));
	jdff dff_A_CSmNRdhO9_1(.dout(w_dff_A_DHeldumB4_1),.din(w_dff_A_CSmNRdhO9_1),.clk(gclk));
	jdff dff_A_NlcaFYkA4_0(.dout(w_n422_0[0]),.din(w_dff_A_NlcaFYkA4_0),.clk(gclk));
	jdff dff_A_LlyypmAA3_0(.dout(w_dff_A_NlcaFYkA4_0),.din(w_dff_A_LlyypmAA3_0),.clk(gclk));
	jdff dff_B_zfCEdJOT5_0(.din(G153),.dout(w_dff_B_zfCEdJOT5_0),.clk(gclk));
	jdff dff_A_BhsS0mFn0_1(.dout(w_n421_0[1]),.din(w_dff_A_BhsS0mFn0_1),.clk(gclk));
	jdff dff_A_AczDAVgJ8_1(.dout(w_dff_A_BhsS0mFn0_1),.din(w_dff_A_AczDAVgJ8_1),.clk(gclk));
	jdff dff_A_7rlPCFmP0_2(.dout(w_n421_0[2]),.din(w_dff_A_7rlPCFmP0_2),.clk(gclk));
	jdff dff_A_0BKpP0JF3_2(.dout(w_dff_A_7rlPCFmP0_2),.din(w_dff_A_0BKpP0JF3_2),.clk(gclk));
	jdff dff_A_iyFxE0WN7_1(.dout(w_n416_0[1]),.din(w_dff_A_iyFxE0WN7_1),.clk(gclk));
	jdff dff_A_0p0bLv4h5_1(.dout(w_dff_A_iyFxE0WN7_1),.din(w_dff_A_0p0bLv4h5_1),.clk(gclk));
	jdff dff_A_rTrW1eUT5_1(.dout(w_dff_A_0p0bLv4h5_1),.din(w_dff_A_rTrW1eUT5_1),.clk(gclk));
	jdff dff_A_4GrWIc1s1_1(.dout(w_dff_A_rTrW1eUT5_1),.din(w_dff_A_4GrWIc1s1_1),.clk(gclk));
	jdff dff_A_NTQ1reO15_1(.dout(w_dff_A_4GrWIc1s1_1),.din(w_dff_A_NTQ1reO15_1),.clk(gclk));
	jdff dff_A_IiPd0a298_1(.dout(w_dff_A_NTQ1reO15_1),.din(w_dff_A_IiPd0a298_1),.clk(gclk));
	jdff dff_A_u0Xv4gTN7_1(.dout(w_dff_A_IiPd0a298_1),.din(w_dff_A_u0Xv4gTN7_1),.clk(gclk));
	jdff dff_A_7nLFGb9G2_1(.dout(w_dff_A_u0Xv4gTN7_1),.din(w_dff_A_7nLFGb9G2_1),.clk(gclk));
	jdff dff_A_PXQxivjl1_1(.dout(w_dff_A_7nLFGb9G2_1),.din(w_dff_A_PXQxivjl1_1),.clk(gclk));
	jdff dff_A_NNCNc2w56_1(.dout(w_dff_A_PXQxivjl1_1),.din(w_dff_A_NNCNc2w56_1),.clk(gclk));
	jdff dff_A_jcUFpHuc8_1(.dout(w_dff_A_NNCNc2w56_1),.din(w_dff_A_jcUFpHuc8_1),.clk(gclk));
	jdff dff_A_WDfCFM9k1_1(.dout(w_dff_A_jcUFpHuc8_1),.din(w_dff_A_WDfCFM9k1_1),.clk(gclk));
	jdff dff_A_v1AG3zii7_1(.dout(w_dff_A_WDfCFM9k1_1),.din(w_dff_A_v1AG3zii7_1),.clk(gclk));
	jdff dff_A_EoMrbiIW1_1(.dout(w_dff_A_v1AG3zii7_1),.din(w_dff_A_EoMrbiIW1_1),.clk(gclk));
	jdff dff_A_IkXlJV928_1(.dout(w_dff_A_EoMrbiIW1_1),.din(w_dff_A_IkXlJV928_1),.clk(gclk));
	jdff dff_A_TdtnEfxh9_1(.dout(w_dff_A_IkXlJV928_1),.din(w_dff_A_TdtnEfxh9_1),.clk(gclk));
	jdff dff_A_jHgTChG39_1(.dout(w_dff_A_TdtnEfxh9_1),.din(w_dff_A_jHgTChG39_1),.clk(gclk));
	jdff dff_A_5NzEaXDh7_1(.dout(w_dff_A_jHgTChG39_1),.din(w_dff_A_5NzEaXDh7_1),.clk(gclk));
	jdff dff_A_nEagDW6k0_1(.dout(w_dff_A_5NzEaXDh7_1),.din(w_dff_A_nEagDW6k0_1),.clk(gclk));
	jdff dff_A_AjcqR7Yg2_1(.dout(w_dff_A_nEagDW6k0_1),.din(w_dff_A_AjcqR7Yg2_1),.clk(gclk));
	jdff dff_A_JDaC1WEL3_1(.dout(w_dff_A_AjcqR7Yg2_1),.din(w_dff_A_JDaC1WEL3_1),.clk(gclk));
	jdff dff_A_Q1QpMwcF1_1(.dout(w_dff_A_JDaC1WEL3_1),.din(w_dff_A_Q1QpMwcF1_1),.clk(gclk));
	jdff dff_A_ClCaIhFk2_1(.dout(w_dff_A_Q1QpMwcF1_1),.din(w_dff_A_ClCaIhFk2_1),.clk(gclk));
	jdff dff_A_1yihF3513_1(.dout(w_dff_A_ClCaIhFk2_1),.din(w_dff_A_1yihF3513_1),.clk(gclk));
	jdff dff_A_xn5aMBvj8_1(.dout(w_dff_A_1yihF3513_1),.din(w_dff_A_xn5aMBvj8_1),.clk(gclk));
	jdff dff_A_6esJE98D4_1(.dout(w_dff_A_xn5aMBvj8_1),.din(w_dff_A_6esJE98D4_1),.clk(gclk));
	jdff dff_A_O2Q6WSYo9_1(.dout(w_dff_A_6esJE98D4_1),.din(w_dff_A_O2Q6WSYo9_1),.clk(gclk));
	jdff dff_A_5LsLCVbA5_1(.dout(w_dff_A_O2Q6WSYo9_1),.din(w_dff_A_5LsLCVbA5_1),.clk(gclk));
	jdff dff_A_ZZDoLTrp5_1(.dout(w_dff_A_5LsLCVbA5_1),.din(w_dff_A_ZZDoLTrp5_1),.clk(gclk));
	jdff dff_A_f4VrnYDr7_1(.dout(w_dff_A_ZZDoLTrp5_1),.din(w_dff_A_f4VrnYDr7_1),.clk(gclk));
	jdff dff_A_ton5okTs8_1(.dout(w_dff_A_f4VrnYDr7_1),.din(w_dff_A_ton5okTs8_1),.clk(gclk));
	jdff dff_A_alS2OU0O7_1(.dout(w_dff_A_ton5okTs8_1),.din(w_dff_A_alS2OU0O7_1),.clk(gclk));
	jdff dff_A_NIIPZnVf3_0(.dout(w_n378_0[0]),.din(w_dff_A_NIIPZnVf3_0),.clk(gclk));
	jdff dff_A_e43K4zLq2_0(.dout(w_dff_A_NIIPZnVf3_0),.din(w_dff_A_e43K4zLq2_0),.clk(gclk));
	jdff dff_B_l5zNm9Gi9_0(.din(G214),.dout(w_dff_B_l5zNm9Gi9_0),.clk(gclk));
	jdff dff_A_Ifa0eeTd3_1(.dout(w_n383_0[1]),.din(w_dff_A_Ifa0eeTd3_1),.clk(gclk));
	jdff dff_A_Dr6I3zdZ5_1(.dout(w_dff_A_Ifa0eeTd3_1),.din(w_dff_A_Dr6I3zdZ5_1),.clk(gclk));
	jdff dff_A_NewWcorh8_2(.dout(w_n383_0[2]),.din(w_dff_A_NewWcorh8_2),.clk(gclk));
	jdff dff_A_6dGCM4iH7_2(.dout(w_dff_A_NewWcorh8_2),.din(w_dff_A_6dGCM4iH7_2),.clk(gclk));
	jdff dff_A_DY1kktFA4_2(.dout(w_G1480_0[2]),.din(w_dff_A_DY1kktFA4_2),.clk(gclk));
	jdff dff_A_Mwxo8oJu9_2(.dout(w_dff_A_DY1kktFA4_2),.din(w_dff_A_Mwxo8oJu9_2),.clk(gclk));
	jdff dff_A_QK14DYwA1_2(.dout(w_dff_A_Mwxo8oJu9_2),.din(w_dff_A_QK14DYwA1_2),.clk(gclk));
	jdff dff_A_rB8GOIbM9_2(.dout(w_dff_A_QK14DYwA1_2),.din(w_dff_A_rB8GOIbM9_2),.clk(gclk));
	jdff dff_B_A4tUEeHk1_0(.din(G215),.dout(w_dff_B_A4tUEeHk1_0),.clk(gclk));
	jdff dff_B_DmC11cly1_2(.din(n385),.dout(w_dff_B_DmC11cly1_2),.clk(gclk));
	jdff dff_B_RleEmAtv9_2(.din(w_dff_B_DmC11cly1_2),.dout(w_dff_B_RleEmAtv9_2),.clk(gclk));
	jdff dff_A_hpoEgCU05_0(.dout(w_G106_1[0]),.din(w_dff_A_hpoEgCU05_0),.clk(gclk));
	jdff dff_A_7eMha8en1_0(.dout(w_dff_A_hpoEgCU05_0),.din(w_dff_A_7eMha8en1_0),.clk(gclk));
	jdff dff_A_RvVpfsPN9_0(.dout(w_dff_A_7eMha8en1_0),.din(w_dff_A_RvVpfsPN9_0),.clk(gclk));
	jdff dff_A_hwt4BvMM2_0(.dout(w_dff_A_RvVpfsPN9_0),.din(w_dff_A_hwt4BvMM2_0),.clk(gclk));
	jdff dff_B_103VmZWn5_1(.din(n1551),.dout(w_dff_B_103VmZWn5_1),.clk(gclk));
	jdff dff_B_agReMxmj6_1(.din(n1552),.dout(w_dff_B_agReMxmj6_1),.clk(gclk));
	jdff dff_B_93yrlnIL7_1(.din(w_dff_B_agReMxmj6_1),.dout(w_dff_B_93yrlnIL7_1),.clk(gclk));
	jdff dff_B_plq1XYuG0_1(.din(w_dff_B_93yrlnIL7_1),.dout(w_dff_B_plq1XYuG0_1),.clk(gclk));
	jdff dff_B_zgrmvCJ14_1(.din(w_dff_B_plq1XYuG0_1),.dout(w_dff_B_zgrmvCJ14_1),.clk(gclk));
	jdff dff_B_aAFM1OFQ8_1(.din(w_dff_B_zgrmvCJ14_1),.dout(w_dff_B_aAFM1OFQ8_1),.clk(gclk));
	jdff dff_B_FbAYhA0K9_1(.din(w_dff_B_aAFM1OFQ8_1),.dout(w_dff_B_FbAYhA0K9_1),.clk(gclk));
	jdff dff_B_rmoIH8jC0_1(.din(w_dff_B_FbAYhA0K9_1),.dout(w_dff_B_rmoIH8jC0_1),.clk(gclk));
	jdff dff_B_sPOB1pyl2_1(.din(w_dff_B_rmoIH8jC0_1),.dout(w_dff_B_sPOB1pyl2_1),.clk(gclk));
	jdff dff_B_6uk0RQrf1_1(.din(w_dff_B_sPOB1pyl2_1),.dout(w_dff_B_6uk0RQrf1_1),.clk(gclk));
	jdff dff_B_Kvf6QrTG2_1(.din(w_dff_B_6uk0RQrf1_1),.dout(w_dff_B_Kvf6QrTG2_1),.clk(gclk));
	jdff dff_B_NUAUviSo4_1(.din(w_dff_B_Kvf6QrTG2_1),.dout(w_dff_B_NUAUviSo4_1),.clk(gclk));
	jdff dff_B_3oV9plvU5_1(.din(w_dff_B_NUAUviSo4_1),.dout(w_dff_B_3oV9plvU5_1),.clk(gclk));
	jdff dff_B_mDdB53xk4_1(.din(w_dff_B_3oV9plvU5_1),.dout(w_dff_B_mDdB53xk4_1),.clk(gclk));
	jdff dff_B_UjeyhpaG1_1(.din(w_dff_B_mDdB53xk4_1),.dout(w_dff_B_UjeyhpaG1_1),.clk(gclk));
	jdff dff_B_IwQzJvZb6_0(.din(n1576),.dout(w_dff_B_IwQzJvZb6_0),.clk(gclk));
	jdff dff_B_aT7TYaF82_0(.din(w_dff_B_IwQzJvZb6_0),.dout(w_dff_B_aT7TYaF82_0),.clk(gclk));
	jdff dff_B_yjpXPO2h6_0(.din(w_dff_B_aT7TYaF82_0),.dout(w_dff_B_yjpXPO2h6_0),.clk(gclk));
	jdff dff_B_uPo0wcI66_0(.din(w_dff_B_yjpXPO2h6_0),.dout(w_dff_B_uPo0wcI66_0),.clk(gclk));
	jdff dff_B_z66APjTh5_0(.din(n1575),.dout(w_dff_B_z66APjTh5_0),.clk(gclk));
	jdff dff_B_C8X1P6Dm0_0(.din(w_dff_B_z66APjTh5_0),.dout(w_dff_B_C8X1P6Dm0_0),.clk(gclk));
	jdff dff_B_jYtn8H0s7_0(.din(n1572),.dout(w_dff_B_jYtn8H0s7_0),.clk(gclk));
	jdff dff_B_mJfFUkk79_0(.din(w_dff_B_jYtn8H0s7_0),.dout(w_dff_B_mJfFUkk79_0),.clk(gclk));
	jdff dff_B_fXaCUOCl5_0(.din(w_dff_B_mJfFUkk79_0),.dout(w_dff_B_fXaCUOCl5_0),.clk(gclk));
	jdff dff_B_moMo4PEw5_0(.din(n1568),.dout(w_dff_B_moMo4PEw5_0),.clk(gclk));
	jdff dff_B_CCxRpgky9_0(.din(w_dff_B_moMo4PEw5_0),.dout(w_dff_B_CCxRpgky9_0),.clk(gclk));
	jdff dff_B_vAnRDzCG8_1(.din(n1560),.dout(w_dff_B_vAnRDzCG8_1),.clk(gclk));
	jdff dff_B_tHfsW3vq4_1(.din(w_dff_B_vAnRDzCG8_1),.dout(w_dff_B_tHfsW3vq4_1),.clk(gclk));
	jdff dff_B_YY2AIPKe1_0(.din(n1563),.dout(w_dff_B_YY2AIPKe1_0),.clk(gclk));
	jdff dff_B_X6ducswn4_0(.din(w_dff_B_YY2AIPKe1_0),.dout(w_dff_B_X6ducswn4_0),.clk(gclk));
	jdff dff_B_kTVk2DZi1_0(.din(w_dff_B_X6ducswn4_0),.dout(w_dff_B_kTVk2DZi1_0),.clk(gclk));
	jdff dff_B_TDlfsMvs7_0(.din(w_dff_B_kTVk2DZi1_0),.dout(w_dff_B_TDlfsMvs7_0),.clk(gclk));
	jdff dff_B_4oBtaw2G0_0(.din(w_dff_B_TDlfsMvs7_0),.dout(w_dff_B_4oBtaw2G0_0),.clk(gclk));
	jdff dff_B_IlZDseQj4_0(.din(w_dff_B_4oBtaw2G0_0),.dout(w_dff_B_IlZDseQj4_0),.clk(gclk));
	jdff dff_B_fc44wMvx8_0(.din(w_dff_B_IlZDseQj4_0),.dout(w_dff_B_fc44wMvx8_0),.clk(gclk));
	jdff dff_A_TT291i8o6_0(.dout(w_n1562_0[0]),.din(w_dff_A_TT291i8o6_0),.clk(gclk));
	jdff dff_A_VhyWcYjA2_0(.dout(w_dff_A_TT291i8o6_0),.din(w_dff_A_VhyWcYjA2_0),.clk(gclk));
	jdff dff_A_sziBKZFJ9_0(.dout(w_dff_A_VhyWcYjA2_0),.din(w_dff_A_sziBKZFJ9_0),.clk(gclk));
	jdff dff_A_zUERrm125_0(.dout(w_dff_A_sziBKZFJ9_0),.din(w_dff_A_zUERrm125_0),.clk(gclk));
	jdff dff_A_b1SzQC9W3_0(.dout(w_dff_A_zUERrm125_0),.din(w_dff_A_b1SzQC9W3_0),.clk(gclk));
	jdff dff_A_732wFWfy2_0(.dout(w_dff_A_b1SzQC9W3_0),.din(w_dff_A_732wFWfy2_0),.clk(gclk));
	jdff dff_A_y1uIFPlM4_0(.dout(w_dff_A_732wFWfy2_0),.din(w_dff_A_y1uIFPlM4_0),.clk(gclk));
	jdff dff_A_GgwafJLG3_1(.dout(w_n1562_0[1]),.din(w_dff_A_GgwafJLG3_1),.clk(gclk));
	jdff dff_A_NXy2NtW05_1(.dout(w_dff_A_GgwafJLG3_1),.din(w_dff_A_NXy2NtW05_1),.clk(gclk));
	jdff dff_A_FD2nd6Wv3_1(.dout(w_dff_A_NXy2NtW05_1),.din(w_dff_A_FD2nd6Wv3_1),.clk(gclk));
	jdff dff_A_8TwFusgJ7_1(.dout(w_dff_A_FD2nd6Wv3_1),.din(w_dff_A_8TwFusgJ7_1),.clk(gclk));
	jdff dff_A_KCyGJCE62_1(.dout(w_dff_A_8TwFusgJ7_1),.din(w_dff_A_KCyGJCE62_1),.clk(gclk));
	jdff dff_A_kaQ6s8Sg9_1(.dout(w_dff_A_KCyGJCE62_1),.din(w_dff_A_kaQ6s8Sg9_1),.clk(gclk));
	jdff dff_A_7W0PCMHr4_1(.dout(w_dff_A_kaQ6s8Sg9_1),.din(w_dff_A_7W0PCMHr4_1),.clk(gclk));
	jdff dff_B_m84ttWlY6_0(.din(n1559),.dout(w_dff_B_m84ttWlY6_0),.clk(gclk));
	jdff dff_B_bt5CqlH54_0(.din(w_dff_B_m84ttWlY6_0),.dout(w_dff_B_bt5CqlH54_0),.clk(gclk));
	jdff dff_B_anNSMSO76_0(.din(w_dff_B_bt5CqlH54_0),.dout(w_dff_B_anNSMSO76_0),.clk(gclk));
	jdff dff_B_uz5JdEPA2_0(.din(n1557),.dout(w_dff_B_uz5JdEPA2_0),.clk(gclk));
	jdff dff_A_G5VoCGkp6_1(.dout(w_n1408_0[1]),.din(w_dff_A_G5VoCGkp6_1),.clk(gclk));
	jdff dff_A_J7u78SKN9_1(.dout(w_dff_A_G5VoCGkp6_1),.din(w_dff_A_J7u78SKN9_1),.clk(gclk));
	jdff dff_A_UyfMFkSm2_1(.dout(w_dff_A_J7u78SKN9_1),.din(w_dff_A_UyfMFkSm2_1),.clk(gclk));
	jdff dff_A_HgLKnW4C8_1(.dout(w_dff_A_UyfMFkSm2_1),.din(w_dff_A_HgLKnW4C8_1),.clk(gclk));
	jdff dff_A_oAA3E9by7_1(.dout(w_dff_A_HgLKnW4C8_1),.din(w_dff_A_oAA3E9by7_1),.clk(gclk));
	jdff dff_A_lfbYJuDe3_1(.dout(w_dff_A_oAA3E9by7_1),.din(w_dff_A_lfbYJuDe3_1),.clk(gclk));
	jdff dff_A_TKUk1gsn4_1(.dout(w_dff_A_lfbYJuDe3_1),.din(w_dff_A_TKUk1gsn4_1),.clk(gclk));
	jdff dff_B_8KIOEasC4_1(.din(n1403),.dout(w_dff_B_8KIOEasC4_1),.clk(gclk));
	jdff dff_B_waw4KLp83_1(.din(w_dff_B_8KIOEasC4_1),.dout(w_dff_B_waw4KLp83_1),.clk(gclk));
	jdff dff_B_hDLAAMvA5_1(.din(w_dff_B_waw4KLp83_1),.dout(w_dff_B_hDLAAMvA5_1),.clk(gclk));
	jdff dff_B_KVrrMNTG3_1(.din(w_dff_B_hDLAAMvA5_1),.dout(w_dff_B_KVrrMNTG3_1),.clk(gclk));
	jdff dff_B_in5wwlVu7_1(.din(w_dff_B_KVrrMNTG3_1),.dout(w_dff_B_in5wwlVu7_1),.clk(gclk));
	jdff dff_B_YuPztimZ1_1(.din(w_dff_B_in5wwlVu7_1),.dout(w_dff_B_YuPztimZ1_1),.clk(gclk));
	jdff dff_B_QRt6WBdp0_0(.din(n1405),.dout(w_dff_B_QRt6WBdp0_0),.clk(gclk));
	jdff dff_B_One0Agdz9_0(.din(w_dff_B_QRt6WBdp0_0),.dout(w_dff_B_One0Agdz9_0),.clk(gclk));
	jdff dff_B_cX7DX5Th0_0(.din(w_dff_B_One0Agdz9_0),.dout(w_dff_B_cX7DX5Th0_0),.clk(gclk));
	jdff dff_A_ecD2UVhc6_1(.dout(w_n1402_0[1]),.din(w_dff_A_ecD2UVhc6_1),.clk(gclk));
	jdff dff_A_cOHiFweG9_1(.dout(w_dff_A_ecD2UVhc6_1),.din(w_dff_A_cOHiFweG9_1),.clk(gclk));
	jdff dff_A_FekR1ssV9_1(.dout(w_dff_A_cOHiFweG9_1),.din(w_dff_A_FekR1ssV9_1),.clk(gclk));
	jdff dff_A_Q9SO47pB3_1(.dout(w_dff_A_FekR1ssV9_1),.din(w_dff_A_Q9SO47pB3_1),.clk(gclk));
	jdff dff_A_aIS6u4cB4_1(.dout(w_dff_A_Q9SO47pB3_1),.din(w_dff_A_aIS6u4cB4_1),.clk(gclk));
	jdff dff_A_OvrM5F6E5_1(.dout(w_dff_A_aIS6u4cB4_1),.din(w_dff_A_OvrM5F6E5_1),.clk(gclk));
	jdff dff_A_02qyTdDV4_1(.dout(w_dff_A_OvrM5F6E5_1),.din(w_dff_A_02qyTdDV4_1),.clk(gclk));
	jdff dff_A_EWnY6QVI2_1(.dout(w_dff_A_02qyTdDV4_1),.din(w_dff_A_EWnY6QVI2_1),.clk(gclk));
	jdff dff_A_Wi9IFu6e2_1(.dout(w_dff_A_EWnY6QVI2_1),.din(w_dff_A_Wi9IFu6e2_1),.clk(gclk));
	jdff dff_A_x9ng5r8N3_1(.dout(w_dff_A_Wi9IFu6e2_1),.din(w_dff_A_x9ng5r8N3_1),.clk(gclk));
	jdff dff_A_JTN3oEue1_1(.dout(w_dff_A_x9ng5r8N3_1),.din(w_dff_A_JTN3oEue1_1),.clk(gclk));
	jdff dff_A_rS5PolOt7_1(.dout(w_dff_A_JTN3oEue1_1),.din(w_dff_A_rS5PolOt7_1),.clk(gclk));
	jdff dff_A_agESjHom7_1(.dout(w_dff_A_rS5PolOt7_1),.din(w_dff_A_agESjHom7_1),.clk(gclk));
	jdff dff_A_Lbuzz2I51_1(.dout(w_dff_A_agESjHom7_1),.din(w_dff_A_Lbuzz2I51_1),.clk(gclk));
	jdff dff_A_GpqMXNZU8_1(.dout(w_dff_A_Lbuzz2I51_1),.din(w_dff_A_GpqMXNZU8_1),.clk(gclk));
	jdff dff_B_pTgNxzNA1_0(.din(n1549),.dout(w_dff_B_pTgNxzNA1_0),.clk(gclk));
	jdff dff_B_JwPkVB3w4_0(.din(n1548),.dout(w_dff_B_JwPkVB3w4_0),.clk(gclk));
	jdff dff_B_FYsF2bfK2_1(.din(n1311),.dout(w_dff_B_FYsF2bfK2_1),.clk(gclk));
	jdff dff_B_gCAW2DAF2_1(.din(w_dff_B_FYsF2bfK2_1),.dout(w_dff_B_gCAW2DAF2_1),.clk(gclk));
	jdff dff_B_CFxhFbna6_1(.din(w_dff_B_gCAW2DAF2_1),.dout(w_dff_B_CFxhFbna6_1),.clk(gclk));
	jdff dff_B_58RorVq24_1(.din(w_dff_B_CFxhFbna6_1),.dout(w_dff_B_58RorVq24_1),.clk(gclk));
	jdff dff_B_cIwl27WB0_1(.din(w_dff_B_58RorVq24_1),.dout(w_dff_B_cIwl27WB0_1),.clk(gclk));
	jdff dff_B_hLttKi5x0_1(.din(w_dff_B_cIwl27WB0_1),.dout(w_dff_B_hLttKi5x0_1),.clk(gclk));
	jdff dff_B_iO8JwX4U0_1(.din(w_dff_B_hLttKi5x0_1),.dout(w_dff_B_iO8JwX4U0_1),.clk(gclk));
	jdff dff_B_1kx18BGy0_1(.din(w_dff_B_iO8JwX4U0_1),.dout(w_dff_B_1kx18BGy0_1),.clk(gclk));
	jdff dff_B_odRQHQ3C6_1(.din(w_dff_B_1kx18BGy0_1),.dout(w_dff_B_odRQHQ3C6_1),.clk(gclk));
	jdff dff_B_LXOtIWEn4_1(.din(w_dff_B_odRQHQ3C6_1),.dout(w_dff_B_LXOtIWEn4_1),.clk(gclk));
	jdff dff_B_UiFwSTNy9_1(.din(w_dff_B_LXOtIWEn4_1),.dout(w_dff_B_UiFwSTNy9_1),.clk(gclk));
	jdff dff_B_nRC0Yr099_1(.din(w_dff_B_UiFwSTNy9_1),.dout(w_dff_B_nRC0Yr099_1),.clk(gclk));
	jdff dff_B_TmRP1p7q3_0(.din(n1545),.dout(w_dff_B_TmRP1p7q3_0),.clk(gclk));
	jdff dff_A_nIsRN38t6_1(.dout(w_n1543_0[1]),.din(w_dff_A_nIsRN38t6_1),.clk(gclk));
	jdff dff_B_d2XB5cjq2_2(.din(n1543),.dout(w_dff_B_d2XB5cjq2_2),.clk(gclk));
	jdff dff_B_B4ZEY8c77_2(.din(w_dff_B_d2XB5cjq2_2),.dout(w_dff_B_B4ZEY8c77_2),.clk(gclk));
	jdff dff_B_LTthsse71_0(.din(n1542),.dout(w_dff_B_LTthsse71_0),.clk(gclk));
	jdff dff_B_WdonE3CV6_0(.din(w_dff_B_LTthsse71_0),.dout(w_dff_B_WdonE3CV6_0),.clk(gclk));
	jdff dff_B_KphS10fo0_0(.din(w_dff_B_WdonE3CV6_0),.dout(w_dff_B_KphS10fo0_0),.clk(gclk));
	jdff dff_B_kAHKnmBg9_0(.din(w_dff_B_KphS10fo0_0),.dout(w_dff_B_kAHKnmBg9_0),.clk(gclk));
	jdff dff_B_jn8IgKiS4_0(.din(n1541),.dout(w_dff_B_jn8IgKiS4_0),.clk(gclk));
	jdff dff_B_Xh53Gc1B2_1(.din(n1538),.dout(w_dff_B_Xh53Gc1B2_1),.clk(gclk));
	jdff dff_B_4MLFFKzK1_1(.din(w_dff_B_Xh53Gc1B2_1),.dout(w_dff_B_4MLFFKzK1_1),.clk(gclk));
	jdff dff_B_vpfiJFkd0_1(.din(w_dff_B_4MLFFKzK1_1),.dout(w_dff_B_vpfiJFkd0_1),.clk(gclk));
	jdff dff_A_iAdNOIPv3_0(.dout(w_n1536_0[0]),.din(w_dff_A_iAdNOIPv3_0),.clk(gclk));
	jdff dff_A_JoU9a7Oq1_0(.dout(w_dff_A_iAdNOIPv3_0),.din(w_dff_A_JoU9a7Oq1_0),.clk(gclk));
	jdff dff_A_9uE2buWy8_0(.dout(w_dff_A_JoU9a7Oq1_0),.din(w_dff_A_9uE2buWy8_0),.clk(gclk));
	jdff dff_A_z6sf7Fkn6_0(.dout(w_dff_A_9uE2buWy8_0),.din(w_dff_A_z6sf7Fkn6_0),.clk(gclk));
	jdff dff_A_EAxVI1FH9_1(.dout(w_n1426_0[1]),.din(w_dff_A_EAxVI1FH9_1),.clk(gclk));
	jdff dff_A_eGotZmrQ3_1(.dout(w_dff_A_EAxVI1FH9_1),.din(w_dff_A_eGotZmrQ3_1),.clk(gclk));
	jdff dff_A_NNu9KYcg2_1(.dout(w_dff_A_eGotZmrQ3_1),.din(w_dff_A_NNu9KYcg2_1),.clk(gclk));
	jdff dff_A_D1LYb21k7_1(.dout(w_dff_A_NNu9KYcg2_1),.din(w_dff_A_D1LYb21k7_1),.clk(gclk));
	jdff dff_A_pSgudIjE3_1(.dout(w_dff_A_D1LYb21k7_1),.din(w_dff_A_pSgudIjE3_1),.clk(gclk));
	jdff dff_A_1wY814jb9_1(.dout(w_dff_A_pSgudIjE3_1),.din(w_dff_A_1wY814jb9_1),.clk(gclk));
	jdff dff_A_ZryUnmGD4_1(.dout(w_dff_A_1wY814jb9_1),.din(w_dff_A_ZryUnmGD4_1),.clk(gclk));
	jdff dff_A_36IVZN5a9_1(.dout(w_dff_A_ZryUnmGD4_1),.din(w_dff_A_36IVZN5a9_1),.clk(gclk));
	jdff dff_A_yPI8eKWu7_1(.dout(w_dff_A_36IVZN5a9_1),.din(w_dff_A_yPI8eKWu7_1),.clk(gclk));
	jdff dff_A_63KGx8rG5_1(.dout(w_dff_A_yPI8eKWu7_1),.din(w_dff_A_63KGx8rG5_1),.clk(gclk));
	jdff dff_A_8SRdCOxw0_1(.dout(w_dff_A_63KGx8rG5_1),.din(w_dff_A_8SRdCOxw0_1),.clk(gclk));
	jdff dff_A_q3UANLk35_1(.dout(w_dff_A_8SRdCOxw0_1),.din(w_dff_A_q3UANLk35_1),.clk(gclk));
	jdff dff_A_hEif0nC70_1(.dout(w_dff_A_q3UANLk35_1),.din(w_dff_A_hEif0nC70_1),.clk(gclk));
	jdff dff_A_AmjgDKJK9_1(.dout(w_dff_A_hEif0nC70_1),.din(w_dff_A_AmjgDKJK9_1),.clk(gclk));
	jdff dff_A_OLJlUU8w0_1(.dout(w_dff_A_AmjgDKJK9_1),.din(w_dff_A_OLJlUU8w0_1),.clk(gclk));
	jdff dff_A_ZZCWqlCV2_1(.dout(w_dff_A_OLJlUU8w0_1),.din(w_dff_A_ZZCWqlCV2_1),.clk(gclk));
	jdff dff_B_FCmJPHfS7_0(.din(n1533),.dout(w_dff_B_FCmJPHfS7_0),.clk(gclk));
	jdff dff_B_td1CobWD0_0(.din(w_dff_B_FCmJPHfS7_0),.dout(w_dff_B_td1CobWD0_0),.clk(gclk));
	jdff dff_B_x6SATIH07_0(.din(w_dff_B_td1CobWD0_0),.dout(w_dff_B_x6SATIH07_0),.clk(gclk));
	jdff dff_B_ryPHwt8F6_0(.din(w_dff_B_x6SATIH07_0),.dout(w_dff_B_ryPHwt8F6_0),.clk(gclk));
	jdff dff_B_d2U7s5oQ6_0(.din(n1532),.dout(w_dff_B_d2U7s5oQ6_0),.clk(gclk));
	jdff dff_B_oaIbomvf7_0(.din(w_dff_B_d2U7s5oQ6_0),.dout(w_dff_B_oaIbomvf7_0),.clk(gclk));
	jdff dff_B_aaz4RO4F3_0(.din(w_dff_B_oaIbomvf7_0),.dout(w_dff_B_aaz4RO4F3_0),.clk(gclk));
	jdff dff_A_Wi6E2LJo4_1(.dout(w_n1419_0[1]),.din(w_dff_A_Wi6E2LJo4_1),.clk(gclk));
	jdff dff_A_9nftVOMq4_1(.dout(w_dff_A_Wi6E2LJo4_1),.din(w_dff_A_9nftVOMq4_1),.clk(gclk));
	jdff dff_A_cyHA4Zav3_1(.dout(w_dff_A_9nftVOMq4_1),.din(w_dff_A_cyHA4Zav3_1),.clk(gclk));
	jdff dff_A_Qg8qfCDN1_1(.dout(w_dff_A_cyHA4Zav3_1),.din(w_dff_A_Qg8qfCDN1_1),.clk(gclk));
	jdff dff_A_pLDhhI3T2_1(.dout(w_dff_A_Qg8qfCDN1_1),.din(w_dff_A_pLDhhI3T2_1),.clk(gclk));
	jdff dff_A_g2n6lwlj0_1(.dout(w_dff_A_pLDhhI3T2_1),.din(w_dff_A_g2n6lwlj0_1),.clk(gclk));
	jdff dff_A_fPjZS4nm8_1(.dout(w_dff_A_g2n6lwlj0_1),.din(w_dff_A_fPjZS4nm8_1),.clk(gclk));
	jdff dff_A_3utLmtf54_1(.dout(w_dff_A_fPjZS4nm8_1),.din(w_dff_A_3utLmtf54_1),.clk(gclk));
	jdff dff_A_WPovrqbZ6_1(.dout(w_dff_A_3utLmtf54_1),.din(w_dff_A_WPovrqbZ6_1),.clk(gclk));
	jdff dff_A_5CgJH34Z8_1(.dout(w_dff_A_WPovrqbZ6_1),.din(w_dff_A_5CgJH34Z8_1),.clk(gclk));
	jdff dff_A_px9vcTcr0_1(.dout(w_dff_A_5CgJH34Z8_1),.din(w_dff_A_px9vcTcr0_1),.clk(gclk));
	jdff dff_A_OEHqpfUh9_1(.dout(w_dff_A_px9vcTcr0_1),.din(w_dff_A_OEHqpfUh9_1),.clk(gclk));
	jdff dff_A_v1SmNGQr8_1(.dout(w_dff_A_OEHqpfUh9_1),.din(w_dff_A_v1SmNGQr8_1),.clk(gclk));
	jdff dff_A_IgszziJX7_1(.dout(w_dff_A_v1SmNGQr8_1),.din(w_dff_A_IgszziJX7_1),.clk(gclk));
	jdff dff_A_3vVToo9h8_1(.dout(w_dff_A_IgszziJX7_1),.din(w_dff_A_3vVToo9h8_1),.clk(gclk));
	jdff dff_A_67SlbUFS4_1(.dout(w_dff_A_3vVToo9h8_1),.din(w_dff_A_67SlbUFS4_1),.clk(gclk));
	jdff dff_A_GSGGZwE50_1(.dout(w_dff_A_67SlbUFS4_1),.din(w_dff_A_GSGGZwE50_1),.clk(gclk));
	jdff dff_A_mN7i3Yrl0_1(.dout(w_dff_A_GSGGZwE50_1),.din(w_dff_A_mN7i3Yrl0_1),.clk(gclk));
	jdff dff_A_DFF7w8UG3_1(.dout(w_dff_A_mN7i3Yrl0_1),.din(w_dff_A_DFF7w8UG3_1),.clk(gclk));
	jdff dff_A_9ELLg1NZ1_1(.dout(w_dff_A_DFF7w8UG3_1),.din(w_dff_A_9ELLg1NZ1_1),.clk(gclk));
	jdff dff_B_XYDuZhvK7_2(.din(n1419),.dout(w_dff_B_XYDuZhvK7_2),.clk(gclk));
	jdff dff_A_9g2qfnBI4_2(.dout(w_n504_0[2]),.din(w_dff_A_9g2qfnBI4_2),.clk(gclk));
	jdff dff_B_OjPSi83b8_1(.din(n502),.dout(w_dff_B_OjPSi83b8_1),.clk(gclk));
	jdff dff_B_hevlZQKt0_0(.din(G66),.dout(w_dff_B_hevlZQKt0_0),.clk(gclk));
	jdff dff_A_AZjeSlZO9_0(.dout(w_n501_0[0]),.din(w_dff_A_AZjeSlZO9_0),.clk(gclk));
	jdff dff_A_jggx32xI4_0(.dout(w_dff_A_AZjeSlZO9_0),.din(w_dff_A_jggx32xI4_0),.clk(gclk));
	jdff dff_A_Tuk0jMnd9_2(.dout(w_n501_0[2]),.din(w_dff_A_Tuk0jMnd9_2),.clk(gclk));
	jdff dff_A_2cU5pr8u4_2(.dout(w_dff_A_Tuk0jMnd9_2),.din(w_dff_A_2cU5pr8u4_2),.clk(gclk));
	jdff dff_A_7yLK3So26_1(.dout(w_G4437_0[1]),.din(w_dff_A_7yLK3So26_1),.clk(gclk));
	jdff dff_A_akYgauwP8_1(.dout(w_dff_A_7yLK3So26_1),.din(w_dff_A_akYgauwP8_1),.clk(gclk));
	jdff dff_A_1s9AXgTT6_1(.dout(w_dff_A_akYgauwP8_1),.din(w_dff_A_1s9AXgTT6_1),.clk(gclk));
	jdff dff_A_4CLa4k1Y8_1(.dout(w_dff_A_1s9AXgTT6_1),.din(w_dff_A_4CLa4k1Y8_1),.clk(gclk));
	jdff dff_A_0KLLPL4s9_1(.dout(w_n1308_0[1]),.din(w_dff_A_0KLLPL4s9_1),.clk(gclk));
	jdff dff_A_pvdZHmJR1_1(.dout(w_dff_A_0KLLPL4s9_1),.din(w_dff_A_pvdZHmJR1_1),.clk(gclk));
	jdff dff_A_8YpAQu4S6_1(.dout(w_dff_A_pvdZHmJR1_1),.din(w_dff_A_8YpAQu4S6_1),.clk(gclk));
	jdff dff_A_S3pMlIGa0_1(.dout(w_dff_A_8YpAQu4S6_1),.din(w_dff_A_S3pMlIGa0_1),.clk(gclk));
	jdff dff_A_EXrf9peh3_1(.dout(w_dff_A_S3pMlIGa0_1),.din(w_dff_A_EXrf9peh3_1),.clk(gclk));
	jdff dff_A_NILS2dXM9_1(.dout(w_dff_A_EXrf9peh3_1),.din(w_dff_A_NILS2dXM9_1),.clk(gclk));
	jdff dff_A_rMlBMTFf2_1(.dout(w_dff_A_NILS2dXM9_1),.din(w_dff_A_rMlBMTFf2_1),.clk(gclk));
	jdff dff_A_NCqt1J6M7_1(.dout(w_dff_A_rMlBMTFf2_1),.din(w_dff_A_NCqt1J6M7_1),.clk(gclk));
	jdff dff_A_7c2tpUQI9_1(.dout(w_dff_A_NCqt1J6M7_1),.din(w_dff_A_7c2tpUQI9_1),.clk(gclk));
	jdff dff_A_p8haoUJq4_1(.dout(w_dff_A_7c2tpUQI9_1),.din(w_dff_A_p8haoUJq4_1),.clk(gclk));
	jdff dff_A_lmL2Uuze4_1(.dout(w_dff_A_p8haoUJq4_1),.din(w_dff_A_lmL2Uuze4_1),.clk(gclk));
	jdff dff_A_PDstxXkQ3_1(.dout(w_dff_A_lmL2Uuze4_1),.din(w_dff_A_PDstxXkQ3_1),.clk(gclk));
	jdff dff_A_gUul2mw15_1(.dout(w_dff_A_PDstxXkQ3_1),.din(w_dff_A_gUul2mw15_1),.clk(gclk));
	jdff dff_A_voPurD9a3_1(.dout(w_dff_A_gUul2mw15_1),.din(w_dff_A_voPurD9a3_1),.clk(gclk));
	jdff dff_A_Rdj7FWHn1_1(.dout(w_dff_A_voPurD9a3_1),.din(w_dff_A_Rdj7FWHn1_1),.clk(gclk));
	jdff dff_A_zlS3VSDO0_1(.dout(w_dff_A_Rdj7FWHn1_1),.din(w_dff_A_zlS3VSDO0_1),.clk(gclk));
	jdff dff_A_powAz74V9_0(.dout(w_n526_0[0]),.din(w_dff_A_powAz74V9_0),.clk(gclk));
	jdff dff_A_PbcLaPLQ3_1(.dout(w_n526_0[1]),.din(w_dff_A_PbcLaPLQ3_1),.clk(gclk));
	jdff dff_A_RExE2HPu3_1(.dout(w_dff_A_PbcLaPLQ3_1),.din(w_dff_A_RExE2HPu3_1),.clk(gclk));
	jdff dff_A_prtf9rx73_1(.dout(w_dff_A_RExE2HPu3_1),.din(w_dff_A_prtf9rx73_1),.clk(gclk));
	jdff dff_A_YMpjr2zA1_1(.dout(w_dff_A_prtf9rx73_1),.din(w_dff_A_YMpjr2zA1_1),.clk(gclk));
	jdff dff_A_pytR5S3c5_1(.dout(w_dff_A_YMpjr2zA1_1),.din(w_dff_A_pytR5S3c5_1),.clk(gclk));
	jdff dff_A_gj1an2Kd8_1(.dout(w_dff_A_pytR5S3c5_1),.din(w_dff_A_gj1an2Kd8_1),.clk(gclk));
	jdff dff_A_NDBWt4Gi7_1(.dout(w_dff_A_gj1an2Kd8_1),.din(w_dff_A_NDBWt4Gi7_1),.clk(gclk));
	jdff dff_A_x0vXnbmk4_1(.dout(w_dff_A_NDBWt4Gi7_1),.din(w_dff_A_x0vXnbmk4_1),.clk(gclk));
	jdff dff_A_gjE7Cwl60_1(.dout(w_dff_A_x0vXnbmk4_1),.din(w_dff_A_gjE7Cwl60_1),.clk(gclk));
	jdff dff_A_EWvrhSlB1_1(.dout(w_dff_A_gjE7Cwl60_1),.din(w_dff_A_EWvrhSlB1_1),.clk(gclk));
	jdff dff_A_d3yFPxrF5_1(.dout(w_dff_A_EWvrhSlB1_1),.din(w_dff_A_d3yFPxrF5_1),.clk(gclk));
	jdff dff_A_gk5TTWpK9_1(.dout(w_dff_A_d3yFPxrF5_1),.din(w_dff_A_gk5TTWpK9_1),.clk(gclk));
	jdff dff_A_alYCBDb98_1(.dout(w_dff_A_gk5TTWpK9_1),.din(w_dff_A_alYCBDb98_1),.clk(gclk));
	jdff dff_A_zcKipE6K2_1(.dout(w_dff_A_alYCBDb98_1),.din(w_dff_A_zcKipE6K2_1),.clk(gclk));
	jdff dff_A_6ToQmENd2_1(.dout(w_dff_A_zcKipE6K2_1),.din(w_dff_A_6ToQmENd2_1),.clk(gclk));
	jdff dff_B_mkdFzHJL4_0(.din(n1528),.dout(w_dff_B_mkdFzHJL4_0),.clk(gclk));
	jdff dff_A_xgd73YNd1_0(.dout(w_n687_0[0]),.din(w_dff_A_xgd73YNd1_0),.clk(gclk));
	jdff dff_A_EwimlYRb6_0(.dout(w_dff_A_xgd73YNd1_0),.din(w_dff_A_EwimlYRb6_0),.clk(gclk));
	jdff dff_A_IojLoow58_0(.dout(w_n694_0[0]),.din(w_dff_A_IojLoow58_0),.clk(gclk));
	jdff dff_A_KWRn9VrQ3_0(.dout(w_dff_A_IojLoow58_0),.din(w_dff_A_KWRn9VrQ3_0),.clk(gclk));
	jdff dff_A_Bg8ECj7Q6_0(.dout(w_dff_A_KWRn9VrQ3_0),.din(w_dff_A_Bg8ECj7Q6_0),.clk(gclk));
	jdff dff_A_J61Cz9ao4_0(.dout(w_dff_A_Bg8ECj7Q6_0),.din(w_dff_A_J61Cz9ao4_0),.clk(gclk));
	jdff dff_A_pDZnYLP57_0(.dout(w_dff_A_J61Cz9ao4_0),.din(w_dff_A_pDZnYLP57_0),.clk(gclk));
	jdff dff_A_QjDMdVsT3_0(.dout(w_dff_A_pDZnYLP57_0),.din(w_dff_A_QjDMdVsT3_0),.clk(gclk));
	jdff dff_A_MqXFakvJ1_0(.dout(w_dff_A_QjDMdVsT3_0),.din(w_dff_A_MqXFakvJ1_0),.clk(gclk));
	jdff dff_A_9JHRMoDA2_0(.dout(w_dff_A_MqXFakvJ1_0),.din(w_dff_A_9JHRMoDA2_0),.clk(gclk));
	jdff dff_A_SybwssI75_0(.dout(w_dff_A_9JHRMoDA2_0),.din(w_dff_A_SybwssI75_0),.clk(gclk));
	jdff dff_A_8KsBEpC97_0(.dout(w_dff_A_SybwssI75_0),.din(w_dff_A_8KsBEpC97_0),.clk(gclk));
	jdff dff_A_bPfJXG0X2_0(.dout(w_dff_A_8KsBEpC97_0),.din(w_dff_A_bPfJXG0X2_0),.clk(gclk));
	jdff dff_A_euClOofw5_0(.dout(w_dff_A_bPfJXG0X2_0),.din(w_dff_A_euClOofw5_0),.clk(gclk));
	jdff dff_A_xOFp0yv78_0(.dout(w_dff_A_euClOofw5_0),.din(w_dff_A_xOFp0yv78_0),.clk(gclk));
	jdff dff_A_35YdLmI60_0(.dout(w_dff_A_xOFp0yv78_0),.din(w_dff_A_35YdLmI60_0),.clk(gclk));
	jdff dff_A_s4tbPafp6_0(.dout(w_dff_A_35YdLmI60_0),.din(w_dff_A_s4tbPafp6_0),.clk(gclk));
	jdff dff_A_q5tRPNSs9_0(.dout(w_dff_A_s4tbPafp6_0),.din(w_dff_A_q5tRPNSs9_0),.clk(gclk));
	jdff dff_B_zif2k5jg5_1(.din(n691),.dout(w_dff_B_zif2k5jg5_1),.clk(gclk));
	jdff dff_A_Dj3DA7wv9_2(.dout(w_n524_1[2]),.din(w_dff_A_Dj3DA7wv9_2),.clk(gclk));
	jdff dff_A_7Tau7gTA6_2(.dout(w_dff_A_Dj3DA7wv9_2),.din(w_dff_A_7Tau7gTA6_2),.clk(gclk));
	jdff dff_A_gicobGyc3_2(.dout(w_dff_A_7Tau7gTA6_2),.din(w_dff_A_gicobGyc3_2),.clk(gclk));
	jdff dff_A_w1ybD9kK7_2(.dout(w_dff_A_gicobGyc3_2),.din(w_dff_A_w1ybD9kK7_2),.clk(gclk));
	jdff dff_A_ds8IdZiz7_2(.dout(w_dff_A_w1ybD9kK7_2),.din(w_dff_A_ds8IdZiz7_2),.clk(gclk));
	jdff dff_A_0cnjByHZ7_2(.dout(w_dff_A_ds8IdZiz7_2),.din(w_dff_A_0cnjByHZ7_2),.clk(gclk));
	jdff dff_A_zOr7Kzy26_2(.dout(w_dff_A_0cnjByHZ7_2),.din(w_dff_A_zOr7Kzy26_2),.clk(gclk));
	jdff dff_A_rZ8T6MVo3_2(.dout(w_dff_A_zOr7Kzy26_2),.din(w_dff_A_rZ8T6MVo3_2),.clk(gclk));
	jdff dff_A_fwufgFKK9_2(.dout(w_dff_A_rZ8T6MVo3_2),.din(w_dff_A_fwufgFKK9_2),.clk(gclk));
	jdff dff_A_8eEiDzOi0_2(.dout(w_dff_A_fwufgFKK9_2),.din(w_dff_A_8eEiDzOi0_2),.clk(gclk));
	jdff dff_A_eveQR6kS6_2(.dout(w_dff_A_8eEiDzOi0_2),.din(w_dff_A_eveQR6kS6_2),.clk(gclk));
	jdff dff_A_q3PuDnq04_2(.dout(w_dff_A_eveQR6kS6_2),.din(w_dff_A_q3PuDnq04_2),.clk(gclk));
	jdff dff_A_u52IRCK89_2(.dout(w_dff_A_q3PuDnq04_2),.din(w_dff_A_u52IRCK89_2),.clk(gclk));
	jdff dff_A_9eJ9HbSg4_2(.dout(w_dff_A_u52IRCK89_2),.din(w_dff_A_9eJ9HbSg4_2),.clk(gclk));
	jdff dff_A_vSC06nqv4_2(.dout(w_dff_A_9eJ9HbSg4_2),.din(w_dff_A_vSC06nqv4_2),.clk(gclk));
	jdff dff_A_hafLcM778_2(.dout(w_dff_A_vSC06nqv4_2),.din(w_dff_A_hafLcM778_2),.clk(gclk));
	jdff dff_A_E8kYfVRo1_2(.dout(w_dff_A_hafLcM778_2),.din(w_dff_A_E8kYfVRo1_2),.clk(gclk));
	jdff dff_A_ijuTNTL78_0(.dout(w_n518_1[0]),.din(w_dff_A_ijuTNTL78_0),.clk(gclk));
	jdff dff_A_6Z1d3v7H1_0(.dout(w_dff_A_ijuTNTL78_0),.din(w_dff_A_6Z1d3v7H1_0),.clk(gclk));
	jdff dff_A_BXjGEBES7_0(.dout(w_dff_A_6Z1d3v7H1_0),.din(w_dff_A_BXjGEBES7_0),.clk(gclk));
	jdff dff_A_fdpv6NKn2_0(.dout(w_dff_A_BXjGEBES7_0),.din(w_dff_A_fdpv6NKn2_0),.clk(gclk));
	jdff dff_A_HRaddUvR5_0(.dout(w_dff_A_fdpv6NKn2_0),.din(w_dff_A_HRaddUvR5_0),.clk(gclk));
	jdff dff_A_sENznjUR7_0(.dout(w_dff_A_HRaddUvR5_0),.din(w_dff_A_sENznjUR7_0),.clk(gclk));
	jdff dff_A_6ITc35Vn3_0(.dout(w_dff_A_sENznjUR7_0),.din(w_dff_A_6ITc35Vn3_0),.clk(gclk));
	jdff dff_A_jvKDct7U9_0(.dout(w_dff_A_6ITc35Vn3_0),.din(w_dff_A_jvKDct7U9_0),.clk(gclk));
	jdff dff_A_66c7i4qM5_0(.dout(w_dff_A_jvKDct7U9_0),.din(w_dff_A_66c7i4qM5_0),.clk(gclk));
	jdff dff_A_P7wMnUqo9_0(.dout(w_dff_A_66c7i4qM5_0),.din(w_dff_A_P7wMnUqo9_0),.clk(gclk));
	jdff dff_A_JbXlZfCK4_0(.dout(w_dff_A_P7wMnUqo9_0),.din(w_dff_A_JbXlZfCK4_0),.clk(gclk));
	jdff dff_A_RLwTPzdA1_0(.dout(w_dff_A_JbXlZfCK4_0),.din(w_dff_A_RLwTPzdA1_0),.clk(gclk));
	jdff dff_A_BouNLdYb9_0(.dout(w_dff_A_RLwTPzdA1_0),.din(w_dff_A_BouNLdYb9_0),.clk(gclk));
	jdff dff_A_9M46Ac4o7_0(.dout(w_dff_A_BouNLdYb9_0),.din(w_dff_A_9M46Ac4o7_0),.clk(gclk));
	jdff dff_A_B8cVVLXC0_0(.dout(w_dff_A_9M46Ac4o7_0),.din(w_dff_A_B8cVVLXC0_0),.clk(gclk));
	jdff dff_A_rITaSCkS6_0(.dout(w_dff_A_B8cVVLXC0_0),.din(w_dff_A_rITaSCkS6_0),.clk(gclk));
	jdff dff_A_ndPhYgKa6_0(.dout(w_dff_A_rITaSCkS6_0),.din(w_dff_A_ndPhYgKa6_0),.clk(gclk));
	jdff dff_A_5oso5I1j9_0(.dout(w_dff_A_ndPhYgKa6_0),.din(w_dff_A_5oso5I1j9_0),.clk(gclk));
	jdff dff_B_kgtB5zK48_1(.din(n515),.dout(w_dff_B_kgtB5zK48_1),.clk(gclk));
	jdff dff_B_6Hnef3P70_0(.din(G35),.dout(w_dff_B_6Hnef3P70_0),.clk(gclk));
	jdff dff_B_qEqpUElT1_2(.din(n514),.dout(w_dff_B_qEqpUElT1_2),.clk(gclk));
	jdff dff_B_V2dp9oao7_2(.din(w_dff_B_qEqpUElT1_2),.dout(w_dff_B_V2dp9oao7_2),.clk(gclk));
	jdff dff_A_O38cRWwB9_0(.dout(w_G4420_1[0]),.din(w_dff_A_O38cRWwB9_0),.clk(gclk));
	jdff dff_A_bqzeMAZm9_0(.dout(w_dff_A_O38cRWwB9_0),.din(w_dff_A_bqzeMAZm9_0),.clk(gclk));
	jdff dff_A_b5cgMnwu5_0(.dout(w_dff_A_bqzeMAZm9_0),.din(w_dff_A_b5cgMnwu5_0),.clk(gclk));
	jdff dff_A_HBJIOJCi0_0(.dout(w_dff_A_b5cgMnwu5_0),.din(w_dff_A_HBJIOJCi0_0),.clk(gclk));
	jdff dff_B_1uxc9meZ2_1(.din(n521),.dout(w_dff_B_1uxc9meZ2_1),.clk(gclk));
	jdff dff_B_FI8IhTCi2_0(.din(G32),.dout(w_dff_B_FI8IhTCi2_0),.clk(gclk));
	jdff dff_B_Ku9p1LZk8_2(.din(n520),.dout(w_dff_B_Ku9p1LZk8_2),.clk(gclk));
	jdff dff_B_9w2r0qCf1_2(.din(w_dff_B_Ku9p1LZk8_2),.dout(w_dff_B_9w2r0qCf1_2),.clk(gclk));
	jdff dff_A_cBpxTyuL7_1(.dout(w_n690_0[1]),.din(w_dff_A_cBpxTyuL7_1),.clk(gclk));
	jdff dff_B_stDaMQtR2_2(.din(n690),.dout(w_dff_B_stDaMQtR2_2),.clk(gclk));
	jdff dff_A_JOmmXEPd3_2(.dout(w_n513_0[2]),.din(w_dff_A_JOmmXEPd3_2),.clk(gclk));
	jdff dff_A_lvSU19PP7_2(.dout(w_dff_A_JOmmXEPd3_2),.din(w_dff_A_lvSU19PP7_2),.clk(gclk));
	jdff dff_A_Z9nIQoCp2_2(.dout(w_dff_A_lvSU19PP7_2),.din(w_dff_A_Z9nIQoCp2_2),.clk(gclk));
	jdff dff_A_H8YYUOsO4_2(.dout(w_dff_A_Z9nIQoCp2_2),.din(w_dff_A_H8YYUOsO4_2),.clk(gclk));
	jdff dff_A_mEQNs6C42_2(.dout(w_dff_A_H8YYUOsO4_2),.din(w_dff_A_mEQNs6C42_2),.clk(gclk));
	jdff dff_B_eprve7413_1(.din(n510),.dout(w_dff_B_eprve7413_1),.clk(gclk));
	jdff dff_B_kh9eKsd88_0(.din(G50),.dout(w_dff_B_kh9eKsd88_0),.clk(gclk));
	jdff dff_A_5S4Af8175_1(.dout(w_n509_0[1]),.din(w_dff_A_5S4Af8175_1),.clk(gclk));
	jdff dff_A_iDCFiOTb3_1(.dout(w_dff_A_5S4Af8175_1),.din(w_dff_A_iDCFiOTb3_1),.clk(gclk));
	jdff dff_A_KCLPAnYJ7_2(.dout(w_n509_0[2]),.din(w_dff_A_KCLPAnYJ7_2),.clk(gclk));
	jdff dff_A_eBZdL6T88_2(.dout(w_dff_A_KCLPAnYJ7_2),.din(w_dff_A_eBZdL6T88_2),.clk(gclk));
	jdff dff_A_nRpXKqVf5_1(.dout(w_G4432_0[1]),.din(w_dff_A_nRpXKqVf5_1),.clk(gclk));
	jdff dff_A_etaTxasj8_1(.dout(w_dff_A_nRpXKqVf5_1),.din(w_dff_A_etaTxasj8_1),.clk(gclk));
	jdff dff_A_6hNQKIf72_1(.dout(w_dff_A_etaTxasj8_1),.din(w_dff_A_6hNQKIf72_1),.clk(gclk));
	jdff dff_A_7nXfocmh8_1(.dout(w_dff_A_6hNQKIf72_1),.din(w_dff_A_7nXfocmh8_1),.clk(gclk));
	jdff dff_A_tTzWUmWD5_1(.dout(w_n1309_0[1]),.din(w_dff_A_tTzWUmWD5_1),.clk(gclk));
	jdff dff_A_JQtcVcW30_1(.dout(w_dff_A_tTzWUmWD5_1),.din(w_dff_A_JQtcVcW30_1),.clk(gclk));
	jdff dff_A_GUwOCB6M5_1(.dout(w_dff_A_JQtcVcW30_1),.din(w_dff_A_GUwOCB6M5_1),.clk(gclk));
	jdff dff_A_HnVWsxJd4_1(.dout(w_dff_A_GUwOCB6M5_1),.din(w_dff_A_HnVWsxJd4_1),.clk(gclk));
	jdff dff_A_ckG5mk5n5_1(.dout(w_n572_1[1]),.din(w_dff_A_ckG5mk5n5_1),.clk(gclk));
	jdff dff_A_cBVGppdq7_1(.dout(w_dff_A_ckG5mk5n5_1),.din(w_dff_A_cBVGppdq7_1),.clk(gclk));
	jdff dff_A_b5O9x9WL1_1(.dout(w_dff_A_cBVGppdq7_1),.din(w_dff_A_b5O9x9WL1_1),.clk(gclk));
	jdff dff_A_ChrPDoUt9_1(.dout(w_dff_A_b5O9x9WL1_1),.din(w_dff_A_ChrPDoUt9_1),.clk(gclk));
	jdff dff_A_kxNOyO7N4_1(.dout(w_dff_A_ChrPDoUt9_1),.din(w_dff_A_kxNOyO7N4_1),.clk(gclk));
	jdff dff_B_Ik4vbIEX3_1(.din(n532),.dout(w_dff_B_Ik4vbIEX3_1),.clk(gclk));
	jdff dff_B_QQ6alOl00_1(.din(w_dff_B_Ik4vbIEX3_1),.dout(w_dff_B_QQ6alOl00_1),.clk(gclk));
	jdff dff_B_X2FDpMm36_1(.din(w_dff_B_QQ6alOl00_1),.dout(w_dff_B_X2FDpMm36_1),.clk(gclk));
	jdff dff_B_MHByK6Eq9_1(.din(w_dff_B_X2FDpMm36_1),.dout(w_dff_B_MHByK6Eq9_1),.clk(gclk));
	jdff dff_B_iYETiQbB5_1(.din(w_dff_B_MHByK6Eq9_1),.dout(w_dff_B_iYETiQbB5_1),.clk(gclk));
	jdff dff_B_Venm6auk9_1(.din(w_dff_B_iYETiQbB5_1),.dout(w_dff_B_Venm6auk9_1),.clk(gclk));
	jdff dff_B_qb6YZBQ74_1(.din(w_dff_B_Venm6auk9_1),.dout(w_dff_B_qb6YZBQ74_1),.clk(gclk));
	jdff dff_B_NzvuBmVy4_1(.din(w_dff_B_qb6YZBQ74_1),.dout(w_dff_B_NzvuBmVy4_1),.clk(gclk));
	jdff dff_B_BEuDBo4u4_1(.din(w_dff_B_NzvuBmVy4_1),.dout(w_dff_B_BEuDBo4u4_1),.clk(gclk));
	jdff dff_B_0kqVoX2y3_1(.din(n535),.dout(w_dff_B_0kqVoX2y3_1),.clk(gclk));
	jdff dff_B_vNMvTpCU8_1(.din(w_dff_B_0kqVoX2y3_1),.dout(w_dff_B_vNMvTpCU8_1),.clk(gclk));
	jdff dff_B_Nlt59Phy8_1(.din(w_dff_B_vNMvTpCU8_1),.dout(w_dff_B_Nlt59Phy8_1),.clk(gclk));
	jdff dff_B_RyXZpfk67_1(.din(w_dff_B_Nlt59Phy8_1),.dout(w_dff_B_RyXZpfk67_1),.clk(gclk));
	jdff dff_B_4PI7nKJX5_1(.din(w_dff_B_RyXZpfk67_1),.dout(w_dff_B_4PI7nKJX5_1),.clk(gclk));
	jdff dff_B_DkdIHtIg6_1(.din(w_dff_B_4PI7nKJX5_1),.dout(w_dff_B_DkdIHtIg6_1),.clk(gclk));
	jdff dff_A_PMlK8EoZ3_1(.dout(w_n570_1[1]),.din(w_dff_A_PMlK8EoZ3_1),.clk(gclk));
	jdff dff_A_NNm5HebY3_1(.dout(w_dff_A_PMlK8EoZ3_1),.din(w_dff_A_NNm5HebY3_1),.clk(gclk));
	jdff dff_A_vFPzkZcD1_1(.dout(w_dff_A_NNm5HebY3_1),.din(w_dff_A_vFPzkZcD1_1),.clk(gclk));
	jdff dff_A_IRf6ExwL3_1(.dout(w_dff_A_vFPzkZcD1_1),.din(w_dff_A_IRf6ExwL3_1),.clk(gclk));
	jdff dff_A_rNK7SLuU1_1(.dout(w_dff_A_IRf6ExwL3_1),.din(w_dff_A_rNK7SLuU1_1),.clk(gclk));
	jdff dff_A_CE8TZrZ11_1(.dout(w_dff_A_rNK7SLuU1_1),.din(w_dff_A_CE8TZrZ11_1),.clk(gclk));
	jdff dff_A_vtLg4Pz35_1(.dout(w_dff_A_CE8TZrZ11_1),.din(w_dff_A_vtLg4Pz35_1),.clk(gclk));
	jdff dff_B_YrCqxNbT4_1(.din(n540),.dout(w_dff_B_YrCqxNbT4_1),.clk(gclk));
	jdff dff_B_SB8hL7Ki5_1(.din(w_dff_B_YrCqxNbT4_1),.dout(w_dff_B_SB8hL7Ki5_1),.clk(gclk));
	jdff dff_B_gUpevgBD3_1(.din(w_dff_B_SB8hL7Ki5_1),.dout(w_dff_B_gUpevgBD3_1),.clk(gclk));
	jdff dff_B_HE2ZpfZg5_1(.din(w_dff_B_gUpevgBD3_1),.dout(w_dff_B_HE2ZpfZg5_1),.clk(gclk));
	jdff dff_B_UcisGcxM6_1(.din(w_dff_B_HE2ZpfZg5_1),.dout(w_dff_B_UcisGcxM6_1),.clk(gclk));
	jdff dff_B_N4pNtpjI3_1(.din(w_dff_B_UcisGcxM6_1),.dout(w_dff_B_N4pNtpjI3_1),.clk(gclk));
	jdff dff_B_iu005BEr3_1(.din(w_dff_B_N4pNtpjI3_1),.dout(w_dff_B_iu005BEr3_1),.clk(gclk));
	jdff dff_B_RA7GSw6j4_1(.din(n543),.dout(w_dff_B_RA7GSw6j4_1),.clk(gclk));
	jdff dff_B_gopcol739_1(.din(w_dff_B_RA7GSw6j4_1),.dout(w_dff_B_gopcol739_1),.clk(gclk));
	jdff dff_B_wxZYj8iP6_1(.din(w_dff_B_gopcol739_1),.dout(w_dff_B_wxZYj8iP6_1),.clk(gclk));
	jdff dff_B_FeOV8fMy1_1(.din(w_dff_B_wxZYj8iP6_1),.dout(w_dff_B_FeOV8fMy1_1),.clk(gclk));
	jdff dff_B_QAni6bGw5_1(.din(n551),.dout(w_dff_B_QAni6bGw5_1),.clk(gclk));
	jdff dff_B_M54LwU609_1(.din(w_dff_B_QAni6bGw5_1),.dout(w_dff_B_M54LwU609_1),.clk(gclk));
	jdff dff_A_vJugByyt6_0(.dout(w_n566_0[0]),.din(w_dff_A_vJugByyt6_0),.clk(gclk));
	jdff dff_A_BaT3VEvH7_0(.dout(w_dff_A_vJugByyt6_0),.din(w_dff_A_BaT3VEvH7_0),.clk(gclk));
	jdff dff_A_0ZUkzLIF1_0(.dout(w_dff_A_BaT3VEvH7_0),.din(w_dff_A_0ZUkzLIF1_0),.clk(gclk));
	jdff dff_A_blumDytY3_0(.dout(w_dff_A_0ZUkzLIF1_0),.din(w_dff_A_blumDytY3_0),.clk(gclk));
	jdff dff_A_Kd3z0hum8_0(.dout(w_dff_A_blumDytY3_0),.din(w_dff_A_Kd3z0hum8_0),.clk(gclk));
	jdff dff_A_V6ue6u8k0_0(.dout(w_dff_A_Kd3z0hum8_0),.din(w_dff_A_V6ue6u8k0_0),.clk(gclk));
	jdff dff_A_ebunmQqZ3_0(.dout(w_dff_A_V6ue6u8k0_0),.din(w_dff_A_ebunmQqZ3_0),.clk(gclk));
	jdff dff_A_LjYP9uA77_0(.dout(w_dff_A_ebunmQqZ3_0),.din(w_dff_A_LjYP9uA77_0),.clk(gclk));
	jdff dff_A_SzYy73Gq8_0(.dout(w_dff_A_LjYP9uA77_0),.din(w_dff_A_SzYy73Gq8_0),.clk(gclk));
	jdff dff_A_vXJCbXxc0_0(.dout(w_dff_A_SzYy73Gq8_0),.din(w_dff_A_vXJCbXxc0_0),.clk(gclk));
	jdff dff_A_SFSrMxs73_0(.dout(w_dff_A_vXJCbXxc0_0),.din(w_dff_A_SFSrMxs73_0),.clk(gclk));
	jdff dff_A_N94m8ke02_1(.dout(w_n564_0[1]),.din(w_dff_A_N94m8ke02_1),.clk(gclk));
	jdff dff_A_8SPwT7SL5_1(.dout(w_dff_A_N94m8ke02_1),.din(w_dff_A_8SPwT7SL5_1),.clk(gclk));
	jdff dff_A_AlL3C5b40_1(.dout(w_dff_A_8SPwT7SL5_1),.din(w_dff_A_AlL3C5b40_1),.clk(gclk));
	jdff dff_A_G5mp3rok0_1(.dout(w_dff_A_AlL3C5b40_1),.din(w_dff_A_G5mp3rok0_1),.clk(gclk));
	jdff dff_A_DxZAQzaO9_1(.dout(w_dff_A_G5mp3rok0_1),.din(w_dff_A_DxZAQzaO9_1),.clk(gclk));
	jdff dff_A_YMitZxPN7_1(.dout(w_dff_A_DxZAQzaO9_1),.din(w_dff_A_YMitZxPN7_1),.clk(gclk));
	jdff dff_A_tc6v9mLJ2_1(.dout(w_dff_A_YMitZxPN7_1),.din(w_dff_A_tc6v9mLJ2_1),.clk(gclk));
	jdff dff_A_D7MDysKd6_1(.dout(w_dff_A_tc6v9mLJ2_1),.din(w_dff_A_D7MDysKd6_1),.clk(gclk));
	jdff dff_A_4a1uEYYr2_1(.dout(w_dff_A_D7MDysKd6_1),.din(w_dff_A_4a1uEYYr2_1),.clk(gclk));
	jdff dff_A_3oJZCltt9_1(.dout(w_dff_A_4a1uEYYr2_1),.din(w_dff_A_3oJZCltt9_1),.clk(gclk));
	jdff dff_A_LQDSPVtc1_1(.dout(w_dff_A_3oJZCltt9_1),.din(w_dff_A_LQDSPVtc1_1),.clk(gclk));
	jdff dff_A_iGsFYc2f1_1(.dout(w_dff_A_LQDSPVtc1_1),.din(w_dff_A_iGsFYc2f1_1),.clk(gclk));
	jdff dff_A_8ygS51Vp9_1(.dout(w_dff_A_iGsFYc2f1_1),.din(w_dff_A_8ygS51Vp9_1),.clk(gclk));
	jdff dff_A_tZIMvvsQ3_1(.dout(w_dff_A_8ygS51Vp9_1),.din(w_dff_A_tZIMvvsQ3_1),.clk(gclk));
	jdff dff_A_9eFk9Aht4_1(.dout(w_dff_A_tZIMvvsQ3_1),.din(w_dff_A_9eFk9Aht4_1),.clk(gclk));
	jdff dff_A_bvENYMJC6_2(.dout(w_n564_0[2]),.din(w_dff_A_bvENYMJC6_2),.clk(gclk));
	jdff dff_A_8HZhCT4c0_2(.dout(w_dff_A_bvENYMJC6_2),.din(w_dff_A_8HZhCT4c0_2),.clk(gclk));
	jdff dff_A_QLaHShLO6_0(.dout(w_n558_0[0]),.din(w_dff_A_QLaHShLO6_0),.clk(gclk));
	jdff dff_A_wYCagy7e1_1(.dout(w_n556_0[1]),.din(w_dff_A_wYCagy7e1_1),.clk(gclk));
	jdff dff_A_BA1F0Zgy1_2(.dout(w_n556_0[2]),.din(w_dff_A_BA1F0Zgy1_2),.clk(gclk));
	jdff dff_A_EzDBjIMm5_2(.dout(w_dff_A_BA1F0Zgy1_2),.din(w_dff_A_EzDBjIMm5_2),.clk(gclk));
	jdff dff_A_JTbuxVf88_2(.dout(w_dff_A_EzDBjIMm5_2),.din(w_dff_A_JTbuxVf88_2),.clk(gclk));
	jdff dff_A_dPBMJ54I4_0(.dout(w_n550_0[0]),.din(w_dff_A_dPBMJ54I4_0),.clk(gclk));
	jdff dff_A_6RKzcdbo6_0(.dout(w_dff_A_dPBMJ54I4_0),.din(w_dff_A_6RKzcdbo6_0),.clk(gclk));
	jdff dff_A_3cuPesp66_0(.dout(w_dff_A_6RKzcdbo6_0),.din(w_dff_A_3cuPesp66_0),.clk(gclk));
	jdff dff_A_Z193WOGo5_0(.dout(w_dff_A_3cuPesp66_0),.din(w_dff_A_Z193WOGo5_0),.clk(gclk));
	jdff dff_A_KhFQ59lS2_0(.dout(w_dff_A_Z193WOGo5_0),.din(w_dff_A_KhFQ59lS2_0),.clk(gclk));
	jdff dff_A_C08UO7vJ2_1(.dout(w_n548_0[1]),.din(w_dff_A_C08UO7vJ2_1),.clk(gclk));
	jdff dff_A_p8TbQbTy4_1(.dout(w_dff_A_C08UO7vJ2_1),.din(w_dff_A_p8TbQbTy4_1),.clk(gclk));
	jdff dff_A_4S11vnnI9_1(.dout(w_dff_A_p8TbQbTy4_1),.din(w_dff_A_4S11vnnI9_1),.clk(gclk));
	jdff dff_A_TZznZrcF6_1(.dout(w_dff_A_4S11vnnI9_1),.din(w_dff_A_TZznZrcF6_1),.clk(gclk));
	jdff dff_A_VK935xeR7_1(.dout(w_dff_A_TZznZrcF6_1),.din(w_dff_A_VK935xeR7_1),.clk(gclk));
	jdff dff_A_Lsy9KzB41_1(.dout(w_n1310_0[1]),.din(w_dff_A_Lsy9KzB41_1),.clk(gclk));
	jdff dff_A_7hPF4fB09_1(.dout(w_dff_A_Lsy9KzB41_1),.din(w_dff_A_7hPF4fB09_1),.clk(gclk));
	jdff dff_B_KJ16u6mD3_2(.din(n1310),.dout(w_dff_B_KJ16u6mD3_2),.clk(gclk));
	jdff dff_B_CVqjWA7C4_2(.din(w_dff_B_KJ16u6mD3_2),.dout(w_dff_B_CVqjWA7C4_2),.clk(gclk));
	jdff dff_B_7Y9ChrHQ0_2(.din(w_dff_B_CVqjWA7C4_2),.dout(w_dff_B_7Y9ChrHQ0_2),.clk(gclk));
	jdff dff_B_aHyXyoDH8_2(.din(w_dff_B_7Y9ChrHQ0_2),.dout(w_dff_B_aHyXyoDH8_2),.clk(gclk));
	jdff dff_B_iZ6gBjLr1_2(.din(w_dff_B_aHyXyoDH8_2),.dout(w_dff_B_iZ6gBjLr1_2),.clk(gclk));
	jdff dff_B_E97Us8X46_2(.din(w_dff_B_iZ6gBjLr1_2),.dout(w_dff_B_E97Us8X46_2),.clk(gclk));
	jdff dff_B_K5x5SohI6_2(.din(w_dff_B_E97Us8X46_2),.dout(w_dff_B_K5x5SohI6_2),.clk(gclk));
	jdff dff_B_cMRHQBCL1_2(.din(w_dff_B_K5x5SohI6_2),.dout(w_dff_B_cMRHQBCL1_2),.clk(gclk));
	jdff dff_A_ysMVdwFZ3_0(.dout(w_n581_0[0]),.din(w_dff_A_ysMVdwFZ3_0),.clk(gclk));
	jdff dff_A_gPzslvf37_0(.dout(w_dff_A_ysMVdwFZ3_0),.din(w_dff_A_gPzslvf37_0),.clk(gclk));
	jdff dff_A_vuvPEHOq4_0(.dout(w_dff_A_gPzslvf37_0),.din(w_dff_A_vuvPEHOq4_0),.clk(gclk));
	jdff dff_A_6AioAxSI3_0(.dout(w_dff_A_vuvPEHOq4_0),.din(w_dff_A_6AioAxSI3_0),.clk(gclk));
	jdff dff_A_PWTQCgE72_0(.dout(w_dff_A_6AioAxSI3_0),.din(w_dff_A_PWTQCgE72_0),.clk(gclk));
	jdff dff_A_vCz0QbXB2_0(.dout(w_dff_A_PWTQCgE72_0),.din(w_dff_A_vCz0QbXB2_0),.clk(gclk));
	jdff dff_A_kU1oxVam1_0(.dout(w_dff_A_vCz0QbXB2_0),.din(w_dff_A_kU1oxVam1_0),.clk(gclk));
	jdff dff_A_71DzBzYo3_2(.dout(w_n581_0[2]),.din(w_dff_A_71DzBzYo3_2),.clk(gclk));
	jdff dff_A_3sBOF4St6_2(.dout(w_dff_A_71DzBzYo3_2),.din(w_dff_A_3sBOF4St6_2),.clk(gclk));
	jdff dff_A_dB2iJaPX3_2(.dout(w_dff_A_3sBOF4St6_2),.din(w_dff_A_dB2iJaPX3_2),.clk(gclk));
	jdff dff_A_p9pMCzO73_2(.dout(w_dff_A_dB2iJaPX3_2),.din(w_dff_A_p9pMCzO73_2),.clk(gclk));
	jdff dff_A_p3KhwOOd0_2(.dout(w_dff_A_p9pMCzO73_2),.din(w_dff_A_p3KhwOOd0_2),.clk(gclk));
	jdff dff_A_W2jkEVHY0_2(.dout(w_dff_A_p3KhwOOd0_2),.din(w_dff_A_W2jkEVHY0_2),.clk(gclk));
	jdff dff_A_oTKXff7P4_2(.dout(w_dff_A_W2jkEVHY0_2),.din(w_dff_A_oTKXff7P4_2),.clk(gclk));
	jdff dff_A_miJ4WaIk0_2(.dout(w_dff_A_oTKXff7P4_2),.din(w_dff_A_miJ4WaIk0_2),.clk(gclk));
	jdff dff_A_IZiN2qeO5_2(.dout(w_dff_A_miJ4WaIk0_2),.din(w_dff_A_IZiN2qeO5_2),.clk(gclk));
	jdff dff_A_GY5bjR3s4_2(.dout(w_dff_A_IZiN2qeO5_2),.din(w_dff_A_GY5bjR3s4_2),.clk(gclk));
	jdff dff_A_GXXDDDUQ5_2(.dout(w_dff_A_GY5bjR3s4_2),.din(w_dff_A_GXXDDDUQ5_2),.clk(gclk));
	jdff dff_A_2Cawg4TM3_0(.dout(w_n580_0[0]),.din(w_dff_A_2Cawg4TM3_0),.clk(gclk));
	jdff dff_A_xgz65GIG9_0(.dout(w_dff_A_2Cawg4TM3_0),.din(w_dff_A_xgz65GIG9_0),.clk(gclk));
	jdff dff_A_Wfs2Q56b3_0(.dout(w_dff_A_xgz65GIG9_0),.din(w_dff_A_Wfs2Q56b3_0),.clk(gclk));
	jdff dff_A_t67qWl7n1_0(.dout(w_dff_A_Wfs2Q56b3_0),.din(w_dff_A_t67qWl7n1_0),.clk(gclk));
	jdff dff_A_kCaYLmSo8_0(.dout(w_dff_A_t67qWl7n1_0),.din(w_dff_A_kCaYLmSo8_0),.clk(gclk));
	jdff dff_A_CugJAFDh4_0(.dout(w_dff_A_kCaYLmSo8_0),.din(w_dff_A_CugJAFDh4_0),.clk(gclk));
	jdff dff_A_l2nWqKwK2_0(.dout(w_dff_A_CugJAFDh4_0),.din(w_dff_A_l2nWqKwK2_0),.clk(gclk));
	jdff dff_A_IAVF5e637_1(.dout(w_n580_0[1]),.din(w_dff_A_IAVF5e637_1),.clk(gclk));
	jdff dff_A_pkWrhgyj1_1(.dout(w_dff_A_IAVF5e637_1),.din(w_dff_A_pkWrhgyj1_1),.clk(gclk));
	jdff dff_A_azkasoZy5_1(.dout(w_dff_A_pkWrhgyj1_1),.din(w_dff_A_azkasoZy5_1),.clk(gclk));
	jdff dff_A_6d1kYrZC2_1(.dout(w_dff_A_azkasoZy5_1),.din(w_dff_A_6d1kYrZC2_1),.clk(gclk));
	jdff dff_A_BvaK4DRU8_1(.dout(w_dff_A_6d1kYrZC2_1),.din(w_dff_A_BvaK4DRU8_1),.clk(gclk));
	jdff dff_A_M2QEomtA6_1(.dout(w_dff_A_BvaK4DRU8_1),.din(w_dff_A_M2QEomtA6_1),.clk(gclk));
	jdff dff_A_CZEXJRqe6_1(.dout(w_dff_A_M2QEomtA6_1),.din(w_dff_A_CZEXJRqe6_1),.clk(gclk));
	jdff dff_A_4esIxRVH1_1(.dout(w_dff_A_CZEXJRqe6_1),.din(w_dff_A_4esIxRVH1_1),.clk(gclk));
	jdff dff_A_5xWiSkwM3_1(.dout(w_dff_A_4esIxRVH1_1),.din(w_dff_A_5xWiSkwM3_1),.clk(gclk));
	jdff dff_A_L9qQU0RR2_1(.dout(w_dff_A_5xWiSkwM3_1),.din(w_dff_A_L9qQU0RR2_1),.clk(gclk));
	jdff dff_A_k2kAb4RG9_1(.dout(w_dff_A_L9qQU0RR2_1),.din(w_dff_A_k2kAb4RG9_1),.clk(gclk));
	jdff dff_A_mon5JnRv2_1(.dout(w_dff_A_k2kAb4RG9_1),.din(w_dff_A_mon5JnRv2_1),.clk(gclk));
	jdff dff_A_lqffWO2G4_0(.dout(w_n578_0[0]),.din(w_dff_A_lqffWO2G4_0),.clk(gclk));
	jdff dff_A_acD5kKi72_1(.dout(w_n578_0[1]),.din(w_dff_A_acD5kKi72_1),.clk(gclk));
	jdff dff_A_B8ZxuV172_1(.dout(w_dff_A_acD5kKi72_1),.din(w_dff_A_B8ZxuV172_1),.clk(gclk));
	jdff dff_A_Au93wacp1_1(.dout(w_dff_A_B8ZxuV172_1),.din(w_dff_A_Au93wacp1_1),.clk(gclk));
	jdff dff_A_3gxpf3SG0_1(.dout(w_dff_A_Au93wacp1_1),.din(w_dff_A_3gxpf3SG0_1),.clk(gclk));
	jdff dff_A_CUgKotio2_1(.dout(w_dff_A_3gxpf3SG0_1),.din(w_dff_A_CUgKotio2_1),.clk(gclk));
	jdff dff_A_JmJgEfVy3_1(.dout(w_dff_A_CUgKotio2_1),.din(w_dff_A_JmJgEfVy3_1),.clk(gclk));
	jdff dff_A_9j9WAkp86_1(.dout(w_dff_A_JmJgEfVy3_1),.din(w_dff_A_9j9WAkp86_1),.clk(gclk));
	jdff dff_A_UhJAmNbx4_1(.dout(w_dff_A_9j9WAkp86_1),.din(w_dff_A_UhJAmNbx4_1),.clk(gclk));
	jdff dff_A_W0e2XS114_1(.dout(w_dff_A_UhJAmNbx4_1),.din(w_dff_A_W0e2XS114_1),.clk(gclk));
	jdff dff_A_SJvgTQ1q5_1(.dout(w_dff_A_W0e2XS114_1),.din(w_dff_A_SJvgTQ1q5_1),.clk(gclk));
	jdff dff_A_kOxryNfs6_1(.dout(w_dff_A_SJvgTQ1q5_1),.din(w_dff_A_kOxryNfs6_1),.clk(gclk));
	jdff dff_A_OpJIBC5E1_1(.dout(w_dff_A_kOxryNfs6_1),.din(w_dff_A_OpJIBC5E1_1),.clk(gclk));
	jdff dff_A_zYOezuNr4_1(.dout(w_dff_A_OpJIBC5E1_1),.din(w_dff_A_zYOezuNr4_1),.clk(gclk));
	jdff dff_A_tXO1PP5z8_1(.dout(w_dff_A_zYOezuNr4_1),.din(w_dff_A_tXO1PP5z8_1),.clk(gclk));
	jdff dff_A_yeAsge4y4_1(.dout(w_dff_A_tXO1PP5z8_1),.din(w_dff_A_yeAsge4y4_1),.clk(gclk));
	jdff dff_A_0TdKwvQd0_1(.dout(w_dff_A_yeAsge4y4_1),.din(w_dff_A_0TdKwvQd0_1),.clk(gclk));
	jdff dff_B_qIPZoZRM4_1(.din(n545),.dout(w_dff_B_qIPZoZRM4_1),.clk(gclk));
	jdff dff_B_Riboc5A53_0(.din(G94),.dout(w_dff_B_Riboc5A53_0),.clk(gclk));
	jdff dff_B_XccfJ9tn6_2(.din(n544),.dout(w_dff_B_XccfJ9tn6_2),.clk(gclk));
	jdff dff_B_ihvAxHVv3_2(.din(w_dff_B_XccfJ9tn6_2),.dout(w_dff_B_ihvAxHVv3_2),.clk(gclk));
	jdff dff_A_xgTb31pd1_0(.dout(w_G4405_1[0]),.din(w_dff_A_xgTb31pd1_0),.clk(gclk));
	jdff dff_A_v88eWpYU9_0(.dout(w_dff_A_xgTb31pd1_0),.din(w_dff_A_v88eWpYU9_0),.clk(gclk));
	jdff dff_A_1WAWknsy7_0(.dout(w_dff_A_v88eWpYU9_0),.din(w_dff_A_1WAWknsy7_0),.clk(gclk));
	jdff dff_A_lTrelQPG1_0(.dout(w_dff_A_1WAWknsy7_0),.din(w_dff_A_lTrelQPG1_0),.clk(gclk));
	jdff dff_B_dQ2S0xJ08_1(.din(n537),.dout(w_dff_B_dQ2S0xJ08_1),.clk(gclk));
	jdff dff_B_p60qXJgH6_0(.din(G121),.dout(w_dff_B_p60qXJgH6_0),.clk(gclk));
	jdff dff_A_f9O9ovBw2_1(.dout(w_n536_0[1]),.din(w_dff_A_f9O9ovBw2_1),.clk(gclk));
	jdff dff_A_dLMjmZVF5_1(.dout(w_dff_A_f9O9ovBw2_1),.din(w_dff_A_dLMjmZVF5_1),.clk(gclk));
	jdff dff_A_1px5iE7k2_2(.dout(w_n536_0[2]),.din(w_dff_A_1px5iE7k2_2),.clk(gclk));
	jdff dff_A_TgcstwJn7_2(.dout(w_dff_A_1px5iE7k2_2),.din(w_dff_A_TgcstwJn7_2),.clk(gclk));
	jdff dff_A_jCIFrJNW2_1(.dout(w_G4410_0[1]),.din(w_dff_A_jCIFrJNW2_1),.clk(gclk));
	jdff dff_A_7Htipfr83_1(.dout(w_dff_A_jCIFrJNW2_1),.din(w_dff_A_7Htipfr83_1),.clk(gclk));
	jdff dff_A_XpHdLBPY4_1(.dout(w_dff_A_7Htipfr83_1),.din(w_dff_A_XpHdLBPY4_1),.clk(gclk));
	jdff dff_A_9wSeb58Q6_1(.dout(w_dff_A_XpHdLBPY4_1),.din(w_dff_A_9wSeb58Q6_1),.clk(gclk));
	jdff dff_A_N3WShLZG1_0(.dout(w_n576_0[0]),.din(w_dff_A_N3WShLZG1_0),.clk(gclk));
	jdff dff_A_DvtYQeO81_0(.dout(w_dff_A_N3WShLZG1_0),.din(w_dff_A_DvtYQeO81_0),.clk(gclk));
	jdff dff_A_4FiJ6Abm9_0(.dout(w_dff_A_DvtYQeO81_0),.din(w_dff_A_4FiJ6Abm9_0),.clk(gclk));
	jdff dff_A_kabXAEER0_0(.dout(w_dff_A_4FiJ6Abm9_0),.din(w_dff_A_kabXAEER0_0),.clk(gclk));
	jdff dff_A_PPGF0MwR1_0(.dout(w_dff_A_kabXAEER0_0),.din(w_dff_A_PPGF0MwR1_0),.clk(gclk));
	jdff dff_A_PNH8FUOz4_0(.dout(w_dff_A_PPGF0MwR1_0),.din(w_dff_A_PNH8FUOz4_0),.clk(gclk));
	jdff dff_A_sNYJcCNi8_0(.dout(w_dff_A_PNH8FUOz4_0),.din(w_dff_A_sNYJcCNi8_0),.clk(gclk));
	jdff dff_A_kB8hMKWp6_0(.dout(w_dff_A_sNYJcCNi8_0),.din(w_dff_A_kB8hMKWp6_0),.clk(gclk));
	jdff dff_A_u3019IJd7_0(.dout(w_dff_A_kB8hMKWp6_0),.din(w_dff_A_u3019IJd7_0),.clk(gclk));
	jdff dff_A_wcaFuKEE8_0(.dout(w_dff_A_u3019IJd7_0),.din(w_dff_A_wcaFuKEE8_0),.clk(gclk));
	jdff dff_A_bGViTR6f4_0(.dout(w_dff_A_wcaFuKEE8_0),.din(w_dff_A_bGViTR6f4_0),.clk(gclk));
	jdff dff_A_a9XS4HMB7_0(.dout(w_dff_A_bGViTR6f4_0),.din(w_dff_A_a9XS4HMB7_0),.clk(gclk));
	jdff dff_A_hz18Lgjr9_0(.dout(w_dff_A_a9XS4HMB7_0),.din(w_dff_A_hz18Lgjr9_0),.clk(gclk));
	jdff dff_A_NvpZ0mFy4_0(.dout(w_n575_1[0]),.din(w_dff_A_NvpZ0mFy4_0),.clk(gclk));
	jdff dff_A_WVd6taLi7_0(.dout(w_dff_A_NvpZ0mFy4_0),.din(w_dff_A_WVd6taLi7_0),.clk(gclk));
	jdff dff_A_UHRhb0km1_0(.dout(w_dff_A_WVd6taLi7_0),.din(w_dff_A_UHRhb0km1_0),.clk(gclk));
	jdff dff_A_8o1EvQQ89_0(.dout(w_dff_A_UHRhb0km1_0),.din(w_dff_A_8o1EvQQ89_0),.clk(gclk));
	jdff dff_A_DPHt0NE36_0(.dout(w_dff_A_8o1EvQQ89_0),.din(w_dff_A_DPHt0NE36_0),.clk(gclk));
	jdff dff_A_amYwbKsM0_0(.dout(w_dff_A_DPHt0NE36_0),.din(w_dff_A_amYwbKsM0_0),.clk(gclk));
	jdff dff_A_Wq2N3hnR2_0(.dout(w_dff_A_amYwbKsM0_0),.din(w_dff_A_Wq2N3hnR2_0),.clk(gclk));
	jdff dff_A_V1PNa2iC3_0(.dout(w_dff_A_Wq2N3hnR2_0),.din(w_dff_A_V1PNa2iC3_0),.clk(gclk));
	jdff dff_A_IkU1o7ym0_0(.dout(w_dff_A_V1PNa2iC3_0),.din(w_dff_A_IkU1o7ym0_0),.clk(gclk));
	jdff dff_A_fwOiAooC4_0(.dout(w_dff_A_IkU1o7ym0_0),.din(w_dff_A_fwOiAooC4_0),.clk(gclk));
	jdff dff_A_OvfXvPDW2_0(.dout(w_dff_A_fwOiAooC4_0),.din(w_dff_A_OvfXvPDW2_0),.clk(gclk));
	jdff dff_A_D2ClmSTB0_0(.dout(w_dff_A_OvfXvPDW2_0),.din(w_dff_A_D2ClmSTB0_0),.clk(gclk));
	jdff dff_A_BEQMLTWM3_0(.dout(w_dff_A_D2ClmSTB0_0),.din(w_dff_A_BEQMLTWM3_0),.clk(gclk));
	jdff dff_A_8x3bmntu0_0(.dout(w_dff_A_BEQMLTWM3_0),.din(w_dff_A_8x3bmntu0_0),.clk(gclk));
	jdff dff_A_p4US44f95_2(.dout(w_n575_0[2]),.din(w_dff_A_p4US44f95_2),.clk(gclk));
	jdff dff_A_u22XtAVW7_2(.dout(w_dff_A_p4US44f95_2),.din(w_dff_A_u22XtAVW7_2),.clk(gclk));
	jdff dff_A_736VvCll4_2(.dout(w_dff_A_u22XtAVW7_2),.din(w_dff_A_736VvCll4_2),.clk(gclk));
	jdff dff_A_nlQeMzFL1_2(.dout(w_dff_A_736VvCll4_2),.din(w_dff_A_nlQeMzFL1_2),.clk(gclk));
	jdff dff_A_pundBuOL3_2(.dout(w_dff_A_nlQeMzFL1_2),.din(w_dff_A_pundBuOL3_2),.clk(gclk));
	jdff dff_A_rSR9TcK67_2(.dout(w_dff_A_pundBuOL3_2),.din(w_dff_A_rSR9TcK67_2),.clk(gclk));
	jdff dff_A_uweABs4V3_2(.dout(w_dff_A_rSR9TcK67_2),.din(w_dff_A_uweABs4V3_2),.clk(gclk));
	jdff dff_A_Jnt2VpNM3_2(.dout(w_dff_A_uweABs4V3_2),.din(w_dff_A_Jnt2VpNM3_2),.clk(gclk));
	jdff dff_A_hUGxjfsN8_2(.dout(w_dff_A_Jnt2VpNM3_2),.din(w_dff_A_hUGxjfsN8_2),.clk(gclk));
	jdff dff_A_2HpiObd17_2(.dout(w_dff_A_hUGxjfsN8_2),.din(w_dff_A_2HpiObd17_2),.clk(gclk));
	jdff dff_A_xAiIsYas7_2(.dout(w_dff_A_2HpiObd17_2),.din(w_dff_A_xAiIsYas7_2),.clk(gclk));
	jdff dff_A_atlK1W1j0_2(.dout(w_dff_A_xAiIsYas7_2),.din(w_dff_A_atlK1W1j0_2),.clk(gclk));
	jdff dff_A_YRz67tca0_2(.dout(w_dff_A_atlK1W1j0_2),.din(w_dff_A_YRz67tca0_2),.clk(gclk));
	jdff dff_A_7r7a95wO4_2(.dout(w_dff_A_YRz67tca0_2),.din(w_dff_A_7r7a95wO4_2),.clk(gclk));
	jdff dff_B_5J78YsqT1_1(.din(n561),.dout(w_dff_B_5J78YsqT1_1),.clk(gclk));
	jdff dff_B_3iz5PsYf1_0(.din(G118),.dout(w_dff_B_3iz5PsYf1_0),.clk(gclk));
	jdff dff_B_VwWmTBK90_2(.din(n560),.dout(w_dff_B_VwWmTBK90_2),.clk(gclk));
	jdff dff_B_7TqLiHyu6_2(.din(w_dff_B_VwWmTBK90_2),.dout(w_dff_B_7TqLiHyu6_2),.clk(gclk));
	jdff dff_A_Pkfnl6f13_2(.dout(w_G4394_0[2]),.din(w_dff_A_Pkfnl6f13_2),.clk(gclk));
	jdff dff_A_iuaibS5Y5_2(.dout(w_dff_A_Pkfnl6f13_2),.din(w_dff_A_iuaibS5Y5_2),.clk(gclk));
	jdff dff_A_yzUKPOdA1_2(.dout(w_dff_A_iuaibS5Y5_2),.din(w_dff_A_yzUKPOdA1_2),.clk(gclk));
	jdff dff_A_IutNNJpv4_2(.dout(w_dff_A_yzUKPOdA1_2),.din(w_dff_A_IutNNJpv4_2),.clk(gclk));
	jdff dff_A_OC50sEMX8_1(.dout(w_n574_0[1]),.din(w_dff_A_OC50sEMX8_1),.clk(gclk));
	jdff dff_A_jAzB48uU8_1(.dout(w_dff_A_OC50sEMX8_1),.din(w_dff_A_jAzB48uU8_1),.clk(gclk));
	jdff dff_A_Av1rnJiU2_1(.dout(w_dff_A_jAzB48uU8_1),.din(w_dff_A_Av1rnJiU2_1),.clk(gclk));
	jdff dff_A_RaQj24hW2_1(.dout(w_dff_A_Av1rnJiU2_1),.din(w_dff_A_RaQj24hW2_1),.clk(gclk));
	jdff dff_A_bW3y7cdp8_1(.dout(w_dff_A_RaQj24hW2_1),.din(w_dff_A_bW3y7cdp8_1),.clk(gclk));
	jdff dff_A_e4WQQvfR9_1(.dout(w_dff_A_bW3y7cdp8_1),.din(w_dff_A_e4WQQvfR9_1),.clk(gclk));
	jdff dff_A_MVe4SJEJ1_1(.dout(w_dff_A_e4WQQvfR9_1),.din(w_dff_A_MVe4SJEJ1_1),.clk(gclk));
	jdff dff_A_B2WhMACO0_1(.dout(w_dff_A_MVe4SJEJ1_1),.din(w_dff_A_B2WhMACO0_1),.clk(gclk));
	jdff dff_A_SZ5m0Uam4_1(.dout(w_dff_A_B2WhMACO0_1),.din(w_dff_A_SZ5m0Uam4_1),.clk(gclk));
	jdff dff_A_sOGc9nEV3_1(.dout(w_dff_A_SZ5m0Uam4_1),.din(w_dff_A_sOGc9nEV3_1),.clk(gclk));
	jdff dff_A_S9zR2MoY0_1(.dout(w_dff_A_sOGc9nEV3_1),.din(w_dff_A_S9zR2MoY0_1),.clk(gclk));
	jdff dff_A_DxrbamLN8_1(.dout(w_dff_A_S9zR2MoY0_1),.din(w_dff_A_DxrbamLN8_1),.clk(gclk));
	jdff dff_A_ddPo7jrP3_1(.dout(w_dff_A_DxrbamLN8_1),.din(w_dff_A_ddPo7jrP3_1),.clk(gclk));
	jdff dff_A_fVl5iCD92_1(.dout(w_dff_A_ddPo7jrP3_1),.din(w_dff_A_fVl5iCD92_1),.clk(gclk));
	jdff dff_A_b6AGPVkI5_1(.dout(w_dff_A_fVl5iCD92_1),.din(w_dff_A_b6AGPVkI5_1),.clk(gclk));
	jdff dff_A_ygwklOHH0_1(.dout(w_dff_A_b6AGPVkI5_1),.din(w_dff_A_ygwklOHH0_1),.clk(gclk));
	jdff dff_B_38xGnxtj6_1(.din(n553),.dout(w_dff_B_38xGnxtj6_1),.clk(gclk));
	jdff dff_B_7tTp421h9_0(.din(G97),.dout(w_dff_B_7tTp421h9_0),.clk(gclk));
	jdff dff_B_PVbhmyMo4_2(.din(n552),.dout(w_dff_B_PVbhmyMo4_2),.clk(gclk));
	jdff dff_B_BCtcMeMM9_2(.din(w_dff_B_PVbhmyMo4_2),.dout(w_dff_B_BCtcMeMM9_2),.clk(gclk));
	jdff dff_A_xmQWixmU5_0(.dout(w_G4400_1[0]),.din(w_dff_A_xmQWixmU5_0),.clk(gclk));
	jdff dff_A_jNF1ql180_0(.dout(w_dff_A_xmQWixmU5_0),.din(w_dff_A_jNF1ql180_0),.clk(gclk));
	jdff dff_A_Og3rJbXB4_0(.dout(w_dff_A_jNF1ql180_0),.din(w_dff_A_Og3rJbXB4_0),.clk(gclk));
	jdff dff_A_sFIkmB0G0_0(.dout(w_dff_A_Og3rJbXB4_0),.din(w_dff_A_sFIkmB0G0_0),.clk(gclk));
	jdff dff_A_7fuK7RtU0_0(.dout(w_n573_1[0]),.din(w_dff_A_7fuK7RtU0_0),.clk(gclk));
	jdff dff_A_6izLRkuO9_0(.dout(w_dff_A_7fuK7RtU0_0),.din(w_dff_A_6izLRkuO9_0),.clk(gclk));
	jdff dff_A_rXlwLnIN3_0(.dout(w_dff_A_6izLRkuO9_0),.din(w_dff_A_rXlwLnIN3_0),.clk(gclk));
	jdff dff_A_T1k0BBKT5_0(.dout(w_dff_A_rXlwLnIN3_0),.din(w_dff_A_T1k0BBKT5_0),.clk(gclk));
	jdff dff_A_E6ImUlFE7_0(.dout(w_dff_A_T1k0BBKT5_0),.din(w_dff_A_E6ImUlFE7_0),.clk(gclk));
	jdff dff_A_yPefPCJk6_0(.dout(w_dff_A_E6ImUlFE7_0),.din(w_dff_A_yPefPCJk6_0),.clk(gclk));
	jdff dff_A_tz40ulXB7_0(.dout(w_dff_A_yPefPCJk6_0),.din(w_dff_A_tz40ulXB7_0),.clk(gclk));
	jdff dff_A_42BOIvwl5_0(.dout(w_dff_A_tz40ulXB7_0),.din(w_dff_A_42BOIvwl5_0),.clk(gclk));
	jdff dff_A_fuCPdAOi6_0(.dout(w_dff_A_42BOIvwl5_0),.din(w_dff_A_fuCPdAOi6_0),.clk(gclk));
	jdff dff_A_kEQhtFmE3_0(.dout(w_dff_A_fuCPdAOi6_0),.din(w_dff_A_kEQhtFmE3_0),.clk(gclk));
	jdff dff_A_Glr05qO79_0(.dout(w_dff_A_kEQhtFmE3_0),.din(w_dff_A_Glr05qO79_0),.clk(gclk));
	jdff dff_A_C08EW8Rb1_0(.dout(w_dff_A_Glr05qO79_0),.din(w_dff_A_C08EW8Rb1_0),.clk(gclk));
	jdff dff_A_qittnX8T7_0(.dout(w_dff_A_C08EW8Rb1_0),.din(w_dff_A_qittnX8T7_0),.clk(gclk));
	jdff dff_A_LvjM02uI6_0(.dout(w_dff_A_qittnX8T7_0),.din(w_dff_A_LvjM02uI6_0),.clk(gclk));
	jdff dff_A_hLOoceXz1_1(.dout(w_n573_0[1]),.din(w_dff_A_hLOoceXz1_1),.clk(gclk));
	jdff dff_A_oYqyl08q4_1(.dout(w_dff_A_hLOoceXz1_1),.din(w_dff_A_oYqyl08q4_1),.clk(gclk));
	jdff dff_A_MNSi9QRU8_1(.dout(w_dff_A_oYqyl08q4_1),.din(w_dff_A_MNSi9QRU8_1),.clk(gclk));
	jdff dff_A_mvKoU86b7_2(.dout(w_n573_0[2]),.din(w_dff_A_mvKoU86b7_2),.clk(gclk));
	jdff dff_A_tuR61V1o1_2(.dout(w_dff_A_mvKoU86b7_2),.din(w_dff_A_tuR61V1o1_2),.clk(gclk));
	jdff dff_B_9C4K4mYd5_3(.din(n573),.dout(w_dff_B_9C4K4mYd5_3),.clk(gclk));
	jdff dff_B_8mpWh9QD7_3(.din(w_dff_B_9C4K4mYd5_3),.dout(w_dff_B_8mpWh9QD7_3),.clk(gclk));
	jdff dff_B_t9qFBe8s0_1(.din(n529),.dout(w_dff_B_t9qFBe8s0_1),.clk(gclk));
	jdff dff_B_kRuWr5Ze3_0(.din(G47),.dout(w_dff_B_kRuWr5Ze3_0),.clk(gclk));
	jdff dff_B_N7qyj0SS7_2(.din(n528),.dout(w_dff_B_N7qyj0SS7_2),.clk(gclk));
	jdff dff_B_O4P7ekHV9_2(.din(w_dff_B_N7qyj0SS7_2),.dout(w_dff_B_O4P7ekHV9_2),.clk(gclk));
	jdff dff_A_0KBxwsSj2_0(.dout(w_G4415_1[0]),.din(w_dff_A_0KBxwsSj2_0),.clk(gclk));
	jdff dff_A_aLmk8uKN5_0(.dout(w_dff_A_0KBxwsSj2_0),.din(w_dff_A_aLmk8uKN5_0),.clk(gclk));
	jdff dff_A_jyj8FSGN1_0(.dout(w_dff_A_aLmk8uKN5_0),.din(w_dff_A_jyj8FSGN1_0),.clk(gclk));
	jdff dff_A_lnZFptbP4_0(.dout(w_dff_A_jyj8FSGN1_0),.din(w_dff_A_lnZFptbP4_0),.clk(gclk));
	jdff dff_B_1MnPFWTn6_1(.din(n589),.dout(w_dff_B_1MnPFWTn6_1),.clk(gclk));
	jdff dff_B_CzRc0bBz7_1(.din(w_dff_B_1MnPFWTn6_1),.dout(w_dff_B_CzRc0bBz7_1),.clk(gclk));
	jdff dff_B_e2BLbAhW4_1(.din(w_dff_B_CzRc0bBz7_1),.dout(w_dff_B_e2BLbAhW4_1),.clk(gclk));
	jdff dff_B_UDhXF6iJ1_1(.din(w_dff_B_e2BLbAhW4_1),.dout(w_dff_B_UDhXF6iJ1_1),.clk(gclk));
	jdff dff_B_BEhZtLA78_1(.din(w_dff_B_UDhXF6iJ1_1),.dout(w_dff_B_BEhZtLA78_1),.clk(gclk));
	jdff dff_B_BoOkr2Ex8_1(.din(w_dff_B_BEhZtLA78_1),.dout(w_dff_B_BoOkr2Ex8_1),.clk(gclk));
	jdff dff_B_kc1tfybA7_1(.din(w_dff_B_BoOkr2Ex8_1),.dout(w_dff_B_kc1tfybA7_1),.clk(gclk));
	jdff dff_B_O1q6X0h10_1(.din(w_dff_B_kc1tfybA7_1),.dout(w_dff_B_O1q6X0h10_1),.clk(gclk));
	jdff dff_B_jdSfgv1h5_1(.din(w_dff_B_O1q6X0h10_1),.dout(w_dff_B_jdSfgv1h5_1),.clk(gclk));
	jdff dff_B_88xv0lQT3_1(.din(w_dff_B_jdSfgv1h5_1),.dout(w_dff_B_88xv0lQT3_1),.clk(gclk));
	jdff dff_B_ldq4NBgL5_1(.din(n620),.dout(w_dff_B_ldq4NBgL5_1),.clk(gclk));
	jdff dff_B_xycWIFKM6_1(.din(w_dff_B_ldq4NBgL5_1),.dout(w_dff_B_xycWIFKM6_1),.clk(gclk));
	jdff dff_B_WyXqx9GF2_1(.din(w_dff_B_xycWIFKM6_1),.dout(w_dff_B_WyXqx9GF2_1),.clk(gclk));
	jdff dff_B_Sf0ECSPo6_1(.din(w_dff_B_WyXqx9GF2_1),.dout(w_dff_B_Sf0ECSPo6_1),.clk(gclk));
	jdff dff_B_eVzLRdWj1_1(.din(n621),.dout(w_dff_B_eVzLRdWj1_1),.clk(gclk));
	jdff dff_B_1qfAXtC86_1(.din(w_dff_B_eVzLRdWj1_1),.dout(w_dff_B_1qfAXtC86_1),.clk(gclk));
	jdff dff_B_nguaJ4fU0_1(.din(w_dff_B_1qfAXtC86_1),.dout(w_dff_B_nguaJ4fU0_1),.clk(gclk));
	jdff dff_B_Ok5coIGX5_1(.din(w_dff_B_nguaJ4fU0_1),.dout(w_dff_B_Ok5coIGX5_1),.clk(gclk));
	jdff dff_A_FBA4pPba7_0(.dout(w_G4526_2[0]),.din(w_dff_A_FBA4pPba7_0),.clk(gclk));
	jdff dff_A_SMOczHxq3_0(.dout(w_dff_A_FBA4pPba7_0),.din(w_dff_A_SMOczHxq3_0),.clk(gclk));
	jdff dff_A_BzVI7Hmc4_0(.dout(w_dff_A_SMOczHxq3_0),.din(w_dff_A_BzVI7Hmc4_0),.clk(gclk));
	jdff dff_A_otTBf6UK0_1(.dout(w_G4526_2[1]),.din(w_dff_A_otTBf6UK0_1),.clk(gclk));
	jdff dff_A_t8eUGYfF0_1(.dout(w_dff_A_otTBf6UK0_1),.din(w_dff_A_t8eUGYfF0_1),.clk(gclk));
	jdff dff_A_mFwHVCmR1_1(.dout(w_dff_A_t8eUGYfF0_1),.din(w_dff_A_mFwHVCmR1_1),.clk(gclk));
	jdff dff_A_B4YaPbWH1_1(.dout(w_dff_A_mFwHVCmR1_1),.din(w_dff_A_B4YaPbWH1_1),.clk(gclk));
	jdff dff_A_EaGWucWr5_1(.dout(w_dff_A_B4YaPbWH1_1),.din(w_dff_A_EaGWucWr5_1),.clk(gclk));
	jdff dff_A_1g1knSvq5_1(.dout(w_dff_A_EaGWucWr5_1),.din(w_dff_A_1g1knSvq5_1),.clk(gclk));
	jdff dff_A_KEpOUmLI6_1(.dout(w_dff_A_1g1knSvq5_1),.din(w_dff_A_KEpOUmLI6_1),.clk(gclk));
	jdff dff_A_Z9KREoSp5_0(.dout(w_n588_0[0]),.din(w_dff_A_Z9KREoSp5_0),.clk(gclk));
	jdff dff_A_cQ64OiLb2_0(.dout(w_dff_A_Z9KREoSp5_0),.din(w_dff_A_cQ64OiLb2_0),.clk(gclk));
	jdff dff_A_jwrJUxZu5_0(.dout(w_dff_A_cQ64OiLb2_0),.din(w_dff_A_jwrJUxZu5_0),.clk(gclk));
	jdff dff_A_YAzPImYi1_0(.dout(w_dff_A_jwrJUxZu5_0),.din(w_dff_A_YAzPImYi1_0),.clk(gclk));
	jdff dff_A_0D7DRRfH4_0(.dout(w_dff_A_YAzPImYi1_0),.din(w_dff_A_0D7DRRfH4_0),.clk(gclk));
	jdff dff_A_qSCmXCoz6_0(.dout(w_dff_A_0D7DRRfH4_0),.din(w_dff_A_qSCmXCoz6_0),.clk(gclk));
	jdff dff_A_9ieRz2IT8_0(.dout(w_dff_A_qSCmXCoz6_0),.din(w_dff_A_9ieRz2IT8_0),.clk(gclk));
	jdff dff_A_ulwkfI8V2_0(.dout(w_dff_A_9ieRz2IT8_0),.din(w_dff_A_ulwkfI8V2_0),.clk(gclk));
	jdff dff_A_I9cviMoA4_0(.dout(w_dff_A_ulwkfI8V2_0),.din(w_dff_A_I9cviMoA4_0),.clk(gclk));
	jdff dff_A_rE0JRAc74_0(.dout(w_dff_A_I9cviMoA4_0),.din(w_dff_A_rE0JRAc74_0),.clk(gclk));
	jdff dff_A_RjDBOhul3_0(.dout(w_dff_A_rE0JRAc74_0),.din(w_dff_A_RjDBOhul3_0),.clk(gclk));
	jdff dff_A_KNCJspG11_1(.dout(w_n586_0[1]),.din(w_dff_A_KNCJspG11_1),.clk(gclk));
	jdff dff_A_Rb3tevW70_1(.dout(w_dff_A_KNCJspG11_1),.din(w_dff_A_Rb3tevW70_1),.clk(gclk));
	jdff dff_A_YLKPixlB3_1(.dout(w_dff_A_Rb3tevW70_1),.din(w_dff_A_YLKPixlB3_1),.clk(gclk));
	jdff dff_A_2EbvKKd93_1(.dout(w_dff_A_YLKPixlB3_1),.din(w_dff_A_2EbvKKd93_1),.clk(gclk));
	jdff dff_A_hxTGiEPx4_1(.dout(w_dff_A_2EbvKKd93_1),.din(w_dff_A_hxTGiEPx4_1),.clk(gclk));
	jdff dff_A_GiUdOuoH4_1(.dout(w_dff_A_hxTGiEPx4_1),.din(w_dff_A_GiUdOuoH4_1),.clk(gclk));
	jdff dff_A_ZO06GEhO5_1(.dout(w_dff_A_GiUdOuoH4_1),.din(w_dff_A_ZO06GEhO5_1),.clk(gclk));
	jdff dff_A_OJGNnBwV2_1(.dout(w_dff_A_ZO06GEhO5_1),.din(w_dff_A_OJGNnBwV2_1),.clk(gclk));
	jdff dff_A_7qzebuRD8_1(.dout(w_dff_A_OJGNnBwV2_1),.din(w_dff_A_7qzebuRD8_1),.clk(gclk));
	jdff dff_A_vsLeinxy3_1(.dout(w_dff_A_7qzebuRD8_1),.din(w_dff_A_vsLeinxy3_1),.clk(gclk));
	jdff dff_A_FUS7ZetH6_1(.dout(w_dff_A_vsLeinxy3_1),.din(w_dff_A_FUS7ZetH6_1),.clk(gclk));
	jdff dff_A_wcIRTCIK3_1(.dout(w_dff_A_FUS7ZetH6_1),.din(w_dff_A_wcIRTCIK3_1),.clk(gclk));
	jdff dff_A_2tPgZb2z2_1(.dout(w_dff_A_wcIRTCIK3_1),.din(w_dff_A_2tPgZb2z2_1),.clk(gclk));
	jdff dff_A_McxqYnwG5_2(.dout(w_n586_0[2]),.din(w_dff_A_McxqYnwG5_2),.clk(gclk));
	jdff dff_A_eXL2fdfm5_2(.dout(w_dff_A_McxqYnwG5_2),.din(w_dff_A_eXL2fdfm5_2),.clk(gclk));
	jdff dff_A_WDwcHOGF9_2(.dout(w_dff_A_eXL2fdfm5_2),.din(w_dff_A_WDwcHOGF9_2),.clk(gclk));
	jdff dff_A_Oc5dMlRx2_2(.dout(w_dff_A_WDwcHOGF9_2),.din(w_dff_A_Oc5dMlRx2_2),.clk(gclk));
	jdff dff_A_aKAJ4X310_2(.dout(w_dff_A_Oc5dMlRx2_2),.din(w_dff_A_aKAJ4X310_2),.clk(gclk));
	jdff dff_A_hU48JwK29_2(.dout(w_dff_A_aKAJ4X310_2),.din(w_dff_A_hU48JwK29_2),.clk(gclk));
	jdff dff_A_Cn0Vxd4t7_2(.dout(w_dff_A_hU48JwK29_2),.din(w_dff_A_Cn0Vxd4t7_2),.clk(gclk));
	jdff dff_A_t8LjUqfe9_2(.dout(w_dff_A_Cn0Vxd4t7_2),.din(w_dff_A_t8LjUqfe9_2),.clk(gclk));
	jdff dff_A_RqBsZQBk7_2(.dout(w_dff_A_t8LjUqfe9_2),.din(w_dff_A_RqBsZQBk7_2),.clk(gclk));
	jdff dff_A_i9EFuq3a5_2(.dout(w_dff_A_RqBsZQBk7_2),.din(w_dff_A_i9EFuq3a5_2),.clk(gclk));
	jdff dff_A_45OF1Ef03_2(.dout(w_dff_A_i9EFuq3a5_2),.din(w_dff_A_45OF1Ef03_2),.clk(gclk));
	jdff dff_A_CYddlKxF6_2(.dout(w_dff_A_45OF1Ef03_2),.din(w_dff_A_CYddlKxF6_2),.clk(gclk));
	jdff dff_A_WKfWzS9X7_2(.dout(w_dff_A_CYddlKxF6_2),.din(w_dff_A_WKfWzS9X7_2),.clk(gclk));
	jdff dff_B_a7EzQSxI7_0(.din(n1631),.dout(w_dff_B_a7EzQSxI7_0),.clk(gclk));
	jdff dff_B_T3gQHh6T4_0(.din(w_dff_B_a7EzQSxI7_0),.dout(w_dff_B_T3gQHh6T4_0),.clk(gclk));
	jdff dff_B_CfL1mf701_0(.din(w_dff_B_T3gQHh6T4_0),.dout(w_dff_B_CfL1mf701_0),.clk(gclk));
	jdff dff_B_96jNs8Ki9_0(.din(w_dff_B_CfL1mf701_0),.dout(w_dff_B_96jNs8Ki9_0),.clk(gclk));
	jdff dff_B_BJI2hD937_0(.din(w_dff_B_96jNs8Ki9_0),.dout(w_dff_B_BJI2hD937_0),.clk(gclk));
	jdff dff_B_6qVgfeOH7_0(.din(w_dff_B_BJI2hD937_0),.dout(w_dff_B_6qVgfeOH7_0),.clk(gclk));
	jdff dff_B_8AUtE38n6_0(.din(w_dff_B_6qVgfeOH7_0),.dout(w_dff_B_8AUtE38n6_0),.clk(gclk));
	jdff dff_B_mNlrzDub2_0(.din(w_dff_B_8AUtE38n6_0),.dout(w_dff_B_mNlrzDub2_0),.clk(gclk));
	jdff dff_B_CuGglQsX9_0(.din(w_dff_B_mNlrzDub2_0),.dout(w_dff_B_CuGglQsX9_0),.clk(gclk));
	jdff dff_B_yktIWuvJ8_0(.din(w_dff_B_CuGglQsX9_0),.dout(w_dff_B_yktIWuvJ8_0),.clk(gclk));
	jdff dff_B_3p4fg0Jy6_0(.din(w_dff_B_yktIWuvJ8_0),.dout(w_dff_B_3p4fg0Jy6_0),.clk(gclk));
	jdff dff_B_HUTbIaS43_1(.din(n1621),.dout(w_dff_B_HUTbIaS43_1),.clk(gclk));
	jdff dff_B_ngg18DwO4_1(.din(w_dff_B_HUTbIaS43_1),.dout(w_dff_B_ngg18DwO4_1),.clk(gclk));
	jdff dff_B_rJyFWDR91_1(.din(n1622),.dout(w_dff_B_rJyFWDR91_1),.clk(gclk));
	jdff dff_A_KF6NnfZB2_0(.dout(w_n1620_0[0]),.din(w_dff_A_KF6NnfZB2_0),.clk(gclk));
	jdff dff_A_tNhpBkgq5_0(.dout(w_dff_A_KF6NnfZB2_0),.din(w_dff_A_tNhpBkgq5_0),.clk(gclk));
	jdff dff_B_zRmf5Vmx7_0(.din(n1617),.dout(w_dff_B_zRmf5Vmx7_0),.clk(gclk));
	jdff dff_B_0ZuZZlVW5_0(.din(w_dff_B_zRmf5Vmx7_0),.dout(w_dff_B_0ZuZZlVW5_0),.clk(gclk));
	jdff dff_B_kradYcl35_1(.din(n1611),.dout(w_dff_B_kradYcl35_1),.clk(gclk));
	jdff dff_B_R2AitHJL1_1(.din(w_dff_B_kradYcl35_1),.dout(w_dff_B_R2AitHJL1_1),.clk(gclk));
	jdff dff_B_Ak1eFJ806_1(.din(n1608),.dout(w_dff_B_Ak1eFJ806_1),.clk(gclk));
	jdff dff_B_uud4iB130_0(.din(n1609),.dout(w_dff_B_uud4iB130_0),.clk(gclk));
	jdff dff_B_XkQg6ELH9_0(.din(w_dff_B_uud4iB130_0),.dout(w_dff_B_XkQg6ELH9_0),.clk(gclk));
	jdff dff_B_oGy0A1gd7_0(.din(w_dff_B_XkQg6ELH9_0),.dout(w_dff_B_oGy0A1gd7_0),.clk(gclk));
	jdff dff_B_DeW867u91_0(.din(w_dff_B_oGy0A1gd7_0),.dout(w_dff_B_DeW867u91_0),.clk(gclk));
	jdff dff_B_YhKwkhYb7_0(.din(w_dff_B_DeW867u91_0),.dout(w_dff_B_YhKwkhYb7_0),.clk(gclk));
	jdff dff_A_4kWqaBCf0_0(.dout(w_n1607_0[0]),.din(w_dff_A_4kWqaBCf0_0),.clk(gclk));
	jdff dff_A_zAzTDnyc4_0(.dout(w_dff_A_4kWqaBCf0_0),.din(w_dff_A_zAzTDnyc4_0),.clk(gclk));
	jdff dff_A_WUvdjBcC0_0(.dout(w_dff_A_zAzTDnyc4_0),.din(w_dff_A_WUvdjBcC0_0),.clk(gclk));
	jdff dff_B_2Jgxhcxe8_0(.din(n1606),.dout(w_dff_B_2Jgxhcxe8_0),.clk(gclk));
	jdff dff_A_bDMyFFig2_0(.dout(w_n1605_0[0]),.din(w_dff_A_bDMyFFig2_0),.clk(gclk));
	jdff dff_A_feYm9Cay4_0(.dout(w_dff_A_bDMyFFig2_0),.din(w_dff_A_feYm9Cay4_0),.clk(gclk));
	jdff dff_A_6n6nbIef7_0(.dout(w_dff_A_feYm9Cay4_0),.din(w_dff_A_6n6nbIef7_0),.clk(gclk));
	jdff dff_A_TuTJ2ZQJ1_0(.dout(w_dff_A_6n6nbIef7_0),.din(w_dff_A_TuTJ2ZQJ1_0),.clk(gclk));
	jdff dff_A_qHTQzuGI7_0(.dout(w_dff_A_TuTJ2ZQJ1_0),.din(w_dff_A_qHTQzuGI7_0),.clk(gclk));
	jdff dff_B_oHa9ooEO4_0(.din(n1603),.dout(w_dff_B_oHa9ooEO4_0),.clk(gclk));
	jdff dff_B_AkmfGLxS3_1(.din(n1588),.dout(w_dff_B_AkmfGLxS3_1),.clk(gclk));
	jdff dff_A_bu5l24mo1_1(.dout(w_n1597_0[1]),.din(w_dff_A_bu5l24mo1_1),.clk(gclk));
	jdff dff_B_2qDZexht2_2(.din(n1597),.dout(w_dff_B_2qDZexht2_2),.clk(gclk));
	jdff dff_B_wFidWInp6_0(.din(n1596),.dout(w_dff_B_wFidWInp6_0),.clk(gclk));
	jdff dff_B_2hPWlplO9_0(.din(n1595),.dout(w_dff_B_2hPWlplO9_0),.clk(gclk));
	jdff dff_B_BZvg9vHT9_0(.din(w_dff_B_2hPWlplO9_0),.dout(w_dff_B_BZvg9vHT9_0),.clk(gclk));
	jdff dff_B_kzPwRbqB8_0(.din(w_dff_B_BZvg9vHT9_0),.dout(w_dff_B_kzPwRbqB8_0),.clk(gclk));
	jdff dff_B_veFixvxm7_0(.din(n1592),.dout(w_dff_B_veFixvxm7_0),.clk(gclk));
	jdff dff_A_xbYiXmtF2_1(.dout(w_n1106_0[1]),.din(w_dff_A_xbYiXmtF2_1),.clk(gclk));
	jdff dff_A_TjyU1OXs3_1(.dout(w_dff_A_xbYiXmtF2_1),.din(w_dff_A_TjyU1OXs3_1),.clk(gclk));
	jdff dff_A_oB7sxDnQ9_1(.dout(w_dff_A_TjyU1OXs3_1),.din(w_dff_A_oB7sxDnQ9_1),.clk(gclk));
	jdff dff_A_8sBd1jj22_1(.dout(w_dff_A_oB7sxDnQ9_1),.din(w_dff_A_8sBd1jj22_1),.clk(gclk));
	jdff dff_A_ZXN5ixdo4_1(.dout(w_dff_A_8sBd1jj22_1),.din(w_dff_A_ZXN5ixdo4_1),.clk(gclk));
	jdff dff_A_BWNUhscW4_1(.dout(w_dff_A_ZXN5ixdo4_1),.din(w_dff_A_BWNUhscW4_1),.clk(gclk));
	jdff dff_A_LXIdQTAd3_1(.dout(w_dff_A_BWNUhscW4_1),.din(w_dff_A_LXIdQTAd3_1),.clk(gclk));
	jdff dff_A_DhEd4Yhf6_1(.dout(w_dff_A_LXIdQTAd3_1),.din(w_dff_A_DhEd4Yhf6_1),.clk(gclk));
	jdff dff_A_YPCb7Y197_1(.dout(w_dff_A_DhEd4Yhf6_1),.din(w_dff_A_YPCb7Y197_1),.clk(gclk));
	jdff dff_A_7QPIrrcj9_1(.dout(w_dff_A_YPCb7Y197_1),.din(w_dff_A_7QPIrrcj9_1),.clk(gclk));
	jdff dff_A_i5KSLdrG3_1(.dout(w_n619_0[1]),.din(w_dff_A_i5KSLdrG3_1),.clk(gclk));
	jdff dff_A_sSgBY74Z6_1(.dout(w_dff_A_i5KSLdrG3_1),.din(w_dff_A_sSgBY74Z6_1),.clk(gclk));
	jdff dff_A_hoDPsrQ82_1(.dout(w_dff_A_sSgBY74Z6_1),.din(w_dff_A_hoDPsrQ82_1),.clk(gclk));
	jdff dff_A_tp6F6lUs4_1(.dout(w_dff_A_hoDPsrQ82_1),.din(w_dff_A_tp6F6lUs4_1),.clk(gclk));
	jdff dff_A_nT099fAz5_1(.dout(w_dff_A_tp6F6lUs4_1),.din(w_dff_A_nT099fAz5_1),.clk(gclk));
	jdff dff_B_eZX0uqCU7_1(.din(n607),.dout(w_dff_B_eZX0uqCU7_1),.clk(gclk));
	jdff dff_B_ZbK3sXt04_1(.din(w_dff_B_eZX0uqCU7_1),.dout(w_dff_B_ZbK3sXt04_1),.clk(gclk));
	jdff dff_A_XiAuJxIm0_0(.dout(w_n618_0[0]),.din(w_dff_A_XiAuJxIm0_0),.clk(gclk));
	jdff dff_A_y5kFTxXt5_0(.dout(w_dff_A_XiAuJxIm0_0),.din(w_dff_A_y5kFTxXt5_0),.clk(gclk));
	jdff dff_A_FxK24AHN5_0(.dout(w_dff_A_y5kFTxXt5_0),.din(w_dff_A_FxK24AHN5_0),.clk(gclk));
	jdff dff_A_6EreClJn7_0(.dout(w_dff_A_FxK24AHN5_0),.din(w_dff_A_6EreClJn7_0),.clk(gclk));
	jdff dff_A_Kz2uNPy41_0(.dout(w_dff_A_6EreClJn7_0),.din(w_dff_A_Kz2uNPy41_0),.clk(gclk));
	jdff dff_B_0UPOrKaP0_1(.din(n611),.dout(w_dff_B_0UPOrKaP0_1),.clk(gclk));
	jdff dff_B_hy0ml6fJ9_1(.din(w_dff_B_0UPOrKaP0_1),.dout(w_dff_B_hy0ml6fJ9_1),.clk(gclk));
	jdff dff_A_eBmxvIUd3_0(.dout(w_n605_0[0]),.din(w_dff_A_eBmxvIUd3_0),.clk(gclk));
	jdff dff_A_VLtttGbJ4_0(.dout(w_dff_A_eBmxvIUd3_0),.din(w_dff_A_VLtttGbJ4_0),.clk(gclk));
	jdff dff_A_mzrBUT0E4_1(.dout(w_n605_0[1]),.din(w_dff_A_mzrBUT0E4_1),.clk(gclk));
	jdff dff_A_9XOtSCNm2_1(.dout(w_dff_A_mzrBUT0E4_1),.din(w_dff_A_9XOtSCNm2_1),.clk(gclk));
	jdff dff_A_njp2cFh33_1(.dout(w_dff_A_9XOtSCNm2_1),.din(w_dff_A_njp2cFh33_1),.clk(gclk));
	jdff dff_A_0PcztyWg5_1(.dout(w_dff_A_njp2cFh33_1),.din(w_dff_A_0PcztyWg5_1),.clk(gclk));
	jdff dff_A_AX8YAVEV9_1(.dout(w_dff_A_0PcztyWg5_1),.din(w_dff_A_AX8YAVEV9_1),.clk(gclk));
	jdff dff_A_QO3Ew3Hl7_1(.dout(w_dff_A_AX8YAVEV9_1),.din(w_dff_A_QO3Ew3Hl7_1),.clk(gclk));
	jdff dff_A_qsGsNXAh3_1(.dout(w_dff_A_QO3Ew3Hl7_1),.din(w_dff_A_qsGsNXAh3_1),.clk(gclk));
	jdff dff_A_n6YmIM1H6_1(.dout(w_dff_A_qsGsNXAh3_1),.din(w_dff_A_n6YmIM1H6_1),.clk(gclk));
	jdff dff_A_lUsHpICq5_1(.dout(w_dff_A_n6YmIM1H6_1),.din(w_dff_A_lUsHpICq5_1),.clk(gclk));
	jdff dff_A_C2x1klrX5_0(.dout(w_n604_0[0]),.din(w_dff_A_C2x1klrX5_0),.clk(gclk));
	jdff dff_A_rMM9sWQL4_0(.dout(w_dff_A_C2x1klrX5_0),.din(w_dff_A_rMM9sWQL4_0),.clk(gclk));
	jdff dff_A_3b07Xonv3_0(.dout(w_dff_A_rMM9sWQL4_0),.din(w_dff_A_3b07Xonv3_0),.clk(gclk));
	jdff dff_A_MqzgzvAT4_0(.dout(w_dff_A_3b07Xonv3_0),.din(w_dff_A_MqzgzvAT4_0),.clk(gclk));
	jdff dff_A_WYCJ9KX06_0(.dout(w_dff_A_MqzgzvAT4_0),.din(w_dff_A_WYCJ9KX06_0),.clk(gclk));
	jdff dff_A_GzP3BLua7_0(.dout(w_dff_A_WYCJ9KX06_0),.din(w_dff_A_GzP3BLua7_0),.clk(gclk));
	jdff dff_A_tKkvh8lj4_0(.dout(w_dff_A_GzP3BLua7_0),.din(w_dff_A_tKkvh8lj4_0),.clk(gclk));
	jdff dff_A_v394gfxm8_0(.dout(w_dff_A_tKkvh8lj4_0),.din(w_dff_A_v394gfxm8_0),.clk(gclk));
	jdff dff_A_EusGPNz78_0(.dout(w_dff_A_v394gfxm8_0),.din(w_dff_A_EusGPNz78_0),.clk(gclk));
	jdff dff_A_fpwKEp9r3_0(.dout(w_dff_A_EusGPNz78_0),.din(w_dff_A_fpwKEp9r3_0),.clk(gclk));
	jdff dff_A_MqdtD7bv8_1(.dout(w_n594_0[1]),.din(w_dff_A_MqdtD7bv8_1),.clk(gclk));
	jdff dff_A_HL4xyrhO9_1(.dout(w_dff_A_MqdtD7bv8_1),.din(w_dff_A_HL4xyrhO9_1),.clk(gclk));
	jdff dff_A_am7P2UTf1_1(.dout(w_dff_A_HL4xyrhO9_1),.din(w_dff_A_am7P2UTf1_1),.clk(gclk));
	jdff dff_A_3ZRPYQxP9_1(.dout(w_dff_A_am7P2UTf1_1),.din(w_dff_A_3ZRPYQxP9_1),.clk(gclk));
	jdff dff_A_2l3z9mCJ6_1(.dout(w_dff_A_3ZRPYQxP9_1),.din(w_dff_A_2l3z9mCJ6_1),.clk(gclk));
	jdff dff_A_zcN8Ytqm3_1(.dout(w_dff_A_2l3z9mCJ6_1),.din(w_dff_A_zcN8Ytqm3_1),.clk(gclk));
	jdff dff_A_ZeXlIfVU6_1(.dout(w_dff_A_zcN8Ytqm3_1),.din(w_dff_A_ZeXlIfVU6_1),.clk(gclk));
	jdff dff_A_IYz19oPn3_1(.dout(w_dff_A_ZeXlIfVU6_1),.din(w_dff_A_IYz19oPn3_1),.clk(gclk));
	jdff dff_A_OCLlUMon3_1(.dout(w_dff_A_IYz19oPn3_1),.din(w_dff_A_OCLlUMon3_1),.clk(gclk));
	jdff dff_A_OziQOkLQ4_1(.dout(w_dff_A_OCLlUMon3_1),.din(w_dff_A_OziQOkLQ4_1),.clk(gclk));
	jdff dff_A_Xv9SHgSe6_1(.dout(w_dff_A_OziQOkLQ4_1),.din(w_dff_A_Xv9SHgSe6_1),.clk(gclk));
	jdff dff_A_hJkd0q0H7_1(.dout(w_dff_A_Xv9SHgSe6_1),.din(w_dff_A_hJkd0q0H7_1),.clk(gclk));
	jdff dff_A_uLJhR1De9_2(.dout(w_n594_0[2]),.din(w_dff_A_uLJhR1De9_2),.clk(gclk));
	jdff dff_B_bFXeCJWI1_1(.din(n650),.dout(w_dff_B_bFXeCJWI1_1),.clk(gclk));
	jdff dff_B_P2NvOeP18_1(.din(w_dff_B_bFXeCJWI1_1),.dout(w_dff_B_P2NvOeP18_1),.clk(gclk));
	jdff dff_B_SPEF7vWy2_1(.din(w_dff_B_P2NvOeP18_1),.dout(w_dff_B_SPEF7vWy2_1),.clk(gclk));
	jdff dff_B_C1GdZ4kY1_1(.din(w_dff_B_SPEF7vWy2_1),.dout(w_dff_B_C1GdZ4kY1_1),.clk(gclk));
	jdff dff_A_Bwd6QaoA3_0(.dout(w_n666_0[0]),.din(w_dff_A_Bwd6QaoA3_0),.clk(gclk));
	jdff dff_A_S7RxhA6h0_0(.dout(w_n664_0[0]),.din(w_dff_A_S7RxhA6h0_0),.clk(gclk));
	jdff dff_A_k4tZXlm27_0(.dout(w_dff_A_S7RxhA6h0_0),.din(w_dff_A_k4tZXlm27_0),.clk(gclk));
	jdff dff_B_okLIaUll6_2(.din(n664),.dout(w_dff_B_okLIaUll6_2),.clk(gclk));
	jdff dff_A_g3iSUOi77_1(.dout(w_n662_0[1]),.din(w_dff_A_g3iSUOi77_1),.clk(gclk));
	jdff dff_A_g47FT1Sz5_1(.dout(w_n661_0[1]),.din(w_dff_A_g47FT1Sz5_1),.clk(gclk));
	jdff dff_A_R2bpxslN8_1(.dout(w_dff_A_g47FT1Sz5_1),.din(w_dff_A_R2bpxslN8_1),.clk(gclk));
	jdff dff_A_fUruxAvU7_1(.dout(w_dff_A_R2bpxslN8_1),.din(w_dff_A_fUruxAvU7_1),.clk(gclk));
	jdff dff_A_lqYBdj6U0_2(.dout(w_n661_0[2]),.din(w_dff_A_lqYBdj6U0_2),.clk(gclk));
	jdff dff_B_QnNTBcV28_1(.din(n658),.dout(w_dff_B_QnNTBcV28_1),.clk(gclk));
	jdff dff_A_eMdK6NeO2_1(.dout(w_n657_0[1]),.din(w_dff_A_eMdK6NeO2_1),.clk(gclk));
	jdff dff_A_T6DH3wwq8_1(.dout(w_dff_A_eMdK6NeO2_1),.din(w_dff_A_T6DH3wwq8_1),.clk(gclk));
	jdff dff_A_KrLgufYI9_2(.dout(w_n657_0[2]),.din(w_dff_A_KrLgufYI9_2),.clk(gclk));
	jdff dff_A_mb2OTymV4_2(.dout(w_dff_A_KrLgufYI9_2),.din(w_dff_A_mb2OTymV4_2),.clk(gclk));
	jdff dff_A_SLcNwMxy7_0(.dout(w_n653_0[0]),.din(w_dff_A_SLcNwMxy7_0),.clk(gclk));
	jdff dff_A_lC4qb3jX0_0(.dout(w_dff_A_SLcNwMxy7_0),.din(w_dff_A_lC4qb3jX0_0),.clk(gclk));
	jdff dff_A_lZXB9Ylo4_0(.dout(w_dff_A_lC4qb3jX0_0),.din(w_dff_A_lZXB9Ylo4_0),.clk(gclk));
	jdff dff_B_9jMRwUAO9_2(.din(n653),.dout(w_dff_B_9jMRwUAO9_2),.clk(gclk));
	jdff dff_B_kPkQ15z64_2(.din(w_dff_B_9jMRwUAO9_2),.dout(w_dff_B_kPkQ15z64_2),.clk(gclk));
	jdff dff_B_kKtfS4rA8_2(.din(w_dff_B_kPkQ15z64_2),.dout(w_dff_B_kKtfS4rA8_2),.clk(gclk));
	jdff dff_A_jX290eNI2_0(.dout(w_n1094_0[0]),.din(w_dff_A_jX290eNI2_0),.clk(gclk));
	jdff dff_A_s8xnPzOq5_1(.dout(w_n1094_0[1]),.din(w_dff_A_s8xnPzOq5_1),.clk(gclk));
	jdff dff_A_SxvGIu5g6_1(.dout(w_dff_A_s8xnPzOq5_1),.din(w_dff_A_SxvGIu5g6_1),.clk(gclk));
	jdff dff_B_W9vLfPdA9_3(.din(n1094),.dout(w_dff_B_W9vLfPdA9_3),.clk(gclk));
	jdff dff_B_uwGCQ1Gp5_3(.din(w_dff_B_W9vLfPdA9_3),.dout(w_dff_B_uwGCQ1Gp5_3),.clk(gclk));
	jdff dff_B_RgcyJSHo2_3(.din(w_dff_B_uwGCQ1Gp5_3),.dout(w_dff_B_RgcyJSHo2_3),.clk(gclk));
	jdff dff_B_bzl0gWHi7_3(.din(w_dff_B_RgcyJSHo2_3),.dout(w_dff_B_bzl0gWHi7_3),.clk(gclk));
	jdff dff_B_yRq3ZuRu6_3(.din(w_dff_B_bzl0gWHi7_3),.dout(w_dff_B_yRq3ZuRu6_3),.clk(gclk));
	jdff dff_B_zJt5tn4C4_3(.din(w_dff_B_yRq3ZuRu6_3),.dout(w_dff_B_zJt5tn4C4_3),.clk(gclk));
	jdff dff_B_baY7IJcr3_3(.din(w_dff_B_zJt5tn4C4_3),.dout(w_dff_B_baY7IJcr3_3),.clk(gclk));
	jdff dff_B_GA7pTdUZ8_3(.din(w_dff_B_baY7IJcr3_3),.dout(w_dff_B_GA7pTdUZ8_3),.clk(gclk));
	jdff dff_B_T8FdJU7K8_3(.din(w_dff_B_GA7pTdUZ8_3),.dout(w_dff_B_T8FdJU7K8_3),.clk(gclk));
	jdff dff_B_5RF7sKrM0_3(.din(w_dff_B_T8FdJU7K8_3),.dout(w_dff_B_5RF7sKrM0_3),.clk(gclk));
	jdff dff_B_ldnKndYB2_3(.din(w_dff_B_5RF7sKrM0_3),.dout(w_dff_B_ldnKndYB2_3),.clk(gclk));
	jdff dff_A_F0MUBJYi3_0(.dout(w_G4526_1[0]),.din(w_dff_A_F0MUBJYi3_0),.clk(gclk));
	jdff dff_A_WzpvETxh7_0(.dout(w_dff_A_F0MUBJYi3_0),.din(w_dff_A_WzpvETxh7_0),.clk(gclk));
	jdff dff_A_NvDLcwJC7_0(.dout(w_dff_A_WzpvETxh7_0),.din(w_dff_A_NvDLcwJC7_0),.clk(gclk));
	jdff dff_A_6afAvTiA1_0(.dout(w_dff_A_NvDLcwJC7_0),.din(w_dff_A_6afAvTiA1_0),.clk(gclk));
	jdff dff_A_AWdn3BLB4_0(.dout(w_dff_A_6afAvTiA1_0),.din(w_dff_A_AWdn3BLB4_0),.clk(gclk));
	jdff dff_A_Avu9ZOkc3_0(.dout(w_dff_A_AWdn3BLB4_0),.din(w_dff_A_Avu9ZOkc3_0),.clk(gclk));
	jdff dff_A_0begA1fN1_0(.dout(w_dff_A_Avu9ZOkc3_0),.din(w_dff_A_0begA1fN1_0),.clk(gclk));
	jdff dff_A_ffGYkaM04_0(.dout(w_dff_A_0begA1fN1_0),.din(w_dff_A_ffGYkaM04_0),.clk(gclk));
	jdff dff_A_R7Bcrq286_0(.dout(w_dff_A_ffGYkaM04_0),.din(w_dff_A_R7Bcrq286_0),.clk(gclk));
	jdff dff_A_QsS64q9h6_0(.dout(w_dff_A_R7Bcrq286_0),.din(w_dff_A_QsS64q9h6_0),.clk(gclk));
	jdff dff_A_N02OklIP5_0(.dout(w_dff_A_QsS64q9h6_0),.din(w_dff_A_N02OklIP5_0),.clk(gclk));
	jdff dff_A_zFcb95415_0(.dout(w_dff_A_N02OklIP5_0),.din(w_dff_A_zFcb95415_0),.clk(gclk));
	jdff dff_A_D0l4WvQv4_0(.dout(w_dff_A_zFcb95415_0),.din(w_dff_A_D0l4WvQv4_0),.clk(gclk));
	jdff dff_A_ehAwgVB08_0(.dout(w_dff_A_D0l4WvQv4_0),.din(w_dff_A_ehAwgVB08_0),.clk(gclk));
	jdff dff_A_yBL0tugy4_2(.dout(w_G4526_1[2]),.din(w_dff_A_yBL0tugy4_2),.clk(gclk));
	jdff dff_A_gm1J99Qc7_2(.dout(w_dff_A_yBL0tugy4_2),.din(w_dff_A_gm1J99Qc7_2),.clk(gclk));
	jdff dff_A_HXkUXqia7_2(.dout(w_dff_A_gm1J99Qc7_2),.din(w_dff_A_HXkUXqia7_2),.clk(gclk));
	jdff dff_A_rFBNmaJz8_2(.dout(w_dff_A_HXkUXqia7_2),.din(w_dff_A_rFBNmaJz8_2),.clk(gclk));
	jdff dff_A_M7wVrncw9_2(.dout(w_dff_A_rFBNmaJz8_2),.din(w_dff_A_M7wVrncw9_2),.clk(gclk));
	jdff dff_A_G0fSlt6T2_1(.dout(w_G4526_0[1]),.din(w_dff_A_G0fSlt6T2_1),.clk(gclk));
	jdff dff_A_bXAyjwwu1_1(.dout(w_dff_A_G0fSlt6T2_1),.din(w_dff_A_bXAyjwwu1_1),.clk(gclk));
	jdff dff_A_Fw08xDqB0_1(.dout(w_dff_A_bXAyjwwu1_1),.din(w_dff_A_Fw08xDqB0_1),.clk(gclk));
	jdff dff_A_ehkbIuDh9_1(.dout(w_dff_A_Fw08xDqB0_1),.din(w_dff_A_ehkbIuDh9_1),.clk(gclk));
	jdff dff_A_pSxPcOGY3_1(.dout(w_dff_A_ehkbIuDh9_1),.din(w_dff_A_pSxPcOGY3_1),.clk(gclk));
	jdff dff_A_XCpN15Zn1_2(.dout(w_G4526_0[2]),.din(w_dff_A_XCpN15Zn1_2),.clk(gclk));
	jdff dff_A_3jDpRkMg1_2(.dout(w_dff_A_XCpN15Zn1_2),.din(w_dff_A_3jDpRkMg1_2),.clk(gclk));
	jdff dff_A_MmY3BLUr3_2(.dout(w_dff_A_3jDpRkMg1_2),.din(w_dff_A_MmY3BLUr3_2),.clk(gclk));
	jdff dff_A_uHvhsYT62_2(.dout(w_dff_A_MmY3BLUr3_2),.din(w_dff_A_uHvhsYT62_2),.clk(gclk));
	jdff dff_A_geXDWWpj9_2(.dout(w_dff_A_uHvhsYT62_2),.din(w_dff_A_geXDWWpj9_2),.clk(gclk));
	jdff dff_A_2cAierZb3_2(.dout(w_dff_A_geXDWWpj9_2),.din(w_dff_A_2cAierZb3_2),.clk(gclk));
	jdff dff_A_Jg55DGE26_2(.dout(w_dff_A_2cAierZb3_2),.din(w_dff_A_Jg55DGE26_2),.clk(gclk));
	jdff dff_A_lQlJXt8t3_2(.dout(w_dff_A_Jg55DGE26_2),.din(w_dff_A_lQlJXt8t3_2),.clk(gclk));
	jdff dff_A_RiQyqCRg9_2(.dout(w_dff_A_lQlJXt8t3_2),.din(w_dff_A_RiQyqCRg9_2),.clk(gclk));
	jdff dff_A_hphdq8121_2(.dout(w_dff_A_RiQyqCRg9_2),.din(w_dff_A_hphdq8121_2),.clk(gclk));
	jdff dff_A_qtSG9lwf5_2(.dout(w_dff_A_hphdq8121_2),.din(w_dff_A_qtSG9lwf5_2),.clk(gclk));
	jdff dff_A_XLa1vGuz1_2(.dout(w_dff_A_qtSG9lwf5_2),.din(w_dff_A_XLa1vGuz1_2),.clk(gclk));
	jdff dff_A_1RvgfV2T7_2(.dout(w_dff_A_XLa1vGuz1_2),.din(w_dff_A_1RvgfV2T7_2),.clk(gclk));
	jdff dff_B_cI4nzNZ88_0(.din(n1586),.dout(w_dff_B_cI4nzNZ88_0),.clk(gclk));
	jdff dff_B_L2qPwmGX6_0(.din(w_dff_B_cI4nzNZ88_0),.dout(w_dff_B_L2qPwmGX6_0),.clk(gclk));
	jdff dff_B_9P2eLogb0_1(.din(n1582),.dout(w_dff_B_9P2eLogb0_1),.clk(gclk));
	jdff dff_B_GtBINyod8_1(.din(w_dff_B_9P2eLogb0_1),.dout(w_dff_B_GtBINyod8_1),.clk(gclk));
	jdff dff_B_FekjwbPH0_0(.din(n1584),.dout(w_dff_B_FekjwbPH0_0),.clk(gclk));
	jdff dff_A_yC57tngl3_0(.dout(w_n610_0[0]),.din(w_dff_A_yC57tngl3_0),.clk(gclk));
	jdff dff_A_oEs2wZ5J3_0(.dout(w_dff_A_yC57tngl3_0),.din(w_dff_A_oEs2wZ5J3_0),.clk(gclk));
	jdff dff_A_zXTFClyW9_1(.dout(w_n590_0[1]),.din(w_dff_A_zXTFClyW9_1),.clk(gclk));
	jdff dff_A_ekkaAfHZ3_1(.dout(w_dff_A_zXTFClyW9_1),.din(w_dff_A_ekkaAfHZ3_1),.clk(gclk));
	jdff dff_A_MNZ06QkH1_2(.dout(w_n590_0[2]),.din(w_dff_A_MNZ06QkH1_2),.clk(gclk));
	jdff dff_A_LqdujMuD7_2(.dout(w_dff_A_MNZ06QkH1_2),.din(w_dff_A_LqdujMuD7_2),.clk(gclk));
	jdff dff_A_qWObL3q60_1(.dout(w_n615_0[1]),.din(w_dff_A_qWObL3q60_1),.clk(gclk));
	jdff dff_A_EC2x0mWa3_1(.dout(w_dff_A_qWObL3q60_1),.din(w_dff_A_EC2x0mWa3_1),.clk(gclk));
	jdff dff_A_xWPT1tlm4_1(.dout(w_dff_A_EC2x0mWa3_1),.din(w_dff_A_xWPT1tlm4_1),.clk(gclk));
	jdff dff_A_WmoD18nh9_1(.dout(w_dff_A_xWPT1tlm4_1),.din(w_dff_A_WmoD18nh9_1),.clk(gclk));
	jdff dff_A_UpOGuhrs6_1(.dout(w_dff_A_WmoD18nh9_1),.din(w_dff_A_UpOGuhrs6_1),.clk(gclk));
	jdff dff_A_OtXKASWw2_1(.dout(w_dff_A_UpOGuhrs6_1),.din(w_dff_A_OtXKASWw2_1),.clk(gclk));
	jdff dff_A_0OPGAQxC3_1(.dout(w_dff_A_OtXKASWw2_1),.din(w_dff_A_0OPGAQxC3_1),.clk(gclk));
	jdff dff_A_Ym2u3F2I1_1(.dout(w_dff_A_0OPGAQxC3_1),.din(w_dff_A_Ym2u3F2I1_1),.clk(gclk));
	jdff dff_A_QJDwRvtH6_1(.dout(w_dff_A_Ym2u3F2I1_1),.din(w_dff_A_QJDwRvtH6_1),.clk(gclk));
	jdff dff_B_txm5M3Xs0_2(.din(n600),.dout(w_dff_B_txm5M3Xs0_2),.clk(gclk));
	jdff dff_B_TNGCVpEa1_2(.din(w_dff_B_txm5M3Xs0_2),.dout(w_dff_B_TNGCVpEa1_2),.clk(gclk));
	jdff dff_A_wLnESNMi5_1(.dout(w_n612_0[1]),.din(w_dff_A_wLnESNMi5_1),.clk(gclk));
	jdff dff_A_f82UZDuO2_1(.dout(w_n609_0[1]),.din(w_dff_A_f82UZDuO2_1),.clk(gclk));
	jdff dff_B_0P5kGAq49_2(.din(n609),.dout(w_dff_B_0P5kGAq49_2),.clk(gclk));
	jdff dff_B_n6OpHj769_2(.din(w_dff_B_0P5kGAq49_2),.dout(w_dff_B_n6OpHj769_2),.clk(gclk));
	jdff dff_B_wfvo8goK1_1(.din(n591),.dout(w_dff_B_wfvo8goK1_1),.clk(gclk));
	jdff dff_B_s7RfLXDr5_0(.din(G124),.dout(w_dff_B_s7RfLXDr5_0),.clk(gclk));
	jdff dff_A_SUobC3IH6_1(.dout(w_G3743_0[1]),.din(w_dff_A_SUobC3IH6_1),.clk(gclk));
	jdff dff_A_DlWciL399_1(.dout(w_dff_A_SUobC3IH6_1),.din(w_dff_A_DlWciL399_1),.clk(gclk));
	jdff dff_A_v7RoWmpE5_1(.dout(w_dff_A_DlWciL399_1),.din(w_dff_A_v7RoWmpE5_1),.clk(gclk));
	jdff dff_A_h7Gae4JC6_1(.dout(w_dff_A_v7RoWmpE5_1),.din(w_dff_A_h7Gae4JC6_1),.clk(gclk));
	jdff dff_A_T2l5DZtf0_1(.dout(w_n1084_0[1]),.din(w_dff_A_T2l5DZtf0_1),.clk(gclk));
	jdff dff_A_ZWMNnxvV5_2(.dout(w_n1084_0[2]),.din(w_dff_A_ZWMNnxvV5_2),.clk(gclk));
	jdff dff_A_vKGARMXT5_2(.dout(w_dff_A_ZWMNnxvV5_2),.din(w_dff_A_vKGARMXT5_2),.clk(gclk));
	jdff dff_A_51wQeFao0_2(.dout(w_dff_A_vKGARMXT5_2),.din(w_dff_A_51wQeFao0_2),.clk(gclk));
	jdff dff_A_erKoI9zu3_2(.dout(w_dff_A_51wQeFao0_2),.din(w_dff_A_erKoI9zu3_2),.clk(gclk));
	jdff dff_A_27MsNwcw0_2(.dout(w_dff_A_erKoI9zu3_2),.din(w_dff_A_27MsNwcw0_2),.clk(gclk));
	jdff dff_A_8FAGhlia4_2(.dout(w_dff_A_27MsNwcw0_2),.din(w_dff_A_8FAGhlia4_2),.clk(gclk));
	jdff dff_A_9C1hqSRx7_2(.dout(w_dff_A_8FAGhlia4_2),.din(w_dff_A_9C1hqSRx7_2),.clk(gclk));
	jdff dff_A_GbsbaBAM0_2(.dout(w_dff_A_9C1hqSRx7_2),.din(w_dff_A_GbsbaBAM0_2),.clk(gclk));
	jdff dff_A_6BvlZLHM4_2(.dout(w_dff_A_GbsbaBAM0_2),.din(w_dff_A_6BvlZLHM4_2),.clk(gclk));
	jdff dff_A_3WkyXO8q5_2(.dout(w_dff_A_6BvlZLHM4_2),.din(w_dff_A_3WkyXO8q5_2),.clk(gclk));
	jdff dff_A_D6zaqLRz9_2(.dout(w_dff_A_3WkyXO8q5_2),.din(w_dff_A_D6zaqLRz9_2),.clk(gclk));
	jdff dff_A_9nPoXgzs7_2(.dout(w_dff_A_D6zaqLRz9_2),.din(w_dff_A_9nPoXgzs7_2),.clk(gclk));
	jdff dff_B_8cvNMGpq8_1(.din(n583),.dout(w_dff_B_8cvNMGpq8_1),.clk(gclk));
	jdff dff_B_M6rCd2HD1_0(.din(G100),.dout(w_dff_B_M6rCd2HD1_0),.clk(gclk));
	jdff dff_A_mz1xwCoR0_0(.dout(w_n582_0[0]),.din(w_dff_A_mz1xwCoR0_0),.clk(gclk));
	jdff dff_A_Tr8DNePw2_0(.dout(w_dff_A_mz1xwCoR0_0),.din(w_dff_A_Tr8DNePw2_0),.clk(gclk));
	jdff dff_A_W2sQknpv5_2(.dout(w_n582_0[2]),.din(w_dff_A_W2sQknpv5_2),.clk(gclk));
	jdff dff_A_fwUXfxUZ0_2(.dout(w_dff_A_W2sQknpv5_2),.din(w_dff_A_fwUXfxUZ0_2),.clk(gclk));
	jdff dff_A_DJ3DCg119_1(.dout(w_G3749_0[1]),.din(w_dff_A_DJ3DCg119_1),.clk(gclk));
	jdff dff_A_10wQNGWj8_1(.dout(w_dff_A_DJ3DCg119_1),.din(w_dff_A_10wQNGWj8_1),.clk(gclk));
	jdff dff_A_q9efD5AW6_1(.dout(w_dff_A_10wQNGWj8_1),.din(w_dff_A_q9efD5AW6_1),.clk(gclk));
	jdff dff_A_grsjDkSy3_1(.dout(w_dff_A_q9efD5AW6_1),.din(w_dff_A_grsjDkSy3_1),.clk(gclk));
	jdff dff_A_CpakcBnU6_1(.dout(w_n1108_0[1]),.din(w_dff_A_CpakcBnU6_1),.clk(gclk));
	jdff dff_A_4WvY5A2k1_1(.dout(w_dff_A_CpakcBnU6_1),.din(w_dff_A_4WvY5A2k1_1),.clk(gclk));
	jdff dff_A_2PIS5woK2_1(.dout(w_dff_A_4WvY5A2k1_1),.din(w_dff_A_2PIS5woK2_1),.clk(gclk));
	jdff dff_A_vwftn3eC3_1(.dout(w_dff_A_2PIS5woK2_1),.din(w_dff_A_vwftn3eC3_1),.clk(gclk));
	jdff dff_A_3dPNGlx54_1(.dout(w_dff_A_vwftn3eC3_1),.din(w_dff_A_3dPNGlx54_1),.clk(gclk));
	jdff dff_A_z9Is80aF2_1(.dout(w_dff_A_3dPNGlx54_1),.din(w_dff_A_z9Is80aF2_1),.clk(gclk));
	jdff dff_A_vMJgKACb1_1(.dout(w_dff_A_z9Is80aF2_1),.din(w_dff_A_vMJgKACb1_1),.clk(gclk));
	jdff dff_A_cQUJLcfI9_1(.dout(w_dff_A_vMJgKACb1_1),.din(w_dff_A_cQUJLcfI9_1),.clk(gclk));
	jdff dff_A_dju4lfQv3_1(.dout(w_dff_A_cQUJLcfI9_1),.din(w_dff_A_dju4lfQv3_1),.clk(gclk));
	jdff dff_B_a2pNsB9Y1_1(.din(n601),.dout(w_dff_B_a2pNsB9Y1_1),.clk(gclk));
	jdff dff_B_7QV1unCt1_0(.din(G130),.dout(w_dff_B_7QV1unCt1_0),.clk(gclk));
	jdff dff_A_bNwzzcrN2_2(.dout(w_G3729_0[2]),.din(w_dff_A_bNwzzcrN2_2),.clk(gclk));
	jdff dff_A_C8AfzeSp8_2(.dout(w_dff_A_bNwzzcrN2_2),.din(w_dff_A_C8AfzeSp8_2),.clk(gclk));
	jdff dff_A_kepke5qS6_2(.dout(w_dff_A_C8AfzeSp8_2),.din(w_dff_A_kepke5qS6_2),.clk(gclk));
	jdff dff_A_d6USlwJ36_2(.dout(w_dff_A_kepke5qS6_2),.din(w_dff_A_d6USlwJ36_2),.clk(gclk));
	jdff dff_A_DB2Wrj6J1_1(.dout(w_n1105_0[1]),.din(w_dff_A_DB2Wrj6J1_1),.clk(gclk));
	jdff dff_A_Olvsr9NF6_1(.dout(w_dff_A_DB2Wrj6J1_1),.din(w_dff_A_Olvsr9NF6_1),.clk(gclk));
	jdff dff_A_RWSabYOR2_1(.dout(w_dff_A_Olvsr9NF6_1),.din(w_dff_A_RWSabYOR2_1),.clk(gclk));
	jdff dff_A_0St775YA1_1(.dout(w_dff_A_RWSabYOR2_1),.din(w_dff_A_0St775YA1_1),.clk(gclk));
	jdff dff_A_IM7OfCDf7_1(.dout(w_dff_A_0St775YA1_1),.din(w_dff_A_IM7OfCDf7_1),.clk(gclk));
	jdff dff_A_AaWoBz0U8_1(.dout(w_dff_A_IM7OfCDf7_1),.din(w_dff_A_AaWoBz0U8_1),.clk(gclk));
	jdff dff_A_eRNhunRI9_1(.dout(w_dff_A_AaWoBz0U8_1),.din(w_dff_A_eRNhunRI9_1),.clk(gclk));
	jdff dff_A_4qWlNzCh6_1(.dout(w_dff_A_eRNhunRI9_1),.din(w_dff_A_4qWlNzCh6_1),.clk(gclk));
	jdff dff_A_qjV563ti3_1(.dout(w_dff_A_4qWlNzCh6_1),.din(w_dff_A_qjV563ti3_1),.clk(gclk));
	jdff dff_A_0FiDF4Wn0_1(.dout(w_dff_A_qjV563ti3_1),.din(w_dff_A_0FiDF4Wn0_1),.clk(gclk));
	jdff dff_B_50ilp20S7_2(.din(n1105),.dout(w_dff_B_50ilp20S7_2),.clk(gclk));
	jdff dff_B_xjUMoG9V3_1(.din(n596),.dout(w_dff_B_xjUMoG9V3_1),.clk(gclk));
	jdff dff_B_fE0qDrAB4_0(.din(G127),.dout(w_dff_B_fE0qDrAB4_0),.clk(gclk));
	jdff dff_A_lQ3831J44_1(.dout(w_n595_0[1]),.din(w_dff_A_lQ3831J44_1),.clk(gclk));
	jdff dff_A_JBmjHym93_1(.dout(w_dff_A_lQ3831J44_1),.din(w_dff_A_JBmjHym93_1),.clk(gclk));
	jdff dff_A_97Q6vCgf6_2(.dout(w_n595_0[2]),.din(w_dff_A_97Q6vCgf6_2),.clk(gclk));
	jdff dff_A_lw13vdjv0_2(.dout(w_dff_A_97Q6vCgf6_2),.din(w_dff_A_lw13vdjv0_2),.clk(gclk));
	jdff dff_A_m6ftOYds0_1(.dout(w_G3737_0[1]),.din(w_dff_A_m6ftOYds0_1),.clk(gclk));
	jdff dff_A_FTlmgWLO4_1(.dout(w_dff_A_m6ftOYds0_1),.din(w_dff_A_FTlmgWLO4_1),.clk(gclk));
	jdff dff_A_udDzy56d3_1(.dout(w_dff_A_FTlmgWLO4_1),.din(w_dff_A_udDzy56d3_1),.clk(gclk));
	jdff dff_A_5JKO9HUY8_1(.dout(w_dff_A_udDzy56d3_1),.din(w_dff_A_5JKO9HUY8_1),.clk(gclk));
	jdff dff_B_L7ehRztw8_1(.din(n1087),.dout(w_dff_B_L7ehRztw8_1),.clk(gclk));
	jdff dff_B_P7u6YAzT2_1(.din(w_dff_B_L7ehRztw8_1),.dout(w_dff_B_P7u6YAzT2_1),.clk(gclk));
	jdff dff_B_NtNfFnlQ6_1(.din(w_dff_B_P7u6YAzT2_1),.dout(w_dff_B_NtNfFnlQ6_1),.clk(gclk));
	jdff dff_B_FWwsQ1OX3_1(.din(w_dff_B_NtNfFnlQ6_1),.dout(w_dff_B_FWwsQ1OX3_1),.clk(gclk));
	jdff dff_B_7GV5nmRp3_1(.din(w_dff_B_FWwsQ1OX3_1),.dout(w_dff_B_7GV5nmRp3_1),.clk(gclk));
	jdff dff_B_APXEe3xc8_1(.din(w_dff_B_7GV5nmRp3_1),.dout(w_dff_B_APXEe3xc8_1),.clk(gclk));
	jdff dff_B_bb6ohPrX4_1(.din(n1088),.dout(w_dff_B_bb6ohPrX4_1),.clk(gclk));
	jdff dff_B_0ty9xCX39_1(.din(w_dff_B_bb6ohPrX4_1),.dout(w_dff_B_0ty9xCX39_1),.clk(gclk));
	jdff dff_B_C1fNn5vN1_1(.din(w_dff_B_0ty9xCX39_1),.dout(w_dff_B_C1fNn5vN1_1),.clk(gclk));
	jdff dff_B_PyqZRoxv3_1(.din(n1062),.dout(w_dff_B_PyqZRoxv3_1),.clk(gclk));
	jdff dff_B_8ReLGgYj4_1(.din(w_dff_B_PyqZRoxv3_1),.dout(w_dff_B_8ReLGgYj4_1),.clk(gclk));
	jdff dff_B_Dn49nIRW9_1(.din(n1063),.dout(w_dff_B_Dn49nIRW9_1),.clk(gclk));
	jdff dff_B_sYlCGmio9_1(.din(n1064),.dout(w_dff_B_sYlCGmio9_1),.clk(gclk));
	jdff dff_A_tVHP3ub39_1(.dout(w_n656_0[1]),.din(w_dff_A_tVHP3ub39_1),.clk(gclk));
	jdff dff_A_We4CQKko3_1(.dout(w_dff_A_tVHP3ub39_1),.din(w_dff_A_We4CQKko3_1),.clk(gclk));
	jdff dff_A_OLYZPrwD4_1(.dout(w_n655_0[1]),.din(w_dff_A_OLYZPrwD4_1),.clk(gclk));
	jdff dff_A_2MoRzi234_1(.dout(w_dff_A_OLYZPrwD4_1),.din(w_dff_A_2MoRzi234_1),.clk(gclk));
	jdff dff_A_pjFj03hC5_1(.dout(w_dff_A_2MoRzi234_1),.din(w_dff_A_pjFj03hC5_1),.clk(gclk));
	jdff dff_A_i2BNmNkV7_1(.dout(w_n654_0[1]),.din(w_dff_A_i2BNmNkV7_1),.clk(gclk));
	jdff dff_A_rkCiUCNi9_1(.dout(w_dff_A_i2BNmNkV7_1),.din(w_dff_A_rkCiUCNi9_1),.clk(gclk));
	jdff dff_A_jmIQUttQ0_1(.dout(w_dff_A_rkCiUCNi9_1),.din(w_dff_A_jmIQUttQ0_1),.clk(gclk));
	jdff dff_A_VAADDw1t6_1(.dout(w_dff_A_jmIQUttQ0_1),.din(w_dff_A_VAADDw1t6_1),.clk(gclk));
	jdff dff_A_4ffNxxmu7_1(.dout(w_dff_A_VAADDw1t6_1),.din(w_dff_A_4ffNxxmu7_1),.clk(gclk));
	jdff dff_A_o6MVf1uf5_1(.dout(w_dff_A_4ffNxxmu7_1),.din(w_dff_A_o6MVf1uf5_1),.clk(gclk));
	jdff dff_A_uPsZQYsd5_1(.dout(w_dff_A_o6MVf1uf5_1),.din(w_dff_A_uPsZQYsd5_1),.clk(gclk));
	jdff dff_A_wxbAMaeY6_2(.dout(w_n654_0[2]),.din(w_dff_A_wxbAMaeY6_2),.clk(gclk));
	jdff dff_A_u55ca3qf7_2(.dout(w_dff_A_wxbAMaeY6_2),.din(w_dff_A_u55ca3qf7_2),.clk(gclk));
	jdff dff_A_4V5MLa2f1_2(.dout(w_dff_A_u55ca3qf7_2),.din(w_dff_A_4V5MLa2f1_2),.clk(gclk));
	jdff dff_A_RzDvUsnI8_2(.dout(w_dff_A_4V5MLa2f1_2),.din(w_dff_A_RzDvUsnI8_2),.clk(gclk));
	jdff dff_A_wFuCSSMj3_0(.dout(w_n652_0[0]),.din(w_dff_A_wFuCSSMj3_0),.clk(gclk));
	jdff dff_A_1fbhWlmc2_0(.dout(w_dff_A_wFuCSSMj3_0),.din(w_dff_A_1fbhWlmc2_0),.clk(gclk));
	jdff dff_A_HIs4Qe9V0_0(.dout(w_dff_A_1fbhWlmc2_0),.din(w_dff_A_HIs4Qe9V0_0),.clk(gclk));
	jdff dff_A_QcjPCR3s1_0(.dout(w_dff_A_HIs4Qe9V0_0),.din(w_dff_A_QcjPCR3s1_0),.clk(gclk));
	jdff dff_A_eytVzZhE5_0(.dout(w_n649_0[0]),.din(w_dff_A_eytVzZhE5_0),.clk(gclk));
	jdff dff_A_TnK07E4D0_0(.dout(w_dff_A_eytVzZhE5_0),.din(w_dff_A_TnK07E4D0_0),.clk(gclk));
	jdff dff_A_Dnw5UdAG5_0(.dout(w_dff_A_TnK07E4D0_0),.din(w_dff_A_Dnw5UdAG5_0),.clk(gclk));
	jdff dff_A_l9F1dX233_0(.dout(w_dff_A_Dnw5UdAG5_0),.din(w_dff_A_l9F1dX233_0),.clk(gclk));
	jdff dff_A_CQBBE4km1_0(.dout(w_dff_A_l9F1dX233_0),.din(w_dff_A_CQBBE4km1_0),.clk(gclk));
	jdff dff_A_aUNklMmy4_1(.dout(w_n647_0[1]),.din(w_dff_A_aUNklMmy4_1),.clk(gclk));
	jdff dff_A_mnGL5ekG2_1(.dout(w_dff_A_aUNklMmy4_1),.din(w_dff_A_mnGL5ekG2_1),.clk(gclk));
	jdff dff_A_a31CDdwQ9_1(.dout(w_dff_A_mnGL5ekG2_1),.din(w_dff_A_a31CDdwQ9_1),.clk(gclk));
	jdff dff_A_tYeMHNTp3_1(.dout(w_dff_A_a31CDdwQ9_1),.din(w_dff_A_tYeMHNTp3_1),.clk(gclk));
	jdff dff_A_wdpgfduw9_1(.dout(w_dff_A_tYeMHNTp3_1),.din(w_dff_A_wdpgfduw9_1),.clk(gclk));
	jdff dff_A_dijHIl8Y2_1(.dout(w_dff_A_wdpgfduw9_1),.din(w_dff_A_dijHIl8Y2_1),.clk(gclk));
	jdff dff_A_u7CR8iOw3_1(.dout(w_dff_A_dijHIl8Y2_1),.din(w_dff_A_u7CR8iOw3_1),.clk(gclk));
	jdff dff_A_HwbULfST9_0(.dout(w_n1086_0[0]),.din(w_dff_A_HwbULfST9_0),.clk(gclk));
	jdff dff_B_rBPl433c7_2(.din(n1086),.dout(w_dff_B_rBPl433c7_2),.clk(gclk));
	jdff dff_B_IL6LlgCz6_2(.din(w_dff_B_rBPl433c7_2),.dout(w_dff_B_IL6LlgCz6_2),.clk(gclk));
	jdff dff_A_QSMjHyq86_1(.dout(w_n646_0[1]),.din(w_dff_A_QSMjHyq86_1),.clk(gclk));
	jdff dff_A_R5PM2Q5y9_1(.dout(w_dff_A_QSMjHyq86_1),.din(w_dff_A_R5PM2Q5y9_1),.clk(gclk));
	jdff dff_A_G23F854o3_1(.dout(w_dff_A_R5PM2Q5y9_1),.din(w_dff_A_G23F854o3_1),.clk(gclk));
	jdff dff_A_2MAJkVPS5_1(.dout(w_n642_0[1]),.din(w_dff_A_2MAJkVPS5_1),.clk(gclk));
	jdff dff_A_rNwQE5Az1_1(.dout(w_dff_A_2MAJkVPS5_1),.din(w_dff_A_rNwQE5Az1_1),.clk(gclk));
	jdff dff_B_iivay0ji0_3(.din(n642),.dout(w_dff_B_iivay0ji0_3),.clk(gclk));
	jdff dff_A_TcgSIRFV1_0(.dout(w_G29_0[0]),.din(w_dff_A_TcgSIRFV1_0),.clk(gclk));
	jdff dff_A_8kUJOeFo4_0(.dout(w_G3705_1[0]),.din(w_dff_A_8kUJOeFo4_0),.clk(gclk));
	jdff dff_A_EVwhCroP0_0(.dout(w_dff_A_8kUJOeFo4_0),.din(w_dff_A_EVwhCroP0_0),.clk(gclk));
	jdff dff_A_0ekPl5pE5_0(.dout(w_dff_A_EVwhCroP0_0),.din(w_dff_A_0ekPl5pE5_0),.clk(gclk));
	jdff dff_A_pk4VvjxV7_2(.dout(w_G3705_1[2]),.din(w_dff_A_pk4VvjxV7_2),.clk(gclk));
	jdff dff_A_8VRlv9Ky3_2(.dout(w_dff_A_pk4VvjxV7_2),.din(w_dff_A_8VRlv9Ky3_2),.clk(gclk));
	jdff dff_A_JJz8ZuTB3_2(.dout(w_dff_A_8VRlv9Ky3_2),.din(w_dff_A_JJz8ZuTB3_2),.clk(gclk));
	jdff dff_A_lEOyIBCx6_2(.dout(w_G3705_0[2]),.din(w_dff_A_lEOyIBCx6_2),.clk(gclk));
	jdff dff_A_JeMr8D3h9_2(.dout(w_dff_A_lEOyIBCx6_2),.din(w_dff_A_JeMr8D3h9_2),.clk(gclk));
	jdff dff_A_BtE9KoFR5_2(.dout(w_dff_A_JeMr8D3h9_2),.din(w_dff_A_BtE9KoFR5_2),.clk(gclk));
	jdff dff_A_GIscOO4y1_0(.dout(w_n357_0[0]),.din(w_dff_A_GIscOO4y1_0),.clk(gclk));
	jdff dff_A_AA1GIeGo7_0(.dout(w_dff_A_GIscOO4y1_0),.din(w_dff_A_AA1GIeGo7_0),.clk(gclk));
	jdff dff_A_6OPMGmh60_0(.dout(w_dff_A_AA1GIeGo7_0),.din(w_dff_A_6OPMGmh60_0),.clk(gclk));
	jdff dff_B_oEDRfFsY6_3(.din(n354),.dout(w_dff_B_oEDRfFsY6_3),.clk(gclk));
	jdff dff_A_lQtzHlbT7_0(.dout(w_G41_0[0]),.din(w_dff_A_lQtzHlbT7_0),.clk(gclk));
	jdff dff_A_8gH7ZCXd4_1(.dout(w_G3701_1[1]),.din(w_dff_A_8gH7ZCXd4_1),.clk(gclk));
	jdff dff_A_abmFYAEM6_0(.dout(w_G3701_0[0]),.din(w_dff_A_abmFYAEM6_0),.clk(gclk));
	jdff dff_A_OUvp96IM3_1(.dout(w_n636_0[1]),.din(w_dff_A_OUvp96IM3_1),.clk(gclk));
	jdff dff_A_hfbqRdsU0_1(.dout(w_dff_A_OUvp96IM3_1),.din(w_dff_A_hfbqRdsU0_1),.clk(gclk));
	jdff dff_A_4yJLPBI18_1(.dout(w_dff_A_hfbqRdsU0_1),.din(w_dff_A_4yJLPBI18_1),.clk(gclk));
	jdff dff_A_fMw4awqK4_1(.dout(w_dff_A_4yJLPBI18_1),.din(w_dff_A_fMw4awqK4_1),.clk(gclk));
	jdff dff_A_G5JbCDNA5_2(.dout(w_n636_0[2]),.din(w_dff_A_G5JbCDNA5_2),.clk(gclk));
	jdff dff_A_qhiPFY6g6_2(.dout(w_dff_A_G5JbCDNA5_2),.din(w_dff_A_qhiPFY6g6_2),.clk(gclk));
	jdff dff_B_1i2SLdk65_1(.din(n633),.dout(w_dff_B_1i2SLdk65_1),.clk(gclk));
	jdff dff_B_ELLLUtH34_0(.din(G26),.dout(w_dff_B_ELLLUtH34_0),.clk(gclk));
	jdff dff_A_jCHUc5Ti2_1(.dout(w_G18_42[1]),.din(w_dff_A_jCHUc5Ti2_1),.clk(gclk));
	jdff dff_A_k5oACphD2_0(.dout(w_n632_0[0]),.din(w_dff_A_k5oACphD2_0),.clk(gclk));
	jdff dff_A_xecZ0YzB1_0(.dout(w_dff_A_k5oACphD2_0),.din(w_dff_A_xecZ0YzB1_0),.clk(gclk));
	jdff dff_A_FIyIO9se7_2(.dout(w_n632_0[2]),.din(w_dff_A_FIyIO9se7_2),.clk(gclk));
	jdff dff_A_XWBOdunm4_2(.dout(w_dff_A_FIyIO9se7_2),.din(w_dff_A_XWBOdunm4_2),.clk(gclk));
	jdff dff_A_uabqrrnq4_1(.dout(w_n631_0[1]),.din(w_dff_A_uabqrrnq4_1),.clk(gclk));
	jdff dff_A_nAghyw0R2_1(.dout(w_dff_A_uabqrrnq4_1),.din(w_dff_A_nAghyw0R2_1),.clk(gclk));
	jdff dff_A_v1DPICNN5_1(.dout(w_dff_A_nAghyw0R2_1),.din(w_dff_A_v1DPICNN5_1),.clk(gclk));
	jdff dff_A_EBj3uFbd5_1(.dout(w_dff_A_v1DPICNN5_1),.din(w_dff_A_EBj3uFbd5_1),.clk(gclk));
	jdff dff_A_726Qwzzu5_1(.dout(w_dff_A_EBj3uFbd5_1),.din(w_dff_A_726Qwzzu5_1),.clk(gclk));
	jdff dff_A_4jEPWjE13_1(.dout(w_dff_A_726Qwzzu5_1),.din(w_dff_A_4jEPWjE13_1),.clk(gclk));
	jdff dff_A_WZmF5jrl7_1(.dout(w_dff_A_4jEPWjE13_1),.din(w_dff_A_WZmF5jrl7_1),.clk(gclk));
	jdff dff_A_ZCmzAjkn2_2(.dout(w_n631_0[2]),.din(w_dff_A_ZCmzAjkn2_2),.clk(gclk));
	jdff dff_A_1wCTM7hN2_2(.dout(w_dff_A_ZCmzAjkn2_2),.din(w_dff_A_1wCTM7hN2_2),.clk(gclk));
	jdff dff_A_LKOjZSAq4_2(.dout(w_dff_A_1wCTM7hN2_2),.din(w_dff_A_LKOjZSAq4_2),.clk(gclk));
	jdff dff_B_pxBIfhne4_1(.din(n628),.dout(w_dff_B_pxBIfhne4_1),.clk(gclk));
	jdff dff_B_q1q8bvml7_0(.din(G23),.dout(w_dff_B_q1q8bvml7_0),.clk(gclk));
	jdff dff_A_byP7oCMA1_1(.dout(w_n627_0[1]),.din(w_dff_A_byP7oCMA1_1),.clk(gclk));
	jdff dff_A_3QSoSmmK1_1(.dout(w_dff_A_byP7oCMA1_1),.din(w_dff_A_3QSoSmmK1_1),.clk(gclk));
	jdff dff_A_VAhCKBDb7_2(.dout(w_n627_0[2]),.din(w_dff_A_VAhCKBDb7_2),.clk(gclk));
	jdff dff_A_MQZwyx2v6_2(.dout(w_dff_A_VAhCKBDb7_2),.din(w_dff_A_MQZwyx2v6_2),.clk(gclk));
	jdff dff_A_rw8FVwEy8_1(.dout(w_G3717_0[1]),.din(w_dff_A_rw8FVwEy8_1),.clk(gclk));
	jdff dff_A_AhzntgmX8_1(.dout(w_dff_A_rw8FVwEy8_1),.din(w_dff_A_AhzntgmX8_1),.clk(gclk));
	jdff dff_A_HOmbI2og8_1(.dout(w_dff_A_AhzntgmX8_1),.din(w_dff_A_HOmbI2og8_1),.clk(gclk));
	jdff dff_A_ky1Zb9sY5_1(.dout(w_dff_A_HOmbI2og8_1),.din(w_dff_A_ky1Zb9sY5_1),.clk(gclk));
	jdff dff_A_Ifwq6ZIh7_0(.dout(w_n626_1[0]),.din(w_dff_A_Ifwq6ZIh7_0),.clk(gclk));
	jdff dff_A_NutrcOz82_0(.dout(w_dff_A_Ifwq6ZIh7_0),.din(w_dff_A_NutrcOz82_0),.clk(gclk));
	jdff dff_A_eVsK6hWb2_0(.dout(w_dff_A_NutrcOz82_0),.din(w_dff_A_eVsK6hWb2_0),.clk(gclk));
	jdff dff_A_XDICiVpS9_0(.dout(w_dff_A_eVsK6hWb2_0),.din(w_dff_A_XDICiVpS9_0),.clk(gclk));
	jdff dff_A_RoLXqBJa7_0(.dout(w_dff_A_XDICiVpS9_0),.din(w_dff_A_RoLXqBJa7_0),.clk(gclk));
	jdff dff_A_ZnXxb8QY4_0(.dout(w_n626_0[0]),.din(w_dff_A_ZnXxb8QY4_0),.clk(gclk));
	jdff dff_A_kpVQThfN9_0(.dout(w_dff_A_ZnXxb8QY4_0),.din(w_dff_A_kpVQThfN9_0),.clk(gclk));
	jdff dff_A_r2JoQ3I74_0(.dout(w_dff_A_kpVQThfN9_0),.din(w_dff_A_r2JoQ3I74_0),.clk(gclk));
	jdff dff_A_lEWmyDbc0_0(.dout(w_dff_A_r2JoQ3I74_0),.din(w_dff_A_lEWmyDbc0_0),.clk(gclk));
	jdff dff_A_pumRDhR26_1(.dout(w_n626_0[1]),.din(w_dff_A_pumRDhR26_1),.clk(gclk));
	jdff dff_A_KfabqNKi2_1(.dout(w_dff_A_pumRDhR26_1),.din(w_dff_A_KfabqNKi2_1),.clk(gclk));
	jdff dff_A_sWU4GC0H7_1(.dout(w_dff_A_KfabqNKi2_1),.din(w_dff_A_sWU4GC0H7_1),.clk(gclk));
	jdff dff_A_ZNiXlFuF1_1(.dout(w_dff_A_sWU4GC0H7_1),.din(w_dff_A_ZNiXlFuF1_1),.clk(gclk));
	jdff dff_B_9E1ofxPW9_1(.din(n623),.dout(w_dff_B_9E1ofxPW9_1),.clk(gclk));
	jdff dff_B_xFCehTzh4_0(.din(G103),.dout(w_dff_B_xFCehTzh4_0),.clk(gclk));
	jdff dff_A_9oWdtRfv0_2(.dout(w_G18_49[2]),.din(w_dff_A_9oWdtRfv0_2),.clk(gclk));
	jdff dff_A_ghbSHbT54_1(.dout(w_n622_0[1]),.din(w_dff_A_ghbSHbT54_1),.clk(gclk));
	jdff dff_A_6JY6j7Qz2_1(.dout(w_dff_A_ghbSHbT54_1),.din(w_dff_A_6JY6j7Qz2_1),.clk(gclk));
	jdff dff_A_nFnDtmKI9_2(.dout(w_n622_0[2]),.din(w_dff_A_nFnDtmKI9_2),.clk(gclk));
	jdff dff_A_f2nqb3SF5_2(.dout(w_dff_A_nFnDtmKI9_2),.din(w_dff_A_f2nqb3SF5_2),.clk(gclk));
	jdff dff_A_cxdFok9Y7_1(.dout(w_G3723_0[1]),.din(w_dff_A_cxdFok9Y7_1),.clk(gclk));
	jdff dff_A_K1Y39WDO9_1(.dout(w_dff_A_cxdFok9Y7_1),.din(w_dff_A_K1Y39WDO9_1),.clk(gclk));
	jdff dff_A_1mrJC09w4_1(.dout(w_dff_A_K1Y39WDO9_1),.din(w_dff_A_1mrJC09w4_1),.clk(gclk));
	jdff dff_A_EXeMCmjT5_1(.dout(w_dff_A_1mrJC09w4_1),.din(w_dff_A_EXeMCmjT5_1),.clk(gclk));
	jdff dff_A_22M6stkl3_1(.dout(w_dff_A_S4BFoTEg6_0),.din(w_dff_A_22M6stkl3_1),.clk(gclk));
	jdff dff_A_S4BFoTEg6_0(.dout(w_dff_A_cUjB2sxD9_0),.din(w_dff_A_S4BFoTEg6_0),.clk(gclk));
	jdff dff_A_cUjB2sxD9_0(.dout(w_dff_A_2FGcljJN8_0),.din(w_dff_A_cUjB2sxD9_0),.clk(gclk));
	jdff dff_A_2FGcljJN8_0(.dout(w_dff_A_Q0WvdquK7_0),.din(w_dff_A_2FGcljJN8_0),.clk(gclk));
	jdff dff_A_Q0WvdquK7_0(.dout(w_dff_A_WgqfywFy7_0),.din(w_dff_A_Q0WvdquK7_0),.clk(gclk));
	jdff dff_A_WgqfywFy7_0(.dout(w_dff_A_ooOM0ng85_0),.din(w_dff_A_WgqfywFy7_0),.clk(gclk));
	jdff dff_A_ooOM0ng85_0(.dout(w_dff_A_iG3EWeGa5_0),.din(w_dff_A_ooOM0ng85_0),.clk(gclk));
	jdff dff_A_iG3EWeGa5_0(.dout(w_dff_A_jshj2HiV8_0),.din(w_dff_A_iG3EWeGa5_0),.clk(gclk));
	jdff dff_A_jshj2HiV8_0(.dout(w_dff_A_tW6X4tx01_0),.din(w_dff_A_jshj2HiV8_0),.clk(gclk));
	jdff dff_A_tW6X4tx01_0(.dout(w_dff_A_J9C4wcfI8_0),.din(w_dff_A_tW6X4tx01_0),.clk(gclk));
	jdff dff_A_J9C4wcfI8_0(.dout(w_dff_A_qysSZoJr1_0),.din(w_dff_A_J9C4wcfI8_0),.clk(gclk));
	jdff dff_A_qysSZoJr1_0(.dout(w_dff_A_yU5Vka497_0),.din(w_dff_A_qysSZoJr1_0),.clk(gclk));
	jdff dff_A_yU5Vka497_0(.dout(w_dff_A_Ph4Tfi194_0),.din(w_dff_A_yU5Vka497_0),.clk(gclk));
	jdff dff_A_Ph4Tfi194_0(.dout(w_dff_A_5QfYp62S4_0),.din(w_dff_A_Ph4Tfi194_0),.clk(gclk));
	jdff dff_A_5QfYp62S4_0(.dout(w_dff_A_l4sKdUgq2_0),.din(w_dff_A_5QfYp62S4_0),.clk(gclk));
	jdff dff_A_l4sKdUgq2_0(.dout(w_dff_A_9kWW4kCv6_0),.din(w_dff_A_l4sKdUgq2_0),.clk(gclk));
	jdff dff_A_9kWW4kCv6_0(.dout(w_dff_A_8ALYuyfL6_0),.din(w_dff_A_9kWW4kCv6_0),.clk(gclk));
	jdff dff_A_8ALYuyfL6_0(.dout(w_dff_A_FAb7LJJY5_0),.din(w_dff_A_8ALYuyfL6_0),.clk(gclk));
	jdff dff_A_FAb7LJJY5_0(.dout(w_dff_A_Fv2hj1QM1_0),.din(w_dff_A_FAb7LJJY5_0),.clk(gclk));
	jdff dff_A_Fv2hj1QM1_0(.dout(w_dff_A_XKd3H5AC1_0),.din(w_dff_A_Fv2hj1QM1_0),.clk(gclk));
	jdff dff_A_XKd3H5AC1_0(.dout(w_dff_A_o5d3wDgu8_0),.din(w_dff_A_XKd3H5AC1_0),.clk(gclk));
	jdff dff_A_o5d3wDgu8_0(.dout(w_dff_A_zeVGAt1I0_0),.din(w_dff_A_o5d3wDgu8_0),.clk(gclk));
	jdff dff_A_zeVGAt1I0_0(.dout(w_dff_A_eXbbmxP21_0),.din(w_dff_A_zeVGAt1I0_0),.clk(gclk));
	jdff dff_A_eXbbmxP21_0(.dout(w_dff_A_RmA6BJyc6_0),.din(w_dff_A_eXbbmxP21_0),.clk(gclk));
	jdff dff_A_RmA6BJyc6_0(.dout(w_dff_A_hMn7lFQn0_0),.din(w_dff_A_RmA6BJyc6_0),.clk(gclk));
	jdff dff_A_hMn7lFQn0_0(.dout(w_dff_A_oaFdoqsV7_0),.din(w_dff_A_hMn7lFQn0_0),.clk(gclk));
	jdff dff_A_oaFdoqsV7_0(.dout(w_dff_A_LUm5Lnf42_0),.din(w_dff_A_oaFdoqsV7_0),.clk(gclk));
	jdff dff_A_LUm5Lnf42_0(.dout(w_dff_A_hXiG1aqj1_0),.din(w_dff_A_LUm5Lnf42_0),.clk(gclk));
	jdff dff_A_hXiG1aqj1_0(.dout(w_dff_A_amNfyYye3_0),.din(w_dff_A_hXiG1aqj1_0),.clk(gclk));
	jdff dff_A_amNfyYye3_0(.dout(w_dff_A_dySuGVcc0_0),.din(w_dff_A_amNfyYye3_0),.clk(gclk));
	jdff dff_A_dySuGVcc0_0(.dout(w_dff_A_ESk33UDh2_0),.din(w_dff_A_dySuGVcc0_0),.clk(gclk));
	jdff dff_A_ESk33UDh2_0(.dout(w_dff_A_HBJBjulU5_0),.din(w_dff_A_ESk33UDh2_0),.clk(gclk));
	jdff dff_A_HBJBjulU5_0(.dout(w_dff_A_wKp5vQlJ0_0),.din(w_dff_A_HBJBjulU5_0),.clk(gclk));
	jdff dff_A_wKp5vQlJ0_0(.dout(w_dff_A_TYsgP5zn3_0),.din(w_dff_A_wKp5vQlJ0_0),.clk(gclk));
	jdff dff_A_TYsgP5zn3_0(.dout(w_dff_A_J41lkMAy3_0),.din(w_dff_A_TYsgP5zn3_0),.clk(gclk));
	jdff dff_A_J41lkMAy3_0(.dout(w_dff_A_PgBZ7IZV6_0),.din(w_dff_A_J41lkMAy3_0),.clk(gclk));
	jdff dff_A_PgBZ7IZV6_0(.dout(w_dff_A_aowgxbNX0_0),.din(w_dff_A_PgBZ7IZV6_0),.clk(gclk));
	jdff dff_A_aowgxbNX0_0(.dout(w_dff_A_HVDuQ0YC1_0),.din(w_dff_A_aowgxbNX0_0),.clk(gclk));
	jdff dff_A_HVDuQ0YC1_0(.dout(G2),.din(w_dff_A_HVDuQ0YC1_0),.clk(gclk));
	jdff dff_A_FXX2zFPh3_1(.dout(w_dff_A_kb1Jqb6t5_0),.din(w_dff_A_FXX2zFPh3_1),.clk(gclk));
	jdff dff_A_kb1Jqb6t5_0(.dout(w_dff_A_ESnj91XR7_0),.din(w_dff_A_kb1Jqb6t5_0),.clk(gclk));
	jdff dff_A_ESnj91XR7_0(.dout(w_dff_A_uP4QCxyX4_0),.din(w_dff_A_ESnj91XR7_0),.clk(gclk));
	jdff dff_A_uP4QCxyX4_0(.dout(w_dff_A_96M8kcMJ0_0),.din(w_dff_A_uP4QCxyX4_0),.clk(gclk));
	jdff dff_A_96M8kcMJ0_0(.dout(w_dff_A_GVrsSbyC8_0),.din(w_dff_A_96M8kcMJ0_0),.clk(gclk));
	jdff dff_A_GVrsSbyC8_0(.dout(w_dff_A_Yvn67Gvx1_0),.din(w_dff_A_GVrsSbyC8_0),.clk(gclk));
	jdff dff_A_Yvn67Gvx1_0(.dout(w_dff_A_WAnU2WVe6_0),.din(w_dff_A_Yvn67Gvx1_0),.clk(gclk));
	jdff dff_A_WAnU2WVe6_0(.dout(w_dff_A_Ak3wK5Nx7_0),.din(w_dff_A_WAnU2WVe6_0),.clk(gclk));
	jdff dff_A_Ak3wK5Nx7_0(.dout(w_dff_A_wdjaViia8_0),.din(w_dff_A_Ak3wK5Nx7_0),.clk(gclk));
	jdff dff_A_wdjaViia8_0(.dout(w_dff_A_YdebARPe6_0),.din(w_dff_A_wdjaViia8_0),.clk(gclk));
	jdff dff_A_YdebARPe6_0(.dout(w_dff_A_Ca4iiYRE3_0),.din(w_dff_A_YdebARPe6_0),.clk(gclk));
	jdff dff_A_Ca4iiYRE3_0(.dout(w_dff_A_2bRzvp8s6_0),.din(w_dff_A_Ca4iiYRE3_0),.clk(gclk));
	jdff dff_A_2bRzvp8s6_0(.dout(w_dff_A_tDHIY1q45_0),.din(w_dff_A_2bRzvp8s6_0),.clk(gclk));
	jdff dff_A_tDHIY1q45_0(.dout(w_dff_A_Tki5cdCZ2_0),.din(w_dff_A_tDHIY1q45_0),.clk(gclk));
	jdff dff_A_Tki5cdCZ2_0(.dout(w_dff_A_8wxorWK81_0),.din(w_dff_A_Tki5cdCZ2_0),.clk(gclk));
	jdff dff_A_8wxorWK81_0(.dout(w_dff_A_BkjYdNYj3_0),.din(w_dff_A_8wxorWK81_0),.clk(gclk));
	jdff dff_A_BkjYdNYj3_0(.dout(w_dff_A_8VhYLVrL6_0),.din(w_dff_A_BkjYdNYj3_0),.clk(gclk));
	jdff dff_A_8VhYLVrL6_0(.dout(w_dff_A_pYU1CmHc1_0),.din(w_dff_A_8VhYLVrL6_0),.clk(gclk));
	jdff dff_A_pYU1CmHc1_0(.dout(w_dff_A_GWI359iE7_0),.din(w_dff_A_pYU1CmHc1_0),.clk(gclk));
	jdff dff_A_GWI359iE7_0(.dout(w_dff_A_1x7sEI0E9_0),.din(w_dff_A_GWI359iE7_0),.clk(gclk));
	jdff dff_A_1x7sEI0E9_0(.dout(w_dff_A_FuxWOYa01_0),.din(w_dff_A_1x7sEI0E9_0),.clk(gclk));
	jdff dff_A_FuxWOYa01_0(.dout(w_dff_A_bRszjOR23_0),.din(w_dff_A_FuxWOYa01_0),.clk(gclk));
	jdff dff_A_bRszjOR23_0(.dout(w_dff_A_bRuHXpf80_0),.din(w_dff_A_bRszjOR23_0),.clk(gclk));
	jdff dff_A_bRuHXpf80_0(.dout(w_dff_A_KpBloNhI2_0),.din(w_dff_A_bRuHXpf80_0),.clk(gclk));
	jdff dff_A_KpBloNhI2_0(.dout(w_dff_A_7PtS6bqi0_0),.din(w_dff_A_KpBloNhI2_0),.clk(gclk));
	jdff dff_A_7PtS6bqi0_0(.dout(w_dff_A_7t5sQ2k68_0),.din(w_dff_A_7PtS6bqi0_0),.clk(gclk));
	jdff dff_A_7t5sQ2k68_0(.dout(w_dff_A_ErKWJn080_0),.din(w_dff_A_7t5sQ2k68_0),.clk(gclk));
	jdff dff_A_ErKWJn080_0(.dout(w_dff_A_WgoReFDp1_0),.din(w_dff_A_ErKWJn080_0),.clk(gclk));
	jdff dff_A_WgoReFDp1_0(.dout(w_dff_A_qS46TXoT6_0),.din(w_dff_A_WgoReFDp1_0),.clk(gclk));
	jdff dff_A_qS46TXoT6_0(.dout(w_dff_A_gdDr2Rt98_0),.din(w_dff_A_qS46TXoT6_0),.clk(gclk));
	jdff dff_A_gdDr2Rt98_0(.dout(w_dff_A_Z8a0uKeH2_0),.din(w_dff_A_gdDr2Rt98_0),.clk(gclk));
	jdff dff_A_Z8a0uKeH2_0(.dout(w_dff_A_dKOU73DZ5_0),.din(w_dff_A_Z8a0uKeH2_0),.clk(gclk));
	jdff dff_A_dKOU73DZ5_0(.dout(w_dff_A_S0bU80Qj9_0),.din(w_dff_A_dKOU73DZ5_0),.clk(gclk));
	jdff dff_A_S0bU80Qj9_0(.dout(w_dff_A_0ouWjXHq3_0),.din(w_dff_A_S0bU80Qj9_0),.clk(gclk));
	jdff dff_A_0ouWjXHq3_0(.dout(w_dff_A_2asVuN543_0),.din(w_dff_A_0ouWjXHq3_0),.clk(gclk));
	jdff dff_A_2asVuN543_0(.dout(w_dff_A_VzLzMeMV6_0),.din(w_dff_A_2asVuN543_0),.clk(gclk));
	jdff dff_A_VzLzMeMV6_0(.dout(w_dff_A_pN6dqDnS3_0),.din(w_dff_A_VzLzMeMV6_0),.clk(gclk));
	jdff dff_A_pN6dqDnS3_0(.dout(w_dff_A_2rLl3HX90_0),.din(w_dff_A_pN6dqDnS3_0),.clk(gclk));
	jdff dff_A_2rLl3HX90_0(.dout(G3),.din(w_dff_A_2rLl3HX90_0),.clk(gclk));
	jdff dff_A_APRPgR7j9_1(.dout(w_dff_A_joyYYdNZ9_0),.din(w_dff_A_APRPgR7j9_1),.clk(gclk));
	jdff dff_A_joyYYdNZ9_0(.dout(w_dff_A_Jf93922w9_0),.din(w_dff_A_joyYYdNZ9_0),.clk(gclk));
	jdff dff_A_Jf93922w9_0(.dout(w_dff_A_Gr38YLUF1_0),.din(w_dff_A_Jf93922w9_0),.clk(gclk));
	jdff dff_A_Gr38YLUF1_0(.dout(w_dff_A_7f7gfzmx5_0),.din(w_dff_A_Gr38YLUF1_0),.clk(gclk));
	jdff dff_A_7f7gfzmx5_0(.dout(w_dff_A_9e0u9XDq2_0),.din(w_dff_A_7f7gfzmx5_0),.clk(gclk));
	jdff dff_A_9e0u9XDq2_0(.dout(w_dff_A_jxaGMBcM1_0),.din(w_dff_A_9e0u9XDq2_0),.clk(gclk));
	jdff dff_A_jxaGMBcM1_0(.dout(w_dff_A_A4CM5ywT6_0),.din(w_dff_A_jxaGMBcM1_0),.clk(gclk));
	jdff dff_A_A4CM5ywT6_0(.dout(w_dff_A_PeUX5KYj9_0),.din(w_dff_A_A4CM5ywT6_0),.clk(gclk));
	jdff dff_A_PeUX5KYj9_0(.dout(w_dff_A_1SIO7G3m7_0),.din(w_dff_A_PeUX5KYj9_0),.clk(gclk));
	jdff dff_A_1SIO7G3m7_0(.dout(w_dff_A_vseIl3hp2_0),.din(w_dff_A_1SIO7G3m7_0),.clk(gclk));
	jdff dff_A_vseIl3hp2_0(.dout(w_dff_A_cJ6w0haZ7_0),.din(w_dff_A_vseIl3hp2_0),.clk(gclk));
	jdff dff_A_cJ6w0haZ7_0(.dout(w_dff_A_NJQndC2a4_0),.din(w_dff_A_cJ6w0haZ7_0),.clk(gclk));
	jdff dff_A_NJQndC2a4_0(.dout(w_dff_A_TGfx6qn55_0),.din(w_dff_A_NJQndC2a4_0),.clk(gclk));
	jdff dff_A_TGfx6qn55_0(.dout(w_dff_A_lhQJjV5B4_0),.din(w_dff_A_TGfx6qn55_0),.clk(gclk));
	jdff dff_A_lhQJjV5B4_0(.dout(w_dff_A_t1E4pHzx1_0),.din(w_dff_A_lhQJjV5B4_0),.clk(gclk));
	jdff dff_A_t1E4pHzx1_0(.dout(w_dff_A_GCmU1yjW9_0),.din(w_dff_A_t1E4pHzx1_0),.clk(gclk));
	jdff dff_A_GCmU1yjW9_0(.dout(w_dff_A_4ePGndEy2_0),.din(w_dff_A_GCmU1yjW9_0),.clk(gclk));
	jdff dff_A_4ePGndEy2_0(.dout(w_dff_A_deH99ELa8_0),.din(w_dff_A_4ePGndEy2_0),.clk(gclk));
	jdff dff_A_deH99ELa8_0(.dout(w_dff_A_EhrpGzo54_0),.din(w_dff_A_deH99ELa8_0),.clk(gclk));
	jdff dff_A_EhrpGzo54_0(.dout(w_dff_A_Pb2Rtkhx1_0),.din(w_dff_A_EhrpGzo54_0),.clk(gclk));
	jdff dff_A_Pb2Rtkhx1_0(.dout(w_dff_A_hikMJNge3_0),.din(w_dff_A_Pb2Rtkhx1_0),.clk(gclk));
	jdff dff_A_hikMJNge3_0(.dout(w_dff_A_ReDCaeiz6_0),.din(w_dff_A_hikMJNge3_0),.clk(gclk));
	jdff dff_A_ReDCaeiz6_0(.dout(w_dff_A_rPRVe1h62_0),.din(w_dff_A_ReDCaeiz6_0),.clk(gclk));
	jdff dff_A_rPRVe1h62_0(.dout(w_dff_A_4zA1Yrov6_0),.din(w_dff_A_rPRVe1h62_0),.clk(gclk));
	jdff dff_A_4zA1Yrov6_0(.dout(w_dff_A_7SFxjS3U8_0),.din(w_dff_A_4zA1Yrov6_0),.clk(gclk));
	jdff dff_A_7SFxjS3U8_0(.dout(w_dff_A_atmgDZ0b6_0),.din(w_dff_A_7SFxjS3U8_0),.clk(gclk));
	jdff dff_A_atmgDZ0b6_0(.dout(w_dff_A_E5BsM33q3_0),.din(w_dff_A_atmgDZ0b6_0),.clk(gclk));
	jdff dff_A_E5BsM33q3_0(.dout(w_dff_A_jEDbpPey0_0),.din(w_dff_A_E5BsM33q3_0),.clk(gclk));
	jdff dff_A_jEDbpPey0_0(.dout(w_dff_A_LHPxXMxu9_0),.din(w_dff_A_jEDbpPey0_0),.clk(gclk));
	jdff dff_A_LHPxXMxu9_0(.dout(w_dff_A_HFeGHG6V1_0),.din(w_dff_A_LHPxXMxu9_0),.clk(gclk));
	jdff dff_A_HFeGHG6V1_0(.dout(w_dff_A_9ymznQRo8_0),.din(w_dff_A_HFeGHG6V1_0),.clk(gclk));
	jdff dff_A_9ymznQRo8_0(.dout(w_dff_A_VOfRLEwm1_0),.din(w_dff_A_9ymznQRo8_0),.clk(gclk));
	jdff dff_A_VOfRLEwm1_0(.dout(w_dff_A_FsAWgeSX1_0),.din(w_dff_A_VOfRLEwm1_0),.clk(gclk));
	jdff dff_A_FsAWgeSX1_0(.dout(w_dff_A_ruaAMZbA3_0),.din(w_dff_A_FsAWgeSX1_0),.clk(gclk));
	jdff dff_A_ruaAMZbA3_0(.dout(w_dff_A_yy8WFVP23_0),.din(w_dff_A_ruaAMZbA3_0),.clk(gclk));
	jdff dff_A_yy8WFVP23_0(.dout(w_dff_A_GLO2zFsA6_0),.din(w_dff_A_yy8WFVP23_0),.clk(gclk));
	jdff dff_A_GLO2zFsA6_0(.dout(w_dff_A_2DVGfjUz6_0),.din(w_dff_A_GLO2zFsA6_0),.clk(gclk));
	jdff dff_A_2DVGfjUz6_0(.dout(w_dff_A_Kpoxo9Ac0_0),.din(w_dff_A_2DVGfjUz6_0),.clk(gclk));
	jdff dff_A_Kpoxo9Ac0_0(.dout(G450),.din(w_dff_A_Kpoxo9Ac0_0),.clk(gclk));
	jdff dff_A_NJEEXzqd5_1(.dout(w_dff_A_pLDhAxMW8_0),.din(w_dff_A_NJEEXzqd5_1),.clk(gclk));
	jdff dff_A_pLDhAxMW8_0(.dout(w_dff_A_HrgcHspM1_0),.din(w_dff_A_pLDhAxMW8_0),.clk(gclk));
	jdff dff_A_HrgcHspM1_0(.dout(w_dff_A_vItZSYUu0_0),.din(w_dff_A_HrgcHspM1_0),.clk(gclk));
	jdff dff_A_vItZSYUu0_0(.dout(w_dff_A_C2s8FxDV2_0),.din(w_dff_A_vItZSYUu0_0),.clk(gclk));
	jdff dff_A_C2s8FxDV2_0(.dout(w_dff_A_50huoxlO8_0),.din(w_dff_A_C2s8FxDV2_0),.clk(gclk));
	jdff dff_A_50huoxlO8_0(.dout(w_dff_A_ymn8d7Ed9_0),.din(w_dff_A_50huoxlO8_0),.clk(gclk));
	jdff dff_A_ymn8d7Ed9_0(.dout(w_dff_A_N2s6VMqI2_0),.din(w_dff_A_ymn8d7Ed9_0),.clk(gclk));
	jdff dff_A_N2s6VMqI2_0(.dout(w_dff_A_4x2ySOQx5_0),.din(w_dff_A_N2s6VMqI2_0),.clk(gclk));
	jdff dff_A_4x2ySOQx5_0(.dout(w_dff_A_rJQDC5Ul8_0),.din(w_dff_A_4x2ySOQx5_0),.clk(gclk));
	jdff dff_A_rJQDC5Ul8_0(.dout(w_dff_A_lzE6P0r60_0),.din(w_dff_A_rJQDC5Ul8_0),.clk(gclk));
	jdff dff_A_lzE6P0r60_0(.dout(w_dff_A_Kvpt5Jz93_0),.din(w_dff_A_lzE6P0r60_0),.clk(gclk));
	jdff dff_A_Kvpt5Jz93_0(.dout(w_dff_A_rR3p43uK6_0),.din(w_dff_A_Kvpt5Jz93_0),.clk(gclk));
	jdff dff_A_rR3p43uK6_0(.dout(w_dff_A_qvSXeoiA3_0),.din(w_dff_A_rR3p43uK6_0),.clk(gclk));
	jdff dff_A_qvSXeoiA3_0(.dout(w_dff_A_EpUsK3Ox6_0),.din(w_dff_A_qvSXeoiA3_0),.clk(gclk));
	jdff dff_A_EpUsK3Ox6_0(.dout(w_dff_A_qIxks7bg9_0),.din(w_dff_A_EpUsK3Ox6_0),.clk(gclk));
	jdff dff_A_qIxks7bg9_0(.dout(w_dff_A_hw0WMDrl4_0),.din(w_dff_A_qIxks7bg9_0),.clk(gclk));
	jdff dff_A_hw0WMDrl4_0(.dout(w_dff_A_JMjM0Poi2_0),.din(w_dff_A_hw0WMDrl4_0),.clk(gclk));
	jdff dff_A_JMjM0Poi2_0(.dout(w_dff_A_1oOQQzJq1_0),.din(w_dff_A_JMjM0Poi2_0),.clk(gclk));
	jdff dff_A_1oOQQzJq1_0(.dout(w_dff_A_YYIfwsKE6_0),.din(w_dff_A_1oOQQzJq1_0),.clk(gclk));
	jdff dff_A_YYIfwsKE6_0(.dout(w_dff_A_7cCxsnQj9_0),.din(w_dff_A_YYIfwsKE6_0),.clk(gclk));
	jdff dff_A_7cCxsnQj9_0(.dout(w_dff_A_V0sMGLOD2_0),.din(w_dff_A_7cCxsnQj9_0),.clk(gclk));
	jdff dff_A_V0sMGLOD2_0(.dout(w_dff_A_JZ9MfmNk1_0),.din(w_dff_A_V0sMGLOD2_0),.clk(gclk));
	jdff dff_A_JZ9MfmNk1_0(.dout(w_dff_A_bLjutzPT2_0),.din(w_dff_A_JZ9MfmNk1_0),.clk(gclk));
	jdff dff_A_bLjutzPT2_0(.dout(w_dff_A_19OpLNiN2_0),.din(w_dff_A_bLjutzPT2_0),.clk(gclk));
	jdff dff_A_19OpLNiN2_0(.dout(w_dff_A_ozZ9DEEF6_0),.din(w_dff_A_19OpLNiN2_0),.clk(gclk));
	jdff dff_A_ozZ9DEEF6_0(.dout(w_dff_A_Nrvh4t3X0_0),.din(w_dff_A_ozZ9DEEF6_0),.clk(gclk));
	jdff dff_A_Nrvh4t3X0_0(.dout(w_dff_A_psu5GN3F5_0),.din(w_dff_A_Nrvh4t3X0_0),.clk(gclk));
	jdff dff_A_psu5GN3F5_0(.dout(w_dff_A_BMjsK2cp1_0),.din(w_dff_A_psu5GN3F5_0),.clk(gclk));
	jdff dff_A_BMjsK2cp1_0(.dout(w_dff_A_hFHxa1pX2_0),.din(w_dff_A_BMjsK2cp1_0),.clk(gclk));
	jdff dff_A_hFHxa1pX2_0(.dout(w_dff_A_swjjkuwg7_0),.din(w_dff_A_hFHxa1pX2_0),.clk(gclk));
	jdff dff_A_swjjkuwg7_0(.dout(w_dff_A_DPx1y6bV7_0),.din(w_dff_A_swjjkuwg7_0),.clk(gclk));
	jdff dff_A_DPx1y6bV7_0(.dout(w_dff_A_2gyv21uI6_0),.din(w_dff_A_DPx1y6bV7_0),.clk(gclk));
	jdff dff_A_2gyv21uI6_0(.dout(w_dff_A_TK11w9Mu1_0),.din(w_dff_A_2gyv21uI6_0),.clk(gclk));
	jdff dff_A_TK11w9Mu1_0(.dout(w_dff_A_UsPHTIis6_0),.din(w_dff_A_TK11w9Mu1_0),.clk(gclk));
	jdff dff_A_UsPHTIis6_0(.dout(w_dff_A_ePDkRL1W0_0),.din(w_dff_A_UsPHTIis6_0),.clk(gclk));
	jdff dff_A_ePDkRL1W0_0(.dout(w_dff_A_mM7rX9mh2_0),.din(w_dff_A_ePDkRL1W0_0),.clk(gclk));
	jdff dff_A_mM7rX9mh2_0(.dout(w_dff_A_lMMfu7Xz6_0),.din(w_dff_A_mM7rX9mh2_0),.clk(gclk));
	jdff dff_A_lMMfu7Xz6_0(.dout(w_dff_A_iLl64GnQ8_0),.din(w_dff_A_lMMfu7Xz6_0),.clk(gclk));
	jdff dff_A_iLl64GnQ8_0(.dout(G448),.din(w_dff_A_iLl64GnQ8_0),.clk(gclk));
	jdff dff_A_pjeMTmIZ9_1(.dout(w_dff_A_5VHOhAeF2_0),.din(w_dff_A_pjeMTmIZ9_1),.clk(gclk));
	jdff dff_A_5VHOhAeF2_0(.dout(w_dff_A_U9QzQQ9X1_0),.din(w_dff_A_5VHOhAeF2_0),.clk(gclk));
	jdff dff_A_U9QzQQ9X1_0(.dout(w_dff_A_VQFCUgMN2_0),.din(w_dff_A_U9QzQQ9X1_0),.clk(gclk));
	jdff dff_A_VQFCUgMN2_0(.dout(w_dff_A_zIT6kIx26_0),.din(w_dff_A_VQFCUgMN2_0),.clk(gclk));
	jdff dff_A_zIT6kIx26_0(.dout(w_dff_A_XMBCQbZP8_0),.din(w_dff_A_zIT6kIx26_0),.clk(gclk));
	jdff dff_A_XMBCQbZP8_0(.dout(w_dff_A_cr8nApi83_0),.din(w_dff_A_XMBCQbZP8_0),.clk(gclk));
	jdff dff_A_cr8nApi83_0(.dout(w_dff_A_HUnZAv1t8_0),.din(w_dff_A_cr8nApi83_0),.clk(gclk));
	jdff dff_A_HUnZAv1t8_0(.dout(w_dff_A_DS8rsTnH4_0),.din(w_dff_A_HUnZAv1t8_0),.clk(gclk));
	jdff dff_A_DS8rsTnH4_0(.dout(w_dff_A_RUxLkkNd4_0),.din(w_dff_A_DS8rsTnH4_0),.clk(gclk));
	jdff dff_A_RUxLkkNd4_0(.dout(w_dff_A_De5hgCDX4_0),.din(w_dff_A_RUxLkkNd4_0),.clk(gclk));
	jdff dff_A_De5hgCDX4_0(.dout(w_dff_A_VPO65Toq8_0),.din(w_dff_A_De5hgCDX4_0),.clk(gclk));
	jdff dff_A_VPO65Toq8_0(.dout(w_dff_A_KpwmRhmd8_0),.din(w_dff_A_VPO65Toq8_0),.clk(gclk));
	jdff dff_A_KpwmRhmd8_0(.dout(w_dff_A_HZKXD9XM7_0),.din(w_dff_A_KpwmRhmd8_0),.clk(gclk));
	jdff dff_A_HZKXD9XM7_0(.dout(w_dff_A_UpxB5qYb2_0),.din(w_dff_A_HZKXD9XM7_0),.clk(gclk));
	jdff dff_A_UpxB5qYb2_0(.dout(w_dff_A_hbYWN6iI1_0),.din(w_dff_A_UpxB5qYb2_0),.clk(gclk));
	jdff dff_A_hbYWN6iI1_0(.dout(w_dff_A_sulSAXgm5_0),.din(w_dff_A_hbYWN6iI1_0),.clk(gclk));
	jdff dff_A_sulSAXgm5_0(.dout(w_dff_A_TFdCJt3D0_0),.din(w_dff_A_sulSAXgm5_0),.clk(gclk));
	jdff dff_A_TFdCJt3D0_0(.dout(w_dff_A_aD0Xtqq53_0),.din(w_dff_A_TFdCJt3D0_0),.clk(gclk));
	jdff dff_A_aD0Xtqq53_0(.dout(w_dff_A_qXy8SuO81_0),.din(w_dff_A_aD0Xtqq53_0),.clk(gclk));
	jdff dff_A_qXy8SuO81_0(.dout(w_dff_A_N3PHSIqS1_0),.din(w_dff_A_qXy8SuO81_0),.clk(gclk));
	jdff dff_A_N3PHSIqS1_0(.dout(w_dff_A_sqfIr7R24_0),.din(w_dff_A_N3PHSIqS1_0),.clk(gclk));
	jdff dff_A_sqfIr7R24_0(.dout(w_dff_A_0fVAjGjA0_0),.din(w_dff_A_sqfIr7R24_0),.clk(gclk));
	jdff dff_A_0fVAjGjA0_0(.dout(w_dff_A_GE8rLY793_0),.din(w_dff_A_0fVAjGjA0_0),.clk(gclk));
	jdff dff_A_GE8rLY793_0(.dout(w_dff_A_NtiNDVCG5_0),.din(w_dff_A_GE8rLY793_0),.clk(gclk));
	jdff dff_A_NtiNDVCG5_0(.dout(w_dff_A_7xeFGeCz4_0),.din(w_dff_A_NtiNDVCG5_0),.clk(gclk));
	jdff dff_A_7xeFGeCz4_0(.dout(w_dff_A_eGcgMxIJ4_0),.din(w_dff_A_7xeFGeCz4_0),.clk(gclk));
	jdff dff_A_eGcgMxIJ4_0(.dout(w_dff_A_C5PEqtWi0_0),.din(w_dff_A_eGcgMxIJ4_0),.clk(gclk));
	jdff dff_A_C5PEqtWi0_0(.dout(w_dff_A_rxe9sFe13_0),.din(w_dff_A_C5PEqtWi0_0),.clk(gclk));
	jdff dff_A_rxe9sFe13_0(.dout(w_dff_A_XNvkBDgL3_0),.din(w_dff_A_rxe9sFe13_0),.clk(gclk));
	jdff dff_A_XNvkBDgL3_0(.dout(w_dff_A_IJNGve9L7_0),.din(w_dff_A_XNvkBDgL3_0),.clk(gclk));
	jdff dff_A_IJNGve9L7_0(.dout(w_dff_A_Nsd9QtNA2_0),.din(w_dff_A_IJNGve9L7_0),.clk(gclk));
	jdff dff_A_Nsd9QtNA2_0(.dout(w_dff_A_YaqgMtqt4_0),.din(w_dff_A_Nsd9QtNA2_0),.clk(gclk));
	jdff dff_A_YaqgMtqt4_0(.dout(w_dff_A_ieI7m9dX1_0),.din(w_dff_A_YaqgMtqt4_0),.clk(gclk));
	jdff dff_A_ieI7m9dX1_0(.dout(w_dff_A_YHyu4QRf7_0),.din(w_dff_A_ieI7m9dX1_0),.clk(gclk));
	jdff dff_A_YHyu4QRf7_0(.dout(w_dff_A_Rp9Mh0v21_0),.din(w_dff_A_YHyu4QRf7_0),.clk(gclk));
	jdff dff_A_Rp9Mh0v21_0(.dout(w_dff_A_tc341b1e3_0),.din(w_dff_A_Rp9Mh0v21_0),.clk(gclk));
	jdff dff_A_tc341b1e3_0(.dout(w_dff_A_H0i7A5Jk0_0),.din(w_dff_A_tc341b1e3_0),.clk(gclk));
	jdff dff_A_H0i7A5Jk0_0(.dout(w_dff_A_R6NsU4lJ8_0),.din(w_dff_A_H0i7A5Jk0_0),.clk(gclk));
	jdff dff_A_R6NsU4lJ8_0(.dout(G444),.din(w_dff_A_R6NsU4lJ8_0),.clk(gclk));
	jdff dff_A_wpKXgQFK7_1(.dout(w_dff_A_NRfkR5Rg5_0),.din(w_dff_A_wpKXgQFK7_1),.clk(gclk));
	jdff dff_A_NRfkR5Rg5_0(.dout(w_dff_A_aSrchFsx3_0),.din(w_dff_A_NRfkR5Rg5_0),.clk(gclk));
	jdff dff_A_aSrchFsx3_0(.dout(w_dff_A_1uZ6WErQ9_0),.din(w_dff_A_aSrchFsx3_0),.clk(gclk));
	jdff dff_A_1uZ6WErQ9_0(.dout(w_dff_A_T7iW3xuc1_0),.din(w_dff_A_1uZ6WErQ9_0),.clk(gclk));
	jdff dff_A_T7iW3xuc1_0(.dout(w_dff_A_MooRyZOh2_0),.din(w_dff_A_T7iW3xuc1_0),.clk(gclk));
	jdff dff_A_MooRyZOh2_0(.dout(w_dff_A_w5D30tJ44_0),.din(w_dff_A_MooRyZOh2_0),.clk(gclk));
	jdff dff_A_w5D30tJ44_0(.dout(w_dff_A_YJxLTvYM8_0),.din(w_dff_A_w5D30tJ44_0),.clk(gclk));
	jdff dff_A_YJxLTvYM8_0(.dout(w_dff_A_rSipwpsY5_0),.din(w_dff_A_YJxLTvYM8_0),.clk(gclk));
	jdff dff_A_rSipwpsY5_0(.dout(w_dff_A_ZBXtti1C9_0),.din(w_dff_A_rSipwpsY5_0),.clk(gclk));
	jdff dff_A_ZBXtti1C9_0(.dout(w_dff_A_MVqZHUEl9_0),.din(w_dff_A_ZBXtti1C9_0),.clk(gclk));
	jdff dff_A_MVqZHUEl9_0(.dout(w_dff_A_yI3eLD4U0_0),.din(w_dff_A_MVqZHUEl9_0),.clk(gclk));
	jdff dff_A_yI3eLD4U0_0(.dout(w_dff_A_S25IkXfV5_0),.din(w_dff_A_yI3eLD4U0_0),.clk(gclk));
	jdff dff_A_S25IkXfV5_0(.dout(w_dff_A_r3ahwtRx7_0),.din(w_dff_A_S25IkXfV5_0),.clk(gclk));
	jdff dff_A_r3ahwtRx7_0(.dout(w_dff_A_VsEkdvk80_0),.din(w_dff_A_r3ahwtRx7_0),.clk(gclk));
	jdff dff_A_VsEkdvk80_0(.dout(w_dff_A_BRkNOJsf7_0),.din(w_dff_A_VsEkdvk80_0),.clk(gclk));
	jdff dff_A_BRkNOJsf7_0(.dout(w_dff_A_iiKzEKlV2_0),.din(w_dff_A_BRkNOJsf7_0),.clk(gclk));
	jdff dff_A_iiKzEKlV2_0(.dout(w_dff_A_k9Irk9G35_0),.din(w_dff_A_iiKzEKlV2_0),.clk(gclk));
	jdff dff_A_k9Irk9G35_0(.dout(w_dff_A_jOe8RLtg7_0),.din(w_dff_A_k9Irk9G35_0),.clk(gclk));
	jdff dff_A_jOe8RLtg7_0(.dout(w_dff_A_V3hm9Lmh5_0),.din(w_dff_A_jOe8RLtg7_0),.clk(gclk));
	jdff dff_A_V3hm9Lmh5_0(.dout(w_dff_A_X8aFoeJu3_0),.din(w_dff_A_V3hm9Lmh5_0),.clk(gclk));
	jdff dff_A_X8aFoeJu3_0(.dout(w_dff_A_X9wJXq9V7_0),.din(w_dff_A_X8aFoeJu3_0),.clk(gclk));
	jdff dff_A_X9wJXq9V7_0(.dout(w_dff_A_9oMvkVNg9_0),.din(w_dff_A_X9wJXq9V7_0),.clk(gclk));
	jdff dff_A_9oMvkVNg9_0(.dout(w_dff_A_2weA3CNg6_0),.din(w_dff_A_9oMvkVNg9_0),.clk(gclk));
	jdff dff_A_2weA3CNg6_0(.dout(w_dff_A_9vnvz8Io1_0),.din(w_dff_A_2weA3CNg6_0),.clk(gclk));
	jdff dff_A_9vnvz8Io1_0(.dout(w_dff_A_oCtwRTgz3_0),.din(w_dff_A_9vnvz8Io1_0),.clk(gclk));
	jdff dff_A_oCtwRTgz3_0(.dout(w_dff_A_jG079AtQ9_0),.din(w_dff_A_oCtwRTgz3_0),.clk(gclk));
	jdff dff_A_jG079AtQ9_0(.dout(w_dff_A_LGRfUNvg7_0),.din(w_dff_A_jG079AtQ9_0),.clk(gclk));
	jdff dff_A_LGRfUNvg7_0(.dout(w_dff_A_S2o33HEF5_0),.din(w_dff_A_LGRfUNvg7_0),.clk(gclk));
	jdff dff_A_S2o33HEF5_0(.dout(w_dff_A_0vdKzqsL4_0),.din(w_dff_A_S2o33HEF5_0),.clk(gclk));
	jdff dff_A_0vdKzqsL4_0(.dout(w_dff_A_UtkowifO0_0),.din(w_dff_A_0vdKzqsL4_0),.clk(gclk));
	jdff dff_A_UtkowifO0_0(.dout(w_dff_A_8QSAcOa86_0),.din(w_dff_A_UtkowifO0_0),.clk(gclk));
	jdff dff_A_8QSAcOa86_0(.dout(w_dff_A_YMEXzMq00_0),.din(w_dff_A_8QSAcOa86_0),.clk(gclk));
	jdff dff_A_YMEXzMq00_0(.dout(w_dff_A_uHVHlb2t0_0),.din(w_dff_A_YMEXzMq00_0),.clk(gclk));
	jdff dff_A_uHVHlb2t0_0(.dout(w_dff_A_dxfDkiid8_0),.din(w_dff_A_uHVHlb2t0_0),.clk(gclk));
	jdff dff_A_dxfDkiid8_0(.dout(w_dff_A_WRg3cFNA0_0),.din(w_dff_A_dxfDkiid8_0),.clk(gclk));
	jdff dff_A_WRg3cFNA0_0(.dout(w_dff_A_mv9TeVLQ0_0),.din(w_dff_A_WRg3cFNA0_0),.clk(gclk));
	jdff dff_A_mv9TeVLQ0_0(.dout(w_dff_A_N4kyoXmk4_0),.din(w_dff_A_mv9TeVLQ0_0),.clk(gclk));
	jdff dff_A_N4kyoXmk4_0(.dout(w_dff_A_T5ewH2rZ8_0),.din(w_dff_A_N4kyoXmk4_0),.clk(gclk));
	jdff dff_A_T5ewH2rZ8_0(.dout(G442),.din(w_dff_A_T5ewH2rZ8_0),.clk(gclk));
	jdff dff_A_anzn7UR03_1(.dout(w_dff_A_v6uTtzOE0_0),.din(w_dff_A_anzn7UR03_1),.clk(gclk));
	jdff dff_A_v6uTtzOE0_0(.dout(w_dff_A_2eVirea68_0),.din(w_dff_A_v6uTtzOE0_0),.clk(gclk));
	jdff dff_A_2eVirea68_0(.dout(w_dff_A_OlmaOuYn5_0),.din(w_dff_A_2eVirea68_0),.clk(gclk));
	jdff dff_A_OlmaOuYn5_0(.dout(w_dff_A_adIBZ9nD8_0),.din(w_dff_A_OlmaOuYn5_0),.clk(gclk));
	jdff dff_A_adIBZ9nD8_0(.dout(w_dff_A_a8gVUd2g9_0),.din(w_dff_A_adIBZ9nD8_0),.clk(gclk));
	jdff dff_A_a8gVUd2g9_0(.dout(w_dff_A_39vzzhvZ8_0),.din(w_dff_A_a8gVUd2g9_0),.clk(gclk));
	jdff dff_A_39vzzhvZ8_0(.dout(w_dff_A_EQM940HP3_0),.din(w_dff_A_39vzzhvZ8_0),.clk(gclk));
	jdff dff_A_EQM940HP3_0(.dout(w_dff_A_FlIdlKtr1_0),.din(w_dff_A_EQM940HP3_0),.clk(gclk));
	jdff dff_A_FlIdlKtr1_0(.dout(w_dff_A_Ecx36kOV9_0),.din(w_dff_A_FlIdlKtr1_0),.clk(gclk));
	jdff dff_A_Ecx36kOV9_0(.dout(w_dff_A_2ENfJecH1_0),.din(w_dff_A_Ecx36kOV9_0),.clk(gclk));
	jdff dff_A_2ENfJecH1_0(.dout(w_dff_A_l6Op9T8j6_0),.din(w_dff_A_2ENfJecH1_0),.clk(gclk));
	jdff dff_A_l6Op9T8j6_0(.dout(w_dff_A_gZOGycUB6_0),.din(w_dff_A_l6Op9T8j6_0),.clk(gclk));
	jdff dff_A_gZOGycUB6_0(.dout(w_dff_A_wClD1ypr4_0),.din(w_dff_A_gZOGycUB6_0),.clk(gclk));
	jdff dff_A_wClD1ypr4_0(.dout(w_dff_A_FxuEfVco8_0),.din(w_dff_A_wClD1ypr4_0),.clk(gclk));
	jdff dff_A_FxuEfVco8_0(.dout(w_dff_A_oJZOEiA06_0),.din(w_dff_A_FxuEfVco8_0),.clk(gclk));
	jdff dff_A_oJZOEiA06_0(.dout(w_dff_A_HBxp9Q4m2_0),.din(w_dff_A_oJZOEiA06_0),.clk(gclk));
	jdff dff_A_HBxp9Q4m2_0(.dout(w_dff_A_FKBI3KL28_0),.din(w_dff_A_HBxp9Q4m2_0),.clk(gclk));
	jdff dff_A_FKBI3KL28_0(.dout(w_dff_A_uYj6YSfL4_0),.din(w_dff_A_FKBI3KL28_0),.clk(gclk));
	jdff dff_A_uYj6YSfL4_0(.dout(w_dff_A_QfirL6wC1_0),.din(w_dff_A_uYj6YSfL4_0),.clk(gclk));
	jdff dff_A_QfirL6wC1_0(.dout(w_dff_A_pibm4Z2y9_0),.din(w_dff_A_QfirL6wC1_0),.clk(gclk));
	jdff dff_A_pibm4Z2y9_0(.dout(w_dff_A_DLSmdPvn1_0),.din(w_dff_A_pibm4Z2y9_0),.clk(gclk));
	jdff dff_A_DLSmdPvn1_0(.dout(w_dff_A_0BWT3AG56_0),.din(w_dff_A_DLSmdPvn1_0),.clk(gclk));
	jdff dff_A_0BWT3AG56_0(.dout(w_dff_A_gd1pvYuj4_0),.din(w_dff_A_0BWT3AG56_0),.clk(gclk));
	jdff dff_A_gd1pvYuj4_0(.dout(w_dff_A_UDJaqCAE2_0),.din(w_dff_A_gd1pvYuj4_0),.clk(gclk));
	jdff dff_A_UDJaqCAE2_0(.dout(w_dff_A_tW2S6lpC2_0),.din(w_dff_A_UDJaqCAE2_0),.clk(gclk));
	jdff dff_A_tW2S6lpC2_0(.dout(w_dff_A_bGAxGVPH0_0),.din(w_dff_A_tW2S6lpC2_0),.clk(gclk));
	jdff dff_A_bGAxGVPH0_0(.dout(w_dff_A_3MM7oVWi2_0),.din(w_dff_A_bGAxGVPH0_0),.clk(gclk));
	jdff dff_A_3MM7oVWi2_0(.dout(w_dff_A_fF2TI0ro4_0),.din(w_dff_A_3MM7oVWi2_0),.clk(gclk));
	jdff dff_A_fF2TI0ro4_0(.dout(w_dff_A_1kksXPnv6_0),.din(w_dff_A_fF2TI0ro4_0),.clk(gclk));
	jdff dff_A_1kksXPnv6_0(.dout(w_dff_A_2N90lZmI6_0),.din(w_dff_A_1kksXPnv6_0),.clk(gclk));
	jdff dff_A_2N90lZmI6_0(.dout(w_dff_A_6CPn6VuH5_0),.din(w_dff_A_2N90lZmI6_0),.clk(gclk));
	jdff dff_A_6CPn6VuH5_0(.dout(w_dff_A_oKpCBGvs8_0),.din(w_dff_A_6CPn6VuH5_0),.clk(gclk));
	jdff dff_A_oKpCBGvs8_0(.dout(w_dff_A_prIP4twm0_0),.din(w_dff_A_oKpCBGvs8_0),.clk(gclk));
	jdff dff_A_prIP4twm0_0(.dout(w_dff_A_hXNc79B47_0),.din(w_dff_A_prIP4twm0_0),.clk(gclk));
	jdff dff_A_hXNc79B47_0(.dout(w_dff_A_mMTCwnvF9_0),.din(w_dff_A_hXNc79B47_0),.clk(gclk));
	jdff dff_A_mMTCwnvF9_0(.dout(w_dff_A_zRJ58SpW8_0),.din(w_dff_A_mMTCwnvF9_0),.clk(gclk));
	jdff dff_A_zRJ58SpW8_0(.dout(w_dff_A_emxznUEz5_0),.din(w_dff_A_zRJ58SpW8_0),.clk(gclk));
	jdff dff_A_emxznUEz5_0(.dout(w_dff_A_w4IbDKxW6_0),.din(w_dff_A_emxznUEz5_0),.clk(gclk));
	jdff dff_A_w4IbDKxW6_0(.dout(G440),.din(w_dff_A_w4IbDKxW6_0),.clk(gclk));
	jdff dff_A_SmHHSwBU9_1(.dout(w_dff_A_IllnQw2i3_0),.din(w_dff_A_SmHHSwBU9_1),.clk(gclk));
	jdff dff_A_IllnQw2i3_0(.dout(w_dff_A_MoIg7aE97_0),.din(w_dff_A_IllnQw2i3_0),.clk(gclk));
	jdff dff_A_MoIg7aE97_0(.dout(w_dff_A_RTuxeuop9_0),.din(w_dff_A_MoIg7aE97_0),.clk(gclk));
	jdff dff_A_RTuxeuop9_0(.dout(w_dff_A_cs9yoYxh6_0),.din(w_dff_A_RTuxeuop9_0),.clk(gclk));
	jdff dff_A_cs9yoYxh6_0(.dout(w_dff_A_9vD9Msxf3_0),.din(w_dff_A_cs9yoYxh6_0),.clk(gclk));
	jdff dff_A_9vD9Msxf3_0(.dout(w_dff_A_YE8pMHkq1_0),.din(w_dff_A_9vD9Msxf3_0),.clk(gclk));
	jdff dff_A_YE8pMHkq1_0(.dout(w_dff_A_vmCRhtlb3_0),.din(w_dff_A_YE8pMHkq1_0),.clk(gclk));
	jdff dff_A_vmCRhtlb3_0(.dout(w_dff_A_bksCjaE00_0),.din(w_dff_A_vmCRhtlb3_0),.clk(gclk));
	jdff dff_A_bksCjaE00_0(.dout(w_dff_A_8XGRIX9H7_0),.din(w_dff_A_bksCjaE00_0),.clk(gclk));
	jdff dff_A_8XGRIX9H7_0(.dout(w_dff_A_aDQZd3382_0),.din(w_dff_A_8XGRIX9H7_0),.clk(gclk));
	jdff dff_A_aDQZd3382_0(.dout(w_dff_A_8Y9VSXqN9_0),.din(w_dff_A_aDQZd3382_0),.clk(gclk));
	jdff dff_A_8Y9VSXqN9_0(.dout(w_dff_A_fO4se0o44_0),.din(w_dff_A_8Y9VSXqN9_0),.clk(gclk));
	jdff dff_A_fO4se0o44_0(.dout(w_dff_A_tR5P0jYG9_0),.din(w_dff_A_fO4se0o44_0),.clk(gclk));
	jdff dff_A_tR5P0jYG9_0(.dout(w_dff_A_B1PheY4K2_0),.din(w_dff_A_tR5P0jYG9_0),.clk(gclk));
	jdff dff_A_B1PheY4K2_0(.dout(w_dff_A_O1scLa9C1_0),.din(w_dff_A_B1PheY4K2_0),.clk(gclk));
	jdff dff_A_O1scLa9C1_0(.dout(w_dff_A_I7VUaWfu0_0),.din(w_dff_A_O1scLa9C1_0),.clk(gclk));
	jdff dff_A_I7VUaWfu0_0(.dout(w_dff_A_X8IZP3vW9_0),.din(w_dff_A_I7VUaWfu0_0),.clk(gclk));
	jdff dff_A_X8IZP3vW9_0(.dout(w_dff_A_pmSQrNhR3_0),.din(w_dff_A_X8IZP3vW9_0),.clk(gclk));
	jdff dff_A_pmSQrNhR3_0(.dout(w_dff_A_zTi8jiHI0_0),.din(w_dff_A_pmSQrNhR3_0),.clk(gclk));
	jdff dff_A_zTi8jiHI0_0(.dout(w_dff_A_GnmzxZgJ0_0),.din(w_dff_A_zTi8jiHI0_0),.clk(gclk));
	jdff dff_A_GnmzxZgJ0_0(.dout(w_dff_A_Wfdp2Woa9_0),.din(w_dff_A_GnmzxZgJ0_0),.clk(gclk));
	jdff dff_A_Wfdp2Woa9_0(.dout(w_dff_A_NiBiFuvV6_0),.din(w_dff_A_Wfdp2Woa9_0),.clk(gclk));
	jdff dff_A_NiBiFuvV6_0(.dout(w_dff_A_GBKZmWoa2_0),.din(w_dff_A_NiBiFuvV6_0),.clk(gclk));
	jdff dff_A_GBKZmWoa2_0(.dout(w_dff_A_9RgFqwdU7_0),.din(w_dff_A_GBKZmWoa2_0),.clk(gclk));
	jdff dff_A_9RgFqwdU7_0(.dout(w_dff_A_kMmQEkZV6_0),.din(w_dff_A_9RgFqwdU7_0),.clk(gclk));
	jdff dff_A_kMmQEkZV6_0(.dout(w_dff_A_IfwIk9Mo6_0),.din(w_dff_A_kMmQEkZV6_0),.clk(gclk));
	jdff dff_A_IfwIk9Mo6_0(.dout(w_dff_A_qFwxWb6H9_0),.din(w_dff_A_IfwIk9Mo6_0),.clk(gclk));
	jdff dff_A_qFwxWb6H9_0(.dout(w_dff_A_9T4GLeUL7_0),.din(w_dff_A_qFwxWb6H9_0),.clk(gclk));
	jdff dff_A_9T4GLeUL7_0(.dout(w_dff_A_pnPsdKjh3_0),.din(w_dff_A_9T4GLeUL7_0),.clk(gclk));
	jdff dff_A_pnPsdKjh3_0(.dout(w_dff_A_7IIicVW07_0),.din(w_dff_A_pnPsdKjh3_0),.clk(gclk));
	jdff dff_A_7IIicVW07_0(.dout(w_dff_A_KQoFEcxO5_0),.din(w_dff_A_7IIicVW07_0),.clk(gclk));
	jdff dff_A_KQoFEcxO5_0(.dout(w_dff_A_vx3J51w74_0),.din(w_dff_A_KQoFEcxO5_0),.clk(gclk));
	jdff dff_A_vx3J51w74_0(.dout(w_dff_A_XJDpRknC7_0),.din(w_dff_A_vx3J51w74_0),.clk(gclk));
	jdff dff_A_XJDpRknC7_0(.dout(w_dff_A_AdZ9fheF7_0),.din(w_dff_A_XJDpRknC7_0),.clk(gclk));
	jdff dff_A_AdZ9fheF7_0(.dout(w_dff_A_5KNDTQtG6_0),.din(w_dff_A_AdZ9fheF7_0),.clk(gclk));
	jdff dff_A_5KNDTQtG6_0(.dout(w_dff_A_id4zQhtR6_0),.din(w_dff_A_5KNDTQtG6_0),.clk(gclk));
	jdff dff_A_id4zQhtR6_0(.dout(w_dff_A_0YQTmjmN1_0),.din(w_dff_A_id4zQhtR6_0),.clk(gclk));
	jdff dff_A_0YQTmjmN1_0(.dout(w_dff_A_OSb0Z9x99_0),.din(w_dff_A_0YQTmjmN1_0),.clk(gclk));
	jdff dff_A_OSb0Z9x99_0(.dout(G438),.din(w_dff_A_OSb0Z9x99_0),.clk(gclk));
	jdff dff_A_80xgeO6u2_1(.dout(w_dff_A_ezgQ9NYB2_0),.din(w_dff_A_80xgeO6u2_1),.clk(gclk));
	jdff dff_A_ezgQ9NYB2_0(.dout(w_dff_A_biwJmZpO0_0),.din(w_dff_A_ezgQ9NYB2_0),.clk(gclk));
	jdff dff_A_biwJmZpO0_0(.dout(w_dff_A_JkUfybyo6_0),.din(w_dff_A_biwJmZpO0_0),.clk(gclk));
	jdff dff_A_JkUfybyo6_0(.dout(w_dff_A_v58gaw6T7_0),.din(w_dff_A_JkUfybyo6_0),.clk(gclk));
	jdff dff_A_v58gaw6T7_0(.dout(w_dff_A_bzeXVAKH7_0),.din(w_dff_A_v58gaw6T7_0),.clk(gclk));
	jdff dff_A_bzeXVAKH7_0(.dout(w_dff_A_z3P9eGGF9_0),.din(w_dff_A_bzeXVAKH7_0),.clk(gclk));
	jdff dff_A_z3P9eGGF9_0(.dout(w_dff_A_APjyFnb33_0),.din(w_dff_A_z3P9eGGF9_0),.clk(gclk));
	jdff dff_A_APjyFnb33_0(.dout(w_dff_A_YWuP8LU71_0),.din(w_dff_A_APjyFnb33_0),.clk(gclk));
	jdff dff_A_YWuP8LU71_0(.dout(w_dff_A_5dRQYwzG2_0),.din(w_dff_A_YWuP8LU71_0),.clk(gclk));
	jdff dff_A_5dRQYwzG2_0(.dout(w_dff_A_0llwhG3y7_0),.din(w_dff_A_5dRQYwzG2_0),.clk(gclk));
	jdff dff_A_0llwhG3y7_0(.dout(w_dff_A_FYuuIKS63_0),.din(w_dff_A_0llwhG3y7_0),.clk(gclk));
	jdff dff_A_FYuuIKS63_0(.dout(w_dff_A_6dW1B7MK5_0),.din(w_dff_A_FYuuIKS63_0),.clk(gclk));
	jdff dff_A_6dW1B7MK5_0(.dout(w_dff_A_nOmjzmaC0_0),.din(w_dff_A_6dW1B7MK5_0),.clk(gclk));
	jdff dff_A_nOmjzmaC0_0(.dout(w_dff_A_8plihuOL8_0),.din(w_dff_A_nOmjzmaC0_0),.clk(gclk));
	jdff dff_A_8plihuOL8_0(.dout(w_dff_A_LNIor2Xf0_0),.din(w_dff_A_8plihuOL8_0),.clk(gclk));
	jdff dff_A_LNIor2Xf0_0(.dout(w_dff_A_CEBDPqtw5_0),.din(w_dff_A_LNIor2Xf0_0),.clk(gclk));
	jdff dff_A_CEBDPqtw5_0(.dout(w_dff_A_16OuaOQH2_0),.din(w_dff_A_CEBDPqtw5_0),.clk(gclk));
	jdff dff_A_16OuaOQH2_0(.dout(w_dff_A_AVimHYPv4_0),.din(w_dff_A_16OuaOQH2_0),.clk(gclk));
	jdff dff_A_AVimHYPv4_0(.dout(w_dff_A_vvESrzoA1_0),.din(w_dff_A_AVimHYPv4_0),.clk(gclk));
	jdff dff_A_vvESrzoA1_0(.dout(w_dff_A_yATOE5Va9_0),.din(w_dff_A_vvESrzoA1_0),.clk(gclk));
	jdff dff_A_yATOE5Va9_0(.dout(w_dff_A_EcludsJw6_0),.din(w_dff_A_yATOE5Va9_0),.clk(gclk));
	jdff dff_A_EcludsJw6_0(.dout(w_dff_A_pY3RRJxD2_0),.din(w_dff_A_EcludsJw6_0),.clk(gclk));
	jdff dff_A_pY3RRJxD2_0(.dout(w_dff_A_WFNoR3kn7_0),.din(w_dff_A_pY3RRJxD2_0),.clk(gclk));
	jdff dff_A_WFNoR3kn7_0(.dout(w_dff_A_MHpEk0p79_0),.din(w_dff_A_WFNoR3kn7_0),.clk(gclk));
	jdff dff_A_MHpEk0p79_0(.dout(w_dff_A_WOmtw4fb2_0),.din(w_dff_A_MHpEk0p79_0),.clk(gclk));
	jdff dff_A_WOmtw4fb2_0(.dout(w_dff_A_ZmMtlInh1_0),.din(w_dff_A_WOmtw4fb2_0),.clk(gclk));
	jdff dff_A_ZmMtlInh1_0(.dout(w_dff_A_RHUMRomJ5_0),.din(w_dff_A_ZmMtlInh1_0),.clk(gclk));
	jdff dff_A_RHUMRomJ5_0(.dout(w_dff_A_dJNh6HjZ3_0),.din(w_dff_A_RHUMRomJ5_0),.clk(gclk));
	jdff dff_A_dJNh6HjZ3_0(.dout(w_dff_A_RbrVPB010_0),.din(w_dff_A_dJNh6HjZ3_0),.clk(gclk));
	jdff dff_A_RbrVPB010_0(.dout(w_dff_A_g0nl9VDs2_0),.din(w_dff_A_RbrVPB010_0),.clk(gclk));
	jdff dff_A_g0nl9VDs2_0(.dout(w_dff_A_9IjAxkMp3_0),.din(w_dff_A_g0nl9VDs2_0),.clk(gclk));
	jdff dff_A_9IjAxkMp3_0(.dout(w_dff_A_SuYkeoy75_0),.din(w_dff_A_9IjAxkMp3_0),.clk(gclk));
	jdff dff_A_SuYkeoy75_0(.dout(w_dff_A_pxcwxjmd6_0),.din(w_dff_A_SuYkeoy75_0),.clk(gclk));
	jdff dff_A_pxcwxjmd6_0(.dout(w_dff_A_ec3ctuvZ9_0),.din(w_dff_A_pxcwxjmd6_0),.clk(gclk));
	jdff dff_A_ec3ctuvZ9_0(.dout(w_dff_A_Tf1nq2nt0_0),.din(w_dff_A_ec3ctuvZ9_0),.clk(gclk));
	jdff dff_A_Tf1nq2nt0_0(.dout(w_dff_A_cRrTHZtY5_0),.din(w_dff_A_Tf1nq2nt0_0),.clk(gclk));
	jdff dff_A_cRrTHZtY5_0(.dout(w_dff_A_mxSh4hRX4_0),.din(w_dff_A_cRrTHZtY5_0),.clk(gclk));
	jdff dff_A_mxSh4hRX4_0(.dout(w_dff_A_8yyeYsUc3_0),.din(w_dff_A_mxSh4hRX4_0),.clk(gclk));
	jdff dff_A_8yyeYsUc3_0(.dout(G496),.din(w_dff_A_8yyeYsUc3_0),.clk(gclk));
	jdff dff_A_YVg7X2Az1_1(.dout(w_dff_A_MXaWD79m3_0),.din(w_dff_A_YVg7X2Az1_1),.clk(gclk));
	jdff dff_A_MXaWD79m3_0(.dout(w_dff_A_jLdr1f5V8_0),.din(w_dff_A_MXaWD79m3_0),.clk(gclk));
	jdff dff_A_jLdr1f5V8_0(.dout(w_dff_A_UFyh85405_0),.din(w_dff_A_jLdr1f5V8_0),.clk(gclk));
	jdff dff_A_UFyh85405_0(.dout(w_dff_A_p1eiRlI63_0),.din(w_dff_A_UFyh85405_0),.clk(gclk));
	jdff dff_A_p1eiRlI63_0(.dout(w_dff_A_FNKxDVsY5_0),.din(w_dff_A_p1eiRlI63_0),.clk(gclk));
	jdff dff_A_FNKxDVsY5_0(.dout(w_dff_A_GpjnpPWB6_0),.din(w_dff_A_FNKxDVsY5_0),.clk(gclk));
	jdff dff_A_GpjnpPWB6_0(.dout(w_dff_A_WRkQc04j3_0),.din(w_dff_A_GpjnpPWB6_0),.clk(gclk));
	jdff dff_A_WRkQc04j3_0(.dout(w_dff_A_t4dCEtDO0_0),.din(w_dff_A_WRkQc04j3_0),.clk(gclk));
	jdff dff_A_t4dCEtDO0_0(.dout(w_dff_A_GbRewRmk2_0),.din(w_dff_A_t4dCEtDO0_0),.clk(gclk));
	jdff dff_A_GbRewRmk2_0(.dout(w_dff_A_AO0R8pZt7_0),.din(w_dff_A_GbRewRmk2_0),.clk(gclk));
	jdff dff_A_AO0R8pZt7_0(.dout(w_dff_A_Sd5Okzlu6_0),.din(w_dff_A_AO0R8pZt7_0),.clk(gclk));
	jdff dff_A_Sd5Okzlu6_0(.dout(w_dff_A_utuPAZp03_0),.din(w_dff_A_Sd5Okzlu6_0),.clk(gclk));
	jdff dff_A_utuPAZp03_0(.dout(w_dff_A_i314Kx4Z4_0),.din(w_dff_A_utuPAZp03_0),.clk(gclk));
	jdff dff_A_i314Kx4Z4_0(.dout(w_dff_A_8cMlb01G5_0),.din(w_dff_A_i314Kx4Z4_0),.clk(gclk));
	jdff dff_A_8cMlb01G5_0(.dout(w_dff_A_aeMYdjSe5_0),.din(w_dff_A_8cMlb01G5_0),.clk(gclk));
	jdff dff_A_aeMYdjSe5_0(.dout(w_dff_A_VYRWkyGi3_0),.din(w_dff_A_aeMYdjSe5_0),.clk(gclk));
	jdff dff_A_VYRWkyGi3_0(.dout(w_dff_A_CiJDJtQR6_0),.din(w_dff_A_VYRWkyGi3_0),.clk(gclk));
	jdff dff_A_CiJDJtQR6_0(.dout(w_dff_A_KW1APJHx1_0),.din(w_dff_A_CiJDJtQR6_0),.clk(gclk));
	jdff dff_A_KW1APJHx1_0(.dout(w_dff_A_8FTIaBrG0_0),.din(w_dff_A_KW1APJHx1_0),.clk(gclk));
	jdff dff_A_8FTIaBrG0_0(.dout(w_dff_A_cEPE2HEn9_0),.din(w_dff_A_8FTIaBrG0_0),.clk(gclk));
	jdff dff_A_cEPE2HEn9_0(.dout(w_dff_A_fGni8lWD1_0),.din(w_dff_A_cEPE2HEn9_0),.clk(gclk));
	jdff dff_A_fGni8lWD1_0(.dout(w_dff_A_UXajtxwi9_0),.din(w_dff_A_fGni8lWD1_0),.clk(gclk));
	jdff dff_A_UXajtxwi9_0(.dout(w_dff_A_AOieRl762_0),.din(w_dff_A_UXajtxwi9_0),.clk(gclk));
	jdff dff_A_AOieRl762_0(.dout(w_dff_A_e9d9JLwp0_0),.din(w_dff_A_AOieRl762_0),.clk(gclk));
	jdff dff_A_e9d9JLwp0_0(.dout(w_dff_A_gQNRETQP8_0),.din(w_dff_A_e9d9JLwp0_0),.clk(gclk));
	jdff dff_A_gQNRETQP8_0(.dout(w_dff_A_1IKU9MDR5_0),.din(w_dff_A_gQNRETQP8_0),.clk(gclk));
	jdff dff_A_1IKU9MDR5_0(.dout(w_dff_A_YtYnKT9c6_0),.din(w_dff_A_1IKU9MDR5_0),.clk(gclk));
	jdff dff_A_YtYnKT9c6_0(.dout(w_dff_A_lhyrcOQn2_0),.din(w_dff_A_YtYnKT9c6_0),.clk(gclk));
	jdff dff_A_lhyrcOQn2_0(.dout(w_dff_A_xUhD7t390_0),.din(w_dff_A_lhyrcOQn2_0),.clk(gclk));
	jdff dff_A_xUhD7t390_0(.dout(w_dff_A_nkJ6LJve5_0),.din(w_dff_A_xUhD7t390_0),.clk(gclk));
	jdff dff_A_nkJ6LJve5_0(.dout(w_dff_A_xznqdVAg2_0),.din(w_dff_A_nkJ6LJve5_0),.clk(gclk));
	jdff dff_A_xznqdVAg2_0(.dout(w_dff_A_SCLFNjAf3_0),.din(w_dff_A_xznqdVAg2_0),.clk(gclk));
	jdff dff_A_SCLFNjAf3_0(.dout(w_dff_A_lmcW9Wyn7_0),.din(w_dff_A_SCLFNjAf3_0),.clk(gclk));
	jdff dff_A_lmcW9Wyn7_0(.dout(w_dff_A_vlXgyy7X4_0),.din(w_dff_A_lmcW9Wyn7_0),.clk(gclk));
	jdff dff_A_vlXgyy7X4_0(.dout(w_dff_A_lKgm11G57_0),.din(w_dff_A_vlXgyy7X4_0),.clk(gclk));
	jdff dff_A_lKgm11G57_0(.dout(w_dff_A_4uC7qwO28_0),.din(w_dff_A_lKgm11G57_0),.clk(gclk));
	jdff dff_A_4uC7qwO28_0(.dout(w_dff_A_JYBOTeNq5_0),.din(w_dff_A_4uC7qwO28_0),.clk(gclk));
	jdff dff_A_JYBOTeNq5_0(.dout(w_dff_A_cRtgBYsu5_0),.din(w_dff_A_JYBOTeNq5_0),.clk(gclk));
	jdff dff_A_cRtgBYsu5_0(.dout(G494),.din(w_dff_A_cRtgBYsu5_0),.clk(gclk));
	jdff dff_A_mpaoxbKU2_1(.dout(w_dff_A_cYZ2IKGn7_0),.din(w_dff_A_mpaoxbKU2_1),.clk(gclk));
	jdff dff_A_cYZ2IKGn7_0(.dout(w_dff_A_cycveu3Z7_0),.din(w_dff_A_cYZ2IKGn7_0),.clk(gclk));
	jdff dff_A_cycveu3Z7_0(.dout(w_dff_A_CIoCGSL70_0),.din(w_dff_A_cycveu3Z7_0),.clk(gclk));
	jdff dff_A_CIoCGSL70_0(.dout(w_dff_A_J2ionYCO1_0),.din(w_dff_A_CIoCGSL70_0),.clk(gclk));
	jdff dff_A_J2ionYCO1_0(.dout(w_dff_A_K2yjXhet7_0),.din(w_dff_A_J2ionYCO1_0),.clk(gclk));
	jdff dff_A_K2yjXhet7_0(.dout(w_dff_A_anAyCNaC6_0),.din(w_dff_A_K2yjXhet7_0),.clk(gclk));
	jdff dff_A_anAyCNaC6_0(.dout(w_dff_A_zJlDiPSJ3_0),.din(w_dff_A_anAyCNaC6_0),.clk(gclk));
	jdff dff_A_zJlDiPSJ3_0(.dout(w_dff_A_g9kp4wvI9_0),.din(w_dff_A_zJlDiPSJ3_0),.clk(gclk));
	jdff dff_A_g9kp4wvI9_0(.dout(w_dff_A_omvzH8zG3_0),.din(w_dff_A_g9kp4wvI9_0),.clk(gclk));
	jdff dff_A_omvzH8zG3_0(.dout(w_dff_A_ccqN55Ia5_0),.din(w_dff_A_omvzH8zG3_0),.clk(gclk));
	jdff dff_A_ccqN55Ia5_0(.dout(w_dff_A_6gbjhOCs0_0),.din(w_dff_A_ccqN55Ia5_0),.clk(gclk));
	jdff dff_A_6gbjhOCs0_0(.dout(w_dff_A_4MBoiJ1d1_0),.din(w_dff_A_6gbjhOCs0_0),.clk(gclk));
	jdff dff_A_4MBoiJ1d1_0(.dout(w_dff_A_O8VjdEiG0_0),.din(w_dff_A_4MBoiJ1d1_0),.clk(gclk));
	jdff dff_A_O8VjdEiG0_0(.dout(w_dff_A_xioW0aD39_0),.din(w_dff_A_O8VjdEiG0_0),.clk(gclk));
	jdff dff_A_xioW0aD39_0(.dout(w_dff_A_1CvV8QTk9_0),.din(w_dff_A_xioW0aD39_0),.clk(gclk));
	jdff dff_A_1CvV8QTk9_0(.dout(w_dff_A_tR8aNwGo7_0),.din(w_dff_A_1CvV8QTk9_0),.clk(gclk));
	jdff dff_A_tR8aNwGo7_0(.dout(w_dff_A_nBYRpbld3_0),.din(w_dff_A_tR8aNwGo7_0),.clk(gclk));
	jdff dff_A_nBYRpbld3_0(.dout(w_dff_A_kvRiJ8q16_0),.din(w_dff_A_nBYRpbld3_0),.clk(gclk));
	jdff dff_A_kvRiJ8q16_0(.dout(w_dff_A_qWhhbW5h1_0),.din(w_dff_A_kvRiJ8q16_0),.clk(gclk));
	jdff dff_A_qWhhbW5h1_0(.dout(w_dff_A_dfq6BZrT7_0),.din(w_dff_A_qWhhbW5h1_0),.clk(gclk));
	jdff dff_A_dfq6BZrT7_0(.dout(w_dff_A_VyTe9x7Q3_0),.din(w_dff_A_dfq6BZrT7_0),.clk(gclk));
	jdff dff_A_VyTe9x7Q3_0(.dout(w_dff_A_vJ6wse6q6_0),.din(w_dff_A_VyTe9x7Q3_0),.clk(gclk));
	jdff dff_A_vJ6wse6q6_0(.dout(w_dff_A_XbiUDmNj9_0),.din(w_dff_A_vJ6wse6q6_0),.clk(gclk));
	jdff dff_A_XbiUDmNj9_0(.dout(w_dff_A_r2vlyFyq6_0),.din(w_dff_A_XbiUDmNj9_0),.clk(gclk));
	jdff dff_A_r2vlyFyq6_0(.dout(w_dff_A_uPjsHCum6_0),.din(w_dff_A_r2vlyFyq6_0),.clk(gclk));
	jdff dff_A_uPjsHCum6_0(.dout(w_dff_A_KJTLbru53_0),.din(w_dff_A_uPjsHCum6_0),.clk(gclk));
	jdff dff_A_KJTLbru53_0(.dout(w_dff_A_bfFVPh7U2_0),.din(w_dff_A_KJTLbru53_0),.clk(gclk));
	jdff dff_A_bfFVPh7U2_0(.dout(w_dff_A_g2brIlxC0_0),.din(w_dff_A_bfFVPh7U2_0),.clk(gclk));
	jdff dff_A_g2brIlxC0_0(.dout(w_dff_A_nCLp73rZ4_0),.din(w_dff_A_g2brIlxC0_0),.clk(gclk));
	jdff dff_A_nCLp73rZ4_0(.dout(w_dff_A_5XSOq4r64_0),.din(w_dff_A_nCLp73rZ4_0),.clk(gclk));
	jdff dff_A_5XSOq4r64_0(.dout(w_dff_A_j5H86hvk2_0),.din(w_dff_A_5XSOq4r64_0),.clk(gclk));
	jdff dff_A_j5H86hvk2_0(.dout(w_dff_A_m4SKr0up3_0),.din(w_dff_A_j5H86hvk2_0),.clk(gclk));
	jdff dff_A_m4SKr0up3_0(.dout(w_dff_A_4Eq57y9q2_0),.din(w_dff_A_m4SKr0up3_0),.clk(gclk));
	jdff dff_A_4Eq57y9q2_0(.dout(w_dff_A_TNHctidh2_0),.din(w_dff_A_4Eq57y9q2_0),.clk(gclk));
	jdff dff_A_TNHctidh2_0(.dout(w_dff_A_YOpylAWh6_0),.din(w_dff_A_TNHctidh2_0),.clk(gclk));
	jdff dff_A_YOpylAWh6_0(.dout(w_dff_A_X8mRE8At2_0),.din(w_dff_A_YOpylAWh6_0),.clk(gclk));
	jdff dff_A_X8mRE8At2_0(.dout(w_dff_A_TFZIlna89_0),.din(w_dff_A_X8mRE8At2_0),.clk(gclk));
	jdff dff_A_TFZIlna89_0(.dout(w_dff_A_NG80fwJf3_0),.din(w_dff_A_TFZIlna89_0),.clk(gclk));
	jdff dff_A_NG80fwJf3_0(.dout(G492),.din(w_dff_A_NG80fwJf3_0),.clk(gclk));
	jdff dff_A_gICE3Ix18_1(.dout(w_dff_A_hAy73yhW6_0),.din(w_dff_A_gICE3Ix18_1),.clk(gclk));
	jdff dff_A_hAy73yhW6_0(.dout(w_dff_A_mIioMXJ75_0),.din(w_dff_A_hAy73yhW6_0),.clk(gclk));
	jdff dff_A_mIioMXJ75_0(.dout(w_dff_A_OkALlnOw5_0),.din(w_dff_A_mIioMXJ75_0),.clk(gclk));
	jdff dff_A_OkALlnOw5_0(.dout(w_dff_A_UhZFbW2Y2_0),.din(w_dff_A_OkALlnOw5_0),.clk(gclk));
	jdff dff_A_UhZFbW2Y2_0(.dout(w_dff_A_JS6anSuB8_0),.din(w_dff_A_UhZFbW2Y2_0),.clk(gclk));
	jdff dff_A_JS6anSuB8_0(.dout(w_dff_A_bhDUjaVG7_0),.din(w_dff_A_JS6anSuB8_0),.clk(gclk));
	jdff dff_A_bhDUjaVG7_0(.dout(w_dff_A_qk8ezBHH1_0),.din(w_dff_A_bhDUjaVG7_0),.clk(gclk));
	jdff dff_A_qk8ezBHH1_0(.dout(w_dff_A_jftG65BW3_0),.din(w_dff_A_qk8ezBHH1_0),.clk(gclk));
	jdff dff_A_jftG65BW3_0(.dout(w_dff_A_W60Ja46K7_0),.din(w_dff_A_jftG65BW3_0),.clk(gclk));
	jdff dff_A_W60Ja46K7_0(.dout(w_dff_A_aRka5JIz5_0),.din(w_dff_A_W60Ja46K7_0),.clk(gclk));
	jdff dff_A_aRka5JIz5_0(.dout(w_dff_A_jlLkGC4H5_0),.din(w_dff_A_aRka5JIz5_0),.clk(gclk));
	jdff dff_A_jlLkGC4H5_0(.dout(w_dff_A_RkGwdNfh5_0),.din(w_dff_A_jlLkGC4H5_0),.clk(gclk));
	jdff dff_A_RkGwdNfh5_0(.dout(w_dff_A_XvFD3BqM1_0),.din(w_dff_A_RkGwdNfh5_0),.clk(gclk));
	jdff dff_A_XvFD3BqM1_0(.dout(w_dff_A_NgdQUWgm4_0),.din(w_dff_A_XvFD3BqM1_0),.clk(gclk));
	jdff dff_A_NgdQUWgm4_0(.dout(w_dff_A_gMMartza4_0),.din(w_dff_A_NgdQUWgm4_0),.clk(gclk));
	jdff dff_A_gMMartza4_0(.dout(w_dff_A_3NpBXOue6_0),.din(w_dff_A_gMMartza4_0),.clk(gclk));
	jdff dff_A_3NpBXOue6_0(.dout(w_dff_A_yBAykUBv1_0),.din(w_dff_A_3NpBXOue6_0),.clk(gclk));
	jdff dff_A_yBAykUBv1_0(.dout(w_dff_A_rStL3uCh5_0),.din(w_dff_A_yBAykUBv1_0),.clk(gclk));
	jdff dff_A_rStL3uCh5_0(.dout(w_dff_A_pY3iuBvZ6_0),.din(w_dff_A_rStL3uCh5_0),.clk(gclk));
	jdff dff_A_pY3iuBvZ6_0(.dout(w_dff_A_2v8gQzCh1_0),.din(w_dff_A_pY3iuBvZ6_0),.clk(gclk));
	jdff dff_A_2v8gQzCh1_0(.dout(w_dff_A_7iOw09Wk2_0),.din(w_dff_A_2v8gQzCh1_0),.clk(gclk));
	jdff dff_A_7iOw09Wk2_0(.dout(w_dff_A_3EDjtkm78_0),.din(w_dff_A_7iOw09Wk2_0),.clk(gclk));
	jdff dff_A_3EDjtkm78_0(.dout(w_dff_A_LpddJ1ql4_0),.din(w_dff_A_3EDjtkm78_0),.clk(gclk));
	jdff dff_A_LpddJ1ql4_0(.dout(w_dff_A_AERKqKoX2_0),.din(w_dff_A_LpddJ1ql4_0),.clk(gclk));
	jdff dff_A_AERKqKoX2_0(.dout(w_dff_A_Q0Nw8LDx6_0),.din(w_dff_A_AERKqKoX2_0),.clk(gclk));
	jdff dff_A_Q0Nw8LDx6_0(.dout(w_dff_A_NxLKSlcU2_0),.din(w_dff_A_Q0Nw8LDx6_0),.clk(gclk));
	jdff dff_A_NxLKSlcU2_0(.dout(w_dff_A_rJYzxeyq1_0),.din(w_dff_A_NxLKSlcU2_0),.clk(gclk));
	jdff dff_A_rJYzxeyq1_0(.dout(w_dff_A_qWbwLqEz2_0),.din(w_dff_A_rJYzxeyq1_0),.clk(gclk));
	jdff dff_A_qWbwLqEz2_0(.dout(w_dff_A_Ck2igJu86_0),.din(w_dff_A_qWbwLqEz2_0),.clk(gclk));
	jdff dff_A_Ck2igJu86_0(.dout(w_dff_A_ASAKMGb29_0),.din(w_dff_A_Ck2igJu86_0),.clk(gclk));
	jdff dff_A_ASAKMGb29_0(.dout(w_dff_A_APh0v85o0_0),.din(w_dff_A_ASAKMGb29_0),.clk(gclk));
	jdff dff_A_APh0v85o0_0(.dout(w_dff_A_cfYMOmt40_0),.din(w_dff_A_APh0v85o0_0),.clk(gclk));
	jdff dff_A_cfYMOmt40_0(.dout(w_dff_A_lDPvVcJx8_0),.din(w_dff_A_cfYMOmt40_0),.clk(gclk));
	jdff dff_A_lDPvVcJx8_0(.dout(w_dff_A_0gcyLViY4_0),.din(w_dff_A_lDPvVcJx8_0),.clk(gclk));
	jdff dff_A_0gcyLViY4_0(.dout(w_dff_A_7sM2PFdl2_0),.din(w_dff_A_0gcyLViY4_0),.clk(gclk));
	jdff dff_A_7sM2PFdl2_0(.dout(w_dff_A_Gkt4wVHe7_0),.din(w_dff_A_7sM2PFdl2_0),.clk(gclk));
	jdff dff_A_Gkt4wVHe7_0(.dout(w_dff_A_wZMYVtAT5_0),.din(w_dff_A_Gkt4wVHe7_0),.clk(gclk));
	jdff dff_A_wZMYVtAT5_0(.dout(w_dff_A_dR862AWT0_0),.din(w_dff_A_wZMYVtAT5_0),.clk(gclk));
	jdff dff_A_dR862AWT0_0(.dout(G490),.din(w_dff_A_dR862AWT0_0),.clk(gclk));
	jdff dff_A_m3c6GcYD1_1(.dout(w_dff_A_neS8Pgns2_0),.din(w_dff_A_m3c6GcYD1_1),.clk(gclk));
	jdff dff_A_neS8Pgns2_0(.dout(w_dff_A_rdz9Xd5D5_0),.din(w_dff_A_neS8Pgns2_0),.clk(gclk));
	jdff dff_A_rdz9Xd5D5_0(.dout(w_dff_A_ztTt08Oi4_0),.din(w_dff_A_rdz9Xd5D5_0),.clk(gclk));
	jdff dff_A_ztTt08Oi4_0(.dout(w_dff_A_943GbJWl9_0),.din(w_dff_A_ztTt08Oi4_0),.clk(gclk));
	jdff dff_A_943GbJWl9_0(.dout(w_dff_A_xTFEDmBO1_0),.din(w_dff_A_943GbJWl9_0),.clk(gclk));
	jdff dff_A_xTFEDmBO1_0(.dout(w_dff_A_nPOe1cdb0_0),.din(w_dff_A_xTFEDmBO1_0),.clk(gclk));
	jdff dff_A_nPOe1cdb0_0(.dout(w_dff_A_rXh3dXAu9_0),.din(w_dff_A_nPOe1cdb0_0),.clk(gclk));
	jdff dff_A_rXh3dXAu9_0(.dout(w_dff_A_9PXEMyFt7_0),.din(w_dff_A_rXh3dXAu9_0),.clk(gclk));
	jdff dff_A_9PXEMyFt7_0(.dout(w_dff_A_UwqongY06_0),.din(w_dff_A_9PXEMyFt7_0),.clk(gclk));
	jdff dff_A_UwqongY06_0(.dout(w_dff_A_w0K9tAnF1_0),.din(w_dff_A_UwqongY06_0),.clk(gclk));
	jdff dff_A_w0K9tAnF1_0(.dout(w_dff_A_Fb82YPe71_0),.din(w_dff_A_w0K9tAnF1_0),.clk(gclk));
	jdff dff_A_Fb82YPe71_0(.dout(w_dff_A_mstaH5dM2_0),.din(w_dff_A_Fb82YPe71_0),.clk(gclk));
	jdff dff_A_mstaH5dM2_0(.dout(w_dff_A_S8OODCLB7_0),.din(w_dff_A_mstaH5dM2_0),.clk(gclk));
	jdff dff_A_S8OODCLB7_0(.dout(w_dff_A_js3HKh461_0),.din(w_dff_A_S8OODCLB7_0),.clk(gclk));
	jdff dff_A_js3HKh461_0(.dout(w_dff_A_oKqEzSjx9_0),.din(w_dff_A_js3HKh461_0),.clk(gclk));
	jdff dff_A_oKqEzSjx9_0(.dout(w_dff_A_QJVmFa2Y6_0),.din(w_dff_A_oKqEzSjx9_0),.clk(gclk));
	jdff dff_A_QJVmFa2Y6_0(.dout(w_dff_A_f87hGuYl5_0),.din(w_dff_A_QJVmFa2Y6_0),.clk(gclk));
	jdff dff_A_f87hGuYl5_0(.dout(w_dff_A_XG7333ai6_0),.din(w_dff_A_f87hGuYl5_0),.clk(gclk));
	jdff dff_A_XG7333ai6_0(.dout(w_dff_A_cxYubjPU6_0),.din(w_dff_A_XG7333ai6_0),.clk(gclk));
	jdff dff_A_cxYubjPU6_0(.dout(w_dff_A_j34uCqX86_0),.din(w_dff_A_cxYubjPU6_0),.clk(gclk));
	jdff dff_A_j34uCqX86_0(.dout(w_dff_A_luFbhypQ6_0),.din(w_dff_A_j34uCqX86_0),.clk(gclk));
	jdff dff_A_luFbhypQ6_0(.dout(w_dff_A_sM0bIXdM6_0),.din(w_dff_A_luFbhypQ6_0),.clk(gclk));
	jdff dff_A_sM0bIXdM6_0(.dout(w_dff_A_HwhAxqBb0_0),.din(w_dff_A_sM0bIXdM6_0),.clk(gclk));
	jdff dff_A_HwhAxqBb0_0(.dout(w_dff_A_vNnowdhk0_0),.din(w_dff_A_HwhAxqBb0_0),.clk(gclk));
	jdff dff_A_vNnowdhk0_0(.dout(w_dff_A_MWNV53vX6_0),.din(w_dff_A_vNnowdhk0_0),.clk(gclk));
	jdff dff_A_MWNV53vX6_0(.dout(w_dff_A_oLMKUFjx2_0),.din(w_dff_A_MWNV53vX6_0),.clk(gclk));
	jdff dff_A_oLMKUFjx2_0(.dout(w_dff_A_8kp5LDLQ8_0),.din(w_dff_A_oLMKUFjx2_0),.clk(gclk));
	jdff dff_A_8kp5LDLQ8_0(.dout(w_dff_A_qfQRVDYx2_0),.din(w_dff_A_8kp5LDLQ8_0),.clk(gclk));
	jdff dff_A_qfQRVDYx2_0(.dout(w_dff_A_m1mERx9q2_0),.din(w_dff_A_qfQRVDYx2_0),.clk(gclk));
	jdff dff_A_m1mERx9q2_0(.dout(w_dff_A_N7UUOuJD4_0),.din(w_dff_A_m1mERx9q2_0),.clk(gclk));
	jdff dff_A_N7UUOuJD4_0(.dout(w_dff_A_Tng41wUW5_0),.din(w_dff_A_N7UUOuJD4_0),.clk(gclk));
	jdff dff_A_Tng41wUW5_0(.dout(w_dff_A_lhCvl2OA6_0),.din(w_dff_A_Tng41wUW5_0),.clk(gclk));
	jdff dff_A_lhCvl2OA6_0(.dout(w_dff_A_2N58DUVH5_0),.din(w_dff_A_lhCvl2OA6_0),.clk(gclk));
	jdff dff_A_2N58DUVH5_0(.dout(w_dff_A_49fNHbAV5_0),.din(w_dff_A_2N58DUVH5_0),.clk(gclk));
	jdff dff_A_49fNHbAV5_0(.dout(w_dff_A_tvUAzi222_0),.din(w_dff_A_49fNHbAV5_0),.clk(gclk));
	jdff dff_A_tvUAzi222_0(.dout(w_dff_A_JnVh7jBS1_0),.din(w_dff_A_tvUAzi222_0),.clk(gclk));
	jdff dff_A_JnVh7jBS1_0(.dout(w_dff_A_23cXEvfi6_0),.din(w_dff_A_JnVh7jBS1_0),.clk(gclk));
	jdff dff_A_23cXEvfi6_0(.dout(w_dff_A_veXBQrut6_0),.din(w_dff_A_23cXEvfi6_0),.clk(gclk));
	jdff dff_A_veXBQrut6_0(.dout(G488),.din(w_dff_A_veXBQrut6_0),.clk(gclk));
	jdff dff_A_DbjIJw5y8_1(.dout(w_dff_A_QYSelc0D7_0),.din(w_dff_A_DbjIJw5y8_1),.clk(gclk));
	jdff dff_A_QYSelc0D7_0(.dout(w_dff_A_Tq1uZKXt2_0),.din(w_dff_A_QYSelc0D7_0),.clk(gclk));
	jdff dff_A_Tq1uZKXt2_0(.dout(w_dff_A_97EzWTwg3_0),.din(w_dff_A_Tq1uZKXt2_0),.clk(gclk));
	jdff dff_A_97EzWTwg3_0(.dout(w_dff_A_FWtycdES8_0),.din(w_dff_A_97EzWTwg3_0),.clk(gclk));
	jdff dff_A_FWtycdES8_0(.dout(w_dff_A_R0yC1cZQ9_0),.din(w_dff_A_FWtycdES8_0),.clk(gclk));
	jdff dff_A_R0yC1cZQ9_0(.dout(w_dff_A_Rhv9BR7e1_0),.din(w_dff_A_R0yC1cZQ9_0),.clk(gclk));
	jdff dff_A_Rhv9BR7e1_0(.dout(w_dff_A_dhGNVNjb8_0),.din(w_dff_A_Rhv9BR7e1_0),.clk(gclk));
	jdff dff_A_dhGNVNjb8_0(.dout(w_dff_A_cmhEXjT05_0),.din(w_dff_A_dhGNVNjb8_0),.clk(gclk));
	jdff dff_A_cmhEXjT05_0(.dout(w_dff_A_UtPqRUnd7_0),.din(w_dff_A_cmhEXjT05_0),.clk(gclk));
	jdff dff_A_UtPqRUnd7_0(.dout(w_dff_A_TRUcJJt18_0),.din(w_dff_A_UtPqRUnd7_0),.clk(gclk));
	jdff dff_A_TRUcJJt18_0(.dout(w_dff_A_64Xz9RBk9_0),.din(w_dff_A_TRUcJJt18_0),.clk(gclk));
	jdff dff_A_64Xz9RBk9_0(.dout(w_dff_A_0l3uT3AI1_0),.din(w_dff_A_64Xz9RBk9_0),.clk(gclk));
	jdff dff_A_0l3uT3AI1_0(.dout(w_dff_A_2Ty6CJTh4_0),.din(w_dff_A_0l3uT3AI1_0),.clk(gclk));
	jdff dff_A_2Ty6CJTh4_0(.dout(w_dff_A_RZ7SBawl7_0),.din(w_dff_A_2Ty6CJTh4_0),.clk(gclk));
	jdff dff_A_RZ7SBawl7_0(.dout(w_dff_A_Y3wCbXW99_0),.din(w_dff_A_RZ7SBawl7_0),.clk(gclk));
	jdff dff_A_Y3wCbXW99_0(.dout(w_dff_A_aqLYkpf27_0),.din(w_dff_A_Y3wCbXW99_0),.clk(gclk));
	jdff dff_A_aqLYkpf27_0(.dout(w_dff_A_Ydp6s5eV0_0),.din(w_dff_A_aqLYkpf27_0),.clk(gclk));
	jdff dff_A_Ydp6s5eV0_0(.dout(w_dff_A_vV0R2ADP3_0),.din(w_dff_A_Ydp6s5eV0_0),.clk(gclk));
	jdff dff_A_vV0R2ADP3_0(.dout(w_dff_A_xz0c9TPD2_0),.din(w_dff_A_vV0R2ADP3_0),.clk(gclk));
	jdff dff_A_xz0c9TPD2_0(.dout(w_dff_A_kVaBKblE5_0),.din(w_dff_A_xz0c9TPD2_0),.clk(gclk));
	jdff dff_A_kVaBKblE5_0(.dout(w_dff_A_JzBG10k53_0),.din(w_dff_A_kVaBKblE5_0),.clk(gclk));
	jdff dff_A_JzBG10k53_0(.dout(w_dff_A_0QyNtdmT3_0),.din(w_dff_A_JzBG10k53_0),.clk(gclk));
	jdff dff_A_0QyNtdmT3_0(.dout(w_dff_A_PnpAtMP68_0),.din(w_dff_A_0QyNtdmT3_0),.clk(gclk));
	jdff dff_A_PnpAtMP68_0(.dout(w_dff_A_3zeNyRdK4_0),.din(w_dff_A_PnpAtMP68_0),.clk(gclk));
	jdff dff_A_3zeNyRdK4_0(.dout(w_dff_A_PfcutuxV2_0),.din(w_dff_A_3zeNyRdK4_0),.clk(gclk));
	jdff dff_A_PfcutuxV2_0(.dout(w_dff_A_q7AOk8wm3_0),.din(w_dff_A_PfcutuxV2_0),.clk(gclk));
	jdff dff_A_q7AOk8wm3_0(.dout(w_dff_A_313SaAKf7_0),.din(w_dff_A_q7AOk8wm3_0),.clk(gclk));
	jdff dff_A_313SaAKf7_0(.dout(w_dff_A_5ST6FeWs7_0),.din(w_dff_A_313SaAKf7_0),.clk(gclk));
	jdff dff_A_5ST6FeWs7_0(.dout(w_dff_A_VcOPj1xB5_0),.din(w_dff_A_5ST6FeWs7_0),.clk(gclk));
	jdff dff_A_VcOPj1xB5_0(.dout(w_dff_A_XrKAWLTg1_0),.din(w_dff_A_VcOPj1xB5_0),.clk(gclk));
	jdff dff_A_XrKAWLTg1_0(.dout(w_dff_A_fS3KHqaN9_0),.din(w_dff_A_XrKAWLTg1_0),.clk(gclk));
	jdff dff_A_fS3KHqaN9_0(.dout(w_dff_A_dXsAKbSW6_0),.din(w_dff_A_fS3KHqaN9_0),.clk(gclk));
	jdff dff_A_dXsAKbSW6_0(.dout(w_dff_A_GcSKwiS31_0),.din(w_dff_A_dXsAKbSW6_0),.clk(gclk));
	jdff dff_A_GcSKwiS31_0(.dout(w_dff_A_hOyQfFMB6_0),.din(w_dff_A_GcSKwiS31_0),.clk(gclk));
	jdff dff_A_hOyQfFMB6_0(.dout(w_dff_A_DFrt3KYs7_0),.din(w_dff_A_hOyQfFMB6_0),.clk(gclk));
	jdff dff_A_DFrt3KYs7_0(.dout(w_dff_A_5X3ERRQL3_0),.din(w_dff_A_DFrt3KYs7_0),.clk(gclk));
	jdff dff_A_5X3ERRQL3_0(.dout(w_dff_A_4rFzbcav9_0),.din(w_dff_A_5X3ERRQL3_0),.clk(gclk));
	jdff dff_A_4rFzbcav9_0(.dout(w_dff_A_P2HSYyjk1_0),.din(w_dff_A_4rFzbcav9_0),.clk(gclk));
	jdff dff_A_P2HSYyjk1_0(.dout(G486),.din(w_dff_A_P2HSYyjk1_0),.clk(gclk));
	jdff dff_A_b76irSqt9_1(.dout(w_dff_A_reT6XF4V4_0),.din(w_dff_A_b76irSqt9_1),.clk(gclk));
	jdff dff_A_reT6XF4V4_0(.dout(w_dff_A_kXX141018_0),.din(w_dff_A_reT6XF4V4_0),.clk(gclk));
	jdff dff_A_kXX141018_0(.dout(w_dff_A_S3KLaESd4_0),.din(w_dff_A_kXX141018_0),.clk(gclk));
	jdff dff_A_S3KLaESd4_0(.dout(w_dff_A_P7ViR7n67_0),.din(w_dff_A_S3KLaESd4_0),.clk(gclk));
	jdff dff_A_P7ViR7n67_0(.dout(w_dff_A_yQLnTgxJ9_0),.din(w_dff_A_P7ViR7n67_0),.clk(gclk));
	jdff dff_A_yQLnTgxJ9_0(.dout(w_dff_A_NZ7CLybj4_0),.din(w_dff_A_yQLnTgxJ9_0),.clk(gclk));
	jdff dff_A_NZ7CLybj4_0(.dout(w_dff_A_cpmCXHgA6_0),.din(w_dff_A_NZ7CLybj4_0),.clk(gclk));
	jdff dff_A_cpmCXHgA6_0(.dout(w_dff_A_ILKfShA53_0),.din(w_dff_A_cpmCXHgA6_0),.clk(gclk));
	jdff dff_A_ILKfShA53_0(.dout(w_dff_A_kzQ9x1E33_0),.din(w_dff_A_ILKfShA53_0),.clk(gclk));
	jdff dff_A_kzQ9x1E33_0(.dout(w_dff_A_T3Fq2j7j1_0),.din(w_dff_A_kzQ9x1E33_0),.clk(gclk));
	jdff dff_A_T3Fq2j7j1_0(.dout(w_dff_A_oUahWUZq1_0),.din(w_dff_A_T3Fq2j7j1_0),.clk(gclk));
	jdff dff_A_oUahWUZq1_0(.dout(w_dff_A_h4gozfmx1_0),.din(w_dff_A_oUahWUZq1_0),.clk(gclk));
	jdff dff_A_h4gozfmx1_0(.dout(w_dff_A_Wt2eAbIB6_0),.din(w_dff_A_h4gozfmx1_0),.clk(gclk));
	jdff dff_A_Wt2eAbIB6_0(.dout(w_dff_A_bYX0Rqqi9_0),.din(w_dff_A_Wt2eAbIB6_0),.clk(gclk));
	jdff dff_A_bYX0Rqqi9_0(.dout(w_dff_A_a3awiYBU0_0),.din(w_dff_A_bYX0Rqqi9_0),.clk(gclk));
	jdff dff_A_a3awiYBU0_0(.dout(w_dff_A_DFBPr1fE6_0),.din(w_dff_A_a3awiYBU0_0),.clk(gclk));
	jdff dff_A_DFBPr1fE6_0(.dout(w_dff_A_lYij1PQv5_0),.din(w_dff_A_DFBPr1fE6_0),.clk(gclk));
	jdff dff_A_lYij1PQv5_0(.dout(w_dff_A_Nz1EZmFF7_0),.din(w_dff_A_lYij1PQv5_0),.clk(gclk));
	jdff dff_A_Nz1EZmFF7_0(.dout(w_dff_A_8WRbKEq50_0),.din(w_dff_A_Nz1EZmFF7_0),.clk(gclk));
	jdff dff_A_8WRbKEq50_0(.dout(w_dff_A_cvG73VD89_0),.din(w_dff_A_8WRbKEq50_0),.clk(gclk));
	jdff dff_A_cvG73VD89_0(.dout(w_dff_A_OUkmg86w7_0),.din(w_dff_A_cvG73VD89_0),.clk(gclk));
	jdff dff_A_OUkmg86w7_0(.dout(w_dff_A_CNqfQS2a6_0),.din(w_dff_A_OUkmg86w7_0),.clk(gclk));
	jdff dff_A_CNqfQS2a6_0(.dout(w_dff_A_BdPQEPs52_0),.din(w_dff_A_CNqfQS2a6_0),.clk(gclk));
	jdff dff_A_BdPQEPs52_0(.dout(w_dff_A_EOBdxKmj9_0),.din(w_dff_A_BdPQEPs52_0),.clk(gclk));
	jdff dff_A_EOBdxKmj9_0(.dout(w_dff_A_VwxVqiaW2_0),.din(w_dff_A_EOBdxKmj9_0),.clk(gclk));
	jdff dff_A_VwxVqiaW2_0(.dout(w_dff_A_vkFrLgkq8_0),.din(w_dff_A_VwxVqiaW2_0),.clk(gclk));
	jdff dff_A_vkFrLgkq8_0(.dout(w_dff_A_DK06YMd55_0),.din(w_dff_A_vkFrLgkq8_0),.clk(gclk));
	jdff dff_A_DK06YMd55_0(.dout(w_dff_A_bZTLqbwK9_0),.din(w_dff_A_DK06YMd55_0),.clk(gclk));
	jdff dff_A_bZTLqbwK9_0(.dout(w_dff_A_0FG6J8lp3_0),.din(w_dff_A_bZTLqbwK9_0),.clk(gclk));
	jdff dff_A_0FG6J8lp3_0(.dout(w_dff_A_qVey2nH26_0),.din(w_dff_A_0FG6J8lp3_0),.clk(gclk));
	jdff dff_A_qVey2nH26_0(.dout(w_dff_A_o7YYdPZb8_0),.din(w_dff_A_qVey2nH26_0),.clk(gclk));
	jdff dff_A_o7YYdPZb8_0(.dout(w_dff_A_8e3NSgGz4_0),.din(w_dff_A_o7YYdPZb8_0),.clk(gclk));
	jdff dff_A_8e3NSgGz4_0(.dout(w_dff_A_ZdajZTpo7_0),.din(w_dff_A_8e3NSgGz4_0),.clk(gclk));
	jdff dff_A_ZdajZTpo7_0(.dout(w_dff_A_G7pNbg3o5_0),.din(w_dff_A_ZdajZTpo7_0),.clk(gclk));
	jdff dff_A_G7pNbg3o5_0(.dout(w_dff_A_t15XqLDb6_0),.din(w_dff_A_G7pNbg3o5_0),.clk(gclk));
	jdff dff_A_t15XqLDb6_0(.dout(w_dff_A_i0uMMR9k8_0),.din(w_dff_A_t15XqLDb6_0),.clk(gclk));
	jdff dff_A_i0uMMR9k8_0(.dout(w_dff_A_RNq0drEK1_0),.din(w_dff_A_i0uMMR9k8_0),.clk(gclk));
	jdff dff_A_RNq0drEK1_0(.dout(w_dff_A_hp9W9RQd6_0),.din(w_dff_A_RNq0drEK1_0),.clk(gclk));
	jdff dff_A_hp9W9RQd6_0(.dout(G484),.din(w_dff_A_hp9W9RQd6_0),.clk(gclk));
	jdff dff_A_TsLfMgku7_1(.dout(w_dff_A_f1O61jzJ1_0),.din(w_dff_A_TsLfMgku7_1),.clk(gclk));
	jdff dff_A_f1O61jzJ1_0(.dout(w_dff_A_Lg3biNeC0_0),.din(w_dff_A_f1O61jzJ1_0),.clk(gclk));
	jdff dff_A_Lg3biNeC0_0(.dout(w_dff_A_PCzP35HW3_0),.din(w_dff_A_Lg3biNeC0_0),.clk(gclk));
	jdff dff_A_PCzP35HW3_0(.dout(w_dff_A_X7bcaziw6_0),.din(w_dff_A_PCzP35HW3_0),.clk(gclk));
	jdff dff_A_X7bcaziw6_0(.dout(w_dff_A_Ew4NW7Qv0_0),.din(w_dff_A_X7bcaziw6_0),.clk(gclk));
	jdff dff_A_Ew4NW7Qv0_0(.dout(w_dff_A_HR0ph5xB1_0),.din(w_dff_A_Ew4NW7Qv0_0),.clk(gclk));
	jdff dff_A_HR0ph5xB1_0(.dout(w_dff_A_hvp87gTd3_0),.din(w_dff_A_HR0ph5xB1_0),.clk(gclk));
	jdff dff_A_hvp87gTd3_0(.dout(w_dff_A_SnrefMJk4_0),.din(w_dff_A_hvp87gTd3_0),.clk(gclk));
	jdff dff_A_SnrefMJk4_0(.dout(w_dff_A_3j0jRYW06_0),.din(w_dff_A_SnrefMJk4_0),.clk(gclk));
	jdff dff_A_3j0jRYW06_0(.dout(w_dff_A_6uMRXNgg4_0),.din(w_dff_A_3j0jRYW06_0),.clk(gclk));
	jdff dff_A_6uMRXNgg4_0(.dout(w_dff_A_6ZoRoiwh3_0),.din(w_dff_A_6uMRXNgg4_0),.clk(gclk));
	jdff dff_A_6ZoRoiwh3_0(.dout(w_dff_A_YPFnoJnQ3_0),.din(w_dff_A_6ZoRoiwh3_0),.clk(gclk));
	jdff dff_A_YPFnoJnQ3_0(.dout(w_dff_A_fHfI0eZM9_0),.din(w_dff_A_YPFnoJnQ3_0),.clk(gclk));
	jdff dff_A_fHfI0eZM9_0(.dout(w_dff_A_gRuPA4TU2_0),.din(w_dff_A_fHfI0eZM9_0),.clk(gclk));
	jdff dff_A_gRuPA4TU2_0(.dout(w_dff_A_XOH9Vxbi6_0),.din(w_dff_A_gRuPA4TU2_0),.clk(gclk));
	jdff dff_A_XOH9Vxbi6_0(.dout(w_dff_A_cxzg8MLS7_0),.din(w_dff_A_XOH9Vxbi6_0),.clk(gclk));
	jdff dff_A_cxzg8MLS7_0(.dout(w_dff_A_IIkQb37F3_0),.din(w_dff_A_cxzg8MLS7_0),.clk(gclk));
	jdff dff_A_IIkQb37F3_0(.dout(w_dff_A_3SrfgKcy4_0),.din(w_dff_A_IIkQb37F3_0),.clk(gclk));
	jdff dff_A_3SrfgKcy4_0(.dout(w_dff_A_H0zE0MqB5_0),.din(w_dff_A_3SrfgKcy4_0),.clk(gclk));
	jdff dff_A_H0zE0MqB5_0(.dout(w_dff_A_jEJsBPDI2_0),.din(w_dff_A_H0zE0MqB5_0),.clk(gclk));
	jdff dff_A_jEJsBPDI2_0(.dout(w_dff_A_lwdGFB0M9_0),.din(w_dff_A_jEJsBPDI2_0),.clk(gclk));
	jdff dff_A_lwdGFB0M9_0(.dout(w_dff_A_E43OOoqb7_0),.din(w_dff_A_lwdGFB0M9_0),.clk(gclk));
	jdff dff_A_E43OOoqb7_0(.dout(w_dff_A_ExYbjIgL7_0),.din(w_dff_A_E43OOoqb7_0),.clk(gclk));
	jdff dff_A_ExYbjIgL7_0(.dout(w_dff_A_N99zULwH4_0),.din(w_dff_A_ExYbjIgL7_0),.clk(gclk));
	jdff dff_A_N99zULwH4_0(.dout(w_dff_A_Q7DsiNFS6_0),.din(w_dff_A_N99zULwH4_0),.clk(gclk));
	jdff dff_A_Q7DsiNFS6_0(.dout(w_dff_A_Bp9PA9I03_0),.din(w_dff_A_Q7DsiNFS6_0),.clk(gclk));
	jdff dff_A_Bp9PA9I03_0(.dout(w_dff_A_WHA63cDu3_0),.din(w_dff_A_Bp9PA9I03_0),.clk(gclk));
	jdff dff_A_WHA63cDu3_0(.dout(w_dff_A_88bYetJ04_0),.din(w_dff_A_WHA63cDu3_0),.clk(gclk));
	jdff dff_A_88bYetJ04_0(.dout(w_dff_A_aYKkb3F38_0),.din(w_dff_A_88bYetJ04_0),.clk(gclk));
	jdff dff_A_aYKkb3F38_0(.dout(w_dff_A_yvuYe1cI1_0),.din(w_dff_A_aYKkb3F38_0),.clk(gclk));
	jdff dff_A_yvuYe1cI1_0(.dout(w_dff_A_ecqAn2cX8_0),.din(w_dff_A_yvuYe1cI1_0),.clk(gclk));
	jdff dff_A_ecqAn2cX8_0(.dout(w_dff_A_Qx3u5Vze8_0),.din(w_dff_A_ecqAn2cX8_0),.clk(gclk));
	jdff dff_A_Qx3u5Vze8_0(.dout(w_dff_A_yLz1uhqc8_0),.din(w_dff_A_Qx3u5Vze8_0),.clk(gclk));
	jdff dff_A_yLz1uhqc8_0(.dout(w_dff_A_Ec1mXMq14_0),.din(w_dff_A_yLz1uhqc8_0),.clk(gclk));
	jdff dff_A_Ec1mXMq14_0(.dout(w_dff_A_Tw0LEMIy5_0),.din(w_dff_A_Ec1mXMq14_0),.clk(gclk));
	jdff dff_A_Tw0LEMIy5_0(.dout(w_dff_A_eZMBy8LW3_0),.din(w_dff_A_Tw0LEMIy5_0),.clk(gclk));
	jdff dff_A_eZMBy8LW3_0(.dout(w_dff_A_1VKNnZiP6_0),.din(w_dff_A_eZMBy8LW3_0),.clk(gclk));
	jdff dff_A_1VKNnZiP6_0(.dout(w_dff_A_53yowiEy8_0),.din(w_dff_A_1VKNnZiP6_0),.clk(gclk));
	jdff dff_A_53yowiEy8_0(.dout(G482),.din(w_dff_A_53yowiEy8_0),.clk(gclk));
	jdff dff_A_2530MqCy4_1(.dout(w_dff_A_u3ZY1c3w1_0),.din(w_dff_A_2530MqCy4_1),.clk(gclk));
	jdff dff_A_u3ZY1c3w1_0(.dout(w_dff_A_FKw4GYPd0_0),.din(w_dff_A_u3ZY1c3w1_0),.clk(gclk));
	jdff dff_A_FKw4GYPd0_0(.dout(w_dff_A_2dWXPccF2_0),.din(w_dff_A_FKw4GYPd0_0),.clk(gclk));
	jdff dff_A_2dWXPccF2_0(.dout(w_dff_A_Mxelbxml5_0),.din(w_dff_A_2dWXPccF2_0),.clk(gclk));
	jdff dff_A_Mxelbxml5_0(.dout(w_dff_A_2HIeRP1a8_0),.din(w_dff_A_Mxelbxml5_0),.clk(gclk));
	jdff dff_A_2HIeRP1a8_0(.dout(w_dff_A_YSnFNhfn7_0),.din(w_dff_A_2HIeRP1a8_0),.clk(gclk));
	jdff dff_A_YSnFNhfn7_0(.dout(w_dff_A_dGIOdedb0_0),.din(w_dff_A_YSnFNhfn7_0),.clk(gclk));
	jdff dff_A_dGIOdedb0_0(.dout(w_dff_A_5G15qr067_0),.din(w_dff_A_dGIOdedb0_0),.clk(gclk));
	jdff dff_A_5G15qr067_0(.dout(w_dff_A_m6Kg4wvX6_0),.din(w_dff_A_5G15qr067_0),.clk(gclk));
	jdff dff_A_m6Kg4wvX6_0(.dout(w_dff_A_9xIV4Aai7_0),.din(w_dff_A_m6Kg4wvX6_0),.clk(gclk));
	jdff dff_A_9xIV4Aai7_0(.dout(w_dff_A_hP868HXy7_0),.din(w_dff_A_9xIV4Aai7_0),.clk(gclk));
	jdff dff_A_hP868HXy7_0(.dout(w_dff_A_PmkPx5z52_0),.din(w_dff_A_hP868HXy7_0),.clk(gclk));
	jdff dff_A_PmkPx5z52_0(.dout(w_dff_A_7pZIGqW44_0),.din(w_dff_A_PmkPx5z52_0),.clk(gclk));
	jdff dff_A_7pZIGqW44_0(.dout(w_dff_A_8IEzc5wK7_0),.din(w_dff_A_7pZIGqW44_0),.clk(gclk));
	jdff dff_A_8IEzc5wK7_0(.dout(w_dff_A_SUYVqbea4_0),.din(w_dff_A_8IEzc5wK7_0),.clk(gclk));
	jdff dff_A_SUYVqbea4_0(.dout(w_dff_A_yf7d9Imp7_0),.din(w_dff_A_SUYVqbea4_0),.clk(gclk));
	jdff dff_A_yf7d9Imp7_0(.dout(w_dff_A_sRS5qING4_0),.din(w_dff_A_yf7d9Imp7_0),.clk(gclk));
	jdff dff_A_sRS5qING4_0(.dout(w_dff_A_T6eia1x64_0),.din(w_dff_A_sRS5qING4_0),.clk(gclk));
	jdff dff_A_T6eia1x64_0(.dout(w_dff_A_rofsiZJc8_0),.din(w_dff_A_T6eia1x64_0),.clk(gclk));
	jdff dff_A_rofsiZJc8_0(.dout(w_dff_A_ACNn2aBM3_0),.din(w_dff_A_rofsiZJc8_0),.clk(gclk));
	jdff dff_A_ACNn2aBM3_0(.dout(w_dff_A_uMhffgGd6_0),.din(w_dff_A_ACNn2aBM3_0),.clk(gclk));
	jdff dff_A_uMhffgGd6_0(.dout(w_dff_A_AhsZBdRY8_0),.din(w_dff_A_uMhffgGd6_0),.clk(gclk));
	jdff dff_A_AhsZBdRY8_0(.dout(w_dff_A_iv2h2Ekl5_0),.din(w_dff_A_AhsZBdRY8_0),.clk(gclk));
	jdff dff_A_iv2h2Ekl5_0(.dout(w_dff_A_lchCOYYE6_0),.din(w_dff_A_iv2h2Ekl5_0),.clk(gclk));
	jdff dff_A_lchCOYYE6_0(.dout(w_dff_A_QyxtzM7w5_0),.din(w_dff_A_lchCOYYE6_0),.clk(gclk));
	jdff dff_A_QyxtzM7w5_0(.dout(w_dff_A_pgBbFTUJ7_0),.din(w_dff_A_QyxtzM7w5_0),.clk(gclk));
	jdff dff_A_pgBbFTUJ7_0(.dout(w_dff_A_VE8bT0ec1_0),.din(w_dff_A_pgBbFTUJ7_0),.clk(gclk));
	jdff dff_A_VE8bT0ec1_0(.dout(w_dff_A_ULACfosk9_0),.din(w_dff_A_VE8bT0ec1_0),.clk(gclk));
	jdff dff_A_ULACfosk9_0(.dout(w_dff_A_W8pp6NW67_0),.din(w_dff_A_ULACfosk9_0),.clk(gclk));
	jdff dff_A_W8pp6NW67_0(.dout(w_dff_A_5ojiMLSw4_0),.din(w_dff_A_W8pp6NW67_0),.clk(gclk));
	jdff dff_A_5ojiMLSw4_0(.dout(w_dff_A_7kMqU2V71_0),.din(w_dff_A_5ojiMLSw4_0),.clk(gclk));
	jdff dff_A_7kMqU2V71_0(.dout(w_dff_A_bazroMft3_0),.din(w_dff_A_7kMqU2V71_0),.clk(gclk));
	jdff dff_A_bazroMft3_0(.dout(w_dff_A_hI6L4BFx2_0),.din(w_dff_A_bazroMft3_0),.clk(gclk));
	jdff dff_A_hI6L4BFx2_0(.dout(w_dff_A_S71oothp2_0),.din(w_dff_A_hI6L4BFx2_0),.clk(gclk));
	jdff dff_A_S71oothp2_0(.dout(w_dff_A_1au17JYi4_0),.din(w_dff_A_S71oothp2_0),.clk(gclk));
	jdff dff_A_1au17JYi4_0(.dout(w_dff_A_ge44J7sP0_0),.din(w_dff_A_1au17JYi4_0),.clk(gclk));
	jdff dff_A_ge44J7sP0_0(.dout(w_dff_A_7uUriDOv6_0),.din(w_dff_A_ge44J7sP0_0),.clk(gclk));
	jdff dff_A_7uUriDOv6_0(.dout(w_dff_A_8sQcEexO1_0),.din(w_dff_A_7uUriDOv6_0),.clk(gclk));
	jdff dff_A_8sQcEexO1_0(.dout(G480),.din(w_dff_A_8sQcEexO1_0),.clk(gclk));
	jdff dff_A_LItvViFw0_1(.dout(w_dff_A_hEONwuQo9_0),.din(w_dff_A_LItvViFw0_1),.clk(gclk));
	jdff dff_A_hEONwuQo9_0(.dout(w_dff_A_Sup9vN4O5_0),.din(w_dff_A_hEONwuQo9_0),.clk(gclk));
	jdff dff_A_Sup9vN4O5_0(.dout(w_dff_A_owix1sHB2_0),.din(w_dff_A_Sup9vN4O5_0),.clk(gclk));
	jdff dff_A_owix1sHB2_0(.dout(w_dff_A_RzDwBfp12_0),.din(w_dff_A_owix1sHB2_0),.clk(gclk));
	jdff dff_A_RzDwBfp12_0(.dout(w_dff_A_m5KEiS5a3_0),.din(w_dff_A_RzDwBfp12_0),.clk(gclk));
	jdff dff_A_m5KEiS5a3_0(.dout(w_dff_A_T6Tluu1o6_0),.din(w_dff_A_m5KEiS5a3_0),.clk(gclk));
	jdff dff_A_T6Tluu1o6_0(.dout(w_dff_A_82rB9WJf6_0),.din(w_dff_A_T6Tluu1o6_0),.clk(gclk));
	jdff dff_A_82rB9WJf6_0(.dout(w_dff_A_JfPR4Bnq9_0),.din(w_dff_A_82rB9WJf6_0),.clk(gclk));
	jdff dff_A_JfPR4Bnq9_0(.dout(w_dff_A_KrnNDBXj2_0),.din(w_dff_A_JfPR4Bnq9_0),.clk(gclk));
	jdff dff_A_KrnNDBXj2_0(.dout(w_dff_A_HKzJ4Kr05_0),.din(w_dff_A_KrnNDBXj2_0),.clk(gclk));
	jdff dff_A_HKzJ4Kr05_0(.dout(w_dff_A_2z7kxOfK8_0),.din(w_dff_A_HKzJ4Kr05_0),.clk(gclk));
	jdff dff_A_2z7kxOfK8_0(.dout(w_dff_A_tXpRaclm5_0),.din(w_dff_A_2z7kxOfK8_0),.clk(gclk));
	jdff dff_A_tXpRaclm5_0(.dout(w_dff_A_56rCdv0G7_0),.din(w_dff_A_tXpRaclm5_0),.clk(gclk));
	jdff dff_A_56rCdv0G7_0(.dout(w_dff_A_idQtLsYp5_0),.din(w_dff_A_56rCdv0G7_0),.clk(gclk));
	jdff dff_A_idQtLsYp5_0(.dout(w_dff_A_PTbWvBUr4_0),.din(w_dff_A_idQtLsYp5_0),.clk(gclk));
	jdff dff_A_PTbWvBUr4_0(.dout(w_dff_A_oiwUN3C77_0),.din(w_dff_A_PTbWvBUr4_0),.clk(gclk));
	jdff dff_A_oiwUN3C77_0(.dout(w_dff_A_EKyhdG104_0),.din(w_dff_A_oiwUN3C77_0),.clk(gclk));
	jdff dff_A_EKyhdG104_0(.dout(w_dff_A_HteDVVk90_0),.din(w_dff_A_EKyhdG104_0),.clk(gclk));
	jdff dff_A_HteDVVk90_0(.dout(w_dff_A_PjyJv4ia5_0),.din(w_dff_A_HteDVVk90_0),.clk(gclk));
	jdff dff_A_PjyJv4ia5_0(.dout(w_dff_A_qsz4TLkT1_0),.din(w_dff_A_PjyJv4ia5_0),.clk(gclk));
	jdff dff_A_qsz4TLkT1_0(.dout(w_dff_A_TBilviF56_0),.din(w_dff_A_qsz4TLkT1_0),.clk(gclk));
	jdff dff_A_TBilviF56_0(.dout(w_dff_A_5Hc8v8rE9_0),.din(w_dff_A_TBilviF56_0),.clk(gclk));
	jdff dff_A_5Hc8v8rE9_0(.dout(w_dff_A_ew6xvEHu8_0),.din(w_dff_A_5Hc8v8rE9_0),.clk(gclk));
	jdff dff_A_ew6xvEHu8_0(.dout(w_dff_A_NxL9531h2_0),.din(w_dff_A_ew6xvEHu8_0),.clk(gclk));
	jdff dff_A_NxL9531h2_0(.dout(w_dff_A_W2Baw9qX6_0),.din(w_dff_A_NxL9531h2_0),.clk(gclk));
	jdff dff_A_W2Baw9qX6_0(.dout(w_dff_A_hV6JXWaV1_0),.din(w_dff_A_W2Baw9qX6_0),.clk(gclk));
	jdff dff_A_hV6JXWaV1_0(.dout(w_dff_A_SFVzwpxV7_0),.din(w_dff_A_hV6JXWaV1_0),.clk(gclk));
	jdff dff_A_SFVzwpxV7_0(.dout(w_dff_A_fioC63og8_0),.din(w_dff_A_SFVzwpxV7_0),.clk(gclk));
	jdff dff_A_fioC63og8_0(.dout(w_dff_A_2D4uhXIu5_0),.din(w_dff_A_fioC63og8_0),.clk(gclk));
	jdff dff_A_2D4uhXIu5_0(.dout(w_dff_A_SeTkpVWa2_0),.din(w_dff_A_2D4uhXIu5_0),.clk(gclk));
	jdff dff_A_SeTkpVWa2_0(.dout(w_dff_A_gTkDgGKf8_0),.din(w_dff_A_SeTkpVWa2_0),.clk(gclk));
	jdff dff_A_gTkDgGKf8_0(.dout(w_dff_A_6Zc7PEBQ8_0),.din(w_dff_A_gTkDgGKf8_0),.clk(gclk));
	jdff dff_A_6Zc7PEBQ8_0(.dout(w_dff_A_XsDY4orp4_0),.din(w_dff_A_6Zc7PEBQ8_0),.clk(gclk));
	jdff dff_A_XsDY4orp4_0(.dout(w_dff_A_edTETl5E2_0),.din(w_dff_A_XsDY4orp4_0),.clk(gclk));
	jdff dff_A_edTETl5E2_0(.dout(w_dff_A_RbL5fwkj5_0),.din(w_dff_A_edTETl5E2_0),.clk(gclk));
	jdff dff_A_RbL5fwkj5_0(.dout(w_dff_A_U06ymaAX7_0),.din(w_dff_A_RbL5fwkj5_0),.clk(gclk));
	jdff dff_A_U06ymaAX7_0(.dout(w_dff_A_pnwIKx1Y2_0),.din(w_dff_A_U06ymaAX7_0),.clk(gclk));
	jdff dff_A_pnwIKx1Y2_0(.dout(w_dff_A_YjjJQKyr1_0),.din(w_dff_A_pnwIKx1Y2_0),.clk(gclk));
	jdff dff_A_YjjJQKyr1_0(.dout(G560),.din(w_dff_A_YjjJQKyr1_0),.clk(gclk));
	jdff dff_A_vnhaT5SN9_1(.dout(w_dff_A_G9tMNoQa9_0),.din(w_dff_A_vnhaT5SN9_1),.clk(gclk));
	jdff dff_A_G9tMNoQa9_0(.dout(w_dff_A_omjDHzPE6_0),.din(w_dff_A_G9tMNoQa9_0),.clk(gclk));
	jdff dff_A_omjDHzPE6_0(.dout(w_dff_A_eLKOlVg81_0),.din(w_dff_A_omjDHzPE6_0),.clk(gclk));
	jdff dff_A_eLKOlVg81_0(.dout(w_dff_A_oNeJbNLr0_0),.din(w_dff_A_eLKOlVg81_0),.clk(gclk));
	jdff dff_A_oNeJbNLr0_0(.dout(w_dff_A_w8jiqpA43_0),.din(w_dff_A_oNeJbNLr0_0),.clk(gclk));
	jdff dff_A_w8jiqpA43_0(.dout(w_dff_A_L9fEAcTQ1_0),.din(w_dff_A_w8jiqpA43_0),.clk(gclk));
	jdff dff_A_L9fEAcTQ1_0(.dout(w_dff_A_Wuql2Nan2_0),.din(w_dff_A_L9fEAcTQ1_0),.clk(gclk));
	jdff dff_A_Wuql2Nan2_0(.dout(w_dff_A_c5Cq1KLm0_0),.din(w_dff_A_Wuql2Nan2_0),.clk(gclk));
	jdff dff_A_c5Cq1KLm0_0(.dout(w_dff_A_FtI0Pbei6_0),.din(w_dff_A_c5Cq1KLm0_0),.clk(gclk));
	jdff dff_A_FtI0Pbei6_0(.dout(w_dff_A_PmH1NPZn3_0),.din(w_dff_A_FtI0Pbei6_0),.clk(gclk));
	jdff dff_A_PmH1NPZn3_0(.dout(w_dff_A_qBjKAfGX9_0),.din(w_dff_A_PmH1NPZn3_0),.clk(gclk));
	jdff dff_A_qBjKAfGX9_0(.dout(w_dff_A_Wad7dzZ72_0),.din(w_dff_A_qBjKAfGX9_0),.clk(gclk));
	jdff dff_A_Wad7dzZ72_0(.dout(w_dff_A_LEBHHY8y6_0),.din(w_dff_A_Wad7dzZ72_0),.clk(gclk));
	jdff dff_A_LEBHHY8y6_0(.dout(w_dff_A_7VEdD81l7_0),.din(w_dff_A_LEBHHY8y6_0),.clk(gclk));
	jdff dff_A_7VEdD81l7_0(.dout(w_dff_A_Hes6odD83_0),.din(w_dff_A_7VEdD81l7_0),.clk(gclk));
	jdff dff_A_Hes6odD83_0(.dout(w_dff_A_ewM9UXo09_0),.din(w_dff_A_Hes6odD83_0),.clk(gclk));
	jdff dff_A_ewM9UXo09_0(.dout(w_dff_A_6EZDpP983_0),.din(w_dff_A_ewM9UXo09_0),.clk(gclk));
	jdff dff_A_6EZDpP983_0(.dout(w_dff_A_lPteOT4K6_0),.din(w_dff_A_6EZDpP983_0),.clk(gclk));
	jdff dff_A_lPteOT4K6_0(.dout(w_dff_A_G0J0sIXi6_0),.din(w_dff_A_lPteOT4K6_0),.clk(gclk));
	jdff dff_A_G0J0sIXi6_0(.dout(w_dff_A_M4Q3ZGpu8_0),.din(w_dff_A_G0J0sIXi6_0),.clk(gclk));
	jdff dff_A_M4Q3ZGpu8_0(.dout(w_dff_A_68M00IZ28_0),.din(w_dff_A_M4Q3ZGpu8_0),.clk(gclk));
	jdff dff_A_68M00IZ28_0(.dout(w_dff_A_1QHzNTzL8_0),.din(w_dff_A_68M00IZ28_0),.clk(gclk));
	jdff dff_A_1QHzNTzL8_0(.dout(w_dff_A_ZMmhDyv55_0),.din(w_dff_A_1QHzNTzL8_0),.clk(gclk));
	jdff dff_A_ZMmhDyv55_0(.dout(w_dff_A_pi1Tr7P82_0),.din(w_dff_A_ZMmhDyv55_0),.clk(gclk));
	jdff dff_A_pi1Tr7P82_0(.dout(w_dff_A_ip5Ey8nq0_0),.din(w_dff_A_pi1Tr7P82_0),.clk(gclk));
	jdff dff_A_ip5Ey8nq0_0(.dout(w_dff_A_j5kHKfiM9_0),.din(w_dff_A_ip5Ey8nq0_0),.clk(gclk));
	jdff dff_A_j5kHKfiM9_0(.dout(w_dff_A_eLn2iFOw5_0),.din(w_dff_A_j5kHKfiM9_0),.clk(gclk));
	jdff dff_A_eLn2iFOw5_0(.dout(w_dff_A_LSff1cIb9_0),.din(w_dff_A_eLn2iFOw5_0),.clk(gclk));
	jdff dff_A_LSff1cIb9_0(.dout(w_dff_A_XCbC5SHI0_0),.din(w_dff_A_LSff1cIb9_0),.clk(gclk));
	jdff dff_A_XCbC5SHI0_0(.dout(w_dff_A_z3hAff878_0),.din(w_dff_A_XCbC5SHI0_0),.clk(gclk));
	jdff dff_A_z3hAff878_0(.dout(w_dff_A_QGjGK16B2_0),.din(w_dff_A_z3hAff878_0),.clk(gclk));
	jdff dff_A_QGjGK16B2_0(.dout(w_dff_A_brRFeKfR2_0),.din(w_dff_A_QGjGK16B2_0),.clk(gclk));
	jdff dff_A_brRFeKfR2_0(.dout(w_dff_A_KkmY2knc5_0),.din(w_dff_A_brRFeKfR2_0),.clk(gclk));
	jdff dff_A_KkmY2knc5_0(.dout(w_dff_A_BaWrWveG5_0),.din(w_dff_A_KkmY2knc5_0),.clk(gclk));
	jdff dff_A_BaWrWveG5_0(.dout(w_dff_A_NZQMJ2Hb8_0),.din(w_dff_A_BaWrWveG5_0),.clk(gclk));
	jdff dff_A_NZQMJ2Hb8_0(.dout(w_dff_A_BAMtfML29_0),.din(w_dff_A_NZQMJ2Hb8_0),.clk(gclk));
	jdff dff_A_BAMtfML29_0(.dout(w_dff_A_7MQyo9mS8_0),.din(w_dff_A_BAMtfML29_0),.clk(gclk));
	jdff dff_A_7MQyo9mS8_0(.dout(w_dff_A_IKXSTLAS2_0),.din(w_dff_A_7MQyo9mS8_0),.clk(gclk));
	jdff dff_A_IKXSTLAS2_0(.dout(G542),.din(w_dff_A_IKXSTLAS2_0),.clk(gclk));
	jdff dff_A_LUDcVW948_1(.dout(w_dff_A_X9YYyhJt4_0),.din(w_dff_A_LUDcVW948_1),.clk(gclk));
	jdff dff_A_X9YYyhJt4_0(.dout(w_dff_A_dfLPMELM5_0),.din(w_dff_A_X9YYyhJt4_0),.clk(gclk));
	jdff dff_A_dfLPMELM5_0(.dout(w_dff_A_WBm55wzQ7_0),.din(w_dff_A_dfLPMELM5_0),.clk(gclk));
	jdff dff_A_WBm55wzQ7_0(.dout(w_dff_A_qund6fSy6_0),.din(w_dff_A_WBm55wzQ7_0),.clk(gclk));
	jdff dff_A_qund6fSy6_0(.dout(w_dff_A_kbMK0lRx7_0),.din(w_dff_A_qund6fSy6_0),.clk(gclk));
	jdff dff_A_kbMK0lRx7_0(.dout(w_dff_A_jfdW6br75_0),.din(w_dff_A_kbMK0lRx7_0),.clk(gclk));
	jdff dff_A_jfdW6br75_0(.dout(w_dff_A_bTQNog3I2_0),.din(w_dff_A_jfdW6br75_0),.clk(gclk));
	jdff dff_A_bTQNog3I2_0(.dout(w_dff_A_8pSMHK1a6_0),.din(w_dff_A_bTQNog3I2_0),.clk(gclk));
	jdff dff_A_8pSMHK1a6_0(.dout(w_dff_A_xgzBJHGm1_0),.din(w_dff_A_8pSMHK1a6_0),.clk(gclk));
	jdff dff_A_xgzBJHGm1_0(.dout(w_dff_A_hU2l9HEg1_0),.din(w_dff_A_xgzBJHGm1_0),.clk(gclk));
	jdff dff_A_hU2l9HEg1_0(.dout(w_dff_A_D3qznDfe4_0),.din(w_dff_A_hU2l9HEg1_0),.clk(gclk));
	jdff dff_A_D3qznDfe4_0(.dout(w_dff_A_JTWzKiJT7_0),.din(w_dff_A_D3qznDfe4_0),.clk(gclk));
	jdff dff_A_JTWzKiJT7_0(.dout(w_dff_A_sRxDq0wE5_0),.din(w_dff_A_JTWzKiJT7_0),.clk(gclk));
	jdff dff_A_sRxDq0wE5_0(.dout(w_dff_A_xu2u7iYx8_0),.din(w_dff_A_sRxDq0wE5_0),.clk(gclk));
	jdff dff_A_xu2u7iYx8_0(.dout(w_dff_A_HX08QI1R4_0),.din(w_dff_A_xu2u7iYx8_0),.clk(gclk));
	jdff dff_A_HX08QI1R4_0(.dout(w_dff_A_W7tll8Kn7_0),.din(w_dff_A_HX08QI1R4_0),.clk(gclk));
	jdff dff_A_W7tll8Kn7_0(.dout(w_dff_A_w6Uqyi141_0),.din(w_dff_A_W7tll8Kn7_0),.clk(gclk));
	jdff dff_A_w6Uqyi141_0(.dout(w_dff_A_UxCJXwjV5_0),.din(w_dff_A_w6Uqyi141_0),.clk(gclk));
	jdff dff_A_UxCJXwjV5_0(.dout(w_dff_A_znO0lCOk1_0),.din(w_dff_A_UxCJXwjV5_0),.clk(gclk));
	jdff dff_A_znO0lCOk1_0(.dout(w_dff_A_05UaASIe7_0),.din(w_dff_A_znO0lCOk1_0),.clk(gclk));
	jdff dff_A_05UaASIe7_0(.dout(w_dff_A_Yb3OQUze3_0),.din(w_dff_A_05UaASIe7_0),.clk(gclk));
	jdff dff_A_Yb3OQUze3_0(.dout(w_dff_A_MLoAZUGu2_0),.din(w_dff_A_Yb3OQUze3_0),.clk(gclk));
	jdff dff_A_MLoAZUGu2_0(.dout(w_dff_A_HGdACXJw5_0),.din(w_dff_A_MLoAZUGu2_0),.clk(gclk));
	jdff dff_A_HGdACXJw5_0(.dout(w_dff_A_wAlFokZx2_0),.din(w_dff_A_HGdACXJw5_0),.clk(gclk));
	jdff dff_A_wAlFokZx2_0(.dout(w_dff_A_84w4AuBQ4_0),.din(w_dff_A_wAlFokZx2_0),.clk(gclk));
	jdff dff_A_84w4AuBQ4_0(.dout(w_dff_A_v8wXJQ4y2_0),.din(w_dff_A_84w4AuBQ4_0),.clk(gclk));
	jdff dff_A_v8wXJQ4y2_0(.dout(w_dff_A_F5wxTxZB3_0),.din(w_dff_A_v8wXJQ4y2_0),.clk(gclk));
	jdff dff_A_F5wxTxZB3_0(.dout(w_dff_A_wk8UXeRf8_0),.din(w_dff_A_F5wxTxZB3_0),.clk(gclk));
	jdff dff_A_wk8UXeRf8_0(.dout(w_dff_A_HS9Bc7a39_0),.din(w_dff_A_wk8UXeRf8_0),.clk(gclk));
	jdff dff_A_HS9Bc7a39_0(.dout(w_dff_A_2TsYyfjP2_0),.din(w_dff_A_HS9Bc7a39_0),.clk(gclk));
	jdff dff_A_2TsYyfjP2_0(.dout(w_dff_A_a4Pl5pdD8_0),.din(w_dff_A_2TsYyfjP2_0),.clk(gclk));
	jdff dff_A_a4Pl5pdD8_0(.dout(w_dff_A_rJrvrkpQ6_0),.din(w_dff_A_a4Pl5pdD8_0),.clk(gclk));
	jdff dff_A_rJrvrkpQ6_0(.dout(w_dff_A_7hE47G178_0),.din(w_dff_A_rJrvrkpQ6_0),.clk(gclk));
	jdff dff_A_7hE47G178_0(.dout(w_dff_A_Dzu1FWcg0_0),.din(w_dff_A_7hE47G178_0),.clk(gclk));
	jdff dff_A_Dzu1FWcg0_0(.dout(w_dff_A_WKTmC0dz8_0),.din(w_dff_A_Dzu1FWcg0_0),.clk(gclk));
	jdff dff_A_WKTmC0dz8_0(.dout(w_dff_A_GS4gIo068_0),.din(w_dff_A_WKTmC0dz8_0),.clk(gclk));
	jdff dff_A_GS4gIo068_0(.dout(w_dff_A_klrKteQO1_0),.din(w_dff_A_GS4gIo068_0),.clk(gclk));
	jdff dff_A_klrKteQO1_0(.dout(w_dff_A_i2I4SPfK6_0),.din(w_dff_A_klrKteQO1_0),.clk(gclk));
	jdff dff_A_i2I4SPfK6_0(.dout(G558),.din(w_dff_A_i2I4SPfK6_0),.clk(gclk));
	jdff dff_A_YgGp9OAD8_1(.dout(w_dff_A_0QlK25Ds0_0),.din(w_dff_A_YgGp9OAD8_1),.clk(gclk));
	jdff dff_A_0QlK25Ds0_0(.dout(w_dff_A_zIPE5OUr0_0),.din(w_dff_A_0QlK25Ds0_0),.clk(gclk));
	jdff dff_A_zIPE5OUr0_0(.dout(w_dff_A_uaGCy09q6_0),.din(w_dff_A_zIPE5OUr0_0),.clk(gclk));
	jdff dff_A_uaGCy09q6_0(.dout(w_dff_A_GwBIRKze0_0),.din(w_dff_A_uaGCy09q6_0),.clk(gclk));
	jdff dff_A_GwBIRKze0_0(.dout(w_dff_A_EE7qzUBt2_0),.din(w_dff_A_GwBIRKze0_0),.clk(gclk));
	jdff dff_A_EE7qzUBt2_0(.dout(w_dff_A_3Sn0e4Ym4_0),.din(w_dff_A_EE7qzUBt2_0),.clk(gclk));
	jdff dff_A_3Sn0e4Ym4_0(.dout(w_dff_A_i515ZKvw2_0),.din(w_dff_A_3Sn0e4Ym4_0),.clk(gclk));
	jdff dff_A_i515ZKvw2_0(.dout(w_dff_A_Bf7dUFB88_0),.din(w_dff_A_i515ZKvw2_0),.clk(gclk));
	jdff dff_A_Bf7dUFB88_0(.dout(w_dff_A_LQzbzHAh7_0),.din(w_dff_A_Bf7dUFB88_0),.clk(gclk));
	jdff dff_A_LQzbzHAh7_0(.dout(w_dff_A_3kC3B4rI8_0),.din(w_dff_A_LQzbzHAh7_0),.clk(gclk));
	jdff dff_A_3kC3B4rI8_0(.dout(w_dff_A_NQmCufV21_0),.din(w_dff_A_3kC3B4rI8_0),.clk(gclk));
	jdff dff_A_NQmCufV21_0(.dout(w_dff_A_iT40sNiM0_0),.din(w_dff_A_NQmCufV21_0),.clk(gclk));
	jdff dff_A_iT40sNiM0_0(.dout(w_dff_A_gkCiHrCh7_0),.din(w_dff_A_iT40sNiM0_0),.clk(gclk));
	jdff dff_A_gkCiHrCh7_0(.dout(w_dff_A_BKY44R154_0),.din(w_dff_A_gkCiHrCh7_0),.clk(gclk));
	jdff dff_A_BKY44R154_0(.dout(w_dff_A_zb4o4c8M6_0),.din(w_dff_A_BKY44R154_0),.clk(gclk));
	jdff dff_A_zb4o4c8M6_0(.dout(w_dff_A_SJtMSAf81_0),.din(w_dff_A_zb4o4c8M6_0),.clk(gclk));
	jdff dff_A_SJtMSAf81_0(.dout(w_dff_A_KflnuDOR8_0),.din(w_dff_A_SJtMSAf81_0),.clk(gclk));
	jdff dff_A_KflnuDOR8_0(.dout(w_dff_A_i8eqpaAh1_0),.din(w_dff_A_KflnuDOR8_0),.clk(gclk));
	jdff dff_A_i8eqpaAh1_0(.dout(w_dff_A_UXEqZ9wj2_0),.din(w_dff_A_i8eqpaAh1_0),.clk(gclk));
	jdff dff_A_UXEqZ9wj2_0(.dout(w_dff_A_ySpLjSze5_0),.din(w_dff_A_UXEqZ9wj2_0),.clk(gclk));
	jdff dff_A_ySpLjSze5_0(.dout(w_dff_A_05agX0Ev1_0),.din(w_dff_A_ySpLjSze5_0),.clk(gclk));
	jdff dff_A_05agX0Ev1_0(.dout(w_dff_A_F5elunu49_0),.din(w_dff_A_05agX0Ev1_0),.clk(gclk));
	jdff dff_A_F5elunu49_0(.dout(w_dff_A_XtB4WoBz8_0),.din(w_dff_A_F5elunu49_0),.clk(gclk));
	jdff dff_A_XtB4WoBz8_0(.dout(w_dff_A_S6EMwAXX9_0),.din(w_dff_A_XtB4WoBz8_0),.clk(gclk));
	jdff dff_A_S6EMwAXX9_0(.dout(w_dff_A_nGSzjTJM9_0),.din(w_dff_A_S6EMwAXX9_0),.clk(gclk));
	jdff dff_A_nGSzjTJM9_0(.dout(w_dff_A_emgDBOkS0_0),.din(w_dff_A_nGSzjTJM9_0),.clk(gclk));
	jdff dff_A_emgDBOkS0_0(.dout(w_dff_A_ecjFM3G38_0),.din(w_dff_A_emgDBOkS0_0),.clk(gclk));
	jdff dff_A_ecjFM3G38_0(.dout(w_dff_A_nhhOIW3N3_0),.din(w_dff_A_ecjFM3G38_0),.clk(gclk));
	jdff dff_A_nhhOIW3N3_0(.dout(w_dff_A_Ag1zIeCj0_0),.din(w_dff_A_nhhOIW3N3_0),.clk(gclk));
	jdff dff_A_Ag1zIeCj0_0(.dout(w_dff_A_1VwfO0Fo5_0),.din(w_dff_A_Ag1zIeCj0_0),.clk(gclk));
	jdff dff_A_1VwfO0Fo5_0(.dout(w_dff_A_45jw5LT38_0),.din(w_dff_A_1VwfO0Fo5_0),.clk(gclk));
	jdff dff_A_45jw5LT38_0(.dout(w_dff_A_FmChxGpk6_0),.din(w_dff_A_45jw5LT38_0),.clk(gclk));
	jdff dff_A_FmChxGpk6_0(.dout(w_dff_A_JCxyAt8p3_0),.din(w_dff_A_FmChxGpk6_0),.clk(gclk));
	jdff dff_A_JCxyAt8p3_0(.dout(w_dff_A_4SCFmmLB0_0),.din(w_dff_A_JCxyAt8p3_0),.clk(gclk));
	jdff dff_A_4SCFmmLB0_0(.dout(w_dff_A_eMK9UIsO4_0),.din(w_dff_A_4SCFmmLB0_0),.clk(gclk));
	jdff dff_A_eMK9UIsO4_0(.dout(w_dff_A_6UmeON7q0_0),.din(w_dff_A_eMK9UIsO4_0),.clk(gclk));
	jdff dff_A_6UmeON7q0_0(.dout(w_dff_A_0nYxeyv95_0),.din(w_dff_A_6UmeON7q0_0),.clk(gclk));
	jdff dff_A_0nYxeyv95_0(.dout(w_dff_A_GY6VqlmW0_0),.din(w_dff_A_0nYxeyv95_0),.clk(gclk));
	jdff dff_A_GY6VqlmW0_0(.dout(G556),.din(w_dff_A_GY6VqlmW0_0),.clk(gclk));
	jdff dff_A_0NogE0yY4_1(.dout(w_dff_A_Nvdx9tAO0_0),.din(w_dff_A_0NogE0yY4_1),.clk(gclk));
	jdff dff_A_Nvdx9tAO0_0(.dout(w_dff_A_Ott9JlcE6_0),.din(w_dff_A_Nvdx9tAO0_0),.clk(gclk));
	jdff dff_A_Ott9JlcE6_0(.dout(w_dff_A_kzTENg772_0),.din(w_dff_A_Ott9JlcE6_0),.clk(gclk));
	jdff dff_A_kzTENg772_0(.dout(w_dff_A_LCANN16k2_0),.din(w_dff_A_kzTENg772_0),.clk(gclk));
	jdff dff_A_LCANN16k2_0(.dout(w_dff_A_Lkyqgqbx3_0),.din(w_dff_A_LCANN16k2_0),.clk(gclk));
	jdff dff_A_Lkyqgqbx3_0(.dout(w_dff_A_zu0QWtS43_0),.din(w_dff_A_Lkyqgqbx3_0),.clk(gclk));
	jdff dff_A_zu0QWtS43_0(.dout(w_dff_A_OGLDDCL70_0),.din(w_dff_A_zu0QWtS43_0),.clk(gclk));
	jdff dff_A_OGLDDCL70_0(.dout(w_dff_A_z6yUUIVR2_0),.din(w_dff_A_OGLDDCL70_0),.clk(gclk));
	jdff dff_A_z6yUUIVR2_0(.dout(w_dff_A_GBbJVQwi5_0),.din(w_dff_A_z6yUUIVR2_0),.clk(gclk));
	jdff dff_A_GBbJVQwi5_0(.dout(w_dff_A_8DZfy4kQ5_0),.din(w_dff_A_GBbJVQwi5_0),.clk(gclk));
	jdff dff_A_8DZfy4kQ5_0(.dout(w_dff_A_RjhtBDwM8_0),.din(w_dff_A_8DZfy4kQ5_0),.clk(gclk));
	jdff dff_A_RjhtBDwM8_0(.dout(w_dff_A_CdEYTqNb2_0),.din(w_dff_A_RjhtBDwM8_0),.clk(gclk));
	jdff dff_A_CdEYTqNb2_0(.dout(w_dff_A_evSR5vPu2_0),.din(w_dff_A_CdEYTqNb2_0),.clk(gclk));
	jdff dff_A_evSR5vPu2_0(.dout(w_dff_A_0gEGOtzx8_0),.din(w_dff_A_evSR5vPu2_0),.clk(gclk));
	jdff dff_A_0gEGOtzx8_0(.dout(w_dff_A_bFOhM57K2_0),.din(w_dff_A_0gEGOtzx8_0),.clk(gclk));
	jdff dff_A_bFOhM57K2_0(.dout(w_dff_A_IwRwMLat5_0),.din(w_dff_A_bFOhM57K2_0),.clk(gclk));
	jdff dff_A_IwRwMLat5_0(.dout(w_dff_A_FafZDnee1_0),.din(w_dff_A_IwRwMLat5_0),.clk(gclk));
	jdff dff_A_FafZDnee1_0(.dout(w_dff_A_Hzm2QZ7G8_0),.din(w_dff_A_FafZDnee1_0),.clk(gclk));
	jdff dff_A_Hzm2QZ7G8_0(.dout(w_dff_A_VKymOSal2_0),.din(w_dff_A_Hzm2QZ7G8_0),.clk(gclk));
	jdff dff_A_VKymOSal2_0(.dout(w_dff_A_PorutfbF3_0),.din(w_dff_A_VKymOSal2_0),.clk(gclk));
	jdff dff_A_PorutfbF3_0(.dout(w_dff_A_qJeIaSCR4_0),.din(w_dff_A_PorutfbF3_0),.clk(gclk));
	jdff dff_A_qJeIaSCR4_0(.dout(w_dff_A_234ifCIy2_0),.din(w_dff_A_qJeIaSCR4_0),.clk(gclk));
	jdff dff_A_234ifCIy2_0(.dout(w_dff_A_3zfAX6XL4_0),.din(w_dff_A_234ifCIy2_0),.clk(gclk));
	jdff dff_A_3zfAX6XL4_0(.dout(w_dff_A_9a46uQbX8_0),.din(w_dff_A_3zfAX6XL4_0),.clk(gclk));
	jdff dff_A_9a46uQbX8_0(.dout(w_dff_A_fgPiidmh7_0),.din(w_dff_A_9a46uQbX8_0),.clk(gclk));
	jdff dff_A_fgPiidmh7_0(.dout(w_dff_A_knJEV6iV6_0),.din(w_dff_A_fgPiidmh7_0),.clk(gclk));
	jdff dff_A_knJEV6iV6_0(.dout(w_dff_A_ZDYYDH1t9_0),.din(w_dff_A_knJEV6iV6_0),.clk(gclk));
	jdff dff_A_ZDYYDH1t9_0(.dout(w_dff_A_PeQX62QY1_0),.din(w_dff_A_ZDYYDH1t9_0),.clk(gclk));
	jdff dff_A_PeQX62QY1_0(.dout(w_dff_A_16dSxHqO9_0),.din(w_dff_A_PeQX62QY1_0),.clk(gclk));
	jdff dff_A_16dSxHqO9_0(.dout(w_dff_A_xOsVZGl18_0),.din(w_dff_A_16dSxHqO9_0),.clk(gclk));
	jdff dff_A_xOsVZGl18_0(.dout(w_dff_A_0BcjZkzi9_0),.din(w_dff_A_xOsVZGl18_0),.clk(gclk));
	jdff dff_A_0BcjZkzi9_0(.dout(w_dff_A_gFbqdkQx3_0),.din(w_dff_A_0BcjZkzi9_0),.clk(gclk));
	jdff dff_A_gFbqdkQx3_0(.dout(w_dff_A_bRh5qoeL9_0),.din(w_dff_A_gFbqdkQx3_0),.clk(gclk));
	jdff dff_A_bRh5qoeL9_0(.dout(w_dff_A_nhbAUFk49_0),.din(w_dff_A_bRh5qoeL9_0),.clk(gclk));
	jdff dff_A_nhbAUFk49_0(.dout(w_dff_A_WZGRpOHd1_0),.din(w_dff_A_nhbAUFk49_0),.clk(gclk));
	jdff dff_A_WZGRpOHd1_0(.dout(w_dff_A_P9H4QUlG4_0),.din(w_dff_A_WZGRpOHd1_0),.clk(gclk));
	jdff dff_A_P9H4QUlG4_0(.dout(w_dff_A_zkyjy38M1_0),.din(w_dff_A_P9H4QUlG4_0),.clk(gclk));
	jdff dff_A_zkyjy38M1_0(.dout(w_dff_A_yETswr8r4_0),.din(w_dff_A_zkyjy38M1_0),.clk(gclk));
	jdff dff_A_yETswr8r4_0(.dout(G554),.din(w_dff_A_yETswr8r4_0),.clk(gclk));
	jdff dff_A_B1CtAN1E0_1(.dout(w_dff_A_x0z06xRE3_0),.din(w_dff_A_B1CtAN1E0_1),.clk(gclk));
	jdff dff_A_x0z06xRE3_0(.dout(w_dff_A_RFDGyIYF6_0),.din(w_dff_A_x0z06xRE3_0),.clk(gclk));
	jdff dff_A_RFDGyIYF6_0(.dout(w_dff_A_QEehQPA88_0),.din(w_dff_A_RFDGyIYF6_0),.clk(gclk));
	jdff dff_A_QEehQPA88_0(.dout(w_dff_A_qrPugM7A5_0),.din(w_dff_A_QEehQPA88_0),.clk(gclk));
	jdff dff_A_qrPugM7A5_0(.dout(w_dff_A_UAMn1Up06_0),.din(w_dff_A_qrPugM7A5_0),.clk(gclk));
	jdff dff_A_UAMn1Up06_0(.dout(w_dff_A_gMuqVDUc9_0),.din(w_dff_A_UAMn1Up06_0),.clk(gclk));
	jdff dff_A_gMuqVDUc9_0(.dout(w_dff_A_aUGvikyU2_0),.din(w_dff_A_gMuqVDUc9_0),.clk(gclk));
	jdff dff_A_aUGvikyU2_0(.dout(w_dff_A_FiS1OJIh8_0),.din(w_dff_A_aUGvikyU2_0),.clk(gclk));
	jdff dff_A_FiS1OJIh8_0(.dout(w_dff_A_Zl9N27pS1_0),.din(w_dff_A_FiS1OJIh8_0),.clk(gclk));
	jdff dff_A_Zl9N27pS1_0(.dout(w_dff_A_6a4R9skz6_0),.din(w_dff_A_Zl9N27pS1_0),.clk(gclk));
	jdff dff_A_6a4R9skz6_0(.dout(w_dff_A_ysZsao199_0),.din(w_dff_A_6a4R9skz6_0),.clk(gclk));
	jdff dff_A_ysZsao199_0(.dout(w_dff_A_C2rjcaTl9_0),.din(w_dff_A_ysZsao199_0),.clk(gclk));
	jdff dff_A_C2rjcaTl9_0(.dout(w_dff_A_jeNX7dG11_0),.din(w_dff_A_C2rjcaTl9_0),.clk(gclk));
	jdff dff_A_jeNX7dG11_0(.dout(w_dff_A_7xhBNyUp1_0),.din(w_dff_A_jeNX7dG11_0),.clk(gclk));
	jdff dff_A_7xhBNyUp1_0(.dout(w_dff_A_190ctC065_0),.din(w_dff_A_7xhBNyUp1_0),.clk(gclk));
	jdff dff_A_190ctC065_0(.dout(w_dff_A_eTZUHcvB5_0),.din(w_dff_A_190ctC065_0),.clk(gclk));
	jdff dff_A_eTZUHcvB5_0(.dout(w_dff_A_5mB3WdhG2_0),.din(w_dff_A_eTZUHcvB5_0),.clk(gclk));
	jdff dff_A_5mB3WdhG2_0(.dout(w_dff_A_geMJTZzl9_0),.din(w_dff_A_5mB3WdhG2_0),.clk(gclk));
	jdff dff_A_geMJTZzl9_0(.dout(w_dff_A_s3bH4qku5_0),.din(w_dff_A_geMJTZzl9_0),.clk(gclk));
	jdff dff_A_s3bH4qku5_0(.dout(w_dff_A_1ce1HdOi2_0),.din(w_dff_A_s3bH4qku5_0),.clk(gclk));
	jdff dff_A_1ce1HdOi2_0(.dout(w_dff_A_ADOZWDe22_0),.din(w_dff_A_1ce1HdOi2_0),.clk(gclk));
	jdff dff_A_ADOZWDe22_0(.dout(w_dff_A_WvcocX5X9_0),.din(w_dff_A_ADOZWDe22_0),.clk(gclk));
	jdff dff_A_WvcocX5X9_0(.dout(w_dff_A_SbKRXqAB1_0),.din(w_dff_A_WvcocX5X9_0),.clk(gclk));
	jdff dff_A_SbKRXqAB1_0(.dout(w_dff_A_wLr2L8Pe8_0),.din(w_dff_A_SbKRXqAB1_0),.clk(gclk));
	jdff dff_A_wLr2L8Pe8_0(.dout(w_dff_A_aVeR2SgY8_0),.din(w_dff_A_wLr2L8Pe8_0),.clk(gclk));
	jdff dff_A_aVeR2SgY8_0(.dout(w_dff_A_qN2rgI7h4_0),.din(w_dff_A_aVeR2SgY8_0),.clk(gclk));
	jdff dff_A_qN2rgI7h4_0(.dout(w_dff_A_d2Leqkyp2_0),.din(w_dff_A_qN2rgI7h4_0),.clk(gclk));
	jdff dff_A_d2Leqkyp2_0(.dout(w_dff_A_bGGfmgPl6_0),.din(w_dff_A_d2Leqkyp2_0),.clk(gclk));
	jdff dff_A_bGGfmgPl6_0(.dout(w_dff_A_go56ikbc7_0),.din(w_dff_A_bGGfmgPl6_0),.clk(gclk));
	jdff dff_A_go56ikbc7_0(.dout(w_dff_A_f3CHvaWl7_0),.din(w_dff_A_go56ikbc7_0),.clk(gclk));
	jdff dff_A_f3CHvaWl7_0(.dout(w_dff_A_jqQC6r8m8_0),.din(w_dff_A_f3CHvaWl7_0),.clk(gclk));
	jdff dff_A_jqQC6r8m8_0(.dout(w_dff_A_aBGzrkyQ3_0),.din(w_dff_A_jqQC6r8m8_0),.clk(gclk));
	jdff dff_A_aBGzrkyQ3_0(.dout(w_dff_A_Za1zlMD60_0),.din(w_dff_A_aBGzrkyQ3_0),.clk(gclk));
	jdff dff_A_Za1zlMD60_0(.dout(w_dff_A_qzfSJFPC9_0),.din(w_dff_A_Za1zlMD60_0),.clk(gclk));
	jdff dff_A_qzfSJFPC9_0(.dout(w_dff_A_rT8MbJeM2_0),.din(w_dff_A_qzfSJFPC9_0),.clk(gclk));
	jdff dff_A_rT8MbJeM2_0(.dout(w_dff_A_gJXzCv1j1_0),.din(w_dff_A_rT8MbJeM2_0),.clk(gclk));
	jdff dff_A_gJXzCv1j1_0(.dout(w_dff_A_Vi5XxNHS2_0),.din(w_dff_A_gJXzCv1j1_0),.clk(gclk));
	jdff dff_A_Vi5XxNHS2_0(.dout(w_dff_A_L53p63RB4_0),.din(w_dff_A_Vi5XxNHS2_0),.clk(gclk));
	jdff dff_A_L53p63RB4_0(.dout(G552),.din(w_dff_A_L53p63RB4_0),.clk(gclk));
	jdff dff_A_OfvxdAZI9_1(.dout(w_dff_A_u6w11RdQ8_0),.din(w_dff_A_OfvxdAZI9_1),.clk(gclk));
	jdff dff_A_u6w11RdQ8_0(.dout(w_dff_A_gVfvJfFu9_0),.din(w_dff_A_u6w11RdQ8_0),.clk(gclk));
	jdff dff_A_gVfvJfFu9_0(.dout(w_dff_A_6qP8pnkO8_0),.din(w_dff_A_gVfvJfFu9_0),.clk(gclk));
	jdff dff_A_6qP8pnkO8_0(.dout(w_dff_A_0evuJGdV0_0),.din(w_dff_A_6qP8pnkO8_0),.clk(gclk));
	jdff dff_A_0evuJGdV0_0(.dout(w_dff_A_gQNLP9a55_0),.din(w_dff_A_0evuJGdV0_0),.clk(gclk));
	jdff dff_A_gQNLP9a55_0(.dout(w_dff_A_WguEMg0S5_0),.din(w_dff_A_gQNLP9a55_0),.clk(gclk));
	jdff dff_A_WguEMg0S5_0(.dout(w_dff_A_3kZrnrwH9_0),.din(w_dff_A_WguEMg0S5_0),.clk(gclk));
	jdff dff_A_3kZrnrwH9_0(.dout(w_dff_A_72MKYkRT3_0),.din(w_dff_A_3kZrnrwH9_0),.clk(gclk));
	jdff dff_A_72MKYkRT3_0(.dout(w_dff_A_oQxkLytR8_0),.din(w_dff_A_72MKYkRT3_0),.clk(gclk));
	jdff dff_A_oQxkLytR8_0(.dout(w_dff_A_OnQOin4c2_0),.din(w_dff_A_oQxkLytR8_0),.clk(gclk));
	jdff dff_A_OnQOin4c2_0(.dout(w_dff_A_mAzHswCT5_0),.din(w_dff_A_OnQOin4c2_0),.clk(gclk));
	jdff dff_A_mAzHswCT5_0(.dout(w_dff_A_O64vvKgi2_0),.din(w_dff_A_mAzHswCT5_0),.clk(gclk));
	jdff dff_A_O64vvKgi2_0(.dout(w_dff_A_r6ffcCki1_0),.din(w_dff_A_O64vvKgi2_0),.clk(gclk));
	jdff dff_A_r6ffcCki1_0(.dout(w_dff_A_UMKyvzuM8_0),.din(w_dff_A_r6ffcCki1_0),.clk(gclk));
	jdff dff_A_UMKyvzuM8_0(.dout(w_dff_A_AyJ4YQeu2_0),.din(w_dff_A_UMKyvzuM8_0),.clk(gclk));
	jdff dff_A_AyJ4YQeu2_0(.dout(w_dff_A_0RHyS6RY9_0),.din(w_dff_A_AyJ4YQeu2_0),.clk(gclk));
	jdff dff_A_0RHyS6RY9_0(.dout(w_dff_A_lN8WtdiX8_0),.din(w_dff_A_0RHyS6RY9_0),.clk(gclk));
	jdff dff_A_lN8WtdiX8_0(.dout(w_dff_A_09I1zbWa9_0),.din(w_dff_A_lN8WtdiX8_0),.clk(gclk));
	jdff dff_A_09I1zbWa9_0(.dout(w_dff_A_zX5IKqPQ7_0),.din(w_dff_A_09I1zbWa9_0),.clk(gclk));
	jdff dff_A_zX5IKqPQ7_0(.dout(w_dff_A_lhmmAC7S3_0),.din(w_dff_A_zX5IKqPQ7_0),.clk(gclk));
	jdff dff_A_lhmmAC7S3_0(.dout(w_dff_A_4auHpJRm7_0),.din(w_dff_A_lhmmAC7S3_0),.clk(gclk));
	jdff dff_A_4auHpJRm7_0(.dout(w_dff_A_2i9WPWth9_0),.din(w_dff_A_4auHpJRm7_0),.clk(gclk));
	jdff dff_A_2i9WPWth9_0(.dout(w_dff_A_aPEbTLQu3_0),.din(w_dff_A_2i9WPWth9_0),.clk(gclk));
	jdff dff_A_aPEbTLQu3_0(.dout(w_dff_A_K4uzrSny2_0),.din(w_dff_A_aPEbTLQu3_0),.clk(gclk));
	jdff dff_A_K4uzrSny2_0(.dout(w_dff_A_Y16NZxXz7_0),.din(w_dff_A_K4uzrSny2_0),.clk(gclk));
	jdff dff_A_Y16NZxXz7_0(.dout(w_dff_A_Kz7a0dJK3_0),.din(w_dff_A_Y16NZxXz7_0),.clk(gclk));
	jdff dff_A_Kz7a0dJK3_0(.dout(w_dff_A_Qxtx3XIQ0_0),.din(w_dff_A_Kz7a0dJK3_0),.clk(gclk));
	jdff dff_A_Qxtx3XIQ0_0(.dout(w_dff_A_F6jp2qLA6_0),.din(w_dff_A_Qxtx3XIQ0_0),.clk(gclk));
	jdff dff_A_F6jp2qLA6_0(.dout(w_dff_A_h61LNy6v1_0),.din(w_dff_A_F6jp2qLA6_0),.clk(gclk));
	jdff dff_A_h61LNy6v1_0(.dout(w_dff_A_n7aRZqte7_0),.din(w_dff_A_h61LNy6v1_0),.clk(gclk));
	jdff dff_A_n7aRZqte7_0(.dout(w_dff_A_1wnQql9o7_0),.din(w_dff_A_n7aRZqte7_0),.clk(gclk));
	jdff dff_A_1wnQql9o7_0(.dout(w_dff_A_Geec7v7P3_0),.din(w_dff_A_1wnQql9o7_0),.clk(gclk));
	jdff dff_A_Geec7v7P3_0(.dout(w_dff_A_BSKXJ16d3_0),.din(w_dff_A_Geec7v7P3_0),.clk(gclk));
	jdff dff_A_BSKXJ16d3_0(.dout(w_dff_A_3nrr3Pyi6_0),.din(w_dff_A_BSKXJ16d3_0),.clk(gclk));
	jdff dff_A_3nrr3Pyi6_0(.dout(w_dff_A_c6DmA7c72_0),.din(w_dff_A_3nrr3Pyi6_0),.clk(gclk));
	jdff dff_A_c6DmA7c72_0(.dout(w_dff_A_seyxrpUW8_0),.din(w_dff_A_c6DmA7c72_0),.clk(gclk));
	jdff dff_A_seyxrpUW8_0(.dout(w_dff_A_KVv70fzu6_0),.din(w_dff_A_seyxrpUW8_0),.clk(gclk));
	jdff dff_A_KVv70fzu6_0(.dout(w_dff_A_cWBRYjaq1_0),.din(w_dff_A_KVv70fzu6_0),.clk(gclk));
	jdff dff_A_cWBRYjaq1_0(.dout(G550),.din(w_dff_A_cWBRYjaq1_0),.clk(gclk));
	jdff dff_A_raA4ZSOf6_1(.dout(w_dff_A_JsonzD2n9_0),.din(w_dff_A_raA4ZSOf6_1),.clk(gclk));
	jdff dff_A_JsonzD2n9_0(.dout(w_dff_A_1FEFb6k40_0),.din(w_dff_A_JsonzD2n9_0),.clk(gclk));
	jdff dff_A_1FEFb6k40_0(.dout(w_dff_A_27xWi6MH1_0),.din(w_dff_A_1FEFb6k40_0),.clk(gclk));
	jdff dff_A_27xWi6MH1_0(.dout(w_dff_A_RRigINkF0_0),.din(w_dff_A_27xWi6MH1_0),.clk(gclk));
	jdff dff_A_RRigINkF0_0(.dout(w_dff_A_dNvhmzVZ6_0),.din(w_dff_A_RRigINkF0_0),.clk(gclk));
	jdff dff_A_dNvhmzVZ6_0(.dout(w_dff_A_YifYED4m2_0),.din(w_dff_A_dNvhmzVZ6_0),.clk(gclk));
	jdff dff_A_YifYED4m2_0(.dout(w_dff_A_YwG0u98N9_0),.din(w_dff_A_YifYED4m2_0),.clk(gclk));
	jdff dff_A_YwG0u98N9_0(.dout(w_dff_A_agu1s1IU2_0),.din(w_dff_A_YwG0u98N9_0),.clk(gclk));
	jdff dff_A_agu1s1IU2_0(.dout(w_dff_A_H8w1aGhe8_0),.din(w_dff_A_agu1s1IU2_0),.clk(gclk));
	jdff dff_A_H8w1aGhe8_0(.dout(w_dff_A_b20fpsaN7_0),.din(w_dff_A_H8w1aGhe8_0),.clk(gclk));
	jdff dff_A_b20fpsaN7_0(.dout(w_dff_A_6o3FVUH64_0),.din(w_dff_A_b20fpsaN7_0),.clk(gclk));
	jdff dff_A_6o3FVUH64_0(.dout(w_dff_A_6YCWbd2H3_0),.din(w_dff_A_6o3FVUH64_0),.clk(gclk));
	jdff dff_A_6YCWbd2H3_0(.dout(w_dff_A_JXZK6Gig5_0),.din(w_dff_A_6YCWbd2H3_0),.clk(gclk));
	jdff dff_A_JXZK6Gig5_0(.dout(w_dff_A_u4giKg3J1_0),.din(w_dff_A_JXZK6Gig5_0),.clk(gclk));
	jdff dff_A_u4giKg3J1_0(.dout(w_dff_A_tnzplJ4T0_0),.din(w_dff_A_u4giKg3J1_0),.clk(gclk));
	jdff dff_A_tnzplJ4T0_0(.dout(w_dff_A_CIdePGpv1_0),.din(w_dff_A_tnzplJ4T0_0),.clk(gclk));
	jdff dff_A_CIdePGpv1_0(.dout(w_dff_A_xYfrSgnN8_0),.din(w_dff_A_CIdePGpv1_0),.clk(gclk));
	jdff dff_A_xYfrSgnN8_0(.dout(w_dff_A_8c83QNxC2_0),.din(w_dff_A_xYfrSgnN8_0),.clk(gclk));
	jdff dff_A_8c83QNxC2_0(.dout(w_dff_A_JTDxKvRv8_0),.din(w_dff_A_8c83QNxC2_0),.clk(gclk));
	jdff dff_A_JTDxKvRv8_0(.dout(w_dff_A_UnKXg5GR2_0),.din(w_dff_A_JTDxKvRv8_0),.clk(gclk));
	jdff dff_A_UnKXg5GR2_0(.dout(w_dff_A_aZvQrLwx4_0),.din(w_dff_A_UnKXg5GR2_0),.clk(gclk));
	jdff dff_A_aZvQrLwx4_0(.dout(w_dff_A_3LWuqz2S5_0),.din(w_dff_A_aZvQrLwx4_0),.clk(gclk));
	jdff dff_A_3LWuqz2S5_0(.dout(w_dff_A_5NwHhuGE2_0),.din(w_dff_A_3LWuqz2S5_0),.clk(gclk));
	jdff dff_A_5NwHhuGE2_0(.dout(w_dff_A_NKpto9AQ6_0),.din(w_dff_A_5NwHhuGE2_0),.clk(gclk));
	jdff dff_A_NKpto9AQ6_0(.dout(w_dff_A_PhVbRa9F6_0),.din(w_dff_A_NKpto9AQ6_0),.clk(gclk));
	jdff dff_A_PhVbRa9F6_0(.dout(w_dff_A_vJ3Libtc0_0),.din(w_dff_A_PhVbRa9F6_0),.clk(gclk));
	jdff dff_A_vJ3Libtc0_0(.dout(w_dff_A_jJSL0Y978_0),.din(w_dff_A_vJ3Libtc0_0),.clk(gclk));
	jdff dff_A_jJSL0Y978_0(.dout(w_dff_A_fPdXwmPX5_0),.din(w_dff_A_jJSL0Y978_0),.clk(gclk));
	jdff dff_A_fPdXwmPX5_0(.dout(w_dff_A_rQPHKf2f9_0),.din(w_dff_A_fPdXwmPX5_0),.clk(gclk));
	jdff dff_A_rQPHKf2f9_0(.dout(w_dff_A_2uHhfrbJ5_0),.din(w_dff_A_rQPHKf2f9_0),.clk(gclk));
	jdff dff_A_2uHhfrbJ5_0(.dout(w_dff_A_H7igYsBG8_0),.din(w_dff_A_2uHhfrbJ5_0),.clk(gclk));
	jdff dff_A_H7igYsBG8_0(.dout(w_dff_A_PCJQs6Ti8_0),.din(w_dff_A_H7igYsBG8_0),.clk(gclk));
	jdff dff_A_PCJQs6Ti8_0(.dout(w_dff_A_ZLxdT2nR1_0),.din(w_dff_A_PCJQs6Ti8_0),.clk(gclk));
	jdff dff_A_ZLxdT2nR1_0(.dout(w_dff_A_1WBCEbt64_0),.din(w_dff_A_ZLxdT2nR1_0),.clk(gclk));
	jdff dff_A_1WBCEbt64_0(.dout(w_dff_A_qEqrCszF4_0),.din(w_dff_A_1WBCEbt64_0),.clk(gclk));
	jdff dff_A_qEqrCszF4_0(.dout(w_dff_A_D1bRoyE32_0),.din(w_dff_A_qEqrCszF4_0),.clk(gclk));
	jdff dff_A_D1bRoyE32_0(.dout(w_dff_A_zl51YVJi4_0),.din(w_dff_A_D1bRoyE32_0),.clk(gclk));
	jdff dff_A_zl51YVJi4_0(.dout(w_dff_A_AYvTdkIM1_0),.din(w_dff_A_zl51YVJi4_0),.clk(gclk));
	jdff dff_A_AYvTdkIM1_0(.dout(G548),.din(w_dff_A_AYvTdkIM1_0),.clk(gclk));
	jdff dff_A_cdzx6Owo0_1(.dout(w_dff_A_Q2vYo6iT3_0),.din(w_dff_A_cdzx6Owo0_1),.clk(gclk));
	jdff dff_A_Q2vYo6iT3_0(.dout(w_dff_A_I2nAqOy29_0),.din(w_dff_A_Q2vYo6iT3_0),.clk(gclk));
	jdff dff_A_I2nAqOy29_0(.dout(w_dff_A_hEW80LHj8_0),.din(w_dff_A_I2nAqOy29_0),.clk(gclk));
	jdff dff_A_hEW80LHj8_0(.dout(w_dff_A_5AqO0yc54_0),.din(w_dff_A_hEW80LHj8_0),.clk(gclk));
	jdff dff_A_5AqO0yc54_0(.dout(w_dff_A_sFVRGxik1_0),.din(w_dff_A_5AqO0yc54_0),.clk(gclk));
	jdff dff_A_sFVRGxik1_0(.dout(w_dff_A_fBSuky5A1_0),.din(w_dff_A_sFVRGxik1_0),.clk(gclk));
	jdff dff_A_fBSuky5A1_0(.dout(w_dff_A_78wQVgxb4_0),.din(w_dff_A_fBSuky5A1_0),.clk(gclk));
	jdff dff_A_78wQVgxb4_0(.dout(w_dff_A_uRcIAe7U4_0),.din(w_dff_A_78wQVgxb4_0),.clk(gclk));
	jdff dff_A_uRcIAe7U4_0(.dout(w_dff_A_XopxEOvI9_0),.din(w_dff_A_uRcIAe7U4_0),.clk(gclk));
	jdff dff_A_XopxEOvI9_0(.dout(w_dff_A_DQ2lfse11_0),.din(w_dff_A_XopxEOvI9_0),.clk(gclk));
	jdff dff_A_DQ2lfse11_0(.dout(w_dff_A_rlQG7AFW3_0),.din(w_dff_A_DQ2lfse11_0),.clk(gclk));
	jdff dff_A_rlQG7AFW3_0(.dout(w_dff_A_FmaAT13e0_0),.din(w_dff_A_rlQG7AFW3_0),.clk(gclk));
	jdff dff_A_FmaAT13e0_0(.dout(w_dff_A_lYEkRAoq4_0),.din(w_dff_A_FmaAT13e0_0),.clk(gclk));
	jdff dff_A_lYEkRAoq4_0(.dout(w_dff_A_3K9slGGc9_0),.din(w_dff_A_lYEkRAoq4_0),.clk(gclk));
	jdff dff_A_3K9slGGc9_0(.dout(w_dff_A_8Lc4IL521_0),.din(w_dff_A_3K9slGGc9_0),.clk(gclk));
	jdff dff_A_8Lc4IL521_0(.dout(w_dff_A_10MirRNo9_0),.din(w_dff_A_8Lc4IL521_0),.clk(gclk));
	jdff dff_A_10MirRNo9_0(.dout(w_dff_A_4ZLUGN9Y2_0),.din(w_dff_A_10MirRNo9_0),.clk(gclk));
	jdff dff_A_4ZLUGN9Y2_0(.dout(w_dff_A_CIYjPe135_0),.din(w_dff_A_4ZLUGN9Y2_0),.clk(gclk));
	jdff dff_A_CIYjPe135_0(.dout(w_dff_A_lRt2hjzH2_0),.din(w_dff_A_CIYjPe135_0),.clk(gclk));
	jdff dff_A_lRt2hjzH2_0(.dout(w_dff_A_HYYqvbGz5_0),.din(w_dff_A_lRt2hjzH2_0),.clk(gclk));
	jdff dff_A_HYYqvbGz5_0(.dout(w_dff_A_fNzDb7rS7_0),.din(w_dff_A_HYYqvbGz5_0),.clk(gclk));
	jdff dff_A_fNzDb7rS7_0(.dout(w_dff_A_h4oIc3Mn2_0),.din(w_dff_A_fNzDb7rS7_0),.clk(gclk));
	jdff dff_A_h4oIc3Mn2_0(.dout(w_dff_A_tX8PkE9y2_0),.din(w_dff_A_h4oIc3Mn2_0),.clk(gclk));
	jdff dff_A_tX8PkE9y2_0(.dout(w_dff_A_BOgF5B9s8_0),.din(w_dff_A_tX8PkE9y2_0),.clk(gclk));
	jdff dff_A_BOgF5B9s8_0(.dout(w_dff_A_uV0C22BX2_0),.din(w_dff_A_BOgF5B9s8_0),.clk(gclk));
	jdff dff_A_uV0C22BX2_0(.dout(w_dff_A_GZxWhTm66_0),.din(w_dff_A_uV0C22BX2_0),.clk(gclk));
	jdff dff_A_GZxWhTm66_0(.dout(w_dff_A_azJgPFh68_0),.din(w_dff_A_GZxWhTm66_0),.clk(gclk));
	jdff dff_A_azJgPFh68_0(.dout(w_dff_A_Gf4MZAsF8_0),.din(w_dff_A_azJgPFh68_0),.clk(gclk));
	jdff dff_A_Gf4MZAsF8_0(.dout(w_dff_A_AfH548px0_0),.din(w_dff_A_Gf4MZAsF8_0),.clk(gclk));
	jdff dff_A_AfH548px0_0(.dout(w_dff_A_12qmTvYC5_0),.din(w_dff_A_AfH548px0_0),.clk(gclk));
	jdff dff_A_12qmTvYC5_0(.dout(w_dff_A_zOE9RhDo4_0),.din(w_dff_A_12qmTvYC5_0),.clk(gclk));
	jdff dff_A_zOE9RhDo4_0(.dout(w_dff_A_nT8oR8Zy9_0),.din(w_dff_A_zOE9RhDo4_0),.clk(gclk));
	jdff dff_A_nT8oR8Zy9_0(.dout(w_dff_A_wdPlmwse4_0),.din(w_dff_A_nT8oR8Zy9_0),.clk(gclk));
	jdff dff_A_wdPlmwse4_0(.dout(w_dff_A_0iLuSKBQ0_0),.din(w_dff_A_wdPlmwse4_0),.clk(gclk));
	jdff dff_A_0iLuSKBQ0_0(.dout(w_dff_A_c4LIxd3n2_0),.din(w_dff_A_0iLuSKBQ0_0),.clk(gclk));
	jdff dff_A_c4LIxd3n2_0(.dout(w_dff_A_QgJWroce0_0),.din(w_dff_A_c4LIxd3n2_0),.clk(gclk));
	jdff dff_A_QgJWroce0_0(.dout(w_dff_A_nbgJAfPH5_0),.din(w_dff_A_QgJWroce0_0),.clk(gclk));
	jdff dff_A_nbgJAfPH5_0(.dout(w_dff_A_RHmuEuxu0_0),.din(w_dff_A_nbgJAfPH5_0),.clk(gclk));
	jdff dff_A_RHmuEuxu0_0(.dout(G546),.din(w_dff_A_RHmuEuxu0_0),.clk(gclk));
	jdff dff_A_34A5K7yA7_1(.dout(w_dff_A_YYy4sqko7_0),.din(w_dff_A_34A5K7yA7_1),.clk(gclk));
	jdff dff_A_YYy4sqko7_0(.dout(w_dff_A_O6WxUSNV2_0),.din(w_dff_A_YYy4sqko7_0),.clk(gclk));
	jdff dff_A_O6WxUSNV2_0(.dout(w_dff_A_Hww3Vx2F3_0),.din(w_dff_A_O6WxUSNV2_0),.clk(gclk));
	jdff dff_A_Hww3Vx2F3_0(.dout(w_dff_A_nZ8o2BWI4_0),.din(w_dff_A_Hww3Vx2F3_0),.clk(gclk));
	jdff dff_A_nZ8o2BWI4_0(.dout(w_dff_A_wn9mJYof6_0),.din(w_dff_A_nZ8o2BWI4_0),.clk(gclk));
	jdff dff_A_wn9mJYof6_0(.dout(w_dff_A_pjOWfvd54_0),.din(w_dff_A_wn9mJYof6_0),.clk(gclk));
	jdff dff_A_pjOWfvd54_0(.dout(w_dff_A_Kr9kCJOH5_0),.din(w_dff_A_pjOWfvd54_0),.clk(gclk));
	jdff dff_A_Kr9kCJOH5_0(.dout(w_dff_A_wg2BCycD8_0),.din(w_dff_A_Kr9kCJOH5_0),.clk(gclk));
	jdff dff_A_wg2BCycD8_0(.dout(w_dff_A_MYe3cHNE2_0),.din(w_dff_A_wg2BCycD8_0),.clk(gclk));
	jdff dff_A_MYe3cHNE2_0(.dout(w_dff_A_w9IBA8XL6_0),.din(w_dff_A_MYe3cHNE2_0),.clk(gclk));
	jdff dff_A_w9IBA8XL6_0(.dout(w_dff_A_2nDwcplW4_0),.din(w_dff_A_w9IBA8XL6_0),.clk(gclk));
	jdff dff_A_2nDwcplW4_0(.dout(w_dff_A_h535TGIq5_0),.din(w_dff_A_2nDwcplW4_0),.clk(gclk));
	jdff dff_A_h535TGIq5_0(.dout(w_dff_A_rOou0g5I4_0),.din(w_dff_A_h535TGIq5_0),.clk(gclk));
	jdff dff_A_rOou0g5I4_0(.dout(w_dff_A_cgo5ybVO1_0),.din(w_dff_A_rOou0g5I4_0),.clk(gclk));
	jdff dff_A_cgo5ybVO1_0(.dout(w_dff_A_AI6EbtoA9_0),.din(w_dff_A_cgo5ybVO1_0),.clk(gclk));
	jdff dff_A_AI6EbtoA9_0(.dout(w_dff_A_YDJNwgpP5_0),.din(w_dff_A_AI6EbtoA9_0),.clk(gclk));
	jdff dff_A_YDJNwgpP5_0(.dout(w_dff_A_QPrX51YL7_0),.din(w_dff_A_YDJNwgpP5_0),.clk(gclk));
	jdff dff_A_QPrX51YL7_0(.dout(w_dff_A_Es8ZUgLv8_0),.din(w_dff_A_QPrX51YL7_0),.clk(gclk));
	jdff dff_A_Es8ZUgLv8_0(.dout(w_dff_A_0GRQwzjl4_0),.din(w_dff_A_Es8ZUgLv8_0),.clk(gclk));
	jdff dff_A_0GRQwzjl4_0(.dout(w_dff_A_mLHrelrP7_0),.din(w_dff_A_0GRQwzjl4_0),.clk(gclk));
	jdff dff_A_mLHrelrP7_0(.dout(w_dff_A_8cuvPt7V1_0),.din(w_dff_A_mLHrelrP7_0),.clk(gclk));
	jdff dff_A_8cuvPt7V1_0(.dout(w_dff_A_NwBWVVcX1_0),.din(w_dff_A_8cuvPt7V1_0),.clk(gclk));
	jdff dff_A_NwBWVVcX1_0(.dout(w_dff_A_Dx9qxdNX2_0),.din(w_dff_A_NwBWVVcX1_0),.clk(gclk));
	jdff dff_A_Dx9qxdNX2_0(.dout(w_dff_A_F4ma6W6j2_0),.din(w_dff_A_Dx9qxdNX2_0),.clk(gclk));
	jdff dff_A_F4ma6W6j2_0(.dout(w_dff_A_rEMHaQ3A4_0),.din(w_dff_A_F4ma6W6j2_0),.clk(gclk));
	jdff dff_A_rEMHaQ3A4_0(.dout(w_dff_A_6Fu8ZWVr2_0),.din(w_dff_A_rEMHaQ3A4_0),.clk(gclk));
	jdff dff_A_6Fu8ZWVr2_0(.dout(w_dff_A_NAg3yQwV2_0),.din(w_dff_A_6Fu8ZWVr2_0),.clk(gclk));
	jdff dff_A_NAg3yQwV2_0(.dout(w_dff_A_bWPxweDt0_0),.din(w_dff_A_NAg3yQwV2_0),.clk(gclk));
	jdff dff_A_bWPxweDt0_0(.dout(w_dff_A_FZEVdlcS9_0),.din(w_dff_A_bWPxweDt0_0),.clk(gclk));
	jdff dff_A_FZEVdlcS9_0(.dout(w_dff_A_JxgndWWk8_0),.din(w_dff_A_FZEVdlcS9_0),.clk(gclk));
	jdff dff_A_JxgndWWk8_0(.dout(w_dff_A_0cIJTg6E1_0),.din(w_dff_A_JxgndWWk8_0),.clk(gclk));
	jdff dff_A_0cIJTg6E1_0(.dout(w_dff_A_2DR5c3VK1_0),.din(w_dff_A_0cIJTg6E1_0),.clk(gclk));
	jdff dff_A_2DR5c3VK1_0(.dout(w_dff_A_YJoPn7qq5_0),.din(w_dff_A_2DR5c3VK1_0),.clk(gclk));
	jdff dff_A_YJoPn7qq5_0(.dout(w_dff_A_Ixrh25oI7_0),.din(w_dff_A_YJoPn7qq5_0),.clk(gclk));
	jdff dff_A_Ixrh25oI7_0(.dout(w_dff_A_XvcRrPbp4_0),.din(w_dff_A_Ixrh25oI7_0),.clk(gclk));
	jdff dff_A_XvcRrPbp4_0(.dout(w_dff_A_2AAweAFa4_0),.din(w_dff_A_XvcRrPbp4_0),.clk(gclk));
	jdff dff_A_2AAweAFa4_0(.dout(w_dff_A_KKwDUADl4_0),.din(w_dff_A_2AAweAFa4_0),.clk(gclk));
	jdff dff_A_KKwDUADl4_0(.dout(w_dff_A_tCT5eKfd3_0),.din(w_dff_A_KKwDUADl4_0),.clk(gclk));
	jdff dff_A_tCT5eKfd3_0(.dout(G544),.din(w_dff_A_tCT5eKfd3_0),.clk(gclk));
	jdff dff_A_kb3quiGP8_1(.dout(w_dff_A_sws1mcak6_0),.din(w_dff_A_kb3quiGP8_1),.clk(gclk));
	jdff dff_A_sws1mcak6_0(.dout(w_dff_A_eHVzY1QB8_0),.din(w_dff_A_sws1mcak6_0),.clk(gclk));
	jdff dff_A_eHVzY1QB8_0(.dout(w_dff_A_7T5N5bgl5_0),.din(w_dff_A_eHVzY1QB8_0),.clk(gclk));
	jdff dff_A_7T5N5bgl5_0(.dout(w_dff_A_YN3Svbd34_0),.din(w_dff_A_7T5N5bgl5_0),.clk(gclk));
	jdff dff_A_YN3Svbd34_0(.dout(w_dff_A_tWWm99yc8_0),.din(w_dff_A_YN3Svbd34_0),.clk(gclk));
	jdff dff_A_tWWm99yc8_0(.dout(w_dff_A_t2wWbrph2_0),.din(w_dff_A_tWWm99yc8_0),.clk(gclk));
	jdff dff_A_t2wWbrph2_0(.dout(w_dff_A_4Z18cAcd1_0),.din(w_dff_A_t2wWbrph2_0),.clk(gclk));
	jdff dff_A_4Z18cAcd1_0(.dout(w_dff_A_YRGoSWNz9_0),.din(w_dff_A_4Z18cAcd1_0),.clk(gclk));
	jdff dff_A_YRGoSWNz9_0(.dout(w_dff_A_jGCQWyix8_0),.din(w_dff_A_YRGoSWNz9_0),.clk(gclk));
	jdff dff_A_jGCQWyix8_0(.dout(w_dff_A_jgC289Hi2_0),.din(w_dff_A_jGCQWyix8_0),.clk(gclk));
	jdff dff_A_jgC289Hi2_0(.dout(w_dff_A_dno8tfrB2_0),.din(w_dff_A_jgC289Hi2_0),.clk(gclk));
	jdff dff_A_dno8tfrB2_0(.dout(w_dff_A_4i6coCeV3_0),.din(w_dff_A_dno8tfrB2_0),.clk(gclk));
	jdff dff_A_4i6coCeV3_0(.dout(w_dff_A_jzC4GcB65_0),.din(w_dff_A_4i6coCeV3_0),.clk(gclk));
	jdff dff_A_jzC4GcB65_0(.dout(w_dff_A_XACZ4ObN1_0),.din(w_dff_A_jzC4GcB65_0),.clk(gclk));
	jdff dff_A_XACZ4ObN1_0(.dout(w_dff_A_8unOYwrm5_0),.din(w_dff_A_XACZ4ObN1_0),.clk(gclk));
	jdff dff_A_8unOYwrm5_0(.dout(w_dff_A_JZ8Zvg5O6_0),.din(w_dff_A_8unOYwrm5_0),.clk(gclk));
	jdff dff_A_JZ8Zvg5O6_0(.dout(w_dff_A_qZ7Ldncm9_0),.din(w_dff_A_JZ8Zvg5O6_0),.clk(gclk));
	jdff dff_A_qZ7Ldncm9_0(.dout(w_dff_A_LbQ70CBp4_0),.din(w_dff_A_qZ7Ldncm9_0),.clk(gclk));
	jdff dff_A_LbQ70CBp4_0(.dout(w_dff_A_815YWJ2x8_0),.din(w_dff_A_LbQ70CBp4_0),.clk(gclk));
	jdff dff_A_815YWJ2x8_0(.dout(w_dff_A_vH264ND87_0),.din(w_dff_A_815YWJ2x8_0),.clk(gclk));
	jdff dff_A_vH264ND87_0(.dout(w_dff_A_flJHiBxc1_0),.din(w_dff_A_vH264ND87_0),.clk(gclk));
	jdff dff_A_flJHiBxc1_0(.dout(w_dff_A_G0wH6e5i3_0),.din(w_dff_A_flJHiBxc1_0),.clk(gclk));
	jdff dff_A_G0wH6e5i3_0(.dout(w_dff_A_DltdmxHx7_0),.din(w_dff_A_G0wH6e5i3_0),.clk(gclk));
	jdff dff_A_DltdmxHx7_0(.dout(w_dff_A_ByPB2ARu6_0),.din(w_dff_A_DltdmxHx7_0),.clk(gclk));
	jdff dff_A_ByPB2ARu6_0(.dout(w_dff_A_Olq6KVgr2_0),.din(w_dff_A_ByPB2ARu6_0),.clk(gclk));
	jdff dff_A_Olq6KVgr2_0(.dout(w_dff_A_vs1JXJ5y8_0),.din(w_dff_A_Olq6KVgr2_0),.clk(gclk));
	jdff dff_A_vs1JXJ5y8_0(.dout(w_dff_A_Xfkpeue67_0),.din(w_dff_A_vs1JXJ5y8_0),.clk(gclk));
	jdff dff_A_Xfkpeue67_0(.dout(w_dff_A_aR3Sna410_0),.din(w_dff_A_Xfkpeue67_0),.clk(gclk));
	jdff dff_A_aR3Sna410_0(.dout(w_dff_A_6VorzEux4_0),.din(w_dff_A_aR3Sna410_0),.clk(gclk));
	jdff dff_A_6VorzEux4_0(.dout(w_dff_A_ELM2bTzb3_0),.din(w_dff_A_6VorzEux4_0),.clk(gclk));
	jdff dff_A_ELM2bTzb3_0(.dout(w_dff_A_YJuaxuA56_0),.din(w_dff_A_ELM2bTzb3_0),.clk(gclk));
	jdff dff_A_YJuaxuA56_0(.dout(w_dff_A_7PtTTNbd7_0),.din(w_dff_A_YJuaxuA56_0),.clk(gclk));
	jdff dff_A_7PtTTNbd7_0(.dout(w_dff_A_blD2RiJn5_0),.din(w_dff_A_7PtTTNbd7_0),.clk(gclk));
	jdff dff_A_blD2RiJn5_0(.dout(w_dff_A_nVDlxkkq5_0),.din(w_dff_A_blD2RiJn5_0),.clk(gclk));
	jdff dff_A_nVDlxkkq5_0(.dout(w_dff_A_yGDEcFTE9_0),.din(w_dff_A_nVDlxkkq5_0),.clk(gclk));
	jdff dff_A_yGDEcFTE9_0(.dout(w_dff_A_lx6OzEzQ5_0),.din(w_dff_A_yGDEcFTE9_0),.clk(gclk));
	jdff dff_A_lx6OzEzQ5_0(.dout(w_dff_A_mbyBwvos9_0),.din(w_dff_A_lx6OzEzQ5_0),.clk(gclk));
	jdff dff_A_mbyBwvos9_0(.dout(w_dff_A_Vj1kNBeA7_0),.din(w_dff_A_mbyBwvos9_0),.clk(gclk));
	jdff dff_A_Vj1kNBeA7_0(.dout(G540),.din(w_dff_A_Vj1kNBeA7_0),.clk(gclk));
	jdff dff_A_5GiWzOQF0_1(.dout(w_dff_A_aEpl5dPU0_0),.din(w_dff_A_5GiWzOQF0_1),.clk(gclk));
	jdff dff_A_aEpl5dPU0_0(.dout(w_dff_A_5oSoT8jO1_0),.din(w_dff_A_aEpl5dPU0_0),.clk(gclk));
	jdff dff_A_5oSoT8jO1_0(.dout(w_dff_A_rwVjqHsJ6_0),.din(w_dff_A_5oSoT8jO1_0),.clk(gclk));
	jdff dff_A_rwVjqHsJ6_0(.dout(w_dff_A_dp23amMn5_0),.din(w_dff_A_rwVjqHsJ6_0),.clk(gclk));
	jdff dff_A_dp23amMn5_0(.dout(w_dff_A_WJcD30dT3_0),.din(w_dff_A_dp23amMn5_0),.clk(gclk));
	jdff dff_A_WJcD30dT3_0(.dout(w_dff_A_scoYqcGf7_0),.din(w_dff_A_WJcD30dT3_0),.clk(gclk));
	jdff dff_A_scoYqcGf7_0(.dout(w_dff_A_jBFjaZrK3_0),.din(w_dff_A_scoYqcGf7_0),.clk(gclk));
	jdff dff_A_jBFjaZrK3_0(.dout(w_dff_A_hZNQNLVY3_0),.din(w_dff_A_jBFjaZrK3_0),.clk(gclk));
	jdff dff_A_hZNQNLVY3_0(.dout(w_dff_A_1ahuj7sp4_0),.din(w_dff_A_hZNQNLVY3_0),.clk(gclk));
	jdff dff_A_1ahuj7sp4_0(.dout(w_dff_A_eC30xmAe9_0),.din(w_dff_A_1ahuj7sp4_0),.clk(gclk));
	jdff dff_A_eC30xmAe9_0(.dout(w_dff_A_aEG3ns3P3_0),.din(w_dff_A_eC30xmAe9_0),.clk(gclk));
	jdff dff_A_aEG3ns3P3_0(.dout(w_dff_A_EWZHG3wT8_0),.din(w_dff_A_aEG3ns3P3_0),.clk(gclk));
	jdff dff_A_EWZHG3wT8_0(.dout(w_dff_A_WXYRMgKc2_0),.din(w_dff_A_EWZHG3wT8_0),.clk(gclk));
	jdff dff_A_WXYRMgKc2_0(.dout(w_dff_A_WqG2lU4F2_0),.din(w_dff_A_WXYRMgKc2_0),.clk(gclk));
	jdff dff_A_WqG2lU4F2_0(.dout(w_dff_A_n2XbPuEm2_0),.din(w_dff_A_WqG2lU4F2_0),.clk(gclk));
	jdff dff_A_n2XbPuEm2_0(.dout(w_dff_A_dodAIOqs3_0),.din(w_dff_A_n2XbPuEm2_0),.clk(gclk));
	jdff dff_A_dodAIOqs3_0(.dout(w_dff_A_5eikFxYu7_0),.din(w_dff_A_dodAIOqs3_0),.clk(gclk));
	jdff dff_A_5eikFxYu7_0(.dout(w_dff_A_aFKANECi0_0),.din(w_dff_A_5eikFxYu7_0),.clk(gclk));
	jdff dff_A_aFKANECi0_0(.dout(w_dff_A_MeBg5q7G5_0),.din(w_dff_A_aFKANECi0_0),.clk(gclk));
	jdff dff_A_MeBg5q7G5_0(.dout(w_dff_A_sMTyoztj8_0),.din(w_dff_A_MeBg5q7G5_0),.clk(gclk));
	jdff dff_A_sMTyoztj8_0(.dout(w_dff_A_MZSXbWH45_0),.din(w_dff_A_sMTyoztj8_0),.clk(gclk));
	jdff dff_A_MZSXbWH45_0(.dout(w_dff_A_749LB0Xs8_0),.din(w_dff_A_MZSXbWH45_0),.clk(gclk));
	jdff dff_A_749LB0Xs8_0(.dout(w_dff_A_pudogwcz5_0),.din(w_dff_A_749LB0Xs8_0),.clk(gclk));
	jdff dff_A_pudogwcz5_0(.dout(w_dff_A_Tj3pnvvU6_0),.din(w_dff_A_pudogwcz5_0),.clk(gclk));
	jdff dff_A_Tj3pnvvU6_0(.dout(w_dff_A_Aioi3WAO4_0),.din(w_dff_A_Tj3pnvvU6_0),.clk(gclk));
	jdff dff_A_Aioi3WAO4_0(.dout(w_dff_A_00lnqNId7_0),.din(w_dff_A_Aioi3WAO4_0),.clk(gclk));
	jdff dff_A_00lnqNId7_0(.dout(w_dff_A_yNqaZA5K5_0),.din(w_dff_A_00lnqNId7_0),.clk(gclk));
	jdff dff_A_yNqaZA5K5_0(.dout(w_dff_A_Jt4d8DcT6_0),.din(w_dff_A_yNqaZA5K5_0),.clk(gclk));
	jdff dff_A_Jt4d8DcT6_0(.dout(w_dff_A_Ag6yEwyO8_0),.din(w_dff_A_Jt4d8DcT6_0),.clk(gclk));
	jdff dff_A_Ag6yEwyO8_0(.dout(w_dff_A_GgSRjkx82_0),.din(w_dff_A_Ag6yEwyO8_0),.clk(gclk));
	jdff dff_A_GgSRjkx82_0(.dout(w_dff_A_ghQsRmtn1_0),.din(w_dff_A_GgSRjkx82_0),.clk(gclk));
	jdff dff_A_ghQsRmtn1_0(.dout(w_dff_A_SvIOz8Nl1_0),.din(w_dff_A_ghQsRmtn1_0),.clk(gclk));
	jdff dff_A_SvIOz8Nl1_0(.dout(w_dff_A_ZItLgTyd3_0),.din(w_dff_A_SvIOz8Nl1_0),.clk(gclk));
	jdff dff_A_ZItLgTyd3_0(.dout(w_dff_A_8rHoO3FM4_0),.din(w_dff_A_ZItLgTyd3_0),.clk(gclk));
	jdff dff_A_8rHoO3FM4_0(.dout(w_dff_A_kld8f9Z77_0),.din(w_dff_A_8rHoO3FM4_0),.clk(gclk));
	jdff dff_A_kld8f9Z77_0(.dout(w_dff_A_Kj5KJFDM7_0),.din(w_dff_A_kld8f9Z77_0),.clk(gclk));
	jdff dff_A_Kj5KJFDM7_0(.dout(w_dff_A_2KX31jHY6_0),.din(w_dff_A_Kj5KJFDM7_0),.clk(gclk));
	jdff dff_A_2KX31jHY6_0(.dout(w_dff_A_0nfS8F1I7_0),.din(w_dff_A_2KX31jHY6_0),.clk(gclk));
	jdff dff_A_0nfS8F1I7_0(.dout(G538),.din(w_dff_A_0nfS8F1I7_0),.clk(gclk));
	jdff dff_A_vkEKZ9tY8_1(.dout(w_dff_A_3Hga92oZ0_0),.din(w_dff_A_vkEKZ9tY8_1),.clk(gclk));
	jdff dff_A_3Hga92oZ0_0(.dout(w_dff_A_khtVPgM78_0),.din(w_dff_A_3Hga92oZ0_0),.clk(gclk));
	jdff dff_A_khtVPgM78_0(.dout(w_dff_A_11Wyybou4_0),.din(w_dff_A_khtVPgM78_0),.clk(gclk));
	jdff dff_A_11Wyybou4_0(.dout(w_dff_A_WoMGRrGq8_0),.din(w_dff_A_11Wyybou4_0),.clk(gclk));
	jdff dff_A_WoMGRrGq8_0(.dout(w_dff_A_M3jD6m6m0_0),.din(w_dff_A_WoMGRrGq8_0),.clk(gclk));
	jdff dff_A_M3jD6m6m0_0(.dout(w_dff_A_dp2iTbNE4_0),.din(w_dff_A_M3jD6m6m0_0),.clk(gclk));
	jdff dff_A_dp2iTbNE4_0(.dout(w_dff_A_2zauRqPv3_0),.din(w_dff_A_dp2iTbNE4_0),.clk(gclk));
	jdff dff_A_2zauRqPv3_0(.dout(w_dff_A_Iv07XKB11_0),.din(w_dff_A_2zauRqPv3_0),.clk(gclk));
	jdff dff_A_Iv07XKB11_0(.dout(w_dff_A_AYcvrKBm4_0),.din(w_dff_A_Iv07XKB11_0),.clk(gclk));
	jdff dff_A_AYcvrKBm4_0(.dout(w_dff_A_USkBZdhj3_0),.din(w_dff_A_AYcvrKBm4_0),.clk(gclk));
	jdff dff_A_USkBZdhj3_0(.dout(w_dff_A_Hl6BNh9y6_0),.din(w_dff_A_USkBZdhj3_0),.clk(gclk));
	jdff dff_A_Hl6BNh9y6_0(.dout(w_dff_A_gq3eAXEG8_0),.din(w_dff_A_Hl6BNh9y6_0),.clk(gclk));
	jdff dff_A_gq3eAXEG8_0(.dout(w_dff_A_qNoK2uQk1_0),.din(w_dff_A_gq3eAXEG8_0),.clk(gclk));
	jdff dff_A_qNoK2uQk1_0(.dout(w_dff_A_1SmrEwel9_0),.din(w_dff_A_qNoK2uQk1_0),.clk(gclk));
	jdff dff_A_1SmrEwel9_0(.dout(w_dff_A_YydFjzVM7_0),.din(w_dff_A_1SmrEwel9_0),.clk(gclk));
	jdff dff_A_YydFjzVM7_0(.dout(w_dff_A_W2mIK5yg7_0),.din(w_dff_A_YydFjzVM7_0),.clk(gclk));
	jdff dff_A_W2mIK5yg7_0(.dout(w_dff_A_03IhAZp77_0),.din(w_dff_A_W2mIK5yg7_0),.clk(gclk));
	jdff dff_A_03IhAZp77_0(.dout(w_dff_A_aB6KPaFm9_0),.din(w_dff_A_03IhAZp77_0),.clk(gclk));
	jdff dff_A_aB6KPaFm9_0(.dout(w_dff_A_skQ4Dmx88_0),.din(w_dff_A_aB6KPaFm9_0),.clk(gclk));
	jdff dff_A_skQ4Dmx88_0(.dout(w_dff_A_YWqL8S1h1_0),.din(w_dff_A_skQ4Dmx88_0),.clk(gclk));
	jdff dff_A_YWqL8S1h1_0(.dout(w_dff_A_AKbjk9nv2_0),.din(w_dff_A_YWqL8S1h1_0),.clk(gclk));
	jdff dff_A_AKbjk9nv2_0(.dout(w_dff_A_F8RXZ21P3_0),.din(w_dff_A_AKbjk9nv2_0),.clk(gclk));
	jdff dff_A_F8RXZ21P3_0(.dout(w_dff_A_T8jB2xNd3_0),.din(w_dff_A_F8RXZ21P3_0),.clk(gclk));
	jdff dff_A_T8jB2xNd3_0(.dout(w_dff_A_dJsbkDX95_0),.din(w_dff_A_T8jB2xNd3_0),.clk(gclk));
	jdff dff_A_dJsbkDX95_0(.dout(w_dff_A_axCQjWg46_0),.din(w_dff_A_dJsbkDX95_0),.clk(gclk));
	jdff dff_A_axCQjWg46_0(.dout(w_dff_A_FjIr2JJr1_0),.din(w_dff_A_axCQjWg46_0),.clk(gclk));
	jdff dff_A_FjIr2JJr1_0(.dout(w_dff_A_zInnHBRp3_0),.din(w_dff_A_FjIr2JJr1_0),.clk(gclk));
	jdff dff_A_zInnHBRp3_0(.dout(w_dff_A_yBWDkHuo3_0),.din(w_dff_A_zInnHBRp3_0),.clk(gclk));
	jdff dff_A_yBWDkHuo3_0(.dout(w_dff_A_xuEmGywE2_0),.din(w_dff_A_yBWDkHuo3_0),.clk(gclk));
	jdff dff_A_xuEmGywE2_0(.dout(w_dff_A_5OVNLf8I4_0),.din(w_dff_A_xuEmGywE2_0),.clk(gclk));
	jdff dff_A_5OVNLf8I4_0(.dout(w_dff_A_oHn3GFpu5_0),.din(w_dff_A_5OVNLf8I4_0),.clk(gclk));
	jdff dff_A_oHn3GFpu5_0(.dout(w_dff_A_zEXVDgTy4_0),.din(w_dff_A_oHn3GFpu5_0),.clk(gclk));
	jdff dff_A_zEXVDgTy4_0(.dout(w_dff_A_0fTmNK6w1_0),.din(w_dff_A_zEXVDgTy4_0),.clk(gclk));
	jdff dff_A_0fTmNK6w1_0(.dout(w_dff_A_PW9dBE841_0),.din(w_dff_A_0fTmNK6w1_0),.clk(gclk));
	jdff dff_A_PW9dBE841_0(.dout(w_dff_A_h5mQSizS4_0),.din(w_dff_A_PW9dBE841_0),.clk(gclk));
	jdff dff_A_h5mQSizS4_0(.dout(w_dff_A_cROyc4D50_0),.din(w_dff_A_h5mQSizS4_0),.clk(gclk));
	jdff dff_A_cROyc4D50_0(.dout(w_dff_A_ZInPEIfL0_0),.din(w_dff_A_cROyc4D50_0),.clk(gclk));
	jdff dff_A_ZInPEIfL0_0(.dout(w_dff_A_5DMb0lvz5_0),.din(w_dff_A_ZInPEIfL0_0),.clk(gclk));
	jdff dff_A_5DMb0lvz5_0(.dout(G536),.din(w_dff_A_5DMb0lvz5_0),.clk(gclk));
	jdff dff_A_Y0XsnTNc9_1(.dout(w_dff_A_T7a8vy667_0),.din(w_dff_A_Y0XsnTNc9_1),.clk(gclk));
	jdff dff_A_T7a8vy667_0(.dout(w_dff_A_QjisMclL7_0),.din(w_dff_A_T7a8vy667_0),.clk(gclk));
	jdff dff_A_QjisMclL7_0(.dout(w_dff_A_V1nFNSGM9_0),.din(w_dff_A_QjisMclL7_0),.clk(gclk));
	jdff dff_A_V1nFNSGM9_0(.dout(w_dff_A_l7ShLEp08_0),.din(w_dff_A_V1nFNSGM9_0),.clk(gclk));
	jdff dff_A_l7ShLEp08_0(.dout(w_dff_A_ogvvfXQc4_0),.din(w_dff_A_l7ShLEp08_0),.clk(gclk));
	jdff dff_A_ogvvfXQc4_0(.dout(w_dff_A_daaCWMT53_0),.din(w_dff_A_ogvvfXQc4_0),.clk(gclk));
	jdff dff_A_daaCWMT53_0(.dout(w_dff_A_cbH8fffg2_0),.din(w_dff_A_daaCWMT53_0),.clk(gclk));
	jdff dff_A_cbH8fffg2_0(.dout(w_dff_A_YKAcz1qg2_0),.din(w_dff_A_cbH8fffg2_0),.clk(gclk));
	jdff dff_A_YKAcz1qg2_0(.dout(w_dff_A_YYzpSPer0_0),.din(w_dff_A_YKAcz1qg2_0),.clk(gclk));
	jdff dff_A_YYzpSPer0_0(.dout(w_dff_A_WbSzd5fG5_0),.din(w_dff_A_YYzpSPer0_0),.clk(gclk));
	jdff dff_A_WbSzd5fG5_0(.dout(w_dff_A_Vxafupq79_0),.din(w_dff_A_WbSzd5fG5_0),.clk(gclk));
	jdff dff_A_Vxafupq79_0(.dout(w_dff_A_obNLe7ck8_0),.din(w_dff_A_Vxafupq79_0),.clk(gclk));
	jdff dff_A_obNLe7ck8_0(.dout(w_dff_A_RRVBhwzk0_0),.din(w_dff_A_obNLe7ck8_0),.clk(gclk));
	jdff dff_A_RRVBhwzk0_0(.dout(w_dff_A_sZ87DjIv2_0),.din(w_dff_A_RRVBhwzk0_0),.clk(gclk));
	jdff dff_A_sZ87DjIv2_0(.dout(w_dff_A_7vDfyxsn6_0),.din(w_dff_A_sZ87DjIv2_0),.clk(gclk));
	jdff dff_A_7vDfyxsn6_0(.dout(w_dff_A_puks27fJ6_0),.din(w_dff_A_7vDfyxsn6_0),.clk(gclk));
	jdff dff_A_puks27fJ6_0(.dout(w_dff_A_TCDd4YRd4_0),.din(w_dff_A_puks27fJ6_0),.clk(gclk));
	jdff dff_A_TCDd4YRd4_0(.dout(w_dff_A_gopMhbKD8_0),.din(w_dff_A_TCDd4YRd4_0),.clk(gclk));
	jdff dff_A_gopMhbKD8_0(.dout(w_dff_A_ZX7d4pxK9_0),.din(w_dff_A_gopMhbKD8_0),.clk(gclk));
	jdff dff_A_ZX7d4pxK9_0(.dout(w_dff_A_fPIXqN9E5_0),.din(w_dff_A_ZX7d4pxK9_0),.clk(gclk));
	jdff dff_A_fPIXqN9E5_0(.dout(w_dff_A_LSPT52hn1_0),.din(w_dff_A_fPIXqN9E5_0),.clk(gclk));
	jdff dff_A_LSPT52hn1_0(.dout(w_dff_A_GqLBgOHo7_0),.din(w_dff_A_LSPT52hn1_0),.clk(gclk));
	jdff dff_A_GqLBgOHo7_0(.dout(w_dff_A_j42bWZsS5_0),.din(w_dff_A_GqLBgOHo7_0),.clk(gclk));
	jdff dff_A_j42bWZsS5_0(.dout(w_dff_A_M8vHD1Ac8_0),.din(w_dff_A_j42bWZsS5_0),.clk(gclk));
	jdff dff_A_M8vHD1Ac8_0(.dout(w_dff_A_O4HCTYPZ1_0),.din(w_dff_A_M8vHD1Ac8_0),.clk(gclk));
	jdff dff_A_O4HCTYPZ1_0(.dout(w_dff_A_pd5eUize2_0),.din(w_dff_A_O4HCTYPZ1_0),.clk(gclk));
	jdff dff_A_pd5eUize2_0(.dout(w_dff_A_y6qSF2Ev1_0),.din(w_dff_A_pd5eUize2_0),.clk(gclk));
	jdff dff_A_y6qSF2Ev1_0(.dout(w_dff_A_w3E732Vl5_0),.din(w_dff_A_y6qSF2Ev1_0),.clk(gclk));
	jdff dff_A_w3E732Vl5_0(.dout(w_dff_A_D5suDTaQ3_0),.din(w_dff_A_w3E732Vl5_0),.clk(gclk));
	jdff dff_A_D5suDTaQ3_0(.dout(w_dff_A_bu96vTmr7_0),.din(w_dff_A_D5suDTaQ3_0),.clk(gclk));
	jdff dff_A_bu96vTmr7_0(.dout(w_dff_A_5rZ717lo4_0),.din(w_dff_A_bu96vTmr7_0),.clk(gclk));
	jdff dff_A_5rZ717lo4_0(.dout(w_dff_A_2toj0yy12_0),.din(w_dff_A_5rZ717lo4_0),.clk(gclk));
	jdff dff_A_2toj0yy12_0(.dout(w_dff_A_vcT4gfum4_0),.din(w_dff_A_2toj0yy12_0),.clk(gclk));
	jdff dff_A_vcT4gfum4_0(.dout(w_dff_A_xovUDJzy7_0),.din(w_dff_A_vcT4gfum4_0),.clk(gclk));
	jdff dff_A_xovUDJzy7_0(.dout(w_dff_A_2Pbeh5Cg0_0),.din(w_dff_A_xovUDJzy7_0),.clk(gclk));
	jdff dff_A_2Pbeh5Cg0_0(.dout(w_dff_A_aPMfGfWe8_0),.din(w_dff_A_2Pbeh5Cg0_0),.clk(gclk));
	jdff dff_A_aPMfGfWe8_0(.dout(w_dff_A_P0SWuub67_0),.din(w_dff_A_aPMfGfWe8_0),.clk(gclk));
	jdff dff_A_P0SWuub67_0(.dout(w_dff_A_yVsYAMKi6_0),.din(w_dff_A_P0SWuub67_0),.clk(gclk));
	jdff dff_A_yVsYAMKi6_0(.dout(G534),.din(w_dff_A_yVsYAMKi6_0),.clk(gclk));
	jdff dff_A_o22oslEs2_1(.dout(w_dff_A_SWudl3fH6_0),.din(w_dff_A_o22oslEs2_1),.clk(gclk));
	jdff dff_A_SWudl3fH6_0(.dout(w_dff_A_kFYwmWPx8_0),.din(w_dff_A_SWudl3fH6_0),.clk(gclk));
	jdff dff_A_kFYwmWPx8_0(.dout(w_dff_A_GjjemOjO5_0),.din(w_dff_A_kFYwmWPx8_0),.clk(gclk));
	jdff dff_A_GjjemOjO5_0(.dout(w_dff_A_Wd24Repo5_0),.din(w_dff_A_GjjemOjO5_0),.clk(gclk));
	jdff dff_A_Wd24Repo5_0(.dout(w_dff_A_mcIabQoo0_0),.din(w_dff_A_Wd24Repo5_0),.clk(gclk));
	jdff dff_A_mcIabQoo0_0(.dout(w_dff_A_vNWVtsxY0_0),.din(w_dff_A_mcIabQoo0_0),.clk(gclk));
	jdff dff_A_vNWVtsxY0_0(.dout(w_dff_A_LbyYWF4Z8_0),.din(w_dff_A_vNWVtsxY0_0),.clk(gclk));
	jdff dff_A_LbyYWF4Z8_0(.dout(w_dff_A_SNaNUHVy7_0),.din(w_dff_A_LbyYWF4Z8_0),.clk(gclk));
	jdff dff_A_SNaNUHVy7_0(.dout(w_dff_A_iLDs1PeX6_0),.din(w_dff_A_SNaNUHVy7_0),.clk(gclk));
	jdff dff_A_iLDs1PeX6_0(.dout(w_dff_A_icN3eGbN8_0),.din(w_dff_A_iLDs1PeX6_0),.clk(gclk));
	jdff dff_A_icN3eGbN8_0(.dout(w_dff_A_3qNU8Oj16_0),.din(w_dff_A_icN3eGbN8_0),.clk(gclk));
	jdff dff_A_3qNU8Oj16_0(.dout(w_dff_A_iGRTyvPk4_0),.din(w_dff_A_3qNU8Oj16_0),.clk(gclk));
	jdff dff_A_iGRTyvPk4_0(.dout(w_dff_A_lrSiQmtD4_0),.din(w_dff_A_iGRTyvPk4_0),.clk(gclk));
	jdff dff_A_lrSiQmtD4_0(.dout(w_dff_A_yN2i2zPk7_0),.din(w_dff_A_lrSiQmtD4_0),.clk(gclk));
	jdff dff_A_yN2i2zPk7_0(.dout(w_dff_A_Lt70lOct4_0),.din(w_dff_A_yN2i2zPk7_0),.clk(gclk));
	jdff dff_A_Lt70lOct4_0(.dout(w_dff_A_UE6mAHTh1_0),.din(w_dff_A_Lt70lOct4_0),.clk(gclk));
	jdff dff_A_UE6mAHTh1_0(.dout(w_dff_A_MvkKaeaj4_0),.din(w_dff_A_UE6mAHTh1_0),.clk(gclk));
	jdff dff_A_MvkKaeaj4_0(.dout(w_dff_A_tgX9iR9T3_0),.din(w_dff_A_MvkKaeaj4_0),.clk(gclk));
	jdff dff_A_tgX9iR9T3_0(.dout(w_dff_A_OmA1Ya523_0),.din(w_dff_A_tgX9iR9T3_0),.clk(gclk));
	jdff dff_A_OmA1Ya523_0(.dout(w_dff_A_aw5W9kgK5_0),.din(w_dff_A_OmA1Ya523_0),.clk(gclk));
	jdff dff_A_aw5W9kgK5_0(.dout(w_dff_A_QxQyy5JU8_0),.din(w_dff_A_aw5W9kgK5_0),.clk(gclk));
	jdff dff_A_QxQyy5JU8_0(.dout(w_dff_A_mVzhrwoW5_0),.din(w_dff_A_QxQyy5JU8_0),.clk(gclk));
	jdff dff_A_mVzhrwoW5_0(.dout(w_dff_A_fBcNLUnm6_0),.din(w_dff_A_mVzhrwoW5_0),.clk(gclk));
	jdff dff_A_fBcNLUnm6_0(.dout(w_dff_A_v2B4HLeQ0_0),.din(w_dff_A_fBcNLUnm6_0),.clk(gclk));
	jdff dff_A_v2B4HLeQ0_0(.dout(w_dff_A_4IbIkKsT0_0),.din(w_dff_A_v2B4HLeQ0_0),.clk(gclk));
	jdff dff_A_4IbIkKsT0_0(.dout(w_dff_A_Hg0LsFs22_0),.din(w_dff_A_4IbIkKsT0_0),.clk(gclk));
	jdff dff_A_Hg0LsFs22_0(.dout(w_dff_A_jxZF3BAR8_0),.din(w_dff_A_Hg0LsFs22_0),.clk(gclk));
	jdff dff_A_jxZF3BAR8_0(.dout(w_dff_A_PSWajxFq8_0),.din(w_dff_A_jxZF3BAR8_0),.clk(gclk));
	jdff dff_A_PSWajxFq8_0(.dout(w_dff_A_3cptEHxw6_0),.din(w_dff_A_PSWajxFq8_0),.clk(gclk));
	jdff dff_A_3cptEHxw6_0(.dout(w_dff_A_DNGDY2Ph1_0),.din(w_dff_A_3cptEHxw6_0),.clk(gclk));
	jdff dff_A_DNGDY2Ph1_0(.dout(w_dff_A_FCCMkWCz6_0),.din(w_dff_A_DNGDY2Ph1_0),.clk(gclk));
	jdff dff_A_FCCMkWCz6_0(.dout(w_dff_A_suDbfMfF5_0),.din(w_dff_A_FCCMkWCz6_0),.clk(gclk));
	jdff dff_A_suDbfMfF5_0(.dout(w_dff_A_BIMIoinK2_0),.din(w_dff_A_suDbfMfF5_0),.clk(gclk));
	jdff dff_A_BIMIoinK2_0(.dout(w_dff_A_Qmvh1YgZ5_0),.din(w_dff_A_BIMIoinK2_0),.clk(gclk));
	jdff dff_A_Qmvh1YgZ5_0(.dout(w_dff_A_ma8oUp8w2_0),.din(w_dff_A_Qmvh1YgZ5_0),.clk(gclk));
	jdff dff_A_ma8oUp8w2_0(.dout(w_dff_A_ODou38dY2_0),.din(w_dff_A_ma8oUp8w2_0),.clk(gclk));
	jdff dff_A_ODou38dY2_0(.dout(w_dff_A_krEJdneQ4_0),.din(w_dff_A_ODou38dY2_0),.clk(gclk));
	jdff dff_A_krEJdneQ4_0(.dout(w_dff_A_Hf7d0RiV9_0),.din(w_dff_A_krEJdneQ4_0),.clk(gclk));
	jdff dff_A_Hf7d0RiV9_0(.dout(G532),.din(w_dff_A_Hf7d0RiV9_0),.clk(gclk));
	jdff dff_A_HR72Rhmh8_1(.dout(w_dff_A_L4mAU5u48_0),.din(w_dff_A_HR72Rhmh8_1),.clk(gclk));
	jdff dff_A_L4mAU5u48_0(.dout(w_dff_A_Up0ZXbfK1_0),.din(w_dff_A_L4mAU5u48_0),.clk(gclk));
	jdff dff_A_Up0ZXbfK1_0(.dout(w_dff_A_aCiQFfaL4_0),.din(w_dff_A_Up0ZXbfK1_0),.clk(gclk));
	jdff dff_A_aCiQFfaL4_0(.dout(w_dff_A_NOXl3xAN5_0),.din(w_dff_A_aCiQFfaL4_0),.clk(gclk));
	jdff dff_A_NOXl3xAN5_0(.dout(w_dff_A_JXLM4iq89_0),.din(w_dff_A_NOXl3xAN5_0),.clk(gclk));
	jdff dff_A_JXLM4iq89_0(.dout(w_dff_A_UaeNUpip8_0),.din(w_dff_A_JXLM4iq89_0),.clk(gclk));
	jdff dff_A_UaeNUpip8_0(.dout(w_dff_A_HjgzRhnt0_0),.din(w_dff_A_UaeNUpip8_0),.clk(gclk));
	jdff dff_A_HjgzRhnt0_0(.dout(w_dff_A_6lXovPbp7_0),.din(w_dff_A_HjgzRhnt0_0),.clk(gclk));
	jdff dff_A_6lXovPbp7_0(.dout(w_dff_A_O9BjyBi62_0),.din(w_dff_A_6lXovPbp7_0),.clk(gclk));
	jdff dff_A_O9BjyBi62_0(.dout(w_dff_A_ltnuCPoY6_0),.din(w_dff_A_O9BjyBi62_0),.clk(gclk));
	jdff dff_A_ltnuCPoY6_0(.dout(w_dff_A_1dPmnWAJ4_0),.din(w_dff_A_ltnuCPoY6_0),.clk(gclk));
	jdff dff_A_1dPmnWAJ4_0(.dout(w_dff_A_mljuEguS8_0),.din(w_dff_A_1dPmnWAJ4_0),.clk(gclk));
	jdff dff_A_mljuEguS8_0(.dout(w_dff_A_T7uqPioX1_0),.din(w_dff_A_mljuEguS8_0),.clk(gclk));
	jdff dff_A_T7uqPioX1_0(.dout(w_dff_A_lsku68HW7_0),.din(w_dff_A_T7uqPioX1_0),.clk(gclk));
	jdff dff_A_lsku68HW7_0(.dout(w_dff_A_p1O28qaI2_0),.din(w_dff_A_lsku68HW7_0),.clk(gclk));
	jdff dff_A_p1O28qaI2_0(.dout(w_dff_A_YVGVUQl08_0),.din(w_dff_A_p1O28qaI2_0),.clk(gclk));
	jdff dff_A_YVGVUQl08_0(.dout(w_dff_A_xGPAdEvR3_0),.din(w_dff_A_YVGVUQl08_0),.clk(gclk));
	jdff dff_A_xGPAdEvR3_0(.dout(w_dff_A_gH1sdyky3_0),.din(w_dff_A_xGPAdEvR3_0),.clk(gclk));
	jdff dff_A_gH1sdyky3_0(.dout(w_dff_A_JSSzHHmi4_0),.din(w_dff_A_gH1sdyky3_0),.clk(gclk));
	jdff dff_A_JSSzHHmi4_0(.dout(w_dff_A_o9yy6nCv3_0),.din(w_dff_A_JSSzHHmi4_0),.clk(gclk));
	jdff dff_A_o9yy6nCv3_0(.dout(w_dff_A_LNP5akWZ2_0),.din(w_dff_A_o9yy6nCv3_0),.clk(gclk));
	jdff dff_A_LNP5akWZ2_0(.dout(w_dff_A_q0fcwMf04_0),.din(w_dff_A_LNP5akWZ2_0),.clk(gclk));
	jdff dff_A_q0fcwMf04_0(.dout(w_dff_A_bfcZ9Axs7_0),.din(w_dff_A_q0fcwMf04_0),.clk(gclk));
	jdff dff_A_bfcZ9Axs7_0(.dout(w_dff_A_kwuIIMe07_0),.din(w_dff_A_bfcZ9Axs7_0),.clk(gclk));
	jdff dff_A_kwuIIMe07_0(.dout(w_dff_A_2tNBqF4j3_0),.din(w_dff_A_kwuIIMe07_0),.clk(gclk));
	jdff dff_A_2tNBqF4j3_0(.dout(w_dff_A_ifLkofgn5_0),.din(w_dff_A_2tNBqF4j3_0),.clk(gclk));
	jdff dff_A_ifLkofgn5_0(.dout(w_dff_A_17OsI95U8_0),.din(w_dff_A_ifLkofgn5_0),.clk(gclk));
	jdff dff_A_17OsI95U8_0(.dout(w_dff_A_Bhm3YoXP9_0),.din(w_dff_A_17OsI95U8_0),.clk(gclk));
	jdff dff_A_Bhm3YoXP9_0(.dout(w_dff_A_UD468PUo7_0),.din(w_dff_A_Bhm3YoXP9_0),.clk(gclk));
	jdff dff_A_UD468PUo7_0(.dout(w_dff_A_uWKsv6AY7_0),.din(w_dff_A_UD468PUo7_0),.clk(gclk));
	jdff dff_A_uWKsv6AY7_0(.dout(w_dff_A_fJGcvVX29_0),.din(w_dff_A_uWKsv6AY7_0),.clk(gclk));
	jdff dff_A_fJGcvVX29_0(.dout(w_dff_A_UlHOXTTj5_0),.din(w_dff_A_fJGcvVX29_0),.clk(gclk));
	jdff dff_A_UlHOXTTj5_0(.dout(w_dff_A_0qOKb5Iz9_0),.din(w_dff_A_UlHOXTTj5_0),.clk(gclk));
	jdff dff_A_0qOKb5Iz9_0(.dout(w_dff_A_HSPwinYF8_0),.din(w_dff_A_0qOKb5Iz9_0),.clk(gclk));
	jdff dff_A_HSPwinYF8_0(.dout(w_dff_A_vnHQNcEU3_0),.din(w_dff_A_HSPwinYF8_0),.clk(gclk));
	jdff dff_A_vnHQNcEU3_0(.dout(w_dff_A_I4409HAU4_0),.din(w_dff_A_vnHQNcEU3_0),.clk(gclk));
	jdff dff_A_I4409HAU4_0(.dout(w_dff_A_CWbfRxkb1_0),.din(w_dff_A_I4409HAU4_0),.clk(gclk));
	jdff dff_A_CWbfRxkb1_0(.dout(w_dff_A_Lh4jv2Bj5_0),.din(w_dff_A_CWbfRxkb1_0),.clk(gclk));
	jdff dff_A_Lh4jv2Bj5_0(.dout(G530),.din(w_dff_A_Lh4jv2Bj5_0),.clk(gclk));
	jdff dff_A_p7sM1NwD4_1(.dout(w_dff_A_ZwzT2qxk8_0),.din(w_dff_A_p7sM1NwD4_1),.clk(gclk));
	jdff dff_A_ZwzT2qxk8_0(.dout(w_dff_A_60tzlkKa4_0),.din(w_dff_A_ZwzT2qxk8_0),.clk(gclk));
	jdff dff_A_60tzlkKa4_0(.dout(w_dff_A_M8i6pD6M0_0),.din(w_dff_A_60tzlkKa4_0),.clk(gclk));
	jdff dff_A_M8i6pD6M0_0(.dout(w_dff_A_DJpZwrAq2_0),.din(w_dff_A_M8i6pD6M0_0),.clk(gclk));
	jdff dff_A_DJpZwrAq2_0(.dout(w_dff_A_BV8BsgHy2_0),.din(w_dff_A_DJpZwrAq2_0),.clk(gclk));
	jdff dff_A_BV8BsgHy2_0(.dout(w_dff_A_XOhjJSgs0_0),.din(w_dff_A_BV8BsgHy2_0),.clk(gclk));
	jdff dff_A_XOhjJSgs0_0(.dout(w_dff_A_3nNodtXk4_0),.din(w_dff_A_XOhjJSgs0_0),.clk(gclk));
	jdff dff_A_3nNodtXk4_0(.dout(w_dff_A_CdQnmaiK3_0),.din(w_dff_A_3nNodtXk4_0),.clk(gclk));
	jdff dff_A_CdQnmaiK3_0(.dout(w_dff_A_34PWiVlI1_0),.din(w_dff_A_CdQnmaiK3_0),.clk(gclk));
	jdff dff_A_34PWiVlI1_0(.dout(w_dff_A_5Be4p3Dh1_0),.din(w_dff_A_34PWiVlI1_0),.clk(gclk));
	jdff dff_A_5Be4p3Dh1_0(.dout(w_dff_A_36NETdFm6_0),.din(w_dff_A_5Be4p3Dh1_0),.clk(gclk));
	jdff dff_A_36NETdFm6_0(.dout(w_dff_A_Q8eqRP257_0),.din(w_dff_A_36NETdFm6_0),.clk(gclk));
	jdff dff_A_Q8eqRP257_0(.dout(w_dff_A_iWGNhWis4_0),.din(w_dff_A_Q8eqRP257_0),.clk(gclk));
	jdff dff_A_iWGNhWis4_0(.dout(w_dff_A_qsE37HYN4_0),.din(w_dff_A_iWGNhWis4_0),.clk(gclk));
	jdff dff_A_qsE37HYN4_0(.dout(w_dff_A_PsNvbgbS2_0),.din(w_dff_A_qsE37HYN4_0),.clk(gclk));
	jdff dff_A_PsNvbgbS2_0(.dout(w_dff_A_A8yPce9r5_0),.din(w_dff_A_PsNvbgbS2_0),.clk(gclk));
	jdff dff_A_A8yPce9r5_0(.dout(w_dff_A_DSKIPWAX9_0),.din(w_dff_A_A8yPce9r5_0),.clk(gclk));
	jdff dff_A_DSKIPWAX9_0(.dout(w_dff_A_5I0lhWkl6_0),.din(w_dff_A_DSKIPWAX9_0),.clk(gclk));
	jdff dff_A_5I0lhWkl6_0(.dout(w_dff_A_hHgjl12u8_0),.din(w_dff_A_5I0lhWkl6_0),.clk(gclk));
	jdff dff_A_hHgjl12u8_0(.dout(w_dff_A_tS3kruGW0_0),.din(w_dff_A_hHgjl12u8_0),.clk(gclk));
	jdff dff_A_tS3kruGW0_0(.dout(w_dff_A_G6YL1vPH1_0),.din(w_dff_A_tS3kruGW0_0),.clk(gclk));
	jdff dff_A_G6YL1vPH1_0(.dout(w_dff_A_DEhrCFrZ9_0),.din(w_dff_A_G6YL1vPH1_0),.clk(gclk));
	jdff dff_A_DEhrCFrZ9_0(.dout(w_dff_A_dXGZVzsO6_0),.din(w_dff_A_DEhrCFrZ9_0),.clk(gclk));
	jdff dff_A_dXGZVzsO6_0(.dout(w_dff_A_rSHqQfRY7_0),.din(w_dff_A_dXGZVzsO6_0),.clk(gclk));
	jdff dff_A_rSHqQfRY7_0(.dout(w_dff_A_ZOlQ0VHj1_0),.din(w_dff_A_rSHqQfRY7_0),.clk(gclk));
	jdff dff_A_ZOlQ0VHj1_0(.dout(w_dff_A_k866hyE98_0),.din(w_dff_A_ZOlQ0VHj1_0),.clk(gclk));
	jdff dff_A_k866hyE98_0(.dout(w_dff_A_woUojX6s0_0),.din(w_dff_A_k866hyE98_0),.clk(gclk));
	jdff dff_A_woUojX6s0_0(.dout(w_dff_A_LKGX8AmU1_0),.din(w_dff_A_woUojX6s0_0),.clk(gclk));
	jdff dff_A_LKGX8AmU1_0(.dout(w_dff_A_dgIvbyZM9_0),.din(w_dff_A_LKGX8AmU1_0),.clk(gclk));
	jdff dff_A_dgIvbyZM9_0(.dout(w_dff_A_mhqGb4EO9_0),.din(w_dff_A_dgIvbyZM9_0),.clk(gclk));
	jdff dff_A_mhqGb4EO9_0(.dout(w_dff_A_CijkUDh53_0),.din(w_dff_A_mhqGb4EO9_0),.clk(gclk));
	jdff dff_A_CijkUDh53_0(.dout(w_dff_A_vAxk4ePj9_0),.din(w_dff_A_CijkUDh53_0),.clk(gclk));
	jdff dff_A_vAxk4ePj9_0(.dout(w_dff_A_VyuPYwbb9_0),.din(w_dff_A_vAxk4ePj9_0),.clk(gclk));
	jdff dff_A_VyuPYwbb9_0(.dout(w_dff_A_hWwlbegk8_0),.din(w_dff_A_VyuPYwbb9_0),.clk(gclk));
	jdff dff_A_hWwlbegk8_0(.dout(w_dff_A_JByeqisy2_0),.din(w_dff_A_hWwlbegk8_0),.clk(gclk));
	jdff dff_A_JByeqisy2_0(.dout(w_dff_A_a1bUKP9I2_0),.din(w_dff_A_JByeqisy2_0),.clk(gclk));
	jdff dff_A_a1bUKP9I2_0(.dout(w_dff_A_4hl7L4aQ1_0),.din(w_dff_A_a1bUKP9I2_0),.clk(gclk));
	jdff dff_A_4hl7L4aQ1_0(.dout(w_dff_A_eHE9IdWZ8_0),.din(w_dff_A_4hl7L4aQ1_0),.clk(gclk));
	jdff dff_A_eHE9IdWZ8_0(.dout(G528),.din(w_dff_A_eHE9IdWZ8_0),.clk(gclk));
	jdff dff_A_vAZbA4Z74_1(.dout(w_dff_A_2MMp62kH6_0),.din(w_dff_A_vAZbA4Z74_1),.clk(gclk));
	jdff dff_A_2MMp62kH6_0(.dout(w_dff_A_Uezq7o1B3_0),.din(w_dff_A_2MMp62kH6_0),.clk(gclk));
	jdff dff_A_Uezq7o1B3_0(.dout(w_dff_A_BhLPUd8a5_0),.din(w_dff_A_Uezq7o1B3_0),.clk(gclk));
	jdff dff_A_BhLPUd8a5_0(.dout(w_dff_A_DjgBeDDH9_0),.din(w_dff_A_BhLPUd8a5_0),.clk(gclk));
	jdff dff_A_DjgBeDDH9_0(.dout(w_dff_A_PGkMPdFJ2_0),.din(w_dff_A_DjgBeDDH9_0),.clk(gclk));
	jdff dff_A_PGkMPdFJ2_0(.dout(w_dff_A_yEbciAXi2_0),.din(w_dff_A_PGkMPdFJ2_0),.clk(gclk));
	jdff dff_A_yEbciAXi2_0(.dout(w_dff_A_dbq3GH680_0),.din(w_dff_A_yEbciAXi2_0),.clk(gclk));
	jdff dff_A_dbq3GH680_0(.dout(w_dff_A_xEQ4c4kd0_0),.din(w_dff_A_dbq3GH680_0),.clk(gclk));
	jdff dff_A_xEQ4c4kd0_0(.dout(w_dff_A_4M4XRUCz6_0),.din(w_dff_A_xEQ4c4kd0_0),.clk(gclk));
	jdff dff_A_4M4XRUCz6_0(.dout(w_dff_A_SgUjyxAP9_0),.din(w_dff_A_4M4XRUCz6_0),.clk(gclk));
	jdff dff_A_SgUjyxAP9_0(.dout(w_dff_A_vrW4C4ix7_0),.din(w_dff_A_SgUjyxAP9_0),.clk(gclk));
	jdff dff_A_vrW4C4ix7_0(.dout(w_dff_A_m7BdAZj59_0),.din(w_dff_A_vrW4C4ix7_0),.clk(gclk));
	jdff dff_A_m7BdAZj59_0(.dout(w_dff_A_3kbH9r0a1_0),.din(w_dff_A_m7BdAZj59_0),.clk(gclk));
	jdff dff_A_3kbH9r0a1_0(.dout(w_dff_A_0AAUV0yJ2_0),.din(w_dff_A_3kbH9r0a1_0),.clk(gclk));
	jdff dff_A_0AAUV0yJ2_0(.dout(w_dff_A_pjfqcciz7_0),.din(w_dff_A_0AAUV0yJ2_0),.clk(gclk));
	jdff dff_A_pjfqcciz7_0(.dout(w_dff_A_8wtueMno8_0),.din(w_dff_A_pjfqcciz7_0),.clk(gclk));
	jdff dff_A_8wtueMno8_0(.dout(w_dff_A_WB0DWFEg4_0),.din(w_dff_A_8wtueMno8_0),.clk(gclk));
	jdff dff_A_WB0DWFEg4_0(.dout(w_dff_A_gjvpN5Wr2_0),.din(w_dff_A_WB0DWFEg4_0),.clk(gclk));
	jdff dff_A_gjvpN5Wr2_0(.dout(w_dff_A_QbzNtfmz9_0),.din(w_dff_A_gjvpN5Wr2_0),.clk(gclk));
	jdff dff_A_QbzNtfmz9_0(.dout(w_dff_A_Pugu3RvD2_0),.din(w_dff_A_QbzNtfmz9_0),.clk(gclk));
	jdff dff_A_Pugu3RvD2_0(.dout(w_dff_A_dw9GOxEv1_0),.din(w_dff_A_Pugu3RvD2_0),.clk(gclk));
	jdff dff_A_dw9GOxEv1_0(.dout(w_dff_A_AR1CtIRJ8_0),.din(w_dff_A_dw9GOxEv1_0),.clk(gclk));
	jdff dff_A_AR1CtIRJ8_0(.dout(w_dff_A_lh3xLDUg4_0),.din(w_dff_A_AR1CtIRJ8_0),.clk(gclk));
	jdff dff_A_lh3xLDUg4_0(.dout(w_dff_A_CwQlRBn45_0),.din(w_dff_A_lh3xLDUg4_0),.clk(gclk));
	jdff dff_A_CwQlRBn45_0(.dout(w_dff_A_UUSNmJRB2_0),.din(w_dff_A_CwQlRBn45_0),.clk(gclk));
	jdff dff_A_UUSNmJRB2_0(.dout(w_dff_A_RxD0gh791_0),.din(w_dff_A_UUSNmJRB2_0),.clk(gclk));
	jdff dff_A_RxD0gh791_0(.dout(w_dff_A_GU26L0L16_0),.din(w_dff_A_RxD0gh791_0),.clk(gclk));
	jdff dff_A_GU26L0L16_0(.dout(w_dff_A_Q8SU1OhR9_0),.din(w_dff_A_GU26L0L16_0),.clk(gclk));
	jdff dff_A_Q8SU1OhR9_0(.dout(w_dff_A_7YbTRTcE1_0),.din(w_dff_A_Q8SU1OhR9_0),.clk(gclk));
	jdff dff_A_7YbTRTcE1_0(.dout(w_dff_A_UKvk0YiI1_0),.din(w_dff_A_7YbTRTcE1_0),.clk(gclk));
	jdff dff_A_UKvk0YiI1_0(.dout(w_dff_A_kpItN9ID0_0),.din(w_dff_A_UKvk0YiI1_0),.clk(gclk));
	jdff dff_A_kpItN9ID0_0(.dout(w_dff_A_KwL4tTzp8_0),.din(w_dff_A_kpItN9ID0_0),.clk(gclk));
	jdff dff_A_KwL4tTzp8_0(.dout(w_dff_A_zxTDcH0z3_0),.din(w_dff_A_KwL4tTzp8_0),.clk(gclk));
	jdff dff_A_zxTDcH0z3_0(.dout(w_dff_A_70CmHYck2_0),.din(w_dff_A_zxTDcH0z3_0),.clk(gclk));
	jdff dff_A_70CmHYck2_0(.dout(w_dff_A_fJ82zzi54_0),.din(w_dff_A_70CmHYck2_0),.clk(gclk));
	jdff dff_A_fJ82zzi54_0(.dout(w_dff_A_zAl7ihCX2_0),.din(w_dff_A_fJ82zzi54_0),.clk(gclk));
	jdff dff_A_zAl7ihCX2_0(.dout(w_dff_A_HZt1AhWg5_0),.din(w_dff_A_zAl7ihCX2_0),.clk(gclk));
	jdff dff_A_HZt1AhWg5_0(.dout(w_dff_A_sFNRtXSA0_0),.din(w_dff_A_HZt1AhWg5_0),.clk(gclk));
	jdff dff_A_sFNRtXSA0_0(.dout(G526),.din(w_dff_A_sFNRtXSA0_0),.clk(gclk));
	jdff dff_A_mt2rqSeK3_1(.dout(w_dff_A_xbmFH1iK5_0),.din(w_dff_A_mt2rqSeK3_1),.clk(gclk));
	jdff dff_A_xbmFH1iK5_0(.dout(w_dff_A_xbiJKr2Z6_0),.din(w_dff_A_xbmFH1iK5_0),.clk(gclk));
	jdff dff_A_xbiJKr2Z6_0(.dout(w_dff_A_ofcDf6b19_0),.din(w_dff_A_xbiJKr2Z6_0),.clk(gclk));
	jdff dff_A_ofcDf6b19_0(.dout(w_dff_A_qpW2n5U76_0),.din(w_dff_A_ofcDf6b19_0),.clk(gclk));
	jdff dff_A_qpW2n5U76_0(.dout(w_dff_A_LFeS4H0z5_0),.din(w_dff_A_qpW2n5U76_0),.clk(gclk));
	jdff dff_A_LFeS4H0z5_0(.dout(w_dff_A_qGOcPXK40_0),.din(w_dff_A_LFeS4H0z5_0),.clk(gclk));
	jdff dff_A_qGOcPXK40_0(.dout(w_dff_A_C734e5R69_0),.din(w_dff_A_qGOcPXK40_0),.clk(gclk));
	jdff dff_A_C734e5R69_0(.dout(w_dff_A_ZaUUDSYa3_0),.din(w_dff_A_C734e5R69_0),.clk(gclk));
	jdff dff_A_ZaUUDSYa3_0(.dout(w_dff_A_l3d6zRP65_0),.din(w_dff_A_ZaUUDSYa3_0),.clk(gclk));
	jdff dff_A_l3d6zRP65_0(.dout(w_dff_A_YbJHumxK4_0),.din(w_dff_A_l3d6zRP65_0),.clk(gclk));
	jdff dff_A_YbJHumxK4_0(.dout(w_dff_A_sFKswxqH0_0),.din(w_dff_A_YbJHumxK4_0),.clk(gclk));
	jdff dff_A_sFKswxqH0_0(.dout(w_dff_A_xv7CYBWv2_0),.din(w_dff_A_sFKswxqH0_0),.clk(gclk));
	jdff dff_A_xv7CYBWv2_0(.dout(w_dff_A_79wXGOJO1_0),.din(w_dff_A_xv7CYBWv2_0),.clk(gclk));
	jdff dff_A_79wXGOJO1_0(.dout(w_dff_A_fMCP0aMa3_0),.din(w_dff_A_79wXGOJO1_0),.clk(gclk));
	jdff dff_A_fMCP0aMa3_0(.dout(w_dff_A_VSwDGCem0_0),.din(w_dff_A_fMCP0aMa3_0),.clk(gclk));
	jdff dff_A_VSwDGCem0_0(.dout(w_dff_A_1pvS7Uzg9_0),.din(w_dff_A_VSwDGCem0_0),.clk(gclk));
	jdff dff_A_1pvS7Uzg9_0(.dout(w_dff_A_Tl4ODZsD9_0),.din(w_dff_A_1pvS7Uzg9_0),.clk(gclk));
	jdff dff_A_Tl4ODZsD9_0(.dout(w_dff_A_typFEyuf4_0),.din(w_dff_A_Tl4ODZsD9_0),.clk(gclk));
	jdff dff_A_typFEyuf4_0(.dout(w_dff_A_2tOivj167_0),.din(w_dff_A_typFEyuf4_0),.clk(gclk));
	jdff dff_A_2tOivj167_0(.dout(w_dff_A_lToGJ2b27_0),.din(w_dff_A_2tOivj167_0),.clk(gclk));
	jdff dff_A_lToGJ2b27_0(.dout(w_dff_A_0o5o424W3_0),.din(w_dff_A_lToGJ2b27_0),.clk(gclk));
	jdff dff_A_0o5o424W3_0(.dout(w_dff_A_YOz7mk6i7_0),.din(w_dff_A_0o5o424W3_0),.clk(gclk));
	jdff dff_A_YOz7mk6i7_0(.dout(w_dff_A_rORy3Q6Z9_0),.din(w_dff_A_YOz7mk6i7_0),.clk(gclk));
	jdff dff_A_rORy3Q6Z9_0(.dout(w_dff_A_S9ryIOuu0_0),.din(w_dff_A_rORy3Q6Z9_0),.clk(gclk));
	jdff dff_A_S9ryIOuu0_0(.dout(w_dff_A_YPgn7Exi0_0),.din(w_dff_A_S9ryIOuu0_0),.clk(gclk));
	jdff dff_A_YPgn7Exi0_0(.dout(w_dff_A_dsE7BO5X6_0),.din(w_dff_A_YPgn7Exi0_0),.clk(gclk));
	jdff dff_A_dsE7BO5X6_0(.dout(w_dff_A_rfFe7aCU5_0),.din(w_dff_A_dsE7BO5X6_0),.clk(gclk));
	jdff dff_A_rfFe7aCU5_0(.dout(w_dff_A_a6mlJYpW4_0),.din(w_dff_A_rfFe7aCU5_0),.clk(gclk));
	jdff dff_A_a6mlJYpW4_0(.dout(w_dff_A_MbLrLki79_0),.din(w_dff_A_a6mlJYpW4_0),.clk(gclk));
	jdff dff_A_MbLrLki79_0(.dout(w_dff_A_7XMwCsdi2_0),.din(w_dff_A_MbLrLki79_0),.clk(gclk));
	jdff dff_A_7XMwCsdi2_0(.dout(w_dff_A_KCKSzwGq7_0),.din(w_dff_A_7XMwCsdi2_0),.clk(gclk));
	jdff dff_A_KCKSzwGq7_0(.dout(w_dff_A_zshp0VFt3_0),.din(w_dff_A_KCKSzwGq7_0),.clk(gclk));
	jdff dff_A_zshp0VFt3_0(.dout(w_dff_A_DMiGRzAQ7_0),.din(w_dff_A_zshp0VFt3_0),.clk(gclk));
	jdff dff_A_DMiGRzAQ7_0(.dout(w_dff_A_mtQZz3yC9_0),.din(w_dff_A_DMiGRzAQ7_0),.clk(gclk));
	jdff dff_A_mtQZz3yC9_0(.dout(w_dff_A_ov4lPmoW6_0),.din(w_dff_A_mtQZz3yC9_0),.clk(gclk));
	jdff dff_A_ov4lPmoW6_0(.dout(w_dff_A_KyCXR99V6_0),.din(w_dff_A_ov4lPmoW6_0),.clk(gclk));
	jdff dff_A_KyCXR99V6_0(.dout(w_dff_A_VvZqcXFo5_0),.din(w_dff_A_KyCXR99V6_0),.clk(gclk));
	jdff dff_A_VvZqcXFo5_0(.dout(w_dff_A_PHcpn06L7_0),.din(w_dff_A_VvZqcXFo5_0),.clk(gclk));
	jdff dff_A_PHcpn06L7_0(.dout(G524),.din(w_dff_A_PHcpn06L7_0),.clk(gclk));
	jdff dff_A_TSybH3fu9_1(.dout(w_dff_A_wUfJfbab4_0),.din(w_dff_A_TSybH3fu9_1),.clk(gclk));
	jdff dff_A_wUfJfbab4_0(.dout(w_dff_A_dxnGsKwm7_0),.din(w_dff_A_wUfJfbab4_0),.clk(gclk));
	jdff dff_A_dxnGsKwm7_0(.dout(w_dff_A_111G5MnE0_0),.din(w_dff_A_dxnGsKwm7_0),.clk(gclk));
	jdff dff_A_111G5MnE0_0(.dout(w_dff_A_ruUpCu2q4_0),.din(w_dff_A_111G5MnE0_0),.clk(gclk));
	jdff dff_A_ruUpCu2q4_0(.dout(w_dff_A_iviRMjc33_0),.din(w_dff_A_ruUpCu2q4_0),.clk(gclk));
	jdff dff_A_iviRMjc33_0(.dout(w_dff_A_YM5RG50y9_0),.din(w_dff_A_iviRMjc33_0),.clk(gclk));
	jdff dff_A_YM5RG50y9_0(.dout(w_dff_A_ueBud0cC9_0),.din(w_dff_A_YM5RG50y9_0),.clk(gclk));
	jdff dff_A_ueBud0cC9_0(.dout(w_dff_A_k6wISBbL2_0),.din(w_dff_A_ueBud0cC9_0),.clk(gclk));
	jdff dff_A_k6wISBbL2_0(.dout(w_dff_A_0IzXZe2J3_0),.din(w_dff_A_k6wISBbL2_0),.clk(gclk));
	jdff dff_A_0IzXZe2J3_0(.dout(w_dff_A_dGVSNvSl7_0),.din(w_dff_A_0IzXZe2J3_0),.clk(gclk));
	jdff dff_A_dGVSNvSl7_0(.dout(w_dff_A_O5oDpgQH9_0),.din(w_dff_A_dGVSNvSl7_0),.clk(gclk));
	jdff dff_A_O5oDpgQH9_0(.dout(w_dff_A_0b6JbqDN7_0),.din(w_dff_A_O5oDpgQH9_0),.clk(gclk));
	jdff dff_A_0b6JbqDN7_0(.dout(w_dff_A_vgVSCNHd1_0),.din(w_dff_A_0b6JbqDN7_0),.clk(gclk));
	jdff dff_A_vgVSCNHd1_0(.dout(w_dff_A_Pv71OZNk7_0),.din(w_dff_A_vgVSCNHd1_0),.clk(gclk));
	jdff dff_A_Pv71OZNk7_0(.dout(w_dff_A_NhKCvbut6_0),.din(w_dff_A_Pv71OZNk7_0),.clk(gclk));
	jdff dff_A_NhKCvbut6_0(.dout(w_dff_A_C3Qvz7a30_0),.din(w_dff_A_NhKCvbut6_0),.clk(gclk));
	jdff dff_A_C3Qvz7a30_0(.dout(w_dff_A_LC7wDpGe7_0),.din(w_dff_A_C3Qvz7a30_0),.clk(gclk));
	jdff dff_A_LC7wDpGe7_0(.dout(w_dff_A_6BkqTbXD3_0),.din(w_dff_A_LC7wDpGe7_0),.clk(gclk));
	jdff dff_A_6BkqTbXD3_0(.dout(w_dff_A_NFdnTzuk7_0),.din(w_dff_A_6BkqTbXD3_0),.clk(gclk));
	jdff dff_A_NFdnTzuk7_0(.dout(w_dff_A_p78Ohcai2_0),.din(w_dff_A_NFdnTzuk7_0),.clk(gclk));
	jdff dff_A_p78Ohcai2_0(.dout(w_dff_A_zvbxpQgT1_0),.din(w_dff_A_p78Ohcai2_0),.clk(gclk));
	jdff dff_A_zvbxpQgT1_0(.dout(w_dff_A_voC7HsMn0_0),.din(w_dff_A_zvbxpQgT1_0),.clk(gclk));
	jdff dff_A_voC7HsMn0_0(.dout(w_dff_A_7BzzUeIZ2_0),.din(w_dff_A_voC7HsMn0_0),.clk(gclk));
	jdff dff_A_7BzzUeIZ2_0(.dout(w_dff_A_qz6BamNr6_0),.din(w_dff_A_7BzzUeIZ2_0),.clk(gclk));
	jdff dff_A_qz6BamNr6_0(.dout(w_dff_A_4uXHtAva8_0),.din(w_dff_A_qz6BamNr6_0),.clk(gclk));
	jdff dff_A_4uXHtAva8_0(.dout(w_dff_A_DMAjX8Vy8_0),.din(w_dff_A_4uXHtAva8_0),.clk(gclk));
	jdff dff_A_DMAjX8Vy8_0(.dout(w_dff_A_K06MPBqo0_0),.din(w_dff_A_DMAjX8Vy8_0),.clk(gclk));
	jdff dff_A_K06MPBqo0_0(.dout(w_dff_A_cpZusPVZ8_0),.din(w_dff_A_K06MPBqo0_0),.clk(gclk));
	jdff dff_A_cpZusPVZ8_0(.dout(w_dff_A_hX9yW4Hs7_0),.din(w_dff_A_cpZusPVZ8_0),.clk(gclk));
	jdff dff_A_hX9yW4Hs7_0(.dout(w_dff_A_17jpNigM5_0),.din(w_dff_A_hX9yW4Hs7_0),.clk(gclk));
	jdff dff_A_17jpNigM5_0(.dout(w_dff_A_PABwR32d7_0),.din(w_dff_A_17jpNigM5_0),.clk(gclk));
	jdff dff_A_PABwR32d7_0(.dout(w_dff_A_EHAb92WK2_0),.din(w_dff_A_PABwR32d7_0),.clk(gclk));
	jdff dff_A_EHAb92WK2_0(.dout(w_dff_A_nsGyaO1J4_0),.din(w_dff_A_EHAb92WK2_0),.clk(gclk));
	jdff dff_A_nsGyaO1J4_0(.dout(w_dff_A_yiwkFo8X6_0),.din(w_dff_A_nsGyaO1J4_0),.clk(gclk));
	jdff dff_A_yiwkFo8X6_0(.dout(w_dff_A_Ii6OrUsK4_0),.din(w_dff_A_yiwkFo8X6_0),.clk(gclk));
	jdff dff_A_Ii6OrUsK4_0(.dout(w_dff_A_iuSd4yFD0_0),.din(w_dff_A_Ii6OrUsK4_0),.clk(gclk));
	jdff dff_A_iuSd4yFD0_0(.dout(w_dff_A_F8U0IhfW5_0),.din(w_dff_A_iuSd4yFD0_0),.clk(gclk));
	jdff dff_A_F8U0IhfW5_0(.dout(G279),.din(w_dff_A_F8U0IhfW5_0),.clk(gclk));
	jdff dff_A_l1LtiW1L5_1(.dout(w_dff_A_n2eZmFw13_0),.din(w_dff_A_l1LtiW1L5_1),.clk(gclk));
	jdff dff_A_n2eZmFw13_0(.dout(w_dff_A_VD6nyx6i9_0),.din(w_dff_A_n2eZmFw13_0),.clk(gclk));
	jdff dff_A_VD6nyx6i9_0(.dout(w_dff_A_0ZU42tqb6_0),.din(w_dff_A_VD6nyx6i9_0),.clk(gclk));
	jdff dff_A_0ZU42tqb6_0(.dout(w_dff_A_oHR3riFy7_0),.din(w_dff_A_0ZU42tqb6_0),.clk(gclk));
	jdff dff_A_oHR3riFy7_0(.dout(w_dff_A_fyxfenTr9_0),.din(w_dff_A_oHR3riFy7_0),.clk(gclk));
	jdff dff_A_fyxfenTr9_0(.dout(w_dff_A_c8uAtUer9_0),.din(w_dff_A_fyxfenTr9_0),.clk(gclk));
	jdff dff_A_c8uAtUer9_0(.dout(w_dff_A_hItoQ4gS7_0),.din(w_dff_A_c8uAtUer9_0),.clk(gclk));
	jdff dff_A_hItoQ4gS7_0(.dout(w_dff_A_sWW8MIeX3_0),.din(w_dff_A_hItoQ4gS7_0),.clk(gclk));
	jdff dff_A_sWW8MIeX3_0(.dout(w_dff_A_z7J0neZo6_0),.din(w_dff_A_sWW8MIeX3_0),.clk(gclk));
	jdff dff_A_z7J0neZo6_0(.dout(w_dff_A_aSMoqDED7_0),.din(w_dff_A_z7J0neZo6_0),.clk(gclk));
	jdff dff_A_aSMoqDED7_0(.dout(w_dff_A_zCw2bg9x2_0),.din(w_dff_A_aSMoqDED7_0),.clk(gclk));
	jdff dff_A_zCw2bg9x2_0(.dout(w_dff_A_oJswhKXS1_0),.din(w_dff_A_zCw2bg9x2_0),.clk(gclk));
	jdff dff_A_oJswhKXS1_0(.dout(w_dff_A_lnHBadhK4_0),.din(w_dff_A_oJswhKXS1_0),.clk(gclk));
	jdff dff_A_lnHBadhK4_0(.dout(w_dff_A_eK7qKMgm7_0),.din(w_dff_A_lnHBadhK4_0),.clk(gclk));
	jdff dff_A_eK7qKMgm7_0(.dout(w_dff_A_ON5FvVXy1_0),.din(w_dff_A_eK7qKMgm7_0),.clk(gclk));
	jdff dff_A_ON5FvVXy1_0(.dout(w_dff_A_gRqDjITU4_0),.din(w_dff_A_ON5FvVXy1_0),.clk(gclk));
	jdff dff_A_gRqDjITU4_0(.dout(w_dff_A_9rkra2Mh0_0),.din(w_dff_A_gRqDjITU4_0),.clk(gclk));
	jdff dff_A_9rkra2Mh0_0(.dout(w_dff_A_hwZxyIz79_0),.din(w_dff_A_9rkra2Mh0_0),.clk(gclk));
	jdff dff_A_hwZxyIz79_0(.dout(w_dff_A_jE3CuK5s3_0),.din(w_dff_A_hwZxyIz79_0),.clk(gclk));
	jdff dff_A_jE3CuK5s3_0(.dout(w_dff_A_r74hzztW8_0),.din(w_dff_A_jE3CuK5s3_0),.clk(gclk));
	jdff dff_A_r74hzztW8_0(.dout(w_dff_A_6Kr9jzom6_0),.din(w_dff_A_r74hzztW8_0),.clk(gclk));
	jdff dff_A_6Kr9jzom6_0(.dout(w_dff_A_Z4OIoiN49_0),.din(w_dff_A_6Kr9jzom6_0),.clk(gclk));
	jdff dff_A_Z4OIoiN49_0(.dout(w_dff_A_6ntirba20_0),.din(w_dff_A_Z4OIoiN49_0),.clk(gclk));
	jdff dff_A_6ntirba20_0(.dout(w_dff_A_gAa2w9kM6_0),.din(w_dff_A_6ntirba20_0),.clk(gclk));
	jdff dff_A_gAa2w9kM6_0(.dout(w_dff_A_awoxwtPU7_0),.din(w_dff_A_gAa2w9kM6_0),.clk(gclk));
	jdff dff_A_awoxwtPU7_0(.dout(w_dff_A_GceHtWRX7_0),.din(w_dff_A_awoxwtPU7_0),.clk(gclk));
	jdff dff_A_GceHtWRX7_0(.dout(w_dff_A_q2X91lZv2_0),.din(w_dff_A_GceHtWRX7_0),.clk(gclk));
	jdff dff_A_q2X91lZv2_0(.dout(w_dff_A_9W89dofE4_0),.din(w_dff_A_q2X91lZv2_0),.clk(gclk));
	jdff dff_A_9W89dofE4_0(.dout(w_dff_A_SzKoG7Nf0_0),.din(w_dff_A_9W89dofE4_0),.clk(gclk));
	jdff dff_A_SzKoG7Nf0_0(.dout(w_dff_A_Vqyhnwny2_0),.din(w_dff_A_SzKoG7Nf0_0),.clk(gclk));
	jdff dff_A_Vqyhnwny2_0(.dout(w_dff_A_x5mplucE6_0),.din(w_dff_A_Vqyhnwny2_0),.clk(gclk));
	jdff dff_A_x5mplucE6_0(.dout(w_dff_A_t6Eg007H0_0),.din(w_dff_A_x5mplucE6_0),.clk(gclk));
	jdff dff_A_t6Eg007H0_0(.dout(w_dff_A_npW94Dfe7_0),.din(w_dff_A_t6Eg007H0_0),.clk(gclk));
	jdff dff_A_npW94Dfe7_0(.dout(w_dff_A_e8DteCl24_0),.din(w_dff_A_npW94Dfe7_0),.clk(gclk));
	jdff dff_A_e8DteCl24_0(.dout(w_dff_A_nXOA6hWi9_0),.din(w_dff_A_e8DteCl24_0),.clk(gclk));
	jdff dff_A_nXOA6hWi9_0(.dout(w_dff_A_t2C4BIya5_0),.din(w_dff_A_nXOA6hWi9_0),.clk(gclk));
	jdff dff_A_t2C4BIya5_0(.dout(w_dff_A_yd6bdb4p1_0),.din(w_dff_A_t2C4BIya5_0),.clk(gclk));
	jdff dff_A_yd6bdb4p1_0(.dout(w_dff_A_5XalOgPE1_0),.din(w_dff_A_yd6bdb4p1_0),.clk(gclk));
	jdff dff_A_5XalOgPE1_0(.dout(G436),.din(w_dff_A_5XalOgPE1_0),.clk(gclk));
	jdff dff_A_gDU3XBye5_1(.dout(w_dff_A_XaqKY3Uv8_0),.din(w_dff_A_gDU3XBye5_1),.clk(gclk));
	jdff dff_A_XaqKY3Uv8_0(.dout(w_dff_A_HT7RyJrq9_0),.din(w_dff_A_XaqKY3Uv8_0),.clk(gclk));
	jdff dff_A_HT7RyJrq9_0(.dout(w_dff_A_uKdcXXce1_0),.din(w_dff_A_HT7RyJrq9_0),.clk(gclk));
	jdff dff_A_uKdcXXce1_0(.dout(w_dff_A_S55DiAsQ2_0),.din(w_dff_A_uKdcXXce1_0),.clk(gclk));
	jdff dff_A_S55DiAsQ2_0(.dout(w_dff_A_14iiDsQQ6_0),.din(w_dff_A_S55DiAsQ2_0),.clk(gclk));
	jdff dff_A_14iiDsQQ6_0(.dout(w_dff_A_2ERLpZRJ8_0),.din(w_dff_A_14iiDsQQ6_0),.clk(gclk));
	jdff dff_A_2ERLpZRJ8_0(.dout(w_dff_A_ZOuhXUfD9_0),.din(w_dff_A_2ERLpZRJ8_0),.clk(gclk));
	jdff dff_A_ZOuhXUfD9_0(.dout(w_dff_A_VPTkTMMH5_0),.din(w_dff_A_ZOuhXUfD9_0),.clk(gclk));
	jdff dff_A_VPTkTMMH5_0(.dout(w_dff_A_bUiwIDly7_0),.din(w_dff_A_VPTkTMMH5_0),.clk(gclk));
	jdff dff_A_bUiwIDly7_0(.dout(w_dff_A_KLJ1kaQ70_0),.din(w_dff_A_bUiwIDly7_0),.clk(gclk));
	jdff dff_A_KLJ1kaQ70_0(.dout(w_dff_A_ycUmO0n55_0),.din(w_dff_A_KLJ1kaQ70_0),.clk(gclk));
	jdff dff_A_ycUmO0n55_0(.dout(w_dff_A_c5ukUARk7_0),.din(w_dff_A_ycUmO0n55_0),.clk(gclk));
	jdff dff_A_c5ukUARk7_0(.dout(w_dff_A_p1RpYnfq1_0),.din(w_dff_A_c5ukUARk7_0),.clk(gclk));
	jdff dff_A_p1RpYnfq1_0(.dout(w_dff_A_T0MSFy8n7_0),.din(w_dff_A_p1RpYnfq1_0),.clk(gclk));
	jdff dff_A_T0MSFy8n7_0(.dout(w_dff_A_5OZjwaVm4_0),.din(w_dff_A_T0MSFy8n7_0),.clk(gclk));
	jdff dff_A_5OZjwaVm4_0(.dout(w_dff_A_iQbagzNJ7_0),.din(w_dff_A_5OZjwaVm4_0),.clk(gclk));
	jdff dff_A_iQbagzNJ7_0(.dout(w_dff_A_Om19IT620_0),.din(w_dff_A_iQbagzNJ7_0),.clk(gclk));
	jdff dff_A_Om19IT620_0(.dout(w_dff_A_GqV94TZb7_0),.din(w_dff_A_Om19IT620_0),.clk(gclk));
	jdff dff_A_GqV94TZb7_0(.dout(w_dff_A_C8BBNJca9_0),.din(w_dff_A_GqV94TZb7_0),.clk(gclk));
	jdff dff_A_C8BBNJca9_0(.dout(w_dff_A_DQPdZpQ47_0),.din(w_dff_A_C8BBNJca9_0),.clk(gclk));
	jdff dff_A_DQPdZpQ47_0(.dout(w_dff_A_36kNi4lH9_0),.din(w_dff_A_DQPdZpQ47_0),.clk(gclk));
	jdff dff_A_36kNi4lH9_0(.dout(w_dff_A_nrs4xXtW1_0),.din(w_dff_A_36kNi4lH9_0),.clk(gclk));
	jdff dff_A_nrs4xXtW1_0(.dout(w_dff_A_RoCASpEY7_0),.din(w_dff_A_nrs4xXtW1_0),.clk(gclk));
	jdff dff_A_RoCASpEY7_0(.dout(w_dff_A_N94buLv33_0),.din(w_dff_A_RoCASpEY7_0),.clk(gclk));
	jdff dff_A_N94buLv33_0(.dout(w_dff_A_iHESPorf3_0),.din(w_dff_A_N94buLv33_0),.clk(gclk));
	jdff dff_A_iHESPorf3_0(.dout(w_dff_A_uwyn9o5o1_0),.din(w_dff_A_iHESPorf3_0),.clk(gclk));
	jdff dff_A_uwyn9o5o1_0(.dout(w_dff_A_BjG5g2wx7_0),.din(w_dff_A_uwyn9o5o1_0),.clk(gclk));
	jdff dff_A_BjG5g2wx7_0(.dout(w_dff_A_0UFCBU9A4_0),.din(w_dff_A_BjG5g2wx7_0),.clk(gclk));
	jdff dff_A_0UFCBU9A4_0(.dout(w_dff_A_dIPEFoYA6_0),.din(w_dff_A_0UFCBU9A4_0),.clk(gclk));
	jdff dff_A_dIPEFoYA6_0(.dout(w_dff_A_In1Y5C103_0),.din(w_dff_A_dIPEFoYA6_0),.clk(gclk));
	jdff dff_A_In1Y5C103_0(.dout(w_dff_A_sl6JrQzi9_0),.din(w_dff_A_In1Y5C103_0),.clk(gclk));
	jdff dff_A_sl6JrQzi9_0(.dout(w_dff_A_RKaIDixn2_0),.din(w_dff_A_sl6JrQzi9_0),.clk(gclk));
	jdff dff_A_RKaIDixn2_0(.dout(w_dff_A_oi7ybY5V9_0),.din(w_dff_A_RKaIDixn2_0),.clk(gclk));
	jdff dff_A_oi7ybY5V9_0(.dout(w_dff_A_Stah2Cq73_0),.din(w_dff_A_oi7ybY5V9_0),.clk(gclk));
	jdff dff_A_Stah2Cq73_0(.dout(w_dff_A_1oAPG64a6_0),.din(w_dff_A_Stah2Cq73_0),.clk(gclk));
	jdff dff_A_1oAPG64a6_0(.dout(w_dff_A_GGRN8gwU6_0),.din(w_dff_A_1oAPG64a6_0),.clk(gclk));
	jdff dff_A_GGRN8gwU6_0(.dout(w_dff_A_ocRhdTu39_0),.din(w_dff_A_GGRN8gwU6_0),.clk(gclk));
	jdff dff_A_ocRhdTu39_0(.dout(w_dff_A_j5NQvppo7_0),.din(w_dff_A_ocRhdTu39_0),.clk(gclk));
	jdff dff_A_j5NQvppo7_0(.dout(G478),.din(w_dff_A_j5NQvppo7_0),.clk(gclk));
	jdff dff_A_A1UvnyQh2_1(.dout(w_dff_A_juuvXi4i5_0),.din(w_dff_A_A1UvnyQh2_1),.clk(gclk));
	jdff dff_A_juuvXi4i5_0(.dout(w_dff_A_r73q4xdv6_0),.din(w_dff_A_juuvXi4i5_0),.clk(gclk));
	jdff dff_A_r73q4xdv6_0(.dout(w_dff_A_aAZO6Nog0_0),.din(w_dff_A_r73q4xdv6_0),.clk(gclk));
	jdff dff_A_aAZO6Nog0_0(.dout(w_dff_A_ER8IkTw92_0),.din(w_dff_A_aAZO6Nog0_0),.clk(gclk));
	jdff dff_A_ER8IkTw92_0(.dout(w_dff_A_o4IQMRov5_0),.din(w_dff_A_ER8IkTw92_0),.clk(gclk));
	jdff dff_A_o4IQMRov5_0(.dout(w_dff_A_r3uHDbat4_0),.din(w_dff_A_o4IQMRov5_0),.clk(gclk));
	jdff dff_A_r3uHDbat4_0(.dout(w_dff_A_kRzEGgJu7_0),.din(w_dff_A_r3uHDbat4_0),.clk(gclk));
	jdff dff_A_kRzEGgJu7_0(.dout(w_dff_A_qf4wB7cb9_0),.din(w_dff_A_kRzEGgJu7_0),.clk(gclk));
	jdff dff_A_qf4wB7cb9_0(.dout(w_dff_A_Y8vkjRUW5_0),.din(w_dff_A_qf4wB7cb9_0),.clk(gclk));
	jdff dff_A_Y8vkjRUW5_0(.dout(w_dff_A_cXCYdfaI5_0),.din(w_dff_A_Y8vkjRUW5_0),.clk(gclk));
	jdff dff_A_cXCYdfaI5_0(.dout(w_dff_A_i97WNmP72_0),.din(w_dff_A_cXCYdfaI5_0),.clk(gclk));
	jdff dff_A_i97WNmP72_0(.dout(w_dff_A_NC1IORo18_0),.din(w_dff_A_i97WNmP72_0),.clk(gclk));
	jdff dff_A_NC1IORo18_0(.dout(w_dff_A_8K3toON05_0),.din(w_dff_A_NC1IORo18_0),.clk(gclk));
	jdff dff_A_8K3toON05_0(.dout(w_dff_A_VlbAE4hi5_0),.din(w_dff_A_8K3toON05_0),.clk(gclk));
	jdff dff_A_VlbAE4hi5_0(.dout(w_dff_A_1ZcrHtIr3_0),.din(w_dff_A_VlbAE4hi5_0),.clk(gclk));
	jdff dff_A_1ZcrHtIr3_0(.dout(w_dff_A_1C1ZgeCE3_0),.din(w_dff_A_1ZcrHtIr3_0),.clk(gclk));
	jdff dff_A_1C1ZgeCE3_0(.dout(w_dff_A_cPO6wbOn0_0),.din(w_dff_A_1C1ZgeCE3_0),.clk(gclk));
	jdff dff_A_cPO6wbOn0_0(.dout(w_dff_A_wQdq0cQ51_0),.din(w_dff_A_cPO6wbOn0_0),.clk(gclk));
	jdff dff_A_wQdq0cQ51_0(.dout(w_dff_A_HecgiphY4_0),.din(w_dff_A_wQdq0cQ51_0),.clk(gclk));
	jdff dff_A_HecgiphY4_0(.dout(w_dff_A_F0iMQwZu7_0),.din(w_dff_A_HecgiphY4_0),.clk(gclk));
	jdff dff_A_F0iMQwZu7_0(.dout(w_dff_A_QKYiXZuG4_0),.din(w_dff_A_F0iMQwZu7_0),.clk(gclk));
	jdff dff_A_QKYiXZuG4_0(.dout(w_dff_A_kbNUKgLM4_0),.din(w_dff_A_QKYiXZuG4_0),.clk(gclk));
	jdff dff_A_kbNUKgLM4_0(.dout(w_dff_A_jQFjtW4i1_0),.din(w_dff_A_kbNUKgLM4_0),.clk(gclk));
	jdff dff_A_jQFjtW4i1_0(.dout(w_dff_A_tvsClI7Q6_0),.din(w_dff_A_jQFjtW4i1_0),.clk(gclk));
	jdff dff_A_tvsClI7Q6_0(.dout(w_dff_A_wG3InMlT3_0),.din(w_dff_A_tvsClI7Q6_0),.clk(gclk));
	jdff dff_A_wG3InMlT3_0(.dout(w_dff_A_8jX9fUtF4_0),.din(w_dff_A_wG3InMlT3_0),.clk(gclk));
	jdff dff_A_8jX9fUtF4_0(.dout(w_dff_A_tgINGoiR5_0),.din(w_dff_A_8jX9fUtF4_0),.clk(gclk));
	jdff dff_A_tgINGoiR5_0(.dout(w_dff_A_aglNXVMK6_0),.din(w_dff_A_tgINGoiR5_0),.clk(gclk));
	jdff dff_A_aglNXVMK6_0(.dout(w_dff_A_YqUCq5HW9_0),.din(w_dff_A_aglNXVMK6_0),.clk(gclk));
	jdff dff_A_YqUCq5HW9_0(.dout(w_dff_A_asljbY750_0),.din(w_dff_A_YqUCq5HW9_0),.clk(gclk));
	jdff dff_A_asljbY750_0(.dout(w_dff_A_m4NMEdVN7_0),.din(w_dff_A_asljbY750_0),.clk(gclk));
	jdff dff_A_m4NMEdVN7_0(.dout(w_dff_A_rQfQiJ3b0_0),.din(w_dff_A_m4NMEdVN7_0),.clk(gclk));
	jdff dff_A_rQfQiJ3b0_0(.dout(w_dff_A_oxLrrY4h2_0),.din(w_dff_A_rQfQiJ3b0_0),.clk(gclk));
	jdff dff_A_oxLrrY4h2_0(.dout(w_dff_A_2fnleoYj8_0),.din(w_dff_A_oxLrrY4h2_0),.clk(gclk));
	jdff dff_A_2fnleoYj8_0(.dout(w_dff_A_QKaa79P86_0),.din(w_dff_A_2fnleoYj8_0),.clk(gclk));
	jdff dff_A_QKaa79P86_0(.dout(w_dff_A_y6VYdPWv5_0),.din(w_dff_A_QKaa79P86_0),.clk(gclk));
	jdff dff_A_y6VYdPWv5_0(.dout(w_dff_A_F6Zd8z8H0_0),.din(w_dff_A_y6VYdPWv5_0),.clk(gclk));
	jdff dff_A_F6Zd8z8H0_0(.dout(w_dff_A_7xpMx7Hg3_0),.din(w_dff_A_F6Zd8z8H0_0),.clk(gclk));
	jdff dff_A_7xpMx7Hg3_0(.dout(G522),.din(w_dff_A_7xpMx7Hg3_0),.clk(gclk));
	jdff dff_A_ytKocOgQ9_2(.dout(w_dff_A_u5xFHdfj4_0),.din(w_dff_A_ytKocOgQ9_2),.clk(gclk));
	jdff dff_A_u5xFHdfj4_0(.dout(w_dff_A_WjhAFeTN3_0),.din(w_dff_A_u5xFHdfj4_0),.clk(gclk));
	jdff dff_A_WjhAFeTN3_0(.dout(w_dff_A_i0Qe0xZI2_0),.din(w_dff_A_WjhAFeTN3_0),.clk(gclk));
	jdff dff_A_i0Qe0xZI2_0(.dout(w_dff_A_uu0dqjlh6_0),.din(w_dff_A_i0Qe0xZI2_0),.clk(gclk));
	jdff dff_A_uu0dqjlh6_0(.dout(w_dff_A_MUSNqhkS9_0),.din(w_dff_A_uu0dqjlh6_0),.clk(gclk));
	jdff dff_A_MUSNqhkS9_0(.dout(w_dff_A_CdTwKHOO1_0),.din(w_dff_A_MUSNqhkS9_0),.clk(gclk));
	jdff dff_A_CdTwKHOO1_0(.dout(w_dff_A_zDHfvWjw4_0),.din(w_dff_A_CdTwKHOO1_0),.clk(gclk));
	jdff dff_A_zDHfvWjw4_0(.dout(w_dff_A_REomNbKK3_0),.din(w_dff_A_zDHfvWjw4_0),.clk(gclk));
	jdff dff_A_REomNbKK3_0(.dout(w_dff_A_1PiOxjdb9_0),.din(w_dff_A_REomNbKK3_0),.clk(gclk));
	jdff dff_A_1PiOxjdb9_0(.dout(w_dff_A_lVT4Lv2J2_0),.din(w_dff_A_1PiOxjdb9_0),.clk(gclk));
	jdff dff_A_lVT4Lv2J2_0(.dout(w_dff_A_17kDSziH4_0),.din(w_dff_A_lVT4Lv2J2_0),.clk(gclk));
	jdff dff_A_17kDSziH4_0(.dout(w_dff_A_PseaJE7S1_0),.din(w_dff_A_17kDSziH4_0),.clk(gclk));
	jdff dff_A_PseaJE7S1_0(.dout(w_dff_A_kt8TGQsx6_0),.din(w_dff_A_PseaJE7S1_0),.clk(gclk));
	jdff dff_A_kt8TGQsx6_0(.dout(w_dff_A_9VH95EMP3_0),.din(w_dff_A_kt8TGQsx6_0),.clk(gclk));
	jdff dff_A_9VH95EMP3_0(.dout(w_dff_A_m7SZCh5R7_0),.din(w_dff_A_9VH95EMP3_0),.clk(gclk));
	jdff dff_A_m7SZCh5R7_0(.dout(w_dff_A_HLy6FROn2_0),.din(w_dff_A_m7SZCh5R7_0),.clk(gclk));
	jdff dff_A_HLy6FROn2_0(.dout(w_dff_A_vVOcTRRB1_0),.din(w_dff_A_HLy6FROn2_0),.clk(gclk));
	jdff dff_A_vVOcTRRB1_0(.dout(w_dff_A_qxxy23fn0_0),.din(w_dff_A_vVOcTRRB1_0),.clk(gclk));
	jdff dff_A_qxxy23fn0_0(.dout(w_dff_A_LUMijow94_0),.din(w_dff_A_qxxy23fn0_0),.clk(gclk));
	jdff dff_A_LUMijow94_0(.dout(w_dff_A_QcqMtWdv5_0),.din(w_dff_A_LUMijow94_0),.clk(gclk));
	jdff dff_A_QcqMtWdv5_0(.dout(w_dff_A_BU6FsyXU0_0),.din(w_dff_A_QcqMtWdv5_0),.clk(gclk));
	jdff dff_A_BU6FsyXU0_0(.dout(w_dff_A_iYOqQ03s6_0),.din(w_dff_A_BU6FsyXU0_0),.clk(gclk));
	jdff dff_A_iYOqQ03s6_0(.dout(w_dff_A_F17JKdJi0_0),.din(w_dff_A_iYOqQ03s6_0),.clk(gclk));
	jdff dff_A_F17JKdJi0_0(.dout(w_dff_A_zcTBT6Mo7_0),.din(w_dff_A_F17JKdJi0_0),.clk(gclk));
	jdff dff_A_zcTBT6Mo7_0(.dout(w_dff_A_aCEpFAws8_0),.din(w_dff_A_zcTBT6Mo7_0),.clk(gclk));
	jdff dff_A_aCEpFAws8_0(.dout(w_dff_A_hYJjWxaU4_0),.din(w_dff_A_aCEpFAws8_0),.clk(gclk));
	jdff dff_A_hYJjWxaU4_0(.dout(w_dff_A_edeUIN8j2_0),.din(w_dff_A_hYJjWxaU4_0),.clk(gclk));
	jdff dff_A_edeUIN8j2_0(.dout(w_dff_A_oRNrh9pK4_0),.din(w_dff_A_edeUIN8j2_0),.clk(gclk));
	jdff dff_A_oRNrh9pK4_0(.dout(w_dff_A_ADmdLgf23_0),.din(w_dff_A_oRNrh9pK4_0),.clk(gclk));
	jdff dff_A_ADmdLgf23_0(.dout(w_dff_A_SmSVMTgY7_0),.din(w_dff_A_ADmdLgf23_0),.clk(gclk));
	jdff dff_A_SmSVMTgY7_0(.dout(w_dff_A_sgXfAoIJ8_0),.din(w_dff_A_SmSVMTgY7_0),.clk(gclk));
	jdff dff_A_sgXfAoIJ8_0(.dout(w_dff_A_IfOjwXXJ5_0),.din(w_dff_A_sgXfAoIJ8_0),.clk(gclk));
	jdff dff_A_IfOjwXXJ5_0(.dout(w_dff_A_MZSXz5CL7_0),.din(w_dff_A_IfOjwXXJ5_0),.clk(gclk));
	jdff dff_A_MZSXz5CL7_0(.dout(w_dff_A_nwL4j4is7_0),.din(w_dff_A_MZSXz5CL7_0),.clk(gclk));
	jdff dff_A_nwL4j4is7_0(.dout(w_dff_A_NOAIjAV92_0),.din(w_dff_A_nwL4j4is7_0),.clk(gclk));
	jdff dff_A_NOAIjAV92_0(.dout(w_dff_A_i8ISFjqi3_0),.din(w_dff_A_NOAIjAV92_0),.clk(gclk));
	jdff dff_A_i8ISFjqi3_0(.dout(w_dff_A_lap6QBdo1_0),.din(w_dff_A_i8ISFjqi3_0),.clk(gclk));
	jdff dff_A_lap6QBdo1_0(.dout(G402),.din(w_dff_A_lap6QBdo1_0),.clk(gclk));
	jdff dff_A_J1N7OnNX3_1(.dout(w_dff_A_cZlyu6Op5_0),.din(w_dff_A_J1N7OnNX3_1),.clk(gclk));
	jdff dff_A_cZlyu6Op5_0(.dout(w_dff_A_2iWyQBWE1_0),.din(w_dff_A_cZlyu6Op5_0),.clk(gclk));
	jdff dff_A_2iWyQBWE1_0(.dout(w_dff_A_WQuOi4cU9_0),.din(w_dff_A_2iWyQBWE1_0),.clk(gclk));
	jdff dff_A_WQuOi4cU9_0(.dout(w_dff_A_GYvyVxEJ1_0),.din(w_dff_A_WQuOi4cU9_0),.clk(gclk));
	jdff dff_A_GYvyVxEJ1_0(.dout(w_dff_A_z4eYSgZB9_0),.din(w_dff_A_GYvyVxEJ1_0),.clk(gclk));
	jdff dff_A_z4eYSgZB9_0(.dout(w_dff_A_G22fjfJg1_0),.din(w_dff_A_z4eYSgZB9_0),.clk(gclk));
	jdff dff_A_G22fjfJg1_0(.dout(w_dff_A_0BtYIAYk7_0),.din(w_dff_A_G22fjfJg1_0),.clk(gclk));
	jdff dff_A_0BtYIAYk7_0(.dout(w_dff_A_c0Qgxy8h0_0),.din(w_dff_A_0BtYIAYk7_0),.clk(gclk));
	jdff dff_A_c0Qgxy8h0_0(.dout(w_dff_A_ZlbS6m6V5_0),.din(w_dff_A_c0Qgxy8h0_0),.clk(gclk));
	jdff dff_A_ZlbS6m6V5_0(.dout(w_dff_A_3fKf1FqW7_0),.din(w_dff_A_ZlbS6m6V5_0),.clk(gclk));
	jdff dff_A_3fKf1FqW7_0(.dout(w_dff_A_m6vayyXN6_0),.din(w_dff_A_3fKf1FqW7_0),.clk(gclk));
	jdff dff_A_m6vayyXN6_0(.dout(w_dff_A_zHOyvh6I5_0),.din(w_dff_A_m6vayyXN6_0),.clk(gclk));
	jdff dff_A_zHOyvh6I5_0(.dout(w_dff_A_3xsB2VpR0_0),.din(w_dff_A_zHOyvh6I5_0),.clk(gclk));
	jdff dff_A_3xsB2VpR0_0(.dout(w_dff_A_F6GOwVeM8_0),.din(w_dff_A_3xsB2VpR0_0),.clk(gclk));
	jdff dff_A_F6GOwVeM8_0(.dout(w_dff_A_qFyn40Y37_0),.din(w_dff_A_F6GOwVeM8_0),.clk(gclk));
	jdff dff_A_qFyn40Y37_0(.dout(w_dff_A_KheC66zi1_0),.din(w_dff_A_qFyn40Y37_0),.clk(gclk));
	jdff dff_A_KheC66zi1_0(.dout(w_dff_A_FThAYanL2_0),.din(w_dff_A_KheC66zi1_0),.clk(gclk));
	jdff dff_A_FThAYanL2_0(.dout(w_dff_A_FxhLIXlx9_0),.din(w_dff_A_FThAYanL2_0),.clk(gclk));
	jdff dff_A_FxhLIXlx9_0(.dout(w_dff_A_kMh4pZ8s4_0),.din(w_dff_A_FxhLIXlx9_0),.clk(gclk));
	jdff dff_A_kMh4pZ8s4_0(.dout(w_dff_A_xER7NfyN8_0),.din(w_dff_A_kMh4pZ8s4_0),.clk(gclk));
	jdff dff_A_xER7NfyN8_0(.dout(w_dff_A_6CAWJEE01_0),.din(w_dff_A_xER7NfyN8_0),.clk(gclk));
	jdff dff_A_6CAWJEE01_0(.dout(w_dff_A_1TxotZe58_0),.din(w_dff_A_6CAWJEE01_0),.clk(gclk));
	jdff dff_A_1TxotZe58_0(.dout(w_dff_A_0vSiCIxz0_0),.din(w_dff_A_1TxotZe58_0),.clk(gclk));
	jdff dff_A_0vSiCIxz0_0(.dout(w_dff_A_ONIgy8xa7_0),.din(w_dff_A_0vSiCIxz0_0),.clk(gclk));
	jdff dff_A_ONIgy8xa7_0(.dout(w_dff_A_sAWWlxPQ1_0),.din(w_dff_A_ONIgy8xa7_0),.clk(gclk));
	jdff dff_A_sAWWlxPQ1_0(.dout(w_dff_A_K6eae1RU0_0),.din(w_dff_A_sAWWlxPQ1_0),.clk(gclk));
	jdff dff_A_K6eae1RU0_0(.dout(w_dff_A_39OMQxVR5_0),.din(w_dff_A_K6eae1RU0_0),.clk(gclk));
	jdff dff_A_39OMQxVR5_0(.dout(w_dff_A_ryC3YZ0i3_0),.din(w_dff_A_39OMQxVR5_0),.clk(gclk));
	jdff dff_A_ryC3YZ0i3_0(.dout(w_dff_A_RcZpSoEr1_0),.din(w_dff_A_ryC3YZ0i3_0),.clk(gclk));
	jdff dff_A_RcZpSoEr1_0(.dout(w_dff_A_Qj9Fo3y39_0),.din(w_dff_A_RcZpSoEr1_0),.clk(gclk));
	jdff dff_A_Qj9Fo3y39_0(.dout(w_dff_A_I02JL7wp8_0),.din(w_dff_A_Qj9Fo3y39_0),.clk(gclk));
	jdff dff_A_I02JL7wp8_0(.dout(w_dff_A_XnvXlk3W7_0),.din(w_dff_A_I02JL7wp8_0),.clk(gclk));
	jdff dff_A_XnvXlk3W7_0(.dout(w_dff_A_SBLRncLt0_0),.din(w_dff_A_XnvXlk3W7_0),.clk(gclk));
	jdff dff_A_SBLRncLt0_0(.dout(w_dff_A_kGAyADmM3_0),.din(w_dff_A_SBLRncLt0_0),.clk(gclk));
	jdff dff_A_kGAyADmM3_0(.dout(w_dff_A_4JNmywKz3_0),.din(w_dff_A_kGAyADmM3_0),.clk(gclk));
	jdff dff_A_4JNmywKz3_0(.dout(G404),.din(w_dff_A_4JNmywKz3_0),.clk(gclk));
	jdff dff_A_vKZYkuMo0_1(.dout(w_dff_A_y1wWVzf25_0),.din(w_dff_A_vKZYkuMo0_1),.clk(gclk));
	jdff dff_A_y1wWVzf25_0(.dout(w_dff_A_xJ6PQyQB2_0),.din(w_dff_A_y1wWVzf25_0),.clk(gclk));
	jdff dff_A_xJ6PQyQB2_0(.dout(w_dff_A_9fONwAQG3_0),.din(w_dff_A_xJ6PQyQB2_0),.clk(gclk));
	jdff dff_A_9fONwAQG3_0(.dout(w_dff_A_NVCuZiQI8_0),.din(w_dff_A_9fONwAQG3_0),.clk(gclk));
	jdff dff_A_NVCuZiQI8_0(.dout(w_dff_A_k0TrAN6J8_0),.din(w_dff_A_NVCuZiQI8_0),.clk(gclk));
	jdff dff_A_k0TrAN6J8_0(.dout(w_dff_A_BNaTlAM82_0),.din(w_dff_A_k0TrAN6J8_0),.clk(gclk));
	jdff dff_A_BNaTlAM82_0(.dout(w_dff_A_L0AVxZpo7_0),.din(w_dff_A_BNaTlAM82_0),.clk(gclk));
	jdff dff_A_L0AVxZpo7_0(.dout(w_dff_A_iqtFYjiF8_0),.din(w_dff_A_L0AVxZpo7_0),.clk(gclk));
	jdff dff_A_iqtFYjiF8_0(.dout(w_dff_A_gnHKDHsb3_0),.din(w_dff_A_iqtFYjiF8_0),.clk(gclk));
	jdff dff_A_gnHKDHsb3_0(.dout(w_dff_A_IjITfvdX3_0),.din(w_dff_A_gnHKDHsb3_0),.clk(gclk));
	jdff dff_A_IjITfvdX3_0(.dout(w_dff_A_9zsa2Fmy4_0),.din(w_dff_A_IjITfvdX3_0),.clk(gclk));
	jdff dff_A_9zsa2Fmy4_0(.dout(w_dff_A_qLyNy7Xk7_0),.din(w_dff_A_9zsa2Fmy4_0),.clk(gclk));
	jdff dff_A_qLyNy7Xk7_0(.dout(w_dff_A_ADjBySD68_0),.din(w_dff_A_qLyNy7Xk7_0),.clk(gclk));
	jdff dff_A_ADjBySD68_0(.dout(w_dff_A_P0c72Ign7_0),.din(w_dff_A_ADjBySD68_0),.clk(gclk));
	jdff dff_A_P0c72Ign7_0(.dout(w_dff_A_y0rhxQyx4_0),.din(w_dff_A_P0c72Ign7_0),.clk(gclk));
	jdff dff_A_y0rhxQyx4_0(.dout(w_dff_A_N1tgLf6D6_0),.din(w_dff_A_y0rhxQyx4_0),.clk(gclk));
	jdff dff_A_N1tgLf6D6_0(.dout(w_dff_A_D96EK0Sb7_0),.din(w_dff_A_N1tgLf6D6_0),.clk(gclk));
	jdff dff_A_D96EK0Sb7_0(.dout(w_dff_A_Jm0BlKwW1_0),.din(w_dff_A_D96EK0Sb7_0),.clk(gclk));
	jdff dff_A_Jm0BlKwW1_0(.dout(w_dff_A_p335ytl93_0),.din(w_dff_A_Jm0BlKwW1_0),.clk(gclk));
	jdff dff_A_p335ytl93_0(.dout(w_dff_A_sOloWGCk6_0),.din(w_dff_A_p335ytl93_0),.clk(gclk));
	jdff dff_A_sOloWGCk6_0(.dout(w_dff_A_mIMorqH67_0),.din(w_dff_A_sOloWGCk6_0),.clk(gclk));
	jdff dff_A_mIMorqH67_0(.dout(w_dff_A_HS6lVqRg9_0),.din(w_dff_A_mIMorqH67_0),.clk(gclk));
	jdff dff_A_HS6lVqRg9_0(.dout(w_dff_A_BHAdBjoz8_0),.din(w_dff_A_HS6lVqRg9_0),.clk(gclk));
	jdff dff_A_BHAdBjoz8_0(.dout(w_dff_A_w7EP3kX83_0),.din(w_dff_A_BHAdBjoz8_0),.clk(gclk));
	jdff dff_A_w7EP3kX83_0(.dout(w_dff_A_efElcyDT8_0),.din(w_dff_A_w7EP3kX83_0),.clk(gclk));
	jdff dff_A_efElcyDT8_0(.dout(w_dff_A_nBnFMORK2_0),.din(w_dff_A_efElcyDT8_0),.clk(gclk));
	jdff dff_A_nBnFMORK2_0(.dout(w_dff_A_vAcffl565_0),.din(w_dff_A_nBnFMORK2_0),.clk(gclk));
	jdff dff_A_vAcffl565_0(.dout(w_dff_A_MnEcJrgw4_0),.din(w_dff_A_vAcffl565_0),.clk(gclk));
	jdff dff_A_MnEcJrgw4_0(.dout(w_dff_A_iRZ7G1i57_0),.din(w_dff_A_MnEcJrgw4_0),.clk(gclk));
	jdff dff_A_iRZ7G1i57_0(.dout(w_dff_A_9JtKrjYg0_0),.din(w_dff_A_iRZ7G1i57_0),.clk(gclk));
	jdff dff_A_9JtKrjYg0_0(.dout(w_dff_A_4VhiGOsD6_0),.din(w_dff_A_9JtKrjYg0_0),.clk(gclk));
	jdff dff_A_4VhiGOsD6_0(.dout(w_dff_A_RkOevjGX8_0),.din(w_dff_A_4VhiGOsD6_0),.clk(gclk));
	jdff dff_A_RkOevjGX8_0(.dout(w_dff_A_bX2iq0xp7_0),.din(w_dff_A_RkOevjGX8_0),.clk(gclk));
	jdff dff_A_bX2iq0xp7_0(.dout(w_dff_A_Mm3jRJD58_0),.din(w_dff_A_bX2iq0xp7_0),.clk(gclk));
	jdff dff_A_Mm3jRJD58_0(.dout(w_dff_A_UO7Ui96n4_0),.din(w_dff_A_Mm3jRJD58_0),.clk(gclk));
	jdff dff_A_UO7Ui96n4_0(.dout(G406),.din(w_dff_A_UO7Ui96n4_0),.clk(gclk));
	jdff dff_A_pWywJuT40_1(.dout(w_dff_A_OmcSt8XA9_0),.din(w_dff_A_pWywJuT40_1),.clk(gclk));
	jdff dff_A_OmcSt8XA9_0(.dout(w_dff_A_G3whShqi9_0),.din(w_dff_A_OmcSt8XA9_0),.clk(gclk));
	jdff dff_A_G3whShqi9_0(.dout(w_dff_A_CZWnj7yt0_0),.din(w_dff_A_G3whShqi9_0),.clk(gclk));
	jdff dff_A_CZWnj7yt0_0(.dout(w_dff_A_WKcQ9D6q1_0),.din(w_dff_A_CZWnj7yt0_0),.clk(gclk));
	jdff dff_A_WKcQ9D6q1_0(.dout(w_dff_A_SuqlomHn0_0),.din(w_dff_A_WKcQ9D6q1_0),.clk(gclk));
	jdff dff_A_SuqlomHn0_0(.dout(w_dff_A_52SSafLD6_0),.din(w_dff_A_SuqlomHn0_0),.clk(gclk));
	jdff dff_A_52SSafLD6_0(.dout(w_dff_A_rhyFH44k0_0),.din(w_dff_A_52SSafLD6_0),.clk(gclk));
	jdff dff_A_rhyFH44k0_0(.dout(w_dff_A_Jvz11xS98_0),.din(w_dff_A_rhyFH44k0_0),.clk(gclk));
	jdff dff_A_Jvz11xS98_0(.dout(w_dff_A_ohBE1dOx0_0),.din(w_dff_A_Jvz11xS98_0),.clk(gclk));
	jdff dff_A_ohBE1dOx0_0(.dout(w_dff_A_YcrqZh111_0),.din(w_dff_A_ohBE1dOx0_0),.clk(gclk));
	jdff dff_A_YcrqZh111_0(.dout(w_dff_A_z2qtqzGQ5_0),.din(w_dff_A_YcrqZh111_0),.clk(gclk));
	jdff dff_A_z2qtqzGQ5_0(.dout(w_dff_A_BYl4qxk40_0),.din(w_dff_A_z2qtqzGQ5_0),.clk(gclk));
	jdff dff_A_BYl4qxk40_0(.dout(w_dff_A_pNKDWu4z1_0),.din(w_dff_A_BYl4qxk40_0),.clk(gclk));
	jdff dff_A_pNKDWu4z1_0(.dout(w_dff_A_J3a95Kom8_0),.din(w_dff_A_pNKDWu4z1_0),.clk(gclk));
	jdff dff_A_J3a95Kom8_0(.dout(w_dff_A_EsWQiaez5_0),.din(w_dff_A_J3a95Kom8_0),.clk(gclk));
	jdff dff_A_EsWQiaez5_0(.dout(w_dff_A_fGLI1hom9_0),.din(w_dff_A_EsWQiaez5_0),.clk(gclk));
	jdff dff_A_fGLI1hom9_0(.dout(w_dff_A_lqZ1YNqm0_0),.din(w_dff_A_fGLI1hom9_0),.clk(gclk));
	jdff dff_A_lqZ1YNqm0_0(.dout(w_dff_A_aES1XdRl7_0),.din(w_dff_A_lqZ1YNqm0_0),.clk(gclk));
	jdff dff_A_aES1XdRl7_0(.dout(w_dff_A_XezniCnN2_0),.din(w_dff_A_aES1XdRl7_0),.clk(gclk));
	jdff dff_A_XezniCnN2_0(.dout(w_dff_A_G1qFyNAM7_0),.din(w_dff_A_XezniCnN2_0),.clk(gclk));
	jdff dff_A_G1qFyNAM7_0(.dout(w_dff_A_77v2BGaR4_0),.din(w_dff_A_G1qFyNAM7_0),.clk(gclk));
	jdff dff_A_77v2BGaR4_0(.dout(w_dff_A_imZMvE2Z6_0),.din(w_dff_A_77v2BGaR4_0),.clk(gclk));
	jdff dff_A_imZMvE2Z6_0(.dout(w_dff_A_90aUtIOG5_0),.din(w_dff_A_imZMvE2Z6_0),.clk(gclk));
	jdff dff_A_90aUtIOG5_0(.dout(w_dff_A_0v7KErAQ1_0),.din(w_dff_A_90aUtIOG5_0),.clk(gclk));
	jdff dff_A_0v7KErAQ1_0(.dout(w_dff_A_nx3FjhIU3_0),.din(w_dff_A_0v7KErAQ1_0),.clk(gclk));
	jdff dff_A_nx3FjhIU3_0(.dout(w_dff_A_s9cDMHhc8_0),.din(w_dff_A_nx3FjhIU3_0),.clk(gclk));
	jdff dff_A_s9cDMHhc8_0(.dout(w_dff_A_hE3LesJc5_0),.din(w_dff_A_s9cDMHhc8_0),.clk(gclk));
	jdff dff_A_hE3LesJc5_0(.dout(w_dff_A_VqfrfqeV1_0),.din(w_dff_A_hE3LesJc5_0),.clk(gclk));
	jdff dff_A_VqfrfqeV1_0(.dout(w_dff_A_L7xPMk6m2_0),.din(w_dff_A_VqfrfqeV1_0),.clk(gclk));
	jdff dff_A_L7xPMk6m2_0(.dout(w_dff_A_oxMLrf1v5_0),.din(w_dff_A_L7xPMk6m2_0),.clk(gclk));
	jdff dff_A_oxMLrf1v5_0(.dout(w_dff_A_BNGkmhFq8_0),.din(w_dff_A_oxMLrf1v5_0),.clk(gclk));
	jdff dff_A_BNGkmhFq8_0(.dout(w_dff_A_LIqfwZBR1_0),.din(w_dff_A_BNGkmhFq8_0),.clk(gclk));
	jdff dff_A_LIqfwZBR1_0(.dout(w_dff_A_4Vgnq3KN2_0),.din(w_dff_A_LIqfwZBR1_0),.clk(gclk));
	jdff dff_A_4Vgnq3KN2_0(.dout(w_dff_A_B2VwcZ5K1_0),.din(w_dff_A_4Vgnq3KN2_0),.clk(gclk));
	jdff dff_A_B2VwcZ5K1_0(.dout(w_dff_A_tswiLVgG9_0),.din(w_dff_A_B2VwcZ5K1_0),.clk(gclk));
	jdff dff_A_tswiLVgG9_0(.dout(G408),.din(w_dff_A_tswiLVgG9_0),.clk(gclk));
	jdff dff_A_4rlRYtVI6_1(.dout(w_dff_A_lVJCs9ZF4_0),.din(w_dff_A_4rlRYtVI6_1),.clk(gclk));
	jdff dff_A_lVJCs9ZF4_0(.dout(w_dff_A_BzvzbFi90_0),.din(w_dff_A_lVJCs9ZF4_0),.clk(gclk));
	jdff dff_A_BzvzbFi90_0(.dout(w_dff_A_8ApUZZPu5_0),.din(w_dff_A_BzvzbFi90_0),.clk(gclk));
	jdff dff_A_8ApUZZPu5_0(.dout(w_dff_A_5p3tVPcr1_0),.din(w_dff_A_8ApUZZPu5_0),.clk(gclk));
	jdff dff_A_5p3tVPcr1_0(.dout(w_dff_A_9nnseZvV1_0),.din(w_dff_A_5p3tVPcr1_0),.clk(gclk));
	jdff dff_A_9nnseZvV1_0(.dout(w_dff_A_J3LHzdNO5_0),.din(w_dff_A_9nnseZvV1_0),.clk(gclk));
	jdff dff_A_J3LHzdNO5_0(.dout(w_dff_A_xUbCm4fK5_0),.din(w_dff_A_J3LHzdNO5_0),.clk(gclk));
	jdff dff_A_xUbCm4fK5_0(.dout(w_dff_A_FGV63dXO2_0),.din(w_dff_A_xUbCm4fK5_0),.clk(gclk));
	jdff dff_A_FGV63dXO2_0(.dout(w_dff_A_3dJgQMh64_0),.din(w_dff_A_FGV63dXO2_0),.clk(gclk));
	jdff dff_A_3dJgQMh64_0(.dout(w_dff_A_V0NOh91S7_0),.din(w_dff_A_3dJgQMh64_0),.clk(gclk));
	jdff dff_A_V0NOh91S7_0(.dout(w_dff_A_9ujKsLdH3_0),.din(w_dff_A_V0NOh91S7_0),.clk(gclk));
	jdff dff_A_9ujKsLdH3_0(.dout(w_dff_A_czrNmvtQ8_0),.din(w_dff_A_9ujKsLdH3_0),.clk(gclk));
	jdff dff_A_czrNmvtQ8_0(.dout(w_dff_A_kYBm0jpd5_0),.din(w_dff_A_czrNmvtQ8_0),.clk(gclk));
	jdff dff_A_kYBm0jpd5_0(.dout(w_dff_A_NNGpHLtA3_0),.din(w_dff_A_kYBm0jpd5_0),.clk(gclk));
	jdff dff_A_NNGpHLtA3_0(.dout(w_dff_A_NK0zeahi0_0),.din(w_dff_A_NNGpHLtA3_0),.clk(gclk));
	jdff dff_A_NK0zeahi0_0(.dout(w_dff_A_vrxORiO87_0),.din(w_dff_A_NK0zeahi0_0),.clk(gclk));
	jdff dff_A_vrxORiO87_0(.dout(w_dff_A_iRnrcSFN8_0),.din(w_dff_A_vrxORiO87_0),.clk(gclk));
	jdff dff_A_iRnrcSFN8_0(.dout(w_dff_A_vRfM4m8o0_0),.din(w_dff_A_iRnrcSFN8_0),.clk(gclk));
	jdff dff_A_vRfM4m8o0_0(.dout(w_dff_A_wWnhpshe5_0),.din(w_dff_A_vRfM4m8o0_0),.clk(gclk));
	jdff dff_A_wWnhpshe5_0(.dout(w_dff_A_JzeHmLeB7_0),.din(w_dff_A_wWnhpshe5_0),.clk(gclk));
	jdff dff_A_JzeHmLeB7_0(.dout(w_dff_A_6UzM0ipI4_0),.din(w_dff_A_JzeHmLeB7_0),.clk(gclk));
	jdff dff_A_6UzM0ipI4_0(.dout(w_dff_A_Z4IxsRvl0_0),.din(w_dff_A_6UzM0ipI4_0),.clk(gclk));
	jdff dff_A_Z4IxsRvl0_0(.dout(w_dff_A_hemLPamn5_0),.din(w_dff_A_Z4IxsRvl0_0),.clk(gclk));
	jdff dff_A_hemLPamn5_0(.dout(w_dff_A_K8mVxuH75_0),.din(w_dff_A_hemLPamn5_0),.clk(gclk));
	jdff dff_A_K8mVxuH75_0(.dout(w_dff_A_RPtz7jam2_0),.din(w_dff_A_K8mVxuH75_0),.clk(gclk));
	jdff dff_A_RPtz7jam2_0(.dout(w_dff_A_hgm0GLFr8_0),.din(w_dff_A_RPtz7jam2_0),.clk(gclk));
	jdff dff_A_hgm0GLFr8_0(.dout(w_dff_A_cEMixir65_0),.din(w_dff_A_hgm0GLFr8_0),.clk(gclk));
	jdff dff_A_cEMixir65_0(.dout(w_dff_A_lHSRB4If0_0),.din(w_dff_A_cEMixir65_0),.clk(gclk));
	jdff dff_A_lHSRB4If0_0(.dout(w_dff_A_7DiyNd2U7_0),.din(w_dff_A_lHSRB4If0_0),.clk(gclk));
	jdff dff_A_7DiyNd2U7_0(.dout(w_dff_A_NEKHCgtP6_0),.din(w_dff_A_7DiyNd2U7_0),.clk(gclk));
	jdff dff_A_NEKHCgtP6_0(.dout(w_dff_A_fJ9wCbnK3_0),.din(w_dff_A_NEKHCgtP6_0),.clk(gclk));
	jdff dff_A_fJ9wCbnK3_0(.dout(w_dff_A_PBtBLRCE7_0),.din(w_dff_A_fJ9wCbnK3_0),.clk(gclk));
	jdff dff_A_PBtBLRCE7_0(.dout(w_dff_A_2sK6pDFq1_0),.din(w_dff_A_PBtBLRCE7_0),.clk(gclk));
	jdff dff_A_2sK6pDFq1_0(.dout(w_dff_A_zKLxZxQ44_0),.din(w_dff_A_2sK6pDFq1_0),.clk(gclk));
	jdff dff_A_zKLxZxQ44_0(.dout(w_dff_A_jA7dYkxF0_0),.din(w_dff_A_zKLxZxQ44_0),.clk(gclk));
	jdff dff_A_jA7dYkxF0_0(.dout(G410),.din(w_dff_A_jA7dYkxF0_0),.clk(gclk));
	jdff dff_A_Vu8cR4Jp7_1(.dout(w_dff_A_5i8cpLHb5_0),.din(w_dff_A_Vu8cR4Jp7_1),.clk(gclk));
	jdff dff_A_5i8cpLHb5_0(.dout(w_dff_A_DMpA8Top1_0),.din(w_dff_A_5i8cpLHb5_0),.clk(gclk));
	jdff dff_A_DMpA8Top1_0(.dout(w_dff_A_qwTR4BgR4_0),.din(w_dff_A_DMpA8Top1_0),.clk(gclk));
	jdff dff_A_qwTR4BgR4_0(.dout(w_dff_A_dmW5sze64_0),.din(w_dff_A_qwTR4BgR4_0),.clk(gclk));
	jdff dff_A_dmW5sze64_0(.dout(w_dff_A_nyK44cbR3_0),.din(w_dff_A_dmW5sze64_0),.clk(gclk));
	jdff dff_A_nyK44cbR3_0(.dout(w_dff_A_wStYp6HT4_0),.din(w_dff_A_nyK44cbR3_0),.clk(gclk));
	jdff dff_A_wStYp6HT4_0(.dout(w_dff_A_VaIU62lX1_0),.din(w_dff_A_wStYp6HT4_0),.clk(gclk));
	jdff dff_A_VaIU62lX1_0(.dout(w_dff_A_s3ZZiT9V0_0),.din(w_dff_A_VaIU62lX1_0),.clk(gclk));
	jdff dff_A_s3ZZiT9V0_0(.dout(w_dff_A_fcSOBhbo1_0),.din(w_dff_A_s3ZZiT9V0_0),.clk(gclk));
	jdff dff_A_fcSOBhbo1_0(.dout(w_dff_A_64DurM4V4_0),.din(w_dff_A_fcSOBhbo1_0),.clk(gclk));
	jdff dff_A_64DurM4V4_0(.dout(w_dff_A_ZHpPe69W6_0),.din(w_dff_A_64DurM4V4_0),.clk(gclk));
	jdff dff_A_ZHpPe69W6_0(.dout(w_dff_A_jKtpQYMP9_0),.din(w_dff_A_ZHpPe69W6_0),.clk(gclk));
	jdff dff_A_jKtpQYMP9_0(.dout(w_dff_A_gPhuUl9e5_0),.din(w_dff_A_jKtpQYMP9_0),.clk(gclk));
	jdff dff_A_gPhuUl9e5_0(.dout(w_dff_A_rdnhWoVd3_0),.din(w_dff_A_gPhuUl9e5_0),.clk(gclk));
	jdff dff_A_rdnhWoVd3_0(.dout(w_dff_A_kaewQR4S1_0),.din(w_dff_A_rdnhWoVd3_0),.clk(gclk));
	jdff dff_A_kaewQR4S1_0(.dout(w_dff_A_K3hv1RBr7_0),.din(w_dff_A_kaewQR4S1_0),.clk(gclk));
	jdff dff_A_K3hv1RBr7_0(.dout(w_dff_A_VVggvK314_0),.din(w_dff_A_K3hv1RBr7_0),.clk(gclk));
	jdff dff_A_VVggvK314_0(.dout(w_dff_A_TYQzpptT9_0),.din(w_dff_A_VVggvK314_0),.clk(gclk));
	jdff dff_A_TYQzpptT9_0(.dout(w_dff_A_5nTvMQDm1_0),.din(w_dff_A_TYQzpptT9_0),.clk(gclk));
	jdff dff_A_5nTvMQDm1_0(.dout(w_dff_A_Rd1xvNJk0_0),.din(w_dff_A_5nTvMQDm1_0),.clk(gclk));
	jdff dff_A_Rd1xvNJk0_0(.dout(w_dff_A_lpTnLFOU4_0),.din(w_dff_A_Rd1xvNJk0_0),.clk(gclk));
	jdff dff_A_lpTnLFOU4_0(.dout(w_dff_A_Kdortbxs2_0),.din(w_dff_A_lpTnLFOU4_0),.clk(gclk));
	jdff dff_A_Kdortbxs2_0(.dout(w_dff_A_jF6WUCVy7_0),.din(w_dff_A_Kdortbxs2_0),.clk(gclk));
	jdff dff_A_jF6WUCVy7_0(.dout(w_dff_A_fknDQMDx4_0),.din(w_dff_A_jF6WUCVy7_0),.clk(gclk));
	jdff dff_A_fknDQMDx4_0(.dout(w_dff_A_tmDtVvh60_0),.din(w_dff_A_fknDQMDx4_0),.clk(gclk));
	jdff dff_A_tmDtVvh60_0(.dout(w_dff_A_AP9pPwuU0_0),.din(w_dff_A_tmDtVvh60_0),.clk(gclk));
	jdff dff_A_AP9pPwuU0_0(.dout(w_dff_A_qEDjwCFU2_0),.din(w_dff_A_AP9pPwuU0_0),.clk(gclk));
	jdff dff_A_qEDjwCFU2_0(.dout(w_dff_A_ZxQnCWNX0_0),.din(w_dff_A_qEDjwCFU2_0),.clk(gclk));
	jdff dff_A_ZxQnCWNX0_0(.dout(w_dff_A_N3niM0mL6_0),.din(w_dff_A_ZxQnCWNX0_0),.clk(gclk));
	jdff dff_A_N3niM0mL6_0(.dout(w_dff_A_MESrp0w46_0),.din(w_dff_A_N3niM0mL6_0),.clk(gclk));
	jdff dff_A_MESrp0w46_0(.dout(w_dff_A_VydHrt5f2_0),.din(w_dff_A_MESrp0w46_0),.clk(gclk));
	jdff dff_A_VydHrt5f2_0(.dout(w_dff_A_KwPWcltU3_0),.din(w_dff_A_VydHrt5f2_0),.clk(gclk));
	jdff dff_A_KwPWcltU3_0(.dout(w_dff_A_O6iDQXGb4_0),.din(w_dff_A_KwPWcltU3_0),.clk(gclk));
	jdff dff_A_O6iDQXGb4_0(.dout(w_dff_A_pK8l7x282_0),.din(w_dff_A_O6iDQXGb4_0),.clk(gclk));
	jdff dff_A_pK8l7x282_0(.dout(w_dff_A_oZ17SNP94_0),.din(w_dff_A_pK8l7x282_0),.clk(gclk));
	jdff dff_A_oZ17SNP94_0(.dout(w_dff_A_3k3A0XI34_0),.din(w_dff_A_oZ17SNP94_0),.clk(gclk));
	jdff dff_A_3k3A0XI34_0(.dout(w_dff_A_B6U3A0sW5_0),.din(w_dff_A_3k3A0XI34_0),.clk(gclk));
	jdff dff_A_B6U3A0sW5_0(.dout(w_dff_A_cUs6tElO5_0),.din(w_dff_A_B6U3A0sW5_0),.clk(gclk));
	jdff dff_A_cUs6tElO5_0(.dout(G432),.din(w_dff_A_cUs6tElO5_0),.clk(gclk));
	jdff dff_A_5vq1NzK46_1(.dout(w_dff_A_RWhZPeyn5_0),.din(w_dff_A_5vq1NzK46_1),.clk(gclk));
	jdff dff_A_RWhZPeyn5_0(.dout(w_dff_A_69t1KPyU5_0),.din(w_dff_A_RWhZPeyn5_0),.clk(gclk));
	jdff dff_A_69t1KPyU5_0(.dout(w_dff_A_oRLo3DGd9_0),.din(w_dff_A_69t1KPyU5_0),.clk(gclk));
	jdff dff_A_oRLo3DGd9_0(.dout(w_dff_A_bG0dqtIO2_0),.din(w_dff_A_oRLo3DGd9_0),.clk(gclk));
	jdff dff_A_bG0dqtIO2_0(.dout(w_dff_A_4d62k3gL4_0),.din(w_dff_A_bG0dqtIO2_0),.clk(gclk));
	jdff dff_A_4d62k3gL4_0(.dout(w_dff_A_AqzIaTTa0_0),.din(w_dff_A_4d62k3gL4_0),.clk(gclk));
	jdff dff_A_AqzIaTTa0_0(.dout(w_dff_A_LrVSuCY69_0),.din(w_dff_A_AqzIaTTa0_0),.clk(gclk));
	jdff dff_A_LrVSuCY69_0(.dout(w_dff_A_ZTk8f71O4_0),.din(w_dff_A_LrVSuCY69_0),.clk(gclk));
	jdff dff_A_ZTk8f71O4_0(.dout(w_dff_A_DzSrgD5D8_0),.din(w_dff_A_ZTk8f71O4_0),.clk(gclk));
	jdff dff_A_DzSrgD5D8_0(.dout(w_dff_A_J5bLCuQa5_0),.din(w_dff_A_DzSrgD5D8_0),.clk(gclk));
	jdff dff_A_J5bLCuQa5_0(.dout(w_dff_A_HKjWBDn83_0),.din(w_dff_A_J5bLCuQa5_0),.clk(gclk));
	jdff dff_A_HKjWBDn83_0(.dout(w_dff_A_kyJOby1d8_0),.din(w_dff_A_HKjWBDn83_0),.clk(gclk));
	jdff dff_A_kyJOby1d8_0(.dout(w_dff_A_EtL645nO0_0),.din(w_dff_A_kyJOby1d8_0),.clk(gclk));
	jdff dff_A_EtL645nO0_0(.dout(w_dff_A_R05f0I603_0),.din(w_dff_A_EtL645nO0_0),.clk(gclk));
	jdff dff_A_R05f0I603_0(.dout(w_dff_A_lNBHcHsV8_0),.din(w_dff_A_R05f0I603_0),.clk(gclk));
	jdff dff_A_lNBHcHsV8_0(.dout(w_dff_A_nfPGEAUK3_0),.din(w_dff_A_lNBHcHsV8_0),.clk(gclk));
	jdff dff_A_nfPGEAUK3_0(.dout(w_dff_A_PNtiR7ui6_0),.din(w_dff_A_nfPGEAUK3_0),.clk(gclk));
	jdff dff_A_PNtiR7ui6_0(.dout(w_dff_A_4w1V4leJ9_0),.din(w_dff_A_PNtiR7ui6_0),.clk(gclk));
	jdff dff_A_4w1V4leJ9_0(.dout(w_dff_A_xTQhv5cJ1_0),.din(w_dff_A_4w1V4leJ9_0),.clk(gclk));
	jdff dff_A_xTQhv5cJ1_0(.dout(w_dff_A_d9pzY2252_0),.din(w_dff_A_xTQhv5cJ1_0),.clk(gclk));
	jdff dff_A_d9pzY2252_0(.dout(w_dff_A_ZXUZEbvX1_0),.din(w_dff_A_d9pzY2252_0),.clk(gclk));
	jdff dff_A_ZXUZEbvX1_0(.dout(w_dff_A_tFuMzwrz1_0),.din(w_dff_A_ZXUZEbvX1_0),.clk(gclk));
	jdff dff_A_tFuMzwrz1_0(.dout(w_dff_A_fnFz8lJJ6_0),.din(w_dff_A_tFuMzwrz1_0),.clk(gclk));
	jdff dff_A_fnFz8lJJ6_0(.dout(w_dff_A_YX0uaIbB1_0),.din(w_dff_A_fnFz8lJJ6_0),.clk(gclk));
	jdff dff_A_YX0uaIbB1_0(.dout(w_dff_A_cE95QgSE5_0),.din(w_dff_A_YX0uaIbB1_0),.clk(gclk));
	jdff dff_A_cE95QgSE5_0(.dout(w_dff_A_ATLcBc094_0),.din(w_dff_A_cE95QgSE5_0),.clk(gclk));
	jdff dff_A_ATLcBc094_0(.dout(w_dff_A_OyHI66Sc8_0),.din(w_dff_A_ATLcBc094_0),.clk(gclk));
	jdff dff_A_OyHI66Sc8_0(.dout(w_dff_A_v9n2gnZu9_0),.din(w_dff_A_OyHI66Sc8_0),.clk(gclk));
	jdff dff_A_v9n2gnZu9_0(.dout(w_dff_A_3HL1oRR98_0),.din(w_dff_A_v9n2gnZu9_0),.clk(gclk));
	jdff dff_A_3HL1oRR98_0(.dout(w_dff_A_RBvs5vBl3_0),.din(w_dff_A_3HL1oRR98_0),.clk(gclk));
	jdff dff_A_RBvs5vBl3_0(.dout(w_dff_A_9UTDv1vd6_0),.din(w_dff_A_RBvs5vBl3_0),.clk(gclk));
	jdff dff_A_9UTDv1vd6_0(.dout(w_dff_A_BWBcdv017_0),.din(w_dff_A_9UTDv1vd6_0),.clk(gclk));
	jdff dff_A_BWBcdv017_0(.dout(w_dff_A_eyrzJ9co8_0),.din(w_dff_A_BWBcdv017_0),.clk(gclk));
	jdff dff_A_eyrzJ9co8_0(.dout(w_dff_A_HUPnCAvo6_0),.din(w_dff_A_eyrzJ9co8_0),.clk(gclk));
	jdff dff_A_HUPnCAvo6_0(.dout(w_dff_A_Q1owd4z01_0),.din(w_dff_A_HUPnCAvo6_0),.clk(gclk));
	jdff dff_A_Q1owd4z01_0(.dout(w_dff_A_N90zrYVj4_0),.din(w_dff_A_Q1owd4z01_0),.clk(gclk));
	jdff dff_A_N90zrYVj4_0(.dout(w_dff_A_xgtMHEqH5_0),.din(w_dff_A_N90zrYVj4_0),.clk(gclk));
	jdff dff_A_xgtMHEqH5_0(.dout(w_dff_A_7DFVRbGw8_0),.din(w_dff_A_xgtMHEqH5_0),.clk(gclk));
	jdff dff_A_7DFVRbGw8_0(.dout(G446),.din(w_dff_A_7DFVRbGw8_0),.clk(gclk));
	jdff dff_A_wmykSRR86_2(.dout(w_dff_A_Z51GU5HB7_0),.din(w_dff_A_wmykSRR86_2),.clk(gclk));
	jdff dff_A_Z51GU5HB7_0(.dout(w_dff_A_zGrKeZqZ5_0),.din(w_dff_A_Z51GU5HB7_0),.clk(gclk));
	jdff dff_A_zGrKeZqZ5_0(.dout(w_dff_A_PXuxDnnM5_0),.din(w_dff_A_zGrKeZqZ5_0),.clk(gclk));
	jdff dff_A_PXuxDnnM5_0(.dout(w_dff_A_ol68DJzv4_0),.din(w_dff_A_PXuxDnnM5_0),.clk(gclk));
	jdff dff_A_ol68DJzv4_0(.dout(w_dff_A_AOORy8nP5_0),.din(w_dff_A_ol68DJzv4_0),.clk(gclk));
	jdff dff_A_AOORy8nP5_0(.dout(w_dff_A_XCwxvokX3_0),.din(w_dff_A_AOORy8nP5_0),.clk(gclk));
	jdff dff_A_XCwxvokX3_0(.dout(w_dff_A_F6HjEGE46_0),.din(w_dff_A_XCwxvokX3_0),.clk(gclk));
	jdff dff_A_F6HjEGE46_0(.dout(w_dff_A_5lelyWJW0_0),.din(w_dff_A_F6HjEGE46_0),.clk(gclk));
	jdff dff_A_5lelyWJW0_0(.dout(w_dff_A_YIzQye5Q8_0),.din(w_dff_A_5lelyWJW0_0),.clk(gclk));
	jdff dff_A_YIzQye5Q8_0(.dout(w_dff_A_imD8Z55Y9_0),.din(w_dff_A_YIzQye5Q8_0),.clk(gclk));
	jdff dff_A_imD8Z55Y9_0(.dout(w_dff_A_OHJsVG1g2_0),.din(w_dff_A_imD8Z55Y9_0),.clk(gclk));
	jdff dff_A_OHJsVG1g2_0(.dout(w_dff_A_GHJmHHPj3_0),.din(w_dff_A_OHJsVG1g2_0),.clk(gclk));
	jdff dff_A_GHJmHHPj3_0(.dout(w_dff_A_WpU0gC1M2_0),.din(w_dff_A_GHJmHHPj3_0),.clk(gclk));
	jdff dff_A_WpU0gC1M2_0(.dout(w_dff_A_C3w5BKHM3_0),.din(w_dff_A_WpU0gC1M2_0),.clk(gclk));
	jdff dff_A_C3w5BKHM3_0(.dout(w_dff_A_WhEpmYTP2_0),.din(w_dff_A_C3w5BKHM3_0),.clk(gclk));
	jdff dff_A_WhEpmYTP2_0(.dout(w_dff_A_T97Vuu3R3_0),.din(w_dff_A_WhEpmYTP2_0),.clk(gclk));
	jdff dff_A_T97Vuu3R3_0(.dout(w_dff_A_GRGcX3AD1_0),.din(w_dff_A_T97Vuu3R3_0),.clk(gclk));
	jdff dff_A_GRGcX3AD1_0(.dout(w_dff_A_8A0qKjGt6_0),.din(w_dff_A_GRGcX3AD1_0),.clk(gclk));
	jdff dff_A_8A0qKjGt6_0(.dout(w_dff_A_Vkh5GnhK1_0),.din(w_dff_A_8A0qKjGt6_0),.clk(gclk));
	jdff dff_A_Vkh5GnhK1_0(.dout(w_dff_A_5B6xlWj57_0),.din(w_dff_A_Vkh5GnhK1_0),.clk(gclk));
	jdff dff_A_5B6xlWj57_0(.dout(w_dff_A_Dx3Vfwf22_0),.din(w_dff_A_5B6xlWj57_0),.clk(gclk));
	jdff dff_A_Dx3Vfwf22_0(.dout(w_dff_A_MZjFnhSg8_0),.din(w_dff_A_Dx3Vfwf22_0),.clk(gclk));
	jdff dff_A_MZjFnhSg8_0(.dout(w_dff_A_gtXoUYHa9_0),.din(w_dff_A_MZjFnhSg8_0),.clk(gclk));
	jdff dff_A_gtXoUYHa9_0(.dout(w_dff_A_fS6QIagt1_0),.din(w_dff_A_gtXoUYHa9_0),.clk(gclk));
	jdff dff_A_fS6QIagt1_0(.dout(w_dff_A_VjFsIsaQ0_0),.din(w_dff_A_fS6QIagt1_0),.clk(gclk));
	jdff dff_A_VjFsIsaQ0_0(.dout(w_dff_A_uRNgKGz43_0),.din(w_dff_A_VjFsIsaQ0_0),.clk(gclk));
	jdff dff_A_uRNgKGz43_0(.dout(w_dff_A_lggBUf2K4_0),.din(w_dff_A_uRNgKGz43_0),.clk(gclk));
	jdff dff_A_lggBUf2K4_0(.dout(w_dff_A_eGhgYgQh1_0),.din(w_dff_A_lggBUf2K4_0),.clk(gclk));
	jdff dff_A_eGhgYgQh1_0(.dout(w_dff_A_Ffwg5ycn5_0),.din(w_dff_A_eGhgYgQh1_0),.clk(gclk));
	jdff dff_A_Ffwg5ycn5_0(.dout(w_dff_A_3F30JImT4_0),.din(w_dff_A_Ffwg5ycn5_0),.clk(gclk));
	jdff dff_A_3F30JImT4_0(.dout(w_dff_A_VUe7KyNH7_0),.din(w_dff_A_3F30JImT4_0),.clk(gclk));
	jdff dff_A_VUe7KyNH7_0(.dout(w_dff_A_7TtxzLVg4_0),.din(w_dff_A_VUe7KyNH7_0),.clk(gclk));
	jdff dff_A_7TtxzLVg4_0(.dout(w_dff_A_cus4gAfG4_0),.din(w_dff_A_7TtxzLVg4_0),.clk(gclk));
	jdff dff_A_cus4gAfG4_0(.dout(w_dff_A_WQRpURD65_0),.din(w_dff_A_cus4gAfG4_0),.clk(gclk));
	jdff dff_A_WQRpURD65_0(.dout(w_dff_A_lyW3cX1Q4_0),.din(w_dff_A_WQRpURD65_0),.clk(gclk));
	jdff dff_A_lyW3cX1Q4_0(.dout(w_dff_A_Kr8Zppao6_0),.din(w_dff_A_lyW3cX1Q4_0),.clk(gclk));
	jdff dff_A_Kr8Zppao6_0(.dout(G284),.din(w_dff_A_Kr8Zppao6_0),.clk(gclk));
	jdff dff_A_LK3Lj7IW8_1(.dout(w_dff_A_vv713Bvq1_0),.din(w_dff_A_LK3Lj7IW8_1),.clk(gclk));
	jdff dff_A_vv713Bvq1_0(.dout(w_dff_A_zEbL5uDi0_0),.din(w_dff_A_vv713Bvq1_0),.clk(gclk));
	jdff dff_A_zEbL5uDi0_0(.dout(w_dff_A_SQp6LKnd4_0),.din(w_dff_A_zEbL5uDi0_0),.clk(gclk));
	jdff dff_A_SQp6LKnd4_0(.dout(w_dff_A_PQYNnWu59_0),.din(w_dff_A_SQp6LKnd4_0),.clk(gclk));
	jdff dff_A_PQYNnWu59_0(.dout(w_dff_A_ZyBpAdI46_0),.din(w_dff_A_PQYNnWu59_0),.clk(gclk));
	jdff dff_A_ZyBpAdI46_0(.dout(w_dff_A_YTqWs3Sx5_0),.din(w_dff_A_ZyBpAdI46_0),.clk(gclk));
	jdff dff_A_YTqWs3Sx5_0(.dout(w_dff_A_Nyh6K99J5_0),.din(w_dff_A_YTqWs3Sx5_0),.clk(gclk));
	jdff dff_A_Nyh6K99J5_0(.dout(w_dff_A_vbwYQ40B2_0),.din(w_dff_A_Nyh6K99J5_0),.clk(gclk));
	jdff dff_A_vbwYQ40B2_0(.dout(w_dff_A_fm3Ygbhl8_0),.din(w_dff_A_vbwYQ40B2_0),.clk(gclk));
	jdff dff_A_fm3Ygbhl8_0(.dout(w_dff_A_nGFsQlsp1_0),.din(w_dff_A_fm3Ygbhl8_0),.clk(gclk));
	jdff dff_A_nGFsQlsp1_0(.dout(w_dff_A_0EKOTzA42_0),.din(w_dff_A_nGFsQlsp1_0),.clk(gclk));
	jdff dff_A_0EKOTzA42_0(.dout(w_dff_A_D2xOMZRz9_0),.din(w_dff_A_0EKOTzA42_0),.clk(gclk));
	jdff dff_A_D2xOMZRz9_0(.dout(w_dff_A_KgnTolMr3_0),.din(w_dff_A_D2xOMZRz9_0),.clk(gclk));
	jdff dff_A_KgnTolMr3_0(.dout(w_dff_A_lJp42sc29_0),.din(w_dff_A_KgnTolMr3_0),.clk(gclk));
	jdff dff_A_lJp42sc29_0(.dout(w_dff_A_ghXbvJ1f8_0),.din(w_dff_A_lJp42sc29_0),.clk(gclk));
	jdff dff_A_ghXbvJ1f8_0(.dout(w_dff_A_uy9TUzlO2_0),.din(w_dff_A_ghXbvJ1f8_0),.clk(gclk));
	jdff dff_A_uy9TUzlO2_0(.dout(w_dff_A_2hZ8ETyn4_0),.din(w_dff_A_uy9TUzlO2_0),.clk(gclk));
	jdff dff_A_2hZ8ETyn4_0(.dout(w_dff_A_7jQfeHko0_0),.din(w_dff_A_2hZ8ETyn4_0),.clk(gclk));
	jdff dff_A_7jQfeHko0_0(.dout(w_dff_A_A8HAJWnj9_0),.din(w_dff_A_7jQfeHko0_0),.clk(gclk));
	jdff dff_A_A8HAJWnj9_0(.dout(w_dff_A_HVcHDPwV4_0),.din(w_dff_A_A8HAJWnj9_0),.clk(gclk));
	jdff dff_A_HVcHDPwV4_0(.dout(w_dff_A_SMhDs7gf6_0),.din(w_dff_A_HVcHDPwV4_0),.clk(gclk));
	jdff dff_A_SMhDs7gf6_0(.dout(w_dff_A_af1a85sD4_0),.din(w_dff_A_SMhDs7gf6_0),.clk(gclk));
	jdff dff_A_af1a85sD4_0(.dout(w_dff_A_fqstAJLj5_0),.din(w_dff_A_af1a85sD4_0),.clk(gclk));
	jdff dff_A_fqstAJLj5_0(.dout(w_dff_A_bJdLdHTK8_0),.din(w_dff_A_fqstAJLj5_0),.clk(gclk));
	jdff dff_A_bJdLdHTK8_0(.dout(w_dff_A_3tPXQOIt0_0),.din(w_dff_A_bJdLdHTK8_0),.clk(gclk));
	jdff dff_A_3tPXQOIt0_0(.dout(w_dff_A_UJc8fYiZ0_0),.din(w_dff_A_3tPXQOIt0_0),.clk(gclk));
	jdff dff_A_UJc8fYiZ0_0(.dout(w_dff_A_TERPNisl1_0),.din(w_dff_A_UJc8fYiZ0_0),.clk(gclk));
	jdff dff_A_TERPNisl1_0(.dout(w_dff_A_8RV9zaeB0_0),.din(w_dff_A_TERPNisl1_0),.clk(gclk));
	jdff dff_A_8RV9zaeB0_0(.dout(w_dff_A_Fq8lh1uI3_0),.din(w_dff_A_8RV9zaeB0_0),.clk(gclk));
	jdff dff_A_Fq8lh1uI3_0(.dout(w_dff_A_PLbobi7e6_0),.din(w_dff_A_Fq8lh1uI3_0),.clk(gclk));
	jdff dff_A_PLbobi7e6_0(.dout(w_dff_A_gAWdG71D4_0),.din(w_dff_A_PLbobi7e6_0),.clk(gclk));
	jdff dff_A_gAWdG71D4_0(.dout(w_dff_A_YQMTkIYH3_0),.din(w_dff_A_gAWdG71D4_0),.clk(gclk));
	jdff dff_A_YQMTkIYH3_0(.dout(w_dff_A_x8BFfMcg6_0),.din(w_dff_A_YQMTkIYH3_0),.clk(gclk));
	jdff dff_A_x8BFfMcg6_0(.dout(w_dff_A_c0YvDkVh3_0),.din(w_dff_A_x8BFfMcg6_0),.clk(gclk));
	jdff dff_A_c0YvDkVh3_0(.dout(w_dff_A_bZSNPdQs8_0),.din(w_dff_A_c0YvDkVh3_0),.clk(gclk));
	jdff dff_A_bZSNPdQs8_0(.dout(w_dff_A_xcQwQ9SM8_0),.din(w_dff_A_bZSNPdQs8_0),.clk(gclk));
	jdff dff_A_xcQwQ9SM8_0(.dout(w_dff_A_m9WXrRFw4_0),.din(w_dff_A_xcQwQ9SM8_0),.clk(gclk));
	jdff dff_A_m9WXrRFw4_0(.dout(G286),.din(w_dff_A_m9WXrRFw4_0),.clk(gclk));
	jdff dff_A_Zda8mllT3_2(.dout(w_dff_A_ANWSoPVe0_0),.din(w_dff_A_Zda8mllT3_2),.clk(gclk));
	jdff dff_A_ANWSoPVe0_0(.dout(w_dff_A_ENPSlR9V8_0),.din(w_dff_A_ANWSoPVe0_0),.clk(gclk));
	jdff dff_A_ENPSlR9V8_0(.dout(w_dff_A_tr6UedhH1_0),.din(w_dff_A_ENPSlR9V8_0),.clk(gclk));
	jdff dff_A_tr6UedhH1_0(.dout(w_dff_A_o2mxWgGN3_0),.din(w_dff_A_tr6UedhH1_0),.clk(gclk));
	jdff dff_A_o2mxWgGN3_0(.dout(w_dff_A_fPCIrz2y1_0),.din(w_dff_A_o2mxWgGN3_0),.clk(gclk));
	jdff dff_A_fPCIrz2y1_0(.dout(w_dff_A_DZkV7ReE7_0),.din(w_dff_A_fPCIrz2y1_0),.clk(gclk));
	jdff dff_A_DZkV7ReE7_0(.dout(w_dff_A_S5GL391M7_0),.din(w_dff_A_DZkV7ReE7_0),.clk(gclk));
	jdff dff_A_S5GL391M7_0(.dout(w_dff_A_wlig9YlB9_0),.din(w_dff_A_S5GL391M7_0),.clk(gclk));
	jdff dff_A_wlig9YlB9_0(.dout(w_dff_A_c84YCPeC5_0),.din(w_dff_A_wlig9YlB9_0),.clk(gclk));
	jdff dff_A_c84YCPeC5_0(.dout(w_dff_A_kT4Seda37_0),.din(w_dff_A_c84YCPeC5_0),.clk(gclk));
	jdff dff_A_kT4Seda37_0(.dout(w_dff_A_feMNgSdp0_0),.din(w_dff_A_kT4Seda37_0),.clk(gclk));
	jdff dff_A_feMNgSdp0_0(.dout(w_dff_A_I0Tdke2j5_0),.din(w_dff_A_feMNgSdp0_0),.clk(gclk));
	jdff dff_A_I0Tdke2j5_0(.dout(w_dff_A_CT9V92q39_0),.din(w_dff_A_I0Tdke2j5_0),.clk(gclk));
	jdff dff_A_CT9V92q39_0(.dout(w_dff_A_rWJd1lxd0_0),.din(w_dff_A_CT9V92q39_0),.clk(gclk));
	jdff dff_A_rWJd1lxd0_0(.dout(w_dff_A_xmgpYhAA6_0),.din(w_dff_A_rWJd1lxd0_0),.clk(gclk));
	jdff dff_A_xmgpYhAA6_0(.dout(w_dff_A_ysMsFMnY4_0),.din(w_dff_A_xmgpYhAA6_0),.clk(gclk));
	jdff dff_A_ysMsFMnY4_0(.dout(w_dff_A_CxL67Ksl0_0),.din(w_dff_A_ysMsFMnY4_0),.clk(gclk));
	jdff dff_A_CxL67Ksl0_0(.dout(w_dff_A_GXVuplTV8_0),.din(w_dff_A_CxL67Ksl0_0),.clk(gclk));
	jdff dff_A_GXVuplTV8_0(.dout(w_dff_A_rlfxZZjm3_0),.din(w_dff_A_GXVuplTV8_0),.clk(gclk));
	jdff dff_A_rlfxZZjm3_0(.dout(w_dff_A_HR6Im4lF0_0),.din(w_dff_A_rlfxZZjm3_0),.clk(gclk));
	jdff dff_A_HR6Im4lF0_0(.dout(w_dff_A_GTRhtGmT5_0),.din(w_dff_A_HR6Im4lF0_0),.clk(gclk));
	jdff dff_A_GTRhtGmT5_0(.dout(w_dff_A_9sztd85p7_0),.din(w_dff_A_GTRhtGmT5_0),.clk(gclk));
	jdff dff_A_9sztd85p7_0(.dout(w_dff_A_bDzlcFXt1_0),.din(w_dff_A_9sztd85p7_0),.clk(gclk));
	jdff dff_A_bDzlcFXt1_0(.dout(w_dff_A_mpb3HOcT8_0),.din(w_dff_A_bDzlcFXt1_0),.clk(gclk));
	jdff dff_A_mpb3HOcT8_0(.dout(w_dff_A_B7fRJPiM1_0),.din(w_dff_A_mpb3HOcT8_0),.clk(gclk));
	jdff dff_A_B7fRJPiM1_0(.dout(w_dff_A_olsAFkr41_0),.din(w_dff_A_B7fRJPiM1_0),.clk(gclk));
	jdff dff_A_olsAFkr41_0(.dout(w_dff_A_u7o8P4pA6_0),.din(w_dff_A_olsAFkr41_0),.clk(gclk));
	jdff dff_A_u7o8P4pA6_0(.dout(w_dff_A_LEKUdH8H6_0),.din(w_dff_A_u7o8P4pA6_0),.clk(gclk));
	jdff dff_A_LEKUdH8H6_0(.dout(w_dff_A_VjIfLl0q2_0),.din(w_dff_A_LEKUdH8H6_0),.clk(gclk));
	jdff dff_A_VjIfLl0q2_0(.dout(w_dff_A_AtfvshBG0_0),.din(w_dff_A_VjIfLl0q2_0),.clk(gclk));
	jdff dff_A_AtfvshBG0_0(.dout(w_dff_A_yVvlo2nG3_0),.din(w_dff_A_AtfvshBG0_0),.clk(gclk));
	jdff dff_A_yVvlo2nG3_0(.dout(w_dff_A_amVJRz0l2_0),.din(w_dff_A_yVvlo2nG3_0),.clk(gclk));
	jdff dff_A_amVJRz0l2_0(.dout(w_dff_A_kgUi1bYH3_0),.din(w_dff_A_amVJRz0l2_0),.clk(gclk));
	jdff dff_A_kgUi1bYH3_0(.dout(w_dff_A_VkzLy2zk9_0),.din(w_dff_A_kgUi1bYH3_0),.clk(gclk));
	jdff dff_A_VkzLy2zk9_0(.dout(w_dff_A_1Q23ub1H0_0),.din(w_dff_A_VkzLy2zk9_0),.clk(gclk));
	jdff dff_A_1Q23ub1H0_0(.dout(w_dff_A_9KmSwSEi9_0),.din(w_dff_A_1Q23ub1H0_0),.clk(gclk));
	jdff dff_A_9KmSwSEi9_0(.dout(G289),.din(w_dff_A_9KmSwSEi9_0),.clk(gclk));
	jdff dff_A_D8xH8Oi22_2(.dout(w_dff_A_QeaqzpoA3_0),.din(w_dff_A_D8xH8Oi22_2),.clk(gclk));
	jdff dff_A_QeaqzpoA3_0(.dout(w_dff_A_UlKbVGnf9_0),.din(w_dff_A_QeaqzpoA3_0),.clk(gclk));
	jdff dff_A_UlKbVGnf9_0(.dout(w_dff_A_RUH0X1aq1_0),.din(w_dff_A_UlKbVGnf9_0),.clk(gclk));
	jdff dff_A_RUH0X1aq1_0(.dout(w_dff_A_LTjQI9qp2_0),.din(w_dff_A_RUH0X1aq1_0),.clk(gclk));
	jdff dff_A_LTjQI9qp2_0(.dout(w_dff_A_EFgoXyTb1_0),.din(w_dff_A_LTjQI9qp2_0),.clk(gclk));
	jdff dff_A_EFgoXyTb1_0(.dout(w_dff_A_TQYILxmN6_0),.din(w_dff_A_EFgoXyTb1_0),.clk(gclk));
	jdff dff_A_TQYILxmN6_0(.dout(w_dff_A_EV6b3my62_0),.din(w_dff_A_TQYILxmN6_0),.clk(gclk));
	jdff dff_A_EV6b3my62_0(.dout(w_dff_A_c4hGrQpA7_0),.din(w_dff_A_EV6b3my62_0),.clk(gclk));
	jdff dff_A_c4hGrQpA7_0(.dout(w_dff_A_wrxJuxDE4_0),.din(w_dff_A_c4hGrQpA7_0),.clk(gclk));
	jdff dff_A_wrxJuxDE4_0(.dout(w_dff_A_16Mm9h3l1_0),.din(w_dff_A_wrxJuxDE4_0),.clk(gclk));
	jdff dff_A_16Mm9h3l1_0(.dout(w_dff_A_I8wEl9ob2_0),.din(w_dff_A_16Mm9h3l1_0),.clk(gclk));
	jdff dff_A_I8wEl9ob2_0(.dout(w_dff_A_1wzQhIEN6_0),.din(w_dff_A_I8wEl9ob2_0),.clk(gclk));
	jdff dff_A_1wzQhIEN6_0(.dout(w_dff_A_Xqd6tnkC1_0),.din(w_dff_A_1wzQhIEN6_0),.clk(gclk));
	jdff dff_A_Xqd6tnkC1_0(.dout(w_dff_A_RLLruLqB2_0),.din(w_dff_A_Xqd6tnkC1_0),.clk(gclk));
	jdff dff_A_RLLruLqB2_0(.dout(w_dff_A_nJtGxlW45_0),.din(w_dff_A_RLLruLqB2_0),.clk(gclk));
	jdff dff_A_nJtGxlW45_0(.dout(w_dff_A_J17VpB8y7_0),.din(w_dff_A_nJtGxlW45_0),.clk(gclk));
	jdff dff_A_J17VpB8y7_0(.dout(w_dff_A_3KaJR61b6_0),.din(w_dff_A_J17VpB8y7_0),.clk(gclk));
	jdff dff_A_3KaJR61b6_0(.dout(w_dff_A_ImVMVU8X4_0),.din(w_dff_A_3KaJR61b6_0),.clk(gclk));
	jdff dff_A_ImVMVU8X4_0(.dout(w_dff_A_UvYnuncs2_0),.din(w_dff_A_ImVMVU8X4_0),.clk(gclk));
	jdff dff_A_UvYnuncs2_0(.dout(w_dff_A_FmvigApb9_0),.din(w_dff_A_UvYnuncs2_0),.clk(gclk));
	jdff dff_A_FmvigApb9_0(.dout(w_dff_A_JoVMRdbh2_0),.din(w_dff_A_FmvigApb9_0),.clk(gclk));
	jdff dff_A_JoVMRdbh2_0(.dout(w_dff_A_NsS6ZsxL4_0),.din(w_dff_A_JoVMRdbh2_0),.clk(gclk));
	jdff dff_A_NsS6ZsxL4_0(.dout(w_dff_A_GQLbrFlD0_0),.din(w_dff_A_NsS6ZsxL4_0),.clk(gclk));
	jdff dff_A_GQLbrFlD0_0(.dout(w_dff_A_tFinVVOt8_0),.din(w_dff_A_GQLbrFlD0_0),.clk(gclk));
	jdff dff_A_tFinVVOt8_0(.dout(w_dff_A_qsDEeN3N2_0),.din(w_dff_A_tFinVVOt8_0),.clk(gclk));
	jdff dff_A_qsDEeN3N2_0(.dout(w_dff_A_7tya0M0h9_0),.din(w_dff_A_qsDEeN3N2_0),.clk(gclk));
	jdff dff_A_7tya0M0h9_0(.dout(w_dff_A_hwszIDsf6_0),.din(w_dff_A_7tya0M0h9_0),.clk(gclk));
	jdff dff_A_hwszIDsf6_0(.dout(w_dff_A_NKkSuLOP3_0),.din(w_dff_A_hwszIDsf6_0),.clk(gclk));
	jdff dff_A_NKkSuLOP3_0(.dout(w_dff_A_lKQqMRGc9_0),.din(w_dff_A_NKkSuLOP3_0),.clk(gclk));
	jdff dff_A_lKQqMRGc9_0(.dout(w_dff_A_1yF2FMkm4_0),.din(w_dff_A_lKQqMRGc9_0),.clk(gclk));
	jdff dff_A_1yF2FMkm4_0(.dout(w_dff_A_UEzsUctU8_0),.din(w_dff_A_1yF2FMkm4_0),.clk(gclk));
	jdff dff_A_UEzsUctU8_0(.dout(w_dff_A_fgRZTT0e8_0),.din(w_dff_A_UEzsUctU8_0),.clk(gclk));
	jdff dff_A_fgRZTT0e8_0(.dout(w_dff_A_hvkTvSRV7_0),.din(w_dff_A_fgRZTT0e8_0),.clk(gclk));
	jdff dff_A_hvkTvSRV7_0(.dout(w_dff_A_guDGb1dG0_0),.din(w_dff_A_hvkTvSRV7_0),.clk(gclk));
	jdff dff_A_guDGb1dG0_0(.dout(w_dff_A_2lOuxi4F3_0),.din(w_dff_A_guDGb1dG0_0),.clk(gclk));
	jdff dff_A_2lOuxi4F3_0(.dout(G292),.din(w_dff_A_2lOuxi4F3_0),.clk(gclk));
	jdff dff_A_GbPQfCGT0_1(.dout(w_dff_A_irDydLFs4_0),.din(w_dff_A_GbPQfCGT0_1),.clk(gclk));
	jdff dff_A_irDydLFs4_0(.dout(w_dff_A_cDmpTu5Y2_0),.din(w_dff_A_irDydLFs4_0),.clk(gclk));
	jdff dff_A_cDmpTu5Y2_0(.dout(w_dff_A_kNrv0VxV9_0),.din(w_dff_A_cDmpTu5Y2_0),.clk(gclk));
	jdff dff_A_kNrv0VxV9_0(.dout(w_dff_A_tWLpSJRW1_0),.din(w_dff_A_kNrv0VxV9_0),.clk(gclk));
	jdff dff_A_tWLpSJRW1_0(.dout(w_dff_A_u55keSlm9_0),.din(w_dff_A_tWLpSJRW1_0),.clk(gclk));
	jdff dff_A_u55keSlm9_0(.dout(w_dff_A_Q8wsBj6h9_0),.din(w_dff_A_u55keSlm9_0),.clk(gclk));
	jdff dff_A_Q8wsBj6h9_0(.dout(w_dff_A_tplCoRQI2_0),.din(w_dff_A_Q8wsBj6h9_0),.clk(gclk));
	jdff dff_A_tplCoRQI2_0(.dout(w_dff_A_I7o8meEr5_0),.din(w_dff_A_tplCoRQI2_0),.clk(gclk));
	jdff dff_A_I7o8meEr5_0(.dout(w_dff_A_TLkILGK99_0),.din(w_dff_A_I7o8meEr5_0),.clk(gclk));
	jdff dff_A_TLkILGK99_0(.dout(w_dff_A_J2LBPLHi3_0),.din(w_dff_A_TLkILGK99_0),.clk(gclk));
	jdff dff_A_J2LBPLHi3_0(.dout(w_dff_A_Rf6o4KNF3_0),.din(w_dff_A_J2LBPLHi3_0),.clk(gclk));
	jdff dff_A_Rf6o4KNF3_0(.dout(w_dff_A_LV1LWeau9_0),.din(w_dff_A_Rf6o4KNF3_0),.clk(gclk));
	jdff dff_A_LV1LWeau9_0(.dout(w_dff_A_bamJNO4J8_0),.din(w_dff_A_LV1LWeau9_0),.clk(gclk));
	jdff dff_A_bamJNO4J8_0(.dout(w_dff_A_Dk3ozH7T4_0),.din(w_dff_A_bamJNO4J8_0),.clk(gclk));
	jdff dff_A_Dk3ozH7T4_0(.dout(w_dff_A_gbygC4fj8_0),.din(w_dff_A_Dk3ozH7T4_0),.clk(gclk));
	jdff dff_A_gbygC4fj8_0(.dout(w_dff_A_qtCeMX6g6_0),.din(w_dff_A_gbygC4fj8_0),.clk(gclk));
	jdff dff_A_qtCeMX6g6_0(.dout(w_dff_A_3lANmBzG1_0),.din(w_dff_A_qtCeMX6g6_0),.clk(gclk));
	jdff dff_A_3lANmBzG1_0(.dout(w_dff_A_Hp2aH8Te5_0),.din(w_dff_A_3lANmBzG1_0),.clk(gclk));
	jdff dff_A_Hp2aH8Te5_0(.dout(w_dff_A_5EEAs0TA0_0),.din(w_dff_A_Hp2aH8Te5_0),.clk(gclk));
	jdff dff_A_5EEAs0TA0_0(.dout(w_dff_A_vQZG6WeP3_0),.din(w_dff_A_5EEAs0TA0_0),.clk(gclk));
	jdff dff_A_vQZG6WeP3_0(.dout(w_dff_A_53xjXXvi9_0),.din(w_dff_A_vQZG6WeP3_0),.clk(gclk));
	jdff dff_A_53xjXXvi9_0(.dout(w_dff_A_DTKax7gg9_0),.din(w_dff_A_53xjXXvi9_0),.clk(gclk));
	jdff dff_A_DTKax7gg9_0(.dout(w_dff_A_1bQCAe5l2_0),.din(w_dff_A_DTKax7gg9_0),.clk(gclk));
	jdff dff_A_1bQCAe5l2_0(.dout(w_dff_A_ad9ZMT4Z0_0),.din(w_dff_A_1bQCAe5l2_0),.clk(gclk));
	jdff dff_A_ad9ZMT4Z0_0(.dout(w_dff_A_H6MSNFsM6_0),.din(w_dff_A_ad9ZMT4Z0_0),.clk(gclk));
	jdff dff_A_H6MSNFsM6_0(.dout(w_dff_A_SdmCZUZD1_0),.din(w_dff_A_H6MSNFsM6_0),.clk(gclk));
	jdff dff_A_SdmCZUZD1_0(.dout(w_dff_A_1N1Kpv939_0),.din(w_dff_A_SdmCZUZD1_0),.clk(gclk));
	jdff dff_A_1N1Kpv939_0(.dout(w_dff_A_qUdhMDYJ4_0),.din(w_dff_A_1N1Kpv939_0),.clk(gclk));
	jdff dff_A_qUdhMDYJ4_0(.dout(w_dff_A_HCAzTAlZ3_0),.din(w_dff_A_qUdhMDYJ4_0),.clk(gclk));
	jdff dff_A_HCAzTAlZ3_0(.dout(w_dff_A_lsPXM3Wn5_0),.din(w_dff_A_HCAzTAlZ3_0),.clk(gclk));
	jdff dff_A_lsPXM3Wn5_0(.dout(w_dff_A_e0E61vYZ3_0),.din(w_dff_A_lsPXM3Wn5_0),.clk(gclk));
	jdff dff_A_e0E61vYZ3_0(.dout(w_dff_A_ApsbvxKn4_0),.din(w_dff_A_e0E61vYZ3_0),.clk(gclk));
	jdff dff_A_ApsbvxKn4_0(.dout(w_dff_A_pnoAOqv47_0),.din(w_dff_A_ApsbvxKn4_0),.clk(gclk));
	jdff dff_A_pnoAOqv47_0(.dout(w_dff_A_QMTuUWtV1_0),.din(w_dff_A_pnoAOqv47_0),.clk(gclk));
	jdff dff_A_QMTuUWtV1_0(.dout(w_dff_A_SnxHDgde9_0),.din(w_dff_A_QMTuUWtV1_0),.clk(gclk));
	jdff dff_A_SnxHDgde9_0(.dout(w_dff_A_c9brB2b12_0),.din(w_dff_A_SnxHDgde9_0),.clk(gclk));
	jdff dff_A_c9brB2b12_0(.dout(w_dff_A_f2PAfZVx0_0),.din(w_dff_A_c9brB2b12_0),.clk(gclk));
	jdff dff_A_f2PAfZVx0_0(.dout(G341),.din(w_dff_A_f2PAfZVx0_0),.clk(gclk));
	jdff dff_A_9eF0pr3b7_2(.dout(w_dff_A_U5aihzHX7_0),.din(w_dff_A_9eF0pr3b7_2),.clk(gclk));
	jdff dff_A_U5aihzHX7_0(.dout(w_dff_A_Ebt2Dh5G4_0),.din(w_dff_A_U5aihzHX7_0),.clk(gclk));
	jdff dff_A_Ebt2Dh5G4_0(.dout(w_dff_A_UOIeNXiL8_0),.din(w_dff_A_Ebt2Dh5G4_0),.clk(gclk));
	jdff dff_A_UOIeNXiL8_0(.dout(w_dff_A_igtWn4hb3_0),.din(w_dff_A_UOIeNXiL8_0),.clk(gclk));
	jdff dff_A_igtWn4hb3_0(.dout(w_dff_A_U5APrh1d1_0),.din(w_dff_A_igtWn4hb3_0),.clk(gclk));
	jdff dff_A_U5APrh1d1_0(.dout(w_dff_A_vP9pbXTf6_0),.din(w_dff_A_U5APrh1d1_0),.clk(gclk));
	jdff dff_A_vP9pbXTf6_0(.dout(w_dff_A_dHhyIdd24_0),.din(w_dff_A_vP9pbXTf6_0),.clk(gclk));
	jdff dff_A_dHhyIdd24_0(.dout(w_dff_A_57JAJ3C18_0),.din(w_dff_A_dHhyIdd24_0),.clk(gclk));
	jdff dff_A_57JAJ3C18_0(.dout(w_dff_A_WK4SPcEo0_0),.din(w_dff_A_57JAJ3C18_0),.clk(gclk));
	jdff dff_A_WK4SPcEo0_0(.dout(w_dff_A_fMxxyZX77_0),.din(w_dff_A_WK4SPcEo0_0),.clk(gclk));
	jdff dff_A_fMxxyZX77_0(.dout(w_dff_A_YqKXUNoP6_0),.din(w_dff_A_fMxxyZX77_0),.clk(gclk));
	jdff dff_A_YqKXUNoP6_0(.dout(w_dff_A_alhtDkAp7_0),.din(w_dff_A_YqKXUNoP6_0),.clk(gclk));
	jdff dff_A_alhtDkAp7_0(.dout(w_dff_A_F3hDwAHE7_0),.din(w_dff_A_alhtDkAp7_0),.clk(gclk));
	jdff dff_A_F3hDwAHE7_0(.dout(w_dff_A_AhqxXLdX3_0),.din(w_dff_A_F3hDwAHE7_0),.clk(gclk));
	jdff dff_A_AhqxXLdX3_0(.dout(w_dff_A_m9g9MC1d9_0),.din(w_dff_A_AhqxXLdX3_0),.clk(gclk));
	jdff dff_A_m9g9MC1d9_0(.dout(w_dff_A_pj3aacqR7_0),.din(w_dff_A_m9g9MC1d9_0),.clk(gclk));
	jdff dff_A_pj3aacqR7_0(.dout(w_dff_A_aghY5Z0G6_0),.din(w_dff_A_pj3aacqR7_0),.clk(gclk));
	jdff dff_A_aghY5Z0G6_0(.dout(w_dff_A_ylHZq5le6_0),.din(w_dff_A_aghY5Z0G6_0),.clk(gclk));
	jdff dff_A_ylHZq5le6_0(.dout(w_dff_A_Jl4jzpA91_0),.din(w_dff_A_ylHZq5le6_0),.clk(gclk));
	jdff dff_A_Jl4jzpA91_0(.dout(w_dff_A_K7RRo5073_0),.din(w_dff_A_Jl4jzpA91_0),.clk(gclk));
	jdff dff_A_K7RRo5073_0(.dout(w_dff_A_ETH7nLvz9_0),.din(w_dff_A_K7RRo5073_0),.clk(gclk));
	jdff dff_A_ETH7nLvz9_0(.dout(w_dff_A_yWt2LeYO8_0),.din(w_dff_A_ETH7nLvz9_0),.clk(gclk));
	jdff dff_A_yWt2LeYO8_0(.dout(w_dff_A_HBWfBKkJ9_0),.din(w_dff_A_yWt2LeYO8_0),.clk(gclk));
	jdff dff_A_HBWfBKkJ9_0(.dout(w_dff_A_Y2KUgy323_0),.din(w_dff_A_HBWfBKkJ9_0),.clk(gclk));
	jdff dff_A_Y2KUgy323_0(.dout(w_dff_A_y9BS71jB9_0),.din(w_dff_A_Y2KUgy323_0),.clk(gclk));
	jdff dff_A_y9BS71jB9_0(.dout(w_dff_A_KJ5YL3Fu2_0),.din(w_dff_A_y9BS71jB9_0),.clk(gclk));
	jdff dff_A_KJ5YL3Fu2_0(.dout(w_dff_A_esaUVrAh2_0),.din(w_dff_A_KJ5YL3Fu2_0),.clk(gclk));
	jdff dff_A_esaUVrAh2_0(.dout(w_dff_A_ozpON0Wj9_0),.din(w_dff_A_esaUVrAh2_0),.clk(gclk));
	jdff dff_A_ozpON0Wj9_0(.dout(w_dff_A_H5pdPkaq8_0),.din(w_dff_A_ozpON0Wj9_0),.clk(gclk));
	jdff dff_A_H5pdPkaq8_0(.dout(w_dff_A_s8gxRBU05_0),.din(w_dff_A_H5pdPkaq8_0),.clk(gclk));
	jdff dff_A_s8gxRBU05_0(.dout(w_dff_A_0XLYwrdL8_0),.din(w_dff_A_s8gxRBU05_0),.clk(gclk));
	jdff dff_A_0XLYwrdL8_0(.dout(w_dff_A_CF594JrW0_0),.din(w_dff_A_0XLYwrdL8_0),.clk(gclk));
	jdff dff_A_CF594JrW0_0(.dout(w_dff_A_Z2hBtZLw1_0),.din(w_dff_A_CF594JrW0_0),.clk(gclk));
	jdff dff_A_Z2hBtZLw1_0(.dout(w_dff_A_IWgvaZ752_0),.din(w_dff_A_Z2hBtZLw1_0),.clk(gclk));
	jdff dff_A_IWgvaZ752_0(.dout(w_dff_A_4HyqLyIS7_0),.din(w_dff_A_IWgvaZ752_0),.clk(gclk));
	jdff dff_A_4HyqLyIS7_0(.dout(G281),.din(w_dff_A_4HyqLyIS7_0),.clk(gclk));
	jdff dff_A_VajKcQKi2_1(.dout(w_dff_A_iGg4Nv891_0),.din(w_dff_A_VajKcQKi2_1),.clk(gclk));
	jdff dff_A_iGg4Nv891_0(.dout(w_dff_A_25goQeuA9_0),.din(w_dff_A_iGg4Nv891_0),.clk(gclk));
	jdff dff_A_25goQeuA9_0(.dout(w_dff_A_HatPLPWP1_0),.din(w_dff_A_25goQeuA9_0),.clk(gclk));
	jdff dff_A_HatPLPWP1_0(.dout(w_dff_A_qzThAfp04_0),.din(w_dff_A_HatPLPWP1_0),.clk(gclk));
	jdff dff_A_qzThAfp04_0(.dout(w_dff_A_AhGh7UAO2_0),.din(w_dff_A_qzThAfp04_0),.clk(gclk));
	jdff dff_A_AhGh7UAO2_0(.dout(w_dff_A_ibjJ9Hns4_0),.din(w_dff_A_AhGh7UAO2_0),.clk(gclk));
	jdff dff_A_ibjJ9Hns4_0(.dout(w_dff_A_BCoYnTiM9_0),.din(w_dff_A_ibjJ9Hns4_0),.clk(gclk));
	jdff dff_A_BCoYnTiM9_0(.dout(w_dff_A_26Aud73p7_0),.din(w_dff_A_BCoYnTiM9_0),.clk(gclk));
	jdff dff_A_26Aud73p7_0(.dout(w_dff_A_TfnDFASo2_0),.din(w_dff_A_26Aud73p7_0),.clk(gclk));
	jdff dff_A_TfnDFASo2_0(.dout(w_dff_A_v2o9LzU17_0),.din(w_dff_A_TfnDFASo2_0),.clk(gclk));
	jdff dff_A_v2o9LzU17_0(.dout(w_dff_A_N9P4dUAr8_0),.din(w_dff_A_v2o9LzU17_0),.clk(gclk));
	jdff dff_A_N9P4dUAr8_0(.dout(w_dff_A_tGlkqVm22_0),.din(w_dff_A_N9P4dUAr8_0),.clk(gclk));
	jdff dff_A_tGlkqVm22_0(.dout(w_dff_A_VjHpNReM8_0),.din(w_dff_A_tGlkqVm22_0),.clk(gclk));
	jdff dff_A_VjHpNReM8_0(.dout(w_dff_A_2j0VGHDN6_0),.din(w_dff_A_VjHpNReM8_0),.clk(gclk));
	jdff dff_A_2j0VGHDN6_0(.dout(w_dff_A_IzYZAoVZ8_0),.din(w_dff_A_2j0VGHDN6_0),.clk(gclk));
	jdff dff_A_IzYZAoVZ8_0(.dout(w_dff_A_0nnwbXVY7_0),.din(w_dff_A_IzYZAoVZ8_0),.clk(gclk));
	jdff dff_A_0nnwbXVY7_0(.dout(w_dff_A_KEowFla87_0),.din(w_dff_A_0nnwbXVY7_0),.clk(gclk));
	jdff dff_A_KEowFla87_0(.dout(w_dff_A_Tpchak8d5_0),.din(w_dff_A_KEowFla87_0),.clk(gclk));
	jdff dff_A_Tpchak8d5_0(.dout(w_dff_A_av91L8Q51_0),.din(w_dff_A_Tpchak8d5_0),.clk(gclk));
	jdff dff_A_av91L8Q51_0(.dout(w_dff_A_SZXiAgwB9_0),.din(w_dff_A_av91L8Q51_0),.clk(gclk));
	jdff dff_A_SZXiAgwB9_0(.dout(w_dff_A_eucxQIuR4_0),.din(w_dff_A_SZXiAgwB9_0),.clk(gclk));
	jdff dff_A_eucxQIuR4_0(.dout(w_dff_A_uMrkjlE98_0),.din(w_dff_A_eucxQIuR4_0),.clk(gclk));
	jdff dff_A_uMrkjlE98_0(.dout(w_dff_A_PZEL2WM43_0),.din(w_dff_A_uMrkjlE98_0),.clk(gclk));
	jdff dff_A_PZEL2WM43_0(.dout(w_dff_A_eko1wODP7_0),.din(w_dff_A_PZEL2WM43_0),.clk(gclk));
	jdff dff_A_eko1wODP7_0(.dout(w_dff_A_KAN9EA0y5_0),.din(w_dff_A_eko1wODP7_0),.clk(gclk));
	jdff dff_A_KAN9EA0y5_0(.dout(w_dff_A_Bv3P9Ohy5_0),.din(w_dff_A_KAN9EA0y5_0),.clk(gclk));
	jdff dff_A_Bv3P9Ohy5_0(.dout(w_dff_A_7viZ92165_0),.din(w_dff_A_Bv3P9Ohy5_0),.clk(gclk));
	jdff dff_A_7viZ92165_0(.dout(w_dff_A_vXMDM2cu8_0),.din(w_dff_A_7viZ92165_0),.clk(gclk));
	jdff dff_A_vXMDM2cu8_0(.dout(w_dff_A_ij20ieMK5_0),.din(w_dff_A_vXMDM2cu8_0),.clk(gclk));
	jdff dff_A_ij20ieMK5_0(.dout(w_dff_A_QygmYoyv5_0),.din(w_dff_A_ij20ieMK5_0),.clk(gclk));
	jdff dff_A_QygmYoyv5_0(.dout(w_dff_A_bL4S26bH5_0),.din(w_dff_A_QygmYoyv5_0),.clk(gclk));
	jdff dff_A_bL4S26bH5_0(.dout(w_dff_A_Cg2zNbpT6_0),.din(w_dff_A_bL4S26bH5_0),.clk(gclk));
	jdff dff_A_Cg2zNbpT6_0(.dout(w_dff_A_FGeTxGOj4_0),.din(w_dff_A_Cg2zNbpT6_0),.clk(gclk));
	jdff dff_A_FGeTxGOj4_0(.dout(w_dff_A_OPflZcUf0_0),.din(w_dff_A_FGeTxGOj4_0),.clk(gclk));
	jdff dff_A_OPflZcUf0_0(.dout(w_dff_A_pCjmLV2F7_0),.din(w_dff_A_OPflZcUf0_0),.clk(gclk));
	jdff dff_A_pCjmLV2F7_0(.dout(w_dff_A_RYBntYTO7_0),.din(w_dff_A_pCjmLV2F7_0),.clk(gclk));
	jdff dff_A_RYBntYTO7_0(.dout(w_dff_A_3y7xPflI7_0),.din(w_dff_A_RYBntYTO7_0),.clk(gclk));
	jdff dff_A_3y7xPflI7_0(.dout(w_dff_A_iliYjplN9_0),.din(w_dff_A_3y7xPflI7_0),.clk(gclk));
	jdff dff_A_iliYjplN9_0(.dout(G453),.din(w_dff_A_iliYjplN9_0),.clk(gclk));
	jdff dff_A_yJxiPeRD1_2(.dout(w_dff_A_iHVGdYtC5_0),.din(w_dff_A_yJxiPeRD1_2),.clk(gclk));
	jdff dff_A_iHVGdYtC5_0(.dout(w_dff_A_Z8YN3F5L8_0),.din(w_dff_A_iHVGdYtC5_0),.clk(gclk));
	jdff dff_A_Z8YN3F5L8_0(.dout(w_dff_A_rGU61j2x4_0),.din(w_dff_A_Z8YN3F5L8_0),.clk(gclk));
	jdff dff_A_rGU61j2x4_0(.dout(w_dff_A_EUtMwiv20_0),.din(w_dff_A_rGU61j2x4_0),.clk(gclk));
	jdff dff_A_EUtMwiv20_0(.dout(w_dff_A_JK7lKOAd9_0),.din(w_dff_A_EUtMwiv20_0),.clk(gclk));
	jdff dff_A_JK7lKOAd9_0(.dout(w_dff_A_u0WiDjz06_0),.din(w_dff_A_JK7lKOAd9_0),.clk(gclk));
	jdff dff_A_u0WiDjz06_0(.dout(w_dff_A_fGrgpTCd4_0),.din(w_dff_A_u0WiDjz06_0),.clk(gclk));
	jdff dff_A_fGrgpTCd4_0(.dout(w_dff_A_cMg4yR6h7_0),.din(w_dff_A_fGrgpTCd4_0),.clk(gclk));
	jdff dff_A_cMg4yR6h7_0(.dout(w_dff_A_VcRvXCnt1_0),.din(w_dff_A_cMg4yR6h7_0),.clk(gclk));
	jdff dff_A_VcRvXCnt1_0(.dout(w_dff_A_ppGeXKRj7_0),.din(w_dff_A_VcRvXCnt1_0),.clk(gclk));
	jdff dff_A_ppGeXKRj7_0(.dout(w_dff_A_uUrkPgJd2_0),.din(w_dff_A_ppGeXKRj7_0),.clk(gclk));
	jdff dff_A_uUrkPgJd2_0(.dout(w_dff_A_gwWwRlz55_0),.din(w_dff_A_uUrkPgJd2_0),.clk(gclk));
	jdff dff_A_gwWwRlz55_0(.dout(w_dff_A_8885U0Yd4_0),.din(w_dff_A_gwWwRlz55_0),.clk(gclk));
	jdff dff_A_8885U0Yd4_0(.dout(w_dff_A_z6AFslYN4_0),.din(w_dff_A_8885U0Yd4_0),.clk(gclk));
	jdff dff_A_z6AFslYN4_0(.dout(w_dff_A_HAPUPDnJ5_0),.din(w_dff_A_z6AFslYN4_0),.clk(gclk));
	jdff dff_A_HAPUPDnJ5_0(.dout(w_dff_A_ifnRkYcn9_0),.din(w_dff_A_HAPUPDnJ5_0),.clk(gclk));
	jdff dff_A_ifnRkYcn9_0(.dout(w_dff_A_PUCYaq8L6_0),.din(w_dff_A_ifnRkYcn9_0),.clk(gclk));
	jdff dff_A_PUCYaq8L6_0(.dout(w_dff_A_q5YU6Sbn5_0),.din(w_dff_A_PUCYaq8L6_0),.clk(gclk));
	jdff dff_A_q5YU6Sbn5_0(.dout(w_dff_A_bojcxAPn8_0),.din(w_dff_A_q5YU6Sbn5_0),.clk(gclk));
	jdff dff_A_bojcxAPn8_0(.dout(w_dff_A_fnS28SFh7_0),.din(w_dff_A_bojcxAPn8_0),.clk(gclk));
	jdff dff_A_fnS28SFh7_0(.dout(w_dff_A_fK8fBM9u7_0),.din(w_dff_A_fnS28SFh7_0),.clk(gclk));
	jdff dff_A_fK8fBM9u7_0(.dout(w_dff_A_xW1zuY2b6_0),.din(w_dff_A_fK8fBM9u7_0),.clk(gclk));
	jdff dff_A_xW1zuY2b6_0(.dout(w_dff_A_4oh8RdhF9_0),.din(w_dff_A_xW1zuY2b6_0),.clk(gclk));
	jdff dff_A_4oh8RdhF9_0(.dout(w_dff_A_E2dOlFAB5_0),.din(w_dff_A_4oh8RdhF9_0),.clk(gclk));
	jdff dff_A_E2dOlFAB5_0(.dout(w_dff_A_5eKDupkb3_0),.din(w_dff_A_E2dOlFAB5_0),.clk(gclk));
	jdff dff_A_5eKDupkb3_0(.dout(w_dff_A_L0tboVp27_0),.din(w_dff_A_5eKDupkb3_0),.clk(gclk));
	jdff dff_A_L0tboVp27_0(.dout(w_dff_A_0aDugl4U4_0),.din(w_dff_A_L0tboVp27_0),.clk(gclk));
	jdff dff_A_0aDugl4U4_0(.dout(w_dff_A_qlUrri2u5_0),.din(w_dff_A_0aDugl4U4_0),.clk(gclk));
	jdff dff_A_qlUrri2u5_0(.dout(w_dff_A_ZrAVO2IU7_0),.din(w_dff_A_qlUrri2u5_0),.clk(gclk));
	jdff dff_A_ZrAVO2IU7_0(.dout(w_dff_A_4LD1nPrA5_0),.din(w_dff_A_ZrAVO2IU7_0),.clk(gclk));
	jdff dff_A_4LD1nPrA5_0(.dout(w_dff_A_MlgP1iY98_0),.din(w_dff_A_4LD1nPrA5_0),.clk(gclk));
	jdff dff_A_MlgP1iY98_0(.dout(w_dff_A_fvKcz1on6_0),.din(w_dff_A_MlgP1iY98_0),.clk(gclk));
	jdff dff_A_fvKcz1on6_0(.dout(w_dff_A_9iFHD7mZ9_0),.din(w_dff_A_fvKcz1on6_0),.clk(gclk));
	jdff dff_A_9iFHD7mZ9_0(.dout(w_dff_A_W9gYILl37_0),.din(w_dff_A_9iFHD7mZ9_0),.clk(gclk));
	jdff dff_A_W9gYILl37_0(.dout(w_dff_A_kviH5ehM8_0),.din(w_dff_A_W9gYILl37_0),.clk(gclk));
	jdff dff_A_kviH5ehM8_0(.dout(w_dff_A_kp2e2jZt0_0),.din(w_dff_A_kviH5ehM8_0),.clk(gclk));
	jdff dff_A_kp2e2jZt0_0(.dout(w_dff_A_MC5uGbXK2_0),.din(w_dff_A_kp2e2jZt0_0),.clk(gclk));
	jdff dff_A_MC5uGbXK2_0(.dout(G278),.din(w_dff_A_MC5uGbXK2_0),.clk(gclk));
	jdff dff_A_62FaZpmK6_2(.dout(w_dff_A_g69OA2CD8_0),.din(w_dff_A_62FaZpmK6_2),.clk(gclk));
	jdff dff_A_g69OA2CD8_0(.dout(w_dff_A_QuiRtBwq1_0),.din(w_dff_A_g69OA2CD8_0),.clk(gclk));
	jdff dff_A_QuiRtBwq1_0(.dout(w_dff_A_TlIzQDNG4_0),.din(w_dff_A_QuiRtBwq1_0),.clk(gclk));
	jdff dff_A_TlIzQDNG4_0(.dout(w_dff_A_Z7FljO0j8_0),.din(w_dff_A_TlIzQDNG4_0),.clk(gclk));
	jdff dff_A_Z7FljO0j8_0(.dout(w_dff_A_1jhYuCaq9_0),.din(w_dff_A_Z7FljO0j8_0),.clk(gclk));
	jdff dff_A_1jhYuCaq9_0(.dout(w_dff_A_a04esJpm8_0),.din(w_dff_A_1jhYuCaq9_0),.clk(gclk));
	jdff dff_A_a04esJpm8_0(.dout(w_dff_A_wf0HrOHu5_0),.din(w_dff_A_a04esJpm8_0),.clk(gclk));
	jdff dff_A_wf0HrOHu5_0(.dout(w_dff_A_p28Vpuyy9_0),.din(w_dff_A_wf0HrOHu5_0),.clk(gclk));
	jdff dff_A_p28Vpuyy9_0(.dout(w_dff_A_aRu70x720_0),.din(w_dff_A_p28Vpuyy9_0),.clk(gclk));
	jdff dff_A_aRu70x720_0(.dout(w_dff_A_Y0bK5UJ64_0),.din(w_dff_A_aRu70x720_0),.clk(gclk));
	jdff dff_A_Y0bK5UJ64_0(.dout(w_dff_A_LFn6pe3n6_0),.din(w_dff_A_Y0bK5UJ64_0),.clk(gclk));
	jdff dff_A_LFn6pe3n6_0(.dout(w_dff_A_sutW7no98_0),.din(w_dff_A_LFn6pe3n6_0),.clk(gclk));
	jdff dff_A_sutW7no98_0(.dout(w_dff_A_lmvuzq220_0),.din(w_dff_A_sutW7no98_0),.clk(gclk));
	jdff dff_A_lmvuzq220_0(.dout(w_dff_A_KCalkvOR0_0),.din(w_dff_A_lmvuzq220_0),.clk(gclk));
	jdff dff_A_KCalkvOR0_0(.dout(w_dff_A_Tmn7GQBH2_0),.din(w_dff_A_KCalkvOR0_0),.clk(gclk));
	jdff dff_A_Tmn7GQBH2_0(.dout(w_dff_A_BvtVsQ6g7_0),.din(w_dff_A_Tmn7GQBH2_0),.clk(gclk));
	jdff dff_A_BvtVsQ6g7_0(.dout(w_dff_A_hWK0YZrx1_0),.din(w_dff_A_BvtVsQ6g7_0),.clk(gclk));
	jdff dff_A_hWK0YZrx1_0(.dout(w_dff_A_xOLgtix93_0),.din(w_dff_A_hWK0YZrx1_0),.clk(gclk));
	jdff dff_A_xOLgtix93_0(.dout(w_dff_A_EkoUja323_0),.din(w_dff_A_xOLgtix93_0),.clk(gclk));
	jdff dff_A_EkoUja323_0(.dout(w_dff_A_hZjZiFLp0_0),.din(w_dff_A_EkoUja323_0),.clk(gclk));
	jdff dff_A_hZjZiFLp0_0(.dout(w_dff_A_rccexe282_0),.din(w_dff_A_hZjZiFLp0_0),.clk(gclk));
	jdff dff_A_rccexe282_0(.dout(w_dff_A_tSTR4kib9_0),.din(w_dff_A_rccexe282_0),.clk(gclk));
	jdff dff_A_tSTR4kib9_0(.dout(w_dff_A_taBGw0sO5_0),.din(w_dff_A_tSTR4kib9_0),.clk(gclk));
	jdff dff_A_taBGw0sO5_0(.dout(w_dff_A_LFuVQOqR2_0),.din(w_dff_A_taBGw0sO5_0),.clk(gclk));
	jdff dff_A_LFuVQOqR2_0(.dout(w_dff_A_99dDVmuY5_0),.din(w_dff_A_LFuVQOqR2_0),.clk(gclk));
	jdff dff_A_99dDVmuY5_0(.dout(w_dff_A_cUEa9D5Z8_0),.din(w_dff_A_99dDVmuY5_0),.clk(gclk));
	jdff dff_A_cUEa9D5Z8_0(.dout(w_dff_A_46SttGKm0_0),.din(w_dff_A_cUEa9D5Z8_0),.clk(gclk));
	jdff dff_A_46SttGKm0_0(.dout(w_dff_A_38FWKvTq4_0),.din(w_dff_A_46SttGKm0_0),.clk(gclk));
	jdff dff_A_38FWKvTq4_0(.dout(w_dff_A_XYDVWFAH6_0),.din(w_dff_A_38FWKvTq4_0),.clk(gclk));
	jdff dff_A_XYDVWFAH6_0(.dout(w_dff_A_scyCPkrx4_0),.din(w_dff_A_XYDVWFAH6_0),.clk(gclk));
	jdff dff_A_scyCPkrx4_0(.dout(w_dff_A_Wiugym454_0),.din(w_dff_A_scyCPkrx4_0),.clk(gclk));
	jdff dff_A_Wiugym454_0(.dout(w_dff_A_fDL61mJj8_0),.din(w_dff_A_Wiugym454_0),.clk(gclk));
	jdff dff_A_fDL61mJj8_0(.dout(G373),.din(w_dff_A_fDL61mJj8_0),.clk(gclk));
	jdff dff_A_ajNjXzv73_2(.dout(w_dff_A_TT4aLrxh8_0),.din(w_dff_A_ajNjXzv73_2),.clk(gclk));
	jdff dff_A_TT4aLrxh8_0(.dout(w_dff_A_b0mGOHEG0_0),.din(w_dff_A_TT4aLrxh8_0),.clk(gclk));
	jdff dff_A_b0mGOHEG0_0(.dout(w_dff_A_OnzrlcE83_0),.din(w_dff_A_b0mGOHEG0_0),.clk(gclk));
	jdff dff_A_OnzrlcE83_0(.dout(w_dff_A_Ni1LBTDx6_0),.din(w_dff_A_OnzrlcE83_0),.clk(gclk));
	jdff dff_A_Ni1LBTDx6_0(.dout(w_dff_A_51H5h98E4_0),.din(w_dff_A_Ni1LBTDx6_0),.clk(gclk));
	jdff dff_A_51H5h98E4_0(.dout(w_dff_A_IQtwMLvQ3_0),.din(w_dff_A_51H5h98E4_0),.clk(gclk));
	jdff dff_A_IQtwMLvQ3_0(.dout(w_dff_A_AT6yNBzT9_0),.din(w_dff_A_IQtwMLvQ3_0),.clk(gclk));
	jdff dff_A_AT6yNBzT9_0(.dout(w_dff_A_YHG8H1Bh1_0),.din(w_dff_A_AT6yNBzT9_0),.clk(gclk));
	jdff dff_A_YHG8H1Bh1_0(.dout(w_dff_A_3hIjCyoX8_0),.din(w_dff_A_YHG8H1Bh1_0),.clk(gclk));
	jdff dff_A_3hIjCyoX8_0(.dout(w_dff_A_AVEnn40H0_0),.din(w_dff_A_3hIjCyoX8_0),.clk(gclk));
	jdff dff_A_AVEnn40H0_0(.dout(G258),.din(w_dff_A_AVEnn40H0_0),.clk(gclk));
	jdff dff_A_Q0KcgJhF3_2(.dout(w_dff_A_KOl0W78C0_0),.din(w_dff_A_Q0KcgJhF3_2),.clk(gclk));
	jdff dff_A_KOl0W78C0_0(.dout(w_dff_A_Z3KaIGIt9_0),.din(w_dff_A_KOl0W78C0_0),.clk(gclk));
	jdff dff_A_Z3KaIGIt9_0(.dout(w_dff_A_kh0fWH8s9_0),.din(w_dff_A_Z3KaIGIt9_0),.clk(gclk));
	jdff dff_A_kh0fWH8s9_0(.dout(w_dff_A_RIu0V3s05_0),.din(w_dff_A_kh0fWH8s9_0),.clk(gclk));
	jdff dff_A_RIu0V3s05_0(.dout(w_dff_A_L2FBgBar5_0),.din(w_dff_A_RIu0V3s05_0),.clk(gclk));
	jdff dff_A_L2FBgBar5_0(.dout(w_dff_A_os08S9Zl1_0),.din(w_dff_A_L2FBgBar5_0),.clk(gclk));
	jdff dff_A_os08S9Zl1_0(.dout(w_dff_A_s9YsBpMv2_0),.din(w_dff_A_os08S9Zl1_0),.clk(gclk));
	jdff dff_A_s9YsBpMv2_0(.dout(w_dff_A_nrhjltUI8_0),.din(w_dff_A_s9YsBpMv2_0),.clk(gclk));
	jdff dff_A_nrhjltUI8_0(.dout(w_dff_A_ZpScyhoT6_0),.din(w_dff_A_nrhjltUI8_0),.clk(gclk));
	jdff dff_A_ZpScyhoT6_0(.dout(w_dff_A_Mdo2LnXM0_0),.din(w_dff_A_ZpScyhoT6_0),.clk(gclk));
	jdff dff_A_Mdo2LnXM0_0(.dout(G264),.din(w_dff_A_Mdo2LnXM0_0),.clk(gclk));
	jdff dff_A_x51Q2GgN5_2(.dout(w_dff_A_QXfTuB9g2_0),.din(w_dff_A_x51Q2GgN5_2),.clk(gclk));
	jdff dff_A_QXfTuB9g2_0(.dout(w_dff_A_8AmfZoAq5_0),.din(w_dff_A_QXfTuB9g2_0),.clk(gclk));
	jdff dff_A_8AmfZoAq5_0(.dout(w_dff_A_IbzWtfJ57_0),.din(w_dff_A_8AmfZoAq5_0),.clk(gclk));
	jdff dff_A_IbzWtfJ57_0(.dout(w_dff_A_nQDqItJ52_0),.din(w_dff_A_IbzWtfJ57_0),.clk(gclk));
	jdff dff_A_nQDqItJ52_0(.dout(w_dff_A_1A2juYv22_0),.din(w_dff_A_nQDqItJ52_0),.clk(gclk));
	jdff dff_A_1A2juYv22_0(.dout(w_dff_A_7kVhfNGW5_0),.din(w_dff_A_1A2juYv22_0),.clk(gclk));
	jdff dff_A_7kVhfNGW5_0(.dout(w_dff_A_4FGNoSC30_0),.din(w_dff_A_7kVhfNGW5_0),.clk(gclk));
	jdff dff_A_4FGNoSC30_0(.dout(w_dff_A_XsqEqve71_0),.din(w_dff_A_4FGNoSC30_0),.clk(gclk));
	jdff dff_A_XsqEqve71_0(.dout(w_dff_A_6XKQXWdV0_0),.din(w_dff_A_XsqEqve71_0),.clk(gclk));
	jdff dff_A_6XKQXWdV0_0(.dout(w_dff_A_axiQnByq7_0),.din(w_dff_A_6XKQXWdV0_0),.clk(gclk));
	jdff dff_A_axiQnByq7_0(.dout(w_dff_A_1zmDcDJv6_0),.din(w_dff_A_axiQnByq7_0),.clk(gclk));
	jdff dff_A_1zmDcDJv6_0(.dout(w_dff_A_2JzmCsOe5_0),.din(w_dff_A_1zmDcDJv6_0),.clk(gclk));
	jdff dff_A_2JzmCsOe5_0(.dout(w_dff_A_m5nnqRn43_0),.din(w_dff_A_2JzmCsOe5_0),.clk(gclk));
	jdff dff_A_m5nnqRn43_0(.dout(w_dff_A_bZxY0xT66_0),.din(w_dff_A_m5nnqRn43_0),.clk(gclk));
	jdff dff_A_bZxY0xT66_0(.dout(w_dff_A_HtTAx8rO5_0),.din(w_dff_A_bZxY0xT66_0),.clk(gclk));
	jdff dff_A_HtTAx8rO5_0(.dout(w_dff_A_PobgbFdN5_0),.din(w_dff_A_HtTAx8rO5_0),.clk(gclk));
	jdff dff_A_PobgbFdN5_0(.dout(w_dff_A_1D3r5Csv8_0),.din(w_dff_A_PobgbFdN5_0),.clk(gclk));
	jdff dff_A_1D3r5Csv8_0(.dout(w_dff_A_zP4AdlFR4_0),.din(w_dff_A_1D3r5Csv8_0),.clk(gclk));
	jdff dff_A_zP4AdlFR4_0(.dout(w_dff_A_R5K8hbGX9_0),.din(w_dff_A_zP4AdlFR4_0),.clk(gclk));
	jdff dff_A_R5K8hbGX9_0(.dout(w_dff_A_YzPpywWF1_0),.din(w_dff_A_R5K8hbGX9_0),.clk(gclk));
	jdff dff_A_YzPpywWF1_0(.dout(w_dff_A_IqpCznLV2_0),.din(w_dff_A_YzPpywWF1_0),.clk(gclk));
	jdff dff_A_IqpCznLV2_0(.dout(w_dff_A_74miDqLV3_0),.din(w_dff_A_IqpCznLV2_0),.clk(gclk));
	jdff dff_A_74miDqLV3_0(.dout(w_dff_A_cnOsFqtO4_0),.din(w_dff_A_74miDqLV3_0),.clk(gclk));
	jdff dff_A_cnOsFqtO4_0(.dout(w_dff_A_w1xkvhtt2_0),.din(w_dff_A_cnOsFqtO4_0),.clk(gclk));
	jdff dff_A_w1xkvhtt2_0(.dout(G388),.din(w_dff_A_w1xkvhtt2_0),.clk(gclk));
	jdff dff_A_tgXJYLwI4_2(.dout(w_dff_A_e8n7Ar3U3_0),.din(w_dff_A_tgXJYLwI4_2),.clk(gclk));
	jdff dff_A_e8n7Ar3U3_0(.dout(w_dff_A_wv5xUv0L1_0),.din(w_dff_A_e8n7Ar3U3_0),.clk(gclk));
	jdff dff_A_wv5xUv0L1_0(.dout(w_dff_A_shkJdoO66_0),.din(w_dff_A_wv5xUv0L1_0),.clk(gclk));
	jdff dff_A_shkJdoO66_0(.dout(w_dff_A_lDZ4pdgI4_0),.din(w_dff_A_shkJdoO66_0),.clk(gclk));
	jdff dff_A_lDZ4pdgI4_0(.dout(w_dff_A_e8Lf7LST4_0),.din(w_dff_A_lDZ4pdgI4_0),.clk(gclk));
	jdff dff_A_e8Lf7LST4_0(.dout(w_dff_A_TTlPoZiz7_0),.din(w_dff_A_e8Lf7LST4_0),.clk(gclk));
	jdff dff_A_TTlPoZiz7_0(.dout(w_dff_A_8DBmWNwx2_0),.din(w_dff_A_TTlPoZiz7_0),.clk(gclk));
	jdff dff_A_8DBmWNwx2_0(.dout(w_dff_A_QYoWCk942_0),.din(w_dff_A_8DBmWNwx2_0),.clk(gclk));
	jdff dff_A_QYoWCk942_0(.dout(w_dff_A_qwXBWzUf1_0),.din(w_dff_A_QYoWCk942_0),.clk(gclk));
	jdff dff_A_qwXBWzUf1_0(.dout(w_dff_A_J92Njuev3_0),.din(w_dff_A_qwXBWzUf1_0),.clk(gclk));
	jdff dff_A_J92Njuev3_0(.dout(w_dff_A_lF18xUBi2_0),.din(w_dff_A_J92Njuev3_0),.clk(gclk));
	jdff dff_A_lF18xUBi2_0(.dout(w_dff_A_PbYKugJO5_0),.din(w_dff_A_lF18xUBi2_0),.clk(gclk));
	jdff dff_A_PbYKugJO5_0(.dout(w_dff_A_MFIzeAoe9_0),.din(w_dff_A_PbYKugJO5_0),.clk(gclk));
	jdff dff_A_MFIzeAoe9_0(.dout(w_dff_A_zTlAwahR5_0),.din(w_dff_A_MFIzeAoe9_0),.clk(gclk));
	jdff dff_A_zTlAwahR5_0(.dout(w_dff_A_Cjn9rNU64_0),.din(w_dff_A_zTlAwahR5_0),.clk(gclk));
	jdff dff_A_Cjn9rNU64_0(.dout(w_dff_A_WR4UX0mG1_0),.din(w_dff_A_Cjn9rNU64_0),.clk(gclk));
	jdff dff_A_WR4UX0mG1_0(.dout(w_dff_A_SjN8FEkV4_0),.din(w_dff_A_WR4UX0mG1_0),.clk(gclk));
	jdff dff_A_SjN8FEkV4_0(.dout(w_dff_A_nVanINLU6_0),.din(w_dff_A_SjN8FEkV4_0),.clk(gclk));
	jdff dff_A_nVanINLU6_0(.dout(w_dff_A_KdBdRfhE9_0),.din(w_dff_A_nVanINLU6_0),.clk(gclk));
	jdff dff_A_KdBdRfhE9_0(.dout(w_dff_A_64vzetlD5_0),.din(w_dff_A_KdBdRfhE9_0),.clk(gclk));
	jdff dff_A_64vzetlD5_0(.dout(w_dff_A_KB6jdD1o0_0),.din(w_dff_A_64vzetlD5_0),.clk(gclk));
	jdff dff_A_KB6jdD1o0_0(.dout(w_dff_A_gyCzG5ON0_0),.din(w_dff_A_KB6jdD1o0_0),.clk(gclk));
	jdff dff_A_gyCzG5ON0_0(.dout(w_dff_A_Vn7EchJy1_0),.din(w_dff_A_gyCzG5ON0_0),.clk(gclk));
	jdff dff_A_Vn7EchJy1_0(.dout(w_dff_A_AZGuGxhX2_0),.din(w_dff_A_Vn7EchJy1_0),.clk(gclk));
	jdff dff_A_AZGuGxhX2_0(.dout(w_dff_A_4NLTdJkF2_0),.din(w_dff_A_AZGuGxhX2_0),.clk(gclk));
	jdff dff_A_4NLTdJkF2_0(.dout(w_dff_A_zOyK1N2d6_0),.din(w_dff_A_4NLTdJkF2_0),.clk(gclk));
	jdff dff_A_zOyK1N2d6_0(.dout(G391),.din(w_dff_A_zOyK1N2d6_0),.clk(gclk));
	jdff dff_A_hkO5sPZ89_2(.dout(w_dff_A_hDf1sSif9_0),.din(w_dff_A_hkO5sPZ89_2),.clk(gclk));
	jdff dff_A_hDf1sSif9_0(.dout(w_dff_A_FKu6O3aV5_0),.din(w_dff_A_hDf1sSif9_0),.clk(gclk));
	jdff dff_A_FKu6O3aV5_0(.dout(w_dff_A_rcWQz1U65_0),.din(w_dff_A_FKu6O3aV5_0),.clk(gclk));
	jdff dff_A_rcWQz1U65_0(.dout(w_dff_A_uFpE2Po36_0),.din(w_dff_A_rcWQz1U65_0),.clk(gclk));
	jdff dff_A_uFpE2Po36_0(.dout(w_dff_A_keeOhkK75_0),.din(w_dff_A_uFpE2Po36_0),.clk(gclk));
	jdff dff_A_keeOhkK75_0(.dout(w_dff_A_MsShcQ7S4_0),.din(w_dff_A_keeOhkK75_0),.clk(gclk));
	jdff dff_A_MsShcQ7S4_0(.dout(w_dff_A_oNjxtp9A8_0),.din(w_dff_A_MsShcQ7S4_0),.clk(gclk));
	jdff dff_A_oNjxtp9A8_0(.dout(w_dff_A_rC0muEOt1_0),.din(w_dff_A_oNjxtp9A8_0),.clk(gclk));
	jdff dff_A_rC0muEOt1_0(.dout(w_dff_A_erigIFGs7_0),.din(w_dff_A_rC0muEOt1_0),.clk(gclk));
	jdff dff_A_erigIFGs7_0(.dout(w_dff_A_8NSbKSdI9_0),.din(w_dff_A_erigIFGs7_0),.clk(gclk));
	jdff dff_A_8NSbKSdI9_0(.dout(w_dff_A_IR4XtSOk8_0),.din(w_dff_A_8NSbKSdI9_0),.clk(gclk));
	jdff dff_A_IR4XtSOk8_0(.dout(w_dff_A_y9o18sIB9_0),.din(w_dff_A_IR4XtSOk8_0),.clk(gclk));
	jdff dff_A_y9o18sIB9_0(.dout(w_dff_A_TEolZjW42_0),.din(w_dff_A_y9o18sIB9_0),.clk(gclk));
	jdff dff_A_TEolZjW42_0(.dout(w_dff_A_DqLLjM5I8_0),.din(w_dff_A_TEolZjW42_0),.clk(gclk));
	jdff dff_A_DqLLjM5I8_0(.dout(w_dff_A_EIhcovon5_0),.din(w_dff_A_DqLLjM5I8_0),.clk(gclk));
	jdff dff_A_EIhcovon5_0(.dout(w_dff_A_XqDFxfmS0_0),.din(w_dff_A_EIhcovon5_0),.clk(gclk));
	jdff dff_A_XqDFxfmS0_0(.dout(w_dff_A_fxpMamxY8_0),.din(w_dff_A_XqDFxfmS0_0),.clk(gclk));
	jdff dff_A_fxpMamxY8_0(.dout(w_dff_A_2lMCaGUg2_0),.din(w_dff_A_fxpMamxY8_0),.clk(gclk));
	jdff dff_A_2lMCaGUg2_0(.dout(w_dff_A_B7BVzTId6_0),.din(w_dff_A_2lMCaGUg2_0),.clk(gclk));
	jdff dff_A_B7BVzTId6_0(.dout(w_dff_A_9Hiq8nFQ8_0),.din(w_dff_A_B7BVzTId6_0),.clk(gclk));
	jdff dff_A_9Hiq8nFQ8_0(.dout(w_dff_A_M2FgQ2rq9_0),.din(w_dff_A_9Hiq8nFQ8_0),.clk(gclk));
	jdff dff_A_M2FgQ2rq9_0(.dout(w_dff_A_dEMzwWWl4_0),.din(w_dff_A_M2FgQ2rq9_0),.clk(gclk));
	jdff dff_A_dEMzwWWl4_0(.dout(w_dff_A_G2oBSjtg8_0),.din(w_dff_A_dEMzwWWl4_0),.clk(gclk));
	jdff dff_A_G2oBSjtg8_0(.dout(w_dff_A_8LK18O1Z3_0),.din(w_dff_A_G2oBSjtg8_0),.clk(gclk));
	jdff dff_A_8LK18O1Z3_0(.dout(w_dff_A_LQJK2jlo1_0),.din(w_dff_A_8LK18O1Z3_0),.clk(gclk));
	jdff dff_A_LQJK2jlo1_0(.dout(w_dff_A_MA2zVwB88_0),.din(w_dff_A_LQJK2jlo1_0),.clk(gclk));
	jdff dff_A_MA2zVwB88_0(.dout(w_dff_A_4vkxo6Gj6_0),.din(w_dff_A_MA2zVwB88_0),.clk(gclk));
	jdff dff_A_4vkxo6Gj6_0(.dout(w_dff_A_8RB6P5rK6_0),.din(w_dff_A_4vkxo6Gj6_0),.clk(gclk));
	jdff dff_A_8RB6P5rK6_0(.dout(w_dff_A_aT2yF8k26_0),.din(w_dff_A_8RB6P5rK6_0),.clk(gclk));
	jdff dff_A_aT2yF8k26_0(.dout(G394),.din(w_dff_A_aT2yF8k26_0),.clk(gclk));
	jdff dff_A_pvUyVpXg5_2(.dout(w_dff_A_aQnNbj4A1_0),.din(w_dff_A_pvUyVpXg5_2),.clk(gclk));
	jdff dff_A_aQnNbj4A1_0(.dout(w_dff_A_GM2XjGwi6_0),.din(w_dff_A_aQnNbj4A1_0),.clk(gclk));
	jdff dff_A_GM2XjGwi6_0(.dout(w_dff_A_afYCStxr6_0),.din(w_dff_A_GM2XjGwi6_0),.clk(gclk));
	jdff dff_A_afYCStxr6_0(.dout(w_dff_A_ArzSCmgO4_0),.din(w_dff_A_afYCStxr6_0),.clk(gclk));
	jdff dff_A_ArzSCmgO4_0(.dout(w_dff_A_ANBeOubi5_0),.din(w_dff_A_ArzSCmgO4_0),.clk(gclk));
	jdff dff_A_ANBeOubi5_0(.dout(w_dff_A_PirPFoVG9_0),.din(w_dff_A_ANBeOubi5_0),.clk(gclk));
	jdff dff_A_PirPFoVG9_0(.dout(w_dff_A_6Km1af7F4_0),.din(w_dff_A_PirPFoVG9_0),.clk(gclk));
	jdff dff_A_6Km1af7F4_0(.dout(w_dff_A_1AOz8bgR5_0),.din(w_dff_A_6Km1af7F4_0),.clk(gclk));
	jdff dff_A_1AOz8bgR5_0(.dout(w_dff_A_TQyB4yGi6_0),.din(w_dff_A_1AOz8bgR5_0),.clk(gclk));
	jdff dff_A_TQyB4yGi6_0(.dout(w_dff_A_JPi4u3Gg9_0),.din(w_dff_A_TQyB4yGi6_0),.clk(gclk));
	jdff dff_A_JPi4u3Gg9_0(.dout(w_dff_A_XgAjAylE0_0),.din(w_dff_A_JPi4u3Gg9_0),.clk(gclk));
	jdff dff_A_XgAjAylE0_0(.dout(w_dff_A_R8HW4Iw66_0),.din(w_dff_A_XgAjAylE0_0),.clk(gclk));
	jdff dff_A_R8HW4Iw66_0(.dout(w_dff_A_AMDfN9IF8_0),.din(w_dff_A_R8HW4Iw66_0),.clk(gclk));
	jdff dff_A_AMDfN9IF8_0(.dout(w_dff_A_bG1X534F1_0),.din(w_dff_A_AMDfN9IF8_0),.clk(gclk));
	jdff dff_A_bG1X534F1_0(.dout(w_dff_A_Olh0tCaK3_0),.din(w_dff_A_bG1X534F1_0),.clk(gclk));
	jdff dff_A_Olh0tCaK3_0(.dout(w_dff_A_ICOjzVrE7_0),.din(w_dff_A_Olh0tCaK3_0),.clk(gclk));
	jdff dff_A_ICOjzVrE7_0(.dout(w_dff_A_V4d4Pfi78_0),.din(w_dff_A_ICOjzVrE7_0),.clk(gclk));
	jdff dff_A_V4d4Pfi78_0(.dout(w_dff_A_U9Mlowu36_0),.din(w_dff_A_V4d4Pfi78_0),.clk(gclk));
	jdff dff_A_U9Mlowu36_0(.dout(w_dff_A_o7ACEmcQ1_0),.din(w_dff_A_U9Mlowu36_0),.clk(gclk));
	jdff dff_A_o7ACEmcQ1_0(.dout(w_dff_A_ByUSFJiO5_0),.din(w_dff_A_o7ACEmcQ1_0),.clk(gclk));
	jdff dff_A_ByUSFJiO5_0(.dout(w_dff_A_cEuF0Rzi9_0),.din(w_dff_A_ByUSFJiO5_0),.clk(gclk));
	jdff dff_A_cEuF0Rzi9_0(.dout(w_dff_A_9957mxCD8_0),.din(w_dff_A_cEuF0Rzi9_0),.clk(gclk));
	jdff dff_A_9957mxCD8_0(.dout(w_dff_A_HFWFTiPj0_0),.din(w_dff_A_9957mxCD8_0),.clk(gclk));
	jdff dff_A_HFWFTiPj0_0(.dout(w_dff_A_HlwiP6gc5_0),.din(w_dff_A_HFWFTiPj0_0),.clk(gclk));
	jdff dff_A_HlwiP6gc5_0(.dout(w_dff_A_5oN3giQS6_0),.din(w_dff_A_HlwiP6gc5_0),.clk(gclk));
	jdff dff_A_5oN3giQS6_0(.dout(w_dff_A_K0kl6G7I1_0),.din(w_dff_A_5oN3giQS6_0),.clk(gclk));
	jdff dff_A_K0kl6G7I1_0(.dout(w_dff_A_Y37qaQCu8_0),.din(w_dff_A_K0kl6G7I1_0),.clk(gclk));
	jdff dff_A_Y37qaQCu8_0(.dout(w_dff_A_GWYdknZy7_0),.din(w_dff_A_Y37qaQCu8_0),.clk(gclk));
	jdff dff_A_GWYdknZy7_0(.dout(w_dff_A_CoNVsJtZ1_0),.din(w_dff_A_GWYdknZy7_0),.clk(gclk));
	jdff dff_A_CoNVsJtZ1_0(.dout(w_dff_A_663F91Cz0_0),.din(w_dff_A_CoNVsJtZ1_0),.clk(gclk));
	jdff dff_A_663F91Cz0_0(.dout(G397),.din(w_dff_A_663F91Cz0_0),.clk(gclk));
	jdff dff_A_GuechTS56_2(.dout(w_dff_A_DreT6W6u5_0),.din(w_dff_A_GuechTS56_2),.clk(gclk));
	jdff dff_A_DreT6W6u5_0(.dout(w_dff_A_YOm0inDL0_0),.din(w_dff_A_DreT6W6u5_0),.clk(gclk));
	jdff dff_A_YOm0inDL0_0(.dout(w_dff_A_e4jPZs2m6_0),.din(w_dff_A_YOm0inDL0_0),.clk(gclk));
	jdff dff_A_e4jPZs2m6_0(.dout(w_dff_A_Vr572Rtv1_0),.din(w_dff_A_e4jPZs2m6_0),.clk(gclk));
	jdff dff_A_Vr572Rtv1_0(.dout(w_dff_A_DOUAVlbY7_0),.din(w_dff_A_Vr572Rtv1_0),.clk(gclk));
	jdff dff_A_DOUAVlbY7_0(.dout(w_dff_A_FcKAJZuq1_0),.din(w_dff_A_DOUAVlbY7_0),.clk(gclk));
	jdff dff_A_FcKAJZuq1_0(.dout(w_dff_A_fJ3zIYMN2_0),.din(w_dff_A_FcKAJZuq1_0),.clk(gclk));
	jdff dff_A_fJ3zIYMN2_0(.dout(w_dff_A_6S90kLS13_0),.din(w_dff_A_fJ3zIYMN2_0),.clk(gclk));
	jdff dff_A_6S90kLS13_0(.dout(w_dff_A_kdPz2qcZ8_0),.din(w_dff_A_6S90kLS13_0),.clk(gclk));
	jdff dff_A_kdPz2qcZ8_0(.dout(w_dff_A_Vm79z5F93_0),.din(w_dff_A_kdPz2qcZ8_0),.clk(gclk));
	jdff dff_A_Vm79z5F93_0(.dout(w_dff_A_AWdaB3Ec6_0),.din(w_dff_A_Vm79z5F93_0),.clk(gclk));
	jdff dff_A_AWdaB3Ec6_0(.dout(w_dff_A_zaIDG96W8_0),.din(w_dff_A_AWdaB3Ec6_0),.clk(gclk));
	jdff dff_A_zaIDG96W8_0(.dout(w_dff_A_gZJ7ln329_0),.din(w_dff_A_zaIDG96W8_0),.clk(gclk));
	jdff dff_A_gZJ7ln329_0(.dout(w_dff_A_KUkinsFk0_0),.din(w_dff_A_gZJ7ln329_0),.clk(gclk));
	jdff dff_A_KUkinsFk0_0(.dout(w_dff_A_Ype3lJny5_0),.din(w_dff_A_KUkinsFk0_0),.clk(gclk));
	jdff dff_A_Ype3lJny5_0(.dout(w_dff_A_C3XdZN2U6_0),.din(w_dff_A_Ype3lJny5_0),.clk(gclk));
	jdff dff_A_C3XdZN2U6_0(.dout(w_dff_A_Z9f3GqZY4_0),.din(w_dff_A_C3XdZN2U6_0),.clk(gclk));
	jdff dff_A_Z9f3GqZY4_0(.dout(w_dff_A_VhDx769O3_0),.din(w_dff_A_Z9f3GqZY4_0),.clk(gclk));
	jdff dff_A_VhDx769O3_0(.dout(w_dff_A_l23cfTzy2_0),.din(w_dff_A_VhDx769O3_0),.clk(gclk));
	jdff dff_A_l23cfTzy2_0(.dout(G376),.din(w_dff_A_l23cfTzy2_0),.clk(gclk));
	jdff dff_A_ZvFxzFFl6_2(.dout(w_dff_A_yl4c68K17_0),.din(w_dff_A_ZvFxzFFl6_2),.clk(gclk));
	jdff dff_A_yl4c68K17_0(.dout(w_dff_A_BWACLAwZ7_0),.din(w_dff_A_yl4c68K17_0),.clk(gclk));
	jdff dff_A_BWACLAwZ7_0(.dout(w_dff_A_pYW6OGzw3_0),.din(w_dff_A_BWACLAwZ7_0),.clk(gclk));
	jdff dff_A_pYW6OGzw3_0(.dout(w_dff_A_HByCGAtg4_0),.din(w_dff_A_pYW6OGzw3_0),.clk(gclk));
	jdff dff_A_HByCGAtg4_0(.dout(w_dff_A_7yPhfK087_0),.din(w_dff_A_HByCGAtg4_0),.clk(gclk));
	jdff dff_A_7yPhfK087_0(.dout(w_dff_A_nzCs7fQd0_0),.din(w_dff_A_7yPhfK087_0),.clk(gclk));
	jdff dff_A_nzCs7fQd0_0(.dout(w_dff_A_mM4BEOBM8_0),.din(w_dff_A_nzCs7fQd0_0),.clk(gclk));
	jdff dff_A_mM4BEOBM8_0(.dout(w_dff_A_vW1ke1cG7_0),.din(w_dff_A_mM4BEOBM8_0),.clk(gclk));
	jdff dff_A_vW1ke1cG7_0(.dout(w_dff_A_rGreo9cd6_0),.din(w_dff_A_vW1ke1cG7_0),.clk(gclk));
	jdff dff_A_rGreo9cd6_0(.dout(w_dff_A_eJJTBJwz2_0),.din(w_dff_A_rGreo9cd6_0),.clk(gclk));
	jdff dff_A_eJJTBJwz2_0(.dout(w_dff_A_6YfKyfQg2_0),.din(w_dff_A_eJJTBJwz2_0),.clk(gclk));
	jdff dff_A_6YfKyfQg2_0(.dout(w_dff_A_eMGdGFOn4_0),.din(w_dff_A_6YfKyfQg2_0),.clk(gclk));
	jdff dff_A_eMGdGFOn4_0(.dout(w_dff_A_x134uNko5_0),.din(w_dff_A_eMGdGFOn4_0),.clk(gclk));
	jdff dff_A_x134uNko5_0(.dout(w_dff_A_nU6I5wxd2_0),.din(w_dff_A_x134uNko5_0),.clk(gclk));
	jdff dff_A_nU6I5wxd2_0(.dout(w_dff_A_l6yd9qmU7_0),.din(w_dff_A_nU6I5wxd2_0),.clk(gclk));
	jdff dff_A_l6yd9qmU7_0(.dout(w_dff_A_EcGTPUBE1_0),.din(w_dff_A_l6yd9qmU7_0),.clk(gclk));
	jdff dff_A_EcGTPUBE1_0(.dout(w_dff_A_1kgivv1n3_0),.din(w_dff_A_EcGTPUBE1_0),.clk(gclk));
	jdff dff_A_1kgivv1n3_0(.dout(w_dff_A_H0wMBfXf4_0),.din(w_dff_A_1kgivv1n3_0),.clk(gclk));
	jdff dff_A_H0wMBfXf4_0(.dout(w_dff_A_dEMtNCfJ5_0),.din(w_dff_A_H0wMBfXf4_0),.clk(gclk));
	jdff dff_A_dEMtNCfJ5_0(.dout(w_dff_A_zKLkmPlr7_0),.din(w_dff_A_dEMtNCfJ5_0),.clk(gclk));
	jdff dff_A_zKLkmPlr7_0(.dout(w_dff_A_YqoFysBa9_0),.din(w_dff_A_zKLkmPlr7_0),.clk(gclk));
	jdff dff_A_YqoFysBa9_0(.dout(G379),.din(w_dff_A_YqoFysBa9_0),.clk(gclk));
	jdff dff_A_5w4VshfQ8_2(.dout(w_dff_A_q7n93WK18_0),.din(w_dff_A_5w4VshfQ8_2),.clk(gclk));
	jdff dff_A_q7n93WK18_0(.dout(w_dff_A_lvbsOgSD4_0),.din(w_dff_A_q7n93WK18_0),.clk(gclk));
	jdff dff_A_lvbsOgSD4_0(.dout(w_dff_A_wFHhGfu92_0),.din(w_dff_A_lvbsOgSD4_0),.clk(gclk));
	jdff dff_A_wFHhGfu92_0(.dout(w_dff_A_Tu5a0fAV7_0),.din(w_dff_A_wFHhGfu92_0),.clk(gclk));
	jdff dff_A_Tu5a0fAV7_0(.dout(w_dff_A_3St9h9bx2_0),.din(w_dff_A_Tu5a0fAV7_0),.clk(gclk));
	jdff dff_A_3St9h9bx2_0(.dout(w_dff_A_NyrB6F5Q5_0),.din(w_dff_A_3St9h9bx2_0),.clk(gclk));
	jdff dff_A_NyrB6F5Q5_0(.dout(w_dff_A_0f8N24lP9_0),.din(w_dff_A_NyrB6F5Q5_0),.clk(gclk));
	jdff dff_A_0f8N24lP9_0(.dout(w_dff_A_b621w5zO5_0),.din(w_dff_A_0f8N24lP9_0),.clk(gclk));
	jdff dff_A_b621w5zO5_0(.dout(w_dff_A_XRs9b6JG2_0),.din(w_dff_A_b621w5zO5_0),.clk(gclk));
	jdff dff_A_XRs9b6JG2_0(.dout(w_dff_A_TjQF7fUR9_0),.din(w_dff_A_XRs9b6JG2_0),.clk(gclk));
	jdff dff_A_TjQF7fUR9_0(.dout(w_dff_A_mY6ane3F4_0),.din(w_dff_A_TjQF7fUR9_0),.clk(gclk));
	jdff dff_A_mY6ane3F4_0(.dout(w_dff_A_fxNW82Go9_0),.din(w_dff_A_mY6ane3F4_0),.clk(gclk));
	jdff dff_A_fxNW82Go9_0(.dout(w_dff_A_DFuXy87B4_0),.din(w_dff_A_fxNW82Go9_0),.clk(gclk));
	jdff dff_A_DFuXy87B4_0(.dout(w_dff_A_O5b2Z5p05_0),.din(w_dff_A_DFuXy87B4_0),.clk(gclk));
	jdff dff_A_O5b2Z5p05_0(.dout(w_dff_A_VrUYWFm31_0),.din(w_dff_A_O5b2Z5p05_0),.clk(gclk));
	jdff dff_A_VrUYWFm31_0(.dout(w_dff_A_imV7IoPg4_0),.din(w_dff_A_VrUYWFm31_0),.clk(gclk));
	jdff dff_A_imV7IoPg4_0(.dout(w_dff_A_Wb9TkMDO0_0),.din(w_dff_A_imV7IoPg4_0),.clk(gclk));
	jdff dff_A_Wb9TkMDO0_0(.dout(w_dff_A_6Lsfjqr59_0),.din(w_dff_A_Wb9TkMDO0_0),.clk(gclk));
	jdff dff_A_6Lsfjqr59_0(.dout(w_dff_A_8wj6Wm7R1_0),.din(w_dff_A_6Lsfjqr59_0),.clk(gclk));
	jdff dff_A_8wj6Wm7R1_0(.dout(w_dff_A_vdQfoMTJ6_0),.din(w_dff_A_8wj6Wm7R1_0),.clk(gclk));
	jdff dff_A_vdQfoMTJ6_0(.dout(w_dff_A_kL0ot33z2_0),.din(w_dff_A_vdQfoMTJ6_0),.clk(gclk));
	jdff dff_A_kL0ot33z2_0(.dout(G382),.din(w_dff_A_kL0ot33z2_0),.clk(gclk));
	jdff dff_A_DUPrbXiE4_2(.dout(w_dff_A_2ivTuG0o4_0),.din(w_dff_A_DUPrbXiE4_2),.clk(gclk));
	jdff dff_A_2ivTuG0o4_0(.dout(w_dff_A_Quh7QA6X1_0),.din(w_dff_A_2ivTuG0o4_0),.clk(gclk));
	jdff dff_A_Quh7QA6X1_0(.dout(w_dff_A_4yJtbFSK1_0),.din(w_dff_A_Quh7QA6X1_0),.clk(gclk));
	jdff dff_A_4yJtbFSK1_0(.dout(w_dff_A_N5r2sCJW6_0),.din(w_dff_A_4yJtbFSK1_0),.clk(gclk));
	jdff dff_A_N5r2sCJW6_0(.dout(w_dff_A_41HNgVQJ9_0),.din(w_dff_A_N5r2sCJW6_0),.clk(gclk));
	jdff dff_A_41HNgVQJ9_0(.dout(w_dff_A_ZiYWAXPU8_0),.din(w_dff_A_41HNgVQJ9_0),.clk(gclk));
	jdff dff_A_ZiYWAXPU8_0(.dout(w_dff_A_khwVr4Ex7_0),.din(w_dff_A_ZiYWAXPU8_0),.clk(gclk));
	jdff dff_A_khwVr4Ex7_0(.dout(w_dff_A_B0hqfcLv2_0),.din(w_dff_A_khwVr4Ex7_0),.clk(gclk));
	jdff dff_A_B0hqfcLv2_0(.dout(w_dff_A_oNali3mg7_0),.din(w_dff_A_B0hqfcLv2_0),.clk(gclk));
	jdff dff_A_oNali3mg7_0(.dout(w_dff_A_DgZ3Dx7Y1_0),.din(w_dff_A_oNali3mg7_0),.clk(gclk));
	jdff dff_A_DgZ3Dx7Y1_0(.dout(w_dff_A_7KBxL5iM3_0),.din(w_dff_A_DgZ3Dx7Y1_0),.clk(gclk));
	jdff dff_A_7KBxL5iM3_0(.dout(w_dff_A_wm5El60a6_0),.din(w_dff_A_7KBxL5iM3_0),.clk(gclk));
	jdff dff_A_wm5El60a6_0(.dout(w_dff_A_EfTPYhTn4_0),.din(w_dff_A_wm5El60a6_0),.clk(gclk));
	jdff dff_A_EfTPYhTn4_0(.dout(w_dff_A_zxSMasvo1_0),.din(w_dff_A_EfTPYhTn4_0),.clk(gclk));
	jdff dff_A_zxSMasvo1_0(.dout(w_dff_A_hZVaN7bZ1_0),.din(w_dff_A_zxSMasvo1_0),.clk(gclk));
	jdff dff_A_hZVaN7bZ1_0(.dout(w_dff_A_ulTVmNjv0_0),.din(w_dff_A_hZVaN7bZ1_0),.clk(gclk));
	jdff dff_A_ulTVmNjv0_0(.dout(w_dff_A_ZhR5ERnX7_0),.din(w_dff_A_ulTVmNjv0_0),.clk(gclk));
	jdff dff_A_ZhR5ERnX7_0(.dout(w_dff_A_UiJ7KuGz5_0),.din(w_dff_A_ZhR5ERnX7_0),.clk(gclk));
	jdff dff_A_UiJ7KuGz5_0(.dout(w_dff_A_1LaUYo8R6_0),.din(w_dff_A_UiJ7KuGz5_0),.clk(gclk));
	jdff dff_A_1LaUYo8R6_0(.dout(w_dff_A_I61dxXyN6_0),.din(w_dff_A_1LaUYo8R6_0),.clk(gclk));
	jdff dff_A_I61dxXyN6_0(.dout(w_dff_A_mtaQzUXW4_0),.din(w_dff_A_I61dxXyN6_0),.clk(gclk));
	jdff dff_A_mtaQzUXW4_0(.dout(w_dff_A_lLR2aZWF8_0),.din(w_dff_A_mtaQzUXW4_0),.clk(gclk));
	jdff dff_A_lLR2aZWF8_0(.dout(w_dff_A_uEdtUAss8_0),.din(w_dff_A_lLR2aZWF8_0),.clk(gclk));
	jdff dff_A_uEdtUAss8_0(.dout(G385),.din(w_dff_A_uEdtUAss8_0),.clk(gclk));
	jdff dff_A_CNbvXIlX4_1(.dout(w_dff_A_8LJshTeN7_0),.din(w_dff_A_CNbvXIlX4_1),.clk(gclk));
	jdff dff_A_8LJshTeN7_0(.dout(w_dff_A_cmvwVrDb7_0),.din(w_dff_A_8LJshTeN7_0),.clk(gclk));
	jdff dff_A_cmvwVrDb7_0(.dout(w_dff_A_7D5mA9my9_0),.din(w_dff_A_cmvwVrDb7_0),.clk(gclk));
	jdff dff_A_7D5mA9my9_0(.dout(w_dff_A_C5C6CeiH3_0),.din(w_dff_A_7D5mA9my9_0),.clk(gclk));
	jdff dff_A_C5C6CeiH3_0(.dout(w_dff_A_vmR9uS2j2_0),.din(w_dff_A_C5C6CeiH3_0),.clk(gclk));
	jdff dff_A_vmR9uS2j2_0(.dout(w_dff_A_NRrrW3Nn8_0),.din(w_dff_A_vmR9uS2j2_0),.clk(gclk));
	jdff dff_A_NRrrW3Nn8_0(.dout(w_dff_A_Gixi2GFr1_0),.din(w_dff_A_NRrrW3Nn8_0),.clk(gclk));
	jdff dff_A_Gixi2GFr1_0(.dout(w_dff_A_BLTyQRrj2_0),.din(w_dff_A_Gixi2GFr1_0),.clk(gclk));
	jdff dff_A_BLTyQRrj2_0(.dout(w_dff_A_L4MvBRI58_0),.din(w_dff_A_BLTyQRrj2_0),.clk(gclk));
	jdff dff_A_L4MvBRI58_0(.dout(w_dff_A_NoZQupbt3_0),.din(w_dff_A_L4MvBRI58_0),.clk(gclk));
	jdff dff_A_NoZQupbt3_0(.dout(w_dff_A_WfXEtKLE8_0),.din(w_dff_A_NoZQupbt3_0),.clk(gclk));
	jdff dff_A_WfXEtKLE8_0(.dout(w_dff_A_rClWGEqo3_0),.din(w_dff_A_WfXEtKLE8_0),.clk(gclk));
	jdff dff_A_rClWGEqo3_0(.dout(w_dff_A_ZjEpd6U45_0),.din(w_dff_A_rClWGEqo3_0),.clk(gclk));
	jdff dff_A_ZjEpd6U45_0(.dout(w_dff_A_voZF0aPA0_0),.din(w_dff_A_ZjEpd6U45_0),.clk(gclk));
	jdff dff_A_voZF0aPA0_0(.dout(w_dff_A_MJm2m4Ol4_0),.din(w_dff_A_voZF0aPA0_0),.clk(gclk));
	jdff dff_A_MJm2m4Ol4_0(.dout(w_dff_A_IXPfjlOj1_0),.din(w_dff_A_MJm2m4Ol4_0),.clk(gclk));
	jdff dff_A_IXPfjlOj1_0(.dout(w_dff_A_bJTur37y6_0),.din(w_dff_A_IXPfjlOj1_0),.clk(gclk));
	jdff dff_A_bJTur37y6_0(.dout(w_dff_A_Gv9xqr5e8_0),.din(w_dff_A_bJTur37y6_0),.clk(gclk));
	jdff dff_A_Gv9xqr5e8_0(.dout(w_dff_A_T6kEokzt6_0),.din(w_dff_A_Gv9xqr5e8_0),.clk(gclk));
	jdff dff_A_T6kEokzt6_0(.dout(w_dff_A_Sj8e0U7L1_0),.din(w_dff_A_T6kEokzt6_0),.clk(gclk));
	jdff dff_A_Sj8e0U7L1_0(.dout(w_dff_A_bFkTP5Xb4_0),.din(w_dff_A_Sj8e0U7L1_0),.clk(gclk));
	jdff dff_A_bFkTP5Xb4_0(.dout(w_dff_A_EOVDFatY7_0),.din(w_dff_A_bFkTP5Xb4_0),.clk(gclk));
	jdff dff_A_EOVDFatY7_0(.dout(w_dff_A_lMf3jntd4_0),.din(w_dff_A_EOVDFatY7_0),.clk(gclk));
	jdff dff_A_lMf3jntd4_0(.dout(w_dff_A_JTfPbw8A4_0),.din(w_dff_A_lMf3jntd4_0),.clk(gclk));
	jdff dff_A_JTfPbw8A4_0(.dout(w_dff_A_w0Bp0l8X8_0),.din(w_dff_A_JTfPbw8A4_0),.clk(gclk));
	jdff dff_A_w0Bp0l8X8_0(.dout(w_dff_A_ZhHw2eDs6_0),.din(w_dff_A_w0Bp0l8X8_0),.clk(gclk));
	jdff dff_A_ZhHw2eDs6_0(.dout(w_dff_A_CbgiTCht4_0),.din(w_dff_A_ZhHw2eDs6_0),.clk(gclk));
	jdff dff_A_CbgiTCht4_0(.dout(G412),.din(w_dff_A_CbgiTCht4_0),.clk(gclk));
	jdff dff_A_UmDLHC9r2_1(.dout(w_dff_A_fpzQTFJ88_0),.din(w_dff_A_UmDLHC9r2_1),.clk(gclk));
	jdff dff_A_fpzQTFJ88_0(.dout(w_dff_A_apvPFEcu1_0),.din(w_dff_A_fpzQTFJ88_0),.clk(gclk));
	jdff dff_A_apvPFEcu1_0(.dout(w_dff_A_NKZ9uYqh1_0),.din(w_dff_A_apvPFEcu1_0),.clk(gclk));
	jdff dff_A_NKZ9uYqh1_0(.dout(w_dff_A_tb2fT9FA9_0),.din(w_dff_A_NKZ9uYqh1_0),.clk(gclk));
	jdff dff_A_tb2fT9FA9_0(.dout(w_dff_A_cS7YiuoZ3_0),.din(w_dff_A_tb2fT9FA9_0),.clk(gclk));
	jdff dff_A_cS7YiuoZ3_0(.dout(w_dff_A_2djp1TUH2_0),.din(w_dff_A_cS7YiuoZ3_0),.clk(gclk));
	jdff dff_A_2djp1TUH2_0(.dout(w_dff_A_54QTNkBY3_0),.din(w_dff_A_2djp1TUH2_0),.clk(gclk));
	jdff dff_A_54QTNkBY3_0(.dout(w_dff_A_PHxgHErl7_0),.din(w_dff_A_54QTNkBY3_0),.clk(gclk));
	jdff dff_A_PHxgHErl7_0(.dout(w_dff_A_TTVQ65Tf8_0),.din(w_dff_A_PHxgHErl7_0),.clk(gclk));
	jdff dff_A_TTVQ65Tf8_0(.dout(w_dff_A_6Tm1qKK22_0),.din(w_dff_A_TTVQ65Tf8_0),.clk(gclk));
	jdff dff_A_6Tm1qKK22_0(.dout(w_dff_A_gRYMJjOw4_0),.din(w_dff_A_6Tm1qKK22_0),.clk(gclk));
	jdff dff_A_gRYMJjOw4_0(.dout(w_dff_A_JhLcErlz3_0),.din(w_dff_A_gRYMJjOw4_0),.clk(gclk));
	jdff dff_A_JhLcErlz3_0(.dout(w_dff_A_S8VLBB1r3_0),.din(w_dff_A_JhLcErlz3_0),.clk(gclk));
	jdff dff_A_S8VLBB1r3_0(.dout(w_dff_A_1MEE1oU61_0),.din(w_dff_A_S8VLBB1r3_0),.clk(gclk));
	jdff dff_A_1MEE1oU61_0(.dout(w_dff_A_Xq4Wyqyy4_0),.din(w_dff_A_1MEE1oU61_0),.clk(gclk));
	jdff dff_A_Xq4Wyqyy4_0(.dout(w_dff_A_yue0ZhoI1_0),.din(w_dff_A_Xq4Wyqyy4_0),.clk(gclk));
	jdff dff_A_yue0ZhoI1_0(.dout(w_dff_A_eNDQTfor1_0),.din(w_dff_A_yue0ZhoI1_0),.clk(gclk));
	jdff dff_A_eNDQTfor1_0(.dout(w_dff_A_jACVARD91_0),.din(w_dff_A_eNDQTfor1_0),.clk(gclk));
	jdff dff_A_jACVARD91_0(.dout(w_dff_A_ZEp5Uszh1_0),.din(w_dff_A_jACVARD91_0),.clk(gclk));
	jdff dff_A_ZEp5Uszh1_0(.dout(w_dff_A_SseCrQIB5_0),.din(w_dff_A_ZEp5Uszh1_0),.clk(gclk));
	jdff dff_A_SseCrQIB5_0(.dout(w_dff_A_9lLQRbp46_0),.din(w_dff_A_SseCrQIB5_0),.clk(gclk));
	jdff dff_A_9lLQRbp46_0(.dout(w_dff_A_L5Jy556h1_0),.din(w_dff_A_9lLQRbp46_0),.clk(gclk));
	jdff dff_A_L5Jy556h1_0(.dout(w_dff_A_3nug4nro5_0),.din(w_dff_A_L5Jy556h1_0),.clk(gclk));
	jdff dff_A_3nug4nro5_0(.dout(w_dff_A_yRGTWnt00_0),.din(w_dff_A_3nug4nro5_0),.clk(gclk));
	jdff dff_A_yRGTWnt00_0(.dout(w_dff_A_lSvp8Sbu1_0),.din(w_dff_A_yRGTWnt00_0),.clk(gclk));
	jdff dff_A_lSvp8Sbu1_0(.dout(w_dff_A_udFZ3Dq62_0),.din(w_dff_A_lSvp8Sbu1_0),.clk(gclk));
	jdff dff_A_udFZ3Dq62_0(.dout(w_dff_A_BsUIBrL06_0),.din(w_dff_A_udFZ3Dq62_0),.clk(gclk));
	jdff dff_A_BsUIBrL06_0(.dout(w_dff_A_XdoZMduP1_0),.din(w_dff_A_BsUIBrL06_0),.clk(gclk));
	jdff dff_A_XdoZMduP1_0(.dout(w_dff_A_x2zyQsxn2_0),.din(w_dff_A_XdoZMduP1_0),.clk(gclk));
	jdff dff_A_x2zyQsxn2_0(.dout(G414),.din(w_dff_A_x2zyQsxn2_0),.clk(gclk));
	jdff dff_A_R88Dkp5e7_1(.dout(w_dff_A_PgfZ5iMz1_0),.din(w_dff_A_R88Dkp5e7_1),.clk(gclk));
	jdff dff_A_PgfZ5iMz1_0(.dout(w_dff_A_5ar995Zr9_0),.din(w_dff_A_PgfZ5iMz1_0),.clk(gclk));
	jdff dff_A_5ar995Zr9_0(.dout(w_dff_A_bvX4qXK23_0),.din(w_dff_A_5ar995Zr9_0),.clk(gclk));
	jdff dff_A_bvX4qXK23_0(.dout(w_dff_A_ygLL3ad08_0),.din(w_dff_A_bvX4qXK23_0),.clk(gclk));
	jdff dff_A_ygLL3ad08_0(.dout(w_dff_A_jKnj2jlE8_0),.din(w_dff_A_ygLL3ad08_0),.clk(gclk));
	jdff dff_A_jKnj2jlE8_0(.dout(w_dff_A_RtyD8z916_0),.din(w_dff_A_jKnj2jlE8_0),.clk(gclk));
	jdff dff_A_RtyD8z916_0(.dout(w_dff_A_fRKrrvAt0_0),.din(w_dff_A_RtyD8z916_0),.clk(gclk));
	jdff dff_A_fRKrrvAt0_0(.dout(w_dff_A_Z9UaPxn51_0),.din(w_dff_A_fRKrrvAt0_0),.clk(gclk));
	jdff dff_A_Z9UaPxn51_0(.dout(w_dff_A_nSMqXAOa3_0),.din(w_dff_A_Z9UaPxn51_0),.clk(gclk));
	jdff dff_A_nSMqXAOa3_0(.dout(w_dff_A_iYlIXvBp6_0),.din(w_dff_A_nSMqXAOa3_0),.clk(gclk));
	jdff dff_A_iYlIXvBp6_0(.dout(w_dff_A_OPtxso7F4_0),.din(w_dff_A_iYlIXvBp6_0),.clk(gclk));
	jdff dff_A_OPtxso7F4_0(.dout(w_dff_A_donPucLe5_0),.din(w_dff_A_OPtxso7F4_0),.clk(gclk));
	jdff dff_A_donPucLe5_0(.dout(w_dff_A_S39SYTDx8_0),.din(w_dff_A_donPucLe5_0),.clk(gclk));
	jdff dff_A_S39SYTDx8_0(.dout(w_dff_A_KTChpuad1_0),.din(w_dff_A_S39SYTDx8_0),.clk(gclk));
	jdff dff_A_KTChpuad1_0(.dout(w_dff_A_ElT9XbFR7_0),.din(w_dff_A_KTChpuad1_0),.clk(gclk));
	jdff dff_A_ElT9XbFR7_0(.dout(w_dff_A_5D3gpbdx6_0),.din(w_dff_A_ElT9XbFR7_0),.clk(gclk));
	jdff dff_A_5D3gpbdx6_0(.dout(w_dff_A_SUhHr1jl9_0),.din(w_dff_A_5D3gpbdx6_0),.clk(gclk));
	jdff dff_A_SUhHr1jl9_0(.dout(w_dff_A_rViJZvoT5_0),.din(w_dff_A_SUhHr1jl9_0),.clk(gclk));
	jdff dff_A_rViJZvoT5_0(.dout(w_dff_A_cSgCoskL8_0),.din(w_dff_A_rViJZvoT5_0),.clk(gclk));
	jdff dff_A_cSgCoskL8_0(.dout(w_dff_A_V478lIvK7_0),.din(w_dff_A_cSgCoskL8_0),.clk(gclk));
	jdff dff_A_V478lIvK7_0(.dout(w_dff_A_s8s7KUzL3_0),.din(w_dff_A_V478lIvK7_0),.clk(gclk));
	jdff dff_A_s8s7KUzL3_0(.dout(w_dff_A_imoyar1A6_0),.din(w_dff_A_s8s7KUzL3_0),.clk(gclk));
	jdff dff_A_imoyar1A6_0(.dout(w_dff_A_scCGR20z6_0),.din(w_dff_A_imoyar1A6_0),.clk(gclk));
	jdff dff_A_scCGR20z6_0(.dout(w_dff_A_VshQyyec1_0),.din(w_dff_A_scCGR20z6_0),.clk(gclk));
	jdff dff_A_VshQyyec1_0(.dout(w_dff_A_ZrAtgBOy7_0),.din(w_dff_A_VshQyyec1_0),.clk(gclk));
	jdff dff_A_ZrAtgBOy7_0(.dout(w_dff_A_iwnZEO5h9_0),.din(w_dff_A_ZrAtgBOy7_0),.clk(gclk));
	jdff dff_A_iwnZEO5h9_0(.dout(w_dff_A_VdZczkdE1_0),.din(w_dff_A_iwnZEO5h9_0),.clk(gclk));
	jdff dff_A_VdZczkdE1_0(.dout(w_dff_A_eEEDelEM6_0),.din(w_dff_A_VdZczkdE1_0),.clk(gclk));
	jdff dff_A_eEEDelEM6_0(.dout(G416),.din(w_dff_A_eEEDelEM6_0),.clk(gclk));
	jdff dff_A_5fdEYc6z9_2(.dout(w_dff_A_EORhwlQA5_0),.din(w_dff_A_5fdEYc6z9_2),.clk(gclk));
	jdff dff_A_EORhwlQA5_0(.dout(w_dff_A_BCtXgJXy4_0),.din(w_dff_A_EORhwlQA5_0),.clk(gclk));
	jdff dff_A_BCtXgJXy4_0(.dout(w_dff_A_HpSA6GNa2_0),.din(w_dff_A_BCtXgJXy4_0),.clk(gclk));
	jdff dff_A_HpSA6GNa2_0(.dout(w_dff_A_Z6W0c00I9_0),.din(w_dff_A_HpSA6GNa2_0),.clk(gclk));
	jdff dff_A_Z6W0c00I9_0(.dout(w_dff_A_iHS23Xyr0_0),.din(w_dff_A_Z6W0c00I9_0),.clk(gclk));
	jdff dff_A_iHS23Xyr0_0(.dout(w_dff_A_JTPkDerP5_0),.din(w_dff_A_iHS23Xyr0_0),.clk(gclk));
	jdff dff_A_JTPkDerP5_0(.dout(w_dff_A_vVBTWctA0_0),.din(w_dff_A_JTPkDerP5_0),.clk(gclk));
	jdff dff_A_vVBTWctA0_0(.dout(w_dff_A_CIEdHvQv7_0),.din(w_dff_A_vVBTWctA0_0),.clk(gclk));
	jdff dff_A_CIEdHvQv7_0(.dout(w_dff_A_7tpVCytZ9_0),.din(w_dff_A_CIEdHvQv7_0),.clk(gclk));
	jdff dff_A_7tpVCytZ9_0(.dout(w_dff_A_hO2CJKlI2_0),.din(w_dff_A_7tpVCytZ9_0),.clk(gclk));
	jdff dff_A_hO2CJKlI2_0(.dout(G249),.din(w_dff_A_hO2CJKlI2_0),.clk(gclk));
	jdff dff_A_3zfTOB0e0_2(.dout(w_dff_A_lSxQCspR5_0),.din(w_dff_A_3zfTOB0e0_2),.clk(gclk));
	jdff dff_A_lSxQCspR5_0(.dout(w_dff_A_X4Ne4JLj5_0),.din(w_dff_A_lSxQCspR5_0),.clk(gclk));
	jdff dff_A_X4Ne4JLj5_0(.dout(w_dff_A_1OHz36ns6_0),.din(w_dff_A_X4Ne4JLj5_0),.clk(gclk));
	jdff dff_A_1OHz36ns6_0(.dout(w_dff_A_WYSgW46M0_0),.din(w_dff_A_1OHz36ns6_0),.clk(gclk));
	jdff dff_A_WYSgW46M0_0(.dout(w_dff_A_z71eXQPj8_0),.din(w_dff_A_WYSgW46M0_0),.clk(gclk));
	jdff dff_A_z71eXQPj8_0(.dout(w_dff_A_6RbivZWz4_0),.din(w_dff_A_z71eXQPj8_0),.clk(gclk));
	jdff dff_A_6RbivZWz4_0(.dout(w_dff_A_4LaOOQ7W1_0),.din(w_dff_A_6RbivZWz4_0),.clk(gclk));
	jdff dff_A_4LaOOQ7W1_0(.dout(w_dff_A_FovQvqSJ1_0),.din(w_dff_A_4LaOOQ7W1_0),.clk(gclk));
	jdff dff_A_FovQvqSJ1_0(.dout(w_dff_A_fS9GxS7v6_0),.din(w_dff_A_FovQvqSJ1_0),.clk(gclk));
	jdff dff_A_fS9GxS7v6_0(.dout(w_dff_A_k5zg3SHu2_0),.din(w_dff_A_fS9GxS7v6_0),.clk(gclk));
	jdff dff_A_k5zg3SHu2_0(.dout(G295),.din(w_dff_A_k5zg3SHu2_0),.clk(gclk));
	jdff dff_A_fKN3Ov279_2(.dout(w_dff_A_kLygOFrb5_0),.din(w_dff_A_fKN3Ov279_2),.clk(gclk));
	jdff dff_A_kLygOFrb5_0(.dout(w_dff_A_A8k1YTxs7_0),.din(w_dff_A_kLygOFrb5_0),.clk(gclk));
	jdff dff_A_A8k1YTxs7_0(.dout(w_dff_A_fWYw82rE4_0),.din(w_dff_A_A8k1YTxs7_0),.clk(gclk));
	jdff dff_A_fWYw82rE4_0(.dout(G324),.din(w_dff_A_fWYw82rE4_0),.clk(gclk));
	jdff dff_A_0iaYpmVK7_1(.dout(w_dff_A_nd7AJyg36_0),.din(w_dff_A_0iaYpmVK7_1),.clk(gclk));
	jdff dff_A_nd7AJyg36_0(.dout(w_dff_A_f2JQRMEI9_0),.din(w_dff_A_nd7AJyg36_0),.clk(gclk));
	jdff dff_A_f2JQRMEI9_0(.dout(w_dff_A_9moGAJdc7_0),.din(w_dff_A_f2JQRMEI9_0),.clk(gclk));
	jdff dff_A_9moGAJdc7_0(.dout(w_dff_A_074rv2Fs0_0),.din(w_dff_A_9moGAJdc7_0),.clk(gclk));
	jdff dff_A_074rv2Fs0_0(.dout(w_dff_A_AfXj7ETA8_0),.din(w_dff_A_074rv2Fs0_0),.clk(gclk));
	jdff dff_A_AfXj7ETA8_0(.dout(w_dff_A_YekKFm1z6_0),.din(w_dff_A_AfXj7ETA8_0),.clk(gclk));
	jdff dff_A_YekKFm1z6_0(.dout(w_dff_A_kU9ikpeo2_0),.din(w_dff_A_YekKFm1z6_0),.clk(gclk));
	jdff dff_A_kU9ikpeo2_0(.dout(w_dff_A_zLDth2L44_0),.din(w_dff_A_kU9ikpeo2_0),.clk(gclk));
	jdff dff_A_zLDth2L44_0(.dout(w_dff_A_CrMRH2oI7_0),.din(w_dff_A_zLDth2L44_0),.clk(gclk));
	jdff dff_A_CrMRH2oI7_0(.dout(w_dff_A_lE2sFZxr7_0),.din(w_dff_A_CrMRH2oI7_0),.clk(gclk));
	jdff dff_A_lE2sFZxr7_0(.dout(w_dff_A_4b11MPkO2_0),.din(w_dff_A_lE2sFZxr7_0),.clk(gclk));
	jdff dff_A_4b11MPkO2_0(.dout(w_dff_A_AqDBN58x7_0),.din(w_dff_A_4b11MPkO2_0),.clk(gclk));
	jdff dff_A_AqDBN58x7_0(.dout(w_dff_A_055wRPif3_0),.din(w_dff_A_AqDBN58x7_0),.clk(gclk));
	jdff dff_A_055wRPif3_0(.dout(w_dff_A_RevDtGVB1_0),.din(w_dff_A_055wRPif3_0),.clk(gclk));
	jdff dff_A_RevDtGVB1_0(.dout(w_dff_A_4L3ylKuf4_0),.din(w_dff_A_RevDtGVB1_0),.clk(gclk));
	jdff dff_A_4L3ylKuf4_0(.dout(w_dff_A_mQpxvKvk7_0),.din(w_dff_A_4L3ylKuf4_0),.clk(gclk));
	jdff dff_A_mQpxvKvk7_0(.dout(w_dff_A_Na6gBKa89_0),.din(w_dff_A_mQpxvKvk7_0),.clk(gclk));
	jdff dff_A_Na6gBKa89_0(.dout(w_dff_A_xZ5XmhYy0_0),.din(w_dff_A_Na6gBKa89_0),.clk(gclk));
	jdff dff_A_xZ5XmhYy0_0(.dout(w_dff_A_N22YiHxz7_0),.din(w_dff_A_xZ5XmhYy0_0),.clk(gclk));
	jdff dff_A_N22YiHxz7_0(.dout(w_dff_A_8x1oYZfP3_0),.din(w_dff_A_N22YiHxz7_0),.clk(gclk));
	jdff dff_A_8x1oYZfP3_0(.dout(G252),.din(w_dff_A_8x1oYZfP3_0),.clk(gclk));
	jdff dff_A_BYw8wZjg9_2(.dout(w_dff_A_V6aVPXsc1_0),.din(w_dff_A_BYw8wZjg9_2),.clk(gclk));
	jdff dff_A_V6aVPXsc1_0(.dout(w_dff_A_Bd28jUTQ4_0),.din(w_dff_A_V6aVPXsc1_0),.clk(gclk));
	jdff dff_A_Bd28jUTQ4_0(.dout(w_dff_A_QMYkzvZA8_0),.din(w_dff_A_Bd28jUTQ4_0),.clk(gclk));
	jdff dff_A_QMYkzvZA8_0(.dout(w_dff_A_VLQlYb5f8_0),.din(w_dff_A_QMYkzvZA8_0),.clk(gclk));
	jdff dff_A_VLQlYb5f8_0(.dout(w_dff_A_xPeoULhC5_0),.din(w_dff_A_VLQlYb5f8_0),.clk(gclk));
	jdff dff_A_xPeoULhC5_0(.dout(G310),.din(w_dff_A_xPeoULhC5_0),.clk(gclk));
	jdff dff_A_3tjmx9Te0_2(.dout(w_dff_A_EtOCEjPl6_0),.din(w_dff_A_3tjmx9Te0_2),.clk(gclk));
	jdff dff_A_EtOCEjPl6_0(.dout(w_dff_A_Bd5eKFnI8_0),.din(w_dff_A_EtOCEjPl6_0),.clk(gclk));
	jdff dff_A_Bd5eKFnI8_0(.dout(w_dff_A_3N0DEjoK4_0),.din(w_dff_A_Bd5eKFnI8_0),.clk(gclk));
	jdff dff_A_3N0DEjoK4_0(.dout(w_dff_A_hygaRTBY6_0),.din(w_dff_A_3N0DEjoK4_0),.clk(gclk));
	jdff dff_A_hygaRTBY6_0(.dout(G313),.din(w_dff_A_hygaRTBY6_0),.clk(gclk));
	jdff dff_A_gZ1v9epB1_2(.dout(w_dff_A_D7ucvZLP8_0),.din(w_dff_A_gZ1v9epB1_2),.clk(gclk));
	jdff dff_A_D7ucvZLP8_0(.dout(w_dff_A_5bO1MY4L3_0),.din(w_dff_A_D7ucvZLP8_0),.clk(gclk));
	jdff dff_A_5bO1MY4L3_0(.dout(w_dff_A_dvDrvt444_0),.din(w_dff_A_5bO1MY4L3_0),.clk(gclk));
	jdff dff_A_dvDrvt444_0(.dout(w_dff_A_2FUZ899C1_0),.din(w_dff_A_dvDrvt444_0),.clk(gclk));
	jdff dff_A_2FUZ899C1_0(.dout(w_dff_A_XUGEsEnh5_0),.din(w_dff_A_2FUZ899C1_0),.clk(gclk));
	jdff dff_A_XUGEsEnh5_0(.dout(w_dff_A_DNmFV2Mc1_0),.din(w_dff_A_XUGEsEnh5_0),.clk(gclk));
	jdff dff_A_DNmFV2Mc1_0(.dout(w_dff_A_wP1tavFb2_0),.din(w_dff_A_DNmFV2Mc1_0),.clk(gclk));
	jdff dff_A_wP1tavFb2_0(.dout(w_dff_A_Tp7fuB0T8_0),.din(w_dff_A_wP1tavFb2_0),.clk(gclk));
	jdff dff_A_Tp7fuB0T8_0(.dout(G316),.din(w_dff_A_Tp7fuB0T8_0),.clk(gclk));
	jdff dff_A_F2Gv4zZ05_2(.dout(w_dff_A_gy11JA5I7_0),.din(w_dff_A_F2Gv4zZ05_2),.clk(gclk));
	jdff dff_A_gy11JA5I7_0(.dout(w_dff_A_s76ba72r2_0),.din(w_dff_A_gy11JA5I7_0),.clk(gclk));
	jdff dff_A_s76ba72r2_0(.dout(w_dff_A_ldh5CQJd0_0),.din(w_dff_A_s76ba72r2_0),.clk(gclk));
	jdff dff_A_ldh5CQJd0_0(.dout(w_dff_A_jwyxDsZy2_0),.din(w_dff_A_ldh5CQJd0_0),.clk(gclk));
	jdff dff_A_jwyxDsZy2_0(.dout(w_dff_A_7rEevuaQ2_0),.din(w_dff_A_jwyxDsZy2_0),.clk(gclk));
	jdff dff_A_7rEevuaQ2_0(.dout(w_dff_A_ffhrifTG8_0),.din(w_dff_A_7rEevuaQ2_0),.clk(gclk));
	jdff dff_A_ffhrifTG8_0(.dout(w_dff_A_iu1Ysb078_0),.din(w_dff_A_ffhrifTG8_0),.clk(gclk));
	jdff dff_A_iu1Ysb078_0(.dout(w_dff_A_YhiS2eGY6_0),.din(w_dff_A_iu1Ysb078_0),.clk(gclk));
	jdff dff_A_YhiS2eGY6_0(.dout(G319),.din(w_dff_A_YhiS2eGY6_0),.clk(gclk));
	jdff dff_A_7obnZiGZ1_2(.dout(w_dff_A_FE5QoXE37_0),.din(w_dff_A_7obnZiGZ1_2),.clk(gclk));
	jdff dff_A_FE5QoXE37_0(.dout(G327),.din(w_dff_A_FE5QoXE37_0),.clk(gclk));
	jdff dff_A_UdtblJ0F2_2(.dout(w_dff_A_6NY2N59Y3_0),.din(w_dff_A_UdtblJ0F2_2),.clk(gclk));
	jdff dff_A_6NY2N59Y3_0(.dout(G330),.din(w_dff_A_6NY2N59Y3_0),.clk(gclk));
	jdff dff_A_PsLnarY76_2(.dout(w_dff_A_xYPcZIYe7_0),.din(w_dff_A_PsLnarY76_2),.clk(gclk));
	jdff dff_A_xYPcZIYe7_0(.dout(G336),.din(w_dff_A_xYPcZIYe7_0),.clk(gclk));
	jdff dff_A_YlBNGGZi2_2(.dout(w_dff_A_8nPXRQOf6_0),.din(w_dff_A_YlBNGGZi2_2),.clk(gclk));
	jdff dff_A_8nPXRQOf6_0(.dout(w_dff_A_exSyuo865_0),.din(w_dff_A_8nPXRQOf6_0),.clk(gclk));
	jdff dff_A_exSyuo865_0(.dout(w_dff_A_jtwMi6hO8_0),.din(w_dff_A_exSyuo865_0),.clk(gclk));
	jdff dff_A_jtwMi6hO8_0(.dout(w_dff_A_QR7dOgq43_0),.din(w_dff_A_jtwMi6hO8_0),.clk(gclk));
	jdff dff_A_QR7dOgq43_0(.dout(w_dff_A_Kk5KURfM1_0),.din(w_dff_A_QR7dOgq43_0),.clk(gclk));
	jdff dff_A_Kk5KURfM1_0(.dout(w_dff_A_crNFTGrv7_0),.din(w_dff_A_Kk5KURfM1_0),.clk(gclk));
	jdff dff_A_crNFTGrv7_0(.dout(w_dff_A_1BREmXEr6_0),.din(w_dff_A_crNFTGrv7_0),.clk(gclk));
	jdff dff_A_1BREmXEr6_0(.dout(w_dff_A_qJ50bqhN4_0),.din(w_dff_A_1BREmXEr6_0),.clk(gclk));
	jdff dff_A_qJ50bqhN4_0(.dout(w_dff_A_BjosxPRc4_0),.din(w_dff_A_qJ50bqhN4_0),.clk(gclk));
	jdff dff_A_BjosxPRc4_0(.dout(w_dff_A_4Ad49jj66_0),.din(w_dff_A_BjosxPRc4_0),.clk(gclk));
	jdff dff_A_4Ad49jj66_0(.dout(w_dff_A_8z8uGJbX4_0),.din(w_dff_A_4Ad49jj66_0),.clk(gclk));
	jdff dff_A_8z8uGJbX4_0(.dout(w_dff_A_1Glriinb3_0),.din(w_dff_A_8z8uGJbX4_0),.clk(gclk));
	jdff dff_A_1Glriinb3_0(.dout(w_dff_A_LC1YCvD15_0),.din(w_dff_A_1Glriinb3_0),.clk(gclk));
	jdff dff_A_LC1YCvD15_0(.dout(w_dff_A_gmEY2Ycu3_0),.din(w_dff_A_LC1YCvD15_0),.clk(gclk));
	jdff dff_A_gmEY2Ycu3_0(.dout(w_dff_A_wI6qLgtO3_0),.din(w_dff_A_gmEY2Ycu3_0),.clk(gclk));
	jdff dff_A_wI6qLgtO3_0(.dout(w_dff_A_p0wxxp632_0),.din(w_dff_A_wI6qLgtO3_0),.clk(gclk));
	jdff dff_A_p0wxxp632_0(.dout(w_dff_A_9nSFi8Nl6_0),.din(w_dff_A_p0wxxp632_0),.clk(gclk));
	jdff dff_A_9nSFi8Nl6_0(.dout(w_dff_A_CD2gKyok9_0),.din(w_dff_A_9nSFi8Nl6_0),.clk(gclk));
	jdff dff_A_CD2gKyok9_0(.dout(w_dff_A_mzpcjNh41_0),.din(w_dff_A_CD2gKyok9_0),.clk(gclk));
	jdff dff_A_mzpcjNh41_0(.dout(w_dff_A_MXOMLNmN4_0),.din(w_dff_A_mzpcjNh41_0),.clk(gclk));
	jdff dff_A_MXOMLNmN4_0(.dout(w_dff_A_tXdazhKJ0_0),.din(w_dff_A_MXOMLNmN4_0),.clk(gclk));
	jdff dff_A_tXdazhKJ0_0(.dout(w_dff_A_gkBkkFd59_0),.din(w_dff_A_tXdazhKJ0_0),.clk(gclk));
	jdff dff_A_gkBkkFd59_0(.dout(w_dff_A_wdOZv0zc9_0),.din(w_dff_A_gkBkkFd59_0),.clk(gclk));
	jdff dff_A_wdOZv0zc9_0(.dout(w_dff_A_XcZolYWe6_0),.din(w_dff_A_wdOZv0zc9_0),.clk(gclk));
	jdff dff_A_XcZolYWe6_0(.dout(G418),.din(w_dff_A_XcZolYWe6_0),.clk(gclk));
	jdff dff_A_PSGSlOxf2_2(.dout(w_dff_A_yyOA2ltG6_0),.din(w_dff_A_PSGSlOxf2_2),.clk(gclk));
	jdff dff_A_yyOA2ltG6_0(.dout(w_dff_A_tgoJ9R3q8_0),.din(w_dff_A_yyOA2ltG6_0),.clk(gclk));
	jdff dff_A_tgoJ9R3q8_0(.dout(w_dff_A_nRmN2kCU9_0),.din(w_dff_A_tgoJ9R3q8_0),.clk(gclk));
	jdff dff_A_nRmN2kCU9_0(.dout(w_dff_A_kZHY9oCh1_0),.din(w_dff_A_nRmN2kCU9_0),.clk(gclk));
	jdff dff_A_kZHY9oCh1_0(.dout(w_dff_A_hZVgUNuc6_0),.din(w_dff_A_kZHY9oCh1_0),.clk(gclk));
	jdff dff_A_hZVgUNuc6_0(.dout(G298),.din(w_dff_A_hZVgUNuc6_0),.clk(gclk));
	jdff dff_A_FicGj5tX6_2(.dout(w_dff_A_VbWxeYIa1_0),.din(w_dff_A_FicGj5tX6_2),.clk(gclk));
	jdff dff_A_VbWxeYIa1_0(.dout(w_dff_A_2btqfOnt3_0),.din(w_dff_A_VbWxeYIa1_0),.clk(gclk));
	jdff dff_A_2btqfOnt3_0(.dout(w_dff_A_pY1t3G7j6_0),.din(w_dff_A_2btqfOnt3_0),.clk(gclk));
	jdff dff_A_pY1t3G7j6_0(.dout(w_dff_A_4TrwIiOk1_0),.din(w_dff_A_pY1t3G7j6_0),.clk(gclk));
	jdff dff_A_4TrwIiOk1_0(.dout(w_dff_A_I9bGlMmw8_0),.din(w_dff_A_4TrwIiOk1_0),.clk(gclk));
	jdff dff_A_I9bGlMmw8_0(.dout(G301),.din(w_dff_A_I9bGlMmw8_0),.clk(gclk));
	jdff dff_A_IHdVYUXP2_2(.dout(w_dff_A_n66B77iq3_0),.din(w_dff_A_IHdVYUXP2_2),.clk(gclk));
	jdff dff_A_n66B77iq3_0(.dout(w_dff_A_h3tYHDBo0_0),.din(w_dff_A_n66B77iq3_0),.clk(gclk));
	jdff dff_A_h3tYHDBo0_0(.dout(w_dff_A_uCdvdXR31_0),.din(w_dff_A_h3tYHDBo0_0),.clk(gclk));
	jdff dff_A_uCdvdXR31_0(.dout(w_dff_A_ThQPVUZP2_0),.din(w_dff_A_uCdvdXR31_0),.clk(gclk));
	jdff dff_A_ThQPVUZP2_0(.dout(w_dff_A_LPZCpK0T7_0),.din(w_dff_A_ThQPVUZP2_0),.clk(gclk));
	jdff dff_A_LPZCpK0T7_0(.dout(G304),.din(w_dff_A_LPZCpK0T7_0),.clk(gclk));
	jdff dff_A_aKlzg0Oe8_2(.dout(w_dff_A_XKCHa7yq9_0),.din(w_dff_A_aKlzg0Oe8_2),.clk(gclk));
	jdff dff_A_XKCHa7yq9_0(.dout(w_dff_A_9lGyOzaR7_0),.din(w_dff_A_XKCHa7yq9_0),.clk(gclk));
	jdff dff_A_9lGyOzaR7_0(.dout(w_dff_A_hbCd1HdE8_0),.din(w_dff_A_9lGyOzaR7_0),.clk(gclk));
	jdff dff_A_hbCd1HdE8_0(.dout(w_dff_A_yh5GrPfm0_0),.din(w_dff_A_hbCd1HdE8_0),.clk(gclk));
	jdff dff_A_yh5GrPfm0_0(.dout(w_dff_A_2uPZWpXo8_0),.din(w_dff_A_yh5GrPfm0_0),.clk(gclk));
	jdff dff_A_2uPZWpXo8_0(.dout(w_dff_A_LKzkoi9k2_0),.din(w_dff_A_2uPZWpXo8_0),.clk(gclk));
	jdff dff_A_LKzkoi9k2_0(.dout(w_dff_A_DgiL5ows8_0),.din(w_dff_A_LKzkoi9k2_0),.clk(gclk));
	jdff dff_A_DgiL5ows8_0(.dout(G307),.din(w_dff_A_DgiL5ows8_0),.clk(gclk));
	jdff dff_A_6BxXv4053_2(.dout(w_dff_A_T7FLFExf7_0),.din(w_dff_A_6BxXv4053_2),.clk(gclk));
	jdff dff_A_T7FLFExf7_0(.dout(w_dff_A_gxXrxuWL9_0),.din(w_dff_A_T7FLFExf7_0),.clk(gclk));
	jdff dff_A_gxXrxuWL9_0(.dout(w_dff_A_CUaJcXwy6_0),.din(w_dff_A_gxXrxuWL9_0),.clk(gclk));
	jdff dff_A_CUaJcXwy6_0(.dout(w_dff_A_rj3gX9H63_0),.din(w_dff_A_CUaJcXwy6_0),.clk(gclk));
	jdff dff_A_rj3gX9H63_0(.dout(w_dff_A_LR5uCdEj9_0),.din(w_dff_A_rj3gX9H63_0),.clk(gclk));
	jdff dff_A_LR5uCdEj9_0(.dout(w_dff_A_stHxCVM24_0),.din(w_dff_A_LR5uCdEj9_0),.clk(gclk));
	jdff dff_A_stHxCVM24_0(.dout(w_dff_A_KtULCR773_0),.din(w_dff_A_stHxCVM24_0),.clk(gclk));
	jdff dff_A_KtULCR773_0(.dout(w_dff_A_4IIErU4q7_0),.din(w_dff_A_KtULCR773_0),.clk(gclk));
	jdff dff_A_4IIErU4q7_0(.dout(w_dff_A_h8jLWbDh0_0),.din(w_dff_A_4IIErU4q7_0),.clk(gclk));
	jdff dff_A_h8jLWbDh0_0(.dout(w_dff_A_bFHILsoQ2_0),.din(w_dff_A_h8jLWbDh0_0),.clk(gclk));
	jdff dff_A_bFHILsoQ2_0(.dout(w_dff_A_uJlXdGCo4_0),.din(w_dff_A_bFHILsoQ2_0),.clk(gclk));
	jdff dff_A_uJlXdGCo4_0(.dout(w_dff_A_OA4O4XbX5_0),.din(w_dff_A_uJlXdGCo4_0),.clk(gclk));
	jdff dff_A_OA4O4XbX5_0(.dout(w_dff_A_mV9ksafz0_0),.din(w_dff_A_OA4O4XbX5_0),.clk(gclk));
	jdff dff_A_mV9ksafz0_0(.dout(w_dff_A_EPDQAWEU0_0),.din(w_dff_A_mV9ksafz0_0),.clk(gclk));
	jdff dff_A_EPDQAWEU0_0(.dout(w_dff_A_LQYxvjbz1_0),.din(w_dff_A_EPDQAWEU0_0),.clk(gclk));
	jdff dff_A_LQYxvjbz1_0(.dout(w_dff_A_O7a0owzQ8_0),.din(w_dff_A_LQYxvjbz1_0),.clk(gclk));
	jdff dff_A_O7a0owzQ8_0(.dout(w_dff_A_zp7is1dU1_0),.din(w_dff_A_O7a0owzQ8_0),.clk(gclk));
	jdff dff_A_zp7is1dU1_0(.dout(w_dff_A_evLEjbNM1_0),.din(w_dff_A_zp7is1dU1_0),.clk(gclk));
	jdff dff_A_evLEjbNM1_0(.dout(w_dff_A_V10yD3eU5_0),.din(w_dff_A_evLEjbNM1_0),.clk(gclk));
	jdff dff_A_V10yD3eU5_0(.dout(G344),.din(w_dff_A_V10yD3eU5_0),.clk(gclk));
	jdff dff_A_3gY2Zx692_2(.dout(w_dff_A_YEfry8FO8_0),.din(w_dff_A_3gY2Zx692_2),.clk(gclk));
	jdff dff_A_YEfry8FO8_0(.dout(G419),.din(w_dff_A_YEfry8FO8_0),.clk(gclk));
	jdff dff_A_aRxRy8Qx1_2(.dout(w_dff_A_M26jmssu0_0),.din(w_dff_A_aRxRy8Qx1_2),.clk(gclk));
	jdff dff_A_M26jmssu0_0(.dout(G471),.din(w_dff_A_M26jmssu0_0),.clk(gclk));
	jdff dff_A_pGz0TzDp7_2(.dout(w_dff_A_1Ze2UWsQ7_0),.din(w_dff_A_pGz0TzDp7_2),.clk(gclk));
	jdff dff_A_1Ze2UWsQ7_0(.dout(w_dff_A_tRBRv4QH4_0),.din(w_dff_A_1Ze2UWsQ7_0),.clk(gclk));
	jdff dff_A_tRBRv4QH4_0(.dout(w_dff_A_ArwEOjAo5_0),.din(w_dff_A_tRBRv4QH4_0),.clk(gclk));
	jdff dff_A_ArwEOjAo5_0(.dout(w_dff_A_K1LKraZY5_0),.din(w_dff_A_ArwEOjAo5_0),.clk(gclk));
	jdff dff_A_K1LKraZY5_0(.dout(w_dff_A_FnHRRYsr4_0),.din(w_dff_A_K1LKraZY5_0),.clk(gclk));
	jdff dff_A_FnHRRYsr4_0(.dout(w_dff_A_mGv8qgAs6_0),.din(w_dff_A_FnHRRYsr4_0),.clk(gclk));
	jdff dff_A_mGv8qgAs6_0(.dout(w_dff_A_1iNBjEtb2_0),.din(w_dff_A_mGv8qgAs6_0),.clk(gclk));
	jdff dff_A_1iNBjEtb2_0(.dout(w_dff_A_TZUlzPwn3_0),.din(w_dff_A_1iNBjEtb2_0),.clk(gclk));
	jdff dff_A_TZUlzPwn3_0(.dout(w_dff_A_0bS4kFjy0_0),.din(w_dff_A_TZUlzPwn3_0),.clk(gclk));
	jdff dff_A_0bS4kFjy0_0(.dout(w_dff_A_n88kCQf22_0),.din(w_dff_A_0bS4kFjy0_0),.clk(gclk));
	jdff dff_A_n88kCQf22_0(.dout(w_dff_A_rvnlIuCq0_0),.din(w_dff_A_n88kCQf22_0),.clk(gclk));
	jdff dff_A_rvnlIuCq0_0(.dout(w_dff_A_cbZfSeR66_0),.din(w_dff_A_rvnlIuCq0_0),.clk(gclk));
	jdff dff_A_cbZfSeR66_0(.dout(w_dff_A_4RSug8h85_0),.din(w_dff_A_cbZfSeR66_0),.clk(gclk));
	jdff dff_A_4RSug8h85_0(.dout(w_dff_A_Cuc6i5YH6_0),.din(w_dff_A_4RSug8h85_0),.clk(gclk));
	jdff dff_A_Cuc6i5YH6_0(.dout(w_dff_A_bC7cKcKa8_0),.din(w_dff_A_Cuc6i5YH6_0),.clk(gclk));
	jdff dff_A_bC7cKcKa8_0(.dout(w_dff_A_jXnLANAr8_0),.din(w_dff_A_bC7cKcKa8_0),.clk(gclk));
	jdff dff_A_jXnLANAr8_0(.dout(w_dff_A_f6XPnz5h0_0),.din(w_dff_A_jXnLANAr8_0),.clk(gclk));
	jdff dff_A_f6XPnz5h0_0(.dout(G359),.din(w_dff_A_f6XPnz5h0_0),.clk(gclk));
	jdff dff_A_39LSarcR8_2(.dout(w_dff_A_Or38g4ww3_0),.din(w_dff_A_39LSarcR8_2),.clk(gclk));
	jdff dff_A_Or38g4ww3_0(.dout(w_dff_A_frBTXjWn8_0),.din(w_dff_A_Or38g4ww3_0),.clk(gclk));
	jdff dff_A_frBTXjWn8_0(.dout(w_dff_A_wCld7PdR6_0),.din(w_dff_A_frBTXjWn8_0),.clk(gclk));
	jdff dff_A_wCld7PdR6_0(.dout(w_dff_A_Dk1DG5NK1_0),.din(w_dff_A_wCld7PdR6_0),.clk(gclk));
	jdff dff_A_Dk1DG5NK1_0(.dout(w_dff_A_NDIquvQZ6_0),.din(w_dff_A_Dk1DG5NK1_0),.clk(gclk));
	jdff dff_A_NDIquvQZ6_0(.dout(w_dff_A_lpfcRF452_0),.din(w_dff_A_NDIquvQZ6_0),.clk(gclk));
	jdff dff_A_lpfcRF452_0(.dout(w_dff_A_hTgLSKpD6_0),.din(w_dff_A_lpfcRF452_0),.clk(gclk));
	jdff dff_A_hTgLSKpD6_0(.dout(w_dff_A_eshq81ff7_0),.din(w_dff_A_hTgLSKpD6_0),.clk(gclk));
	jdff dff_A_eshq81ff7_0(.dout(w_dff_A_oeDvoZ4n8_0),.din(w_dff_A_eshq81ff7_0),.clk(gclk));
	jdff dff_A_oeDvoZ4n8_0(.dout(w_dff_A_KXMEQTyr6_0),.din(w_dff_A_oeDvoZ4n8_0),.clk(gclk));
	jdff dff_A_KXMEQTyr6_0(.dout(w_dff_A_XPTkbgQm6_0),.din(w_dff_A_KXMEQTyr6_0),.clk(gclk));
	jdff dff_A_XPTkbgQm6_0(.dout(w_dff_A_IJAOBrqm7_0),.din(w_dff_A_XPTkbgQm6_0),.clk(gclk));
	jdff dff_A_IJAOBrqm7_0(.dout(w_dff_A_E1DccclB9_0),.din(w_dff_A_IJAOBrqm7_0),.clk(gclk));
	jdff dff_A_E1DccclB9_0(.dout(w_dff_A_R2ygSeKK7_0),.din(w_dff_A_E1DccclB9_0),.clk(gclk));
	jdff dff_A_R2ygSeKK7_0(.dout(w_dff_A_aQ9HZ5sN7_0),.din(w_dff_A_R2ygSeKK7_0),.clk(gclk));
	jdff dff_A_aQ9HZ5sN7_0(.dout(w_dff_A_uzccgCpY4_0),.din(w_dff_A_aQ9HZ5sN7_0),.clk(gclk));
	jdff dff_A_uzccgCpY4_0(.dout(w_dff_A_WEZgCqLO8_0),.din(w_dff_A_uzccgCpY4_0),.clk(gclk));
	jdff dff_A_WEZgCqLO8_0(.dout(G362),.din(w_dff_A_WEZgCqLO8_0),.clk(gclk));
	jdff dff_A_Ok6uAbWN4_2(.dout(w_dff_A_0ayCAdl21_0),.din(w_dff_A_Ok6uAbWN4_2),.clk(gclk));
	jdff dff_A_0ayCAdl21_0(.dout(w_dff_A_Hai4Bxo74_0),.din(w_dff_A_0ayCAdl21_0),.clk(gclk));
	jdff dff_A_Hai4Bxo74_0(.dout(w_dff_A_fUvfw16W8_0),.din(w_dff_A_Hai4Bxo74_0),.clk(gclk));
	jdff dff_A_fUvfw16W8_0(.dout(w_dff_A_cWyOtGep6_0),.din(w_dff_A_fUvfw16W8_0),.clk(gclk));
	jdff dff_A_cWyOtGep6_0(.dout(w_dff_A_IHHwLxq40_0),.din(w_dff_A_cWyOtGep6_0),.clk(gclk));
	jdff dff_A_IHHwLxq40_0(.dout(w_dff_A_hrMgtwa86_0),.din(w_dff_A_IHHwLxq40_0),.clk(gclk));
	jdff dff_A_hrMgtwa86_0(.dout(w_dff_A_F4nXchMr5_0),.din(w_dff_A_hrMgtwa86_0),.clk(gclk));
	jdff dff_A_F4nXchMr5_0(.dout(w_dff_A_kZcCp9ng2_0),.din(w_dff_A_F4nXchMr5_0),.clk(gclk));
	jdff dff_A_kZcCp9ng2_0(.dout(w_dff_A_l4l0kOFP9_0),.din(w_dff_A_kZcCp9ng2_0),.clk(gclk));
	jdff dff_A_l4l0kOFP9_0(.dout(w_dff_A_9vqlPN4g2_0),.din(w_dff_A_l4l0kOFP9_0),.clk(gclk));
	jdff dff_A_9vqlPN4g2_0(.dout(w_dff_A_GLPquVQM1_0),.din(w_dff_A_9vqlPN4g2_0),.clk(gclk));
	jdff dff_A_GLPquVQM1_0(.dout(w_dff_A_e8yGQNQJ4_0),.din(w_dff_A_GLPquVQM1_0),.clk(gclk));
	jdff dff_A_e8yGQNQJ4_0(.dout(w_dff_A_RqlPRQDE2_0),.din(w_dff_A_e8yGQNQJ4_0),.clk(gclk));
	jdff dff_A_RqlPRQDE2_0(.dout(w_dff_A_VBz0642q7_0),.din(w_dff_A_RqlPRQDE2_0),.clk(gclk));
	jdff dff_A_VBz0642q7_0(.dout(w_dff_A_1tUKpQca0_0),.din(w_dff_A_VBz0642q7_0),.clk(gclk));
	jdff dff_A_1tUKpQca0_0(.dout(w_dff_A_QUQ54itN9_0),.din(w_dff_A_1tUKpQca0_0),.clk(gclk));
	jdff dff_A_QUQ54itN9_0(.dout(w_dff_A_Bmbl6rZ65_0),.din(w_dff_A_QUQ54itN9_0),.clk(gclk));
	jdff dff_A_Bmbl6rZ65_0(.dout(G365),.din(w_dff_A_Bmbl6rZ65_0),.clk(gclk));
	jdff dff_A_N1mAsmmi2_2(.dout(w_dff_A_e86IiVHH3_0),.din(w_dff_A_N1mAsmmi2_2),.clk(gclk));
	jdff dff_A_e86IiVHH3_0(.dout(w_dff_A_M36832ah7_0),.din(w_dff_A_e86IiVHH3_0),.clk(gclk));
	jdff dff_A_M36832ah7_0(.dout(w_dff_A_e0Orb4lA6_0),.din(w_dff_A_M36832ah7_0),.clk(gclk));
	jdff dff_A_e0Orb4lA6_0(.dout(w_dff_A_5eBgw1Tk2_0),.din(w_dff_A_e0Orb4lA6_0),.clk(gclk));
	jdff dff_A_5eBgw1Tk2_0(.dout(w_dff_A_JcuY7N3g4_0),.din(w_dff_A_5eBgw1Tk2_0),.clk(gclk));
	jdff dff_A_JcuY7N3g4_0(.dout(w_dff_A_zPNojqUB6_0),.din(w_dff_A_JcuY7N3g4_0),.clk(gclk));
	jdff dff_A_zPNojqUB6_0(.dout(w_dff_A_BrEpKekj3_0),.din(w_dff_A_zPNojqUB6_0),.clk(gclk));
	jdff dff_A_BrEpKekj3_0(.dout(w_dff_A_encOh2s40_0),.din(w_dff_A_BrEpKekj3_0),.clk(gclk));
	jdff dff_A_encOh2s40_0(.dout(w_dff_A_9cJOMgqh0_0),.din(w_dff_A_encOh2s40_0),.clk(gclk));
	jdff dff_A_9cJOMgqh0_0(.dout(w_dff_A_fRd1r4RP4_0),.din(w_dff_A_9cJOMgqh0_0),.clk(gclk));
	jdff dff_A_fRd1r4RP4_0(.dout(w_dff_A_CZbadehM3_0),.din(w_dff_A_fRd1r4RP4_0),.clk(gclk));
	jdff dff_A_CZbadehM3_0(.dout(w_dff_A_lswNp0EP2_0),.din(w_dff_A_CZbadehM3_0),.clk(gclk));
	jdff dff_A_lswNp0EP2_0(.dout(w_dff_A_qlGniEvj2_0),.din(w_dff_A_lswNp0EP2_0),.clk(gclk));
	jdff dff_A_qlGniEvj2_0(.dout(w_dff_A_N007mEEt9_0),.din(w_dff_A_qlGniEvj2_0),.clk(gclk));
	jdff dff_A_N007mEEt9_0(.dout(w_dff_A_DS3zjS1V5_0),.din(w_dff_A_N007mEEt9_0),.clk(gclk));
	jdff dff_A_DS3zjS1V5_0(.dout(w_dff_A_b5ZoaKfv0_0),.din(w_dff_A_DS3zjS1V5_0),.clk(gclk));
	jdff dff_A_b5ZoaKfv0_0(.dout(w_dff_A_Z8oRwTuK9_0),.din(w_dff_A_b5ZoaKfv0_0),.clk(gclk));
	jdff dff_A_Z8oRwTuK9_0(.dout(G368),.din(w_dff_A_Z8oRwTuK9_0),.clk(gclk));
	jdff dff_A_HerJdIIO9_2(.dout(w_dff_A_Zw4k2O9c9_0),.din(w_dff_A_HerJdIIO9_2),.clk(gclk));
	jdff dff_A_Zw4k2O9c9_0(.dout(w_dff_A_ORQZ0sdf8_0),.din(w_dff_A_Zw4k2O9c9_0),.clk(gclk));
	jdff dff_A_ORQZ0sdf8_0(.dout(w_dff_A_T46XX8Qa8_0),.din(w_dff_A_ORQZ0sdf8_0),.clk(gclk));
	jdff dff_A_T46XX8Qa8_0(.dout(w_dff_A_erjosBMk0_0),.din(w_dff_A_T46XX8Qa8_0),.clk(gclk));
	jdff dff_A_erjosBMk0_0(.dout(w_dff_A_fuPWfSGP0_0),.din(w_dff_A_erjosBMk0_0),.clk(gclk));
	jdff dff_A_fuPWfSGP0_0(.dout(w_dff_A_YvaQSWAJ8_0),.din(w_dff_A_fuPWfSGP0_0),.clk(gclk));
	jdff dff_A_YvaQSWAJ8_0(.dout(w_dff_A_7bjsJIrq2_0),.din(w_dff_A_YvaQSWAJ8_0),.clk(gclk));
	jdff dff_A_7bjsJIrq2_0(.dout(w_dff_A_D9Te1xWZ6_0),.din(w_dff_A_7bjsJIrq2_0),.clk(gclk));
	jdff dff_A_D9Te1xWZ6_0(.dout(w_dff_A_PhUca8Jx0_0),.din(w_dff_A_D9Te1xWZ6_0),.clk(gclk));
	jdff dff_A_PhUca8Jx0_0(.dout(w_dff_A_aWMShC4i6_0),.din(w_dff_A_PhUca8Jx0_0),.clk(gclk));
	jdff dff_A_aWMShC4i6_0(.dout(w_dff_A_WbEsNmol1_0),.din(w_dff_A_aWMShC4i6_0),.clk(gclk));
	jdff dff_A_WbEsNmol1_0(.dout(w_dff_A_szg5BwvA8_0),.din(w_dff_A_WbEsNmol1_0),.clk(gclk));
	jdff dff_A_szg5BwvA8_0(.dout(G347),.din(w_dff_A_szg5BwvA8_0),.clk(gclk));
	jdff dff_A_cmrFAdAy7_2(.dout(w_dff_A_JJeTwaYA8_0),.din(w_dff_A_cmrFAdAy7_2),.clk(gclk));
	jdff dff_A_JJeTwaYA8_0(.dout(w_dff_A_dii8jI0N8_0),.din(w_dff_A_JJeTwaYA8_0),.clk(gclk));
	jdff dff_A_dii8jI0N8_0(.dout(w_dff_A_ubCvPUdn0_0),.din(w_dff_A_dii8jI0N8_0),.clk(gclk));
	jdff dff_A_ubCvPUdn0_0(.dout(w_dff_A_3LMAsPgj4_0),.din(w_dff_A_ubCvPUdn0_0),.clk(gclk));
	jdff dff_A_3LMAsPgj4_0(.dout(w_dff_A_6j41Zqs12_0),.din(w_dff_A_3LMAsPgj4_0),.clk(gclk));
	jdff dff_A_6j41Zqs12_0(.dout(w_dff_A_73sxFhUA2_0),.din(w_dff_A_6j41Zqs12_0),.clk(gclk));
	jdff dff_A_73sxFhUA2_0(.dout(w_dff_A_9b2rEQ9O6_0),.din(w_dff_A_73sxFhUA2_0),.clk(gclk));
	jdff dff_A_9b2rEQ9O6_0(.dout(w_dff_A_opntaJuZ7_0),.din(w_dff_A_9b2rEQ9O6_0),.clk(gclk));
	jdff dff_A_opntaJuZ7_0(.dout(w_dff_A_ftHqaEUe4_0),.din(w_dff_A_opntaJuZ7_0),.clk(gclk));
	jdff dff_A_ftHqaEUe4_0(.dout(w_dff_A_JTd57Y9V7_0),.din(w_dff_A_ftHqaEUe4_0),.clk(gclk));
	jdff dff_A_JTd57Y9V7_0(.dout(w_dff_A_fZnjr7TN2_0),.din(w_dff_A_JTd57Y9V7_0),.clk(gclk));
	jdff dff_A_fZnjr7TN2_0(.dout(w_dff_A_8MpDjeCt8_0),.din(w_dff_A_fZnjr7TN2_0),.clk(gclk));
	jdff dff_A_8MpDjeCt8_0(.dout(w_dff_A_7kOYqbgg5_0),.din(w_dff_A_8MpDjeCt8_0),.clk(gclk));
	jdff dff_A_7kOYqbgg5_0(.dout(G350),.din(w_dff_A_7kOYqbgg5_0),.clk(gclk));
	jdff dff_A_zYA4qFmc0_2(.dout(w_dff_A_xCaeHS7k4_0),.din(w_dff_A_zYA4qFmc0_2),.clk(gclk));
	jdff dff_A_xCaeHS7k4_0(.dout(w_dff_A_91RMdsVf8_0),.din(w_dff_A_xCaeHS7k4_0),.clk(gclk));
	jdff dff_A_91RMdsVf8_0(.dout(w_dff_A_buf0kbXX3_0),.din(w_dff_A_91RMdsVf8_0),.clk(gclk));
	jdff dff_A_buf0kbXX3_0(.dout(w_dff_A_kfjrNXJh5_0),.din(w_dff_A_buf0kbXX3_0),.clk(gclk));
	jdff dff_A_kfjrNXJh5_0(.dout(w_dff_A_BLuQR1Qx7_0),.din(w_dff_A_kfjrNXJh5_0),.clk(gclk));
	jdff dff_A_BLuQR1Qx7_0(.dout(w_dff_A_HYhVbmDM8_0),.din(w_dff_A_BLuQR1Qx7_0),.clk(gclk));
	jdff dff_A_HYhVbmDM8_0(.dout(w_dff_A_FkCRMnaE6_0),.din(w_dff_A_HYhVbmDM8_0),.clk(gclk));
	jdff dff_A_FkCRMnaE6_0(.dout(w_dff_A_uRo3uB4I6_0),.din(w_dff_A_FkCRMnaE6_0),.clk(gclk));
	jdff dff_A_uRo3uB4I6_0(.dout(w_dff_A_rdB7BPKt8_0),.din(w_dff_A_uRo3uB4I6_0),.clk(gclk));
	jdff dff_A_rdB7BPKt8_0(.dout(w_dff_A_UbmbXZi94_0),.din(w_dff_A_rdB7BPKt8_0),.clk(gclk));
	jdff dff_A_UbmbXZi94_0(.dout(w_dff_A_3Wdne82Z6_0),.din(w_dff_A_UbmbXZi94_0),.clk(gclk));
	jdff dff_A_3Wdne82Z6_0(.dout(w_dff_A_4roMcrxw9_0),.din(w_dff_A_3Wdne82Z6_0),.clk(gclk));
	jdff dff_A_4roMcrxw9_0(.dout(w_dff_A_8fCtJaLk4_0),.din(w_dff_A_4roMcrxw9_0),.clk(gclk));
	jdff dff_A_8fCtJaLk4_0(.dout(w_dff_A_KNA2aBHr1_0),.din(w_dff_A_8fCtJaLk4_0),.clk(gclk));
	jdff dff_A_KNA2aBHr1_0(.dout(w_dff_A_FNRnCz2S2_0),.din(w_dff_A_KNA2aBHr1_0),.clk(gclk));
	jdff dff_A_FNRnCz2S2_0(.dout(G353),.din(w_dff_A_FNRnCz2S2_0),.clk(gclk));
	jdff dff_A_IpwnXTLg0_2(.dout(w_dff_A_1KQy76900_0),.din(w_dff_A_IpwnXTLg0_2),.clk(gclk));
	jdff dff_A_1KQy76900_0(.dout(w_dff_A_NNJdX76P6_0),.din(w_dff_A_1KQy76900_0),.clk(gclk));
	jdff dff_A_NNJdX76P6_0(.dout(w_dff_A_LtTshqNf1_0),.din(w_dff_A_NNJdX76P6_0),.clk(gclk));
	jdff dff_A_LtTshqNf1_0(.dout(w_dff_A_2YNl0r4s9_0),.din(w_dff_A_LtTshqNf1_0),.clk(gclk));
	jdff dff_A_2YNl0r4s9_0(.dout(w_dff_A_HDpytnws8_0),.din(w_dff_A_2YNl0r4s9_0),.clk(gclk));
	jdff dff_A_HDpytnws8_0(.dout(w_dff_A_LEfRcKZu6_0),.din(w_dff_A_HDpytnws8_0),.clk(gclk));
	jdff dff_A_LEfRcKZu6_0(.dout(w_dff_A_kQQnB38u1_0),.din(w_dff_A_LEfRcKZu6_0),.clk(gclk));
	jdff dff_A_kQQnB38u1_0(.dout(w_dff_A_EfBYDn0W6_0),.din(w_dff_A_kQQnB38u1_0),.clk(gclk));
	jdff dff_A_EfBYDn0W6_0(.dout(w_dff_A_5rgiUtMz3_0),.din(w_dff_A_EfBYDn0W6_0),.clk(gclk));
	jdff dff_A_5rgiUtMz3_0(.dout(w_dff_A_bDmVCKah5_0),.din(w_dff_A_5rgiUtMz3_0),.clk(gclk));
	jdff dff_A_bDmVCKah5_0(.dout(w_dff_A_4UV6Aa7P7_0),.din(w_dff_A_bDmVCKah5_0),.clk(gclk));
	jdff dff_A_4UV6Aa7P7_0(.dout(w_dff_A_Kh6KxNtQ8_0),.din(w_dff_A_4UV6Aa7P7_0),.clk(gclk));
	jdff dff_A_Kh6KxNtQ8_0(.dout(w_dff_A_HhDMNim98_0),.din(w_dff_A_Kh6KxNtQ8_0),.clk(gclk));
	jdff dff_A_HhDMNim98_0(.dout(w_dff_A_UZQTJyrc7_0),.din(w_dff_A_HhDMNim98_0),.clk(gclk));
	jdff dff_A_UZQTJyrc7_0(.dout(w_dff_A_KGm3qQhT2_0),.din(w_dff_A_UZQTJyrc7_0),.clk(gclk));
	jdff dff_A_KGm3qQhT2_0(.dout(w_dff_A_CJf3sWow9_0),.din(w_dff_A_KGm3qQhT2_0),.clk(gclk));
	jdff dff_A_CJf3sWow9_0(.dout(w_dff_A_wIhJ1ELX0_0),.din(w_dff_A_CJf3sWow9_0),.clk(gclk));
	jdff dff_A_wIhJ1ELX0_0(.dout(G356),.din(w_dff_A_wIhJ1ELX0_0),.clk(gclk));
	jdff dff_A_DxbKqrBV1_2(.dout(w_dff_A_BsORI0N07_0),.din(w_dff_A_DxbKqrBV1_2),.clk(gclk));
	jdff dff_A_BsORI0N07_0(.dout(w_dff_A_RdRs7Zcf0_0),.din(w_dff_A_BsORI0N07_0),.clk(gclk));
	jdff dff_A_RdRs7Zcf0_0(.dout(w_dff_A_74jZjFLF0_0),.din(w_dff_A_RdRs7Zcf0_0),.clk(gclk));
	jdff dff_A_74jZjFLF0_0(.dout(w_dff_A_ZVxD6Kul4_0),.din(w_dff_A_74jZjFLF0_0),.clk(gclk));
	jdff dff_A_ZVxD6Kul4_0(.dout(w_dff_A_ihJQiTas3_0),.din(w_dff_A_ZVxD6Kul4_0),.clk(gclk));
	jdff dff_A_ihJQiTas3_0(.dout(G321),.din(w_dff_A_ihJQiTas3_0),.clk(gclk));
	jdff dff_A_SofaJqix2_2(.dout(G338),.din(w_dff_A_SofaJqix2_2),.clk(gclk));
	jdff dff_A_jT5X6nYq2_2(.dout(w_dff_A_T7aJU2ej9_0),.din(w_dff_A_jT5X6nYq2_2),.clk(gclk));
	jdff dff_A_T7aJU2ej9_0(.dout(w_dff_A_TfS78Cxh5_0),.din(w_dff_A_T7aJU2ej9_0),.clk(gclk));
	jdff dff_A_TfS78Cxh5_0(.dout(w_dff_A_52IkDmef8_0),.din(w_dff_A_TfS78Cxh5_0),.clk(gclk));
	jdff dff_A_52IkDmef8_0(.dout(w_dff_A_AHIN5y2A5_0),.din(w_dff_A_52IkDmef8_0),.clk(gclk));
	jdff dff_A_AHIN5y2A5_0(.dout(w_dff_A_87HskYOj1_0),.din(w_dff_A_AHIN5y2A5_0),.clk(gclk));
	jdff dff_A_87HskYOj1_0(.dout(w_dff_A_koxF0wgk2_0),.din(w_dff_A_87HskYOj1_0),.clk(gclk));
	jdff dff_A_koxF0wgk2_0(.dout(w_dff_A_JuP36eVp6_0),.din(w_dff_A_koxF0wgk2_0),.clk(gclk));
	jdff dff_A_JuP36eVp6_0(.dout(w_dff_A_pe6aqDYz1_0),.din(w_dff_A_JuP36eVp6_0),.clk(gclk));
	jdff dff_A_pe6aqDYz1_0(.dout(w_dff_A_dQ9g9yfS3_0),.din(w_dff_A_pe6aqDYz1_0),.clk(gclk));
	jdff dff_A_dQ9g9yfS3_0(.dout(w_dff_A_1jKm0Lkr1_0),.din(w_dff_A_dQ9g9yfS3_0),.clk(gclk));
	jdff dff_A_1jKm0Lkr1_0(.dout(w_dff_A_l9tCs6TB9_0),.din(w_dff_A_1jKm0Lkr1_0),.clk(gclk));
	jdff dff_A_l9tCs6TB9_0(.dout(w_dff_A_q059EdLg0_0),.din(w_dff_A_l9tCs6TB9_0),.clk(gclk));
	jdff dff_A_q059EdLg0_0(.dout(w_dff_A_3lC6Xhkx8_0),.din(w_dff_A_q059EdLg0_0),.clk(gclk));
	jdff dff_A_3lC6Xhkx8_0(.dout(w_dff_A_d6aRNQxc8_0),.din(w_dff_A_3lC6Xhkx8_0),.clk(gclk));
	jdff dff_A_d6aRNQxc8_0(.dout(w_dff_A_xxupOa4X3_0),.din(w_dff_A_d6aRNQxc8_0),.clk(gclk));
	jdff dff_A_xxupOa4X3_0(.dout(w_dff_A_U4owkrqr3_0),.din(w_dff_A_xxupOa4X3_0),.clk(gclk));
	jdff dff_A_U4owkrqr3_0(.dout(G370),.din(w_dff_A_U4owkrqr3_0),.clk(gclk));
	jdff dff_A_3UnuSp1X4_2(.dout(w_dff_A_K8LeKm9Q2_0),.din(w_dff_A_3UnuSp1X4_2),.clk(gclk));
	jdff dff_A_K8LeKm9Q2_0(.dout(w_dff_A_GC3ghFZB9_0),.din(w_dff_A_K8LeKm9Q2_0),.clk(gclk));
	jdff dff_A_GC3ghFZB9_0(.dout(w_dff_A_ESuSZBGM1_0),.din(w_dff_A_GC3ghFZB9_0),.clk(gclk));
	jdff dff_A_ESuSZBGM1_0(.dout(w_dff_A_uTtzCnn51_0),.din(w_dff_A_ESuSZBGM1_0),.clk(gclk));
	jdff dff_A_uTtzCnn51_0(.dout(w_dff_A_yEjBOBBS7_0),.din(w_dff_A_uTtzCnn51_0),.clk(gclk));
	jdff dff_A_yEjBOBBS7_0(.dout(w_dff_A_nbJmh1Ss8_0),.din(w_dff_A_yEjBOBBS7_0),.clk(gclk));
	jdff dff_A_nbJmh1Ss8_0(.dout(w_dff_A_ynywxUvS5_0),.din(w_dff_A_nbJmh1Ss8_0),.clk(gclk));
	jdff dff_A_ynywxUvS5_0(.dout(w_dff_A_NKEk5aAE6_0),.din(w_dff_A_ynywxUvS5_0),.clk(gclk));
	jdff dff_A_NKEk5aAE6_0(.dout(w_dff_A_TNlNeo4I2_0),.din(w_dff_A_NKEk5aAE6_0),.clk(gclk));
	jdff dff_A_TNlNeo4I2_0(.dout(w_dff_A_cZ4FOvJs2_0),.din(w_dff_A_TNlNeo4I2_0),.clk(gclk));
	jdff dff_A_cZ4FOvJs2_0(.dout(w_dff_A_IiVWy0E29_0),.din(w_dff_A_cZ4FOvJs2_0),.clk(gclk));
	jdff dff_A_IiVWy0E29_0(.dout(w_dff_A_3m5eUpMJ9_0),.din(w_dff_A_IiVWy0E29_0),.clk(gclk));
	jdff dff_A_3m5eUpMJ9_0(.dout(w_dff_A_8HyNi9Vr8_0),.din(w_dff_A_3m5eUpMJ9_0),.clk(gclk));
	jdff dff_A_8HyNi9Vr8_0(.dout(w_dff_A_QzauXjnj9_0),.din(w_dff_A_8HyNi9Vr8_0),.clk(gclk));
	jdff dff_A_QzauXjnj9_0(.dout(w_dff_A_QHuSf2Ia6_0),.din(w_dff_A_QzauXjnj9_0),.clk(gclk));
	jdff dff_A_QHuSf2Ia6_0(.dout(w_dff_A_zS6HEnMW4_0),.din(w_dff_A_QHuSf2Ia6_0),.clk(gclk));
	jdff dff_A_zS6HEnMW4_0(.dout(w_dff_A_wyp349xj3_0),.din(w_dff_A_zS6HEnMW4_0),.clk(gclk));
	jdff dff_A_wyp349xj3_0(.dout(w_dff_A_OSd91su29_0),.din(w_dff_A_wyp349xj3_0),.clk(gclk));
	jdff dff_A_OSd91su29_0(.dout(w_dff_A_yCUoTRVp8_0),.din(w_dff_A_OSd91su29_0),.clk(gclk));
	jdff dff_A_yCUoTRVp8_0(.dout(w_dff_A_iKhB3adl6_0),.din(w_dff_A_yCUoTRVp8_0),.clk(gclk));
	jdff dff_A_iKhB3adl6_0(.dout(G399),.din(w_dff_A_iKhB3adl6_0),.clk(gclk));
endmodule

