/*

c3540:
	jxor: 52
	jspl: 225
	jspl3: 338
	jnot: 188
	jdff: 2183
	jand: 525
	jor: 352

Summary:
	jxor: 52
	jspl: 225
	jspl3: 338
	jnot: 188
	jdff: 2183
	jand: 525
	jor: 352
*/

module c3540(gclk, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698, G2897, G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402);
	input gclk;
	input G1;
	input G13;
	input G20;
	input G33;
	input G41;
	input G45;
	input G50;
	input G58;
	input G68;
	input G77;
	input G87;
	input G97;
	input G107;
	input G116;
	input G124;
	input G125;
	input G128;
	input G132;
	input G137;
	input G143;
	input G150;
	input G159;
	input G169;
	input G179;
	input G190;
	input G200;
	input G213;
	input G222;
	input G223;
	input G226;
	input G232;
	input G238;
	input G244;
	input G250;
	input G257;
	input G264;
	input G270;
	input G274;
	input G283;
	input G294;
	input G303;
	input G311;
	input G317;
	input G322;
	input G326;
	input G329;
	input G330;
	input G343;
	input G1698;
	input G2897;
	output G353;
	output G355;
	output G361;
	output G358;
	output G351;
	output G372;
	output G369;
	output G399;
	output G364;
	output G396;
	output G384;
	output G367;
	output G387;
	output G393;
	output G390;
	output G378;
	output G375;
	output G381;
	output G407;
	output G409;
	output G405;
	output G402;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire [2:0] w_G1_0;
	wire [2:0] w_G1_1;
	wire [1:0] w_G1_2;
	wire [2:0] w_G13_0;
	wire [2:0] w_G13_1;
	wire [1:0] w_G13_2;
	wire [2:0] w_G20_0;
	wire [2:0] w_G20_1;
	wire [2:0] w_G20_2;
	wire [2:0] w_G20_3;
	wire [2:0] w_G20_4;
	wire [2:0] w_G20_5;
	wire [2:0] w_G20_6;
	wire [2:0] w_G33_0;
	wire [2:0] w_G33_1;
	wire [2:0] w_G33_2;
	wire [2:0] w_G33_3;
	wire [2:0] w_G33_4;
	wire [2:0] w_G33_5;
	wire [2:0] w_G33_6;
	wire [2:0] w_G33_7;
	wire [2:0] w_G33_8;
	wire [2:0] w_G33_9;
	wire [2:0] w_G33_10;
	wire [2:0] w_G33_11;
	wire [2:0] w_G33_12;
	wire [2:0] w_G41_0;
	wire [2:0] w_G45_0;
	wire [1:0] w_G45_1;
	wire [2:0] w_G50_0;
	wire [2:0] w_G50_1;
	wire [2:0] w_G50_2;
	wire [2:0] w_G50_3;
	wire [2:0] w_G50_4;
	wire [2:0] w_G50_5;
	wire [2:0] w_G58_0;
	wire [2:0] w_G58_1;
	wire [2:0] w_G58_2;
	wire [2:0] w_G58_3;
	wire [2:0] w_G58_4;
	wire [2:0] w_G58_5;
	wire [2:0] w_G68_0;
	wire [2:0] w_G68_1;
	wire [2:0] w_G68_2;
	wire [2:0] w_G68_3;
	wire [2:0] w_G68_4;
	wire [2:0] w_G68_5;
	wire [2:0] w_G77_0;
	wire [2:0] w_G77_1;
	wire [2:0] w_G77_2;
	wire [2:0] w_G77_3;
	wire [2:0] w_G77_4;
	wire [2:0] w_G87_0;
	wire [2:0] w_G87_1;
	wire [2:0] w_G87_2;
	wire [2:0] w_G87_3;
	wire [2:0] w_G97_0;
	wire [2:0] w_G97_1;
	wire [2:0] w_G97_2;
	wire [2:0] w_G97_3;
	wire [2:0] w_G97_4;
	wire [2:0] w_G107_0;
	wire [2:0] w_G107_1;
	wire [2:0] w_G107_2;
	wire [2:0] w_G107_3;
	wire [1:0] w_G107_4;
	wire [2:0] w_G116_0;
	wire [2:0] w_G116_1;
	wire [2:0] w_G116_2;
	wire [2:0] w_G116_3;
	wire [2:0] w_G116_4;
	wire [2:0] w_G116_5;
	wire [1:0] w_G125_0;
	wire [2:0] w_G128_0;
	wire [2:0] w_G132_0;
	wire [1:0] w_G132_1;
	wire [2:0] w_G137_0;
	wire [2:0] w_G137_1;
	wire [2:0] w_G143_0;
	wire [2:0] w_G143_1;
	wire [1:0] w_G143_2;
	wire [2:0] w_G150_0;
	wire [2:0] w_G150_1;
	wire [2:0] w_G150_2;
	wire [1:0] w_G150_3;
	wire [2:0] w_G159_0;
	wire [2:0] w_G159_1;
	wire [2:0] w_G159_2;
	wire [2:0] w_G159_3;
	wire [2:0] w_G169_0;
	wire [2:0] w_G169_1;
	wire [2:0] w_G169_2;
	wire [1:0] w_G169_3;
	wire [2:0] w_G179_0;
	wire [2:0] w_G179_1;
	wire [2:0] w_G179_2;
	wire [2:0] w_G190_0;
	wire [2:0] w_G190_1;
	wire [2:0] w_G190_2;
	wire [2:0] w_G190_3;
	wire [2:0] w_G190_4;
	wire [2:0] w_G200_0;
	wire [2:0] w_G200_1;
	wire [2:0] w_G200_2;
	wire [1:0] w_G200_3;
	wire [2:0] w_G213_0;
	wire [1:0] w_G223_0;
	wire [2:0] w_G226_0;
	wire [2:0] w_G226_1;
	wire [2:0] w_G232_0;
	wire [2:0] w_G232_1;
	wire [2:0] w_G238_0;
	wire [2:0] w_G244_0;
	wire [1:0] w_G244_1;
	wire [2:0] w_G250_0;
	wire [2:0] w_G257_0;
	wire [2:0] w_G257_1;
	wire [2:0] w_G264_0;
	wire [2:0] w_G270_0;
	wire [2:0] w_G274_0;
	wire [2:0] w_G283_0;
	wire [2:0] w_G283_1;
	wire [2:0] w_G283_2;
	wire [2:0] w_G283_3;
	wire [2:0] w_G294_0;
	wire [2:0] w_G294_1;
	wire [2:0] w_G294_2;
	wire [1:0] w_G294_3;
	wire [2:0] w_G303_0;
	wire [2:0] w_G303_1;
	wire [2:0] w_G303_2;
	wire [2:0] w_G311_0;
	wire [2:0] w_G311_1;
	wire [2:0] w_G317_0;
	wire [1:0] w_G317_1;
	wire [2:0] w_G322_0;
	wire [1:0] w_G326_0;
	wire [2:0] w_G330_0;
	wire [1:0] w_G343_0;
	wire [2:0] w_G1698_0;
	wire w_G355_0;
	wire G355_fa_;
	wire w_G396_0;
	wire G396_fa_;
	wire w_G384_0;
	wire G384_fa_;
	wire [2:0] w_n72_0;
	wire [2:0] w_n72_1;
	wire [2:0] w_n73_0;
	wire [2:0] w_n73_1;
	wire [2:0] w_n73_2;
	wire [2:0] w_n74_0;
	wire [2:0] w_n74_1;
	wire [1:0] w_n74_2;
	wire [2:0] w_n75_0;
	wire [2:0] w_n75_1;
	wire [1:0] w_n75_2;
	wire [1:0] w_n76_0;
	wire [1:0] w_n77_0;
	wire [2:0] w_n79_0;
	wire [2:0] w_n79_1;
	wire [2:0] w_n80_0;
	wire [2:0] w_n80_1;
	wire [2:0] w_n81_0;
	wire [2:0] w_n81_1;
	wire [1:0] w_n81_2;
	wire [2:0] w_n84_0;
	wire [2:0] w_n84_1;
	wire [1:0] w_n85_0;
	wire [2:0] w_n86_0;
	wire [1:0] w_n89_0;
	wire [2:0] w_n90_0;
	wire [2:0] w_n91_0;
	wire [2:0] w_n91_1;
	wire [2:0] w_n94_0;
	wire [2:0] w_n96_0;
	wire [2:0] w_n105_0;
	wire [1:0] w_n105_1;
	wire [2:0] w_n111_0;
	wire [1:0] w_n112_0;
	wire [2:0] w_n118_0;
	wire [1:0] w_n120_0;
	wire [1:0] w_n126_0;
	wire [1:0] w_n130_0;
	wire [1:0] w_n134_0;
	wire [1:0] w_n137_0;
	wire [2:0] w_n139_0;
	wire [2:0] w_n139_1;
	wire [1:0] w_n140_0;
	wire [2:0] w_n141_0;
	wire [2:0] w_n141_1;
	wire [2:0] w_n141_2;
	wire [1:0] w_n141_3;
	wire [2:0] w_n142_0;
	wire [2:0] w_n142_1;
	wire [1:0] w_n142_2;
	wire [1:0] w_n143_0;
	wire [2:0] w_n144_0;
	wire [2:0] w_n144_1;
	wire [1:0] w_n144_2;
	wire [2:0] w_n147_0;
	wire [1:0] w_n148_0;
	wire [2:0] w_n151_0;
	wire [2:0] w_n151_1;
	wire [2:0] w_n151_2;
	wire [2:0] w_n151_3;
	wire [2:0] w_n151_4;
	wire [2:0] w_n151_5;
	wire [1:0] w_n151_6;
	wire [2:0] w_n152_0;
	wire [2:0] w_n153_0;
	wire [2:0] w_n153_1;
	wire [2:0] w_n153_2;
	wire [2:0] w_n153_3;
	wire [2:0] w_n153_4;
	wire [2:0] w_n153_5;
	wire [2:0] w_n153_6;
	wire [2:0] w_n153_7;
	wire [1:0] w_n153_8;
	wire [2:0] w_n161_0;
	wire [2:0] w_n163_0;
	wire [1:0] w_n163_1;
	wire [2:0] w_n164_0;
	wire [1:0] w_n165_0;
	wire [1:0] w_n167_0;
	wire [2:0] w_n168_0;
	wire [2:0] w_n168_1;
	wire [2:0] w_n168_2;
	wire [2:0] w_n168_3;
	wire [2:0] w_n168_4;
	wire [1:0] w_n168_5;
	wire [1:0] w_n169_0;
	wire [2:0] w_n170_0;
	wire [2:0] w_n172_0;
	wire [2:0] w_n172_1;
	wire [2:0] w_n172_2;
	wire [2:0] w_n172_3;
	wire [2:0] w_n172_4;
	wire [2:0] w_n173_0;
	wire [2:0] w_n173_1;
	wire [2:0] w_n173_2;
	wire [1:0] w_n173_3;
	wire [1:0] w_n176_0;
	wire [2:0] w_n177_0;
	wire [2:0] w_n177_1;
	wire [2:0] w_n182_0;
	wire [1:0] w_n182_1;
	wire [2:0] w_n186_0;
	wire [2:0] w_n186_1;
	wire [2:0] w_n189_0;
	wire [2:0] w_n189_1;
	wire [2:0] w_n189_2;
	wire [1:0] w_n190_0;
	wire [2:0] w_n192_0;
	wire [2:0] w_n198_0;
	wire [2:0] w_n199_0;
	wire [1:0] w_n201_0;
	wire [1:0] w_n202_0;
	wire [2:0] w_n205_0;
	wire [1:0] w_n205_1;
	wire [1:0] w_n207_0;
	wire [2:0] w_n212_0;
	wire [1:0] w_n212_1;
	wire [1:0] w_n213_0;
	wire [1:0] w_n215_0;
	wire [1:0] w_n218_0;
	wire [2:0] w_n224_0;
	wire [1:0] w_n224_1;
	wire [1:0] w_n225_0;
	wire [1:0] w_n229_0;
	wire [2:0] w_n234_0;
	wire [1:0] w_n234_1;
	wire [2:0] w_n237_0;
	wire [1:0] w_n238_0;
	wire [2:0] w_n242_0;
	wire [1:0] w_n243_0;
	wire [1:0] w_n247_0;
	wire [1:0] w_n250_0;
	wire [1:0] w_n251_0;
	wire [2:0] w_n255_0;
	wire [1:0] w_n255_1;
	wire [1:0] w_n256_0;
	wire [1:0] w_n257_0;
	wire [1:0] w_n259_0;
	wire [1:0] w_n260_0;
	wire [2:0] w_n261_0;
	wire [2:0] w_n261_1;
	wire [2:0] w_n262_0;
	wire [1:0] w_n269_0;
	wire [1:0] w_n272_0;
	wire [2:0] w_n279_0;
	wire [1:0] w_n279_1;
	wire [1:0] w_n282_0;
	wire [1:0] w_n283_0;
	wire [2:0] w_n292_0;
	wire [1:0] w_n298_0;
	wire [2:0] w_n308_0;
	wire [2:0] w_n308_1;
	wire [1:0] w_n309_0;
	wire [1:0] w_n310_0;
	wire [1:0] w_n312_0;
	wire [1:0] w_n313_0;
	wire [2:0] w_n315_0;
	wire [1:0] w_n321_0;
	wire [2:0] w_n323_0;
	wire [2:0] w_n330_0;
	wire [1:0] w_n333_0;
	wire [1:0] w_n334_0;
	wire [1:0] w_n344_0;
	wire [1:0] w_n347_0;
	wire [1:0] w_n348_0;
	wire [1:0] w_n349_0;
	wire [1:0] w_n350_0;
	wire [1:0] w_n351_0;
	wire [2:0] w_n352_0;
	wire [1:0] w_n352_1;
	wire [2:0] w_n354_0;
	wire [1:0] w_n354_1;
	wire [1:0] w_n355_0;
	wire [2:0] w_n356_0;
	wire [1:0] w_n356_1;
	wire [1:0] w_n357_0;
	wire [2:0] w_n367_0;
	wire [1:0] w_n367_1;
	wire [1:0] w_n370_0;
	wire [1:0] w_n375_0;
	wire [1:0] w_n378_0;
	wire [2:0] w_n383_0;
	wire [2:0] w_n387_0;
	wire [2:0] w_n388_0;
	wire [2:0] w_n388_1;
	wire [1:0] w_n388_2;
	wire [1:0] w_n394_0;
	wire [1:0] w_n395_0;
	wire [2:0] w_n404_0;
	wire [1:0] w_n405_0;
	wire [1:0] w_n407_0;
	wire [2:0] w_n414_0;
	wire [2:0] w_n417_0;
	wire [1:0] w_n420_0;
	wire [1:0] w_n425_0;
	wire [1:0] w_n426_0;
	wire [1:0] w_n428_0;
	wire [1:0] w_n430_0;
	wire [1:0] w_n435_0;
	wire [2:0] w_n439_0;
	wire [1:0] w_n441_0;
	wire [1:0] w_n445_0;
	wire [1:0] w_n450_0;
	wire [1:0] w_n452_0;
	wire [1:0] w_n456_0;
	wire [1:0] w_n457_0;
	wire [1:0] w_n465_0;
	wire [1:0] w_n472_0;
	wire [1:0] w_n473_0;
	wire [2:0] w_n482_0;
	wire [1:0] w_n483_0;
	wire [1:0] w_n494_0;
	wire [1:0] w_n499_0;
	wire [1:0] w_n500_0;
	wire [2:0] w_n503_0;
	wire [2:0] w_n507_0;
	wire [2:0] w_n507_1;
	wire [1:0] w_n507_2;
	wire [1:0] w_n511_0;
	wire [1:0] w_n512_0;
	wire [2:0] w_n514_0;
	wire [1:0] w_n514_1;
	wire [1:0] w_n520_0;
	wire [1:0] w_n533_0;
	wire [1:0] w_n534_0;
	wire [1:0] w_n541_0;
	wire [1:0] w_n542_0;
	wire [1:0] w_n543_0;
	wire [1:0] w_n544_0;
	wire [1:0] w_n548_0;
	wire [1:0] w_n550_0;
	wire [1:0] w_n551_0;
	wire [1:0] w_n559_0;
	wire [1:0] w_n562_0;
	wire [2:0] w_n566_0;
	wire [1:0] w_n566_1;
	wire [2:0] w_n567_0;
	wire [2:0] w_n567_1;
	wire [2:0] w_n567_2;
	wire [2:0] w_n567_3;
	wire [2:0] w_n567_4;
	wire [1:0] w_n567_5;
	wire [1:0] w_n569_0;
	wire [1:0] w_n570_0;
	wire [2:0] w_n571_0;
	wire [2:0] w_n571_1;
	wire [1:0] w_n571_2;
	wire [2:0] w_n572_0;
	wire [1:0] w_n573_0;
	wire [1:0] w_n574_0;
	wire [2:0] w_n576_0;
	wire [1:0] w_n577_0;
	wire [2:0] w_n579_0;
	wire [1:0] w_n579_1;
	wire [2:0] w_n580_0;
	wire [1:0] w_n582_0;
	wire [1:0] w_n584_0;
	wire [1:0] w_n598_0;
	wire [2:0] w_n600_0;
	wire [2:0] w_n600_1;
	wire [2:0] w_n601_0;
	wire [1:0] w_n602_0;
	wire [2:0] w_n604_0;
	wire [2:0] w_n604_1;
	wire [2:0] w_n604_2;
	wire [2:0] w_n605_0;
	wire [2:0] w_n613_0;
	wire [2:0] w_n613_1;
	wire [2:0] w_n614_0;
	wire [2:0] w_n614_1;
	wire [2:0] w_n614_2;
	wire [2:0] w_n614_3;
	wire [2:0] w_n614_4;
	wire [1:0] w_n614_5;
	wire [2:0] w_n618_0;
	wire [2:0] w_n618_1;
	wire [1:0] w_n618_2;
	wire [2:0] w_n619_0;
	wire [2:0] w_n620_0;
	wire [1:0] w_n622_0;
	wire [1:0] w_n624_0;
	wire [2:0] w_n626_0;
	wire [1:0] w_n628_0;
	wire [2:0] w_n629_0;
	wire [2:0] w_n629_1;
	wire [2:0] w_n629_2;
	wire [2:0] w_n629_3;
	wire [2:0] w_n629_4;
	wire [1:0] w_n629_5;
	wire [1:0] w_n630_0;
	wire [1:0] w_n632_0;
	wire [2:0] w_n633_0;
	wire [2:0] w_n633_1;
	wire [2:0] w_n633_2;
	wire [2:0] w_n633_3;
	wire [2:0] w_n633_4;
	wire [2:0] w_n633_5;
	wire [1:0] w_n633_6;
	wire [1:0] w_n634_0;
	wire [1:0] w_n637_0;
	wire [2:0] w_n638_0;
	wire [2:0] w_n638_1;
	wire [2:0] w_n638_2;
	wire [2:0] w_n638_3;
	wire [2:0] w_n638_4;
	wire [2:0] w_n638_5;
	wire [2:0] w_n638_6;
	wire [1:0] w_n638_7;
	wire [2:0] w_n640_0;
	wire [2:0] w_n640_1;
	wire [2:0] w_n640_2;
	wire [2:0] w_n640_3;
	wire [2:0] w_n640_4;
	wire [2:0] w_n640_5;
	wire [2:0] w_n640_6;
	wire [1:0] w_n640_7;
	wire [2:0] w_n646_0;
	wire [2:0] w_n646_1;
	wire [2:0] w_n646_2;
	wire [2:0] w_n646_3;
	wire [2:0] w_n646_4;
	wire [2:0] w_n646_5;
	wire [2:0] w_n646_6;
	wire [1:0] w_n646_7;
	wire [2:0] w_n648_0;
	wire [2:0] w_n648_1;
	wire [2:0] w_n648_2;
	wire [2:0] w_n648_3;
	wire [1:0] w_n648_4;
	wire [1:0] w_n649_0;
	wire [1:0] w_n650_0;
	wire [2:0] w_n651_0;
	wire [2:0] w_n651_1;
	wire [2:0] w_n651_2;
	wire [2:0] w_n651_3;
	wire [2:0] w_n651_4;
	wire [2:0] w_n651_5;
	wire [2:0] w_n651_6;
	wire [1:0] w_n651_7;
	wire [2:0] w_n653_0;
	wire [2:0] w_n653_1;
	wire [2:0] w_n653_2;
	wire [2:0] w_n653_3;
	wire [2:0] w_n653_4;
	wire [2:0] w_n653_5;
	wire [2:0] w_n653_6;
	wire [1:0] w_n653_7;
	wire [2:0] w_n680_0;
	wire [2:0] w_n680_1;
	wire [2:0] w_n680_2;
	wire [2:0] w_n680_3;
	wire [1:0] w_n680_4;
	wire [1:0] w_n682_0;
	wire [2:0] w_n684_0;
	wire [1:0] w_n685_0;
	wire [2:0] w_n690_0;
	wire [1:0] w_n690_1;
	wire [1:0] w_n692_0;
	wire [2:0] w_n703_0;
	wire [1:0] w_n703_1;
	wire [1:0] w_n704_0;
	wire [1:0] w_n718_0;
	wire [1:0] w_n733_0;
	wire [2:0] w_n741_0;
	wire [1:0] w_n741_1;
	wire [1:0] w_n748_0;
	wire [1:0] w_n754_0;
	wire [1:0] w_n759_0;
	wire [1:0] w_n766_0;
	wire [2:0] w_n767_0;
	wire [1:0] w_n767_1;
	wire [2:0] w_n771_0;
	wire [1:0] w_n771_1;
	wire [1:0] w_n772_0;
	wire [1:0] w_n773_0;
	wire [1:0] w_n775_0;
	wire [1:0] w_n777_0;
	wire [1:0] w_n782_0;
	wire [1:0] w_n798_0;
	wire [2:0] w_n802_0;
	wire [1:0] w_n817_0;
	wire [1:0] w_n830_0;
	wire [1:0] w_n833_0;
	wire [2:0] w_n845_0;
	wire [1:0] w_n855_0;
	wire [1:0] w_n860_0;
	wire [1:0] w_n861_0;
	wire [2:0] w_n863_0;
	wire [2:0] w_n869_0;
	wire [1:0] w_n873_0;
	wire [1:0] w_n875_0;
	wire [1:0] w_n884_0;
	wire [1:0] w_n887_0;
	wire [2:0] w_n937_0;
	wire [1:0] w_n959_0;
	wire [2:0] w_n987_0;
	wire [2:0] w_n1029_0;
	wire [1:0] w_n1033_0;
	wire [1:0] w_n1036_0;
	wire [1:0] w_n1039_0;
	wire [1:0] w_n1040_0;
	wire [1:0] w_n1041_0;
	wire [1:0] w_n1043_0;
	wire [1:0] w_n1044_0;
	wire [1:0] w_n1045_0;
	wire [1:0] w_n1048_0;
	wire [2:0] w_n1053_0;
	wire [1:0] w_n1056_0;
	wire [1:0] w_n1062_0;
	wire [1:0] w_n1091_0;
	wire [2:0] w_n1114_0;
	wire [2:0] w_n1159_0;
	wire [1:0] w_n1161_0;
	wire [1:0] w_n1164_0;
	wire [1:0] w_n1168_0;
	wire [1:0] w_n1170_0;
	wire [1:0] w_n1177_0;
	wire [1:0] w_n1178_0;
	wire [1:0] w_n1179_0;
	wire [1:0] w_n1184_0;
	wire w_dff_B_FisDzS2G3_1;
	wire w_dff_B_6qk4aTx82_1;
	wire w_dff_B_JvinlRL29_1;
	wire w_dff_B_TDSDGv6d9_0;
	wire w_dff_B_Ihv2Jms46_0;
	wire w_dff_B_C6ZHnywj8_1;
	wire w_dff_B_hMorE4od6_1;
	wire w_dff_B_EGuQuSgs1_0;
	wire w_dff_B_TASNkIqq7_1;
	wire w_dff_B_Woaokfvf6_1;
	wire w_dff_B_QTLoulrx0_1;
	wire w_dff_B_08OolUYY8_1;
	wire w_dff_B_GrXsNCMJ1_1;
	wire w_dff_B_BEAgXbjz7_1;
	wire w_dff_B_Bvb69Xmu7_1;
	wire w_dff_B_8zPPKHFI8_1;
	wire w_dff_B_0wR6m3aT5_1;
	wire w_dff_B_uwdEgYRk7_1;
	wire w_dff_B_AcMmPzkD8_1;
	wire w_dff_B_FyC6zzOK0_1;
	wire w_dff_B_tvCErOkh9_1;
	wire w_dff_B_IiicwIpp4_1;
	wire w_dff_B_bhqxOEXJ8_1;
	wire w_dff_B_EQCVdU6e3_1;
	wire w_dff_B_tkqstEIK6_0;
	wire w_dff_B_tNVLTYxr0_0;
	wire w_dff_B_QSMvEAzn2_0;
	wire w_dff_B_N8qLehVz8_0;
	wire w_dff_B_iTzdb2r78_0;
	wire w_dff_B_irI9PjkJ7_0;
	wire w_dff_B_nZgEs5t84_0;
	wire w_dff_B_ni6t9HIS6_0;
	wire w_dff_B_mtzlxig94_0;
	wire w_dff_B_BzfrBKk04_0;
	wire w_dff_B_8L2g9nce6_0;
	wire w_dff_B_0QPvJRGD3_0;
	wire w_dff_B_lnBonCWs7_0;
	wire w_dff_B_UReCyPV51_0;
	wire w_dff_B_Kwxh1Sr80_0;
	wire w_dff_B_6wTKYiMy6_0;
	wire w_dff_B_HNxUzeNO3_0;
	wire w_dff_B_8y5Qywf70_0;
	wire w_dff_B_qz0yT4u13_0;
	wire w_dff_B_ujE6Yytb4_0;
	wire w_dff_B_Jgozzp5O5_0;
	wire w_dff_B_Ij2wRnEv9_0;
	wire w_dff_B_sVx04yGb5_0;
	wire w_dff_B_yxPDP1Hg4_0;
	wire w_dff_B_PQqpOgbm4_0;
	wire w_dff_B_IW7K4Xhv7_0;
	wire w_dff_B_Xk7HAGc29_0;
	wire w_dff_B_VXjQKKOq0_0;
	wire w_dff_B_pzOzuQKD8_0;
	wire w_dff_B_aXgPwDHK0_0;
	wire w_dff_B_tv2ZYgBB6_0;
	wire w_dff_B_YjUwNIFM7_0;
	wire w_dff_A_DQoYhr6W3_1;
	wire w_dff_A_TyPS3WoP1_1;
	wire w_dff_A_UDU0rIU67_1;
	wire w_dff_B_1OBZCMhy3_0;
	wire w_dff_B_tSx2xLMj3_1;
	wire w_dff_B_C8rCXM4B9_1;
	wire w_dff_B_G0UMSRUW8_1;
	wire w_dff_B_BkJ0qat38_1;
	wire w_dff_B_fUV0KDod1_1;
	wire w_dff_B_666hIiDX3_1;
	wire w_dff_B_Xmye5mS34_1;
	wire w_dff_B_xVzKSrU77_1;
	wire w_dff_B_d7gv71Hn9_1;
	wire w_dff_B_C5TkIlfG6_1;
	wire w_dff_B_PWsTpzww3_1;
	wire w_dff_B_CJ0tkKYS7_1;
	wire w_dff_B_t7byUmWW0_1;
	wire w_dff_B_71Z0PtaJ2_1;
	wire w_dff_B_GUTpCPzJ4_1;
	wire w_dff_B_80BwfMuo1_1;
	wire w_dff_B_lKf6zE3u4_1;
	wire w_dff_B_XEYBo1O55_1;
	wire w_dff_B_L1sWVBgv2_0;
	wire w_dff_A_l0vAzSjO1_0;
	wire w_dff_B_O0pQzvgJ1_1;
	wire w_dff_B_frMcGxgf5_1;
	wire w_dff_B_jqOtryg55_1;
	wire w_dff_B_oOkU1t0k3_1;
	wire w_dff_B_rExM3eu09_1;
	wire w_dff_B_VO0XmfdD9_1;
	wire w_dff_B_tm5M35OS1_1;
	wire w_dff_B_G1cOep062_1;
	wire w_dff_B_MQS5xDSO2_1;
	wire w_dff_B_CNW9yy9e7_1;
	wire w_dff_B_r4uPlvMp9_1;
	wire w_dff_B_E5Je6U2n4_1;
	wire w_dff_B_Cy6THfc74_1;
	wire w_dff_B_8n8mkhmR1_1;
	wire w_dff_B_sCyau8fA4_1;
	wire w_dff_B_n6B4OGTu7_1;
	wire w_dff_B_hWlgKtWM3_1;
	wire w_dff_B_iL5VXfsp1_1;
	wire w_dff_B_BdE3Le4u3_1;
	wire w_dff_B_e0Gwb0W57_1;
	wire w_dff_B_Ie3d7nLS0_1;
	wire w_dff_B_CacUVfs86_1;
	wire w_dff_B_x4oHjoEA8_1;
	wire w_dff_B_yTxwHFCj4_1;
	wire w_dff_B_dKsDdogj7_1;
	wire w_dff_B_BhqnfbyR0_1;
	wire w_dff_B_KQ6GFgsG1_1;
	wire w_dff_B_MknqKfFr2_1;
	wire w_dff_B_8HFEJnXu5_1;
	wire w_dff_B_FwJFZ6BF6_1;
	wire w_dff_B_AmjHcgx98_0;
	wire w_dff_B_48cNaTjh5_0;
	wire w_dff_A_bIPlIXri0_1;
	wire w_dff_B_aG3jgnq64_1;
	wire w_dff_B_ZAzMLZjE2_1;
	wire w_dff_B_743ovYwE6_1;
	wire w_dff_B_4dxmTCCL6_1;
	wire w_dff_B_Tr26cAK27_1;
	wire w_dff_B_p3kTBsde8_1;
	wire w_dff_B_ENVTFoNk4_1;
	wire w_dff_B_K0pcvSBU0_1;
	wire w_dff_B_LbYXLk3t8_1;
	wire w_dff_B_mRcD0r6B8_1;
	wire w_dff_B_ifODZ0W21_1;
	wire w_dff_B_C8Byw6xg1_1;
	wire w_dff_B_jIOcnVBj3_1;
	wire w_dff_B_kTZ06aED6_1;
	wire w_dff_B_0l7va75j8_1;
	wire w_dff_B_Af02HnkB5_1;
	wire w_dff_B_5ed415NZ0_1;
	wire w_dff_B_46wcFXb09_1;
	wire w_dff_B_haq2xpEC6_1;
	wire w_dff_B_HiuuKYU86_1;
	wire w_dff_B_2EP0XXjU0_1;
	wire w_dff_B_6vypaYpT5_1;
	wire w_dff_B_Su3dtXyJ0_1;
	wire w_dff_B_IDtFmd019_1;
	wire w_dff_B_lY2Ax7b13_1;
	wire w_dff_B_PpUIfjdo0_1;
	wire w_dff_B_kWRWoWwz2_1;
	wire w_dff_B_YEK212ql2_1;
	wire w_dff_B_cNXx9oAG3_1;
	wire w_dff_B_k27Nc5al7_1;
	wire w_dff_B_gdKSErvz3_1;
	wire w_dff_B_3YqxDNy86_1;
	wire w_dff_B_VOogdegQ3_1;
	wire w_dff_B_TrqHHWcp0_1;
	wire w_dff_B_Nv92AX2s3_1;
	wire w_dff_B_6O3fuYLp3_1;
	wire w_dff_B_z6hslOBF1_1;
	wire w_dff_B_yYF6DQEQ6_1;
	wire w_dff_B_nV7xsVl07_1;
	wire w_dff_B_3noChfJt3_1;
	wire w_dff_B_8u2om3fQ9_1;
	wire w_dff_B_gfaZYkfb7_1;
	wire w_dff_B_QfVH3H3o5_1;
	wire w_dff_B_GBSecZs41_1;
	wire w_dff_B_nJa0Ckn88_1;
	wire w_dff_B_4xK9j6Kk4_1;
	wire w_dff_B_DDcZLK1K1_1;
	wire w_dff_B_WxdgpjY17_1;
	wire w_dff_B_HE9qHSVP8_1;
	wire w_dff_B_IU7mi6NF8_1;
	wire w_dff_B_nVelMIe07_1;
	wire w_dff_B_fhFDzsU53_1;
	wire w_dff_A_oEkZzEYX3_1;
	wire w_dff_A_2aSPumVB0_1;
	wire w_dff_A_nc9pRLfW0_1;
	wire w_dff_A_ymO1q5WJ9_1;
	wire w_dff_A_97gF6N6G5_1;
	wire w_dff_A_DGqvrLS62_1;
	wire w_dff_A_xuAxr93G4_1;
	wire w_dff_A_uMceIChW0_1;
	wire w_dff_A_OJgpjU1k7_1;
	wire w_dff_A_sKgk3hIT5_1;
	wire w_dff_A_x8Ypizl98_1;
	wire w_dff_A_WTIedmAo2_1;
	wire w_dff_A_TIJGeD1Z6_1;
	wire w_dff_A_6zUO43MB8_1;
	wire w_dff_A_89fyoYdW2_1;
	wire w_dff_A_BtXQrUYB8_1;
	wire w_dff_A_DQGQIvbH8_1;
	wire w_dff_A_fC6BJDS77_1;
	wire w_dff_A_iv679SmZ3_1;
	wire w_dff_A_g74wpa3S6_1;
	wire w_dff_A_Q6aavcP76_1;
	wire w_dff_A_1ykcvOfP0_1;
	wire w_dff_A_Tv9wjDeq9_1;
	wire w_dff_A_oUsiejR33_1;
	wire w_dff_A_LHYgxu1A5_1;
	wire w_dff_A_632WFSdJ0_1;
	wire w_dff_A_dkfYjhzC3_1;
	wire w_dff_A_e1I1FwBw6_1;
	wire w_dff_A_EaGAQYq91_1;
	wire w_dff_A_TUSdV0av9_1;
	wire w_dff_A_R3xkoru75_1;
	wire w_dff_A_XoITSO2M6_1;
	wire w_dff_A_GEHe4JQR6_1;
	wire w_dff_A_6mCe0wye9_1;
	wire w_dff_A_MT7vUpff4_1;
	wire w_dff_A_HxieEi5Q0_1;
	wire w_dff_A_KzrAGZO89_1;
	wire w_dff_A_gsDHJLme9_1;
	wire w_dff_A_lFJsCO5g3_1;
	wire w_dff_A_yz6Ci5FY0_1;
	wire w_dff_A_l7UgMVOv0_1;
	wire w_dff_A_gmbyOslU0_1;
	wire w_dff_A_6WUQ2ZRA2_1;
	wire w_dff_A_J2vkXNR49_1;
	wire w_dff_A_zPe37f148_1;
	wire w_dff_A_GejfoAzr1_1;
	wire w_dff_A_ztItkpuL0_1;
	wire w_dff_A_ucWO2dQd1_1;
	wire w_dff_A_RBuzc3PJ3_1;
	wire w_dff_A_WE3vj2CX5_1;
	wire w_dff_A_lyWdlucm2_1;
	wire w_dff_A_ZQl9FZJa0_1;
	wire w_dff_B_xWGvZ6jQ1_0;
	wire w_dff_B_ig3HG5L75_0;
	wire w_dff_B_80ts38i57_0;
	wire w_dff_B_CjsrJNf85_0;
	wire w_dff_B_RtZjEUoh5_0;
	wire w_dff_B_NAj0O6MK7_0;
	wire w_dff_B_ZBwqG1ji1_0;
	wire w_dff_B_lJfyTnvH0_0;
	wire w_dff_B_1uOPiDZv0_0;
	wire w_dff_B_MNfomTFq9_0;
	wire w_dff_B_U8KLbiZe2_0;
	wire w_dff_B_qNxgxsmg8_0;
	wire w_dff_B_BLEwuBJe3_0;
	wire w_dff_B_YoznAWsr8_0;
	wire w_dff_B_Y1rcZzZB7_1;
	wire w_dff_B_LkeHFOvD2_1;
	wire w_dff_B_6QTp5PQ74_1;
	wire w_dff_B_i8UZeDtG7_1;
	wire w_dff_B_tR9yNUqP8_1;
	wire w_dff_B_CSSbkLuy4_1;
	wire w_dff_B_pSvqTTRd7_1;
	wire w_dff_B_mBKeCzen2_1;
	wire w_dff_B_oYNtwwoa6_1;
	wire w_dff_B_5RuyAYUz8_1;
	wire w_dff_B_6IigKEW58_1;
	wire w_dff_B_gUOa6haK3_0;
	wire w_dff_B_0idgkjQN3_1;
	wire w_dff_B_BK1PEsdO6_1;
	wire w_dff_B_LgGx67mV7_0;
	wire w_dff_B_qQIrSnQJ5_1;
	wire w_dff_B_x85OuUaa8_0;
	wire w_dff_B_m4XxvndL2_1;
	wire w_dff_B_Qxf9hIPF6_1;
	wire w_dff_B_H61T9q7t9_1;
	wire w_dff_B_RAbVov9X1_1;
	wire w_dff_B_cQ8DBxlb8_1;
	wire w_dff_B_pEDu6DlF5_0;
	wire w_dff_B_kXRsGkfF4_0;
	wire w_dff_B_QoyuoMYs5_0;
	wire w_dff_B_wqi3mgeV4_1;
	wire w_dff_A_HI2lnYjI5_1;
	wire w_dff_A_jLgJwv0p4_1;
	wire w_dff_A_nmBo6tOR0_1;
	wire w_dff_A_0rdu9bIW9_1;
	wire w_dff_A_Cr2CoSXm3_1;
	wire w_dff_A_EpSeeTrY9_1;
	wire w_dff_A_FKDTVBOb4_1;
	wire w_dff_A_siV6TsMS4_1;
	wire w_dff_B_fosDWTk39_0;
	wire w_dff_B_ZjAM4XCm8_0;
	wire w_dff_B_GkoJ5LLd8_1;
	wire w_dff_B_qN9kuMNm7_1;
	wire w_dff_B_UajQjeRI7_1;
	wire w_dff_B_677kXUgA3_1;
	wire w_dff_B_z4YEo8u39_1;
	wire w_dff_B_9j17tiSc0_1;
	wire w_dff_B_49cFV0nF6_1;
	wire w_dff_B_7Cxjwifc4_1;
	wire w_dff_A_Lx5EfmK91_1;
	wire w_dff_A_JfapGmZe9_1;
	wire w_dff_A_K39VnRtC5_1;
	wire w_dff_B_c5F11mB04_0;
	wire w_dff_B_1OmdDj2w7_0;
	wire w_dff_B_wEulYuc23_0;
	wire w_dff_B_BQmU4Cyx9_0;
	wire w_dff_B_EH72ZePG7_0;
	wire w_dff_B_QanFgOYD7_0;
	wire w_dff_B_zeMOrs7R0_0;
	wire w_dff_B_w1V2tbQf1_1;
	wire w_dff_B_jP4u0LC54_1;
	wire w_dff_B_MpNgiRne8_1;
	wire w_dff_B_IxRQbdCt3_1;
	wire w_dff_B_FPvrbdE18_1;
	wire w_dff_B_IWf6MZfP4_1;
	wire w_dff_B_Cdqyq45c9_1;
	wire w_dff_B_rMuyGdqc6_1;
	wire w_dff_B_fIWXbCll5_0;
	wire w_dff_A_FRgHQq6A9_1;
	wire w_dff_A_6YUtQTR05_1;
	wire w_dff_B_eEPnibS64_1;
	wire w_dff_B_6lVSt8ed3_1;
	wire w_dff_A_TA13gUh84_1;
	wire w_dff_A_kZIueL6h2_1;
	wire w_dff_A_NRLBxT1t3_1;
	wire w_dff_A_EyzfIyiW1_1;
	wire w_dff_A_fdpzGfW16_1;
	wire w_dff_A_YktNIekQ9_2;
	wire w_dff_A_Z9sBJwWm2_2;
	wire w_dff_A_rKBlyUaW6_2;
	wire w_dff_B_oOwqTsSo4_3;
	wire w_dff_B_gWNyL8z93_3;
	wire w_dff_A_pHISlmdY7_1;
	wire w_dff_B_4I3jzZeY7_0;
	wire w_dff_B_iiwKL2hO2_0;
	wire w_dff_B_6bHBSDGV1_0;
	wire w_dff_B_BiuoirYW2_0;
	wire w_dff_B_dlBr8R3K6_0;
	wire w_dff_B_sjjFa77P5_0;
	wire w_dff_B_mgULKXz23_1;
	wire w_dff_B_XudOkgBB5_1;
	wire w_dff_B_Gl0g4FKD0_0;
	wire w_dff_B_fYOfFF587_1;
	wire w_dff_B_zxYraqje1_1;
	wire w_dff_B_wzqu9s0k8_1;
	wire w_dff_B_GZqDTNiB8_1;
	wire w_dff_B_zHp34f0p2_1;
	wire w_dff_B_dv2uFe8e2_1;
	wire w_dff_B_77O0B9s62_1;
	wire w_dff_B_3LiZdvJa5_1;
	wire w_dff_B_ZSMIrfLb0_0;
	wire w_dff_B_Ijayki2N9_1;
	wire w_dff_A_OAACL1iP1_1;
	wire w_dff_B_zerNUWn88_2;
	wire w_dff_B_r6X535Li1_2;
	wire w_dff_B_NXq1WUpR1_2;
	wire w_dff_A_30wqftnc0_0;
	wire w_dff_A_CCYaXbSh6_0;
	wire w_dff_A_dLJ03ZvW5_0;
	wire w_dff_A_a8uuI0z37_1;
	wire w_dff_A_N746gYgC1_1;
	wire w_dff_A_cTD5tyEA5_1;
	wire w_dff_A_FMSR0ZCj0_1;
	wire w_dff_A_I4CaDGW37_1;
	wire w_dff_A_kVQKTSbv0_1;
	wire w_dff_A_rdz1rvvg2_1;
	wire w_dff_A_fXYDABUs7_1;
	wire w_dff_A_YHZ9rSjz4_1;
	wire w_dff_A_8oeDgHHV2_1;
	wire w_dff_A_POL1wn4v6_1;
	wire w_dff_B_1QEF5TMg9_0;
	wire w_dff_B_Y3vRi9GH1_0;
	wire w_dff_B_36qOmuvW2_1;
	wire w_dff_B_VHTaDOFl1_1;
	wire w_dff_B_zvs1keRG1_1;
	wire w_dff_B_n8p0L0ug4_1;
	wire w_dff_B_FdkCw2n75_1;
	wire w_dff_B_LHKZR8h56_1;
	wire w_dff_B_3mkVTSnB2_0;
	wire w_dff_B_kjZSD6wT0_1;
	wire w_dff_B_ukbYK3mL7_0;
	wire w_dff_A_MvoiZR3U7_0;
	wire w_dff_A_EGrOcpeG1_1;
	wire w_dff_A_hhoYO9hg9_1;
	wire w_dff_A_HT9a3MaW1_2;
	wire w_dff_A_v1McfurO5_2;
	wire w_dff_A_FRkws6Vl4_0;
	wire w_dff_B_vix8ijZT3_1;
	wire w_dff_B_d2AqgI6h4_1;
	wire w_dff_B_t9FRZKtK5_1;
	wire w_dff_B_RJARQDl49_1;
	wire w_dff_B_xhe3WgjF4_1;
	wire w_dff_B_AibjIE2U8_1;
	wire w_dff_A_iTgn9Xz62_0;
	wire w_dff_B_K4FHGxx43_1;
	wire w_dff_A_DNdT5Ak99_1;
	wire w_dff_A_HCXleRxp7_1;
	wire w_dff_A_KV5z3AXq7_1;
	wire w_dff_A_OxPTfjlh4_1;
	wire w_dff_A_bFCQX2iL3_1;
	wire w_dff_A_eaHt07N52_1;
	wire w_dff_A_BGJNNgD99_2;
	wire w_dff_A_JaMkopz46_2;
	wire w_dff_A_Cx0w8QtE6_2;
	wire w_dff_A_3GyNeKS69_0;
	wire w_dff_B_61EjpAtY1_1;
	wire w_dff_B_0SZdy8yD4_1;
	wire w_dff_B_XwAHOEav0_1;
	wire w_dff_B_Ubi5PWTg3_1;
	wire w_dff_B_vkJ7ryfr0_1;
	wire w_dff_B_CqwipQjJ2_1;
	wire w_dff_B_uIKuRZbo0_1;
	wire w_dff_B_kJhu1W4f8_1;
	wire w_dff_A_Ydbojq200_1;
	wire w_dff_A_NCw5ISe29_0;
	wire w_dff_B_EV0oZ51Q6_1;
	wire w_dff_A_fM9TVJlP3_0;
	wire w_dff_A_4toUY6Qz0_0;
	wire w_dff_A_d5tGjkKH7_0;
	wire w_dff_A_SGTn5YJd4_2;
	wire w_dff_A_PqZgsTd56_2;
	wire w_dff_A_8lVb8cug4_2;
	wire w_dff_B_2nIrxPWo3_1;
	wire w_dff_A_b7shwyO36_1;
	wire w_dff_A_c23foJsE2_0;
	wire w_dff_B_bbh4JCIm1_2;
	wire w_dff_B_F2IAu7YI9_2;
	wire w_dff_A_4YrgVHni8_0;
	wire w_dff_A_RFNPLB650_0;
	wire w_dff_A_XhzSou9P1_0;
	wire w_dff_A_EwJdGVxo2_0;
	wire w_dff_B_AjqoEEW30_2;
	wire w_dff_A_5vTYak7O9_1;
	wire w_dff_A_9305tNKF3_0;
	wire w_dff_A_Zmg066ZD5_0;
	wire w_dff_A_KNoPRY6W5_0;
	wire w_dff_A_7JEsw6sy5_0;
	wire w_dff_A_mXsJ5cto9_0;
	wire w_dff_A_89d5J4bx4_0;
	wire w_dff_A_SWu8eWN90_0;
	wire w_dff_B_5VUEyggF9_0;
	wire w_dff_B_0AwsjEXO5_0;
	wire w_dff_B_5q9U8p1K7_0;
	wire w_dff_B_2zIANsAj2_0;
	wire w_dff_B_BwhTBNMm1_0;
	wire w_dff_B_48tfzXcl0_0;
	wire w_dff_B_psmvs0JI6_0;
	wire w_dff_B_lT5Ns2Yr0_0;
	wire w_dff_B_4HbUW6mA5_0;
	wire w_dff_B_pPIEZ9EV1_0;
	wire w_dff_B_LQeloxLE6_0;
	wire w_dff_B_eaKMHYqK0_1;
	wire w_dff_B_NlD4pxdV4_1;
	wire w_dff_B_pds4Bk8m8_1;
	wire w_dff_B_F4vkc31U9_1;
	wire w_dff_B_wKM8UG592_1;
	wire w_dff_B_sE2vD7Q96_1;
	wire w_dff_B_mKbZNNwd7_1;
	wire w_dff_B_oazDjgne2_1;
	wire w_dff_B_D74Jixrd2_1;
	wire w_dff_B_TQMJOALO8_1;
	wire w_dff_B_mdsd82Yu5_1;
	wire w_dff_A_UshgANoK0_0;
	wire w_dff_B_J67n9Fgl9_3;
	wire w_dff_B_yr1c9DKG0_3;
	wire w_dff_B_5uutoYik1_3;
	wire w_dff_A_6WtM1vEI3_0;
	wire w_dff_A_H3r4BdW72_1;
	wire w_dff_A_9GG5FGtY4_1;
	wire w_dff_A_8hjcKo8F0_1;
	wire w_dff_A_0zdnIMgX1_1;
	wire w_dff_B_26OSP5554_1;
	wire w_dff_B_vMDHdvrG4_1;
	wire w_dff_A_9reIYKkx5_0;
	wire w_dff_A_vt49kmHw4_1;
	wire w_dff_A_2Jr8D4s51_2;
	wire w_dff_B_HwTHqegq0_1;
	wire w_dff_B_xpsKkW372_1;
	wire w_dff_A_b6RVrugm3_1;
	wire w_dff_A_7pDiKzB21_2;
	wire w_dff_A_yblqBuNC5_2;
	wire w_dff_A_avRL46u46_2;
	wire w_dff_A_1d6IbwNh2_2;
	wire w_dff_B_Opz9X0i83_0;
	wire w_dff_B_10PqCySC3_0;
	wire w_dff_B_CYWKAXAg8_0;
	wire w_dff_B_toa3xpjP1_0;
	wire w_dff_A_T8uo1aQq5_1;
	wire w_dff_A_Xi4JRTa49_1;
	wire w_dff_A_vcxg1qYh8_2;
	wire w_dff_B_rECt16696_1;
	wire w_dff_B_ss6wQMSM1_1;
	wire w_dff_B_eRaeAqzx5_1;
	wire w_dff_B_REqKySol5_1;
	wire w_dff_A_awADi5dy0_0;
	wire w_dff_A_DRU23pch3_0;
	wire w_dff_A_ErTh8wLX2_2;
	wire w_dff_A_QR5cJbr74_2;
	wire w_dff_A_MadWnhvV5_2;
	wire w_dff_A_yLA6kELO7_2;
	wire w_dff_A_9NFBB2sh2_2;
	wire w_dff_B_cQDb0x8w8_0;
	wire w_dff_A_Td2GGZBJ4_1;
	wire w_dff_B_WSAyDDDI9_1;
	wire w_dff_B_A0x9HqyM7_1;
	wire w_dff_B_yaVOpD0p0_1;
	wire w_dff_A_Cf3iR7zw1_0;
	wire w_dff_A_IfVgLIMX6_0;
	wire w_dff_A_kk0bhBUK1_0;
	wire w_dff_A_CEzkFtCv3_0;
	wire w_dff_A_KkTi9hGO7_0;
	wire w_dff_A_72xvU02r3_0;
	wire w_dff_A_PF283EE86_0;
	wire w_dff_A_H0XydCmF2_0;
	wire w_dff_A_ZZIjx8KE4_0;
	wire w_dff_B_Xt38zowO9_1;
	wire w_dff_B_VnAYDJq25_1;
	wire w_dff_B_b6ipeSB23_0;
	wire w_dff_B_wffm9AH96_1;
	wire w_dff_A_RtYubszG9_0;
	wire w_dff_A_VN574AsW8_0;
	wire w_dff_A_aPNn3EpD9_0;
	wire w_dff_B_9JCi7FQT0_0;
	wire w_dff_B_WxuNFnKF1_0;
	wire w_dff_B_AGGp1nRs5_0;
	wire w_dff_B_UN52YtQS4_0;
	wire w_dff_B_vWa9fJa06_0;
	wire w_dff_B_YwhNRbe39_0;
	wire w_dff_B_zPEJRzuL7_0;
	wire w_dff_B_GFUvPOFf8_0;
	wire w_dff_B_XYEEje5n4_1;
	wire w_dff_A_Rh403l8r6_0;
	wire w_dff_A_vaJNcwWB3_0;
	wire w_dff_A_5Ty3TnsM0_0;
	wire w_dff_A_2AzRzcU75_0;
	wire w_dff_A_vW7RpPeh6_0;
	wire w_dff_A_Uldg6yWl3_0;
	wire w_dff_A_ZrG1LffZ7_0;
	wire w_dff_A_AkhiEvVQ8_0;
	wire w_dff_A_9Co6SrCG3_0;
	wire w_dff_A_yo2xpoMC5_0;
	wire w_dff_A_ocxPA7mX1_0;
	wire w_dff_A_tS7MsuFi0_1;
	wire w_dff_A_AA3gEA2K1_1;
	wire w_dff_A_NH8R1pZz6_1;
	wire w_dff_A_Moh5KKKy7_1;
	wire w_dff_A_ydAqYyKh0_1;
	wire w_dff_A_PCx2iXYg6_1;
	wire w_dff_A_w8cy5tjY3_1;
	wire w_dff_A_GhLDPFKD8_1;
	wire w_dff_A_VJgypklu9_1;
	wire w_dff_A_TePc5rIr7_1;
	wire w_dff_A_1psSUxf49_1;
	wire w_dff_B_5F7UX6Mj8_0;
	wire w_dff_B_hfXWDO4K3_0;
	wire w_dff_B_rFZsDiXU3_1;
	wire w_dff_B_Ien3t5Ck6_1;
	wire w_dff_B_0km3CmbJ7_1;
	wire w_dff_A_zU3v8NVp9_0;
	wire w_dff_A_E8QLvYZR7_0;
	wire w_dff_A_j65Yf79E8_0;
	wire w_dff_A_rKyVvHD16_0;
	wire w_dff_B_ksfw1szy2_2;
	wire w_dff_B_Ct5oodQI2_1;
	wire w_dff_A_uvenekGE3_1;
	wire w_dff_B_hDRpT2tv7_3;
	wire w_dff_B_yS6MQTAQ7_3;
	wire w_dff_B_UP0PQyuR2_3;
	wire w_dff_B_GzK86MKc0_1;
	wire w_dff_B_SFYn7sTX4_1;
	wire w_dff_B_AVdJ0gQA0_0;
	wire w_dff_A_PmkHxSYn8_0;
	wire w_dff_A_1OACN2q06_0;
	wire w_dff_A_ntj8JBwS3_0;
	wire w_dff_A_hRJp7vWr2_0;
	wire w_dff_A_DDmYIJHw9_0;
	wire w_dff_A_ElC4w09o7_0;
	wire w_dff_A_9DxxuXB93_1;
	wire w_dff_A_Ri7ncHCl4_1;
	wire w_dff_A_13LBD0XT5_1;
	wire w_dff_A_TiXB0ib65_2;
	wire w_dff_B_qMMpENxz7_0;
	wire w_dff_B_ojiNcVtd8_0;
	wire w_dff_B_f6176n3t8_0;
	wire w_dff_B_gAgA76Jv1_0;
	wire w_dff_B_mCIk2dZs8_0;
	wire w_dff_A_c60IsobB1_0;
	wire w_dff_A_CZjEQc8K0_1;
	wire w_dff_A_tpiQOmRR1_1;
	wire w_dff_A_dbW3SnzF1_1;
	wire w_dff_A_WrqDm6nI6_1;
	wire w_dff_A_XV4Q8hST0_1;
	wire w_dff_A_XsYOkWAa1_1;
	wire w_dff_A_ZRods4mx6_1;
	wire w_dff_A_oNuluRoW1_1;
	wire w_dff_B_2zO82OCK7_1;
	wire w_dff_B_tHyOvIpT5_1;
	wire w_dff_A_YvrL0TOD8_1;
	wire w_dff_A_i6KgicKk7_1;
	wire w_dff_A_EilZvoQR7_1;
	wire w_dff_B_bxIqVvov8_1;
	wire w_dff_B_eQWyAsEn2_0;
	wire w_dff_B_62Ls3ksn7_1;
	wire w_dff_A_UZUteTL87_0;
	wire w_dff_A_AzQ9Rfkm7_0;
	wire w_dff_B_shsYs3545_2;
	wire w_dff_B_Q1nhhtqB4_0;
	wire w_dff_B_5pQ1P8OX7_1;
	wire w_dff_A_oCDmwxQd4_1;
	wire w_dff_A_r1xFQf2C4_1;
	wire w_dff_A_UjOJvMcG4_0;
	wire w_dff_A_s56N452h0_1;
	wire w_dff_A_2v5adAyr4_2;
	wire w_dff_A_o0jD4GnU1_0;
	wire w_dff_A_5gjoHNAA6_1;
	wire w_dff_A_knkxMSEg2_2;
	wire w_dff_A_0jrw4gfZ6_1;
	wire w_dff_A_R35VlzGe6_1;
	wire w_dff_B_jIhpRT4v7_2;
	wire w_dff_B_6kMIKriX5_2;
	wire w_dff_B_V5R8BYO09_1;
	wire w_dff_B_7nl7DOtC1_1;
	wire w_dff_B_ZN7OJbMQ8_0;
	wire w_dff_B_P3RPMK2f3_0;
	wire w_dff_B_DPEIDd9G1_0;
	wire w_dff_B_UcOqa7wm6_0;
	wire w_dff_B_dBM934nq7_0;
	wire w_dff_B_9KRF2h341_0;
	wire w_dff_B_x2J2RxHQ3_0;
	wire w_dff_B_uSlMZpg44_1;
	wire w_dff_B_gpfmQNdc9_1;
	wire w_dff_B_WEUy2SL86_1;
	wire w_dff_B_mhOjddX57_1;
	wire w_dff_B_FWJMrzgD2_1;
	wire w_dff_B_SLq0e8Kd6_1;
	wire w_dff_A_gsN1zYW38_2;
	wire w_dff_B_xNg1sUQ42_1;
	wire w_dff_A_6ms29Wfm8_1;
	wire w_dff_B_ou8phIP07_1;
	wire w_dff_B_OwepyVfj8_1;
	wire w_dff_B_r8bLlVZ74_1;
	wire w_dff_B_ounUMgFs8_1;
	wire w_dff_B_cnDPdZq33_1;
	wire w_dff_B_hdG0pbbR9_1;
	wire w_dff_A_ImRUhdDb0_0;
	wire w_dff_A_fJJ6n7k51_0;
	wire w_dff_A_Q4XdTMH92_0;
	wire w_dff_A_s0qi0ndp0_2;
	wire w_dff_A_g49N9GbX7_1;
	wire w_dff_A_sPVdBoWT8_1;
	wire w_dff_A_klVsZxkz3_1;
	wire w_dff_A_IfxbrZjd4_2;
	wire w_dff_A_iG6SEfJ78_2;
	wire w_dff_A_uchtVzkm2_2;
	wire w_dff_B_pQFgIYcx9_1;
	wire w_dff_B_Fk6489C09_1;
	wire w_dff_B_qayTBsAn8_0;
	wire w_dff_A_kTfg7kte6_0;
	wire w_dff_B_3sc9Ecjf8_0;
	wire w_dff_B_pL18KfnZ3_1;
	wire w_dff_B_IqFXHgBs6_1;
	wire w_dff_B_wxIrUPRk3_1;
	wire w_dff_B_eBA4zMxn0_1;
	wire w_dff_B_Fxf59Ko60_1;
	wire w_dff_B_kPb1VbpD9_1;
	wire w_dff_B_YMfXw1AN3_1;
	wire w_dff_B_wmhtPQGZ2_1;
	wire w_dff_B_ApcI78CP0_1;
	wire w_dff_B_a7sBk9jl0_1;
	wire w_dff_B_ySXOopji0_0;
	wire w_dff_A_uuXYZh7f9_0;
	wire w_dff_A_aeBcOHkp3_0;
	wire w_dff_A_nI7djk5b5_0;
	wire w_dff_A_Gt3uamDq6_2;
	wire w_dff_B_orJoUx8x2_1;
	wire w_dff_B_b8Fn2muT3_1;
	wire w_dff_B_hiwWDqOG1_1;
	wire w_dff_B_In3jeXyT8_1;
	wire w_dff_B_VjYy4XQB0_1;
	wire w_dff_B_7fAGyRMk1_0;
	wire w_dff_A_3aHxw2DG4_1;
	wire w_dff_A_7Mu1Dhco8_1;
	wire w_dff_A_lFUaObDu7_0;
	wire w_dff_A_DdNK124j6_0;
	wire w_dff_A_6VGMMbyj4_0;
	wire w_dff_B_cWK7IIex0_0;
	wire w_dff_B_FDvsbCPd3_0;
	wire w_dff_A_P5A958rJ9_1;
	wire w_dff_A_0QAog1zj5_1;
	wire w_dff_A_PJ6xGTsY9_1;
	wire w_dff_A_gGJ6Bts46_1;
	wire w_dff_B_4U45jzSB5_0;
	wire w_dff_B_PJ66t5yM2_0;
	wire w_dff_B_Uf0XxWAg0_0;
	wire w_dff_A_fGNBHnwj8_1;
	wire w_dff_A_nnTQgwfk1_1;
	wire w_dff_B_XjXOnsmf3_0;
	wire w_dff_B_6esktB4V4_1;
	wire w_dff_B_dDHsSDnA9_1;
	wire w_dff_B_zT8eHC0d9_1;
	wire w_dff_B_hjXK9s2E9_1;
	wire w_dff_B_1bIJ8zSE5_1;
	wire w_dff_B_ufJdp9e54_1;
	wire w_dff_B_RQ0tSwua1_1;
	wire w_dff_B_VQ8gnLiz2_0;
	wire w_dff_A_t8N1d5Pb7_0;
	wire w_dff_B_YSJ6bEhz9_1;
	wire w_dff_A_bKy6J2rE7_0;
	wire w_dff_A_gM5IJcWt1_0;
	wire w_dff_A_xkJlU7Il1_0;
	wire w_dff_A_2QxankVB8_2;
	wire w_dff_A_9qQuyDoI6_2;
	wire w_dff_A_quOWGrrx4_2;
	wire w_dff_A_0y1D0MhM1_2;
	wire w_dff_B_CF3vVTP54_3;
	wire w_dff_B_57chmTx82_3;
	wire w_dff_B_1WN0ZySe4_3;
	wire w_dff_B_BdpCwJC28_1;
	wire w_dff_A_zT8TQK0W9_1;
	wire w_dff_B_ThHvDAIp5_3;
	wire w_dff_B_ArM46iT91_3;
	wire w_dff_B_szlZOZXh5_3;
	wire w_dff_B_MpMlUWve7_1;
	wire w_dff_B_rU4T2go71_1;
	wire w_dff_B_tmSYz4yx9_1;
	wire w_dff_B_5iAuwOLi4_1;
	wire w_dff_B_1IAQThCU0_1;
	wire w_dff_A_HEyFGdAl1_1;
	wire w_dff_B_T5V9d2Bh4_1;
	wire w_dff_A_N8zkPk2V5_0;
	wire w_dff_A_v8vdYEFd9_0;
	wire w_dff_A_4UGmj34i8_0;
	wire w_dff_A_f7y5WgPL4_0;
	wire w_dff_A_nXgID33p2_0;
	wire w_dff_A_pzRQG86f7_0;
	wire w_dff_A_hW8AAyM75_0;
	wire w_dff_A_k6m6EGB75_2;
	wire w_dff_A_0EEZjhwS3_2;
	wire w_dff_A_odTVlco66_2;
	wire w_dff_A_kQVuwrPh6_2;
	wire w_dff_A_SuGQnfHG3_2;
	wire w_dff_A_0etCkqs48_2;
	wire w_dff_B_fW4BpqX15_1;
	wire w_dff_B_2ANOq5n72_1;
	wire w_dff_B_Fxsrb80G4_0;
	wire w_dff_A_S3wOPQv49_0;
	wire w_dff_B_Xy3Tfcgg6_0;
	wire w_dff_A_EQTcbEZH4_1;
	wire w_dff_A_8vmb2NwO7_1;
	wire w_dff_A_e0QIJYxy9_1;
	wire w_dff_A_cetJO7la0_1;
	wire w_dff_A_07Ru6seW5_1;
	wire w_dff_A_zrrb1dWY3_1;
	wire w_dff_A_jzGcGysS2_1;
	wire w_dff_A_NMgCCs5d2_1;
	wire w_dff_A_YNwvWcum7_1;
	wire w_dff_A_JsZ5AxpJ8_1;
	wire w_dff_A_h4H1DHsB8_1;
	wire w_dff_A_HfBoGHCo1_1;
	wire w_dff_A_edMqENaC1_2;
	wire w_dff_A_dPPxc8oq7_2;
	wire w_dff_A_FYxxkD401_2;
	wire w_dff_A_oZO6c03a0_2;
	wire w_dff_A_7ljpYLmB9_0;
	wire w_dff_A_dXgb7lB73_0;
	wire w_dff_A_3AJGYNJi7_0;
	wire w_dff_A_8e3u4AU77_0;
	wire w_dff_A_VCu3sJlL1_0;
	wire w_dff_B_nKDuQ6uv3_0;
	wire w_dff_B_8GrNoiK39_0;
	wire w_dff_A_CAZW4RVx2_2;
	wire w_dff_A_qAWZsXJr4_2;
	wire w_dff_A_eTQddzzA9_2;
	wire w_dff_A_PVE1CDEL4_2;
	wire w_dff_A_F23E7Z5V8_2;
	wire w_dff_A_rPtILABT7_2;
	wire w_dff_A_pgcBG5UC7_2;
	wire w_dff_A_OghlpeEH0_2;
	wire w_dff_A_BcrQTTm06_2;
	wire w_dff_B_Y8wnFUcd0_0;
	wire w_dff_B_1ymcwVnc5_0;
	wire w_dff_B_bnEJzStn0_0;
	wire w_dff_B_01GKseaG2_0;
	wire w_dff_B_kBTgxbTc6_0;
	wire w_dff_B_ThDjJH2c2_0;
	wire w_dff_B_lRcnW8Hx2_0;
	wire w_dff_B_ZuP8Rk7Z9_1;
	wire w_dff_B_N8VLJqyG2_1;
	wire w_dff_B_VkhJlcVA1_1;
	wire w_dff_B_9sPCvJLp1_0;
	wire w_dff_B_qpxD3fEa0_0;
	wire w_dff_B_3E0Ul3YV3_0;
	wire w_dff_A_V6O6VTJa3_1;
	wire w_dff_A_Ye7xy3Ka0_1;
	wire w_dff_A_ujABWE8i1_2;
	wire w_dff_A_G8EXsN8I4_2;
	wire w_dff_A_AqxmzgaN0_2;
	wire w_dff_A_hCY0c5F84_2;
	wire w_dff_A_4csDuuaN6_2;
	wire w_dff_A_R8bxaq8C7_2;
	wire w_dff_A_kBcCz6HL9_2;
	wire w_dff_A_tF8vX1f22_2;
	wire w_dff_B_Ln9ZbyCK9_0;
	wire w_dff_B_f9OO8QL00_0;
	wire w_dff_A_sGUw0pmT6_1;
	wire w_dff_B_dVKmhsVS6_0;
	wire w_dff_A_6b1FezRd7_0;
	wire w_dff_A_Gus10aQ47_0;
	wire w_dff_A_8DYJNc5I8_1;
	wire w_dff_A_aFrgECxh2_1;
	wire w_dff_A_sM4oKHqN0_1;
	wire w_dff_A_eoF0XVMH7_2;
	wire w_dff_A_73qoDkLk9_2;
	wire w_dff_A_OnZNoG9q7_0;
	wire w_dff_A_SpIpFv3q9_0;
	wire w_dff_A_72t6ETG10_1;
	wire w_dff_A_X1tZQeR31_1;
	wire w_dff_A_Og5MRb3q7_2;
	wire w_dff_A_L5KZjV4q2_2;
	wire w_dff_A_sEVsS5Ua6_2;
	wire w_dff_A_pGqw67Fc1_1;
	wire w_dff_A_sAcMoqNB6_1;
	wire w_dff_A_FH96tEjZ0_1;
	wire w_dff_A_VMOJjKVJ3_1;
	wire w_dff_B_CdPONrv61_0;
	wire w_dff_B_Lc4vOZKj4_0;
	wire w_dff_B_BxPg4YKO0_1;
	wire w_dff_B_7ENqnbhr4_1;
	wire w_dff_B_wjSu0zAU3_1;
	wire w_dff_B_hVb0CsHc0_1;
	wire w_dff_B_5iePj3C97_0;
	wire w_dff_A_ymCLt7bK8_1;
	wire w_dff_A_gqd75nBO0_1;
	wire w_dff_A_maskZQOy6_1;
	wire w_dff_A_qCiB9QtQ7_1;
	wire w_dff_A_EjlM9Hnm1_1;
	wire w_dff_A_M6yMn2DP4_2;
	wire w_dff_A_V4Oy8Dsb1_2;
	wire w_dff_B_VPxtV2Dm3_1;
	wire w_dff_B_RSXJqNCL9_1;
	wire w_dff_A_VexwC1p14_1;
	wire w_dff_B_9z8F1Thl9_1;
	wire w_dff_B_DDUoAJAO2_1;
	wire w_dff_B_ml9GC6oQ8_0;
	wire w_dff_B_7bU8Sqr96_0;
	wire w_dff_B_HALy3Khn7_1;
	wire w_dff_A_67XSxAJS6_1;
	wire w_dff_A_YVUJFrSK3_0;
	wire w_dff_A_cZPzdJwJ2_1;
	wire w_dff_B_yVxTtLLJ4_3;
	wire w_dff_B_fxZ7pw9z2_3;
	wire w_dff_A_u86Ibo975_0;
	wire w_dff_A_6bLnyUtW9_0;
	wire w_dff_A_AU5f9WES5_0;
	wire w_dff_A_OeXoWeOW9_1;
	wire w_dff_A_TttI0QSF7_1;
	wire w_dff_A_tzRFdULo5_1;
	wire w_dff_A_BcUIqjLa9_1;
	wire w_dff_A_GJ0JER405_0;
	wire w_dff_A_8PYxwOD49_1;
	wire w_dff_A_z1JNQAMu2_1;
	wire w_dff_A_QAlOaucd4_2;
	wire w_dff_B_S1TWYexl9_1;
	wire w_dff_B_qO6l6Hji1_1;
	wire w_dff_A_TE9mGCgW0_1;
	wire w_dff_A_4lNsKam10_1;
	wire w_dff_A_NG3RrSe38_1;
	wire w_dff_A_jJQgm6LR5_2;
	wire w_dff_A_XElAkDnA6_2;
	wire w_dff_A_sKmGXIaU0_2;
	wire w_dff_A_9LWVJ9J94_2;
	wire w_dff_A_RMo9H0qy0_1;
	wire w_dff_A_VOJ3Gx0C6_1;
	wire w_dff_A_XF5SPZMu9_1;
	wire w_dff_A_w4f6Aana9_1;
	wire w_dff_A_CzPuB0WY5_1;
	wire w_dff_A_SmDPUhHV2_0;
	wire w_dff_A_F1LSShtC4_0;
	wire w_dff_A_vXOkiJ2b4_2;
	wire w_dff_A_E72xmQJQ7_2;
	wire w_dff_A_7L8arQuy9_0;
	wire w_dff_A_zQ0aq7wq3_0;
	wire w_dff_A_X4weM8Cq6_2;
	wire w_dff_A_IQpk0kVG8_2;
	wire w_dff_A_7lY5Beui3_2;
	wire w_dff_A_4zFnBeeD1_1;
	wire w_dff_A_XsDSl20W7_1;
	wire w_dff_A_DB0ardjG5_1;
	wire w_dff_A_VRH3paYD6_1;
	wire w_dff_A_9YxXXqlF6_2;
	wire w_dff_A_krrjJfzj6_2;
	wire w_dff_A_vViKNCfp1_2;
	wire w_dff_A_VrIy1Jep0_2;
	wire w_dff_A_1poxb7it2_2;
	wire w_dff_A_C1NEEAJW6_2;
	wire w_dff_A_toS1cSfk5_2;
	wire w_dff_A_W2tX3q3y2_2;
	wire w_dff_A_3NM5qXvP7_2;
	wire w_dff_A_bVZSU6GH8_1;
	wire w_dff_A_1JsX1pGC1_1;
	wire w_dff_A_mG4NQv9y8_0;
	wire w_dff_A_lFlKgL0f6_1;
	wire w_dff_A_AD8s80ZX9_1;
	wire w_dff_B_lsLzXNMs1_0;
	wire w_dff_A_XqsxgXkg9_0;
	wire w_dff_A_qiJW42G68_0;
	wire w_dff_A_3xum2mTS6_1;
	wire w_dff_A_Hi8ULcd96_1;
	wire w_dff_A_FA6PyYmV0_1;
	wire w_dff_A_DAWbyz9E8_1;
	wire w_dff_A_i4C8CJMS1_1;
	wire w_dff_B_mRBBmtHJ5_0;
	wire w_dff_B_dlM9eFUA4_0;
	wire w_dff_A_PDfB6XMd4_1;
	wire w_dff_A_uiIIcp3f6_1;
	wire w_dff_A_25sVWHOy3_1;
	wire w_dff_A_H4ms9W386_1;
	wire w_dff_A_7dtRq2NS9_1;
	wire w_dff_A_yrHzOZpB0_0;
	wire w_dff_B_F4cGoxfX8_1;
	wire w_dff_B_ei1IRPYu3_1;
	wire w_dff_B_O8VhvD2i9_1;
	wire w_dff_A_SG9uoOXf1_1;
	wire w_dff_A_rDmAkkS04_2;
	wire w_dff_B_1RzhudOz1_1;
	wire w_dff_B_llEH8sKq5_1;
	wire w_dff_A_gRveNVBj0_2;
	wire w_dff_A_QfY9ycPs7_1;
	wire w_dff_A_nNSVdi6V0_2;
	wire w_dff_A_rxnjzVgC9_0;
	wire w_dff_A_xSMk7Iu53_0;
	wire w_dff_A_Qsh7UEam8_0;
	wire w_dff_A_LS8Kd3zY6_1;
	wire w_dff_A_NH0586Nw4_1;
	wire w_dff_B_uHyrMRuq9_0;
	wire w_dff_A_Mfoln7al3_1;
	wire w_dff_A_JD62UApS0_1;
	wire w_dff_B_BKOW30cU3_1;
	wire w_dff_A_xSfVpV0A9_2;
	wire w_dff_A_PPac0J2D5_2;
	wire w_dff_A_jOenf4jn0_1;
	wire w_dff_A_jFkwn7bH5_1;
	wire w_dff_A_PfwbTdmM6_1;
	wire w_dff_A_BXQjOJiv0_1;
	wire w_dff_A_Deq1UrMn3_2;
	wire w_dff_A_AZmo76qN7_2;
	wire w_dff_A_PxFH9qKR2_0;
	wire w_dff_A_JSngJh1o7_0;
	wire w_dff_A_lbfPEgwu3_2;
	wire w_dff_A_aUuFFNoZ0_2;
	wire w_dff_A_C6fhdDYB1_1;
	wire w_dff_A_vSQVX5kt8_0;
	wire w_dff_A_kHyPVeGO3_0;
	wire w_dff_A_eHGMUOgQ9_0;
	wire w_dff_A_bXF8Ko468_0;
	wire w_dff_A_v2s6uZoF7_0;
	wire w_dff_A_tnk2iPlc2_1;
	wire w_dff_A_66o4pQgu8_1;
	wire w_dff_A_gH22s1fJ8_0;
	wire w_dff_A_nKjGZzcD3_0;
	wire w_dff_A_9TorVuzk2_0;
	wire w_dff_A_A8RKeC036_0;
	wire w_dff_A_STf4gIso3_0;
	wire w_dff_A_VRn3UZHx9_0;
	wire w_dff_A_3gRB1EJk6_0;
	wire w_dff_A_78XtRBs74_0;
	wire w_dff_A_NC3D814C8_1;
	wire w_dff_A_5hmUbngm0_1;
	wire w_dff_A_r7coMN1H0_1;
	wire w_dff_A_uDbIhnhQ0_1;
	wire w_dff_B_Z5BUScwi0_0;
	wire w_dff_B_teAz4mHt2_1;
	wire w_dff_A_tbzq0ca04_0;
	wire w_dff_A_WZhaYv5b6_1;
	wire w_dff_A_QrqwqCbg4_1;
	wire w_dff_A_jWhzem8v7_2;
	wire w_dff_A_k0Hrm9on7_2;
	wire w_dff_A_1YteJ72n8_1;
	wire w_dff_A_Ae8V3D2h6_0;
	wire w_dff_A_F49VzkO16_2;
	wire w_dff_A_ibTsKWpo0_2;
	wire w_dff_A_NUaPsx8q7_0;
	wire w_dff_A_us0AcsJW6_0;
	wire w_dff_A_ZwN0FY9s9_0;
	wire w_dff_A_PhnE6QKk6_0;
	wire w_dff_A_oaqMv60T3_1;
	wire w_dff_A_gsERAYf14_1;
	wire w_dff_A_ZW7DFe3L2_0;
	wire w_dff_A_kt8vfdUT2_1;
	wire w_dff_A_EgbFodsF6_1;
	wire w_dff_A_Bn1ER3N95_1;
	wire w_dff_A_IWTwbYrN4_2;
	wire w_dff_A_aSoHVQ5s5_2;
	wire w_dff_A_h7ftODI60_1;
	wire w_dff_A_U3CmrLaq8_1;
	wire w_dff_A_HOhlGm5x4_0;
	wire w_dff_A_UjEXtY9A0_1;
	wire w_dff_A_93Zd3l2g8_1;
	wire w_dff_A_tgNieMpj3_0;
	wire w_dff_A_Ns6FvkDn8_0;
	wire w_dff_A_aXlyl3Fd0_0;
	wire w_dff_A_xYXY8fqB5_1;
	wire w_dff_A_AwnHk9988_1;
	wire w_dff_A_YcSEk4u81_0;
	wire w_dff_A_2yVxaMzY3_1;
	wire w_dff_A_oRkKDqT53_1;
	wire w_dff_A_7U1UTgYe7_2;
	wire w_dff_A_NS8jNmWs2_2;
	wire w_dff_A_O7ejGNVk3_1;
	wire w_dff_A_CecK2pIg7_2;
	wire w_dff_A_upzh20eh1_2;
	wire w_dff_A_CAWMciHy2_0;
	wire w_dff_A_Q2LPEikI5_0;
	wire w_dff_A_b1wPHBan4_0;
	wire w_dff_A_LsbrMTkE4_0;
	wire w_dff_A_60vNIaI08_1;
	wire w_dff_A_WxdUJPLt4_1;
	wire w_dff_A_hDEczb3X8_0;
	wire w_dff_B_vHNzx2Rh3_0;
	wire w_dff_A_9bQoZvaZ9_2;
	wire w_dff_B_FIelMW6t1_0;
	wire w_dff_B_2DsSV5zE4_0;
	wire w_dff_B_w9d2YWfE9_0;
	wire w_dff_A_7UwZUzIm3_0;
	wire w_dff_A_iQuhWqzD7_0;
	wire w_dff_A_Ild9kzuP5_1;
	wire w_dff_A_eM79DCKB4_1;
	wire w_dff_A_96MVLQZu7_2;
	wire w_dff_A_Jz9hUAx84_2;
	wire w_dff_B_7cE0JC4U6_3;
	wire w_dff_B_i6tp0XE54_3;
	wire w_dff_B_Q838d2J84_3;
	wire w_dff_B_xJUEBMqN3_3;
	wire w_dff_B_kxKU4Zyf9_3;
	wire w_dff_A_0qCPDfMR7_1;
	wire w_dff_A_APNkAsNs8_1;
	wire w_dff_A_TRlDMbyE9_1;
	wire w_dff_A_OzLmUVZf7_1;
	wire w_dff_A_FurO07le1_1;
	wire w_dff_A_ogos4tL26_1;
	wire w_dff_A_Me1fhYuZ2_0;
	wire w_dff_A_uNIKy0Cp2_1;
	wire w_dff_A_ZMKhAMUR0_1;
	wire w_dff_A_HDWYnpOB9_2;
	wire w_dff_A_1279TGH46_1;
	wire w_dff_A_TfJltKmd2_1;
	wire w_dff_A_9a3Em77c0_1;
	wire w_dff_A_gBaa83Ed2_1;
	wire w_dff_A_fS0LlvZK6_1;
	wire w_dff_A_2WoCuG5J3_1;
	wire w_dff_B_VZM5CY1Z9_1;
	wire w_dff_A_5HXFfcAo9_1;
	wire w_dff_B_yMYeWhuq7_1;
	wire w_dff_B_mypaOipd7_1;
	wire w_dff_A_OlooEsLk1_0;
	wire w_dff_A_MDqOfozP8_2;
	wire w_dff_B_AiBGyhXP0_0;
	wire w_dff_B_8kuGAAZk2_1;
	wire w_dff_A_qAdhCfa83_1;
	wire w_dff_A_zY3WHwLO9_0;
	wire w_dff_B_LiSmy9oS4_0;
	wire w_dff_A_vevyfFaW1_0;
	wire w_dff_A_UYDQdNuH7_1;
	wire w_dff_A_E8cAH0dG6_1;
	wire w_dff_A_bRRjJPyT6_1;
	wire w_dff_A_REIo9ffo7_0;
	wire w_dff_A_Z1rKLJEN2_2;
	wire w_dff_A_c6nYiNQz8_1;
	wire w_dff_A_oAkhjJVX7_2;
	wire w_dff_A_T7sl5B3r6_0;
	wire w_dff_A_O35QWYi73_0;
	wire w_dff_A_WdejfyvY0_1;
	wire w_dff_A_aaQzLjKd6_1;
	wire w_dff_A_nANvYK136_1;
	wire w_dff_A_38YAPIYS1_0;
	wire w_dff_A_TIDzhtUv3_0;
	wire w_dff_A_TwV63DNe3_1;
	wire w_dff_A_J55No7Ox2_1;
	wire w_dff_A_iqzJtzSj0_0;
	wire w_dff_A_aLVZsU2V1_0;
	wire w_dff_A_b8n47nWS4_0;
	wire w_dff_A_GRRwwvD30_2;
	wire w_dff_B_wjJvFzl57_3;
	wire w_dff_B_bN40Ll332_3;
	wire w_dff_B_vmS78ivG2_3;
	wire w_dff_B_H7cRpZho8_3;
	wire w_dff_B_By5IOUUi6_3;
	wire w_dff_B_KU0nt64i4_3;
	wire w_dff_A_ihw0ivVJ5_0;
	wire w_dff_A_C61XykJj3_0;
	wire w_dff_B_JgsaM3to7_2;
	wire w_dff_B_Ig6Xmlhb8_2;
	wire w_dff_B_EwQVB6tX8_2;
	wire w_dff_B_DqFvCkPD9_2;
	wire w_dff_B_0I1CikA97_1;
	wire w_dff_B_gI3qsLLX6_0;
	wire w_dff_B_VRcvTawS5_0;
	wire w_dff_B_kPQnTKnU7_0;
	wire w_dff_B_cEH9gJjW1_0;
	wire w_dff_B_DDLmV1sL9_0;
	wire w_dff_A_mBfYHKxY7_0;
	wire w_dff_A_SmwWHC6v9_0;
	wire w_dff_A_Zg11fxW30_0;
	wire w_dff_A_vkCkv83m6_0;
	wire w_dff_A_aRrmc5Aj4_0;
	wire w_dff_A_QedZhUyP9_0;
	wire w_dff_A_PMwywllJ0_0;
	wire w_dff_A_5yT7bRBN7_1;
	wire w_dff_A_QZArltnf9_1;
	wire w_dff_A_BXgTb1ev9_1;
	wire w_dff_A_PGw1wZYf4_1;
	wire w_dff_A_z7nYyzmH2_1;
	wire w_dff_A_3oPoLBjJ4_0;
	wire w_dff_A_h1B3mJfH4_2;
	wire w_dff_A_LdOBTXp65_2;
	wire w_dff_A_VjANystY2_2;
	wire w_dff_A_TZCEIUvz2_0;
	wire w_dff_A_hHIrK42a3_0;
	wire w_dff_A_z5eoBffp8_0;
	wire w_dff_A_ykQuhNr48_0;
	wire w_dff_A_Ga9HDaAh5_0;
	wire w_dff_A_LArgObzU8_0;
	wire w_dff_A_kB4WD2uz7_1;
	wire w_dff_A_XEMYXWQY2_1;
	wire w_dff_A_so2b6Mk06_1;
	wire w_dff_A_Jw4UgDiI5_2;
	wire w_dff_A_8EDbM3VO1_2;
	wire w_dff_A_YdIp8JhS8_2;
	wire w_dff_A_Tev3nFhw1_1;
	wire w_dff_A_hIrgyG9Q4_1;
	wire w_dff_A_eqyl31wS2_2;
	wire w_dff_A_n1QeoCI66_2;
	wire w_dff_A_V8PP1KKa7_2;
	wire w_dff_A_nmcIZyGl1_2;
	wire w_dff_A_8SqCKDX28_0;
	wire w_dff_A_Yu5PzgA72_0;
	wire w_dff_A_kVVVfSmH2_0;
	wire w_dff_A_ObjgFuti1_0;
	wire w_dff_A_98rMngqj2_2;
	wire w_dff_A_0BCjYyTD0_1;
	wire w_dff_A_yOUXbtIP7_1;
	wire w_dff_A_1FSyIZIT2_0;
	wire w_dff_B_bMygN5jQ5_1;
	wire w_dff_B_eXnXffhz6_1;
	wire w_dff_B_NI5hjL856_1;
	wire w_dff_B_wHCIhoNy1_1;
	wire w_dff_A_UKI5si2f1_2;
	wire w_dff_A_Qo9GQida4_2;
	wire w_dff_A_4dQJKf2J1_2;
	wire w_dff_A_EhOeGe6S7_2;
	wire w_dff_A_SxkNvj3H7_2;
	wire w_dff_A_j14lyMv84_2;
	wire w_dff_A_GYJ1jS5R7_2;
	wire w_dff_A_KgkWMurd5_2;
	wire w_dff_A_D9G1yZ2a1_0;
	wire w_dff_A_SIvmIlwI9_0;
	wire w_dff_A_UFHF0I219_0;
	wire w_dff_A_9KKD5hdf2_0;
	wire w_dff_A_MZfX7DFR6_0;
	wire w_dff_A_57ZRTMa09_0;
	wire w_dff_A_PVZi9aMd7_1;
	wire w_dff_A_a4I94ztY4_1;
	wire w_dff_A_ZslAtP5G6_1;
	wire w_dff_A_iVfLRPJb5_0;
	wire w_dff_A_3Ekhpmm29_0;
	wire w_dff_A_LPoGvtSe4_1;
	wire w_dff_A_wUc9r8FB4_1;
	wire w_dff_A_acbnPoFk7_1;
	wire w_dff_A_165wfq2N1_0;
	wire w_dff_A_KkFJ5Hfk9_1;
	wire w_dff_A_Ukt0XTUJ4_1;
	wire w_dff_A_EiFIn5iG2_1;
	wire w_dff_A_aC0WX6qI9_1;
	wire w_dff_A_54F53hGA1_0;
	wire w_dff_A_fXJA9ANq0_2;
	wire w_dff_A_0ZrkUSCb5_2;
	wire w_dff_A_pbAlY6TH8_2;
	wire w_dff_A_vd9Cswqp1_0;
	wire w_dff_A_zHuTCMKi6_1;
	wire w_dff_A_bqMO1Dy82_1;
	wire w_dff_A_XaU3ZVoN5_1;
	wire w_dff_A_VxkHbEoJ1_0;
	wire w_dff_A_9v9LOQ0m0_1;
	wire w_dff_A_jTYMQv605_1;
	wire w_dff_A_vAwRVnA50_1;
	wire w_dff_A_6yFqqlZp9_1;
	wire w_dff_A_9wmDGhK17_2;
	wire w_dff_A_OgC0qXEc7_2;
	wire w_dff_A_h72eUwTZ4_2;
	wire w_dff_A_kCrYY3sM9_1;
	wire w_dff_A_9KiZmsk92_1;
	wire w_dff_A_6Trf0unK8_1;
	wire w_dff_A_UECuCKLI4_1;
	wire w_dff_A_bm8Y9ewL9_1;
	wire w_dff_A_d3NLE3HZ0_1;
	wire w_dff_A_zVBPWxrM0_1;
	wire w_dff_A_6mxnApiT3_1;
	wire w_dff_A_5qPU88WJ5_1;
	wire w_dff_A_xLUenMFY1_1;
	wire w_dff_A_ygevY0Ts1_1;
	wire w_dff_A_XlRzNeBV1_1;
	wire w_dff_A_PA2EIylc3_1;
	wire w_dff_A_YpPsNNyi0_1;
	wire w_dff_A_KHRD8akD2_1;
	wire w_dff_A_0f2aY4Fl4_1;
	wire w_dff_A_kzmIfMe73_1;
	wire w_dff_A_UpoNaDfn7_1;
	wire w_dff_A_eXb4slFv4_1;
	wire w_dff_A_0vEhVMaq7_1;
	wire w_dff_A_1t4dqa8B4_1;
	wire w_dff_A_ofAzEnEg9_1;
	wire w_dff_A_SQbxlJ3h6_1;
	wire w_dff_A_1y3mWi0F2_1;
	wire w_dff_A_cl3wp3JZ1_1;
	wire w_dff_A_a77xGqki2_1;
	wire w_dff_A_CLpnZf594_1;
	wire w_dff_A_CHwOrggI4_1;
	wire w_dff_A_1t47kqJw6_1;
	wire w_dff_A_RVQRq0Pq2_1;
	wire w_dff_A_Pog6FL2u0_2;
	wire w_dff_A_VILqyT0n7_2;
	wire w_dff_A_KDRBfgLl1_2;
	wire w_dff_A_3tiSyFd27_2;
	wire w_dff_A_DIw65otO6_2;
	wire w_dff_A_74qqsdmk8_2;
	wire w_dff_A_BKSTxEcr2_2;
	wire w_dff_A_3krxqJlc2_2;
	wire w_dff_A_aVbwgv255_1;
	wire w_dff_A_gKi8yo9w2_1;
	wire w_dff_A_fGufZ8pH1_1;
	wire w_dff_B_Yr1JPm3o5_0;
	wire w_dff_B_ICvUMYKM8_0;
	wire w_dff_B_BFrZPIXe7_1;
	wire w_dff_B_RP6BSa9O4_1;
	wire w_dff_B_HHMlweB50_1;
	wire w_dff_B_vPFDHvJh1_1;
	wire w_dff_B_fjFwbOIT9_0;
	wire w_dff_A_FScjjiaP9_0;
	wire w_dff_B_kxpliCxs7_3;
	wire w_dff_B_ANkkWsD70_3;
	wire w_dff_B_lCwqRcNN5_3;
	wire w_dff_A_uHrmcmKh9_1;
	wire w_dff_B_iemHjl6C8_3;
	wire w_dff_B_ZpoKtMzY1_3;
	wire w_dff_B_WJf49pZb6_3;
	wire w_dff_B_6hP6nKcU1_1;
	wire w_dff_B_BHujTII25_1;
	wire w_dff_B_5q32YLO21_1;
	wire w_dff_B_X2gvFluv2_1;
	wire w_dff_B_J2PbBJUE9_0;
	wire w_dff_B_4OPNyqaq3_0;
	wire w_dff_A_3oePydcL6_0;
	wire w_dff_B_I8F6JcTl3_2;
	wire w_dff_B_UgFMn3Bk1_2;
	wire w_dff_B_lMmWfDJV8_2;
	wire w_dff_B_yj2II1H15_1;
	wire w_dff_A_7ieWbLck8_0;
	wire w_dff_A_zCo5Gg825_0;
	wire w_dff_A_cnxeaZtt8_0;
	wire w_dff_A_OzvO7sgZ4_0;
	wire w_dff_A_4gnjVid50_0;
	wire w_dff_A_NmBoDBTE5_0;
	wire w_dff_A_mOudWFRR2_0;
	wire w_dff_A_52VXOKlF3_1;
	wire w_dff_A_NbmQmMQd6_1;
	wire w_dff_A_ighade174_1;
	wire w_dff_A_eumKDIYD0_0;
	wire w_dff_B_27uRssiL8_3;
	wire w_dff_B_EjMYS9bm4_3;
	wire w_dff_B_SsOHuoV00_3;
	wire w_dff_B_myZ2XzXV4_0;
	wire w_dff_B_mqqainCH2_1;
	wire w_dff_B_PnhJcXFb8_1;
	wire w_dff_A_70XTfknm0_1;
	wire w_dff_A_toJ0YaT87_1;
	wire w_dff_A_zlDsV8Ur1_2;
	wire w_dff_A_5JEDc2PT9_2;
	wire w_dff_A_MoPl1Dqo0_2;
	wire w_dff_A_lRzML6Mb2_0;
	wire w_dff_A_mmRpLKz87_0;
	wire w_dff_A_RbkvkLIx2_1;
	wire w_dff_A_3CWmlWEH5_1;
	wire w_dff_A_X3FU8xLS8_0;
	wire w_dff_A_8LbIGvRR0_2;
	wire w_dff_A_j2vEdCQF4_2;
	wire w_dff_A_5I8oE4Ae9_2;
	wire w_dff_A_hpXedVji2_2;
	wire w_dff_A_Hd7FvtnU2_1;
	wire w_dff_A_SI4ahCmL4_0;
	wire w_dff_A_g8wPMPOg8_0;
	wire w_dff_A_BBf4G9ah5_0;
	wire w_dff_A_lz046jDm0_1;
	wire w_dff_A_tGrfnBzK0_1;
	wire w_dff_A_pPVzhuRw2_1;
	wire w_dff_A_lpyZ4Tfq1_0;
	wire w_dff_A_v4KsQ1He7_0;
	wire w_dff_A_uVJ5F7Xq3_0;
	wire w_dff_A_L4WK5rxH3_2;
	wire w_dff_A_vIZPcx7T9_2;
	wire w_dff_A_FnySFvXJ1_2;
	wire w_dff_A_FLFFGcne8_2;
	wire w_dff_A_9njr8Asa5_2;
	wire w_dff_A_4sD7ZGpF7_1;
	wire w_dff_B_X7YjN2rJ7_1;
	wire w_dff_B_gCWrTEup1_1;
	wire w_dff_A_Yzeoj65M9_0;
	wire w_dff_A_DHqjW4NS9_0;
	wire w_dff_A_F3hCORgC0_0;
	wire w_dff_A_8PNDLNEK5_1;
	wire w_dff_A_bQxUdfq12_1;
	wire w_dff_A_nVvevhsn6_1;
	wire w_dff_A_oXxWy2579_1;
	wire w_dff_A_8723l0Ow7_0;
	wire w_dff_A_YXvWWlFI9_0;
	wire w_dff_A_HlTdhWGI7_0;
	wire w_dff_A_c5YuD6Qa7_1;
	wire w_dff_A_bCRGNL845_1;
	wire w_dff_A_icJRTxbs6_1;
	wire w_dff_A_bgXHxdSP6_0;
	wire w_dff_A_ZPhdqEDj4_0;
	wire w_dff_A_YY8hlWwA5_0;
	wire w_dff_A_Rc1R6jDI9_0;
	wire w_dff_A_oo5FkNuM5_0;
	wire w_dff_A_ivs22P1q2_0;
	wire w_dff_A_BJRX0yQT4_1;
	wire w_dff_A_kNhp2yBW2_1;
	wire w_dff_A_712ULcCv3_1;
	wire w_dff_A_sdSmB09l4_1;
	wire w_dff_A_mbAwSa6M3_1;
	wire w_dff_A_FaeAKi4W3_1;
	wire w_dff_A_GaxknGMP0_1;
	wire w_dff_A_mQ3qDXyH4_1;
	wire w_dff_A_yWfi02f91_1;
	wire w_dff_A_TaJ9Tvf54_1;
	wire w_dff_A_ri80zXZg9_1;
	wire w_dff_A_HYv2t2Sc3_1;
	wire w_dff_A_Sg9pd1EJ4_1;
	wire w_dff_A_8Wqz2aeg8_1;
	wire w_dff_A_5fvJvEOG9_1;
	wire w_dff_A_muz11URF6_2;
	wire w_dff_A_YCDcsEIS3_2;
	wire w_dff_A_KrU73EEJ6_2;
	wire w_dff_A_pZOaYuK99_2;
	wire w_dff_A_ZID46GEC5_2;
	wire w_dff_A_Bts8WQCO4_2;
	wire w_dff_A_KRBhaKoL6_2;
	wire w_dff_A_bcvv62SF1_0;
	wire w_dff_A_erMOcKIW6_0;
	wire w_dff_A_XdFUXiYj2_0;
	wire w_dff_A_4FcJkg507_2;
	wire w_dff_A_IIdbkcLz0_2;
	wire w_dff_A_SSQAyeQo5_2;
	wire w_dff_A_14rTpuBW4_1;
	wire w_dff_A_vDc3UwJq2_1;
	wire w_dff_A_fMqTtTDq2_0;
	wire w_dff_A_MQ4TaRnf0_0;
	wire w_dff_A_astzEWJ06_0;
	wire w_dff_A_qGb9CV3y4_0;
	wire w_dff_A_m3yRD9YY2_0;
	wire w_dff_A_C9Ok3oI29_0;
	wire w_dff_A_Ilws0PQQ1_1;
	wire w_dff_B_kt5ToKu03_0;
	wire w_dff_A_9AWUBrYy9_0;
	wire w_dff_A_us1sAlX99_0;
	wire w_dff_A_8KS8086U1_0;
	wire w_dff_A_hgsEczfJ6_1;
	wire w_dff_A_9IFLZ5XQ2_1;
	wire w_dff_A_Z5pizf2f2_1;
	wire w_dff_A_lO8NRHu24_0;
	wire w_dff_A_P4E7cyLt3_0;
	wire w_dff_A_MFLTO2Ch3_0;
	wire w_dff_A_JtIPGaNL4_0;
	wire w_dff_A_f3OZvj1Y3_2;
	wire w_dff_A_kXDMht8p9_2;
	wire w_dff_A_VHghzJcb7_2;
	wire w_dff_A_2aXEwhUq6_2;
	wire w_dff_A_zMiLK88G4_2;
	wire w_dff_A_7atZrdQS0_2;
	wire w_dff_A_J4XvV5vL2_2;
	wire w_dff_A_9DcS5XPD4_2;
	wire w_dff_A_IGkdb4hj6_0;
	wire w_dff_A_LNiO5wDO0_0;
	wire w_dff_A_dBe52Yhh4_1;
	wire w_dff_A_MnIkuD4d6_1;
	wire w_dff_A_tGd31CWb0_1;
	wire w_dff_A_xWlsNxxd9_1;
	wire w_dff_A_xvzK95Pw1_1;
	wire w_dff_A_dYMqDWDe6_1;
	wire w_dff_A_M1oOOEom0_1;
	wire w_dff_A_Sy4bVevd0_2;
	wire w_dff_A_iHds2Ppo4_0;
	wire w_dff_A_JQqvRTx24_0;
	wire w_dff_A_ruYeLqrG0_2;
	wire w_dff_A_mLE1O6VH1_2;
	wire w_dff_A_ZQEm9SnP6_2;
	wire w_dff_A_ejOX0Npw7_2;
	wire w_dff_A_h7pu5H8W1_2;
	wire w_dff_A_pSgOUg0m4_2;
	wire w_dff_A_yr7TgXcb7_2;
	wire w_dff_A_5eVJVE8F5_2;
	wire w_dff_A_kYWp7nK21_2;
	wire w_dff_A_vloAHOvc1_0;
	wire w_dff_A_fE8K8uMx9_0;
	wire w_dff_A_5H7DAu1C4_0;
	wire w_dff_A_4Ryte8mL2_0;
	wire w_dff_A_xDLcMC0L3_0;
	wire w_dff_A_tl2aQEaD1_0;
	wire w_dff_A_mVzC57TR9_0;
	wire w_dff_A_F0l7AFWz3_0;
	wire w_dff_A_PBbAEb990_0;
	wire w_dff_A_SeG4EnS90_0;
	wire w_dff_A_ElGLvhAj1_0;
	wire w_dff_A_5EPsDdxo5_0;
	wire w_dff_A_LxUlK06f0_0;
	wire w_dff_A_lCzPaocn8_2;
	wire w_dff_A_iueAX1qg8_2;
	wire w_dff_A_Zu6j4K7T0_2;
	wire w_dff_A_3Kmfi5V94_2;
	wire w_dff_A_BJcyh7Br9_2;
	wire w_dff_A_UPbk3OGX8_2;
	wire w_dff_A_KdhLW2a17_2;
	wire w_dff_A_YMrjh7iP6_2;
	wire w_dff_A_M2eNuPQZ2_2;
	wire w_dff_A_9HYA86y12_2;
	wire w_dff_A_NMyEOfkP3_0;
	wire w_dff_A_sBDXXBtF8_0;
	wire w_dff_A_92Ak7KAc8_0;
	wire w_dff_A_7g01XhgD9_0;
	wire w_dff_A_zzmjPlyV1_0;
	wire w_dff_A_QrKTtc2A1_0;
	wire w_dff_A_tiFSzDKt6_0;
	wire w_dff_A_2ls2bfCR5_0;
	wire w_dff_A_qzftM5jx2_0;
	wire w_dff_A_kItzOBoR2_0;
	wire w_dff_A_PftzUIhx2_1;
	wire w_dff_A_Ciucv7ih8_1;
	wire w_dff_A_uxKwg3TH2_1;
	wire w_dff_A_7Y8Bwgiw5_1;
	wire w_dff_A_XrQnTngF8_1;
	wire w_dff_A_2z9xH6HH0_1;
	wire w_dff_A_HS47RF610_1;
	wire w_dff_A_xbD5Qbtu0_1;
	wire w_dff_A_N9SE4bwk6_1;
	wire w_dff_A_4sqRfDi83_0;
	wire w_dff_A_L7vwNtPl9_0;
	wire w_dff_A_E8HCYfYS5_0;
	wire w_dff_A_VvPpyrV11_0;
	wire w_dff_A_yOhTKhzB7_0;
	wire w_dff_A_CAtdGYKT0_0;
	wire w_dff_A_Srq3KN5m2_0;
	wire w_dff_A_9rBs5DuH8_0;
	wire w_dff_A_OKjONHKc8_0;
	wire w_dff_A_pzy8VVvM5_0;
	wire w_dff_A_udHnopOJ6_0;
	wire w_dff_A_aDqx3MgK9_0;
	wire w_dff_A_TOm96VmT0_0;
	wire w_dff_A_OYAX7tzg9_2;
	wire w_dff_A_yhkUkvuk4_2;
	wire w_dff_A_M7r6AIJo1_2;
	wire w_dff_A_CWhbu3dK4_2;
	wire w_dff_A_X0Scy0Mx6_2;
	wire w_dff_A_hYjqc3Uq2_2;
	wire w_dff_A_FCCJcO7k9_2;
	wire w_dff_A_T0cGMJoL3_2;
	wire w_dff_A_GQjFCc4r9_2;
	wire w_dff_A_rKuDsEIW0_2;
	wire w_dff_A_oAapYwWF8_2;
	wire w_dff_A_leBPYbM77_2;
	wire w_dff_A_eY5S2s1i4_0;
	wire w_dff_A_kWQ85yIV8_0;
	wire w_dff_A_3ZEeqlf08_0;
	wire w_dff_A_BrvxRotp4_0;
	wire w_dff_A_StcY7TdP4_0;
	wire w_dff_A_vePoAHTu0_0;
	wire w_dff_B_p246Exej3_1;
	wire w_dff_B_khDhyt378_1;
	wire w_dff_B_SoTVFqOj6_1;
	wire w_dff_B_E42CMBiT4_1;
	wire w_dff_B_QIveM39a7_1;
	wire w_dff_B_J0G1r0Mf6_1;
	wire w_dff_B_BY8Aebhw8_1;
	wire w_dff_B_mecUk3Q59_1;
	wire w_dff_B_oBRmApze4_0;
	wire w_dff_B_XmTbCIly1_0;
	wire w_dff_B_KKMEIeZg9_0;
	wire w_dff_B_QAuHnfYV8_0;
	wire w_dff_A_cBzamRCz6_0;
	wire w_dff_A_KDzKgusz2_0;
	wire w_dff_A_p7REkyA23_0;
	wire w_dff_A_J5JKGTJv5_0;
	wire w_dff_A_CCZIbur15_0;
	wire w_dff_A_bp3UPr9D4_0;
	wire w_dff_A_bgtWyCku0_0;
	wire w_dff_A_Zs0Q64kA6_0;
	wire w_dff_A_pgQqVXZC5_0;
	wire w_dff_A_HziYoL3O0_0;
	wire w_dff_A_hLHVdNtW3_0;
	wire w_dff_A_KB4MxrlC1_2;
	wire w_dff_A_hwYlgUYn7_2;
	wire w_dff_A_6WZiKHKH9_2;
	wire w_dff_A_iXmpsiu60_2;
	wire w_dff_A_YnVsCIew1_2;
	wire w_dff_A_F3nGzQEX1_2;
	wire w_dff_A_8GIHkBZ16_2;
	wire w_dff_A_spQo6kNC4_2;
	wire w_dff_A_8dvVbGxP0_2;
	wire w_dff_A_SebHfa9a5_2;
	wire w_dff_A_tz7qKgnZ4_1;
	wire w_dff_A_5gHDYrhf4_1;
	wire w_dff_A_nulbQinz5_1;
	wire w_dff_A_ReHVIFOI4_2;
	wire w_dff_A_ZmqweskX2_2;
	wire w_dff_A_BQoRkNuz7_1;
	wire w_dff_A_gna1lane3_1;
	wire w_dff_A_6HSQCE8g2_1;
	wire w_dff_A_ACrTOCto7_1;
	wire w_dff_A_SaBZhgma6_1;
	wire w_dff_A_FvSoSi5H3_2;
	wire w_dff_A_ayT2PZaO5_2;
	wire w_dff_A_4EdfMcyJ7_2;
	wire w_dff_A_QDiCPetD4_2;
	wire w_dff_A_a77PsJUx4_2;
	wire w_dff_A_rUnl0ppz2_0;
	wire w_dff_A_skkI8VF88_2;
	wire w_dff_A_YSi94fau9_2;
	wire w_dff_A_AuzAKPCc6_1;
	wire w_dff_A_hM3THRsg9_1;
	wire w_dff_A_JmW3Ihxc8_1;
	wire w_dff_A_WVSrChD69_1;
	wire w_dff_A_bnC8QV0j7_2;
	wire w_dff_B_YnaDh83O0_1;
	wire w_dff_B_cuojKOfz4_1;
	wire w_dff_A_Su0dW8rr4_1;
	wire w_dff_A_0yhDhK1R7_2;
	wire w_dff_A_R3WQr2sD2_2;
	wire w_dff_A_ijVSSTmt9_0;
	wire w_dff_A_tpmf8KZl1_0;
	wire w_dff_A_3YjxHHOi9_0;
	wire w_dff_A_JWCzRV0Q8_0;
	wire w_dff_A_naQTATWe7_0;
	wire w_dff_A_ZoHb93cZ1_0;
	wire w_dff_A_vQANGHd58_0;
	wire w_dff_A_bMsbkEkt6_2;
	wire w_dff_A_GQPiGC388_2;
	wire w_dff_A_NOvU5JuC3_2;
	wire w_dff_A_x3XqxMef9_2;
	wire w_dff_A_lTn0LJ062_2;
	wire w_dff_A_TZ7yFRSH9_2;
	wire w_dff_A_ew18bozs6_2;
	wire w_dff_A_cepuc8ky3_2;
	wire w_dff_A_DZ2umtH22_2;
	wire w_dff_A_8FFohwbb2_2;
	wire w_dff_A_5EsIkV012_2;
	wire w_dff_A_PRPk6bvs1_2;
	wire w_dff_A_jb9Wwk7I8_2;
	wire w_dff_A_m8AjJmOU7_2;
	wire w_dff_A_gXQuaMnl3_2;
	wire w_dff_A_ZypU1M0j6_1;
	wire w_dff_A_KNfRQKVM6_1;
	wire w_dff_B_Ji80iO3W0_1;
	wire w_dff_B_OEsLG4yF6_1;
	wire w_dff_A_A6Ofxp4u6_1;
	wire w_dff_A_ZN1HbWSE0_1;
	wire w_dff_A_WxnTA56b3_2;
	wire w_dff_A_udFISggS8_0;
	wire w_dff_A_Z6NkXakE9_0;
	wire w_dff_A_hhute4kg0_0;
	wire w_dff_A_Kqjde74b7_0;
	wire w_dff_A_UtHLjOxk6_0;
	wire w_dff_A_b53XyEOm5_0;
	wire w_dff_A_PB8t3Hvz9_1;
	wire w_dff_A_H0zqYxPy1_1;
	wire w_dff_A_Er0bsRYb9_1;
	wire w_dff_A_udnaR6Ee8_1;
	wire w_dff_A_eU84hw6U8_1;
	wire w_dff_A_OGcwN2MC2_1;
	wire w_dff_A_N0BEEMJX4_0;
	wire w_dff_A_DjXYqC9V1_0;
	wire w_dff_A_xkG9Hc0j8_0;
	wire w_dff_A_yP34O01m9_0;
	wire w_dff_A_ecswXMSM3_0;
	wire w_dff_A_TMEXgCiV3_0;
	wire w_dff_A_LCUuEBXe0_0;
	wire w_dff_A_RKSuQUOB6_0;
	wire w_dff_A_1UgETKAM2_1;
	wire w_dff_A_1LD0OQSW4_1;
	wire w_dff_A_5IjsnvRM4_1;
	wire w_dff_A_faN238Rh5_1;
	wire w_dff_A_9WTQOPrW0_1;
	wire w_dff_A_81qg6Jm97_1;
	wire w_dff_A_r0X3Rd9Y4_1;
	wire w_dff_A_2EJuJVo33_1;
	wire w_dff_A_ElvWcEP37_0;
	wire w_dff_A_v2CFLhBw2_0;
	wire w_dff_A_zq8Txwaj5_0;
	wire w_dff_A_ubxbXNuN4_0;
	wire w_dff_A_28Uh1vw04_0;
	wire w_dff_A_PLkSvc9g4_0;
	wire w_dff_A_belxD7F03_0;
	wire w_dff_A_oNI79irw8_0;
	wire w_dff_A_g9nn8Zc14_1;
	wire w_dff_B_Tqm4dI2w6_0;
	wire w_dff_A_8z1FTl5P0_0;
	wire w_dff_A_aKkaL1z45_0;
	wire w_dff_A_oU1nba1o6_0;
	wire w_dff_A_TgPEKW4v9_1;
	wire w_dff_B_RrvFTnon4_1;
	wire w_dff_B_PzI6ITzR8_1;
	wire w_dff_B_Qf4tPweB9_1;
	wire w_dff_A_9umbvbKS6_0;
	wire w_dff_A_Qvpf57IH7_0;
	wire w_dff_A_XszD7M3c5_1;
	wire w_dff_A_AC2I0mRQ3_1;
	wire w_dff_A_kuQLI3Vo2_1;
	wire w_dff_A_HVUG87jc0_2;
	wire w_dff_A_7LBgXwEW5_2;
	wire w_dff_A_mLm1PJlt2_0;
	wire w_dff_A_HeBLclxv7_0;
	wire w_dff_A_y9csACmr9_0;
	wire w_dff_A_qmCoNXiI4_1;
	wire w_dff_A_nKLqndak4_1;
	wire w_dff_A_tGoKlo0V2_1;
	wire w_dff_A_uwjvYkAu9_0;
	wire w_dff_A_wreUxZbJ9_0;
	wire w_dff_A_cftYHiFH1_0;
	wire w_dff_A_dZ7D7Tmw4_2;
	wire w_dff_A_pfWE9oTo5_2;
	wire w_dff_A_Fw7xNyJB7_2;
	wire w_dff_A_Az6zVtTd4_2;
	wire w_dff_A_vjQCyBhw6_2;
	wire w_dff_A_gnrdzkWR0_0;
	wire w_dff_A_WCp84g3m6_0;
	wire w_dff_A_UybTJBfR0_0;
	wire w_dff_A_vj4kD5vR4_1;
	wire w_dff_A_wW8gMsRw4_1;
	wire w_dff_A_pMvMwwFC3_1;
	wire w_dff_A_vga5hyTG0_1;
	wire w_dff_A_GKGGy3Mq8_2;
	wire w_dff_A_nvMEuQpG9_2;
	wire w_dff_A_dOZL61cq6_1;
	wire w_dff_A_7tTiqfhT6_1;
	wire w_dff_A_8o0l8bfO3_2;
	wire w_dff_A_3AAwax0a6_2;
	wire w_dff_A_M86Y64q06_1;
	wire w_dff_A_IxbcIBxm6_1;
	wire w_dff_A_Jo7k03HD9_2;
	wire w_dff_A_hSgxQEJA9_2;
	wire w_dff_A_b1EAzkv06_2;
	wire w_dff_B_WnJKDA8q3_3;
	wire w_dff_A_QPcPdCI90_1;
	wire w_dff_A_Rb3AcJSg6_0;
	wire w_dff_A_YNlKx5VQ6_0;
	wire w_dff_A_GCs8Nm6Y4_2;
	wire w_dff_A_yqzXBbLR1_2;
	wire w_dff_A_ZYdtO75G0_2;
	wire w_dff_A_QCW8hcPI2_1;
	wire w_dff_A_iD4J6MS45_1;
	wire w_dff_A_JXJGeXc22_0;
	wire w_dff_A_1Pahpig79_0;
	wire w_dff_A_4Yknphgw5_0;
	wire w_dff_A_jvI5Dpa70_0;
	wire w_dff_A_8MA6hMpj0_0;
	wire w_dff_A_cWKHglpW6_0;
	wire w_dff_A_RFIN0BPS2_0;
	wire w_dff_A_B9Pl3UY61_0;
	wire w_dff_A_mXN2Xjw79_0;
	wire w_dff_A_amIHWbpj5_0;
	wire w_dff_A_2NR8m91N7_0;
	wire w_dff_A_3sbJ8hsb1_0;
	wire w_dff_A_v6RcmkOt3_0;
	wire w_dff_A_oHxxIHUn5_0;
	wire w_dff_A_FjzdyPWx7_0;
	wire w_dff_A_rpg1F2RK8_0;
	wire w_dff_A_ZszvsuPY6_0;
	wire w_dff_A_lhYU8i2i5_0;
	wire w_dff_A_EwrqlWyp2_1;
	wire w_dff_A_2sAm4jEc0_1;
	wire w_dff_A_wabDsVEP0_1;
	wire w_dff_A_m6esQfdP1_1;
	wire w_dff_A_R06S8aZw0_1;
	wire w_dff_A_lIULxlXG7_1;
	wire w_dff_A_W1E9wiDD9_1;
	wire w_dff_A_HzEUQJyU0_1;
	wire w_dff_A_gNdOfnno1_1;
	wire w_dff_A_q2xWHlDq8_0;
	wire w_dff_A_rTxpwddn3_1;
	wire w_dff_A_wuTDcEKF8_1;
	wire w_dff_A_2XCjO6Ip1_1;
	wire w_dff_A_LNEZeKsk8_1;
	wire w_dff_A_GYbrrVB18_1;
	wire w_dff_A_XsW0EsCf7_1;
	wire w_dff_A_Dy3TAhzW2_1;
	wire w_dff_A_OUi7JFIo4_1;
	wire w_dff_A_Kmx4IvMP5_1;
	wire w_dff_B_WZdnyJp83_0;
	wire w_dff_B_hEwfdFJC4_0;
	wire w_dff_A_X07PXF714_0;
	wire w_dff_A_5Bk3phfE6_0;
	wire w_dff_A_ILUERALf3_1;
	wire w_dff_A_Xp4JgKbh6_1;
	wire w_dff_A_Ik8vCPxA0_1;
	wire w_dff_A_Hx5Huinu0_2;
	wire w_dff_A_55jDWv245_2;
	wire w_dff_B_O5lDCoGi9_1;
	wire w_dff_B_6s69clhL3_1;
	wire w_dff_B_ThrNonlU3_1;
	wire w_dff_A_E5wgSxP68_0;
	wire w_dff_A_zZy4bo4X3_1;
	wire w_dff_A_SZoFlOny9_1;
	wire w_dff_A_jZz3IHDG8_1;
	wire w_dff_A_CfHpfQCw4_2;
	wire w_dff_A_77fyP2ar1_2;
	wire w_dff_A_2dNZana21_2;
	wire w_dff_A_WhbXSYJK8_1;
	wire w_dff_A_Hz8IvoM91_1;
	wire w_dff_A_4EL6Kdd02_1;
	wire w_dff_A_jAqQNxKk1_2;
	wire w_dff_A_t6R5PWtB3_2;
	wire w_dff_A_twm6ZtqJ4_2;
	wire w_dff_A_dZWH8cyL6_2;
	wire w_dff_A_oBcMi1la7_2;
	wire w_dff_A_zvQa7yxe5_2;
	wire w_dff_A_xZyeqGsy9_2;
	wire w_dff_A_2EJxM0j54_0;
	wire w_dff_A_3QeCQqy86_0;
	wire w_dff_A_dfW7T59s0_2;
	wire w_dff_A_pDj358Ch0_0;
	wire w_dff_A_C1G414EV2_0;
	wire w_dff_A_M3o1gwDr0_0;
	wire w_dff_A_gPqY2UvA5_1;
	wire w_dff_A_UEp8HpzD5_1;
	wire w_dff_A_YSKr3QoK9_1;
	wire w_dff_A_jMOKjR4O9_0;
	wire w_dff_A_s1QWKw7V6_0;
	wire w_dff_A_4FvfAcLi4_0;
	wire w_dff_A_MHD1ok412_1;
	wire w_dff_A_XyTCi7xB9_1;
	wire w_dff_A_u11qo1Wn5_1;
	wire w_dff_A_Q5xQh3CZ8_0;
	wire w_dff_A_wFaGRlsO1_1;
	wire w_dff_A_myOFtcpJ7_2;
	wire w_dff_A_kKS7HTiK1_2;
	wire w_dff_A_FvBhCFCY3_0;
	wire w_dff_A_dOsjTESK6_0;
	wire w_dff_A_hiFDXRRs9_0;
	wire w_dff_B_uJ3xOORm6_0;
	wire w_dff_B_l2pSoTrH7_0;
	wire w_dff_A_G2a5RTLJ1_0;
	wire w_dff_A_Qu1KcUFZ3_0;
	wire w_dff_A_y5QVgwBk6_1;
	wire w_dff_A_2A6upE0W0_2;
	wire w_dff_A_PWJAmKAm3_0;
	wire w_dff_A_eWawSKNL7_0;
	wire w_dff_A_x0xr0h3r0_0;
	wire w_dff_A_Nx08apME8_0;
	wire w_dff_A_cQeHUXR74_2;
	wire w_dff_A_nt1bhD358_0;
	wire w_dff_A_X78oElrO3_0;
	wire w_dff_A_XMenjuw07_1;
	wire w_dff_A_9bPYAUYV5_0;
	wire w_dff_A_TlLqHoIT8_0;
	wire w_dff_A_kOZD6D7K7_0;
	wire w_dff_A_sitw6DNQ1_0;
	wire w_dff_A_BcLcGbZ95_0;
	wire w_dff_A_cPT0Uvut7_0;
	wire w_dff_A_xm7aeCbx9_1;
	wire w_dff_A_CgkkcF1d8_2;
	wire w_dff_A_dSGRiRnu7_2;
	wire w_dff_A_BHeSO7qT3_2;
	wire w_dff_A_2miAVqjQ8_1;
	wire w_dff_A_uuSGeSRB5_1;
	wire w_dff_A_K6dqxKfC2_1;
	wire w_dff_A_CqsrBYPW0_2;
	wire w_dff_A_0q8OseDv1_2;
	wire w_dff_A_YMOYBBOY5_2;
	wire w_dff_A_2czuDZR02_0;
	wire w_dff_A_TSdrlmcq5_2;
	wire w_dff_B_JYUQ1Fpi1_3;
	wire w_dff_B_pUTUUMiT7_3;
	wire w_dff_B_pnGVR7CE7_3;
	wire w_dff_B_sD7AOtzq4_3;
	wire w_dff_B_TEVwNqdr1_3;
	wire w_dff_B_KMQGD8eI4_3;
	wire w_dff_B_q7cY9u6B8_3;
	wire w_dff_B_fPAlwEwd1_3;
	wire w_dff_B_40nn1Lwz9_3;
	wire w_dff_B_sBT8MF3N1_3;
	wire w_dff_B_XgAtqVZK0_3;
	wire w_dff_B_xtK22yGs4_3;
	wire w_dff_B_C95NgCdz3_3;
	wire w_dff_A_hgtqga5P4_0;
	wire w_dff_A_uUwQnBy62_0;
	wire w_dff_A_RisR2R3J7_0;
	wire w_dff_A_tjPHyHJn9_0;
	wire w_dff_A_lgHh6aBg8_0;
	wire w_dff_A_Ekp2IG5W4_0;
	wire w_dff_A_p0cEIKKC8_0;
	wire w_dff_A_hfEkKlwp6_0;
	wire w_dff_A_Ry1rX72q4_0;
	wire w_dff_A_F3IObSgd7_0;
	wire w_dff_A_IMLKiumh3_0;
	wire w_dff_A_Sl5uowRH7_0;
	wire w_dff_A_6ly3l6PO0_2;
	wire w_dff_A_jHpiulKy1_2;
	wire w_dff_A_0H6vXaff9_2;
	wire w_dff_A_LyjjHCk80_2;
	wire w_dff_A_JpVKkyZd2_2;
	wire w_dff_A_ZXPClYE07_2;
	wire w_dff_A_CmrXkvrz6_2;
	wire w_dff_A_QbbBYFjq7_2;
	wire w_dff_A_jBEXj34q3_2;
	wire w_dff_A_lLMrfQwz0_2;
	wire w_dff_A_I9tN8kjN3_2;
	wire w_dff_A_CMbgeeVU9_1;
	wire w_dff_A_FdAIvIHk9_1;
	wire w_dff_A_xbIFYLSo9_1;
	wire w_dff_A_8wFEYYyP1_1;
	wire w_dff_A_Q1KQFFFf3_1;
	wire w_dff_A_PxRhIh5L4_1;
	wire w_dff_A_hdzvul4H2_1;
	wire w_dff_A_LlBPJ9I44_2;
	wire w_dff_A_Zjy67xRR6_2;
	wire w_dff_A_NOPBrzRH5_2;
	wire w_dff_A_mf1f6WvQ6_2;
	wire w_dff_A_DLFXdhd73_2;
	wire w_dff_A_1R9Si16O6_0;
	wire w_dff_A_obybAHqW1_0;
	wire w_dff_A_Qc3xcAoD7_0;
	wire w_dff_A_FXKyyztp3_0;
	wire w_dff_A_3uKSBR5i7_0;
	wire w_dff_A_sWTMSEHn0_0;
	wire w_dff_A_12WjBE4m9_0;
	wire w_dff_A_qYB9Dq1x9_0;
	wire w_dff_A_GWni51SR5_0;
	wire w_dff_A_UlhBziJO7_0;
	wire w_dff_A_rTeRCFc31_0;
	wire w_dff_A_IvWnj4Wv1_0;
	wire w_dff_A_AqgmJPPZ1_0;
	wire w_dff_A_wfZHBpMz4_0;
	wire w_dff_A_0xhGggqU0_1;
	wire w_dff_A_QefcfXOk7_1;
	wire w_dff_A_4NiS6VyX1_1;
	wire w_dff_A_FRc0Ilhy3_1;
	wire w_dff_A_3wM92rCX6_1;
	wire w_dff_A_IGQnP4ks6_1;
	wire w_dff_A_nVb6Ejce5_1;
	wire w_dff_A_tppcESnG0_1;
	wire w_dff_A_kEuUguBW8_1;
	wire w_dff_A_BIZ6vh7c2_1;
	wire w_dff_A_4HbW5Xy46_1;
	wire w_dff_A_A2BL1Dqj5_1;
	wire w_dff_A_8rU6N7RT9_1;
	wire w_dff_A_MagKJvnV4_1;
	wire w_dff_A_3dAvlS0C4_1;
	wire w_dff_A_LDI5uEvl8_1;
	wire w_dff_A_wgx6Rqqe4_1;
	wire w_dff_A_yL92aNsz9_1;
	wire w_dff_A_GTI0iPQO3_1;
	wire w_dff_A_FjQWOwTT2_1;
	wire w_dff_A_uRAYGopk5_1;
	wire w_dff_A_WZu9qbWm8_1;
	wire w_dff_A_8dtSbyEy9_1;
	wire w_dff_A_WSlqBq2Q4_1;
	wire w_dff_A_ZThLgVBk1_1;
	wire w_dff_A_gLfYp3ZM8_1;
	wire w_dff_A_pdliC2tE7_1;
	wire w_dff_A_oKM9GWo78_1;
	wire w_dff_A_PZ0LGSYx0_1;
	wire w_dff_A_Oglos4Ku8_2;
	wire w_dff_A_Ya9hip4R8_2;
	wire w_dff_A_d0Thoz854_2;
	wire w_dff_A_QrPAXaBb6_2;
	wire w_dff_A_EmCbQ7yN5_2;
	wire w_dff_A_i3JSTl7Z2_2;
	wire w_dff_A_H7XOka0E0_2;
	wire w_dff_A_ECridoI04_2;
	wire w_dff_A_lrCOda6n4_2;
	wire w_dff_A_CHTE9K1c1_2;
	wire w_dff_A_GgC3TkUe9_2;
	wire w_dff_A_u9yvO9bL3_2;
	wire w_dff_A_nsfrGHtl6_2;
	wire w_dff_A_JxrKfOgy3_2;
	wire w_dff_A_KFHMGHX69_2;
	wire w_dff_A_PI2cxiYp5_2;
	wire w_dff_A_4pvAQzxU1_2;
	wire w_dff_B_1Lv68ur21_3;
	wire w_dff_A_JwdWPdBz1_1;
	wire w_dff_A_ix5lpmXU0_1;
	wire w_dff_A_WlqT3q5V3_1;
	wire w_dff_A_QqWgiOB68_0;
	wire w_dff_A_d48y1CTs7_2;
	wire w_dff_A_shuBNnAO4_2;
	wire w_dff_A_DjzwFZwv6_0;
	wire w_dff_A_BqhNtu9n3_2;
	wire w_dff_A_5LV0ZNYi7_0;
	wire w_dff_A_yWAHEjrD4_0;
	wire w_dff_A_C0Y1nxKr5_0;
	wire w_dff_A_N8uUEA564_0;
	wire w_dff_A_FC1iz72s0_0;
	wire w_dff_A_mYU0z91q4_0;
	wire w_dff_A_xgDM7dwZ7_0;
	wire w_dff_A_PWK2Wi2W5_0;
	wire w_dff_A_OcU4o0PY9_0;
	wire w_dff_A_6iuFEKGn1_0;
	wire w_dff_A_fa7POqnd3_0;
	wire w_dff_A_eA3Hz6G88_0;
	wire w_dff_A_QNi4j1dS1_0;
	wire w_dff_A_RJcwQIOp0_0;
	wire w_dff_A_7FQombol2_0;
	wire w_dff_A_R9Tb3AaW0_0;
	wire w_dff_A_WIoQs0wk6_0;
	wire w_dff_A_PjYVHhuR2_0;
	wire w_dff_A_fWHv26iz4_0;
	wire w_dff_A_99Pg9m6g2_0;
	wire w_dff_A_AHJMJUka6_0;
	wire w_dff_A_zvrsVdck8_0;
	wire w_dff_A_NZyLzJFy7_0;
	wire w_dff_A_tviPC0cg8_0;
	wire w_dff_A_gVbHCnsA3_0;
	wire w_dff_A_egO8b8PU9_0;
	wire w_dff_A_bhftzGJH2_0;
	wire w_dff_A_rTq4C2s82_0;
	wire w_dff_A_QgXvcrKk2_0;
	wire w_dff_A_wO4aJOgl9_0;
	wire w_dff_A_DSBhHVGb0_2;
	wire w_dff_A_sOs4v8DJ5_2;
	wire w_dff_A_BUFbwBqi6_2;
	wire w_dff_A_kEcJPfP69_2;
	wire w_dff_A_vMKfo7I57_2;
	wire w_dff_A_SsWESpZx2_2;
	wire w_dff_A_E0A4jplz8_2;
	wire w_dff_A_1ll4yG0V1_2;
	wire w_dff_A_B3QQj4Ub4_2;
	wire w_dff_A_qXc8K7HE9_2;
	wire w_dff_A_kae52u6T9_2;
	wire w_dff_A_74MvuWDk0_2;
	wire w_dff_A_ZTuxilk38_2;
	wire w_dff_A_qBD6oLY86_2;
	wire w_dff_A_kOpgo1hg4_2;
	wire w_dff_A_WIx6MBO00_2;
	wire w_dff_A_qgnPfh6H0_0;
	wire w_dff_A_rJrIH5jY5_1;
	wire w_dff_A_C3AB7ibC0_2;
	wire w_dff_A_Q46LP6PO3_2;
	wire w_dff_A_G1WJMjkL0_2;
	wire w_dff_A_7986Ijkt6_2;
	wire w_dff_A_5x6ZmtxS3_0;
	wire w_dff_A_7JrKyfu22_0;
	wire w_dff_A_Y8WSD0v91_2;
	wire w_dff_A_smLdoHTq5_2;
	wire w_dff_A_8uDIUc495_0;
	wire w_dff_A_IRLX5wUz8_2;
	wire w_dff_A_CHib6UZM2_1;
	wire w_dff_A_lI6RmWBc9_1;
	wire w_dff_A_I7yF9JIC0_1;
	wire w_dff_A_IEut3ixz5_1;
	wire w_dff_A_0sJdbqaP8_1;
	wire w_dff_A_jeojB7IL6_1;
	wire w_dff_A_sIpatig60_1;
	wire w_dff_A_gMBPaD9G2_1;
	wire w_dff_A_O2bBxmb51_1;
	wire w_dff_A_uoPZYNJ70_1;
	wire w_dff_A_PB3oHri44_1;
	wire w_dff_A_NdEaSX8R9_2;
	wire w_dff_A_7HilQhhT0_2;
	wire w_dff_A_dvfHxH6U7_2;
	wire w_dff_A_lQD0TU6M9_0;
	wire w_dff_A_FXipZlDr0_0;
	wire w_dff_A_ViIZUB9l5_0;
	wire w_dff_A_2akBU97p0_0;
	wire w_dff_A_yvX93bRn9_0;
	wire w_dff_A_mvXyFqv12_0;
	wire w_dff_A_2pL9S8xB2_0;
	wire w_dff_A_vrS3NHSZ1_0;
	wire w_dff_A_sVWFZwx82_0;
	wire w_dff_A_SCcE3mM90_0;
	wire w_dff_A_ZxMMe4fR3_0;
	wire w_dff_A_0WhpOIuC2_0;
	wire w_dff_A_m1CnoXj26_0;
	wire w_dff_A_g5H1H4El9_0;
	wire w_dff_A_yfPBnnf84_0;
	wire w_dff_A_ufkPlikO5_0;
	wire w_dff_A_RLJVZK2G8_0;
	wire w_dff_A_BaOeCvDH3_0;
	wire w_dff_A_OKumeTud6_0;
	wire w_dff_A_YlHksyqL1_0;
	wire w_dff_A_JwsvjUze0_0;
	wire w_dff_A_8VYXWAyJ9_0;
	wire w_dff_A_n9C3awQk2_0;
	wire w_dff_A_YkZB4vyM3_0;
	wire w_dff_A_I7A3yWWS5_0;
	wire w_dff_A_wCCyFw6L0_0;
	wire w_dff_A_jteEvgx45_1;
	wire w_dff_A_X67LN1Bf4_0;
	wire w_dff_A_jMdOBbu30_0;
	wire w_dff_A_XJfZkCo89_0;
	wire w_dff_A_WlyUcA2o3_0;
	wire w_dff_A_ZLuIMkLz5_0;
	wire w_dff_A_IQZCiqyM2_0;
	wire w_dff_A_7Bxq12E40_0;
	wire w_dff_A_Oh6VSvYU0_0;
	wire w_dff_A_pgFRIrOs0_0;
	wire w_dff_A_70xqkUAe6_0;
	wire w_dff_A_3p3GpOYP7_0;
	wire w_dff_A_54q4HlXO8_0;
	wire w_dff_A_wkE7jZiQ1_0;
	wire w_dff_A_UioTpEI78_0;
	wire w_dff_A_g8xwiyng7_0;
	wire w_dff_A_BKhw5jh21_0;
	wire w_dff_A_VetyY1zY4_0;
	wire w_dff_A_eHSwebds9_0;
	wire w_dff_A_2w49CTng6_0;
	wire w_dff_A_7X90HefZ6_0;
	wire w_dff_A_0GD5q4Eq8_0;
	wire w_dff_A_nNCInwRr4_0;
	wire w_dff_A_f78lEgGc0_0;
	wire w_dff_A_MAFvvJ157_0;
	wire w_dff_A_yqhI50uz1_0;
	wire w_dff_A_Hf1wkeAO0_0;
	wire w_dff_A_qOUGhVbK5_0;
	wire w_dff_A_JOEDEGQA0_2;
	wire w_dff_A_rYz2HKC41_0;
	wire w_dff_A_1YTb7ARq9_0;
	wire w_dff_A_5O2kPZzG2_0;
	wire w_dff_A_APvWXbhT4_0;
	wire w_dff_A_qO3YfwMZ8_0;
	wire w_dff_A_4lztVejE9_0;
	wire w_dff_A_l0UyLx583_0;
	wire w_dff_A_v8k0iaiU6_0;
	wire w_dff_A_DihRufN79_0;
	wire w_dff_A_lIXyRskE8_0;
	wire w_dff_A_bPbxL5fV0_0;
	wire w_dff_A_mmRqkyfv9_0;
	wire w_dff_A_cZ5LdLCG5_0;
	wire w_dff_A_Vxg88BlP0_0;
	wire w_dff_A_LefBbsUQ1_0;
	wire w_dff_A_hDdd8gJf2_0;
	wire w_dff_A_hB0ERWBs1_0;
	wire w_dff_A_KG9hLs979_0;
	wire w_dff_A_eLKBOjPD9_0;
	wire w_dff_A_zC8URcQ80_0;
	wire w_dff_A_NqXqbQbd6_0;
	wire w_dff_A_G8WT6kR23_0;
	wire w_dff_A_IRozgalU2_2;
	wire w_dff_A_6EuHXGSU2_0;
	wire w_dff_A_jUpMeuZt8_0;
	wire w_dff_A_OhViaEMp3_0;
	wire w_dff_A_jtHrDZij6_0;
	wire w_dff_A_NEi4l9kO4_0;
	wire w_dff_A_KmcwJAqm2_0;
	wire w_dff_A_xkNIAmfP4_0;
	wire w_dff_A_AGjpLRWf3_0;
	wire w_dff_A_yNoHbPBA8_0;
	wire w_dff_A_NhLXKGeP9_0;
	wire w_dff_A_SgFdvEgU6_0;
	wire w_dff_A_lLYoPJk01_0;
	wire w_dff_A_t3l7K1vH2_0;
	wire w_dff_A_ygHS9l900_0;
	wire w_dff_A_PCmF4Sys9_0;
	wire w_dff_A_uRItRhdz3_0;
	wire w_dff_A_16p9pGa21_0;
	wire w_dff_A_BtAV4KZf3_0;
	wire w_dff_A_bajZLfm07_0;
	wire w_dff_A_fRu6qHu15_0;
	wire w_dff_A_OQp68ksv5_0;
	wire w_dff_A_z1k4NQFU1_0;
	wire w_dff_A_Kpjv5gdY0_0;
	wire w_dff_A_nQIK8Zit8_0;
	wire w_dff_A_T0ChLpHK4_0;
	wire w_dff_A_rJIYourm4_2;
	wire w_dff_A_TOumBzkK2_0;
	wire w_dff_A_bjhIJXWY0_0;
	wire w_dff_A_XpghVJi75_0;
	wire w_dff_A_u3iZTuj79_0;
	wire w_dff_A_Lvb23Mf41_0;
	wire w_dff_A_SRgK80nf5_0;
	wire w_dff_A_SSh2RfLE9_0;
	wire w_dff_A_6omLeoJL4_0;
	wire w_dff_A_UqBhDRfT9_0;
	wire w_dff_A_ENrCIkFF9_0;
	wire w_dff_A_ptCoTQtI9_0;
	wire w_dff_A_A0GQ3z722_0;
	wire w_dff_A_pDPzjMxa5_0;
	wire w_dff_A_sUXIRc6K2_0;
	wire w_dff_A_xUBjtKW42_0;
	wire w_dff_A_VVge2dm36_0;
	wire w_dff_A_awm6kvCg6_0;
	wire w_dff_A_CaLOVrzE3_0;
	wire w_dff_A_lrij1AOu6_0;
	wire w_dff_A_AUbvzYts2_0;
	wire w_dff_A_T1ZfaDTv1_0;
	wire w_dff_A_iBxk3XZc2_0;
	wire w_dff_A_C1kxaIbC2_0;
	wire w_dff_A_iSpF9Bqd8_0;
	wire w_dff_A_9CN4yY6f6_0;
	wire w_dff_A_l5NPhoxX4_0;
	wire w_dff_A_8Q6yYxeC8_2;
	wire w_dff_A_WryAIHdl9_0;
	wire w_dff_A_Ns2Rn6eP8_0;
	wire w_dff_A_PMnLeR4T5_0;
	wire w_dff_A_UcateCLQ6_0;
	wire w_dff_A_8mJTbhwH7_0;
	wire w_dff_A_pFxc3PwR3_0;
	wire w_dff_A_fO3yNdQP8_0;
	wire w_dff_A_6i5VrFKt7_0;
	wire w_dff_A_eu8WA5MA7_0;
	wire w_dff_A_03dKo0OU5_0;
	wire w_dff_A_ogyD4tfk5_0;
	wire w_dff_A_uO2oNi8c1_0;
	wire w_dff_A_QxrJEAvT4_0;
	wire w_dff_A_cLFUR3629_2;
	wire w_dff_A_TE1fgRoX5_0;
	wire w_dff_A_QduNW8g18_0;
	wire w_dff_A_BAQ5CWZM6_0;
	wire w_dff_A_mB2QYAqB5_0;
	wire w_dff_A_Rz2uBJNn8_0;
	wire w_dff_A_ziIlOHJp2_0;
	wire w_dff_A_ryW1PJWv3_0;
	wire w_dff_A_RxKSzTvT1_0;
	wire w_dff_A_ZLCaXi6H5_0;
	wire w_dff_A_P68wLghG5_0;
	wire w_dff_A_tmYKP9X75_0;
	wire w_dff_A_dB0sU7VX1_2;
	wire w_dff_A_MxtLPZu36_0;
	wire w_dff_A_HotI6sFd3_0;
	wire w_dff_A_ubLH2ZY53_0;
	wire w_dff_A_mp4Cxt8K0_0;
	wire w_dff_A_3cpAejMl5_0;
	wire w_dff_A_KsaeLJyy1_0;
	wire w_dff_A_W8BEe51M6_0;
	wire w_dff_A_SjPffqPZ2_0;
	wire w_dff_A_cd2AsH7w8_0;
	wire w_dff_A_TSaMQ2GW2_0;
	wire w_dff_A_QIJzC3fc7_0;
	wire w_dff_A_Aew9ff5B4_0;
	wire w_dff_A_yhA4RyZz4_0;
	wire w_dff_A_pYXSlu0u3_2;
	wire w_dff_A_cyy8OSOT3_0;
	wire w_dff_A_1c7FcxnV5_0;
	wire w_dff_A_5kO10u8s0_0;
	wire w_dff_A_3BBkXED38_0;
	wire w_dff_A_KwwakGil9_0;
	wire w_dff_A_VcxXrr4O6_0;
	wire w_dff_A_NdrhWOkV6_0;
	wire w_dff_A_MsZJIKpq4_0;
	wire w_dff_A_7VLwJoOx0_1;
	wire w_dff_A_PssIiQXc0_0;
	wire w_dff_A_ePdVpKv11_0;
	wire w_dff_A_ctvXemYK2_0;
	wire w_dff_A_l6ymKFxy6_0;
	wire w_dff_A_JF0rtjhO4_0;
	wire w_dff_A_dYO5zxbJ5_0;
	wire w_dff_A_mEcX5aBD7_0;
	wire w_dff_A_gsv9fq2T7_0;
	wire w_dff_A_pVLj9Wzt1_0;
	wire w_dff_A_lIpENpu48_0;
	wire w_dff_A_aE38d95m6_0;
	wire w_dff_A_ARHG76Xk0_0;
	wire w_dff_A_cMTHFec67_1;
	wire w_dff_A_rfD6WCBD7_0;
	wire w_dff_A_aG5zNwq98_0;
	wire w_dff_A_5vo19zre5_0;
	wire w_dff_A_yiMVGmsJ9_0;
	wire w_dff_A_SuASy8FB1_0;
	wire w_dff_A_KaTjYwsO0_0;
	wire w_dff_A_igJmY0qZ1_0;
	wire w_dff_A_tne6B1924_2;
	wire w_dff_A_bsRgQ6HQ9_0;
	wire w_dff_A_BbNo7saQ6_0;
	wire w_dff_A_7rhlFlZj9_0;
	wire w_dff_A_eBfPA8zD8_0;
	wire w_dff_A_QlyGS8GL6_0;
	wire w_dff_A_uqG9iPFp0_0;
	wire w_dff_A_vfRDkQlW9_1;
	wire w_dff_A_nNRWStQ55_0;
	wire w_dff_A_XPIeNpRI4_0;
	wire w_dff_A_zoC0sDli6_0;
	wire w_dff_A_KukjoOi82_0;
	wire w_dff_A_SL9TcYRZ1_0;
	wire w_dff_A_ywVOaL5R9_1;
	wire w_dff_A_EPAaCQJU2_0;
	wire w_dff_A_iAa84ZRP0_0;
	wire w_dff_A_S8cpcl4d3_0;
	wire w_dff_A_eKIaLvsK6_0;
	wire w_dff_A_r4TZM15t1_0;
	wire w_dff_A_NaAXIQL28_0;
	wire w_dff_A_Ezxpsepx8_1;
	wire w_dff_A_PGrXCgsV6_0;
	wire w_dff_A_k8QWObmZ5_0;
	wire w_dff_A_PWmGEvrn1_0;
	wire w_dff_A_it6GNzsI2_0;
	wire w_dff_A_dY0mTyTs3_0;
	wire w_dff_A_XSgKg9OT8_1;
	wire w_dff_A_aY5NSo1j9_0;
	wire w_dff_A_i549ZAOL4_0;
	wire w_dff_A_sx55JEQH2_0;
	wire w_dff_A_lw3JEhUA7_1;
	wire w_dff_A_viqP63LY9_0;
	wire w_dff_A_yVUWWQzq4_0;
	wire w_dff_A_jCTZi0uI1_0;
	wire w_dff_A_qbIctODl9_1;
	wire w_dff_A_BnZP0qRU9_0;
	wire w_dff_A_ndrSBHWg4_0;
	wire w_dff_A_4DmmGz8o2_0;
	wire w_dff_A_0IWw5YRT1_1;
	wire w_dff_A_A80hFMiP3_2;
	wire w_dff_A_GxCQ8ad60_0;
	jnot g0000(.din(w_G77_4[2]),.dout(n72),.clk(gclk));
	jnot g0001(.din(w_G50_5[2]),.dout(n73),.clk(gclk));
	jnot g0002(.din(w_G58_5[2]),.dout(n74),.clk(gclk));
	jnot g0003(.din(w_G68_5[2]),.dout(n75),.clk(gclk));
	jand g0004(.dina(w_n75_2[1]),.dinb(w_n74_2[1]),.dout(n76),.clk(gclk));
	jand g0005(.dina(w_n76_0[1]),.dinb(w_n73_2[2]),.dout(n77),.clk(gclk));
	jand g0006(.dina(w_n77_0[1]),.dinb(w_n72_1[2]),.dout(w_dff_A_dvfHxH6U7_2),.clk(gclk));
	jnot g0007(.din(w_G87_3[2]),.dout(n79),.clk(gclk));
	jnot g0008(.din(w_G97_4[2]),.dout(n80),.clk(gclk));
	jnot g0009(.din(w_G107_4[1]),.dout(n81),.clk(gclk));
	jand g0010(.dina(w_n81_2[1]),.dinb(w_n80_1[2]),.dout(n82),.clk(gclk));
	jor g0011(.dina(n82),.dinb(w_n79_1[2]),.dout(G355_fa_),.clk(gclk));
	jnot g0012(.din(w_G250_0[2]),.dout(n84),.clk(gclk));
	jnot g0013(.din(w_G257_1[2]),.dout(n85),.clk(gclk));
	jnot g0014(.din(w_G264_0[2]),.dout(n86),.clk(gclk));
	jand g0015(.dina(w_n86_0[2]),.dinb(w_n85_0[1]),.dout(n87),.clk(gclk));
	jor g0016(.dina(n87),.dinb(w_n84_1[2]),.dout(n88),.clk(gclk));
	jnot g0017(.din(w_G13_2[1]),.dout(n89),.clk(gclk));
	jand g0018(.dina(w_n89_0[1]),.dinb(w_G1_2[1]),.dout(n90),.clk(gclk));
	jand g0019(.dina(w_n90_0[2]),.dinb(w_G20_6[2]),.dout(n91),.clk(gclk));
	jand g0020(.dina(w_n91_1[2]),.dinb(n88),.dout(n92),.clk(gclk));
	jor g0021(.dina(w_n85_0[0]),.dinb(w_n80_1[1]),.dout(n93),.clk(gclk));
	jnot g0022(.din(w_G244_1[1]),.dout(n94),.clk(gclk));
	jor g0023(.dina(w_n94_0[2]),.dinb(w_n72_1[1]),.dout(n95),.clk(gclk));
	jnot g0024(.din(w_G238_0[2]),.dout(n96),.clk(gclk));
	jor g0025(.dina(w_n96_0[2]),.dinb(w_n75_2[0]),.dout(n97),.clk(gclk));
	jand g0026(.dina(n97),.dinb(n95),.dout(n98),.clk(gclk));
	jnot g0027(.din(w_G226_1[2]),.dout(n99),.clk(gclk));
	jor g0028(.dina(n99),.dinb(w_n73_2[1]),.dout(n100),.clk(gclk));
	jand g0029(.dina(w_dff_B_EGuQuSgs1_0),.dinb(n98),.dout(n101),.clk(gclk));
	jand g0030(.dina(n101),.dinb(w_dff_B_hMorE4od6_1),.dout(n102),.clk(gclk));
	jnot g0031(.din(w_G232_1[2]),.dout(n103),.clk(gclk));
	jor g0032(.dina(n103),.dinb(w_n74_2[0]),.dout(n104),.clk(gclk));
	jnot g0033(.din(w_G116_5[2]),.dout(n105),.clk(gclk));
	jnot g0034(.din(w_G270_0[2]),.dout(n106),.clk(gclk));
	jor g0035(.dina(n106),.dinb(w_n105_1[1]),.dout(n107),.clk(gclk));
	jand g0036(.dina(n107),.dinb(n104),.dout(n108),.clk(gclk));
	jor g0037(.dina(w_n86_0[1]),.dinb(w_n81_2[0]),.dout(n109),.clk(gclk));
	jand g0038(.dina(w_dff_B_Ihv2Jms46_0),.dinb(n108),.dout(n110),.clk(gclk));
	jand g0039(.dina(w_G20_6[1]),.dinb(w_G1_2[0]),.dout(n111),.clk(gclk));
	jnot g0040(.din(w_n111_0[2]),.dout(n112),.clk(gclk));
	jor g0041(.dina(w_n84_1[1]),.dinb(w_n79_1[1]),.dout(n113),.clk(gclk));
	jand g0042(.dina(n113),.dinb(w_n112_0[1]),.dout(n114),.clk(gclk));
	jand g0043(.dina(w_dff_B_TDSDGv6d9_0),.dinb(n110),.dout(n115),.clk(gclk));
	jand g0044(.dina(n115),.dinb(n102),.dout(n116),.clk(gclk));
	jnot g0045(.din(w_n76_0[0]),.dout(n117),.clk(gclk));
	jand g0046(.dina(n117),.dinb(w_G50_5[1]),.dout(n118),.clk(gclk));
	jnot g0047(.din(w_n118_0[2]),.dout(n119),.clk(gclk));
	jand g0048(.dina(w_n111_0[1]),.dinb(w_G13_2[0]),.dout(n120),.clk(gclk));
	jand g0049(.dina(w_n120_0[1]),.dinb(n119),.dout(n121),.clk(gclk));
	jor g0050(.dina(n121),.dinb(n116),.dout(n122),.clk(gclk));
	jor g0051(.dina(n122),.dinb(w_dff_B_JvinlRL29_1),.dout(w_dff_A_JOEDEGQA0_2),.clk(gclk));
	jxor g0052(.dina(w_G270_0[1]),.dinb(w_n86_0[0]),.dout(n124),.clk(gclk));
	jxor g0053(.dina(w_G257_1[1]),.dinb(w_G250_0[1]),.dout(n125),.clk(gclk));
	jxor g0054(.dina(w_dff_B_Xy3Tfcgg6_0),.dinb(n124),.dout(n126),.clk(gclk));
	jnot g0055(.din(w_n126_0[1]),.dout(n127),.clk(gclk));
	jxor g0056(.dina(w_G244_1[0]),.dinb(w_n96_0[1]),.dout(n128),.clk(gclk));
	jxor g0057(.dina(w_G232_1[1]),.dinb(w_G226_1[1]),.dout(n129),.clk(gclk));
	jxor g0058(.dina(w_dff_B_dVKmhsVS6_0),.dinb(n128),.dout(n130),.clk(gclk));
	jxor g0059(.dina(w_n130_0[1]),.dinb(n127),.dout(w_dff_A_IRozgalU2_2),.clk(gclk));
	jxor g0060(.dina(w_G58_5[1]),.dinb(w_G50_5[0]),.dout(n132),.clk(gclk));
	jxor g0061(.dina(w_G77_4[1]),.dinb(w_G68_5[1]),.dout(n133),.clk(gclk));
	jxor g0062(.dina(n133),.dinb(n132),.dout(n134),.clk(gclk));
	jxor g0063(.dina(w_G116_5[1]),.dinb(w_n81_1[2]),.dout(n135),.clk(gclk));
	jxor g0064(.dina(w_G97_4[1]),.dinb(w_G87_3[1]),.dout(n136),.clk(gclk));
	jxor g0065(.dina(w_dff_B_3sc9Ecjf8_0),.dinb(n135),.dout(n137),.clk(gclk));
	jxor g0066(.dina(w_n137_0[1]),.dinb(w_n134_0[1]),.dout(w_dff_A_rJIYourm4_2),.clk(gclk));
	jand g0067(.dina(w_G13_1[2]),.dinb(w_G1_1[2]),.dout(n139),.clk(gclk));
	jand g0068(.dina(w_n111_0[0]),.dinb(w_G33_12[2]),.dout(n140),.clk(gclk));
	jor g0069(.dina(w_n140_0[1]),.dinb(w_n139_1[2]),.dout(n141),.clk(gclk));
	jnot g0070(.din(w_G1_1[1]),.dout(n142),.clk(gclk));
	jand g0071(.dina(w_G13_1[1]),.dinb(w_n142_2[1]),.dout(n143),.clk(gclk));
	jand g0072(.dina(w_n143_0[1]),.dinb(w_G20_6[0]),.dout(n144),.clk(gclk));
	jor g0073(.dina(w_n144_2[1]),.dinb(w_n141_3[1]),.dout(n145),.clk(gclk));
	jand g0074(.dina(w_G33_12[1]),.dinb(w_n142_2[0]),.dout(n146),.clk(gclk));
	jor g0075(.dina(w_dff_B_l2pSoTrH7_0),.dinb(n145),.dout(n147),.clk(gclk));
	jnot g0076(.din(w_n147_0[2]),.dout(n148),.clk(gclk));
	jand g0077(.dina(w_n148_0[1]),.dinb(w_G116_5[0]),.dout(n149),.clk(gclk));
	jand g0078(.dina(w_G116_4[2]),.dinb(w_G20_5[2]),.dout(n150),.clk(gclk));
	jnot g0079(.din(w_G20_5[1]),.dout(n151),.clk(gclk));
	jand g0080(.dina(w_G283_3[2]),.dinb(w_G33_12[0]),.dout(n152),.clk(gclk));
	jnot g0081(.din(w_G33_11[2]),.dout(n153),.clk(gclk));
	jand g0082(.dina(w_G97_4[0]),.dinb(w_n153_8[1]),.dout(n154),.clk(gclk));
	jor g0083(.dina(n154),.dinb(w_n152_0[2]),.dout(n155),.clk(gclk));
	jand g0084(.dina(n155),.dinb(w_n151_6[1]),.dout(n156),.clk(gclk));
	jor g0085(.dina(n156),.dinb(w_dff_B_ThrNonlU3_1),.dout(n157),.clk(gclk));
	jand g0086(.dina(n157),.dinb(w_n141_3[0]),.dout(n158),.clk(gclk));
	jand g0087(.dina(w_n144_2[0]),.dinb(w_n105_1[0]),.dout(n159),.clk(gclk));
	jor g0088(.dina(w_dff_B_hEwfdFJC4_0),.dinb(n158),.dout(n160),.clk(gclk));
	jor g0089(.dina(n160),.dinb(n149),.dout(n161),.clk(gclk));
	jnot g0090(.din(w_n161_0[2]),.dout(n162),.clk(gclk));
	jnot g0091(.din(w_G41_0[2]),.dout(n163),.clk(gclk));
	jand g0092(.dina(w_G45_1[1]),.dinb(w_n142_1[2]),.dout(n164),.clk(gclk));
	jand g0093(.dina(w_n164_0[2]),.dinb(w_n163_1[1]),.dout(n165),.clk(gclk));
	jnot g0094(.din(w_n139_1[1]),.dout(n166),.clk(gclk));
	jand g0095(.dina(w_G41_0[1]),.dinb(w_G33_11[1]),.dout(n167),.clk(gclk));
	jor g0096(.dina(w_n167_0[1]),.dinb(n166),.dout(n168),.clk(gclk));
	jand g0097(.dina(w_n168_5[1]),.dinb(w_G274_0[2]),.dout(n169),.clk(gclk));
	jand g0098(.dina(w_n169_0[1]),.dinb(w_n165_0[1]),.dout(n170),.clk(gclk));
	jnot g0099(.din(w_n167_0[0]),.dout(n171),.clk(gclk));
	jand g0100(.dina(n171),.dinb(w_n139_1[0]),.dout(n172),.clk(gclk));
	jand g0101(.dina(w_G1698_0[2]),.dinb(w_n153_8[0]),.dout(n173),.clk(gclk));
	jand g0102(.dina(w_n173_3[1]),.dinb(w_G264_0[1]),.dout(n174),.clk(gclk));
	jand g0103(.dina(w_G303_2[2]),.dinb(w_G33_11[0]),.dout(n175),.clk(gclk));
	jnot g0104(.din(w_G1698_0[1]),.dout(n176),.clk(gclk));
	jand g0105(.dina(w_n176_0[1]),.dinb(w_n153_7[2]),.dout(n177),.clk(gclk));
	jand g0106(.dina(w_n177_1[2]),.dinb(w_G257_1[0]),.dout(n178),.clk(gclk));
	jor g0107(.dina(n178),.dinb(w_dff_B_Qf4tPweB9_1),.dout(n179),.clk(gclk));
	jor g0108(.dina(n179),.dinb(w_dff_B_RrvFTnon4_1),.dout(n180),.clk(gclk));
	jand g0109(.dina(n180),.dinb(w_n172_4[2]),.dout(n181),.clk(gclk));
	jnot g0110(.din(w_n165_0[0]),.dout(n182),.clk(gclk));
	jand g0111(.dina(w_n168_5[0]),.dinb(w_G270_0[0]),.dout(n183),.clk(gclk));
	jand g0112(.dina(n183),.dinb(w_n182_1[1]),.dout(n184),.clk(gclk));
	jor g0113(.dina(w_dff_B_Tqm4dI2w6_0),.dinb(n181),.dout(n185),.clk(gclk));
	jor g0114(.dina(n185),.dinb(w_n170_0[2]),.dout(n186),.clk(gclk));
	jand g0115(.dina(w_n186_1[2]),.dinb(w_G169_3[1]),.dout(n187),.clk(gclk));
	jnot g0116(.din(n187),.dout(n188),.clk(gclk));
	jnot g0117(.din(w_G179_2[2]),.dout(n189),.clk(gclk));
	jor g0118(.dina(w_n186_1[1]),.dinb(w_n189_2[2]),.dout(n190),.clk(gclk));
	jand g0119(.dina(w_n190_0[1]),.dinb(n188),.dout(n191),.clk(gclk));
	jor g0120(.dina(n191),.dinb(w_dff_B_OEsLG4yF6_1),.dout(n192),.clk(gclk));
	jand g0121(.dina(w_n186_1[0]),.dinb(w_G200_3[1]),.dout(n193),.clk(gclk));
	jnot g0122(.din(w_n186_0[2]),.dout(n194),.clk(gclk));
	jand g0123(.dina(n194),.dinb(w_G190_4[2]),.dout(n195),.clk(gclk));
	jor g0124(.dina(n195),.dinb(w_n161_0[1]),.dout(n196),.clk(gclk));
	jor g0125(.dina(n196),.dinb(w_dff_B_cuojKOfz4_1),.dout(n197),.clk(gclk));
	jand g0126(.dina(n197),.dinb(w_n192_0[2]),.dout(n198),.clk(gclk));
	jnot g0127(.din(w_G169_3[0]),.dout(n199),.clk(gclk));
	jand g0128(.dina(w_n168_4[2]),.dinb(w_G264_0[0]),.dout(n200),.clk(gclk));
	jand g0129(.dina(n200),.dinb(w_n182_1[0]),.dout(n201),.clk(gclk));
	jand g0130(.dina(w_n173_3[0]),.dinb(w_G257_0[2]),.dout(n202),.clk(gclk));
	jand g0131(.dina(w_G294_3[1]),.dinb(w_G33_10[2]),.dout(n203),.clk(gclk));
	jnot g0132(.din(n203),.dout(n204),.clk(gclk));
	jor g0133(.dina(w_G1698_0[0]),.dinb(w_G33_10[1]),.dout(n205),.clk(gclk));
	jor g0134(.dina(w_n205_1[1]),.dinb(w_n84_1[0]),.dout(n206),.clk(gclk));
	jand g0135(.dina(n206),.dinb(n204),.dout(n207),.clk(gclk));
	jnot g0136(.din(w_n207_0[1]),.dout(n208),.clk(gclk));
	jor g0137(.dina(n208),.dinb(w_n202_0[1]),.dout(n209),.clk(gclk));
	jand g0138(.dina(n209),.dinb(w_n172_4[1]),.dout(n210),.clk(gclk));
	jor g0139(.dina(n210),.dinb(w_n170_0[1]),.dout(n211),.clk(gclk));
	jor g0140(.dina(n211),.dinb(w_n201_0[1]),.dout(n212),.clk(gclk));
	jand g0141(.dina(w_n212_1[1]),.dinb(w_n199_0[2]),.dout(n213),.clk(gclk));
	jand g0142(.dina(w_n148_0[0]),.dinb(w_G107_4[0]),.dout(n214),.clk(gclk));
	jor g0143(.dina(w_n140_0[0]),.dinb(w_G13_1[0]),.dout(n215),.clk(gclk));
	jand g0144(.dina(w_n81_1[1]),.dinb(w_G20_5[0]),.dout(n216),.clk(gclk));
	jand g0145(.dina(w_dff_B_LiSmy9oS4_0),.dinb(w_n215_0[1]),.dout(n217),.clk(gclk));
	jand g0146(.dina(w_G116_4[1]),.dinb(w_G33_10[0]),.dout(n218),.clk(gclk));
	jand g0147(.dina(w_G87_3[0]),.dinb(w_n153_7[1]),.dout(n219),.clk(gclk));
	jor g0148(.dina(n219),.dinb(w_n218_0[1]),.dout(n220),.clk(gclk));
	jand g0149(.dina(n220),.dinb(w_n141_2[2]),.dout(n221),.clk(gclk));
	jand g0150(.dina(n221),.dinb(w_n151_6[0]),.dout(n222),.clk(gclk));
	jor g0151(.dina(n222),.dinb(w_dff_B_8kuGAAZk2_1),.dout(n223),.clk(gclk));
	jor g0152(.dina(w_dff_B_AiBGyhXP0_0),.dinb(n214),.dout(n224),.clk(gclk));
	jnot g0153(.din(w_n224_1[1]),.dout(n225),.clk(gclk));
	jnot g0154(.din(w_n201_0[0]),.dout(n226),.clk(gclk));
	jnot g0155(.din(w_G274_0[1]),.dout(n227),.clk(gclk));
	jor g0156(.dina(w_n172_4[0]),.dinb(w_dff_B_mypaOipd7_1),.dout(n228),.clk(gclk));
	jor g0157(.dina(n228),.dinb(w_n182_0[2]),.dout(n229),.clk(gclk));
	jnot g0158(.din(w_n202_0[0]),.dout(n230),.clk(gclk));
	jand g0159(.dina(w_n207_0[0]),.dinb(n230),.dout(n231),.clk(gclk));
	jor g0160(.dina(n231),.dinb(w_n168_4[1]),.dout(n232),.clk(gclk));
	jand g0161(.dina(n232),.dinb(w_n229_0[1]),.dout(n233),.clk(gclk));
	jand g0162(.dina(n233),.dinb(w_dff_B_VZM5CY1Z9_1),.dout(n234),.clk(gclk));
	jand g0163(.dina(w_n234_1[1]),.dinb(w_n189_2[1]),.dout(n235),.clk(gclk));
	jor g0164(.dina(n235),.dinb(w_n225_0[1]),.dout(n236),.clk(gclk));
	jor g0165(.dina(n236),.dinb(w_n213_0[1]),.dout(n237),.clk(gclk));
	jand g0166(.dina(w_n234_1[0]),.dinb(w_G190_4[1]),.dout(n238),.clk(gclk));
	jand g0167(.dina(w_n212_1[0]),.dinb(w_G200_3[0]),.dout(n239),.clk(gclk));
	jor g0168(.dina(n239),.dinb(w_n224_1[0]),.dout(n240),.clk(gclk));
	jor g0169(.dina(n240),.dinb(w_n238_0[1]),.dout(n241),.clk(gclk));
	jand g0170(.dina(n241),.dinb(w_n237_0[2]),.dout(n242),.clk(gclk));
	jand g0171(.dina(w_n173_2[2]),.dinb(w_G244_0[2]),.dout(n243),.clk(gclk));
	jnot g0172(.din(w_n243_0[1]),.dout(n244),.clk(gclk));
	jnot g0173(.din(w_n218_0[0]),.dout(n245),.clk(gclk));
	jor g0174(.dina(w_n205_1[0]),.dinb(w_n96_0[0]),.dout(n246),.clk(gclk));
	jand g0175(.dina(n246),.dinb(n245),.dout(n247),.clk(gclk));
	jand g0176(.dina(w_n247_0[1]),.dinb(n244),.dout(n248),.clk(gclk));
	jand g0177(.dina(n248),.dinb(w_n172_3[2]),.dout(n249),.clk(gclk));
	jor g0178(.dina(w_n164_0[1]),.dinb(w_n84_0[2]),.dout(n250),.clk(gclk));
	jand g0179(.dina(w_n164_0[0]),.dinb(w_G274_0[0]),.dout(n251),.clk(gclk));
	jnot g0180(.din(w_n251_0[1]),.dout(n252),.clk(gclk));
	jand g0181(.dina(n252),.dinb(w_n250_0[1]),.dout(n253),.clk(gclk));
	jand g0182(.dina(n253),.dinb(w_n168_4[0]),.dout(n254),.clk(gclk));
	jor g0183(.dina(n254),.dinb(n249),.dout(n255),.clk(gclk));
	jand g0184(.dina(w_n255_1[1]),.dinb(w_n189_2[0]),.dout(n256),.clk(gclk));
	jor g0185(.dina(w_n147_0[1]),.dinb(w_n79_1[0]),.dout(n257),.clk(gclk));
	jand g0186(.dina(w_n80_1[0]),.dinb(w_n79_0[2]),.dout(n258),.clk(gclk));
	jand g0187(.dina(n258),.dinb(w_n81_1[0]),.dout(n259),.clk(gclk));
	jand g0188(.dina(w_n259_0[1]),.dinb(w_G20_4[2]),.dout(n260),.clk(gclk));
	jnot g0189(.din(w_n141_2[1]),.dout(n261),.clk(gclk));
	jand g0190(.dina(w_G97_3[2]),.dinb(w_G33_9[2]),.dout(n262),.clk(gclk));
	jnot g0191(.din(w_n262_0[2]),.dout(n263),.clk(gclk));
	jor g0192(.dina(w_n75_1[2]),.dinb(w_G33_9[1]),.dout(n264),.clk(gclk));
	jand g0193(.dina(n264),.dinb(w_n151_5[2]),.dout(n265),.clk(gclk));
	jand g0194(.dina(n265),.dinb(w_dff_B_teAz4mHt2_1),.dout(n266),.clk(gclk));
	jor g0195(.dina(n266),.dinb(w_n261_1[2]),.dout(n267),.clk(gclk));
	jor g0196(.dina(n267),.dinb(w_n260_0[1]),.dout(n268),.clk(gclk));
	jand g0197(.dina(w_n144_1[2]),.dinb(w_n79_0[1]),.dout(n269),.clk(gclk));
	jnot g0198(.din(w_n269_0[1]),.dout(n270),.clk(gclk));
	jand g0199(.dina(w_dff_B_Z5BUScwi0_0),.dinb(n268),.dout(n271),.clk(gclk));
	jand g0200(.dina(n271),.dinb(w_n257_0[1]),.dout(n272),.clk(gclk));
	jnot g0201(.din(w_n247_0[0]),.dout(n273),.clk(gclk));
	jor g0202(.dina(n273),.dinb(w_n243_0[0]),.dout(n274),.clk(gclk));
	jor g0203(.dina(n274),.dinb(w_n168_3[2]),.dout(n275),.clk(gclk));
	jnot g0204(.din(w_n250_0[0]),.dout(n276),.clk(gclk));
	jor g0205(.dina(w_n251_0[0]),.dinb(n276),.dout(n277),.clk(gclk));
	jor g0206(.dina(n277),.dinb(w_n172_3[1]),.dout(n278),.clk(gclk));
	jand g0207(.dina(n278),.dinb(n275),.dout(n279),.clk(gclk));
	jand g0208(.dina(w_n279_1[1]),.dinb(w_n199_0[1]),.dout(n280),.clk(gclk));
	jor g0209(.dina(n280),.dinb(w_n272_0[1]),.dout(n281),.clk(gclk));
	jor g0210(.dina(n281),.dinb(w_n256_0[1]),.dout(n282),.clk(gclk));
	jand g0211(.dina(w_n279_1[0]),.dinb(w_G200_2[2]),.dout(n283),.clk(gclk));
	jnot g0212(.din(w_n257_0[0]),.dout(n284),.clk(gclk));
	jnot g0213(.din(w_n260_0[0]),.dout(n285),.clk(gclk));
	jand g0214(.dina(w_G68_5[0]),.dinb(w_n153_7[0]),.dout(n286),.clk(gclk));
	jor g0215(.dina(n286),.dinb(w_G20_4[1]),.dout(n287),.clk(gclk));
	jor g0216(.dina(n287),.dinb(w_n262_0[1]),.dout(n288),.clk(gclk));
	jand g0217(.dina(n288),.dinb(w_n141_2[0]),.dout(n289),.clk(gclk));
	jand g0218(.dina(n289),.dinb(n285),.dout(n290),.clk(gclk));
	jor g0219(.dina(w_n269_0[0]),.dinb(n290),.dout(n291),.clk(gclk));
	jor g0220(.dina(n291),.dinb(n284),.dout(n292),.clk(gclk));
	jand g0221(.dina(w_n255_1[0]),.dinb(w_G190_4[0]),.dout(n293),.clk(gclk));
	jor g0222(.dina(n293),.dinb(w_n292_0[2]),.dout(n294),.clk(gclk));
	jor g0223(.dina(n294),.dinb(w_n283_0[1]),.dout(n295),.clk(gclk));
	jand g0224(.dina(n295),.dinb(w_n282_0[1]),.dout(n296),.clk(gclk));
	jand g0225(.dina(w_n168_3[1]),.dinb(w_G257_0[1]),.dout(n297),.clk(gclk));
	jand g0226(.dina(n297),.dinb(w_n182_0[1]),.dout(n298),.clk(gclk));
	jnot g0227(.din(w_n298_0[1]),.dout(n299),.clk(gclk));
	jor g0228(.dina(w_n176_0[0]),.dinb(w_G33_9[0]),.dout(n300),.clk(gclk));
	jor g0229(.dina(n300),.dinb(w_n84_0[1]),.dout(n301),.clk(gclk));
	jnot g0230(.din(w_n152_0[1]),.dout(n302),.clk(gclk));
	jor g0231(.dina(w_n205_0[2]),.dinb(w_n94_0[1]),.dout(n303),.clk(gclk));
	jand g0232(.dina(n303),.dinb(n302),.dout(n304),.clk(gclk));
	jand g0233(.dina(n304),.dinb(n301),.dout(n305),.clk(gclk));
	jor g0234(.dina(n305),.dinb(w_n168_3[0]),.dout(n306),.clk(gclk));
	jand g0235(.dina(n306),.dinb(w_n229_0[0]),.dout(n307),.clk(gclk));
	jand g0236(.dina(n307),.dinb(n299),.dout(n308),.clk(gclk));
	jand g0237(.dina(w_n308_1[2]),.dinb(w_G190_3[2]),.dout(n309),.clk(gclk));
	jor g0238(.dina(w_n147_0[0]),.dinb(w_n80_0[2]),.dout(n310),.clk(gclk));
	jnot g0239(.din(w_n310_0[1]),.dout(n311),.clk(gclk));
	jxor g0240(.dina(w_G107_3[2]),.dinb(w_G97_3[1]),.dout(n312),.clk(gclk));
	jand g0241(.dina(w_n312_0[1]),.dinb(w_G20_4[0]),.dout(n313),.clk(gclk));
	jnot g0242(.din(w_n313_0[1]),.dout(n314),.clk(gclk));
	jand g0243(.dina(w_G107_3[1]),.dinb(w_G33_8[2]),.dout(n315),.clk(gclk));
	jand g0244(.dina(w_G77_4[0]),.dinb(w_n153_6[2]),.dout(n316),.clk(gclk));
	jor g0245(.dina(n316),.dinb(w_G20_3[2]),.dout(n317),.clk(gclk));
	jor g0246(.dina(n317),.dinb(w_n315_0[2]),.dout(n318),.clk(gclk));
	jand g0247(.dina(n318),.dinb(w_n141_1[2]),.dout(n319),.clk(gclk));
	jand g0248(.dina(n319),.dinb(w_dff_B_llEH8sKq5_1),.dout(n320),.clk(gclk));
	jand g0249(.dina(w_n144_1[1]),.dinb(w_n80_0[1]),.dout(n321),.clk(gclk));
	jor g0250(.dina(w_n321_0[1]),.dinb(n320),.dout(n322),.clk(gclk));
	jor g0251(.dina(n322),.dinb(n311),.dout(n323),.clk(gclk));
	jand g0252(.dina(w_n173_2[1]),.dinb(w_G250_0[0]),.dout(n324),.clk(gclk));
	jand g0253(.dina(w_n177_1[1]),.dinb(w_G244_0[1]),.dout(n325),.clk(gclk));
	jor g0254(.dina(n325),.dinb(w_n152_0[0]),.dout(n326),.clk(gclk));
	jor g0255(.dina(n326),.dinb(w_dff_B_O8VhvD2i9_1),.dout(n327),.clk(gclk));
	jand g0256(.dina(n327),.dinb(w_n172_3[0]),.dout(n328),.clk(gclk));
	jor g0257(.dina(n328),.dinb(w_n170_0[0]),.dout(n329),.clk(gclk));
	jor g0258(.dina(n329),.dinb(w_n298_0[0]),.dout(n330),.clk(gclk));
	jand g0259(.dina(w_n330_0[2]),.dinb(w_G200_2[1]),.dout(n331),.clk(gclk));
	jor g0260(.dina(n331),.dinb(w_n323_0[2]),.dout(n332),.clk(gclk));
	jor g0261(.dina(n332),.dinb(w_n309_0[1]),.dout(n333),.clk(gclk));
	jor g0262(.dina(w_n308_1[1]),.dinb(w_G169_2[2]),.dout(n334),.clk(gclk));
	jnot g0263(.din(w_n334_0[1]),.dout(n335),.clk(gclk));
	jnot g0264(.din(w_n315_0[1]),.dout(n336),.clk(gclk));
	jor g0265(.dina(w_n72_1[0]),.dinb(w_G33_8[1]),.dout(n337),.clk(gclk));
	jand g0266(.dina(n337),.dinb(w_n151_5[1]),.dout(n338),.clk(gclk));
	jand g0267(.dina(n338),.dinb(w_dff_B_BKOW30cU3_1),.dout(n339),.clk(gclk));
	jor g0268(.dina(n339),.dinb(w_n261_1[1]),.dout(n340),.clk(gclk));
	jor g0269(.dina(n340),.dinb(w_n313_0[0]),.dout(n341),.clk(gclk));
	jnot g0270(.din(w_n321_0[0]),.dout(n342),.clk(gclk));
	jand g0271(.dina(w_dff_B_uHyrMRuq9_0),.dinb(n341),.dout(n343),.clk(gclk));
	jand g0272(.dina(n343),.dinb(w_n310_0[0]),.dout(n344),.clk(gclk));
	jand g0273(.dina(w_n308_1[0]),.dinb(w_n189_1[2]),.dout(n345),.clk(gclk));
	jor g0274(.dina(n345),.dinb(w_n344_0[1]),.dout(n346),.clk(gclk));
	jor g0275(.dina(n346),.dinb(n335),.dout(n347),.clk(gclk));
	jand g0276(.dina(w_n347_0[1]),.dinb(w_n333_0[1]),.dout(n348),.clk(gclk));
	jand g0277(.dina(w_n348_0[1]),.dinb(w_dff_B_wffm9AH96_1),.dout(n349),.clk(gclk));
	jand g0278(.dina(w_n349_0[1]),.dinb(w_n242_0[2]),.dout(n350),.clk(gclk));
	jand g0279(.dina(w_n350_0[1]),.dinb(w_n198_0[2]),.dout(n351),.clk(gclk));
	jnot g0280(.din(w_G45_1[0]),.dout(n352),.clk(gclk));
	jand g0281(.dina(w_n352_1[1]),.dinb(w_n163_1[0]),.dout(n353),.clk(gclk));
	jor g0282(.dina(n353),.dinb(w_G1_1[0]),.dout(n354),.clk(gclk));
	jnot g0283(.din(w_n354_1[1]),.dout(n355),.clk(gclk));
	jand g0284(.dina(w_n355_0[1]),.dinb(w_n169_0[0]),.dout(n356),.clk(gclk));
	jnot g0285(.din(w_n356_1[1]),.dout(n357),.clk(gclk));
	jand g0286(.dina(w_n173_2[0]),.dinb(w_G238_0[1]),.dout(n358),.clk(gclk));
	jand g0287(.dina(w_n177_1[0]),.dinb(w_G232_1[0]),.dout(n359),.clk(gclk));
	jor g0288(.dina(n359),.dinb(w_n315_0[0]),.dout(n360),.clk(gclk));
	jor g0289(.dina(n360),.dinb(w_dff_B_5pQ1P8OX7_1),.dout(n361),.clk(gclk));
	jand g0290(.dina(n361),.dinb(w_n172_2[2]),.dout(n362),.clk(gclk));
	jnot g0291(.din(n362),.dout(n363),.clk(gclk));
	jor g0292(.dina(w_n355_0[0]),.dinb(w_n94_0[0]),.dout(n364),.clk(gclk));
	jor g0293(.dina(n364),.dinb(w_n172_2[1]),.dout(n365),.clk(gclk));
	jand g0294(.dina(w_dff_B_Q1nhhtqB4_0),.dinb(n363),.dout(n366),.clk(gclk));
	jand g0295(.dina(n366),.dinb(w_n357_0[1]),.dout(n367),.clk(gclk));
	jnot g0296(.din(w_n367_1[1]),.dout(n368),.clk(gclk));
	jand g0297(.dina(n368),.dinb(w_n199_0[0]),.dout(n369),.clk(gclk));
	jand g0298(.dina(w_G87_2[2]),.dinb(w_G33_8[0]),.dout(n370),.clk(gclk));
	jand g0299(.dina(w_G58_5[0]),.dinb(w_n153_6[1]),.dout(n371),.clk(gclk));
	jor g0300(.dina(n371),.dinb(w_n370_0[1]),.dout(n372),.clk(gclk));
	jand g0301(.dina(n372),.dinb(w_n151_5[0]),.dout(n373),.clk(gclk));
	jand g0302(.dina(n373),.dinb(w_n141_1[1]),.dout(n374),.clk(gclk));
	jand g0303(.dina(w_n139_0[2]),.dinb(w_n151_4[2]),.dout(n375),.clk(gclk));
	jnot g0304(.din(w_n375_0[1]),.dout(n376),.clk(gclk));
	jand g0305(.dina(w_G20_3[1]),.dinb(w_n142_1[1]),.dout(n377),.clk(gclk));
	jnot g0306(.din(n377),.dout(n378),.clk(gclk));
	jand g0307(.dina(w_n378_0[1]),.dinb(w_G77_3[2]),.dout(n379),.clk(gclk));
	jand g0308(.dina(n379),.dinb(w_dff_B_62Ls3ksn7_1),.dout(n380),.clk(gclk));
	jand g0309(.dina(w_n144_1[0]),.dinb(w_n72_0[2]),.dout(n381),.clk(gclk));
	jor g0310(.dina(w_dff_B_eQWyAsEn2_0),.dinb(n380),.dout(n382),.clk(gclk));
	jor g0311(.dina(n382),.dinb(w_dff_B_bxIqVvov8_1),.dout(n383),.clk(gclk));
	jnot g0312(.din(w_n383_0[2]),.dout(n384),.clk(gclk));
	jand g0313(.dina(w_n367_1[0]),.dinb(w_n189_1[1]),.dout(n385),.clk(gclk));
	jor g0314(.dina(n385),.dinb(w_dff_B_tHyOvIpT5_1),.dout(n386),.clk(gclk));
	jor g0315(.dina(n386),.dinb(n369),.dout(n387),.clk(gclk));
	jnot g0316(.din(w_G200_2[0]),.dout(n388),.clk(gclk));
	jor g0317(.dina(w_n367_0[2]),.dinb(w_n388_2[1]),.dout(n389),.clk(gclk));
	jnot g0318(.din(n389),.dout(n390),.clk(gclk));
	jand g0319(.dina(w_n367_0[1]),.dinb(w_G190_3[1]),.dout(n391),.clk(gclk));
	jor g0320(.dina(n391),.dinb(w_n383_0[1]),.dout(n392),.clk(gclk));
	jor g0321(.dina(n392),.dinb(n390),.dout(n393),.clk(gclk));
	jand g0322(.dina(n393),.dinb(w_n387_0[2]),.dout(n394),.clk(gclk));
	jnot g0323(.din(w_n394_0[1]),.dout(n395),.clk(gclk));
	jand g0324(.dina(w_n168_2[2]),.dinb(w_G238_0[0]),.dout(n396),.clk(gclk));
	jand g0325(.dina(n396),.dinb(w_n354_1[0]),.dout(n397),.clk(gclk));
	jand g0326(.dina(w_n173_1[2]),.dinb(w_G232_0[2]),.dout(n398),.clk(gclk));
	jand g0327(.dina(w_n177_0[2]),.dinb(w_G226_1[0]),.dout(n399),.clk(gclk));
	jor g0328(.dina(n399),.dinb(w_n262_0[0]),.dout(n400),.clk(gclk));
	jor g0329(.dina(n400),.dinb(w_dff_B_yaVOpD0p0_1),.dout(n401),.clk(gclk));
	jand g0330(.dina(n401),.dinb(w_n172_2[0]),.dout(n402),.clk(gclk));
	jor g0331(.dina(n402),.dinb(w_n356_1[0]),.dout(n403),.clk(gclk));
	jor g0332(.dina(n403),.dinb(w_dff_B_A0x9HqyM7_1),.dout(n404),.clk(gclk));
	jnot g0333(.din(w_n404_0[2]),.dout(n405),.clk(gclk));
	jor g0334(.dina(w_n405_0[1]),.dinb(w_G169_2[1]),.dout(n406),.clk(gclk));
	jand g0335(.dina(w_G77_3[1]),.dinb(w_G33_7[2]),.dout(n407),.clk(gclk));
	jand g0336(.dina(w_G50_4[2]),.dinb(w_n153_6[0]),.dout(n408),.clk(gclk));
	jor g0337(.dina(n408),.dinb(w_n407_0[1]),.dout(n409),.clk(gclk));
	jand g0338(.dina(n409),.dinb(w_n141_1[0]),.dout(n410),.clk(gclk));
	jand g0339(.dina(n410),.dinb(w_n151_4[1]),.dout(n411),.clk(gclk));
	jand g0340(.dina(w_n75_1[1]),.dinb(w_G20_3[0]),.dout(n412),.clk(gclk));
	jand g0341(.dina(w_dff_B_cQDb0x8w8_0),.dinb(w_n215_0[0]),.dout(n413),.clk(gclk));
	jand g0342(.dina(w_n378_0[0]),.dinb(w_n261_1[0]),.dout(n414),.clk(gclk));
	jand g0343(.dina(w_n414_0[2]),.dinb(w_G68_4[2]),.dout(n415),.clk(gclk));
	jor g0344(.dina(n415),.dinb(w_dff_B_REqKySol5_1),.dout(n416),.clk(gclk));
	jor g0345(.dina(n416),.dinb(w_dff_B_ss6wQMSM1_1),.dout(n417),.clk(gclk));
	jor g0346(.dina(w_n404_0[1]),.dinb(w_G179_2[1]),.dout(n418),.clk(gclk));
	jand g0347(.dina(n418),.dinb(w_n417_0[2]),.dout(n419),.clk(gclk));
	jand g0348(.dina(n419),.dinb(n406),.dout(n420),.clk(gclk));
	jand g0349(.dina(w_n405_0[0]),.dinb(w_G190_3[0]),.dout(n421),.clk(gclk));
	jand g0350(.dina(w_n404_0[0]),.dinb(w_G200_1[2]),.dout(n422),.clk(gclk));
	jor g0351(.dina(n422),.dinb(w_n417_0[1]),.dout(n423),.clk(gclk));
	jor g0352(.dina(n423),.dinb(n421),.dout(n424),.clk(gclk));
	jnot g0353(.din(n424),.dout(n425),.clk(gclk));
	jor g0354(.dina(w_n425_0[1]),.dinb(w_n420_0[1]),.dout(n426),.clk(gclk));
	jand g0355(.dina(w_n168_2[1]),.dinb(w_G226_0[2]),.dout(n427),.clk(gclk));
	jand g0356(.dina(n427),.dinb(w_n354_0[2]),.dout(n428),.clk(gclk));
	jnot g0357(.din(w_n428_0[1]),.dout(n429),.clk(gclk));
	jand g0358(.dina(w_n173_1[1]),.dinb(w_G223_0[1]),.dout(n430),.clk(gclk));
	jnot g0359(.din(w_n430_0[1]),.dout(n431),.clk(gclk));
	jnot g0360(.din(w_n407_0[0]),.dout(n432),.clk(gclk));
	jnot g0361(.din(G222),.dout(n433),.clk(gclk));
	jor g0362(.dina(w_n205_0[1]),.dinb(n433),.dout(n434),.clk(gclk));
	jand g0363(.dina(n434),.dinb(n432),.dout(n435),.clk(gclk));
	jand g0364(.dina(w_n435_0[1]),.dinb(n431),.dout(n436),.clk(gclk));
	jor g0365(.dina(n436),.dinb(w_n168_2[0]),.dout(n437),.clk(gclk));
	jand g0366(.dina(n437),.dinb(w_n357_0[0]),.dout(n438),.clk(gclk));
	jand g0367(.dina(n438),.dinb(w_dff_B_2nIrxPWo3_1),.dout(n439),.clk(gclk));
	jor g0368(.dina(w_n439_0[2]),.dinb(w_G169_2[0]),.dout(n440),.clk(gclk));
	jand g0369(.dina(w_G33_7[1]),.dinb(w_n151_4[0]),.dout(n441),.clk(gclk));
	jand g0370(.dina(w_n441_0[1]),.dinb(w_G58_4[2]),.dout(n442),.clk(gclk));
	jnot g0371(.din(n442),.dout(n443),.clk(gclk));
	jor g0372(.dina(w_n77_0[0]),.dinb(w_n151_3[2]),.dout(n444),.clk(gclk));
	jand g0373(.dina(w_n153_5[2]),.dinb(w_n151_3[1]),.dout(n445),.clk(gclk));
	jand g0374(.dina(w_n445_0[1]),.dinb(w_G150_3[1]),.dout(n446),.clk(gclk));
	jnot g0375(.din(n446),.dout(n447),.clk(gclk));
	jand g0376(.dina(n447),.dinb(n444),.dout(n448),.clk(gclk));
	jand g0377(.dina(n448),.dinb(w_dff_B_EV0oZ51Q6_1),.dout(n449),.clk(gclk));
	jor g0378(.dina(n449),.dinb(w_n261_0[2]),.dout(n450),.clk(gclk));
	jnot g0379(.din(w_n450_0[1]),.dout(n451),.clk(gclk));
	jnot g0380(.din(w_n144_0[2]),.dout(n452),.clk(gclk));
	jand g0381(.dina(w_n452_0[1]),.dinb(w_n73_2[0]),.dout(n453),.clk(gclk));
	jnot g0382(.din(n453),.dout(n454),.clk(gclk));
	jor g0383(.dina(w_n414_0[1]),.dinb(w_n73_1[2]),.dout(n455),.clk(gclk));
	jand g0384(.dina(n455),.dinb(n454),.dout(n456),.clk(gclk));
	jor g0385(.dina(w_n456_0[1]),.dinb(n451),.dout(n457),.clk(gclk));
	jnot g0386(.din(w_n435_0[0]),.dout(n458),.clk(gclk));
	jor g0387(.dina(n458),.dinb(w_n430_0[0]),.dout(n459),.clk(gclk));
	jand g0388(.dina(n459),.dinb(w_n172_1[2]),.dout(n460),.clk(gclk));
	jor g0389(.dina(n460),.dinb(w_n356_0[2]),.dout(n461),.clk(gclk));
	jor g0390(.dina(n461),.dinb(w_n428_0[0]),.dout(n462),.clk(gclk));
	jor g0391(.dina(n462),.dinb(w_G179_2[0]),.dout(n463),.clk(gclk));
	jand g0392(.dina(n463),.dinb(w_n457_0[1]),.dout(n464),.clk(gclk));
	jand g0393(.dina(n464),.dinb(w_dff_B_K4FHGxx43_1),.dout(n465),.clk(gclk));
	jand g0394(.dina(w_n439_0[1]),.dinb(w_G190_2[2]),.dout(n466),.clk(gclk));
	jnot g0395(.din(n466),.dout(n467),.clk(gclk));
	jnot g0396(.din(w_n456_0[0]),.dout(n468),.clk(gclk));
	jand g0397(.dina(n468),.dinb(w_n450_0[0]),.dout(n469),.clk(gclk));
	jor g0398(.dina(w_n439_0[0]),.dinb(w_n388_2[0]),.dout(n470),.clk(gclk));
	jand g0399(.dina(n470),.dinb(n469),.dout(n471),.clk(gclk));
	jand g0400(.dina(n471),.dinb(n467),.dout(n472),.clk(gclk));
	jor g0401(.dina(w_n472_0[1]),.dinb(w_n465_0[1]),.dout(n473),.clk(gclk));
	jand g0402(.dina(w_n168_1[2]),.dinb(w_G232_0[1]),.dout(n474),.clk(gclk));
	jand g0403(.dina(n474),.dinb(w_n354_0[1]),.dout(n475),.clk(gclk));
	jand g0404(.dina(w_n173_1[0]),.dinb(w_G226_0[1]),.dout(n476),.clk(gclk));
	jand g0405(.dina(w_n177_0[1]),.dinb(w_G223_0[0]),.dout(n477),.clk(gclk));
	jor g0406(.dina(n477),.dinb(w_n370_0[0]),.dout(n478),.clk(gclk));
	jor g0407(.dina(n478),.dinb(w_dff_B_kJhu1W4f8_1),.dout(n479),.clk(gclk));
	jand g0408(.dina(n479),.dinb(w_n172_1[1]),.dout(n480),.clk(gclk));
	jor g0409(.dina(n480),.dinb(w_n356_0[1]),.dout(n481),.clk(gclk));
	jor g0410(.dina(n481),.dinb(w_dff_B_uIKuRZbo0_1),.dout(n482),.clk(gclk));
	jnot g0411(.din(w_n482_0[2]),.dout(n483),.clk(gclk));
	jor g0412(.dina(w_n483_0[1]),.dinb(w_G169_1[2]),.dout(n484),.clk(gclk));
	jnot g0413(.din(w_G159_3[2]),.dout(n485),.clk(gclk));
	jnot g0414(.din(w_n445_0[0]),.dout(n486),.clk(gclk));
	jor g0415(.dina(n486),.dinb(w_dff_B_vkJ7ryfr0_1),.dout(n487),.clk(gclk));
	jxor g0416(.dina(w_G68_4[1]),.dinb(w_G58_4[1]),.dout(n488),.clk(gclk));
	jor g0417(.dina(n488),.dinb(w_n151_3[0]),.dout(n489),.clk(gclk));
	jand g0418(.dina(w_n441_0[0]),.dinb(w_G68_4[0]),.dout(n490),.clk(gclk));
	jnot g0419(.din(n490),.dout(n491),.clk(gclk));
	jand g0420(.dina(n491),.dinb(w_dff_B_XwAHOEav0_1),.dout(n492),.clk(gclk));
	jand g0421(.dina(n492),.dinb(w_dff_B_61EjpAtY1_1),.dout(n493),.clk(gclk));
	jor g0422(.dina(n493),.dinb(w_n261_0[1]),.dout(n494),.clk(gclk));
	jnot g0423(.din(w_n494_0[1]),.dout(n495),.clk(gclk));
	jand g0424(.dina(w_n452_0[0]),.dinb(w_n74_1[2]),.dout(n496),.clk(gclk));
	jnot g0425(.din(n496),.dout(n497),.clk(gclk));
	jor g0426(.dina(w_n414_0[0]),.dinb(w_n74_1[1]),.dout(n498),.clk(gclk));
	jand g0427(.dina(n498),.dinb(n497),.dout(n499),.clk(gclk));
	jor g0428(.dina(w_n499_0[1]),.dinb(n495),.dout(n500),.clk(gclk));
	jor g0429(.dina(w_n482_0[1]),.dinb(w_G179_1[2]),.dout(n501),.clk(gclk));
	jand g0430(.dina(n501),.dinb(w_n500_0[1]),.dout(n502),.clk(gclk));
	jand g0431(.dina(n502),.dinb(n484),.dout(n503),.clk(gclk));
	jor g0432(.dina(w_n483_0[0]),.dinb(w_n388_1[2]),.dout(n504),.clk(gclk));
	jnot g0433(.din(w_n499_0[0]),.dout(n505),.clk(gclk));
	jand g0434(.dina(n505),.dinb(w_n494_0[0]),.dout(n506),.clk(gclk));
	jnot g0435(.din(w_G190_2[1]),.dout(n507),.clk(gclk));
	jor g0436(.dina(w_n482_0[0]),.dinb(w_n507_2[1]),.dout(n508),.clk(gclk));
	jand g0437(.dina(n508),.dinb(n506),.dout(n509),.clk(gclk));
	jand g0438(.dina(n509),.dinb(n504),.dout(n510),.clk(gclk));
	jor g0439(.dina(n510),.dinb(w_n503_0[2]),.dout(n511),.clk(gclk));
	jor g0440(.dina(w_n511_0[1]),.dinb(w_n473_0[1]),.dout(n512),.clk(gclk));
	jor g0441(.dina(w_n512_0[1]),.dinb(w_n426_0[1]),.dout(n513),.clk(gclk));
	jor g0442(.dina(n513),.dinb(w_n395_0[1]),.dout(n514),.clk(gclk));
	jnot g0443(.din(w_n514_1[1]),.dout(n515),.clk(gclk));
	jand g0444(.dina(n515),.dinb(w_n351_0[1]),.dout(w_dff_A_8Q6yYxeC8_2),.clk(gclk));
	jnot g0445(.din(w_n213_0[0]),.dout(n517),.clk(gclk));
	jor g0446(.dina(w_n212_0[2]),.dinb(w_G179_1[1]),.dout(n518),.clk(gclk));
	jand g0447(.dina(n518),.dinb(w_n224_0[2]),.dout(n519),.clk(gclk));
	jand g0448(.dina(n519),.dinb(n517),.dout(n520),.clk(gclk));
	jnot g0449(.din(w_n238_0[0]),.dout(n521),.clk(gclk));
	jor g0450(.dina(w_n234_0[2]),.dinb(w_n388_1[1]),.dout(n522),.clk(gclk));
	jand g0451(.dina(n522),.dinb(w_n225_0[0]),.dout(n523),.clk(gclk));
	jand g0452(.dina(n523),.dinb(n521),.dout(n524),.clk(gclk));
	jor g0453(.dina(n524),.dinb(w_n520_0[1]),.dout(n525),.clk(gclk));
	jnot g0454(.din(w_n256_0[0]),.dout(n526),.clk(gclk));
	jor g0455(.dina(w_n255_0[2]),.dinb(w_G169_1[1]),.dout(n527),.clk(gclk));
	jand g0456(.dina(n527),.dinb(w_n292_0[1]),.dout(n528),.clk(gclk));
	jand g0457(.dina(n528),.dinb(n526),.dout(n529),.clk(gclk));
	jnot g0458(.din(w_n283_0[0]),.dout(n530),.clk(gclk));
	jor g0459(.dina(w_n279_0[2]),.dinb(w_n507_2[0]),.dout(n531),.clk(gclk));
	jand g0460(.dina(n531),.dinb(w_n272_0[0]),.dout(n532),.clk(gclk));
	jand g0461(.dina(n532),.dinb(n530),.dout(n533),.clk(gclk));
	jor g0462(.dina(w_n533_0[1]),.dinb(n529),.dout(n534),.clk(gclk));
	jnot g0463(.din(w_n309_0[0]),.dout(n535),.clk(gclk));
	jor g0464(.dina(w_n308_0[2]),.dinb(w_n388_1[0]),.dout(n536),.clk(gclk));
	jand g0465(.dina(n536),.dinb(w_n344_0[0]),.dout(n537),.clk(gclk));
	jand g0466(.dina(n537),.dinb(n535),.dout(n538),.clk(gclk));
	jor g0467(.dina(w_n330_0[1]),.dinb(w_G179_1[0]),.dout(n539),.clk(gclk));
	jand g0468(.dina(n539),.dinb(w_n323_0[1]),.dout(n540),.clk(gclk));
	jand g0469(.dina(n540),.dinb(w_n334_0[0]),.dout(n541),.clk(gclk));
	jor g0470(.dina(w_n541_0[1]),.dinb(w_dff_B_ei1IRPYu3_1),.dout(n542),.clk(gclk));
	jor g0471(.dina(w_n542_0[1]),.dinb(w_n534_0[1]),.dout(n543),.clk(gclk));
	jor g0472(.dina(w_n543_0[1]),.dinb(w_dff_B_F4cGoxfX8_1),.dout(n544),.clk(gclk));
	jor g0473(.dina(w_n544_0[1]),.dinb(w_n192_0[1]),.dout(n545),.clk(gclk));
	jor g0474(.dina(w_n543_0[0]),.dinb(w_n237_0[1]),.dout(n546),.clk(gclk));
	jor g0475(.dina(w_n347_0[0]),.dinb(w_n533_0[0]),.dout(n547),.clk(gclk));
	jand g0476(.dina(n547),.dinb(w_n282_0[0]),.dout(n548),.clk(gclk));
	jand g0477(.dina(w_n548_0[1]),.dinb(n546),.dout(n549),.clk(gclk));
	jand g0478(.dina(n549),.dinb(n545),.dout(n550),.clk(gclk));
	jor g0479(.dina(w_n550_0[1]),.dinb(w_n514_1[0]),.dout(n551),.clk(gclk));
	jnot g0480(.din(w_n551_0[1]),.dout(n552),.clk(gclk));
	jnot g0481(.din(w_n472_0[0]),.dout(n553),.clk(gclk));
	jand g0482(.dina(w_n503_0[1]),.dinb(n553),.dout(n554),.clk(gclk));
	jnot g0483(.din(n554),.dout(n555),.clk(gclk));
	jnot g0484(.din(w_n465_0[0]),.dout(n556),.clk(gclk));
	jnot g0485(.din(w_n420_0[0]),.dout(n557),.clk(gclk));
	jor g0486(.dina(w_n425_0[0]),.dinb(w_n387_0[1]),.dout(n558),.clk(gclk));
	jand g0487(.dina(n558),.dinb(w_dff_B_AibjIE2U8_1),.dout(n559),.clk(gclk));
	jor g0488(.dina(w_n559_0[1]),.dinb(w_n512_0[0]),.dout(n560),.clk(gclk));
	jand g0489(.dina(n560),.dinb(w_dff_B_xhe3WgjF4_1),.dout(n561),.clk(gclk));
	jand g0490(.dina(n561),.dinb(w_dff_B_d2AqgI6h4_1),.dout(n562),.clk(gclk));
	jnot g0491(.din(w_n562_0[1]),.dout(n563),.clk(gclk));
	jor g0492(.dina(n563),.dinb(n552),.dout(w_dff_A_cLFUR3629_2),.clk(gclk));
	jand g0493(.dina(w_n143_0[0]),.dinb(w_G213_0[2]),.dout(n565),.clk(gclk));
	jand g0494(.dina(n565),.dinb(w_n151_2[2]),.dout(n566),.clk(gclk));
	jand g0495(.dina(w_n566_1[1]),.dinb(w_G343_0[1]),.dout(n567),.clk(gclk));
	jor g0496(.dina(w_n567_5[1]),.dinb(w_n237_0[0]),.dout(n568),.clk(gclk));
	jnot g0497(.din(n568),.dout(n569),.clk(gclk));
	jnot g0498(.din(w_n192_0[0]),.dout(n570),.clk(gclk));
	jnot g0499(.din(w_n567_5[0]),.dout(n571),.clk(gclk));
	jand g0500(.dina(w_n571_2[1]),.dinb(w_n570_0[1]),.dout(n572),.clk(gclk));
	jand g0501(.dina(w_n572_0[2]),.dinb(w_n242_0[1]),.dout(n573),.clk(gclk));
	jor g0502(.dina(w_n573_0[1]),.dinb(w_n569_0[1]),.dout(n574),.clk(gclk));
	jand g0503(.dina(w_n567_4[2]),.dinb(w_n161_0[0]),.dout(n575),.clk(gclk));
	jxor g0504(.dina(w_dff_B_QAuHnfYV8_0),.dinb(w_n198_0[1]),.dout(n576),.clk(gclk));
	jand g0505(.dina(w_n576_0[2]),.dinb(w_G330_0[2]),.dout(n577),.clk(gclk));
	jand g0506(.dina(w_n567_4[1]),.dinb(w_n224_0[1]),.dout(n578),.clk(gclk));
	jxor g0507(.dina(w_dff_B_w9d2YWfE9_0),.dinb(w_n242_0[0]),.dout(n579),.clk(gclk));
	jand g0508(.dina(w_n579_1[1]),.dinb(w_n577_0[1]),.dout(n580),.clk(gclk));
	jor g0509(.dina(w_n580_0[2]),.dinb(w_n574_0[1]),.dout(w_dff_A_dB0sU7VX1_2),.clk(gclk));
	jand g0510(.dina(w_n91_1[1]),.dinb(w_n163_0[2]),.dout(n582),.clk(gclk));
	jand g0511(.dina(w_n582_0[1]),.dinb(w_n118_0[1]),.dout(n583),.clk(gclk));
	jor g0512(.dina(w_n567_4[0]),.dinb(w_n550_0[0]),.dout(n584),.clk(gclk));
	jnot g0513(.din(w_n198_0[0]),.dout(n585),.clk(gclk));
	jor g0514(.dina(w_n544_0[0]),.dinb(n585),.dout(n586),.clk(gclk));
	jand g0515(.dina(w_n571_2[0]),.dinb(n586),.dout(n587),.clk(gclk));
	jnot g0516(.din(w_n190_0[0]),.dout(n588),.clk(gclk));
	jand g0517(.dina(w_n308_0[1]),.dinb(w_n255_0[1]),.dout(n589),.clk(gclk));
	jand g0518(.dina(w_dff_B_dlM9eFUA4_0),.dinb(n588),.dout(n590),.clk(gclk));
	jand g0519(.dina(n590),.dinb(w_n234_0[1]),.dout(n591),.clk(gclk));
	jand g0520(.dina(w_n279_0[1]),.dinb(w_n189_1[0]),.dout(n592),.clk(gclk));
	jand g0521(.dina(n592),.dinb(w_n330_0[0]),.dout(n593),.clk(gclk));
	jand g0522(.dina(n593),.dinb(w_n186_0[1]),.dout(n594),.clk(gclk));
	jand g0523(.dina(n594),.dinb(w_n212_0[1]),.dout(n595),.clk(gclk));
	jor g0524(.dina(n595),.dinb(w_n571_1[2]),.dout(n596),.clk(gclk));
	jor g0525(.dina(n596),.dinb(n591),.dout(n597),.clk(gclk));
	jand g0526(.dina(n597),.dinb(w_G330_0[1]),.dout(n598),.clk(gclk));
	jnot g0527(.din(w_n598_0[1]),.dout(n599),.clk(gclk));
	jor g0528(.dina(w_dff_B_lsLzXNMs1_0),.dinb(n587),.dout(n600),.clk(gclk));
	jand g0529(.dina(w_n600_1[2]),.dinb(w_n584_0[1]),.dout(n601),.clk(gclk));
	jnot g0530(.din(w_n601_0[2]),.dout(n602),.clk(gclk));
	jand g0531(.dina(w_n602_0[1]),.dinb(w_n142_1[0]),.dout(n603),.clk(gclk));
	jnot g0532(.din(w_n582_0[0]),.dout(n604),.clk(gclk));
	jand g0533(.dina(w_n259_0[0]),.dinb(w_n105_0[2]),.dout(n605),.clk(gclk));
	jand g0534(.dina(w_n605_0[2]),.dinb(w_G1_0[2]),.dout(n606),.clk(gclk));
	jand g0535(.dina(n606),.dinb(w_n604_2[2]),.dout(n607),.clk(gclk));
	jor g0536(.dina(w_dff_B_UReCyPV51_0),.dinb(n603),.dout(n608),.clk(gclk));
	jor g0537(.dina(n608),.dinb(w_dff_B_EQCVdU6e3_1),.dout(w_dff_A_pYXSlu0u3_2),.clk(gclk));
	jand g0538(.dina(w_G45_0[2]),.dinb(w_G13_0[2]),.dout(n610),.clk(gclk));
	jand g0539(.dina(n610),.dinb(w_n151_2[1]),.dout(n611),.clk(gclk));
	jor g0540(.dina(n611),.dinb(w_n142_0[2]),.dout(n612),.clk(gclk));
	jnot g0541(.din(n612),.dout(n613),.clk(gclk));
	jand g0542(.dina(w_n613_1[2]),.dinb(w_n604_2[1]),.dout(n614),.clk(gclk));
	jnot g0543(.din(w_n614_5[1]),.dout(n615),.clk(gclk));
	jxor g0544(.dina(w_n576_0[1]),.dinb(w_G330_0[0]),.dout(n616),.clk(gclk));
	jand g0545(.dina(n616),.dinb(w_dff_B_mecUk3Q59_1),.dout(n617),.clk(gclk));
	jand g0546(.dina(w_n153_5[1]),.dinb(w_n89_0[0]),.dout(n618),.clk(gclk));
	jand g0547(.dina(w_n618_2[1]),.dinb(w_n151_2[0]),.dout(n619),.clk(gclk));
	jnot g0548(.din(w_n619_0[2]),.dout(n620),.clk(gclk));
	jor g0549(.dina(w_n620_0[2]),.dinb(w_n576_0[0]),.dout(n621),.clk(gclk));
	jand g0550(.dina(w_n507_1[2]),.dinb(w_G20_2[2]),.dout(n622),.clk(gclk));
	jnot g0551(.din(w_n622_0[1]),.dout(n623),.clk(gclk));
	jand g0552(.dina(w_G200_1[1]),.dinb(w_G20_2[1]),.dout(n624),.clk(gclk));
	jnot g0553(.din(w_n624_0[1]),.dout(n625),.clk(gclk));
	jand g0554(.dina(w_G179_0[2]),.dinb(w_G20_2[0]),.dout(n626),.clk(gclk));
	jnot g0555(.din(w_n626_0[2]),.dout(n627),.clk(gclk));
	jand g0556(.dina(n627),.dinb(n625),.dout(n628),.clk(gclk));
	jand g0557(.dina(w_n628_0[1]),.dinb(n623),.dout(n629),.clk(gclk));
	jand g0558(.dina(w_n629_5[1]),.dinb(w_G97_3[0]),.dout(n630),.clk(gclk));
	jnot g0559(.din(w_n630_0[1]),.dout(n631),.clk(gclk));
	jand g0560(.dina(w_n624_0[0]),.dinb(w_n189_0[2]),.dout(n632),.clk(gclk));
	jand g0561(.dina(w_n632_0[1]),.dinb(w_G190_2[0]),.dout(n633),.clk(gclk));
	jand g0562(.dina(w_n633_6[1]),.dinb(w_G87_2[1]),.dout(n634),.clk(gclk));
	jnot g0563(.din(w_n634_0[1]),.dout(n635),.clk(gclk));
	jand g0564(.dina(w_dff_B_kt5ToKu03_0),.dinb(n631),.dout(n636),.clk(gclk));
	jand g0565(.dina(w_n626_0[1]),.dinb(w_n388_0[2]),.dout(n637),.clk(gclk));
	jand g0566(.dina(w_n637_0[1]),.dinb(w_n507_1[1]),.dout(n638),.clk(gclk));
	jand g0567(.dina(w_n638_7[1]),.dinb(w_G77_3[0]),.dout(n639),.clk(gclk));
	jand g0568(.dina(w_n628_0[0]),.dinb(w_n622_0[0]),.dout(n640),.clk(gclk));
	jand g0569(.dina(w_n640_7[1]),.dinb(w_G159_3[1]),.dout(n641),.clk(gclk));
	jor g0570(.dina(n641),.dinb(w_dff_B_gCWrTEup1_1),.dout(n642),.clk(gclk));
	jor g0571(.dina(n642),.dinb(w_G33_7[0]),.dout(n643),.clk(gclk));
	jnot g0572(.din(n643),.dout(n644),.clk(gclk));
	jand g0573(.dina(n644),.dinb(w_dff_B_X7YjN2rJ7_1),.dout(n645),.clk(gclk));
	jand g0574(.dina(w_n637_0[0]),.dinb(w_G190_1[2]),.dout(n646),.clk(gclk));
	jand g0575(.dina(w_n646_7[1]),.dinb(w_G58_4[0]),.dout(n647),.clk(gclk));
	jand g0576(.dina(w_n632_0[0]),.dinb(w_n507_1[0]),.dout(n648),.clk(gclk));
	jand g0577(.dina(w_n648_4[1]),.dinb(w_G107_3[0]),.dout(n649),.clk(gclk));
	jand g0578(.dina(w_n626_0[0]),.dinb(w_G200_1[0]),.dout(n650),.clk(gclk));
	jand g0579(.dina(w_n650_0[1]),.dinb(w_G190_1[1]),.dout(n651),.clk(gclk));
	jand g0580(.dina(w_n651_7[1]),.dinb(w_G50_4[1]),.dout(n652),.clk(gclk));
	jand g0581(.dina(w_n650_0[0]),.dinb(w_n507_0[2]),.dout(n653),.clk(gclk));
	jand g0582(.dina(w_n653_7[1]),.dinb(w_G68_3[2]),.dout(n654),.clk(gclk));
	jor g0583(.dina(n654),.dinb(n652),.dout(n655),.clk(gclk));
	jor g0584(.dina(n655),.dinb(w_n649_0[1]),.dout(n656),.clk(gclk));
	jor g0585(.dina(n656),.dinb(w_dff_B_PnhJcXFb8_1),.dout(n657),.clk(gclk));
	jnot g0586(.din(n657),.dout(n658),.clk(gclk));
	jand g0587(.dina(w_dff_B_myZ2XzXV4_0),.dinb(n645),.dout(n659),.clk(gclk));
	jnot g0588(.din(n659),.dout(n660),.clk(gclk));
	jand g0589(.dina(w_n646_7[0]),.dinb(w_G322_0[2]),.dout(n661),.clk(gclk));
	jand g0590(.dina(w_n633_6[0]),.dinb(w_G303_2[1]),.dout(n662),.clk(gclk));
	jand g0591(.dina(w_n629_5[0]),.dinb(w_G294_3[0]),.dout(n663),.clk(gclk));
	jor g0592(.dina(n663),.dinb(w_dff_B_yj2II1H15_1),.dout(n664),.clk(gclk));
	jand g0593(.dina(w_n651_7[0]),.dinb(w_G326_0[1]),.dout(n665),.clk(gclk));
	jor g0594(.dina(w_dff_B_4OPNyqaq3_0),.dinb(n664),.dout(n666),.clk(gclk));
	jand g0595(.dina(w_n640_7[0]),.dinb(w_dff_B_X2gvFluv2_1),.dout(n667),.clk(gclk));
	jor g0596(.dina(n667),.dinb(w_n153_5[0]),.dout(n668),.clk(gclk));
	jand g0597(.dina(w_n638_7[0]),.dinb(w_G311_1[2]),.dout(n669),.clk(gclk));
	jand g0598(.dina(w_n653_7[0]),.dinb(w_G317_1[1]),.dout(n670),.clk(gclk));
	jor g0599(.dina(n670),.dinb(n669),.dout(n671),.clk(gclk));
	jand g0600(.dina(w_n648_4[0]),.dinb(w_G283_3[1]),.dout(n672),.clk(gclk));
	jor g0601(.dina(w_dff_B_fjFwbOIT9_0),.dinb(n671),.dout(n673),.clk(gclk));
	jor g0602(.dina(n673),.dinb(n668),.dout(n674),.clk(gclk));
	jor g0603(.dina(n674),.dinb(n666),.dout(n675),.clk(gclk));
	jor g0604(.dina(n675),.dinb(w_dff_B_vPFDHvJh1_1),.dout(n676),.clk(gclk));
	jand g0605(.dina(w_dff_B_ICvUMYKM8_0),.dinb(n660),.dout(n677),.clk(gclk));
	jand g0606(.dina(w_n139_0[1]),.dinb(w_G169_1[0]),.dout(n678),.clk(gclk));
	jor g0607(.dina(n678),.dinb(w_n375_0[0]),.dout(n679),.clk(gclk));
	jnot g0608(.din(n679),.dout(n680),.clk(gclk));
	jor g0609(.dina(w_n680_4[1]),.dinb(n677),.dout(n681),.clk(gclk));
	jand g0610(.dina(w_n680_4[0]),.dinb(w_n620_0[1]),.dout(n682),.clk(gclk));
	jor g0611(.dina(w_n134_0[0]),.dinb(w_n352_1[0]),.dout(n683),.clk(gclk));
	jand g0612(.dina(w_n91_1[0]),.dinb(w_G33_6[2]),.dout(n684),.clk(gclk));
	jnot g0613(.din(w_n684_0[2]),.dout(n685),.clk(gclk));
	jand g0614(.dina(w_n118_0[0]),.dinb(w_n352_0[2]),.dout(n686),.clk(gclk));
	jor g0615(.dina(n686),.dinb(w_n685_0[1]),.dout(n687),.clk(gclk));
	jnot g0616(.din(n687),.dout(n688),.clk(gclk));
	jand g0617(.dina(n688),.dinb(w_dff_B_wHCIhoNy1_1),.dout(n689),.clk(gclk));
	jnot g0618(.din(w_n91_0[2]),.dout(n690),.clk(gclk));
	jand g0619(.dina(w_n690_1[1]),.dinb(w_n105_0[1]),.dout(n691),.clk(gclk));
	jand g0620(.dina(w_n91_0[1]),.dinb(w_n153_4[2]),.dout(n692),.clk(gclk));
	jand g0621(.dina(w_n692_0[1]),.dinb(w_G355_0),.dout(n693),.clk(gclk));
	jor g0622(.dina(n693),.dinb(n691),.dout(n694),.clk(gclk));
	jor g0623(.dina(w_dff_B_DDLmV1sL9_0),.dinb(n689),.dout(n695),.clk(gclk));
	jand g0624(.dina(n695),.dinb(w_n682_0[1]),.dout(n696),.clk(gclk));
	jnot g0625(.din(n696),.dout(n697),.clk(gclk));
	jand g0626(.dina(w_dff_B_kPQnTKnU7_0),.dinb(n681),.dout(n698),.clk(gclk));
	jand g0627(.dina(w_dff_B_gI3qsLLX6_0),.dinb(n621),.dout(n699),.clk(gclk));
	jand g0628(.dina(n699),.dinb(w_n614_5[0]),.dout(n700),.clk(gclk));
	jor g0629(.dina(n700),.dinb(w_dff_B_0I1CikA97_1),.dout(G396_fa_),.clk(gclk));
	jand g0630(.dina(w_n567_3[2]),.dinb(w_n383_0[0]),.dout(n702),.clk(gclk));
	jxor g0631(.dina(w_dff_B_mCIk2dZs8_0),.dinb(w_n394_0[0]),.dout(n703),.clk(gclk));
	jnot g0632(.din(w_n703_1[1]),.dout(n704),.clk(gclk));
	jand g0633(.dina(w_n704_0[1]),.dinb(w_n618_2[0]),.dout(n705),.clk(gclk));
	jnot g0634(.din(n705),.dout(n706),.clk(gclk));
	jand g0635(.dina(w_n653_6[2]),.dinb(w_G150_3[0]),.dout(n707),.clk(gclk));
	jand g0636(.dina(w_n651_6[2]),.dinb(w_G137_1[2]),.dout(n708),.clk(gclk));
	jand g0637(.dina(w_n633_5[2]),.dinb(w_G50_4[0]),.dout(n709),.clk(gclk));
	jor g0638(.dina(n709),.dinb(n708),.dout(n710),.clk(gclk));
	jand g0639(.dina(w_n646_6[2]),.dinb(w_G143_2[1]),.dout(n711),.clk(gclk));
	jor g0640(.dina(w_dff_B_AVdJ0gQA0_0),.dinb(n710),.dout(n712),.clk(gclk));
	jor g0641(.dina(n712),.dinb(w_dff_B_SFYn7sTX4_1),.dout(n713),.clk(gclk));
	jand g0642(.dina(w_n638_6[2]),.dinb(w_G159_3[0]),.dout(n714),.clk(gclk));
	jand g0643(.dina(w_n640_6[2]),.dinb(w_G132_1[1]),.dout(n715),.clk(gclk));
	jor g0644(.dina(n715),.dinb(w_dff_B_Ct5oodQI2_1),.dout(n716),.clk(gclk));
	jand g0645(.dina(w_n629_4[2]),.dinb(w_G58_3[2]),.dout(n717),.clk(gclk));
	jand g0646(.dina(w_n648_3[2]),.dinb(w_G68_3[1]),.dout(n718),.clk(gclk));
	jor g0647(.dina(w_n718_0[1]),.dinb(n717),.dout(n719),.clk(gclk));
	jor g0648(.dina(n719),.dinb(w_G33_6[1]),.dout(n720),.clk(gclk));
	jor g0649(.dina(n720),.dinb(w_dff_B_0km3CmbJ7_1),.dout(n721),.clk(gclk));
	jor g0650(.dina(n721),.dinb(w_dff_B_Ien3t5Ck6_1),.dout(n722),.clk(gclk));
	jand g0651(.dina(w_n653_6[1]),.dinb(w_G283_3[0]),.dout(n723),.clk(gclk));
	jand g0652(.dina(w_n640_6[1]),.dinb(w_G311_1[1]),.dout(n724),.clk(gclk));
	jor g0653(.dina(n724),.dinb(w_dff_B_rFZsDiXU3_1),.dout(n725),.clk(gclk));
	jand g0654(.dina(w_n633_5[1]),.dinb(w_G107_2[2]),.dout(n726),.clk(gclk));
	jor g0655(.dina(w_dff_B_hfXWDO4K3_0),.dinb(w_n630_0[0]),.dout(n727),.clk(gclk));
	jor g0656(.dina(n727),.dinb(n725),.dout(n728),.clk(gclk));
	jand g0657(.dina(w_n646_6[1]),.dinb(w_G294_2[2]),.dout(n729),.clk(gclk));
	jand g0658(.dina(w_n638_6[1]),.dinb(w_G116_4[0]),.dout(n730),.clk(gclk));
	jor g0659(.dina(n730),.dinb(n729),.dout(n731),.clk(gclk));
	jand g0660(.dina(w_n651_6[1]),.dinb(w_G303_2[0]),.dout(n732),.clk(gclk));
	jand g0661(.dina(w_n648_3[1]),.dinb(w_G87_2[0]),.dout(n733),.clk(gclk));
	jor g0662(.dina(w_n733_0[1]),.dinb(n732),.dout(n734),.clk(gclk));
	jor g0663(.dina(n734),.dinb(n731),.dout(n735),.clk(gclk));
	jor g0664(.dina(w_dff_B_5F7UX6Mj8_0),.dinb(n728),.dout(n736),.clk(gclk));
	jor g0665(.dina(n736),.dinb(w_n153_4[1]),.dout(n737),.clk(gclk));
	jand g0666(.dina(n737),.dinb(n722),.dout(n738),.clk(gclk));
	jor g0667(.dina(n738),.dinb(w_n680_3[2]),.dout(n739),.clk(gclk));
	jnot g0668(.din(w_n618_1[2]),.dout(n740),.clk(gclk));
	jand g0669(.dina(w_n680_3[1]),.dinb(w_dff_B_XYEEje5n4_1),.dout(n741),.clk(gclk));
	jand g0670(.dina(w_n741_1[1]),.dinb(w_n72_0[1]),.dout(n742),.clk(gclk));
	jnot g0671(.din(n742),.dout(n743),.clk(gclk));
	jand g0672(.dina(w_dff_B_GFUvPOFf8_0),.dinb(n739),.dout(n744),.clk(gclk));
	jand g0673(.dina(n744),.dinb(w_n614_4[2]),.dout(n745),.clk(gclk));
	jand g0674(.dina(w_dff_B_UN52YtQS4_0),.dinb(n706),.dout(n746),.clk(gclk));
	jnot g0675(.din(n746),.dout(n747),.clk(gclk));
	jor g0676(.dina(w_n584_0[0]),.dinb(w_n395_0[0]),.dout(n748),.clk(gclk));
	jand g0677(.dina(w_n350_0[0]),.dinb(w_n570_0[0]),.dout(n749),.clk(gclk));
	jand g0678(.dina(w_n349_0[0]),.dinb(w_n520_0[0]),.dout(n750),.clk(gclk));
	jnot g0679(.din(w_n548_0[0]),.dout(n751),.clk(gclk));
	jor g0680(.dina(w_dff_B_b6ipeSB23_0),.dinb(n750),.dout(n752),.clk(gclk));
	jor g0681(.dina(n752),.dinb(n749),.dout(n753),.clk(gclk));
	jand g0682(.dina(w_n571_1[1]),.dinb(n753),.dout(n754),.clk(gclk));
	jor g0683(.dina(w_n703_1[0]),.dinb(w_n754_0[1]),.dout(n755),.clk(gclk));
	jand g0684(.dina(n755),.dinb(w_n748_0[1]),.dout(n756),.clk(gclk));
	jxor g0685(.dina(n756),.dinb(w_n600_1[1]),.dout(n757),.clk(gclk));
	jor g0686(.dina(n757),.dinb(w_n614_4[1]),.dout(n758),.clk(gclk));
	jand g0687(.dina(n758),.dinb(w_dff_B_VnAYDJq25_1),.dout(n759),.clk(gclk));
	jnot g0688(.din(w_n759_0[1]),.dout(G384_fa_),.clk(gclk));
	jnot g0689(.din(w_n90_0[1]),.dout(n761),.clk(gclk));
	jand g0690(.dina(w_n112_0[0]),.dinb(n761),.dout(n762),.clk(gclk));
	jnot g0691(.din(w_n566_1[0]),.dout(n763),.clk(gclk));
	jand g0692(.dina(w_dff_B_QanFgOYD7_0),.dinb(w_n503_0[0]),.dout(n764),.clk(gclk));
	jand g0693(.dina(w_n566_0[2]),.dinb(w_n500_0[0]),.dout(n765),.clk(gclk));
	jxor g0694(.dina(w_dff_B_Y3vRi9GH1_0),.dinb(w_n511_0[0]),.dout(n766),.clk(gclk));
	jnot g0695(.din(w_n766_0[1]),.dout(n767),.clk(gclk));
	jor g0696(.dina(w_n567_3[1]),.dinb(w_n559_0[0]),.dout(n768),.clk(gclk));
	jnot g0697(.din(n768),.dout(n769),.clk(gclk));
	jand g0698(.dina(w_n567_3[0]),.dinb(w_n417_0[0]),.dout(n770),.clk(gclk));
	jxor g0699(.dina(w_dff_B_toa3xpjP1_0),.dinb(w_n426_0[0]),.dout(n771),.clk(gclk));
	jnot g0700(.din(w_n771_1[1]),.dout(n772),.clk(gclk));
	jand g0701(.dina(w_n772_0[1]),.dinb(w_n703_0[2]),.dout(n773),.clk(gclk));
	jand g0702(.dina(w_n773_0[1]),.dinb(w_n754_0[0]),.dout(n774),.clk(gclk));
	jor g0703(.dina(n774),.dinb(w_dff_B_6lVSt8ed3_1),.dout(n775),.clk(gclk));
	jand g0704(.dina(w_n775_0[1]),.dinb(w_n767_1[1]),.dout(n776),.clk(gclk));
	jor g0705(.dina(n776),.dinb(w_dff_B_7Cxjwifc4_1),.dout(n777),.clk(gclk));
	jand g0706(.dina(w_n773_0[0]),.dinb(w_n767_1[0]),.dout(n778),.clk(gclk));
	jxor g0707(.dina(n778),.dinb(w_n514_0[2]),.dout(n779),.clk(gclk));
	jor g0708(.dina(n779),.dinb(w_n600_1[0]),.dout(n780),.clk(gclk));
	jor g0709(.dina(w_n567_2[2]),.dinb(w_n551_0[0]),.dout(n781),.clk(gclk));
	jand g0710(.dina(n781),.dinb(w_n562_0[0]),.dout(n782),.clk(gclk));
	jxor g0711(.dina(w_n782_0[1]),.dinb(n780),.dout(n783),.clk(gclk));
	jxor g0712(.dina(w_dff_B_L1sWVBgv2_0),.dinb(w_n777_0[1]),.dout(n784),.clk(gclk));
	jand g0713(.dina(n784),.dinb(w_dff_B_XEYBo1O55_1),.dout(n785),.clk(gclk));
	jor g0714(.dina(w_n75_1[0]),.dinb(w_n74_1[0]),.dout(n786),.clk(gclk));
	jand g0715(.dina(n786),.dinb(w_G77_2[2]),.dout(n787),.clk(gclk));
	jor g0716(.dina(n787),.dinb(w_n73_1[1]),.dout(n788),.clk(gclk));
	jand g0717(.dina(w_G58_3[1]),.dinb(w_G50_3[2]),.dout(n789),.clk(gclk));
	jor g0718(.dina(n789),.dinb(w_G68_3[0]),.dout(n790),.clk(gclk));
	jand g0719(.dina(n790),.dinb(w_n90_0[0]),.dout(n791),.clk(gclk));
	jand g0720(.dina(w_dff_B_1OBZCMhy3_0),.dinb(n788),.dout(n792),.clk(gclk));
	jand g0721(.dina(w_n312_0[0]),.dinb(w_n120_0[0]),.dout(n793),.clk(gclk));
	jand g0722(.dina(n793),.dinb(w_G116_3[2]),.dout(n794),.clk(gclk));
	jor g0723(.dina(w_dff_B_YjUwNIFM7_0),.dinb(n792),.dout(n795),.clk(gclk));
	jor g0724(.dina(w_dff_B_tv2ZYgBB6_0),.dinb(n785),.dout(w_dff_A_tne6B1924_2),.clk(gclk));
	jand g0725(.dina(w_n567_2[1]),.dinb(w_n292_0[0]),.dout(n797),.clk(gclk));
	jxor g0726(.dina(w_dff_B_8GrNoiK39_0),.dinb(w_n534_0[0]),.dout(n798),.clk(gclk));
	jand g0727(.dina(w_n798_0[1]),.dinb(w_n619_0[1]),.dout(n799),.clk(gclk));
	jnot g0728(.din(n799),.dout(n800),.clk(gclk));
	jand g0729(.dina(w_n684_0[1]),.dinb(w_n126_0[0]),.dout(n801),.clk(gclk));
	jnot g0730(.din(w_n682_0[0]),.dout(n802),.clk(gclk));
	jand g0731(.dina(w_n690_1[0]),.dinb(w_G87_1[2]),.dout(n803),.clk(gclk));
	jor g0732(.dina(w_dff_B_Fxsrb80G4_0),.dinb(w_n802_0[2]),.dout(n804),.clk(gclk));
	jor g0733(.dina(n804),.dinb(w_dff_B_2ANOq5n72_1),.dout(n805),.clk(gclk));
	jand g0734(.dina(n805),.dinb(w_n614_4[0]),.dout(n806),.clk(gclk));
	jand g0735(.dina(w_n646_6[0]),.dinb(w_G303_1[2]),.dout(n807),.clk(gclk));
	jand g0736(.dina(w_n638_6[0]),.dinb(w_G283_2[2]),.dout(n808),.clk(gclk));
	jor g0737(.dina(n808),.dinb(n807),.dout(n809),.clk(gclk));
	jand g0738(.dina(w_n651_6[0]),.dinb(w_G311_1[0]),.dout(n810),.clk(gclk));
	jand g0739(.dina(w_n633_5[0]),.dinb(w_G116_3[1]),.dout(n811),.clk(gclk));
	jor g0740(.dina(n811),.dinb(n810),.dout(n812),.clk(gclk));
	jand g0741(.dina(w_n653_6[0]),.dinb(w_G294_2[1]),.dout(n813),.clk(gclk));
	jand g0742(.dina(w_n640_6[0]),.dinb(w_G317_1[0]),.dout(n814),.clk(gclk));
	jor g0743(.dina(n814),.dinb(w_dff_B_T5V9d2Bh4_1),.dout(n815),.clk(gclk));
	jand g0744(.dina(w_n629_4[1]),.dinb(w_G107_2[1]),.dout(n816),.clk(gclk));
	jand g0745(.dina(w_n648_3[0]),.dinb(w_G97_2[2]),.dout(n817),.clk(gclk));
	jor g0746(.dina(w_n817_0[1]),.dinb(n816),.dout(n818),.clk(gclk));
	jor g0747(.dina(n818),.dinb(n815),.dout(n819),.clk(gclk));
	jor g0748(.dina(n819),.dinb(w_dff_B_1IAQThCU0_1),.dout(n820),.clk(gclk));
	jor g0749(.dina(n820),.dinb(w_dff_B_tmSYz4yx9_1),.dout(n821),.clk(gclk));
	jand g0750(.dina(n821),.dinb(w_G33_6[0]),.dout(n822),.clk(gclk));
	jand g0751(.dina(w_n638_5[2]),.dinb(w_G50_3[1]),.dout(n823),.clk(gclk));
	jand g0752(.dina(w_n640_5[2]),.dinb(w_G137_1[1]),.dout(n824),.clk(gclk));
	jor g0753(.dina(n824),.dinb(w_dff_B_BdpCwJC28_1),.dout(n825),.clk(gclk));
	jand g0754(.dina(w_n651_5[2]),.dinb(w_G143_2[0]),.dout(n826),.clk(gclk));
	jand g0755(.dina(w_n653_5[2]),.dinb(w_G159_2[2]),.dout(n827),.clk(gclk));
	jor g0756(.dina(n827),.dinb(n826),.dout(n828),.clk(gclk));
	jand g0757(.dina(w_n633_4[2]),.dinb(w_G58_3[0]),.dout(n829),.clk(gclk));
	jand g0758(.dina(w_n629_4[0]),.dinb(w_G68_2[2]),.dout(n830),.clk(gclk));
	jor g0759(.dina(w_n830_0[1]),.dinb(w_dff_B_YSJ6bEhz9_1),.dout(n831),.clk(gclk));
	jand g0760(.dina(w_n646_5[2]),.dinb(w_G150_2[2]),.dout(n832),.clk(gclk));
	jand g0761(.dina(w_n648_2[2]),.dinb(w_G77_2[1]),.dout(n833),.clk(gclk));
	jor g0762(.dina(w_n833_0[1]),.dinb(n832),.dout(n834),.clk(gclk));
	jor g0763(.dina(w_dff_B_VQ8gnLiz2_0),.dinb(n831),.dout(n835),.clk(gclk));
	jor g0764(.dina(n835),.dinb(w_dff_B_RQ0tSwua1_1),.dout(n836),.clk(gclk));
	jor g0765(.dina(n836),.dinb(w_dff_B_1bIJ8zSE5_1),.dout(n837),.clk(gclk));
	jand g0766(.dina(n837),.dinb(w_n153_4[0]),.dout(n838),.clk(gclk));
	jor g0767(.dina(n838),.dinb(n822),.dout(n839),.clk(gclk));
	jor g0768(.dina(n839),.dinb(w_n680_3[0]),.dout(n840),.clk(gclk));
	jand g0769(.dina(n840),.dinb(w_dff_B_zT8eHC0d9_1),.dout(n841),.clk(gclk));
	jand g0770(.dina(w_dff_B_XjXOnsmf3_0),.dinb(n800),.dout(n842),.clk(gclk));
	jnot g0771(.din(n842),.dout(n843),.clk(gclk));
	jand g0772(.dina(w_n567_2[0]),.dinb(w_n323_0[0]),.dout(n844),.clk(gclk));
	jxor g0773(.dina(w_dff_B_Uf0XxWAg0_0),.dinb(w_n542_0[0]),.dout(n845),.clk(gclk));
	jnot g0774(.din(w_n845_0[2]),.dout(n846),.clk(gclk));
	jand g0775(.dina(w_dff_B_FDvsbCPd3_0),.dinb(w_n580_0[1]),.dout(n847),.clk(gclk));
	jand g0776(.dina(w_n571_1[0]),.dinb(w_n541_0[0]),.dout(n848),.clk(gclk));
	jand g0777(.dina(w_n579_1[0]),.dinb(w_n348_0[0]),.dout(n849),.clk(gclk));
	jand g0778(.dina(n849),.dinb(w_n572_0[1]),.dout(n850),.clk(gclk));
	jand g0779(.dina(w_n569_0[0]),.dinb(w_n333_0[0]),.dout(n851),.clk(gclk));
	jor g0780(.dina(w_dff_B_7fAGyRMk1_0),.dinb(n850),.dout(n852),.clk(gclk));
	jor g0781(.dina(n852),.dinb(w_dff_B_VjYy4XQB0_1),.dout(n853),.clk(gclk));
	jxor g0782(.dina(n853),.dinb(w_n798_0[0]),.dout(n854),.clk(gclk));
	jxor g0783(.dina(n854),.dinb(w_dff_B_orJoUx8x2_1),.dout(n855),.clk(gclk));
	jor g0784(.dina(w_n855_0[1]),.dinb(w_n613_1[1]),.dout(n856),.clk(gclk));
	jnot g0785(.din(w_n573_0[0]),.dout(n857),.clk(gclk));
	jor g0786(.dina(w_n579_0[2]),.dinb(w_n572_0[0]),.dout(n858),.clk(gclk));
	jand g0787(.dina(w_dff_B_vHNzx2Rh3_0),.dinb(n857),.dout(n859),.clk(gclk));
	jxor g0788(.dina(n859),.dinb(w_n577_0[0]),.dout(n860),.clk(gclk));
	jnot g0789(.din(w_n860_0[1]),.dout(n861),.clk(gclk));
	jxor g0790(.dina(w_n580_0[0]),.dinb(w_n574_0[0]),.dout(n862),.clk(gclk));
	jxor g0791(.dina(n862),.dinb(w_n845_0[1]),.dout(n863),.clk(gclk));
	jor g0792(.dina(w_n863_0[2]),.dinb(w_n861_0[1]),.dout(n864),.clk(gclk));
	jand g0793(.dina(n864),.dinb(w_n601_0[1]),.dout(n865),.clk(gclk));
	jor g0794(.dina(w_n855_0[0]),.dinb(w_n604_2[0]),.dout(n866),.clk(gclk));
	jor g0795(.dina(w_dff_B_ySXOopji0_0),.dinb(n865),.dout(n867),.clk(gclk));
	jand g0796(.dina(n867),.dinb(w_dff_B_a7sBk9jl0_1),.dout(n868),.clk(gclk));
	jand g0797(.dina(n868),.dinb(w_dff_B_wmhtPQGZ2_1),.dout(n869),.clk(gclk));
	jnot g0798(.din(w_n869_0[2]),.dout(w_dff_A_vfRDkQlW9_1),.clk(gclk));
	jor g0799(.dina(w_n602_0[0]),.dinb(w_n604_1[2]),.dout(n871),.clk(gclk));
	jand g0800(.dina(n871),.dinb(w_n861_0[0]),.dout(n872),.clk(gclk));
	jand g0801(.dina(w_n860_0[0]),.dinb(w_n601_0[0]),.dout(n873),.clk(gclk));
	jand g0802(.dina(w_n873_0[1]),.dinb(w_n613_1[0]),.dout(n874),.clk(gclk));
	jor g0803(.dina(n874),.dinb(w_n614_3[2]),.dout(n875),.clk(gclk));
	jor g0804(.dina(w_n875_0[1]),.dinb(n872),.dout(n876),.clk(gclk));
	jor g0805(.dina(w_n620_0[0]),.dinb(w_n579_0[1]),.dout(n877),.clk(gclk));
	jand g0806(.dina(w_n653_5[1]),.dinb(w_G58_2[2]),.dout(n878),.clk(gclk));
	jand g0807(.dina(w_n638_5[1]),.dinb(w_G68_2[1]),.dout(n879),.clk(gclk));
	jor g0808(.dina(n879),.dinb(w_n817_0[0]),.dout(n880),.clk(gclk));
	jor g0809(.dina(n880),.dinb(w_G33_5[2]),.dout(n881),.clk(gclk));
	jor g0810(.dina(n881),.dinb(w_dff_B_qO6l6Hji1_1),.dout(n882),.clk(gclk));
	jnot g0811(.din(n882),.dout(n883),.clk(gclk));
	jand g0812(.dina(w_n629_3[2]),.dinb(w_G87_1[1]),.dout(n884),.clk(gclk));
	jnot g0813(.din(w_n884_0[1]),.dout(n885),.clk(gclk));
	jand g0814(.dina(w_n633_4[1]),.dinb(w_G77_2[0]),.dout(n886),.clk(gclk));
	jnot g0815(.din(n886),.dout(n887),.clk(gclk));
	jand g0816(.dina(w_n887_0[1]),.dinb(n885),.dout(n888),.clk(gclk));
	jand g0817(.dina(w_n646_5[1]),.dinb(w_G50_3[0]),.dout(n889),.clk(gclk));
	jand g0818(.dina(w_n640_5[1]),.dinb(w_G150_2[1]),.dout(n890),.clk(gclk));
	jor g0819(.dina(n890),.dinb(w_dff_B_HALy3Khn7_1),.dout(n891),.clk(gclk));
	jand g0820(.dina(w_n651_5[1]),.dinb(w_G159_2[1]),.dout(n892),.clk(gclk));
	jor g0821(.dina(w_dff_B_7bU8Sqr96_0),.dinb(n891),.dout(n893),.clk(gclk));
	jnot g0822(.din(n893),.dout(n894),.clk(gclk));
	jand g0823(.dina(n894),.dinb(w_dff_B_DDUoAJAO2_1),.dout(n895),.clk(gclk));
	jand g0824(.dina(n895),.dinb(w_dff_B_9z8F1Thl9_1),.dout(n896),.clk(gclk));
	jnot g0825(.din(n896),.dout(n897),.clk(gclk));
	jand g0826(.dina(w_n653_5[0]),.dinb(w_G311_0[2]),.dout(n898),.clk(gclk));
	jand g0827(.dina(w_n633_4[0]),.dinb(w_G294_2[0]),.dout(n899),.clk(gclk));
	jand g0828(.dina(w_n629_3[1]),.dinb(w_G283_2[1]),.dout(n900),.clk(gclk));
	jor g0829(.dina(n900),.dinb(w_dff_B_RSXJqNCL9_1),.dout(n901),.clk(gclk));
	jand g0830(.dina(w_n651_5[0]),.dinb(w_G322_0[1]),.dout(n902),.clk(gclk));
	jand g0831(.dina(w_n640_5[0]),.dinb(w_G326_0[0]),.dout(n903),.clk(gclk));
	jor g0832(.dina(n903),.dinb(w_dff_B_VPxtV2Dm3_1),.dout(n904),.clk(gclk));
	jor g0833(.dina(n904),.dinb(n901),.dout(n905),.clk(gclk));
	jand g0834(.dina(w_n638_5[0]),.dinb(w_G303_1[1]),.dout(n906),.clk(gclk));
	jand g0835(.dina(w_n648_2[1]),.dinb(w_G116_3[0]),.dout(n907),.clk(gclk));
	jor g0836(.dina(n907),.dinb(n906),.dout(n908),.clk(gclk));
	jand g0837(.dina(w_n646_5[0]),.dinb(w_G317_0[2]),.dout(n909),.clk(gclk));
	jor g0838(.dina(w_dff_B_5iePj3C97_0),.dinb(n908),.dout(n910),.clk(gclk));
	jor g0839(.dina(n910),.dinb(w_n153_3[2]),.dout(n911),.clk(gclk));
	jor g0840(.dina(n911),.dinb(n905),.dout(n912),.clk(gclk));
	jor g0841(.dina(n912),.dinb(w_dff_B_hVb0CsHc0_1),.dout(n913),.clk(gclk));
	jand g0842(.dina(w_dff_B_Lc4vOZKj4_0),.dinb(n897),.dout(n914),.clk(gclk));
	jor g0843(.dina(n914),.dinb(w_n680_2[2]),.dout(n915),.clk(gclk));
	jand g0844(.dina(w_n690_0[2]),.dinb(w_n81_0[2]),.dout(n916),.clk(gclk));
	jnot g0845(.din(n916),.dout(n917),.clk(gclk));
	jnot g0846(.din(w_n605_0[1]),.dout(n918),.clk(gclk));
	jand g0847(.dina(w_n692_0[0]),.dinb(n918),.dout(n919),.clk(gclk));
	jnot g0848(.din(n919),.dout(n920),.clk(gclk));
	jand g0849(.dina(w_n130_0[0]),.dinb(w_G45_0[1]),.dout(n921),.clk(gclk));
	jor g0850(.dina(w_dff_B_f9OO8QL00_0),.dinb(w_n685_0[0]),.dout(n922),.clk(gclk));
	jand g0851(.dina(w_dff_B_Ln9ZbyCK9_0),.dinb(n920),.dout(n923),.clk(gclk));
	jand g0852(.dina(w_G77_1[2]),.dinb(w_G68_2[0]),.dout(n924),.clk(gclk));
	jnot g0853(.din(n924),.dout(n925),.clk(gclk));
	jand g0854(.dina(w_G58_2[1]),.dinb(w_n73_1[0]),.dout(n926),.clk(gclk));
	jand g0855(.dina(n926),.dinb(n925),.dout(n927),.clk(gclk));
	jand g0856(.dina(w_dff_B_3E0Ul3YV3_0),.dinb(w_n605_0[0]),.dout(n928),.clk(gclk));
	jand g0857(.dina(n928),.dinb(w_n352_0[1]),.dout(n929),.clk(gclk));
	jor g0858(.dina(w_dff_B_qpxD3fEa0_0),.dinb(n923),.dout(n930),.clk(gclk));
	jand g0859(.dina(n930),.dinb(w_dff_B_VkhJlcVA1_1),.dout(n931),.clk(gclk));
	jor g0860(.dina(n931),.dinb(w_n802_0[1]),.dout(n932),.clk(gclk));
	jand g0861(.dina(w_dff_B_lRcnW8Hx2_0),.dinb(n915),.dout(n933),.clk(gclk));
	jand g0862(.dina(n933),.dinb(n877),.dout(n934),.clk(gclk));
	jand g0863(.dina(n934),.dinb(w_n614_3[1]),.dout(n935),.clk(gclk));
	jnot g0864(.din(n935),.dout(n936),.clk(gclk));
	jand g0865(.dina(w_dff_B_kBTgxbTc6_0),.dinb(n876),.dout(n937),.clk(gclk));
	jnot g0866(.din(w_n937_0[2]),.dout(w_dff_A_ywVOaL5R9_1),.clk(gclk));
	jnot g0867(.din(w_n863_0[1]),.dout(n939),.clk(gclk));
	jnot g0868(.din(w_n873_0[0]),.dout(n940),.clk(gclk));
	jor g0869(.dina(n940),.dinb(w_dff_B_pL18KfnZ3_1),.dout(n941),.clk(gclk));
	jor g0870(.dina(n941),.dinb(w_n604_1[1]),.dout(n942),.clk(gclk));
	jor g0871(.dina(w_n875_0[0]),.dinb(w_n863_0[0]),.dout(n943),.clk(gclk));
	jand g0872(.dina(w_n845_0[0]),.dinb(w_n619_0[0]),.dout(n944),.clk(gclk));
	jnot g0873(.din(n944),.dout(n945),.clk(gclk));
	jand g0874(.dina(w_n690_0[1]),.dinb(w_G97_2[1]),.dout(n946),.clk(gclk));
	jand g0875(.dina(w_n684_0[0]),.dinb(w_n137_0[0]),.dout(n947),.clk(gclk));
	jor g0876(.dina(w_dff_B_qayTBsAn8_0),.dinb(w_n802_0[0]),.dout(n948),.clk(gclk));
	jor g0877(.dina(n948),.dinb(w_dff_B_Fk6489C09_1),.dout(n949),.clk(gclk));
	jand g0878(.dina(w_n653_4[2]),.dinb(w_G50_2[2]),.dout(n950),.clk(gclk));
	jand g0879(.dina(w_n638_4[2]),.dinb(w_G58_2[0]),.dout(n951),.clk(gclk));
	jor g0880(.dina(n951),.dinb(n950),.dout(n952),.clk(gclk));
	jand g0881(.dina(w_n646_4[2]),.dinb(w_G159_2[0]),.dout(n953),.clk(gclk));
	jand g0882(.dina(w_n633_3[2]),.dinb(w_G68_1[2]),.dout(n954),.clk(gclk));
	jor g0883(.dina(n954),.dinb(n953),.dout(n955),.clk(gclk));
	jand g0884(.dina(w_n651_4[2]),.dinb(w_G150_2[0]),.dout(n956),.clk(gclk));
	jor g0885(.dina(n956),.dinb(w_n733_0[0]),.dout(n957),.clk(gclk));
	jand g0886(.dina(w_n640_4[2]),.dinb(w_G143_1[2]),.dout(n958),.clk(gclk));
	jand g0887(.dina(w_n629_3[0]),.dinb(w_G77_1[1]),.dout(n959),.clk(gclk));
	jor g0888(.dina(w_n959_0[1]),.dinb(n958),.dout(n960),.clk(gclk));
	jor g0889(.dina(n960),.dinb(w_dff_B_hdG0pbbR9_1),.dout(n961),.clk(gclk));
	jor g0890(.dina(n961),.dinb(w_dff_B_cnDPdZq33_1),.dout(n962),.clk(gclk));
	jor g0891(.dina(n962),.dinb(w_dff_B_r8bLlVZ74_1),.dout(n963),.clk(gclk));
	jand g0892(.dina(n963),.dinb(w_n153_3[1]),.dout(n964),.clk(gclk));
	jand g0893(.dina(w_n638_4[1]),.dinb(w_G294_1[2]),.dout(n965),.clk(gclk));
	jand g0894(.dina(w_n640_4[1]),.dinb(w_G322_0[0]),.dout(n966),.clk(gclk));
	jor g0895(.dina(n966),.dinb(w_dff_B_xNg1sUQ42_1),.dout(n967),.clk(gclk));
	jand g0896(.dina(w_n646_4[1]),.dinb(w_G311_0[1]),.dout(n968),.clk(gclk));
	jand g0897(.dina(w_n651_4[1]),.dinb(w_G317_0[1]),.dout(n969),.clk(gclk));
	jor g0898(.dina(n969),.dinb(n968),.dout(n970),.clk(gclk));
	jand g0899(.dina(w_n653_4[1]),.dinb(w_G303_1[0]),.dout(n971),.clk(gclk));
	jor g0900(.dina(n971),.dinb(w_n649_0[0]),.dout(n972),.clk(gclk));
	jor g0901(.dina(n972),.dinb(n970),.dout(n973),.clk(gclk));
	jand g0902(.dina(w_n633_3[1]),.dinb(w_G283_2[0]),.dout(n974),.clk(gclk));
	jand g0903(.dina(w_n629_2[2]),.dinb(w_G116_2[2]),.dout(n975),.clk(gclk));
	jor g0904(.dina(n975),.dinb(w_dff_B_SLq0e8Kd6_1),.dout(n976),.clk(gclk));
	jor g0905(.dina(n976),.dinb(n973),.dout(n977),.clk(gclk));
	jor g0906(.dina(n977),.dinb(w_dff_B_FWJMrzgD2_1),.dout(n978),.clk(gclk));
	jand g0907(.dina(n978),.dinb(w_G33_5[1]),.dout(n979),.clk(gclk));
	jor g0908(.dina(n979),.dinb(w_n680_2[1]),.dout(n980),.clk(gclk));
	jor g0909(.dina(n980),.dinb(n964),.dout(n981),.clk(gclk));
	jand g0910(.dina(n981),.dinb(w_n614_3[0]),.dout(n982),.clk(gclk));
	jand g0911(.dina(n982),.dinb(w_dff_B_mhOjddX57_1),.dout(n983),.clk(gclk));
	jand g0912(.dina(w_dff_B_x2J2RxHQ3_0),.dinb(n945),.dout(n984),.clk(gclk));
	jnot g0913(.din(n984),.dout(n985),.clk(gclk));
	jand g0914(.dina(w_dff_B_dBM934nq7_0),.dinb(n943),.dout(n986),.clk(gclk));
	jand g0915(.dina(n986),.dinb(w_dff_B_7nl7DOtC1_1),.dout(n987),.clk(gclk));
	jnot g0916(.din(w_n987_0[2]),.dout(w_dff_A_Ezxpsepx8_1),.clk(gclk));
	jand g0917(.dina(w_n766_0[0]),.dinb(w_n618_1[1]),.dout(n989),.clk(gclk));
	jnot g0918(.din(n989),.dout(n990),.clk(gclk));
	jand g0919(.dina(w_n651_4[0]),.dinb(w_G128_0[2]),.dout(n991),.clk(gclk));
	jand g0920(.dina(w_n640_4[0]),.dinb(w_G125_0[1]),.dout(n992),.clk(gclk));
	jor g0921(.dina(n992),.dinb(w_dff_B_Ijayki2N9_1),.dout(n993),.clk(gclk));
	jand g0922(.dina(w_n648_2[0]),.dinb(w_G50_2[1]),.dout(n994),.clk(gclk));
	jand g0923(.dina(w_n653_4[0]),.dinb(w_G137_1[0]),.dout(n995),.clk(gclk));
	jor g0924(.dina(n995),.dinb(n994),.dout(n996),.clk(gclk));
	jor g0925(.dina(n996),.dinb(w_G33_5[0]),.dout(n997),.clk(gclk));
	jor g0926(.dina(n997),.dinb(n993),.dout(n998),.clk(gclk));
	jand g0927(.dina(w_n638_4[0]),.dinb(w_G143_1[1]),.dout(n999),.clk(gclk));
	jand g0928(.dina(w_n633_3[0]),.dinb(w_G150_1[2]),.dout(n1000),.clk(gclk));
	jand g0929(.dina(w_n629_2[1]),.dinb(w_G159_1[2]),.dout(n1001),.clk(gclk));
	jand g0930(.dina(w_n646_4[0]),.dinb(w_G132_1[0]),.dout(n1002),.clk(gclk));
	jor g0931(.dina(w_dff_B_ZSMIrfLb0_0),.dinb(n1001),.dout(n1003),.clk(gclk));
	jor g0932(.dina(n1003),.dinb(w_dff_B_3LiZdvJa5_1),.dout(n1004),.clk(gclk));
	jor g0933(.dina(n1004),.dinb(w_dff_B_dv2uFe8e2_1),.dout(n1005),.clk(gclk));
	jor g0934(.dina(n1005),.dinb(w_dff_B_wzqu9s0k8_1),.dout(n1006),.clk(gclk));
	jand g0935(.dina(w_n651_3[2]),.dinb(w_G283_1[2]),.dout(n1007),.clk(gclk));
	jand g0936(.dina(w_n638_3[2]),.dinb(w_G97_2[0]),.dout(n1008),.clk(gclk));
	jor g0937(.dina(n1008),.dinb(w_n153_3[0]),.dout(n1009),.clk(gclk));
	jor g0938(.dina(n1009),.dinb(w_dff_B_zxYraqje1_1),.dout(n1010),.clk(gclk));
	jand g0939(.dina(w_n646_3[2]),.dinb(w_G116_2[1]),.dout(n1011),.clk(gclk));
	jand g0940(.dina(w_n640_3[2]),.dinb(w_G294_1[1]),.dout(n1012),.clk(gclk));
	jor g0941(.dina(n1012),.dinb(w_dff_B_fYOfFF587_1),.dout(n1013),.clk(gclk));
	jand g0942(.dina(w_n653_3[2]),.dinb(w_G107_2[0]),.dout(n1014),.clk(gclk));
	jor g0943(.dina(n1014),.dinb(w_n634_0[0]),.dout(n1015),.clk(gclk));
	jor g0944(.dina(w_dff_B_Gl0g4FKD0_0),.dinb(n1013),.dout(n1016),.clk(gclk));
	jor g0945(.dina(n1016),.dinb(w_dff_B_XudOkgBB5_1),.dout(n1017),.clk(gclk));
	jor g0946(.dina(n1017),.dinb(w_n959_0[0]),.dout(n1018),.clk(gclk));
	jor g0947(.dina(n1018),.dinb(w_n718_0[0]),.dout(n1019),.clk(gclk));
	jand g0948(.dina(n1019),.dinb(w_dff_B_mgULKXz23_1),.dout(n1020),.clk(gclk));
	jor g0949(.dina(n1020),.dinb(w_n680_2[0]),.dout(n1021),.clk(gclk));
	jand g0950(.dina(w_n741_1[0]),.dinb(w_n74_0[2]),.dout(n1022),.clk(gclk));
	jnot g0951(.din(n1022),.dout(n1023),.clk(gclk));
	jand g0952(.dina(w_dff_B_sjjFa77P5_0),.dinb(n1021),.dout(n1024),.clk(gclk));
	jand g0953(.dina(n1024),.dinb(w_n614_2[2]),.dout(n1025),.clk(gclk));
	jand g0954(.dina(w_dff_B_4I3jzZeY7_0),.dinb(n990),.dout(n1026),.clk(gclk));
	jnot g0955(.din(n1026),.dout(n1027),.clk(gclk));
	jor g0956(.dina(w_n600_0[2]),.dinb(w_n514_0[1]),.dout(n1028),.clk(gclk));
	jand g0957(.dina(w_dff_B_ukbYK3mL7_0),.dinb(w_n782_0[0]),.dout(n1029),.clk(gclk));
	jnot g0958(.din(w_n387_0[0]),.dout(n1030),.clk(gclk));
	jand g0959(.dina(w_n571_0[2]),.dinb(n1030),.dout(n1031),.clk(gclk));
	jnot g0960(.din(n1031),.dout(n1032),.clk(gclk));
	jand g0961(.dina(w_dff_B_5q9U8p1K7_0),.dinb(w_n748_0[0]),.dout(n1033),.clk(gclk));
	jor g0962(.dina(w_n567_1[2]),.dinb(w_n351_0[0]),.dout(n1034),.clk(gclk));
	jand g0963(.dina(w_n598_0[0]),.dinb(n1034),.dout(n1035),.clk(gclk));
	jand g0964(.dina(w_n703_0[1]),.dinb(n1035),.dout(n1036),.clk(gclk));
	jxor g0965(.dina(w_n1036_0[1]),.dinb(w_n771_1[0]),.dout(n1037),.clk(gclk));
	jxor g0966(.dina(n1037),.dinb(w_n1033_0[1]),.dout(n1038),.clk(gclk));
	jand g0967(.dina(n1038),.dinb(w_n1029_0[2]),.dout(n1039),.clk(gclk));
	jor g0968(.dina(w_n1039_0[1]),.dinb(w_n604_1[0]),.dout(n1040),.clk(gclk));
	jand g0969(.dina(w_n1040_0[1]),.dinb(w_n613_0[2]),.dout(n1041),.clk(gclk));
	jor g0970(.dina(w_n704_0[0]),.dinb(w_n600_0[1]),.dout(n1042),.clk(gclk));
	jor g0971(.dina(n1042),.dinb(w_n771_0[2]),.dout(n1043),.clk(gclk));
	jxor g0972(.dina(w_n775_0[0]),.dinb(w_n767_0[2]),.dout(n1044),.clk(gclk));
	jxor g0973(.dina(w_n1044_0[1]),.dinb(w_n1043_0[1]),.dout(n1045),.clk(gclk));
	jor g0974(.dina(w_n1045_0[1]),.dinb(w_n1041_0[1]),.dout(n1046),.clk(gclk));
	jnot g0975(.din(w_n1039_0[0]),.dout(n1047),.clk(gclk));
	jnot g0976(.din(w_n1043_0[0]),.dout(n1048),.clk(gclk));
	jxor g0977(.dina(w_n1044_0[0]),.dinb(w_n1048_0[1]),.dout(n1049),.clk(gclk));
	jor g0978(.dina(n1049),.dinb(w_n604_0[2]),.dout(n1050),.clk(gclk));
	jor g0979(.dina(n1050),.dinb(n1047),.dout(n1051),.clk(gclk));
	jand g0980(.dina(w_dff_B_fIWXbCll5_0),.dinb(n1046),.dout(n1052),.clk(gclk));
	jand g0981(.dina(n1052),.dinb(w_dff_B_rMuyGdqc6_1),.dout(n1053),.clk(gclk));
	jnot g0982(.din(w_n1053_0[2]),.dout(w_dff_A_XSgKg9OT8_1),.clk(gclk));
	jxor g0983(.dina(w_n1036_0[0]),.dinb(w_n772_0[0]),.dout(n1055),.clk(gclk));
	jxor g0984(.dina(n1055),.dinb(w_n1033_0[0]),.dout(n1056),.clk(gclk));
	jor g0985(.dina(w_n1045_0[0]),.dinb(w_n1056_0[1]),.dout(n1057),.clk(gclk));
	jand g0986(.dina(w_n1029_0[1]),.dinb(w_n613_0[1]),.dout(n1058),.clk(gclk));
	jand g0987(.dina(w_dff_B_zeMOrs7R0_0),.dinb(n1057),.dout(n1059),.clk(gclk));
	jand g0988(.dina(w_n1048_0[0]),.dinb(w_n767_0[1]),.dout(n1060),.clk(gclk));
	jand g0989(.dina(w_n566_0[1]),.dinb(w_n457_0[0]),.dout(n1061),.clk(gclk));
	jxor g0990(.dina(w_dff_B_ZjAM4XCm8_0),.dinb(w_n473_0[0]),.dout(n1062),.clk(gclk));
	jxor g0991(.dina(w_n1062_0[1]),.dinb(w_n777_0[0]),.dout(n1063),.clk(gclk));
	jxor g0992(.dina(n1063),.dinb(w_dff_B_wqi3mgeV4_1),.dout(n1064),.clk(gclk));
	jor g0993(.dina(n1064),.dinb(n1059),.dout(n1065),.clk(gclk));
	jor g0994(.dina(n1065),.dinb(w_n614_2[1]),.dout(n1066),.clk(gclk));
	jand g0995(.dina(w_n1062_0[0]),.dinb(w_n618_1[0]),.dout(n1067),.clk(gclk));
	jnot g0996(.din(n1067),.dout(n1068),.clk(gclk));
	jand g0997(.dina(w_G50_2[0]),.dinb(w_G41_0[0]),.dout(n1069),.clk(gclk));
	jor g0998(.dina(w_dff_B_QoyuoMYs5_0),.dinb(w_n680_1[2]),.dout(n1070),.clk(gclk));
	jand g0999(.dina(w_n638_3[1]),.dinb(w_G137_0[2]),.dout(n1071),.clk(gclk));
	jand g1000(.dina(w_n633_2[2]),.dinb(w_G143_1[0]),.dout(n1072),.clk(gclk));
	jand g1001(.dina(w_n651_3[1]),.dinb(w_G125_0[0]),.dout(n1073),.clk(gclk));
	jor g1002(.dina(n1073),.dinb(n1072),.dout(n1074),.clk(gclk));
	jor g1003(.dina(n1074),.dinb(w_dff_B_cQ8DBxlb8_1),.dout(n1075),.clk(gclk));
	jand g1004(.dina(w_n640_3[1]),.dinb(w_dff_B_RAbVov9X1_1),.dout(n1076),.clk(gclk));
	jand g1005(.dina(w_n629_2[0]),.dinb(w_G150_1[1]),.dout(n1077),.clk(gclk));
	jand g1006(.dina(w_n646_3[1]),.dinb(w_G128_0[1]),.dout(n1078),.clk(gclk));
	jor g1007(.dina(w_dff_B_x85OuUaa8_0),.dinb(n1077),.dout(n1079),.clk(gclk));
	jor g1008(.dina(n1079),.dinb(w_dff_B_qQIrSnQJ5_1),.dout(n1080),.clk(gclk));
	jand g1009(.dina(w_n648_1[2]),.dinb(w_G159_1[1]),.dout(n1081),.clk(gclk));
	jand g1010(.dina(w_n653_3[1]),.dinb(w_G132_0[2]),.dout(n1082),.clk(gclk));
	jor g1011(.dina(n1082),.dinb(n1081),.dout(n1083),.clk(gclk));
	jor g1012(.dina(n1083),.dinb(w_G33_4[2]),.dout(n1084),.clk(gclk));
	jor g1013(.dina(w_dff_B_LgGx67mV7_0),.dinb(n1080),.dout(n1085),.clk(gclk));
	jor g1014(.dina(n1085),.dinb(w_dff_B_BK1PEsdO6_1),.dout(n1086),.clk(gclk));
	jand g1015(.dina(w_n653_3[0]),.dinb(w_G97_1[2]),.dout(n1087),.clk(gclk));
	jand g1016(.dina(w_n646_3[0]),.dinb(w_G107_1[2]),.dout(n1088),.clk(gclk));
	jor g1017(.dina(n1088),.dinb(n1087),.dout(n1089),.clk(gclk));
	jnot g1018(.din(n1089),.dout(n1090),.clk(gclk));
	jand g1019(.dina(w_n648_1[1]),.dinb(w_G58_1[2]),.dout(n1091),.clk(gclk));
	jnot g1020(.din(w_n1091_0[1]),.dout(n1092),.clk(gclk));
	jand g1021(.dina(n1092),.dinb(w_n887_0[0]),.dout(n1093),.clk(gclk));
	jand g1022(.dina(n1093),.dinb(n1090),.dout(n1094),.clk(gclk));
	jand g1023(.dina(w_n640_3[0]),.dinb(w_G283_1[1]),.dout(n1095),.clk(gclk));
	jor g1024(.dina(n1095),.dinb(w_n830_0[0]),.dout(n1096),.clk(gclk));
	jand g1025(.dina(w_n651_3[0]),.dinb(w_G116_2[0]),.dout(n1097),.clk(gclk));
	jand g1026(.dina(w_n638_3[0]),.dinb(w_G87_1[0]),.dout(n1098),.clk(gclk));
	jor g1027(.dina(n1098),.dinb(n1097),.dout(n1099),.clk(gclk));
	jor g1028(.dina(w_dff_B_gUOa6haK3_0),.dinb(n1096),.dout(n1100),.clk(gclk));
	jnot g1029(.din(n1100),.dout(n1101),.clk(gclk));
	jand g1030(.dina(n1101),.dinb(w_dff_B_6IigKEW58_1),.dout(n1102),.clk(gclk));
	jand g1031(.dina(n1102),.dinb(w_G33_4[1]),.dout(n1103),.clk(gclk));
	jnot g1032(.din(n1103),.dout(n1104),.clk(gclk));
	jand g1033(.dina(n1104),.dinb(w_dff_B_5RuyAYUz8_1),.dout(n1105),.clk(gclk));
	jand g1034(.dina(n1105),.dinb(w_n163_0[1]),.dout(n1106),.clk(gclk));
	jor g1035(.dina(n1106),.dinb(w_dff_B_mBKeCzen2_1),.dout(n1107),.clk(gclk));
	jand g1036(.dina(w_n741_0[2]),.dinb(w_n73_0[2]),.dout(n1108),.clk(gclk));
	jnot g1037(.din(n1108),.dout(n1109),.clk(gclk));
	jand g1038(.dina(w_dff_B_YoznAWsr8_0),.dinb(n1107),.dout(n1110),.clk(gclk));
	jand g1039(.dina(n1110),.dinb(n1068),.dout(n1111),.clk(gclk));
	jand g1040(.dina(n1111),.dinb(w_n614_2[0]),.dout(n1112),.clk(gclk));
	jnot g1041(.din(n1112),.dout(n1113),.clk(gclk));
	jand g1042(.dina(w_dff_B_ZBwqG1ji1_0),.dinb(n1066),.dout(n1114),.clk(gclk));
	jnot g1043(.din(w_n1114_0[2]),.dout(w_dff_A_lw3JEhUA7_1),.clk(gclk));
	jand g1044(.dina(w_n771_0[1]),.dinb(w_n618_0[2]),.dout(n1116),.clk(gclk));
	jnot g1045(.din(n1116),.dout(n1117),.clk(gclk));
	jand g1046(.dina(w_n646_2[2]),.dinb(w_G283_1[0]),.dout(n1118),.clk(gclk));
	jand g1047(.dina(w_n633_2[1]),.dinb(w_G97_1[1]),.dout(n1119),.clk(gclk));
	jand g1048(.dina(w_n653_2[2]),.dinb(w_G116_1[2]),.dout(n1120),.clk(gclk));
	jor g1049(.dina(n1120),.dinb(n1119),.dout(n1121),.clk(gclk));
	jand g1050(.dina(w_n640_2[2]),.dinb(w_G303_0[2]),.dout(n1122),.clk(gclk));
	jor g1051(.dina(n1122),.dinb(n1121),.dout(n1123),.clk(gclk));
	jor g1052(.dina(n1123),.dinb(w_dff_B_xpsKkW372_1),.dout(n1124),.clk(gclk));
	jor g1053(.dina(w_n884_0[0]),.dinb(w_n833_0[0]),.dout(n1125),.clk(gclk));
	jand g1054(.dina(w_n651_2[2]),.dinb(w_G294_1[0]),.dout(n1126),.clk(gclk));
	jand g1055(.dina(w_n638_2[2]),.dinb(w_G107_1[1]),.dout(n1127),.clk(gclk));
	jor g1056(.dina(n1127),.dinb(n1126),.dout(n1128),.clk(gclk));
	jor g1057(.dina(n1128),.dinb(w_n153_2[2]),.dout(n1129),.clk(gclk));
	jor g1058(.dina(n1129),.dinb(n1125),.dout(n1130),.clk(gclk));
	jor g1059(.dina(n1130),.dinb(n1124),.dout(n1131),.clk(gclk));
	jand g1060(.dina(w_n646_2[1]),.dinb(w_G137_0[1]),.dout(n1132),.clk(gclk));
	jand g1061(.dina(w_n633_2[0]),.dinb(w_G159_1[0]),.dout(n1133),.clk(gclk));
	jand g1062(.dina(w_n638_2[1]),.dinb(w_G150_1[0]),.dout(n1134),.clk(gclk));
	jor g1063(.dina(n1134),.dinb(n1133),.dout(n1135),.clk(gclk));
	jand g1064(.dina(w_n651_2[1]),.dinb(w_G132_0[1]),.dout(n1136),.clk(gclk));
	jand g1065(.dina(w_n629_1[2]),.dinb(w_G50_1[2]),.dout(n1137),.clk(gclk));
	jor g1066(.dina(n1137),.dinb(w_n1091_0[0]),.dout(n1138),.clk(gclk));
	jor g1067(.dina(n1138),.dinb(w_dff_B_vMDHdvrG4_1),.dout(n1139),.clk(gclk));
	jand g1068(.dina(w_n653_2[1]),.dinb(w_G143_0[2]),.dout(n1140),.clk(gclk));
	jand g1069(.dina(w_n640_2[1]),.dinb(w_G128_0[0]),.dout(n1141),.clk(gclk));
	jor g1070(.dina(n1141),.dinb(w_dff_B_mdsd82Yu5_1),.dout(n1142),.clk(gclk));
	jor g1071(.dina(n1142),.dinb(w_G33_4[0]),.dout(n1143),.clk(gclk));
	jor g1072(.dina(n1143),.dinb(n1139),.dout(n1144),.clk(gclk));
	jor g1073(.dina(n1144),.dinb(w_dff_B_TQMJOALO8_1),.dout(n1145),.clk(gclk));
	jor g1074(.dina(n1145),.dinb(w_dff_B_mKbZNNwd7_1),.dout(n1146),.clk(gclk));
	jand g1075(.dina(n1146),.dinb(w_dff_B_NlD4pxdV4_1),.dout(n1147),.clk(gclk));
	jor g1076(.dina(n1147),.dinb(w_n680_1[1]),.dout(n1148),.clk(gclk));
	jand g1077(.dina(w_n741_0[1]),.dinb(w_n75_0[2]),.dout(n1149),.clk(gclk));
	jnot g1078(.din(n1149),.dout(n1150),.clk(gclk));
	jand g1079(.dina(w_dff_B_LQeloxLE6_0),.dinb(n1148),.dout(n1151),.clk(gclk));
	jand g1080(.dina(w_dff_B_48tfzXcl0_0),.dinb(n1117),.dout(n1152),.clk(gclk));
	jand g1081(.dina(n1152),.dinb(w_n614_1[2]),.dout(n1153),.clk(gclk));
	jnot g1082(.din(n1153),.dout(n1154),.clk(gclk));
	jor g1083(.dina(w_n1041_0[0]),.dinb(w_n1056_0[0]),.dout(n1155),.clk(gclk));
	jnot g1084(.din(w_n1029_0[0]),.dout(n1156),.clk(gclk));
	jor g1085(.dina(w_n1040_0[0]),.dinb(w_dff_B_kjZSD6wT0_1),.dout(n1157),.clk(gclk));
	jand g1086(.dina(w_dff_B_3mkVTSnB2_0),.dinb(n1155),.dout(n1158),.clk(gclk));
	jand g1087(.dina(n1158),.dinb(w_dff_B_LHKZR8h56_1),.dout(n1159),.clk(gclk));
	jnot g1088(.din(w_n1159_0[2]),.dout(w_dff_A_qbIctODl9_1),.clk(gclk));
	jand g1089(.dina(w_n1114_0[1]),.dinb(w_n1053_0[1]),.dout(n1161),.clk(gclk));
	jand g1090(.dina(w_n1159_0[1]),.dinb(w_n759_0[0]),.dout(n1162),.clk(gclk));
	jand g1091(.dina(w_n987_0[1]),.dinb(w_n869_0[1]),.dout(n1163),.clk(gclk));
	jnot g1092(.din(w_G396_0),.dout(n1164),.clk(gclk));
	jand g1093(.dina(w_n937_0[1]),.dinb(w_n1164_0[1]),.dout(n1165),.clk(gclk));
	jand g1094(.dina(w_dff_B_48cNaTjh5_0),.dinb(n1163),.dout(n1166),.clk(gclk));
	jand g1095(.dina(w_dff_B_AmjHcgx98_0),.dinb(n1162),.dout(n1167),.clk(gclk));
	jand g1096(.dina(n1167),.dinb(w_n1161_0[1]),.dout(n1168),.clk(gclk));
	jnot g1097(.din(w_n1168_0[1]),.dout(w_dff_A_0IWw5YRT1_1),.clk(gclk));
	jnot g1098(.din(w_G343_0[0]),.dout(n1170),.clk(gclk));
	jand g1099(.dina(w_n1161_0[0]),.dinb(w_n1170_0[1]),.dout(n1171),.clk(gclk));
	jnot g1100(.din(w_G213_0[1]),.dout(n1172),.clk(gclk));
	jor g1101(.dina(w_n1168_0[0]),.dinb(w_dff_B_FwJFZ6BF6_1),.dout(n1173),.clk(gclk));
	jor g1102(.dina(n1173),.dinb(w_dff_B_frMcGxgf5_1),.dout(G409),.clk(gclk));
	jxor g1103(.dina(w_n937_0[0]),.dinb(w_n1164_0[0]),.dout(n1175),.clk(gclk));
	jxor g1104(.dina(w_n987_0[0]),.dinb(w_n869_0[0]),.dout(n1176),.clk(gclk));
	jxor g1105(.dina(n1176),.dinb(w_dff_B_V5R8BYO09_1),.dout(n1177),.clk(gclk));
	jand g1106(.dina(w_n1170_0[0]),.dinb(w_G213_0[0]),.dout(n1178),.clk(gclk));
	jxor g1107(.dina(w_n1159_0[0]),.dinb(w_G384_0),.dout(n1179),.clk(gclk));
	jxor g1108(.dina(w_n1179_0[1]),.dinb(w_dff_B_fhFDzsU53_1),.dout(n1180),.clk(gclk));
	jand g1109(.dina(n1180),.dinb(w_n1178_0[1]),.dout(n1181),.clk(gclk));
	jnot g1110(.din(w_n1178_0[0]),.dout(n1182),.clk(gclk));
	jxor g1111(.dina(w_n1114_0[0]),.dinb(w_n1053_0[0]),.dout(n1183),.clk(gclk));
	jxor g1112(.dina(n1183),.dinb(w_n1179_0[0]),.dout(n1184),.clk(gclk));
	jand g1113(.dina(w_n1184_0[1]),.dinb(w_dff_B_lY2Ax7b13_1),.dout(n1185),.clk(gclk));
	jor g1114(.dina(n1185),.dinb(n1181),.dout(n1186),.clk(gclk));
	jxor g1115(.dina(n1186),.dinb(w_n1177_0[1]),.dout(G405),.clk(gclk));
	jxor g1116(.dina(w_n1184_0[0]),.dinb(w_n1177_0[0]),.dout(w_dff_A_A80hFMiP3_2),.clk(gclk));
	jspl3 jspl3_w_G1_0(.douta(w_G1_0[0]),.doutb(w_G1_0[1]),.doutc(w_dff_A_7986Ijkt6_2),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_dff_A_yWAHEjrD4_0),.doutb(w_G1_1[1]),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl jspl_w_G1_2(.douta(w_G1_2[0]),.doutb(w_dff_A_rJrIH5jY5_1),.din(w_G1_0[1]));
	jspl3 jspl3_w_G13_0(.douta(w_G13_0[0]),.doutb(w_G13_0[1]),.doutc(w_G13_0[2]),.din(G13));
	jspl3 jspl3_w_G13_1(.douta(w_dff_A_X78oElrO3_0),.doutb(w_dff_A_XMenjuw07_1),.doutc(w_G13_1[2]),.din(w_G13_0[0]));
	jspl jspl_w_G13_2(.douta(w_dff_A_qgnPfh6H0_0),.doutb(w_G13_2[1]),.din(w_G13_0[1]));
	jspl3 jspl3_w_G20_0(.douta(w_G20_0[0]),.doutb(w_G20_0[1]),.doutc(w_dff_A_IRLX5wUz8_2),.din(G20));
	jspl3 jspl3_w_G20_1(.douta(w_dff_A_8uDIUc495_0),.doutb(w_G20_1[1]),.doutc(w_G20_1[2]),.din(w_G20_0[0]));
	jspl3 jspl3_w_G20_2(.douta(w_G20_2[0]),.doutb(w_G20_2[1]),.doutc(w_dff_A_kYWp7nK21_2),.din(w_G20_0[1]));
	jspl3 jspl3_w_G20_3(.douta(w_G20_3[0]),.doutb(w_G20_3[1]),.doutc(w_dff_A_gRveNVBj0_2),.din(w_G20_0[2]));
	jspl3 jspl3_w_G20_4(.douta(w_G20_4[0]),.doutb(w_dff_A_Bn1ER3N95_1),.doutc(w_dff_A_aSoHVQ5s5_2),.din(w_G20_1[0]));
	jspl3 jspl3_w_G20_5(.douta(w_dff_A_DjzwFZwv6_0),.doutb(w_G20_5[1]),.doutc(w_G20_5[2]),.din(w_G20_1[1]));
	jspl3 jspl3_w_G20_6(.douta(w_dff_A_7JrKyfu22_0),.doutb(w_G20_6[1]),.doutc(w_dff_A_smLdoHTq5_2),.din(w_G20_1[2]));
	jspl3 jspl3_w_G33_0(.douta(w_dff_A_x0xr0h3r0_0),.doutb(w_G33_0[1]),.doutc(w_G33_0[2]),.din(G33));
	jspl3 jspl3_w_G33_1(.douta(w_dff_A_3Ekhpmm29_0),.doutb(w_dff_A_wUc9r8FB4_1),.doutc(w_G33_1[2]),.din(w_G33_0[0]));
	jspl3 jspl3_w_G33_2(.douta(w_G33_2[0]),.doutb(w_G33_2[1]),.doutc(w_G33_2[2]),.din(w_G33_0[1]));
	jspl3 jspl3_w_G33_3(.douta(w_G33_3[0]),.doutb(w_G33_3[1]),.doutc(w_G33_3[2]),.din(w_G33_0[2]));
	jspl3 jspl3_w_G33_4(.douta(w_dff_A_6WtM1vEI3_0),.doutb(w_dff_A_0zdnIMgX1_1),.doutc(w_G33_4[2]),.din(w_G33_1[0]));
	jspl3 jspl3_w_G33_5(.douta(w_G33_5[0]),.doutb(w_dff_A_CzPuB0WY5_1),.doutc(w_G33_5[2]),.din(w_G33_1[1]));
	jspl3 jspl3_w_G33_6(.douta(w_dff_A_57ZRTMa09_0),.doutb(w_dff_A_ZslAtP5G6_1),.doutc(w_G33_6[2]),.din(w_G33_1[2]));
	jspl3 jspl3_w_G33_7(.douta(w_dff_A_C9Ok3oI29_0),.doutb(w_dff_A_Ilws0PQQ1_1),.doutc(w_G33_7[2]),.din(w_G33_2[0]));
	jspl3 jspl3_w_G33_8(.douta(w_G33_8[0]),.doutb(w_dff_A_C6fhdDYB1_1),.doutc(w_G33_8[2]),.din(w_G33_2[1]));
	jspl3 jspl3_w_G33_9(.douta(w_dff_A_ZW7DFe3L2_0),.doutb(w_dff_A_kt8vfdUT2_1),.doutc(w_G33_9[2]),.din(w_G33_2[2]));
	jspl3 jspl3_w_G33_10(.douta(w_G33_10[0]),.doutb(w_G33_10[1]),.doutc(w_G33_10[2]),.din(w_G33_3[0]));
	jspl3 jspl3_w_G33_11(.douta(w_G33_11[0]),.doutb(w_G33_11[1]),.doutc(w_G33_11[2]),.din(w_G33_3[1]));
	jspl3 jspl3_w_G33_12(.douta(w_G33_12[0]),.doutb(w_dff_A_y5QVgwBk6_1),.doutc(w_dff_A_2A6upE0W0_2),.din(w_G33_3[2]));
	jspl3 jspl3_w_G41_0(.douta(w_G41_0[0]),.doutb(w_G41_0[1]),.doutc(w_G41_0[2]),.din(G41));
	jspl3 jspl3_w_G45_0(.douta(w_G45_0[0]),.doutb(w_dff_A_WlqT3q5V3_1),.doutc(w_G45_0[2]),.din(G45));
	jspl jspl_w_G45_1(.douta(w_G45_1[0]),.doutb(w_dff_A_iD4J6MS45_1),.din(w_G45_0[0]));
	jspl3 jspl3_w_G50_0(.douta(w_G50_0[0]),.doutb(w_G50_0[1]),.doutc(w_G50_0[2]),.din(G50));
	jspl3 jspl3_w_G50_1(.douta(w_dff_A_X3FU8xLS8_0),.doutb(w_G50_1[1]),.doutc(w_dff_A_hpXedVji2_2),.din(w_G50_0[0]));
	jspl3 jspl3_w_G50_2(.douta(w_G50_2[0]),.doutb(w_dff_A_klVsZxkz3_1),.doutc(w_dff_A_uchtVzkm2_2),.din(w_G50_0[1]));
	jspl3 jspl3_w_G50_3(.douta(w_dff_A_AU5f9WES5_0),.doutb(w_dff_A_tzRFdULo5_1),.doutc(w_G50_3[2]),.din(w_G50_0[2]));
	jspl3 jspl3_w_G50_4(.douta(w_dff_A_mmRpLKz87_0),.doutb(w_dff_A_3CWmlWEH5_1),.doutc(w_G50_4[2]),.din(w_G50_1[0]));
	jspl3 jspl3_w_G50_5(.douta(w_G50_5[0]),.doutb(w_dff_A_XaU3ZVoN5_1),.doutc(w_G50_5[2]),.din(w_G50_1[1]));
	jspl3 jspl3_w_G58_0(.douta(w_G58_0[0]),.doutb(w_dff_A_4sD7ZGpF7_1),.doutc(w_G58_0[2]),.din(G58));
	jspl3 jspl3_w_G58_1(.douta(w_G58_1[0]),.doutb(w_G58_1[1]),.doutc(w_dff_A_9njr8Asa5_2),.din(w_G58_0[0]));
	jspl3 jspl3_w_G58_2(.douta(w_dff_A_F1LSShtC4_0),.doutb(w_G58_2[1]),.doutc(w_dff_A_E72xmQJQ7_2),.din(w_G58_0[1]));
	jspl3 jspl3_w_G58_3(.douta(w_dff_A_xkJlU7Il1_0),.doutb(w_G58_3[1]),.doutc(w_dff_A_0y1D0MhM1_2),.din(w_G58_0[2]));
	jspl3 jspl3_w_G58_4(.douta(w_dff_A_uVJ5F7Xq3_0),.doutb(w_G58_4[1]),.doutc(w_dff_A_vIZPcx7T9_2),.din(w_G58_1[0]));
	jspl3 jspl3_w_G58_5(.douta(w_dff_A_vd9Cswqp1_0),.doutb(w_G58_5[1]),.doutc(w_G58_5[2]),.din(w_G58_1[1]));
	jspl3 jspl3_w_G68_0(.douta(w_G68_0[0]),.doutb(w_G68_0[1]),.doutc(w_dff_A_MoPl1Dqo0_2),.din(G68));
	jspl3 jspl3_w_G68_1(.douta(w_G68_1[0]),.doutb(w_G68_1[1]),.doutc(w_dff_A_pbAlY6TH8_2),.din(w_G68_0[0]));
	jspl3 jspl3_w_G68_2(.douta(w_G68_2[0]),.doutb(w_dff_A_NG3RrSe38_1),.doutc(w_dff_A_9LWVJ9J94_2),.din(w_G68_0[1]));
	jspl3 jspl3_w_G68_3(.douta(w_G68_3[0]),.doutb(w_dff_A_toJ0YaT87_1),.doutc(w_dff_A_5JEDc2PT9_2),.din(w_G68_0[2]));
	jspl3 jspl3_w_G68_4(.douta(w_dff_A_DRU23pch3_0),.doutb(w_G68_4[1]),.doutc(w_dff_A_9NFBB2sh2_2),.din(w_G68_1[0]));
	jspl3 jspl3_w_G68_5(.douta(w_dff_A_54F53hGA1_0),.doutb(w_G68_5[1]),.doutc(w_G68_5[2]),.din(w_G68_1[1]));
	jspl3 jspl3_w_G77_0(.douta(w_G77_0[0]),.doutb(w_dff_A_vDc3UwJq2_1),.doutc(w_G77_0[2]),.din(G77));
	jspl3 jspl3_w_G77_1(.douta(w_G77_1[0]),.doutb(w_dff_A_aC0WX6qI9_1),.doutc(w_G77_1[2]),.din(w_G77_0[0]));
	jspl3 jspl3_w_G77_2(.douta(w_dff_A_GJ0JER405_0),.doutb(w_dff_A_8PYxwOD49_1),.doutc(w_G77_2[2]),.din(w_G77_0[1]));
	jspl3 jspl3_w_G77_3(.douta(w_dff_A_XdFUXiYj2_0),.doutb(w_G77_3[1]),.doutc(w_dff_A_SSQAyeQo5_2),.din(w_G77_0[2]));
	jspl3 jspl3_w_G77_4(.douta(w_dff_A_165wfq2N1_0),.doutb(w_G77_4[1]),.doutc(w_G77_4[2]),.din(w_G77_1[0]));
	jspl3 jspl3_w_G87_0(.douta(w_dff_A_MFLTO2Ch3_0),.doutb(w_G87_0[1]),.doutc(w_G87_0[2]),.din(G87));
	jspl3 jspl3_w_G87_1(.douta(w_G87_1[0]),.doutb(w_dff_A_z1JNQAMu2_1),.doutc(w_dff_A_QAlOaucd4_2),.din(w_G87_0[0]));
	jspl3 jspl3_w_G87_2(.douta(w_dff_A_8KS8086U1_0),.doutb(w_dff_A_Z5pizf2f2_1),.doutc(w_G87_2[2]),.din(w_G87_0[1]));
	jspl3 jspl3_w_G87_3(.douta(w_dff_A_1FSyIZIT2_0),.doutb(w_G87_3[1]),.doutc(w_G87_3[2]),.din(w_G87_0[2]));
	jspl3 jspl3_w_G97_0(.douta(w_G97_0[0]),.doutb(w_dff_A_4EL6Kdd02_1),.doutc(w_G97_0[2]),.din(G97));
	jspl3 jspl3_w_G97_1(.douta(w_G97_1[0]),.doutb(w_dff_A_jZz3IHDG8_1),.doutc(w_dff_A_2dNZana21_2),.din(w_G97_0[0]));
	jspl3 jspl3_w_G97_2(.douta(w_G97_2[0]),.doutb(w_dff_A_VOJ3Gx0C6_1),.doutc(w_G97_2[2]),.din(w_G97_0[1]));
	jspl3 jspl3_w_G97_3(.douta(w_dff_A_4Ryte8mL2_0),.doutb(w_G97_3[1]),.doutc(w_G97_3[2]),.din(w_G97_0[2]));
	jspl3 jspl3_w_G97_4(.douta(w_dff_A_E5wgSxP68_0),.doutb(w_G97_4[1]),.doutc(w_G97_4[2]),.din(w_G97_1[0]));
	jspl3 jspl3_w_G107_0(.douta(w_G107_0[0]),.doutb(w_dff_A_pPVzhuRw2_1),.doutc(w_G107_0[2]),.din(G107));
	jspl3 jspl3_w_G107_1(.douta(w_G107_1[0]),.doutb(w_dff_A_so2b6Mk06_1),.doutc(w_dff_A_YdIp8JhS8_2),.din(w_G107_0[0]));
	jspl3 jspl3_w_G107_2(.douta(w_G107_2[0]),.doutb(w_dff_A_HEyFGdAl1_1),.doutc(w_G107_2[2]),.din(w_G107_0[1]));
	jspl3 jspl3_w_G107_3(.douta(w_dff_A_BBf4G9ah5_0),.doutb(w_G107_3[1]),.doutc(w_G107_3[2]),.din(w_G107_0[2]));
	jspl jspl_w_G107_4(.douta(w_dff_A_LArgObzU8_0),.doutb(w_G107_4[1]),.din(w_G107_1[0]));
	jspl3 jspl3_w_G116_0(.douta(w_G116_0[0]),.doutb(w_dff_A_K6dqxKfC2_1),.doutc(w_dff_A_YMOYBBOY5_2),.din(G116));
	jspl3 jspl3_w_G116_1(.douta(w_G116_1[0]),.doutb(w_G116_1[1]),.doutc(w_dff_A_BHeSO7qT3_2),.din(w_G116_0[0]));
	jspl3 jspl3_w_G116_2(.douta(w_G116_2[0]),.doutb(w_G116_2[1]),.doutc(w_dff_A_gsN1zYW38_2),.din(w_G116_0[1]));
	jspl3 jspl3_w_G116_3(.douta(w_G116_3[0]),.doutb(w_G116_3[1]),.doutc(w_G116_3[2]),.din(w_G116_0[2]));
	jspl3 jspl3_w_G116_4(.douta(w_dff_A_hiFDXRRs9_0),.doutb(w_G116_4[1]),.doutc(w_G116_4[2]),.din(w_G116_1[0]));
	jspl3 jspl3_w_G116_5(.douta(w_dff_A_cPT0Uvut7_0),.doutb(w_dff_A_xm7aeCbx9_1),.doutc(w_G116_5[2]),.din(w_G116_1[1]));
	jspl jspl_w_G125_0(.douta(w_G125_0[0]),.doutb(w_dff_A_OAACL1iP1_1),.din(w_dff_B_NXq1WUpR1_2));
	jspl3 jspl3_w_G128_0(.douta(w_dff_A_UshgANoK0_0),.doutb(w_G128_0[1]),.doutc(w_G128_0[2]),.din(w_dff_B_5uutoYik1_3));
	jspl3 jspl3_w_G132_0(.douta(w_G132_0[0]),.doutb(w_G132_0[1]),.doutc(w_G132_0[2]),.din(w_dff_B_UP0PQyuR2_3));
	jspl jspl_w_G132_1(.douta(w_G132_1[0]),.doutb(w_dff_A_uvenekGE3_1),.din(w_G132_0[0]));
	jspl3 jspl3_w_G137_0(.douta(w_G137_0[0]),.doutb(w_G137_0[1]),.doutc(w_G137_0[2]),.din(w_dff_B_szlZOZXh5_3));
	jspl3 jspl3_w_G137_1(.douta(w_G137_1[0]),.doutb(w_dff_A_zT8TQK0W9_1),.doutc(w_G137_1[2]),.din(w_G137_0[0]));
	jspl3 jspl3_w_G143_0(.douta(w_G143_0[0]),.doutb(w_G143_0[1]),.doutc(w_G143_0[2]),.din(w_dff_B_1WN0ZySe4_3));
	jspl3 jspl3_w_G143_1(.douta(w_G143_1[0]),.doutb(w_G143_1[1]),.doutc(w_dff_A_s0qi0ndp0_2),.din(w_G143_0[0]));
	jspl jspl_w_G143_2(.douta(w_G143_2[0]),.doutb(w_G143_2[1]),.din(w_G143_0[1]));
	jspl3 jspl3_w_G150_0(.douta(w_dff_A_YVUJFrSK3_0),.doutb(w_dff_A_cZPzdJwJ2_1),.doutc(w_G150_0[2]),.din(w_dff_B_fxZ7pw9z2_3));
	jspl3 jspl3_w_G150_1(.douta(w_G150_1[0]),.doutb(w_dff_A_vt49kmHw4_1),.doutc(w_G150_1[2]),.din(w_G150_0[0]));
	jspl3 jspl3_w_G150_2(.douta(w_G150_2[0]),.doutb(w_dff_A_67XSxAJS6_1),.doutc(w_G150_2[2]),.din(w_G150_0[1]));
	jspl jspl_w_G150_3(.douta(w_dff_A_PmkHxSYn8_0),.doutb(w_G150_3[1]),.din(w_G150_0[2]));
	jspl3 jspl3_w_G159_0(.douta(w_dff_A_HlTdhWGI7_0),.doutb(w_dff_A_icJRTxbs6_1),.doutc(w_G159_0[2]),.din(G159));
	jspl3 jspl3_w_G159_1(.douta(w_G159_1[0]),.doutb(w_G159_1[1]),.doutc(w_dff_A_2Jr8D4s51_2),.din(w_G159_0[0]));
	jspl3 jspl3_w_G159_2(.douta(w_G159_2[0]),.doutb(w_G159_2[1]),.doutc(w_G159_2[2]),.din(w_G159_0[1]));
	jspl3 jspl3_w_G159_3(.douta(w_dff_A_F3hCORgC0_0),.doutb(w_dff_A_oXxWy2579_1),.doutc(w_G159_3[2]),.din(w_G159_0[2]));
	jspl3 jspl3_w_G169_0(.douta(w_dff_A_q2xWHlDq8_0),.doutb(w_dff_A_Dy3TAhzW2_1),.doutc(w_G169_0[2]),.din(G169));
	jspl3 jspl3_w_G169_1(.douta(w_G169_1[0]),.doutb(w_dff_A_RVQRq0Pq2_1),.doutc(w_dff_A_3krxqJlc2_2),.din(w_G169_0[0]));
	jspl3 jspl3_w_G169_2(.douta(w_dff_A_Qsh7UEam8_0),.doutb(w_dff_A_NH0586Nw4_1),.doutc(w_G169_2[2]),.din(w_G169_0[1]));
	jspl jspl_w_G169_3(.douta(w_G169_3[0]),.doutb(w_dff_A_gNdOfnno1_1),.din(w_G169_0[2]));
	jspl3 jspl3_w_G179_0(.douta(w_dff_A_oNI79irw8_0),.doutb(w_G179_0[1]),.doutc(w_G179_0[2]),.din(G179));
	jspl3 jspl3_w_G179_1(.douta(w_G179_1[0]),.doutb(w_G179_1[1]),.doutc(w_G179_1[2]),.din(w_G179_0[0]));
	jspl3 jspl3_w_G179_2(.douta(w_dff_A_RKSuQUOB6_0),.doutb(w_dff_A_2EJuJVo33_1),.doutc(w_G179_2[2]),.din(w_G179_0[1]));
	jspl3 jspl3_w_G190_0(.douta(w_dff_A_vQANGHd58_0),.doutb(w_G190_0[1]),.doutc(w_dff_A_ew18bozs6_2),.din(G190));
	jspl3 jspl3_w_G190_1(.douta(w_dff_A_naQTATWe7_0),.doutb(w_G190_1[1]),.doutc(w_G190_1[2]),.din(w_G190_0[0]));
	jspl3 jspl3_w_G190_2(.douta(w_dff_A_JQqvRTx24_0),.doutb(w_G190_2[1]),.doutc(w_dff_A_5eVJVE8F5_2),.din(w_G190_0[1]));
	jspl3 jspl3_w_G190_3(.douta(w_dff_A_78XtRBs74_0),.doutb(w_dff_A_5hmUbngm0_1),.doutc(w_G190_3[2]),.din(w_G190_0[2]));
	jspl3 jspl3_w_G190_4(.douta(w_G190_4[0]),.doutb(w_dff_A_Su0dW8rr4_1),.doutc(w_dff_A_R3WQr2sD2_2),.din(w_G190_1[0]));
	jspl3 jspl3_w_G200_0(.douta(w_G200_0[0]),.doutb(w_G200_0[1]),.doutc(w_dff_A_gXQuaMnl3_2),.din(G200));
	jspl3 jspl3_w_G200_1(.douta(w_dff_A_JtIPGaNL4_0),.doutb(w_G200_1[1]),.doutc(w_dff_A_9DcS5XPD4_2),.din(w_G200_0[0]));
	jspl3 jspl3_w_G200_2(.douta(w_G200_2[0]),.doutb(w_dff_A_5fvJvEOG9_1),.doutc(w_dff_A_KRBhaKoL6_2),.din(w_G200_0[1]));
	jspl jspl_w_G200_3(.douta(w_G200_3[0]),.doutb(w_G200_3[1]),.din(w_G200_0[2]));
	jspl3 jspl3_w_G213_0(.douta(w_dff_A_rUnl0ppz2_0),.doutb(w_G213_0[1]),.doutc(w_dff_A_YSi94fau9_2),.din(G213));
	jspl jspl_w_G223_0(.douta(w_G223_0[0]),.doutb(w_G223_0[1]),.din(w_dff_B_F2IAu7YI9_2));
	jspl3 jspl3_w_G226_0(.douta(w_G226_0[0]),.doutb(w_dff_A_X1tZQeR31_1),.doutc(w_dff_A_sEVsS5Ua6_2),.din(G226));
	jspl3 jspl3_w_G226_1(.douta(w_dff_A_SpIpFv3q9_0),.doutb(w_G226_1[1]),.doutc(w_G226_1[2]),.din(w_G226_0[0]));
	jspl3 jspl3_w_G232_0(.douta(w_G232_0[0]),.doutb(w_dff_A_sM4oKHqN0_1),.doutc(w_dff_A_73qoDkLk9_2),.din(G232));
	jspl3 jspl3_w_G232_1(.douta(w_dff_A_Gus10aQ47_0),.doutb(w_G232_1[1]),.doutc(w_G232_1[2]),.din(w_G232_0[0]));
	jspl3 jspl3_w_G238_0(.douta(w_dff_A_aXlyl3Fd0_0),.doutb(w_dff_A_AwnHk9988_1),.doutc(w_G238_0[2]),.din(G238));
	jspl3 jspl3_w_G244_0(.douta(w_G244_0[0]),.doutb(w_dff_A_oRkKDqT53_1),.doutc(w_dff_A_NS8jNmWs2_2),.din(G244));
	jspl jspl_w_G244_1(.douta(w_dff_A_A8RKeC036_0),.doutb(w_G244_1[1]),.din(w_G244_0[0]));
	jspl3 jspl3_w_G250_0(.douta(w_dff_A_O35QWYi73_0),.doutb(w_G250_0[1]),.doutc(w_G250_0[2]),.din(G250));
	jspl3 jspl3_w_G257_0(.douta(w_G257_0[0]),.doutb(w_dff_A_kuQLI3Vo2_1),.doutc(w_dff_A_7LBgXwEW5_2),.din(G257));
	jspl3 jspl3_w_G257_1(.douta(w_dff_A_Qvpf57IH7_0),.doutb(w_G257_1[1]),.doutc(w_G257_1[2]),.din(w_G257_0[0]));
	jspl3 jspl3_w_G264_0(.douta(w_dff_A_UybTJBfR0_0),.doutb(w_dff_A_wW8gMsRw4_1),.doutc(w_G264_0[2]),.din(G264));
	jspl3 jspl3_w_G270_0(.douta(w_dff_A_oU1nba1o6_0),.doutb(w_dff_A_TgPEKW4v9_1),.doutc(w_G270_0[2]),.din(G270));
	jspl3 jspl3_w_G274_0(.douta(w_dff_A_YNlKx5VQ6_0),.doutb(w_G274_0[1]),.doutc(w_dff_A_ZYdtO75G0_2),.din(G274));
	jspl3 jspl3_w_G283_0(.douta(w_dff_A_4FvfAcLi4_0),.doutb(w_dff_A_u11qo1Wn5_1),.doutc(w_G283_0[2]),.din(G283));
	jspl3 jspl3_w_G283_1(.douta(w_G283_1[0]),.doutb(w_dff_A_b6RVrugm3_1),.doutc(w_G283_1[2]),.din(w_G283_0[0]));
	jspl3 jspl3_w_G283_2(.douta(w_G283_2[0]),.doutb(w_dff_A_VexwC1p14_1),.doutc(w_G283_2[2]),.din(w_G283_0[1]));
	jspl3 jspl3_w_G283_3(.douta(w_dff_A_M3o1gwDr0_0),.doutb(w_dff_A_YSKr3QoK9_1),.doutc(w_G283_3[2]),.din(w_G283_0[2]));
	jspl3 jspl3_w_G294_0(.douta(w_dff_A_mOudWFRR2_0),.doutb(w_dff_A_ighade174_1),.doutc(w_G294_0[2]),.din(G294));
	jspl3 jspl3_w_G294_1(.douta(w_G294_1[0]),.doutb(w_dff_A_6ms29Wfm8_1),.doutc(w_G294_1[2]),.din(w_G294_0[0]));
	jspl3 jspl3_w_G294_2(.douta(w_G294_2[0]),.doutb(w_G294_2[1]),.doutc(w_G294_2[2]),.din(w_G294_0[1]));
	jspl jspl_w_G294_3(.douta(w_dff_A_OzvO7sgZ4_0),.doutb(w_G294_3[1]),.din(w_G294_0[2]));
	jspl3 jspl3_w_G303_0(.douta(w_dff_A_cftYHiFH1_0),.doutb(w_G303_0[1]),.doutc(w_dff_A_Az6zVtTd4_2),.din(G303));
	jspl3 jspl3_w_G303_1(.douta(w_G303_1[0]),.doutb(w_G303_1[1]),.doutc(w_G303_1[2]),.din(w_G303_0[0]));
	jspl3 jspl3_w_G303_2(.douta(w_dff_A_y9csACmr9_0),.doutb(w_dff_A_tGoKlo0V2_1),.doutc(w_G303_2[2]),.din(w_G303_0[1]));
	jspl3 jspl3_w_G311_0(.douta(w_G311_0[0]),.doutb(w_G311_0[1]),.doutc(w_G311_0[2]),.din(w_dff_B_WJf49pZb6_3));
	jspl3 jspl3_w_G311_1(.douta(w_G311_1[0]),.doutb(w_dff_A_uHrmcmKh9_1),.doutc(w_G311_1[2]),.din(w_G311_0[0]));
	jspl3 jspl3_w_G317_0(.douta(w_G317_0[0]),.doutb(w_G317_0[1]),.doutc(w_G317_0[2]),.din(w_dff_B_lCwqRcNN5_3));
	jspl jspl_w_G317_1(.douta(w_dff_A_FScjjiaP9_0),.doutb(w_G317_1[1]),.din(w_G317_0[0]));
	jspl3 jspl3_w_G322_0(.douta(w_dff_A_eumKDIYD0_0),.doutb(w_G322_0[1]),.doutc(w_G322_0[2]),.din(w_dff_B_SsOHuoV00_3));
	jspl jspl_w_G326_0(.douta(w_dff_A_3oePydcL6_0),.doutb(w_G326_0[1]),.din(w_dff_B_lMmWfDJV8_2));
	jspl3 jspl3_w_G330_0(.douta(w_dff_A_2czuDZR02_0),.doutb(w_G330_0[1]),.doutc(w_dff_A_TSdrlmcq5_2),.din(w_dff_B_C95NgCdz3_3));
	jspl jspl_w_G343_0(.douta(w_G343_0[0]),.doutb(w_dff_A_WVSrChD69_1),.din(G343));
	jspl3 jspl3_w_G1698_0(.douta(w_G1698_0[0]),.doutb(w_G1698_0[1]),.doutc(w_dff_A_vjQCyBhw6_2),.din(G1698));
	jspl jspl_w_G355_0(.douta(w_dff_A_3oPoLBjJ4_0),.doutb(w_dff_A_jteEvgx45_1),.din(G355_fa_));
	jspl jspl_w_G396_0(.douta(w_G396_0),.doutb(w_dff_A_7VLwJoOx0_1),.din(G396_fa_));
	jspl jspl_w_G384_0(.douta(w_dff_A_KkTi9hGO7_0),.doutb(w_dff_A_cMTHFec67_1),.din(G384_fa_));
	jspl3 jspl3_w_n72_0(.douta(w_n72_0[0]),.doutb(w_dff_A_BXQjOJiv0_1),.doutc(w_dff_A_AZmo76qN7_2),.din(n72));
	jspl3 jspl3_w_n72_1(.douta(w_n72_1[0]),.doutb(w_n72_1[1]),.doutc(w_dff_A_PPac0J2D5_2),.din(w_n72_0[0]));
	jspl3 jspl3_w_n73_0(.douta(w_n73_0[0]),.doutb(w_n73_0[1]),.doutc(w_dff_A_tF8vX1f22_2),.din(n73));
	jspl3 jspl3_w_n73_1(.douta(w_n73_1[0]),.doutb(w_dff_A_Ye7xy3Ka0_1),.doutc(w_dff_A_hCY0c5F84_2),.din(w_n73_0[0]));
	jspl3 jspl3_w_n73_2(.douta(w_dff_A_d5tGjkKH7_0),.doutb(w_n73_2[1]),.doutc(w_dff_A_SGTn5YJd4_2),.din(w_n73_0[1]));
	jspl3 jspl3_w_n74_0(.douta(w_n74_0[0]),.doutb(w_n74_0[1]),.doutc(w_dff_A_KgkWMurd5_2),.din(n74));
	jspl3 jspl3_w_n74_1(.douta(w_n74_1[0]),.doutb(w_dff_A_eaHt07N52_1),.doutc(w_dff_A_Cx0w8QtE6_2),.din(w_n74_0[0]));
	jspl jspl_w_n74_2(.douta(w_n74_2[0]),.doutb(w_n74_2[1]),.din(w_n74_0[1]));
	jspl3 jspl3_w_n75_0(.douta(w_n75_0[0]),.doutb(w_n75_0[1]),.doutc(w_dff_A_EhOeGe6S7_2),.din(n75));
	jspl3 jspl3_w_n75_1(.douta(w_n75_1[0]),.doutb(w_n75_1[1]),.doutc(w_n75_1[2]),.din(w_n75_0[0]));
	jspl jspl_w_n75_2(.douta(w_n75_2[0]),.doutb(w_n75_2[1]),.din(w_n75_0[1]));
	jspl jspl_w_n76_0(.douta(w_n76_0[0]),.doutb(w_n76_0[1]),.din(n76));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl3 jspl3_w_n79_0(.douta(w_n79_0[0]),.doutb(w_dff_A_yOUXbtIP7_1),.doutc(w_n79_0[2]),.din(n79));
	jspl3 jspl3_w_n79_1(.douta(w_dff_A_ObjgFuti1_0),.doutb(w_n79_1[1]),.doutc(w_dff_A_98rMngqj2_2),.din(w_n79_0[0]));
	jspl3 jspl3_w_n80_0(.douta(w_n80_0[0]),.doutb(w_dff_A_hIrgyG9Q4_1),.doutc(w_dff_A_nmcIZyGl1_2),.din(n80));
	jspl3 jspl3_w_n80_1(.douta(w_n80_1[0]),.doutb(w_n80_1[1]),.doutc(w_n80_1[2]),.din(w_n80_0[0]));
	jspl3 jspl3_w_n81_0(.douta(w_n81_0[0]),.doutb(w_n81_0[1]),.doutc(w_dff_A_VjANystY2_2),.din(n81));
	jspl3 jspl3_w_n81_1(.douta(w_dff_A_vevyfFaW1_0),.doutb(w_n81_1[1]),.doutc(w_n81_1[2]),.din(w_n81_0[0]));
	jspl jspl_w_n81_2(.douta(w_n81_2[0]),.doutb(w_n81_2[1]),.din(w_n81_0[1]));
	jspl3 jspl3_w_n84_0(.douta(w_n84_0[0]),.doutb(w_dff_A_c6nYiNQz8_1),.doutc(w_dff_A_oAkhjJVX7_2),.din(n84));
	jspl3 jspl3_w_n84_1(.douta(w_n84_1[0]),.doutb(w_n84_1[1]),.doutc(w_dff_A_Z1rKLJEN2_2),.din(w_n84_0[0]));
	jspl jspl_w_n85_0(.douta(w_n85_0[0]),.doutb(w_n85_0[1]),.din(n85));
	jspl3 jspl3_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.doutc(w_n86_0[2]),.din(n86));
	jspl jspl_w_n89_0(.douta(w_n89_0[0]),.doutb(w_n89_0[1]),.din(n89));
	jspl3 jspl3_w_n90_0(.douta(w_n90_0[0]),.doutb(w_n90_0[1]),.doutc(w_n90_0[2]),.din(n90));
	jspl3 jspl3_w_n91_0(.douta(w_n91_0[0]),.doutb(w_n91_0[1]),.doutc(w_n91_0[2]),.din(n91));
	jspl3 jspl3_w_n91_1(.douta(w_n91_1[0]),.doutb(w_n91_1[1]),.doutc(w_n91_1[2]),.din(w_n91_0[0]));
	jspl3 jspl3_w_n94_0(.douta(w_dff_A_9TorVuzk2_0),.doutb(w_n94_0[1]),.doutc(w_n94_0[2]),.din(n94));
	jspl3 jspl3_w_n96_0(.douta(w_n96_0[0]),.doutb(w_n96_0[1]),.doutc(w_n96_0[2]),.din(n96));
	jspl3 jspl3_w_n105_0(.douta(w_n105_0[0]),.doutb(w_dff_A_Ik8vCPxA0_1),.doutc(w_dff_A_55jDWv245_2),.din(n105));
	jspl jspl_w_n105_1(.douta(w_dff_A_5Bk3phfE6_0),.doutb(w_n105_1[1]),.din(w_n105_0[0]));
	jspl3 jspl3_w_n111_0(.douta(w_n111_0[0]),.doutb(w_n111_0[1]),.doutc(w_n111_0[2]),.din(n111));
	jspl jspl_w_n112_0(.douta(w_dff_A_l0vAzSjO1_0),.doutb(w_n112_0[1]),.din(n112));
	jspl3 jspl3_w_n118_0(.douta(w_n118_0[0]),.doutb(w_n118_0[1]),.doutc(w_n118_0[2]),.din(n118));
	jspl jspl_w_n120_0(.douta(w_n120_0[0]),.doutb(w_dff_A_UDU0rIU67_1),.din(n120));
	jspl jspl_w_n126_0(.douta(w_dff_A_S3wOPQv49_0),.doutb(w_n126_0[1]),.din(n126));
	jspl jspl_w_n130_0(.douta(w_n130_0[0]),.doutb(w_dff_A_sGUw0pmT6_1),.din(n130));
	jspl jspl_w_n134_0(.douta(w_n134_0[0]),.doutb(w_dff_A_acbnPoFk7_1),.din(n134));
	jspl jspl_w_n137_0(.douta(w_dff_A_kTfg7kte6_0),.doutb(w_n137_0[1]),.din(n137));
	jspl3 jspl3_w_n139_0(.douta(w_n139_0[0]),.doutb(w_n139_0[1]),.doutc(w_n139_0[2]),.din(n139));
	jspl3 jspl3_w_n139_1(.douta(w_dff_A_Nx08apME8_0),.doutb(w_n139_1[1]),.doutc(w_dff_A_cQeHUXR74_2),.din(w_n139_0[0]));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl3 jspl3_w_n141_0(.douta(w_n141_0[0]),.doutb(w_n141_0[1]),.doutc(w_n141_0[2]),.din(n141));
	jspl3 jspl3_w_n141_1(.douta(w_n141_1[0]),.doutb(w_dff_A_QfY9ycPs7_1),.doutc(w_dff_A_nNSVdi6V0_2),.din(w_n141_0[0]));
	jspl3 jspl3_w_n141_2(.douta(w_dff_A_zY3WHwLO9_0),.doutb(w_n141_2[1]),.doutc(w_n141_2[2]),.din(w_n141_0[1]));
	jspl jspl_w_n141_3(.douta(w_dff_A_Qu1KcUFZ3_0),.doutb(w_n141_3[1]),.din(w_n141_0[2]));
	jspl3 jspl3_w_n142_0(.douta(w_n142_0[0]),.doutb(w_n142_0[1]),.doutc(w_dff_A_BqhNtu9n3_2),.din(n142));
	jspl3 jspl3_w_n142_1(.douta(w_dff_A_lhYU8i2i5_0),.doutb(w_n142_1[1]),.doutc(w_n142_1[2]),.din(w_n142_0[0]));
	jspl jspl_w_n142_2(.douta(w_n142_2[0]),.doutb(w_n142_2[1]),.din(w_n142_0[1]));
	jspl jspl_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.din(n143));
	jspl3 jspl3_w_n144_0(.douta(w_n144_0[0]),.doutb(w_n144_0[1]),.doutc(w_n144_0[2]),.din(n144));
	jspl3 jspl3_w_n144_1(.douta(w_n144_1[0]),.doutb(w_n144_1[1]),.doutc(w_n144_1[2]),.din(w_n144_0[0]));
	jspl jspl_w_n144_2(.douta(w_n144_2[0]),.doutb(w_n144_2[1]),.din(w_n144_0[1]));
	jspl3 jspl3_w_n147_0(.douta(w_n147_0[0]),.doutb(w_n147_0[1]),.doutc(w_n147_0[2]),.din(n147));
	jspl jspl_w_n148_0(.douta(w_n148_0[0]),.doutb(w_n148_0[1]),.din(n148));
	jspl3 jspl3_w_n151_0(.douta(w_n151_0[0]),.doutb(w_n151_0[1]),.doutc(w_n151_0[2]),.din(n151));
	jspl3 jspl3_w_n151_1(.douta(w_n151_1[0]),.doutb(w_dff_A_wFaGRlsO1_1),.doutc(w_dff_A_kKS7HTiK1_2),.din(w_n151_0[0]));
	jspl3 jspl3_w_n151_2(.douta(w_dff_A_QqWgiOB68_0),.doutb(w_n151_2[1]),.doutc(w_dff_A_shuBNnAO4_2),.din(w_n151_0[1]));
	jspl3 jspl3_w_n151_3(.douta(w_n151_3[0]),.doutb(w_n151_3[1]),.doutc(w_dff_A_8lVb8cug4_2),.din(w_n151_0[2]));
	jspl3 jspl3_w_n151_4(.douta(w_n151_4[0]),.doutb(w_dff_A_fGufZ8pH1_1),.doutc(w_n151_4[2]),.din(w_n151_1[0]));
	jspl3 jspl3_w_n151_5(.douta(w_dff_A_tbzq0ca04_0),.doutb(w_n151_5[1]),.doutc(w_n151_5[2]),.din(w_n151_1[1]));
	jspl jspl_w_n151_6(.douta(w_dff_A_Q5xQh3CZ8_0),.doutb(w_n151_6[1]),.din(w_n151_1[2]));
	jspl3 jspl3_w_n152_0(.douta(w_dff_A_3QeCQqy86_0),.doutb(w_n152_0[1]),.doutc(w_dff_A_dfW7T59s0_2),.din(n152));
	jspl3 jspl3_w_n153_0(.douta(w_n153_0[0]),.doutb(w_n153_0[1]),.doutc(w_dff_A_xZyeqGsy9_2),.din(n153));
	jspl3 jspl3_w_n153_1(.douta(w_dff_A_vePoAHTu0_0),.doutb(w_n153_1[1]),.doutc(w_n153_1[2]),.din(w_n153_0[0]));
	jspl3 jspl3_w_n153_2(.douta(w_n153_2[0]),.doutb(w_n153_2[1]),.doutc(w_dff_A_dZWH8cyL6_2),.din(w_n153_0[1]));
	jspl3 jspl3_w_n153_3(.douta(w_n153_3[0]),.doutb(w_dff_A_EjlM9Hnm1_1),.doutc(w_dff_A_V4Oy8Dsb1_2),.din(w_n153_0[2]));
	jspl3 jspl3_w_n153_4(.douta(w_dff_A_PMwywllJ0_0),.doutb(w_dff_A_z7nYyzmH2_1),.doutc(w_n153_4[2]),.din(w_n153_1[0]));
	jspl3 jspl3_w_n153_5(.douta(w_dff_A_BrvxRotp4_0),.doutb(w_n153_5[1]),.doutc(w_n153_5[2]),.din(w_n153_1[1]));
	jspl3 jspl3_w_n153_6(.douta(w_n153_6[0]),.doutb(w_n153_6[1]),.doutc(w_n153_6[2]),.din(w_n153_1[2]));
	jspl3 jspl3_w_n153_7(.douta(w_n153_7[0]),.doutb(w_n153_7[1]),.doutc(w_n153_7[2]),.din(w_n153_2[0]));
	jspl jspl_w_n153_8(.douta(w_n153_8[0]),.doutb(w_n153_8[1]),.din(w_n153_2[1]));
	jspl3 jspl3_w_n161_0(.douta(w_n161_0[0]),.doutb(w_dff_A_Kmx4IvMP5_1),.doutc(w_n161_0[2]),.din(n161));
	jspl3 jspl3_w_n163_0(.douta(w_n163_0[0]),.doutb(w_dff_A_PB3oHri44_1),.doutc(w_dff_A_7HilQhhT0_2),.din(n163));
	jspl jspl_w_n163_1(.douta(w_n163_1[0]),.doutb(w_dff_A_EwrqlWyp2_1),.din(w_n163_0[0]));
	jspl3 jspl3_w_n164_0(.douta(w_n164_0[0]),.doutb(w_n164_0[1]),.doutc(w_n164_0[2]),.din(n164));
	jspl jspl_w_n165_0(.douta(w_n165_0[0]),.doutb(w_dff_A_QCW8hcPI2_1),.din(n165));
	jspl jspl_w_n167_0(.douta(w_n167_0[0]),.doutb(w_dff_A_QPcPdCI90_1),.din(n167));
	jspl3 jspl3_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.doutc(w_n168_0[2]),.din(n168));
	jspl3 jspl3_w_n168_1(.douta(w_n168_1[0]),.doutb(w_n168_1[1]),.doutc(w_n168_1[2]),.din(w_n168_0[0]));
	jspl3 jspl3_w_n168_2(.douta(w_dff_A_IfVgLIMX6_0),.doutb(w_n168_2[1]),.doutc(w_n168_2[2]),.din(w_n168_0[1]));
	jspl3 jspl3_w_n168_3(.douta(w_dff_A_Ae8V3D2h6_0),.doutb(w_n168_3[1]),.doutc(w_dff_A_ibTsKWpo0_2),.din(w_n168_0[2]));
	jspl3 jspl3_w_n168_4(.douta(w_dff_A_TIDzhtUv3_0),.doutb(w_dff_A_J55No7Ox2_1),.doutc(w_n168_4[2]),.din(w_n168_1[0]));
	jspl jspl_w_n168_5(.douta(w_n168_5[0]),.doutb(w_n168_5[1]),.din(w_n168_1[1]));
	jspl jspl_w_n169_0(.douta(w_n169_0[0]),.doutb(w_n169_0[1]),.din(n169));
	jspl3 jspl3_w_n170_0(.douta(w_n170_0[0]),.doutb(w_n170_0[1]),.doutc(w_dff_A_b1EAzkv06_2),.din(w_dff_B_WnJKDA8q3_3));
	jspl3 jspl3_w_n172_0(.douta(w_n172_0[0]),.doutb(w_dff_A_IxbcIBxm6_1),.doutc(w_dff_A_hSgxQEJA9_2),.din(n172));
	jspl3 jspl3_w_n172_1(.douta(w_n172_1[0]),.doutb(w_dff_A_7tTiqfhT6_1),.doutc(w_dff_A_3AAwax0a6_2),.din(w_n172_0[0]));
	jspl3 jspl3_w_n172_2(.douta(w_n172_2[0]),.doutb(w_n172_2[1]),.doutc(w_n172_2[2]),.din(w_n172_0[1]));
	jspl3 jspl3_w_n172_3(.douta(w_n172_3[0]),.doutb(w_n172_3[1]),.doutc(w_n172_3[2]),.din(w_n172_0[2]));
	jspl3 jspl3_w_n172_4(.douta(w_n172_4[0]),.doutb(w_dff_A_vga5hyTG0_1),.doutc(w_dff_A_nvMEuQpG9_2),.din(w_n172_1[0]));
	jspl3 jspl3_w_n173_0(.douta(w_n173_0[0]),.doutb(w_n173_0[1]),.doutc(w_n173_0[2]),.din(n173));
	jspl3 jspl3_w_n173_1(.douta(w_n173_1[0]),.doutb(w_n173_1[1]),.doutc(w_n173_1[2]),.din(w_n173_0[0]));
	jspl3 jspl3_w_n173_2(.douta(w_n173_2[0]),.doutb(w_n173_2[1]),.doutc(w_n173_2[2]),.din(w_n173_0[1]));
	jspl jspl_w_n173_3(.douta(w_n173_3[0]),.doutb(w_n173_3[1]),.din(w_n173_0[2]));
	jspl jspl_w_n176_0(.douta(w_n176_0[0]),.doutb(w_n176_0[1]),.din(n176));
	jspl3 jspl3_w_n177_0(.douta(w_n177_0[0]),.doutb(w_n177_0[1]),.doutc(w_n177_0[2]),.din(n177));
	jspl3 jspl3_w_n177_1(.douta(w_n177_1[0]),.doutb(w_n177_1[1]),.doutc(w_n177_1[2]),.din(w_n177_0[0]));
	jspl3 jspl3_w_n182_0(.douta(w_n182_0[0]),.doutb(w_n182_0[1]),.doutc(w_n182_0[2]),.din(n182));
	jspl jspl_w_n182_1(.douta(w_n182_1[0]),.doutb(w_n182_1[1]),.din(w_n182_0[0]));
	jspl3 jspl3_w_n186_0(.douta(w_n186_0[0]),.doutb(w_dff_A_g9nn8Zc14_1),.doutc(w_n186_0[2]),.din(n186));
	jspl3 jspl3_w_n186_1(.douta(w_n186_1[0]),.doutb(w_n186_1[1]),.doutc(w_n186_1[2]),.din(w_n186_0[0]));
	jspl3 jspl3_w_n189_0(.douta(w_dff_A_b53XyEOm5_0),.doutb(w_dff_A_OGcwN2MC2_1),.doutc(w_n189_0[2]),.din(n189));
	jspl3 jspl3_w_n189_1(.douta(w_n189_1[0]),.doutb(w_dff_A_7dtRq2NS9_1),.doutc(w_n189_1[2]),.din(w_n189_0[0]));
	jspl3 jspl3_w_n189_2(.douta(w_n189_2[0]),.doutb(w_dff_A_ZN1HbWSE0_1),.doutc(w_dff_A_WxnTA56b3_2),.din(w_n189_0[1]));
	jspl jspl_w_n190_0(.douta(w_n190_0[0]),.doutb(w_dff_A_A6Ofxp4u6_1),.din(n190));
	jspl3 jspl3_w_n192_0(.douta(w_n192_0[0]),.doutb(w_dff_A_KNfRQKVM6_1),.doutc(w_n192_0[2]),.din(n192));
	jspl3 jspl3_w_n198_0(.douta(w_n198_0[0]),.doutb(w_n198_0[1]),.doutc(w_dff_A_bnC8QV0j7_2),.din(n198));
	jspl3 jspl3_w_n199_0(.douta(w_dff_A_b8n47nWS4_0),.doutb(w_n199_0[1]),.doutc(w_dff_A_GRRwwvD30_2),.din(w_dff_B_KU0nt64i4_3));
	jspl jspl_w_n201_0(.douta(w_n201_0[0]),.doutb(w_dff_A_nANvYK136_1),.din(n201));
	jspl jspl_w_n202_0(.douta(w_n202_0[0]),.doutb(w_dff_A_WdejfyvY0_1),.din(n202));
	jspl3 jspl3_w_n205_0(.douta(w_n205_0[0]),.doutb(w_n205_0[1]),.doutc(w_n205_0[2]),.din(n205));
	jspl jspl_w_n205_1(.douta(w_n205_1[0]),.doutb(w_n205_1[1]),.din(w_n205_0[0]));
	jspl jspl_w_n207_0(.douta(w_dff_A_REIo9ffo7_0),.doutb(w_n207_0[1]),.din(n207));
	jspl3 jspl3_w_n212_0(.douta(w_n212_0[0]),.doutb(w_dff_A_bRRjJPyT6_1),.doutc(w_n212_0[2]),.din(n212));
	jspl jspl_w_n212_1(.douta(w_n212_1[0]),.doutb(w_n212_1[1]),.din(w_n212_0[0]));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_dff_A_UYDQdNuH7_1),.din(n213));
	jspl jspl_w_n215_0(.douta(w_n215_0[0]),.doutb(w_n215_0[1]),.din(n215));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_dff_A_qAdhCfa83_1),.din(n218));
	jspl3 jspl3_w_n224_0(.douta(w_n224_0[0]),.doutb(w_n224_0[1]),.doutc(w_dff_A_MDqOfozP8_2),.din(n224));
	jspl jspl_w_n224_1(.douta(w_dff_A_OlooEsLk1_0),.doutb(w_n224_1[1]),.din(w_n224_0[0]));
	jspl jspl_w_n225_0(.douta(w_n225_0[0]),.doutb(w_n225_0[1]),.din(n225));
	jspl jspl_w_n229_0(.douta(w_n229_0[0]),.doutb(w_dff_A_5HXFfcAo9_1),.din(n229));
	jspl3 jspl3_w_n234_0(.douta(w_n234_0[0]),.doutb(w_dff_A_2WoCuG5J3_1),.doutc(w_n234_0[2]),.din(n234));
	jspl jspl_w_n234_1(.douta(w_n234_1[0]),.doutb(w_n234_1[1]),.din(w_n234_0[0]));
	jspl3 jspl3_w_n237_0(.douta(w_n237_0[0]),.doutb(w_dff_A_9a3Em77c0_1),.doutc(w_n237_0[2]),.din(n237));
	jspl jspl_w_n238_0(.douta(w_n238_0[0]),.doutb(w_dff_A_1279TGH46_1),.din(n238));
	jspl3 jspl3_w_n242_0(.douta(w_n242_0[0]),.doutb(w_dff_A_ZMKhAMUR0_1),.doutc(w_dff_A_HDWYnpOB9_2),.din(n242));
	jspl jspl_w_n243_0(.douta(w_dff_A_YcSEk4u81_0),.doutb(w_n243_0[1]),.din(n243));
	jspl jspl_w_n247_0(.douta(w_n247_0[0]),.doutb(w_dff_A_93Zd3l2g8_1),.din(n247));
	jspl jspl_w_n250_0(.douta(w_n250_0[0]),.doutb(w_dff_A_UjEXtY9A0_1),.din(n250));
	jspl jspl_w_n251_0(.douta(w_dff_A_HOhlGm5x4_0),.doutb(w_n251_0[1]),.din(n251));
	jspl3 jspl3_w_n255_0(.douta(w_n255_0[0]),.doutb(w_n255_0[1]),.doutc(w_n255_0[2]),.din(n255));
	jspl jspl_w_n255_1(.douta(w_n255_1[0]),.doutb(w_n255_1[1]),.din(w_n255_0[0]));
	jspl jspl_w_n256_0(.douta(w_n256_0[0]),.doutb(w_dff_A_U3CmrLaq8_1),.din(n256));
	jspl jspl_w_n257_0(.douta(w_n257_0[0]),.doutb(w_dff_A_h7ftODI60_1),.din(n257));
	jspl jspl_w_n259_0(.douta(w_n259_0[0]),.doutb(w_n259_0[1]),.din(n259));
	jspl jspl_w_n260_0(.douta(w_n260_0[0]),.doutb(w_dff_A_EgbFodsF6_1),.din(n260));
	jspl3 jspl3_w_n261_0(.douta(w_n261_0[0]),.doutb(w_dff_A_QrqwqCbg4_1),.doutc(w_dff_A_k0Hrm9on7_2),.din(n261));
	jspl3 jspl3_w_n261_1(.douta(w_n261_1[0]),.doutb(w_n261_1[1]),.doutc(w_n261_1[2]),.din(w_n261_0[0]));
	jspl3 jspl3_w_n262_0(.douta(w_dff_A_PhnE6QKk6_0),.doutb(w_dff_A_gsERAYf14_1),.doutc(w_n262_0[2]),.din(n262));
	jspl jspl_w_n269_0(.douta(w_dff_A_us0AcsJW6_0),.doutb(w_n269_0[1]),.din(n269));
	jspl jspl_w_n272_0(.douta(w_n272_0[0]),.doutb(w_n272_0[1]),.din(n272));
	jspl3 jspl3_w_n279_0(.douta(w_n279_0[0]),.doutb(w_n279_0[1]),.doutc(w_n279_0[2]),.din(n279));
	jspl jspl_w_n279_1(.douta(w_n279_1[0]),.doutb(w_n279_1[1]),.din(w_n279_0[0]));
	jspl jspl_w_n282_0(.douta(w_dff_A_yrHzOZpB0_0),.doutb(w_n282_0[1]),.din(n282));
	jspl jspl_w_n283_0(.douta(w_n283_0[0]),.doutb(w_dff_A_1YteJ72n8_1),.din(n283));
	jspl3 jspl3_w_n292_0(.douta(w_n292_0[0]),.doutb(w_n292_0[1]),.doutc(w_n292_0[2]),.din(n292));
	jspl jspl_w_n298_0(.douta(w_dff_A_VRn3UZHx9_0),.doutb(w_n298_0[1]),.din(n298));
	jspl3 jspl3_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.doutc(w_n308_0[2]),.din(n308));
	jspl3 jspl3_w_n308_1(.douta(w_n308_1[0]),.doutb(w_n308_1[1]),.doutc(w_n308_1[2]),.din(w_n308_0[0]));
	jspl jspl_w_n309_0(.douta(w_n309_0[0]),.doutb(w_dff_A_66o4pQgu8_1),.din(n309));
	jspl jspl_w_n310_0(.douta(w_dff_A_v2s6uZoF7_0),.doutb(w_n310_0[1]),.din(n310));
	jspl jspl_w_n312_0(.douta(w_dff_A_bXF8Ko468_0),.doutb(w_n312_0[1]),.din(n312));
	jspl jspl_w_n313_0(.douta(w_dff_A_eHGMUOgQ9_0),.doutb(w_n313_0[1]),.din(n313));
	jspl3 jspl3_w_n315_0(.douta(w_dff_A_JSngJh1o7_0),.doutb(w_n315_0[1]),.doutc(w_dff_A_aUuFFNoZ0_2),.din(n315));
	jspl jspl_w_n321_0(.douta(w_n321_0[0]),.doutb(w_dff_A_JD62UApS0_1),.din(n321));
	jspl3 jspl3_w_n323_0(.douta(w_n323_0[0]),.doutb(w_dff_A_SG9uoOXf1_1),.doutc(w_dff_A_rDmAkkS04_2),.din(n323));
	jspl3 jspl3_w_n330_0(.douta(w_n330_0[0]),.doutb(w_n330_0[1]),.doutc(w_n330_0[2]),.din(n330));
	jspl jspl_w_n333_0(.douta(w_dff_A_6VGMMbyj4_0),.doutb(w_n333_0[1]),.din(n333));
	jspl jspl_w_n334_0(.douta(w_dff_A_xSMk7Iu53_0),.doutb(w_n334_0[1]),.din(n334));
	jspl jspl_w_n344_0(.douta(w_n344_0[0]),.doutb(w_n344_0[1]),.din(n344));
	jspl jspl_w_n347_0(.douta(w_n347_0[0]),.doutb(w_dff_A_25sVWHOy3_1),.din(n347));
	jspl jspl_w_n348_0(.douta(w_dff_A_lFUaObDu7_0),.doutb(w_n348_0[1]),.din(n348));
	jspl jspl_w_n349_0(.douta(w_n349_0[0]),.doutb(w_n349_0[1]),.din(n349));
	jspl jspl_w_n350_0(.douta(w_n350_0[0]),.doutb(w_n350_0[1]),.din(n350));
	jspl jspl_w_n351_0(.douta(w_n351_0[0]),.doutb(w_dff_A_5vTYak7O9_1),.din(n351));
	jspl3 jspl3_w_n352_0(.douta(w_n352_0[0]),.doutb(w_dff_A_6yFqqlZp9_1),.doutc(w_dff_A_h72eUwTZ4_2),.din(n352));
	jspl jspl_w_n352_1(.douta(w_dff_A_VxkHbEoJ1_0),.doutb(w_n352_1[1]),.din(w_n352_0[0]));
	jspl3 jspl3_w_n354_0(.douta(w_n354_0[0]),.doutb(w_dff_A_5gjoHNAA6_1),.doutc(w_dff_A_knkxMSEg2_2),.din(n354));
	jspl jspl_w_n354_1(.douta(w_dff_A_o0jD4GnU1_0),.doutb(w_n354_1[1]),.din(w_n354_0[0]));
	jspl jspl_w_n355_0(.douta(w_n355_0[0]),.doutb(w_n355_0[1]),.din(n355));
	jspl3 jspl3_w_n356_0(.douta(w_n356_0[0]),.doutb(w_dff_A_s56N452h0_1),.doutc(w_dff_A_2v5adAyr4_2),.din(n356));
	jspl jspl_w_n356_1(.douta(w_dff_A_UjOJvMcG4_0),.doutb(w_n356_1[1]),.din(w_n356_0[0]));
	jspl jspl_w_n357_0(.douta(w_n357_0[0]),.doutb(w_dff_A_r1xFQf2C4_1),.din(n357));
	jspl3 jspl3_w_n367_0(.douta(w_n367_0[0]),.doutb(w_n367_0[1]),.doutc(w_n367_0[2]),.din(n367));
	jspl jspl_w_n367_1(.douta(w_n367_1[0]),.doutb(w_n367_1[1]),.din(w_n367_0[0]));
	jspl jspl_w_n370_0(.douta(w_dff_A_AzQ9Rfkm7_0),.doutb(w_n370_0[1]),.din(w_dff_B_shsYs3545_2));
	jspl jspl_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.din(n375));
	jspl jspl_w_n378_0(.douta(w_dff_A_UZUteTL87_0),.doutb(w_n378_0[1]),.din(n378));
	jspl3 jspl3_w_n383_0(.douta(w_n383_0[0]),.doutb(w_dff_A_EilZvoQR7_1),.doutc(w_n383_0[2]),.din(n383));
	jspl3 jspl3_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.doutc(w_n387_0[2]),.din(n387));
	jspl3 jspl3_w_n388_0(.douta(w_dff_A_ivs22P1q2_0),.doutb(w_dff_A_GaxknGMP0_1),.doutc(w_n388_0[2]),.din(n388));
	jspl3 jspl3_w_n388_1(.douta(w_n388_1[0]),.doutb(w_dff_A_O7ejGNVk3_1),.doutc(w_dff_A_upzh20eh1_2),.din(w_n388_0[0]));
	jspl jspl_w_n388_2(.douta(w_n388_2[0]),.doutb(w_dff_A_oNuluRoW1_1),.din(w_n388_0[1]));
	jspl jspl_w_n394_0(.douta(w_n394_0[0]),.doutb(w_n394_0[1]),.din(n394));
	jspl jspl_w_n395_0(.douta(w_dff_A_aPNn3EpD9_0),.doutb(w_n395_0[1]),.din(n395));
	jspl3 jspl3_w_n404_0(.douta(w_n404_0[0]),.doutb(w_n404_0[1]),.doutc(w_n404_0[2]),.din(n404));
	jspl jspl_w_n405_0(.douta(w_n405_0[0]),.doutb(w_n405_0[1]),.din(n405));
	jspl jspl_w_n407_0(.douta(w_n407_0[0]),.doutb(w_dff_A_Td2GGZBJ4_1),.din(n407));
	jspl3 jspl3_w_n414_0(.douta(w_n414_0[0]),.doutb(w_n414_0[1]),.doutc(w_n414_0[2]),.din(n414));
	jspl3 jspl3_w_n417_0(.douta(w_n417_0[0]),.doutb(w_dff_A_Xi4JRTa49_1),.doutc(w_dff_A_vcxg1qYh8_2),.din(n417));
	jspl jspl_w_n420_0(.douta(w_n420_0[0]),.doutb(w_dff_A_T8uo1aQq5_1),.din(n420));
	jspl jspl_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.din(n425));
	jspl jspl_w_n426_0(.douta(w_n426_0[0]),.doutb(w_n426_0[1]),.din(n426));
	jspl jspl_w_n428_0(.douta(w_dff_A_RFNPLB650_0),.doutb(w_n428_0[1]),.din(n428));
	jspl jspl_w_n430_0(.douta(w_dff_A_c23foJsE2_0),.doutb(w_n430_0[1]),.din(n430));
	jspl jspl_w_n435_0(.douta(w_n435_0[0]),.doutb(w_dff_A_b7shwyO36_1),.din(n435));
	jspl3 jspl3_w_n439_0(.douta(w_n439_0[0]),.doutb(w_n439_0[1]),.doutc(w_n439_0[2]),.din(n439));
	jspl jspl_w_n441_0(.douta(w_n441_0[0]),.doutb(w_n441_0[1]),.din(n441));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl jspl_w_n450_0(.douta(w_dff_A_NCw5ISe29_0),.doutb(w_n450_0[1]),.din(n450));
	jspl jspl_w_n452_0(.douta(w_n452_0[0]),.doutb(w_n452_0[1]),.din(n452));
	jspl jspl_w_n456_0(.douta(w_n456_0[0]),.doutb(w_dff_A_Ydbojq200_1),.din(n456));
	jspl jspl_w_n457_0(.douta(w_n457_0[0]),.doutb(w_n457_0[1]),.din(n457));
	jspl jspl_w_n465_0(.douta(w_n465_0[0]),.doutb(w_n465_0[1]),.din(n465));
	jspl jspl_w_n472_0(.douta(w_n472_0[0]),.doutb(w_n472_0[1]),.din(n472));
	jspl jspl_w_n473_0(.douta(w_n473_0[0]),.doutb(w_n473_0[1]),.din(n473));
	jspl3 jspl3_w_n482_0(.douta(w_n482_0[0]),.doutb(w_n482_0[1]),.doutc(w_n482_0[2]),.din(n482));
	jspl jspl_w_n483_0(.douta(w_n483_0[0]),.doutb(w_n483_0[1]),.din(n483));
	jspl jspl_w_n494_0(.douta(w_dff_A_3GyNeKS69_0),.doutb(w_n494_0[1]),.din(n494));
	jspl jspl_w_n499_0(.douta(w_n499_0[0]),.doutb(w_dff_A_HCXleRxp7_1),.din(n499));
	jspl jspl_w_n500_0(.douta(w_n500_0[0]),.doutb(w_n500_0[1]),.din(n500));
	jspl3 jspl3_w_n503_0(.douta(w_n503_0[0]),.doutb(w_dff_A_DNdT5Ak99_1),.doutc(w_n503_0[2]),.din(n503));
	jspl3 jspl3_w_n507_0(.douta(w_n507_0[0]),.doutb(w_dff_A_M1oOOEom0_1),.doutc(w_dff_A_Sy4bVevd0_2),.din(n507));
	jspl3 jspl3_w_n507_1(.douta(w_dff_A_LNiO5wDO0_0),.doutb(w_dff_A_dBe52Yhh4_1),.doutc(w_n507_1[2]),.din(w_n507_0[0]));
	jspl jspl_w_n507_2(.douta(w_n507_2[0]),.doutb(w_dff_A_uDbIhnhQ0_1),.din(w_n507_0[1]));
	jspl jspl_w_n511_0(.douta(w_n511_0[0]),.doutb(w_n511_0[1]),.din(n511));
	jspl jspl_w_n512_0(.douta(w_dff_A_iTgn9Xz62_0),.doutb(w_n512_0[1]),.din(n512));
	jspl3 jspl3_w_n514_0(.douta(w_n514_0[0]),.doutb(w_dff_A_hhoYO9hg9_1),.doutc(w_dff_A_v1McfurO5_2),.din(n514));
	jspl jspl_w_n514_1(.douta(w_dff_A_MvoiZR3U7_0),.doutb(w_n514_1[1]),.din(w_n514_0[0]));
	jspl jspl_w_n520_0(.douta(w_dff_A_Q2LPEikI5_0),.doutb(w_n520_0[1]),.din(n520));
	jspl jspl_w_n533_0(.douta(w_n533_0[0]),.doutb(w_n533_0[1]),.din(n533));
	jspl jspl_w_n534_0(.douta(w_n534_0[0]),.doutb(w_dff_A_r7coMN1H0_1),.din(n534));
	jspl jspl_w_n541_0(.douta(w_n541_0[0]),.doutb(w_n541_0[1]),.din(n541));
	jspl jspl_w_n542_0(.douta(w_n542_0[0]),.doutb(w_n542_0[1]),.din(n542));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_n543_0[1]),.din(n543));
	jspl jspl_w_n544_0(.douta(w_n544_0[0]),.doutb(w_n544_0[1]),.din(n544));
	jspl jspl_w_n548_0(.douta(w_n548_0[0]),.doutb(w_dff_A_uiIIcp3f6_1),.din(n548));
	jspl jspl_w_n550_0(.douta(w_n550_0[0]),.doutb(w_n550_0[1]),.din(n550));
	jspl jspl_w_n551_0(.douta(w_n551_0[0]),.doutb(w_n551_0[1]),.din(n551));
	jspl jspl_w_n559_0(.douta(w_n559_0[0]),.doutb(w_n559_0[1]),.din(n559));
	jspl jspl_w_n562_0(.douta(w_dff_A_FRkws6Vl4_0),.doutb(w_n562_0[1]),.din(n562));
	jspl3 jspl3_w_n566_0(.douta(w_n566_0[0]),.doutb(w_dff_A_SaBZhgma6_1),.doutc(w_dff_A_a77PsJUx4_2),.din(n566));
	jspl jspl_w_n566_1(.douta(w_n566_1[0]),.doutb(w_n566_1[1]),.din(w_n566_0[0]));
	jspl3 jspl3_w_n567_0(.douta(w_n567_0[0]),.doutb(w_dff_A_nulbQinz5_1),.doutc(w_dff_A_ZmqweskX2_2),.din(n567));
	jspl3 jspl3_w_n567_1(.douta(w_dff_A_hLHVdNtW3_0),.doutb(w_n567_1[1]),.doutc(w_dff_A_SebHfa9a5_2),.din(w_n567_0[0]));
	jspl3 jspl3_w_n567_2(.douta(w_n567_2[0]),.doutb(w_n567_2[1]),.doutc(w_dff_A_BcrQTTm06_2),.din(w_n567_0[1]));
	jspl3 jspl3_w_n567_3(.douta(w_dff_A_c60IsobB1_0),.doutb(w_dff_A_ZRods4mx6_1),.doutc(w_n567_3[2]),.din(w_n567_0[2]));
	jspl3 jspl3_w_n567_4(.douta(w_dff_A_Zs0Q64kA6_0),.doutb(w_n567_4[1]),.doutc(w_n567_4[2]),.din(w_n567_1[0]));
	jspl jspl_w_n567_5(.douta(w_n567_5[0]),.doutb(w_dff_A_ogos4tL26_1),.din(w_n567_1[1]));
	jspl jspl_w_n569_0(.douta(w_n569_0[0]),.doutb(w_dff_A_7Mu1Dhco8_1),.din(n569));
	jspl jspl_w_n570_0(.douta(w_dff_A_Me1fhYuZ2_0),.doutb(w_n570_0[1]),.din(n570));
	jspl3 jspl3_w_n571_0(.douta(w_n571_0[0]),.doutb(w_dff_A_eM79DCKB4_1),.doutc(w_dff_A_Jz9hUAx84_2),.din(w_dff_B_kxKU4Zyf9_3));
	jspl3 jspl3_w_n571_1(.douta(w_n571_1[0]),.doutb(w_dff_A_i4C8CJMS1_1),.doutc(w_n571_1[2]),.din(w_n571_0[0]));
	jspl jspl_w_n571_2(.douta(w_dff_A_iQuhWqzD7_0),.doutb(w_n571_2[1]),.din(w_n571_0[1]));
	jspl3 jspl3_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.doutc(w_n572_0[2]),.din(n572));
	jspl jspl_w_n573_0(.douta(w_n573_0[0]),.doutb(w_n573_0[1]),.din(n573));
	jspl jspl_w_n574_0(.douta(w_n574_0[0]),.doutb(w_n574_0[1]),.din(n574));
	jspl3 jspl3_w_n576_0(.douta(w_n576_0[0]),.doutb(w_n576_0[1]),.doutc(w_n576_0[2]),.din(n576));
	jspl jspl_w_n577_0(.douta(w_dff_A_C61XykJj3_0),.doutb(w_n577_0[1]),.din(n577));
	jspl3 jspl3_w_n579_0(.douta(w_n579_0[0]),.doutb(w_n579_0[1]),.doutc(w_dff_A_9bQoZvaZ9_2),.din(n579));
	jspl jspl_w_n579_1(.douta(w_n579_1[0]),.doutb(w_dff_A_nnTQgwfk1_1),.din(w_n579_0[0]));
	jspl3 jspl3_w_n580_0(.douta(w_n580_0[0]),.doutb(w_n580_0[1]),.doutc(w_n580_0[2]),.din(n580));
	jspl jspl_w_n582_0(.douta(w_n582_0[0]),.doutb(w_n582_0[1]),.din(n582));
	jspl jspl_w_n584_0(.douta(w_n584_0[0]),.doutb(w_n584_0[1]),.din(n584));
	jspl jspl_w_n598_0(.douta(w_dff_A_qiJW42G68_0),.doutb(w_n598_0[1]),.din(n598));
	jspl3 jspl3_w_n600_0(.douta(w_n600_0[0]),.doutb(w_n600_0[1]),.doutc(w_n600_0[2]),.din(n600));
	jspl3 jspl3_w_n600_1(.douta(w_dff_A_mG4NQv9y8_0),.doutb(w_dff_A_AD8s80ZX9_1),.doutc(w_n600_1[2]),.din(w_n600_0[0]));
	jspl3 jspl3_w_n601_0(.douta(w_n601_0[0]),.doutb(w_dff_A_1JsX1pGC1_1),.doutc(w_n601_0[2]),.din(n601));
	jspl jspl_w_n602_0(.douta(w_n602_0[0]),.doutb(w_n602_0[1]),.din(n602));
	jspl3 jspl3_w_n604_0(.douta(w_dff_A_wO4aJOgl9_0),.doutb(w_n604_0[1]),.doutc(w_dff_A_WIx6MBO00_2),.din(n604));
	jspl3 jspl3_w_n604_1(.douta(w_dff_A_LsbrMTkE4_0),.doutb(w_dff_A_WxdUJPLt4_1),.doutc(w_n604_1[2]),.din(w_n604_0[0]));
	jspl3 jspl3_w_n604_2(.douta(w_dff_A_R9Tb3AaW0_0),.doutb(w_n604_2[1]),.doutc(w_n604_2[2]),.din(w_n604_0[1]));
	jspl3 jspl3_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.doutc(w_n605_0[2]),.din(n605));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_dff_A_PZ0LGSYx0_1),.doutc(w_dff_A_4pvAQzxU1_2),.din(w_dff_B_1Lv68ur21_3));
	jspl3 jspl3_w_n613_1(.douta(w_dff_A_wfZHBpMz4_0),.doutb(w_dff_A_MagKJvnV4_1),.doutc(w_n613_1[2]),.din(w_n613_0[0]));
	jspl3 jspl3_w_n614_0(.douta(w_n614_0[0]),.doutb(w_dff_A_hdzvul4H2_1),.doutc(w_dff_A_DLFXdhd73_2),.din(n614));
	jspl3 jspl3_w_n614_1(.douta(w_dff_A_Sl5uowRH7_0),.doutb(w_n614_1[1]),.doutc(w_dff_A_I9tN8kjN3_2),.din(w_n614_0[0]));
	jspl3 jspl3_w_n614_2(.douta(w_dff_A_dLJ03ZvW5_0),.doutb(w_dff_A_POL1wn4v6_1),.doutc(w_n614_2[2]),.din(w_n614_0[1]));
	jspl3 jspl3_w_n614_3(.douta(w_n614_3[0]),.doutb(w_dff_A_VRH3paYD6_1),.doutc(w_dff_A_3NM5qXvP7_2),.din(w_n614_0[2]));
	jspl3 jspl3_w_n614_4(.douta(w_n614_4[0]),.doutb(w_dff_A_HfBoGHCo1_1),.doutc(w_dff_A_oZO6c03a0_2),.din(w_n614_1[0]));
	jspl jspl_w_n614_5(.douta(w_dff_A_F3IObSgd7_0),.doutb(w_n614_5[1]),.din(w_n614_1[1]));
	jspl3 jspl3_w_n618_0(.douta(w_n618_0[0]),.doutb(w_n618_0[1]),.doutc(w_dff_A_leBPYbM77_2),.din(n618));
	jspl3 jspl3_w_n618_1(.douta(w_dff_A_ocxPA7mX1_0),.doutb(w_dff_A_1psSUxf49_1),.doutc(w_n618_1[2]),.din(w_n618_0[0]));
	jspl jspl_w_n618_2(.douta(w_dff_A_TOm96VmT0_0),.doutb(w_n618_2[1]),.din(w_n618_0[1]));
	jspl3 jspl3_w_n619_0(.douta(w_dff_A_kItzOBoR2_0),.doutb(w_dff_A_N9SE4bwk6_1),.doutc(w_n619_0[2]),.din(n619));
	jspl3 jspl3_w_n620_0(.douta(w_dff_A_LxUlK06f0_0),.doutb(w_n620_0[1]),.doutc(w_dff_A_9HYA86y12_2),.din(n620));
	jspl jspl_w_n622_0(.douta(w_dff_A_IGkdb4hj6_0),.doutb(w_n622_0[1]),.din(n622));
	jspl jspl_w_n624_0(.douta(w_n624_0[0]),.doutb(w_n624_0[1]),.din(n624));
	jspl3 jspl3_w_n626_0(.douta(w_n626_0[0]),.doutb(w_n626_0[1]),.doutc(w_n626_0[2]),.din(n626));
	jspl jspl_w_n628_0(.douta(w_n628_0[0]),.doutb(w_n628_0[1]),.din(n628));
	jspl3 jspl3_w_n629_0(.douta(w_n629_0[0]),.doutb(w_n629_0[1]),.doutc(w_n629_0[2]),.din(n629));
	jspl3 jspl3_w_n629_1(.douta(w_n629_1[0]),.doutb(w_n629_1[1]),.doutc(w_n629_1[2]),.din(w_n629_0[0]));
	jspl3 jspl3_w_n629_2(.douta(w_n629_2[0]),.doutb(w_n629_2[1]),.doutc(w_n629_2[2]),.din(w_n629_0[1]));
	jspl3 jspl3_w_n629_3(.douta(w_n629_3[0]),.doutb(w_n629_3[1]),.doutc(w_n629_3[2]),.din(w_n629_0[2]));
	jspl3 jspl3_w_n629_4(.douta(w_n629_4[0]),.doutb(w_n629_4[1]),.doutc(w_n629_4[2]),.din(w_n629_1[0]));
	jspl jspl_w_n629_5(.douta(w_n629_5[0]),.doutb(w_n629_5[1]),.din(w_n629_1[1]));
	jspl jspl_w_n630_0(.douta(w_n630_0[0]),.doutb(w_n630_0[1]),.din(n630));
	jspl jspl_w_n632_0(.douta(w_n632_0[0]),.doutb(w_n632_0[1]),.din(n632));
	jspl3 jspl3_w_n633_0(.douta(w_n633_0[0]),.doutb(w_n633_0[1]),.doutc(w_n633_0[2]),.din(n633));
	jspl3 jspl3_w_n633_1(.douta(w_n633_1[0]),.doutb(w_n633_1[1]),.doutc(w_n633_1[2]),.din(w_n633_0[0]));
	jspl3 jspl3_w_n633_2(.douta(w_n633_2[0]),.doutb(w_n633_2[1]),.doutc(w_n633_2[2]),.din(w_n633_0[1]));
	jspl3 jspl3_w_n633_3(.douta(w_n633_3[0]),.doutb(w_n633_3[1]),.doutc(w_n633_3[2]),.din(w_n633_0[2]));
	jspl3 jspl3_w_n633_4(.douta(w_n633_4[0]),.doutb(w_n633_4[1]),.doutc(w_n633_4[2]),.din(w_n633_1[0]));
	jspl3 jspl3_w_n633_5(.douta(w_n633_5[0]),.doutb(w_n633_5[1]),.doutc(w_n633_5[2]),.din(w_n633_1[1]));
	jspl jspl_w_n633_6(.douta(w_n633_6[0]),.doutb(w_n633_6[1]),.din(w_n633_1[2]));
	jspl jspl_w_n634_0(.douta(w_n634_0[0]),.doutb(w_n634_0[1]),.din(n634));
	jspl jspl_w_n637_0(.douta(w_n637_0[0]),.doutb(w_n637_0[1]),.din(n637));
	jspl3 jspl3_w_n638_0(.douta(w_n638_0[0]),.doutb(w_n638_0[1]),.doutc(w_n638_0[2]),.din(n638));
	jspl3 jspl3_w_n638_1(.douta(w_n638_1[0]),.doutb(w_n638_1[1]),.doutc(w_n638_1[2]),.din(w_n638_0[0]));
	jspl3 jspl3_w_n638_2(.douta(w_n638_2[0]),.doutb(w_n638_2[1]),.doutc(w_n638_2[2]),.din(w_n638_0[1]));
	jspl3 jspl3_w_n638_3(.douta(w_n638_3[0]),.doutb(w_n638_3[1]),.doutc(w_n638_3[2]),.din(w_n638_0[2]));
	jspl3 jspl3_w_n638_4(.douta(w_n638_4[0]),.doutb(w_n638_4[1]),.doutc(w_n638_4[2]),.din(w_n638_1[0]));
	jspl3 jspl3_w_n638_5(.douta(w_n638_5[0]),.doutb(w_n638_5[1]),.doutc(w_n638_5[2]),.din(w_n638_1[1]));
	jspl3 jspl3_w_n638_6(.douta(w_n638_6[0]),.doutb(w_n638_6[1]),.doutc(w_n638_6[2]),.din(w_n638_1[2]));
	jspl jspl_w_n638_7(.douta(w_n638_7[0]),.doutb(w_n638_7[1]),.din(w_n638_2[0]));
	jspl3 jspl3_w_n640_0(.douta(w_n640_0[0]),.doutb(w_n640_0[1]),.doutc(w_n640_0[2]),.din(n640));
	jspl3 jspl3_w_n640_1(.douta(w_n640_1[0]),.doutb(w_n640_1[1]),.doutc(w_n640_1[2]),.din(w_n640_0[0]));
	jspl3 jspl3_w_n640_2(.douta(w_n640_2[0]),.doutb(w_n640_2[1]),.doutc(w_n640_2[2]),.din(w_n640_0[1]));
	jspl3 jspl3_w_n640_3(.douta(w_n640_3[0]),.doutb(w_n640_3[1]),.doutc(w_n640_3[2]),.din(w_n640_0[2]));
	jspl3 jspl3_w_n640_4(.douta(w_n640_4[0]),.doutb(w_n640_4[1]),.doutc(w_n640_4[2]),.din(w_n640_1[0]));
	jspl3 jspl3_w_n640_5(.douta(w_n640_5[0]),.doutb(w_n640_5[1]),.doutc(w_n640_5[2]),.din(w_n640_1[1]));
	jspl3 jspl3_w_n640_6(.douta(w_n640_6[0]),.doutb(w_n640_6[1]),.doutc(w_n640_6[2]),.din(w_n640_1[2]));
	jspl jspl_w_n640_7(.douta(w_n640_7[0]),.doutb(w_n640_7[1]),.din(w_n640_2[0]));
	jspl3 jspl3_w_n646_0(.douta(w_n646_0[0]),.doutb(w_n646_0[1]),.doutc(w_n646_0[2]),.din(n646));
	jspl3 jspl3_w_n646_1(.douta(w_n646_1[0]),.doutb(w_n646_1[1]),.doutc(w_n646_1[2]),.din(w_n646_0[0]));
	jspl3 jspl3_w_n646_2(.douta(w_n646_2[0]),.doutb(w_n646_2[1]),.doutc(w_n646_2[2]),.din(w_n646_0[1]));
	jspl3 jspl3_w_n646_3(.douta(w_n646_3[0]),.doutb(w_n646_3[1]),.doutc(w_n646_3[2]),.din(w_n646_0[2]));
	jspl3 jspl3_w_n646_4(.douta(w_n646_4[0]),.doutb(w_n646_4[1]),.doutc(w_n646_4[2]),.din(w_n646_1[0]));
	jspl3 jspl3_w_n646_5(.douta(w_n646_5[0]),.doutb(w_n646_5[1]),.doutc(w_n646_5[2]),.din(w_n646_1[1]));
	jspl3 jspl3_w_n646_6(.douta(w_n646_6[0]),.doutb(w_n646_6[1]),.doutc(w_n646_6[2]),.din(w_n646_1[2]));
	jspl jspl_w_n646_7(.douta(w_n646_7[0]),.doutb(w_n646_7[1]),.din(w_n646_2[0]));
	jspl3 jspl3_w_n648_0(.douta(w_n648_0[0]),.doutb(w_n648_0[1]),.doutc(w_n648_0[2]),.din(n648));
	jspl3 jspl3_w_n648_1(.douta(w_n648_1[0]),.doutb(w_n648_1[1]),.doutc(w_n648_1[2]),.din(w_n648_0[0]));
	jspl3 jspl3_w_n648_2(.douta(w_n648_2[0]),.doutb(w_n648_2[1]),.doutc(w_n648_2[2]),.din(w_n648_0[1]));
	jspl3 jspl3_w_n648_3(.douta(w_n648_3[0]),.doutb(w_n648_3[1]),.doutc(w_n648_3[2]),.din(w_n648_0[2]));
	jspl jspl_w_n648_4(.douta(w_n648_4[0]),.doutb(w_n648_4[1]),.din(w_n648_1[0]));
	jspl jspl_w_n649_0(.douta(w_n649_0[0]),.doutb(w_dff_A_Hd7FvtnU2_1),.din(n649));
	jspl jspl_w_n650_0(.douta(w_n650_0[0]),.doutb(w_n650_0[1]),.din(n650));
	jspl3 jspl3_w_n651_0(.douta(w_n651_0[0]),.doutb(w_n651_0[1]),.doutc(w_n651_0[2]),.din(n651));
	jspl3 jspl3_w_n651_1(.douta(w_n651_1[0]),.doutb(w_n651_1[1]),.doutc(w_n651_1[2]),.din(w_n651_0[0]));
	jspl3 jspl3_w_n651_2(.douta(w_n651_2[0]),.doutb(w_n651_2[1]),.doutc(w_n651_2[2]),.din(w_n651_0[1]));
	jspl3 jspl3_w_n651_3(.douta(w_n651_3[0]),.doutb(w_n651_3[1]),.doutc(w_n651_3[2]),.din(w_n651_0[2]));
	jspl3 jspl3_w_n651_4(.douta(w_n651_4[0]),.doutb(w_n651_4[1]),.doutc(w_n651_4[2]),.din(w_n651_1[0]));
	jspl3 jspl3_w_n651_5(.douta(w_n651_5[0]),.doutb(w_n651_5[1]),.doutc(w_n651_5[2]),.din(w_n651_1[1]));
	jspl3 jspl3_w_n651_6(.douta(w_n651_6[0]),.doutb(w_n651_6[1]),.doutc(w_n651_6[2]),.din(w_n651_1[2]));
	jspl jspl_w_n651_7(.douta(w_n651_7[0]),.doutb(w_n651_7[1]),.din(w_n651_2[0]));
	jspl3 jspl3_w_n653_0(.douta(w_n653_0[0]),.doutb(w_n653_0[1]),.doutc(w_n653_0[2]),.din(n653));
	jspl3 jspl3_w_n653_1(.douta(w_n653_1[0]),.doutb(w_n653_1[1]),.doutc(w_n653_1[2]),.din(w_n653_0[0]));
	jspl3 jspl3_w_n653_2(.douta(w_n653_2[0]),.doutb(w_n653_2[1]),.doutc(w_n653_2[2]),.din(w_n653_0[1]));
	jspl3 jspl3_w_n653_3(.douta(w_n653_3[0]),.doutb(w_n653_3[1]),.doutc(w_n653_3[2]),.din(w_n653_0[2]));
	jspl3 jspl3_w_n653_4(.douta(w_n653_4[0]),.doutb(w_n653_4[1]),.doutc(w_n653_4[2]),.din(w_n653_1[0]));
	jspl3 jspl3_w_n653_5(.douta(w_n653_5[0]),.doutb(w_n653_5[1]),.doutc(w_n653_5[2]),.din(w_n653_1[1]));
	jspl3 jspl3_w_n653_6(.douta(w_n653_6[0]),.doutb(w_n653_6[1]),.doutc(w_n653_6[2]),.din(w_n653_1[2]));
	jspl jspl_w_n653_7(.douta(w_n653_7[0]),.doutb(w_n653_7[1]),.din(w_n653_2[0]));
	jspl3 jspl3_w_n680_0(.douta(w_n680_0[0]),.doutb(w_dff_A_1y3mWi0F2_1),.doutc(w_n680_0[2]),.din(n680));
	jspl3 jspl3_w_n680_1(.douta(w_n680_1[0]),.doutb(w_dff_A_eXb4slFv4_1),.doutc(w_n680_1[2]),.din(w_n680_0[0]));
	jspl3 jspl3_w_n680_2(.douta(w_dff_A_zQ0aq7wq3_0),.doutb(w_n680_2[1]),.doutc(w_dff_A_7lY5Beui3_2),.din(w_n680_0[1]));
	jspl3 jspl3_w_n680_3(.douta(w_dff_A_hW8AAyM75_0),.doutb(w_n680_3[1]),.doutc(w_dff_A_0etCkqs48_2),.din(w_n680_0[2]));
	jspl jspl_w_n680_4(.douta(w_n680_4[0]),.doutb(w_dff_A_XlRzNeBV1_1),.din(w_n680_1[0]));
	jspl jspl_w_n682_0(.douta(w_n682_0[0]),.doutb(w_dff_A_UECuCKLI4_1),.din(n682));
	jspl3 jspl3_w_n684_0(.douta(w_n684_0[0]),.doutb(w_n684_0[1]),.doutc(w_n684_0[2]),.din(n684));
	jspl jspl_w_n685_0(.douta(w_n685_0[0]),.doutb(w_n685_0[1]),.din(n685));
	jspl3 jspl3_w_n690_0(.douta(w_n690_0[0]),.doutb(w_n690_0[1]),.doutc(w_n690_0[2]),.din(n690));
	jspl jspl_w_n690_1(.douta(w_n690_1[0]),.doutb(w_n690_1[1]),.din(w_n690_0[0]));
	jspl jspl_w_n692_0(.douta(w_dff_A_mBfYHKxY7_0),.doutb(w_n692_0[1]),.din(n692));
	jspl3 jspl3_w_n703_0(.douta(w_n703_0[0]),.doutb(w_dff_A_13LBD0XT5_1),.doutc(w_dff_A_TiXB0ib65_2),.din(n703));
	jspl jspl_w_n703_1(.douta(w_dff_A_ElC4w09o7_0),.doutb(w_n703_1[1]),.din(w_n703_0[0]));
	jspl jspl_w_n704_0(.douta(w_dff_A_ntj8JBwS3_0),.doutb(w_n704_0[1]),.din(n704));
	jspl jspl_w_n718_0(.douta(w_dff_A_rKyVvHD16_0),.doutb(w_n718_0[1]),.din(w_dff_B_ksfw1szy2_2));
	jspl jspl_w_n733_0(.douta(w_n733_0[0]),.doutb(w_n733_0[1]),.din(n733));
	jspl3 jspl3_w_n741_0(.douta(w_n741_0[0]),.doutb(w_n741_0[1]),.doutc(w_n741_0[2]),.din(n741));
	jspl jspl_w_n741_1(.douta(w_n741_1[0]),.doutb(w_n741_1[1]),.din(w_n741_0[0]));
	jspl jspl_w_n748_0(.douta(w_n748_0[0]),.doutb(w_n748_0[1]),.din(n748));
	jspl jspl_w_n754_0(.douta(w_n754_0[0]),.doutb(w_n754_0[1]),.din(n754));
	jspl jspl_w_n759_0(.douta(w_dff_A_ZZIjx8KE4_0),.doutb(w_n759_0[1]),.din(n759));
	jspl jspl_w_n766_0(.douta(w_n766_0[0]),.doutb(w_n766_0[1]),.din(n766));
	jspl3 jspl3_w_n767_0(.douta(w_n767_0[0]),.doutb(w_dff_A_fdpzGfW16_1),.doutc(w_dff_A_rKBlyUaW6_2),.din(w_dff_B_gWNyL8z93_3));
	jspl jspl_w_n767_1(.douta(w_n767_1[0]),.doutb(w_dff_A_K39VnRtC5_1),.din(w_n767_0[0]));
	jspl3 jspl3_w_n771_0(.douta(w_n771_0[0]),.doutb(w_n771_0[1]),.doutc(w_dff_A_1d6IbwNh2_2),.din(n771));
	jspl jspl_w_n771_1(.douta(w_dff_A_SWu8eWN90_0),.doutb(w_n771_1[1]),.din(w_n771_0[0]));
	jspl jspl_w_n772_0(.douta(w_dff_A_KNoPRY6W5_0),.doutb(w_n772_0[1]),.din(n772));
	jspl jspl_w_n773_0(.douta(w_n773_0[0]),.doutb(w_dff_A_TA13gUh84_1),.din(n773));
	jspl jspl_w_n775_0(.douta(w_n775_0[0]),.doutb(w_n775_0[1]),.din(n775));
	jspl jspl_w_n777_0(.douta(w_n777_0[0]),.doutb(w_n777_0[1]),.din(n777));
	jspl jspl_w_n782_0(.douta(w_n782_0[0]),.doutb(w_n782_0[1]),.din(n782));
	jspl jspl_w_n798_0(.douta(w_dff_A_VCu3sJlL1_0),.doutb(w_n798_0[1]),.din(n798));
	jspl3 jspl3_w_n802_0(.douta(w_n802_0[0]),.doutb(w_dff_A_VMOJjKVJ3_1),.doutc(w_n802_0[2]),.din(n802));
	jspl jspl_w_n817_0(.douta(w_n817_0[0]),.doutb(w_dff_A_RMo9H0qy0_1),.din(n817));
	jspl jspl_w_n830_0(.douta(w_n830_0[0]),.doutb(w_n830_0[1]),.din(n830));
	jspl jspl_w_n833_0(.douta(w_dff_A_t8N1d5Pb7_0),.doutb(w_n833_0[1]),.din(n833));
	jspl3 jspl3_w_n845_0(.douta(w_n845_0[0]),.doutb(w_dff_A_gGJ6Bts46_1),.doutc(w_n845_0[2]),.din(n845));
	jspl jspl_w_n855_0(.douta(w_n855_0[0]),.doutb(w_n855_0[1]),.din(n855));
	jspl jspl_w_n860_0(.douta(w_n860_0[0]),.doutb(w_n860_0[1]),.din(n860));
	jspl jspl_w_n861_0(.douta(w_dff_A_hDEczb3X8_0),.doutb(w_n861_0[1]),.din(n861));
	jspl3 jspl3_w_n863_0(.douta(w_dff_A_nI7djk5b5_0),.doutb(w_n863_0[1]),.doutc(w_dff_A_Gt3uamDq6_2),.din(n863));
	jspl3 jspl3_w_n869_0(.douta(w_n869_0[0]),.doutb(w_n869_0[1]),.doutc(w_n869_0[2]),.din(n869));
	jspl jspl_w_n873_0(.douta(w_n873_0[0]),.doutb(w_n873_0[1]),.din(n873));
	jspl jspl_w_n875_0(.douta(w_n875_0[0]),.doutb(w_n875_0[1]),.din(n875));
	jspl jspl_w_n884_0(.douta(w_n884_0[0]),.doutb(w_n884_0[1]),.din(n884));
	jspl jspl_w_n887_0(.douta(w_n887_0[0]),.doutb(w_dff_A_BcUIqjLa9_1),.din(n887));
	jspl3 jspl3_w_n937_0(.douta(w_n937_0[0]),.doutb(w_n937_0[1]),.doutc(w_n937_0[2]),.din(n937));
	jspl jspl_w_n959_0(.douta(w_dff_A_Q4XdTMH92_0),.doutb(w_n959_0[1]),.din(n959));
	jspl3 jspl3_w_n987_0(.douta(w_n987_0[0]),.doutb(w_n987_0[1]),.doutc(w_n987_0[2]),.din(n987));
	jspl3 jspl3_w_n1029_0(.douta(w_n1029_0[0]),.doutb(w_n1029_0[1]),.doutc(w_n1029_0[2]),.din(n1029));
	jspl jspl_w_n1033_0(.douta(w_n1033_0[0]),.doutb(w_n1033_0[1]),.din(n1033));
	jspl jspl_w_n1036_0(.douta(w_n1036_0[0]),.doutb(w_n1036_0[1]),.din(n1036));
	jspl jspl_w_n1039_0(.douta(w_n1039_0[0]),.doutb(w_n1039_0[1]),.din(n1039));
	jspl jspl_w_n1040_0(.douta(w_n1040_0[0]),.doutb(w_n1040_0[1]),.din(n1040));
	jspl jspl_w_n1041_0(.douta(w_n1041_0[0]),.doutb(w_n1041_0[1]),.din(n1041));
	jspl jspl_w_n1043_0(.douta(w_n1043_0[0]),.doutb(w_dff_A_pHISlmdY7_1),.din(n1043));
	jspl jspl_w_n1044_0(.douta(w_n1044_0[0]),.doutb(w_n1044_0[1]),.din(n1044));
	jspl jspl_w_n1045_0(.douta(w_n1045_0[0]),.doutb(w_dff_A_6YUtQTR05_1),.din(n1045));
	jspl jspl_w_n1048_0(.douta(w_n1048_0[0]),.doutb(w_n1048_0[1]),.din(n1048));
	jspl3 jspl3_w_n1053_0(.douta(w_n1053_0[0]),.doutb(w_n1053_0[1]),.doutc(w_n1053_0[2]),.din(n1053));
	jspl jspl_w_n1056_0(.douta(w_dff_A_EwJdGVxo2_0),.doutb(w_n1056_0[1]),.din(w_dff_B_AjqoEEW30_2));
	jspl jspl_w_n1062_0(.douta(w_n1062_0[0]),.doutb(w_dff_A_siV6TsMS4_1),.din(n1062));
	jspl jspl_w_n1091_0(.douta(w_dff_A_9reIYKkx5_0),.doutb(w_n1091_0[1]),.din(n1091));
	jspl3 jspl3_w_n1114_0(.douta(w_n1114_0[0]),.doutb(w_n1114_0[1]),.doutc(w_n1114_0[2]),.din(n1114));
	jspl3 jspl3_w_n1159_0(.douta(w_n1159_0[0]),.doutb(w_n1159_0[1]),.doutc(w_n1159_0[2]),.din(n1159));
	jspl jspl_w_n1161_0(.douta(w_n1161_0[0]),.doutb(w_dff_A_bIPlIXri0_1),.din(n1161));
	jspl jspl_w_n1164_0(.douta(w_n1164_0[0]),.doutb(w_n1164_0[1]),.din(w_dff_B_DqFvCkPD9_2));
	jspl jspl_w_n1168_0(.douta(w_n1168_0[0]),.doutb(w_n1168_0[1]),.din(n1168));
	jspl jspl_w_n1170_0(.douta(w_n1170_0[0]),.doutb(w_dff_A_ZQl9FZJa0_1),.din(n1170));
	jspl jspl_w_n1177_0(.douta(w_n1177_0[0]),.doutb(w_dff_A_R35VlzGe6_1),.din(w_dff_B_6kMIKriX5_2));
	jspl jspl_w_n1178_0(.douta(w_n1178_0[0]),.doutb(w_dff_A_632WFSdJ0_1),.din(n1178));
	jspl jspl_w_n1179_0(.douta(w_n1179_0[0]),.doutb(w_n1179_0[1]),.din(n1179));
	jspl jspl_w_n1184_0(.douta(w_n1184_0[0]),.doutb(w_n1184_0[1]),.din(n1184));
	jdff dff_B_FisDzS2G3_1(.din(n92),.dout(w_dff_B_FisDzS2G3_1),.clk(gclk));
	jdff dff_B_6qk4aTx82_1(.din(w_dff_B_FisDzS2G3_1),.dout(w_dff_B_6qk4aTx82_1),.clk(gclk));
	jdff dff_B_JvinlRL29_1(.din(w_dff_B_6qk4aTx82_1),.dout(w_dff_B_JvinlRL29_1),.clk(gclk));
	jdff dff_B_TDSDGv6d9_0(.din(n114),.dout(w_dff_B_TDSDGv6d9_0),.clk(gclk));
	jdff dff_B_Ihv2Jms46_0(.din(n109),.dout(w_dff_B_Ihv2Jms46_0),.clk(gclk));
	jdff dff_B_C6ZHnywj8_1(.din(n93),.dout(w_dff_B_C6ZHnywj8_1),.clk(gclk));
	jdff dff_B_hMorE4od6_1(.din(w_dff_B_C6ZHnywj8_1),.dout(w_dff_B_hMorE4od6_1),.clk(gclk));
	jdff dff_B_EGuQuSgs1_0(.din(n100),.dout(w_dff_B_EGuQuSgs1_0),.clk(gclk));
	jdff dff_B_TASNkIqq7_1(.din(n583),.dout(w_dff_B_TASNkIqq7_1),.clk(gclk));
	jdff dff_B_Woaokfvf6_1(.din(w_dff_B_TASNkIqq7_1),.dout(w_dff_B_Woaokfvf6_1),.clk(gclk));
	jdff dff_B_QTLoulrx0_1(.din(w_dff_B_Woaokfvf6_1),.dout(w_dff_B_QTLoulrx0_1),.clk(gclk));
	jdff dff_B_08OolUYY8_1(.din(w_dff_B_QTLoulrx0_1),.dout(w_dff_B_08OolUYY8_1),.clk(gclk));
	jdff dff_B_GrXsNCMJ1_1(.din(w_dff_B_08OolUYY8_1),.dout(w_dff_B_GrXsNCMJ1_1),.clk(gclk));
	jdff dff_B_BEAgXbjz7_1(.din(w_dff_B_GrXsNCMJ1_1),.dout(w_dff_B_BEAgXbjz7_1),.clk(gclk));
	jdff dff_B_Bvb69Xmu7_1(.din(w_dff_B_BEAgXbjz7_1),.dout(w_dff_B_Bvb69Xmu7_1),.clk(gclk));
	jdff dff_B_8zPPKHFI8_1(.din(w_dff_B_Bvb69Xmu7_1),.dout(w_dff_B_8zPPKHFI8_1),.clk(gclk));
	jdff dff_B_0wR6m3aT5_1(.din(w_dff_B_8zPPKHFI8_1),.dout(w_dff_B_0wR6m3aT5_1),.clk(gclk));
	jdff dff_B_uwdEgYRk7_1(.din(w_dff_B_0wR6m3aT5_1),.dout(w_dff_B_uwdEgYRk7_1),.clk(gclk));
	jdff dff_B_AcMmPzkD8_1(.din(w_dff_B_uwdEgYRk7_1),.dout(w_dff_B_AcMmPzkD8_1),.clk(gclk));
	jdff dff_B_FyC6zzOK0_1(.din(w_dff_B_AcMmPzkD8_1),.dout(w_dff_B_FyC6zzOK0_1),.clk(gclk));
	jdff dff_B_tvCErOkh9_1(.din(w_dff_B_FyC6zzOK0_1),.dout(w_dff_B_tvCErOkh9_1),.clk(gclk));
	jdff dff_B_IiicwIpp4_1(.din(w_dff_B_tvCErOkh9_1),.dout(w_dff_B_IiicwIpp4_1),.clk(gclk));
	jdff dff_B_bhqxOEXJ8_1(.din(w_dff_B_IiicwIpp4_1),.dout(w_dff_B_bhqxOEXJ8_1),.clk(gclk));
	jdff dff_B_EQCVdU6e3_1(.din(w_dff_B_bhqxOEXJ8_1),.dout(w_dff_B_EQCVdU6e3_1),.clk(gclk));
	jdff dff_B_tkqstEIK6_0(.din(n607),.dout(w_dff_B_tkqstEIK6_0),.clk(gclk));
	jdff dff_B_tNVLTYxr0_0(.din(w_dff_B_tkqstEIK6_0),.dout(w_dff_B_tNVLTYxr0_0),.clk(gclk));
	jdff dff_B_QSMvEAzn2_0(.din(w_dff_B_tNVLTYxr0_0),.dout(w_dff_B_QSMvEAzn2_0),.clk(gclk));
	jdff dff_B_N8qLehVz8_0(.din(w_dff_B_QSMvEAzn2_0),.dout(w_dff_B_N8qLehVz8_0),.clk(gclk));
	jdff dff_B_iTzdb2r78_0(.din(w_dff_B_N8qLehVz8_0),.dout(w_dff_B_iTzdb2r78_0),.clk(gclk));
	jdff dff_B_irI9PjkJ7_0(.din(w_dff_B_iTzdb2r78_0),.dout(w_dff_B_irI9PjkJ7_0),.clk(gclk));
	jdff dff_B_nZgEs5t84_0(.din(w_dff_B_irI9PjkJ7_0),.dout(w_dff_B_nZgEs5t84_0),.clk(gclk));
	jdff dff_B_ni6t9HIS6_0(.din(w_dff_B_nZgEs5t84_0),.dout(w_dff_B_ni6t9HIS6_0),.clk(gclk));
	jdff dff_B_mtzlxig94_0(.din(w_dff_B_ni6t9HIS6_0),.dout(w_dff_B_mtzlxig94_0),.clk(gclk));
	jdff dff_B_BzfrBKk04_0(.din(w_dff_B_mtzlxig94_0),.dout(w_dff_B_BzfrBKk04_0),.clk(gclk));
	jdff dff_B_8L2g9nce6_0(.din(w_dff_B_BzfrBKk04_0),.dout(w_dff_B_8L2g9nce6_0),.clk(gclk));
	jdff dff_B_0QPvJRGD3_0(.din(w_dff_B_8L2g9nce6_0),.dout(w_dff_B_0QPvJRGD3_0),.clk(gclk));
	jdff dff_B_lnBonCWs7_0(.din(w_dff_B_0QPvJRGD3_0),.dout(w_dff_B_lnBonCWs7_0),.clk(gclk));
	jdff dff_B_UReCyPV51_0(.din(w_dff_B_lnBonCWs7_0),.dout(w_dff_B_UReCyPV51_0),.clk(gclk));
	jdff dff_B_Kwxh1Sr80_0(.din(n795),.dout(w_dff_B_Kwxh1Sr80_0),.clk(gclk));
	jdff dff_B_6wTKYiMy6_0(.din(w_dff_B_Kwxh1Sr80_0),.dout(w_dff_B_6wTKYiMy6_0),.clk(gclk));
	jdff dff_B_HNxUzeNO3_0(.din(w_dff_B_6wTKYiMy6_0),.dout(w_dff_B_HNxUzeNO3_0),.clk(gclk));
	jdff dff_B_8y5Qywf70_0(.din(w_dff_B_HNxUzeNO3_0),.dout(w_dff_B_8y5Qywf70_0),.clk(gclk));
	jdff dff_B_qz0yT4u13_0(.din(w_dff_B_8y5Qywf70_0),.dout(w_dff_B_qz0yT4u13_0),.clk(gclk));
	jdff dff_B_ujE6Yytb4_0(.din(w_dff_B_qz0yT4u13_0),.dout(w_dff_B_ujE6Yytb4_0),.clk(gclk));
	jdff dff_B_Jgozzp5O5_0(.din(w_dff_B_ujE6Yytb4_0),.dout(w_dff_B_Jgozzp5O5_0),.clk(gclk));
	jdff dff_B_Ij2wRnEv9_0(.din(w_dff_B_Jgozzp5O5_0),.dout(w_dff_B_Ij2wRnEv9_0),.clk(gclk));
	jdff dff_B_sVx04yGb5_0(.din(w_dff_B_Ij2wRnEv9_0),.dout(w_dff_B_sVx04yGb5_0),.clk(gclk));
	jdff dff_B_yxPDP1Hg4_0(.din(w_dff_B_sVx04yGb5_0),.dout(w_dff_B_yxPDP1Hg4_0),.clk(gclk));
	jdff dff_B_PQqpOgbm4_0(.din(w_dff_B_yxPDP1Hg4_0),.dout(w_dff_B_PQqpOgbm4_0),.clk(gclk));
	jdff dff_B_IW7K4Xhv7_0(.din(w_dff_B_PQqpOgbm4_0),.dout(w_dff_B_IW7K4Xhv7_0),.clk(gclk));
	jdff dff_B_Xk7HAGc29_0(.din(w_dff_B_IW7K4Xhv7_0),.dout(w_dff_B_Xk7HAGc29_0),.clk(gclk));
	jdff dff_B_VXjQKKOq0_0(.din(w_dff_B_Xk7HAGc29_0),.dout(w_dff_B_VXjQKKOq0_0),.clk(gclk));
	jdff dff_B_pzOzuQKD8_0(.din(w_dff_B_VXjQKKOq0_0),.dout(w_dff_B_pzOzuQKD8_0),.clk(gclk));
	jdff dff_B_aXgPwDHK0_0(.din(w_dff_B_pzOzuQKD8_0),.dout(w_dff_B_aXgPwDHK0_0),.clk(gclk));
	jdff dff_B_tv2ZYgBB6_0(.din(w_dff_B_aXgPwDHK0_0),.dout(w_dff_B_tv2ZYgBB6_0),.clk(gclk));
	jdff dff_B_YjUwNIFM7_0(.din(n794),.dout(w_dff_B_YjUwNIFM7_0),.clk(gclk));
	jdff dff_A_DQoYhr6W3_1(.dout(w_n120_0[1]),.din(w_dff_A_DQoYhr6W3_1),.clk(gclk));
	jdff dff_A_TyPS3WoP1_1(.dout(w_dff_A_DQoYhr6W3_1),.din(w_dff_A_TyPS3WoP1_1),.clk(gclk));
	jdff dff_A_UDU0rIU67_1(.dout(w_dff_A_TyPS3WoP1_1),.din(w_dff_A_UDU0rIU67_1),.clk(gclk));
	jdff dff_B_1OBZCMhy3_0(.din(n791),.dout(w_dff_B_1OBZCMhy3_0),.clk(gclk));
	jdff dff_B_tSx2xLMj3_1(.din(n762),.dout(w_dff_B_tSx2xLMj3_1),.clk(gclk));
	jdff dff_B_C8rCXM4B9_1(.din(w_dff_B_tSx2xLMj3_1),.dout(w_dff_B_C8rCXM4B9_1),.clk(gclk));
	jdff dff_B_G0UMSRUW8_1(.din(w_dff_B_C8rCXM4B9_1),.dout(w_dff_B_G0UMSRUW8_1),.clk(gclk));
	jdff dff_B_BkJ0qat38_1(.din(w_dff_B_G0UMSRUW8_1),.dout(w_dff_B_BkJ0qat38_1),.clk(gclk));
	jdff dff_B_fUV0KDod1_1(.din(w_dff_B_BkJ0qat38_1),.dout(w_dff_B_fUV0KDod1_1),.clk(gclk));
	jdff dff_B_666hIiDX3_1(.din(w_dff_B_fUV0KDod1_1),.dout(w_dff_B_666hIiDX3_1),.clk(gclk));
	jdff dff_B_Xmye5mS34_1(.din(w_dff_B_666hIiDX3_1),.dout(w_dff_B_Xmye5mS34_1),.clk(gclk));
	jdff dff_B_xVzKSrU77_1(.din(w_dff_B_Xmye5mS34_1),.dout(w_dff_B_xVzKSrU77_1),.clk(gclk));
	jdff dff_B_d7gv71Hn9_1(.din(w_dff_B_xVzKSrU77_1),.dout(w_dff_B_d7gv71Hn9_1),.clk(gclk));
	jdff dff_B_C5TkIlfG6_1(.din(w_dff_B_d7gv71Hn9_1),.dout(w_dff_B_C5TkIlfG6_1),.clk(gclk));
	jdff dff_B_PWsTpzww3_1(.din(w_dff_B_C5TkIlfG6_1),.dout(w_dff_B_PWsTpzww3_1),.clk(gclk));
	jdff dff_B_CJ0tkKYS7_1(.din(w_dff_B_PWsTpzww3_1),.dout(w_dff_B_CJ0tkKYS7_1),.clk(gclk));
	jdff dff_B_t7byUmWW0_1(.din(w_dff_B_CJ0tkKYS7_1),.dout(w_dff_B_t7byUmWW0_1),.clk(gclk));
	jdff dff_B_71Z0PtaJ2_1(.din(w_dff_B_t7byUmWW0_1),.dout(w_dff_B_71Z0PtaJ2_1),.clk(gclk));
	jdff dff_B_GUTpCPzJ4_1(.din(w_dff_B_71Z0PtaJ2_1),.dout(w_dff_B_GUTpCPzJ4_1),.clk(gclk));
	jdff dff_B_80BwfMuo1_1(.din(w_dff_B_GUTpCPzJ4_1),.dout(w_dff_B_80BwfMuo1_1),.clk(gclk));
	jdff dff_B_lKf6zE3u4_1(.din(w_dff_B_80BwfMuo1_1),.dout(w_dff_B_lKf6zE3u4_1),.clk(gclk));
	jdff dff_B_XEYBo1O55_1(.din(w_dff_B_lKf6zE3u4_1),.dout(w_dff_B_XEYBo1O55_1),.clk(gclk));
	jdff dff_B_L1sWVBgv2_0(.din(n783),.dout(w_dff_B_L1sWVBgv2_0),.clk(gclk));
	jdff dff_A_l0vAzSjO1_0(.dout(w_n112_0[0]),.din(w_dff_A_l0vAzSjO1_0),.clk(gclk));
	jdff dff_B_O0pQzvgJ1_1(.din(n1171),.dout(w_dff_B_O0pQzvgJ1_1),.clk(gclk));
	jdff dff_B_frMcGxgf5_1(.din(w_dff_B_O0pQzvgJ1_1),.dout(w_dff_B_frMcGxgf5_1),.clk(gclk));
	jdff dff_B_jqOtryg55_1(.din(n1172),.dout(w_dff_B_jqOtryg55_1),.clk(gclk));
	jdff dff_B_oOkU1t0k3_1(.din(w_dff_B_jqOtryg55_1),.dout(w_dff_B_oOkU1t0k3_1),.clk(gclk));
	jdff dff_B_rExM3eu09_1(.din(w_dff_B_oOkU1t0k3_1),.dout(w_dff_B_rExM3eu09_1),.clk(gclk));
	jdff dff_B_VO0XmfdD9_1(.din(w_dff_B_rExM3eu09_1),.dout(w_dff_B_VO0XmfdD9_1),.clk(gclk));
	jdff dff_B_tm5M35OS1_1(.din(w_dff_B_VO0XmfdD9_1),.dout(w_dff_B_tm5M35OS1_1),.clk(gclk));
	jdff dff_B_G1cOep062_1(.din(w_dff_B_tm5M35OS1_1),.dout(w_dff_B_G1cOep062_1),.clk(gclk));
	jdff dff_B_MQS5xDSO2_1(.din(w_dff_B_G1cOep062_1),.dout(w_dff_B_MQS5xDSO2_1),.clk(gclk));
	jdff dff_B_CNW9yy9e7_1(.din(w_dff_B_MQS5xDSO2_1),.dout(w_dff_B_CNW9yy9e7_1),.clk(gclk));
	jdff dff_B_r4uPlvMp9_1(.din(w_dff_B_CNW9yy9e7_1),.dout(w_dff_B_r4uPlvMp9_1),.clk(gclk));
	jdff dff_B_E5Je6U2n4_1(.din(w_dff_B_r4uPlvMp9_1),.dout(w_dff_B_E5Je6U2n4_1),.clk(gclk));
	jdff dff_B_Cy6THfc74_1(.din(w_dff_B_E5Je6U2n4_1),.dout(w_dff_B_Cy6THfc74_1),.clk(gclk));
	jdff dff_B_8n8mkhmR1_1(.din(w_dff_B_Cy6THfc74_1),.dout(w_dff_B_8n8mkhmR1_1),.clk(gclk));
	jdff dff_B_sCyau8fA4_1(.din(w_dff_B_8n8mkhmR1_1),.dout(w_dff_B_sCyau8fA4_1),.clk(gclk));
	jdff dff_B_n6B4OGTu7_1(.din(w_dff_B_sCyau8fA4_1),.dout(w_dff_B_n6B4OGTu7_1),.clk(gclk));
	jdff dff_B_hWlgKtWM3_1(.din(w_dff_B_n6B4OGTu7_1),.dout(w_dff_B_hWlgKtWM3_1),.clk(gclk));
	jdff dff_B_iL5VXfsp1_1(.din(w_dff_B_hWlgKtWM3_1),.dout(w_dff_B_iL5VXfsp1_1),.clk(gclk));
	jdff dff_B_BdE3Le4u3_1(.din(w_dff_B_iL5VXfsp1_1),.dout(w_dff_B_BdE3Le4u3_1),.clk(gclk));
	jdff dff_B_e0Gwb0W57_1(.din(w_dff_B_BdE3Le4u3_1),.dout(w_dff_B_e0Gwb0W57_1),.clk(gclk));
	jdff dff_B_Ie3d7nLS0_1(.din(w_dff_B_e0Gwb0W57_1),.dout(w_dff_B_Ie3d7nLS0_1),.clk(gclk));
	jdff dff_B_CacUVfs86_1(.din(w_dff_B_Ie3d7nLS0_1),.dout(w_dff_B_CacUVfs86_1),.clk(gclk));
	jdff dff_B_x4oHjoEA8_1(.din(w_dff_B_CacUVfs86_1),.dout(w_dff_B_x4oHjoEA8_1),.clk(gclk));
	jdff dff_B_yTxwHFCj4_1(.din(w_dff_B_x4oHjoEA8_1),.dout(w_dff_B_yTxwHFCj4_1),.clk(gclk));
	jdff dff_B_dKsDdogj7_1(.din(w_dff_B_yTxwHFCj4_1),.dout(w_dff_B_dKsDdogj7_1),.clk(gclk));
	jdff dff_B_BhqnfbyR0_1(.din(w_dff_B_dKsDdogj7_1),.dout(w_dff_B_BhqnfbyR0_1),.clk(gclk));
	jdff dff_B_KQ6GFgsG1_1(.din(w_dff_B_BhqnfbyR0_1),.dout(w_dff_B_KQ6GFgsG1_1),.clk(gclk));
	jdff dff_B_MknqKfFr2_1(.din(w_dff_B_KQ6GFgsG1_1),.dout(w_dff_B_MknqKfFr2_1),.clk(gclk));
	jdff dff_B_8HFEJnXu5_1(.din(w_dff_B_MknqKfFr2_1),.dout(w_dff_B_8HFEJnXu5_1),.clk(gclk));
	jdff dff_B_FwJFZ6BF6_1(.din(w_dff_B_8HFEJnXu5_1),.dout(w_dff_B_FwJFZ6BF6_1),.clk(gclk));
	jdff dff_B_AmjHcgx98_0(.din(n1166),.dout(w_dff_B_AmjHcgx98_0),.clk(gclk));
	jdff dff_B_48cNaTjh5_0(.din(n1165),.dout(w_dff_B_48cNaTjh5_0),.clk(gclk));
	jdff dff_A_bIPlIXri0_1(.dout(w_n1161_0[1]),.din(w_dff_A_bIPlIXri0_1),.clk(gclk));
	jdff dff_B_aG3jgnq64_1(.din(n1182),.dout(w_dff_B_aG3jgnq64_1),.clk(gclk));
	jdff dff_B_ZAzMLZjE2_1(.din(w_dff_B_aG3jgnq64_1),.dout(w_dff_B_ZAzMLZjE2_1),.clk(gclk));
	jdff dff_B_743ovYwE6_1(.din(w_dff_B_ZAzMLZjE2_1),.dout(w_dff_B_743ovYwE6_1),.clk(gclk));
	jdff dff_B_4dxmTCCL6_1(.din(w_dff_B_743ovYwE6_1),.dout(w_dff_B_4dxmTCCL6_1),.clk(gclk));
	jdff dff_B_Tr26cAK27_1(.din(w_dff_B_4dxmTCCL6_1),.dout(w_dff_B_Tr26cAK27_1),.clk(gclk));
	jdff dff_B_p3kTBsde8_1(.din(w_dff_B_Tr26cAK27_1),.dout(w_dff_B_p3kTBsde8_1),.clk(gclk));
	jdff dff_B_ENVTFoNk4_1(.din(w_dff_B_p3kTBsde8_1),.dout(w_dff_B_ENVTFoNk4_1),.clk(gclk));
	jdff dff_B_K0pcvSBU0_1(.din(w_dff_B_ENVTFoNk4_1),.dout(w_dff_B_K0pcvSBU0_1),.clk(gclk));
	jdff dff_B_LbYXLk3t8_1(.din(w_dff_B_K0pcvSBU0_1),.dout(w_dff_B_LbYXLk3t8_1),.clk(gclk));
	jdff dff_B_mRcD0r6B8_1(.din(w_dff_B_LbYXLk3t8_1),.dout(w_dff_B_mRcD0r6B8_1),.clk(gclk));
	jdff dff_B_ifODZ0W21_1(.din(w_dff_B_mRcD0r6B8_1),.dout(w_dff_B_ifODZ0W21_1),.clk(gclk));
	jdff dff_B_C8Byw6xg1_1(.din(w_dff_B_ifODZ0W21_1),.dout(w_dff_B_C8Byw6xg1_1),.clk(gclk));
	jdff dff_B_jIOcnVBj3_1(.din(w_dff_B_C8Byw6xg1_1),.dout(w_dff_B_jIOcnVBj3_1),.clk(gclk));
	jdff dff_B_kTZ06aED6_1(.din(w_dff_B_jIOcnVBj3_1),.dout(w_dff_B_kTZ06aED6_1),.clk(gclk));
	jdff dff_B_0l7va75j8_1(.din(w_dff_B_kTZ06aED6_1),.dout(w_dff_B_0l7va75j8_1),.clk(gclk));
	jdff dff_B_Af02HnkB5_1(.din(w_dff_B_0l7va75j8_1),.dout(w_dff_B_Af02HnkB5_1),.clk(gclk));
	jdff dff_B_5ed415NZ0_1(.din(w_dff_B_Af02HnkB5_1),.dout(w_dff_B_5ed415NZ0_1),.clk(gclk));
	jdff dff_B_46wcFXb09_1(.din(w_dff_B_5ed415NZ0_1),.dout(w_dff_B_46wcFXb09_1),.clk(gclk));
	jdff dff_B_haq2xpEC6_1(.din(w_dff_B_46wcFXb09_1),.dout(w_dff_B_haq2xpEC6_1),.clk(gclk));
	jdff dff_B_HiuuKYU86_1(.din(w_dff_B_haq2xpEC6_1),.dout(w_dff_B_HiuuKYU86_1),.clk(gclk));
	jdff dff_B_2EP0XXjU0_1(.din(w_dff_B_HiuuKYU86_1),.dout(w_dff_B_2EP0XXjU0_1),.clk(gclk));
	jdff dff_B_6vypaYpT5_1(.din(w_dff_B_2EP0XXjU0_1),.dout(w_dff_B_6vypaYpT5_1),.clk(gclk));
	jdff dff_B_Su3dtXyJ0_1(.din(w_dff_B_6vypaYpT5_1),.dout(w_dff_B_Su3dtXyJ0_1),.clk(gclk));
	jdff dff_B_IDtFmd019_1(.din(w_dff_B_Su3dtXyJ0_1),.dout(w_dff_B_IDtFmd019_1),.clk(gclk));
	jdff dff_B_lY2Ax7b13_1(.din(w_dff_B_IDtFmd019_1),.dout(w_dff_B_lY2Ax7b13_1),.clk(gclk));
	jdff dff_B_PpUIfjdo0_1(.din(G2897),.dout(w_dff_B_PpUIfjdo0_1),.clk(gclk));
	jdff dff_B_kWRWoWwz2_1(.din(w_dff_B_PpUIfjdo0_1),.dout(w_dff_B_kWRWoWwz2_1),.clk(gclk));
	jdff dff_B_YEK212ql2_1(.din(w_dff_B_kWRWoWwz2_1),.dout(w_dff_B_YEK212ql2_1),.clk(gclk));
	jdff dff_B_cNXx9oAG3_1(.din(w_dff_B_YEK212ql2_1),.dout(w_dff_B_cNXx9oAG3_1),.clk(gclk));
	jdff dff_B_k27Nc5al7_1(.din(w_dff_B_cNXx9oAG3_1),.dout(w_dff_B_k27Nc5al7_1),.clk(gclk));
	jdff dff_B_gdKSErvz3_1(.din(w_dff_B_k27Nc5al7_1),.dout(w_dff_B_gdKSErvz3_1),.clk(gclk));
	jdff dff_B_3YqxDNy86_1(.din(w_dff_B_gdKSErvz3_1),.dout(w_dff_B_3YqxDNy86_1),.clk(gclk));
	jdff dff_B_VOogdegQ3_1(.din(w_dff_B_3YqxDNy86_1),.dout(w_dff_B_VOogdegQ3_1),.clk(gclk));
	jdff dff_B_TrqHHWcp0_1(.din(w_dff_B_VOogdegQ3_1),.dout(w_dff_B_TrqHHWcp0_1),.clk(gclk));
	jdff dff_B_Nv92AX2s3_1(.din(w_dff_B_TrqHHWcp0_1),.dout(w_dff_B_Nv92AX2s3_1),.clk(gclk));
	jdff dff_B_6O3fuYLp3_1(.din(w_dff_B_Nv92AX2s3_1),.dout(w_dff_B_6O3fuYLp3_1),.clk(gclk));
	jdff dff_B_z6hslOBF1_1(.din(w_dff_B_6O3fuYLp3_1),.dout(w_dff_B_z6hslOBF1_1),.clk(gclk));
	jdff dff_B_yYF6DQEQ6_1(.din(w_dff_B_z6hslOBF1_1),.dout(w_dff_B_yYF6DQEQ6_1),.clk(gclk));
	jdff dff_B_nV7xsVl07_1(.din(w_dff_B_yYF6DQEQ6_1),.dout(w_dff_B_nV7xsVl07_1),.clk(gclk));
	jdff dff_B_3noChfJt3_1(.din(w_dff_B_nV7xsVl07_1),.dout(w_dff_B_3noChfJt3_1),.clk(gclk));
	jdff dff_B_8u2om3fQ9_1(.din(w_dff_B_3noChfJt3_1),.dout(w_dff_B_8u2om3fQ9_1),.clk(gclk));
	jdff dff_B_gfaZYkfb7_1(.din(w_dff_B_8u2om3fQ9_1),.dout(w_dff_B_gfaZYkfb7_1),.clk(gclk));
	jdff dff_B_QfVH3H3o5_1(.din(w_dff_B_gfaZYkfb7_1),.dout(w_dff_B_QfVH3H3o5_1),.clk(gclk));
	jdff dff_B_GBSecZs41_1(.din(w_dff_B_QfVH3H3o5_1),.dout(w_dff_B_GBSecZs41_1),.clk(gclk));
	jdff dff_B_nJa0Ckn88_1(.din(w_dff_B_GBSecZs41_1),.dout(w_dff_B_nJa0Ckn88_1),.clk(gclk));
	jdff dff_B_4xK9j6Kk4_1(.din(w_dff_B_nJa0Ckn88_1),.dout(w_dff_B_4xK9j6Kk4_1),.clk(gclk));
	jdff dff_B_DDcZLK1K1_1(.din(w_dff_B_4xK9j6Kk4_1),.dout(w_dff_B_DDcZLK1K1_1),.clk(gclk));
	jdff dff_B_WxdgpjY17_1(.din(w_dff_B_DDcZLK1K1_1),.dout(w_dff_B_WxdgpjY17_1),.clk(gclk));
	jdff dff_B_HE9qHSVP8_1(.din(w_dff_B_WxdgpjY17_1),.dout(w_dff_B_HE9qHSVP8_1),.clk(gclk));
	jdff dff_B_IU7mi6NF8_1(.din(w_dff_B_HE9qHSVP8_1),.dout(w_dff_B_IU7mi6NF8_1),.clk(gclk));
	jdff dff_B_nVelMIe07_1(.din(w_dff_B_IU7mi6NF8_1),.dout(w_dff_B_nVelMIe07_1),.clk(gclk));
	jdff dff_B_fhFDzsU53_1(.din(w_dff_B_nVelMIe07_1),.dout(w_dff_B_fhFDzsU53_1),.clk(gclk));
	jdff dff_A_oEkZzEYX3_1(.dout(w_n1178_0[1]),.din(w_dff_A_oEkZzEYX3_1),.clk(gclk));
	jdff dff_A_2aSPumVB0_1(.dout(w_dff_A_oEkZzEYX3_1),.din(w_dff_A_2aSPumVB0_1),.clk(gclk));
	jdff dff_A_nc9pRLfW0_1(.dout(w_dff_A_2aSPumVB0_1),.din(w_dff_A_nc9pRLfW0_1),.clk(gclk));
	jdff dff_A_ymO1q5WJ9_1(.dout(w_dff_A_nc9pRLfW0_1),.din(w_dff_A_ymO1q5WJ9_1),.clk(gclk));
	jdff dff_A_97gF6N6G5_1(.dout(w_dff_A_ymO1q5WJ9_1),.din(w_dff_A_97gF6N6G5_1),.clk(gclk));
	jdff dff_A_DGqvrLS62_1(.dout(w_dff_A_97gF6N6G5_1),.din(w_dff_A_DGqvrLS62_1),.clk(gclk));
	jdff dff_A_xuAxr93G4_1(.dout(w_dff_A_DGqvrLS62_1),.din(w_dff_A_xuAxr93G4_1),.clk(gclk));
	jdff dff_A_uMceIChW0_1(.dout(w_dff_A_xuAxr93G4_1),.din(w_dff_A_uMceIChW0_1),.clk(gclk));
	jdff dff_A_OJgpjU1k7_1(.dout(w_dff_A_uMceIChW0_1),.din(w_dff_A_OJgpjU1k7_1),.clk(gclk));
	jdff dff_A_sKgk3hIT5_1(.dout(w_dff_A_OJgpjU1k7_1),.din(w_dff_A_sKgk3hIT5_1),.clk(gclk));
	jdff dff_A_x8Ypizl98_1(.dout(w_dff_A_sKgk3hIT5_1),.din(w_dff_A_x8Ypizl98_1),.clk(gclk));
	jdff dff_A_WTIedmAo2_1(.dout(w_dff_A_x8Ypizl98_1),.din(w_dff_A_WTIedmAo2_1),.clk(gclk));
	jdff dff_A_TIJGeD1Z6_1(.dout(w_dff_A_WTIedmAo2_1),.din(w_dff_A_TIJGeD1Z6_1),.clk(gclk));
	jdff dff_A_6zUO43MB8_1(.dout(w_dff_A_TIJGeD1Z6_1),.din(w_dff_A_6zUO43MB8_1),.clk(gclk));
	jdff dff_A_89fyoYdW2_1(.dout(w_dff_A_6zUO43MB8_1),.din(w_dff_A_89fyoYdW2_1),.clk(gclk));
	jdff dff_A_BtXQrUYB8_1(.dout(w_dff_A_89fyoYdW2_1),.din(w_dff_A_BtXQrUYB8_1),.clk(gclk));
	jdff dff_A_DQGQIvbH8_1(.dout(w_dff_A_BtXQrUYB8_1),.din(w_dff_A_DQGQIvbH8_1),.clk(gclk));
	jdff dff_A_fC6BJDS77_1(.dout(w_dff_A_DQGQIvbH8_1),.din(w_dff_A_fC6BJDS77_1),.clk(gclk));
	jdff dff_A_iv679SmZ3_1(.dout(w_dff_A_fC6BJDS77_1),.din(w_dff_A_iv679SmZ3_1),.clk(gclk));
	jdff dff_A_g74wpa3S6_1(.dout(w_dff_A_iv679SmZ3_1),.din(w_dff_A_g74wpa3S6_1),.clk(gclk));
	jdff dff_A_Q6aavcP76_1(.dout(w_dff_A_g74wpa3S6_1),.din(w_dff_A_Q6aavcP76_1),.clk(gclk));
	jdff dff_A_1ykcvOfP0_1(.dout(w_dff_A_Q6aavcP76_1),.din(w_dff_A_1ykcvOfP0_1),.clk(gclk));
	jdff dff_A_Tv9wjDeq9_1(.dout(w_dff_A_1ykcvOfP0_1),.din(w_dff_A_Tv9wjDeq9_1),.clk(gclk));
	jdff dff_A_oUsiejR33_1(.dout(w_dff_A_Tv9wjDeq9_1),.din(w_dff_A_oUsiejR33_1),.clk(gclk));
	jdff dff_A_LHYgxu1A5_1(.dout(w_dff_A_oUsiejR33_1),.din(w_dff_A_LHYgxu1A5_1),.clk(gclk));
	jdff dff_A_632WFSdJ0_1(.dout(w_dff_A_LHYgxu1A5_1),.din(w_dff_A_632WFSdJ0_1),.clk(gclk));
	jdff dff_A_dkfYjhzC3_1(.dout(w_n1170_0[1]),.din(w_dff_A_dkfYjhzC3_1),.clk(gclk));
	jdff dff_A_e1I1FwBw6_1(.dout(w_dff_A_dkfYjhzC3_1),.din(w_dff_A_e1I1FwBw6_1),.clk(gclk));
	jdff dff_A_EaGAQYq91_1(.dout(w_dff_A_e1I1FwBw6_1),.din(w_dff_A_EaGAQYq91_1),.clk(gclk));
	jdff dff_A_TUSdV0av9_1(.dout(w_dff_A_EaGAQYq91_1),.din(w_dff_A_TUSdV0av9_1),.clk(gclk));
	jdff dff_A_R3xkoru75_1(.dout(w_dff_A_TUSdV0av9_1),.din(w_dff_A_R3xkoru75_1),.clk(gclk));
	jdff dff_A_XoITSO2M6_1(.dout(w_dff_A_R3xkoru75_1),.din(w_dff_A_XoITSO2M6_1),.clk(gclk));
	jdff dff_A_GEHe4JQR6_1(.dout(w_dff_A_XoITSO2M6_1),.din(w_dff_A_GEHe4JQR6_1),.clk(gclk));
	jdff dff_A_6mCe0wye9_1(.dout(w_dff_A_GEHe4JQR6_1),.din(w_dff_A_6mCe0wye9_1),.clk(gclk));
	jdff dff_A_MT7vUpff4_1(.dout(w_dff_A_6mCe0wye9_1),.din(w_dff_A_MT7vUpff4_1),.clk(gclk));
	jdff dff_A_HxieEi5Q0_1(.dout(w_dff_A_MT7vUpff4_1),.din(w_dff_A_HxieEi5Q0_1),.clk(gclk));
	jdff dff_A_KzrAGZO89_1(.dout(w_dff_A_HxieEi5Q0_1),.din(w_dff_A_KzrAGZO89_1),.clk(gclk));
	jdff dff_A_gsDHJLme9_1(.dout(w_dff_A_KzrAGZO89_1),.din(w_dff_A_gsDHJLme9_1),.clk(gclk));
	jdff dff_A_lFJsCO5g3_1(.dout(w_dff_A_gsDHJLme9_1),.din(w_dff_A_lFJsCO5g3_1),.clk(gclk));
	jdff dff_A_yz6Ci5FY0_1(.dout(w_dff_A_lFJsCO5g3_1),.din(w_dff_A_yz6Ci5FY0_1),.clk(gclk));
	jdff dff_A_l7UgMVOv0_1(.dout(w_dff_A_yz6Ci5FY0_1),.din(w_dff_A_l7UgMVOv0_1),.clk(gclk));
	jdff dff_A_gmbyOslU0_1(.dout(w_dff_A_l7UgMVOv0_1),.din(w_dff_A_gmbyOslU0_1),.clk(gclk));
	jdff dff_A_6WUQ2ZRA2_1(.dout(w_dff_A_gmbyOslU0_1),.din(w_dff_A_6WUQ2ZRA2_1),.clk(gclk));
	jdff dff_A_J2vkXNR49_1(.dout(w_dff_A_6WUQ2ZRA2_1),.din(w_dff_A_J2vkXNR49_1),.clk(gclk));
	jdff dff_A_zPe37f148_1(.dout(w_dff_A_J2vkXNR49_1),.din(w_dff_A_zPe37f148_1),.clk(gclk));
	jdff dff_A_GejfoAzr1_1(.dout(w_dff_A_zPe37f148_1),.din(w_dff_A_GejfoAzr1_1),.clk(gclk));
	jdff dff_A_ztItkpuL0_1(.dout(w_dff_A_GejfoAzr1_1),.din(w_dff_A_ztItkpuL0_1),.clk(gclk));
	jdff dff_A_ucWO2dQd1_1(.dout(w_dff_A_ztItkpuL0_1),.din(w_dff_A_ucWO2dQd1_1),.clk(gclk));
	jdff dff_A_RBuzc3PJ3_1(.dout(w_dff_A_ucWO2dQd1_1),.din(w_dff_A_RBuzc3PJ3_1),.clk(gclk));
	jdff dff_A_WE3vj2CX5_1(.dout(w_dff_A_RBuzc3PJ3_1),.din(w_dff_A_WE3vj2CX5_1),.clk(gclk));
	jdff dff_A_lyWdlucm2_1(.dout(w_dff_A_WE3vj2CX5_1),.din(w_dff_A_lyWdlucm2_1),.clk(gclk));
	jdff dff_A_ZQl9FZJa0_1(.dout(w_dff_A_lyWdlucm2_1),.din(w_dff_A_ZQl9FZJa0_1),.clk(gclk));
	jdff dff_B_xWGvZ6jQ1_0(.din(n1113),.dout(w_dff_B_xWGvZ6jQ1_0),.clk(gclk));
	jdff dff_B_ig3HG5L75_0(.din(w_dff_B_xWGvZ6jQ1_0),.dout(w_dff_B_ig3HG5L75_0),.clk(gclk));
	jdff dff_B_80ts38i57_0(.din(w_dff_B_ig3HG5L75_0),.dout(w_dff_B_80ts38i57_0),.clk(gclk));
	jdff dff_B_CjsrJNf85_0(.din(w_dff_B_80ts38i57_0),.dout(w_dff_B_CjsrJNf85_0),.clk(gclk));
	jdff dff_B_RtZjEUoh5_0(.din(w_dff_B_CjsrJNf85_0),.dout(w_dff_B_RtZjEUoh5_0),.clk(gclk));
	jdff dff_B_NAj0O6MK7_0(.din(w_dff_B_RtZjEUoh5_0),.dout(w_dff_B_NAj0O6MK7_0),.clk(gclk));
	jdff dff_B_ZBwqG1ji1_0(.din(w_dff_B_NAj0O6MK7_0),.dout(w_dff_B_ZBwqG1ji1_0),.clk(gclk));
	jdff dff_B_lJfyTnvH0_0(.din(n1109),.dout(w_dff_B_lJfyTnvH0_0),.clk(gclk));
	jdff dff_B_1uOPiDZv0_0(.din(w_dff_B_lJfyTnvH0_0),.dout(w_dff_B_1uOPiDZv0_0),.clk(gclk));
	jdff dff_B_MNfomTFq9_0(.din(w_dff_B_1uOPiDZv0_0),.dout(w_dff_B_MNfomTFq9_0),.clk(gclk));
	jdff dff_B_U8KLbiZe2_0(.din(w_dff_B_MNfomTFq9_0),.dout(w_dff_B_U8KLbiZe2_0),.clk(gclk));
	jdff dff_B_qNxgxsmg8_0(.din(w_dff_B_U8KLbiZe2_0),.dout(w_dff_B_qNxgxsmg8_0),.clk(gclk));
	jdff dff_B_BLEwuBJe3_0(.din(w_dff_B_qNxgxsmg8_0),.dout(w_dff_B_BLEwuBJe3_0),.clk(gclk));
	jdff dff_B_YoznAWsr8_0(.din(w_dff_B_BLEwuBJe3_0),.dout(w_dff_B_YoznAWsr8_0),.clk(gclk));
	jdff dff_B_Y1rcZzZB7_1(.din(n1070),.dout(w_dff_B_Y1rcZzZB7_1),.clk(gclk));
	jdff dff_B_LkeHFOvD2_1(.din(w_dff_B_Y1rcZzZB7_1),.dout(w_dff_B_LkeHFOvD2_1),.clk(gclk));
	jdff dff_B_6QTp5PQ74_1(.din(w_dff_B_LkeHFOvD2_1),.dout(w_dff_B_6QTp5PQ74_1),.clk(gclk));
	jdff dff_B_i8UZeDtG7_1(.din(w_dff_B_6QTp5PQ74_1),.dout(w_dff_B_i8UZeDtG7_1),.clk(gclk));
	jdff dff_B_tR9yNUqP8_1(.din(w_dff_B_i8UZeDtG7_1),.dout(w_dff_B_tR9yNUqP8_1),.clk(gclk));
	jdff dff_B_CSSbkLuy4_1(.din(w_dff_B_tR9yNUqP8_1),.dout(w_dff_B_CSSbkLuy4_1),.clk(gclk));
	jdff dff_B_pSvqTTRd7_1(.din(w_dff_B_CSSbkLuy4_1),.dout(w_dff_B_pSvqTTRd7_1),.clk(gclk));
	jdff dff_B_mBKeCzen2_1(.din(w_dff_B_pSvqTTRd7_1),.dout(w_dff_B_mBKeCzen2_1),.clk(gclk));
	jdff dff_B_oYNtwwoa6_1(.din(n1086),.dout(w_dff_B_oYNtwwoa6_1),.clk(gclk));
	jdff dff_B_5RuyAYUz8_1(.din(w_dff_B_oYNtwwoa6_1),.dout(w_dff_B_5RuyAYUz8_1),.clk(gclk));
	jdff dff_B_6IigKEW58_1(.din(n1094),.dout(w_dff_B_6IigKEW58_1),.clk(gclk));
	jdff dff_B_gUOa6haK3_0(.din(n1099),.dout(w_dff_B_gUOa6haK3_0),.clk(gclk));
	jdff dff_B_0idgkjQN3_1(.din(n1075),.dout(w_dff_B_0idgkjQN3_1),.clk(gclk));
	jdff dff_B_BK1PEsdO6_1(.din(w_dff_B_0idgkjQN3_1),.dout(w_dff_B_BK1PEsdO6_1),.clk(gclk));
	jdff dff_B_LgGx67mV7_0(.din(n1084),.dout(w_dff_B_LgGx67mV7_0),.clk(gclk));
	jdff dff_B_qQIrSnQJ5_1(.din(n1076),.dout(w_dff_B_qQIrSnQJ5_1),.clk(gclk));
	jdff dff_B_x85OuUaa8_0(.din(n1078),.dout(w_dff_B_x85OuUaa8_0),.clk(gclk));
	jdff dff_B_m4XxvndL2_1(.din(G124),.dout(w_dff_B_m4XxvndL2_1),.clk(gclk));
	jdff dff_B_Qxf9hIPF6_1(.din(w_dff_B_m4XxvndL2_1),.dout(w_dff_B_Qxf9hIPF6_1),.clk(gclk));
	jdff dff_B_H61T9q7t9_1(.din(w_dff_B_Qxf9hIPF6_1),.dout(w_dff_B_H61T9q7t9_1),.clk(gclk));
	jdff dff_B_RAbVov9X1_1(.din(w_dff_B_H61T9q7t9_1),.dout(w_dff_B_RAbVov9X1_1),.clk(gclk));
	jdff dff_B_cQ8DBxlb8_1(.din(n1071),.dout(w_dff_B_cQ8DBxlb8_1),.clk(gclk));
	jdff dff_B_pEDu6DlF5_0(.din(n1069),.dout(w_dff_B_pEDu6DlF5_0),.clk(gclk));
	jdff dff_B_kXRsGkfF4_0(.din(w_dff_B_pEDu6DlF5_0),.dout(w_dff_B_kXRsGkfF4_0),.clk(gclk));
	jdff dff_B_QoyuoMYs5_0(.din(w_dff_B_kXRsGkfF4_0),.dout(w_dff_B_QoyuoMYs5_0),.clk(gclk));
	jdff dff_B_wqi3mgeV4_1(.din(n1060),.dout(w_dff_B_wqi3mgeV4_1),.clk(gclk));
	jdff dff_A_HI2lnYjI5_1(.dout(w_n1062_0[1]),.din(w_dff_A_HI2lnYjI5_1),.clk(gclk));
	jdff dff_A_jLgJwv0p4_1(.dout(w_dff_A_HI2lnYjI5_1),.din(w_dff_A_jLgJwv0p4_1),.clk(gclk));
	jdff dff_A_nmBo6tOR0_1(.dout(w_dff_A_jLgJwv0p4_1),.din(w_dff_A_nmBo6tOR0_1),.clk(gclk));
	jdff dff_A_0rdu9bIW9_1(.dout(w_dff_A_nmBo6tOR0_1),.din(w_dff_A_0rdu9bIW9_1),.clk(gclk));
	jdff dff_A_Cr2CoSXm3_1(.dout(w_dff_A_0rdu9bIW9_1),.din(w_dff_A_Cr2CoSXm3_1),.clk(gclk));
	jdff dff_A_EpSeeTrY9_1(.dout(w_dff_A_Cr2CoSXm3_1),.din(w_dff_A_EpSeeTrY9_1),.clk(gclk));
	jdff dff_A_FKDTVBOb4_1(.dout(w_dff_A_EpSeeTrY9_1),.din(w_dff_A_FKDTVBOb4_1),.clk(gclk));
	jdff dff_A_siV6TsMS4_1(.dout(w_dff_A_FKDTVBOb4_1),.din(w_dff_A_siV6TsMS4_1),.clk(gclk));
	jdff dff_B_fosDWTk39_0(.din(n1061),.dout(w_dff_B_fosDWTk39_0),.clk(gclk));
	jdff dff_B_ZjAM4XCm8_0(.din(w_dff_B_fosDWTk39_0),.dout(w_dff_B_ZjAM4XCm8_0),.clk(gclk));
	jdff dff_B_GkoJ5LLd8_1(.din(n764),.dout(w_dff_B_GkoJ5LLd8_1),.clk(gclk));
	jdff dff_B_qN9kuMNm7_1(.din(w_dff_B_GkoJ5LLd8_1),.dout(w_dff_B_qN9kuMNm7_1),.clk(gclk));
	jdff dff_B_UajQjeRI7_1(.din(w_dff_B_qN9kuMNm7_1),.dout(w_dff_B_UajQjeRI7_1),.clk(gclk));
	jdff dff_B_677kXUgA3_1(.din(w_dff_B_UajQjeRI7_1),.dout(w_dff_B_677kXUgA3_1),.clk(gclk));
	jdff dff_B_z4YEo8u39_1(.din(w_dff_B_677kXUgA3_1),.dout(w_dff_B_z4YEo8u39_1),.clk(gclk));
	jdff dff_B_9j17tiSc0_1(.din(w_dff_B_z4YEo8u39_1),.dout(w_dff_B_9j17tiSc0_1),.clk(gclk));
	jdff dff_B_49cFV0nF6_1(.din(w_dff_B_9j17tiSc0_1),.dout(w_dff_B_49cFV0nF6_1),.clk(gclk));
	jdff dff_B_7Cxjwifc4_1(.din(w_dff_B_49cFV0nF6_1),.dout(w_dff_B_7Cxjwifc4_1),.clk(gclk));
	jdff dff_A_Lx5EfmK91_1(.dout(w_n767_1[1]),.din(w_dff_A_Lx5EfmK91_1),.clk(gclk));
	jdff dff_A_JfapGmZe9_1(.dout(w_dff_A_Lx5EfmK91_1),.din(w_dff_A_JfapGmZe9_1),.clk(gclk));
	jdff dff_A_K39VnRtC5_1(.dout(w_dff_A_JfapGmZe9_1),.din(w_dff_A_K39VnRtC5_1),.clk(gclk));
	jdff dff_B_c5F11mB04_0(.din(n763),.dout(w_dff_B_c5F11mB04_0),.clk(gclk));
	jdff dff_B_1OmdDj2w7_0(.din(w_dff_B_c5F11mB04_0),.dout(w_dff_B_1OmdDj2w7_0),.clk(gclk));
	jdff dff_B_wEulYuc23_0(.din(w_dff_B_1OmdDj2w7_0),.dout(w_dff_B_wEulYuc23_0),.clk(gclk));
	jdff dff_B_BQmU4Cyx9_0(.din(w_dff_B_wEulYuc23_0),.dout(w_dff_B_BQmU4Cyx9_0),.clk(gclk));
	jdff dff_B_EH72ZePG7_0(.din(w_dff_B_BQmU4Cyx9_0),.dout(w_dff_B_EH72ZePG7_0),.clk(gclk));
	jdff dff_B_QanFgOYD7_0(.din(w_dff_B_EH72ZePG7_0),.dout(w_dff_B_QanFgOYD7_0),.clk(gclk));
	jdff dff_B_zeMOrs7R0_0(.din(n1058),.dout(w_dff_B_zeMOrs7R0_0),.clk(gclk));
	jdff dff_B_w1V2tbQf1_1(.din(n1027),.dout(w_dff_B_w1V2tbQf1_1),.clk(gclk));
	jdff dff_B_jP4u0LC54_1(.din(w_dff_B_w1V2tbQf1_1),.dout(w_dff_B_jP4u0LC54_1),.clk(gclk));
	jdff dff_B_MpNgiRne8_1(.din(w_dff_B_jP4u0LC54_1),.dout(w_dff_B_MpNgiRne8_1),.clk(gclk));
	jdff dff_B_IxRQbdCt3_1(.din(w_dff_B_MpNgiRne8_1),.dout(w_dff_B_IxRQbdCt3_1),.clk(gclk));
	jdff dff_B_FPvrbdE18_1(.din(w_dff_B_IxRQbdCt3_1),.dout(w_dff_B_FPvrbdE18_1),.clk(gclk));
	jdff dff_B_IWf6MZfP4_1(.din(w_dff_B_FPvrbdE18_1),.dout(w_dff_B_IWf6MZfP4_1),.clk(gclk));
	jdff dff_B_Cdqyq45c9_1(.din(w_dff_B_IWf6MZfP4_1),.dout(w_dff_B_Cdqyq45c9_1),.clk(gclk));
	jdff dff_B_rMuyGdqc6_1(.din(w_dff_B_Cdqyq45c9_1),.dout(w_dff_B_rMuyGdqc6_1),.clk(gclk));
	jdff dff_B_fIWXbCll5_0(.din(n1051),.dout(w_dff_B_fIWXbCll5_0),.clk(gclk));
	jdff dff_A_FRgHQq6A9_1(.dout(w_n1045_0[1]),.din(w_dff_A_FRgHQq6A9_1),.clk(gclk));
	jdff dff_A_6YUtQTR05_1(.dout(w_dff_A_FRgHQq6A9_1),.din(w_dff_A_6YUtQTR05_1),.clk(gclk));
	jdff dff_B_eEPnibS64_1(.din(n769),.dout(w_dff_B_eEPnibS64_1),.clk(gclk));
	jdff dff_B_6lVSt8ed3_1(.din(w_dff_B_eEPnibS64_1),.dout(w_dff_B_6lVSt8ed3_1),.clk(gclk));
	jdff dff_A_TA13gUh84_1(.dout(w_n773_0[1]),.din(w_dff_A_TA13gUh84_1),.clk(gclk));
	jdff dff_A_kZIueL6h2_1(.dout(w_n767_0[1]),.din(w_dff_A_kZIueL6h2_1),.clk(gclk));
	jdff dff_A_NRLBxT1t3_1(.dout(w_dff_A_kZIueL6h2_1),.din(w_dff_A_NRLBxT1t3_1),.clk(gclk));
	jdff dff_A_EyzfIyiW1_1(.dout(w_dff_A_NRLBxT1t3_1),.din(w_dff_A_EyzfIyiW1_1),.clk(gclk));
	jdff dff_A_fdpzGfW16_1(.dout(w_dff_A_EyzfIyiW1_1),.din(w_dff_A_fdpzGfW16_1),.clk(gclk));
	jdff dff_A_YktNIekQ9_2(.dout(w_n767_0[2]),.din(w_dff_A_YktNIekQ9_2),.clk(gclk));
	jdff dff_A_Z9sBJwWm2_2(.dout(w_dff_A_YktNIekQ9_2),.din(w_dff_A_Z9sBJwWm2_2),.clk(gclk));
	jdff dff_A_rKBlyUaW6_2(.dout(w_dff_A_Z9sBJwWm2_2),.din(w_dff_A_rKBlyUaW6_2),.clk(gclk));
	jdff dff_B_oOwqTsSo4_3(.din(n767),.dout(w_dff_B_oOwqTsSo4_3),.clk(gclk));
	jdff dff_B_gWNyL8z93_3(.din(w_dff_B_oOwqTsSo4_3),.dout(w_dff_B_gWNyL8z93_3),.clk(gclk));
	jdff dff_A_pHISlmdY7_1(.dout(w_n1043_0[1]),.din(w_dff_A_pHISlmdY7_1),.clk(gclk));
	jdff dff_B_4I3jzZeY7_0(.din(n1025),.dout(w_dff_B_4I3jzZeY7_0),.clk(gclk));
	jdff dff_B_iiwKL2hO2_0(.din(n1023),.dout(w_dff_B_iiwKL2hO2_0),.clk(gclk));
	jdff dff_B_6bHBSDGV1_0(.din(w_dff_B_iiwKL2hO2_0),.dout(w_dff_B_6bHBSDGV1_0),.clk(gclk));
	jdff dff_B_BiuoirYW2_0(.din(w_dff_B_6bHBSDGV1_0),.dout(w_dff_B_BiuoirYW2_0),.clk(gclk));
	jdff dff_B_dlBr8R3K6_0(.din(w_dff_B_BiuoirYW2_0),.dout(w_dff_B_dlBr8R3K6_0),.clk(gclk));
	jdff dff_B_sjjFa77P5_0(.din(w_dff_B_dlBr8R3K6_0),.dout(w_dff_B_sjjFa77P5_0),.clk(gclk));
	jdff dff_B_mgULKXz23_1(.din(n1006),.dout(w_dff_B_mgULKXz23_1),.clk(gclk));
	jdff dff_B_XudOkgBB5_1(.din(n1010),.dout(w_dff_B_XudOkgBB5_1),.clk(gclk));
	jdff dff_B_Gl0g4FKD0_0(.din(n1015),.dout(w_dff_B_Gl0g4FKD0_0),.clk(gclk));
	jdff dff_B_fYOfFF587_1(.din(n1011),.dout(w_dff_B_fYOfFF587_1),.clk(gclk));
	jdff dff_B_zxYraqje1_1(.din(n1007),.dout(w_dff_B_zxYraqje1_1),.clk(gclk));
	jdff dff_B_wzqu9s0k8_1(.din(n998),.dout(w_dff_B_wzqu9s0k8_1),.clk(gclk));
	jdff dff_B_GZqDTNiB8_1(.din(n999),.dout(w_dff_B_GZqDTNiB8_1),.clk(gclk));
	jdff dff_B_zHp34f0p2_1(.din(w_dff_B_GZqDTNiB8_1),.dout(w_dff_B_zHp34f0p2_1),.clk(gclk));
	jdff dff_B_dv2uFe8e2_1(.din(w_dff_B_zHp34f0p2_1),.dout(w_dff_B_dv2uFe8e2_1),.clk(gclk));
	jdff dff_B_77O0B9s62_1(.din(n1000),.dout(w_dff_B_77O0B9s62_1),.clk(gclk));
	jdff dff_B_3LiZdvJa5_1(.din(w_dff_B_77O0B9s62_1),.dout(w_dff_B_3LiZdvJa5_1),.clk(gclk));
	jdff dff_B_ZSMIrfLb0_0(.din(n1002),.dout(w_dff_B_ZSMIrfLb0_0),.clk(gclk));
	jdff dff_B_Ijayki2N9_1(.din(n991),.dout(w_dff_B_Ijayki2N9_1),.clk(gclk));
	jdff dff_A_OAACL1iP1_1(.dout(w_G125_0[1]),.din(w_dff_A_OAACL1iP1_1),.clk(gclk));
	jdff dff_B_zerNUWn88_2(.din(G125),.dout(w_dff_B_zerNUWn88_2),.clk(gclk));
	jdff dff_B_r6X535Li1_2(.din(w_dff_B_zerNUWn88_2),.dout(w_dff_B_r6X535Li1_2),.clk(gclk));
	jdff dff_B_NXq1WUpR1_2(.din(w_dff_B_r6X535Li1_2),.dout(w_dff_B_NXq1WUpR1_2),.clk(gclk));
	jdff dff_A_30wqftnc0_0(.dout(w_n614_2[0]),.din(w_dff_A_30wqftnc0_0),.clk(gclk));
	jdff dff_A_CCYaXbSh6_0(.dout(w_dff_A_30wqftnc0_0),.din(w_dff_A_CCYaXbSh6_0),.clk(gclk));
	jdff dff_A_dLJ03ZvW5_0(.dout(w_dff_A_CCYaXbSh6_0),.din(w_dff_A_dLJ03ZvW5_0),.clk(gclk));
	jdff dff_A_a8uuI0z37_1(.dout(w_n614_2[1]),.din(w_dff_A_a8uuI0z37_1),.clk(gclk));
	jdff dff_A_N746gYgC1_1(.dout(w_dff_A_a8uuI0z37_1),.din(w_dff_A_N746gYgC1_1),.clk(gclk));
	jdff dff_A_cTD5tyEA5_1(.dout(w_dff_A_N746gYgC1_1),.din(w_dff_A_cTD5tyEA5_1),.clk(gclk));
	jdff dff_A_FMSR0ZCj0_1(.dout(w_dff_A_cTD5tyEA5_1),.din(w_dff_A_FMSR0ZCj0_1),.clk(gclk));
	jdff dff_A_I4CaDGW37_1(.dout(w_dff_A_FMSR0ZCj0_1),.din(w_dff_A_I4CaDGW37_1),.clk(gclk));
	jdff dff_A_kVQKTSbv0_1(.dout(w_dff_A_I4CaDGW37_1),.din(w_dff_A_kVQKTSbv0_1),.clk(gclk));
	jdff dff_A_rdz1rvvg2_1(.dout(w_dff_A_kVQKTSbv0_1),.din(w_dff_A_rdz1rvvg2_1),.clk(gclk));
	jdff dff_A_fXYDABUs7_1(.dout(w_dff_A_rdz1rvvg2_1),.din(w_dff_A_fXYDABUs7_1),.clk(gclk));
	jdff dff_A_YHZ9rSjz4_1(.dout(w_dff_A_fXYDABUs7_1),.din(w_dff_A_YHZ9rSjz4_1),.clk(gclk));
	jdff dff_A_8oeDgHHV2_1(.dout(w_dff_A_YHZ9rSjz4_1),.din(w_dff_A_8oeDgHHV2_1),.clk(gclk));
	jdff dff_A_POL1wn4v6_1(.dout(w_dff_A_8oeDgHHV2_1),.din(w_dff_A_POL1wn4v6_1),.clk(gclk));
	jdff dff_B_1QEF5TMg9_0(.din(n765),.dout(w_dff_B_1QEF5TMg9_0),.clk(gclk));
	jdff dff_B_Y3vRi9GH1_0(.din(w_dff_B_1QEF5TMg9_0),.dout(w_dff_B_Y3vRi9GH1_0),.clk(gclk));
	jdff dff_B_36qOmuvW2_1(.din(n1154),.dout(w_dff_B_36qOmuvW2_1),.clk(gclk));
	jdff dff_B_VHTaDOFl1_1(.din(w_dff_B_36qOmuvW2_1),.dout(w_dff_B_VHTaDOFl1_1),.clk(gclk));
	jdff dff_B_zvs1keRG1_1(.din(w_dff_B_VHTaDOFl1_1),.dout(w_dff_B_zvs1keRG1_1),.clk(gclk));
	jdff dff_B_n8p0L0ug4_1(.din(w_dff_B_zvs1keRG1_1),.dout(w_dff_B_n8p0L0ug4_1),.clk(gclk));
	jdff dff_B_FdkCw2n75_1(.din(w_dff_B_n8p0L0ug4_1),.dout(w_dff_B_FdkCw2n75_1),.clk(gclk));
	jdff dff_B_LHKZR8h56_1(.din(w_dff_B_FdkCw2n75_1),.dout(w_dff_B_LHKZR8h56_1),.clk(gclk));
	jdff dff_B_3mkVTSnB2_0(.din(n1157),.dout(w_dff_B_3mkVTSnB2_0),.clk(gclk));
	jdff dff_B_kjZSD6wT0_1(.din(n1156),.dout(w_dff_B_kjZSD6wT0_1),.clk(gclk));
	jdff dff_B_ukbYK3mL7_0(.din(n1028),.dout(w_dff_B_ukbYK3mL7_0),.clk(gclk));
	jdff dff_A_MvoiZR3U7_0(.dout(w_n514_1[0]),.din(w_dff_A_MvoiZR3U7_0),.clk(gclk));
	jdff dff_A_EGrOcpeG1_1(.dout(w_n514_0[1]),.din(w_dff_A_EGrOcpeG1_1),.clk(gclk));
	jdff dff_A_hhoYO9hg9_1(.dout(w_dff_A_EGrOcpeG1_1),.din(w_dff_A_hhoYO9hg9_1),.clk(gclk));
	jdff dff_A_HT9a3MaW1_2(.dout(w_n514_0[2]),.din(w_dff_A_HT9a3MaW1_2),.clk(gclk));
	jdff dff_A_v1McfurO5_2(.dout(w_dff_A_HT9a3MaW1_2),.din(w_dff_A_v1McfurO5_2),.clk(gclk));
	jdff dff_A_FRkws6Vl4_0(.dout(w_n562_0[0]),.din(w_dff_A_FRkws6Vl4_0),.clk(gclk));
	jdff dff_B_vix8ijZT3_1(.din(n555),.dout(w_dff_B_vix8ijZT3_1),.clk(gclk));
	jdff dff_B_d2AqgI6h4_1(.din(w_dff_B_vix8ijZT3_1),.dout(w_dff_B_d2AqgI6h4_1),.clk(gclk));
	jdff dff_B_t9FRZKtK5_1(.din(n556),.dout(w_dff_B_t9FRZKtK5_1),.clk(gclk));
	jdff dff_B_RJARQDl49_1(.din(w_dff_B_t9FRZKtK5_1),.dout(w_dff_B_RJARQDl49_1),.clk(gclk));
	jdff dff_B_xhe3WgjF4_1(.din(w_dff_B_RJARQDl49_1),.dout(w_dff_B_xhe3WgjF4_1),.clk(gclk));
	jdff dff_B_AibjIE2U8_1(.din(n557),.dout(w_dff_B_AibjIE2U8_1),.clk(gclk));
	jdff dff_A_iTgn9Xz62_0(.dout(w_n512_0[0]),.din(w_dff_A_iTgn9Xz62_0),.clk(gclk));
	jdff dff_B_K4FHGxx43_1(.din(n440),.dout(w_dff_B_K4FHGxx43_1),.clk(gclk));
	jdff dff_A_DNdT5Ak99_1(.dout(w_n503_0[1]),.din(w_dff_A_DNdT5Ak99_1),.clk(gclk));
	jdff dff_A_HCXleRxp7_1(.dout(w_n499_0[1]),.din(w_dff_A_HCXleRxp7_1),.clk(gclk));
	jdff dff_A_KV5z3AXq7_1(.dout(w_n74_1[1]),.din(w_dff_A_KV5z3AXq7_1),.clk(gclk));
	jdff dff_A_OxPTfjlh4_1(.dout(w_dff_A_KV5z3AXq7_1),.din(w_dff_A_OxPTfjlh4_1),.clk(gclk));
	jdff dff_A_bFCQX2iL3_1(.dout(w_dff_A_OxPTfjlh4_1),.din(w_dff_A_bFCQX2iL3_1),.clk(gclk));
	jdff dff_A_eaHt07N52_1(.dout(w_dff_A_bFCQX2iL3_1),.din(w_dff_A_eaHt07N52_1),.clk(gclk));
	jdff dff_A_BGJNNgD99_2(.dout(w_n74_1[2]),.din(w_dff_A_BGJNNgD99_2),.clk(gclk));
	jdff dff_A_JaMkopz46_2(.dout(w_dff_A_BGJNNgD99_2),.din(w_dff_A_JaMkopz46_2),.clk(gclk));
	jdff dff_A_Cx0w8QtE6_2(.dout(w_dff_A_JaMkopz46_2),.din(w_dff_A_Cx0w8QtE6_2),.clk(gclk));
	jdff dff_A_3GyNeKS69_0(.dout(w_n494_0[0]),.din(w_dff_A_3GyNeKS69_0),.clk(gclk));
	jdff dff_B_61EjpAtY1_1(.din(n487),.dout(w_dff_B_61EjpAtY1_1),.clk(gclk));
	jdff dff_B_0SZdy8yD4_1(.din(n489),.dout(w_dff_B_0SZdy8yD4_1),.clk(gclk));
	jdff dff_B_XwAHOEav0_1(.din(w_dff_B_0SZdy8yD4_1),.dout(w_dff_B_XwAHOEav0_1),.clk(gclk));
	jdff dff_B_Ubi5PWTg3_1(.din(n485),.dout(w_dff_B_Ubi5PWTg3_1),.clk(gclk));
	jdff dff_B_vkJ7ryfr0_1(.din(w_dff_B_Ubi5PWTg3_1),.dout(w_dff_B_vkJ7ryfr0_1),.clk(gclk));
	jdff dff_B_CqwipQjJ2_1(.din(n475),.dout(w_dff_B_CqwipQjJ2_1),.clk(gclk));
	jdff dff_B_uIKuRZbo0_1(.din(w_dff_B_CqwipQjJ2_1),.dout(w_dff_B_uIKuRZbo0_1),.clk(gclk));
	jdff dff_B_kJhu1W4f8_1(.din(n476),.dout(w_dff_B_kJhu1W4f8_1),.clk(gclk));
	jdff dff_A_Ydbojq200_1(.dout(w_n456_0[1]),.din(w_dff_A_Ydbojq200_1),.clk(gclk));
	jdff dff_A_NCw5ISe29_0(.dout(w_n450_0[0]),.din(w_dff_A_NCw5ISe29_0),.clk(gclk));
	jdff dff_B_EV0oZ51Q6_1(.din(n443),.dout(w_dff_B_EV0oZ51Q6_1),.clk(gclk));
	jdff dff_A_fM9TVJlP3_0(.dout(w_n73_2[0]),.din(w_dff_A_fM9TVJlP3_0),.clk(gclk));
	jdff dff_A_4toUY6Qz0_0(.dout(w_dff_A_fM9TVJlP3_0),.din(w_dff_A_4toUY6Qz0_0),.clk(gclk));
	jdff dff_A_d5tGjkKH7_0(.dout(w_dff_A_4toUY6Qz0_0),.din(w_dff_A_d5tGjkKH7_0),.clk(gclk));
	jdff dff_A_SGTn5YJd4_2(.dout(w_n73_2[2]),.din(w_dff_A_SGTn5YJd4_2),.clk(gclk));
	jdff dff_A_PqZgsTd56_2(.dout(w_n151_3[2]),.din(w_dff_A_PqZgsTd56_2),.clk(gclk));
	jdff dff_A_8lVb8cug4_2(.dout(w_dff_A_PqZgsTd56_2),.din(w_dff_A_8lVb8cug4_2),.clk(gclk));
	jdff dff_B_2nIrxPWo3_1(.din(n429),.dout(w_dff_B_2nIrxPWo3_1),.clk(gclk));
	jdff dff_A_b7shwyO36_1(.dout(w_n435_0[1]),.din(w_dff_A_b7shwyO36_1),.clk(gclk));
	jdff dff_A_c23foJsE2_0(.dout(w_n430_0[0]),.din(w_dff_A_c23foJsE2_0),.clk(gclk));
	jdff dff_B_bbh4JCIm1_2(.din(G223),.dout(w_dff_B_bbh4JCIm1_2),.clk(gclk));
	jdff dff_B_F2IAu7YI9_2(.din(w_dff_B_bbh4JCIm1_2),.dout(w_dff_B_F2IAu7YI9_2),.clk(gclk));
	jdff dff_A_4YrgVHni8_0(.dout(w_n428_0[0]),.din(w_dff_A_4YrgVHni8_0),.clk(gclk));
	jdff dff_A_RFNPLB650_0(.dout(w_dff_A_4YrgVHni8_0),.din(w_dff_A_RFNPLB650_0),.clk(gclk));
	jdff dff_A_XhzSou9P1_0(.dout(w_n1056_0[0]),.din(w_dff_A_XhzSou9P1_0),.clk(gclk));
	jdff dff_A_EwJdGVxo2_0(.dout(w_dff_A_XhzSou9P1_0),.din(w_dff_A_EwJdGVxo2_0),.clk(gclk));
	jdff dff_B_AjqoEEW30_2(.din(n1056),.dout(w_dff_B_AjqoEEW30_2),.clk(gclk));
	jdff dff_A_5vTYak7O9_1(.dout(w_n351_0[1]),.din(w_dff_A_5vTYak7O9_1),.clk(gclk));
	jdff dff_A_9305tNKF3_0(.dout(w_n772_0[0]),.din(w_dff_A_9305tNKF3_0),.clk(gclk));
	jdff dff_A_Zmg066ZD5_0(.dout(w_dff_A_9305tNKF3_0),.din(w_dff_A_Zmg066ZD5_0),.clk(gclk));
	jdff dff_A_KNoPRY6W5_0(.dout(w_dff_A_Zmg066ZD5_0),.din(w_dff_A_KNoPRY6W5_0),.clk(gclk));
	jdff dff_A_7JEsw6sy5_0(.dout(w_n771_1[0]),.din(w_dff_A_7JEsw6sy5_0),.clk(gclk));
	jdff dff_A_mXsJ5cto9_0(.dout(w_dff_A_7JEsw6sy5_0),.din(w_dff_A_mXsJ5cto9_0),.clk(gclk));
	jdff dff_A_89d5J4bx4_0(.dout(w_dff_A_mXsJ5cto9_0),.din(w_dff_A_89d5J4bx4_0),.clk(gclk));
	jdff dff_A_SWu8eWN90_0(.dout(w_dff_A_89d5J4bx4_0),.din(w_dff_A_SWu8eWN90_0),.clk(gclk));
	jdff dff_B_5VUEyggF9_0(.din(n1032),.dout(w_dff_B_5VUEyggF9_0),.clk(gclk));
	jdff dff_B_0AwsjEXO5_0(.din(w_dff_B_5VUEyggF9_0),.dout(w_dff_B_0AwsjEXO5_0),.clk(gclk));
	jdff dff_B_5q9U8p1K7_0(.din(w_dff_B_0AwsjEXO5_0),.dout(w_dff_B_5q9U8p1K7_0),.clk(gclk));
	jdff dff_B_2zIANsAj2_0(.din(n1151),.dout(w_dff_B_2zIANsAj2_0),.clk(gclk));
	jdff dff_B_BwhTBNMm1_0(.din(w_dff_B_2zIANsAj2_0),.dout(w_dff_B_BwhTBNMm1_0),.clk(gclk));
	jdff dff_B_48tfzXcl0_0(.din(w_dff_B_BwhTBNMm1_0),.dout(w_dff_B_48tfzXcl0_0),.clk(gclk));
	jdff dff_B_psmvs0JI6_0(.din(n1150),.dout(w_dff_B_psmvs0JI6_0),.clk(gclk));
	jdff dff_B_lT5Ns2Yr0_0(.din(w_dff_B_psmvs0JI6_0),.dout(w_dff_B_lT5Ns2Yr0_0),.clk(gclk));
	jdff dff_B_4HbUW6mA5_0(.din(w_dff_B_lT5Ns2Yr0_0),.dout(w_dff_B_4HbUW6mA5_0),.clk(gclk));
	jdff dff_B_pPIEZ9EV1_0(.din(w_dff_B_4HbUW6mA5_0),.dout(w_dff_B_pPIEZ9EV1_0),.clk(gclk));
	jdff dff_B_LQeloxLE6_0(.din(w_dff_B_pPIEZ9EV1_0),.dout(w_dff_B_LQeloxLE6_0),.clk(gclk));
	jdff dff_B_eaKMHYqK0_1(.din(n1131),.dout(w_dff_B_eaKMHYqK0_1),.clk(gclk));
	jdff dff_B_NlD4pxdV4_1(.din(w_dff_B_eaKMHYqK0_1),.dout(w_dff_B_NlD4pxdV4_1),.clk(gclk));
	jdff dff_B_pds4Bk8m8_1(.din(n1132),.dout(w_dff_B_pds4Bk8m8_1),.clk(gclk));
	jdff dff_B_F4vkc31U9_1(.din(w_dff_B_pds4Bk8m8_1),.dout(w_dff_B_F4vkc31U9_1),.clk(gclk));
	jdff dff_B_wKM8UG592_1(.din(w_dff_B_F4vkc31U9_1),.dout(w_dff_B_wKM8UG592_1),.clk(gclk));
	jdff dff_B_sE2vD7Q96_1(.din(w_dff_B_wKM8UG592_1),.dout(w_dff_B_sE2vD7Q96_1),.clk(gclk));
	jdff dff_B_mKbZNNwd7_1(.din(w_dff_B_sE2vD7Q96_1),.dout(w_dff_B_mKbZNNwd7_1),.clk(gclk));
	jdff dff_B_oazDjgne2_1(.din(n1135),.dout(w_dff_B_oazDjgne2_1),.clk(gclk));
	jdff dff_B_D74Jixrd2_1(.din(w_dff_B_oazDjgne2_1),.dout(w_dff_B_D74Jixrd2_1),.clk(gclk));
	jdff dff_B_TQMJOALO8_1(.din(w_dff_B_D74Jixrd2_1),.dout(w_dff_B_TQMJOALO8_1),.clk(gclk));
	jdff dff_B_mdsd82Yu5_1(.din(n1140),.dout(w_dff_B_mdsd82Yu5_1),.clk(gclk));
	jdff dff_A_UshgANoK0_0(.dout(w_G128_0[0]),.din(w_dff_A_UshgANoK0_0),.clk(gclk));
	jdff dff_B_J67n9Fgl9_3(.din(G128),.dout(w_dff_B_J67n9Fgl9_3),.clk(gclk));
	jdff dff_B_yr1c9DKG0_3(.din(w_dff_B_J67n9Fgl9_3),.dout(w_dff_B_yr1c9DKG0_3),.clk(gclk));
	jdff dff_B_5uutoYik1_3(.din(w_dff_B_yr1c9DKG0_3),.dout(w_dff_B_5uutoYik1_3),.clk(gclk));
	jdff dff_A_6WtM1vEI3_0(.dout(w_G33_4[0]),.din(w_dff_A_6WtM1vEI3_0),.clk(gclk));
	jdff dff_A_H3r4BdW72_1(.dout(w_G33_4[1]),.din(w_dff_A_H3r4BdW72_1),.clk(gclk));
	jdff dff_A_9GG5FGtY4_1(.dout(w_dff_A_H3r4BdW72_1),.din(w_dff_A_9GG5FGtY4_1),.clk(gclk));
	jdff dff_A_8hjcKo8F0_1(.dout(w_dff_A_9GG5FGtY4_1),.din(w_dff_A_8hjcKo8F0_1),.clk(gclk));
	jdff dff_A_0zdnIMgX1_1(.dout(w_dff_A_8hjcKo8F0_1),.din(w_dff_A_0zdnIMgX1_1),.clk(gclk));
	jdff dff_B_26OSP5554_1(.din(n1136),.dout(w_dff_B_26OSP5554_1),.clk(gclk));
	jdff dff_B_vMDHdvrG4_1(.din(w_dff_B_26OSP5554_1),.dout(w_dff_B_vMDHdvrG4_1),.clk(gclk));
	jdff dff_A_9reIYKkx5_0(.dout(w_n1091_0[0]),.din(w_dff_A_9reIYKkx5_0),.clk(gclk));
	jdff dff_A_vt49kmHw4_1(.dout(w_G150_1[1]),.din(w_dff_A_vt49kmHw4_1),.clk(gclk));
	jdff dff_A_2Jr8D4s51_2(.dout(w_G159_1[2]),.din(w_dff_A_2Jr8D4s51_2),.clk(gclk));
	jdff dff_B_HwTHqegq0_1(.din(n1118),.dout(w_dff_B_HwTHqegq0_1),.clk(gclk));
	jdff dff_B_xpsKkW372_1(.din(w_dff_B_HwTHqegq0_1),.dout(w_dff_B_xpsKkW372_1),.clk(gclk));
	jdff dff_A_b6RVrugm3_1(.dout(w_G283_1[1]),.din(w_dff_A_b6RVrugm3_1),.clk(gclk));
	jdff dff_A_7pDiKzB21_2(.dout(w_n771_0[2]),.din(w_dff_A_7pDiKzB21_2),.clk(gclk));
	jdff dff_A_yblqBuNC5_2(.dout(w_dff_A_7pDiKzB21_2),.din(w_dff_A_yblqBuNC5_2),.clk(gclk));
	jdff dff_A_avRL46u46_2(.dout(w_dff_A_yblqBuNC5_2),.din(w_dff_A_avRL46u46_2),.clk(gclk));
	jdff dff_A_1d6IbwNh2_2(.dout(w_dff_A_avRL46u46_2),.din(w_dff_A_1d6IbwNh2_2),.clk(gclk));
	jdff dff_B_Opz9X0i83_0(.din(n770),.dout(w_dff_B_Opz9X0i83_0),.clk(gclk));
	jdff dff_B_10PqCySC3_0(.din(w_dff_B_Opz9X0i83_0),.dout(w_dff_B_10PqCySC3_0),.clk(gclk));
	jdff dff_B_CYWKAXAg8_0(.din(w_dff_B_10PqCySC3_0),.dout(w_dff_B_CYWKAXAg8_0),.clk(gclk));
	jdff dff_B_toa3xpjP1_0(.din(w_dff_B_CYWKAXAg8_0),.dout(w_dff_B_toa3xpjP1_0),.clk(gclk));
	jdff dff_A_T8uo1aQq5_1(.dout(w_n420_0[1]),.din(w_dff_A_T8uo1aQq5_1),.clk(gclk));
	jdff dff_A_Xi4JRTa49_1(.dout(w_n417_0[1]),.din(w_dff_A_Xi4JRTa49_1),.clk(gclk));
	jdff dff_A_vcxg1qYh8_2(.dout(w_n417_0[2]),.din(w_dff_A_vcxg1qYh8_2),.clk(gclk));
	jdff dff_B_rECt16696_1(.din(n411),.dout(w_dff_B_rECt16696_1),.clk(gclk));
	jdff dff_B_ss6wQMSM1_1(.din(w_dff_B_rECt16696_1),.dout(w_dff_B_ss6wQMSM1_1),.clk(gclk));
	jdff dff_B_eRaeAqzx5_1(.din(n413),.dout(w_dff_B_eRaeAqzx5_1),.clk(gclk));
	jdff dff_B_REqKySol5_1(.din(w_dff_B_eRaeAqzx5_1),.dout(w_dff_B_REqKySol5_1),.clk(gclk));
	jdff dff_A_awADi5dy0_0(.dout(w_G68_4[0]),.din(w_dff_A_awADi5dy0_0),.clk(gclk));
	jdff dff_A_DRU23pch3_0(.dout(w_dff_A_awADi5dy0_0),.din(w_dff_A_DRU23pch3_0),.clk(gclk));
	jdff dff_A_ErTh8wLX2_2(.dout(w_G68_4[2]),.din(w_dff_A_ErTh8wLX2_2),.clk(gclk));
	jdff dff_A_QR5cJbr74_2(.dout(w_dff_A_ErTh8wLX2_2),.din(w_dff_A_QR5cJbr74_2),.clk(gclk));
	jdff dff_A_MadWnhvV5_2(.dout(w_dff_A_QR5cJbr74_2),.din(w_dff_A_MadWnhvV5_2),.clk(gclk));
	jdff dff_A_yLA6kELO7_2(.dout(w_dff_A_MadWnhvV5_2),.din(w_dff_A_yLA6kELO7_2),.clk(gclk));
	jdff dff_A_9NFBB2sh2_2(.dout(w_dff_A_yLA6kELO7_2),.din(w_dff_A_9NFBB2sh2_2),.clk(gclk));
	jdff dff_B_cQDb0x8w8_0(.din(n412),.dout(w_dff_B_cQDb0x8w8_0),.clk(gclk));
	jdff dff_A_Td2GGZBJ4_1(.dout(w_n407_0[1]),.din(w_dff_A_Td2GGZBJ4_1),.clk(gclk));
	jdff dff_B_WSAyDDDI9_1(.din(n397),.dout(w_dff_B_WSAyDDDI9_1),.clk(gclk));
	jdff dff_B_A0x9HqyM7_1(.din(w_dff_B_WSAyDDDI9_1),.dout(w_dff_B_A0x9HqyM7_1),.clk(gclk));
	jdff dff_B_yaVOpD0p0_1(.din(n398),.dout(w_dff_B_yaVOpD0p0_1),.clk(gclk));
	jdff dff_A_Cf3iR7zw1_0(.dout(w_n168_2[0]),.din(w_dff_A_Cf3iR7zw1_0),.clk(gclk));
	jdff dff_A_IfVgLIMX6_0(.dout(w_dff_A_Cf3iR7zw1_0),.din(w_dff_A_IfVgLIMX6_0),.clk(gclk));
	jdff dff_A_kk0bhBUK1_0(.dout(w_G384_0),.din(w_dff_A_kk0bhBUK1_0),.clk(gclk));
	jdff dff_A_CEzkFtCv3_0(.dout(w_dff_A_kk0bhBUK1_0),.din(w_dff_A_CEzkFtCv3_0),.clk(gclk));
	jdff dff_A_KkTi9hGO7_0(.dout(w_dff_A_CEzkFtCv3_0),.din(w_dff_A_KkTi9hGO7_0),.clk(gclk));
	jdff dff_A_72xvU02r3_0(.dout(w_n759_0[0]),.din(w_dff_A_72xvU02r3_0),.clk(gclk));
	jdff dff_A_PF283EE86_0(.dout(w_dff_A_72xvU02r3_0),.din(w_dff_A_PF283EE86_0),.clk(gclk));
	jdff dff_A_H0XydCmF2_0(.dout(w_dff_A_PF283EE86_0),.din(w_dff_A_H0XydCmF2_0),.clk(gclk));
	jdff dff_A_ZZIjx8KE4_0(.dout(w_dff_A_H0XydCmF2_0),.din(w_dff_A_ZZIjx8KE4_0),.clk(gclk));
	jdff dff_B_Xt38zowO9_1(.din(n747),.dout(w_dff_B_Xt38zowO9_1),.clk(gclk));
	jdff dff_B_VnAYDJq25_1(.din(w_dff_B_Xt38zowO9_1),.dout(w_dff_B_VnAYDJq25_1),.clk(gclk));
	jdff dff_B_b6ipeSB23_0(.din(n751),.dout(w_dff_B_b6ipeSB23_0),.clk(gclk));
	jdff dff_B_wffm9AH96_1(.din(n296),.dout(w_dff_B_wffm9AH96_1),.clk(gclk));
	jdff dff_A_RtYubszG9_0(.dout(w_n395_0[0]),.din(w_dff_A_RtYubszG9_0),.clk(gclk));
	jdff dff_A_VN574AsW8_0(.dout(w_dff_A_RtYubszG9_0),.din(w_dff_A_VN574AsW8_0),.clk(gclk));
	jdff dff_A_aPNn3EpD9_0(.dout(w_dff_A_VN574AsW8_0),.din(w_dff_A_aPNn3EpD9_0),.clk(gclk));
	jdff dff_B_9JCi7FQT0_0(.din(n745),.dout(w_dff_B_9JCi7FQT0_0),.clk(gclk));
	jdff dff_B_WxuNFnKF1_0(.din(w_dff_B_9JCi7FQT0_0),.dout(w_dff_B_WxuNFnKF1_0),.clk(gclk));
	jdff dff_B_AGGp1nRs5_0(.din(w_dff_B_WxuNFnKF1_0),.dout(w_dff_B_AGGp1nRs5_0),.clk(gclk));
	jdff dff_B_UN52YtQS4_0(.din(w_dff_B_AGGp1nRs5_0),.dout(w_dff_B_UN52YtQS4_0),.clk(gclk));
	jdff dff_B_vWa9fJa06_0(.din(n743),.dout(w_dff_B_vWa9fJa06_0),.clk(gclk));
	jdff dff_B_YwhNRbe39_0(.din(w_dff_B_vWa9fJa06_0),.dout(w_dff_B_YwhNRbe39_0),.clk(gclk));
	jdff dff_B_zPEJRzuL7_0(.din(w_dff_B_YwhNRbe39_0),.dout(w_dff_B_zPEJRzuL7_0),.clk(gclk));
	jdff dff_B_GFUvPOFf8_0(.din(w_dff_B_zPEJRzuL7_0),.dout(w_dff_B_GFUvPOFf8_0),.clk(gclk));
	jdff dff_B_XYEEje5n4_1(.din(n740),.dout(w_dff_B_XYEEje5n4_1),.clk(gclk));
	jdff dff_A_Rh403l8r6_0(.dout(w_n618_1[0]),.din(w_dff_A_Rh403l8r6_0),.clk(gclk));
	jdff dff_A_vaJNcwWB3_0(.dout(w_dff_A_Rh403l8r6_0),.din(w_dff_A_vaJNcwWB3_0),.clk(gclk));
	jdff dff_A_5Ty3TnsM0_0(.dout(w_dff_A_vaJNcwWB3_0),.din(w_dff_A_5Ty3TnsM0_0),.clk(gclk));
	jdff dff_A_2AzRzcU75_0(.dout(w_dff_A_5Ty3TnsM0_0),.din(w_dff_A_2AzRzcU75_0),.clk(gclk));
	jdff dff_A_vW7RpPeh6_0(.dout(w_dff_A_2AzRzcU75_0),.din(w_dff_A_vW7RpPeh6_0),.clk(gclk));
	jdff dff_A_Uldg6yWl3_0(.dout(w_dff_A_vW7RpPeh6_0),.din(w_dff_A_Uldg6yWl3_0),.clk(gclk));
	jdff dff_A_ZrG1LffZ7_0(.dout(w_dff_A_Uldg6yWl3_0),.din(w_dff_A_ZrG1LffZ7_0),.clk(gclk));
	jdff dff_A_AkhiEvVQ8_0(.dout(w_dff_A_ZrG1LffZ7_0),.din(w_dff_A_AkhiEvVQ8_0),.clk(gclk));
	jdff dff_A_9Co6SrCG3_0(.dout(w_dff_A_AkhiEvVQ8_0),.din(w_dff_A_9Co6SrCG3_0),.clk(gclk));
	jdff dff_A_yo2xpoMC5_0(.dout(w_dff_A_9Co6SrCG3_0),.din(w_dff_A_yo2xpoMC5_0),.clk(gclk));
	jdff dff_A_ocxPA7mX1_0(.dout(w_dff_A_yo2xpoMC5_0),.din(w_dff_A_ocxPA7mX1_0),.clk(gclk));
	jdff dff_A_tS7MsuFi0_1(.dout(w_n618_1[1]),.din(w_dff_A_tS7MsuFi0_1),.clk(gclk));
	jdff dff_A_AA3gEA2K1_1(.dout(w_dff_A_tS7MsuFi0_1),.din(w_dff_A_AA3gEA2K1_1),.clk(gclk));
	jdff dff_A_NH8R1pZz6_1(.dout(w_dff_A_AA3gEA2K1_1),.din(w_dff_A_NH8R1pZz6_1),.clk(gclk));
	jdff dff_A_Moh5KKKy7_1(.dout(w_dff_A_NH8R1pZz6_1),.din(w_dff_A_Moh5KKKy7_1),.clk(gclk));
	jdff dff_A_ydAqYyKh0_1(.dout(w_dff_A_Moh5KKKy7_1),.din(w_dff_A_ydAqYyKh0_1),.clk(gclk));
	jdff dff_A_PCx2iXYg6_1(.dout(w_dff_A_ydAqYyKh0_1),.din(w_dff_A_PCx2iXYg6_1),.clk(gclk));
	jdff dff_A_w8cy5tjY3_1(.dout(w_dff_A_PCx2iXYg6_1),.din(w_dff_A_w8cy5tjY3_1),.clk(gclk));
	jdff dff_A_GhLDPFKD8_1(.dout(w_dff_A_w8cy5tjY3_1),.din(w_dff_A_GhLDPFKD8_1),.clk(gclk));
	jdff dff_A_VJgypklu9_1(.dout(w_dff_A_GhLDPFKD8_1),.din(w_dff_A_VJgypklu9_1),.clk(gclk));
	jdff dff_A_TePc5rIr7_1(.dout(w_dff_A_VJgypklu9_1),.din(w_dff_A_TePc5rIr7_1),.clk(gclk));
	jdff dff_A_1psSUxf49_1(.dout(w_dff_A_TePc5rIr7_1),.din(w_dff_A_1psSUxf49_1),.clk(gclk));
	jdff dff_B_5F7UX6Mj8_0(.din(n735),.dout(w_dff_B_5F7UX6Mj8_0),.clk(gclk));
	jdff dff_B_hfXWDO4K3_0(.din(n726),.dout(w_dff_B_hfXWDO4K3_0),.clk(gclk));
	jdff dff_B_rFZsDiXU3_1(.din(n723),.dout(w_dff_B_rFZsDiXU3_1),.clk(gclk));
	jdff dff_B_Ien3t5Ck6_1(.din(n713),.dout(w_dff_B_Ien3t5Ck6_1),.clk(gclk));
	jdff dff_B_0km3CmbJ7_1(.din(n716),.dout(w_dff_B_0km3CmbJ7_1),.clk(gclk));
	jdff dff_A_zU3v8NVp9_0(.dout(w_n718_0[0]),.din(w_dff_A_zU3v8NVp9_0),.clk(gclk));
	jdff dff_A_E8QLvYZR7_0(.dout(w_dff_A_zU3v8NVp9_0),.din(w_dff_A_E8QLvYZR7_0),.clk(gclk));
	jdff dff_A_j65Yf79E8_0(.dout(w_dff_A_E8QLvYZR7_0),.din(w_dff_A_j65Yf79E8_0),.clk(gclk));
	jdff dff_A_rKyVvHD16_0(.dout(w_dff_A_j65Yf79E8_0),.din(w_dff_A_rKyVvHD16_0),.clk(gclk));
	jdff dff_B_ksfw1szy2_2(.din(n718),.dout(w_dff_B_ksfw1szy2_2),.clk(gclk));
	jdff dff_B_Ct5oodQI2_1(.din(n714),.dout(w_dff_B_Ct5oodQI2_1),.clk(gclk));
	jdff dff_A_uvenekGE3_1(.dout(w_G132_1[1]),.din(w_dff_A_uvenekGE3_1),.clk(gclk));
	jdff dff_B_hDRpT2tv7_3(.din(G132),.dout(w_dff_B_hDRpT2tv7_3),.clk(gclk));
	jdff dff_B_yS6MQTAQ7_3(.din(w_dff_B_hDRpT2tv7_3),.dout(w_dff_B_yS6MQTAQ7_3),.clk(gclk));
	jdff dff_B_UP0PQyuR2_3(.din(w_dff_B_yS6MQTAQ7_3),.dout(w_dff_B_UP0PQyuR2_3),.clk(gclk));
	jdff dff_B_GzK86MKc0_1(.din(n707),.dout(w_dff_B_GzK86MKc0_1),.clk(gclk));
	jdff dff_B_SFYn7sTX4_1(.din(w_dff_B_GzK86MKc0_1),.dout(w_dff_B_SFYn7sTX4_1),.clk(gclk));
	jdff dff_B_AVdJ0gQA0_0(.din(n711),.dout(w_dff_B_AVdJ0gQA0_0),.clk(gclk));
	jdff dff_A_PmkHxSYn8_0(.dout(w_G150_3[0]),.din(w_dff_A_PmkHxSYn8_0),.clk(gclk));
	jdff dff_A_1OACN2q06_0(.dout(w_n704_0[0]),.din(w_dff_A_1OACN2q06_0),.clk(gclk));
	jdff dff_A_ntj8JBwS3_0(.dout(w_dff_A_1OACN2q06_0),.din(w_dff_A_ntj8JBwS3_0),.clk(gclk));
	jdff dff_A_hRJp7vWr2_0(.dout(w_n703_1[0]),.din(w_dff_A_hRJp7vWr2_0),.clk(gclk));
	jdff dff_A_DDmYIJHw9_0(.dout(w_dff_A_hRJp7vWr2_0),.din(w_dff_A_DDmYIJHw9_0),.clk(gclk));
	jdff dff_A_ElC4w09o7_0(.dout(w_dff_A_DDmYIJHw9_0),.din(w_dff_A_ElC4w09o7_0),.clk(gclk));
	jdff dff_A_9DxxuXB93_1(.dout(w_n703_0[1]),.din(w_dff_A_9DxxuXB93_1),.clk(gclk));
	jdff dff_A_Ri7ncHCl4_1(.dout(w_dff_A_9DxxuXB93_1),.din(w_dff_A_Ri7ncHCl4_1),.clk(gclk));
	jdff dff_A_13LBD0XT5_1(.dout(w_dff_A_Ri7ncHCl4_1),.din(w_dff_A_13LBD0XT5_1),.clk(gclk));
	jdff dff_A_TiXB0ib65_2(.dout(w_n703_0[2]),.din(w_dff_A_TiXB0ib65_2),.clk(gclk));
	jdff dff_B_qMMpENxz7_0(.din(n702),.dout(w_dff_B_qMMpENxz7_0),.clk(gclk));
	jdff dff_B_ojiNcVtd8_0(.din(w_dff_B_qMMpENxz7_0),.dout(w_dff_B_ojiNcVtd8_0),.clk(gclk));
	jdff dff_B_f6176n3t8_0(.din(w_dff_B_ojiNcVtd8_0),.dout(w_dff_B_f6176n3t8_0),.clk(gclk));
	jdff dff_B_gAgA76Jv1_0(.din(w_dff_B_f6176n3t8_0),.dout(w_dff_B_gAgA76Jv1_0),.clk(gclk));
	jdff dff_B_mCIk2dZs8_0(.din(w_dff_B_gAgA76Jv1_0),.dout(w_dff_B_mCIk2dZs8_0),.clk(gclk));
	jdff dff_A_c60IsobB1_0(.dout(w_n567_3[0]),.din(w_dff_A_c60IsobB1_0),.clk(gclk));
	jdff dff_A_CZjEQc8K0_1(.dout(w_n567_3[1]),.din(w_dff_A_CZjEQc8K0_1),.clk(gclk));
	jdff dff_A_tpiQOmRR1_1(.dout(w_dff_A_CZjEQc8K0_1),.din(w_dff_A_tpiQOmRR1_1),.clk(gclk));
	jdff dff_A_dbW3SnzF1_1(.dout(w_dff_A_tpiQOmRR1_1),.din(w_dff_A_dbW3SnzF1_1),.clk(gclk));
	jdff dff_A_WrqDm6nI6_1(.dout(w_dff_A_dbW3SnzF1_1),.din(w_dff_A_WrqDm6nI6_1),.clk(gclk));
	jdff dff_A_XV4Q8hST0_1(.dout(w_dff_A_WrqDm6nI6_1),.din(w_dff_A_XV4Q8hST0_1),.clk(gclk));
	jdff dff_A_XsYOkWAa1_1(.dout(w_dff_A_XV4Q8hST0_1),.din(w_dff_A_XsYOkWAa1_1),.clk(gclk));
	jdff dff_A_ZRods4mx6_1(.dout(w_dff_A_XsYOkWAa1_1),.din(w_dff_A_ZRods4mx6_1),.clk(gclk));
	jdff dff_A_oNuluRoW1_1(.dout(w_n388_2[1]),.din(w_dff_A_oNuluRoW1_1),.clk(gclk));
	jdff dff_B_2zO82OCK7_1(.din(n384),.dout(w_dff_B_2zO82OCK7_1),.clk(gclk));
	jdff dff_B_tHyOvIpT5_1(.din(w_dff_B_2zO82OCK7_1),.dout(w_dff_B_tHyOvIpT5_1),.clk(gclk));
	jdff dff_A_YvrL0TOD8_1(.dout(w_n383_0[1]),.din(w_dff_A_YvrL0TOD8_1),.clk(gclk));
	jdff dff_A_i6KgicKk7_1(.dout(w_dff_A_YvrL0TOD8_1),.din(w_dff_A_i6KgicKk7_1),.clk(gclk));
	jdff dff_A_EilZvoQR7_1(.dout(w_dff_A_i6KgicKk7_1),.din(w_dff_A_EilZvoQR7_1),.clk(gclk));
	jdff dff_B_bxIqVvov8_1(.din(n374),.dout(w_dff_B_bxIqVvov8_1),.clk(gclk));
	jdff dff_B_eQWyAsEn2_0(.din(n381),.dout(w_dff_B_eQWyAsEn2_0),.clk(gclk));
	jdff dff_B_62Ls3ksn7_1(.din(n376),.dout(w_dff_B_62Ls3ksn7_1),.clk(gclk));
	jdff dff_A_UZUteTL87_0(.dout(w_n378_0[0]),.din(w_dff_A_UZUteTL87_0),.clk(gclk));
	jdff dff_A_AzQ9Rfkm7_0(.dout(w_n370_0[0]),.din(w_dff_A_AzQ9Rfkm7_0),.clk(gclk));
	jdff dff_B_shsYs3545_2(.din(n370),.dout(w_dff_B_shsYs3545_2),.clk(gclk));
	jdff dff_B_Q1nhhtqB4_0(.din(n365),.dout(w_dff_B_Q1nhhtqB4_0),.clk(gclk));
	jdff dff_B_5pQ1P8OX7_1(.din(n358),.dout(w_dff_B_5pQ1P8OX7_1),.clk(gclk));
	jdff dff_A_oCDmwxQd4_1(.dout(w_n357_0[1]),.din(w_dff_A_oCDmwxQd4_1),.clk(gclk));
	jdff dff_A_r1xFQf2C4_1(.dout(w_dff_A_oCDmwxQd4_1),.din(w_dff_A_r1xFQf2C4_1),.clk(gclk));
	jdff dff_A_UjOJvMcG4_0(.dout(w_n356_1[0]),.din(w_dff_A_UjOJvMcG4_0),.clk(gclk));
	jdff dff_A_s56N452h0_1(.dout(w_n356_0[1]),.din(w_dff_A_s56N452h0_1),.clk(gclk));
	jdff dff_A_2v5adAyr4_2(.dout(w_n356_0[2]),.din(w_dff_A_2v5adAyr4_2),.clk(gclk));
	jdff dff_A_o0jD4GnU1_0(.dout(w_n354_1[0]),.din(w_dff_A_o0jD4GnU1_0),.clk(gclk));
	jdff dff_A_5gjoHNAA6_1(.dout(w_n354_0[1]),.din(w_dff_A_5gjoHNAA6_1),.clk(gclk));
	jdff dff_A_knkxMSEg2_2(.dout(w_n354_0[2]),.din(w_dff_A_knkxMSEg2_2),.clk(gclk));
	jdff dff_A_0jrw4gfZ6_1(.dout(w_n1177_0[1]),.din(w_dff_A_0jrw4gfZ6_1),.clk(gclk));
	jdff dff_A_R35VlzGe6_1(.dout(w_dff_A_0jrw4gfZ6_1),.din(w_dff_A_R35VlzGe6_1),.clk(gclk));
	jdff dff_B_jIhpRT4v7_2(.din(n1177),.dout(w_dff_B_jIhpRT4v7_2),.clk(gclk));
	jdff dff_B_6kMIKriX5_2(.din(w_dff_B_jIhpRT4v7_2),.dout(w_dff_B_6kMIKriX5_2),.clk(gclk));
	jdff dff_B_V5R8BYO09_1(.din(n1175),.dout(w_dff_B_V5R8BYO09_1),.clk(gclk));
	jdff dff_B_7nl7DOtC1_1(.din(n942),.dout(w_dff_B_7nl7DOtC1_1),.clk(gclk));
	jdff dff_B_ZN7OJbMQ8_0(.din(n985),.dout(w_dff_B_ZN7OJbMQ8_0),.clk(gclk));
	jdff dff_B_P3RPMK2f3_0(.din(w_dff_B_ZN7OJbMQ8_0),.dout(w_dff_B_P3RPMK2f3_0),.clk(gclk));
	jdff dff_B_DPEIDd9G1_0(.din(w_dff_B_P3RPMK2f3_0),.dout(w_dff_B_DPEIDd9G1_0),.clk(gclk));
	jdff dff_B_UcOqa7wm6_0(.din(w_dff_B_DPEIDd9G1_0),.dout(w_dff_B_UcOqa7wm6_0),.clk(gclk));
	jdff dff_B_dBM934nq7_0(.din(w_dff_B_UcOqa7wm6_0),.dout(w_dff_B_dBM934nq7_0),.clk(gclk));
	jdff dff_B_9KRF2h341_0(.din(n983),.dout(w_dff_B_9KRF2h341_0),.clk(gclk));
	jdff dff_B_x2J2RxHQ3_0(.din(w_dff_B_9KRF2h341_0),.dout(w_dff_B_x2J2RxHQ3_0),.clk(gclk));
	jdff dff_B_uSlMZpg44_1(.din(n949),.dout(w_dff_B_uSlMZpg44_1),.clk(gclk));
	jdff dff_B_gpfmQNdc9_1(.din(w_dff_B_uSlMZpg44_1),.dout(w_dff_B_gpfmQNdc9_1),.clk(gclk));
	jdff dff_B_WEUy2SL86_1(.din(w_dff_B_gpfmQNdc9_1),.dout(w_dff_B_WEUy2SL86_1),.clk(gclk));
	jdff dff_B_mhOjddX57_1(.din(w_dff_B_WEUy2SL86_1),.dout(w_dff_B_mhOjddX57_1),.clk(gclk));
	jdff dff_B_FWJMrzgD2_1(.din(n967),.dout(w_dff_B_FWJMrzgD2_1),.clk(gclk));
	jdff dff_B_SLq0e8Kd6_1(.din(n974),.dout(w_dff_B_SLq0e8Kd6_1),.clk(gclk));
	jdff dff_A_gsN1zYW38_2(.dout(w_G116_2[2]),.din(w_dff_A_gsN1zYW38_2),.clk(gclk));
	jdff dff_B_xNg1sUQ42_1(.din(n965),.dout(w_dff_B_xNg1sUQ42_1),.clk(gclk));
	jdff dff_A_6ms29Wfm8_1(.dout(w_G294_1[1]),.din(w_dff_A_6ms29Wfm8_1),.clk(gclk));
	jdff dff_B_ou8phIP07_1(.din(n952),.dout(w_dff_B_ou8phIP07_1),.clk(gclk));
	jdff dff_B_OwepyVfj8_1(.din(w_dff_B_ou8phIP07_1),.dout(w_dff_B_OwepyVfj8_1),.clk(gclk));
	jdff dff_B_r8bLlVZ74_1(.din(w_dff_B_OwepyVfj8_1),.dout(w_dff_B_r8bLlVZ74_1),.clk(gclk));
	jdff dff_B_ounUMgFs8_1(.din(n955),.dout(w_dff_B_ounUMgFs8_1),.clk(gclk));
	jdff dff_B_cnDPdZq33_1(.din(w_dff_B_ounUMgFs8_1),.dout(w_dff_B_cnDPdZq33_1),.clk(gclk));
	jdff dff_B_hdG0pbbR9_1(.din(n957),.dout(w_dff_B_hdG0pbbR9_1),.clk(gclk));
	jdff dff_A_ImRUhdDb0_0(.dout(w_n959_0[0]),.din(w_dff_A_ImRUhdDb0_0),.clk(gclk));
	jdff dff_A_fJJ6n7k51_0(.dout(w_dff_A_ImRUhdDb0_0),.din(w_dff_A_fJJ6n7k51_0),.clk(gclk));
	jdff dff_A_Q4XdTMH92_0(.dout(w_dff_A_fJJ6n7k51_0),.din(w_dff_A_Q4XdTMH92_0),.clk(gclk));
	jdff dff_A_s0qi0ndp0_2(.dout(w_G143_1[2]),.din(w_dff_A_s0qi0ndp0_2),.clk(gclk));
	jdff dff_A_g49N9GbX7_1(.dout(w_G50_2[1]),.din(w_dff_A_g49N9GbX7_1),.clk(gclk));
	jdff dff_A_sPVdBoWT8_1(.dout(w_dff_A_g49N9GbX7_1),.din(w_dff_A_sPVdBoWT8_1),.clk(gclk));
	jdff dff_A_klVsZxkz3_1(.dout(w_dff_A_sPVdBoWT8_1),.din(w_dff_A_klVsZxkz3_1),.clk(gclk));
	jdff dff_A_IfxbrZjd4_2(.dout(w_G50_2[2]),.din(w_dff_A_IfxbrZjd4_2),.clk(gclk));
	jdff dff_A_iG6SEfJ78_2(.dout(w_dff_A_IfxbrZjd4_2),.din(w_dff_A_iG6SEfJ78_2),.clk(gclk));
	jdff dff_A_uchtVzkm2_2(.dout(w_dff_A_iG6SEfJ78_2),.din(w_dff_A_uchtVzkm2_2),.clk(gclk));
	jdff dff_B_pQFgIYcx9_1(.din(n946),.dout(w_dff_B_pQFgIYcx9_1),.clk(gclk));
	jdff dff_B_Fk6489C09_1(.din(w_dff_B_pQFgIYcx9_1),.dout(w_dff_B_Fk6489C09_1),.clk(gclk));
	jdff dff_B_qayTBsAn8_0(.din(n947),.dout(w_dff_B_qayTBsAn8_0),.clk(gclk));
	jdff dff_A_kTfg7kte6_0(.dout(w_n137_0[0]),.din(w_dff_A_kTfg7kte6_0),.clk(gclk));
	jdff dff_B_3sc9Ecjf8_0(.din(n136),.dout(w_dff_B_3sc9Ecjf8_0),.clk(gclk));
	jdff dff_B_pL18KfnZ3_1(.din(n939),.dout(w_dff_B_pL18KfnZ3_1),.clk(gclk));
	jdff dff_B_IqFXHgBs6_1(.din(n843),.dout(w_dff_B_IqFXHgBs6_1),.clk(gclk));
	jdff dff_B_wxIrUPRk3_1(.din(w_dff_B_IqFXHgBs6_1),.dout(w_dff_B_wxIrUPRk3_1),.clk(gclk));
	jdff dff_B_eBA4zMxn0_1(.din(w_dff_B_wxIrUPRk3_1),.dout(w_dff_B_eBA4zMxn0_1),.clk(gclk));
	jdff dff_B_Fxf59Ko60_1(.din(w_dff_B_eBA4zMxn0_1),.dout(w_dff_B_Fxf59Ko60_1),.clk(gclk));
	jdff dff_B_kPb1VbpD9_1(.din(w_dff_B_Fxf59Ko60_1),.dout(w_dff_B_kPb1VbpD9_1),.clk(gclk));
	jdff dff_B_YMfXw1AN3_1(.din(w_dff_B_kPb1VbpD9_1),.dout(w_dff_B_YMfXw1AN3_1),.clk(gclk));
	jdff dff_B_wmhtPQGZ2_1(.din(w_dff_B_YMfXw1AN3_1),.dout(w_dff_B_wmhtPQGZ2_1),.clk(gclk));
	jdff dff_B_ApcI78CP0_1(.din(n856),.dout(w_dff_B_ApcI78CP0_1),.clk(gclk));
	jdff dff_B_a7sBk9jl0_1(.din(w_dff_B_ApcI78CP0_1),.dout(w_dff_B_a7sBk9jl0_1),.clk(gclk));
	jdff dff_B_ySXOopji0_0(.din(n866),.dout(w_dff_B_ySXOopji0_0),.clk(gclk));
	jdff dff_A_uuXYZh7f9_0(.dout(w_n863_0[0]),.din(w_dff_A_uuXYZh7f9_0),.clk(gclk));
	jdff dff_A_aeBcOHkp3_0(.dout(w_dff_A_uuXYZh7f9_0),.din(w_dff_A_aeBcOHkp3_0),.clk(gclk));
	jdff dff_A_nI7djk5b5_0(.dout(w_dff_A_aeBcOHkp3_0),.din(w_dff_A_nI7djk5b5_0),.clk(gclk));
	jdff dff_A_Gt3uamDq6_2(.dout(w_n863_0[2]),.din(w_dff_A_Gt3uamDq6_2),.clk(gclk));
	jdff dff_B_orJoUx8x2_1(.din(n847),.dout(w_dff_B_orJoUx8x2_1),.clk(gclk));
	jdff dff_B_b8Fn2muT3_1(.din(n848),.dout(w_dff_B_b8Fn2muT3_1),.clk(gclk));
	jdff dff_B_hiwWDqOG1_1(.din(w_dff_B_b8Fn2muT3_1),.dout(w_dff_B_hiwWDqOG1_1),.clk(gclk));
	jdff dff_B_In3jeXyT8_1(.din(w_dff_B_hiwWDqOG1_1),.dout(w_dff_B_In3jeXyT8_1),.clk(gclk));
	jdff dff_B_VjYy4XQB0_1(.din(w_dff_B_In3jeXyT8_1),.dout(w_dff_B_VjYy4XQB0_1),.clk(gclk));
	jdff dff_B_7fAGyRMk1_0(.din(n851),.dout(w_dff_B_7fAGyRMk1_0),.clk(gclk));
	jdff dff_A_3aHxw2DG4_1(.dout(w_n569_0[1]),.din(w_dff_A_3aHxw2DG4_1),.clk(gclk));
	jdff dff_A_7Mu1Dhco8_1(.dout(w_dff_A_3aHxw2DG4_1),.din(w_dff_A_7Mu1Dhco8_1),.clk(gclk));
	jdff dff_A_lFUaObDu7_0(.dout(w_n348_0[0]),.din(w_dff_A_lFUaObDu7_0),.clk(gclk));
	jdff dff_A_DdNK124j6_0(.dout(w_n333_0[0]),.din(w_dff_A_DdNK124j6_0),.clk(gclk));
	jdff dff_A_6VGMMbyj4_0(.dout(w_dff_A_DdNK124j6_0),.din(w_dff_A_6VGMMbyj4_0),.clk(gclk));
	jdff dff_B_cWK7IIex0_0(.din(n846),.dout(w_dff_B_cWK7IIex0_0),.clk(gclk));
	jdff dff_B_FDvsbCPd3_0(.din(w_dff_B_cWK7IIex0_0),.dout(w_dff_B_FDvsbCPd3_0),.clk(gclk));
	jdff dff_A_P5A958rJ9_1(.dout(w_n845_0[1]),.din(w_dff_A_P5A958rJ9_1),.clk(gclk));
	jdff dff_A_0QAog1zj5_1(.dout(w_dff_A_P5A958rJ9_1),.din(w_dff_A_0QAog1zj5_1),.clk(gclk));
	jdff dff_A_PJ6xGTsY9_1(.dout(w_dff_A_0QAog1zj5_1),.din(w_dff_A_PJ6xGTsY9_1),.clk(gclk));
	jdff dff_A_gGJ6Bts46_1(.dout(w_dff_A_PJ6xGTsY9_1),.din(w_dff_A_gGJ6Bts46_1),.clk(gclk));
	jdff dff_B_4U45jzSB5_0(.din(n844),.dout(w_dff_B_4U45jzSB5_0),.clk(gclk));
	jdff dff_B_PJ66t5yM2_0(.din(w_dff_B_4U45jzSB5_0),.dout(w_dff_B_PJ66t5yM2_0),.clk(gclk));
	jdff dff_B_Uf0XxWAg0_0(.din(w_dff_B_PJ66t5yM2_0),.dout(w_dff_B_Uf0XxWAg0_0),.clk(gclk));
	jdff dff_A_fGNBHnwj8_1(.dout(w_n579_1[1]),.din(w_dff_A_fGNBHnwj8_1),.clk(gclk));
	jdff dff_A_nnTQgwfk1_1(.dout(w_dff_A_fGNBHnwj8_1),.din(w_dff_A_nnTQgwfk1_1),.clk(gclk));
	jdff dff_B_XjXOnsmf3_0(.din(n841),.dout(w_dff_B_XjXOnsmf3_0),.clk(gclk));
	jdff dff_B_6esktB4V4_1(.din(n806),.dout(w_dff_B_6esktB4V4_1),.clk(gclk));
	jdff dff_B_dDHsSDnA9_1(.din(w_dff_B_6esktB4V4_1),.dout(w_dff_B_dDHsSDnA9_1),.clk(gclk));
	jdff dff_B_zT8eHC0d9_1(.din(w_dff_B_dDHsSDnA9_1),.dout(w_dff_B_zT8eHC0d9_1),.clk(gclk));
	jdff dff_B_hjXK9s2E9_1(.din(n825),.dout(w_dff_B_hjXK9s2E9_1),.clk(gclk));
	jdff dff_B_1bIJ8zSE5_1(.din(w_dff_B_hjXK9s2E9_1),.dout(w_dff_B_1bIJ8zSE5_1),.clk(gclk));
	jdff dff_B_ufJdp9e54_1(.din(n828),.dout(w_dff_B_ufJdp9e54_1),.clk(gclk));
	jdff dff_B_RQ0tSwua1_1(.din(w_dff_B_ufJdp9e54_1),.dout(w_dff_B_RQ0tSwua1_1),.clk(gclk));
	jdff dff_B_VQ8gnLiz2_0(.din(n834),.dout(w_dff_B_VQ8gnLiz2_0),.clk(gclk));
	jdff dff_A_t8N1d5Pb7_0(.dout(w_n833_0[0]),.din(w_dff_A_t8N1d5Pb7_0),.clk(gclk));
	jdff dff_B_YSJ6bEhz9_1(.din(n829),.dout(w_dff_B_YSJ6bEhz9_1),.clk(gclk));
	jdff dff_A_bKy6J2rE7_0(.dout(w_G58_3[0]),.din(w_dff_A_bKy6J2rE7_0),.clk(gclk));
	jdff dff_A_gM5IJcWt1_0(.dout(w_dff_A_bKy6J2rE7_0),.din(w_dff_A_gM5IJcWt1_0),.clk(gclk));
	jdff dff_A_xkJlU7Il1_0(.dout(w_dff_A_gM5IJcWt1_0),.din(w_dff_A_xkJlU7Il1_0),.clk(gclk));
	jdff dff_A_2QxankVB8_2(.dout(w_G58_3[2]),.din(w_dff_A_2QxankVB8_2),.clk(gclk));
	jdff dff_A_9qQuyDoI6_2(.dout(w_dff_A_2QxankVB8_2),.din(w_dff_A_9qQuyDoI6_2),.clk(gclk));
	jdff dff_A_quOWGrrx4_2(.dout(w_dff_A_9qQuyDoI6_2),.din(w_dff_A_quOWGrrx4_2),.clk(gclk));
	jdff dff_A_0y1D0MhM1_2(.dout(w_dff_A_quOWGrrx4_2),.din(w_dff_A_0y1D0MhM1_2),.clk(gclk));
	jdff dff_B_CF3vVTP54_3(.din(G143),.dout(w_dff_B_CF3vVTP54_3),.clk(gclk));
	jdff dff_B_57chmTx82_3(.din(w_dff_B_CF3vVTP54_3),.dout(w_dff_B_57chmTx82_3),.clk(gclk));
	jdff dff_B_1WN0ZySe4_3(.din(w_dff_B_57chmTx82_3),.dout(w_dff_B_1WN0ZySe4_3),.clk(gclk));
	jdff dff_B_BdpCwJC28_1(.din(n823),.dout(w_dff_B_BdpCwJC28_1),.clk(gclk));
	jdff dff_A_zT8TQK0W9_1(.dout(w_G137_1[1]),.din(w_dff_A_zT8TQK0W9_1),.clk(gclk));
	jdff dff_B_ThHvDAIp5_3(.din(G137),.dout(w_dff_B_ThHvDAIp5_3),.clk(gclk));
	jdff dff_B_ArM46iT91_3(.din(w_dff_B_ThHvDAIp5_3),.dout(w_dff_B_ArM46iT91_3),.clk(gclk));
	jdff dff_B_szlZOZXh5_3(.din(w_dff_B_ArM46iT91_3),.dout(w_dff_B_szlZOZXh5_3),.clk(gclk));
	jdff dff_B_MpMlUWve7_1(.din(n809),.dout(w_dff_B_MpMlUWve7_1),.clk(gclk));
	jdff dff_B_rU4T2go71_1(.din(w_dff_B_MpMlUWve7_1),.dout(w_dff_B_rU4T2go71_1),.clk(gclk));
	jdff dff_B_tmSYz4yx9_1(.din(w_dff_B_rU4T2go71_1),.dout(w_dff_B_tmSYz4yx9_1),.clk(gclk));
	jdff dff_B_5iAuwOLi4_1(.din(n812),.dout(w_dff_B_5iAuwOLi4_1),.clk(gclk));
	jdff dff_B_1IAQThCU0_1(.din(w_dff_B_5iAuwOLi4_1),.dout(w_dff_B_1IAQThCU0_1),.clk(gclk));
	jdff dff_A_HEyFGdAl1_1(.dout(w_G107_2[1]),.din(w_dff_A_HEyFGdAl1_1),.clk(gclk));
	jdff dff_B_T5V9d2Bh4_1(.din(n813),.dout(w_dff_B_T5V9d2Bh4_1),.clk(gclk));
	jdff dff_A_N8zkPk2V5_0(.dout(w_n680_3[0]),.din(w_dff_A_N8zkPk2V5_0),.clk(gclk));
	jdff dff_A_v8vdYEFd9_0(.dout(w_dff_A_N8zkPk2V5_0),.din(w_dff_A_v8vdYEFd9_0),.clk(gclk));
	jdff dff_A_4UGmj34i8_0(.dout(w_dff_A_v8vdYEFd9_0),.din(w_dff_A_4UGmj34i8_0),.clk(gclk));
	jdff dff_A_f7y5WgPL4_0(.dout(w_dff_A_4UGmj34i8_0),.din(w_dff_A_f7y5WgPL4_0),.clk(gclk));
	jdff dff_A_nXgID33p2_0(.dout(w_dff_A_f7y5WgPL4_0),.din(w_dff_A_nXgID33p2_0),.clk(gclk));
	jdff dff_A_pzRQG86f7_0(.dout(w_dff_A_nXgID33p2_0),.din(w_dff_A_pzRQG86f7_0),.clk(gclk));
	jdff dff_A_hW8AAyM75_0(.dout(w_dff_A_pzRQG86f7_0),.din(w_dff_A_hW8AAyM75_0),.clk(gclk));
	jdff dff_A_k6m6EGB75_2(.dout(w_n680_3[2]),.din(w_dff_A_k6m6EGB75_2),.clk(gclk));
	jdff dff_A_0EEZjhwS3_2(.dout(w_dff_A_k6m6EGB75_2),.din(w_dff_A_0EEZjhwS3_2),.clk(gclk));
	jdff dff_A_odTVlco66_2(.dout(w_dff_A_0EEZjhwS3_2),.din(w_dff_A_odTVlco66_2),.clk(gclk));
	jdff dff_A_kQVuwrPh6_2(.dout(w_dff_A_odTVlco66_2),.din(w_dff_A_kQVuwrPh6_2),.clk(gclk));
	jdff dff_A_SuGQnfHG3_2(.dout(w_dff_A_kQVuwrPh6_2),.din(w_dff_A_SuGQnfHG3_2),.clk(gclk));
	jdff dff_A_0etCkqs48_2(.dout(w_dff_A_SuGQnfHG3_2),.din(w_dff_A_0etCkqs48_2),.clk(gclk));
	jdff dff_B_fW4BpqX15_1(.din(n801),.dout(w_dff_B_fW4BpqX15_1),.clk(gclk));
	jdff dff_B_2ANOq5n72_1(.din(w_dff_B_fW4BpqX15_1),.dout(w_dff_B_2ANOq5n72_1),.clk(gclk));
	jdff dff_B_Fxsrb80G4_0(.din(n803),.dout(w_dff_B_Fxsrb80G4_0),.clk(gclk));
	jdff dff_A_S3wOPQv49_0(.dout(w_n126_0[0]),.din(w_dff_A_S3wOPQv49_0),.clk(gclk));
	jdff dff_B_Xy3Tfcgg6_0(.din(n125),.dout(w_dff_B_Xy3Tfcgg6_0),.clk(gclk));
	jdff dff_A_EQTcbEZH4_1(.dout(w_n614_4[1]),.din(w_dff_A_EQTcbEZH4_1),.clk(gclk));
	jdff dff_A_8vmb2NwO7_1(.dout(w_dff_A_EQTcbEZH4_1),.din(w_dff_A_8vmb2NwO7_1),.clk(gclk));
	jdff dff_A_e0QIJYxy9_1(.dout(w_dff_A_8vmb2NwO7_1),.din(w_dff_A_e0QIJYxy9_1),.clk(gclk));
	jdff dff_A_cetJO7la0_1(.dout(w_dff_A_e0QIJYxy9_1),.din(w_dff_A_cetJO7la0_1),.clk(gclk));
	jdff dff_A_07Ru6seW5_1(.dout(w_dff_A_cetJO7la0_1),.din(w_dff_A_07Ru6seW5_1),.clk(gclk));
	jdff dff_A_zrrb1dWY3_1(.dout(w_dff_A_07Ru6seW5_1),.din(w_dff_A_zrrb1dWY3_1),.clk(gclk));
	jdff dff_A_jzGcGysS2_1(.dout(w_dff_A_zrrb1dWY3_1),.din(w_dff_A_jzGcGysS2_1),.clk(gclk));
	jdff dff_A_NMgCCs5d2_1(.dout(w_dff_A_jzGcGysS2_1),.din(w_dff_A_NMgCCs5d2_1),.clk(gclk));
	jdff dff_A_YNwvWcum7_1(.dout(w_dff_A_NMgCCs5d2_1),.din(w_dff_A_YNwvWcum7_1),.clk(gclk));
	jdff dff_A_JsZ5AxpJ8_1(.dout(w_dff_A_YNwvWcum7_1),.din(w_dff_A_JsZ5AxpJ8_1),.clk(gclk));
	jdff dff_A_h4H1DHsB8_1(.dout(w_dff_A_JsZ5AxpJ8_1),.din(w_dff_A_h4H1DHsB8_1),.clk(gclk));
	jdff dff_A_HfBoGHCo1_1(.dout(w_dff_A_h4H1DHsB8_1),.din(w_dff_A_HfBoGHCo1_1),.clk(gclk));
	jdff dff_A_edMqENaC1_2(.dout(w_n614_4[2]),.din(w_dff_A_edMqENaC1_2),.clk(gclk));
	jdff dff_A_dPPxc8oq7_2(.dout(w_dff_A_edMqENaC1_2),.din(w_dff_A_dPPxc8oq7_2),.clk(gclk));
	jdff dff_A_FYxxkD401_2(.dout(w_dff_A_dPPxc8oq7_2),.din(w_dff_A_FYxxkD401_2),.clk(gclk));
	jdff dff_A_oZO6c03a0_2(.dout(w_dff_A_FYxxkD401_2),.din(w_dff_A_oZO6c03a0_2),.clk(gclk));
	jdff dff_A_7ljpYLmB9_0(.dout(w_n798_0[0]),.din(w_dff_A_7ljpYLmB9_0),.clk(gclk));
	jdff dff_A_dXgb7lB73_0(.dout(w_dff_A_7ljpYLmB9_0),.din(w_dff_A_dXgb7lB73_0),.clk(gclk));
	jdff dff_A_3AJGYNJi7_0(.dout(w_dff_A_dXgb7lB73_0),.din(w_dff_A_3AJGYNJi7_0),.clk(gclk));
	jdff dff_A_8e3u4AU77_0(.dout(w_dff_A_3AJGYNJi7_0),.din(w_dff_A_8e3u4AU77_0),.clk(gclk));
	jdff dff_A_VCu3sJlL1_0(.dout(w_dff_A_8e3u4AU77_0),.din(w_dff_A_VCu3sJlL1_0),.clk(gclk));
	jdff dff_B_nKDuQ6uv3_0(.din(n797),.dout(w_dff_B_nKDuQ6uv3_0),.clk(gclk));
	jdff dff_B_8GrNoiK39_0(.din(w_dff_B_nKDuQ6uv3_0),.dout(w_dff_B_8GrNoiK39_0),.clk(gclk));
	jdff dff_A_CAZW4RVx2_2(.dout(w_n567_2[2]),.din(w_dff_A_CAZW4RVx2_2),.clk(gclk));
	jdff dff_A_qAWZsXJr4_2(.dout(w_dff_A_CAZW4RVx2_2),.din(w_dff_A_qAWZsXJr4_2),.clk(gclk));
	jdff dff_A_eTQddzzA9_2(.dout(w_dff_A_qAWZsXJr4_2),.din(w_dff_A_eTQddzzA9_2),.clk(gclk));
	jdff dff_A_PVE1CDEL4_2(.dout(w_dff_A_eTQddzzA9_2),.din(w_dff_A_PVE1CDEL4_2),.clk(gclk));
	jdff dff_A_F23E7Z5V8_2(.dout(w_dff_A_PVE1CDEL4_2),.din(w_dff_A_F23E7Z5V8_2),.clk(gclk));
	jdff dff_A_rPtILABT7_2(.dout(w_dff_A_F23E7Z5V8_2),.din(w_dff_A_rPtILABT7_2),.clk(gclk));
	jdff dff_A_pgcBG5UC7_2(.dout(w_dff_A_rPtILABT7_2),.din(w_dff_A_pgcBG5UC7_2),.clk(gclk));
	jdff dff_A_OghlpeEH0_2(.dout(w_dff_A_pgcBG5UC7_2),.din(w_dff_A_OghlpeEH0_2),.clk(gclk));
	jdff dff_A_BcrQTTm06_2(.dout(w_dff_A_OghlpeEH0_2),.din(w_dff_A_BcrQTTm06_2),.clk(gclk));
	jdff dff_B_Y8wnFUcd0_0(.din(n936),.dout(w_dff_B_Y8wnFUcd0_0),.clk(gclk));
	jdff dff_B_1ymcwVnc5_0(.din(w_dff_B_Y8wnFUcd0_0),.dout(w_dff_B_1ymcwVnc5_0),.clk(gclk));
	jdff dff_B_bnEJzStn0_0(.din(w_dff_B_1ymcwVnc5_0),.dout(w_dff_B_bnEJzStn0_0),.clk(gclk));
	jdff dff_B_01GKseaG2_0(.din(w_dff_B_bnEJzStn0_0),.dout(w_dff_B_01GKseaG2_0),.clk(gclk));
	jdff dff_B_kBTgxbTc6_0(.din(w_dff_B_01GKseaG2_0),.dout(w_dff_B_kBTgxbTc6_0),.clk(gclk));
	jdff dff_B_ThDjJH2c2_0(.din(n932),.dout(w_dff_B_ThDjJH2c2_0),.clk(gclk));
	jdff dff_B_lRcnW8Hx2_0(.din(w_dff_B_ThDjJH2c2_0),.dout(w_dff_B_lRcnW8Hx2_0),.clk(gclk));
	jdff dff_B_ZuP8Rk7Z9_1(.din(n917),.dout(w_dff_B_ZuP8Rk7Z9_1),.clk(gclk));
	jdff dff_B_N8VLJqyG2_1(.din(w_dff_B_ZuP8Rk7Z9_1),.dout(w_dff_B_N8VLJqyG2_1),.clk(gclk));
	jdff dff_B_VkhJlcVA1_1(.din(w_dff_B_N8VLJqyG2_1),.dout(w_dff_B_VkhJlcVA1_1),.clk(gclk));
	jdff dff_B_9sPCvJLp1_0(.din(n929),.dout(w_dff_B_9sPCvJLp1_0),.clk(gclk));
	jdff dff_B_qpxD3fEa0_0(.din(w_dff_B_9sPCvJLp1_0),.dout(w_dff_B_qpxD3fEa0_0),.clk(gclk));
	jdff dff_B_3E0Ul3YV3_0(.din(n927),.dout(w_dff_B_3E0Ul3YV3_0),.clk(gclk));
	jdff dff_A_V6O6VTJa3_1(.dout(w_n73_1[1]),.din(w_dff_A_V6O6VTJa3_1),.clk(gclk));
	jdff dff_A_Ye7xy3Ka0_1(.dout(w_dff_A_V6O6VTJa3_1),.din(w_dff_A_Ye7xy3Ka0_1),.clk(gclk));
	jdff dff_A_ujABWE8i1_2(.dout(w_n73_1[2]),.din(w_dff_A_ujABWE8i1_2),.clk(gclk));
	jdff dff_A_G8EXsN8I4_2(.dout(w_dff_A_ujABWE8i1_2),.din(w_dff_A_G8EXsN8I4_2),.clk(gclk));
	jdff dff_A_AqxmzgaN0_2(.dout(w_dff_A_G8EXsN8I4_2),.din(w_dff_A_AqxmzgaN0_2),.clk(gclk));
	jdff dff_A_hCY0c5F84_2(.dout(w_dff_A_AqxmzgaN0_2),.din(w_dff_A_hCY0c5F84_2),.clk(gclk));
	jdff dff_A_4csDuuaN6_2(.dout(w_n73_0[2]),.din(w_dff_A_4csDuuaN6_2),.clk(gclk));
	jdff dff_A_R8bxaq8C7_2(.dout(w_dff_A_4csDuuaN6_2),.din(w_dff_A_R8bxaq8C7_2),.clk(gclk));
	jdff dff_A_kBcCz6HL9_2(.dout(w_dff_A_R8bxaq8C7_2),.din(w_dff_A_kBcCz6HL9_2),.clk(gclk));
	jdff dff_A_tF8vX1f22_2(.dout(w_dff_A_kBcCz6HL9_2),.din(w_dff_A_tF8vX1f22_2),.clk(gclk));
	jdff dff_B_Ln9ZbyCK9_0(.din(n922),.dout(w_dff_B_Ln9ZbyCK9_0),.clk(gclk));
	jdff dff_B_f9OO8QL00_0(.din(n921),.dout(w_dff_B_f9OO8QL00_0),.clk(gclk));
	jdff dff_A_sGUw0pmT6_1(.dout(w_n130_0[1]),.din(w_dff_A_sGUw0pmT6_1),.clk(gclk));
	jdff dff_B_dVKmhsVS6_0(.din(n129),.dout(w_dff_B_dVKmhsVS6_0),.clk(gclk));
	jdff dff_A_6b1FezRd7_0(.dout(w_G232_1[0]),.din(w_dff_A_6b1FezRd7_0),.clk(gclk));
	jdff dff_A_Gus10aQ47_0(.dout(w_dff_A_6b1FezRd7_0),.din(w_dff_A_Gus10aQ47_0),.clk(gclk));
	jdff dff_A_8DYJNc5I8_1(.dout(w_G232_0[1]),.din(w_dff_A_8DYJNc5I8_1),.clk(gclk));
	jdff dff_A_aFrgECxh2_1(.dout(w_dff_A_8DYJNc5I8_1),.din(w_dff_A_aFrgECxh2_1),.clk(gclk));
	jdff dff_A_sM4oKHqN0_1(.dout(w_dff_A_aFrgECxh2_1),.din(w_dff_A_sM4oKHqN0_1),.clk(gclk));
	jdff dff_A_eoF0XVMH7_2(.dout(w_G232_0[2]),.din(w_dff_A_eoF0XVMH7_2),.clk(gclk));
	jdff dff_A_73qoDkLk9_2(.dout(w_dff_A_eoF0XVMH7_2),.din(w_dff_A_73qoDkLk9_2),.clk(gclk));
	jdff dff_A_OnZNoG9q7_0(.dout(w_G226_1[0]),.din(w_dff_A_OnZNoG9q7_0),.clk(gclk));
	jdff dff_A_SpIpFv3q9_0(.dout(w_dff_A_OnZNoG9q7_0),.din(w_dff_A_SpIpFv3q9_0),.clk(gclk));
	jdff dff_A_72t6ETG10_1(.dout(w_G226_0[1]),.din(w_dff_A_72t6ETG10_1),.clk(gclk));
	jdff dff_A_X1tZQeR31_1(.dout(w_dff_A_72t6ETG10_1),.din(w_dff_A_X1tZQeR31_1),.clk(gclk));
	jdff dff_A_Og5MRb3q7_2(.dout(w_G226_0[2]),.din(w_dff_A_Og5MRb3q7_2),.clk(gclk));
	jdff dff_A_L5KZjV4q2_2(.dout(w_dff_A_Og5MRb3q7_2),.din(w_dff_A_L5KZjV4q2_2),.clk(gclk));
	jdff dff_A_sEVsS5Ua6_2(.dout(w_dff_A_L5KZjV4q2_2),.din(w_dff_A_sEVsS5Ua6_2),.clk(gclk));
	jdff dff_A_pGqw67Fc1_1(.dout(w_n802_0[1]),.din(w_dff_A_pGqw67Fc1_1),.clk(gclk));
	jdff dff_A_sAcMoqNB6_1(.dout(w_dff_A_pGqw67Fc1_1),.din(w_dff_A_sAcMoqNB6_1),.clk(gclk));
	jdff dff_A_FH96tEjZ0_1(.dout(w_dff_A_sAcMoqNB6_1),.din(w_dff_A_FH96tEjZ0_1),.clk(gclk));
	jdff dff_A_VMOJjKVJ3_1(.dout(w_dff_A_FH96tEjZ0_1),.din(w_dff_A_VMOJjKVJ3_1),.clk(gclk));
	jdff dff_B_CdPONrv61_0(.din(n913),.dout(w_dff_B_CdPONrv61_0),.clk(gclk));
	jdff dff_B_Lc4vOZKj4_0(.din(w_dff_B_CdPONrv61_0),.dout(w_dff_B_Lc4vOZKj4_0),.clk(gclk));
	jdff dff_B_BxPg4YKO0_1(.din(n898),.dout(w_dff_B_BxPg4YKO0_1),.clk(gclk));
	jdff dff_B_7ENqnbhr4_1(.din(w_dff_B_BxPg4YKO0_1),.dout(w_dff_B_7ENqnbhr4_1),.clk(gclk));
	jdff dff_B_wjSu0zAU3_1(.din(w_dff_B_7ENqnbhr4_1),.dout(w_dff_B_wjSu0zAU3_1),.clk(gclk));
	jdff dff_B_hVb0CsHc0_1(.din(w_dff_B_wjSu0zAU3_1),.dout(w_dff_B_hVb0CsHc0_1),.clk(gclk));
	jdff dff_B_5iePj3C97_0(.din(n909),.dout(w_dff_B_5iePj3C97_0),.clk(gclk));
	jdff dff_A_ymCLt7bK8_1(.dout(w_n153_3[1]),.din(w_dff_A_ymCLt7bK8_1),.clk(gclk));
	jdff dff_A_gqd75nBO0_1(.dout(w_dff_A_ymCLt7bK8_1),.din(w_dff_A_gqd75nBO0_1),.clk(gclk));
	jdff dff_A_maskZQOy6_1(.dout(w_dff_A_gqd75nBO0_1),.din(w_dff_A_maskZQOy6_1),.clk(gclk));
	jdff dff_A_qCiB9QtQ7_1(.dout(w_dff_A_maskZQOy6_1),.din(w_dff_A_qCiB9QtQ7_1),.clk(gclk));
	jdff dff_A_EjlM9Hnm1_1(.dout(w_dff_A_qCiB9QtQ7_1),.din(w_dff_A_EjlM9Hnm1_1),.clk(gclk));
	jdff dff_A_M6yMn2DP4_2(.dout(w_n153_3[2]),.din(w_dff_A_M6yMn2DP4_2),.clk(gclk));
	jdff dff_A_V4Oy8Dsb1_2(.dout(w_dff_A_M6yMn2DP4_2),.din(w_dff_A_V4Oy8Dsb1_2),.clk(gclk));
	jdff dff_B_VPxtV2Dm3_1(.din(n902),.dout(w_dff_B_VPxtV2Dm3_1),.clk(gclk));
	jdff dff_B_RSXJqNCL9_1(.din(n899),.dout(w_dff_B_RSXJqNCL9_1),.clk(gclk));
	jdff dff_A_VexwC1p14_1(.dout(w_G283_2[1]),.din(w_dff_A_VexwC1p14_1),.clk(gclk));
	jdff dff_B_9z8F1Thl9_1(.din(n883),.dout(w_dff_B_9z8F1Thl9_1),.clk(gclk));
	jdff dff_B_DDUoAJAO2_1(.din(n888),.dout(w_dff_B_DDUoAJAO2_1),.clk(gclk));
	jdff dff_B_ml9GC6oQ8_0(.din(n892),.dout(w_dff_B_ml9GC6oQ8_0),.clk(gclk));
	jdff dff_B_7bU8Sqr96_0(.din(w_dff_B_ml9GC6oQ8_0),.dout(w_dff_B_7bU8Sqr96_0),.clk(gclk));
	jdff dff_B_HALy3Khn7_1(.din(n889),.dout(w_dff_B_HALy3Khn7_1),.clk(gclk));
	jdff dff_A_67XSxAJS6_1(.dout(w_G150_2[1]),.din(w_dff_A_67XSxAJS6_1),.clk(gclk));
	jdff dff_A_YVUJFrSK3_0(.dout(w_G150_0[0]),.din(w_dff_A_YVUJFrSK3_0),.clk(gclk));
	jdff dff_A_cZPzdJwJ2_1(.dout(w_G150_0[1]),.din(w_dff_A_cZPzdJwJ2_1),.clk(gclk));
	jdff dff_B_yVxTtLLJ4_3(.din(G150),.dout(w_dff_B_yVxTtLLJ4_3),.clk(gclk));
	jdff dff_B_fxZ7pw9z2_3(.din(w_dff_B_yVxTtLLJ4_3),.dout(w_dff_B_fxZ7pw9z2_3),.clk(gclk));
	jdff dff_A_u86Ibo975_0(.dout(w_G50_3[0]),.din(w_dff_A_u86Ibo975_0),.clk(gclk));
	jdff dff_A_6bLnyUtW9_0(.dout(w_dff_A_u86Ibo975_0),.din(w_dff_A_6bLnyUtW9_0),.clk(gclk));
	jdff dff_A_AU5f9WES5_0(.dout(w_dff_A_6bLnyUtW9_0),.din(w_dff_A_AU5f9WES5_0),.clk(gclk));
	jdff dff_A_OeXoWeOW9_1(.dout(w_G50_3[1]),.din(w_dff_A_OeXoWeOW9_1),.clk(gclk));
	jdff dff_A_TttI0QSF7_1(.dout(w_dff_A_OeXoWeOW9_1),.din(w_dff_A_TttI0QSF7_1),.clk(gclk));
	jdff dff_A_tzRFdULo5_1(.dout(w_dff_A_TttI0QSF7_1),.din(w_dff_A_tzRFdULo5_1),.clk(gclk));
	jdff dff_A_BcUIqjLa9_1(.dout(w_n887_0[1]),.din(w_dff_A_BcUIqjLa9_1),.clk(gclk));
	jdff dff_A_GJ0JER405_0(.dout(w_G77_2[0]),.din(w_dff_A_GJ0JER405_0),.clk(gclk));
	jdff dff_A_8PYxwOD49_1(.dout(w_G77_2[1]),.din(w_dff_A_8PYxwOD49_1),.clk(gclk));
	jdff dff_A_z1JNQAMu2_1(.dout(w_G87_1[1]),.din(w_dff_A_z1JNQAMu2_1),.clk(gclk));
	jdff dff_A_QAlOaucd4_2(.dout(w_G87_1[2]),.din(w_dff_A_QAlOaucd4_2),.clk(gclk));
	jdff dff_B_S1TWYexl9_1(.din(n878),.dout(w_dff_B_S1TWYexl9_1),.clk(gclk));
	jdff dff_B_qO6l6Hji1_1(.din(w_dff_B_S1TWYexl9_1),.dout(w_dff_B_qO6l6Hji1_1),.clk(gclk));
	jdff dff_A_TE9mGCgW0_1(.dout(w_G68_2[1]),.din(w_dff_A_TE9mGCgW0_1),.clk(gclk));
	jdff dff_A_4lNsKam10_1(.dout(w_dff_A_TE9mGCgW0_1),.din(w_dff_A_4lNsKam10_1),.clk(gclk));
	jdff dff_A_NG3RrSe38_1(.dout(w_dff_A_4lNsKam10_1),.din(w_dff_A_NG3RrSe38_1),.clk(gclk));
	jdff dff_A_jJQgm6LR5_2(.dout(w_G68_2[2]),.din(w_dff_A_jJQgm6LR5_2),.clk(gclk));
	jdff dff_A_XElAkDnA6_2(.dout(w_dff_A_jJQgm6LR5_2),.din(w_dff_A_XElAkDnA6_2),.clk(gclk));
	jdff dff_A_sKmGXIaU0_2(.dout(w_dff_A_XElAkDnA6_2),.din(w_dff_A_sKmGXIaU0_2),.clk(gclk));
	jdff dff_A_9LWVJ9J94_2(.dout(w_dff_A_sKmGXIaU0_2),.din(w_dff_A_9LWVJ9J94_2),.clk(gclk));
	jdff dff_A_RMo9H0qy0_1(.dout(w_n817_0[1]),.din(w_dff_A_RMo9H0qy0_1),.clk(gclk));
	jdff dff_A_VOJ3Gx0C6_1(.dout(w_G97_2[1]),.din(w_dff_A_VOJ3Gx0C6_1),.clk(gclk));
	jdff dff_A_XF5SPZMu9_1(.dout(w_G33_5[1]),.din(w_dff_A_XF5SPZMu9_1),.clk(gclk));
	jdff dff_A_w4f6Aana9_1(.dout(w_dff_A_XF5SPZMu9_1),.din(w_dff_A_w4f6Aana9_1),.clk(gclk));
	jdff dff_A_CzPuB0WY5_1(.dout(w_dff_A_w4f6Aana9_1),.din(w_dff_A_CzPuB0WY5_1),.clk(gclk));
	jdff dff_A_SmDPUhHV2_0(.dout(w_G58_2[0]),.din(w_dff_A_SmDPUhHV2_0),.clk(gclk));
	jdff dff_A_F1LSShtC4_0(.dout(w_dff_A_SmDPUhHV2_0),.din(w_dff_A_F1LSShtC4_0),.clk(gclk));
	jdff dff_A_vXOkiJ2b4_2(.dout(w_G58_2[2]),.din(w_dff_A_vXOkiJ2b4_2),.clk(gclk));
	jdff dff_A_E72xmQJQ7_2(.dout(w_dff_A_vXOkiJ2b4_2),.din(w_dff_A_E72xmQJQ7_2),.clk(gclk));
	jdff dff_A_7L8arQuy9_0(.dout(w_n680_2[0]),.din(w_dff_A_7L8arQuy9_0),.clk(gclk));
	jdff dff_A_zQ0aq7wq3_0(.dout(w_dff_A_7L8arQuy9_0),.din(w_dff_A_zQ0aq7wq3_0),.clk(gclk));
	jdff dff_A_X4weM8Cq6_2(.dout(w_n680_2[2]),.din(w_dff_A_X4weM8Cq6_2),.clk(gclk));
	jdff dff_A_IQpk0kVG8_2(.dout(w_dff_A_X4weM8Cq6_2),.din(w_dff_A_IQpk0kVG8_2),.clk(gclk));
	jdff dff_A_7lY5Beui3_2(.dout(w_dff_A_IQpk0kVG8_2),.din(w_dff_A_7lY5Beui3_2),.clk(gclk));
	jdff dff_A_4zFnBeeD1_1(.dout(w_n614_3[1]),.din(w_dff_A_4zFnBeeD1_1),.clk(gclk));
	jdff dff_A_XsDSl20W7_1(.dout(w_dff_A_4zFnBeeD1_1),.din(w_dff_A_XsDSl20W7_1),.clk(gclk));
	jdff dff_A_DB0ardjG5_1(.dout(w_dff_A_XsDSl20W7_1),.din(w_dff_A_DB0ardjG5_1),.clk(gclk));
	jdff dff_A_VRH3paYD6_1(.dout(w_dff_A_DB0ardjG5_1),.din(w_dff_A_VRH3paYD6_1),.clk(gclk));
	jdff dff_A_9YxXXqlF6_2(.dout(w_n614_3[2]),.din(w_dff_A_9YxXXqlF6_2),.clk(gclk));
	jdff dff_A_krrjJfzj6_2(.dout(w_dff_A_9YxXXqlF6_2),.din(w_dff_A_krrjJfzj6_2),.clk(gclk));
	jdff dff_A_vViKNCfp1_2(.dout(w_dff_A_krrjJfzj6_2),.din(w_dff_A_vViKNCfp1_2),.clk(gclk));
	jdff dff_A_VrIy1Jep0_2(.dout(w_dff_A_vViKNCfp1_2),.din(w_dff_A_VrIy1Jep0_2),.clk(gclk));
	jdff dff_A_1poxb7it2_2(.dout(w_dff_A_VrIy1Jep0_2),.din(w_dff_A_1poxb7it2_2),.clk(gclk));
	jdff dff_A_C1NEEAJW6_2(.dout(w_dff_A_1poxb7it2_2),.din(w_dff_A_C1NEEAJW6_2),.clk(gclk));
	jdff dff_A_toS1cSfk5_2(.dout(w_dff_A_C1NEEAJW6_2),.din(w_dff_A_toS1cSfk5_2),.clk(gclk));
	jdff dff_A_W2tX3q3y2_2(.dout(w_dff_A_toS1cSfk5_2),.din(w_dff_A_W2tX3q3y2_2),.clk(gclk));
	jdff dff_A_3NM5qXvP7_2(.dout(w_dff_A_W2tX3q3y2_2),.din(w_dff_A_3NM5qXvP7_2),.clk(gclk));
	jdff dff_A_bVZSU6GH8_1(.dout(w_n601_0[1]),.din(w_dff_A_bVZSU6GH8_1),.clk(gclk));
	jdff dff_A_1JsX1pGC1_1(.dout(w_dff_A_bVZSU6GH8_1),.din(w_dff_A_1JsX1pGC1_1),.clk(gclk));
	jdff dff_A_mG4NQv9y8_0(.dout(w_n600_1[0]),.din(w_dff_A_mG4NQv9y8_0),.clk(gclk));
	jdff dff_A_lFlKgL0f6_1(.dout(w_n600_1[1]),.din(w_dff_A_lFlKgL0f6_1),.clk(gclk));
	jdff dff_A_AD8s80ZX9_1(.dout(w_dff_A_lFlKgL0f6_1),.din(w_dff_A_AD8s80ZX9_1),.clk(gclk));
	jdff dff_B_lsLzXNMs1_0(.din(n599),.dout(w_dff_B_lsLzXNMs1_0),.clk(gclk));
	jdff dff_A_XqsxgXkg9_0(.dout(w_n598_0[0]),.din(w_dff_A_XqsxgXkg9_0),.clk(gclk));
	jdff dff_A_qiJW42G68_0(.dout(w_dff_A_XqsxgXkg9_0),.din(w_dff_A_qiJW42G68_0),.clk(gclk));
	jdff dff_A_3xum2mTS6_1(.dout(w_n571_1[1]),.din(w_dff_A_3xum2mTS6_1),.clk(gclk));
	jdff dff_A_Hi8ULcd96_1(.dout(w_dff_A_3xum2mTS6_1),.din(w_dff_A_Hi8ULcd96_1),.clk(gclk));
	jdff dff_A_FA6PyYmV0_1(.dout(w_dff_A_Hi8ULcd96_1),.din(w_dff_A_FA6PyYmV0_1),.clk(gclk));
	jdff dff_A_DAWbyz9E8_1(.dout(w_dff_A_FA6PyYmV0_1),.din(w_dff_A_DAWbyz9E8_1),.clk(gclk));
	jdff dff_A_i4C8CJMS1_1(.dout(w_dff_A_DAWbyz9E8_1),.din(w_dff_A_i4C8CJMS1_1),.clk(gclk));
	jdff dff_B_mRBBmtHJ5_0(.din(n589),.dout(w_dff_B_mRBBmtHJ5_0),.clk(gclk));
	jdff dff_B_dlM9eFUA4_0(.din(w_dff_B_mRBBmtHJ5_0),.dout(w_dff_B_dlM9eFUA4_0),.clk(gclk));
	jdff dff_A_PDfB6XMd4_1(.dout(w_n548_0[1]),.din(w_dff_A_PDfB6XMd4_1),.clk(gclk));
	jdff dff_A_uiIIcp3f6_1(.dout(w_dff_A_PDfB6XMd4_1),.din(w_dff_A_uiIIcp3f6_1),.clk(gclk));
	jdff dff_A_25sVWHOy3_1(.dout(w_n347_0[1]),.din(w_dff_A_25sVWHOy3_1),.clk(gclk));
	jdff dff_A_H4ms9W386_1(.dout(w_n189_1[1]),.din(w_dff_A_H4ms9W386_1),.clk(gclk));
	jdff dff_A_7dtRq2NS9_1(.dout(w_dff_A_H4ms9W386_1),.din(w_dff_A_7dtRq2NS9_1),.clk(gclk));
	jdff dff_A_yrHzOZpB0_0(.dout(w_n282_0[0]),.din(w_dff_A_yrHzOZpB0_0),.clk(gclk));
	jdff dff_B_F4cGoxfX8_1(.din(n525),.dout(w_dff_B_F4cGoxfX8_1),.clk(gclk));
	jdff dff_B_ei1IRPYu3_1(.din(n538),.dout(w_dff_B_ei1IRPYu3_1),.clk(gclk));
	jdff dff_B_O8VhvD2i9_1(.din(n324),.dout(w_dff_B_O8VhvD2i9_1),.clk(gclk));
	jdff dff_A_SG9uoOXf1_1(.dout(w_n323_0[1]),.din(w_dff_A_SG9uoOXf1_1),.clk(gclk));
	jdff dff_A_rDmAkkS04_2(.dout(w_n323_0[2]),.din(w_dff_A_rDmAkkS04_2),.clk(gclk));
	jdff dff_B_1RzhudOz1_1(.din(n314),.dout(w_dff_B_1RzhudOz1_1),.clk(gclk));
	jdff dff_B_llEH8sKq5_1(.din(w_dff_B_1RzhudOz1_1),.dout(w_dff_B_llEH8sKq5_1),.clk(gclk));
	jdff dff_A_gRveNVBj0_2(.dout(w_G20_3[2]),.din(w_dff_A_gRveNVBj0_2),.clk(gclk));
	jdff dff_A_QfY9ycPs7_1(.dout(w_n141_1[1]),.din(w_dff_A_QfY9ycPs7_1),.clk(gclk));
	jdff dff_A_nNSVdi6V0_2(.dout(w_n141_1[2]),.din(w_dff_A_nNSVdi6V0_2),.clk(gclk));
	jdff dff_A_rxnjzVgC9_0(.dout(w_n334_0[0]),.din(w_dff_A_rxnjzVgC9_0),.clk(gclk));
	jdff dff_A_xSMk7Iu53_0(.dout(w_dff_A_rxnjzVgC9_0),.din(w_dff_A_xSMk7Iu53_0),.clk(gclk));
	jdff dff_A_Qsh7UEam8_0(.dout(w_G169_2[0]),.din(w_dff_A_Qsh7UEam8_0),.clk(gclk));
	jdff dff_A_LS8Kd3zY6_1(.dout(w_G169_2[1]),.din(w_dff_A_LS8Kd3zY6_1),.clk(gclk));
	jdff dff_A_NH0586Nw4_1(.dout(w_dff_A_LS8Kd3zY6_1),.din(w_dff_A_NH0586Nw4_1),.clk(gclk));
	jdff dff_B_uHyrMRuq9_0(.din(n342),.dout(w_dff_B_uHyrMRuq9_0),.clk(gclk));
	jdff dff_A_Mfoln7al3_1(.dout(w_n321_0[1]),.din(w_dff_A_Mfoln7al3_1),.clk(gclk));
	jdff dff_A_JD62UApS0_1(.dout(w_dff_A_Mfoln7al3_1),.din(w_dff_A_JD62UApS0_1),.clk(gclk));
	jdff dff_B_BKOW30cU3_1(.din(n336),.dout(w_dff_B_BKOW30cU3_1),.clk(gclk));
	jdff dff_A_xSfVpV0A9_2(.dout(w_n72_1[2]),.din(w_dff_A_xSfVpV0A9_2),.clk(gclk));
	jdff dff_A_PPac0J2D5_2(.dout(w_dff_A_xSfVpV0A9_2),.din(w_dff_A_PPac0J2D5_2),.clk(gclk));
	jdff dff_A_jOenf4jn0_1(.dout(w_n72_0[1]),.din(w_dff_A_jOenf4jn0_1),.clk(gclk));
	jdff dff_A_jFkwn7bH5_1(.dout(w_dff_A_jOenf4jn0_1),.din(w_dff_A_jFkwn7bH5_1),.clk(gclk));
	jdff dff_A_PfwbTdmM6_1(.dout(w_dff_A_jFkwn7bH5_1),.din(w_dff_A_PfwbTdmM6_1),.clk(gclk));
	jdff dff_A_BXQjOJiv0_1(.dout(w_dff_A_PfwbTdmM6_1),.din(w_dff_A_BXQjOJiv0_1),.clk(gclk));
	jdff dff_A_Deq1UrMn3_2(.dout(w_n72_0[2]),.din(w_dff_A_Deq1UrMn3_2),.clk(gclk));
	jdff dff_A_AZmo76qN7_2(.dout(w_dff_A_Deq1UrMn3_2),.din(w_dff_A_AZmo76qN7_2),.clk(gclk));
	jdff dff_A_PxFH9qKR2_0(.dout(w_n315_0[0]),.din(w_dff_A_PxFH9qKR2_0),.clk(gclk));
	jdff dff_A_JSngJh1o7_0(.dout(w_dff_A_PxFH9qKR2_0),.din(w_dff_A_JSngJh1o7_0),.clk(gclk));
	jdff dff_A_lbfPEgwu3_2(.dout(w_n315_0[2]),.din(w_dff_A_lbfPEgwu3_2),.clk(gclk));
	jdff dff_A_aUuFFNoZ0_2(.dout(w_dff_A_lbfPEgwu3_2),.din(w_dff_A_aUuFFNoZ0_2),.clk(gclk));
	jdff dff_A_C6fhdDYB1_1(.dout(w_G33_8[1]),.din(w_dff_A_C6fhdDYB1_1),.clk(gclk));
	jdff dff_A_vSQVX5kt8_0(.dout(w_n313_0[0]),.din(w_dff_A_vSQVX5kt8_0),.clk(gclk));
	jdff dff_A_kHyPVeGO3_0(.dout(w_dff_A_vSQVX5kt8_0),.din(w_dff_A_kHyPVeGO3_0),.clk(gclk));
	jdff dff_A_eHGMUOgQ9_0(.dout(w_dff_A_kHyPVeGO3_0),.din(w_dff_A_eHGMUOgQ9_0),.clk(gclk));
	jdff dff_A_bXF8Ko468_0(.dout(w_n312_0[0]),.din(w_dff_A_bXF8Ko468_0),.clk(gclk));
	jdff dff_A_v2s6uZoF7_0(.dout(w_n310_0[0]),.din(w_dff_A_v2s6uZoF7_0),.clk(gclk));
	jdff dff_A_tnk2iPlc2_1(.dout(w_n309_0[1]),.din(w_dff_A_tnk2iPlc2_1),.clk(gclk));
	jdff dff_A_66o4pQgu8_1(.dout(w_dff_A_tnk2iPlc2_1),.din(w_dff_A_66o4pQgu8_1),.clk(gclk));
	jdff dff_A_gH22s1fJ8_0(.dout(w_n94_0[0]),.din(w_dff_A_gH22s1fJ8_0),.clk(gclk));
	jdff dff_A_nKjGZzcD3_0(.dout(w_dff_A_gH22s1fJ8_0),.din(w_dff_A_nKjGZzcD3_0),.clk(gclk));
	jdff dff_A_9TorVuzk2_0(.dout(w_dff_A_nKjGZzcD3_0),.din(w_dff_A_9TorVuzk2_0),.clk(gclk));
	jdff dff_A_A8RKeC036_0(.dout(w_G244_1[0]),.din(w_dff_A_A8RKeC036_0),.clk(gclk));
	jdff dff_A_STf4gIso3_0(.dout(w_n298_0[0]),.din(w_dff_A_STf4gIso3_0),.clk(gclk));
	jdff dff_A_VRn3UZHx9_0(.dout(w_dff_A_STf4gIso3_0),.din(w_dff_A_VRn3UZHx9_0),.clk(gclk));
	jdff dff_A_3gRB1EJk6_0(.dout(w_G190_3[0]),.din(w_dff_A_3gRB1EJk6_0),.clk(gclk));
	jdff dff_A_78XtRBs74_0(.dout(w_dff_A_3gRB1EJk6_0),.din(w_dff_A_78XtRBs74_0),.clk(gclk));
	jdff dff_A_NC3D814C8_1(.dout(w_G190_3[1]),.din(w_dff_A_NC3D814C8_1),.clk(gclk));
	jdff dff_A_5hmUbngm0_1(.dout(w_dff_A_NC3D814C8_1),.din(w_dff_A_5hmUbngm0_1),.clk(gclk));
	jdff dff_A_r7coMN1H0_1(.dout(w_n534_0[1]),.din(w_dff_A_r7coMN1H0_1),.clk(gclk));
	jdff dff_A_uDbIhnhQ0_1(.dout(w_n507_2[1]),.din(w_dff_A_uDbIhnhQ0_1),.clk(gclk));
	jdff dff_B_Z5BUScwi0_0(.din(n270),.dout(w_dff_B_Z5BUScwi0_0),.clk(gclk));
	jdff dff_B_teAz4mHt2_1(.din(n263),.dout(w_dff_B_teAz4mHt2_1),.clk(gclk));
	jdff dff_A_tbzq0ca04_0(.dout(w_n151_5[0]),.din(w_dff_A_tbzq0ca04_0),.clk(gclk));
	jdff dff_A_WZhaYv5b6_1(.dout(w_n261_0[1]),.din(w_dff_A_WZhaYv5b6_1),.clk(gclk));
	jdff dff_A_QrqwqCbg4_1(.dout(w_dff_A_WZhaYv5b6_1),.din(w_dff_A_QrqwqCbg4_1),.clk(gclk));
	jdff dff_A_jWhzem8v7_2(.dout(w_n261_0[2]),.din(w_dff_A_jWhzem8v7_2),.clk(gclk));
	jdff dff_A_k0Hrm9on7_2(.dout(w_dff_A_jWhzem8v7_2),.din(w_dff_A_k0Hrm9on7_2),.clk(gclk));
	jdff dff_A_1YteJ72n8_1(.dout(w_n283_0[1]),.din(w_dff_A_1YteJ72n8_1),.clk(gclk));
	jdff dff_A_Ae8V3D2h6_0(.dout(w_n168_3[0]),.din(w_dff_A_Ae8V3D2h6_0),.clk(gclk));
	jdff dff_A_F49VzkO16_2(.dout(w_n168_3[2]),.din(w_dff_A_F49VzkO16_2),.clk(gclk));
	jdff dff_A_ibTsKWpo0_2(.dout(w_dff_A_F49VzkO16_2),.din(w_dff_A_ibTsKWpo0_2),.clk(gclk));
	jdff dff_A_NUaPsx8q7_0(.dout(w_n269_0[0]),.din(w_dff_A_NUaPsx8q7_0),.clk(gclk));
	jdff dff_A_us0AcsJW6_0(.dout(w_dff_A_NUaPsx8q7_0),.din(w_dff_A_us0AcsJW6_0),.clk(gclk));
	jdff dff_A_ZwN0FY9s9_0(.dout(w_n262_0[0]),.din(w_dff_A_ZwN0FY9s9_0),.clk(gclk));
	jdff dff_A_PhnE6QKk6_0(.dout(w_dff_A_ZwN0FY9s9_0),.din(w_dff_A_PhnE6QKk6_0),.clk(gclk));
	jdff dff_A_oaqMv60T3_1(.dout(w_n262_0[1]),.din(w_dff_A_oaqMv60T3_1),.clk(gclk));
	jdff dff_A_gsERAYf14_1(.dout(w_dff_A_oaqMv60T3_1),.din(w_dff_A_gsERAYf14_1),.clk(gclk));
	jdff dff_A_ZW7DFe3L2_0(.dout(w_G33_9[0]),.din(w_dff_A_ZW7DFe3L2_0),.clk(gclk));
	jdff dff_A_kt8vfdUT2_1(.dout(w_G33_9[1]),.din(w_dff_A_kt8vfdUT2_1),.clk(gclk));
	jdff dff_A_EgbFodsF6_1(.dout(w_n260_0[1]),.din(w_dff_A_EgbFodsF6_1),.clk(gclk));
	jdff dff_A_Bn1ER3N95_1(.dout(w_G20_4[1]),.din(w_dff_A_Bn1ER3N95_1),.clk(gclk));
	jdff dff_A_IWTwbYrN4_2(.dout(w_G20_4[2]),.din(w_dff_A_IWTwbYrN4_2),.clk(gclk));
	jdff dff_A_aSoHVQ5s5_2(.dout(w_dff_A_IWTwbYrN4_2),.din(w_dff_A_aSoHVQ5s5_2),.clk(gclk));
	jdff dff_A_h7ftODI60_1(.dout(w_n257_0[1]),.din(w_dff_A_h7ftODI60_1),.clk(gclk));
	jdff dff_A_U3CmrLaq8_1(.dout(w_n256_0[1]),.din(w_dff_A_U3CmrLaq8_1),.clk(gclk));
	jdff dff_A_HOhlGm5x4_0(.dout(w_n251_0[0]),.din(w_dff_A_HOhlGm5x4_0),.clk(gclk));
	jdff dff_A_UjEXtY9A0_1(.dout(w_n250_0[1]),.din(w_dff_A_UjEXtY9A0_1),.clk(gclk));
	jdff dff_A_93Zd3l2g8_1(.dout(w_n247_0[1]),.din(w_dff_A_93Zd3l2g8_1),.clk(gclk));
	jdff dff_A_tgNieMpj3_0(.dout(w_G238_0[0]),.din(w_dff_A_tgNieMpj3_0),.clk(gclk));
	jdff dff_A_Ns6FvkDn8_0(.dout(w_dff_A_tgNieMpj3_0),.din(w_dff_A_Ns6FvkDn8_0),.clk(gclk));
	jdff dff_A_aXlyl3Fd0_0(.dout(w_dff_A_Ns6FvkDn8_0),.din(w_dff_A_aXlyl3Fd0_0),.clk(gclk));
	jdff dff_A_xYXY8fqB5_1(.dout(w_G238_0[1]),.din(w_dff_A_xYXY8fqB5_1),.clk(gclk));
	jdff dff_A_AwnHk9988_1(.dout(w_dff_A_xYXY8fqB5_1),.din(w_dff_A_AwnHk9988_1),.clk(gclk));
	jdff dff_A_YcSEk4u81_0(.dout(w_n243_0[0]),.din(w_dff_A_YcSEk4u81_0),.clk(gclk));
	jdff dff_A_2yVxaMzY3_1(.dout(w_G244_0[1]),.din(w_dff_A_2yVxaMzY3_1),.clk(gclk));
	jdff dff_A_oRkKDqT53_1(.dout(w_dff_A_2yVxaMzY3_1),.din(w_dff_A_oRkKDqT53_1),.clk(gclk));
	jdff dff_A_7U1UTgYe7_2(.dout(w_G244_0[2]),.din(w_dff_A_7U1UTgYe7_2),.clk(gclk));
	jdff dff_A_NS8jNmWs2_2(.dout(w_dff_A_7U1UTgYe7_2),.din(w_dff_A_NS8jNmWs2_2),.clk(gclk));
	jdff dff_A_O7ejGNVk3_1(.dout(w_n388_1[1]),.din(w_dff_A_O7ejGNVk3_1),.clk(gclk));
	jdff dff_A_CecK2pIg7_2(.dout(w_n388_1[2]),.din(w_dff_A_CecK2pIg7_2),.clk(gclk));
	jdff dff_A_upzh20eh1_2(.dout(w_dff_A_CecK2pIg7_2),.din(w_dff_A_upzh20eh1_2),.clk(gclk));
	jdff dff_A_CAWMciHy2_0(.dout(w_n520_0[0]),.din(w_dff_A_CAWMciHy2_0),.clk(gclk));
	jdff dff_A_Q2LPEikI5_0(.dout(w_dff_A_CAWMciHy2_0),.din(w_dff_A_Q2LPEikI5_0),.clk(gclk));
	jdff dff_A_b1wPHBan4_0(.dout(w_n604_1[0]),.din(w_dff_A_b1wPHBan4_0),.clk(gclk));
	jdff dff_A_LsbrMTkE4_0(.dout(w_dff_A_b1wPHBan4_0),.din(w_dff_A_LsbrMTkE4_0),.clk(gclk));
	jdff dff_A_60vNIaI08_1(.dout(w_n604_1[1]),.din(w_dff_A_60vNIaI08_1),.clk(gclk));
	jdff dff_A_WxdUJPLt4_1(.dout(w_dff_A_60vNIaI08_1),.din(w_dff_A_WxdUJPLt4_1),.clk(gclk));
	jdff dff_A_hDEczb3X8_0(.dout(w_n861_0[0]),.din(w_dff_A_hDEczb3X8_0),.clk(gclk));
	jdff dff_B_vHNzx2Rh3_0(.din(n858),.dout(w_dff_B_vHNzx2Rh3_0),.clk(gclk));
	jdff dff_A_9bQoZvaZ9_2(.dout(w_n579_0[2]),.din(w_dff_A_9bQoZvaZ9_2),.clk(gclk));
	jdff dff_B_FIelMW6t1_0(.din(n578),.dout(w_dff_B_FIelMW6t1_0),.clk(gclk));
	jdff dff_B_2DsSV5zE4_0(.din(w_dff_B_FIelMW6t1_0),.dout(w_dff_B_2DsSV5zE4_0),.clk(gclk));
	jdff dff_B_w9d2YWfE9_0(.din(w_dff_B_2DsSV5zE4_0),.dout(w_dff_B_w9d2YWfE9_0),.clk(gclk));
	jdff dff_A_7UwZUzIm3_0(.dout(w_n571_2[0]),.din(w_dff_A_7UwZUzIm3_0),.clk(gclk));
	jdff dff_A_iQuhWqzD7_0(.dout(w_dff_A_7UwZUzIm3_0),.din(w_dff_A_iQuhWqzD7_0),.clk(gclk));
	jdff dff_A_Ild9kzuP5_1(.dout(w_n571_0[1]),.din(w_dff_A_Ild9kzuP5_1),.clk(gclk));
	jdff dff_A_eM79DCKB4_1(.dout(w_dff_A_Ild9kzuP5_1),.din(w_dff_A_eM79DCKB4_1),.clk(gclk));
	jdff dff_A_96MVLQZu7_2(.dout(w_n571_0[2]),.din(w_dff_A_96MVLQZu7_2),.clk(gclk));
	jdff dff_A_Jz9hUAx84_2(.dout(w_dff_A_96MVLQZu7_2),.din(w_dff_A_Jz9hUAx84_2),.clk(gclk));
	jdff dff_B_7cE0JC4U6_3(.din(n571),.dout(w_dff_B_7cE0JC4U6_3),.clk(gclk));
	jdff dff_B_i6tp0XE54_3(.din(w_dff_B_7cE0JC4U6_3),.dout(w_dff_B_i6tp0XE54_3),.clk(gclk));
	jdff dff_B_Q838d2J84_3(.din(w_dff_B_i6tp0XE54_3),.dout(w_dff_B_Q838d2J84_3),.clk(gclk));
	jdff dff_B_xJUEBMqN3_3(.din(w_dff_B_Q838d2J84_3),.dout(w_dff_B_xJUEBMqN3_3),.clk(gclk));
	jdff dff_B_kxKU4Zyf9_3(.din(w_dff_B_xJUEBMqN3_3),.dout(w_dff_B_kxKU4Zyf9_3),.clk(gclk));
	jdff dff_A_0qCPDfMR7_1(.dout(w_n567_5[1]),.din(w_dff_A_0qCPDfMR7_1),.clk(gclk));
	jdff dff_A_APNkAsNs8_1(.dout(w_dff_A_0qCPDfMR7_1),.din(w_dff_A_APNkAsNs8_1),.clk(gclk));
	jdff dff_A_TRlDMbyE9_1(.dout(w_dff_A_APNkAsNs8_1),.din(w_dff_A_TRlDMbyE9_1),.clk(gclk));
	jdff dff_A_OzLmUVZf7_1(.dout(w_dff_A_TRlDMbyE9_1),.din(w_dff_A_OzLmUVZf7_1),.clk(gclk));
	jdff dff_A_FurO07le1_1(.dout(w_dff_A_OzLmUVZf7_1),.din(w_dff_A_FurO07le1_1),.clk(gclk));
	jdff dff_A_ogos4tL26_1(.dout(w_dff_A_FurO07le1_1),.din(w_dff_A_ogos4tL26_1),.clk(gclk));
	jdff dff_A_Me1fhYuZ2_0(.dout(w_n570_0[0]),.din(w_dff_A_Me1fhYuZ2_0),.clk(gclk));
	jdff dff_A_uNIKy0Cp2_1(.dout(w_n242_0[1]),.din(w_dff_A_uNIKy0Cp2_1),.clk(gclk));
	jdff dff_A_ZMKhAMUR0_1(.dout(w_dff_A_uNIKy0Cp2_1),.din(w_dff_A_ZMKhAMUR0_1),.clk(gclk));
	jdff dff_A_HDWYnpOB9_2(.dout(w_n242_0[2]),.din(w_dff_A_HDWYnpOB9_2),.clk(gclk));
	jdff dff_A_1279TGH46_1(.dout(w_n238_0[1]),.din(w_dff_A_1279TGH46_1),.clk(gclk));
	jdff dff_A_TfJltKmd2_1(.dout(w_n237_0[1]),.din(w_dff_A_TfJltKmd2_1),.clk(gclk));
	jdff dff_A_9a3Em77c0_1(.dout(w_dff_A_TfJltKmd2_1),.din(w_dff_A_9a3Em77c0_1),.clk(gclk));
	jdff dff_A_gBaa83Ed2_1(.dout(w_n234_0[1]),.din(w_dff_A_gBaa83Ed2_1),.clk(gclk));
	jdff dff_A_fS0LlvZK6_1(.dout(w_dff_A_gBaa83Ed2_1),.din(w_dff_A_fS0LlvZK6_1),.clk(gclk));
	jdff dff_A_2WoCuG5J3_1(.dout(w_dff_A_fS0LlvZK6_1),.din(w_dff_A_2WoCuG5J3_1),.clk(gclk));
	jdff dff_B_VZM5CY1Z9_1(.din(n226),.dout(w_dff_B_VZM5CY1Z9_1),.clk(gclk));
	jdff dff_A_5HXFfcAo9_1(.dout(w_n229_0[1]),.din(w_dff_A_5HXFfcAo9_1),.clk(gclk));
	jdff dff_B_yMYeWhuq7_1(.din(n227),.dout(w_dff_B_yMYeWhuq7_1),.clk(gclk));
	jdff dff_B_mypaOipd7_1(.din(w_dff_B_yMYeWhuq7_1),.dout(w_dff_B_mypaOipd7_1),.clk(gclk));
	jdff dff_A_OlooEsLk1_0(.dout(w_n224_1[0]),.din(w_dff_A_OlooEsLk1_0),.clk(gclk));
	jdff dff_A_MDqOfozP8_2(.dout(w_n224_0[2]),.din(w_dff_A_MDqOfozP8_2),.clk(gclk));
	jdff dff_B_AiBGyhXP0_0(.din(n223),.dout(w_dff_B_AiBGyhXP0_0),.clk(gclk));
	jdff dff_B_8kuGAAZk2_1(.din(n217),.dout(w_dff_B_8kuGAAZk2_1),.clk(gclk));
	jdff dff_A_qAdhCfa83_1(.dout(w_n218_0[1]),.din(w_dff_A_qAdhCfa83_1),.clk(gclk));
	jdff dff_A_zY3WHwLO9_0(.dout(w_n141_2[0]),.din(w_dff_A_zY3WHwLO9_0),.clk(gclk));
	jdff dff_B_LiSmy9oS4_0(.din(n216),.dout(w_dff_B_LiSmy9oS4_0),.clk(gclk));
	jdff dff_A_vevyfFaW1_0(.dout(w_n81_1[0]),.din(w_dff_A_vevyfFaW1_0),.clk(gclk));
	jdff dff_A_UYDQdNuH7_1(.dout(w_n213_0[1]),.din(w_dff_A_UYDQdNuH7_1),.clk(gclk));
	jdff dff_A_E8cAH0dG6_1(.dout(w_n212_0[1]),.din(w_dff_A_E8cAH0dG6_1),.clk(gclk));
	jdff dff_A_bRRjJPyT6_1(.dout(w_dff_A_E8cAH0dG6_1),.din(w_dff_A_bRRjJPyT6_1),.clk(gclk));
	jdff dff_A_REIo9ffo7_0(.dout(w_n207_0[0]),.din(w_dff_A_REIo9ffo7_0),.clk(gclk));
	jdff dff_A_Z1rKLJEN2_2(.dout(w_n84_1[2]),.din(w_dff_A_Z1rKLJEN2_2),.clk(gclk));
	jdff dff_A_c6nYiNQz8_1(.dout(w_n84_0[1]),.din(w_dff_A_c6nYiNQz8_1),.clk(gclk));
	jdff dff_A_oAkhjJVX7_2(.dout(w_n84_0[2]),.din(w_dff_A_oAkhjJVX7_2),.clk(gclk));
	jdff dff_A_T7sl5B3r6_0(.dout(w_G250_0[0]),.din(w_dff_A_T7sl5B3r6_0),.clk(gclk));
	jdff dff_A_O35QWYi73_0(.dout(w_dff_A_T7sl5B3r6_0),.din(w_dff_A_O35QWYi73_0),.clk(gclk));
	jdff dff_A_WdejfyvY0_1(.dout(w_n202_0[1]),.din(w_dff_A_WdejfyvY0_1),.clk(gclk));
	jdff dff_A_aaQzLjKd6_1(.dout(w_n201_0[1]),.din(w_dff_A_aaQzLjKd6_1),.clk(gclk));
	jdff dff_A_nANvYK136_1(.dout(w_dff_A_aaQzLjKd6_1),.din(w_dff_A_nANvYK136_1),.clk(gclk));
	jdff dff_A_38YAPIYS1_0(.dout(w_n168_4[0]),.din(w_dff_A_38YAPIYS1_0),.clk(gclk));
	jdff dff_A_TIDzhtUv3_0(.dout(w_dff_A_38YAPIYS1_0),.din(w_dff_A_TIDzhtUv3_0),.clk(gclk));
	jdff dff_A_TwV63DNe3_1(.dout(w_n168_4[1]),.din(w_dff_A_TwV63DNe3_1),.clk(gclk));
	jdff dff_A_J55No7Ox2_1(.dout(w_dff_A_TwV63DNe3_1),.din(w_dff_A_J55No7Ox2_1),.clk(gclk));
	jdff dff_A_iqzJtzSj0_0(.dout(w_n199_0[0]),.din(w_dff_A_iqzJtzSj0_0),.clk(gclk));
	jdff dff_A_aLVZsU2V1_0(.dout(w_dff_A_iqzJtzSj0_0),.din(w_dff_A_aLVZsU2V1_0),.clk(gclk));
	jdff dff_A_b8n47nWS4_0(.dout(w_dff_A_aLVZsU2V1_0),.din(w_dff_A_b8n47nWS4_0),.clk(gclk));
	jdff dff_A_GRRwwvD30_2(.dout(w_n199_0[2]),.din(w_dff_A_GRRwwvD30_2),.clk(gclk));
	jdff dff_B_wjJvFzl57_3(.din(n199),.dout(w_dff_B_wjJvFzl57_3),.clk(gclk));
	jdff dff_B_bN40Ll332_3(.din(w_dff_B_wjJvFzl57_3),.dout(w_dff_B_bN40Ll332_3),.clk(gclk));
	jdff dff_B_vmS78ivG2_3(.din(w_dff_B_bN40Ll332_3),.dout(w_dff_B_vmS78ivG2_3),.clk(gclk));
	jdff dff_B_H7cRpZho8_3(.din(w_dff_B_vmS78ivG2_3),.dout(w_dff_B_H7cRpZho8_3),.clk(gclk));
	jdff dff_B_By5IOUUi6_3(.din(w_dff_B_H7cRpZho8_3),.dout(w_dff_B_By5IOUUi6_3),.clk(gclk));
	jdff dff_B_KU0nt64i4_3(.din(w_dff_B_By5IOUUi6_3),.dout(w_dff_B_KU0nt64i4_3),.clk(gclk));
	jdff dff_A_ihw0ivVJ5_0(.dout(w_n577_0[0]),.din(w_dff_A_ihw0ivVJ5_0),.clk(gclk));
	jdff dff_A_C61XykJj3_0(.dout(w_dff_A_ihw0ivVJ5_0),.din(w_dff_A_C61XykJj3_0),.clk(gclk));
	jdff dff_B_JgsaM3to7_2(.din(n1164),.dout(w_dff_B_JgsaM3to7_2),.clk(gclk));
	jdff dff_B_Ig6Xmlhb8_2(.din(w_dff_B_JgsaM3to7_2),.dout(w_dff_B_Ig6Xmlhb8_2),.clk(gclk));
	jdff dff_B_EwQVB6tX8_2(.din(w_dff_B_Ig6Xmlhb8_2),.dout(w_dff_B_EwQVB6tX8_2),.clk(gclk));
	jdff dff_B_DqFvCkPD9_2(.din(w_dff_B_EwQVB6tX8_2),.dout(w_dff_B_DqFvCkPD9_2),.clk(gclk));
	jdff dff_B_0I1CikA97_1(.din(n617),.dout(w_dff_B_0I1CikA97_1),.clk(gclk));
	jdff dff_B_gI3qsLLX6_0(.din(n698),.dout(w_dff_B_gI3qsLLX6_0),.clk(gclk));
	jdff dff_B_VRcvTawS5_0(.din(n697),.dout(w_dff_B_VRcvTawS5_0),.clk(gclk));
	jdff dff_B_kPQnTKnU7_0(.din(w_dff_B_VRcvTawS5_0),.dout(w_dff_B_kPQnTKnU7_0),.clk(gclk));
	jdff dff_B_cEH9gJjW1_0(.din(n694),.dout(w_dff_B_cEH9gJjW1_0),.clk(gclk));
	jdff dff_B_DDLmV1sL9_0(.din(w_dff_B_cEH9gJjW1_0),.dout(w_dff_B_DDLmV1sL9_0),.clk(gclk));
	jdff dff_A_mBfYHKxY7_0(.dout(w_n692_0[0]),.din(w_dff_A_mBfYHKxY7_0),.clk(gclk));
	jdff dff_A_SmwWHC6v9_0(.dout(w_n153_4[0]),.din(w_dff_A_SmwWHC6v9_0),.clk(gclk));
	jdff dff_A_Zg11fxW30_0(.dout(w_dff_A_SmwWHC6v9_0),.din(w_dff_A_Zg11fxW30_0),.clk(gclk));
	jdff dff_A_vkCkv83m6_0(.dout(w_dff_A_Zg11fxW30_0),.din(w_dff_A_vkCkv83m6_0),.clk(gclk));
	jdff dff_A_aRrmc5Aj4_0(.dout(w_dff_A_vkCkv83m6_0),.din(w_dff_A_aRrmc5Aj4_0),.clk(gclk));
	jdff dff_A_QedZhUyP9_0(.dout(w_dff_A_aRrmc5Aj4_0),.din(w_dff_A_QedZhUyP9_0),.clk(gclk));
	jdff dff_A_PMwywllJ0_0(.dout(w_dff_A_QedZhUyP9_0),.din(w_dff_A_PMwywllJ0_0),.clk(gclk));
	jdff dff_A_5yT7bRBN7_1(.dout(w_n153_4[1]),.din(w_dff_A_5yT7bRBN7_1),.clk(gclk));
	jdff dff_A_QZArltnf9_1(.dout(w_dff_A_5yT7bRBN7_1),.din(w_dff_A_QZArltnf9_1),.clk(gclk));
	jdff dff_A_BXgTb1ev9_1(.dout(w_dff_A_QZArltnf9_1),.din(w_dff_A_BXgTb1ev9_1),.clk(gclk));
	jdff dff_A_PGw1wZYf4_1(.dout(w_dff_A_BXgTb1ev9_1),.din(w_dff_A_PGw1wZYf4_1),.clk(gclk));
	jdff dff_A_z7nYyzmH2_1(.dout(w_dff_A_PGw1wZYf4_1),.din(w_dff_A_z7nYyzmH2_1),.clk(gclk));
	jdff dff_A_3oPoLBjJ4_0(.dout(w_G355_0),.din(w_dff_A_3oPoLBjJ4_0),.clk(gclk));
	jdff dff_A_h1B3mJfH4_2(.dout(w_n81_0[2]),.din(w_dff_A_h1B3mJfH4_2),.clk(gclk));
	jdff dff_A_LdOBTXp65_2(.dout(w_dff_A_h1B3mJfH4_2),.din(w_dff_A_LdOBTXp65_2),.clk(gclk));
	jdff dff_A_VjANystY2_2(.dout(w_dff_A_LdOBTXp65_2),.din(w_dff_A_VjANystY2_2),.clk(gclk));
	jdff dff_A_TZCEIUvz2_0(.dout(w_G107_4[0]),.din(w_dff_A_TZCEIUvz2_0),.clk(gclk));
	jdff dff_A_hHIrK42a3_0(.dout(w_dff_A_TZCEIUvz2_0),.din(w_dff_A_hHIrK42a3_0),.clk(gclk));
	jdff dff_A_z5eoBffp8_0(.dout(w_dff_A_hHIrK42a3_0),.din(w_dff_A_z5eoBffp8_0),.clk(gclk));
	jdff dff_A_ykQuhNr48_0(.dout(w_dff_A_z5eoBffp8_0),.din(w_dff_A_ykQuhNr48_0),.clk(gclk));
	jdff dff_A_Ga9HDaAh5_0(.dout(w_dff_A_ykQuhNr48_0),.din(w_dff_A_Ga9HDaAh5_0),.clk(gclk));
	jdff dff_A_LArgObzU8_0(.dout(w_dff_A_Ga9HDaAh5_0),.din(w_dff_A_LArgObzU8_0),.clk(gclk));
	jdff dff_A_kB4WD2uz7_1(.dout(w_G107_1[1]),.din(w_dff_A_kB4WD2uz7_1),.clk(gclk));
	jdff dff_A_XEMYXWQY2_1(.dout(w_dff_A_kB4WD2uz7_1),.din(w_dff_A_XEMYXWQY2_1),.clk(gclk));
	jdff dff_A_so2b6Mk06_1(.dout(w_dff_A_XEMYXWQY2_1),.din(w_dff_A_so2b6Mk06_1),.clk(gclk));
	jdff dff_A_Jw4UgDiI5_2(.dout(w_G107_1[2]),.din(w_dff_A_Jw4UgDiI5_2),.clk(gclk));
	jdff dff_A_8EDbM3VO1_2(.dout(w_dff_A_Jw4UgDiI5_2),.din(w_dff_A_8EDbM3VO1_2),.clk(gclk));
	jdff dff_A_YdIp8JhS8_2(.dout(w_dff_A_8EDbM3VO1_2),.din(w_dff_A_YdIp8JhS8_2),.clk(gclk));
	jdff dff_A_Tev3nFhw1_1(.dout(w_n80_0[1]),.din(w_dff_A_Tev3nFhw1_1),.clk(gclk));
	jdff dff_A_hIrgyG9Q4_1(.dout(w_dff_A_Tev3nFhw1_1),.din(w_dff_A_hIrgyG9Q4_1),.clk(gclk));
	jdff dff_A_eqyl31wS2_2(.dout(w_n80_0[2]),.din(w_dff_A_eqyl31wS2_2),.clk(gclk));
	jdff dff_A_n1QeoCI66_2(.dout(w_dff_A_eqyl31wS2_2),.din(w_dff_A_n1QeoCI66_2),.clk(gclk));
	jdff dff_A_V8PP1KKa7_2(.dout(w_dff_A_n1QeoCI66_2),.din(w_dff_A_V8PP1KKa7_2),.clk(gclk));
	jdff dff_A_nmcIZyGl1_2(.dout(w_dff_A_V8PP1KKa7_2),.din(w_dff_A_nmcIZyGl1_2),.clk(gclk));
	jdff dff_A_8SqCKDX28_0(.dout(w_n79_1[0]),.din(w_dff_A_8SqCKDX28_0),.clk(gclk));
	jdff dff_A_Yu5PzgA72_0(.dout(w_dff_A_8SqCKDX28_0),.din(w_dff_A_Yu5PzgA72_0),.clk(gclk));
	jdff dff_A_kVVVfSmH2_0(.dout(w_dff_A_Yu5PzgA72_0),.din(w_dff_A_kVVVfSmH2_0),.clk(gclk));
	jdff dff_A_ObjgFuti1_0(.dout(w_dff_A_kVVVfSmH2_0),.din(w_dff_A_ObjgFuti1_0),.clk(gclk));
	jdff dff_A_98rMngqj2_2(.dout(w_n79_1[2]),.din(w_dff_A_98rMngqj2_2),.clk(gclk));
	jdff dff_A_0BCjYyTD0_1(.dout(w_n79_0[1]),.din(w_dff_A_0BCjYyTD0_1),.clk(gclk));
	jdff dff_A_yOUXbtIP7_1(.dout(w_dff_A_0BCjYyTD0_1),.din(w_dff_A_yOUXbtIP7_1),.clk(gclk));
	jdff dff_A_1FSyIZIT2_0(.dout(w_G87_3[0]),.din(w_dff_A_1FSyIZIT2_0),.clk(gclk));
	jdff dff_B_bMygN5jQ5_1(.din(n683),.dout(w_dff_B_bMygN5jQ5_1),.clk(gclk));
	jdff dff_B_eXnXffhz6_1(.din(w_dff_B_bMygN5jQ5_1),.dout(w_dff_B_eXnXffhz6_1),.clk(gclk));
	jdff dff_B_NI5hjL856_1(.din(w_dff_B_eXnXffhz6_1),.dout(w_dff_B_NI5hjL856_1),.clk(gclk));
	jdff dff_B_wHCIhoNy1_1(.din(w_dff_B_NI5hjL856_1),.dout(w_dff_B_wHCIhoNy1_1),.clk(gclk));
	jdff dff_A_UKI5si2f1_2(.dout(w_n75_0[2]),.din(w_dff_A_UKI5si2f1_2),.clk(gclk));
	jdff dff_A_Qo9GQida4_2(.dout(w_dff_A_UKI5si2f1_2),.din(w_dff_A_Qo9GQida4_2),.clk(gclk));
	jdff dff_A_4dQJKf2J1_2(.dout(w_dff_A_Qo9GQida4_2),.din(w_dff_A_4dQJKf2J1_2),.clk(gclk));
	jdff dff_A_EhOeGe6S7_2(.dout(w_dff_A_4dQJKf2J1_2),.din(w_dff_A_EhOeGe6S7_2),.clk(gclk));
	jdff dff_A_SxkNvj3H7_2(.dout(w_n74_0[2]),.din(w_dff_A_SxkNvj3H7_2),.clk(gclk));
	jdff dff_A_j14lyMv84_2(.dout(w_dff_A_SxkNvj3H7_2),.din(w_dff_A_j14lyMv84_2),.clk(gclk));
	jdff dff_A_GYJ1jS5R7_2(.dout(w_dff_A_j14lyMv84_2),.din(w_dff_A_GYJ1jS5R7_2),.clk(gclk));
	jdff dff_A_KgkWMurd5_2(.dout(w_dff_A_GYJ1jS5R7_2),.din(w_dff_A_KgkWMurd5_2),.clk(gclk));
	jdff dff_A_D9G1yZ2a1_0(.dout(w_G33_6[0]),.din(w_dff_A_D9G1yZ2a1_0),.clk(gclk));
	jdff dff_A_SIvmIlwI9_0(.dout(w_dff_A_D9G1yZ2a1_0),.din(w_dff_A_SIvmIlwI9_0),.clk(gclk));
	jdff dff_A_UFHF0I219_0(.dout(w_dff_A_SIvmIlwI9_0),.din(w_dff_A_UFHF0I219_0),.clk(gclk));
	jdff dff_A_9KKD5hdf2_0(.dout(w_dff_A_UFHF0I219_0),.din(w_dff_A_9KKD5hdf2_0),.clk(gclk));
	jdff dff_A_MZfX7DFR6_0(.dout(w_dff_A_9KKD5hdf2_0),.din(w_dff_A_MZfX7DFR6_0),.clk(gclk));
	jdff dff_A_57ZRTMa09_0(.dout(w_dff_A_MZfX7DFR6_0),.din(w_dff_A_57ZRTMa09_0),.clk(gclk));
	jdff dff_A_PVZi9aMd7_1(.dout(w_G33_6[1]),.din(w_dff_A_PVZi9aMd7_1),.clk(gclk));
	jdff dff_A_a4I94ztY4_1(.dout(w_dff_A_PVZi9aMd7_1),.din(w_dff_A_a4I94ztY4_1),.clk(gclk));
	jdff dff_A_ZslAtP5G6_1(.dout(w_dff_A_a4I94ztY4_1),.din(w_dff_A_ZslAtP5G6_1),.clk(gclk));
	jdff dff_A_iVfLRPJb5_0(.dout(w_G33_1[0]),.din(w_dff_A_iVfLRPJb5_0),.clk(gclk));
	jdff dff_A_3Ekhpmm29_0(.dout(w_dff_A_iVfLRPJb5_0),.din(w_dff_A_3Ekhpmm29_0),.clk(gclk));
	jdff dff_A_LPoGvtSe4_1(.dout(w_G33_1[1]),.din(w_dff_A_LPoGvtSe4_1),.clk(gclk));
	jdff dff_A_wUc9r8FB4_1(.dout(w_dff_A_LPoGvtSe4_1),.din(w_dff_A_wUc9r8FB4_1),.clk(gclk));
	jdff dff_A_acbnPoFk7_1(.dout(w_n134_0[1]),.din(w_dff_A_acbnPoFk7_1),.clk(gclk));
	jdff dff_A_165wfq2N1_0(.dout(w_G77_4[0]),.din(w_dff_A_165wfq2N1_0),.clk(gclk));
	jdff dff_A_KkFJ5Hfk9_1(.dout(w_G77_1[1]),.din(w_dff_A_KkFJ5Hfk9_1),.clk(gclk));
	jdff dff_A_Ukt0XTUJ4_1(.dout(w_dff_A_KkFJ5Hfk9_1),.din(w_dff_A_Ukt0XTUJ4_1),.clk(gclk));
	jdff dff_A_EiFIn5iG2_1(.dout(w_dff_A_Ukt0XTUJ4_1),.din(w_dff_A_EiFIn5iG2_1),.clk(gclk));
	jdff dff_A_aC0WX6qI9_1(.dout(w_dff_A_EiFIn5iG2_1),.din(w_dff_A_aC0WX6qI9_1),.clk(gclk));
	jdff dff_A_54F53hGA1_0(.dout(w_G68_5[0]),.din(w_dff_A_54F53hGA1_0),.clk(gclk));
	jdff dff_A_fXJA9ANq0_2(.dout(w_G68_1[2]),.din(w_dff_A_fXJA9ANq0_2),.clk(gclk));
	jdff dff_A_0ZrkUSCb5_2(.dout(w_dff_A_fXJA9ANq0_2),.din(w_dff_A_0ZrkUSCb5_2),.clk(gclk));
	jdff dff_A_pbAlY6TH8_2(.dout(w_dff_A_0ZrkUSCb5_2),.din(w_dff_A_pbAlY6TH8_2),.clk(gclk));
	jdff dff_A_vd9Cswqp1_0(.dout(w_G58_5[0]),.din(w_dff_A_vd9Cswqp1_0),.clk(gclk));
	jdff dff_A_zHuTCMKi6_1(.dout(w_G50_5[1]),.din(w_dff_A_zHuTCMKi6_1),.clk(gclk));
	jdff dff_A_bqMO1Dy82_1(.dout(w_dff_A_zHuTCMKi6_1),.din(w_dff_A_bqMO1Dy82_1),.clk(gclk));
	jdff dff_A_XaU3ZVoN5_1(.dout(w_dff_A_bqMO1Dy82_1),.din(w_dff_A_XaU3ZVoN5_1),.clk(gclk));
	jdff dff_A_VxkHbEoJ1_0(.dout(w_n352_1[0]),.din(w_dff_A_VxkHbEoJ1_0),.clk(gclk));
	jdff dff_A_9v9LOQ0m0_1(.dout(w_n352_0[1]),.din(w_dff_A_9v9LOQ0m0_1),.clk(gclk));
	jdff dff_A_jTYMQv605_1(.dout(w_dff_A_9v9LOQ0m0_1),.din(w_dff_A_jTYMQv605_1),.clk(gclk));
	jdff dff_A_vAwRVnA50_1(.dout(w_dff_A_jTYMQv605_1),.din(w_dff_A_vAwRVnA50_1),.clk(gclk));
	jdff dff_A_6yFqqlZp9_1(.dout(w_dff_A_vAwRVnA50_1),.din(w_dff_A_6yFqqlZp9_1),.clk(gclk));
	jdff dff_A_9wmDGhK17_2(.dout(w_n352_0[2]),.din(w_dff_A_9wmDGhK17_2),.clk(gclk));
	jdff dff_A_OgC0qXEc7_2(.dout(w_dff_A_9wmDGhK17_2),.din(w_dff_A_OgC0qXEc7_2),.clk(gclk));
	jdff dff_A_h72eUwTZ4_2(.dout(w_dff_A_OgC0qXEc7_2),.din(w_dff_A_h72eUwTZ4_2),.clk(gclk));
	jdff dff_A_kCrYY3sM9_1(.dout(w_n682_0[1]),.din(w_dff_A_kCrYY3sM9_1),.clk(gclk));
	jdff dff_A_9KiZmsk92_1(.dout(w_dff_A_kCrYY3sM9_1),.din(w_dff_A_9KiZmsk92_1),.clk(gclk));
	jdff dff_A_6Trf0unK8_1(.dout(w_dff_A_9KiZmsk92_1),.din(w_dff_A_6Trf0unK8_1),.clk(gclk));
	jdff dff_A_UECuCKLI4_1(.dout(w_dff_A_6Trf0unK8_1),.din(w_dff_A_UECuCKLI4_1),.clk(gclk));
	jdff dff_A_bm8Y9ewL9_1(.dout(w_n680_4[1]),.din(w_dff_A_bm8Y9ewL9_1),.clk(gclk));
	jdff dff_A_d3NLE3HZ0_1(.dout(w_dff_A_bm8Y9ewL9_1),.din(w_dff_A_d3NLE3HZ0_1),.clk(gclk));
	jdff dff_A_zVBPWxrM0_1(.dout(w_dff_A_d3NLE3HZ0_1),.din(w_dff_A_zVBPWxrM0_1),.clk(gclk));
	jdff dff_A_6mxnApiT3_1(.dout(w_dff_A_zVBPWxrM0_1),.din(w_dff_A_6mxnApiT3_1),.clk(gclk));
	jdff dff_A_5qPU88WJ5_1(.dout(w_dff_A_6mxnApiT3_1),.din(w_dff_A_5qPU88WJ5_1),.clk(gclk));
	jdff dff_A_xLUenMFY1_1(.dout(w_dff_A_5qPU88WJ5_1),.din(w_dff_A_xLUenMFY1_1),.clk(gclk));
	jdff dff_A_ygevY0Ts1_1(.dout(w_dff_A_xLUenMFY1_1),.din(w_dff_A_ygevY0Ts1_1),.clk(gclk));
	jdff dff_A_XlRzNeBV1_1(.dout(w_dff_A_ygevY0Ts1_1),.din(w_dff_A_XlRzNeBV1_1),.clk(gclk));
	jdff dff_A_PA2EIylc3_1(.dout(w_n680_1[1]),.din(w_dff_A_PA2EIylc3_1),.clk(gclk));
	jdff dff_A_YpPsNNyi0_1(.dout(w_dff_A_PA2EIylc3_1),.din(w_dff_A_YpPsNNyi0_1),.clk(gclk));
	jdff dff_A_KHRD8akD2_1(.dout(w_dff_A_YpPsNNyi0_1),.din(w_dff_A_KHRD8akD2_1),.clk(gclk));
	jdff dff_A_0f2aY4Fl4_1(.dout(w_dff_A_KHRD8akD2_1),.din(w_dff_A_0f2aY4Fl4_1),.clk(gclk));
	jdff dff_A_kzmIfMe73_1(.dout(w_dff_A_0f2aY4Fl4_1),.din(w_dff_A_kzmIfMe73_1),.clk(gclk));
	jdff dff_A_UpoNaDfn7_1(.dout(w_dff_A_kzmIfMe73_1),.din(w_dff_A_UpoNaDfn7_1),.clk(gclk));
	jdff dff_A_eXb4slFv4_1(.dout(w_dff_A_UpoNaDfn7_1),.din(w_dff_A_eXb4slFv4_1),.clk(gclk));
	jdff dff_A_0vEhVMaq7_1(.dout(w_n680_0[1]),.din(w_dff_A_0vEhVMaq7_1),.clk(gclk));
	jdff dff_A_1t4dqa8B4_1(.dout(w_dff_A_0vEhVMaq7_1),.din(w_dff_A_1t4dqa8B4_1),.clk(gclk));
	jdff dff_A_ofAzEnEg9_1(.dout(w_dff_A_1t4dqa8B4_1),.din(w_dff_A_ofAzEnEg9_1),.clk(gclk));
	jdff dff_A_SQbxlJ3h6_1(.dout(w_dff_A_ofAzEnEg9_1),.din(w_dff_A_SQbxlJ3h6_1),.clk(gclk));
	jdff dff_A_1y3mWi0F2_1(.dout(w_dff_A_SQbxlJ3h6_1),.din(w_dff_A_1y3mWi0F2_1),.clk(gclk));
	jdff dff_A_cl3wp3JZ1_1(.dout(w_G169_1[1]),.din(w_dff_A_cl3wp3JZ1_1),.clk(gclk));
	jdff dff_A_a77xGqki2_1(.dout(w_dff_A_cl3wp3JZ1_1),.din(w_dff_A_a77xGqki2_1),.clk(gclk));
	jdff dff_A_CLpnZf594_1(.dout(w_dff_A_a77xGqki2_1),.din(w_dff_A_CLpnZf594_1),.clk(gclk));
	jdff dff_A_CHwOrggI4_1(.dout(w_dff_A_CLpnZf594_1),.din(w_dff_A_CHwOrggI4_1),.clk(gclk));
	jdff dff_A_1t47kqJw6_1(.dout(w_dff_A_CHwOrggI4_1),.din(w_dff_A_1t47kqJw6_1),.clk(gclk));
	jdff dff_A_RVQRq0Pq2_1(.dout(w_dff_A_1t47kqJw6_1),.din(w_dff_A_RVQRq0Pq2_1),.clk(gclk));
	jdff dff_A_Pog6FL2u0_2(.dout(w_G169_1[2]),.din(w_dff_A_Pog6FL2u0_2),.clk(gclk));
	jdff dff_A_VILqyT0n7_2(.dout(w_dff_A_Pog6FL2u0_2),.din(w_dff_A_VILqyT0n7_2),.clk(gclk));
	jdff dff_A_KDRBfgLl1_2(.dout(w_dff_A_VILqyT0n7_2),.din(w_dff_A_KDRBfgLl1_2),.clk(gclk));
	jdff dff_A_3tiSyFd27_2(.dout(w_dff_A_KDRBfgLl1_2),.din(w_dff_A_3tiSyFd27_2),.clk(gclk));
	jdff dff_A_DIw65otO6_2(.dout(w_dff_A_3tiSyFd27_2),.din(w_dff_A_DIw65otO6_2),.clk(gclk));
	jdff dff_A_74qqsdmk8_2(.dout(w_dff_A_DIw65otO6_2),.din(w_dff_A_74qqsdmk8_2),.clk(gclk));
	jdff dff_A_BKSTxEcr2_2(.dout(w_dff_A_74qqsdmk8_2),.din(w_dff_A_BKSTxEcr2_2),.clk(gclk));
	jdff dff_A_3krxqJlc2_2(.dout(w_dff_A_BKSTxEcr2_2),.din(w_dff_A_3krxqJlc2_2),.clk(gclk));
	jdff dff_A_aVbwgv255_1(.dout(w_n151_4[1]),.din(w_dff_A_aVbwgv255_1),.clk(gclk));
	jdff dff_A_gKi8yo9w2_1(.dout(w_dff_A_aVbwgv255_1),.din(w_dff_A_gKi8yo9w2_1),.clk(gclk));
	jdff dff_A_fGufZ8pH1_1(.dout(w_dff_A_gKi8yo9w2_1),.din(w_dff_A_fGufZ8pH1_1),.clk(gclk));
	jdff dff_B_Yr1JPm3o5_0(.din(n676),.dout(w_dff_B_Yr1JPm3o5_0),.clk(gclk));
	jdff dff_B_ICvUMYKM8_0(.din(w_dff_B_Yr1JPm3o5_0),.dout(w_dff_B_ICvUMYKM8_0),.clk(gclk));
	jdff dff_B_BFrZPIXe7_1(.din(n661),.dout(w_dff_B_BFrZPIXe7_1),.clk(gclk));
	jdff dff_B_RP6BSa9O4_1(.din(w_dff_B_BFrZPIXe7_1),.dout(w_dff_B_RP6BSa9O4_1),.clk(gclk));
	jdff dff_B_HHMlweB50_1(.din(w_dff_B_RP6BSa9O4_1),.dout(w_dff_B_HHMlweB50_1),.clk(gclk));
	jdff dff_B_vPFDHvJh1_1(.din(w_dff_B_HHMlweB50_1),.dout(w_dff_B_vPFDHvJh1_1),.clk(gclk));
	jdff dff_B_fjFwbOIT9_0(.din(n672),.dout(w_dff_B_fjFwbOIT9_0),.clk(gclk));
	jdff dff_A_FScjjiaP9_0(.dout(w_G317_1[0]),.din(w_dff_A_FScjjiaP9_0),.clk(gclk));
	jdff dff_B_kxpliCxs7_3(.din(G317),.dout(w_dff_B_kxpliCxs7_3),.clk(gclk));
	jdff dff_B_ANkkWsD70_3(.din(w_dff_B_kxpliCxs7_3),.dout(w_dff_B_ANkkWsD70_3),.clk(gclk));
	jdff dff_B_lCwqRcNN5_3(.din(w_dff_B_ANkkWsD70_3),.dout(w_dff_B_lCwqRcNN5_3),.clk(gclk));
	jdff dff_A_uHrmcmKh9_1(.dout(w_G311_1[1]),.din(w_dff_A_uHrmcmKh9_1),.clk(gclk));
	jdff dff_B_iemHjl6C8_3(.din(G311),.dout(w_dff_B_iemHjl6C8_3),.clk(gclk));
	jdff dff_B_ZpoKtMzY1_3(.din(w_dff_B_iemHjl6C8_3),.dout(w_dff_B_ZpoKtMzY1_3),.clk(gclk));
	jdff dff_B_WJf49pZb6_3(.din(w_dff_B_ZpoKtMzY1_3),.dout(w_dff_B_WJf49pZb6_3),.clk(gclk));
	jdff dff_B_6hP6nKcU1_1(.din(G329),.dout(w_dff_B_6hP6nKcU1_1),.clk(gclk));
	jdff dff_B_BHujTII25_1(.din(w_dff_B_6hP6nKcU1_1),.dout(w_dff_B_BHujTII25_1),.clk(gclk));
	jdff dff_B_5q32YLO21_1(.din(w_dff_B_BHujTII25_1),.dout(w_dff_B_5q32YLO21_1),.clk(gclk));
	jdff dff_B_X2gvFluv2_1(.din(w_dff_B_5q32YLO21_1),.dout(w_dff_B_X2gvFluv2_1),.clk(gclk));
	jdff dff_B_J2PbBJUE9_0(.din(n665),.dout(w_dff_B_J2PbBJUE9_0),.clk(gclk));
	jdff dff_B_4OPNyqaq3_0(.din(w_dff_B_J2PbBJUE9_0),.dout(w_dff_B_4OPNyqaq3_0),.clk(gclk));
	jdff dff_A_3oePydcL6_0(.dout(w_G326_0[0]),.din(w_dff_A_3oePydcL6_0),.clk(gclk));
	jdff dff_B_I8F6JcTl3_2(.din(G326),.dout(w_dff_B_I8F6JcTl3_2),.clk(gclk));
	jdff dff_B_UgFMn3Bk1_2(.din(w_dff_B_I8F6JcTl3_2),.dout(w_dff_B_UgFMn3Bk1_2),.clk(gclk));
	jdff dff_B_lMmWfDJV8_2(.din(w_dff_B_UgFMn3Bk1_2),.dout(w_dff_B_lMmWfDJV8_2),.clk(gclk));
	jdff dff_B_yj2II1H15_1(.din(n662),.dout(w_dff_B_yj2II1H15_1),.clk(gclk));
	jdff dff_A_7ieWbLck8_0(.dout(w_G294_3[0]),.din(w_dff_A_7ieWbLck8_0),.clk(gclk));
	jdff dff_A_zCo5Gg825_0(.dout(w_dff_A_7ieWbLck8_0),.din(w_dff_A_zCo5Gg825_0),.clk(gclk));
	jdff dff_A_cnxeaZtt8_0(.dout(w_dff_A_zCo5Gg825_0),.din(w_dff_A_cnxeaZtt8_0),.clk(gclk));
	jdff dff_A_OzvO7sgZ4_0(.dout(w_dff_A_cnxeaZtt8_0),.din(w_dff_A_OzvO7sgZ4_0),.clk(gclk));
	jdff dff_A_4gnjVid50_0(.dout(w_G294_0[0]),.din(w_dff_A_4gnjVid50_0),.clk(gclk));
	jdff dff_A_NmBoDBTE5_0(.dout(w_dff_A_4gnjVid50_0),.din(w_dff_A_NmBoDBTE5_0),.clk(gclk));
	jdff dff_A_mOudWFRR2_0(.dout(w_dff_A_NmBoDBTE5_0),.din(w_dff_A_mOudWFRR2_0),.clk(gclk));
	jdff dff_A_52VXOKlF3_1(.dout(w_G294_0[1]),.din(w_dff_A_52VXOKlF3_1),.clk(gclk));
	jdff dff_A_NbmQmMQd6_1(.dout(w_dff_A_52VXOKlF3_1),.din(w_dff_A_NbmQmMQd6_1),.clk(gclk));
	jdff dff_A_ighade174_1(.dout(w_dff_A_NbmQmMQd6_1),.din(w_dff_A_ighade174_1),.clk(gclk));
	jdff dff_A_eumKDIYD0_0(.dout(w_G322_0[0]),.din(w_dff_A_eumKDIYD0_0),.clk(gclk));
	jdff dff_B_27uRssiL8_3(.din(G322),.dout(w_dff_B_27uRssiL8_3),.clk(gclk));
	jdff dff_B_EjMYS9bm4_3(.din(w_dff_B_27uRssiL8_3),.dout(w_dff_B_EjMYS9bm4_3),.clk(gclk));
	jdff dff_B_SsOHuoV00_3(.din(w_dff_B_EjMYS9bm4_3),.dout(w_dff_B_SsOHuoV00_3),.clk(gclk));
	jdff dff_B_myZ2XzXV4_0(.din(n658),.dout(w_dff_B_myZ2XzXV4_0),.clk(gclk));
	jdff dff_B_mqqainCH2_1(.din(n647),.dout(w_dff_B_mqqainCH2_1),.clk(gclk));
	jdff dff_B_PnhJcXFb8_1(.din(w_dff_B_mqqainCH2_1),.dout(w_dff_B_PnhJcXFb8_1),.clk(gclk));
	jdff dff_A_70XTfknm0_1(.dout(w_G68_3[1]),.din(w_dff_A_70XTfknm0_1),.clk(gclk));
	jdff dff_A_toJ0YaT87_1(.dout(w_dff_A_70XTfknm0_1),.din(w_dff_A_toJ0YaT87_1),.clk(gclk));
	jdff dff_A_zlDsV8Ur1_2(.dout(w_G68_3[2]),.din(w_dff_A_zlDsV8Ur1_2),.clk(gclk));
	jdff dff_A_5JEDc2PT9_2(.dout(w_dff_A_zlDsV8Ur1_2),.din(w_dff_A_5JEDc2PT9_2),.clk(gclk));
	jdff dff_A_MoPl1Dqo0_2(.dout(w_G68_0[2]),.din(w_dff_A_MoPl1Dqo0_2),.clk(gclk));
	jdff dff_A_lRzML6Mb2_0(.dout(w_G50_4[0]),.din(w_dff_A_lRzML6Mb2_0),.clk(gclk));
	jdff dff_A_mmRpLKz87_0(.dout(w_dff_A_lRzML6Mb2_0),.din(w_dff_A_mmRpLKz87_0),.clk(gclk));
	jdff dff_A_RbkvkLIx2_1(.dout(w_G50_4[1]),.din(w_dff_A_RbkvkLIx2_1),.clk(gclk));
	jdff dff_A_3CWmlWEH5_1(.dout(w_dff_A_RbkvkLIx2_1),.din(w_dff_A_3CWmlWEH5_1),.clk(gclk));
	jdff dff_A_X3FU8xLS8_0(.dout(w_G50_1[0]),.din(w_dff_A_X3FU8xLS8_0),.clk(gclk));
	jdff dff_A_8LbIGvRR0_2(.dout(w_G50_1[2]),.din(w_dff_A_8LbIGvRR0_2),.clk(gclk));
	jdff dff_A_j2vEdCQF4_2(.dout(w_dff_A_8LbIGvRR0_2),.din(w_dff_A_j2vEdCQF4_2),.clk(gclk));
	jdff dff_A_5I8oE4Ae9_2(.dout(w_dff_A_j2vEdCQF4_2),.din(w_dff_A_5I8oE4Ae9_2),.clk(gclk));
	jdff dff_A_hpXedVji2_2(.dout(w_dff_A_5I8oE4Ae9_2),.din(w_dff_A_hpXedVji2_2),.clk(gclk));
	jdff dff_A_Hd7FvtnU2_1(.dout(w_n649_0[1]),.din(w_dff_A_Hd7FvtnU2_1),.clk(gclk));
	jdff dff_A_SI4ahCmL4_0(.dout(w_G107_3[0]),.din(w_dff_A_SI4ahCmL4_0),.clk(gclk));
	jdff dff_A_g8wPMPOg8_0(.dout(w_dff_A_SI4ahCmL4_0),.din(w_dff_A_g8wPMPOg8_0),.clk(gclk));
	jdff dff_A_BBf4G9ah5_0(.dout(w_dff_A_g8wPMPOg8_0),.din(w_dff_A_BBf4G9ah5_0),.clk(gclk));
	jdff dff_A_lz046jDm0_1(.dout(w_G107_0[1]),.din(w_dff_A_lz046jDm0_1),.clk(gclk));
	jdff dff_A_tGrfnBzK0_1(.dout(w_dff_A_lz046jDm0_1),.din(w_dff_A_tGrfnBzK0_1),.clk(gclk));
	jdff dff_A_pPVzhuRw2_1(.dout(w_dff_A_tGrfnBzK0_1),.din(w_dff_A_pPVzhuRw2_1),.clk(gclk));
	jdff dff_A_lpyZ4Tfq1_0(.dout(w_G58_4[0]),.din(w_dff_A_lpyZ4Tfq1_0),.clk(gclk));
	jdff dff_A_v4KsQ1He7_0(.dout(w_dff_A_lpyZ4Tfq1_0),.din(w_dff_A_v4KsQ1He7_0),.clk(gclk));
	jdff dff_A_uVJ5F7Xq3_0(.dout(w_dff_A_v4KsQ1He7_0),.din(w_dff_A_uVJ5F7Xq3_0),.clk(gclk));
	jdff dff_A_L4WK5rxH3_2(.dout(w_G58_4[2]),.din(w_dff_A_L4WK5rxH3_2),.clk(gclk));
	jdff dff_A_vIZPcx7T9_2(.dout(w_dff_A_L4WK5rxH3_2),.din(w_dff_A_vIZPcx7T9_2),.clk(gclk));
	jdff dff_A_FnySFvXJ1_2(.dout(w_G58_1[2]),.din(w_dff_A_FnySFvXJ1_2),.clk(gclk));
	jdff dff_A_FLFFGcne8_2(.dout(w_dff_A_FnySFvXJ1_2),.din(w_dff_A_FLFFGcne8_2),.clk(gclk));
	jdff dff_A_9njr8Asa5_2(.dout(w_dff_A_FLFFGcne8_2),.din(w_dff_A_9njr8Asa5_2),.clk(gclk));
	jdff dff_A_4sD7ZGpF7_1(.dout(w_G58_0[1]),.din(w_dff_A_4sD7ZGpF7_1),.clk(gclk));
	jdff dff_B_X7YjN2rJ7_1(.din(n636),.dout(w_dff_B_X7YjN2rJ7_1),.clk(gclk));
	jdff dff_B_gCWrTEup1_1(.din(n639),.dout(w_dff_B_gCWrTEup1_1),.clk(gclk));
	jdff dff_A_Yzeoj65M9_0(.dout(w_G159_3[0]),.din(w_dff_A_Yzeoj65M9_0),.clk(gclk));
	jdff dff_A_DHqjW4NS9_0(.dout(w_dff_A_Yzeoj65M9_0),.din(w_dff_A_DHqjW4NS9_0),.clk(gclk));
	jdff dff_A_F3hCORgC0_0(.dout(w_dff_A_DHqjW4NS9_0),.din(w_dff_A_F3hCORgC0_0),.clk(gclk));
	jdff dff_A_8PNDLNEK5_1(.dout(w_G159_3[1]),.din(w_dff_A_8PNDLNEK5_1),.clk(gclk));
	jdff dff_A_bQxUdfq12_1(.dout(w_dff_A_8PNDLNEK5_1),.din(w_dff_A_bQxUdfq12_1),.clk(gclk));
	jdff dff_A_nVvevhsn6_1(.dout(w_dff_A_bQxUdfq12_1),.din(w_dff_A_nVvevhsn6_1),.clk(gclk));
	jdff dff_A_oXxWy2579_1(.dout(w_dff_A_nVvevhsn6_1),.din(w_dff_A_oXxWy2579_1),.clk(gclk));
	jdff dff_A_8723l0Ow7_0(.dout(w_G159_0[0]),.din(w_dff_A_8723l0Ow7_0),.clk(gclk));
	jdff dff_A_YXvWWlFI9_0(.dout(w_dff_A_8723l0Ow7_0),.din(w_dff_A_YXvWWlFI9_0),.clk(gclk));
	jdff dff_A_HlTdhWGI7_0(.dout(w_dff_A_YXvWWlFI9_0),.din(w_dff_A_HlTdhWGI7_0),.clk(gclk));
	jdff dff_A_c5YuD6Qa7_1(.dout(w_G159_0[1]),.din(w_dff_A_c5YuD6Qa7_1),.clk(gclk));
	jdff dff_A_bCRGNL845_1(.dout(w_dff_A_c5YuD6Qa7_1),.din(w_dff_A_bCRGNL845_1),.clk(gclk));
	jdff dff_A_icJRTxbs6_1(.dout(w_dff_A_bCRGNL845_1),.din(w_dff_A_icJRTxbs6_1),.clk(gclk));
	jdff dff_A_bgXHxdSP6_0(.dout(w_n388_0[0]),.din(w_dff_A_bgXHxdSP6_0),.clk(gclk));
	jdff dff_A_ZPhdqEDj4_0(.dout(w_dff_A_bgXHxdSP6_0),.din(w_dff_A_ZPhdqEDj4_0),.clk(gclk));
	jdff dff_A_YY8hlWwA5_0(.dout(w_dff_A_ZPhdqEDj4_0),.din(w_dff_A_YY8hlWwA5_0),.clk(gclk));
	jdff dff_A_Rc1R6jDI9_0(.dout(w_dff_A_YY8hlWwA5_0),.din(w_dff_A_Rc1R6jDI9_0),.clk(gclk));
	jdff dff_A_oo5FkNuM5_0(.dout(w_dff_A_Rc1R6jDI9_0),.din(w_dff_A_oo5FkNuM5_0),.clk(gclk));
	jdff dff_A_ivs22P1q2_0(.dout(w_dff_A_oo5FkNuM5_0),.din(w_dff_A_ivs22P1q2_0),.clk(gclk));
	jdff dff_A_BJRX0yQT4_1(.dout(w_n388_0[1]),.din(w_dff_A_BJRX0yQT4_1),.clk(gclk));
	jdff dff_A_kNhp2yBW2_1(.dout(w_dff_A_BJRX0yQT4_1),.din(w_dff_A_kNhp2yBW2_1),.clk(gclk));
	jdff dff_A_712ULcCv3_1(.dout(w_dff_A_kNhp2yBW2_1),.din(w_dff_A_712ULcCv3_1),.clk(gclk));
	jdff dff_A_sdSmB09l4_1(.dout(w_dff_A_712ULcCv3_1),.din(w_dff_A_sdSmB09l4_1),.clk(gclk));
	jdff dff_A_mbAwSa6M3_1(.dout(w_dff_A_sdSmB09l4_1),.din(w_dff_A_mbAwSa6M3_1),.clk(gclk));
	jdff dff_A_FaeAKi4W3_1(.dout(w_dff_A_mbAwSa6M3_1),.din(w_dff_A_FaeAKi4W3_1),.clk(gclk));
	jdff dff_A_GaxknGMP0_1(.dout(w_dff_A_FaeAKi4W3_1),.din(w_dff_A_GaxknGMP0_1),.clk(gclk));
	jdff dff_A_mQ3qDXyH4_1(.dout(w_G200_2[1]),.din(w_dff_A_mQ3qDXyH4_1),.clk(gclk));
	jdff dff_A_yWfi02f91_1(.dout(w_dff_A_mQ3qDXyH4_1),.din(w_dff_A_yWfi02f91_1),.clk(gclk));
	jdff dff_A_TaJ9Tvf54_1(.dout(w_dff_A_yWfi02f91_1),.din(w_dff_A_TaJ9Tvf54_1),.clk(gclk));
	jdff dff_A_ri80zXZg9_1(.dout(w_dff_A_TaJ9Tvf54_1),.din(w_dff_A_ri80zXZg9_1),.clk(gclk));
	jdff dff_A_HYv2t2Sc3_1(.dout(w_dff_A_ri80zXZg9_1),.din(w_dff_A_HYv2t2Sc3_1),.clk(gclk));
	jdff dff_A_Sg9pd1EJ4_1(.dout(w_dff_A_HYv2t2Sc3_1),.din(w_dff_A_Sg9pd1EJ4_1),.clk(gclk));
	jdff dff_A_8Wqz2aeg8_1(.dout(w_dff_A_Sg9pd1EJ4_1),.din(w_dff_A_8Wqz2aeg8_1),.clk(gclk));
	jdff dff_A_5fvJvEOG9_1(.dout(w_dff_A_8Wqz2aeg8_1),.din(w_dff_A_5fvJvEOG9_1),.clk(gclk));
	jdff dff_A_muz11URF6_2(.dout(w_G200_2[2]),.din(w_dff_A_muz11URF6_2),.clk(gclk));
	jdff dff_A_YCDcsEIS3_2(.dout(w_dff_A_muz11URF6_2),.din(w_dff_A_YCDcsEIS3_2),.clk(gclk));
	jdff dff_A_KrU73EEJ6_2(.dout(w_dff_A_YCDcsEIS3_2),.din(w_dff_A_KrU73EEJ6_2),.clk(gclk));
	jdff dff_A_pZOaYuK99_2(.dout(w_dff_A_KrU73EEJ6_2),.din(w_dff_A_pZOaYuK99_2),.clk(gclk));
	jdff dff_A_ZID46GEC5_2(.dout(w_dff_A_pZOaYuK99_2),.din(w_dff_A_ZID46GEC5_2),.clk(gclk));
	jdff dff_A_Bts8WQCO4_2(.dout(w_dff_A_ZID46GEC5_2),.din(w_dff_A_Bts8WQCO4_2),.clk(gclk));
	jdff dff_A_KRBhaKoL6_2(.dout(w_dff_A_Bts8WQCO4_2),.din(w_dff_A_KRBhaKoL6_2),.clk(gclk));
	jdff dff_A_bcvv62SF1_0(.dout(w_G77_3[0]),.din(w_dff_A_bcvv62SF1_0),.clk(gclk));
	jdff dff_A_erMOcKIW6_0(.dout(w_dff_A_bcvv62SF1_0),.din(w_dff_A_erMOcKIW6_0),.clk(gclk));
	jdff dff_A_XdFUXiYj2_0(.dout(w_dff_A_erMOcKIW6_0),.din(w_dff_A_XdFUXiYj2_0),.clk(gclk));
	jdff dff_A_4FcJkg507_2(.dout(w_G77_3[2]),.din(w_dff_A_4FcJkg507_2),.clk(gclk));
	jdff dff_A_IIdbkcLz0_2(.dout(w_dff_A_4FcJkg507_2),.din(w_dff_A_IIdbkcLz0_2),.clk(gclk));
	jdff dff_A_SSQAyeQo5_2(.dout(w_dff_A_IIdbkcLz0_2),.din(w_dff_A_SSQAyeQo5_2),.clk(gclk));
	jdff dff_A_14rTpuBW4_1(.dout(w_G77_0[1]),.din(w_dff_A_14rTpuBW4_1),.clk(gclk));
	jdff dff_A_vDc3UwJq2_1(.dout(w_dff_A_14rTpuBW4_1),.din(w_dff_A_vDc3UwJq2_1),.clk(gclk));
	jdff dff_A_fMqTtTDq2_0(.dout(w_G33_7[0]),.din(w_dff_A_fMqTtTDq2_0),.clk(gclk));
	jdff dff_A_MQ4TaRnf0_0(.dout(w_dff_A_fMqTtTDq2_0),.din(w_dff_A_MQ4TaRnf0_0),.clk(gclk));
	jdff dff_A_astzEWJ06_0(.dout(w_dff_A_MQ4TaRnf0_0),.din(w_dff_A_astzEWJ06_0),.clk(gclk));
	jdff dff_A_qGb9CV3y4_0(.dout(w_dff_A_astzEWJ06_0),.din(w_dff_A_qGb9CV3y4_0),.clk(gclk));
	jdff dff_A_m3yRD9YY2_0(.dout(w_dff_A_qGb9CV3y4_0),.din(w_dff_A_m3yRD9YY2_0),.clk(gclk));
	jdff dff_A_C9Ok3oI29_0(.dout(w_dff_A_m3yRD9YY2_0),.din(w_dff_A_C9Ok3oI29_0),.clk(gclk));
	jdff dff_A_Ilws0PQQ1_1(.dout(w_G33_7[1]),.din(w_dff_A_Ilws0PQQ1_1),.clk(gclk));
	jdff dff_B_kt5ToKu03_0(.din(n635),.dout(w_dff_B_kt5ToKu03_0),.clk(gclk));
	jdff dff_A_9AWUBrYy9_0(.dout(w_G87_2[0]),.din(w_dff_A_9AWUBrYy9_0),.clk(gclk));
	jdff dff_A_us1sAlX99_0(.dout(w_dff_A_9AWUBrYy9_0),.din(w_dff_A_us1sAlX99_0),.clk(gclk));
	jdff dff_A_8KS8086U1_0(.dout(w_dff_A_us1sAlX99_0),.din(w_dff_A_8KS8086U1_0),.clk(gclk));
	jdff dff_A_hgsEczfJ6_1(.dout(w_G87_2[1]),.din(w_dff_A_hgsEczfJ6_1),.clk(gclk));
	jdff dff_A_9IFLZ5XQ2_1(.dout(w_dff_A_hgsEczfJ6_1),.din(w_dff_A_9IFLZ5XQ2_1),.clk(gclk));
	jdff dff_A_Z5pizf2f2_1(.dout(w_dff_A_9IFLZ5XQ2_1),.din(w_dff_A_Z5pizf2f2_1),.clk(gclk));
	jdff dff_A_lO8NRHu24_0(.dout(w_G87_0[0]),.din(w_dff_A_lO8NRHu24_0),.clk(gclk));
	jdff dff_A_P4E7cyLt3_0(.dout(w_dff_A_lO8NRHu24_0),.din(w_dff_A_P4E7cyLt3_0),.clk(gclk));
	jdff dff_A_MFLTO2Ch3_0(.dout(w_dff_A_P4E7cyLt3_0),.din(w_dff_A_MFLTO2Ch3_0),.clk(gclk));
	jdff dff_A_JtIPGaNL4_0(.dout(w_G200_1[0]),.din(w_dff_A_JtIPGaNL4_0),.clk(gclk));
	jdff dff_A_f3OZvj1Y3_2(.dout(w_G200_1[2]),.din(w_dff_A_f3OZvj1Y3_2),.clk(gclk));
	jdff dff_A_kXDMht8p9_2(.dout(w_dff_A_f3OZvj1Y3_2),.din(w_dff_A_kXDMht8p9_2),.clk(gclk));
	jdff dff_A_VHghzJcb7_2(.dout(w_dff_A_kXDMht8p9_2),.din(w_dff_A_VHghzJcb7_2),.clk(gclk));
	jdff dff_A_2aXEwhUq6_2(.dout(w_dff_A_VHghzJcb7_2),.din(w_dff_A_2aXEwhUq6_2),.clk(gclk));
	jdff dff_A_zMiLK88G4_2(.dout(w_dff_A_2aXEwhUq6_2),.din(w_dff_A_zMiLK88G4_2),.clk(gclk));
	jdff dff_A_7atZrdQS0_2(.dout(w_dff_A_zMiLK88G4_2),.din(w_dff_A_7atZrdQS0_2),.clk(gclk));
	jdff dff_A_J4XvV5vL2_2(.dout(w_dff_A_7atZrdQS0_2),.din(w_dff_A_J4XvV5vL2_2),.clk(gclk));
	jdff dff_A_9DcS5XPD4_2(.dout(w_dff_A_J4XvV5vL2_2),.din(w_dff_A_9DcS5XPD4_2),.clk(gclk));
	jdff dff_A_IGkdb4hj6_0(.dout(w_n622_0[0]),.din(w_dff_A_IGkdb4hj6_0),.clk(gclk));
	jdff dff_A_LNiO5wDO0_0(.dout(w_n507_1[0]),.din(w_dff_A_LNiO5wDO0_0),.clk(gclk));
	jdff dff_A_dBe52Yhh4_1(.dout(w_n507_1[1]),.din(w_dff_A_dBe52Yhh4_1),.clk(gclk));
	jdff dff_A_MnIkuD4d6_1(.dout(w_n507_0[1]),.din(w_dff_A_MnIkuD4d6_1),.clk(gclk));
	jdff dff_A_tGd31CWb0_1(.dout(w_dff_A_MnIkuD4d6_1),.din(w_dff_A_tGd31CWb0_1),.clk(gclk));
	jdff dff_A_xWlsNxxd9_1(.dout(w_dff_A_tGd31CWb0_1),.din(w_dff_A_xWlsNxxd9_1),.clk(gclk));
	jdff dff_A_xvzK95Pw1_1(.dout(w_dff_A_xWlsNxxd9_1),.din(w_dff_A_xvzK95Pw1_1),.clk(gclk));
	jdff dff_A_dYMqDWDe6_1(.dout(w_dff_A_xvzK95Pw1_1),.din(w_dff_A_dYMqDWDe6_1),.clk(gclk));
	jdff dff_A_M1oOOEom0_1(.dout(w_dff_A_dYMqDWDe6_1),.din(w_dff_A_M1oOOEom0_1),.clk(gclk));
	jdff dff_A_Sy4bVevd0_2(.dout(w_n507_0[2]),.din(w_dff_A_Sy4bVevd0_2),.clk(gclk));
	jdff dff_A_iHds2Ppo4_0(.dout(w_G190_2[0]),.din(w_dff_A_iHds2Ppo4_0),.clk(gclk));
	jdff dff_A_JQqvRTx24_0(.dout(w_dff_A_iHds2Ppo4_0),.din(w_dff_A_JQqvRTx24_0),.clk(gclk));
	jdff dff_A_ruYeLqrG0_2(.dout(w_G190_2[2]),.din(w_dff_A_ruYeLqrG0_2),.clk(gclk));
	jdff dff_A_mLE1O6VH1_2(.dout(w_dff_A_ruYeLqrG0_2),.din(w_dff_A_mLE1O6VH1_2),.clk(gclk));
	jdff dff_A_ZQEm9SnP6_2(.dout(w_dff_A_mLE1O6VH1_2),.din(w_dff_A_ZQEm9SnP6_2),.clk(gclk));
	jdff dff_A_ejOX0Npw7_2(.dout(w_dff_A_ZQEm9SnP6_2),.din(w_dff_A_ejOX0Npw7_2),.clk(gclk));
	jdff dff_A_h7pu5H8W1_2(.dout(w_dff_A_ejOX0Npw7_2),.din(w_dff_A_h7pu5H8W1_2),.clk(gclk));
	jdff dff_A_pSgOUg0m4_2(.dout(w_dff_A_h7pu5H8W1_2),.din(w_dff_A_pSgOUg0m4_2),.clk(gclk));
	jdff dff_A_yr7TgXcb7_2(.dout(w_dff_A_pSgOUg0m4_2),.din(w_dff_A_yr7TgXcb7_2),.clk(gclk));
	jdff dff_A_5eVJVE8F5_2(.dout(w_dff_A_yr7TgXcb7_2),.din(w_dff_A_5eVJVE8F5_2),.clk(gclk));
	jdff dff_A_kYWp7nK21_2(.dout(w_G20_2[2]),.din(w_dff_A_kYWp7nK21_2),.clk(gclk));
	jdff dff_A_vloAHOvc1_0(.dout(w_G97_3[0]),.din(w_dff_A_vloAHOvc1_0),.clk(gclk));
	jdff dff_A_fE8K8uMx9_0(.dout(w_dff_A_vloAHOvc1_0),.din(w_dff_A_fE8K8uMx9_0),.clk(gclk));
	jdff dff_A_5H7DAu1C4_0(.dout(w_dff_A_fE8K8uMx9_0),.din(w_dff_A_5H7DAu1C4_0),.clk(gclk));
	jdff dff_A_4Ryte8mL2_0(.dout(w_dff_A_5H7DAu1C4_0),.din(w_dff_A_4Ryte8mL2_0),.clk(gclk));
	jdff dff_A_xDLcMC0L3_0(.dout(w_n620_0[0]),.din(w_dff_A_xDLcMC0L3_0),.clk(gclk));
	jdff dff_A_tl2aQEaD1_0(.dout(w_dff_A_xDLcMC0L3_0),.din(w_dff_A_tl2aQEaD1_0),.clk(gclk));
	jdff dff_A_mVzC57TR9_0(.dout(w_dff_A_tl2aQEaD1_0),.din(w_dff_A_mVzC57TR9_0),.clk(gclk));
	jdff dff_A_F0l7AFWz3_0(.dout(w_dff_A_mVzC57TR9_0),.din(w_dff_A_F0l7AFWz3_0),.clk(gclk));
	jdff dff_A_PBbAEb990_0(.dout(w_dff_A_F0l7AFWz3_0),.din(w_dff_A_PBbAEb990_0),.clk(gclk));
	jdff dff_A_SeG4EnS90_0(.dout(w_dff_A_PBbAEb990_0),.din(w_dff_A_SeG4EnS90_0),.clk(gclk));
	jdff dff_A_ElGLvhAj1_0(.dout(w_dff_A_SeG4EnS90_0),.din(w_dff_A_ElGLvhAj1_0),.clk(gclk));
	jdff dff_A_5EPsDdxo5_0(.dout(w_dff_A_ElGLvhAj1_0),.din(w_dff_A_5EPsDdxo5_0),.clk(gclk));
	jdff dff_A_LxUlK06f0_0(.dout(w_dff_A_5EPsDdxo5_0),.din(w_dff_A_LxUlK06f0_0),.clk(gclk));
	jdff dff_A_lCzPaocn8_2(.dout(w_n620_0[2]),.din(w_dff_A_lCzPaocn8_2),.clk(gclk));
	jdff dff_A_iueAX1qg8_2(.dout(w_dff_A_lCzPaocn8_2),.din(w_dff_A_iueAX1qg8_2),.clk(gclk));
	jdff dff_A_Zu6j4K7T0_2(.dout(w_dff_A_iueAX1qg8_2),.din(w_dff_A_Zu6j4K7T0_2),.clk(gclk));
	jdff dff_A_3Kmfi5V94_2(.dout(w_dff_A_Zu6j4K7T0_2),.din(w_dff_A_3Kmfi5V94_2),.clk(gclk));
	jdff dff_A_BJcyh7Br9_2(.dout(w_dff_A_3Kmfi5V94_2),.din(w_dff_A_BJcyh7Br9_2),.clk(gclk));
	jdff dff_A_UPbk3OGX8_2(.dout(w_dff_A_BJcyh7Br9_2),.din(w_dff_A_UPbk3OGX8_2),.clk(gclk));
	jdff dff_A_KdhLW2a17_2(.dout(w_dff_A_UPbk3OGX8_2),.din(w_dff_A_KdhLW2a17_2),.clk(gclk));
	jdff dff_A_YMrjh7iP6_2(.dout(w_dff_A_KdhLW2a17_2),.din(w_dff_A_YMrjh7iP6_2),.clk(gclk));
	jdff dff_A_M2eNuPQZ2_2(.dout(w_dff_A_YMrjh7iP6_2),.din(w_dff_A_M2eNuPQZ2_2),.clk(gclk));
	jdff dff_A_9HYA86y12_2(.dout(w_dff_A_M2eNuPQZ2_2),.din(w_dff_A_9HYA86y12_2),.clk(gclk));
	jdff dff_A_NMyEOfkP3_0(.dout(w_n619_0[0]),.din(w_dff_A_NMyEOfkP3_0),.clk(gclk));
	jdff dff_A_sBDXXBtF8_0(.dout(w_dff_A_NMyEOfkP3_0),.din(w_dff_A_sBDXXBtF8_0),.clk(gclk));
	jdff dff_A_92Ak7KAc8_0(.dout(w_dff_A_sBDXXBtF8_0),.din(w_dff_A_92Ak7KAc8_0),.clk(gclk));
	jdff dff_A_7g01XhgD9_0(.dout(w_dff_A_92Ak7KAc8_0),.din(w_dff_A_7g01XhgD9_0),.clk(gclk));
	jdff dff_A_zzmjPlyV1_0(.dout(w_dff_A_7g01XhgD9_0),.din(w_dff_A_zzmjPlyV1_0),.clk(gclk));
	jdff dff_A_QrKTtc2A1_0(.dout(w_dff_A_zzmjPlyV1_0),.din(w_dff_A_QrKTtc2A1_0),.clk(gclk));
	jdff dff_A_tiFSzDKt6_0(.dout(w_dff_A_QrKTtc2A1_0),.din(w_dff_A_tiFSzDKt6_0),.clk(gclk));
	jdff dff_A_2ls2bfCR5_0(.dout(w_dff_A_tiFSzDKt6_0),.din(w_dff_A_2ls2bfCR5_0),.clk(gclk));
	jdff dff_A_qzftM5jx2_0(.dout(w_dff_A_2ls2bfCR5_0),.din(w_dff_A_qzftM5jx2_0),.clk(gclk));
	jdff dff_A_kItzOBoR2_0(.dout(w_dff_A_qzftM5jx2_0),.din(w_dff_A_kItzOBoR2_0),.clk(gclk));
	jdff dff_A_PftzUIhx2_1(.dout(w_n619_0[1]),.din(w_dff_A_PftzUIhx2_1),.clk(gclk));
	jdff dff_A_Ciucv7ih8_1(.dout(w_dff_A_PftzUIhx2_1),.din(w_dff_A_Ciucv7ih8_1),.clk(gclk));
	jdff dff_A_uxKwg3TH2_1(.dout(w_dff_A_Ciucv7ih8_1),.din(w_dff_A_uxKwg3TH2_1),.clk(gclk));
	jdff dff_A_7Y8Bwgiw5_1(.dout(w_dff_A_uxKwg3TH2_1),.din(w_dff_A_7Y8Bwgiw5_1),.clk(gclk));
	jdff dff_A_XrQnTngF8_1(.dout(w_dff_A_7Y8Bwgiw5_1),.din(w_dff_A_XrQnTngF8_1),.clk(gclk));
	jdff dff_A_2z9xH6HH0_1(.dout(w_dff_A_XrQnTngF8_1),.din(w_dff_A_2z9xH6HH0_1),.clk(gclk));
	jdff dff_A_HS47RF610_1(.dout(w_dff_A_2z9xH6HH0_1),.din(w_dff_A_HS47RF610_1),.clk(gclk));
	jdff dff_A_xbD5Qbtu0_1(.dout(w_dff_A_HS47RF610_1),.din(w_dff_A_xbD5Qbtu0_1),.clk(gclk));
	jdff dff_A_N9SE4bwk6_1(.dout(w_dff_A_xbD5Qbtu0_1),.din(w_dff_A_N9SE4bwk6_1),.clk(gclk));
	jdff dff_A_4sqRfDi83_0(.dout(w_n618_2[0]),.din(w_dff_A_4sqRfDi83_0),.clk(gclk));
	jdff dff_A_L7vwNtPl9_0(.dout(w_dff_A_4sqRfDi83_0),.din(w_dff_A_L7vwNtPl9_0),.clk(gclk));
	jdff dff_A_E8HCYfYS5_0(.dout(w_dff_A_L7vwNtPl9_0),.din(w_dff_A_E8HCYfYS5_0),.clk(gclk));
	jdff dff_A_VvPpyrV11_0(.dout(w_dff_A_E8HCYfYS5_0),.din(w_dff_A_VvPpyrV11_0),.clk(gclk));
	jdff dff_A_yOhTKhzB7_0(.dout(w_dff_A_VvPpyrV11_0),.din(w_dff_A_yOhTKhzB7_0),.clk(gclk));
	jdff dff_A_CAtdGYKT0_0(.dout(w_dff_A_yOhTKhzB7_0),.din(w_dff_A_CAtdGYKT0_0),.clk(gclk));
	jdff dff_A_Srq3KN5m2_0(.dout(w_dff_A_CAtdGYKT0_0),.din(w_dff_A_Srq3KN5m2_0),.clk(gclk));
	jdff dff_A_9rBs5DuH8_0(.dout(w_dff_A_Srq3KN5m2_0),.din(w_dff_A_9rBs5DuH8_0),.clk(gclk));
	jdff dff_A_OKjONHKc8_0(.dout(w_dff_A_9rBs5DuH8_0),.din(w_dff_A_OKjONHKc8_0),.clk(gclk));
	jdff dff_A_pzy8VVvM5_0(.dout(w_dff_A_OKjONHKc8_0),.din(w_dff_A_pzy8VVvM5_0),.clk(gclk));
	jdff dff_A_udHnopOJ6_0(.dout(w_dff_A_pzy8VVvM5_0),.din(w_dff_A_udHnopOJ6_0),.clk(gclk));
	jdff dff_A_aDqx3MgK9_0(.dout(w_dff_A_udHnopOJ6_0),.din(w_dff_A_aDqx3MgK9_0),.clk(gclk));
	jdff dff_A_TOm96VmT0_0(.dout(w_dff_A_aDqx3MgK9_0),.din(w_dff_A_TOm96VmT0_0),.clk(gclk));
	jdff dff_A_OYAX7tzg9_2(.dout(w_n618_0[2]),.din(w_dff_A_OYAX7tzg9_2),.clk(gclk));
	jdff dff_A_yhkUkvuk4_2(.dout(w_dff_A_OYAX7tzg9_2),.din(w_dff_A_yhkUkvuk4_2),.clk(gclk));
	jdff dff_A_M7r6AIJo1_2(.dout(w_dff_A_yhkUkvuk4_2),.din(w_dff_A_M7r6AIJo1_2),.clk(gclk));
	jdff dff_A_CWhbu3dK4_2(.dout(w_dff_A_M7r6AIJo1_2),.din(w_dff_A_CWhbu3dK4_2),.clk(gclk));
	jdff dff_A_X0Scy0Mx6_2(.dout(w_dff_A_CWhbu3dK4_2),.din(w_dff_A_X0Scy0Mx6_2),.clk(gclk));
	jdff dff_A_hYjqc3Uq2_2(.dout(w_dff_A_X0Scy0Mx6_2),.din(w_dff_A_hYjqc3Uq2_2),.clk(gclk));
	jdff dff_A_FCCJcO7k9_2(.dout(w_dff_A_hYjqc3Uq2_2),.din(w_dff_A_FCCJcO7k9_2),.clk(gclk));
	jdff dff_A_T0cGMJoL3_2(.dout(w_dff_A_FCCJcO7k9_2),.din(w_dff_A_T0cGMJoL3_2),.clk(gclk));
	jdff dff_A_GQjFCc4r9_2(.dout(w_dff_A_T0cGMJoL3_2),.din(w_dff_A_GQjFCc4r9_2),.clk(gclk));
	jdff dff_A_rKuDsEIW0_2(.dout(w_dff_A_GQjFCc4r9_2),.din(w_dff_A_rKuDsEIW0_2),.clk(gclk));
	jdff dff_A_oAapYwWF8_2(.dout(w_dff_A_rKuDsEIW0_2),.din(w_dff_A_oAapYwWF8_2),.clk(gclk));
	jdff dff_A_leBPYbM77_2(.dout(w_dff_A_oAapYwWF8_2),.din(w_dff_A_leBPYbM77_2),.clk(gclk));
	jdff dff_A_eY5S2s1i4_0(.dout(w_n153_5[0]),.din(w_dff_A_eY5S2s1i4_0),.clk(gclk));
	jdff dff_A_kWQ85yIV8_0(.dout(w_dff_A_eY5S2s1i4_0),.din(w_dff_A_kWQ85yIV8_0),.clk(gclk));
	jdff dff_A_3ZEeqlf08_0(.dout(w_dff_A_kWQ85yIV8_0),.din(w_dff_A_3ZEeqlf08_0),.clk(gclk));
	jdff dff_A_BrvxRotp4_0(.dout(w_dff_A_3ZEeqlf08_0),.din(w_dff_A_BrvxRotp4_0),.clk(gclk));
	jdff dff_A_StcY7TdP4_0(.dout(w_n153_1[0]),.din(w_dff_A_StcY7TdP4_0),.clk(gclk));
	jdff dff_A_vePoAHTu0_0(.dout(w_dff_A_StcY7TdP4_0),.din(w_dff_A_vePoAHTu0_0),.clk(gclk));
	jdff dff_B_p246Exej3_1(.din(n615),.dout(w_dff_B_p246Exej3_1),.clk(gclk));
	jdff dff_B_khDhyt378_1(.din(w_dff_B_p246Exej3_1),.dout(w_dff_B_khDhyt378_1),.clk(gclk));
	jdff dff_B_SoTVFqOj6_1(.din(w_dff_B_khDhyt378_1),.dout(w_dff_B_SoTVFqOj6_1),.clk(gclk));
	jdff dff_B_E42CMBiT4_1(.din(w_dff_B_SoTVFqOj6_1),.dout(w_dff_B_E42CMBiT4_1),.clk(gclk));
	jdff dff_B_QIveM39a7_1(.din(w_dff_B_E42CMBiT4_1),.dout(w_dff_B_QIveM39a7_1),.clk(gclk));
	jdff dff_B_J0G1r0Mf6_1(.din(w_dff_B_QIveM39a7_1),.dout(w_dff_B_J0G1r0Mf6_1),.clk(gclk));
	jdff dff_B_BY8Aebhw8_1(.din(w_dff_B_J0G1r0Mf6_1),.dout(w_dff_B_BY8Aebhw8_1),.clk(gclk));
	jdff dff_B_mecUk3Q59_1(.din(w_dff_B_BY8Aebhw8_1),.dout(w_dff_B_mecUk3Q59_1),.clk(gclk));
	jdff dff_B_oBRmApze4_0(.din(n575),.dout(w_dff_B_oBRmApze4_0),.clk(gclk));
	jdff dff_B_XmTbCIly1_0(.din(w_dff_B_oBRmApze4_0),.dout(w_dff_B_XmTbCIly1_0),.clk(gclk));
	jdff dff_B_KKMEIeZg9_0(.din(w_dff_B_XmTbCIly1_0),.dout(w_dff_B_KKMEIeZg9_0),.clk(gclk));
	jdff dff_B_QAuHnfYV8_0(.din(w_dff_B_KKMEIeZg9_0),.dout(w_dff_B_QAuHnfYV8_0),.clk(gclk));
	jdff dff_A_cBzamRCz6_0(.dout(w_n567_4[0]),.din(w_dff_A_cBzamRCz6_0),.clk(gclk));
	jdff dff_A_KDzKgusz2_0(.dout(w_dff_A_cBzamRCz6_0),.din(w_dff_A_KDzKgusz2_0),.clk(gclk));
	jdff dff_A_p7REkyA23_0(.dout(w_dff_A_KDzKgusz2_0),.din(w_dff_A_p7REkyA23_0),.clk(gclk));
	jdff dff_A_J5JKGTJv5_0(.dout(w_dff_A_p7REkyA23_0),.din(w_dff_A_J5JKGTJv5_0),.clk(gclk));
	jdff dff_A_CCZIbur15_0(.dout(w_dff_A_J5JKGTJv5_0),.din(w_dff_A_CCZIbur15_0),.clk(gclk));
	jdff dff_A_bp3UPr9D4_0(.dout(w_dff_A_CCZIbur15_0),.din(w_dff_A_bp3UPr9D4_0),.clk(gclk));
	jdff dff_A_bgtWyCku0_0(.dout(w_dff_A_bp3UPr9D4_0),.din(w_dff_A_bgtWyCku0_0),.clk(gclk));
	jdff dff_A_Zs0Q64kA6_0(.dout(w_dff_A_bgtWyCku0_0),.din(w_dff_A_Zs0Q64kA6_0),.clk(gclk));
	jdff dff_A_pgQqVXZC5_0(.dout(w_n567_1[0]),.din(w_dff_A_pgQqVXZC5_0),.clk(gclk));
	jdff dff_A_HziYoL3O0_0(.dout(w_dff_A_pgQqVXZC5_0),.din(w_dff_A_HziYoL3O0_0),.clk(gclk));
	jdff dff_A_hLHVdNtW3_0(.dout(w_dff_A_HziYoL3O0_0),.din(w_dff_A_hLHVdNtW3_0),.clk(gclk));
	jdff dff_A_KB4MxrlC1_2(.dout(w_n567_1[2]),.din(w_dff_A_KB4MxrlC1_2),.clk(gclk));
	jdff dff_A_hwYlgUYn7_2(.dout(w_dff_A_KB4MxrlC1_2),.din(w_dff_A_hwYlgUYn7_2),.clk(gclk));
	jdff dff_A_6WZiKHKH9_2(.dout(w_dff_A_hwYlgUYn7_2),.din(w_dff_A_6WZiKHKH9_2),.clk(gclk));
	jdff dff_A_iXmpsiu60_2(.dout(w_dff_A_6WZiKHKH9_2),.din(w_dff_A_iXmpsiu60_2),.clk(gclk));
	jdff dff_A_YnVsCIew1_2(.dout(w_dff_A_iXmpsiu60_2),.din(w_dff_A_YnVsCIew1_2),.clk(gclk));
	jdff dff_A_F3nGzQEX1_2(.dout(w_dff_A_YnVsCIew1_2),.din(w_dff_A_F3nGzQEX1_2),.clk(gclk));
	jdff dff_A_8GIHkBZ16_2(.dout(w_dff_A_F3nGzQEX1_2),.din(w_dff_A_8GIHkBZ16_2),.clk(gclk));
	jdff dff_A_spQo6kNC4_2(.dout(w_dff_A_8GIHkBZ16_2),.din(w_dff_A_spQo6kNC4_2),.clk(gclk));
	jdff dff_A_8dvVbGxP0_2(.dout(w_dff_A_spQo6kNC4_2),.din(w_dff_A_8dvVbGxP0_2),.clk(gclk));
	jdff dff_A_SebHfa9a5_2(.dout(w_dff_A_8dvVbGxP0_2),.din(w_dff_A_SebHfa9a5_2),.clk(gclk));
	jdff dff_A_tz7qKgnZ4_1(.dout(w_n567_0[1]),.din(w_dff_A_tz7qKgnZ4_1),.clk(gclk));
	jdff dff_A_5gHDYrhf4_1(.dout(w_dff_A_tz7qKgnZ4_1),.din(w_dff_A_5gHDYrhf4_1),.clk(gclk));
	jdff dff_A_nulbQinz5_1(.dout(w_dff_A_5gHDYrhf4_1),.din(w_dff_A_nulbQinz5_1),.clk(gclk));
	jdff dff_A_ReHVIFOI4_2(.dout(w_n567_0[2]),.din(w_dff_A_ReHVIFOI4_2),.clk(gclk));
	jdff dff_A_ZmqweskX2_2(.dout(w_dff_A_ReHVIFOI4_2),.din(w_dff_A_ZmqweskX2_2),.clk(gclk));
	jdff dff_A_BQoRkNuz7_1(.dout(w_n566_0[1]),.din(w_dff_A_BQoRkNuz7_1),.clk(gclk));
	jdff dff_A_gna1lane3_1(.dout(w_dff_A_BQoRkNuz7_1),.din(w_dff_A_gna1lane3_1),.clk(gclk));
	jdff dff_A_6HSQCE8g2_1(.dout(w_dff_A_gna1lane3_1),.din(w_dff_A_6HSQCE8g2_1),.clk(gclk));
	jdff dff_A_ACrTOCto7_1(.dout(w_dff_A_6HSQCE8g2_1),.din(w_dff_A_ACrTOCto7_1),.clk(gclk));
	jdff dff_A_SaBZhgma6_1(.dout(w_dff_A_ACrTOCto7_1),.din(w_dff_A_SaBZhgma6_1),.clk(gclk));
	jdff dff_A_FvSoSi5H3_2(.dout(w_n566_0[2]),.din(w_dff_A_FvSoSi5H3_2),.clk(gclk));
	jdff dff_A_ayT2PZaO5_2(.dout(w_dff_A_FvSoSi5H3_2),.din(w_dff_A_ayT2PZaO5_2),.clk(gclk));
	jdff dff_A_4EdfMcyJ7_2(.dout(w_dff_A_ayT2PZaO5_2),.din(w_dff_A_4EdfMcyJ7_2),.clk(gclk));
	jdff dff_A_QDiCPetD4_2(.dout(w_dff_A_4EdfMcyJ7_2),.din(w_dff_A_QDiCPetD4_2),.clk(gclk));
	jdff dff_A_a77PsJUx4_2(.dout(w_dff_A_QDiCPetD4_2),.din(w_dff_A_a77PsJUx4_2),.clk(gclk));
	jdff dff_A_rUnl0ppz2_0(.dout(w_G213_0[0]),.din(w_dff_A_rUnl0ppz2_0),.clk(gclk));
	jdff dff_A_skkI8VF88_2(.dout(w_G213_0[2]),.din(w_dff_A_skkI8VF88_2),.clk(gclk));
	jdff dff_A_YSi94fau9_2(.dout(w_dff_A_skkI8VF88_2),.din(w_dff_A_YSi94fau9_2),.clk(gclk));
	jdff dff_A_AuzAKPCc6_1(.dout(w_G343_0[1]),.din(w_dff_A_AuzAKPCc6_1),.clk(gclk));
	jdff dff_A_hM3THRsg9_1(.dout(w_dff_A_AuzAKPCc6_1),.din(w_dff_A_hM3THRsg9_1),.clk(gclk));
	jdff dff_A_JmW3Ihxc8_1(.dout(w_dff_A_hM3THRsg9_1),.din(w_dff_A_JmW3Ihxc8_1),.clk(gclk));
	jdff dff_A_WVSrChD69_1(.dout(w_dff_A_JmW3Ihxc8_1),.din(w_dff_A_WVSrChD69_1),.clk(gclk));
	jdff dff_A_bnC8QV0j7_2(.dout(w_n198_0[2]),.din(w_dff_A_bnC8QV0j7_2),.clk(gclk));
	jdff dff_B_YnaDh83O0_1(.din(n193),.dout(w_dff_B_YnaDh83O0_1),.clk(gclk));
	jdff dff_B_cuojKOfz4_1(.din(w_dff_B_YnaDh83O0_1),.dout(w_dff_B_cuojKOfz4_1),.clk(gclk));
	jdff dff_A_Su0dW8rr4_1(.dout(w_G190_4[1]),.din(w_dff_A_Su0dW8rr4_1),.clk(gclk));
	jdff dff_A_0yhDhK1R7_2(.dout(w_G190_4[2]),.din(w_dff_A_0yhDhK1R7_2),.clk(gclk));
	jdff dff_A_R3WQr2sD2_2(.dout(w_dff_A_0yhDhK1R7_2),.din(w_dff_A_R3WQr2sD2_2),.clk(gclk));
	jdff dff_A_ijVSSTmt9_0(.dout(w_G190_1[0]),.din(w_dff_A_ijVSSTmt9_0),.clk(gclk));
	jdff dff_A_tpmf8KZl1_0(.dout(w_dff_A_ijVSSTmt9_0),.din(w_dff_A_tpmf8KZl1_0),.clk(gclk));
	jdff dff_A_3YjxHHOi9_0(.dout(w_dff_A_tpmf8KZl1_0),.din(w_dff_A_3YjxHHOi9_0),.clk(gclk));
	jdff dff_A_JWCzRV0Q8_0(.dout(w_dff_A_3YjxHHOi9_0),.din(w_dff_A_JWCzRV0Q8_0),.clk(gclk));
	jdff dff_A_naQTATWe7_0(.dout(w_dff_A_JWCzRV0Q8_0),.din(w_dff_A_naQTATWe7_0),.clk(gclk));
	jdff dff_A_ZoHb93cZ1_0(.dout(w_G190_0[0]),.din(w_dff_A_ZoHb93cZ1_0),.clk(gclk));
	jdff dff_A_vQANGHd58_0(.dout(w_dff_A_ZoHb93cZ1_0),.din(w_dff_A_vQANGHd58_0),.clk(gclk));
	jdff dff_A_bMsbkEkt6_2(.dout(w_G190_0[2]),.din(w_dff_A_bMsbkEkt6_2),.clk(gclk));
	jdff dff_A_GQPiGC388_2(.dout(w_dff_A_bMsbkEkt6_2),.din(w_dff_A_GQPiGC388_2),.clk(gclk));
	jdff dff_A_NOvU5JuC3_2(.dout(w_dff_A_GQPiGC388_2),.din(w_dff_A_NOvU5JuC3_2),.clk(gclk));
	jdff dff_A_x3XqxMef9_2(.dout(w_dff_A_NOvU5JuC3_2),.din(w_dff_A_x3XqxMef9_2),.clk(gclk));
	jdff dff_A_lTn0LJ062_2(.dout(w_dff_A_x3XqxMef9_2),.din(w_dff_A_lTn0LJ062_2),.clk(gclk));
	jdff dff_A_TZ7yFRSH9_2(.dout(w_dff_A_lTn0LJ062_2),.din(w_dff_A_TZ7yFRSH9_2),.clk(gclk));
	jdff dff_A_ew18bozs6_2(.dout(w_dff_A_TZ7yFRSH9_2),.din(w_dff_A_ew18bozs6_2),.clk(gclk));
	jdff dff_A_cepuc8ky3_2(.dout(w_G200_0[2]),.din(w_dff_A_cepuc8ky3_2),.clk(gclk));
	jdff dff_A_DZ2umtH22_2(.dout(w_dff_A_cepuc8ky3_2),.din(w_dff_A_DZ2umtH22_2),.clk(gclk));
	jdff dff_A_8FFohwbb2_2(.dout(w_dff_A_DZ2umtH22_2),.din(w_dff_A_8FFohwbb2_2),.clk(gclk));
	jdff dff_A_5EsIkV012_2(.dout(w_dff_A_8FFohwbb2_2),.din(w_dff_A_5EsIkV012_2),.clk(gclk));
	jdff dff_A_PRPk6bvs1_2(.dout(w_dff_A_5EsIkV012_2),.din(w_dff_A_PRPk6bvs1_2),.clk(gclk));
	jdff dff_A_jb9Wwk7I8_2(.dout(w_dff_A_PRPk6bvs1_2),.din(w_dff_A_jb9Wwk7I8_2),.clk(gclk));
	jdff dff_A_m8AjJmOU7_2(.dout(w_dff_A_jb9Wwk7I8_2),.din(w_dff_A_m8AjJmOU7_2),.clk(gclk));
	jdff dff_A_gXQuaMnl3_2(.dout(w_dff_A_m8AjJmOU7_2),.din(w_dff_A_gXQuaMnl3_2),.clk(gclk));
	jdff dff_A_ZypU1M0j6_1(.dout(w_n192_0[1]),.din(w_dff_A_ZypU1M0j6_1),.clk(gclk));
	jdff dff_A_KNfRQKVM6_1(.dout(w_dff_A_ZypU1M0j6_1),.din(w_dff_A_KNfRQKVM6_1),.clk(gclk));
	jdff dff_B_Ji80iO3W0_1(.din(n162),.dout(w_dff_B_Ji80iO3W0_1),.clk(gclk));
	jdff dff_B_OEsLG4yF6_1(.din(w_dff_B_Ji80iO3W0_1),.dout(w_dff_B_OEsLG4yF6_1),.clk(gclk));
	jdff dff_A_A6Ofxp4u6_1(.dout(w_n190_0[1]),.din(w_dff_A_A6Ofxp4u6_1),.clk(gclk));
	jdff dff_A_ZN1HbWSE0_1(.dout(w_n189_2[1]),.din(w_dff_A_ZN1HbWSE0_1),.clk(gclk));
	jdff dff_A_WxnTA56b3_2(.dout(w_n189_2[2]),.din(w_dff_A_WxnTA56b3_2),.clk(gclk));
	jdff dff_A_udFISggS8_0(.dout(w_n189_0[0]),.din(w_dff_A_udFISggS8_0),.clk(gclk));
	jdff dff_A_Z6NkXakE9_0(.dout(w_dff_A_udFISggS8_0),.din(w_dff_A_Z6NkXakE9_0),.clk(gclk));
	jdff dff_A_hhute4kg0_0(.dout(w_dff_A_Z6NkXakE9_0),.din(w_dff_A_hhute4kg0_0),.clk(gclk));
	jdff dff_A_Kqjde74b7_0(.dout(w_dff_A_hhute4kg0_0),.din(w_dff_A_Kqjde74b7_0),.clk(gclk));
	jdff dff_A_UtHLjOxk6_0(.dout(w_dff_A_Kqjde74b7_0),.din(w_dff_A_UtHLjOxk6_0),.clk(gclk));
	jdff dff_A_b53XyEOm5_0(.dout(w_dff_A_UtHLjOxk6_0),.din(w_dff_A_b53XyEOm5_0),.clk(gclk));
	jdff dff_A_PB8t3Hvz9_1(.dout(w_n189_0[1]),.din(w_dff_A_PB8t3Hvz9_1),.clk(gclk));
	jdff dff_A_H0zqYxPy1_1(.dout(w_dff_A_PB8t3Hvz9_1),.din(w_dff_A_H0zqYxPy1_1),.clk(gclk));
	jdff dff_A_Er0bsRYb9_1(.dout(w_dff_A_H0zqYxPy1_1),.din(w_dff_A_Er0bsRYb9_1),.clk(gclk));
	jdff dff_A_udnaR6Ee8_1(.dout(w_dff_A_Er0bsRYb9_1),.din(w_dff_A_udnaR6Ee8_1),.clk(gclk));
	jdff dff_A_eU84hw6U8_1(.dout(w_dff_A_udnaR6Ee8_1),.din(w_dff_A_eU84hw6U8_1),.clk(gclk));
	jdff dff_A_OGcwN2MC2_1(.dout(w_dff_A_eU84hw6U8_1),.din(w_dff_A_OGcwN2MC2_1),.clk(gclk));
	jdff dff_A_N0BEEMJX4_0(.dout(w_G179_2[0]),.din(w_dff_A_N0BEEMJX4_0),.clk(gclk));
	jdff dff_A_DjXYqC9V1_0(.dout(w_dff_A_N0BEEMJX4_0),.din(w_dff_A_DjXYqC9V1_0),.clk(gclk));
	jdff dff_A_xkG9Hc0j8_0(.dout(w_dff_A_DjXYqC9V1_0),.din(w_dff_A_xkG9Hc0j8_0),.clk(gclk));
	jdff dff_A_yP34O01m9_0(.dout(w_dff_A_xkG9Hc0j8_0),.din(w_dff_A_yP34O01m9_0),.clk(gclk));
	jdff dff_A_ecswXMSM3_0(.dout(w_dff_A_yP34O01m9_0),.din(w_dff_A_ecswXMSM3_0),.clk(gclk));
	jdff dff_A_TMEXgCiV3_0(.dout(w_dff_A_ecswXMSM3_0),.din(w_dff_A_TMEXgCiV3_0),.clk(gclk));
	jdff dff_A_LCUuEBXe0_0(.dout(w_dff_A_TMEXgCiV3_0),.din(w_dff_A_LCUuEBXe0_0),.clk(gclk));
	jdff dff_A_RKSuQUOB6_0(.dout(w_dff_A_LCUuEBXe0_0),.din(w_dff_A_RKSuQUOB6_0),.clk(gclk));
	jdff dff_A_1UgETKAM2_1(.dout(w_G179_2[1]),.din(w_dff_A_1UgETKAM2_1),.clk(gclk));
	jdff dff_A_1LD0OQSW4_1(.dout(w_dff_A_1UgETKAM2_1),.din(w_dff_A_1LD0OQSW4_1),.clk(gclk));
	jdff dff_A_5IjsnvRM4_1(.dout(w_dff_A_1LD0OQSW4_1),.din(w_dff_A_5IjsnvRM4_1),.clk(gclk));
	jdff dff_A_faN238Rh5_1(.dout(w_dff_A_5IjsnvRM4_1),.din(w_dff_A_faN238Rh5_1),.clk(gclk));
	jdff dff_A_9WTQOPrW0_1(.dout(w_dff_A_faN238Rh5_1),.din(w_dff_A_9WTQOPrW0_1),.clk(gclk));
	jdff dff_A_81qg6Jm97_1(.dout(w_dff_A_9WTQOPrW0_1),.din(w_dff_A_81qg6Jm97_1),.clk(gclk));
	jdff dff_A_r0X3Rd9Y4_1(.dout(w_dff_A_81qg6Jm97_1),.din(w_dff_A_r0X3Rd9Y4_1),.clk(gclk));
	jdff dff_A_2EJuJVo33_1(.dout(w_dff_A_r0X3Rd9Y4_1),.din(w_dff_A_2EJuJVo33_1),.clk(gclk));
	jdff dff_A_ElvWcEP37_0(.dout(w_G179_0[0]),.din(w_dff_A_ElvWcEP37_0),.clk(gclk));
	jdff dff_A_v2CFLhBw2_0(.dout(w_dff_A_ElvWcEP37_0),.din(w_dff_A_v2CFLhBw2_0),.clk(gclk));
	jdff dff_A_zq8Txwaj5_0(.dout(w_dff_A_v2CFLhBw2_0),.din(w_dff_A_zq8Txwaj5_0),.clk(gclk));
	jdff dff_A_ubxbXNuN4_0(.dout(w_dff_A_zq8Txwaj5_0),.din(w_dff_A_ubxbXNuN4_0),.clk(gclk));
	jdff dff_A_28Uh1vw04_0(.dout(w_dff_A_ubxbXNuN4_0),.din(w_dff_A_28Uh1vw04_0),.clk(gclk));
	jdff dff_A_PLkSvc9g4_0(.dout(w_dff_A_28Uh1vw04_0),.din(w_dff_A_PLkSvc9g4_0),.clk(gclk));
	jdff dff_A_belxD7F03_0(.dout(w_dff_A_PLkSvc9g4_0),.din(w_dff_A_belxD7F03_0),.clk(gclk));
	jdff dff_A_oNI79irw8_0(.dout(w_dff_A_belxD7F03_0),.din(w_dff_A_oNI79irw8_0),.clk(gclk));
	jdff dff_A_g9nn8Zc14_1(.dout(w_n186_0[1]),.din(w_dff_A_g9nn8Zc14_1),.clk(gclk));
	jdff dff_B_Tqm4dI2w6_0(.din(n184),.dout(w_dff_B_Tqm4dI2w6_0),.clk(gclk));
	jdff dff_A_8z1FTl5P0_0(.dout(w_G270_0[0]),.din(w_dff_A_8z1FTl5P0_0),.clk(gclk));
	jdff dff_A_aKkaL1z45_0(.dout(w_dff_A_8z1FTl5P0_0),.din(w_dff_A_aKkaL1z45_0),.clk(gclk));
	jdff dff_A_oU1nba1o6_0(.dout(w_dff_A_aKkaL1z45_0),.din(w_dff_A_oU1nba1o6_0),.clk(gclk));
	jdff dff_A_TgPEKW4v9_1(.dout(w_G270_0[1]),.din(w_dff_A_TgPEKW4v9_1),.clk(gclk));
	jdff dff_B_RrvFTnon4_1(.din(n174),.dout(w_dff_B_RrvFTnon4_1),.clk(gclk));
	jdff dff_B_PzI6ITzR8_1(.din(n175),.dout(w_dff_B_PzI6ITzR8_1),.clk(gclk));
	jdff dff_B_Qf4tPweB9_1(.din(w_dff_B_PzI6ITzR8_1),.dout(w_dff_B_Qf4tPweB9_1),.clk(gclk));
	jdff dff_A_9umbvbKS6_0(.dout(w_G257_1[0]),.din(w_dff_A_9umbvbKS6_0),.clk(gclk));
	jdff dff_A_Qvpf57IH7_0(.dout(w_dff_A_9umbvbKS6_0),.din(w_dff_A_Qvpf57IH7_0),.clk(gclk));
	jdff dff_A_XszD7M3c5_1(.dout(w_G257_0[1]),.din(w_dff_A_XszD7M3c5_1),.clk(gclk));
	jdff dff_A_AC2I0mRQ3_1(.dout(w_dff_A_XszD7M3c5_1),.din(w_dff_A_AC2I0mRQ3_1),.clk(gclk));
	jdff dff_A_kuQLI3Vo2_1(.dout(w_dff_A_AC2I0mRQ3_1),.din(w_dff_A_kuQLI3Vo2_1),.clk(gclk));
	jdff dff_A_HVUG87jc0_2(.dout(w_G257_0[2]),.din(w_dff_A_HVUG87jc0_2),.clk(gclk));
	jdff dff_A_7LBgXwEW5_2(.dout(w_dff_A_HVUG87jc0_2),.din(w_dff_A_7LBgXwEW5_2),.clk(gclk));
	jdff dff_A_mLm1PJlt2_0(.dout(w_G303_2[0]),.din(w_dff_A_mLm1PJlt2_0),.clk(gclk));
	jdff dff_A_HeBLclxv7_0(.dout(w_dff_A_mLm1PJlt2_0),.din(w_dff_A_HeBLclxv7_0),.clk(gclk));
	jdff dff_A_y9csACmr9_0(.dout(w_dff_A_HeBLclxv7_0),.din(w_dff_A_y9csACmr9_0),.clk(gclk));
	jdff dff_A_qmCoNXiI4_1(.dout(w_G303_2[1]),.din(w_dff_A_qmCoNXiI4_1),.clk(gclk));
	jdff dff_A_nKLqndak4_1(.dout(w_dff_A_qmCoNXiI4_1),.din(w_dff_A_nKLqndak4_1),.clk(gclk));
	jdff dff_A_tGoKlo0V2_1(.dout(w_dff_A_nKLqndak4_1),.din(w_dff_A_tGoKlo0V2_1),.clk(gclk));
	jdff dff_A_uwjvYkAu9_0(.dout(w_G303_0[0]),.din(w_dff_A_uwjvYkAu9_0),.clk(gclk));
	jdff dff_A_wreUxZbJ9_0(.dout(w_dff_A_uwjvYkAu9_0),.din(w_dff_A_wreUxZbJ9_0),.clk(gclk));
	jdff dff_A_cftYHiFH1_0(.dout(w_dff_A_wreUxZbJ9_0),.din(w_dff_A_cftYHiFH1_0),.clk(gclk));
	jdff dff_A_dZ7D7Tmw4_2(.dout(w_G303_0[2]),.din(w_dff_A_dZ7D7Tmw4_2),.clk(gclk));
	jdff dff_A_pfWE9oTo5_2(.dout(w_dff_A_dZ7D7Tmw4_2),.din(w_dff_A_pfWE9oTo5_2),.clk(gclk));
	jdff dff_A_Fw7xNyJB7_2(.dout(w_dff_A_pfWE9oTo5_2),.din(w_dff_A_Fw7xNyJB7_2),.clk(gclk));
	jdff dff_A_Az6zVtTd4_2(.dout(w_dff_A_Fw7xNyJB7_2),.din(w_dff_A_Az6zVtTd4_2),.clk(gclk));
	jdff dff_A_vjQCyBhw6_2(.dout(w_G1698_0[2]),.din(w_dff_A_vjQCyBhw6_2),.clk(gclk));
	jdff dff_A_gnrdzkWR0_0(.dout(w_G264_0[0]),.din(w_dff_A_gnrdzkWR0_0),.clk(gclk));
	jdff dff_A_WCp84g3m6_0(.dout(w_dff_A_gnrdzkWR0_0),.din(w_dff_A_WCp84g3m6_0),.clk(gclk));
	jdff dff_A_UybTJBfR0_0(.dout(w_dff_A_WCp84g3m6_0),.din(w_dff_A_UybTJBfR0_0),.clk(gclk));
	jdff dff_A_vj4kD5vR4_1(.dout(w_G264_0[1]),.din(w_dff_A_vj4kD5vR4_1),.clk(gclk));
	jdff dff_A_wW8gMsRw4_1(.dout(w_dff_A_vj4kD5vR4_1),.din(w_dff_A_wW8gMsRw4_1),.clk(gclk));
	jdff dff_A_pMvMwwFC3_1(.dout(w_n172_4[1]),.din(w_dff_A_pMvMwwFC3_1),.clk(gclk));
	jdff dff_A_vga5hyTG0_1(.dout(w_dff_A_pMvMwwFC3_1),.din(w_dff_A_vga5hyTG0_1),.clk(gclk));
	jdff dff_A_GKGGy3Mq8_2(.dout(w_n172_4[2]),.din(w_dff_A_GKGGy3Mq8_2),.clk(gclk));
	jdff dff_A_nvMEuQpG9_2(.dout(w_dff_A_GKGGy3Mq8_2),.din(w_dff_A_nvMEuQpG9_2),.clk(gclk));
	jdff dff_A_dOZL61cq6_1(.dout(w_n172_1[1]),.din(w_dff_A_dOZL61cq6_1),.clk(gclk));
	jdff dff_A_7tTiqfhT6_1(.dout(w_dff_A_dOZL61cq6_1),.din(w_dff_A_7tTiqfhT6_1),.clk(gclk));
	jdff dff_A_8o0l8bfO3_2(.dout(w_n172_1[2]),.din(w_dff_A_8o0l8bfO3_2),.clk(gclk));
	jdff dff_A_3AAwax0a6_2(.dout(w_dff_A_8o0l8bfO3_2),.din(w_dff_A_3AAwax0a6_2),.clk(gclk));
	jdff dff_A_M86Y64q06_1(.dout(w_n172_0[1]),.din(w_dff_A_M86Y64q06_1),.clk(gclk));
	jdff dff_A_IxbcIBxm6_1(.dout(w_dff_A_M86Y64q06_1),.din(w_dff_A_IxbcIBxm6_1),.clk(gclk));
	jdff dff_A_Jo7k03HD9_2(.dout(w_n172_0[2]),.din(w_dff_A_Jo7k03HD9_2),.clk(gclk));
	jdff dff_A_hSgxQEJA9_2(.dout(w_dff_A_Jo7k03HD9_2),.din(w_dff_A_hSgxQEJA9_2),.clk(gclk));
	jdff dff_A_b1EAzkv06_2(.dout(w_n170_0[2]),.din(w_dff_A_b1EAzkv06_2),.clk(gclk));
	jdff dff_B_WnJKDA8q3_3(.din(n170),.dout(w_dff_B_WnJKDA8q3_3),.clk(gclk));
	jdff dff_A_QPcPdCI90_1(.dout(w_n167_0[1]),.din(w_dff_A_QPcPdCI90_1),.clk(gclk));
	jdff dff_A_Rb3AcJSg6_0(.dout(w_G274_0[0]),.din(w_dff_A_Rb3AcJSg6_0),.clk(gclk));
	jdff dff_A_YNlKx5VQ6_0(.dout(w_dff_A_Rb3AcJSg6_0),.din(w_dff_A_YNlKx5VQ6_0),.clk(gclk));
	jdff dff_A_GCs8Nm6Y4_2(.dout(w_G274_0[2]),.din(w_dff_A_GCs8Nm6Y4_2),.clk(gclk));
	jdff dff_A_yqzXBbLR1_2(.dout(w_dff_A_GCs8Nm6Y4_2),.din(w_dff_A_yqzXBbLR1_2),.clk(gclk));
	jdff dff_A_ZYdtO75G0_2(.dout(w_dff_A_yqzXBbLR1_2),.din(w_dff_A_ZYdtO75G0_2),.clk(gclk));
	jdff dff_A_QCW8hcPI2_1(.dout(w_n165_0[1]),.din(w_dff_A_QCW8hcPI2_1),.clk(gclk));
	jdff dff_A_iD4J6MS45_1(.dout(w_G45_1[1]),.din(w_dff_A_iD4J6MS45_1),.clk(gclk));
	jdff dff_A_JXJGeXc22_0(.dout(w_n142_1[0]),.din(w_dff_A_JXJGeXc22_0),.clk(gclk));
	jdff dff_A_1Pahpig79_0(.dout(w_dff_A_JXJGeXc22_0),.din(w_dff_A_1Pahpig79_0),.clk(gclk));
	jdff dff_A_4Yknphgw5_0(.dout(w_dff_A_1Pahpig79_0),.din(w_dff_A_4Yknphgw5_0),.clk(gclk));
	jdff dff_A_jvI5Dpa70_0(.dout(w_dff_A_4Yknphgw5_0),.din(w_dff_A_jvI5Dpa70_0),.clk(gclk));
	jdff dff_A_8MA6hMpj0_0(.dout(w_dff_A_jvI5Dpa70_0),.din(w_dff_A_8MA6hMpj0_0),.clk(gclk));
	jdff dff_A_cWKHglpW6_0(.dout(w_dff_A_8MA6hMpj0_0),.din(w_dff_A_cWKHglpW6_0),.clk(gclk));
	jdff dff_A_RFIN0BPS2_0(.dout(w_dff_A_cWKHglpW6_0),.din(w_dff_A_RFIN0BPS2_0),.clk(gclk));
	jdff dff_A_B9Pl3UY61_0(.dout(w_dff_A_RFIN0BPS2_0),.din(w_dff_A_B9Pl3UY61_0),.clk(gclk));
	jdff dff_A_mXN2Xjw79_0(.dout(w_dff_A_B9Pl3UY61_0),.din(w_dff_A_mXN2Xjw79_0),.clk(gclk));
	jdff dff_A_amIHWbpj5_0(.dout(w_dff_A_mXN2Xjw79_0),.din(w_dff_A_amIHWbpj5_0),.clk(gclk));
	jdff dff_A_2NR8m91N7_0(.dout(w_dff_A_amIHWbpj5_0),.din(w_dff_A_2NR8m91N7_0),.clk(gclk));
	jdff dff_A_3sbJ8hsb1_0(.dout(w_dff_A_2NR8m91N7_0),.din(w_dff_A_3sbJ8hsb1_0),.clk(gclk));
	jdff dff_A_v6RcmkOt3_0(.dout(w_dff_A_3sbJ8hsb1_0),.din(w_dff_A_v6RcmkOt3_0),.clk(gclk));
	jdff dff_A_oHxxIHUn5_0(.dout(w_dff_A_v6RcmkOt3_0),.din(w_dff_A_oHxxIHUn5_0),.clk(gclk));
	jdff dff_A_FjzdyPWx7_0(.dout(w_dff_A_oHxxIHUn5_0),.din(w_dff_A_FjzdyPWx7_0),.clk(gclk));
	jdff dff_A_rpg1F2RK8_0(.dout(w_dff_A_FjzdyPWx7_0),.din(w_dff_A_rpg1F2RK8_0),.clk(gclk));
	jdff dff_A_ZszvsuPY6_0(.dout(w_dff_A_rpg1F2RK8_0),.din(w_dff_A_ZszvsuPY6_0),.clk(gclk));
	jdff dff_A_lhYU8i2i5_0(.dout(w_dff_A_ZszvsuPY6_0),.din(w_dff_A_lhYU8i2i5_0),.clk(gclk));
	jdff dff_A_EwrqlWyp2_1(.dout(w_n163_1[1]),.din(w_dff_A_EwrqlWyp2_1),.clk(gclk));
	jdff dff_A_2sAm4jEc0_1(.dout(w_G169_3[1]),.din(w_dff_A_2sAm4jEc0_1),.clk(gclk));
	jdff dff_A_wabDsVEP0_1(.dout(w_dff_A_2sAm4jEc0_1),.din(w_dff_A_wabDsVEP0_1),.clk(gclk));
	jdff dff_A_m6esQfdP1_1(.dout(w_dff_A_wabDsVEP0_1),.din(w_dff_A_m6esQfdP1_1),.clk(gclk));
	jdff dff_A_R06S8aZw0_1(.dout(w_dff_A_m6esQfdP1_1),.din(w_dff_A_R06S8aZw0_1),.clk(gclk));
	jdff dff_A_lIULxlXG7_1(.dout(w_dff_A_R06S8aZw0_1),.din(w_dff_A_lIULxlXG7_1),.clk(gclk));
	jdff dff_A_W1E9wiDD9_1(.dout(w_dff_A_lIULxlXG7_1),.din(w_dff_A_W1E9wiDD9_1),.clk(gclk));
	jdff dff_A_HzEUQJyU0_1(.dout(w_dff_A_W1E9wiDD9_1),.din(w_dff_A_HzEUQJyU0_1),.clk(gclk));
	jdff dff_A_gNdOfnno1_1(.dout(w_dff_A_HzEUQJyU0_1),.din(w_dff_A_gNdOfnno1_1),.clk(gclk));
	jdff dff_A_q2xWHlDq8_0(.dout(w_G169_0[0]),.din(w_dff_A_q2xWHlDq8_0),.clk(gclk));
	jdff dff_A_rTxpwddn3_1(.dout(w_G169_0[1]),.din(w_dff_A_rTxpwddn3_1),.clk(gclk));
	jdff dff_A_wuTDcEKF8_1(.dout(w_dff_A_rTxpwddn3_1),.din(w_dff_A_wuTDcEKF8_1),.clk(gclk));
	jdff dff_A_2XCjO6Ip1_1(.dout(w_dff_A_wuTDcEKF8_1),.din(w_dff_A_2XCjO6Ip1_1),.clk(gclk));
	jdff dff_A_LNEZeKsk8_1(.dout(w_dff_A_2XCjO6Ip1_1),.din(w_dff_A_LNEZeKsk8_1),.clk(gclk));
	jdff dff_A_GYbrrVB18_1(.dout(w_dff_A_LNEZeKsk8_1),.din(w_dff_A_GYbrrVB18_1),.clk(gclk));
	jdff dff_A_XsW0EsCf7_1(.dout(w_dff_A_GYbrrVB18_1),.din(w_dff_A_XsW0EsCf7_1),.clk(gclk));
	jdff dff_A_Dy3TAhzW2_1(.dout(w_dff_A_XsW0EsCf7_1),.din(w_dff_A_Dy3TAhzW2_1),.clk(gclk));
	jdff dff_A_OUi7JFIo4_1(.dout(w_n161_0[1]),.din(w_dff_A_OUi7JFIo4_1),.clk(gclk));
	jdff dff_A_Kmx4IvMP5_1(.dout(w_dff_A_OUi7JFIo4_1),.din(w_dff_A_Kmx4IvMP5_1),.clk(gclk));
	jdff dff_B_WZdnyJp83_0(.din(n159),.dout(w_dff_B_WZdnyJp83_0),.clk(gclk));
	jdff dff_B_hEwfdFJC4_0(.din(w_dff_B_WZdnyJp83_0),.dout(w_dff_B_hEwfdFJC4_0),.clk(gclk));
	jdff dff_A_X07PXF714_0(.dout(w_n105_1[0]),.din(w_dff_A_X07PXF714_0),.clk(gclk));
	jdff dff_A_5Bk3phfE6_0(.dout(w_dff_A_X07PXF714_0),.din(w_dff_A_5Bk3phfE6_0),.clk(gclk));
	jdff dff_A_ILUERALf3_1(.dout(w_n105_0[1]),.din(w_dff_A_ILUERALf3_1),.clk(gclk));
	jdff dff_A_Xp4JgKbh6_1(.dout(w_dff_A_ILUERALf3_1),.din(w_dff_A_Xp4JgKbh6_1),.clk(gclk));
	jdff dff_A_Ik8vCPxA0_1(.dout(w_dff_A_Xp4JgKbh6_1),.din(w_dff_A_Ik8vCPxA0_1),.clk(gclk));
	jdff dff_A_Hx5Huinu0_2(.dout(w_n105_0[2]),.din(w_dff_A_Hx5Huinu0_2),.clk(gclk));
	jdff dff_A_55jDWv245_2(.dout(w_dff_A_Hx5Huinu0_2),.din(w_dff_A_55jDWv245_2),.clk(gclk));
	jdff dff_B_O5lDCoGi9_1(.din(n150),.dout(w_dff_B_O5lDCoGi9_1),.clk(gclk));
	jdff dff_B_6s69clhL3_1(.din(w_dff_B_O5lDCoGi9_1),.dout(w_dff_B_6s69clhL3_1),.clk(gclk));
	jdff dff_B_ThrNonlU3_1(.din(w_dff_B_6s69clhL3_1),.dout(w_dff_B_ThrNonlU3_1),.clk(gclk));
	jdff dff_A_E5wgSxP68_0(.dout(w_G97_4[0]),.din(w_dff_A_E5wgSxP68_0),.clk(gclk));
	jdff dff_A_zZy4bo4X3_1(.dout(w_G97_1[1]),.din(w_dff_A_zZy4bo4X3_1),.clk(gclk));
	jdff dff_A_SZoFlOny9_1(.dout(w_dff_A_zZy4bo4X3_1),.din(w_dff_A_SZoFlOny9_1),.clk(gclk));
	jdff dff_A_jZz3IHDG8_1(.dout(w_dff_A_SZoFlOny9_1),.din(w_dff_A_jZz3IHDG8_1),.clk(gclk));
	jdff dff_A_CfHpfQCw4_2(.dout(w_G97_1[2]),.din(w_dff_A_CfHpfQCw4_2),.clk(gclk));
	jdff dff_A_77fyP2ar1_2(.dout(w_dff_A_CfHpfQCw4_2),.din(w_dff_A_77fyP2ar1_2),.clk(gclk));
	jdff dff_A_2dNZana21_2(.dout(w_dff_A_77fyP2ar1_2),.din(w_dff_A_2dNZana21_2),.clk(gclk));
	jdff dff_A_WhbXSYJK8_1(.dout(w_G97_0[1]),.din(w_dff_A_WhbXSYJK8_1),.clk(gclk));
	jdff dff_A_Hz8IvoM91_1(.dout(w_dff_A_WhbXSYJK8_1),.din(w_dff_A_Hz8IvoM91_1),.clk(gclk));
	jdff dff_A_4EL6Kdd02_1(.dout(w_dff_A_Hz8IvoM91_1),.din(w_dff_A_4EL6Kdd02_1),.clk(gclk));
	jdff dff_A_jAqQNxKk1_2(.dout(w_n153_2[2]),.din(w_dff_A_jAqQNxKk1_2),.clk(gclk));
	jdff dff_A_t6R5PWtB3_2(.dout(w_dff_A_jAqQNxKk1_2),.din(w_dff_A_t6R5PWtB3_2),.clk(gclk));
	jdff dff_A_twm6ZtqJ4_2(.dout(w_dff_A_t6R5PWtB3_2),.din(w_dff_A_twm6ZtqJ4_2),.clk(gclk));
	jdff dff_A_dZWH8cyL6_2(.dout(w_dff_A_twm6ZtqJ4_2),.din(w_dff_A_dZWH8cyL6_2),.clk(gclk));
	jdff dff_A_oBcMi1la7_2(.dout(w_n153_0[2]),.din(w_dff_A_oBcMi1la7_2),.clk(gclk));
	jdff dff_A_zvQa7yxe5_2(.dout(w_dff_A_oBcMi1la7_2),.din(w_dff_A_zvQa7yxe5_2),.clk(gclk));
	jdff dff_A_xZyeqGsy9_2(.dout(w_dff_A_zvQa7yxe5_2),.din(w_dff_A_xZyeqGsy9_2),.clk(gclk));
	jdff dff_A_2EJxM0j54_0(.dout(w_n152_0[0]),.din(w_dff_A_2EJxM0j54_0),.clk(gclk));
	jdff dff_A_3QeCQqy86_0(.dout(w_dff_A_2EJxM0j54_0),.din(w_dff_A_3QeCQqy86_0),.clk(gclk));
	jdff dff_A_dfW7T59s0_2(.dout(w_n152_0[2]),.din(w_dff_A_dfW7T59s0_2),.clk(gclk));
	jdff dff_A_pDj358Ch0_0(.dout(w_G283_3[0]),.din(w_dff_A_pDj358Ch0_0),.clk(gclk));
	jdff dff_A_C1G414EV2_0(.dout(w_dff_A_pDj358Ch0_0),.din(w_dff_A_C1G414EV2_0),.clk(gclk));
	jdff dff_A_M3o1gwDr0_0(.dout(w_dff_A_C1G414EV2_0),.din(w_dff_A_M3o1gwDr0_0),.clk(gclk));
	jdff dff_A_gPqY2UvA5_1(.dout(w_G283_3[1]),.din(w_dff_A_gPqY2UvA5_1),.clk(gclk));
	jdff dff_A_UEp8HpzD5_1(.dout(w_dff_A_gPqY2UvA5_1),.din(w_dff_A_UEp8HpzD5_1),.clk(gclk));
	jdff dff_A_YSKr3QoK9_1(.dout(w_dff_A_UEp8HpzD5_1),.din(w_dff_A_YSKr3QoK9_1),.clk(gclk));
	jdff dff_A_jMOKjR4O9_0(.dout(w_G283_0[0]),.din(w_dff_A_jMOKjR4O9_0),.clk(gclk));
	jdff dff_A_s1QWKw7V6_0(.dout(w_dff_A_jMOKjR4O9_0),.din(w_dff_A_s1QWKw7V6_0),.clk(gclk));
	jdff dff_A_4FvfAcLi4_0(.dout(w_dff_A_s1QWKw7V6_0),.din(w_dff_A_4FvfAcLi4_0),.clk(gclk));
	jdff dff_A_MHD1ok412_1(.dout(w_G283_0[1]),.din(w_dff_A_MHD1ok412_1),.clk(gclk));
	jdff dff_A_XyTCi7xB9_1(.dout(w_dff_A_MHD1ok412_1),.din(w_dff_A_XyTCi7xB9_1),.clk(gclk));
	jdff dff_A_u11qo1Wn5_1(.dout(w_dff_A_XyTCi7xB9_1),.din(w_dff_A_u11qo1Wn5_1),.clk(gclk));
	jdff dff_A_Q5xQh3CZ8_0(.dout(w_n151_6[0]),.din(w_dff_A_Q5xQh3CZ8_0),.clk(gclk));
	jdff dff_A_wFaGRlsO1_1(.dout(w_n151_1[1]),.din(w_dff_A_wFaGRlsO1_1),.clk(gclk));
	jdff dff_A_myOFtcpJ7_2(.dout(w_n151_1[2]),.din(w_dff_A_myOFtcpJ7_2),.clk(gclk));
	jdff dff_A_kKS7HTiK1_2(.dout(w_dff_A_myOFtcpJ7_2),.din(w_dff_A_kKS7HTiK1_2),.clk(gclk));
	jdff dff_A_FvBhCFCY3_0(.dout(w_G116_4[0]),.din(w_dff_A_FvBhCFCY3_0),.clk(gclk));
	jdff dff_A_dOsjTESK6_0(.dout(w_dff_A_FvBhCFCY3_0),.din(w_dff_A_dOsjTESK6_0),.clk(gclk));
	jdff dff_A_hiFDXRRs9_0(.dout(w_dff_A_dOsjTESK6_0),.din(w_dff_A_hiFDXRRs9_0),.clk(gclk));
	jdff dff_B_uJ3xOORm6_0(.din(n146),.dout(w_dff_B_uJ3xOORm6_0),.clk(gclk));
	jdff dff_B_l2pSoTrH7_0(.din(w_dff_B_uJ3xOORm6_0),.dout(w_dff_B_l2pSoTrH7_0),.clk(gclk));
	jdff dff_A_G2a5RTLJ1_0(.dout(w_n141_3[0]),.din(w_dff_A_G2a5RTLJ1_0),.clk(gclk));
	jdff dff_A_Qu1KcUFZ3_0(.dout(w_dff_A_G2a5RTLJ1_0),.din(w_dff_A_Qu1KcUFZ3_0),.clk(gclk));
	jdff dff_A_y5QVgwBk6_1(.dout(w_G33_12[1]),.din(w_dff_A_y5QVgwBk6_1),.clk(gclk));
	jdff dff_A_2A6upE0W0_2(.dout(w_G33_12[2]),.din(w_dff_A_2A6upE0W0_2),.clk(gclk));
	jdff dff_A_PWJAmKAm3_0(.dout(w_G33_0[0]),.din(w_dff_A_PWJAmKAm3_0),.clk(gclk));
	jdff dff_A_eWawSKNL7_0(.dout(w_dff_A_PWJAmKAm3_0),.din(w_dff_A_eWawSKNL7_0),.clk(gclk));
	jdff dff_A_x0xr0h3r0_0(.dout(w_dff_A_eWawSKNL7_0),.din(w_dff_A_x0xr0h3r0_0),.clk(gclk));
	jdff dff_A_Nx08apME8_0(.dout(w_n139_1[0]),.din(w_dff_A_Nx08apME8_0),.clk(gclk));
	jdff dff_A_cQeHUXR74_2(.dout(w_n139_1[2]),.din(w_dff_A_cQeHUXR74_2),.clk(gclk));
	jdff dff_A_nt1bhD358_0(.dout(w_G13_1[0]),.din(w_dff_A_nt1bhD358_0),.clk(gclk));
	jdff dff_A_X78oElrO3_0(.dout(w_dff_A_nt1bhD358_0),.din(w_dff_A_X78oElrO3_0),.clk(gclk));
	jdff dff_A_XMenjuw07_1(.dout(w_G13_1[1]),.din(w_dff_A_XMenjuw07_1),.clk(gclk));
	jdff dff_A_9bPYAUYV5_0(.dout(w_G116_5[0]),.din(w_dff_A_9bPYAUYV5_0),.clk(gclk));
	jdff dff_A_TlLqHoIT8_0(.dout(w_dff_A_9bPYAUYV5_0),.din(w_dff_A_TlLqHoIT8_0),.clk(gclk));
	jdff dff_A_kOZD6D7K7_0(.dout(w_dff_A_TlLqHoIT8_0),.din(w_dff_A_kOZD6D7K7_0),.clk(gclk));
	jdff dff_A_sitw6DNQ1_0(.dout(w_dff_A_kOZD6D7K7_0),.din(w_dff_A_sitw6DNQ1_0),.clk(gclk));
	jdff dff_A_BcLcGbZ95_0(.dout(w_dff_A_sitw6DNQ1_0),.din(w_dff_A_BcLcGbZ95_0),.clk(gclk));
	jdff dff_A_cPT0Uvut7_0(.dout(w_dff_A_BcLcGbZ95_0),.din(w_dff_A_cPT0Uvut7_0),.clk(gclk));
	jdff dff_A_xm7aeCbx9_1(.dout(w_G116_5[1]),.din(w_dff_A_xm7aeCbx9_1),.clk(gclk));
	jdff dff_A_CgkkcF1d8_2(.dout(w_G116_1[2]),.din(w_dff_A_CgkkcF1d8_2),.clk(gclk));
	jdff dff_A_dSGRiRnu7_2(.dout(w_dff_A_CgkkcF1d8_2),.din(w_dff_A_dSGRiRnu7_2),.clk(gclk));
	jdff dff_A_BHeSO7qT3_2(.dout(w_dff_A_dSGRiRnu7_2),.din(w_dff_A_BHeSO7qT3_2),.clk(gclk));
	jdff dff_A_2miAVqjQ8_1(.dout(w_G116_0[1]),.din(w_dff_A_2miAVqjQ8_1),.clk(gclk));
	jdff dff_A_uuSGeSRB5_1(.dout(w_dff_A_2miAVqjQ8_1),.din(w_dff_A_uuSGeSRB5_1),.clk(gclk));
	jdff dff_A_K6dqxKfC2_1(.dout(w_dff_A_uuSGeSRB5_1),.din(w_dff_A_K6dqxKfC2_1),.clk(gclk));
	jdff dff_A_CqsrBYPW0_2(.dout(w_G116_0[2]),.din(w_dff_A_CqsrBYPW0_2),.clk(gclk));
	jdff dff_A_0q8OseDv1_2(.dout(w_dff_A_CqsrBYPW0_2),.din(w_dff_A_0q8OseDv1_2),.clk(gclk));
	jdff dff_A_YMOYBBOY5_2(.dout(w_dff_A_0q8OseDv1_2),.din(w_dff_A_YMOYBBOY5_2),.clk(gclk));
	jdff dff_A_2czuDZR02_0(.dout(w_G330_0[0]),.din(w_dff_A_2czuDZR02_0),.clk(gclk));
	jdff dff_A_TSdrlmcq5_2(.dout(w_G330_0[2]),.din(w_dff_A_TSdrlmcq5_2),.clk(gclk));
	jdff dff_B_JYUQ1Fpi1_3(.din(G330),.dout(w_dff_B_JYUQ1Fpi1_3),.clk(gclk));
	jdff dff_B_pUTUUMiT7_3(.din(w_dff_B_JYUQ1Fpi1_3),.dout(w_dff_B_pUTUUMiT7_3),.clk(gclk));
	jdff dff_B_pnGVR7CE7_3(.din(w_dff_B_pUTUUMiT7_3),.dout(w_dff_B_pnGVR7CE7_3),.clk(gclk));
	jdff dff_B_sD7AOtzq4_3(.din(w_dff_B_pnGVR7CE7_3),.dout(w_dff_B_sD7AOtzq4_3),.clk(gclk));
	jdff dff_B_TEVwNqdr1_3(.din(w_dff_B_sD7AOtzq4_3),.dout(w_dff_B_TEVwNqdr1_3),.clk(gclk));
	jdff dff_B_KMQGD8eI4_3(.din(w_dff_B_TEVwNqdr1_3),.dout(w_dff_B_KMQGD8eI4_3),.clk(gclk));
	jdff dff_B_q7cY9u6B8_3(.din(w_dff_B_KMQGD8eI4_3),.dout(w_dff_B_q7cY9u6B8_3),.clk(gclk));
	jdff dff_B_fPAlwEwd1_3(.din(w_dff_B_q7cY9u6B8_3),.dout(w_dff_B_fPAlwEwd1_3),.clk(gclk));
	jdff dff_B_40nn1Lwz9_3(.din(w_dff_B_fPAlwEwd1_3),.dout(w_dff_B_40nn1Lwz9_3),.clk(gclk));
	jdff dff_B_sBT8MF3N1_3(.din(w_dff_B_40nn1Lwz9_3),.dout(w_dff_B_sBT8MF3N1_3),.clk(gclk));
	jdff dff_B_XgAtqVZK0_3(.din(w_dff_B_sBT8MF3N1_3),.dout(w_dff_B_XgAtqVZK0_3),.clk(gclk));
	jdff dff_B_xtK22yGs4_3(.din(w_dff_B_XgAtqVZK0_3),.dout(w_dff_B_xtK22yGs4_3),.clk(gclk));
	jdff dff_B_C95NgCdz3_3(.din(w_dff_B_xtK22yGs4_3),.dout(w_dff_B_C95NgCdz3_3),.clk(gclk));
	jdff dff_A_hgtqga5P4_0(.dout(w_n614_5[0]),.din(w_dff_A_hgtqga5P4_0),.clk(gclk));
	jdff dff_A_uUwQnBy62_0(.dout(w_dff_A_hgtqga5P4_0),.din(w_dff_A_uUwQnBy62_0),.clk(gclk));
	jdff dff_A_RisR2R3J7_0(.dout(w_dff_A_uUwQnBy62_0),.din(w_dff_A_RisR2R3J7_0),.clk(gclk));
	jdff dff_A_tjPHyHJn9_0(.dout(w_dff_A_RisR2R3J7_0),.din(w_dff_A_tjPHyHJn9_0),.clk(gclk));
	jdff dff_A_lgHh6aBg8_0(.dout(w_dff_A_tjPHyHJn9_0),.din(w_dff_A_lgHh6aBg8_0),.clk(gclk));
	jdff dff_A_Ekp2IG5W4_0(.dout(w_dff_A_lgHh6aBg8_0),.din(w_dff_A_Ekp2IG5W4_0),.clk(gclk));
	jdff dff_A_p0cEIKKC8_0(.dout(w_dff_A_Ekp2IG5W4_0),.din(w_dff_A_p0cEIKKC8_0),.clk(gclk));
	jdff dff_A_hfEkKlwp6_0(.dout(w_dff_A_p0cEIKKC8_0),.din(w_dff_A_hfEkKlwp6_0),.clk(gclk));
	jdff dff_A_Ry1rX72q4_0(.dout(w_dff_A_hfEkKlwp6_0),.din(w_dff_A_Ry1rX72q4_0),.clk(gclk));
	jdff dff_A_F3IObSgd7_0(.dout(w_dff_A_Ry1rX72q4_0),.din(w_dff_A_F3IObSgd7_0),.clk(gclk));
	jdff dff_A_IMLKiumh3_0(.dout(w_n614_1[0]),.din(w_dff_A_IMLKiumh3_0),.clk(gclk));
	jdff dff_A_Sl5uowRH7_0(.dout(w_dff_A_IMLKiumh3_0),.din(w_dff_A_Sl5uowRH7_0),.clk(gclk));
	jdff dff_A_6ly3l6PO0_2(.dout(w_n614_1[2]),.din(w_dff_A_6ly3l6PO0_2),.clk(gclk));
	jdff dff_A_jHpiulKy1_2(.dout(w_dff_A_6ly3l6PO0_2),.din(w_dff_A_jHpiulKy1_2),.clk(gclk));
	jdff dff_A_0H6vXaff9_2(.dout(w_dff_A_jHpiulKy1_2),.din(w_dff_A_0H6vXaff9_2),.clk(gclk));
	jdff dff_A_LyjjHCk80_2(.dout(w_dff_A_0H6vXaff9_2),.din(w_dff_A_LyjjHCk80_2),.clk(gclk));
	jdff dff_A_JpVKkyZd2_2(.dout(w_dff_A_LyjjHCk80_2),.din(w_dff_A_JpVKkyZd2_2),.clk(gclk));
	jdff dff_A_ZXPClYE07_2(.dout(w_dff_A_JpVKkyZd2_2),.din(w_dff_A_ZXPClYE07_2),.clk(gclk));
	jdff dff_A_CmrXkvrz6_2(.dout(w_dff_A_ZXPClYE07_2),.din(w_dff_A_CmrXkvrz6_2),.clk(gclk));
	jdff dff_A_QbbBYFjq7_2(.dout(w_dff_A_CmrXkvrz6_2),.din(w_dff_A_QbbBYFjq7_2),.clk(gclk));
	jdff dff_A_jBEXj34q3_2(.dout(w_dff_A_QbbBYFjq7_2),.din(w_dff_A_jBEXj34q3_2),.clk(gclk));
	jdff dff_A_lLMrfQwz0_2(.dout(w_dff_A_jBEXj34q3_2),.din(w_dff_A_lLMrfQwz0_2),.clk(gclk));
	jdff dff_A_I9tN8kjN3_2(.dout(w_dff_A_lLMrfQwz0_2),.din(w_dff_A_I9tN8kjN3_2),.clk(gclk));
	jdff dff_A_CMbgeeVU9_1(.dout(w_n614_0[1]),.din(w_dff_A_CMbgeeVU9_1),.clk(gclk));
	jdff dff_A_FdAIvIHk9_1(.dout(w_dff_A_CMbgeeVU9_1),.din(w_dff_A_FdAIvIHk9_1),.clk(gclk));
	jdff dff_A_xbIFYLSo9_1(.dout(w_dff_A_FdAIvIHk9_1),.din(w_dff_A_xbIFYLSo9_1),.clk(gclk));
	jdff dff_A_8wFEYYyP1_1(.dout(w_dff_A_xbIFYLSo9_1),.din(w_dff_A_8wFEYYyP1_1),.clk(gclk));
	jdff dff_A_Q1KQFFFf3_1(.dout(w_dff_A_8wFEYYyP1_1),.din(w_dff_A_Q1KQFFFf3_1),.clk(gclk));
	jdff dff_A_PxRhIh5L4_1(.dout(w_dff_A_Q1KQFFFf3_1),.din(w_dff_A_PxRhIh5L4_1),.clk(gclk));
	jdff dff_A_hdzvul4H2_1(.dout(w_dff_A_PxRhIh5L4_1),.din(w_dff_A_hdzvul4H2_1),.clk(gclk));
	jdff dff_A_LlBPJ9I44_2(.dout(w_n614_0[2]),.din(w_dff_A_LlBPJ9I44_2),.clk(gclk));
	jdff dff_A_Zjy67xRR6_2(.dout(w_dff_A_LlBPJ9I44_2),.din(w_dff_A_Zjy67xRR6_2),.clk(gclk));
	jdff dff_A_NOPBrzRH5_2(.dout(w_dff_A_Zjy67xRR6_2),.din(w_dff_A_NOPBrzRH5_2),.clk(gclk));
	jdff dff_A_mf1f6WvQ6_2(.dout(w_dff_A_NOPBrzRH5_2),.din(w_dff_A_mf1f6WvQ6_2),.clk(gclk));
	jdff dff_A_DLFXdhd73_2(.dout(w_dff_A_mf1f6WvQ6_2),.din(w_dff_A_DLFXdhd73_2),.clk(gclk));
	jdff dff_A_1R9Si16O6_0(.dout(w_n613_1[0]),.din(w_dff_A_1R9Si16O6_0),.clk(gclk));
	jdff dff_A_obybAHqW1_0(.dout(w_dff_A_1R9Si16O6_0),.din(w_dff_A_obybAHqW1_0),.clk(gclk));
	jdff dff_A_Qc3xcAoD7_0(.dout(w_dff_A_obybAHqW1_0),.din(w_dff_A_Qc3xcAoD7_0),.clk(gclk));
	jdff dff_A_FXKyyztp3_0(.dout(w_dff_A_Qc3xcAoD7_0),.din(w_dff_A_FXKyyztp3_0),.clk(gclk));
	jdff dff_A_3uKSBR5i7_0(.dout(w_dff_A_FXKyyztp3_0),.din(w_dff_A_3uKSBR5i7_0),.clk(gclk));
	jdff dff_A_sWTMSEHn0_0(.dout(w_dff_A_3uKSBR5i7_0),.din(w_dff_A_sWTMSEHn0_0),.clk(gclk));
	jdff dff_A_12WjBE4m9_0(.dout(w_dff_A_sWTMSEHn0_0),.din(w_dff_A_12WjBE4m9_0),.clk(gclk));
	jdff dff_A_qYB9Dq1x9_0(.dout(w_dff_A_12WjBE4m9_0),.din(w_dff_A_qYB9Dq1x9_0),.clk(gclk));
	jdff dff_A_GWni51SR5_0(.dout(w_dff_A_qYB9Dq1x9_0),.din(w_dff_A_GWni51SR5_0),.clk(gclk));
	jdff dff_A_UlhBziJO7_0(.dout(w_dff_A_GWni51SR5_0),.din(w_dff_A_UlhBziJO7_0),.clk(gclk));
	jdff dff_A_rTeRCFc31_0(.dout(w_dff_A_UlhBziJO7_0),.din(w_dff_A_rTeRCFc31_0),.clk(gclk));
	jdff dff_A_IvWnj4Wv1_0(.dout(w_dff_A_rTeRCFc31_0),.din(w_dff_A_IvWnj4Wv1_0),.clk(gclk));
	jdff dff_A_AqgmJPPZ1_0(.dout(w_dff_A_IvWnj4Wv1_0),.din(w_dff_A_AqgmJPPZ1_0),.clk(gclk));
	jdff dff_A_wfZHBpMz4_0(.dout(w_dff_A_AqgmJPPZ1_0),.din(w_dff_A_wfZHBpMz4_0),.clk(gclk));
	jdff dff_A_0xhGggqU0_1(.dout(w_n613_1[1]),.din(w_dff_A_0xhGggqU0_1),.clk(gclk));
	jdff dff_A_QefcfXOk7_1(.dout(w_dff_A_0xhGggqU0_1),.din(w_dff_A_QefcfXOk7_1),.clk(gclk));
	jdff dff_A_4NiS6VyX1_1(.dout(w_dff_A_QefcfXOk7_1),.din(w_dff_A_4NiS6VyX1_1),.clk(gclk));
	jdff dff_A_FRc0Ilhy3_1(.dout(w_dff_A_4NiS6VyX1_1),.din(w_dff_A_FRc0Ilhy3_1),.clk(gclk));
	jdff dff_A_3wM92rCX6_1(.dout(w_dff_A_FRc0Ilhy3_1),.din(w_dff_A_3wM92rCX6_1),.clk(gclk));
	jdff dff_A_IGQnP4ks6_1(.dout(w_dff_A_3wM92rCX6_1),.din(w_dff_A_IGQnP4ks6_1),.clk(gclk));
	jdff dff_A_nVb6Ejce5_1(.dout(w_dff_A_IGQnP4ks6_1),.din(w_dff_A_nVb6Ejce5_1),.clk(gclk));
	jdff dff_A_tppcESnG0_1(.dout(w_dff_A_nVb6Ejce5_1),.din(w_dff_A_tppcESnG0_1),.clk(gclk));
	jdff dff_A_kEuUguBW8_1(.dout(w_dff_A_tppcESnG0_1),.din(w_dff_A_kEuUguBW8_1),.clk(gclk));
	jdff dff_A_BIZ6vh7c2_1(.dout(w_dff_A_kEuUguBW8_1),.din(w_dff_A_BIZ6vh7c2_1),.clk(gclk));
	jdff dff_A_4HbW5Xy46_1(.dout(w_dff_A_BIZ6vh7c2_1),.din(w_dff_A_4HbW5Xy46_1),.clk(gclk));
	jdff dff_A_A2BL1Dqj5_1(.dout(w_dff_A_4HbW5Xy46_1),.din(w_dff_A_A2BL1Dqj5_1),.clk(gclk));
	jdff dff_A_8rU6N7RT9_1(.dout(w_dff_A_A2BL1Dqj5_1),.din(w_dff_A_8rU6N7RT9_1),.clk(gclk));
	jdff dff_A_MagKJvnV4_1(.dout(w_dff_A_8rU6N7RT9_1),.din(w_dff_A_MagKJvnV4_1),.clk(gclk));
	jdff dff_A_3dAvlS0C4_1(.dout(w_n613_0[1]),.din(w_dff_A_3dAvlS0C4_1),.clk(gclk));
	jdff dff_A_LDI5uEvl8_1(.dout(w_dff_A_3dAvlS0C4_1),.din(w_dff_A_LDI5uEvl8_1),.clk(gclk));
	jdff dff_A_wgx6Rqqe4_1(.dout(w_dff_A_LDI5uEvl8_1),.din(w_dff_A_wgx6Rqqe4_1),.clk(gclk));
	jdff dff_A_yL92aNsz9_1(.dout(w_dff_A_wgx6Rqqe4_1),.din(w_dff_A_yL92aNsz9_1),.clk(gclk));
	jdff dff_A_GTI0iPQO3_1(.dout(w_dff_A_yL92aNsz9_1),.din(w_dff_A_GTI0iPQO3_1),.clk(gclk));
	jdff dff_A_FjQWOwTT2_1(.dout(w_dff_A_GTI0iPQO3_1),.din(w_dff_A_FjQWOwTT2_1),.clk(gclk));
	jdff dff_A_uRAYGopk5_1(.dout(w_dff_A_FjQWOwTT2_1),.din(w_dff_A_uRAYGopk5_1),.clk(gclk));
	jdff dff_A_WZu9qbWm8_1(.dout(w_dff_A_uRAYGopk5_1),.din(w_dff_A_WZu9qbWm8_1),.clk(gclk));
	jdff dff_A_8dtSbyEy9_1(.dout(w_dff_A_WZu9qbWm8_1),.din(w_dff_A_8dtSbyEy9_1),.clk(gclk));
	jdff dff_A_WSlqBq2Q4_1(.dout(w_dff_A_8dtSbyEy9_1),.din(w_dff_A_WSlqBq2Q4_1),.clk(gclk));
	jdff dff_A_ZThLgVBk1_1(.dout(w_dff_A_WSlqBq2Q4_1),.din(w_dff_A_ZThLgVBk1_1),.clk(gclk));
	jdff dff_A_gLfYp3ZM8_1(.dout(w_dff_A_ZThLgVBk1_1),.din(w_dff_A_gLfYp3ZM8_1),.clk(gclk));
	jdff dff_A_pdliC2tE7_1(.dout(w_dff_A_gLfYp3ZM8_1),.din(w_dff_A_pdliC2tE7_1),.clk(gclk));
	jdff dff_A_oKM9GWo78_1(.dout(w_dff_A_pdliC2tE7_1),.din(w_dff_A_oKM9GWo78_1),.clk(gclk));
	jdff dff_A_PZ0LGSYx0_1(.dout(w_dff_A_oKM9GWo78_1),.din(w_dff_A_PZ0LGSYx0_1),.clk(gclk));
	jdff dff_A_Oglos4Ku8_2(.dout(w_n613_0[2]),.din(w_dff_A_Oglos4Ku8_2),.clk(gclk));
	jdff dff_A_Ya9hip4R8_2(.dout(w_dff_A_Oglos4Ku8_2),.din(w_dff_A_Ya9hip4R8_2),.clk(gclk));
	jdff dff_A_d0Thoz854_2(.dout(w_dff_A_Ya9hip4R8_2),.din(w_dff_A_d0Thoz854_2),.clk(gclk));
	jdff dff_A_QrPAXaBb6_2(.dout(w_dff_A_d0Thoz854_2),.din(w_dff_A_QrPAXaBb6_2),.clk(gclk));
	jdff dff_A_EmCbQ7yN5_2(.dout(w_dff_A_QrPAXaBb6_2),.din(w_dff_A_EmCbQ7yN5_2),.clk(gclk));
	jdff dff_A_i3JSTl7Z2_2(.dout(w_dff_A_EmCbQ7yN5_2),.din(w_dff_A_i3JSTl7Z2_2),.clk(gclk));
	jdff dff_A_H7XOka0E0_2(.dout(w_dff_A_i3JSTl7Z2_2),.din(w_dff_A_H7XOka0E0_2),.clk(gclk));
	jdff dff_A_ECridoI04_2(.dout(w_dff_A_H7XOka0E0_2),.din(w_dff_A_ECridoI04_2),.clk(gclk));
	jdff dff_A_lrCOda6n4_2(.dout(w_dff_A_ECridoI04_2),.din(w_dff_A_lrCOda6n4_2),.clk(gclk));
	jdff dff_A_CHTE9K1c1_2(.dout(w_dff_A_lrCOda6n4_2),.din(w_dff_A_CHTE9K1c1_2),.clk(gclk));
	jdff dff_A_GgC3TkUe9_2(.dout(w_dff_A_CHTE9K1c1_2),.din(w_dff_A_GgC3TkUe9_2),.clk(gclk));
	jdff dff_A_u9yvO9bL3_2(.dout(w_dff_A_GgC3TkUe9_2),.din(w_dff_A_u9yvO9bL3_2),.clk(gclk));
	jdff dff_A_nsfrGHtl6_2(.dout(w_dff_A_u9yvO9bL3_2),.din(w_dff_A_nsfrGHtl6_2),.clk(gclk));
	jdff dff_A_JxrKfOgy3_2(.dout(w_dff_A_nsfrGHtl6_2),.din(w_dff_A_JxrKfOgy3_2),.clk(gclk));
	jdff dff_A_KFHMGHX69_2(.dout(w_dff_A_JxrKfOgy3_2),.din(w_dff_A_KFHMGHX69_2),.clk(gclk));
	jdff dff_A_PI2cxiYp5_2(.dout(w_dff_A_KFHMGHX69_2),.din(w_dff_A_PI2cxiYp5_2),.clk(gclk));
	jdff dff_A_4pvAQzxU1_2(.dout(w_dff_A_PI2cxiYp5_2),.din(w_dff_A_4pvAQzxU1_2),.clk(gclk));
	jdff dff_B_1Lv68ur21_3(.din(n613),.dout(w_dff_B_1Lv68ur21_3),.clk(gclk));
	jdff dff_A_JwdWPdBz1_1(.dout(w_G45_0[1]),.din(w_dff_A_JwdWPdBz1_1),.clk(gclk));
	jdff dff_A_ix5lpmXU0_1(.dout(w_dff_A_JwdWPdBz1_1),.din(w_dff_A_ix5lpmXU0_1),.clk(gclk));
	jdff dff_A_WlqT3q5V3_1(.dout(w_dff_A_ix5lpmXU0_1),.din(w_dff_A_WlqT3q5V3_1),.clk(gclk));
	jdff dff_A_QqWgiOB68_0(.dout(w_n151_2[0]),.din(w_dff_A_QqWgiOB68_0),.clk(gclk));
	jdff dff_A_d48y1CTs7_2(.dout(w_n151_2[2]),.din(w_dff_A_d48y1CTs7_2),.clk(gclk));
	jdff dff_A_shuBNnAO4_2(.dout(w_dff_A_d48y1CTs7_2),.din(w_dff_A_shuBNnAO4_2),.clk(gclk));
	jdff dff_A_DjzwFZwv6_0(.dout(w_G20_5[0]),.din(w_dff_A_DjzwFZwv6_0),.clk(gclk));
	jdff dff_A_BqhNtu9n3_2(.dout(w_n142_0[2]),.din(w_dff_A_BqhNtu9n3_2),.clk(gclk));
	jdff dff_A_5LV0ZNYi7_0(.dout(w_G1_1[0]),.din(w_dff_A_5LV0ZNYi7_0),.clk(gclk));
	jdff dff_A_yWAHEjrD4_0(.dout(w_dff_A_5LV0ZNYi7_0),.din(w_dff_A_yWAHEjrD4_0),.clk(gclk));
	jdff dff_A_C0Y1nxKr5_0(.dout(w_n604_2[0]),.din(w_dff_A_C0Y1nxKr5_0),.clk(gclk));
	jdff dff_A_N8uUEA564_0(.dout(w_dff_A_C0Y1nxKr5_0),.din(w_dff_A_N8uUEA564_0),.clk(gclk));
	jdff dff_A_FC1iz72s0_0(.dout(w_dff_A_N8uUEA564_0),.din(w_dff_A_FC1iz72s0_0),.clk(gclk));
	jdff dff_A_mYU0z91q4_0(.dout(w_dff_A_FC1iz72s0_0),.din(w_dff_A_mYU0z91q4_0),.clk(gclk));
	jdff dff_A_xgDM7dwZ7_0(.dout(w_dff_A_mYU0z91q4_0),.din(w_dff_A_xgDM7dwZ7_0),.clk(gclk));
	jdff dff_A_PWK2Wi2W5_0(.dout(w_dff_A_xgDM7dwZ7_0),.din(w_dff_A_PWK2Wi2W5_0),.clk(gclk));
	jdff dff_A_OcU4o0PY9_0(.dout(w_dff_A_PWK2Wi2W5_0),.din(w_dff_A_OcU4o0PY9_0),.clk(gclk));
	jdff dff_A_6iuFEKGn1_0(.dout(w_dff_A_OcU4o0PY9_0),.din(w_dff_A_6iuFEKGn1_0),.clk(gclk));
	jdff dff_A_fa7POqnd3_0(.dout(w_dff_A_6iuFEKGn1_0),.din(w_dff_A_fa7POqnd3_0),.clk(gclk));
	jdff dff_A_eA3Hz6G88_0(.dout(w_dff_A_fa7POqnd3_0),.din(w_dff_A_eA3Hz6G88_0),.clk(gclk));
	jdff dff_A_QNi4j1dS1_0(.dout(w_dff_A_eA3Hz6G88_0),.din(w_dff_A_QNi4j1dS1_0),.clk(gclk));
	jdff dff_A_RJcwQIOp0_0(.dout(w_dff_A_QNi4j1dS1_0),.din(w_dff_A_RJcwQIOp0_0),.clk(gclk));
	jdff dff_A_7FQombol2_0(.dout(w_dff_A_RJcwQIOp0_0),.din(w_dff_A_7FQombol2_0),.clk(gclk));
	jdff dff_A_R9Tb3AaW0_0(.dout(w_dff_A_7FQombol2_0),.din(w_dff_A_R9Tb3AaW0_0),.clk(gclk));
	jdff dff_A_WIoQs0wk6_0(.dout(w_n604_0[0]),.din(w_dff_A_WIoQs0wk6_0),.clk(gclk));
	jdff dff_A_PjYVHhuR2_0(.dout(w_dff_A_WIoQs0wk6_0),.din(w_dff_A_PjYVHhuR2_0),.clk(gclk));
	jdff dff_A_fWHv26iz4_0(.dout(w_dff_A_PjYVHhuR2_0),.din(w_dff_A_fWHv26iz4_0),.clk(gclk));
	jdff dff_A_99Pg9m6g2_0(.dout(w_dff_A_fWHv26iz4_0),.din(w_dff_A_99Pg9m6g2_0),.clk(gclk));
	jdff dff_A_AHJMJUka6_0(.dout(w_dff_A_99Pg9m6g2_0),.din(w_dff_A_AHJMJUka6_0),.clk(gclk));
	jdff dff_A_zvrsVdck8_0(.dout(w_dff_A_AHJMJUka6_0),.din(w_dff_A_zvrsVdck8_0),.clk(gclk));
	jdff dff_A_NZyLzJFy7_0(.dout(w_dff_A_zvrsVdck8_0),.din(w_dff_A_NZyLzJFy7_0),.clk(gclk));
	jdff dff_A_tviPC0cg8_0(.dout(w_dff_A_NZyLzJFy7_0),.din(w_dff_A_tviPC0cg8_0),.clk(gclk));
	jdff dff_A_gVbHCnsA3_0(.dout(w_dff_A_tviPC0cg8_0),.din(w_dff_A_gVbHCnsA3_0),.clk(gclk));
	jdff dff_A_egO8b8PU9_0(.dout(w_dff_A_gVbHCnsA3_0),.din(w_dff_A_egO8b8PU9_0),.clk(gclk));
	jdff dff_A_bhftzGJH2_0(.dout(w_dff_A_egO8b8PU9_0),.din(w_dff_A_bhftzGJH2_0),.clk(gclk));
	jdff dff_A_rTq4C2s82_0(.dout(w_dff_A_bhftzGJH2_0),.din(w_dff_A_rTq4C2s82_0),.clk(gclk));
	jdff dff_A_QgXvcrKk2_0(.dout(w_dff_A_rTq4C2s82_0),.din(w_dff_A_QgXvcrKk2_0),.clk(gclk));
	jdff dff_A_wO4aJOgl9_0(.dout(w_dff_A_QgXvcrKk2_0),.din(w_dff_A_wO4aJOgl9_0),.clk(gclk));
	jdff dff_A_DSBhHVGb0_2(.dout(w_n604_0[2]),.din(w_dff_A_DSBhHVGb0_2),.clk(gclk));
	jdff dff_A_sOs4v8DJ5_2(.dout(w_dff_A_DSBhHVGb0_2),.din(w_dff_A_sOs4v8DJ5_2),.clk(gclk));
	jdff dff_A_BUFbwBqi6_2(.dout(w_dff_A_sOs4v8DJ5_2),.din(w_dff_A_BUFbwBqi6_2),.clk(gclk));
	jdff dff_A_kEcJPfP69_2(.dout(w_dff_A_BUFbwBqi6_2),.din(w_dff_A_kEcJPfP69_2),.clk(gclk));
	jdff dff_A_vMKfo7I57_2(.dout(w_dff_A_kEcJPfP69_2),.din(w_dff_A_vMKfo7I57_2),.clk(gclk));
	jdff dff_A_SsWESpZx2_2(.dout(w_dff_A_vMKfo7I57_2),.din(w_dff_A_SsWESpZx2_2),.clk(gclk));
	jdff dff_A_E0A4jplz8_2(.dout(w_dff_A_SsWESpZx2_2),.din(w_dff_A_E0A4jplz8_2),.clk(gclk));
	jdff dff_A_1ll4yG0V1_2(.dout(w_dff_A_E0A4jplz8_2),.din(w_dff_A_1ll4yG0V1_2),.clk(gclk));
	jdff dff_A_B3QQj4Ub4_2(.dout(w_dff_A_1ll4yG0V1_2),.din(w_dff_A_B3QQj4Ub4_2),.clk(gclk));
	jdff dff_A_qXc8K7HE9_2(.dout(w_dff_A_B3QQj4Ub4_2),.din(w_dff_A_qXc8K7HE9_2),.clk(gclk));
	jdff dff_A_kae52u6T9_2(.dout(w_dff_A_qXc8K7HE9_2),.din(w_dff_A_kae52u6T9_2),.clk(gclk));
	jdff dff_A_74MvuWDk0_2(.dout(w_dff_A_kae52u6T9_2),.din(w_dff_A_74MvuWDk0_2),.clk(gclk));
	jdff dff_A_ZTuxilk38_2(.dout(w_dff_A_74MvuWDk0_2),.din(w_dff_A_ZTuxilk38_2),.clk(gclk));
	jdff dff_A_qBD6oLY86_2(.dout(w_dff_A_ZTuxilk38_2),.din(w_dff_A_qBD6oLY86_2),.clk(gclk));
	jdff dff_A_kOpgo1hg4_2(.dout(w_dff_A_qBD6oLY86_2),.din(w_dff_A_kOpgo1hg4_2),.clk(gclk));
	jdff dff_A_WIx6MBO00_2(.dout(w_dff_A_kOpgo1hg4_2),.din(w_dff_A_WIx6MBO00_2),.clk(gclk));
	jdff dff_A_qgnPfh6H0_0(.dout(w_G13_2[0]),.din(w_dff_A_qgnPfh6H0_0),.clk(gclk));
	jdff dff_A_rJrIH5jY5_1(.dout(w_G1_2[1]),.din(w_dff_A_rJrIH5jY5_1),.clk(gclk));
	jdff dff_A_C3AB7ibC0_2(.dout(w_G1_0[2]),.din(w_dff_A_C3AB7ibC0_2),.clk(gclk));
	jdff dff_A_Q46LP6PO3_2(.dout(w_dff_A_C3AB7ibC0_2),.din(w_dff_A_Q46LP6PO3_2),.clk(gclk));
	jdff dff_A_G1WJMjkL0_2(.dout(w_dff_A_Q46LP6PO3_2),.din(w_dff_A_G1WJMjkL0_2),.clk(gclk));
	jdff dff_A_7986Ijkt6_2(.dout(w_dff_A_G1WJMjkL0_2),.din(w_dff_A_7986Ijkt6_2),.clk(gclk));
	jdff dff_A_5x6ZmtxS3_0(.dout(w_G20_6[0]),.din(w_dff_A_5x6ZmtxS3_0),.clk(gclk));
	jdff dff_A_7JrKyfu22_0(.dout(w_dff_A_5x6ZmtxS3_0),.din(w_dff_A_7JrKyfu22_0),.clk(gclk));
	jdff dff_A_Y8WSD0v91_2(.dout(w_G20_6[2]),.din(w_dff_A_Y8WSD0v91_2),.clk(gclk));
	jdff dff_A_smLdoHTq5_2(.dout(w_dff_A_Y8WSD0v91_2),.din(w_dff_A_smLdoHTq5_2),.clk(gclk));
	jdff dff_A_8uDIUc495_0(.dout(w_G20_1[0]),.din(w_dff_A_8uDIUc495_0),.clk(gclk));
	jdff dff_A_IRLX5wUz8_2(.dout(w_G20_0[2]),.din(w_dff_A_IRLX5wUz8_2),.clk(gclk));
	jdff dff_A_CHib6UZM2_1(.dout(w_n163_0[1]),.din(w_dff_A_CHib6UZM2_1),.clk(gclk));
	jdff dff_A_lI6RmWBc9_1(.dout(w_dff_A_CHib6UZM2_1),.din(w_dff_A_lI6RmWBc9_1),.clk(gclk));
	jdff dff_A_I7yF9JIC0_1(.dout(w_dff_A_lI6RmWBc9_1),.din(w_dff_A_I7yF9JIC0_1),.clk(gclk));
	jdff dff_A_IEut3ixz5_1(.dout(w_dff_A_I7yF9JIC0_1),.din(w_dff_A_IEut3ixz5_1),.clk(gclk));
	jdff dff_A_0sJdbqaP8_1(.dout(w_dff_A_IEut3ixz5_1),.din(w_dff_A_0sJdbqaP8_1),.clk(gclk));
	jdff dff_A_jeojB7IL6_1(.dout(w_dff_A_0sJdbqaP8_1),.din(w_dff_A_jeojB7IL6_1),.clk(gclk));
	jdff dff_A_sIpatig60_1(.dout(w_dff_A_jeojB7IL6_1),.din(w_dff_A_sIpatig60_1),.clk(gclk));
	jdff dff_A_gMBPaD9G2_1(.dout(w_dff_A_sIpatig60_1),.din(w_dff_A_gMBPaD9G2_1),.clk(gclk));
	jdff dff_A_O2bBxmb51_1(.dout(w_dff_A_gMBPaD9G2_1),.din(w_dff_A_O2bBxmb51_1),.clk(gclk));
	jdff dff_A_uoPZYNJ70_1(.dout(w_dff_A_O2bBxmb51_1),.din(w_dff_A_uoPZYNJ70_1),.clk(gclk));
	jdff dff_A_PB3oHri44_1(.dout(w_dff_A_uoPZYNJ70_1),.din(w_dff_A_PB3oHri44_1),.clk(gclk));
	jdff dff_A_NdEaSX8R9_2(.dout(w_n163_0[2]),.din(w_dff_A_NdEaSX8R9_2),.clk(gclk));
	jdff dff_A_7HilQhhT0_2(.dout(w_dff_A_NdEaSX8R9_2),.din(w_dff_A_7HilQhhT0_2),.clk(gclk));
	jdff dff_A_dvfHxH6U7_2(.dout(w_dff_A_lQD0TU6M9_0),.din(w_dff_A_dvfHxH6U7_2),.clk(gclk));
	jdff dff_A_lQD0TU6M9_0(.dout(w_dff_A_FXipZlDr0_0),.din(w_dff_A_lQD0TU6M9_0),.clk(gclk));
	jdff dff_A_FXipZlDr0_0(.dout(w_dff_A_ViIZUB9l5_0),.din(w_dff_A_FXipZlDr0_0),.clk(gclk));
	jdff dff_A_ViIZUB9l5_0(.dout(w_dff_A_2akBU97p0_0),.din(w_dff_A_ViIZUB9l5_0),.clk(gclk));
	jdff dff_A_2akBU97p0_0(.dout(w_dff_A_yvX93bRn9_0),.din(w_dff_A_2akBU97p0_0),.clk(gclk));
	jdff dff_A_yvX93bRn9_0(.dout(w_dff_A_mvXyFqv12_0),.din(w_dff_A_yvX93bRn9_0),.clk(gclk));
	jdff dff_A_mvXyFqv12_0(.dout(w_dff_A_2pL9S8xB2_0),.din(w_dff_A_mvXyFqv12_0),.clk(gclk));
	jdff dff_A_2pL9S8xB2_0(.dout(w_dff_A_vrS3NHSZ1_0),.din(w_dff_A_2pL9S8xB2_0),.clk(gclk));
	jdff dff_A_vrS3NHSZ1_0(.dout(w_dff_A_sVWFZwx82_0),.din(w_dff_A_vrS3NHSZ1_0),.clk(gclk));
	jdff dff_A_sVWFZwx82_0(.dout(w_dff_A_SCcE3mM90_0),.din(w_dff_A_sVWFZwx82_0),.clk(gclk));
	jdff dff_A_SCcE3mM90_0(.dout(w_dff_A_ZxMMe4fR3_0),.din(w_dff_A_SCcE3mM90_0),.clk(gclk));
	jdff dff_A_ZxMMe4fR3_0(.dout(w_dff_A_0WhpOIuC2_0),.din(w_dff_A_ZxMMe4fR3_0),.clk(gclk));
	jdff dff_A_0WhpOIuC2_0(.dout(w_dff_A_m1CnoXj26_0),.din(w_dff_A_0WhpOIuC2_0),.clk(gclk));
	jdff dff_A_m1CnoXj26_0(.dout(w_dff_A_g5H1H4El9_0),.din(w_dff_A_m1CnoXj26_0),.clk(gclk));
	jdff dff_A_g5H1H4El9_0(.dout(w_dff_A_yfPBnnf84_0),.din(w_dff_A_g5H1H4El9_0),.clk(gclk));
	jdff dff_A_yfPBnnf84_0(.dout(w_dff_A_ufkPlikO5_0),.din(w_dff_A_yfPBnnf84_0),.clk(gclk));
	jdff dff_A_ufkPlikO5_0(.dout(w_dff_A_RLJVZK2G8_0),.din(w_dff_A_ufkPlikO5_0),.clk(gclk));
	jdff dff_A_RLJVZK2G8_0(.dout(w_dff_A_BaOeCvDH3_0),.din(w_dff_A_RLJVZK2G8_0),.clk(gclk));
	jdff dff_A_BaOeCvDH3_0(.dout(w_dff_A_OKumeTud6_0),.din(w_dff_A_BaOeCvDH3_0),.clk(gclk));
	jdff dff_A_OKumeTud6_0(.dout(w_dff_A_YlHksyqL1_0),.din(w_dff_A_OKumeTud6_0),.clk(gclk));
	jdff dff_A_YlHksyqL1_0(.dout(w_dff_A_JwsvjUze0_0),.din(w_dff_A_YlHksyqL1_0),.clk(gclk));
	jdff dff_A_JwsvjUze0_0(.dout(w_dff_A_8VYXWAyJ9_0),.din(w_dff_A_JwsvjUze0_0),.clk(gclk));
	jdff dff_A_8VYXWAyJ9_0(.dout(w_dff_A_n9C3awQk2_0),.din(w_dff_A_8VYXWAyJ9_0),.clk(gclk));
	jdff dff_A_n9C3awQk2_0(.dout(w_dff_A_YkZB4vyM3_0),.din(w_dff_A_n9C3awQk2_0),.clk(gclk));
	jdff dff_A_YkZB4vyM3_0(.dout(w_dff_A_I7A3yWWS5_0),.din(w_dff_A_YkZB4vyM3_0),.clk(gclk));
	jdff dff_A_I7A3yWWS5_0(.dout(w_dff_A_wCCyFw6L0_0),.din(w_dff_A_I7A3yWWS5_0),.clk(gclk));
	jdff dff_A_wCCyFw6L0_0(.dout(G353),.din(w_dff_A_wCCyFw6L0_0),.clk(gclk));
	jdff dff_A_jteEvgx45_1(.dout(w_dff_A_X67LN1Bf4_0),.din(w_dff_A_jteEvgx45_1),.clk(gclk));
	jdff dff_A_X67LN1Bf4_0(.dout(w_dff_A_jMdOBbu30_0),.din(w_dff_A_X67LN1Bf4_0),.clk(gclk));
	jdff dff_A_jMdOBbu30_0(.dout(w_dff_A_XJfZkCo89_0),.din(w_dff_A_jMdOBbu30_0),.clk(gclk));
	jdff dff_A_XJfZkCo89_0(.dout(w_dff_A_WlyUcA2o3_0),.din(w_dff_A_XJfZkCo89_0),.clk(gclk));
	jdff dff_A_WlyUcA2o3_0(.dout(w_dff_A_ZLuIMkLz5_0),.din(w_dff_A_WlyUcA2o3_0),.clk(gclk));
	jdff dff_A_ZLuIMkLz5_0(.dout(w_dff_A_IQZCiqyM2_0),.din(w_dff_A_ZLuIMkLz5_0),.clk(gclk));
	jdff dff_A_IQZCiqyM2_0(.dout(w_dff_A_7Bxq12E40_0),.din(w_dff_A_IQZCiqyM2_0),.clk(gclk));
	jdff dff_A_7Bxq12E40_0(.dout(w_dff_A_Oh6VSvYU0_0),.din(w_dff_A_7Bxq12E40_0),.clk(gclk));
	jdff dff_A_Oh6VSvYU0_0(.dout(w_dff_A_pgFRIrOs0_0),.din(w_dff_A_Oh6VSvYU0_0),.clk(gclk));
	jdff dff_A_pgFRIrOs0_0(.dout(w_dff_A_70xqkUAe6_0),.din(w_dff_A_pgFRIrOs0_0),.clk(gclk));
	jdff dff_A_70xqkUAe6_0(.dout(w_dff_A_3p3GpOYP7_0),.din(w_dff_A_70xqkUAe6_0),.clk(gclk));
	jdff dff_A_3p3GpOYP7_0(.dout(w_dff_A_54q4HlXO8_0),.din(w_dff_A_3p3GpOYP7_0),.clk(gclk));
	jdff dff_A_54q4HlXO8_0(.dout(w_dff_A_wkE7jZiQ1_0),.din(w_dff_A_54q4HlXO8_0),.clk(gclk));
	jdff dff_A_wkE7jZiQ1_0(.dout(w_dff_A_UioTpEI78_0),.din(w_dff_A_wkE7jZiQ1_0),.clk(gclk));
	jdff dff_A_UioTpEI78_0(.dout(w_dff_A_g8xwiyng7_0),.din(w_dff_A_UioTpEI78_0),.clk(gclk));
	jdff dff_A_g8xwiyng7_0(.dout(w_dff_A_BKhw5jh21_0),.din(w_dff_A_g8xwiyng7_0),.clk(gclk));
	jdff dff_A_BKhw5jh21_0(.dout(w_dff_A_VetyY1zY4_0),.din(w_dff_A_BKhw5jh21_0),.clk(gclk));
	jdff dff_A_VetyY1zY4_0(.dout(w_dff_A_eHSwebds9_0),.din(w_dff_A_VetyY1zY4_0),.clk(gclk));
	jdff dff_A_eHSwebds9_0(.dout(w_dff_A_2w49CTng6_0),.din(w_dff_A_eHSwebds9_0),.clk(gclk));
	jdff dff_A_2w49CTng6_0(.dout(w_dff_A_7X90HefZ6_0),.din(w_dff_A_2w49CTng6_0),.clk(gclk));
	jdff dff_A_7X90HefZ6_0(.dout(w_dff_A_0GD5q4Eq8_0),.din(w_dff_A_7X90HefZ6_0),.clk(gclk));
	jdff dff_A_0GD5q4Eq8_0(.dout(w_dff_A_nNCInwRr4_0),.din(w_dff_A_0GD5q4Eq8_0),.clk(gclk));
	jdff dff_A_nNCInwRr4_0(.dout(w_dff_A_f78lEgGc0_0),.din(w_dff_A_nNCInwRr4_0),.clk(gclk));
	jdff dff_A_f78lEgGc0_0(.dout(w_dff_A_MAFvvJ157_0),.din(w_dff_A_f78lEgGc0_0),.clk(gclk));
	jdff dff_A_MAFvvJ157_0(.dout(w_dff_A_yqhI50uz1_0),.din(w_dff_A_MAFvvJ157_0),.clk(gclk));
	jdff dff_A_yqhI50uz1_0(.dout(w_dff_A_Hf1wkeAO0_0),.din(w_dff_A_yqhI50uz1_0),.clk(gclk));
	jdff dff_A_Hf1wkeAO0_0(.dout(w_dff_A_qOUGhVbK5_0),.din(w_dff_A_Hf1wkeAO0_0),.clk(gclk));
	jdff dff_A_qOUGhVbK5_0(.dout(G355),.din(w_dff_A_qOUGhVbK5_0),.clk(gclk));
	jdff dff_A_JOEDEGQA0_2(.dout(w_dff_A_rYz2HKC41_0),.din(w_dff_A_JOEDEGQA0_2),.clk(gclk));
	jdff dff_A_rYz2HKC41_0(.dout(w_dff_A_1YTb7ARq9_0),.din(w_dff_A_rYz2HKC41_0),.clk(gclk));
	jdff dff_A_1YTb7ARq9_0(.dout(w_dff_A_5O2kPZzG2_0),.din(w_dff_A_1YTb7ARq9_0),.clk(gclk));
	jdff dff_A_5O2kPZzG2_0(.dout(w_dff_A_APvWXbhT4_0),.din(w_dff_A_5O2kPZzG2_0),.clk(gclk));
	jdff dff_A_APvWXbhT4_0(.dout(w_dff_A_qO3YfwMZ8_0),.din(w_dff_A_APvWXbhT4_0),.clk(gclk));
	jdff dff_A_qO3YfwMZ8_0(.dout(w_dff_A_4lztVejE9_0),.din(w_dff_A_qO3YfwMZ8_0),.clk(gclk));
	jdff dff_A_4lztVejE9_0(.dout(w_dff_A_l0UyLx583_0),.din(w_dff_A_4lztVejE9_0),.clk(gclk));
	jdff dff_A_l0UyLx583_0(.dout(w_dff_A_v8k0iaiU6_0),.din(w_dff_A_l0UyLx583_0),.clk(gclk));
	jdff dff_A_v8k0iaiU6_0(.dout(w_dff_A_DihRufN79_0),.din(w_dff_A_v8k0iaiU6_0),.clk(gclk));
	jdff dff_A_DihRufN79_0(.dout(w_dff_A_lIXyRskE8_0),.din(w_dff_A_DihRufN79_0),.clk(gclk));
	jdff dff_A_lIXyRskE8_0(.dout(w_dff_A_bPbxL5fV0_0),.din(w_dff_A_lIXyRskE8_0),.clk(gclk));
	jdff dff_A_bPbxL5fV0_0(.dout(w_dff_A_mmRqkyfv9_0),.din(w_dff_A_bPbxL5fV0_0),.clk(gclk));
	jdff dff_A_mmRqkyfv9_0(.dout(w_dff_A_cZ5LdLCG5_0),.din(w_dff_A_mmRqkyfv9_0),.clk(gclk));
	jdff dff_A_cZ5LdLCG5_0(.dout(w_dff_A_Vxg88BlP0_0),.din(w_dff_A_cZ5LdLCG5_0),.clk(gclk));
	jdff dff_A_Vxg88BlP0_0(.dout(w_dff_A_LefBbsUQ1_0),.din(w_dff_A_Vxg88BlP0_0),.clk(gclk));
	jdff dff_A_LefBbsUQ1_0(.dout(w_dff_A_hDdd8gJf2_0),.din(w_dff_A_LefBbsUQ1_0),.clk(gclk));
	jdff dff_A_hDdd8gJf2_0(.dout(w_dff_A_hB0ERWBs1_0),.din(w_dff_A_hDdd8gJf2_0),.clk(gclk));
	jdff dff_A_hB0ERWBs1_0(.dout(w_dff_A_KG9hLs979_0),.din(w_dff_A_hB0ERWBs1_0),.clk(gclk));
	jdff dff_A_KG9hLs979_0(.dout(w_dff_A_eLKBOjPD9_0),.din(w_dff_A_KG9hLs979_0),.clk(gclk));
	jdff dff_A_eLKBOjPD9_0(.dout(w_dff_A_zC8URcQ80_0),.din(w_dff_A_eLKBOjPD9_0),.clk(gclk));
	jdff dff_A_zC8URcQ80_0(.dout(w_dff_A_NqXqbQbd6_0),.din(w_dff_A_zC8URcQ80_0),.clk(gclk));
	jdff dff_A_NqXqbQbd6_0(.dout(w_dff_A_G8WT6kR23_0),.din(w_dff_A_NqXqbQbd6_0),.clk(gclk));
	jdff dff_A_G8WT6kR23_0(.dout(G361),.din(w_dff_A_G8WT6kR23_0),.clk(gclk));
	jdff dff_A_IRozgalU2_2(.dout(w_dff_A_6EuHXGSU2_0),.din(w_dff_A_IRozgalU2_2),.clk(gclk));
	jdff dff_A_6EuHXGSU2_0(.dout(w_dff_A_jUpMeuZt8_0),.din(w_dff_A_6EuHXGSU2_0),.clk(gclk));
	jdff dff_A_jUpMeuZt8_0(.dout(w_dff_A_OhViaEMp3_0),.din(w_dff_A_jUpMeuZt8_0),.clk(gclk));
	jdff dff_A_OhViaEMp3_0(.dout(w_dff_A_jtHrDZij6_0),.din(w_dff_A_OhViaEMp3_0),.clk(gclk));
	jdff dff_A_jtHrDZij6_0(.dout(w_dff_A_NEi4l9kO4_0),.din(w_dff_A_jtHrDZij6_0),.clk(gclk));
	jdff dff_A_NEi4l9kO4_0(.dout(w_dff_A_KmcwJAqm2_0),.din(w_dff_A_NEi4l9kO4_0),.clk(gclk));
	jdff dff_A_KmcwJAqm2_0(.dout(w_dff_A_xkNIAmfP4_0),.din(w_dff_A_KmcwJAqm2_0),.clk(gclk));
	jdff dff_A_xkNIAmfP4_0(.dout(w_dff_A_AGjpLRWf3_0),.din(w_dff_A_xkNIAmfP4_0),.clk(gclk));
	jdff dff_A_AGjpLRWf3_0(.dout(w_dff_A_yNoHbPBA8_0),.din(w_dff_A_AGjpLRWf3_0),.clk(gclk));
	jdff dff_A_yNoHbPBA8_0(.dout(w_dff_A_NhLXKGeP9_0),.din(w_dff_A_yNoHbPBA8_0),.clk(gclk));
	jdff dff_A_NhLXKGeP9_0(.dout(w_dff_A_SgFdvEgU6_0),.din(w_dff_A_NhLXKGeP9_0),.clk(gclk));
	jdff dff_A_SgFdvEgU6_0(.dout(w_dff_A_lLYoPJk01_0),.din(w_dff_A_SgFdvEgU6_0),.clk(gclk));
	jdff dff_A_lLYoPJk01_0(.dout(w_dff_A_t3l7K1vH2_0),.din(w_dff_A_lLYoPJk01_0),.clk(gclk));
	jdff dff_A_t3l7K1vH2_0(.dout(w_dff_A_ygHS9l900_0),.din(w_dff_A_t3l7K1vH2_0),.clk(gclk));
	jdff dff_A_ygHS9l900_0(.dout(w_dff_A_PCmF4Sys9_0),.din(w_dff_A_ygHS9l900_0),.clk(gclk));
	jdff dff_A_PCmF4Sys9_0(.dout(w_dff_A_uRItRhdz3_0),.din(w_dff_A_PCmF4Sys9_0),.clk(gclk));
	jdff dff_A_uRItRhdz3_0(.dout(w_dff_A_16p9pGa21_0),.din(w_dff_A_uRItRhdz3_0),.clk(gclk));
	jdff dff_A_16p9pGa21_0(.dout(w_dff_A_BtAV4KZf3_0),.din(w_dff_A_16p9pGa21_0),.clk(gclk));
	jdff dff_A_BtAV4KZf3_0(.dout(w_dff_A_bajZLfm07_0),.din(w_dff_A_BtAV4KZf3_0),.clk(gclk));
	jdff dff_A_bajZLfm07_0(.dout(w_dff_A_fRu6qHu15_0),.din(w_dff_A_bajZLfm07_0),.clk(gclk));
	jdff dff_A_fRu6qHu15_0(.dout(w_dff_A_OQp68ksv5_0),.din(w_dff_A_fRu6qHu15_0),.clk(gclk));
	jdff dff_A_OQp68ksv5_0(.dout(w_dff_A_z1k4NQFU1_0),.din(w_dff_A_OQp68ksv5_0),.clk(gclk));
	jdff dff_A_z1k4NQFU1_0(.dout(w_dff_A_Kpjv5gdY0_0),.din(w_dff_A_z1k4NQFU1_0),.clk(gclk));
	jdff dff_A_Kpjv5gdY0_0(.dout(w_dff_A_nQIK8Zit8_0),.din(w_dff_A_Kpjv5gdY0_0),.clk(gclk));
	jdff dff_A_nQIK8Zit8_0(.dout(w_dff_A_T0ChLpHK4_0),.din(w_dff_A_nQIK8Zit8_0),.clk(gclk));
	jdff dff_A_T0ChLpHK4_0(.dout(G358),.din(w_dff_A_T0ChLpHK4_0),.clk(gclk));
	jdff dff_A_rJIYourm4_2(.dout(w_dff_A_TOumBzkK2_0),.din(w_dff_A_rJIYourm4_2),.clk(gclk));
	jdff dff_A_TOumBzkK2_0(.dout(w_dff_A_bjhIJXWY0_0),.din(w_dff_A_TOumBzkK2_0),.clk(gclk));
	jdff dff_A_bjhIJXWY0_0(.dout(w_dff_A_XpghVJi75_0),.din(w_dff_A_bjhIJXWY0_0),.clk(gclk));
	jdff dff_A_XpghVJi75_0(.dout(w_dff_A_u3iZTuj79_0),.din(w_dff_A_XpghVJi75_0),.clk(gclk));
	jdff dff_A_u3iZTuj79_0(.dout(w_dff_A_Lvb23Mf41_0),.din(w_dff_A_u3iZTuj79_0),.clk(gclk));
	jdff dff_A_Lvb23Mf41_0(.dout(w_dff_A_SRgK80nf5_0),.din(w_dff_A_Lvb23Mf41_0),.clk(gclk));
	jdff dff_A_SRgK80nf5_0(.dout(w_dff_A_SSh2RfLE9_0),.din(w_dff_A_SRgK80nf5_0),.clk(gclk));
	jdff dff_A_SSh2RfLE9_0(.dout(w_dff_A_6omLeoJL4_0),.din(w_dff_A_SSh2RfLE9_0),.clk(gclk));
	jdff dff_A_6omLeoJL4_0(.dout(w_dff_A_UqBhDRfT9_0),.din(w_dff_A_6omLeoJL4_0),.clk(gclk));
	jdff dff_A_UqBhDRfT9_0(.dout(w_dff_A_ENrCIkFF9_0),.din(w_dff_A_UqBhDRfT9_0),.clk(gclk));
	jdff dff_A_ENrCIkFF9_0(.dout(w_dff_A_ptCoTQtI9_0),.din(w_dff_A_ENrCIkFF9_0),.clk(gclk));
	jdff dff_A_ptCoTQtI9_0(.dout(w_dff_A_A0GQ3z722_0),.din(w_dff_A_ptCoTQtI9_0),.clk(gclk));
	jdff dff_A_A0GQ3z722_0(.dout(w_dff_A_pDPzjMxa5_0),.din(w_dff_A_A0GQ3z722_0),.clk(gclk));
	jdff dff_A_pDPzjMxa5_0(.dout(w_dff_A_sUXIRc6K2_0),.din(w_dff_A_pDPzjMxa5_0),.clk(gclk));
	jdff dff_A_sUXIRc6K2_0(.dout(w_dff_A_xUBjtKW42_0),.din(w_dff_A_sUXIRc6K2_0),.clk(gclk));
	jdff dff_A_xUBjtKW42_0(.dout(w_dff_A_VVge2dm36_0),.din(w_dff_A_xUBjtKW42_0),.clk(gclk));
	jdff dff_A_VVge2dm36_0(.dout(w_dff_A_awm6kvCg6_0),.din(w_dff_A_VVge2dm36_0),.clk(gclk));
	jdff dff_A_awm6kvCg6_0(.dout(w_dff_A_CaLOVrzE3_0),.din(w_dff_A_awm6kvCg6_0),.clk(gclk));
	jdff dff_A_CaLOVrzE3_0(.dout(w_dff_A_lrij1AOu6_0),.din(w_dff_A_CaLOVrzE3_0),.clk(gclk));
	jdff dff_A_lrij1AOu6_0(.dout(w_dff_A_AUbvzYts2_0),.din(w_dff_A_lrij1AOu6_0),.clk(gclk));
	jdff dff_A_AUbvzYts2_0(.dout(w_dff_A_T1ZfaDTv1_0),.din(w_dff_A_AUbvzYts2_0),.clk(gclk));
	jdff dff_A_T1ZfaDTv1_0(.dout(w_dff_A_iBxk3XZc2_0),.din(w_dff_A_T1ZfaDTv1_0),.clk(gclk));
	jdff dff_A_iBxk3XZc2_0(.dout(w_dff_A_C1kxaIbC2_0),.din(w_dff_A_iBxk3XZc2_0),.clk(gclk));
	jdff dff_A_C1kxaIbC2_0(.dout(w_dff_A_iSpF9Bqd8_0),.din(w_dff_A_C1kxaIbC2_0),.clk(gclk));
	jdff dff_A_iSpF9Bqd8_0(.dout(w_dff_A_9CN4yY6f6_0),.din(w_dff_A_iSpF9Bqd8_0),.clk(gclk));
	jdff dff_A_9CN4yY6f6_0(.dout(w_dff_A_l5NPhoxX4_0),.din(w_dff_A_9CN4yY6f6_0),.clk(gclk));
	jdff dff_A_l5NPhoxX4_0(.dout(G351),.din(w_dff_A_l5NPhoxX4_0),.clk(gclk));
	jdff dff_A_8Q6yYxeC8_2(.dout(w_dff_A_WryAIHdl9_0),.din(w_dff_A_8Q6yYxeC8_2),.clk(gclk));
	jdff dff_A_WryAIHdl9_0(.dout(w_dff_A_Ns2Rn6eP8_0),.din(w_dff_A_WryAIHdl9_0),.clk(gclk));
	jdff dff_A_Ns2Rn6eP8_0(.dout(w_dff_A_PMnLeR4T5_0),.din(w_dff_A_Ns2Rn6eP8_0),.clk(gclk));
	jdff dff_A_PMnLeR4T5_0(.dout(w_dff_A_UcateCLQ6_0),.din(w_dff_A_PMnLeR4T5_0),.clk(gclk));
	jdff dff_A_UcateCLQ6_0(.dout(w_dff_A_8mJTbhwH7_0),.din(w_dff_A_UcateCLQ6_0),.clk(gclk));
	jdff dff_A_8mJTbhwH7_0(.dout(w_dff_A_pFxc3PwR3_0),.din(w_dff_A_8mJTbhwH7_0),.clk(gclk));
	jdff dff_A_pFxc3PwR3_0(.dout(w_dff_A_fO3yNdQP8_0),.din(w_dff_A_pFxc3PwR3_0),.clk(gclk));
	jdff dff_A_fO3yNdQP8_0(.dout(w_dff_A_6i5VrFKt7_0),.din(w_dff_A_fO3yNdQP8_0),.clk(gclk));
	jdff dff_A_6i5VrFKt7_0(.dout(w_dff_A_eu8WA5MA7_0),.din(w_dff_A_6i5VrFKt7_0),.clk(gclk));
	jdff dff_A_eu8WA5MA7_0(.dout(w_dff_A_03dKo0OU5_0),.din(w_dff_A_eu8WA5MA7_0),.clk(gclk));
	jdff dff_A_03dKo0OU5_0(.dout(w_dff_A_ogyD4tfk5_0),.din(w_dff_A_03dKo0OU5_0),.clk(gclk));
	jdff dff_A_ogyD4tfk5_0(.dout(w_dff_A_uO2oNi8c1_0),.din(w_dff_A_ogyD4tfk5_0),.clk(gclk));
	jdff dff_A_uO2oNi8c1_0(.dout(w_dff_A_QxrJEAvT4_0),.din(w_dff_A_uO2oNi8c1_0),.clk(gclk));
	jdff dff_A_QxrJEAvT4_0(.dout(G372),.din(w_dff_A_QxrJEAvT4_0),.clk(gclk));
	jdff dff_A_cLFUR3629_2(.dout(w_dff_A_TE1fgRoX5_0),.din(w_dff_A_cLFUR3629_2),.clk(gclk));
	jdff dff_A_TE1fgRoX5_0(.dout(w_dff_A_QduNW8g18_0),.din(w_dff_A_TE1fgRoX5_0),.clk(gclk));
	jdff dff_A_QduNW8g18_0(.dout(w_dff_A_BAQ5CWZM6_0),.din(w_dff_A_QduNW8g18_0),.clk(gclk));
	jdff dff_A_BAQ5CWZM6_0(.dout(w_dff_A_mB2QYAqB5_0),.din(w_dff_A_BAQ5CWZM6_0),.clk(gclk));
	jdff dff_A_mB2QYAqB5_0(.dout(w_dff_A_Rz2uBJNn8_0),.din(w_dff_A_mB2QYAqB5_0),.clk(gclk));
	jdff dff_A_Rz2uBJNn8_0(.dout(w_dff_A_ziIlOHJp2_0),.din(w_dff_A_Rz2uBJNn8_0),.clk(gclk));
	jdff dff_A_ziIlOHJp2_0(.dout(w_dff_A_ryW1PJWv3_0),.din(w_dff_A_ziIlOHJp2_0),.clk(gclk));
	jdff dff_A_ryW1PJWv3_0(.dout(w_dff_A_RxKSzTvT1_0),.din(w_dff_A_ryW1PJWv3_0),.clk(gclk));
	jdff dff_A_RxKSzTvT1_0(.dout(w_dff_A_ZLCaXi6H5_0),.din(w_dff_A_RxKSzTvT1_0),.clk(gclk));
	jdff dff_A_ZLCaXi6H5_0(.dout(w_dff_A_P68wLghG5_0),.din(w_dff_A_ZLCaXi6H5_0),.clk(gclk));
	jdff dff_A_P68wLghG5_0(.dout(w_dff_A_tmYKP9X75_0),.din(w_dff_A_P68wLghG5_0),.clk(gclk));
	jdff dff_A_tmYKP9X75_0(.dout(G369),.din(w_dff_A_tmYKP9X75_0),.clk(gclk));
	jdff dff_A_dB0sU7VX1_2(.dout(w_dff_A_MxtLPZu36_0),.din(w_dff_A_dB0sU7VX1_2),.clk(gclk));
	jdff dff_A_MxtLPZu36_0(.dout(w_dff_A_HotI6sFd3_0),.din(w_dff_A_MxtLPZu36_0),.clk(gclk));
	jdff dff_A_HotI6sFd3_0(.dout(w_dff_A_ubLH2ZY53_0),.din(w_dff_A_HotI6sFd3_0),.clk(gclk));
	jdff dff_A_ubLH2ZY53_0(.dout(w_dff_A_mp4Cxt8K0_0),.din(w_dff_A_ubLH2ZY53_0),.clk(gclk));
	jdff dff_A_mp4Cxt8K0_0(.dout(w_dff_A_3cpAejMl5_0),.din(w_dff_A_mp4Cxt8K0_0),.clk(gclk));
	jdff dff_A_3cpAejMl5_0(.dout(w_dff_A_KsaeLJyy1_0),.din(w_dff_A_3cpAejMl5_0),.clk(gclk));
	jdff dff_A_KsaeLJyy1_0(.dout(w_dff_A_W8BEe51M6_0),.din(w_dff_A_KsaeLJyy1_0),.clk(gclk));
	jdff dff_A_W8BEe51M6_0(.dout(w_dff_A_SjPffqPZ2_0),.din(w_dff_A_W8BEe51M6_0),.clk(gclk));
	jdff dff_A_SjPffqPZ2_0(.dout(w_dff_A_cd2AsH7w8_0),.din(w_dff_A_SjPffqPZ2_0),.clk(gclk));
	jdff dff_A_cd2AsH7w8_0(.dout(w_dff_A_TSaMQ2GW2_0),.din(w_dff_A_cd2AsH7w8_0),.clk(gclk));
	jdff dff_A_TSaMQ2GW2_0(.dout(w_dff_A_QIJzC3fc7_0),.din(w_dff_A_TSaMQ2GW2_0),.clk(gclk));
	jdff dff_A_QIJzC3fc7_0(.dout(w_dff_A_Aew9ff5B4_0),.din(w_dff_A_QIJzC3fc7_0),.clk(gclk));
	jdff dff_A_Aew9ff5B4_0(.dout(w_dff_A_yhA4RyZz4_0),.din(w_dff_A_Aew9ff5B4_0),.clk(gclk));
	jdff dff_A_yhA4RyZz4_0(.dout(G399),.din(w_dff_A_yhA4RyZz4_0),.clk(gclk));
	jdff dff_A_pYXSlu0u3_2(.dout(w_dff_A_cyy8OSOT3_0),.din(w_dff_A_pYXSlu0u3_2),.clk(gclk));
	jdff dff_A_cyy8OSOT3_0(.dout(w_dff_A_1c7FcxnV5_0),.din(w_dff_A_cyy8OSOT3_0),.clk(gclk));
	jdff dff_A_1c7FcxnV5_0(.dout(w_dff_A_5kO10u8s0_0),.din(w_dff_A_1c7FcxnV5_0),.clk(gclk));
	jdff dff_A_5kO10u8s0_0(.dout(w_dff_A_3BBkXED38_0),.din(w_dff_A_5kO10u8s0_0),.clk(gclk));
	jdff dff_A_3BBkXED38_0(.dout(w_dff_A_KwwakGil9_0),.din(w_dff_A_3BBkXED38_0),.clk(gclk));
	jdff dff_A_KwwakGil9_0(.dout(w_dff_A_VcxXrr4O6_0),.din(w_dff_A_KwwakGil9_0),.clk(gclk));
	jdff dff_A_VcxXrr4O6_0(.dout(w_dff_A_NdrhWOkV6_0),.din(w_dff_A_VcxXrr4O6_0),.clk(gclk));
	jdff dff_A_NdrhWOkV6_0(.dout(w_dff_A_MsZJIKpq4_0),.din(w_dff_A_NdrhWOkV6_0),.clk(gclk));
	jdff dff_A_MsZJIKpq4_0(.dout(G364),.din(w_dff_A_MsZJIKpq4_0),.clk(gclk));
	jdff dff_A_7VLwJoOx0_1(.dout(w_dff_A_PssIiQXc0_0),.din(w_dff_A_7VLwJoOx0_1),.clk(gclk));
	jdff dff_A_PssIiQXc0_0(.dout(w_dff_A_ePdVpKv11_0),.din(w_dff_A_PssIiQXc0_0),.clk(gclk));
	jdff dff_A_ePdVpKv11_0(.dout(w_dff_A_ctvXemYK2_0),.din(w_dff_A_ePdVpKv11_0),.clk(gclk));
	jdff dff_A_ctvXemYK2_0(.dout(w_dff_A_l6ymKFxy6_0),.din(w_dff_A_ctvXemYK2_0),.clk(gclk));
	jdff dff_A_l6ymKFxy6_0(.dout(w_dff_A_JF0rtjhO4_0),.din(w_dff_A_l6ymKFxy6_0),.clk(gclk));
	jdff dff_A_JF0rtjhO4_0(.dout(w_dff_A_dYO5zxbJ5_0),.din(w_dff_A_JF0rtjhO4_0),.clk(gclk));
	jdff dff_A_dYO5zxbJ5_0(.dout(w_dff_A_mEcX5aBD7_0),.din(w_dff_A_dYO5zxbJ5_0),.clk(gclk));
	jdff dff_A_mEcX5aBD7_0(.dout(w_dff_A_gsv9fq2T7_0),.din(w_dff_A_mEcX5aBD7_0),.clk(gclk));
	jdff dff_A_gsv9fq2T7_0(.dout(w_dff_A_pVLj9Wzt1_0),.din(w_dff_A_gsv9fq2T7_0),.clk(gclk));
	jdff dff_A_pVLj9Wzt1_0(.dout(w_dff_A_lIpENpu48_0),.din(w_dff_A_pVLj9Wzt1_0),.clk(gclk));
	jdff dff_A_lIpENpu48_0(.dout(w_dff_A_aE38d95m6_0),.din(w_dff_A_lIpENpu48_0),.clk(gclk));
	jdff dff_A_aE38d95m6_0(.dout(w_dff_A_ARHG76Xk0_0),.din(w_dff_A_aE38d95m6_0),.clk(gclk));
	jdff dff_A_ARHG76Xk0_0(.dout(G396),.din(w_dff_A_ARHG76Xk0_0),.clk(gclk));
	jdff dff_A_cMTHFec67_1(.dout(w_dff_A_rfD6WCBD7_0),.din(w_dff_A_cMTHFec67_1),.clk(gclk));
	jdff dff_A_rfD6WCBD7_0(.dout(w_dff_A_aG5zNwq98_0),.din(w_dff_A_rfD6WCBD7_0),.clk(gclk));
	jdff dff_A_aG5zNwq98_0(.dout(w_dff_A_5vo19zre5_0),.din(w_dff_A_aG5zNwq98_0),.clk(gclk));
	jdff dff_A_5vo19zre5_0(.dout(w_dff_A_yiMVGmsJ9_0),.din(w_dff_A_5vo19zre5_0),.clk(gclk));
	jdff dff_A_yiMVGmsJ9_0(.dout(w_dff_A_SuASy8FB1_0),.din(w_dff_A_yiMVGmsJ9_0),.clk(gclk));
	jdff dff_A_SuASy8FB1_0(.dout(w_dff_A_KaTjYwsO0_0),.din(w_dff_A_SuASy8FB1_0),.clk(gclk));
	jdff dff_A_KaTjYwsO0_0(.dout(w_dff_A_igJmY0qZ1_0),.din(w_dff_A_KaTjYwsO0_0),.clk(gclk));
	jdff dff_A_igJmY0qZ1_0(.dout(G384),.din(w_dff_A_igJmY0qZ1_0),.clk(gclk));
	jdff dff_A_tne6B1924_2(.dout(w_dff_A_bsRgQ6HQ9_0),.din(w_dff_A_tne6B1924_2),.clk(gclk));
	jdff dff_A_bsRgQ6HQ9_0(.dout(w_dff_A_BbNo7saQ6_0),.din(w_dff_A_bsRgQ6HQ9_0),.clk(gclk));
	jdff dff_A_BbNo7saQ6_0(.dout(w_dff_A_7rhlFlZj9_0),.din(w_dff_A_BbNo7saQ6_0),.clk(gclk));
	jdff dff_A_7rhlFlZj9_0(.dout(w_dff_A_eBfPA8zD8_0),.din(w_dff_A_7rhlFlZj9_0),.clk(gclk));
	jdff dff_A_eBfPA8zD8_0(.dout(w_dff_A_QlyGS8GL6_0),.din(w_dff_A_eBfPA8zD8_0),.clk(gclk));
	jdff dff_A_QlyGS8GL6_0(.dout(w_dff_A_uqG9iPFp0_0),.din(w_dff_A_QlyGS8GL6_0),.clk(gclk));
	jdff dff_A_uqG9iPFp0_0(.dout(G367),.din(w_dff_A_uqG9iPFp0_0),.clk(gclk));
	jdff dff_A_vfRDkQlW9_1(.dout(w_dff_A_nNRWStQ55_0),.din(w_dff_A_vfRDkQlW9_1),.clk(gclk));
	jdff dff_A_nNRWStQ55_0(.dout(w_dff_A_XPIeNpRI4_0),.din(w_dff_A_nNRWStQ55_0),.clk(gclk));
	jdff dff_A_XPIeNpRI4_0(.dout(w_dff_A_zoC0sDli6_0),.din(w_dff_A_XPIeNpRI4_0),.clk(gclk));
	jdff dff_A_zoC0sDli6_0(.dout(w_dff_A_KukjoOi82_0),.din(w_dff_A_zoC0sDli6_0),.clk(gclk));
	jdff dff_A_KukjoOi82_0(.dout(w_dff_A_SL9TcYRZ1_0),.din(w_dff_A_KukjoOi82_0),.clk(gclk));
	jdff dff_A_SL9TcYRZ1_0(.dout(G387),.din(w_dff_A_SL9TcYRZ1_0),.clk(gclk));
	jdff dff_A_ywVOaL5R9_1(.dout(w_dff_A_EPAaCQJU2_0),.din(w_dff_A_ywVOaL5R9_1),.clk(gclk));
	jdff dff_A_EPAaCQJU2_0(.dout(w_dff_A_iAa84ZRP0_0),.din(w_dff_A_EPAaCQJU2_0),.clk(gclk));
	jdff dff_A_iAa84ZRP0_0(.dout(w_dff_A_S8cpcl4d3_0),.din(w_dff_A_iAa84ZRP0_0),.clk(gclk));
	jdff dff_A_S8cpcl4d3_0(.dout(w_dff_A_eKIaLvsK6_0),.din(w_dff_A_S8cpcl4d3_0),.clk(gclk));
	jdff dff_A_eKIaLvsK6_0(.dout(w_dff_A_r4TZM15t1_0),.din(w_dff_A_eKIaLvsK6_0),.clk(gclk));
	jdff dff_A_r4TZM15t1_0(.dout(w_dff_A_NaAXIQL28_0),.din(w_dff_A_r4TZM15t1_0),.clk(gclk));
	jdff dff_A_NaAXIQL28_0(.dout(G393),.din(w_dff_A_NaAXIQL28_0),.clk(gclk));
	jdff dff_A_Ezxpsepx8_1(.dout(w_dff_A_PGrXCgsV6_0),.din(w_dff_A_Ezxpsepx8_1),.clk(gclk));
	jdff dff_A_PGrXCgsV6_0(.dout(w_dff_A_k8QWObmZ5_0),.din(w_dff_A_PGrXCgsV6_0),.clk(gclk));
	jdff dff_A_k8QWObmZ5_0(.dout(w_dff_A_PWmGEvrn1_0),.din(w_dff_A_k8QWObmZ5_0),.clk(gclk));
	jdff dff_A_PWmGEvrn1_0(.dout(w_dff_A_it6GNzsI2_0),.din(w_dff_A_PWmGEvrn1_0),.clk(gclk));
	jdff dff_A_it6GNzsI2_0(.dout(w_dff_A_dY0mTyTs3_0),.din(w_dff_A_it6GNzsI2_0),.clk(gclk));
	jdff dff_A_dY0mTyTs3_0(.dout(G390),.din(w_dff_A_dY0mTyTs3_0),.clk(gclk));
	jdff dff_A_XSgKg9OT8_1(.dout(w_dff_A_aY5NSo1j9_0),.din(w_dff_A_XSgKg9OT8_1),.clk(gclk));
	jdff dff_A_aY5NSo1j9_0(.dout(w_dff_A_i549ZAOL4_0),.din(w_dff_A_aY5NSo1j9_0),.clk(gclk));
	jdff dff_A_i549ZAOL4_0(.dout(w_dff_A_sx55JEQH2_0),.din(w_dff_A_i549ZAOL4_0),.clk(gclk));
	jdff dff_A_sx55JEQH2_0(.dout(G378),.din(w_dff_A_sx55JEQH2_0),.clk(gclk));
	jdff dff_A_lw3JEhUA7_1(.dout(w_dff_A_viqP63LY9_0),.din(w_dff_A_lw3JEhUA7_1),.clk(gclk));
	jdff dff_A_viqP63LY9_0(.dout(w_dff_A_yVUWWQzq4_0),.din(w_dff_A_viqP63LY9_0),.clk(gclk));
	jdff dff_A_yVUWWQzq4_0(.dout(w_dff_A_jCTZi0uI1_0),.din(w_dff_A_yVUWWQzq4_0),.clk(gclk));
	jdff dff_A_jCTZi0uI1_0(.dout(G375),.din(w_dff_A_jCTZi0uI1_0),.clk(gclk));
	jdff dff_A_qbIctODl9_1(.dout(w_dff_A_BnZP0qRU9_0),.din(w_dff_A_qbIctODl9_1),.clk(gclk));
	jdff dff_A_BnZP0qRU9_0(.dout(w_dff_A_ndrSBHWg4_0),.din(w_dff_A_BnZP0qRU9_0),.clk(gclk));
	jdff dff_A_ndrSBHWg4_0(.dout(w_dff_A_4DmmGz8o2_0),.din(w_dff_A_ndrSBHWg4_0),.clk(gclk));
	jdff dff_A_4DmmGz8o2_0(.dout(G381),.din(w_dff_A_4DmmGz8o2_0),.clk(gclk));
	jdff dff_A_0IWw5YRT1_1(.dout(G407),.din(w_dff_A_0IWw5YRT1_1),.clk(gclk));
	jdff dff_A_A80hFMiP3_2(.dout(w_dff_A_GxCQ8ad60_0),.din(w_dff_A_A80hFMiP3_2),.clk(gclk));
	jdff dff_A_GxCQ8ad60_0(.dout(G402),.din(w_dff_A_GxCQ8ad60_0),.clk(gclk));
endmodule

