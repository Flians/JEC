module rf_c7552(G4528, G4526, G4432, G4427, G4420, G4410, G4405, G4400, G3743, G3729, G3723, G3717, G3711, G3701, G3698, G3705, G2256, G2253, G2247, G2236, G2230, G2204, G1492, G1486, G1455, G1197, G339, G240, G239, G4393, G238, G234, G231, G228, G2239, G225, G2224, G221, G220, G219, G218, G217, G214, G236, G210, G208, G207, G209, G206, G205, G204, G1496, G203, G111, G202, G152, G100, G2218, G161, G97, G88, G223, G87, G118, G233, G53, G3749, G212, G84, G4415, G5, G222, G83, G226, G81, G82, G144, G227, G79, G64, G159, G94, G211, G66, G127, G230, G15, G61, G110, G196, G26, G23, G63, G4394, G78, G12, G62, G156, G73, G18, G9, G1459, G135, G198, G188, G199, G113, G76, G57, G237, G164, G59, G224, G35, G158, G41, G80, G55, G192, G229, G85, G114, G29, G77, G160, G75, G54, G1469, G153, G232, G194, G106, G65, G109, G216, G115, G121, G167, G124, G138, G130, G186, G4437, G200, G170, G134, G1462, G141, G150, G151, G47, G174, G154, G3737, G215, G155, G133, G185, G162, G58, G163, G165, G60, G166, G1480, G147, G168, G44, G1, G56, G169, G171, G2211, G157, G172, G2208, G193, G197, G173, G86, G175, G89, G50, G189, G213, G176, G38, G178, G179, G74, G180, G181, G69, G182, G183, G177, G184, G103, G32, G187, G112, G191, G235, G190, G195, G70, G201, G399, G370, G338, G321, G368, G362, G359, G471, G422, G344, G307, G304, G301, G273, G336, G333, G419, G327, G310, G276, G252, G295, G249, G416, G412, G382, G319, G379, G376, G365, G397, G353, G347, G394, G391, G388, G281, G330, G552, G316, G534, G554, G546, G530, G438, G270, G450, G432, G540, G418, G3, G448, G350, G484, G558, G482, G480, G404, G550, G494, G469, G524, G522, G298, G538, G442, G246, G258, G492, G548, G556, G440, G486, G544, G536, G313, G490, G542, G292, G414, G560, G528, G496, G532, G279, G526, G436, G488, G478, G324, G444, G402, G453, G278, G410, G2, G284, G408, G446, G373, G406, G264, G385, G286, G289, G356, G341);
    input G4528, G4526, G4432, G4427, G4420, G4410, G4405, G4400, G3743, G3729, G3723, G3717, G3711, G3701, G3698, G3705, G2256, G2253, G2247, G2236, G2230, G2204, G1492, G1486, G1455, G1197, G339, G240, G239, G4393, G238, G234, G231, G228, G2239, G225, G2224, G221, G220, G219, G218, G217, G214, G236, G210, G208, G207, G209, G206, G205, G204, G1496, G203, G111, G202, G152, G100, G2218, G161, G97, G88, G223, G87, G118, G233, G53, G3749, G212, G84, G4415, G5, G222, G83, G226, G81, G82, G144, G227, G79, G64, G159, G94, G211, G66, G127, G230, G15, G61, G110, G196, G26, G23, G63, G4394, G78, G12, G62, G156, G73, G18, G9, G1459, G135, G198, G188, G199, G113, G76, G57, G237, G164, G59, G224, G35, G158, G41, G80, G55, G192, G229, G85, G114, G29, G77, G160, G75, G54, G1469, G153, G232, G194, G106, G65, G109, G216, G115, G121, G167, G124, G138, G130, G186, G4437, G200, G170, G134, G1462, G141, G150, G151, G47, G174, G154, G3737, G215, G155, G133, G185, G162, G58, G163, G165, G60, G166, G1480, G147, G168, G44, G1, G56, G169, G171, G2211, G157, G172, G2208, G193, G197, G173, G86, G175, G89, G50, G189, G213, G176, G38, G178, G179, G74, G180, G181, G69, G182, G183, G177, G184, G103, G32, G187, G112, G191, G235, G190, G195, G70, G201;
    output G399, G370, G338, G321, G368, G362, G359, G471, G422, G344, G307, G304, G301, G273, G336, G333, G419, G327, G310, G276, G252, G295, G249, G416, G412, G382, G319, G379, G376, G365, G397, G353, G347, G394, G391, G388, G281, G330, G552, G316, G534, G554, G546, G530, G438, G270, G450, G432, G540, G418, G3, G448, G350, G484, G558, G482, G480, G404, G550, G494, G469, G524, G522, G298, G538, G442, G246, G258, G492, G548, G556, G440, G486, G544, G536, G313, G490, G542, G292, G414, G560, G528, G496, G532, G279, G526, G436, G488, G478, G324, G444, G402, G453, G278, G410, G2, G284, G408, G446, G373, G406, G264, G385, G286, G289, G356, G341;
    wire n316;
    wire n320;
    wire n323;
    wire n326;
    wire n330;
    wire n333;
    wire n336;
    wire n340;
    wire n344;
    wire n347;
    wire n350;
    wire n354;
    wire n357;
    wire n360;
    wire n364;
    wire n368;
    wire n371;
    wire n374;
    wire n378;
    wire n381;
    wire n384;
    wire n388;
    wire n392;
    wire n395;
    wire n398;
    wire n402;
    wire n405;
    wire n408;
    wire n412;
    wire n416;
    wire n419;
    wire n423;
    wire n426;
    wire n429;
    wire n433;
    wire n437;
    wire n441;
    wire n444;
    wire n448;
    wire n452;
    wire n455;
    wire n459;
    wire n463;
    wire n467;
    wire n471;
    wire n474;
    wire n478;
    wire n482;
    wire n486;
    wire n490;
    wire n494;
    wire n497;
    wire n501;
    wire n504;
    wire n507;
    wire n511;
    wire n515;
    wire n519;
    wire n523;
    wire n526;
    wire n529;
    wire n533;
    wire n537;
    wire n540;
    wire n544;
    wire n548;
    wire n551;
    wire n555;
    wire n558;
    wire n561;
    wire n565;
    wire n569;
    wire n573;
    wire n576;
    wire n579;
    wire n583;
    wire n586;
    wire n590;
    wire n594;
    wire n598;
    wire n602;
    wire n605;
    wire n608;
    wire n612;
    wire n615;
    wire n619;
    wire n623;
    wire n627;
    wire n631;
    wire n635;
    wire n639;
    wire n643;
    wire n647;
    wire n651;
    wire n655;
    wire n659;
    wire n663;
    wire n667;
    wire n671;
    wire n675;
    wire n679;
    wire n683;
    wire n687;
    wire n691;
    wire n695;
    wire n699;
    wire n703;
    wire n707;
    wire n710;
    wire n714;
    wire n717;
    wire n720;
    wire n724;
    wire n728;
    wire n732;
    wire n735;
    wire n739;
    wire n742;
    wire n745;
    wire n749;
    wire n753;
    wire n757;
    wire n761;
    wire n765;
    wire n768;
    wire n771;
    wire n775;
    wire n779;
    wire n783;
    wire n786;
    wire n790;
    wire n794;
    wire n798;
    wire n802;
    wire n806;
    wire n810;
    wire n814;
    wire n818;
    wire n822;
    wire n825;
    wire n829;
    wire n833;
    wire n837;
    wire n841;
    wire n845;
    wire n849;
    wire n853;
    wire n857;
    wire n861;
    wire n865;
    wire n869;
    wire n872;
    wire n876;
    wire n880;
    wire n884;
    wire n888;
    wire n891;
    wire n895;
    wire n899;
    wire n903;
    wire n907;
    wire n911;
    wire n915;
    wire n919;
    wire n922;
    wire n926;
    wire n930;
    wire n933;
    wire n937;
    wire n941;
    wire n945;
    wire n949;
    wire n953;
    wire n957;
    wire n961;
    wire n964;
    wire n968;
    wire n972;
    wire n976;
    wire n980;
    wire n983;
    wire n987;
    wire n990;
    wire n994;
    wire n998;
    wire n1001;
    wire n1005;
    wire n1008;
    wire n1011;
    wire n1015;
    wire n1019;
    wire n1022;
    wire n1026;
    wire n1030;
    wire n1034;
    wire n1037;
    wire n1041;
    wire n1045;
    wire n1049;
    wire n1053;
    wire n1057;
    wire n1061;
    wire n1065;
    wire n1069;
    wire n1073;
    wire n1076;
    wire n1080;
    wire n1084;
    wire n1088;
    wire n1092;
    wire n1095;
    wire n1099;
    wire n1103;
    wire n1107;
    wire n1111;
    wire n1115;
    wire n1118;
    wire n1122;
    wire n1126;
    wire n1130;
    wire n1134;
    wire n1137;
    wire n1141;
    wire n1145;
    wire n1149;
    wire n1153;
    wire n1157;
    wire n1161;
    wire n1164;
    wire n1168;
    wire n1171;
    wire n1175;
    wire n1178;
    wire n1182;
    wire n1186;
    wire n1189;
    wire n1193;
    wire n1196;
    wire n1200;
    wire n1204;
    wire n1208;
    wire n1212;
    wire n1216;
    wire n1220;
    wire n1224;
    wire n1228;
    wire n1231;
    wire n1235;
    wire n1238;
    wire n1242;
    wire n1245;
    wire n1249;
    wire n1253;
    wire n1257;
    wire n1260;
    wire n1264;
    wire n1268;
    wire n1272;
    wire n1276;
    wire n1279;
    wire n1283;
    wire n1287;
    wire n1291;
    wire n1295;
    wire n1299;
    wire n1302;
    wire n1306;
    wire n1310;
    wire n1314;
    wire n1318;
    wire n1321;
    wire n1325;
    wire n1329;
    wire n1333;
    wire n1337;
    wire n1341;
    wire n1345;
    wire n1349;
    wire n1352;
    wire n1356;
    wire n1360;
    wire n1363;
    wire n1366;
    wire n1370;
    wire n1374;
    wire n1377;
    wire n1380;
    wire n1384;
    wire n1387;
    wire n1391;
    wire n1394;
    wire n1398;
    wire n1402;
    wire n1406;
    wire n1410;
    wire n1414;
    wire n1418;
    wire n1422;
    wire n1425;
    wire n1429;
    wire n1433;
    wire n1437;
    wire n1441;
    wire n1445;
    wire n1448;
    wire n1452;
    wire n1456;
    wire n1460;
    wire n1463;
    wire n1467;
    wire n1471;
    wire n1475;
    wire n1479;
    wire n1482;
    wire n1486;
    wire n1490;
    wire n1494;
    wire n1497;
    wire n1501;
    wire n1505;
    wire n1509;
    wire n1513;
    wire n1517;
    wire n1520;
    wire n1524;
    wire n1528;
    wire n1531;
    wire n1535;
    wire n1538;
    wire n1542;
    wire n1546;
    wire n1550;
    wire n1554;
    wire n1557;
    wire n1561;
    wire n1564;
    wire n1568;
    wire n1571;
    wire n1575;
    wire n1579;
    wire n1583;
    wire n1587;
    wire n1591;
    wire n1594;
    wire n1598;
    wire n1602;
    wire n1606;
    wire n1609;
    wire n1613;
    wire n1617;
    wire n1621;
    wire n1624;
    wire n1628;
    wire n1632;
    wire n1636;
    wire n1640;
    wire n1643;
    wire n1647;
    wire n1651;
    wire n1655;
    wire n1658;
    wire n1662;
    wire n1666;
    wire n1670;
    wire n1674;
    wire n1678;
    wire n1682;
    wire n1685;
    wire n1689;
    wire n1693;
    wire n1697;
    wire n1701;
    wire n1704;
    wire n1708;
    wire n1712;
    wire n1715;
    wire n1719;
    wire n1722;
    wire n1725;
    wire n1729;
    wire n1732;
    wire n1736;
    wire n1740;
    wire n1744;
    wire n1748;
    wire n1752;
    wire n1756;
    wire n1760;
    wire n1763;
    wire n1767;
    wire n1770;
    wire n1774;
    wire n1778;
    wire n1781;
    wire n1785;
    wire n1788;
    wire n1792;
    wire n1796;
    wire n1799;
    wire n1803;
    wire n1807;
    wire n1810;
    wire n1813;
    wire n1816;
    wire n1820;
    wire n1824;
    wire n1828;
    wire n1832;
    wire n1836;
    wire n1840;
    wire n1843;
    wire n1847;
    wire n1851;
    wire n1855;
    wire n1859;
    wire n1863;
    wire n1867;
    wire n1870;
    wire n1874;
    wire n1878;
    wire n1882;
    wire n1886;
    wire n1890;
    wire n1894;
    wire n1897;
    wire n1901;
    wire n1905;
    wire n1909;
    wire n1913;
    wire n1917;
    wire n1921;
    wire n1924;
    wire n1928;
    wire n1932;
    wire n1936;
    wire n1940;
    wire n1944;
    wire n1948;
    wire n1952;
    wire n1956;
    wire n1960;
    wire n1963;
    wire n1967;
    wire n1971;
    wire n1975;
    wire n1979;
    wire n1983;
    wire n1987;
    wire n1991;
    wire n1995;
    wire n1999;
    wire n2003;
    wire n2007;
    wire n2011;
    wire n2014;
    wire n2018;
    wire n2021;
    wire n2024;
    wire n2028;
    wire n2032;
    wire n2035;
    wire n2039;
    wire n2043;
    wire n2046;
    wire n2050;
    wire n2054;
    wire n2058;
    wire n2062;
    wire n2066;
    wire n2070;
    wire n2074;
    wire n2078;
    wire n2082;
    wire n2086;
    wire n2090;
    wire n2094;
    wire n2098;
    wire n2102;
    wire n2106;
    wire n2110;
    wire n2114;
    wire n2118;
    wire n2122;
    wire n2126;
    wire n2130;
    wire n2133;
    wire n2137;
    wire n2141;
    wire n2145;
    wire n2149;
    wire n2153;
    wire n2157;
    wire n2161;
    wire n2165;
    wire n2169;
    wire n2173;
    wire n2177;
    wire n2181;
    wire n2185;
    wire n2189;
    wire n2192;
    wire n2196;
    wire n2200;
    wire n2204;
    wire n2208;
    wire n2212;
    wire n2216;
    wire n2219;
    wire n2223;
    wire n2227;
    wire n2231;
    wire n2235;
    wire n2239;
    wire n2243;
    wire n2247;
    wire n2250;
    wire n2254;
    wire n2258;
    wire n2261;
    wire n2265;
    wire n2268;
    wire n2272;
    wire n2276;
    wire n2280;
    wire n2283;
    wire n2287;
    wire n2291;
    wire n2295;
    wire n2299;
    wire n2303;
    wire n2307;
    wire n2310;
    wire n2314;
    wire n2318;
    wire n2321;
    wire n2325;
    wire n2329;
    wire n2333;
    wire n2337;
    wire n2340;
    wire n2344;
    wire n2348;
    wire n2352;
    wire n2356;
    wire n2360;
    wire n2363;
    wire n2367;
    wire n2371;
    wire n2375;
    wire n2379;
    wire n2383;
    wire n2387;
    wire n2390;
    wire n2394;
    wire n2397;
    wire n2401;
    wire n2405;
    wire n2408;
    wire n2412;
    wire n2416;
    wire n2419;
    wire n2422;
    wire n2426;
    wire n2430;
    wire n2434;
    wire n2438;
    wire n2441;
    wire n2445;
    wire n2449;
    wire n2453;
    wire n2457;
    wire n2460;
    wire n2464;
    wire n2468;
    wire n2472;
    wire n2476;
    wire n2480;
    wire n2484;
    wire n2488;
    wire n2491;
    wire n2495;
    wire n2499;
    wire n2502;
    wire n2506;
    wire n2510;
    wire n2514;
    wire n2518;
    wire n2522;
    wire n2526;
    wire n2530;
    wire n2534;
    wire n2537;
    wire n2541;
    wire n2545;
    wire n2549;
    wire n2553;
    wire n2556;
    wire n2560;
    wire n2564;
    wire n2567;
    wire n2571;
    wire n2575;
    wire n2579;
    wire n2583;
    wire n2586;
    wire n2590;
    wire n2594;
    wire n2598;
    wire n2602;
    wire n2605;
    wire n2608;
    wire n2612;
    wire n2616;
    wire n2620;
    wire n2624;
    wire n2627;
    wire n2631;
    wire n2635;
    wire n2639;
    wire n2643;
    wire n2646;
    wire n2650;
    wire n2653;
    wire n2657;
    wire n2661;
    wire n2664;
    wire n2668;
    wire n2672;
    wire n2675;
    wire n2679;
    wire n2683;
    wire n2687;
    wire n2691;
    wire n2695;
    wire n2699;
    wire n2703;
    wire n2706;
    wire n2710;
    wire n2713;
    wire n2717;
    wire n2721;
    wire n2725;
    wire n2729;
    wire n2733;
    wire n2737;
    wire n2741;
    wire n2745;
    wire n2749;
    wire n2753;
    wire n2757;
    wire n2761;
    wire n2765;
    wire n2769;
    wire n2773;
    wire n2777;
    wire n2781;
    wire n2785;
    wire n2789;
    wire n2793;
    wire n2797;
    wire n2801;
    wire n2805;
    wire n2809;
    wire n2813;
    wire n2817;
    wire n2821;
    wire n2825;
    wire n2829;
    wire n2833;
    wire n2837;
    wire n2841;
    wire n2845;
    wire n2849;
    wire n2853;
    wire n2857;
    wire n2860;
    wire n2864;
    wire n2868;
    wire n2872;
    wire n2876;
    wire n2880;
    wire n2884;
    wire n2887;
    wire n2891;
    wire n2895;
    wire n2899;
    wire n2902;
    wire n2906;
    wire n2910;
    wire n2913;
    wire n2917;
    wire n2921;
    wire n2925;
    wire n2929;
    wire n2933;
    wire n2937;
    wire n2940;
    wire n2944;
    wire n2948;
    wire n2952;
    wire n2956;
    wire n2960;
    wire n2964;
    wire n2968;
    wire n2972;
    wire n2976;
    wire n2980;
    wire n2984;
    wire n2988;
    wire n2992;
    wire n2996;
    wire n3000;
    wire n3004;
    wire n3008;
    wire n3012;
    wire n3016;
    wire n3020;
    wire n3024;
    wire n3028;
    wire n3032;
    wire n3036;
    wire n3040;
    wire n3044;
    wire n3048;
    wire n3052;
    wire n3056;
    wire n3060;
    wire n3064;
    wire n3068;
    wire n3072;
    wire n3076;
    wire n3080;
    wire n3084;
    wire n3088;
    wire n3092;
    wire n3096;
    wire n3100;
    wire n3104;
    wire n3108;
    wire n3112;
    wire n3116;
    wire n3120;
    wire n3124;
    wire n3128;
    wire n3132;
    wire n3136;
    wire n3140;
    wire n3144;
    wire n3148;
    wire n3151;
    wire n3155;
    wire n3159;
    wire n3163;
    wire n3167;
    wire n3171;
    wire n3175;
    wire n3178;
    wire n3182;
    wire n3186;
    wire n3190;
    wire n3194;
    wire n3198;
    wire n3202;
    wire n3206;
    wire n3209;
    wire n3213;
    wire n3217;
    wire n3221;
    wire n3225;
    wire n3228;
    wire n3232;
    wire n3236;
    wire n3240;
    wire n3244;
    wire n3248;
    wire n3252;
    wire n3256;
    wire n3260;
    wire n3263;
    wire n3267;
    wire n3271;
    wire n3275;
    wire n3279;
    wire n3282;
    wire n3286;
    wire n3290;
    wire n3294;
    wire n3298;
    wire n3301;
    wire n3305;
    wire n3309;
    wire n3312;
    wire n3316;
    wire n3320;
    wire n3324;
    wire n3328;
    wire n3332;
    wire n3336;
    wire n3340;
    wire n3344;
    wire n3348;
    wire n3351;
    wire n3355;
    wire n3359;
    wire n3363;
    wire n3367;
    wire n3371;
    wire n3375;
    wire n3379;
    wire n3383;
    wire n3387;
    wire n3391;
    wire n3395;
    wire n3399;
    wire n3403;
    wire n3407;
    wire n3411;
    wire n3415;
    wire n3419;
    wire n3423;
    wire n3427;
    wire n3431;
    wire n3435;
    wire n3439;
    wire n3443;
    wire n3447;
    wire n3451;
    wire n3455;
    wire n3459;
    wire n3463;
    wire n3467;
    wire n3471;
    wire n3475;
    wire n3479;
    wire n3483;
    wire n3487;
    wire n3491;
    wire n3495;
    wire n3499;
    wire n3503;
    wire n3507;
    wire n3510;
    wire n3514;
    wire n3517;
    wire n3521;
    wire n3525;
    wire n3529;
    wire n3533;
    wire n3537;
    wire n3541;
    wire n3544;
    wire n3548;
    wire n3551;
    wire n3555;
    wire n3559;
    wire n3563;
    wire n3567;
    wire n3571;
    wire n3575;
    wire n3579;
    wire n3583;
    wire n3587;
    wire n3590;
    wire n3594;
    wire n3597;
    wire n3601;
    wire n3605;
    wire n3609;
    wire n3613;
    wire n3617;
    wire n3621;
    wire n3625;
    wire n3629;
    wire n3633;
    wire n3637;
    wire n3641;
    wire n3645;
    wire n3649;
    wire n3653;
    wire n3657;
    wire n3661;
    wire n3665;
    wire n3669;
    wire n3673;
    wire n3677;
    wire n3681;
    wire n3685;
    wire n3689;
    wire n3693;
    wire n3697;
    wire n3701;
    wire n3705;
    wire n3709;
    wire n3713;
    wire n3717;
    wire n3721;
    wire n3725;
    wire n3729;
    wire n3733;
    wire n3737;
    wire n3741;
    wire n3745;
    wire n3749;
    wire n3753;
    wire n3757;
    wire n3761;
    wire n3765;
    wire n3768;
    wire n3772;
    wire n3776;
    wire n3780;
    wire n3784;
    wire n3788;
    wire n3792;
    wire n3796;
    wire n3799;
    wire n3803;
    wire n3807;
    wire n3811;
    wire n3815;
    wire n3819;
    wire n3823;
    wire n3826;
    wire n3830;
    wire n3833;
    wire n3837;
    wire n3841;
    wire n3845;
    wire n3849;
    wire n3853;
    wire n3856;
    wire n3860;
    wire n3864;
    wire n3868;
    wire n3871;
    wire n3875;
    wire n3879;
    wire n3883;
    wire n3887;
    wire n3891;
    wire n3895;
    wire n3899;
    wire n3903;
    wire n3907;
    wire n3911;
    wire n3915;
    wire n3919;
    wire n3923;
    wire n3927;
    wire n3931;
    wire n3935;
    wire n3939;
    wire n3943;
    wire n3946;
    wire n3950;
    wire n3954;
    wire n3958;
    wire n3962;
    wire n3966;
    wire n3970;
    wire n3974;
    wire n3978;
    wire n3982;
    wire n3986;
    wire n3990;
    wire n3993;
    wire n3996;
    wire n4000;
    wire n4004;
    wire n4007;
    wire n4011;
    wire n4015;
    wire n4019;
    wire n4023;
    wire n4026;
    wire n4030;
    wire n4033;
    wire n4037;
    wire n4041;
    wire n4045;
    wire n4049;
    wire n4053;
    wire n4057;
    wire n4061;
    wire n4065;
    wire n4069;
    wire n4073;
    wire n4077;
    wire n4081;
    wire n4084;
    wire n4088;
    wire n4092;
    wire n4095;
    wire n4099;
    wire n4103;
    wire n4107;
    wire n4111;
    wire n4115;
    wire n4119;
    wire n4123;
    wire n4127;
    wire n4131;
    wire n4135;
    wire n4138;
    wire n4142;
    wire n4146;
    wire n4149;
    wire n4153;
    wire n4157;
    wire n4161;
    wire n4165;
    wire n4169;
    wire n4172;
    wire n4175;
    wire n4179;
    wire n4182;
    wire n4185;
    wire n4189;
    wire n4193;
    wire n4197;
    wire n4201;
    wire n4205;
    wire n4209;
    wire n4213;
    wire n4216;
    wire n4220;
    wire n4223;
    wire n4227;
    wire n4231;
    wire n4234;
    wire n4238;
    wire n4241;
    wire n4245;
    wire n4249;
    wire n4253;
    wire n4256;
    wire n4260;
    wire n4264;
    wire n4268;
    wire n4272;
    wire n4276;
    wire n4280;
    wire n4283;
    wire n4287;
    wire n4291;
    wire n4294;
    wire n4298;
    wire n4302;
    wire n4306;
    wire n4310;
    wire n4314;
    wire n4317;
    wire n4321;
    wire n4325;
    wire n4329;
    wire n4333;
    wire n4336;
    wire n4340;
    wire n4343;
    wire n4347;
    wire n4351;
    wire n4355;
    wire n4358;
    wire n4362;
    wire n4365;
    wire n4369;
    wire n4373;
    wire n4376;
    wire n4380;
    wire n4384;
    wire n4388;
    wire n4392;
    wire n4396;
    wire n4399;
    wire n4403;
    wire n4407;
    wire n4410;
    wire n4414;
    wire n4418;
    wire n4422;
    wire n4426;
    wire n4430;
    wire n4434;
    wire n4438;
    wire n4442;
    wire n4446;
    wire n4449;
    wire n4452;
    wire n4455;
    wire n4458;
    wire n4462;
    wire n4466;
    wire n4470;
    wire n4474;
    wire n4478;
    wire n4482;
    wire n4486;
    wire n4489;
    wire n4492;
    wire n4496;
    wire n4500;
    wire n4504;
    wire n4508;
    wire n4512;
    wire n4516;
    wire n4519;
    wire n4522;
    wire n4525;
    wire n4528;
    wire n4532;
    wire n4536;
    wire n4540;
    wire n4544;
    wire n4548;
    wire n4551;
    wire n4555;
    wire n4559;
    wire n4562;
    wire n4566;
    wire n4570;
    wire n4574;
    wire n4578;
    wire n4582;
    wire n4586;
    wire n4590;
    wire n4594;
    wire n4598;
    wire n4602;
    wire n4606;
    wire n4609;
    wire n4612;
    wire n4616;
    wire n4620;
    wire n4624;
    wire n4628;
    wire n4632;
    wire n4635;
    wire n4639;
    wire n4643;
    wire n4646;
    wire n4650;
    wire n4654;
    wire n4658;
    wire n4662;
    wire n4666;
    wire n4669;
    wire n4672;
    wire n4676;
    wire n4680;
    wire n4683;
    wire n4687;
    wire n4691;
    wire n4695;
    wire n4698;
    wire n4701;
    wire n4704;
    wire n4707;
    wire n4711;
    wire n4715;
    wire n4719;
    wire n4723;
    wire n4727;
    wire n4731;
    wire n4735;
    wire n4739;
    wire n4743;
    wire n4747;
    wire n4750;
    wire n4754;
    wire n4758;
    wire n4762;
    wire n4766;
    wire n4770;
    wire n4774;
    wire n4778;
    wire n4782;
    wire n4786;
    wire n4789;
    wire n4793;
    wire n4796;
    wire n4800;
    wire n4804;
    wire n4808;
    wire n4812;
    wire n4816;
    wire n4820;
    wire n4823;
    wire n4826;
    wire n4830;
    wire n4834;
    wire n4838;
    wire n4842;
    wire n4846;
    wire n4850;
    wire n4854;
    wire n4858;
    wire n4861;
    wire n4865;
    wire n4869;
    wire n4873;
    wire n4877;
    wire n4881;
    wire n4885;
    wire n4889;
    wire n4893;
    wire n4896;
    wire n4900;
    wire n4904;
    wire n4908;
    wire n4912;
    wire n4916;
    wire n4920;
    wire n4924;
    wire n4928;
    wire n4932;
    wire n4936;
    wire n4940;
    wire n4944;
    wire n4948;
    wire n4952;
    wire n4956;
    wire n4960;
    wire n4963;
    wire n4967;
    wire n4970;
    wire n4974;
    wire n4978;
    wire n4982;
    wire n4986;
    wire n4990;
    wire n4994;
    wire n4998;
    wire n5002;
    wire n5006;
    wire n5010;
    wire n5014;
    wire n5017;
    wire n5021;
    wire n5025;
    wire n5029;
    wire n5033;
    wire n5037;
    wire n5041;
    wire n5045;
    wire n5049;
    wire n5053;
    wire n5057;
    wire n5061;
    wire n5065;
    wire n5069;
    wire n5073;
    wire n5077;
    wire n5081;
    wire n5085;
    wire n5089;
    wire n5093;
    wire n5097;
    wire n5101;
    wire n5104;
    wire n5108;
    wire n5112;
    wire n5116;
    wire n5120;
    wire n5124;
    wire n5128;
    wire n5132;
    wire n5136;
    wire n5140;
    wire n5144;
    wire n5148;
    wire n5156;
    wire n5160;
    wire n5163;
    wire n5166;
    wire n5170;
    wire n5174;
    wire n5178;
    wire n5182;
    wire n5186;
    wire n5190;
    wire n5194;
    wire n5198;
    wire n5202;
    wire n5206;
    wire n5209;
    wire n5213;
    wire n5217;
    wire n5221;
    wire n5225;
    wire n5229;
    wire n5233;
    wire n5237;
    wire n5241;
    wire n5245;
    wire n5248;
    wire n5251;
    wire n5255;
    wire n5259;
    wire n5263;
    wire n5267;
    wire n5271;
    wire n5275;
    wire n5279;
    wire n5283;
    wire n5287;
    wire n5291;
    wire n5295;
    wire n5299;
    wire n5303;
    wire n5307;
    wire n5311;
    wire n5314;
    wire n5318;
    wire n5322;
    wire n5326;
    wire n5330;
    wire n5334;
    wire n5338;
    wire n5342;
    wire n5346;
    wire n5350;
    wire n5354;
    wire n5357;
    wire n5360;
    wire n5364;
    wire n5368;
    wire n5372;
    wire n5375;
    wire n5379;
    wire n5382;
    wire n5386;
    wire n5390;
    wire n5394;
    wire n5398;
    wire n5402;
    wire n5406;
    wire n5409;
    wire n5413;
    wire n5417;
    wire n5421;
    wire n5424;
    wire n5427;
    wire n5431;
    wire n5435;
    wire n5439;
    wire n5442;
    wire n5445;
    wire n5449;
    wire n5453;
    wire n5457;
    wire n5461;
    wire n5465;
    wire n5468;
    wire n5472;
    wire n5475;
    wire n5479;
    wire n5483;
    wire n5487;
    wire n5491;
    wire n5495;
    wire n5498;
    wire n5502;
    wire n5506;
    wire n5510;
    wire n5514;
    wire n5517;
    wire n5521;
    wire n5524;
    wire n5528;
    wire n5532;
    wire n5536;
    wire n5540;
    wire n5544;
    wire n5548;
    wire n5552;
    wire n5555;
    wire n5559;
    wire n5563;
    wire n5567;
    wire n5571;
    wire n5575;
    wire n5579;
    wire n5583;
    wire n5587;
    wire n5590;
    wire n5594;
    wire n5597;
    wire n5601;
    wire n5605;
    wire n5609;
    wire n5613;
    wire n5617;
    wire n5621;
    wire n5625;
    wire n5628;
    wire n5631;
    wire n5634;
    wire n5637;
    wire n5640;
    wire n5643;
    wire n5646;
    wire n5649;
    wire n5652;
    wire n5655;
    wire n5658;
    wire n5661;
    wire n5664;
    wire n5667;
    wire n5670;
    wire n5673;
    wire n5676;
    wire n5679;
    wire n5682;
    wire n5685;
    wire n5688;
    wire n5691;
    wire n5694;
    wire n5697;
    wire n5700;
    wire n5703;
    wire n5706;
    wire n5709;
    wire n5712;
    wire n5715;
    wire n5718;
    wire n5721;
    wire n5724;
    wire n5727;
    wire n5730;
    wire n5733;
    wire n5736;
    wire n5739;
    wire n5742;
    wire n5745;
    wire n5748;
    wire n5751;
    wire n5755;
    wire n5758;
    wire n5762;
    wire n5765;
    wire n5769;
    wire n5773;
    wire n5777;
    wire n5781;
    wire n5785;
    wire n5789;
    wire n5793;
    wire n8214;
    wire n8217;
    wire n8220;
    wire n8223;
    wire n8226;
    wire n8229;
    wire n8233;
    wire n8236;
    wire n8239;
    wire n8242;
    wire n8245;
    wire n8248;
    wire n8251;
    wire n8254;
    wire n8257;
    wire n8260;
    wire n8263;
    wire n8266;
    wire n8269;
    wire n8272;
    wire n8275;
    wire n8278;
    wire n8281;
    wire n8284;
    wire n8287;
    wire n8290;
    wire n8293;
    wire n8296;
    wire n8299;
    wire n8302;
    wire n8305;
    wire n8308;
    wire n8311;
    wire n8314;
    wire n8317;
    wire n8320;
    wire n8323;
    wire n8326;
    wire n8329;
    wire n8332;
    wire n8335;
    wire n8338;
    wire n8341;
    wire n8344;
    wire n8347;
    wire n8350;
    wire n8353;
    wire n8356;
    wire n8358;
    wire n8361;
    wire n8364;
    wire n8367;
    wire n8371;
    wire n8374;
    wire n8377;
    wire n8380;
    wire n8383;
    wire n8386;
    wire n8389;
    wire n8392;
    wire n8395;
    wire n8398;
    wire n8400;
    wire n8403;
    wire n8406;
    wire n8409;
    wire n8412;
    wire n8415;
    wire n8419;
    wire n8422;
    wire n8425;
    wire n8428;
    wire n8430;
    wire n8433;
    wire n8436;
    wire n8440;
    wire n8443;
    wire n8446;
    wire n8449;
    wire n8452;
    wire n8455;
    wire n8457;
    wire n8460;
    wire n8463;
    wire n8466;
    wire n8469;
    wire n8473;
    wire n8476;
    wire n8479;
    wire n8482;
    wire n8485;
    wire n8487;
    wire n8490;
    wire n8493;
    wire n8496;
    wire n8499;
    wire n8502;
    wire n8506;
    wire n8508;
    wire n8511;
    wire n8514;
    wire n8517;
    wire n8521;
    wire n8524;
    wire n8527;
    wire n8530;
    wire n8533;
    wire n8536;
    wire n8539;
    wire n8542;
    wire n8545;
    wire n8548;
    wire n8551;
    wire n8554;
    wire n8557;
    wire n8560;
    wire n8563;
    wire n8566;
    wire n8569;
    wire n8572;
    wire n8575;
    wire n8577;
    wire n8581;
    wire n8583;
    wire n8586;
    wire n8590;
    wire n8593;
    wire n8596;
    wire n8598;
    wire n8602;
    wire n8605;
    wire n8608;
    wire n8611;
    wire n8614;
    wire n8617;
    wire n8620;
    wire n8622;
    wire n8626;
    wire n8628;
    wire n8631;
    wire n8634;
    wire n8637;
    wire n8640;
    wire n8643;
    wire n8647;
    wire n8650;
    wire n8653;
    wire n8656;
    wire n8658;
    wire n8661;
    wire n8664;
    wire n8667;
    wire n8670;
    wire n8673;
    wire n8677;
    wire n8679;
    wire n8682;
    wire n8685;
    wire n8688;
    wire n8691;
    wire n8694;
    wire n8697;
    wire n8700;
    wire n8703;
    wire n8706;
    wire n8709;
    wire n8712;
    wire n8716;
    wire n8719;
    wire n8721;
    wire n8724;
    wire n8727;
    wire n8730;
    wire n8733;
    wire n8736;
    wire n8739;
    wire n8743;
    wire n8746;
    wire n8749;
    wire n8752;
    wire n8754;
    wire n8758;
    wire n8761;
    wire n8764;
    wire n8767;
    wire n8770;
    wire n8773;
    wire n8776;
    wire n8779;
    wire n8782;
    wire n8785;
    wire n8788;
    wire n8791;
    wire n8794;
    wire n8796;
    wire n8800;
    wire n8803;
    wire n8806;
    wire n8809;
    wire n8812;
    wire n8815;
    wire n8818;
    wire n8821;
    wire n8824;
    wire n8827;
    wire n8830;
    wire n8833;
    wire n8836;
    wire n8839;
    wire n8842;
    wire n8845;
    wire n8848;
    wire n8851;
    wire n8854;
    wire n8857;
    wire n8860;
    wire n8863;
    wire n8866;
    wire n8869;
    wire n8871;
    wire n8875;
    wire n8878;
    wire n8881;
    wire n8884;
    wire n8887;
    wire n8890;
    wire n8893;
    wire n8896;
    wire n8899;
    wire n8902;
    wire n8905;
    wire n8908;
    wire n8911;
    wire n8914;
    wire n8917;
    wire n8920;
    wire n8923;
    wire n8926;
    wire n8929;
    wire n8932;
    wire n8935;
    wire n8938;
    wire n8941;
    wire n8944;
    wire n8947;
    wire n8950;
    wire n8953;
    wire n8956;
    wire n8959;
    wire n8962;
    wire n8965;
    wire n8968;
    wire n8971;
    wire n8974;
    wire n8977;
    wire n8980;
    wire n8983;
    wire n8986;
    wire n8989;
    wire n8992;
    wire n8995;
    wire n8998;
    wire n9001;
    wire n9004;
    wire n9006;
    wire n9010;
    wire n9013;
    wire n9016;
    wire n9019;
    wire n9022;
    wire n9025;
    wire n9028;
    wire n9031;
    wire n9034;
    wire n9037;
    wire n9040;
    wire n9043;
    wire n9046;
    wire n9049;
    wire n9052;
    wire n9055;
    wire n9058;
    wire n9061;
    wire n9064;
    wire n9067;
    wire n9070;
    wire n9073;
    wire n9076;
    wire n9079;
    wire n9082;
    wire n9085;
    wire n9088;
    wire n9091;
    wire n9094;
    wire n9097;
    wire n9100;
    wire n9103;
    wire n9106;
    wire n9109;
    wire n9112;
    wire n9115;
    wire n9118;
    wire n9121;
    wire n9124;
    wire n9127;
    wire n9130;
    wire n9133;
    wire n9136;
    wire n9139;
    wire n9142;
    wire n9145;
    wire n9148;
    wire n9151;
    wire n9154;
    wire n9157;
    wire n9160;
    wire n9163;
    wire n9166;
    wire n9169;
    wire n9172;
    wire n9175;
    wire n9178;
    wire n9181;
    wire n9184;
    wire n9187;
    wire n9190;
    wire n9193;
    wire n9196;
    wire n9199;
    wire n9202;
    wire n9205;
    wire n9208;
    wire n9211;
    wire n9214;
    wire n9217;
    wire n9220;
    wire n9223;
    wire n9226;
    wire n9229;
    wire n9231;
    wire n9235;
    wire n9238;
    wire n9241;
    wire n9244;
    wire n9247;
    wire n9250;
    wire n9253;
    wire n9256;
    wire n9259;
    wire n9262;
    wire n9265;
    wire n9268;
    wire n9271;
    wire n9274;
    wire n9277;
    wire n9280;
    wire n9283;
    wire n9286;
    wire n9289;
    wire n9292;
    wire n9295;
    wire n9297;
    wire n9301;
    wire n9304;
    wire n9307;
    wire n9310;
    wire n9313;
    wire n9316;
    wire n9319;
    wire n9322;
    wire n9325;
    wire n9328;
    wire n9331;
    wire n9334;
    wire n9337;
    wire n9339;
    wire n9343;
    wire n9346;
    wire n9349;
    wire n9352;
    wire n9354;
    wire n9357;
    wire n9361;
    wire n9364;
    wire n9367;
    wire n9370;
    wire n9373;
    wire n9376;
    wire n9378;
    wire n9381;
    wire n9384;
    wire n9387;
    wire n9391;
    wire n9393;
    wire n9396;
    wire n9400;
    wire n9402;
    wire n9405;
    wire n9409;
    wire n9412;
    wire n9414;
    wire n9418;
    wire n9420;
    wire n9423;
    wire n9426;
    wire n9430;
    wire n9433;
    wire n9436;
    wire n9439;
    wire n9442;
    wire n9445;
    wire n9448;
    wire n9451;
    wire n9453;
    wire n9457;
    wire n9460;
    wire n9463;
    wire n9466;
    wire n9468;
    wire n9471;
    wire n9475;
    wire n9478;
    wire n9481;
    wire n9484;
    wire n9487;
    wire n9489;
    wire n9493;
    wire n9495;
    wire n9499;
    wire n9502;
    wire n9505;
    wire n9508;
    wire n9510;
    wire n9514;
    wire n9517;
    wire n9520;
    wire n9523;
    wire n9526;
    wire n9528;
    wire n9531;
    wire n9535;
    wire n9538;
    wire n9540;
    wire n9543;
    wire n9547;
    wire n9549;
    wire n9552;
    wire n9556;
    wire n9558;
    wire n9561;
    wire n9565;
    wire n9567;
    wire n9570;
    wire n9574;
    wire n9576;
    wire n9579;
    wire n9583;
    wire n9585;
    wire n9588;
    wire n9591;
    wire n9595;
    wire n9598;
    wire n9601;
    wire n9604;
    wire n9607;
    wire n9610;
    wire n9613;
    wire n9616;
    wire n9618;
    wire n9621;
    wire n9625;
    wire n9628;
    wire n9631;
    wire n9634;
    wire n9637;
    wire n9640;
    wire n9642;
    wire n9646;
    wire n9649;
    wire n9652;
    wire n9655;
    wire n9658;
    wire n9661;
    wire n9664;
    wire n9667;
    wire n9670;
    wire n9673;
    wire n9676;
    wire n9679;
    wire n9682;
    wire n9685;
    wire n9688;
    wire n9691;
    wire n9694;
    wire n9697;
    wire n9700;
    wire n9703;
    wire n9706;
    wire n9709;
    wire n9712;
    wire n9715;
    wire n9718;
    wire n9721;
    wire n9724;
    wire n9727;
    wire n9730;
    wire n9733;
    wire n9736;
    wire n9739;
    wire n9742;
    wire n9745;
    wire n9748;
    wire n9751;
    wire n9754;
    wire n9757;
    wire n9760;
    wire n9763;
    wire n9765;
    wire n9768;
    wire n9771;
    wire n9775;
    wire n9778;
    wire n9781;
    wire n9784;
    wire n9787;
    wire n9790;
    wire n9793;
    wire n9796;
    wire n9799;
    wire n9801;
    wire n9805;
    wire n9808;
    wire n9811;
    wire n9814;
    wire n9817;
    wire n9820;
    wire n9823;
    wire n9826;
    wire n9829;
    wire n9832;
    wire n9835;
    wire n9838;
    wire n9841;
    wire n9844;
    wire n9847;
    wire n9850;
    wire n9853;
    wire n9856;
    wire n9859;
    wire n9862;
    wire n9865;
    wire n9868;
    wire n9871;
    wire n9874;
    wire n9877;
    wire n9880;
    wire n9883;
    wire n9886;
    wire n9889;
    wire n9892;
    wire n9895;
    wire n9898;
    wire n9901;
    wire n9904;
    wire n9907;
    wire n9910;
    wire n9913;
    wire n9916;
    wire n9919;
    wire n9922;
    wire n9925;
    wire n9927;
    wire n9930;
    wire n9933;
    wire n9936;
    wire n9939;
    wire n9942;
    wire n9945;
    wire n9948;
    wire n9951;
    wire n9954;
    wire n9958;
    wire n9960;
    wire n9963;
    wire n9966;
    wire n9969;
    wire n9972;
    wire n9975;
    wire n9978;
    wire n9981;
    wire n9984;
    wire n9988;
    wire n9991;
    wire n9994;
    wire n9997;
    wire n10000;
    wire n10003;
    wire n10006;
    wire n10009;
    wire n10012;
    wire n10015;
    wire n10017;
    wire n10020;
    wire n10023;
    wire n10026;
    wire n10029;
    wire n10032;
    wire n10035;
    wire n10038;
    wire n10041;
    wire n10045;
    wire n10048;
    wire n10051;
    wire n10054;
    wire n10057;
    wire n10060;
    wire n10062;
    wire n10066;
    wire n10069;
    wire n10072;
    wire n10075;
    wire n10078;
    wire n10081;
    wire n10084;
    wire n10087;
    wire n10090;
    wire n10093;
    wire n10096;
    wire n10099;
    wire n10101;
    wire n10104;
    wire n10107;
    wire n10110;
    wire n10113;
    wire n10116;
    wire n10119;
    wire n10122;
    wire n10125;
    wire n10128;
    wire n10131;
    wire n10135;
    wire n10138;
    wire n10141;
    wire n10144;
    wire n10147;
    wire n10150;
    wire n10153;
    wire n10156;
    wire n10158;
    wire n10161;
    wire n10164;
    wire n10167;
    wire n10170;
    wire n10173;
    wire n10176;
    wire n10179;
    wire n10182;
    wire n10185;
    wire n10188;
    wire n10191;
    wire n10194;
    wire n10197;
    wire n10200;
    wire n10204;
    wire n10207;
    wire n10210;
    wire n10213;
    wire n10215;
    wire n10218;
    wire n10221;
    wire n10224;
    wire n10227;
    wire n10230;
    wire n10233;
    wire n10236;
    wire n10239;
    wire n10242;
    wire n10245;
    wire n10248;
    wire n10252;
    wire n10255;
    wire n10258;
    wire n10261;
    wire n10264;
    wire n10267;
    wire n10270;
    wire n10273;
    wire n10276;
    wire n10279;
    wire n10282;
    wire n10285;
    wire n10288;
    wire n10291;
    wire n10294;
    wire n10297;
    wire n10300;
    wire n10303;
    wire n10306;
    wire n10309;
    wire n10312;
    wire n10315;
    wire n10318;
    wire n10321;
    wire n10324;
    wire n10327;
    wire n10330;
    wire n10333;
    wire n10336;
    wire n10339;
    wire n10342;
    wire n10345;
    wire n10348;
    wire n10351;
    wire n10354;
    wire n10357;
    wire n10360;
    wire n10363;
    wire n10366;
    wire n10369;
    wire n10372;
    wire n10375;
    wire n10378;
    wire n10381;
    wire n10384;
    wire n10387;
    wire n10390;
    wire n10393;
    wire n10396;
    wire n10399;
    wire n10402;
    wire n10405;
    wire n10408;
    wire n10410;
    wire n10413;
    wire n10416;
    wire n10419;
    wire n10422;
    wire n10425;
    wire n10428;
    wire n10431;
    wire n10434;
    wire n10437;
    wire n10440;
    wire n10443;
    wire n10446;
    wire n10449;
    wire n10452;
    wire n10455;
    wire n10458;
    wire n10461;
    wire n10464;
    wire n10467;
    wire n10471;
    wire n10474;
    wire n10477;
    wire n10480;
    wire n10483;
    wire n10486;
    wire n10489;
    wire n10492;
    wire n10495;
    wire n10498;
    wire n10501;
    wire n10504;
    wire n10507;
    wire n10510;
    wire n10513;
    wire n10515;
    wire n10518;
    wire n10521;
    wire n10524;
    wire n10527;
    wire n10530;
    wire n10533;
    wire n10537;
    wire n10540;
    wire n10543;
    wire n10546;
    wire n10549;
    wire n10552;
    wire n10555;
    wire n10558;
    wire n10561;
    wire n10564;
    wire n10567;
    wire n10570;
    wire n10573;
    wire n10576;
    wire n10579;
    wire n10582;
    wire n10585;
    wire n10588;
    wire n10591;
    wire n10594;
    wire n10597;
    wire n10600;
    wire n10603;
    wire n10606;
    wire n10609;
    wire n10612;
    wire n10615;
    wire n10618;
    wire n10621;
    wire n10624;
    wire n10627;
    wire n10630;
    wire n10633;
    wire n10636;
    wire n10639;
    wire n10642;
    wire n10645;
    wire n10648;
    wire n10651;
    wire n10654;
    wire n10657;
    wire n10660;
    wire n10663;
    wire n10665;
    wire n10668;
    wire n10671;
    wire n10674;
    wire n10677;
    wire n10680;
    wire n10683;
    wire n10686;
    wire n10689;
    wire n10692;
    wire n10695;
    wire n10698;
    wire n10701;
    wire n10704;
    wire n10707;
    wire n10710;
    wire n10713;
    wire n10716;
    wire n10719;
    wire n10722;
    wire n10725;
    wire n10728;
    wire n10731;
    wire n10734;
    wire n10738;
    wire n10741;
    wire n10744;
    wire n10747;
    wire n10750;
    wire n10753;
    wire n10756;
    wire n10759;
    wire n10762;
    wire n10765;
    wire n10768;
    wire n10771;
    wire n10774;
    wire n10777;
    wire n10780;
    wire n10783;
    wire n10786;
    wire n10789;
    wire n10792;
    wire n10794;
    wire n10797;
    wire n10800;
    wire n10803;
    wire n10806;
    wire n10809;
    wire n10812;
    wire n10815;
    wire n10818;
    wire n10821;
    wire n10824;
    wire n10828;
    wire n10831;
    wire n10834;
    wire n10837;
    wire n10840;
    wire n10843;
    wire n10846;
    wire n10849;
    wire n10852;
    wire n10855;
    wire n10857;
    wire n10860;
    wire n10863;
    wire n10866;
    wire n10869;
    wire n10872;
    wire n10875;
    wire n10878;
    wire n10881;
    wire n10884;
    wire n10887;
    wire n10890;
    wire n10893;
    wire n10896;
    wire n10899;
    wire n10902;
    wire n10905;
    wire n10908;
    wire n10911;
    wire n10914;
    wire n10917;
    wire n10920;
    wire n10923;
    wire n10926;
    wire n10929;
    wire n10932;
    wire n10935;
    wire n10938;
    wire n10941;
    wire n10944;
    wire n10947;
    wire n10951;
    wire n10954;
    wire n10957;
    wire n10960;
    wire n10963;
    wire n10965;
    wire n10968;
    wire n10971;
    wire n10974;
    wire n10977;
    wire n10981;
    wire n10984;
    wire n10987;
    wire n10990;
    wire n10993;
    wire n10996;
    wire n10999;
    wire n11002;
    wire n11005;
    wire n11008;
    wire n11011;
    wire n11014;
    wire n11016;
    wire n11019;
    wire n11022;
    wire n11025;
    wire n11028;
    wire n11031;
    wire n11034;
    wire n11037;
    wire n11040;
    wire n11043;
    wire n11046;
    wire n11049;
    wire n11052;
    wire n11055;
    wire n11058;
    wire n11061;
    wire n11064;
    wire n11067;
    wire n11070;
    wire n11073;
    wire n11076;
    wire n11079;
    wire n11082;
    wire n11085;
    wire n11088;
    wire n11091;
    wire n11094;
    wire n11097;
    wire n11100;
    wire n11103;
    wire n11106;
    wire n11109;
    wire n11112;
    wire n11115;
    wire n11118;
    wire n11121;
    wire n11124;
    wire n11127;
    wire n11130;
    wire n11133;
    wire n11137;
    wire n11140;
    wire n11143;
    wire n11145;
    wire n11148;
    wire n11151;
    wire n11154;
    wire n11157;
    wire n11160;
    wire n11163;
    wire n11166;
    wire n11169;
    wire n11172;
    wire n11175;
    wire n11178;
    wire n11181;
    wire n11184;
    wire n11187;
    wire n11190;
    wire n11193;
    wire n11196;
    wire n11199;
    wire n11202;
    wire n11205;
    wire n11208;
    wire n11211;
    wire n11214;
    wire n11217;
    wire n11220;
    wire n11223;
    wire n11226;
    wire n11229;
    wire n11232;
    wire n11235;
    wire n11238;
    wire n11241;
    wire n11245;
    wire n11248;
    wire n11251;
    wire n11253;
    wire n11256;
    wire n11259;
    wire n11262;
    wire n11265;
    wire n11268;
    wire n11272;
    wire n11275;
    wire n11278;
    wire n11280;
    wire n11283;
    wire n11286;
    wire n11289;
    wire n11293;
    wire n11296;
    wire n11299;
    wire n11301;
    wire n11304;
    wire n11308;
    wire n11311;
    wire n11314;
    wire n11316;
    wire n11319;
    wire n11322;
    wire n11325;
    wire n11328;
    wire n11331;
    wire n11334;
    wire n11337;
    wire n11340;
    wire n11344;
    wire n11347;
    wire n11350;
    wire n11353;
    wire n11356;
    wire n11359;
    wire n11361;
    wire n11364;
    wire n11367;
    wire n11370;
    wire n11373;
    wire n11376;
    wire n11379;
    wire n11382;
    wire n11385;
    wire n11388;
    wire n11391;
    wire n11394;
    wire n11397;
    wire n11400;
    wire n11403;
    wire n11406;
    wire n11409;
    wire n11412;
    wire n11415;
    wire n11418;
    wire n11421;
    wire n11424;
    wire n11427;
    wire n11430;
    wire n11433;
    wire n11436;
    wire n11439;
    wire n11442;
    wire n11445;
    wire n11448;
    wire n11452;
    wire n11454;
    wire n11457;
    wire n11460;
    wire n11463;
    wire n11466;
    wire n11469;
    wire n11472;
    wire n11475;
    wire n11478;
    wire n11481;
    wire n11484;
    wire n11487;
    wire n11490;
    wire n11493;
    wire n11496;
    wire n11499;
    wire n11502;
    wire n11505;
    wire n11508;
    wire n11511;
    wire n11514;
    wire n11517;
    wire n11520;
    wire n11523;
    wire n11526;
    wire n11529;
    wire n11532;
    wire n11535;
    wire n11538;
    wire n11541;
    wire n11545;
    wire n11548;
    wire n11550;
    wire n11553;
    wire n11556;
    wire n11559;
    wire n11562;
    wire n11566;
    wire n11569;
    wire n11572;
    wire n11575;
    wire n11578;
    wire n11581;
    wire n11584;
    wire n11587;
    wire n11590;
    wire n11593;
    wire n11596;
    wire n11598;
    wire n11601;
    wire n11604;
    wire n11607;
    wire n11610;
    wire n11613;
    wire n11616;
    wire n11619;
    wire n11622;
    wire n11625;
    wire n11628;
    wire n11631;
    wire n11634;
    wire n11637;
    wire n11640;
    wire n11644;
    wire n11647;
    wire n11650;
    wire n11652;
    wire n11655;
    wire n11658;
    wire n11661;
    wire n11664;
    wire n11667;
    wire n11671;
    wire n11674;
    wire n11677;
    wire n11679;
    wire n11682;
    wire n11685;
    wire n11688;
    wire n11691;
    wire n11694;
    wire n11697;
    wire n11700;
    wire n11703;
    wire n11706;
    wire n11709;
    wire n11712;
    wire n11715;
    wire n11718;
    wire n11721;
    wire n11724;
    wire n11727;
    wire n11730;
    wire n11733;
    wire n11736;
    wire n11740;
    wire n11742;
    wire n11745;
    wire n11748;
    wire n11751;
    wire n11754;
    wire n11757;
    wire n11760;
    wire n11763;
    wire n11766;
    wire n11769;
    wire n11772;
    wire n11775;
    wire n11778;
    wire n11781;
    wire n11784;
    wire n11787;
    wire n11790;
    wire n11793;
    wire n11796;
    wire n11799;
    wire n11802;
    wire n11805;
    wire n11808;
    wire n11811;
    wire n11814;
    wire n11817;
    wire n11821;
    wire n11824;
    wire n11827;
    wire n11829;
    wire n11832;
    wire n11835;
    wire n11838;
    wire n11841;
    wire n11845;
    wire n11848;
    wire n11851;
    wire n11854;
    wire n11857;
    wire n11860;
    wire n11863;
    wire n11866;
    wire n11869;
    wire n11872;
    wire n11875;
    wire n11877;
    wire n11880;
    wire n11883;
    wire n11886;
    wire n11889;
    wire n11892;
    wire n11895;
    wire n11898;
    wire n11901;
    wire n11905;
    wire n11908;
    wire n11911;
    wire n11914;
    wire n11917;
    wire n11920;
    wire n11923;
    wire n11925;
    wire n11928;
    wire n11931;
    wire n11934;
    wire n11937;
    wire n11940;
    wire n11943;
    wire n11946;
    wire n11949;
    wire n11952;
    wire n11955;
    wire n11958;
    wire n11961;
    wire n11964;
    wire n11967;
    wire n11970;
    wire n11973;
    wire n11976;
    wire n11979;
    wire n11982;
    wire n11985;
    wire n11988;
    wire n11991;
    wire n11994;
    wire n11997;
    wire n12000;
    wire n12003;
    wire n12006;
    wire n12009;
    wire n12012;
    wire n12015;
    wire n12018;
    wire n12021;
    wire n12024;
    wire n12027;
    wire n12030;
    wire n12034;
    wire n12037;
    wire n12040;
    wire n12043;
    wire n12046;
    wire n12049;
    wire n12052;
    wire n12055;
    wire n12057;
    wire n12060;
    wire n12063;
    wire n12066;
    wire n12069;
    wire n12072;
    wire n12075;
    wire n12078;
    wire n12081;
    wire n12084;
    wire n12088;
    wire n12091;
    wire n12094;
    wire n12097;
    wire n12099;
    wire n12102;
    wire n12105;
    wire n12108;
    wire n12112;
    wire n12115;
    wire n12118;
    wire n12121;
    wire n12123;
    wire n12126;
    wire n12129;
    wire n12132;
    wire n12135;
    wire n12138;
    wire n12141;
    wire n12144;
    wire n12147;
    wire n12150;
    wire n12153;
    wire n12156;
    wire n12159;
    wire n12162;
    wire n12165;
    wire n12168;
    wire n12171;
    wire n12174;
    wire n12177;
    wire n12180;
    wire n12183;
    wire n12186;
    wire n12189;
    wire n12192;
    wire n12195;
    wire n12198;
    wire n12201;
    wire n12204;
    wire n12207;
    wire n12210;
    wire n12213;
    wire n12216;
    wire n12220;
    wire n12223;
    wire n12226;
    wire n12229;
    wire n12231;
    wire n12234;
    wire n12237;
    wire n12240;
    wire n12243;
    wire n12246;
    wire n12249;
    wire n12252;
    wire n12255;
    wire n12258;
    wire n12261;
    wire n12264;
    wire n12267;
    wire n12270;
    wire n12273;
    wire n12277;
    wire n12280;
    wire n12283;
    wire n12286;
    wire n12288;
    wire n12291;
    wire n12294;
    wire n12297;
    wire n12300;
    wire n12303;
    wire n12307;
    wire n12309;
    wire n12312;
    wire n12315;
    wire n12318;
    wire n12322;
    wire n12325;
    wire n12327;
    wire n12330;
    wire n12333;
    wire n12336;
    wire n12340;
    wire n12343;
    wire n12346;
    wire n12349;
    wire n12351;
    wire n12354;
    wire n12357;
    wire n12360;
    wire n12363;
    wire n12367;
    wire n12370;
    wire n12373;
    wire n12376;
    wire n12379;
    wire n12382;
    wire n12385;
    wire n12388;
    wire n12391;
    wire n12394;
    wire n12397;
    wire n12400;
    wire n12403;
    wire n12406;
    wire n12408;
    wire n12411;
    wire n12414;
    wire n12417;
    wire n12420;
    wire n12423;
    wire n12426;
    wire n12429;
    wire n12432;
    wire n12435;
    wire n12438;
    wire n12441;
    wire n12444;
    wire n12447;
    wire n12450;
    wire n12453;
    wire n12456;
    wire n12459;
    wire n12462;
    wire n12465;
    wire n12468;
    wire n12471;
    wire n12474;
    wire n12477;
    wire n12480;
    wire n12483;
    wire n12486;
    wire n12489;
    wire n12492;
    wire n12495;
    wire n12498;
    wire n12501;
    wire n12504;
    wire n12507;
    wire n12510;
    wire n12513;
    wire n12516;
    wire n12519;
    wire n12522;
    wire n12525;
    wire n12528;
    wire n12531;
    wire n12534;
    wire n12537;
    wire n12540;
    wire n12543;
    wire n12546;
    wire n12549;
    wire n12552;
    wire n12555;
    wire n12558;
    wire n12561;
    wire n12564;
    wire n12567;
    wire n12570;
    wire n12573;
    wire n12576;
    wire n12579;
    wire n12582;
    wire n12585;
    wire n12588;
    wire n12591;
    wire n12594;
    wire n12597;
    wire n12600;
    wire n12603;
    wire n12606;
    wire n12609;
    wire n12612;
    wire n12615;
    wire n12619;
    wire n12621;
    wire n12624;
    wire n12627;
    wire n12630;
    wire n12633;
    wire n12636;
    wire n12639;
    wire n12642;
    wire n12645;
    wire n12648;
    wire n12651;
    wire n12654;
    wire n12657;
    wire n12660;
    wire n12663;
    wire n12666;
    wire n12669;
    wire n12672;
    wire n12675;
    wire n12678;
    wire n12681;
    wire n12684;
    wire n12687;
    wire n12690;
    wire n12693;
    wire n12696;
    wire n12699;
    wire n12702;
    wire n12706;
    wire n12709;
    wire n12712;
    wire n12715;
    wire n12718;
    wire n12721;
    wire n12724;
    wire n12727;
    wire n12730;
    wire n12733;
    wire n12736;
    wire n12739;
    wire n12742;
    wire n12745;
    wire n12748;
    wire n12751;
    wire n12754;
    wire n12757;
    wire n12760;
    wire n12763;
    wire n12766;
    wire n12769;
    wire n12772;
    wire n12775;
    wire n12778;
    wire n12781;
    wire n12784;
    wire n12787;
    wire n12790;
    wire n12793;
    wire n12796;
    wire n12799;
    wire n12802;
    wire n12805;
    wire n12807;
    wire n12810;
    wire n12813;
    wire n12816;
    wire n12819;
    wire n12822;
    wire n12825;
    wire n12828;
    wire n12831;
    wire n12834;
    wire n12837;
    wire n12841;
    wire n12844;
    wire n12847;
    wire n12850;
    wire n12853;
    wire n12856;
    wire n12859;
    wire n12861;
    wire n12864;
    wire n12867;
    wire n12870;
    wire n12873;
    wire n12876;
    wire n12879;
    wire n12882;
    wire n12885;
    wire n12888;
    wire n12891;
    wire n12894;
    wire n12898;
    wire n12901;
    wire n12904;
    wire n12907;
    wire n12910;
    wire n12913;
    wire n12916;
    wire n12919;
    wire n12922;
    wire n12925;
    wire n12928;
    wire n12931;
    wire n12934;
    wire n12937;
    wire n12940;
    wire n12943;
    wire n12945;
    wire n12948;
    wire n12951;
    wire n12954;
    wire n12957;
    wire n12960;
    wire n12963;
    wire n12966;
    wire n12969;
    wire n12972;
    wire n12975;
    wire n12979;
    wire n12982;
    wire n12985;
    wire n12988;
    wire n12991;
    wire n12994;
    wire n12997;
    wire n12999;
    wire n13002;
    wire n13005;
    wire n13008;
    wire n13011;
    wire n13014;
    wire n13017;
    wire n13020;
    wire n13023;
    wire n13026;
    wire n13029;
    wire n13032;
    wire n13035;
    wire n13038;
    wire n13041;
    wire n13044;
    wire n13047;
    wire n13050;
    wire n13053;
    wire n13056;
    wire n13059;
    wire n13062;
    wire n13066;
    wire n13069;
    wire n13072;
    wire n13075;
    wire n13078;
    wire n13080;
    wire n13084;
    wire n13087;
    wire n13089;
    wire n13092;
    wire n13095;
    wire n13098;
    wire n13101;
    wire n13104;
    wire n13107;
    wire n13110;
    wire n13113;
    wire n13116;
    wire n13119;
    wire n13122;
    wire n13125;
    wire n13128;
    wire n13131;
    wire n13134;
    wire n13137;
    wire n13140;
    wire n13143;
    wire n13146;
    wire n13150;
    wire n13153;
    wire n13155;
    wire n13158;
    wire n13161;
    wire n13164;
    wire n13167;
    wire n13170;
    wire n13173;
    wire n13176;
    wire n13179;
    wire n13182;
    wire n13185;
    wire n13188;
    wire n13192;
    wire n13195;
    wire n13198;
    wire n13200;
    wire n13203;
    wire n13206;
    wire n13209;
    wire n13212;
    wire n13215;
    wire n13218;
    wire n13221;
    wire n13224;
    wire n13227;
    wire n13230;
    wire n13233;
    wire n13236;
    wire n13239;
    wire n13242;
    wire n13245;
    wire n13248;
    wire n13252;
    wire n13255;
    wire n13257;
    wire n13260;
    wire n13263;
    wire n13266;
    wire n13269;
    wire n13272;
    wire n13275;
    wire n13278;
    wire n13281;
    wire n13285;
    wire n13288;
    wire n13291;
    wire n13294;
    wire n13297;
    wire n13300;
    wire n13303;
    wire n13306;
    wire n13309;
    wire n13312;
    wire n13315;
    wire n13317;
    wire n13320;
    wire n13323;
    wire n13326;
    wire n13329;
    wire n13333;
    wire n13336;
    wire n13339;
    wire n13341;
    wire n13344;
    wire n13347;
    wire n13350;
    wire n13353;
    wire n13356;
    wire n13359;
    wire n13362;
    wire n13365;
    wire n13368;
    wire n13371;
    wire n13374;
    wire n13377;
    wire n13380;
    wire n13383;
    wire n13387;
    wire n13389;
    wire n13392;
    wire n13396;
    wire n13399;
    wire n13402;
    wire n13405;
    wire n13408;
    wire n13411;
    wire n13414;
    wire n13416;
    wire n13419;
    wire n13422;
    wire n13425;
    wire n13428;
    wire n13431;
    wire n13434;
    wire n13437;
    wire n13440;
    wire n13443;
    wire n13446;
    wire n13449;
    wire n13452;
    wire n13455;
    wire n13458;
    wire n13461;
    wire n13464;
    wire n13467;
    wire n13470;
    wire n13473;
    wire n13476;
    wire n13479;
    wire n13482;
    wire n13485;
    wire n13488;
    wire n13492;
    wire n13495;
    wire n13497;
    wire n13500;
    wire n13503;
    wire n13506;
    wire n13509;
    wire n13512;
    wire n13515;
    wire n13518;
    wire n13521;
    wire n13524;
    wire n13527;
    wire n13530;
    wire n13533;
    wire n13536;
    wire n13539;
    wire n13542;
    wire n13546;
    wire n13549;
    wire n13552;
    wire n13555;
    wire n13557;
    wire n13560;
    wire n13563;
    wire n13566;
    wire n13569;
    wire n13572;
    wire n13575;
    wire n13579;
    wire n13582;
    wire n13585;
    wire n13588;
    wire n13590;
    wire n13593;
    wire n13596;
    wire n13599;
    wire n13602;
    wire n13605;
    wire n13608;
    wire n13611;
    wire n13614;
    wire n13617;
    wire n13620;
    wire n13623;
    wire n13626;
    wire n13629;
    wire n13632;
    wire n13635;
    wire n13638;
    wire n13641;
    wire n13644;
    wire n13647;
    wire n13650;
    wire n13654;
    wire n13657;
    wire n13659;
    wire n13662;
    wire n13665;
    wire n13668;
    wire n13671;
    wire n13674;
    wire n13677;
    wire n13680;
    wire n13683;
    wire n13687;
    wire n13690;
    wire n13692;
    wire n13695;
    wire n13698;
    wire n13701;
    wire n13704;
    wire n13707;
    wire n13711;
    wire n13714;
    wire n13717;
    wire n13720;
    wire n13722;
    wire n13725;
    wire n13728;
    wire n13731;
    wire n13734;
    wire n13737;
    wire n13740;
    wire n13743;
    wire n13746;
    wire n13749;
    wire n13752;
    wire n13755;
    wire n13758;
    wire n13761;
    wire n13764;
    wire n13767;
    wire n13770;
    wire n13773;
    wire n13777;
    wire n13780;
    wire n13783;
    wire n13786;
    wire n13788;
    wire n13791;
    wire n13794;
    wire n13797;
    wire n13801;
    wire n13804;
    wire n13807;
    wire n13810;
    wire n13813;
    wire n13816;
    wire n13819;
    wire n13822;
    wire n13825;
    wire n13828;
    wire n13831;
    wire n13834;
    wire n13837;
    wire n13840;
    wire n13843;
    wire n13846;
    wire n13849;
    wire n13852;
    wire n13855;
    wire n13858;
    wire n13861;
    wire n13864;
    wire n13867;
    wire n13870;
    wire n13873;
    wire n13876;
    wire n13879;
    wire n13882;
    wire n13885;
    wire n13888;
    wire n13891;
    wire n13894;
    wire n13897;
    wire n13900;
    wire n13903;
    wire n13906;
    wire n13909;
    wire n13911;
    wire n13914;
    wire n13917;
    wire n13920;
    wire n13924;
    wire n13926;
    wire n13929;
    wire n13932;
    wire n13936;
    wire n13939;
    wire n13942;
    wire n13945;
    wire n13947;
    wire n13950;
    wire n13953;
    wire n13957;
    wire n13960;
    wire n13963;
    wire n13966;
    wire n13968;
    wire n13971;
    wire n13974;
    wire n13977;
    wire n13981;
    wire n13984;
    wire n13987;
    wire n13990;
    wire n13993;
    wire n13996;
    wire n13999;
    wire n14002;
    wire n14005;
    wire n14008;
    wire n14010;
    wire n14013;
    wire n14016;
    wire n14019;
    wire n14023;
    wire n14025;
    wire n14028;
    wire n14031;
    wire n14034;
    wire n14037;
    wire n14040;
    wire n14043;
    wire n14046;
    wire n14049;
    wire n14052;
    wire n14055;
    wire n14058;
    wire n14062;
    wire n14064;
    wire n14067;
    wire n14070;
    wire n14073;
    wire n14076;
    wire n14080;
    wire n14082;
    wire n14085;
    wire n14088;
    wire n14091;
    wire n14094;
    wire n14097;
    wire n14101;
    wire n14104;
    wire n14107;
    wire n14110;
    wire n14112;
    wire n14115;
    wire n14118;
    wire n14121;
    wire n14124;
    wire n14127;
    wire n14130;
    wire n14133;
    wire n14136;
    wire n14139;
    wire n14142;
    wire n14145;
    wire n14149;
    wire n14151;
    wire n14154;
    wire n14158;
    wire n14160;
    wire n14163;
    wire n14166;
    wire n14169;
    wire n14172;
    wire n14175;
    wire n14178;
    wire n14181;
    wire n14184;
    wire n14187;
    wire n14190;
    wire n14193;
    wire n14196;
    wire n14199;
    wire n14202;
    wire n14205;
    wire n14208;
    wire n14211;
    wire n14214;
    wire n14217;
    wire n14220;
    wire n14223;
    wire n14226;
    wire n14229;
    wire n14232;
    wire n14235;
    wire n14238;
    wire n14241;
    wire n14244;
    wire n14248;
    wire n14250;
    wire n14253;
    wire n14256;
    wire n14259;
    wire n14262;
    wire n14265;
    wire n14268;
    wire n14271;
    wire n14274;
    wire n14277;
    wire n14280;
    wire n14283;
    wire n14286;
    wire n14289;
    wire n14292;
    wire n14296;
    wire n14299;
    wire n14301;
    wire n14304;
    wire n14307;
    wire n14310;
    wire n14313;
    wire n14316;
    wire n14319;
    wire n14322;
    wire n14325;
    wire n14328;
    wire n14331;
    wire n14335;
    wire n14337;
    wire n14340;
    wire n14343;
    wire n14346;
    wire n14349;
    wire n14352;
    wire n14355;
    wire n14358;
    wire n14361;
    wire n14364;
    wire n14367;
    wire n14370;
    wire n14373;
    wire n14376;
    wire n14379;
    wire n14382;
    wire n14385;
    wire n14388;
    wire n14391;
    wire n14395;
    wire n14398;
    wire n14401;
    wire n14404;
    wire n14406;
    wire n14409;
    wire n14412;
    wire n14415;
    wire n14418;
    wire n14421;
    wire n14424;
    wire n14427;
    wire n14430;
    wire n14433;
    wire n14436;
    wire n14439;
    wire n14442;
    wire n14445;
    wire n14448;
    wire n14451;
    wire n14454;
    wire n14457;
    wire n14460;
    wire n14463;
    wire n14466;
    wire n14469;
    wire n14472;
    wire n14475;
    wire n14478;
    wire n14481;
    wire n14484;
    wire n14487;
    wire n14490;
    wire n14493;
    wire n14496;
    wire n14499;
    wire n14502;
    wire n14505;
    wire n14508;
    wire n14511;
    wire n14514;
    wire n14517;
    wire n14520;
    wire n14523;
    wire n14526;
    wire n14529;
    wire n14532;
    wire n14535;
    wire n14538;
    wire n14541;
    wire n14544;
    wire n14547;
    wire n14550;
    wire n14553;
    wire n14556;
    wire n14559;
    wire n14562;
    wire n14565;
    wire n14568;
    wire n14571;
    wire n14574;
    wire n14577;
    wire n14580;
    wire n14583;
    wire n14586;
    wire n14589;
    wire n14592;
    wire n14595;
    wire n14598;
    wire n14601;
    wire n14604;
    wire n14607;
    wire n14610;
    wire n14613;
    wire n14616;
    wire n14619;
    wire n14622;
    wire n14625;
    wire n14628;
    wire n14631;
    wire n14634;
    wire n14637;
    wire n14640;
    wire n14643;
    wire n14646;
    wire n14649;
    wire n14652;
    wire n14655;
    wire n14658;
    wire n14661;
    wire n14664;
    wire n14667;
    wire n14670;
    wire n14673;
    wire n14677;
    wire n14680;
    wire n14683;
    wire n14686;
    wire n14689;
    wire n14691;
    wire n14694;
    wire n14697;
    wire n14700;
    wire n14703;
    wire n14706;
    wire n14709;
    wire n14712;
    wire n14715;
    wire n14718;
    wire n14721;
    wire n14724;
    wire n14727;
    wire n14730;
    wire n14733;
    wire n14736;
    wire n14739;
    wire n14742;
    wire n14745;
    wire n14749;
    wire n14751;
    wire n14754;
    wire n14757;
    wire n14760;
    wire n14763;
    wire n14766;
    wire n14769;
    wire n14772;
    wire n14775;
    wire n14778;
    wire n14781;
    wire n14784;
    wire n14787;
    wire n14790;
    wire n14793;
    wire n14796;
    wire n14799;
    wire n14802;
    wire n14805;
    wire n14808;
    wire n14811;
    wire n14815;
    wire n14818;
    wire n14821;
    wire n14823;
    wire n14826;
    wire n14829;
    wire n14832;
    wire n14835;
    wire n14838;
    wire n14841;
    wire n14844;
    wire n14847;
    wire n14850;
    wire n14853;
    wire n14856;
    wire n14859;
    wire n14862;
    wire n14865;
    wire n14868;
    wire n14871;
    wire n14874;
    wire n14877;
    wire n14881;
    wire n14883;
    wire n14886;
    wire n14889;
    wire n14892;
    wire n14895;
    wire n14898;
    wire n14901;
    wire n14904;
    wire n14907;
    wire n14910;
    wire n14913;
    wire n14916;
    wire n14919;
    wire n14922;
    wire n14925;
    wire n14928;
    wire n14932;
    wire n14935;
    wire n14938;
    wire n14940;
    wire n14943;
    wire n14946;
    wire n14949;
    wire n14952;
    wire n14955;
    wire n14958;
    wire n14961;
    wire n14964;
    wire n14967;
    wire n14970;
    wire n14973;
    wire n14976;
    wire n14979;
    wire n14983;
    wire n14986;
    wire n14988;
    wire n14991;
    wire n14994;
    wire n14997;
    wire n15000;
    wire n15003;
    wire n15006;
    wire n15009;
    wire n15012;
    wire n15015;
    wire n15018;
    wire n15021;
    wire n15024;
    wire n15027;
    wire n15030;
    wire n15033;
    wire n15036;
    wire n15039;
    wire n15042;
    wire n15045;
    wire n15048;
    wire n15051;
    wire n15054;
    wire n15057;
    wire n15060;
    wire n15063;
    wire n15066;
    wire n15069;
    wire n15072;
    wire n15075;
    wire n15081;
    wire n15084;
    wire n15087;
    wire n15090;
    wire n15093;
    wire n15096;
    wire n15099;
    wire n15102;
    wire n15105;
    wire n15108;
    wire n15111;
    wire n15114;
    wire n15117;
    wire n15120;
    wire n15123;
    wire n15126;
    wire n15129;
    wire n15132;
    wire n15135;
    wire n15138;
    wire n15141;
    wire n15144;
    wire n15147;
    wire n15150;
    wire n15153;
    wire n15159;
    wire n15162;
    wire n15165;
    wire n15168;
    wire n15171;
    wire n15174;
    wire n15177;
    wire n15180;
    wire n15183;
    wire n15186;
    wire n15189;
    wire n15192;
    wire n15195;
    wire n15198;
    wire n15201;
    wire n15204;
    wire n15207;
    wire n15210;
    wire n15213;
    wire n15216;
    wire n15219;
    wire n15222;
    wire n15225;
    wire n15228;
    wire n15231;
    wire n15237;
    wire n15240;
    wire n15243;
    wire n15246;
    wire n15249;
    wire n15252;
    wire n15255;
    wire n15258;
    wire n15261;
    wire n15264;
    wire n15267;
    wire n15270;
    wire n15273;
    wire n15276;
    wire n15279;
    wire n15282;
    wire n15285;
    wire n15288;
    wire n15291;
    wire n15294;
    wire n15297;
    wire n15300;
    wire n15303;
    wire n15306;
    wire n15309;
    wire n15315;
    wire n15318;
    wire n15321;
    wire n15324;
    wire n15327;
    wire n15330;
    wire n15333;
    wire n15336;
    wire n15339;
    wire n15342;
    wire n15345;
    wire n15348;
    wire n15351;
    wire n15354;
    wire n15357;
    wire n15360;
    wire n15363;
    wire n15366;
    wire n15369;
    wire n15372;
    wire n15375;
    wire n15378;
    wire n15381;
    wire n15384;
    wire n15387;
    wire n15393;
    wire n15396;
    wire n15399;
    wire n15402;
    wire n15405;
    wire n15408;
    wire n15411;
    wire n15414;
    wire n15417;
    wire n15420;
    wire n15423;
    wire n15426;
    wire n15429;
    wire n15432;
    wire n15435;
    wire n15438;
    wire n15441;
    wire n15444;
    wire n15447;
    wire n15450;
    wire n15453;
    wire n15456;
    wire n15459;
    wire n15462;
    wire n15465;
    wire n15471;
    wire n15474;
    wire n15477;
    wire n15480;
    wire n15483;
    wire n15486;
    wire n15489;
    wire n15492;
    wire n15495;
    wire n15498;
    wire n15501;
    wire n15504;
    wire n15507;
    wire n15510;
    wire n15513;
    wire n15516;
    wire n15519;
    wire n15522;
    wire n15525;
    wire n15528;
    wire n15531;
    wire n15534;
    wire n15537;
    wire n15540;
    wire n15543;
    wire n15549;
    wire n15552;
    wire n15555;
    wire n15558;
    wire n15561;
    wire n15564;
    wire n15567;
    wire n15570;
    wire n15573;
    wire n15576;
    wire n15579;
    wire n15582;
    wire n15585;
    wire n15588;
    wire n15591;
    wire n15594;
    wire n15597;
    wire n15600;
    wire n15603;
    wire n15606;
    wire n15609;
    wire n15612;
    wire n15615;
    wire n15618;
    wire n15621;
    wire n15627;
    wire n15630;
    wire n15633;
    wire n15636;
    wire n15639;
    wire n15642;
    wire n15645;
    wire n15648;
    wire n15651;
    wire n15654;
    wire n15657;
    wire n15660;
    wire n15663;
    wire n15666;
    wire n15669;
    wire n15672;
    wire n15675;
    wire n15678;
    wire n15681;
    wire n15684;
    wire n15687;
    wire n15690;
    wire n15693;
    wire n15696;
    wire n15699;
    wire n15705;
    wire n15708;
    wire n15711;
    wire n15714;
    wire n15717;
    wire n15720;
    wire n15723;
    wire n15726;
    wire n15729;
    wire n15732;
    wire n15735;
    wire n15738;
    wire n15741;
    wire n15744;
    wire n15747;
    wire n15750;
    wire n15753;
    wire n15756;
    wire n15759;
    wire n15762;
    wire n15765;
    wire n15768;
    wire n15771;
    wire n15774;
    wire n15777;
    wire n15783;
    wire n15786;
    wire n15789;
    wire n15792;
    wire n15795;
    wire n15798;
    wire n15801;
    wire n15804;
    wire n15807;
    wire n15810;
    wire n15813;
    wire n15816;
    wire n15819;
    wire n15822;
    wire n15825;
    wire n15828;
    wire n15831;
    wire n15834;
    wire n15837;
    wire n15840;
    wire n15843;
    wire n15846;
    wire n15849;
    wire n15852;
    wire n15855;
    wire n15861;
    wire n15864;
    wire n15867;
    wire n15870;
    wire n15873;
    wire n15876;
    wire n15879;
    wire n15882;
    wire n15885;
    wire n15888;
    wire n15891;
    wire n15894;
    wire n15897;
    wire n15900;
    wire n15903;
    wire n15906;
    wire n15909;
    wire n15912;
    wire n15915;
    wire n15918;
    wire n15921;
    wire n15924;
    wire n15927;
    wire n15930;
    wire n15933;
    wire n15939;
    wire n15942;
    wire n15945;
    wire n15948;
    wire n15951;
    wire n15954;
    wire n15957;
    wire n15960;
    wire n15963;
    wire n15966;
    wire n15969;
    wire n15972;
    wire n15975;
    wire n15978;
    wire n15981;
    wire n15984;
    wire n15987;
    wire n15990;
    wire n15993;
    wire n15996;
    wire n15999;
    wire n16002;
    wire n16005;
    wire n16008;
    wire n16011;
    wire n16017;
    wire n16020;
    wire n16023;
    wire n16026;
    wire n16029;
    wire n16032;
    wire n16035;
    wire n16038;
    wire n16041;
    wire n16044;
    wire n16047;
    wire n16050;
    wire n16053;
    wire n16056;
    wire n16059;
    wire n16062;
    wire n16065;
    wire n16068;
    wire n16071;
    wire n16074;
    wire n16077;
    wire n16080;
    wire n16083;
    wire n16086;
    wire n16089;
    wire n16095;
    wire n16098;
    wire n16101;
    wire n16104;
    wire n16107;
    wire n16110;
    wire n16113;
    wire n16116;
    wire n16119;
    wire n16122;
    wire n16125;
    wire n16128;
    wire n16131;
    wire n16134;
    wire n16137;
    wire n16140;
    wire n16143;
    wire n16146;
    wire n16149;
    wire n16152;
    wire n16155;
    wire n16158;
    wire n16161;
    wire n16164;
    wire n16167;
    wire n16173;
    wire n16176;
    wire n16179;
    wire n16182;
    wire n16185;
    wire n16188;
    wire n16191;
    wire n16194;
    wire n16197;
    wire n16200;
    wire n16203;
    wire n16206;
    wire n16209;
    wire n16212;
    wire n16215;
    wire n16218;
    wire n16221;
    wire n16224;
    wire n16227;
    wire n16230;
    wire n16233;
    wire n16236;
    wire n16239;
    wire n16242;
    wire n16245;
    wire n16251;
    wire n16254;
    wire n16257;
    wire n16260;
    wire n16263;
    wire n16266;
    wire n16269;
    wire n16272;
    wire n16275;
    wire n16278;
    wire n16281;
    wire n16284;
    wire n16287;
    wire n16290;
    wire n16293;
    wire n16296;
    wire n16299;
    wire n16302;
    wire n16305;
    wire n16308;
    wire n16311;
    wire n16314;
    wire n16317;
    wire n16320;
    wire n16323;
    wire n16329;
    wire n16332;
    wire n16335;
    wire n16338;
    wire n16341;
    wire n16344;
    wire n16347;
    wire n16350;
    wire n16353;
    wire n16356;
    wire n16359;
    wire n16362;
    wire n16365;
    wire n16368;
    wire n16371;
    wire n16374;
    wire n16377;
    wire n16380;
    wire n16383;
    wire n16386;
    wire n16389;
    wire n16392;
    wire n16395;
    wire n16398;
    wire n16401;
    wire n16407;
    wire n16410;
    wire n16413;
    wire n16416;
    wire n16419;
    wire n16422;
    wire n16425;
    wire n16428;
    wire n16431;
    wire n16434;
    wire n16437;
    wire n16440;
    wire n16443;
    wire n16446;
    wire n16449;
    wire n16452;
    wire n16455;
    wire n16458;
    wire n16461;
    wire n16464;
    wire n16467;
    wire n16470;
    wire n16473;
    wire n16476;
    wire n16479;
    wire n16485;
    wire n16488;
    wire n16491;
    wire n16494;
    wire n16497;
    wire n16500;
    wire n16503;
    wire n16506;
    wire n16509;
    wire n16512;
    wire n16515;
    wire n16518;
    wire n16521;
    wire n16524;
    wire n16527;
    wire n16530;
    wire n16533;
    wire n16536;
    wire n16539;
    wire n16542;
    wire n16545;
    wire n16548;
    wire n16551;
    wire n16554;
    wire n16557;
    wire n16563;
    wire n16566;
    wire n16569;
    wire n16572;
    wire n16575;
    wire n16578;
    wire n16581;
    wire n16584;
    wire n16587;
    wire n16590;
    wire n16593;
    wire n16596;
    wire n16599;
    wire n16602;
    wire n16605;
    wire n16608;
    wire n16611;
    wire n16614;
    wire n16617;
    wire n16620;
    wire n16623;
    wire n16626;
    wire n16629;
    wire n16632;
    wire n16635;
    wire n16641;
    wire n16644;
    wire n16647;
    wire n16650;
    wire n16653;
    wire n16656;
    wire n16659;
    wire n16662;
    wire n16665;
    wire n16668;
    wire n16671;
    wire n16674;
    wire n16677;
    wire n16680;
    wire n16683;
    wire n16686;
    wire n16689;
    wire n16692;
    wire n16695;
    wire n16698;
    wire n16701;
    wire n16704;
    wire n16707;
    wire n16710;
    wire n16713;
    wire n16719;
    wire n16722;
    wire n16725;
    wire n16728;
    wire n16731;
    wire n16734;
    wire n16737;
    wire n16740;
    wire n16743;
    wire n16746;
    wire n16749;
    wire n16752;
    wire n16755;
    wire n16758;
    wire n16761;
    wire n16764;
    wire n16767;
    wire n16770;
    wire n16773;
    wire n16776;
    wire n16779;
    wire n16782;
    wire n16785;
    wire n16788;
    wire n16791;
    wire n16797;
    wire n16800;
    wire n16803;
    wire n16806;
    wire n16809;
    wire n16812;
    wire n16815;
    wire n16818;
    wire n16821;
    wire n16824;
    wire n16827;
    wire n16830;
    wire n16833;
    wire n16836;
    wire n16839;
    wire n16842;
    wire n16845;
    wire n16848;
    wire n16851;
    wire n16854;
    wire n16857;
    wire n16860;
    wire n16863;
    wire n16866;
    wire n16869;
    wire n16875;
    wire n16878;
    wire n16881;
    wire n16884;
    wire n16887;
    wire n16890;
    wire n16893;
    wire n16896;
    wire n16899;
    wire n16902;
    wire n16905;
    wire n16908;
    wire n16911;
    wire n16914;
    wire n16917;
    wire n16920;
    wire n16923;
    wire n16926;
    wire n16929;
    wire n16932;
    wire n16935;
    wire n16938;
    wire n16941;
    wire n16944;
    wire n16947;
    wire n16953;
    wire n16956;
    wire n16959;
    wire n16962;
    wire n16965;
    wire n16968;
    wire n16971;
    wire n16974;
    wire n16977;
    wire n16980;
    wire n16983;
    wire n16986;
    wire n16989;
    wire n16992;
    wire n16995;
    wire n16998;
    wire n17001;
    wire n17004;
    wire n17007;
    wire n17010;
    wire n17013;
    wire n17016;
    wire n17019;
    wire n17022;
    wire n17025;
    wire n17031;
    wire n17034;
    wire n17037;
    wire n17040;
    wire n17043;
    wire n17046;
    wire n17049;
    wire n17052;
    wire n17055;
    wire n17058;
    wire n17061;
    wire n17064;
    wire n17067;
    wire n17070;
    wire n17073;
    wire n17076;
    wire n17079;
    wire n17082;
    wire n17085;
    wire n17088;
    wire n17091;
    wire n17094;
    wire n17097;
    wire n17100;
    wire n17103;
    wire n17109;
    wire n17112;
    wire n17115;
    wire n17118;
    wire n17121;
    wire n17124;
    wire n17127;
    wire n17130;
    wire n17133;
    wire n17136;
    wire n17139;
    wire n17142;
    wire n17145;
    wire n17148;
    wire n17151;
    wire n17154;
    wire n17157;
    wire n17160;
    wire n17163;
    wire n17166;
    wire n17169;
    wire n17172;
    wire n17175;
    wire n17178;
    wire n17181;
    wire n17187;
    wire n17190;
    wire n17193;
    wire n17196;
    wire n17199;
    wire n17202;
    wire n17205;
    wire n17208;
    wire n17211;
    wire n17214;
    wire n17217;
    wire n17220;
    wire n17223;
    wire n17226;
    wire n17229;
    wire n17232;
    wire n17235;
    wire n17238;
    wire n17241;
    wire n17244;
    wire n17247;
    wire n17250;
    wire n17253;
    wire n17256;
    wire n17259;
    wire n17265;
    wire n17268;
    wire n17271;
    wire n17274;
    wire n17277;
    wire n17280;
    wire n17283;
    wire n17286;
    wire n17289;
    wire n17292;
    wire n17295;
    wire n17298;
    wire n17301;
    wire n17304;
    wire n17307;
    wire n17310;
    wire n17313;
    wire n17316;
    wire n17319;
    wire n17322;
    wire n17325;
    wire n17328;
    wire n17331;
    wire n17334;
    wire n17337;
    wire n17343;
    wire n17346;
    wire n17349;
    wire n17352;
    wire n17355;
    wire n17358;
    wire n17361;
    wire n17364;
    wire n17367;
    wire n17370;
    wire n17373;
    wire n17376;
    wire n17379;
    wire n17382;
    wire n17385;
    wire n17388;
    wire n17391;
    wire n17394;
    wire n17397;
    wire n17400;
    wire n17403;
    wire n17406;
    wire n17409;
    wire n17412;
    wire n17415;
    wire n17421;
    wire n17424;
    wire n17427;
    wire n17430;
    wire n17433;
    wire n17436;
    wire n17439;
    wire n17442;
    wire n17445;
    wire n17448;
    wire n17451;
    wire n17454;
    wire n17457;
    wire n17460;
    wire n17463;
    wire n17466;
    wire n17469;
    wire n17472;
    wire n17475;
    wire n17478;
    wire n17481;
    wire n17484;
    wire n17487;
    wire n17490;
    wire n17493;
    wire n17499;
    wire n17502;
    wire n17505;
    wire n17508;
    wire n17511;
    wire n17514;
    wire n17517;
    wire n17520;
    wire n17523;
    wire n17526;
    wire n17529;
    wire n17532;
    wire n17535;
    wire n17538;
    wire n17541;
    wire n17544;
    wire n17547;
    wire n17550;
    wire n17553;
    wire n17556;
    wire n17559;
    wire n17562;
    wire n17565;
    wire n17568;
    wire n17571;
    wire n17577;
    wire n17580;
    wire n17583;
    wire n17586;
    wire n17589;
    wire n17592;
    wire n17595;
    wire n17598;
    wire n17601;
    wire n17604;
    wire n17607;
    wire n17610;
    wire n17613;
    wire n17616;
    wire n17619;
    wire n17622;
    wire n17625;
    wire n17628;
    wire n17631;
    wire n17634;
    wire n17637;
    wire n17640;
    wire n17643;
    wire n17646;
    wire n17649;
    wire n17655;
    wire n17658;
    wire n17661;
    wire n17664;
    wire n17667;
    wire n17670;
    wire n17673;
    wire n17676;
    wire n17679;
    wire n17682;
    wire n17685;
    wire n17688;
    wire n17691;
    wire n17694;
    wire n17697;
    wire n17700;
    wire n17703;
    wire n17706;
    wire n17709;
    wire n17712;
    wire n17715;
    wire n17718;
    wire n17721;
    wire n17724;
    wire n17727;
    wire n17733;
    wire n17736;
    wire n17739;
    wire n17742;
    wire n17745;
    wire n17748;
    wire n17751;
    wire n17754;
    wire n17757;
    wire n17760;
    wire n17763;
    wire n17766;
    wire n17769;
    wire n17772;
    wire n17775;
    wire n17778;
    wire n17781;
    wire n17784;
    wire n17787;
    wire n17790;
    wire n17793;
    wire n17796;
    wire n17799;
    wire n17802;
    wire n17805;
    wire n17811;
    wire n17814;
    wire n17817;
    wire n17820;
    wire n17823;
    wire n17826;
    wire n17829;
    wire n17832;
    wire n17835;
    wire n17838;
    wire n17841;
    wire n17844;
    wire n17847;
    wire n17850;
    wire n17853;
    wire n17856;
    wire n17859;
    wire n17862;
    wire n17865;
    wire n17868;
    wire n17871;
    wire n17874;
    wire n17877;
    wire n17880;
    wire n17883;
    wire n17889;
    wire n17892;
    wire n17895;
    wire n17898;
    wire n17901;
    wire n17904;
    wire n17907;
    wire n17910;
    wire n17913;
    wire n17916;
    wire n17919;
    wire n17922;
    wire n17925;
    wire n17928;
    wire n17931;
    wire n17934;
    wire n17937;
    wire n17940;
    wire n17943;
    wire n17946;
    wire n17949;
    wire n17952;
    wire n17955;
    wire n17958;
    wire n17961;
    wire n17967;
    wire n17970;
    wire n17973;
    wire n17976;
    wire n17979;
    wire n17982;
    wire n17985;
    wire n17988;
    wire n17991;
    wire n17994;
    wire n17997;
    wire n18000;
    wire n18003;
    wire n18006;
    wire n18009;
    wire n18012;
    wire n18015;
    wire n18018;
    wire n18021;
    wire n18024;
    wire n18027;
    wire n18030;
    wire n18033;
    wire n18036;
    wire n18039;
    wire n18045;
    wire n18048;
    wire n18051;
    wire n18054;
    wire n18057;
    wire n18060;
    wire n18063;
    wire n18066;
    wire n18069;
    wire n18072;
    wire n18075;
    wire n18078;
    wire n18081;
    wire n18084;
    wire n18087;
    wire n18090;
    wire n18093;
    wire n18096;
    wire n18099;
    wire n18102;
    wire n18105;
    wire n18108;
    wire n18111;
    wire n18114;
    wire n18117;
    wire n18123;
    wire n18126;
    wire n18129;
    wire n18132;
    wire n18135;
    wire n18138;
    wire n18141;
    wire n18144;
    wire n18147;
    wire n18150;
    wire n18153;
    wire n18156;
    wire n18159;
    wire n18162;
    wire n18165;
    wire n18168;
    wire n18171;
    wire n18174;
    wire n18177;
    wire n18180;
    wire n18183;
    wire n18186;
    wire n18189;
    wire n18192;
    wire n18195;
    wire n18201;
    wire n18204;
    wire n18207;
    wire n18210;
    wire n18213;
    wire n18216;
    wire n18219;
    wire n18222;
    wire n18225;
    wire n18228;
    wire n18231;
    wire n18234;
    wire n18237;
    wire n18240;
    wire n18243;
    wire n18246;
    wire n18249;
    wire n18252;
    wire n18255;
    wire n18258;
    wire n18261;
    wire n18264;
    wire n18267;
    wire n18273;
    wire n18276;
    wire n18279;
    wire n18282;
    wire n18285;
    wire n18288;
    wire n18291;
    wire n18294;
    wire n18297;
    wire n18300;
    wire n18303;
    wire n18306;
    wire n18309;
    wire n18312;
    wire n18315;
    wire n18318;
    wire n18321;
    wire n18324;
    wire n18327;
    wire n18330;
    wire n18333;
    wire n18336;
    wire n18339;
    wire n18345;
    wire n18348;
    wire n18351;
    wire n18354;
    wire n18357;
    wire n18360;
    wire n18363;
    wire n18366;
    wire n18369;
    wire n18372;
    wire n18375;
    wire n18378;
    wire n18381;
    wire n18384;
    wire n18387;
    wire n18390;
    wire n18393;
    wire n18396;
    wire n18399;
    wire n18402;
    wire n18405;
    wire n18408;
    wire n18411;
    wire n18417;
    wire n18420;
    wire n18423;
    wire n18426;
    wire n18429;
    wire n18432;
    wire n18435;
    wire n18438;
    wire n18441;
    wire n18444;
    wire n18447;
    wire n18450;
    wire n18453;
    wire n18456;
    wire n18459;
    wire n18462;
    wire n18465;
    wire n18468;
    wire n18471;
    wire n18474;
    wire n18477;
    wire n18480;
    wire n18483;
    wire n18489;
    wire n18492;
    wire n18495;
    wire n18498;
    wire n18501;
    wire n18504;
    wire n18507;
    wire n18510;
    wire n18513;
    wire n18516;
    wire n18519;
    wire n18522;
    wire n18525;
    wire n18528;
    wire n18531;
    wire n18534;
    wire n18537;
    wire n18540;
    wire n18543;
    wire n18546;
    wire n18549;
    wire n18552;
    wire n18555;
    wire n18558;
    wire n18561;
    wire n18567;
    wire n18570;
    wire n18573;
    wire n18576;
    wire n18579;
    wire n18582;
    wire n18585;
    wire n18588;
    wire n18591;
    wire n18594;
    wire n18597;
    wire n18600;
    wire n18603;
    wire n18606;
    wire n18609;
    wire n18612;
    wire n18615;
    wire n18618;
    wire n18621;
    wire n18624;
    wire n18627;
    wire n18630;
    wire n18633;
    wire n18636;
    wire n18639;
    wire n18645;
    wire n18648;
    wire n18651;
    wire n18654;
    wire n18657;
    wire n18660;
    wire n18663;
    wire n18666;
    wire n18669;
    wire n18672;
    wire n18675;
    wire n18678;
    wire n18681;
    wire n18684;
    wire n18687;
    wire n18690;
    wire n18693;
    wire n18696;
    wire n18699;
    wire n18702;
    wire n18705;
    wire n18708;
    wire n18711;
    wire n18714;
    wire n18720;
    wire n18723;
    wire n18726;
    wire n18729;
    wire n18732;
    wire n18735;
    wire n18738;
    wire n18741;
    wire n18744;
    wire n18747;
    wire n18750;
    wire n18753;
    wire n18756;
    wire n18759;
    wire n18762;
    wire n18765;
    wire n18768;
    wire n18771;
    wire n18774;
    wire n18777;
    wire n18780;
    wire n18783;
    wire n18786;
    wire n18789;
    wire n18792;
    wire n18798;
    wire n18801;
    wire n18804;
    wire n18807;
    wire n18810;
    wire n18813;
    wire n18816;
    wire n18819;
    wire n18822;
    wire n18825;
    wire n18828;
    wire n18831;
    wire n18834;
    wire n18837;
    wire n18840;
    wire n18843;
    wire n18846;
    wire n18849;
    wire n18852;
    wire n18855;
    wire n18858;
    wire n18861;
    wire n18864;
    wire n18867;
    wire n18873;
    wire n18876;
    wire n18879;
    wire n18882;
    wire n18885;
    wire n18888;
    wire n18891;
    wire n18894;
    wire n18897;
    wire n18900;
    wire n18903;
    wire n18906;
    wire n18909;
    wire n18912;
    wire n18915;
    wire n18918;
    wire n18921;
    wire n18924;
    wire n18927;
    wire n18930;
    wire n18933;
    wire n18936;
    wire n18939;
    wire n18945;
    wire n18948;
    wire n18951;
    wire n18954;
    wire n18957;
    wire n18960;
    wire n18963;
    wire n18966;
    wire n18969;
    wire n18972;
    wire n18975;
    wire n18978;
    wire n18981;
    wire n18984;
    wire n18987;
    wire n18990;
    wire n18993;
    wire n18996;
    wire n18999;
    wire n19002;
    wire n19005;
    wire n19008;
    wire n19011;
    wire n19014;
    wire n19017;
    wire n19023;
    wire n19026;
    wire n19029;
    wire n19032;
    wire n19035;
    wire n19038;
    wire n19041;
    wire n19044;
    wire n19047;
    wire n19050;
    wire n19053;
    wire n19056;
    wire n19059;
    wire n19062;
    wire n19065;
    wire n19068;
    wire n19071;
    wire n19074;
    wire n19077;
    wire n19080;
    wire n19083;
    wire n19086;
    wire n19089;
    wire n19095;
    wire n19098;
    wire n19101;
    wire n19104;
    wire n19107;
    wire n19110;
    wire n19113;
    wire n19116;
    wire n19119;
    wire n19122;
    wire n19125;
    wire n19128;
    wire n19131;
    wire n19134;
    wire n19137;
    wire n19140;
    wire n19143;
    wire n19146;
    wire n19149;
    wire n19152;
    wire n19155;
    wire n19158;
    wire n19161;
    wire n19164;
    wire n19167;
    wire n19173;
    wire n19176;
    wire n19179;
    wire n19182;
    wire n19185;
    wire n19188;
    wire n19191;
    wire n19194;
    wire n19197;
    wire n19200;
    wire n19203;
    wire n19206;
    wire n19209;
    wire n19212;
    wire n19215;
    wire n19218;
    wire n19221;
    wire n19224;
    wire n19227;
    wire n19230;
    wire n19233;
    wire n19236;
    wire n19239;
    wire n19242;
    wire n19245;
    wire n19251;
    wire n19254;
    wire n19257;
    wire n19260;
    wire n19263;
    wire n19266;
    wire n19269;
    wire n19272;
    wire n19275;
    wire n19278;
    wire n19281;
    wire n19284;
    wire n19287;
    wire n19290;
    wire n19293;
    wire n19296;
    wire n19299;
    wire n19302;
    wire n19305;
    wire n19308;
    wire n19317;
    wire n19320;
    wire n19323;
    wire n19326;
    wire n19329;
    wire n19332;
    wire n19338;
    wire n19341;
    wire n19344;
    wire n19347;
    wire n19350;
    wire n19353;
    wire n19362;
    wire n19365;
    wire n19368;
    wire n19371;
    wire n19374;
    wire n19377;
    wire n19380;
    wire n19383;
    wire n19386;
    wire n19389;
    wire n19392;
    wire n19395;
    wire n19398;
    wire n19401;
    wire n19407;
    wire n19410;
    wire n19413;
    wire n19416;
    wire n19419;
    wire n19422;
    wire n19425;
    wire n19428;
    wire n19431;
    wire n19434;
    wire n19437;
    wire n19440;
    wire n19443;
    wire n19446;
    wire n19449;
    wire n19452;
    wire n19458;
    wire n19461;
    wire n19464;
    wire n19467;
    wire n19470;
    wire n19473;
    wire n19476;
    wire n19479;
    wire n19482;
    wire n19485;
    wire n19488;
    wire n19491;
    wire n19494;
    wire n19497;
    wire n19500;
    wire n19503;
    wire n19506;
    wire n19512;
    wire n19515;
    wire n19518;
    wire n19521;
    wire n19524;
    wire n19527;
    wire n19530;
    wire n19533;
    wire n19536;
    wire n19539;
    wire n19542;
    wire n19545;
    wire n19548;
    wire n19551;
    wire n19554;
    wire n19557;
    wire n19560;
    wire n19563;
    wire n19569;
    wire n19572;
    wire n19575;
    wire n19578;
    wire n19581;
    wire n19584;
    wire n19587;
    wire n19590;
    wire n19593;
    wire n19596;
    wire n19599;
    wire n19602;
    wire n19608;
    wire n19611;
    wire n19614;
    wire n19617;
    wire n19620;
    wire n19623;
    wire n19626;
    wire n19629;
    wire n19632;
    wire n19635;
    wire n19638;
    wire n19641;
    wire n19644;
    wire n19650;
    wire n19653;
    wire n19656;
    wire n19659;
    wire n19662;
    wire n19665;
    wire n19668;
    wire n19671;
    wire n19674;
    wire n19677;
    wire n19680;
    wire n19683;
    wire n19686;
    wire n19692;
    wire n19695;
    wire n19698;
    wire n19701;
    wire n19704;
    wire n19707;
    wire n19710;
    wire n19713;
    wire n19716;
    wire n19719;
    wire n19722;
    wire n19725;
    wire n19728;
    wire n19731;
    wire n19734;
    wire n19740;
    wire n19743;
    wire n19746;
    wire n19749;
    wire n19752;
    wire n19755;
    wire n19758;
    wire n19761;
    wire n19764;
    wire n19767;
    wire n19770;
    wire n19773;
    wire n19776;
    wire n19779;
    wire n19782;
    wire n19788;
    wire n19791;
    wire n19794;
    wire n19797;
    wire n19800;
    wire n19803;
    wire n19806;
    wire n19809;
    wire n19812;
    wire n19815;
    wire n19818;
    wire n19821;
    wire n19824;
    wire n19827;
    wire n19830;
    wire n19836;
    wire n19839;
    wire n19842;
    wire n19845;
    wire n19848;
    wire n19851;
    wire n19854;
    wire n19857;
    wire n19860;
    wire n19863;
    wire n19866;
    wire n19869;
    wire n19872;
    wire n19878;
    wire n19881;
    wire n19884;
    wire n19887;
    wire n19890;
    wire n19893;
    wire n19899;
    wire n19902;
    wire n19905;
    wire n19908;
    wire n19911;
    wire n19914;
    wire n19917;
    wire n19920;
    wire n19923;
    wire n19929;
    wire n19932;
    wire n19935;
    wire n19938;
    wire n19941;
    wire n19947;
    wire n19950;
    wire n19953;
    wire n19956;
    wire n19959;
    wire n19962;
    wire n19965;
    wire n19968;
    wire n19971;
    wire n19980;
    wire n19983;
    wire n19986;
    wire n19989;
    wire n19992;
    wire n19998;
    wire n20001;
    wire n20004;
    wire n20007;
    wire n20010;
    wire n20013;
    wire n20019;
    wire n20022;
    wire n20025;
    wire n20028;
    wire n20031;
    wire n20034;
    wire n20037;
    wire n20043;
    wire n20046;
    wire n20049;
    wire n20052;
    wire n20055;
    wire n20058;
    wire n20061;
    wire n20067;
    wire n20073;
    wire n20076;
    wire n20082;
    wire n20085;
    wire n20088;
    wire n20094;
    wire n20097;
    wire n20100;
    wire n20106;
    wire n20109;
    wire n20112;
    wire n20115;
    wire n20118;
    wire n20121;
    wire n20124;
    wire n20127;
    wire n20130;
    wire n20133;
    wire n20136;
    wire n20145;
    wire n20148;
    wire n20151;
    wire n20157;
    wire n20160;
    wire n20163;
    wire n20166;
    wire n20169;
    wire n20175;
    wire n20178;
    wire n20181;
    wire n20184;
    wire n20187;
    wire n20193;
    wire n20196;
    wire n20199;
    wire n20202;
    wire n20205;
    wire n20208;
    wire n20211;
    wire n20217;
    wire n20220;
    wire n20223;
    wire n20226;
    wire n20229;
    wire n20232;
    wire n20235;
    wire n20238;
    wire n20241;
    wire n20244;
    wire n20247;
    wire n20250;
    wire n20253;
    wire n20265;
    wire n20268;
    wire n20271;
    wire n20277;
    wire n20280;
    wire n20283;
    wire n20289;
    wire n20292;
    wire n20295;
    wire n20298;
    wire n20301;
    wire n20304;
    wire n20307;
    wire n20310;
    wire n20313;
    wire n20319;
    wire n20322;
    wire n20325;
    wire n20328;
    wire n20331;
    wire n20334;
    wire n20337;
    wire n20340;
    wire n20343;
    wire n20346;
    wire n20352;
    wire n20355;
    wire n20358;
    wire n20361;
    wire n20364;
    wire n20367;
    wire n20370;
    wire n20373;
    wire n20376;
    wire n20379;
    wire n20382;
    wire n20388;
    wire n20391;
    wire n20394;
    wire n20397;
    wire n20400;
    wire n20403;
    wire n20406;
    wire n20409;
    wire n20412;
    wire n20415;
    wire n20418;
    wire n20424;
    wire n20427;
    wire n20430;
    wire n20433;
    wire n20436;
    wire n20439;
    wire n20442;
    wire n20445;
    wire n20451;
    wire n20454;
    wire n20457;
    wire n20460;
    wire n20463;
    wire n20466;
    wire n20469;
    wire n20472;
    wire n20475;
    wire n20481;
    wire n20484;
    wire n20487;
    wire n20490;
    wire n20493;
    wire n20496;
    wire n20499;
    wire n20502;
    wire n20505;
    wire n20511;
    wire n20514;
    wire n20517;
    wire n20520;
    wire n20523;
    wire n20526;
    wire n20529;
    wire n20532;
    wire n20535;
    wire n20538;
    wire n20541;
    wire n20547;
    wire n20550;
    wire n20553;
    wire n20556;
    wire n20562;
    wire n20565;
    wire n20568;
    wire n20571;
    wire n20574;
    wire n20577;
    wire n20583;
    wire n20586;
    wire n20589;
    wire n20592;
    jnot g0000(.din(G15), .dout(n316));
    jor g0001(.dinb(G5), .dina(G57), .dout(n320));
    jnot g0002(.din(G184), .dout(n323));
    jnot g0003(.din(G228), .dout(n326));
    jor g0004(.dinb(n323), .dina(n326), .dout(n330));
    jnot g0005(.din(G150), .dout(n333));
    jnot g0006(.din(G240), .dout(n336));
    jor g0007(.dinb(n333), .dina(n336), .dout(n340));
    jor g0008(.dinb(n330), .dina(n340), .dout(n344));
    jnot g0009(.din(G210), .dout(n347));
    jnot g0010(.din(G218), .dout(n350));
    jor g0011(.dinb(n347), .dina(n350), .dout(n354));
    jnot g0012(.din(G152), .dout(n357));
    jnot g0013(.din(G230), .dout(n360));
    jor g0014(.dinb(n357), .dina(n360), .dout(n364));
    jor g0015(.dinb(n354), .dina(n364), .dout(n368));
    jnot g0016(.din(G183), .dout(n371));
    jnot g0017(.din(G185), .dout(n374));
    jor g0018(.dinb(n371), .dina(n374), .dout(n378));
    jnot g0019(.din(G182), .dout(n381));
    jnot g0020(.din(G186), .dout(n384));
    jor g0021(.dinb(n381), .dina(n384), .dout(n388));
    jor g0022(.dinb(n378), .dina(n388), .dout(n392));
    jnot g0023(.din(G172), .dout(n395));
    jnot g0024(.din(G188), .dout(n398));
    jor g0025(.dinb(n395), .dina(n398), .dout(n402));
    jnot g0026(.din(G162), .dout(n405));
    jnot g0027(.din(G199), .dout(n408));
    jor g0028(.dinb(n405), .dina(n408), .dout(n412));
    jor g0029(.dinb(n402), .dina(n412), .dout(n416));
    jnot g0030(.din(G1197), .dout(n419));
    jor g0031(.dinb(n8220), .dina(n419), .dout(n423));
    jnot g0032(.din(G133), .dout(n426));
    jnot g0033(.din(G134), .dout(n429));
    jor g0034(.dinb(n426), .dina(n429), .dout(n433));
    jor g0035(.dinb(n8214), .dina(n433), .dout(n437));
    jand g0036(.dinb(G1), .dina(G163), .dout(n441));
    jnot g0037(.din(G41), .dout(n444));
    jor g0038(.dinb(n14940), .dina(n444), .dout(n448));
    jor g0039(.dinb(n14316), .dina(n448), .dout(n452));
    jnot g0040(.din(G18), .dout(n455));
    jand g0041(.dinb(n455), .dina(n14349), .dout(n459));
    jand g0042(.dinb(G18), .dina(G229), .dout(n463));
    jor g0043(.dinb(n459), .dina(n14062), .dout(n467));
    jand g0044(.dinb(n455), .dina(n14355), .dout(n471));
    jnot g0045(.din(n471), .dout(n474));
    jor g0046(.dinb(n467), .dina(n474), .dout(n478));
    jand g0047(.dinb(n14248), .dina(n478), .dout(n482));
    jxor g0048(.dinb(n14406), .dina(n482), .dout(n486));
    jand g0049(.dinb(G1496), .dina(G4528), .dout(n490));
    jxor g0050(.dinb(n12693), .dina(n490), .dout(n494));
    jnot g0051(.din(G3723), .dout(n497));
    jand g0052(.dinb(G18), .dina(G235), .dout(n501));
    jnot g0053(.din(n501), .dout(n504));
    jnot g0054(.din(G103), .dout(n507));
    jor g0055(.dinb(n14649), .dina(n507), .dout(n511));
    jand g0056(.dinb(n504), .dina(n511), .dout(n515));
    jxor g0057(.dinb(n14652), .dina(n515), .dout(n519));
    jand g0058(.dinb(G18), .dina(G236), .dout(n523));
    jnot g0059(.din(n523), .dout(n526));
    jnot g0060(.din(G23), .dout(n529));
    jor g0061(.dinb(n14991), .dina(n529), .dout(n533));
    jand g0062(.dinb(n526), .dina(n533), .dout(n537));
    jnot g0063(.din(n537), .dout(n540));
    jxor g0064(.dinb(n14571), .dina(n540), .dout(n544));
    jor g0065(.dinb(n14604), .dina(n544), .dout(n548));
    jnot g0066(.din(G3711), .dout(n551));
    jand g0067(.dinb(G18), .dina(G237), .dout(n555));
    jnot g0068(.din(n555), .dout(n558));
    jnot g0069(.din(G26), .dout(n561));
    jor g0070(.dinb(n14988), .dina(n561), .dout(n565));
    jand g0071(.dinb(n558), .dina(n565), .dout(n569));
    jxor g0072(.dinb(n14986), .dina(n569), .dout(n573));
    jnot g0073(.din(G4526), .dout(n576));
    jnot g0074(.din(G3701), .dout(n579));
    jand g0075(.dinb(n14352), .dina(n459), .dout(n583));
    jnot g0076(.din(G229), .dout(n586));
    jor g0077(.dinb(n455), .dina(n586), .dout(n590));
    jand g0078(.dinb(n448), .dina(n590), .dout(n594));
    jand g0079(.dinb(n594), .dina(n14313), .dout(n598));
    jor g0080(.dinb(n14335), .dina(n598), .dout(n602));
    jnot g0081(.din(G3705), .dout(n605));
    jnot g0082(.din(G238), .dout(n608));
    jor g0083(.dinb(n455), .dina(n608), .dout(n612));
    jnot g0084(.din(G29), .dout(n615));
    jor g0085(.dinb(n14826), .dina(n615), .dout(n619));
    jand g0086(.dinb(n612), .dina(n619), .dout(n623));
    jxor g0087(.dinb(n14299), .dina(n623), .dout(n627));
    jor g0088(.dinb(n602), .dina(n14256), .dout(n631));
    jor g0089(.dinb(n14391), .dina(n631), .dout(n635));
    jor g0090(.dinb(n14487), .dina(n635), .dout(n639));
    jor g0091(.dinb(n14499), .dina(n639), .dout(n643));
    jor g0092(.dinb(n14994), .dina(n569), .dout(n647));
    jor g0093(.dinb(n14248), .dina(n627), .dout(n651));
    jor g0094(.dinb(n14484), .dina(n651), .dout(n655));
    jand g0095(.dinb(n14250), .dina(n655), .dout(n659));
    jor g0096(.dinb(n14496), .dina(n659), .dout(n663));
    jor g0097(.dinb(n14301), .dina(n623), .dout(n667));
    jor g0098(.dinb(n573), .dina(n667), .dout(n671));
    jor g0099(.dinb(n548), .dina(n14202), .dout(n675));
    jor g0100(.dinb(n14658), .dina(n515), .dout(n679));
    jand g0101(.dinb(n14667), .dina(n515), .dout(n683));
    jor g0102(.dinb(n14574), .dina(n537), .dout(n687));
    jor g0103(.dinb(n683), .dina(n687), .dout(n691));
    jand g0104(.dinb(n14158), .dina(n691), .dout(n695));
    jand g0105(.dinb(n675), .dina(n14154), .dout(n699));
    jand g0106(.dinb(n663), .dina(n699), .dout(n703));
    jand g0107(.dinb(n643), .dina(n703), .dout(n707));
    jnot g0108(.din(G3737), .dout(n710));
    jand g0109(.dinb(G18), .dina(G233), .dout(n714));
    jnot g0110(.din(n714), .dout(n717));
    jnot g0111(.din(G127), .dout(n720));
    jor g0112(.dinb(n14823), .dina(n720), .dout(n724));
    jand g0113(.dinb(n717), .dina(n724), .dout(n728));
    jxor g0114(.dinb(n14818), .dina(n728), .dout(n732));
    jnot g0115(.din(G3729), .dout(n735));
    jand g0116(.dinb(G18), .dina(G234), .dout(n739));
    jnot g0117(.din(n739), .dout(n742));
    jnot g0118(.din(G130), .dout(n745));
    jor g0119(.dinb(n14895), .dina(n745), .dout(n749));
    jand g0120(.dinb(n742), .dina(n749), .dout(n753));
    jxor g0121(.dinb(n13677), .dina(n753), .dout(n757));
    jor g0122(.dinb(n732), .dina(n757), .dout(n761));
    jand g0123(.dinb(G18), .dina(G231), .dout(n765));
    jnot g0124(.din(n765), .dout(n768));
    jnot g0125(.din(G100), .dout(n771));
    jor g0126(.dinb(n14949), .dina(n771), .dout(n775));
    jand g0127(.dinb(n768), .dina(n775), .dout(n779));
    jor g0128(.dinb(n14898), .dina(n779), .dout(n783));
    jnot g0129(.din(n783), .dout(n786));
    jand g0130(.dinb(n14898), .dina(n779), .dout(n790));
    jor g0131(.dinb(n786), .dina(n14881), .dout(n794));
    jand g0132(.dinb(G18), .dina(G232), .dout(n798));
    jand g0133(.dinb(n455), .dina(n14938), .dout(n802));
    jor g0134(.dinb(n14935), .dina(n802), .dout(n806));
    jxor g0135(.dinb(n14958), .dina(n806), .dout(n810));
    jor g0136(.dinb(n794), .dina(n14928), .dout(n814));
    jor g0137(.dinb(n13657), .dina(n814), .dout(n818));
    jor g0138(.dinb(n707), .dina(n13617), .dout(n822));
    jnot g0139(.din(n806), .dout(n825));
    jor g0140(.dinb(n14955), .dina(n825), .dout(n829));
    jand g0141(.dinb(n14952), .dina(n825), .dout(n833));
    jor g0142(.dinb(n14829), .dina(n728), .dout(n837));
    jor g0143(.dinb(n14796), .dina(n753), .dout(n841));
    jor g0144(.dinb(n732), .dina(n841), .dout(n845));
    jand g0145(.dinb(n14821), .dina(n845), .dout(n849));
    jor g0146(.dinb(n14856), .dina(n849), .dout(n853));
    jand g0147(.dinb(n14751), .dina(n853), .dout(n857));
    jand g0148(.dinb(n14883), .dina(n857), .dout(n861));
    jor g0149(.dinb(n14868), .dina(n861), .dout(n865));
    jand g0150(.dinb(n822), .dina(n13614), .dout(n869));
    jnot g0151(.din(G4415), .dout(n872));
    jand g0152(.dinb(G18), .dina(G223), .dout(n876));
    jand g0153(.dinb(n455), .dina(n13582), .dout(n880));
    jor g0154(.dinb(n13579), .dina(n880), .dout(n884));
    jxor g0155(.dinb(n13588), .dina(n884), .dout(n888));
    jnot g0156(.din(G4400), .dout(n891));
    jand g0157(.dinb(G18), .dina(G226), .dout(n895));
    jand g0158(.dinb(n455), .dina(n13549), .dout(n899));
    jor g0159(.dinb(n13546), .dina(n899), .dout(n903));
    jxor g0160(.dinb(n13555), .dina(n903), .dout(n907));
    jand g0161(.dinb(G18), .dina(G217), .dout(n911));
    jand g0162(.dinb(n455), .dina(n13495), .dout(n915));
    jor g0163(.dinb(n13492), .dina(n915), .dout(n919));
    jnot g0164(.din(n919), .dout(n922));
    jxor g0165(.dinb(n13497), .dina(n922), .dout(n926));
    jand g0166(.dinb(n13509), .dina(n926), .dout(n930));
    jnot g0167(.din(G4410), .dout(n933));
    jand g0168(.dinb(G18), .dina(G224), .dout(n937));
    jand g0169(.dinb(n455), .dina(n13714), .dout(n941));
    jor g0170(.dinb(n13711), .dina(n941), .dout(n945));
    jxor g0171(.dinb(n13720), .dina(n945), .dout(n949));
    jand g0172(.dinb(G18), .dina(G225), .dout(n953));
    jand g0173(.dinb(n455), .dina(n13690), .dout(n957));
    jor g0174(.dinb(n13687), .dina(n957), .dout(n961));
    jnot g0175(.din(n961), .dout(n964));
    jxor g0176(.dinb(n13692), .dina(n964), .dout(n968));
    jand g0177(.dinb(n13707), .dina(n968), .dout(n972));
    jand g0178(.dinb(n930), .dina(n972), .dout(n976));
    jand g0179(.dinb(n13569), .dina(n976), .dout(n980));
    jnot g0180(.din(n980), .dout(n983));
    jor g0181(.dinb(n869), .dina(n13414), .dout(n987));
    jnot g0182(.din(n884), .dout(n990));
    jand g0183(.dinb(n13590), .dina(n990), .dout(n994));
    jand g0184(.dinb(n13588), .dina(n884), .dout(n998));
    jnot g0185(.din(n998), .dout(n1001));
    jand g0186(.dinb(n13720), .dina(n945), .dout(n1005));
    jnot g0187(.din(n1005), .dout(n1008));
    jnot g0188(.din(n945), .dout(n1011));
    jand g0189(.dinb(n13722), .dina(n1011), .dout(n1015));
    jand g0190(.dinb(n13692), .dina(n964), .dout(n1019));
    jnot g0191(.din(n907), .dout(n1022));
    jor g0192(.dinb(n13497), .dina(n922), .dout(n1026));
    jor g0193(.dinb(n1022), .dina(n1026), .dout(n1030));
    jand g0194(.dinb(n13555), .dina(n903), .dout(n1034));
    jnot g0195(.din(n1034), .dout(n1037));
    jor g0196(.dinb(n13692), .dina(n964), .dout(n1041));
    jand g0197(.dinb(n1037), .dina(n1041), .dout(n1045));
    jand g0198(.dinb(n1030), .dina(n1045), .dout(n1049));
    jor g0199(.dinb(n13383), .dina(n1049), .dout(n1053));
    jor g0200(.dinb(n13339), .dina(n1053), .dout(n1057));
    jand g0201(.dinb(n13405), .dina(n1057), .dout(n1061));
    jand g0202(.dinb(n13315), .dina(n1061), .dout(n1065));
    jor g0203(.dinb(n13300), .dina(n1065), .dout(n1069));
    jand g0204(.dinb(n987), .dina(n13281), .dout(n1073));
    jnot g0205(.din(G4427), .dout(n1076));
    jand g0206(.dinb(G18), .dina(G221), .dout(n1080));
    jand g0207(.dinb(n455), .dina(n13198), .dout(n1084));
    jor g0208(.dinb(n13195), .dina(n1084), .dout(n1088));
    jxor g0209(.dinb(n13206), .dina(n1088), .dout(n1092));
    jnot g0210(.din(G4420), .dout(n1095));
    jand g0211(.dinb(G18), .dina(G222), .dout(n1099));
    jand g0212(.dinb(n455), .dina(n13153), .dout(n1103));
    jor g0213(.dinb(n13150), .dina(n1103), .dout(n1107));
    jxor g0214(.dinb(n13161), .dina(n1107), .dout(n1111));
    jand g0215(.dinb(n1092), .dina(n1111), .dout(n1115));
    jnot g0216(.din(G4437), .dout(n1118));
    jand g0217(.dinb(G18), .dina(G219), .dout(n1122));
    jand g0218(.dinb(n455), .dina(n13255), .dout(n1126));
    jor g0219(.dinb(n13252), .dina(n1126), .dout(n1130));
    jxor g0220(.dinb(n13263), .dina(n1130), .dout(n1134));
    jnot g0221(.din(G4432), .dout(n1137));
    jand g0222(.dinb(G18), .dina(G220), .dout(n1141));
    jand g0223(.dinb(n455), .dina(n13780), .dout(n1145));
    jor g0224(.dinb(n13777), .dina(n1145), .dout(n1149));
    jxor g0225(.dinb(n13786), .dina(n1149), .dout(n1153));
    jand g0226(.dinb(n1134), .dina(n1153), .dout(n1157));
    jand g0227(.dinb(n1115), .dina(n1157), .dout(n1161));
    jnot g0228(.din(n1161), .dout(n1164));
    jor g0229(.dinb(n1073), .dina(n12406), .dout(n1168));
    jnot g0230(.din(n1130), .dout(n1171));
    jand g0231(.dinb(n13269), .dina(n1171), .dout(n1175));
    jnot g0232(.din(n1175), .dout(n1178));
    jand g0233(.dinb(n13257), .dina(n1130), .dout(n1182));
    jand g0234(.dinb(n13786), .dina(n1149), .dout(n1186));
    jnot g0235(.din(n1149), .dout(n1189));
    jand g0236(.dinb(n13788), .dina(n1189), .dout(n1193));
    jnot g0237(.din(n1193), .dout(n1196));
    jand g0238(.dinb(n13200), .dina(n1088), .dout(n1200));
    jand g0239(.dinb(n13155), .dina(n1107), .dout(n1204));
    jand g0240(.dinb(n1092), .dina(n1204), .dout(n1208));
    jor g0241(.dinb(n13192), .dina(n1208), .dout(n1212));
    jand g0242(.dinb(n1196), .dina(n1212), .dout(n1216));
    jor g0243(.dinb(n13080), .dina(n1216), .dout(n1220));
    jor g0244(.dinb(n12385), .dina(n1220), .dout(n1224));
    jand g0245(.dinb(n12373), .dina(n1224), .dout(n1228));
    jnot g0246(.din(n1228), .dout(n1231));
    jand g0247(.dinb(n1168), .dina(n12349), .dout(n1235));
    jnot g0248(.din(G2236), .dout(n1238));
    jand g0249(.dinb(G9), .dina(G12), .dout(n1242));
    jnot g0250(.din(n1242), .dout(n1245));
    jor g0251(.dinb(n455), .dina(n12307), .dout(n1249));
    jand g0252(.dinb(n1245), .dina(n1249), .dout(n1253));
    jxor g0253(.dinb(n12325), .dina(n1253), .dout(n1257));
    jnot g0254(.din(G2218), .dout(n1260));
    jand g0255(.dinb(n455), .dina(n12280), .dout(n1264));
    jand g0256(.dinb(G18), .dina(G160), .dout(n1268));
    jor g0257(.dinb(n1264), .dina(n12277), .dout(n1272));
    jxor g0258(.dinb(n12286), .dina(n1272), .dout(n1276));
    jnot g0259(.din(G2211), .dout(n1279));
    jand g0260(.dinb(n455), .dina(n12223), .dout(n1283));
    jand g0261(.dinb(G18), .dina(G151), .dout(n1287));
    jor g0262(.dinb(n1283), .dina(n12220), .dout(n1291));
    jxor g0263(.dinb(n12229), .dina(n1291), .dout(n1295));
    jand g0264(.dinb(n1276), .dina(n1295), .dout(n1299));
    jnot g0265(.din(G2230), .dout(n1302));
    jand g0266(.dinb(n455), .dina(n12115), .dout(n1306));
    jand g0267(.dinb(G18), .dina(G158), .dout(n1310));
    jor g0268(.dinb(n1306), .dina(n12112), .dout(n1314));
    jxor g0269(.dinb(n12121), .dina(n1314), .dout(n1318));
    jnot g0270(.din(G2224), .dout(n1321));
    jand g0271(.dinb(n455), .dina(n12091), .dout(n1325));
    jand g0272(.dinb(G18), .dina(G159), .dout(n1329));
    jor g0273(.dinb(n1325), .dina(n12088), .dout(n1333));
    jxor g0274(.dinb(n12097), .dina(n1333), .dout(n1337));
    jand g0275(.dinb(n1318), .dina(n1337), .dout(n1341));
    jand g0276(.dinb(n1299), .dina(n1341), .dout(n1345));
    jand g0277(.dinb(n12300), .dina(n1345), .dout(n1349));
    jnot g0278(.din(n1349), .dout(n1352));
    jor g0279(.dinb(n1235), .dina(n12055), .dout(n1356));
    jand g0280(.dinb(n12325), .dina(n1253), .dout(n1360));
    jnot g0281(.din(n1360), .dout(n1363));
    jnot g0282(.din(n1253), .dout(n1366));
    jand g0283(.dinb(n12327), .dina(n1366), .dout(n1370));
    jand g0284(.dinb(n12121), .dina(n1314), .dout(n1374));
    jnot g0285(.din(n1374), .dout(n1377));
    jnot g0286(.din(n1314), .dout(n1380));
    jand g0287(.dinb(n12123), .dina(n1380), .dout(n1384));
    jnot g0288(.din(n1333), .dout(n1387));
    jand g0289(.dinb(n12099), .dina(n1387), .dout(n1391));
    jnot g0290(.din(n1391), .dout(n1394));
    jand g0291(.dinb(n12229), .dina(n1291), .dout(n1398));
    jand g0292(.dinb(n1276), .dina(n1398), .dout(n1402));
    jand g0293(.dinb(n12286), .dina(n1272), .dout(n1406));
    jand g0294(.dinb(n12097), .dina(n1333), .dout(n1410));
    jor g0295(.dinb(n1406), .dina(n1410), .dout(n1414));
    jor g0296(.dinb(n1402), .dina(n1414), .dout(n1418));
    jand g0297(.dinb(n1394), .dina(n1418), .dout(n1422));
    jnot g0298(.din(n1422), .dout(n1425));
    jor g0299(.dinb(n11923), .dina(n1425), .dout(n1429));
    jand g0300(.dinb(n11914), .dina(n1429), .dout(n1433));
    jor g0301(.dinb(n11875), .dina(n1433), .dout(n1437));
    jand g0302(.dinb(n11860), .dina(n1437), .dout(n1441));
    jand g0303(.dinb(n1356), .dina(n11829), .dout(n1445));
    jnot g0304(.din(G2247), .dout(n1448));
    jor g0305(.dinb(n455), .dina(n11821), .dout(n1452));
    jand g0306(.dinb(n1245), .dina(n1452), .dout(n1456));
    jxor g0307(.dinb(n11827), .dina(n1456), .dout(n1460));
    jnot g0308(.din(G2239), .dout(n1463));
    jor g0309(.dinb(n455), .dina(n11740), .dout(n1467));
    jand g0310(.dinb(n1245), .dina(n1467), .dout(n1471));
    jxor g0311(.dinb(n11748), .dina(n1471), .dout(n1475));
    jand g0312(.dinb(n1460), .dina(n1475), .dout(n1479));
    jnot g0313(.din(G2256), .dout(n1482));
    jor g0314(.dinb(n455), .dina(n11671), .dout(n1486));
    jand g0315(.dinb(n1245), .dina(n1486), .dout(n1490));
    jxor g0316(.dinb(n11677), .dina(n1490), .dout(n1494));
    jnot g0317(.din(G2253), .dout(n1497));
    jor g0318(.dinb(n455), .dina(n11644), .dout(n1501));
    jand g0319(.dinb(n1245), .dina(n1501), .dout(n1505));
    jxor g0320(.dinb(n11650), .dina(n1505), .dout(n1509));
    jand g0321(.dinb(n1494), .dina(n1509), .dout(n1513));
    jand g0322(.dinb(n1479), .dina(n1513), .dout(n1517));
    jnot g0323(.din(n1517), .dout(n1520));
    jor g0324(.dinb(n1445), .dina(n11596), .dout(n1524));
    jand g0325(.dinb(n11677), .dina(n1490), .dout(n1528));
    jnot g0326(.din(n1528), .dout(n1531));
    jand g0327(.dinb(n11650), .dina(n1505), .dout(n1535));
    jnot g0328(.din(n1535), .dout(n1538));
    jand g0329(.dinb(n11827), .dina(n1456), .dout(n1542));
    jand g0330(.dinb(n11742), .dina(n1471), .dout(n1546));
    jand g0331(.dinb(n1460), .dina(n1546), .dout(n1550));
    jor g0332(.dinb(n11452), .dina(n1550), .dout(n1554));
    jnot g0333(.din(n1554), .dout(n1557));
    jand g0334(.dinb(n11548), .dina(n1557), .dout(n1561));
    jnot g0335(.din(n1490), .dout(n1564));
    jand g0336(.dinb(n11679), .dina(n1564), .dout(n1568));
    jnot g0337(.din(n1505), .dout(n1571));
    jand g0338(.dinb(n11652), .dina(n1571), .dout(n1575));
    jor g0339(.dinb(n1568), .dina(n1575), .dout(n1579));
    jor g0340(.dinb(n1561), .dina(n11359), .dout(n1583));
    jand g0341(.dinb(n11353), .dina(n1583), .dout(n1587));
    jand g0342(.dinb(n1524), .dina(n11316), .dout(n1591));
    jnot g0343(.din(G1486), .dout(n1594));
    jor g0344(.dinb(n455), .dina(n11308), .dout(n1598));
    jand g0345(.dinb(n1245), .dina(n1598), .dout(n1602));
    jxor g0346(.dinb(n11314), .dina(n1602), .dout(n1606));
    jnot g0347(.din(G1480), .dout(n1609));
    jor g0348(.dinb(n455), .dina(n11293), .dout(n1613));
    jand g0349(.dinb(n1245), .dina(n1613), .dout(n1617));
    jxor g0350(.dinb(n11299), .dina(n1617), .dout(n1621));
    jnot g0351(.din(G106), .dout(n1624));
    jor g0352(.dinb(n455), .dina(n11272), .dout(n1628));
    jand g0353(.dinb(n1245), .dina(n1628), .dout(n1632));
    jxor g0354(.dinb(n11278), .dina(n1632), .dout(n1636));
    jand g0355(.dinb(n1621), .dina(n1636), .dout(n1640));
    jnot g0356(.din(G1469), .dout(n1643));
    jor g0357(.dinb(n455), .dina(n11245), .dout(n1647));
    jand g0358(.dinb(n1245), .dina(n1647), .dout(n1651));
    jxor g0359(.dinb(n11251), .dina(n1651), .dout(n1655));
    jnot g0360(.din(G1462), .dout(n1658));
    jor g0361(.dinb(n455), .dina(n11137), .dout(n1662));
    jand g0362(.dinb(n1245), .dina(n1662), .dout(n1666));
    jxor g0363(.dinb(n11143), .dina(n1666), .dout(n1670));
    jand g0364(.dinb(n1655), .dina(n1670), .dout(n1674));
    jand g0365(.dinb(n1640), .dina(n1674), .dout(n1678));
    jand g0366(.dinb(n11301), .dina(n1678), .dout(n1682));
    jnot g0367(.din(n1682), .dout(n1685));
    jor g0368(.dinb(n1591), .dina(n11014), .dout(n1689));
    jand g0369(.dinb(n11314), .dina(n1602), .dout(n1693));
    jor g0370(.dinb(n11314), .dina(n1602), .dout(n1697));
    jand g0371(.dinb(n11299), .dina(n1617), .dout(n1701));
    jnot g0372(.din(n1701), .dout(n1704));
    jor g0373(.dinb(n11299), .dina(n1617), .dout(n1708));
    jand g0374(.dinb(n11278), .dina(n1632), .dout(n1712));
    jnot g0375(.din(n1632), .dout(n1715));
    jand g0376(.dinb(n11280), .dina(n1715), .dout(n1719));
    jnot g0377(.din(n1719), .dout(n1722));
    jnot g0378(.din(n1651), .dout(n1725));
    jand g0379(.dinb(n11253), .dina(n1725), .dout(n1729));
    jnot g0380(.din(n1729), .dout(n1732));
    jand g0381(.dinb(n11251), .dina(n1651), .dout(n1736));
    jand g0382(.dinb(n11143), .dina(n1666), .dout(n1740));
    jor g0383(.dinb(n1736), .dina(n1740), .dout(n1744));
    jand g0384(.dinb(n1732), .dina(n10855), .dout(n1748));
    jand g0385(.dinb(n10944), .dina(n1748), .dout(n1752));
    jor g0386(.dinb(n10852), .dina(n1752), .dout(n1756));
    jand g0387(.dinb(n10840), .dina(n1756), .dout(n1760));
    jnot g0388(.din(n1760), .dout(n1763));
    jand g0389(.dinb(n10947), .dina(n1763), .dout(n1767));
    jnot g0390(.din(n1767), .dout(n1770));
    jand g0391(.dinb(n10792), .dina(n1770), .dout(n1774));
    jor g0392(.dinb(n10765), .dina(n1774), .dout(n1778));
    jnot g0393(.din(n1778), .dout(n1781));
    jand g0394(.dinb(n1689), .dina(n10707), .dout(n1785));
    jnot g0395(.din(G38), .dout(n1788));
    jand g0396(.dinb(G1492), .dina(G4528), .dout(n1792));
    jxor g0397(.dinb(n1788), .dina(n1792), .dout(n1796));
    jnot g0398(.din(n1796), .dout(n1799));
    jor g0399(.dinb(n1785), .dina(n10663), .dout(n1803));
    jor g0400(.dinb(n12621), .dina(n1803), .dout(n1807));
    jnot g0401(.din(n1807), .dout(n1810));
    jnot g0402(.din(G1492), .dout(n1813));
    jnot g0403(.din(n490), .dout(n1816));
    jor g0404(.dinb(n9718), .dina(n1816), .dout(n1820));
    jand g0405(.dinb(n12684), .dina(n1820), .dout(n1824));
    jor g0406(.dinb(n1810), .dina(n9715), .dout(n1828));
    jor g0407(.dinb(n455), .dina(n9223), .dout(n1832));
    jand g0408(.dinb(n1245), .dina(n1832), .dout(n1836));
    jand g0409(.dinb(G18), .dina(G2236), .dout(n1840));
    jnot g0410(.din(n1840), .dout(n1843));
    jor g0411(.dinb(G18), .dina(G64), .dout(n1847));
    jand g0412(.dinb(n1843), .dina(n9475), .dout(n1851));
    jor g0413(.dinb(n1836), .dina(n1851), .dout(n1855));
    jand g0414(.dinb(G18), .dina(G178), .dout(n1859));
    jor g0415(.dinb(n1306), .dina(n9229), .dout(n1863));
    jand g0416(.dinb(G18), .dina(G2230), .dout(n1867));
    jnot g0417(.din(n1867), .dout(n1870));
    jor g0418(.dinb(G18), .dina(G85), .dout(n1874));
    jand g0419(.dinb(n1870), .dina(n9442), .dout(n1878));
    jor g0420(.dinb(n1863), .dina(n1878), .dout(n1882));
    jand g0421(.dinb(G18), .dina(G179), .dout(n1886));
    jor g0422(.dinb(n1325), .dina(n9235), .dout(n1890));
    jand g0423(.dinb(G18), .dina(G2224), .dout(n1894));
    jnot g0424(.din(n1894), .dout(n1897));
    jor g0425(.dinb(G18), .dina(G84), .dout(n1901));
    jand g0426(.dinb(n1897), .dina(n9439), .dout(n1905));
    jand g0427(.dinb(n1890), .dina(n1905), .dout(n1909));
    jand g0428(.dinb(G18), .dina(G180), .dout(n1913));
    jor g0429(.dinb(n1264), .dina(n9226), .dout(n1917));
    jand g0430(.dinb(G18), .dina(G2218), .dout(n1921));
    jnot g0431(.din(n1921), .dout(n1924));
    jor g0432(.dinb(G18), .dina(G83), .dout(n1928));
    jand g0433(.dinb(n1924), .dina(n9451), .dout(n1932));
    jor g0434(.dinb(n1917), .dina(n1932), .dout(n1936));
    jor g0435(.dinb(n1890), .dina(n1905), .dout(n1940));
    jand g0436(.dinb(n1936), .dina(n1940), .dout(n1944));
    jand g0437(.dinb(n1917), .dina(n1932), .dout(n1948));
    jand g0438(.dinb(G18), .dina(G171), .dout(n1952));
    jor g0439(.dinb(n1283), .dina(n9220), .dout(n1956));
    jand g0440(.dinb(G18), .dina(G2211), .dout(n1960));
    jnot g0441(.din(n1960), .dout(n1963));
    jor g0442(.dinb(G18), .dina(G65), .dout(n1967));
    jand g0443(.dinb(n1963), .dina(n9448), .dout(n1971));
    jand g0444(.dinb(n1956), .dina(n1971), .dout(n1975));
    jor g0445(.dinb(n1948), .dina(n1975), .dout(n1979));
    jand g0446(.dinb(n1944), .dina(n1979), .dout(n1983));
    jor g0447(.dinb(n8493), .dina(n1983), .dout(n1987));
    jand g0448(.dinb(n8499), .dina(n1987), .dout(n1991));
    jand g0449(.dinb(n1863), .dina(n1878), .dout(n1995));
    jand g0450(.dinb(n1836), .dina(n1851), .dout(n1999));
    jor g0451(.dinb(n1995), .dina(n1999), .dout(n2003));
    jor g0452(.dinb(n1991), .dina(n8485), .dout(n2007));
    jand g0453(.dinb(n8508), .dina(n2007), .dout(n2011));
    jnot g0454(.din(n1948), .dout(n2014));
    jand g0455(.dinb(n8506), .dina(n2014), .dout(n2018));
    jnot g0456(.din(n1909), .dout(n2021));
    jnot g0457(.din(n1975), .dout(n2024));
    jand g0458(.dinb(n2021), .dina(n2024), .dout(n2028));
    jand g0459(.dinb(n2018), .dina(n2028), .dout(n2032));
    jnot g0460(.din(n1999), .dout(n2035));
    jor g0461(.dinb(n1956), .dina(n1971), .dout(n2039));
    jand g0462(.dinb(n2035), .dina(n8476), .dout(n2043));
    jnot g0463(.din(n1995), .dout(n2046));
    jand g0464(.dinb(n8521), .dina(n2046), .dout(n2050));
    jand g0465(.dinb(n2043), .dina(n2050), .dout(n2054));
    jand g0466(.dinb(n8487), .dina(n2054), .dout(n2058));
    jand g0467(.dinb(n8473), .dina(n2058), .dout(n2062));
    jand g0468(.dinb(G18), .dina(G191), .dout(n2066));
    jor g0469(.dinb(n1084), .dina(n9352), .dout(n2070));
    jor g0470(.dinb(G18), .dina(G60), .dout(n2074));
    jor g0471(.dinb(n455), .dina(n1076), .dout(n2078));
    jand g0472(.dinb(n9634), .dina(n2078), .dout(n2082));
    jxor g0473(.dinb(n2070), .dina(n2082), .dout(n2086));
    jand g0474(.dinb(G18), .dina(G189), .dout(n2090));
    jor g0475(.dinb(n1126), .dina(n9349), .dout(n2094));
    jor g0476(.dinb(G18), .dina(G62), .dout(n2098));
    jor g0477(.dinb(n455), .dina(n1118), .dout(n2102));
    jand g0478(.dinb(n9631), .dina(n2102), .dout(n2106));
    jxor g0479(.dinb(n2094), .dina(n2106), .dout(n2110));
    jand g0480(.dinb(n2086), .dina(n2110), .dout(n2114));
    jand g0481(.dinb(G18), .dina(G190), .dout(n2118));
    jor g0482(.dinb(n1145), .dina(n9346), .dout(n2122));
    jor g0483(.dinb(G18), .dina(G61), .dout(n2126));
    jand g0484(.dinb(G18), .dina(G4432), .dout(n2130));
    jnot g0485(.din(n2130), .dout(n2133));
    jand g0486(.dinb(n9628), .dina(n2133), .dout(n2137));
    jxor g0487(.dinb(n2122), .dina(n2137), .dout(n2141));
    jand g0488(.dinb(G18), .dina(G192), .dout(n2145));
    jor g0489(.dinb(n1103), .dina(n9343), .dout(n2149));
    jor g0490(.dinb(G18), .dina(G79), .dout(n2153));
    jor g0491(.dinb(n455), .dina(n1095), .dout(n2157));
    jand g0492(.dinb(n9625), .dina(n2157), .dout(n2161));
    jxor g0493(.dinb(n2149), .dina(n2161), .dout(n2165));
    jand g0494(.dinb(n2141), .dina(n2165), .dout(n2169));
    jand g0495(.dinb(n2114), .dina(n2169), .dout(n2173));
    jand g0496(.dinb(G18), .dina(G196), .dout(n2177));
    jor g0497(.dinb(n899), .dina(n9325), .dout(n2181));
    jor g0498(.dinb(G18), .dina(G78), .dout(n2185));
    jand g0499(.dinb(G18), .dina(G4400), .dout(n2189));
    jnot g0500(.din(n2189), .dout(n2192));
    jand g0501(.dinb(n9640), .dina(n2192), .dout(n2196));
    jor g0502(.dinb(n2181), .dina(n2196), .dout(n2200));
    jand g0503(.dinb(G18), .dina(G195), .dout(n2204));
    jor g0504(.dinb(n957), .dina(n9331), .dout(n2208));
    jor g0505(.dinb(G18), .dina(G59), .dout(n2212));
    jand g0506(.dinb(G18), .dina(G4405), .dout(n2216));
    jnot g0507(.din(n2216), .dout(n2219));
    jand g0508(.dinb(n9652), .dina(n2219), .dout(n2223));
    jor g0509(.dinb(n2208), .dina(n2223), .dout(n2227));
    jand g0510(.dinb(n2200), .dina(n2227), .dout(n2231));
    jand g0511(.dinb(G18), .dina(G187), .dout(n2235));
    jor g0512(.dinb(n915), .dina(n9328), .dout(n2239));
    jor g0513(.dinb(G18), .dina(G77), .dout(n2243));
    jand g0514(.dinb(G18), .dina(G4394), .dout(n2247));
    jnot g0515(.din(n2247), .dout(n2250));
    jand g0516(.dinb(n9649), .dina(n2250), .dout(n2254));
    jand g0517(.dinb(n2239), .dina(n2254), .dout(n2258));
    jnot g0518(.din(n2258), .dout(n2261));
    jand g0519(.dinb(n2208), .dina(n2223), .dout(n2265));
    jnot g0520(.din(n2265), .dout(n2268));
    jand g0521(.dinb(n2261), .dina(n2268), .dout(n2272));
    jand g0522(.dinb(n8656), .dina(n2272), .dout(n2276));
    jand g0523(.dinb(n2181), .dina(n2196), .dout(n2280));
    jnot g0524(.din(n2280), .dout(n2283));
    jor g0525(.dinb(n2239), .dina(n2254), .dout(n2287));
    jand g0526(.dinb(n2283), .dina(n8653), .dout(n2291));
    jand g0527(.dinb(G18), .dina(G193), .dout(n2295));
    jor g0528(.dinb(n880), .dina(n9322), .dout(n2299));
    jor g0529(.dinb(G18), .dina(G80), .dout(n2303));
    jand g0530(.dinb(G18), .dina(G4415), .dout(n2307));
    jnot g0531(.din(n2307), .dout(n2310));
    jand g0532(.dinb(n9637), .dina(n2310), .dout(n2314));
    jand g0533(.dinb(n2299), .dina(n2314), .dout(n2318));
    jnot g0534(.din(n2318), .dout(n2321));
    jand g0535(.dinb(G18), .dina(G194), .dout(n2325));
    jor g0536(.dinb(n941), .dina(n9361), .dout(n2329));
    jor g0537(.dinb(G18), .dina(G81), .dout(n2333));
    jand g0538(.dinb(G18), .dina(G4410), .dout(n2337));
    jnot g0539(.din(n2337), .dout(n2340));
    jand g0540(.dinb(n9646), .dina(n2340), .dout(n2344));
    jor g0541(.dinb(n2329), .dina(n2344), .dout(n2348));
    jand g0542(.dinb(n2321), .dina(n8685), .dout(n2352));
    jor g0543(.dinb(n2299), .dina(n2314), .dout(n2356));
    jand g0544(.dinb(n2329), .dina(n2344), .dout(n2360));
    jnot g0545(.din(n2360), .dout(n2363));
    jand g0546(.dinb(n8682), .dina(n2363), .dout(n2367));
    jand g0547(.dinb(n2352), .dina(n2367), .dout(n2371));
    jand g0548(.dinb(n8650), .dina(n2371), .dout(n2375));
    jand g0549(.dinb(n8647), .dina(n2375), .dout(n2379));
    jand g0550(.dinb(n8712), .dina(n2379), .dout(n2383));
    jand g0551(.dinb(G18), .dina(G200), .dout(n2387));
    jnot g0552(.din(n2387), .dout(n2390));
    jand g0553(.dinb(n775), .dina(n2390), .dout(n2394));
    jnot g0554(.din(n2394), .dout(n2397));
    jor g0555(.dinb(G18), .dina(G56), .dout(n2401));
    jand g0556(.dinb(G18), .dina(G3749), .dout(n2405));
    jnot g0557(.din(n2405), .dout(n2408));
    jand g0558(.dinb(n9556), .dina(n2408), .dout(n2412));
    jand g0559(.dinb(n2397), .dina(n9552), .dout(n2416));
    jnot g0560(.din(n2416), .dout(n2419));
    jnot g0561(.din(n724), .dout(n2422));
    jand g0562(.dinb(G18), .dina(G202), .dout(n2426));
    jor g0563(.dinb(n2422), .dina(n9307), .dout(n2430));
    jor g0564(.dinb(G18), .dina(G54), .dout(n2434));
    jand g0565(.dinb(G18), .dina(G3737), .dout(n2438));
    jnot g0566(.din(n2438), .dout(n2441));
    jand g0567(.dinb(n9547), .dina(n2441), .dout(n2445));
    jor g0568(.dinb(n2430), .dina(n9543), .dout(n2449));
    jand g0569(.dinb(n2419), .dina(n8626), .dout(n2453));
    jand g0570(.dinb(n2430), .dina(n9540), .dout(n2457));
    jnot g0571(.din(n2457), .dout(n2460));
    jor g0572(.dinb(n2397), .dina(n9549), .dout(n2464));
    jand g0573(.dinb(n2460), .dina(n8622), .dout(n2468));
    jand g0574(.dinb(n2453), .dina(n2468), .dout(n2472));
    jand g0575(.dinb(G18), .dina(G201), .dout(n2476));
    jor g0576(.dinb(n802), .dina(n9301), .dout(n2480));
    jor g0577(.dinb(G18), .dina(G55), .dout(n2484));
    jand g0578(.dinb(G18), .dina(G3743), .dout(n2488));
    jnot g0579(.din(n2488), .dout(n2491));
    jand g0580(.dinb(n9538), .dina(n2491), .dout(n2495));
    jxor g0581(.dinb(n2480), .dina(n2495), .dout(n2499));
    jnot g0582(.din(n749), .dout(n2502));
    jand g0583(.dinb(G18), .dina(G203), .dout(n2506));
    jor g0584(.dinb(n2502), .dina(n9295), .dout(n2510));
    jor g0585(.dinb(G18), .dina(G53), .dout(n2514));
    jor g0586(.dinb(n455), .dina(n735), .dout(n2518));
    jand g0587(.dinb(n9535), .dina(n2518), .dout(n2522));
    jxor g0588(.dinb(n2510), .dina(n9531), .dout(n2526));
    jand g0589(.dinb(n8620), .dina(n2526), .dout(n2530));
    jand g0590(.dinb(n2472), .dina(n8596), .dout(n2534));
    jnot g0591(.din(n619), .dout(n2537));
    jand g0592(.dinb(G18), .dina(G207), .dout(n2541));
    jor g0593(.dinb(n2537), .dina(n9262), .dout(n2545));
    jor g0594(.dinb(G18), .dina(G74), .dout(n2549));
    jand g0595(.dinb(G18), .dina(G3705), .dout(n2553));
    jnot g0596(.din(n2553), .dout(n2556));
    jand g0597(.dinb(n9598), .dina(n2556), .dout(n2560));
    jor g0598(.dinb(n2545), .dina(n9595), .dout(n2564));
    jnot g0599(.din(n533), .dout(n2567));
    jand g0600(.dinb(G18), .dina(G205), .dout(n2571));
    jor g0601(.dinb(n2567), .dina(n9280), .dout(n2575));
    jor g0602(.dinb(G18), .dina(G75), .dout(n2579));
    jand g0603(.dinb(G18), .dina(G3717), .dout(n2583));
    jnot g0604(.din(n2583), .dout(n2586));
    jand g0605(.dinb(n9565), .dina(n2586), .dout(n2590));
    jor g0606(.dinb(n2575), .dina(n9561), .dout(n2594));
    jand g0607(.dinb(n2564), .dina(n2594), .dout(n2598));
    jand g0608(.dinb(n2575), .dina(n9558), .dout(n2602));
    jnot g0609(.din(n2602), .dout(n2605));
    jnot g0610(.din(n565), .dout(n2608));
    jand g0611(.dinb(G18), .dina(G206), .dout(n2612));
    jor g0612(.dinb(n2608), .dina(n9274), .dout(n2616));
    jor g0613(.dinb(G18), .dina(G76), .dout(n2620));
    jand g0614(.dinb(G18), .dina(G3711), .dout(n2624));
    jnot g0615(.din(n2624), .dout(n2627));
    jand g0616(.dinb(n9583), .dina(n2627), .dout(n2631));
    jor g0617(.dinb(n2616), .dina(n9579), .dout(n2635));
    jand g0618(.dinb(n2605), .dina(n8583), .dout(n2639));
    jand g0619(.dinb(n8581), .dina(n2639), .dout(n2643));
    jnot g0620(.din(G70), .dout(n2646));
    jand g0621(.dinb(n455), .dina(n2646), .dout(n2650));
    jnot g0622(.din(n2650), .dout(n2653));
    jor g0623(.dinb(n14340), .dina(n2653), .dout(n2657));
    jand g0624(.dinb(n14337), .dina(n2653), .dout(n2661));
    jnot g0625(.din(n2661), .dout(n2664));
    jand g0626(.dinb(n8575), .dina(n2664), .dout(n2668));
    jand g0627(.dinb(n8560), .dina(n2668), .dout(n2672));
    jnot g0628(.din(n511), .dout(n2675));
    jand g0629(.dinb(G18), .dina(G204), .dout(n2679));
    jor g0630(.dinb(n2675), .dina(n9268), .dout(n2683));
    jor g0631(.dinb(G18), .dina(G73), .dout(n2687));
    jor g0632(.dinb(n455), .dina(n497), .dout(n2691));
    jand g0633(.dinb(n9574), .dina(n2691), .dout(n2695));
    jxor g0634(.dinb(n2683), .dina(n9567), .dout(n2699));
    jand g0635(.dinb(n2545), .dina(n9595), .dout(n2703));
    jnot g0636(.din(n2703), .dout(n2706));
    jand g0637(.dinb(n2616), .dina(n9576), .dout(n2710));
    jnot g0638(.din(n2710), .dout(n2713));
    jand g0639(.dinb(n2706), .dina(n2713), .dout(n2717));
    jand g0640(.dinb(n8554), .dina(n2717), .dout(n2721));
    jand g0641(.dinb(n8548), .dina(n2721), .dout(n2725));
    jand g0642(.dinb(n8545), .dina(n2725), .dout(n2729));
    jand g0643(.dinb(n8590), .dina(n2729), .dout(n2733));
    jand g0644(.dinb(n8457), .dina(n2733), .dout(n2737));
    jand g0645(.dinb(n2149), .dina(n2161), .dout(n2741));
    jand g0646(.dinb(n2141), .dina(n2741), .dout(n2745));
    jand g0647(.dinb(n2114), .dina(n2745), .dout(n2749));
    jand g0648(.dinb(n2094), .dina(n2106), .dout(n2753));
    jand g0649(.dinb(n2070), .dina(n2082), .dout(n2757));
    jand g0650(.dinb(n2122), .dina(n2137), .dout(n2761));
    jor g0651(.dinb(n2757), .dina(n2761), .dout(n2765));
    jor g0652(.dinb(n2094), .dina(n2106), .dout(n2769));
    jor g0653(.dinb(n2122), .dina(n2137), .dout(n2773));
    jand g0654(.dinb(n2769), .dina(n2773), .dout(n2777));
    jand g0655(.dinb(n2765), .dina(n2777), .dout(n2781));
    jor g0656(.dinb(n8752), .dina(n2781), .dout(n2785));
    jor g0657(.dinb(n8746), .dina(n2785), .dout(n2789));
    jand g0658(.dinb(n2200), .dina(n2258), .dout(n2793));
    jor g0659(.dinb(n2265), .dina(n2280), .dout(n2797));
    jor g0660(.dinb(n2793), .dina(n2797), .dout(n2801));
    jand g0661(.dinb(n2348), .dina(n2356), .dout(n2805));
    jand g0662(.dinb(n8688), .dina(n2805), .dout(n2809));
    jand g0663(.dinb(n2801), .dina(n2809), .dout(n2813));
    jand g0664(.dinb(n2356), .dina(n2360), .dout(n2817));
    jor g0665(.dinb(n8679), .dina(n2817), .dout(n2821));
    jor g0666(.dinb(n2813), .dina(n8677), .dout(n2825));
    jand g0667(.dinb(n8719), .dina(n2825), .dout(n2829));
    jor g0668(.dinb(n8743), .dina(n2829), .dout(n2833));
    jor g0669(.dinb(n2737), .dina(n8455), .dout(n2837));
    jand g0670(.dinb(n8460), .dina(n2837), .dout(n2841));
    jor g0671(.dinb(n8449), .dina(n2841), .dout(n2845));
    jor g0672(.dinb(n455), .dina(n9211), .dout(n2849));
    jand g0673(.dinb(n1245), .dina(n2849), .dout(n2853));
    jand g0674(.dinb(G18), .dina(G2256), .dout(n2857));
    jnot g0675(.din(n2857), .dout(n2860));
    jor g0676(.dinb(G18), .dina(G110), .dout(n2864));
    jand g0677(.dinb(n2860), .dina(n9466), .dout(n2868));
    jor g0678(.dinb(n2853), .dina(n2868), .dout(n2872));
    jor g0679(.dinb(n455), .dina(n9217), .dout(n2876));
    jand g0680(.dinb(n1245), .dina(n2876), .dout(n2880));
    jand g0681(.dinb(G18), .dina(G2247), .dout(n2884));
    jnot g0682(.din(n2884), .dout(n2887));
    jor g0683(.dinb(G18), .dina(G86), .dout(n2891));
    jand g0684(.dinb(n2887), .dina(n9463), .dout(n2895));
    jand g0685(.dinb(n2880), .dina(n2895), .dout(n2899));
    jnot g0686(.din(n2899), .dout(n2902));
    jand g0687(.dinb(n8436), .dina(n2902), .dout(n2906));
    jand g0688(.dinb(n2853), .dina(n2868), .dout(n2910));
    jnot g0689(.din(n2910), .dout(n2913));
    jor g0690(.dinb(n2880), .dina(n2895), .dout(n2917));
    jand g0691(.dinb(n2913), .dina(n8428), .dout(n2921));
    jand g0692(.dinb(n2906), .dina(n2921), .dout(n2925));
    jor g0693(.dinb(n455), .dina(n9208), .dout(n2929));
    jand g0694(.dinb(n1245), .dina(n2929), .dout(n2933));
    jand g0695(.dinb(G18), .dina(G2253), .dout(n2937));
    jnot g0696(.din(n2937), .dout(n2940));
    jor g0697(.dinb(G18), .dina(G109), .dout(n2944));
    jand g0698(.dinb(n2940), .dina(n9460), .dout(n2948));
    jxor g0699(.dinb(n2933), .dina(n2948), .dout(n2952));
    jor g0700(.dinb(n455), .dina(n9214), .dout(n2956));
    jand g0701(.dinb(n1245), .dina(n2956), .dout(n2960));
    jor g0702(.dinb(n455), .dina(n1463), .dout(n2964));
    jor g0703(.dinb(G18), .dina(G63), .dout(n2968));
    jand g0704(.dinb(n2964), .dina(n9457), .dout(n2972));
    jxor g0705(.dinb(n2960), .dina(n2972), .dout(n2976));
    jand g0706(.dinb(n2952), .dina(n2976), .dout(n2980));
    jand g0707(.dinb(n2925), .dina(n8425), .dout(n2984));
    jand g0708(.dinb(n2845), .dina(n8400), .dout(n2988));
    jand g0709(.dinb(n2683), .dina(n9567), .dout(n2992));
    jor g0710(.dinb(n8577), .dina(n2703), .dout(n2996));
    jand g0711(.dinb(n2564), .dina(n2635), .dout(n3000));
    jand g0712(.dinb(n2996), .dina(n3000), .dout(n3004));
    jor g0713(.dinb(n2602), .dina(n2710), .dout(n3008));
    jor g0714(.dinb(n3004), .dina(n8542), .dout(n3012));
    jor g0715(.dinb(n2683), .dina(n9570), .dout(n3016));
    jand g0716(.dinb(n2594), .dina(n3016), .dout(n3020));
    jand g0717(.dinb(n3012), .dina(n8539), .dout(n3024));
    jor g0718(.dinb(n8533), .dina(n3024), .dout(n3028));
    jand g0719(.dinb(n8590), .dina(n3028), .dout(n3032));
    jand g0720(.dinb(n2510), .dina(n9528), .dout(n3036));
    jand g0721(.dinb(n8620), .dina(n3036), .dout(n3040));
    jand g0722(.dinb(n2472), .dina(n8617), .dout(n3044));
    jand g0723(.dinb(n2480), .dina(n2495), .dout(n3048));
    jor g0724(.dinb(n2457), .dina(n8611), .dout(n3052));
    jor g0725(.dinb(n2480), .dina(n2495), .dout(n3056));
    jand g0726(.dinb(n2464), .dina(n8608), .dout(n3060));
    jand g0727(.dinb(n3052), .dina(n3060), .dout(n3064));
    jor g0728(.dinb(n8628), .dina(n3064), .dout(n3068));
    jor g0729(.dinb(n3044), .dina(n8605), .dout(n3072));
    jor g0730(.dinb(n3032), .dina(n8602), .dout(n3076));
    jand g0731(.dinb(n2062), .dina(n8419), .dout(n3080));
    jand g0732(.dinb(n2383), .dina(n3080), .dout(n3084));
    jand g0733(.dinb(n3076), .dina(n8398), .dout(n3088));
    jand g0734(.dinb(n2960), .dina(n2972), .dout(n3092));
    jand g0735(.dinb(n2952), .dina(n3092), .dout(n3096));
    jand g0736(.dinb(n2925), .dina(n8395), .dout(n3100));
    jand g0737(.dinb(n2933), .dina(n2948), .dout(n3104));
    jor g0738(.dinb(n2899), .dina(n3104), .dout(n3108));
    jor g0739(.dinb(n2933), .dina(n2948), .dout(n3112));
    jand g0740(.dinb(n2872), .dina(n3112), .dout(n3116));
    jand g0741(.dinb(n3108), .dina(n3116), .dout(n3120));
    jor g0742(.dinb(n8430), .dina(n3120), .dout(n3124));
    jor g0743(.dinb(n3100), .dina(n8389), .dout(n3128));
    jor g0744(.dinb(n3088), .dina(n8386), .dout(n3132));
    jor g0745(.dinb(n2988), .dina(n8374), .dout(n3136));
    jor g0746(.dinb(n455), .dina(n9418), .dout(n3140));
    jand g0747(.dinb(n1245), .dina(n3140), .dout(n3144));
    jand g0748(.dinb(G18), .dina(G1480), .dout(n3148));
    jnot g0749(.din(n3148), .dout(n3151));
    jor g0750(.dinb(G18), .dina(G112), .dout(n3155));
    jand g0751(.dinb(n3151), .dina(n9499), .dout(n3159));
    jor g0752(.dinb(n3144), .dina(n3159), .dout(n3163));
    jor g0753(.dinb(n455), .dina(n9412), .dout(n3167));
    jand g0754(.dinb(n1245), .dina(n3167), .dout(n3171));
    jand g0755(.dinb(G18), .dina(G1486), .dout(n3175));
    jnot g0756(.din(n3175), .dout(n3178));
    jor g0757(.dinb(G18), .dina(G88), .dout(n3182));
    jand g0758(.dinb(n3178), .dina(n9493), .dout(n3186));
    jor g0759(.dinb(n3171), .dina(n3186), .dout(n3190));
    jand g0760(.dinb(n3163), .dina(n3190), .dout(n3194));
    jor g0761(.dinb(n455), .dina(n9400), .dout(n3198));
    jand g0762(.dinb(n1245), .dina(n3198), .dout(n3202));
    jand g0763(.dinb(G18), .dina(G1469), .dout(n3206));
    jnot g0764(.din(n3206), .dout(n3209));
    jor g0765(.dinb(G18), .dina(G111), .dout(n3213));
    jand g0766(.dinb(n3209), .dina(n9508), .dout(n3217));
    jor g0767(.dinb(n3202), .dina(n3217), .dout(n3221));
    jand g0768(.dinb(G18), .dina(G1462), .dout(n3225));
    jnot g0769(.din(n3225), .dout(n3228));
    jor g0770(.dinb(G18), .dina(G113), .dout(n3232));
    jand g0771(.dinb(n3228), .dina(n9505), .dout(n3236));
    jor g0772(.dinb(n9405), .dina(n3236), .dout(n3240));
    jand g0773(.dinb(n3221), .dina(n3240), .dout(n3244));
    jand g0774(.dinb(n3194), .dina(n3244), .dout(n3248));
    jand g0775(.dinb(n3202), .dina(n3217), .dout(n3252));
    jand g0776(.dinb(n9402), .dina(n3236), .dout(n3256));
    jor g0777(.dinb(n3252), .dina(n3256), .dout(n3260));
    jnot g0778(.din(n3260), .dout(n3263));
    jand g0779(.dinb(n3144), .dina(n3159), .dout(n3267));
    jor g0780(.dinb(n455), .dina(n9391), .dout(n3271));
    jand g0781(.dinb(n1245), .dina(n3271), .dout(n3275));
    jand g0782(.dinb(G18), .dina(G106), .dout(n3279));
    jnot g0783(.din(n3279), .dout(n3282));
    jor g0784(.dinb(G18), .dina(G87), .dout(n3286));
    jand g0785(.dinb(n3282), .dina(n9487), .dout(n3290));
    jand g0786(.dinb(n3275), .dina(n3290), .dout(n3294));
    jor g0787(.dinb(n3267), .dina(n3294), .dout(n3298));
    jnot g0788(.din(n3298), .dout(n3301));
    jor g0789(.dinb(n3275), .dina(n3290), .dout(n3305));
    jand g0790(.dinb(n3171), .dina(n3186), .dout(n3309));
    jnot g0791(.din(n3309), .dout(n3312));
    jand g0792(.dinb(n8358), .dina(n3312), .dout(n3316));
    jand g0793(.dinb(n3301), .dina(n3316), .dout(n3320));
    jand g0794(.dinb(n8356), .dina(n3320), .dout(n3324));
    jand g0795(.dinb(n8353), .dina(n3324), .dout(n3328));
    jand g0796(.dinb(n3136), .dina(n8347), .dout(n3332));
    jand g0797(.dinb(n3221), .dina(n3305), .dout(n3336));
    jand g0798(.dinb(n3260), .dina(n3336), .dout(n3340));
    jor g0799(.dinb(n8361), .dina(n3340), .dout(n3344));
    jand g0800(.dinb(n8364), .dina(n3344), .dout(n3348));
    jnot g0801(.din(G4528), .dout(n3351));
    jor g0802(.dinb(G1455), .dina(G2204), .dout(n3355));
    jor g0803(.dinb(n3351), .dina(n3355), .dout(n3359));
    jand g0804(.dinb(n12699), .dina(n3359), .dout(n3363));
    jor g0805(.dinb(n3309), .dina(n8323), .dout(n3367));
    jor g0806(.dinb(n3348), .dina(n8320), .dout(n3371));
    jor g0807(.dinb(n3332), .dina(n8311), .dout(n3375));
    jand g0808(.dinb(G1455), .dina(G2204), .dout(n3379));
    jor g0809(.dinb(n12696), .dina(n3351), .dout(n3383));
    jor g0810(.dinb(n8284), .dina(n3383), .dout(n3387));
    jand g0811(.dinb(n3375), .dina(n8281), .dout(n3391));
    jand g0812(.dinb(n14091), .dina(n537), .dout(n3395));
    jand g0813(.dinb(n659), .dina(n14199), .dout(n3399));
    jor g0814(.dinb(n13945), .dina(n3399), .dout(n3403));
    jand g0815(.dinb(n14184), .dina(n3403), .dout(n3407));
    jor g0816(.dinb(n14505), .dina(n639), .dout(n3411));
    jand g0817(.dinb(n3407), .dina(n8233), .dout(n3415));
    jxor g0818(.dinb(n14583), .dina(n3415), .dout(n3419));
    jand g0819(.dinb(n639), .dina(n3399), .dout(n3423));
    jxor g0820(.dinb(n14556), .dina(n3423), .dout(n3427));
    jand g0821(.dinb(n14208), .dina(n651), .dout(n3431));
    jand g0822(.dinb(n635), .dina(n13977), .dout(n3435));
    jxor g0823(.dinb(n14970), .dina(n3435), .dout(n3439));
    jor g0824(.dinb(n14404), .dina(n602), .dout(n3443));
    jand g0825(.dinb(n14211), .dina(n3443), .dout(n3447));
    jxor g0826(.dinb(n14286), .dina(n3447), .dout(n3451));
    jor g0827(.dinb(n707), .dina(n13644), .dout(n3455));
    jor g0828(.dinb(n14838), .dina(n3455), .dout(n3459));
    jand g0829(.dinb(n14121), .dina(n3459), .dout(n3463));
    jxor g0830(.dinb(n13623), .dina(n3463), .dout(n3467));
    jand g0831(.dinb(n14760), .dina(n3455), .dout(n3471));
    jxor g0832(.dinb(n14907), .dina(n3471), .dout(n3475));
    jand g0833(.dinb(n14805), .dina(n753), .dout(n3479));
    jor g0834(.dinb(n707), .dina(n14706), .dout(n3483));
    jand g0835(.dinb(n14775), .dina(n3483), .dout(n3487));
    jxor g0836(.dinb(n14724), .dina(n3487), .dout(n3491));
    jxor g0837(.dinb(n707), .dina(n13659), .dout(n3495));
    jxor g0838(.dinb(n1291), .dina(n1314), .dout(n3499));
    jxor g0839(.dinb(n1253), .dina(n1333), .dout(n3503));
    jxor g0840(.dinb(n12273), .dina(n3503), .dout(n3507));
    jnot g0841(.din(n1471), .dout(n3510));
    jor g0842(.dinb(n11814), .dina(n3510), .dout(n3514));
    jnot g0843(.din(n1456), .dout(n3517));
    jor g0844(.dinb(n3517), .dina(n11733), .dout(n3521));
    jand g0845(.dinb(n3514), .dina(n3521), .dout(n3525));
    jor g0846(.dinb(n11664), .dina(n1571), .dout(n3529));
    jor g0847(.dinb(n1564), .dina(n11637), .dout(n3533));
    jand g0848(.dinb(n3529), .dina(n3533), .dout(n3537));
    jxor g0849(.dinb(n3525), .dina(n3537), .dout(n3541));
    jnot g0850(.din(G141), .dout(n3544));
    jor g0851(.dinb(n9489), .dina(n3544), .dout(n3548));
    jnot g0852(.din(G161), .dout(n3551));
    jor g0853(.dinb(n455), .dina(n3551), .dout(n3555));
    jand g0854(.dinb(n3548), .dina(n3555), .dout(n3559));
    jxor g0855(.dinb(n3541), .dina(n9169), .dout(n3563));
    jxor g0856(.dinb(n9157), .dina(n3563), .dout(n3567));
    jxor g0857(.dinb(n9148), .dina(n3567), .dout(n3571));
    jand g0858(.dinb(n9378), .dina(n1245), .dout(n3575));
    jxor g0859(.dinb(G211), .dina(G212), .dout(n3579));
    jand g0860(.dinb(n3575), .dina(n9133), .dout(n3583));
    jor g0861(.dinb(n12318), .dina(n1662), .dout(n3587));
    jnot g0862(.din(n1598), .dout(n3590));
    jand g0863(.dinb(n3590), .dina(n1617), .dout(n3594));
    jnot g0864(.din(n1613), .dout(n3597));
    jand g0865(.dinb(n1602), .dina(n3597), .dout(n3601));
    jor g0866(.dinb(n3594), .dina(n3601), .dout(n3605));
    jor g0867(.dinb(n11265), .dina(n1725), .dout(n3609));
    jor g0868(.dinb(n1715), .dina(n11238), .dout(n3613));
    jand g0869(.dinb(n3609), .dina(n3613), .dout(n3617));
    jxor g0870(.dinb(n9127), .dina(n3617), .dout(n3621));
    jxor g0871(.dinb(n9124), .dina(n3621), .dout(n3625));
    jxor g0872(.dinb(n9112), .dina(n3625), .dout(n3629));
    jand g0873(.dinb(G18), .dina(G239), .dout(n3633));
    jand g0874(.dinb(n455), .dina(n9313), .dout(n3637));
    jor g0875(.dinb(n9100), .dina(n3637), .dout(n3641));
    jxor g0876(.dinb(n728), .dina(n779), .dout(n3645));
    jxor g0877(.dinb(n753), .dina(n806), .dout(n3649));
    jxor g0878(.dinb(n3645), .dina(n3649), .dout(n3653));
    jxor g0879(.dinb(n9097), .dina(n3653), .dout(n3657));
    jxor g0880(.dinb(n515), .dina(n623), .dout(n3661));
    jxor g0881(.dinb(n14568), .dina(n3661), .dout(n3665));
    jxor g0882(.dinb(n467), .dina(n569), .dout(n3669));
    jxor g0883(.dinb(n3665), .dina(n9091), .dout(n3673));
    jxor g0884(.dinb(n3657), .dina(n3673), .dout(n3677));
    jxor g0885(.dinb(n1088), .dina(n1130), .dout(n3681));
    jxor g0886(.dinb(n1107), .dina(n1149), .dout(n3685));
    jxor g0887(.dinb(n3681), .dina(n3685), .dout(n3689));
    jxor g0888(.dinb(n13389), .dina(n3689), .dout(n3693));
    jand g0889(.dinb(G18), .dina(G227), .dout(n3697));
    jand g0890(.dinb(n455), .dina(n9337), .dout(n3701));
    jor g0891(.dinb(n9088), .dina(n3701), .dout(n3705));
    jxor g0892(.dinb(n919), .dina(n961), .dout(n3709));
    jxor g0893(.dinb(n9085), .dina(n3709), .dout(n3713));
    jxor g0894(.dinb(n884), .dina(n903), .dout(n3717));
    jxor g0895(.dinb(n3713), .dina(n9082), .dout(n3721));
    jxor g0896(.dinb(n3693), .dina(n3721), .dout(n3725));
    jor g0897(.dinb(n3677), .dina(n3725), .dout(n3729));
    jor g0898(.dinb(n3629), .dina(n9079), .dout(n3733));
    jor g0899(.dinb(n3571), .dina(n3733), .dout(n3737));
    jxor g0900(.dinb(n2223), .dina(n2254), .dout(n3741));
    jxor g0901(.dinb(n2196), .dina(n2314), .dout(n3745));
    jxor g0902(.dinb(n9642), .dina(n3745), .dout(n3749));
    jxor g0903(.dinb(n2082), .dina(n2106), .dout(n3753));
    jxor g0904(.dinb(n2137), .dina(n2161), .dout(n3757));
    jxor g0905(.dinb(n3753), .dina(n3757), .dout(n3761));
    jor g0906(.dinb(n455), .dina(n9618), .dout(n3765));
    jnot g0907(.din(G58), .dout(n3768));
    jor g0908(.dinb(n14946), .dina(n3768), .dout(n3772));
    jand g0909(.dinb(n3765), .dina(n3772), .dout(n3776));
    jxor g0910(.dinb(n3761), .dina(n9616), .dout(n3780));
    jxor g0911(.dinb(n9610), .dina(n3780), .dout(n3784));
    jxor g0912(.dinb(n9607), .dina(n3784), .dout(n3788));
    jxor g0913(.dinb(n9591), .dina(n579), .dout(n3792));
    jor g0914(.dinb(n9621), .dina(n3792), .dout(n3796));
    jnot g0915(.din(G69), .dout(n3799));
    jand g0916(.dinb(n3799), .dina(n2646), .dout(n3803));
    jand g0917(.dinb(G69), .dina(G70), .dout(n3807));
    jor g0918(.dinb(n14946), .dina(n3807), .dout(n3811));
    jor g0919(.dinb(n3803), .dina(n3811), .dout(n3815));
    jand g0920(.dinb(n3796), .dina(n3815), .dout(n3819));
    jxor g0921(.dinb(n9595), .dina(n3819), .dout(n3823));
    jnot g0922(.din(n3823), .dout(n3826));
    jxor g0923(.dinb(n2631), .dina(n2695), .dout(n3830));
    jnot g0924(.din(n2590), .dout(n3833));
    jxor g0925(.dinb(n2412), .dina(n2445), .dout(n3837));
    jxor g0926(.dinb(n2495), .dina(n2522), .dout(n3841));
    jxor g0927(.dinb(n3837), .dina(n3841), .dout(n3845));
    jxor g0928(.dinb(n9526), .dina(n3845), .dout(n3849));
    jxor g0929(.dinb(n9523), .dina(n3849), .dout(n3853));
    jnot g0930(.din(n3853), .dout(n3856));
    jand g0931(.dinb(n9517), .dina(n3856), .dout(n3860));
    jand g0932(.dinb(n9585), .dina(n3853), .dout(n3864));
    jor g0933(.dinb(n455), .dina(n9510), .dout(n3868));
    jnot g0934(.din(G114), .dout(n3871));
    jor g0935(.dinb(n14946), .dina(n3871), .dout(n3875));
    jand g0936(.dinb(n3868), .dina(n3875), .dout(n3879));
    jxor g0937(.dinb(n3217), .dina(n3236), .dout(n3883));
    jxor g0938(.dinb(n9502), .dina(n3883), .dout(n3887));
    jxor g0939(.dinb(n3186), .dina(n3290), .dout(n3891));
    jxor g0940(.dinb(n9495), .dina(n3891), .dout(n3895));
    jxor g0941(.dinb(G1492), .dina(G1496), .dout(n3899));
    jor g0942(.dinb(n455), .dina(n3899), .dout(n3903));
    jxor g0943(.dinb(G1455), .dina(G2204), .dout(n3907));
    jor g0944(.dinb(n14943), .dina(n3907), .dout(n3911));
    jand g0945(.dinb(n3903), .dina(n3911), .dout(n3915));
    jxor g0946(.dinb(n3895), .dina(n9484), .dout(n3919));
    jxor g0947(.dinb(n9478), .dina(n3919), .dout(n3923));
    jxor g0948(.dinb(n2868), .dina(n2895), .dout(n3927));
    jxor g0949(.dinb(n2948), .dina(n2972), .dout(n3931));
    jxor g0950(.dinb(n3927), .dina(n3931), .dout(n3935));
    jxor g0951(.dinb(n9468), .dina(n3935), .dout(n3939));
    jor g0952(.dinb(n455), .dina(n9453), .dout(n3943));
    jnot g0953(.din(G82), .dout(n3946));
    jor g0954(.dinb(n14943), .dina(n3946), .dout(n3950));
    jand g0955(.dinb(n3943), .dina(n3950), .dout(n3954));
    jxor g0956(.dinb(n1932), .dina(n1971), .dout(n3958));
    jxor g0957(.dinb(n9445), .dina(n3958), .dout(n3962));
    jxor g0958(.dinb(n1878), .dina(n1905), .dout(n3966));
    jxor g0959(.dinb(n3962), .dina(n9436), .dout(n3970));
    jxor g0960(.dinb(n3939), .dina(n3970), .dout(n3974));
    jor g0961(.dinb(n3923), .dina(n3974), .dout(n3978));
    jor g0962(.dinb(n3864), .dina(n3978), .dout(n3982));
    jor g0963(.dinb(n3860), .dina(n3982), .dout(n3986));
    jor g0964(.dinb(n9433), .dina(n3986), .dout(n3990));
    jnot g0965(.din(n3140), .dout(n3993));
    jnot g0966(.din(G170), .dout(n3996));
    jand g0967(.dinb(n14943), .dina(n3996), .dout(n4000));
    jxor g0968(.dinb(n3167), .dina(n4000), .dout(n4004));
    jnot g0969(.din(n4004), .dout(n4007));
    jand g0970(.dinb(n9409), .dina(n4007), .dout(n4011));
    jand g0971(.dinb(n9414), .dina(n4004), .dout(n4015));
    jor g0972(.dinb(n12309), .dina(n4015), .dout(n4019));
    jor g0973(.dinb(n4011), .dina(n4019), .dout(n4023));
    jnot g0974(.din(n3202), .dout(n4026));
    jor g0975(.dinb(n4026), .dina(n9384), .dout(n4030));
    jnot g0976(.din(n3275), .dout(n4033));
    jor g0977(.dinb(n9393), .dina(n4033), .dout(n4037));
    jand g0978(.dinb(n4030), .dina(n4037), .dout(n4041));
    jxor g0979(.dinb(G164), .dina(G165), .dout(n4045));
    jand g0980(.dinb(n3575), .dina(n9376), .dout(n4049));
    jxor g0981(.dinb(n4041), .dina(n9370), .dout(n4053));
    jxor g0982(.dinb(n9364), .dina(n4053), .dout(n4057));
    jxor g0983(.dinb(n2070), .dina(n2094), .dout(n4061));
    jxor g0984(.dinb(n2122), .dina(n2149), .dout(n4065));
    jxor g0985(.dinb(n4061), .dina(n4065), .dout(n4069));
    jxor g0986(.dinb(n9354), .dina(n4069), .dout(n4073));
    jand g0987(.dinb(G18), .dina(G197), .dout(n4077));
    jor g0988(.dinb(n3701), .dina(n9334), .dout(n4081));
    jnot g0989(.din(n4081), .dout(n4084));
    jxor g0990(.dinb(n2208), .dina(n2239), .dout(n4088));
    jxor g0991(.dinb(n4084), .dina(n4088), .dout(n4092));
    jnot g0992(.din(n4092), .dout(n4095));
    jxor g0993(.dinb(n2181), .dina(n2299), .dout(n4099));
    jxor g0994(.dinb(n4095), .dina(n9319), .dout(n4103));
    jand g0995(.dinb(n9339), .dina(n4103), .dout(n4107));
    jor g0996(.dinb(n4057), .dina(n4107), .dout(n4111));
    jand g0997(.dinb(G18), .dina(G208), .dout(n4115));
    jor g0998(.dinb(n3637), .dina(n9310), .dout(n4119));
    jxor g0999(.dinb(n2397), .dina(n2430), .dout(n4123));
    jxor g1000(.dinb(n9297), .dina(n2510), .dout(n4127));
    jxor g1001(.dinb(n4123), .dina(n4127), .dout(n4131));
    jxor g1002(.dinb(n9289), .dina(n4131), .dout(n4135));
    jnot g1003(.din(n2575), .dout(n4138));
    jxor g1004(.dinb(n2616), .dina(n2683), .dout(n4142));
    jxor g1005(.dinb(n4138), .dina(n4142), .dout(n4146));
    jnot g1006(.din(G198), .dout(n4149));
    jor g1007(.dinb(n455), .dina(n4149), .dout(n4153));
    jand g1008(.dinb(n448), .dina(n4153), .dout(n4157));
    jxor g1009(.dinb(n2545), .dina(n9256), .dout(n4161));
    jxor g1010(.dinb(n4146), .dina(n9253), .dout(n4165));
    jand g1011(.dinb(n4135), .dina(n4165), .dout(n4169));
    jnot g1012(.din(n4073), .dout(n4172));
    jnot g1013(.din(n4103), .dout(n4175));
    jand g1014(.dinb(n9250), .dina(n4175), .dout(n4179));
    jnot g1015(.din(n4135), .dout(n4182));
    jnot g1016(.din(n4165), .dout(n4185));
    jand g1017(.dinb(n4182), .dina(n4185), .dout(n4189));
    jor g1018(.dinb(n4179), .dina(n4189), .dout(n4193));
    jor g1019(.dinb(n9247), .dina(n4193), .dout(n4197));
    jor g1020(.dinb(n9241), .dina(n4197), .dout(n4201));
    jxor g1021(.dinb(n1863), .dina(n1917), .dout(n4205));
    jxor g1022(.dinb(n9231), .dina(n4205), .dout(n4209));
    jxor g1023(.dinb(n1836), .dina(n1956), .dout(n4213));
    jnot g1024(.din(n2876), .dout(n4216));
    jand g1025(.dinb(n4216), .dina(n2960), .dout(n4220));
    jnot g1026(.din(n2956), .dout(n4223));
    jand g1027(.dinb(n2880), .dina(n4223), .dout(n4227));
    jor g1028(.dinb(n4220), .dina(n4227), .dout(n4231));
    jnot g1029(.din(n2849), .dout(n4234));
    jand g1030(.dinb(n4234), .dina(n2933), .dout(n4238));
    jnot g1031(.din(n2929), .dout(n4241));
    jand g1032(.dinb(n2853), .dina(n4241), .dout(n4245));
    jor g1033(.dinb(n4238), .dina(n4245), .dout(n4249));
    jxor g1034(.dinb(n4231), .dina(n4249), .dout(n4253));
    jnot g1035(.din(G181), .dout(n4256));
    jor g1036(.dinb(n455), .dina(n4256), .dout(n4260));
    jand g1037(.dinb(n3548), .dina(n4260), .dout(n4264));
    jxor g1038(.dinb(n4253), .dina(n9205), .dout(n4268));
    jxor g1039(.dinb(n9196), .dina(n4268), .dout(n4272));
    jxor g1040(.dinb(n9187), .dina(n4272), .dout(n4276));
    jor g1041(.dinb(n4201), .dina(n9178), .dout(n4280));
    jnot g1042(.din(n519), .dout(n4283));
    jxor g1043(.dinb(n14082), .dina(n537), .dout(n4287));
    jand g1044(.dinb(n4283), .dina(n14080), .dout(n4291));
    jnot g1045(.din(n573), .dout(n4294));
    jxor g1046(.dinb(n14037), .dina(n623), .dout(n4298));
    jand g1047(.dinb(n482), .dina(n14025), .dout(n4302));
    jand g1048(.dinb(n14466), .dina(n4302), .dout(n4306));
    jand g1049(.dinb(n14064), .dina(n4306), .dout(n4310));
    jand g1050(.dinb(n14073), .dina(n4310), .dout(n4314));
    jnot g1051(.din(n647), .dout(n4317));
    jand g1052(.dinb(n14335), .dina(n4298), .dout(n4321));
    jand g1053(.dinb(n4294), .dina(n4321), .dout(n4325));
    jor g1054(.dinb(n14023), .dina(n4325), .dout(n4329));
    jand g1055(.dinb(n14070), .dina(n4329), .dout(n4333));
    jnot g1056(.din(n671), .dout(n4336));
    jand g1057(.dinb(n4291), .dina(n4336), .dout(n4340));
    jnot g1058(.din(n695), .dout(n4343));
    jor g1059(.dinb(n4340), .dina(n4343), .dout(n4347));
    jor g1060(.dinb(n4333), .dina(n4347), .dout(n4351));
    jor g1061(.dinb(n4314), .dina(n4351), .dout(n4355));
    jnot g1062(.din(n818), .dout(n4358));
    jand g1063(.dinb(n4355), .dina(n12979), .dout(n4362));
    jnot g1064(.din(n865), .dout(n4365));
    jor g1065(.dinb(n4362), .dina(n4365), .dout(n4369));
    jand g1066(.dinb(n4369), .dina(n13416), .dout(n4373));
    jnot g1067(.din(n1069), .dout(n4376));
    jor g1068(.dinb(n4373), .dina(n4376), .dout(n4380));
    jand g1069(.dinb(n4380), .dina(n12408), .dout(n4384));
    jor g1070(.dinb(n4384), .dina(n12351), .dout(n4388));
    jxor g1071(.dinb(n4388), .dina(n12135), .dout(n4392));
    jand g1072(.dinb(n4388), .dina(n12057), .dout(n4396));
    jnot g1073(.din(n1441), .dout(n4399));
    jor g1074(.dinb(n4396), .dina(n10606), .dout(n4403));
    jand g1075(.dinb(n4403), .dina(n11598), .dout(n4407));
    jnot g1076(.din(n1587), .dout(n4410));
    jor g1077(.dinb(n4407), .dina(n10594), .dout(n4414));
    jxor g1078(.dinb(n4414), .dina(n11088), .dout(n4418));
    jor g1079(.dinb(n2729), .dina(n3028), .dout(n4422));
    jand g1080(.dinb(n8586), .dina(n4422), .dout(n4426));
    jor g1081(.dinb(n8598), .dina(n4426), .dout(n4430));
    jand g1082(.dinb(n8634), .dina(n4430), .dout(n4434));
    jor g1083(.dinb(n8658), .dina(n4434), .dout(n4438));
    jand g1084(.dinb(n8691), .dina(n4438), .dout(n4442));
    jor g1085(.dinb(n8721), .dina(n4442), .dout(n4446));
    jnot g1086(.din(n1257), .dout(n4449));
    jnot g1087(.din(n1318), .dout(n4452));
    jnot g1088(.din(n1337), .dout(n4455));
    jnot g1089(.din(n1299), .dout(n4458));
    jor g1090(.dinb(n1235), .dina(n9960), .dout(n4462));
    jor g1091(.dinb(n8833), .dina(n4462), .dout(n4466));
    jor g1092(.dinb(n8794), .dina(n4466), .dout(n4470));
    jand g1093(.dinb(n11877), .dina(n4470), .dout(n4474));
    jxor g1094(.dinb(n10017), .dina(n4474), .dout(n4478));
    jand g1095(.dinb(n11925), .dina(n4466), .dout(n4482));
    jxor g1096(.dinb(n8754), .dina(n4482), .dout(n4486));
    jnot g1097(.din(n1406), .dout(n4489));
    jnot g1098(.din(n1402), .dout(n4492));
    jand g1099(.dinb(n9958), .dina(n4492), .dout(n4496));
    jand g1100(.dinb(n4462), .dina(n9927), .dout(n4500));
    jxor g1101(.dinb(n8796), .dina(n4500), .dout(n4504));
    jand g1102(.dinb(n4388), .dina(n12183), .dout(n4508));
    jor g1103(.dinb(n11979), .dina(n4508), .dout(n4512));
    jxor g1104(.dinb(n12231), .dina(n4512), .dout(n4516));
    jnot g1105(.din(n1606), .dout(n4519));
    jnot g1106(.din(n1621), .dout(n4522));
    jnot g1107(.din(n1636), .dout(n4525));
    jnot g1108(.din(n1674), .dout(n4528));
    jor g1109(.dinb(n1591), .dina(n9004), .dout(n4532));
    jor g1110(.dinb(n9055), .dina(n4532), .dout(n4536));
    jor g1111(.dinb(n8923), .dina(n4536), .dout(n4540));
    jand g1112(.dinb(n10794), .dina(n4540), .dout(n4544));
    jxor g1113(.dinb(n10422), .dina(n4544), .dout(n4548));
    jnot g1114(.din(n1756), .dout(n4551));
    jand g1115(.dinb(n8869), .dina(n4536), .dout(n4555));
    jxor g1116(.dinb(n8871), .dina(n4555), .dout(n4559));
    jnot g1117(.din(n1748), .dout(n4562));
    jand g1118(.dinb(n8962), .dina(n4532), .dout(n4566));
    jxor g1119(.dinb(n9006), .dina(n4566), .dout(n4570));
    jand g1120(.dinb(n4414), .dina(n11040), .dout(n4574));
    jor g1121(.dinb(n10893), .dina(n4574), .dout(n4578));
    jxor g1122(.dinb(n11145), .dina(n4578), .dout(n4582));
    jor g1123(.dinb(n344), .dina(n392), .dout(n4586));
    jor g1124(.dinb(n368), .dina(n416), .dout(n4590));
    jor g1125(.dinb(n4586), .dina(n4590), .dout(n4594));
    jor g1126(.dinb(n3737), .dina(n9076), .dout(n4598));
    jor g1127(.dinb(n4280), .dina(n9058), .dout(n4602));
    jor g1128(.dinb(n9420), .dina(n4602), .dout(n4606));
    jnot g1129(.din(n1494), .dout(n4609));
    jnot g1130(.din(n1479), .dout(n4612));
    jor g1131(.dinb(n1445), .dina(n10101), .dout(n4616));
    jand g1132(.dinb(n11415), .dina(n4616), .dout(n4620));
    jor g1133(.dinb(n11361), .dina(n4620), .dout(n4624));
    jand g1134(.dinb(n11502), .dina(n4624), .dout(n4628));
    jxor g1135(.dinb(n10164), .dina(n4628), .dout(n4632));
    jnot g1136(.din(n1509), .dout(n4635));
    jxor g1137(.dinb(n9763), .dina(n4620), .dout(n4639));
    jand g1138(.dinb(n11754), .dina(n3510), .dout(n4643));
    jnot g1139(.din(n4643), .dout(n4646));
    jand g1140(.dinb(n4403), .dina(n10230), .dout(n4650));
    jor g1141(.dinb(n11457), .dina(n4650), .dout(n4654));
    jxor g1142(.dinb(n11766), .dina(n4654), .dout(n4658));
    jxor g1143(.dinb(n4403), .dina(n11691), .dout(n4662));
    jxor g1144(.dinb(n4369), .dina(n13440), .dout(n4666));
    jnot g1145(.din(n1803), .dout(n4669));
    jnot g1146(.din(n494), .dout(n4672));
    jor g1147(.dinb(n1788), .dina(n1792), .dout(n4676));
    jxor g1148(.dinb(n4672), .dina(n12619), .dout(n4680));
    jnot g1149(.din(n4680), .dout(n4683));
    jor g1150(.dinb(n4669), .dina(n10515), .dout(n4687));
    jand g1151(.dinb(n9768), .dina(n4687), .dout(n4691));
    jxor g1152(.dinb(n1785), .dina(n10663), .dout(n4695));
    jnot g1153(.din(n888), .dout(n4698));
    jnot g1154(.din(n949), .dout(n4701));
    jnot g1155(.din(n968), .dout(n4704));
    jnot g1156(.din(n930), .dout(n4707));
    jor g1157(.dinb(n869), .dina(n12825), .dout(n4711));
    jor g1158(.dinb(n9823), .dina(n4711), .dout(n4715));
    jor g1159(.dinb(n9799), .dina(n4715), .dout(n4719));
    jand g1160(.dinb(n13317), .dina(n4719), .dout(n4723));
    jxor g1161(.dinb(n12882), .dina(n4723), .dout(n4727));
    jand g1162(.dinb(n13341), .dina(n4715), .dout(n4731));
    jxor g1163(.dinb(n9771), .dina(n4731), .dout(n4735));
    jand g1164(.dinb(n13362), .dina(n1030), .dout(n4739));
    jand g1165(.dinb(n4711), .dina(n12807), .dout(n4743));
    jxor g1166(.dinb(n9801), .dina(n4743), .dout(n4747));
    jnot g1167(.din(n1026), .dout(n4750));
    jand g1168(.dinb(n4369), .dina(n13470), .dout(n4754));
    jor g1169(.dinb(n12861), .dina(n4754), .dout(n4758));
    jxor g1170(.dinb(n13515), .dina(n4758), .dout(n4762));
    jand g1171(.dinb(n4380), .dina(n12471), .dout(n4766));
    jand g1172(.dinb(n13212), .dina(n4766), .dout(n4770));
    jor g1173(.dinb(n12948), .dina(n4770), .dout(n4774));
    jxor g1174(.dinb(n12432), .dina(n4774), .dout(n4778));
    jor g1175(.dinb(n13089), .dina(n4766), .dout(n4782));
    jxor g1176(.dinb(n13740), .dina(n4782), .dout(n4786));
    jnot g1177(.din(n1107), .dout(n4789));
    jand g1178(.dinb(n13167), .dina(n4789), .dout(n4793));
    jnot g1179(.din(n4793), .dout(n4796));
    jand g1180(.dinb(n4380), .dina(n12999), .dout(n4800));
    jor g1181(.dinb(n13116), .dina(n4800), .dout(n4804));
    jxor g1182(.dinb(n13029), .dina(n4804), .dout(n4808));
    jxor g1183(.dinb(n4380), .dina(n12498), .dout(n4812));
    jxor g1184(.dinb(n1318), .dina(n1337), .dout(n4816));
    jxor g1185(.dinb(n11634), .dina(n4816), .dout(n4820));
    jnot g1186(.din(n1460), .dout(n4823));
    jnot g1187(.din(n1575), .dout(n4826));
    jand g1188(.dinb(n4826), .dina(n1554), .dout(n4830));
    jor g1189(.dinb(n1561), .dina(n10156), .dout(n4834));
    jxor g1190(.dinb(n10213), .dina(n4834), .dout(n4838));
    jxor g1191(.dinb(n10215), .dina(n4838), .dout(n4842));
    jxor g1192(.dinb(n10264), .dina(n4842), .dout(n4846));
    jand g1193(.dinb(n1445), .dina(n10153), .dout(n4850));
    jxor g1194(.dinb(n4823), .dina(n11454), .dout(n4854));
    jand g1195(.dinb(n10135), .dina(n1557), .dout(n4858));
    jnot g1196(.din(n4858), .dout(n4861));
    jor g1197(.dinb(n11550), .dina(n4861), .dout(n4865));
    jor g1198(.dinb(n11406), .dina(n4858), .dout(n4869));
    jand g1199(.dinb(n4865), .dina(n10099), .dout(n4873));
    jxor g1200(.dinb(n10158), .dina(n4873), .dout(n4877));
    jxor g1201(.dinb(n10096), .dina(n4877), .dout(n4881));
    jand g1202(.dinb(n4403), .dina(n10078), .dout(n4885));
    jor g1203(.dinb(n4850), .dina(n4885), .dout(n4889));
    jand g1204(.dinb(n11967), .dina(n1425), .dout(n4893));
    jnot g1205(.din(n1398), .dout(n4896));
    jand g1206(.dinb(n10062), .dina(n1394), .dout(n4900));
    jand g1207(.dinb(n11955), .dina(n4900), .dout(n4904));
    jxor g1208(.dinb(n12171), .dina(n4904), .dout(n4908));
    jor g1209(.dinb(n4893), .dina(n4908), .dout(n4912));
    jor g1210(.dinb(n12286), .dina(n1272), .dout(n4916));
    jand g1211(.dinb(n10015), .dina(n4896), .dout(n4920));
    jor g1212(.dinb(n11961), .dina(n4920), .dout(n4924));
    jxor g1213(.dinb(n1433), .dina(n10012), .dout(n4928));
    jxor g1214(.dinb(n10060), .dina(n4928), .dout(n4932));
    jxor g1215(.dinb(n10003), .dina(n4932), .dout(n4936));
    jor g1216(.dinb(n4388), .dina(n9997), .dout(n4940));
    jand g1217(.dinb(n9988), .dina(n4496), .dout(n4944));
    jxor g1218(.dinb(n12288), .dina(n4944), .dout(n4948));
    jxor g1219(.dinb(n1276), .dina(n1398), .dout(n4952));
    jand g1220(.dinb(n1299), .dina(n12084), .dout(n4956));
    jor g1221(.dinb(n1422), .dina(n9925), .dout(n4960));
    jnot g1222(.din(n4960), .dout(n4963));
    jand g1223(.dinb(n12018), .dina(n4963), .dout(n4967));
    jnot g1224(.din(n1345), .dout(n4970));
    jand g1225(.dinb(n9922), .dina(n4960), .dout(n4974));
    jand g1226(.dinb(n1433), .dina(n9919), .dout(n4978));
    jor g1227(.dinb(n9916), .dina(n4978), .dout(n4982));
    jxor g1228(.dinb(n9913), .dina(n4982), .dout(n4986));
    jxor g1229(.dinb(n9892), .dina(n4986), .dout(n4990));
    jor g1230(.dinb(n1235), .dina(n9880), .dout(n4994));
    jand g1231(.dinb(n4940), .dina(n4994), .dout(n4998));
    jxor g1232(.dinb(n4889), .dina(n9874), .dout(n5002));
    jxor g1233(.dinb(n9868), .dina(n5002), .dout(n5006));
    jand g1234(.dinb(n1785), .dina(n10663), .dout(n5010));
    jor g1235(.dinb(n12561), .dina(n5010), .dout(n5014));
    jnot g1236(.din(n1689), .dout(n5017));
    jand g1237(.dinb(n4414), .dina(n10722), .dout(n5021));
    jand g1238(.dinb(n1781), .dina(n10665), .dout(n5025));
    jor g1239(.dinb(n10570), .dina(n5025), .dout(n5029));
    jor g1240(.dinb(n5021), .dina(n10513), .dout(n5033));
    jor g1241(.dinb(n5017), .dina(n5033), .dout(n5037));
    jand g1242(.dinb(n5014), .dina(n10504), .dout(n5041));
    jand g1243(.dinb(n1778), .dina(n12528), .dout(n5045));
    jand g1244(.dinb(n1591), .dina(n10501), .dout(n5049));
    jor g1245(.dinb(n5041), .dina(n10489), .dout(n5053));
    jxor g1246(.dinb(n1621), .dina(n1636), .dout(n5057));
    jor g1247(.dinb(n10965), .dina(n1756), .dout(n5061));
    jand g1248(.dinb(n1763), .dina(n10408), .dout(n5065));
    jxor g1249(.dinb(n10410), .dina(n5065), .dout(n5069));
    jor g1250(.dinb(n11143), .dina(n1666), .dout(n5073));
    jxor g1251(.dinb(n1655), .dina(n5073), .dout(n5077));
    jxor g1252(.dinb(n1748), .dina(n10405), .dout(n5081));
    jxor g1253(.dinb(n5069), .dina(n10399), .dout(n5085));
    jand g1254(.dinb(n1591), .dina(n10384), .dout(n5089));
    jand g1255(.dinb(n1722), .dina(n11037), .dout(n5093));
    jor g1256(.dinb(n1756), .dina(n10366), .dout(n5097));
    jor g1257(.dinb(n10963), .dina(n5097), .dout(n5101));
    jnot g1258(.din(n5097), .dout(n5104));
    jor g1259(.dinb(n11016), .dina(n5104), .dout(n5108));
    jor g1260(.dinb(n1770), .dina(n10360), .dout(n5112));
    jand g1261(.dinb(n10357), .dina(n5112), .dout(n5116));
    jor g1262(.dinb(n11031), .dina(n1748), .dout(n5120));
    jxor g1263(.dinb(n10477), .dina(n5120), .dout(n5124));
    jxor g1264(.dinb(n5116), .dina(n10348), .dout(n5128));
    jxor g1265(.dinb(n10857), .dina(n5128), .dout(n5132));
    jxor g1266(.dinb(n11199), .dina(n5132), .dout(n5136));
    jand g1267(.dinb(n4414), .dina(n10330), .dout(n5140));
    jor g1268(.dinb(n5089), .dina(n5140), .dout(n5144));
    jxor g1269(.dinb(n10324), .dina(n5144), .dout(n5148));
    jxor g1270(.dinb(n5053), .dina(n10273), .dout(G338));
    jxor g1271(.dinb(n13704), .dina(n968), .dout(n5156));
    jxor g1272(.dinb(n13734), .dina(n5156), .dout(n5160));
    jnot g1273(.din(n1134), .dout(n5163));
    jnot g1274(.din(n1216), .dout(n5166));
    jor g1275(.dinb(n13087), .dina(n1212), .dout(n5170));
    jand g1276(.dinb(n5166), .dina(n13078), .dout(n5174));
    jxor g1277(.dinb(n13075), .dina(n5174), .dout(n5178));
    jxor g1278(.dinb(n13023), .dina(n4796), .dout(n5182));
    jxor g1279(.dinb(n5178), .dina(n12997), .dout(n5186));
    jand g1280(.dinb(n1073), .dina(n12988), .dout(n5190));
    jxor g1281(.dinb(n1092), .dina(n1204), .dout(n5194));
    jxor g1282(.dinb(n13248), .dina(n5194), .dout(n5198));
    jand g1283(.dinb(n13179), .dina(n4796), .dout(n5202));
    jor g1284(.dinb(n13185), .dina(n5202), .dout(n5206));
    jnot g1285(.din(n5206), .dout(n5209));
    jand g1286(.dinb(n12945), .dina(n5209), .dout(n5213));
    jand g1287(.dinb(n13239), .dina(n5206), .dout(n5217));
    jor g1288(.dinb(n5213), .dina(n12943), .dout(n5221));
    jxor g1289(.dinb(n12940), .dina(n5221), .dout(n5225));
    jand g1290(.dinb(n4380), .dina(n12925), .dout(n5229));
    jor g1291(.dinb(n5190), .dina(n5229), .dout(n5233));
    jor g1292(.dinb(n13555), .dina(n903), .dout(n5237));
    jand g1293(.dinb(n12919), .dina(n1026), .dout(n5241));
    jor g1294(.dinb(n13365), .dina(n5241), .dout(n5245));
    jnot g1295(.din(n1061), .dout(n5248));
    jnot g1296(.din(n1053), .dout(n5251));
    jor g1297(.dinb(n13371), .dina(n5251), .dout(n5255));
    jor g1298(.dinb(n4750), .dina(n13387), .dout(n5259));
    jor g1299(.dinb(n13359), .dina(n5259), .dout(n5263));
    jxor g1300(.dinb(n13461), .dina(n5263), .dout(n5267));
    jand g1301(.dinb(n5255), .dina(n12859), .dout(n5271));
    jxor g1302(.dinb(n12913), .dina(n5271), .dout(n5275));
    jxor g1303(.dinb(n12916), .dina(n5275), .dout(n5279));
    jxor g1304(.dinb(n12856), .dina(n5279), .dout(n5283));
    jor g1305(.dinb(n12972), .dina(n5283), .dout(n5287));
    jand g1306(.dinb(n4707), .dina(n4739), .dout(n5291));
    jxor g1307(.dinb(n13557), .dina(n5291), .dout(n5295));
    jxor g1308(.dinb(n13512), .dina(n1026), .dout(n5299));
    jand g1309(.dinb(n930), .dina(n13683), .dout(n5303));
    jor g1310(.dinb(n5251), .dina(n12805), .dout(n5307));
    jor g1311(.dinb(n13392), .dina(n5307), .dout(n5311));
    jnot g1312(.din(n5307), .dout(n5314));
    jor g1313(.dinb(n13428), .dina(n5314), .dout(n5318));
    jor g1314(.dinb(n12916), .dina(n5318), .dout(n5322));
    jand g1315(.dinb(n12799), .dina(n5322), .dout(n5326));
    jxor g1316(.dinb(n12793), .dina(n5326), .dout(n5330));
    jxor g1317(.dinb(n12769), .dina(n5330), .dout(n5334));
    jor g1318(.dinb(n13602), .dina(n5334), .dout(n5338));
    jand g1319(.dinb(n12751), .dina(n5338), .dout(n5342));
    jxor g1320(.dinb(n12745), .dina(n5342), .dout(n5346));
    jxor g1321(.dinb(n12739), .dina(n5346), .dout(n5350));
    jxor g1322(.dinb(n4294), .dina(n14932), .dout(n5354));
    jnot g1323(.din(n829), .dout(n5357));
    jnot g1324(.din(n849), .dout(n5360));
    jor g1325(.dinb(n14749), .dina(n5360), .dout(n5364));
    jand g1326(.dinb(n14757), .dina(n5364), .dout(n5368));
    jxor g1327(.dinb(n14859), .dina(n5368), .dout(n5372));
    jnot g1328(.din(n5372), .dout(n5375));
    jxor g1329(.dinb(n732), .dina(n3479), .dout(n5379));
    jnot g1330(.din(n5379), .dout(n5382));
    jor g1331(.dinb(n5375), .dina(n14689), .dout(n5386));
    jor g1332(.dinb(n5372), .dina(n14691), .dout(n5390));
    jand g1333(.dinb(n14151), .dina(n5390), .dout(n5394));
    jand g1334(.dinb(n5386), .dina(n5394), .dout(n5398));
    jxor g1335(.dinb(n732), .dina(n841), .dout(n5402));
    jxor g1336(.dinb(n794), .dina(n14149), .dout(n5406));
    jnot g1337(.din(n857), .dout(n5409));
    jor g1338(.dinb(n732), .dina(n3479), .dout(n5413));
    jand g1339(.dinb(n14821), .dina(n5413), .dout(n5417));
    jand g1340(.dinb(n5409), .dina(n14112), .dout(n5421));
    jnot g1341(.din(n5421), .dout(n5424));
    jnot g1342(.din(n833), .dout(n5427));
    jor g1343(.dinb(n5427), .dina(n5417), .dout(n5431));
    jand g1344(.dinb(n5424), .dina(n14110), .dout(n5435));
    jor g1345(.dinb(n14133), .dina(n5435), .dout(n5439));
    jnot g1346(.din(n5406), .dout(n5442));
    jnot g1347(.din(n5435), .dout(n5445));
    jor g1348(.dinb(n14008), .dina(n5445), .dout(n5449));
    jand g1349(.dinb(n14010), .dina(n5449), .dout(n5453));
    jand g1350(.dinb(n13993), .dina(n5453), .dout(n5457));
    jor g1351(.dinb(n13987), .dina(n5457), .dout(n5461));
    jand g1352(.dinb(n631), .dina(n3431), .dout(n5465));
    jnot g1353(.din(n5465), .dout(n5468));
    jor g1354(.dinb(n3399), .dina(n5468), .dout(n5472));
    jnot g1355(.din(n3399), .dout(n5475));
    jand g1356(.dinb(n14967), .dina(n4302), .dout(n5479));
    jor g1357(.dinb(n5475), .dina(n13966), .dout(n5483));
    jor g1358(.dinb(n13968), .dina(n5483), .dout(n5487));
    jand g1359(.dinb(n13960), .dina(n5487), .dout(n5491));
    jxor g1360(.dinb(n14625), .dina(n5491), .dout(n5495));
    jnot g1361(.din(n5483), .dout(n5498));
    jor g1362(.dinb(n13926), .dina(n5498), .dout(n5502));
    jand g1363(.dinb(n14160), .dina(n5502), .dout(n5506));
    jxor g1364(.dinb(n14259), .dina(n5506), .dout(n5510));
    jxor g1365(.dinb(n14217), .dina(n5510), .dout(n5514));
    jnot g1366(.din(n5514), .dout(n5517));
    jand g1367(.dinb(n13947), .dina(n5517), .dout(n5521));
    jnot g1368(.din(n5495), .dout(n5524));
    jand g1369(.dinb(n13924), .dina(n5514), .dout(n5528));
    jor g1370(.dinb(n14358), .dina(n5528), .dout(n5532));
    jor g1371(.dinb(n5521), .dina(n5532), .dout(n5536));
    jxor g1372(.dinb(n14607), .dina(n3407), .dout(n5540));
    jand g1373(.dinb(n14248), .dina(n647), .dout(n5544));
    jand g1374(.dinb(n671), .dina(n5544), .dout(n5548));
    jand g1375(.dinb(n14310), .dina(n5548), .dout(n5552));
    jnot g1376(.din(n5548), .dout(n5555));
    jand g1377(.dinb(n14319), .dina(n5475), .dout(n5559));
    jor g1378(.dinb(n14046), .dina(n5559), .dout(n5563));
    jand g1379(.dinb(n13909), .dina(n5563), .dout(n5567));
    jor g1380(.dinb(n13897), .dina(n5567), .dout(n5571));
    jand g1381(.dinb(n14028), .dina(n623), .dout(n5575));
    jor g1382(.dinb(n14335), .dina(n5575), .dout(n5579));
    jand g1383(.dinb(n14205), .dina(n5579), .dout(n5583));
    jxor g1384(.dinb(n5571), .dina(n13882), .dout(n5587));
    jnot g1385(.din(n5587), .dout(n5590));
    jand g1386(.dinb(n13911), .dina(n5590), .dout(n5594));
    jnot g1387(.din(n5540), .dout(n5597));
    jand g1388(.dinb(n13861), .dina(n5587), .dout(n5601));
    jor g1389(.dinb(n14421), .dina(n5601), .dout(n5605));
    jor g1390(.dinb(n5594), .dina(n5605), .dout(n5609));
    jand g1391(.dinb(n5536), .dina(n13855), .dout(n5613));
    jxor g1392(.dinb(n14514), .dina(n5613), .dout(n5617));
    jxor g1393(.dinb(n13852), .dina(n5617), .dout(n5621));
    jxor g1394(.dinb(n13843), .dina(n5621), .dout(n5625));
    jdff g1395(.din(G1), .dout(n5628));
    jdff g1396(.din(G1), .dout(n5631));
    jdff g1397(.din(G1459), .dout(n5634));
    jdff g1398(.din(G1469), .dout(n5637));
    jdff g1399(.din(G1480), .dout(n5640));
    jdff g1400(.din(G1486), .dout(n5643));
    jdff g1401(.din(G1492), .dout(n5646));
    jdff g1402(.din(G1496), .dout(n5649));
    jdff g1403(.din(G2208), .dout(n5652));
    jdff g1404(.din(G2218), .dout(n5655));
    jdff g1405(.din(G2224), .dout(n5658));
    jdff g1406(.din(G2230), .dout(n5661));
    jdff g1407(.din(G2236), .dout(n5664));
    jdff g1408(.din(G2239), .dout(n5667));
    jdff g1409(.din(G2247), .dout(n5670));
    jdff g1410(.din(G2253), .dout(n5673));
    jdff g1411(.din(G2256), .dout(n5676));
    jdff g1412(.din(G3698), .dout(n5679));
    jdff g1413(.din(G3701), .dout(n5682));
    jdff g1414(.din(G3705), .dout(n5685));
    jdff g1415(.din(G3711), .dout(n5688));
    jdff g1416(.din(G3717), .dout(n5691));
    jdff g1417(.din(G3723), .dout(n5694));
    jdff g1418(.din(G3729), .dout(n5697));
    jdff g1419(.din(G3737), .dout(n5700));
    jdff g1420(.din(G3743), .dout(n5703));
    jdff g1421(.din(G3749), .dout(n5706));
    jdff g1422(.din(G4393), .dout(n5709));
    jdff g1423(.din(G4400), .dout(n5712));
    jdff g1424(.din(G4405), .dout(n5715));
    jdff g1425(.din(G4410), .dout(n5718));
    jdff g1426(.din(G4415), .dout(n5721));
    jdff g1427(.din(G4420), .dout(n5724));
    jdff g1428(.din(G4427), .dout(n5727));
    jdff g1429(.din(G4432), .dout(n5730));
    jdff g1430(.din(G4437), .dout(n5733));
    jdff g1431(.din(G1462), .dout(n5736));
    jdff g1432(.din(G2211), .dout(n5739));
    jdff g1433(.din(G4394), .dout(n5742));
    jdff g1434(.din(G1), .dout(n5745));
    jdff g1435(.din(G106), .dout(n5748));
    jnot g1436(.din(G15), .dout(n5751));
    jor g1437(.dinb(n8229), .dina(n419), .dout(n5755));
    jnot g1438(.din(G15), .dout(n5758));
    jor g1439(.dinb(n8223), .dina(n433), .dout(n5762));
    jdff g1440(.din(G1), .dout(n5765));
    jand g1441(.dinb(n3375), .dina(n8281), .dout(n5769));
    jor g1442(.dinb(n1810), .dina(n9715), .dout(n5773));
    jand g1443(.dinb(n3375), .dina(n8281), .dout(n5777));
    jor g1444(.dinb(n1810), .dina(n9715), .dout(n5781));
    jor g1445(.dinb(n1810), .dina(n9715), .dout(n5785));
    jand g1446(.dinb(n9765), .dina(n4687), .dout(n5789));
    jxor g1447(.dinb(n1785), .dina(n10663), .dout(n5793));
    jdff dff_A_BG2uy8SX9_0(.din(n20592), .dout(G399));
    jdff dff_A_uh82oImW5_0(.din(n20589), .dout(n20592));
    jdff dff_A_tlVoCh1Z5_0(.din(n20586), .dout(n20589));
    jdff dff_A_LeXqoUCC1_0(.din(n20583), .dout(n20586));
    jdff dff_A_neBD5Ml89_2(.din(n5625), .dout(n20583));
    jdff dff_A_T0RPmTc91_0(.din(n20577), .dout(G370));
    jdff dff_A_reD76IVv3_0(.din(n20574), .dout(n20577));
    jdff dff_A_8x9IJLGt1_0(.din(n20571), .dout(n20574));
    jdff dff_A_Y0TP6KzS4_0(.din(n20568), .dout(n20571));
    jdff dff_A_5B511Ywc8_0(.din(n20565), .dout(n20568));
    jdff dff_A_yDtmijmt8_0(.din(n20562), .dout(n20565));
    jdff dff_A_p7vnaGTp4_2(.din(n5350), .dout(n20562));
    jdff dff_A_LEzamXti6_0(.din(n20556), .dout(G321));
    jdff dff_A_jfawbR8f2_0(.din(n20553), .dout(n20556));
    jdff dff_A_IOZH2WS93_0(.din(n20550), .dout(n20553));
    jdff dff_A_PtgjT43b1_0(.din(n20547), .dout(n20550));
    jdff dff_A_O0ichDPW1_2(.din(n5006), .dout(n20547));
    jdff dff_A_nv0Y42PX8_0(.din(n20541), .dout(G356));
    jdff dff_A_y6MjP8Qb8_0(.din(n20538), .dout(n20541));
    jdff dff_A_38FS1zn56_0(.din(n20535), .dout(n20538));
    jdff dff_A_OsqvV3eo7_0(.din(n20532), .dout(n20535));
    jdff dff_A_XiIHYqRH8_0(.din(n20529), .dout(n20532));
    jdff dff_A_E1az6nZ82_0(.din(n20526), .dout(n20529));
    jdff dff_A_QWZOHusX0_0(.din(n20523), .dout(n20526));
    jdff dff_A_dAgHZCA45_0(.din(n20520), .dout(n20523));
    jdff dff_A_7BPlkgWi9_0(.din(n20517), .dout(n20520));
    jdff dff_A_tIzFAeLt4_0(.din(n20514), .dout(n20517));
    jdff dff_A_mOswMUxg3_0(.din(n20511), .dout(n20514));
    jdff dff_A_ypcAw9sg9_2(.din(n4812), .dout(n20511));
    jdff dff_A_rw5qINAa0_0(.din(n20505), .dout(G353));
    jdff dff_A_Z3sOWuaz0_0(.din(n20502), .dout(n20505));
    jdff dff_A_0iF253ta6_0(.din(n20499), .dout(n20502));
    jdff dff_A_ea7jBFts1_0(.din(n20496), .dout(n20499));
    jdff dff_A_ieoW1bNp6_0(.din(n20493), .dout(n20496));
    jdff dff_A_WrKJH55W6_0(.din(n20490), .dout(n20493));
    jdff dff_A_ALy7YhUb2_0(.din(n20487), .dout(n20490));
    jdff dff_A_21VOdRlb4_0(.din(n20484), .dout(n20487));
    jdff dff_A_9ybG1xG72_0(.din(n20481), .dout(n20484));
    jdff dff_A_P8hPtzqU4_2(.din(n4808), .dout(n20481));
    jdff dff_A_CzzP5pjZ0_0(.din(n20475), .dout(G350));
    jdff dff_A_6Y8UhFqg3_0(.din(n20472), .dout(n20475));
    jdff dff_A_GjlOPqmp8_0(.din(n20469), .dout(n20472));
    jdff dff_A_VIktzUjc1_0(.din(n20466), .dout(n20469));
    jdff dff_A_IVFAHnMD3_0(.din(n20463), .dout(n20466));
    jdff dff_A_9iZodpNr8_0(.din(n20460), .dout(n20463));
    jdff dff_A_pZELC5nk3_0(.din(n20457), .dout(n20460));
    jdff dff_A_Ab0KCW1j2_0(.din(n20454), .dout(n20457));
    jdff dff_A_ghteABgK6_0(.din(n20451), .dout(n20454));
    jdff dff_A_djG7tKrZ7_2(.din(n4786), .dout(n20451));
    jdff dff_A_dx0HSNzG9_0(.din(n20445), .dout(G347));
    jdff dff_A_ekUOwAko3_0(.din(n20442), .dout(n20445));
    jdff dff_A_Q58gQSBR2_0(.din(n20439), .dout(n20442));
    jdff dff_A_lxkcQEtM0_0(.din(n20436), .dout(n20439));
    jdff dff_A_psKGp7Cq9_0(.din(n20433), .dout(n20436));
    jdff dff_A_GRpvyfWq5_0(.din(n20430), .dout(n20433));
    jdff dff_A_zXS4Xfyi0_0(.din(n20427), .dout(n20430));
    jdff dff_A_3PbZ1Jbq8_0(.din(n20424), .dout(n20427));
    jdff dff_A_VimgZs4n3_2(.din(n4778), .dout(n20424));
    jdff dff_A_mPaS6Mha1_0(.din(n20418), .dout(G368));
    jdff dff_A_cHjh7vKg0_0(.din(n20415), .dout(n20418));
    jdff dff_A_kJM8BYLq2_0(.din(n20412), .dout(n20415));
    jdff dff_A_0T8uOQtH3_0(.din(n20409), .dout(n20412));
    jdff dff_A_1HCHJbDg8_0(.din(n20406), .dout(n20409));
    jdff dff_A_3e1Lm0s86_0(.din(n20403), .dout(n20406));
    jdff dff_A_AOsmoC2R4_0(.din(n20400), .dout(n20403));
    jdff dff_A_jVXSzJcQ9_0(.din(n20397), .dout(n20400));
    jdff dff_A_RMkVxy4D8_0(.din(n20394), .dout(n20397));
    jdff dff_A_5waj8wW36_0(.din(n20391), .dout(n20394));
    jdff dff_A_bTLj5nNy8_0(.din(n20388), .dout(n20391));
    jdff dff_A_BRr7V1Dd0_2(.din(n4762), .dout(n20388));
    jdff dff_A_LLUDcLli2_0(.din(n20382), .dout(G365));
    jdff dff_A_4YZ7HJAB9_0(.din(n20379), .dout(n20382));
    jdff dff_A_HdHLYKd25_0(.din(n20376), .dout(n20379));
    jdff dff_A_oQuZ9C3o7_0(.din(n20373), .dout(n20376));
    jdff dff_A_Gb0kjhg59_0(.din(n20370), .dout(n20373));
    jdff dff_A_hdHDfOPH7_0(.din(n20367), .dout(n20370));
    jdff dff_A_EklCC1Fx2_0(.din(n20364), .dout(n20367));
    jdff dff_A_ZZ2Y7ZiW0_0(.din(n20361), .dout(n20364));
    jdff dff_A_ugyj3iQ65_0(.din(n20358), .dout(n20361));
    jdff dff_A_73WPHF0a8_0(.din(n20355), .dout(n20358));
    jdff dff_A_FBPSAZrq3_0(.din(n20352), .dout(n20355));
    jdff dff_A_OEN3E7xB2_2(.din(n4747), .dout(n20352));
    jdff dff_A_6FJsb1lw2_0(.din(n20346), .dout(G362));
    jdff dff_A_dqPJ984U6_0(.din(n20343), .dout(n20346));
    jdff dff_A_SphUPevv8_0(.din(n20340), .dout(n20343));
    jdff dff_A_z4W1hAW05_0(.din(n20337), .dout(n20340));
    jdff dff_A_HRaAPMWW8_0(.din(n20334), .dout(n20337));
    jdff dff_A_5dlFzehl4_0(.din(n20331), .dout(n20334));
    jdff dff_A_m5y08wEu6_0(.din(n20328), .dout(n20331));
    jdff dff_A_FiiC9BSW1_0(.din(n20325), .dout(n20328));
    jdff dff_A_aaoXjhMP0_0(.din(n20322), .dout(n20325));
    jdff dff_A_zgWesmuJ1_0(.din(n20319), .dout(n20322));
    jdff dff_A_QxgVD2QB2_2(.din(n4735), .dout(n20319));
    jdff dff_A_Xe1ad79S1_0(.din(n20313), .dout(G359));
    jdff dff_A_AQx62qQL1_0(.din(n20310), .dout(n20313));
    jdff dff_A_i45KJBzy6_0(.din(n20307), .dout(n20310));
    jdff dff_A_J5yOHCRL9_0(.din(n20304), .dout(n20307));
    jdff dff_A_gi4w7YCi8_0(.din(n20301), .dout(n20304));
    jdff dff_A_U7c5MoiX0_0(.din(n20298), .dout(n20301));
    jdff dff_A_bwLEuQlq6_0(.din(n20295), .dout(n20298));
    jdff dff_A_zB9ZqTqK2_0(.din(n20292), .dout(n20295));
    jdff dff_A_j9wtRz0k2_0(.din(n20289), .dout(n20292));
    jdff dff_A_Qutbbi7W3_2(.din(n4727), .dout(n20289));
    jdff dff_A_QzOwvaFh3_0(.din(n20283), .dout(G471));
    jdff dff_A_arKIhtye4_0(.din(n20280), .dout(n20283));
    jdff dff_A_wfUaDLW66_0(.din(n20277), .dout(n20280));
    jdff dff_A_E8jalRTs2_2(.din(n5793), .dout(n20277));
    jdff dff_A_EoeqTSWy8_0(.din(n20271), .dout(G419));
    jdff dff_A_ikIdkQUw3_0(.din(n20268), .dout(n20271));
    jdff dff_A_TeChXTMa7_0(.din(n20265), .dout(n20268));
    jdff dff_A_pN6IxNGh5_2(.din(n4695), .dout(n20265));
    jdff dff_A_KJykaV3M0_2(.din(n5789), .dout(G469));
    jdff dff_A_u8189vHk1_2(.din(n4691), .dout(G422));
    jdff dff_A_d63CencI3_0(.din(n20253), .dout(G344));
    jdff dff_A_dflpMAFK7_0(.din(n20250), .dout(n20253));
    jdff dff_A_dGxuGP4h3_0(.din(n20247), .dout(n20250));
    jdff dff_A_vN0bMFAx7_0(.din(n20244), .dout(n20247));
    jdff dff_A_r2jAo6Mu9_0(.din(n20241), .dout(n20244));
    jdff dff_A_nRWXLRke4_0(.din(n20238), .dout(n20241));
    jdff dff_A_SpyAcNEH9_0(.din(n20235), .dout(n20238));
    jdff dff_A_XGIEQCg10_0(.din(n20232), .dout(n20235));
    jdff dff_A_hgG319v29_0(.din(n20229), .dout(n20232));
    jdff dff_A_PZYJlCxG8_0(.din(n20226), .dout(n20229));
    jdff dff_A_DVNHGDkx9_0(.din(n20223), .dout(n20226));
    jdff dff_A_AmHEvaNU2_0(.din(n20220), .dout(n20223));
    jdff dff_A_0WEmXAVP9_0(.din(n20217), .dout(n20220));
    jdff dff_A_u2VS0eu85_2(.din(n4666), .dout(n20217));
    jdff dff_A_CLY8YUQh0_0(.din(n20211), .dout(G307));
    jdff dff_A_7tF7lrrX4_0(.din(n20208), .dout(n20211));
    jdff dff_A_gmPvQ6Lp0_0(.din(n20205), .dout(n20208));
    jdff dff_A_4at4GPYc7_0(.din(n20202), .dout(n20205));
    jdff dff_A_F74uv20G6_0(.din(n20199), .dout(n20202));
    jdff dff_A_QW7ti7wh7_0(.din(n20196), .dout(n20199));
    jdff dff_A_idBcVgJA1_0(.din(n20193), .dout(n20196));
    jdff dff_A_GtDw502C2_2(.din(n4662), .dout(n20193));
    jdff dff_A_15EPoaaV9_0(.din(n20187), .dout(G304));
    jdff dff_A_JqoY9hF47_0(.din(n20184), .dout(n20187));
    jdff dff_A_wMRy0g015_0(.din(n20181), .dout(n20184));
    jdff dff_A_nVo2cKWp6_0(.din(n20178), .dout(n20181));
    jdff dff_A_eF8HMsmM0_0(.din(n20175), .dout(n20178));
    jdff dff_A_QNPL4Nn99_2(.din(n4658), .dout(n20175));
    jdff dff_A_FQeftoZR1_0(.din(n20169), .dout(G301));
    jdff dff_A_pq520oT52_0(.din(n20166), .dout(n20169));
    jdff dff_A_wI0jkKM02_0(.din(n20163), .dout(n20166));
    jdff dff_A_2e7Pzvlt4_0(.din(n20160), .dout(n20163));
    jdff dff_A_KvSYlQtB0_0(.din(n20157), .dout(n20160));
    jdff dff_A_kO1eFYA95_2(.din(n4639), .dout(n20157));
    jdff dff_A_3ubhS1Ve3_0(.din(n20151), .dout(G298));
    jdff dff_A_9IN6LYZ30_0(.din(n20148), .dout(n20151));
    jdff dff_A_Yexk4taD4_0(.din(n20145), .dout(n20148));
    jdff dff_A_bXHu9UF51_2(.din(n4632), .dout(n20145));
    jdff dff_A_FoWZznBm6_2(.din(n5785), .dout(G273));
    jdff dff_A_8zlm28G46_0(.din(n20136), .dout(G418));
    jdff dff_A_mmQlEfuy6_0(.din(n20133), .dout(n20136));
    jdff dff_A_JZZMLKg54_0(.din(n20130), .dout(n20133));
    jdff dff_A_DmSxY9v33_0(.din(n20127), .dout(n20130));
    jdff dff_A_n4QvVDPh2_0(.din(n20124), .dout(n20127));
    jdff dff_A_yTIIXXdG2_0(.din(n20121), .dout(n20124));
    jdff dff_A_89CIiKXN0_0(.din(n20118), .dout(n20121));
    jdff dff_A_W32TXfhs9_0(.din(n20115), .dout(n20118));
    jdff dff_A_r7pMVeiv4_0(.din(n20112), .dout(n20115));
    jdff dff_A_IydLM9Go8_0(.din(n20109), .dout(n20112));
    jdff dff_A_DOhhlZFY7_0(.din(n20106), .dout(n20109));
    jdff dff_A_jhWvCLTd0_2(.din(n4606), .dout(n20106));
    jdff dff_A_Faa1tfed9_0(.din(n20100), .dout(G336));
    jdff dff_A_MrFmcRjM9_0(.din(n20097), .dout(n20100));
    jdff dff_A_DmiOXxqU7_0(.din(n20094), .dout(n20097));
    jdff dff_A_bmy2DIyV3_2(.din(n4582), .dout(n20094));
    jdff dff_A_jVNl1AUr1_0(.din(n20088), .dout(G333));
    jdff dff_A_eoKninLD1_0(.din(n20085), .dout(n20088));
    jdff dff_A_YMbsQHww3_0(.din(n20082), .dout(n20085));
    jdff dff_A_56MDtBHq7_2(.din(n4570), .dout(n20082));
    jdff dff_A_UgHHmDTh0_0(.din(n20076), .dout(G330));
    jdff dff_A_WZFDRTZ02_0(.din(n20073), .dout(n20076));
    jdff dff_A_HUfgb5F17_2(.din(n4559), .dout(n20073));
    jdff dff_A_NvrgdMKU2_0(.din(n20067), .dout(G327));
    jdff dff_A_IyoCa8wx8_2(.din(n4548), .dout(n20067));
    jdff dff_A_yZTlQUTQ7_0(.din(n20061), .dout(G319));
    jdff dff_A_h8Q04HCz0_0(.din(n20058), .dout(n20061));
    jdff dff_A_xI4IW2bo6_0(.din(n20055), .dout(n20058));
    jdff dff_A_4AYGEmap7_0(.din(n20052), .dout(n20055));
    jdff dff_A_aVSyyIGQ5_0(.din(n20049), .dout(n20052));
    jdff dff_A_j0C65L6g2_0(.din(n20046), .dout(n20049));
    jdff dff_A_KDAv0QYT0_0(.din(n20043), .dout(n20046));
    jdff dff_A_IhK2kk8i6_2(.din(n4516), .dout(n20043));
    jdff dff_A_7WMxIowz2_0(.din(n20037), .dout(G316));
    jdff dff_A_eKNM7vN50_0(.din(n20034), .dout(n20037));
    jdff dff_A_a5BYp71V9_0(.din(n20031), .dout(n20034));
    jdff dff_A_THjpltkp3_0(.din(n20028), .dout(n20031));
    jdff dff_A_t5Uihtn31_0(.din(n20025), .dout(n20028));
    jdff dff_A_RxdP6a0E7_0(.din(n20022), .dout(n20025));
    jdff dff_A_DwVU4p0z8_0(.din(n20019), .dout(n20022));
    jdff dff_A_iJCHvIYW2_2(.din(n4504), .dout(n20019));
    jdff dff_A_S7sW2fzJ2_0(.din(n20013), .dout(G313));
    jdff dff_A_BkSUfK953_0(.din(n20010), .dout(n20013));
    jdff dff_A_IMsKFPMu0_0(.din(n20007), .dout(n20010));
    jdff dff_A_eGCBi7UI3_0(.din(n20004), .dout(n20007));
    jdff dff_A_ruIjEfsc5_0(.din(n20001), .dout(n20004));
    jdff dff_A_7l6AgJFW3_0(.din(n19998), .dout(n20001));
    jdff dff_A_u94kLzpL1_2(.din(n4486), .dout(n19998));
    jdff dff_A_pHtuYwCX5_0(.din(n19992), .dout(G310));
    jdff dff_A_Bo9l5qom6_0(.din(n19989), .dout(n19992));
    jdff dff_A_uw9UyzKk2_0(.din(n19986), .dout(n19989));
    jdff dff_A_kifR7LAe6_0(.din(n19983), .dout(n19986));
    jdff dff_A_Y4t8sdBm8_0(.din(n19980), .dout(n19983));
    jdff dff_A_ACqslBCv7_2(.din(n4478), .dout(n19980));
    jdff dff_A_kfLFkw6M5_2(.din(n5781), .dout(G276));
    jdff dff_A_NfzkrZUl7_0(.din(n19971), .dout(G252));
    jdff dff_A_Tsmut07i4_0(.din(n19968), .dout(n19971));
    jdff dff_A_jsap1kaJ3_0(.din(n19965), .dout(n19968));
    jdff dff_A_lgpTcbSX8_0(.din(n19962), .dout(n19965));
    jdff dff_A_r0NcR0A47_0(.din(n19959), .dout(n19962));
    jdff dff_A_Uy4DScXa9_0(.din(n19956), .dout(n19959));
    jdff dff_A_V1Y6LPsY3_0(.din(n19953), .dout(n19956));
    jdff dff_A_aYv5HA7j9_0(.din(n19950), .dout(n19953));
    jdff dff_A_xV6enaR67_0(.din(n19947), .dout(n19950));
    jdff dff_A_y1lICjJJ6_2(.din(n4446), .dout(n19947));
    jdff dff_A_6x2DiZCh2_0(.din(n19941), .dout(G324));
    jdff dff_A_rf51OD4G6_0(.din(n19938), .dout(n19941));
    jdff dff_A_Cle7SSIO7_0(.din(n19935), .dout(n19938));
    jdff dff_A_zYoIwaxo4_0(.din(n19932), .dout(n19935));
    jdff dff_A_I97Xg4N51_0(.din(n19929), .dout(n19932));
    jdff dff_A_ouDDPZkR1_2(.din(n4418), .dout(n19929));
    jdff dff_A_ncsEIN7l2_0(.din(n19923), .dout(G295));
    jdff dff_A_6if8DXLV5_0(.din(n19920), .dout(n19923));
    jdff dff_A_r89USscb9_0(.din(n19917), .dout(n19920));
    jdff dff_A_kdjx6fiP2_0(.din(n19914), .dout(n19917));
    jdff dff_A_nvdRjiDF3_0(.din(n19911), .dout(n19914));
    jdff dff_A_e9EVMRV11_0(.din(n19908), .dout(n19911));
    jdff dff_A_EZQyUxsP2_0(.din(n19905), .dout(n19908));
    jdff dff_A_Otjvdvdr9_0(.din(n19902), .dout(n19905));
    jdff dff_A_GI0MnWIo1_0(.din(n19899), .dout(n19902));
    jdff dff_A_k8fwsG6X8_2(.din(n4392), .dout(n19899));
    jdff dff_A_oXOkdpwq9_0(.din(n19893), .dout(G249));
    jdff dff_A_dz6pocrP5_0(.din(n19890), .dout(n19893));
    jdff dff_A_AACjyD1C0_0(.din(n19887), .dout(n19890));
    jdff dff_A_IShvtZLt9_0(.din(n19884), .dout(n19887));
    jdff dff_A_HRHixrIo2_0(.din(n19881), .dout(n19884));
    jdff dff_A_7iyGzNrG8_0(.din(n19878), .dout(n19881));
    jdff dff_A_hMJWlTAb8_2(.din(n5777), .dout(n19878));
    jdff dff_A_IFN6ScqP4_0(.din(n19872), .dout(G416));
    jdff dff_A_JgCU2Fav8_0(.din(n19869), .dout(n19872));
    jdff dff_A_eZsSL7no0_0(.din(n19866), .dout(n19869));
    jdff dff_A_gGKKYrL76_0(.din(n19863), .dout(n19866));
    jdff dff_A_RUF0Bp9h5_0(.din(n19860), .dout(n19863));
    jdff dff_A_xtdju5j15_0(.din(n19857), .dout(n19860));
    jdff dff_A_dtQrnXPr1_0(.din(n19854), .dout(n19857));
    jdff dff_A_BLZDHSPz7_0(.din(n19851), .dout(n19854));
    jdff dff_A_Y6Rgkjl59_0(.din(n19848), .dout(n19851));
    jdff dff_A_ZIlnqiwe7_0(.din(n19845), .dout(n19848));
    jdff dff_A_9HxK52q10_0(.din(n19842), .dout(n19845));
    jdff dff_A_IPLLeTBj4_0(.din(n19839), .dout(n19842));
    jdff dff_A_SlpxzlWo9_0(.din(n19836), .dout(n19839));
    jdff dff_A_5Phao2qY9_1(.din(n4280), .dout(n19836));
    jdff dff_A_cJ8tRCMf1_0(.din(n19830), .dout(G414));
    jdff dff_A_7yOlvR0b9_0(.din(n19827), .dout(n19830));
    jdff dff_A_l36IXXuE2_0(.din(n19824), .dout(n19827));
    jdff dff_A_uu30PPq45_0(.din(n19821), .dout(n19824));
    jdff dff_A_AJCzSzAi8_0(.din(n19818), .dout(n19821));
    jdff dff_A_E0G0wta24_0(.din(n19815), .dout(n19818));
    jdff dff_A_f8kk55bC7_0(.din(n19812), .dout(n19815));
    jdff dff_A_2VFTo9823_0(.din(n19809), .dout(n19812));
    jdff dff_A_8I9NFbmK2_0(.din(n19806), .dout(n19809));
    jdff dff_A_KCQfCrxM3_0(.din(n19803), .dout(n19806));
    jdff dff_A_KZ876fa08_0(.din(n19800), .dout(n19803));
    jdff dff_A_ydPQZw6P4_0(.din(n19797), .dout(n19800));
    jdff dff_A_ZHXGwIji4_0(.din(n19794), .dout(n19797));
    jdff dff_A_trM5DOrX7_0(.din(n19791), .dout(n19794));
    jdff dff_A_pkJ0GkZQ3_0(.din(n19788), .dout(n19791));
    jdff dff_A_nyyEt9jd2_1(.din(n3990), .dout(n19788));
    jdff dff_A_tgV96mPK7_0(.din(n19782), .dout(G412));
    jdff dff_A_12cptL5E3_0(.din(n19779), .dout(n19782));
    jdff dff_A_bCsRiVss5_0(.din(n19776), .dout(n19779));
    jdff dff_A_AYx6ANXW1_0(.din(n19773), .dout(n19776));
    jdff dff_A_zoXH8DyH0_0(.din(n19770), .dout(n19773));
    jdff dff_A_AXYOX6if8_0(.din(n19767), .dout(n19770));
    jdff dff_A_lpC5Yjxz4_0(.din(n19764), .dout(n19767));
    jdff dff_A_W2Pe5qtY8_0(.din(n19761), .dout(n19764));
    jdff dff_A_1EZv6f307_0(.din(n19758), .dout(n19761));
    jdff dff_A_fJtPq6tq7_0(.din(n19755), .dout(n19758));
    jdff dff_A_wwXYz9bQ8_0(.din(n19752), .dout(n19755));
    jdff dff_A_JEMkHivD3_0(.din(n19749), .dout(n19752));
    jdff dff_A_KSSYnzCg4_0(.din(n19746), .dout(n19749));
    jdff dff_A_wc9ihYAb6_0(.din(n19743), .dout(n19746));
    jdff dff_A_9zPqFGQz7_0(.din(n19740), .dout(n19743));
    jdff dff_A_wykqDbm08_1(.din(n3737), .dout(n19740));
    jdff dff_A_Z4ta4T7k2_0(.din(n19734), .dout(G385));
    jdff dff_A_G4xBhRH19_0(.din(n19731), .dout(n19734));
    jdff dff_A_DzVLEwtQ3_0(.din(n19728), .dout(n19731));
    jdff dff_A_La0VcisY5_0(.din(n19725), .dout(n19728));
    jdff dff_A_bwfAXsGr4_0(.din(n19722), .dout(n19725));
    jdff dff_A_kT2xvXs51_0(.din(n19719), .dout(n19722));
    jdff dff_A_MmLIGxEI6_0(.din(n19716), .dout(n19719));
    jdff dff_A_3oRT5DHU4_0(.din(n19713), .dout(n19716));
    jdff dff_A_wfrMokYK3_0(.din(n19710), .dout(n19713));
    jdff dff_A_udbXHxti9_0(.din(n19707), .dout(n19710));
    jdff dff_A_19jiPMKQ0_0(.din(n19704), .dout(n19707));
    jdff dff_A_507IISw87_0(.din(n19701), .dout(n19704));
    jdff dff_A_Do8OgmES8_0(.din(n19698), .dout(n19701));
    jdff dff_A_kn56FF7D5_0(.din(n19695), .dout(n19698));
    jdff dff_A_NxRbqHJi1_0(.din(n19692), .dout(n19695));
    jdff dff_A_H03IRAWS8_2(.din(n3495), .dout(n19692));
    jdff dff_A_zOjJnjDn1_0(.din(n19686), .dout(G382));
    jdff dff_A_MZeBBfbI7_0(.din(n19683), .dout(n19686));
    jdff dff_A_E0shbqX76_0(.din(n19680), .dout(n19683));
    jdff dff_A_BbYuBmPy4_0(.din(n19677), .dout(n19680));
    jdff dff_A_Mzv24KvU8_0(.din(n19674), .dout(n19677));
    jdff dff_A_MRYJka3J2_0(.din(n19671), .dout(n19674));
    jdff dff_A_Rz8PGoUa2_0(.din(n19668), .dout(n19671));
    jdff dff_A_mVqDdQf03_0(.din(n19665), .dout(n19668));
    jdff dff_A_SeZHf1mh4_0(.din(n19662), .dout(n19665));
    jdff dff_A_NdYWOdoP6_0(.din(n19659), .dout(n19662));
    jdff dff_A_ao8l4W4i3_0(.din(n19656), .dout(n19659));
    jdff dff_A_8nnZTuLO6_0(.din(n19653), .dout(n19656));
    jdff dff_A_9WmLhrWF7_0(.din(n19650), .dout(n19653));
    jdff dff_A_f3sHIXSK4_2(.din(n3491), .dout(n19650));
    jdff dff_A_M1p3FErj9_0(.din(n19644), .dout(G379));
    jdff dff_A_SJ3isSEu3_0(.din(n19641), .dout(n19644));
    jdff dff_A_57TMX5lc6_0(.din(n19638), .dout(n19641));
    jdff dff_A_I4jCtoFc9_0(.din(n19635), .dout(n19638));
    jdff dff_A_0Bx1f9IE1_0(.din(n19632), .dout(n19635));
    jdff dff_A_aXzsrJp07_0(.din(n19629), .dout(n19632));
    jdff dff_A_p8pYFDhF7_0(.din(n19626), .dout(n19629));
    jdff dff_A_rdtp5aFN2_0(.din(n19623), .dout(n19626));
    jdff dff_A_1wUGljjO2_0(.din(n19620), .dout(n19623));
    jdff dff_A_vsPVKiou5_0(.din(n19617), .dout(n19620));
    jdff dff_A_OMstosv94_0(.din(n19614), .dout(n19617));
    jdff dff_A_FmiXhclr4_0(.din(n19611), .dout(n19614));
    jdff dff_A_dnP6G8TY7_0(.din(n19608), .dout(n19611));
    jdff dff_A_8VidLIuF6_2(.din(n3475), .dout(n19608));
    jdff dff_A_dUxt6AWx7_0(.din(n19602), .dout(G376));
    jdff dff_A_RuO7mcqB9_0(.din(n19599), .dout(n19602));
    jdff dff_A_MqYYqK3a1_0(.din(n19596), .dout(n19599));
    jdff dff_A_MJlkpX5O9_0(.din(n19593), .dout(n19596));
    jdff dff_A_IOOoSHDD5_0(.din(n19590), .dout(n19593));
    jdff dff_A_hMo2T9ni6_0(.din(n19587), .dout(n19590));
    jdff dff_A_Gd6waxCM1_0(.din(n19584), .dout(n19587));
    jdff dff_A_bv59T8UL8_0(.din(n19581), .dout(n19584));
    jdff dff_A_Qfzya5Ze6_0(.din(n19578), .dout(n19581));
    jdff dff_A_hvDXOGaJ2_0(.din(n19575), .dout(n19578));
    jdff dff_A_dBqpDcpe0_0(.din(n19572), .dout(n19575));
    jdff dff_A_q36PlStj3_0(.din(n19569), .dout(n19572));
    jdff dff_A_KMCbaGeF1_2(.din(n3467), .dout(n19569));
    jdff dff_A_2FJp0xsN4_0(.din(n19563), .dout(G397));
    jdff dff_A_STpoYxwp4_0(.din(n19560), .dout(n19563));
    jdff dff_A_paqg3lvO4_0(.din(n19557), .dout(n19560));
    jdff dff_A_nYIGNC6q8_0(.din(n19554), .dout(n19557));
    jdff dff_A_4J9jGk8k2_0(.din(n19551), .dout(n19554));
    jdff dff_A_wXGwjV8M1_0(.din(n19548), .dout(n19551));
    jdff dff_A_yg8BF1l82_0(.din(n19545), .dout(n19548));
    jdff dff_A_xfZCYeKO1_0(.din(n19542), .dout(n19545));
    jdff dff_A_3WbuAF9l4_0(.din(n19539), .dout(n19542));
    jdff dff_A_OSTDsA4W7_0(.din(n19536), .dout(n19539));
    jdff dff_A_z1gzQNb06_0(.din(n19533), .dout(n19536));
    jdff dff_A_GNuP6mjp8_0(.din(n19530), .dout(n19533));
    jdff dff_A_D8skds636_0(.din(n19527), .dout(n19530));
    jdff dff_A_VYie8oKZ4_0(.din(n19524), .dout(n19527));
    jdff dff_A_ZUoOI0BO5_0(.din(n19521), .dout(n19524));
    jdff dff_A_iLpUerIY1_0(.din(n19518), .dout(n19521));
    jdff dff_A_FMvSAZ0R2_0(.din(n19515), .dout(n19518));
    jdff dff_A_vmdaJfph6_0(.din(n19512), .dout(n19515));
    jdff dff_A_vEddeJa75_2(.din(n3451), .dout(n19512));
    jdff dff_A_fqNnckpX0_0(.din(n19506), .dout(G394));
    jdff dff_A_bA3xXtm41_0(.din(n19503), .dout(n19506));
    jdff dff_A_rGQ9rEbx1_0(.din(n19500), .dout(n19503));
    jdff dff_A_b4esieFH2_0(.din(n19497), .dout(n19500));
    jdff dff_A_OvuI36Xm3_0(.din(n19494), .dout(n19497));
    jdff dff_A_r8yX35OL0_0(.din(n19491), .dout(n19494));
    jdff dff_A_Ly7xUSq95_0(.din(n19488), .dout(n19491));
    jdff dff_A_wSkeehsm1_0(.din(n19485), .dout(n19488));
    jdff dff_A_pUlb9P5P1_0(.din(n19482), .dout(n19485));
    jdff dff_A_OcCMQ68y4_0(.din(n19479), .dout(n19482));
    jdff dff_A_JFg8rEiJ6_0(.din(n19476), .dout(n19479));
    jdff dff_A_6pg4YxwW2_0(.din(n19473), .dout(n19476));
    jdff dff_A_Bqrd55ic6_0(.din(n19470), .dout(n19473));
    jdff dff_A_fEJYJaC64_0(.din(n19467), .dout(n19470));
    jdff dff_A_nc2zuewP2_0(.din(n19464), .dout(n19467));
    jdff dff_A_JvoLXZv29_0(.din(n19461), .dout(n19464));
    jdff dff_A_bGy4FE5o1_0(.din(n19458), .dout(n19461));
    jdff dff_A_wd3queQl0_2(.din(n3439), .dout(n19458));
    jdff dff_A_xb28ihKw9_0(.din(n19452), .dout(G391));
    jdff dff_A_ahq94RXh2_0(.din(n19449), .dout(n19452));
    jdff dff_A_hMRbFHPt0_0(.din(n19446), .dout(n19449));
    jdff dff_A_bUZ8UM2f2_0(.din(n19443), .dout(n19446));
    jdff dff_A_mRydFenQ2_0(.din(n19440), .dout(n19443));
    jdff dff_A_B1GN1IsM6_0(.din(n19437), .dout(n19440));
    jdff dff_A_5OJnOWhJ3_0(.din(n19434), .dout(n19437));
    jdff dff_A_RUKf3Paw2_0(.din(n19431), .dout(n19434));
    jdff dff_A_5Dx3uy0W1_0(.din(n19428), .dout(n19431));
    jdff dff_A_fOBBr3vE7_0(.din(n19425), .dout(n19428));
    jdff dff_A_L7xEiLZH9_0(.din(n19422), .dout(n19425));
    jdff dff_A_h9k8PZIV0_0(.din(n19419), .dout(n19422));
    jdff dff_A_nwtmSoKe8_0(.din(n19416), .dout(n19419));
    jdff dff_A_jJkwxnye2_0(.din(n19413), .dout(n19416));
    jdff dff_A_evzt3vR01_0(.din(n19410), .dout(n19413));
    jdff dff_A_YjJZ0vk19_0(.din(n19407), .dout(n19410));
    jdff dff_A_f4MjxiJZ3_2(.din(n3427), .dout(n19407));
    jdff dff_A_iTOYy22w6_0(.din(n19401), .dout(G388));
    jdff dff_A_Uw3YYzYS7_0(.din(n19398), .dout(n19401));
    jdff dff_A_XE6rjJ8Q7_0(.din(n19395), .dout(n19398));
    jdff dff_A_PBnnuB6u7_0(.din(n19392), .dout(n19395));
    jdff dff_A_REsitmqL9_0(.din(n19389), .dout(n19392));
    jdff dff_A_AXXGvaV37_0(.din(n19386), .dout(n19389));
    jdff dff_A_lfTIEuZs4_0(.din(n19383), .dout(n19386));
    jdff dff_A_RL0IalGz4_0(.din(n19380), .dout(n19383));
    jdff dff_A_RgXVgALg9_0(.din(n19377), .dout(n19380));
    jdff dff_A_CRC1ax6O2_0(.din(n19374), .dout(n19377));
    jdff dff_A_DstrArim9_0(.din(n19371), .dout(n19374));
    jdff dff_A_LfJ9L3gi7_0(.din(n19368), .dout(n19371));
    jdff dff_A_cYIudUaM3_0(.din(n19365), .dout(n19368));
    jdff dff_A_kyTaRLFF9_0(.din(n19362), .dout(n19365));
    jdff dff_A_l9LCgxGv9_2(.din(n3419), .dout(n19362));
    jdff dff_A_nl5Rctji5_2(.din(n5773), .dout(G270));
    jdff dff_A_k292zF0g9_0(.din(n19353), .dout(G264));
    jdff dff_A_0qrM3nOe3_0(.din(n19350), .dout(n19353));
    jdff dff_A_B7VaiMwO9_0(.din(n19347), .dout(n19350));
    jdff dff_A_XCW9JrQp7_0(.din(n19344), .dout(n19347));
    jdff dff_A_WaQ6FwW05_0(.din(n19341), .dout(n19344));
    jdff dff_A_NfaO50cd0_0(.din(n19338), .dout(n19341));
    jdff dff_A_A5XS2GlF0_2(.din(n5769), .dout(n19338));
    jdff dff_A_VxpAgs9w9_0(.din(n19332), .dout(G258));
    jdff dff_A_xBLn3BnK2_0(.din(n19329), .dout(n19332));
    jdff dff_A_hqOvNHIe1_0(.din(n19326), .dout(n19329));
    jdff dff_A_mlraThnj5_0(.din(n19323), .dout(n19326));
    jdff dff_A_sC8XpTxb0_0(.din(n19320), .dout(n19323));
    jdff dff_A_EolVQK7x9_0(.din(n19317), .dout(n19320));
    jdff dff_A_Q0JJXQ6q2_2(.din(n3391), .dout(n19317));
    jdff dff_A_R2YdaLCt7_2(.din(n1828), .dout(G246));
    jdff dff_A_Vdzrohec1_0(.din(n19308), .dout(G373));
    jdff dff_A_wt6Hobxm6_0(.din(n19305), .dout(n19308));
    jdff dff_A_AOegXKqA3_0(.din(n19302), .dout(n19305));
    jdff dff_A_aOg81CMv9_0(.din(n19299), .dout(n19302));
    jdff dff_A_tUg9irBn6_0(.din(n19296), .dout(n19299));
    jdff dff_A_IZKCF9bv4_0(.din(n19293), .dout(n19296));
    jdff dff_A_J9CsCj704_0(.din(n19290), .dout(n19293));
    jdff dff_A_duZ6ox7B9_0(.din(n19287), .dout(n19290));
    jdff dff_A_2K8I8pYJ2_0(.din(n19284), .dout(n19287));
    jdff dff_A_rDQulIv00_0(.din(n19281), .dout(n19284));
    jdff dff_A_7lvWxaUV1_0(.din(n19278), .dout(n19281));
    jdff dff_A_ffppzAl97_0(.din(n19275), .dout(n19278));
    jdff dff_A_0FfUMgF40_0(.din(n19272), .dout(n19275));
    jdff dff_A_cRyE3iZd2_0(.din(n19269), .dout(n19272));
    jdff dff_A_UkK3hfsn5_0(.din(n19266), .dout(n19269));
    jdff dff_A_RViSHWIa6_0(.din(n19263), .dout(n19266));
    jdff dff_A_k30oTUpH7_0(.din(n19260), .dout(n19263));
    jdff dff_A_AW4dAvYN2_0(.din(n19257), .dout(n19260));
    jdff dff_A_VHezfZ6H0_0(.din(n19254), .dout(n19257));
    jdff dff_A_7g34HPfj9_0(.din(n19251), .dout(n19254));
    jdff dff_A_CGluyyLx8_2(.din(n486), .dout(n19251));
    jdff dff_A_616RzkKH1_0(.din(n19245), .dout(G278));
    jdff dff_A_FTt1kzgv0_0(.din(n19242), .dout(n19245));
    jdff dff_A_g3TADX9Q0_0(.din(n19239), .dout(n19242));
    jdff dff_A_aRdiGPis4_0(.din(n19236), .dout(n19239));
    jdff dff_A_1KH2B4jk1_0(.din(n19233), .dout(n19236));
    jdff dff_A_6uv0cKzz0_0(.din(n19230), .dout(n19233));
    jdff dff_A_FvC1yZEg1_0(.din(n19227), .dout(n19230));
    jdff dff_A_Kk3CIjBV7_0(.din(n19224), .dout(n19227));
    jdff dff_A_juM6jieX6_0(.din(n19221), .dout(n19224));
    jdff dff_A_hIO7XOSO3_0(.din(n19218), .dout(n19221));
    jdff dff_A_u37X9amP7_0(.din(n19215), .dout(n19218));
    jdff dff_A_NsMAW75Q4_0(.din(n19212), .dout(n19215));
    jdff dff_A_4lu8Ud9g5_0(.din(n19209), .dout(n19212));
    jdff dff_A_rFhaQCry4_0(.din(n19206), .dout(n19209));
    jdff dff_A_EKIfQgUg4_0(.din(n19203), .dout(n19206));
    jdff dff_A_uB2ThT4B7_0(.din(n19200), .dout(n19203));
    jdff dff_A_Vywao6KF8_0(.din(n19197), .dout(n19200));
    jdff dff_A_lpZiuo7Q5_0(.din(n19194), .dout(n19197));
    jdff dff_A_9HW4GkQG2_0(.din(n19191), .dout(n19194));
    jdff dff_A_g855YBmC2_0(.din(n19188), .dout(n19191));
    jdff dff_A_l4jzBRgz9_0(.din(n19185), .dout(n19188));
    jdff dff_A_qnwoH1QE8_0(.din(n19182), .dout(n19185));
    jdff dff_A_12W7fw4g4_0(.din(n19179), .dout(n19182));
    jdff dff_A_5GKxlkRZ6_0(.din(n19176), .dout(n19179));
    jdff dff_A_Ed2rPu1D0_0(.din(n19173), .dout(n19176));
    jdff dff_A_NHAxy8Qq4_2(.din(n441), .dout(n19173));
    jdff dff_A_ZsdjeHLx7_0(.din(n19167), .dout(G453));
    jdff dff_A_LnjKUAvC2_0(.din(n19164), .dout(n19167));
    jdff dff_A_8JYjHguq9_0(.din(n19161), .dout(n19164));
    jdff dff_A_jI5PA4cr5_0(.din(n19158), .dout(n19161));
    jdff dff_A_nJBLzrFr4_0(.din(n19155), .dout(n19158));
    jdff dff_A_6YDxurMj0_0(.din(n19152), .dout(n19155));
    jdff dff_A_rw9JupFW6_0(.din(n19149), .dout(n19152));
    jdff dff_A_kMdQl0sT9_0(.din(n19146), .dout(n19149));
    jdff dff_A_828TThmF2_0(.din(n19143), .dout(n19146));
    jdff dff_A_Pr7Qdmus9_0(.din(n19140), .dout(n19143));
    jdff dff_A_sCvFeNMs8_0(.din(n19137), .dout(n19140));
    jdff dff_A_Ggj6PLQA7_0(.din(n19134), .dout(n19137));
    jdff dff_A_4AJOowQ61_0(.din(n19131), .dout(n19134));
    jdff dff_A_l2yFXSXP9_0(.din(n19128), .dout(n19131));
    jdff dff_A_cWKhQbOq7_0(.din(n19125), .dout(n19128));
    jdff dff_A_jGsiy5Vs4_0(.din(n19122), .dout(n19125));
    jdff dff_A_mJaz4RL47_0(.din(n19119), .dout(n19122));
    jdff dff_A_tmjihczE0_0(.din(n19116), .dout(n19119));
    jdff dff_A_IFbVjk4p0_0(.din(n19113), .dout(n19116));
    jdff dff_A_NtXSZeMD2_0(.din(n19110), .dout(n19113));
    jdff dff_A_8ZxcYVqP1_0(.din(n19107), .dout(n19110));
    jdff dff_A_CtB9QTOK3_0(.din(n19104), .dout(n19107));
    jdff dff_A_azWxccFr5_0(.din(n19101), .dout(n19104));
    jdff dff_A_Gjvg1V2t4_0(.din(n19098), .dout(n19101));
    jdff dff_A_tZyf03n89_0(.din(n19095), .dout(n19098));
    jdff dff_A_WfeN12RN7_1(.din(n5765), .dout(n19095));
    jdff dff_A_iq9tyi289_0(.din(n19089), .dout(G281));
    jdff dff_A_JU682vyY6_0(.din(n19086), .dout(n19089));
    jdff dff_A_ERkJuYSS5_0(.din(n19083), .dout(n19086));
    jdff dff_A_cuKXS15k1_0(.din(n19080), .dout(n19083));
    jdff dff_A_vLeYnClR3_0(.din(n19077), .dout(n19080));
    jdff dff_A_ItvX0lT74_0(.din(n19074), .dout(n19077));
    jdff dff_A_LtRtOvmL0_0(.din(n19071), .dout(n19074));
    jdff dff_A_t8W8UlgB0_0(.din(n19068), .dout(n19071));
    jdff dff_A_WuzeQQ1s7_0(.din(n19065), .dout(n19068));
    jdff dff_A_Vf3PdFCW9_0(.din(n19062), .dout(n19065));
    jdff dff_A_euzOGjlo0_0(.din(n19059), .dout(n19062));
    jdff dff_A_1CjAG2pP2_0(.din(n19056), .dout(n19059));
    jdff dff_A_TGP3O5wA8_0(.din(n19053), .dout(n19056));
    jdff dff_A_aZe4e1ew5_0(.din(n19050), .dout(n19053));
    jdff dff_A_CDgFEVpt9_0(.din(n19047), .dout(n19050));
    jdff dff_A_qdpVz5IX4_0(.din(n19044), .dout(n19047));
    jdff dff_A_mfh1uOZu7_0(.din(n19041), .dout(n19044));
    jdff dff_A_JnR1XVpz2_0(.din(n19038), .dout(n19041));
    jdff dff_A_dd5Lt2ZD9_0(.din(n19035), .dout(n19038));
    jdff dff_A_JBkwmDO49_0(.din(n19032), .dout(n19035));
    jdff dff_A_CCfZjVuf9_0(.din(n19029), .dout(n19032));
    jdff dff_A_OgrGov5P8_0(.din(n19026), .dout(n19029));
    jdff dff_A_mVZ1O6Hg3_0(.din(n19023), .dout(n19026));
    jdff dff_A_KrEOdKkt7_2(.din(n5762), .dout(n19023));
    jdff dff_A_ypRPQATu8_0(.din(n19017), .dout(G341));
    jdff dff_A_TUnYOaP23_0(.din(n19014), .dout(n19017));
    jdff dff_A_jJFIApff5_0(.din(n19011), .dout(n19014));
    jdff dff_A_CHKqgrw39_0(.din(n19008), .dout(n19011));
    jdff dff_A_Rau2rxJ47_0(.din(n19005), .dout(n19008));
    jdff dff_A_IJyfc8eZ7_0(.din(n19002), .dout(n19005));
    jdff dff_A_PDcYMmLt2_0(.din(n18999), .dout(n19002));
    jdff dff_A_Px8UShAx9_0(.din(n18996), .dout(n18999));
    jdff dff_A_qKiuXRsu4_0(.din(n18993), .dout(n18996));
    jdff dff_A_bnM2uTsC1_0(.din(n18990), .dout(n18993));
    jdff dff_A_VFB3a0un3_0(.din(n18987), .dout(n18990));
    jdff dff_A_I6Pd9k5c6_0(.din(n18984), .dout(n18987));
    jdff dff_A_7bf8dao58_0(.din(n18981), .dout(n18984));
    jdff dff_A_oNmloiZZ7_0(.din(n18978), .dout(n18981));
    jdff dff_A_mwV8252j8_0(.din(n18975), .dout(n18978));
    jdff dff_A_re6X1cVW3_0(.din(n18972), .dout(n18975));
    jdff dff_A_Z2Wsc5eu7_0(.din(n18969), .dout(n18972));
    jdff dff_A_frIeChTW7_0(.din(n18966), .dout(n18969));
    jdff dff_A_x2gAadT62_0(.din(n18963), .dout(n18966));
    jdff dff_A_vL7Wn4443_0(.din(n18960), .dout(n18963));
    jdff dff_A_Z58CL2R31_0(.din(n18957), .dout(n18960));
    jdff dff_A_KQ3zL1Bu0_0(.din(n18954), .dout(n18957));
    jdff dff_A_RowHP7Ov6_0(.din(n18951), .dout(n18954));
    jdff dff_A_RGEZTkao7_0(.din(n18948), .dout(n18951));
    jdff dff_A_ZmDIu1cI5_0(.din(n18945), .dout(n18948));
    jdff dff_A_w5MdrG526_1(.din(n5758), .dout(n18945));
    jdff dff_A_sSTDtCZF9_0(.din(n18939), .dout(G292));
    jdff dff_A_tVeKdouP0_0(.din(n18936), .dout(n18939));
    jdff dff_A_4UzhitIC0_0(.din(n18933), .dout(n18936));
    jdff dff_A_mTDUt9HN2_0(.din(n18930), .dout(n18933));
    jdff dff_A_WB6mi2477_0(.din(n18927), .dout(n18930));
    jdff dff_A_uKEtiqzL7_0(.din(n18924), .dout(n18927));
    jdff dff_A_BQ2wGKp42_0(.din(n18921), .dout(n18924));
    jdff dff_A_eCEWwOLG8_0(.din(n18918), .dout(n18921));
    jdff dff_A_3NTHNzxg5_0(.din(n18915), .dout(n18918));
    jdff dff_A_Xr7dG80L3_0(.din(n18912), .dout(n18915));
    jdff dff_A_yq4ktUSW8_0(.din(n18909), .dout(n18912));
    jdff dff_A_WltOxQ4d6_0(.din(n18906), .dout(n18909));
    jdff dff_A_uYEAjJdY3_0(.din(n18903), .dout(n18906));
    jdff dff_A_jbFWPGkK0_0(.din(n18900), .dout(n18903));
    jdff dff_A_atxPUGMS8_0(.din(n18897), .dout(n18900));
    jdff dff_A_DzcVN8oE2_0(.din(n18894), .dout(n18897));
    jdff dff_A_3Q53PGQx6_0(.din(n18891), .dout(n18894));
    jdff dff_A_jYew3Hxd8_0(.din(n18888), .dout(n18891));
    jdff dff_A_0IYeoJO08_0(.din(n18885), .dout(n18888));
    jdff dff_A_HwwT2VBs3_0(.din(n18882), .dout(n18885));
    jdff dff_A_kWDoJ2f79_0(.din(n18879), .dout(n18882));
    jdff dff_A_6uYZIZJe3_0(.din(n18876), .dout(n18879));
    jdff dff_A_XZJSgp7Q0_0(.din(n18873), .dout(n18876));
    jdff dff_A_Ti7Z5XKL2_2(.din(n437), .dout(n18873));
    jdff dff_A_jzj3M23R2_0(.din(n18867), .dout(G289));
    jdff dff_A_r6dNMP9X2_0(.din(n18864), .dout(n18867));
    jdff dff_A_mpA9ibvw3_0(.din(n18861), .dout(n18864));
    jdff dff_A_nPVIIYij4_0(.din(n18858), .dout(n18861));
    jdff dff_A_MQJAntPL9_0(.din(n18855), .dout(n18858));
    jdff dff_A_RVwgB2Tj4_0(.din(n18852), .dout(n18855));
    jdff dff_A_K8MY7GbE9_0(.din(n18849), .dout(n18852));
    jdff dff_A_qO8Kzqhg2_0(.din(n18846), .dout(n18849));
    jdff dff_A_EoD8049A5_0(.din(n18843), .dout(n18846));
    jdff dff_A_PFBddvsS8_0(.din(n18840), .dout(n18843));
    jdff dff_A_ffF48l0z7_0(.din(n18837), .dout(n18840));
    jdff dff_A_jtelvk5G4_0(.din(n18834), .dout(n18837));
    jdff dff_A_uvS5cts93_0(.din(n18831), .dout(n18834));
    jdff dff_A_7i0u7VnG0_0(.din(n18828), .dout(n18831));
    jdff dff_A_B5xA7uuC2_0(.din(n18825), .dout(n18828));
    jdff dff_A_td3SoSxZ4_0(.din(n18822), .dout(n18825));
    jdff dff_A_tqr91HKx9_0(.din(n18819), .dout(n18822));
    jdff dff_A_RiaeiVOj0_0(.din(n18816), .dout(n18819));
    jdff dff_A_9U4sHRSA4_0(.din(n18813), .dout(n18816));
    jdff dff_A_Ys4vWhET0_0(.din(n18810), .dout(n18813));
    jdff dff_A_BjoHQKXg5_0(.din(n18807), .dout(n18810));
    jdff dff_A_SRZrteZt4_0(.din(n18804), .dout(n18807));
    jdff dff_A_Ob68xE3g0_0(.din(n18801), .dout(n18804));
    jdff dff_A_FjlWCj2b4_0(.din(n18798), .dout(n18801));
    jdff dff_A_B1dnqkxZ4_2(.din(n5755), .dout(n18798));
    jdff dff_A_bJdDKUnI4_0(.din(n18792), .dout(G286));
    jdff dff_A_JqeIkt3S9_0(.din(n18789), .dout(n18792));
    jdff dff_A_9t4FJwtc1_0(.din(n18786), .dout(n18789));
    jdff dff_A_vmednM2Z1_0(.din(n18783), .dout(n18786));
    jdff dff_A_AMOmrFv77_0(.din(n18780), .dout(n18783));
    jdff dff_A_YX9ndtTA1_0(.din(n18777), .dout(n18780));
    jdff dff_A_jUh98gZM4_0(.din(n18774), .dout(n18777));
    jdff dff_A_QIAjReQU7_0(.din(n18771), .dout(n18774));
    jdff dff_A_gruBKQpP1_0(.din(n18768), .dout(n18771));
    jdff dff_A_SAgrBDqA8_0(.din(n18765), .dout(n18768));
    jdff dff_A_IVfxt1M71_0(.din(n18762), .dout(n18765));
    jdff dff_A_3tbOnTc90_0(.din(n18759), .dout(n18762));
    jdff dff_A_1Vhkare43_0(.din(n18756), .dout(n18759));
    jdff dff_A_fXXipKZO0_0(.din(n18753), .dout(n18756));
    jdff dff_A_pywCpTOG2_0(.din(n18750), .dout(n18753));
    jdff dff_A_s43xw4uT1_0(.din(n18747), .dout(n18750));
    jdff dff_A_H3DCpLJK0_0(.din(n18744), .dout(n18747));
    jdff dff_A_s9tWOigg2_0(.din(n18741), .dout(n18744));
    jdff dff_A_22z3wZQn7_0(.din(n18738), .dout(n18741));
    jdff dff_A_Dzv8NsPq9_0(.din(n18735), .dout(n18738));
    jdff dff_A_mVvi4glR3_0(.din(n18732), .dout(n18735));
    jdff dff_A_2Nla7SxG5_0(.din(n18729), .dout(n18732));
    jdff dff_A_hPzLgahQ0_0(.din(n18726), .dout(n18729));
    jdff dff_A_bbtb0N6U5_0(.din(n18723), .dout(n18726));
    jdff dff_A_ivQxTsSS9_0(.din(n18720), .dout(n18723));
    jdff dff_A_X70tw3Lb1_1(.din(n5751), .dout(n18720));
    jdff dff_A_X9VjWtUB8_0(.din(n18714), .dout(G284));
    jdff dff_A_N445o3Rm9_0(.din(n18711), .dout(n18714));
    jdff dff_A_8ky1ZFCm5_0(.din(n18708), .dout(n18711));
    jdff dff_A_HEctrAiX7_0(.din(n18705), .dout(n18708));
    jdff dff_A_JZoykD9o0_0(.din(n18702), .dout(n18705));
    jdff dff_A_jQaCBwwH6_0(.din(n18699), .dout(n18702));
    jdff dff_A_wtQeivoA9_0(.din(n18696), .dout(n18699));
    jdff dff_A_bt8591e34_0(.din(n18693), .dout(n18696));
    jdff dff_A_B6PFfiDO5_0(.din(n18690), .dout(n18693));
    jdff dff_A_ehqFbnaG5_0(.din(n18687), .dout(n18690));
    jdff dff_A_JaYtXLZq9_0(.din(n18684), .dout(n18687));
    jdff dff_A_ZDQDla7X1_0(.din(n18681), .dout(n18684));
    jdff dff_A_xcBzd2uN8_0(.din(n18678), .dout(n18681));
    jdff dff_A_nZpA95Uc8_0(.din(n18675), .dout(n18678));
    jdff dff_A_gMYI0Bi43_0(.din(n18672), .dout(n18675));
    jdff dff_A_4GXBB69u9_0(.din(n18669), .dout(n18672));
    jdff dff_A_BkYoCBqS3_0(.din(n18666), .dout(n18669));
    jdff dff_A_08gqP7Sd4_0(.din(n18663), .dout(n18666));
    jdff dff_A_gg64z5bj4_0(.din(n18660), .dout(n18663));
    jdff dff_A_l6Mr2j9G6_0(.din(n18657), .dout(n18660));
    jdff dff_A_c9WI7ptW7_0(.din(n18654), .dout(n18657));
    jdff dff_A_2KxLRPgB1_0(.din(n18651), .dout(n18654));
    jdff dff_A_pwJQ3Uk11_0(.din(n18648), .dout(n18651));
    jdff dff_A_5wY67q0c8_0(.din(n18645), .dout(n18648));
    jdff dff_A_g7IbVewx2_2(.din(n423), .dout(n18645));
    jdff dff_A_nbWEwK1h1_0(.din(n18639), .dout(G446));
    jdff dff_A_BiNXUr146_0(.din(n18636), .dout(n18639));
    jdff dff_A_zWXHBiP27_0(.din(n18633), .dout(n18636));
    jdff dff_A_KqK4n9an8_0(.din(n18630), .dout(n18633));
    jdff dff_A_rR1PNAVS2_0(.din(n18627), .dout(n18630));
    jdff dff_A_Xovkznt48_0(.din(n18624), .dout(n18627));
    jdff dff_A_pDkLOFAW9_0(.din(n18621), .dout(n18624));
    jdff dff_A_2h5znEYC7_0(.din(n18618), .dout(n18621));
    jdff dff_A_INP3Vl365_0(.din(n18615), .dout(n18618));
    jdff dff_A_C3Wea6Qn8_0(.din(n18612), .dout(n18615));
    jdff dff_A_lackjnTj4_0(.din(n18609), .dout(n18612));
    jdff dff_A_uqtJAVxu4_0(.din(n18606), .dout(n18609));
    jdff dff_A_0lDEJ6Vf9_0(.din(n18603), .dout(n18606));
    jdff dff_A_InB5Ribs0_0(.din(n18600), .dout(n18603));
    jdff dff_A_zYfAKsO99_0(.din(n18597), .dout(n18600));
    jdff dff_A_sR8KRVtc9_0(.din(n18594), .dout(n18597));
    jdff dff_A_jVbVynpX2_0(.din(n18591), .dout(n18594));
    jdff dff_A_tF0P8ENf7_0(.din(n18588), .dout(n18591));
    jdff dff_A_yB4gbMmo9_0(.din(n18585), .dout(n18588));
    jdff dff_A_mPT6bhaT9_0(.din(n18582), .dout(n18585));
    jdff dff_A_D2MU0aDz7_0(.din(n18579), .dout(n18582));
    jdff dff_A_BLjghiPx3_0(.din(n18576), .dout(n18579));
    jdff dff_A_FzC9c08i2_0(.din(n18573), .dout(n18576));
    jdff dff_A_Yzq3GCri5_0(.din(n18570), .dout(n18573));
    jdff dff_A_Yf6Mekoh8_0(.din(n18567), .dout(n18570));
    jdff dff_A_VcYMcl4d4_1(.din(n5748), .dout(n18567));
    jdff dff_A_OvPuv0aa0_0(.din(n18561), .dout(G432));
    jdff dff_A_bLpXWvvb6_0(.din(n18558), .dout(n18561));
    jdff dff_A_bFsmNfY29_0(.din(n18555), .dout(n18558));
    jdff dff_A_PoAmZBwf0_0(.din(n18552), .dout(n18555));
    jdff dff_A_7F4X4YAc1_0(.din(n18549), .dout(n18552));
    jdff dff_A_YO1pMBP66_0(.din(n18546), .dout(n18549));
    jdff dff_A_pPf9xNxG2_0(.din(n18543), .dout(n18546));
    jdff dff_A_bZDnzNKi7_0(.din(n18540), .dout(n18543));
    jdff dff_A_s7dAlhV41_0(.din(n18537), .dout(n18540));
    jdff dff_A_M9RJhOXS1_0(.din(n18534), .dout(n18537));
    jdff dff_A_rqv531aD1_0(.din(n18531), .dout(n18534));
    jdff dff_A_1fxqwxrk0_0(.din(n18528), .dout(n18531));
    jdff dff_A_F14rt1un7_0(.din(n18525), .dout(n18528));
    jdff dff_A_zvFqjdZP1_0(.din(n18522), .dout(n18525));
    jdff dff_A_H1x1fNcX7_0(.din(n8217), .dout(n8214));
    jdff dff_A_LJ5eExnU7_0(.din(G5), .dout(n8217));
    jdff dff_A_2Rxoc2Fc8_1(.din(G5), .dout(n8220));
    jdff dff_A_DJsdh6RM2_1(.din(n8226), .dout(n8223));
    jdff dff_A_Csyy1rkH6_1(.din(G5), .dout(n8226));
    jdff dff_A_FaHfh2fO1_2(.din(G5), .dout(n8229));
    jdff dff_B_aOYLngUM6_0(.din(n3411), .dout(n8233));
    jdff dff_B_8GT5GJoe7_3(.din(n3387), .dout(n8236));
    jdff dff_B_Fh6oaYhI2_3(.din(n8236), .dout(n8239));
    jdff dff_B_PdMoONtd1_3(.din(n8239), .dout(n8242));
    jdff dff_B_p4BRydNP0_3(.din(n8242), .dout(n8245));
    jdff dff_B_ZthGTssf3_3(.din(n8245), .dout(n8248));
    jdff dff_B_o9rZ0ppE2_3(.din(n8248), .dout(n8251));
    jdff dff_B_uBKdNDcH8_3(.din(n8251), .dout(n8254));
    jdff dff_B_Obt8tKE48_3(.din(n8254), .dout(n8257));
    jdff dff_B_1hfgjHjp7_3(.din(n8257), .dout(n8260));
    jdff dff_B_pSXeCuZx2_3(.din(n8260), .dout(n8263));
    jdff dff_B_SkkVDdcH5_3(.din(n8263), .dout(n8266));
    jdff dff_B_oos6ncU33_3(.din(n8266), .dout(n8269));
    jdff dff_B_aX6FGgSH8_3(.din(n8269), .dout(n8272));
    jdff dff_B_2zK51HxV0_3(.din(n8272), .dout(n8275));
    jdff dff_B_dPUIaYT13_3(.din(n8275), .dout(n8278));
    jdff dff_B_4GVNBzqu1_3(.din(n8278), .dout(n8281));
    jdff dff_B_nmwzeh3H7_1(.din(n3379), .dout(n8284));
    jdff dff_B_zluYwsbb9_0(.din(n3371), .dout(n8287));
    jdff dff_B_kmsBd3pO9_0(.din(n8287), .dout(n8290));
    jdff dff_B_LJchpJ413_0(.din(n8290), .dout(n8293));
    jdff dff_B_ZknSM7Q69_0(.din(n8293), .dout(n8296));
    jdff dff_B_tPUdWo8h1_0(.din(n8296), .dout(n8299));
    jdff dff_B_Jg7oXZfN3_0(.din(n8299), .dout(n8302));
    jdff dff_B_O9PQ5rko9_0(.din(n8302), .dout(n8305));
    jdff dff_B_IKeI7tOk1_0(.din(n8305), .dout(n8308));
    jdff dff_B_eaos86KW9_0(.din(n8308), .dout(n8311));
    jdff dff_B_CmYdmzaQ9_0(.din(n3367), .dout(n8314));
    jdff dff_B_RqVXRd1E5_0(.din(n8314), .dout(n8317));
    jdff dff_B_PlJ4JVtI2_0(.din(n8317), .dout(n8320));
    jdff dff_B_xZjP3xbI8_0(.din(n3363), .dout(n8323));
    jdff dff_B_rgTnpi6f8_0(.din(n3328), .dout(n8326));
    jdff dff_B_5b8wHGdI0_0(.din(n8326), .dout(n8329));
    jdff dff_B_cx1mKahK3_0(.din(n8329), .dout(n8332));
    jdff dff_B_sOzLRDlF8_0(.din(n8332), .dout(n8335));
    jdff dff_B_RPVfbBDI2_0(.din(n8335), .dout(n8338));
    jdff dff_B_lbPZEWeQ2_0(.din(n8338), .dout(n8341));
    jdff dff_B_YzKhEAQz8_0(.din(n8341), .dout(n8344));
    jdff dff_B_sybW8anM3_0(.din(n8344), .dout(n8347));
    jdff dff_B_LoxfYKrX8_1(.din(n3248), .dout(n8350));
    jdff dff_B_Taz8ROiW9_1(.din(n8350), .dout(n8353));
    jdff dff_B_ucUW0KpF7_1(.din(n3263), .dout(n8356));
    jdff dff_A_dNJIceBS3_1(.din(n3305), .dout(n8358));
    jdff dff_A_W8W1Fbec0_0(.din(n3298), .dout(n8361));
    jdff dff_A_JEJp4n9Z2_0(.din(n8367), .dout(n8364));
    jdff dff_A_wZ1bMUCk5_0(.din(n3194), .dout(n8367));
    jdff dff_B_clBketc26_0(.din(n3132), .dout(n8371));
    jdff dff_B_owubJqtn6_0(.din(n8371), .dout(n8374));
    jdff dff_B_uGdKD9RF0_0(.din(n3128), .dout(n8377));
    jdff dff_B_3YcnjEPM0_0(.din(n8377), .dout(n8380));
    jdff dff_B_Ke6pguCj6_0(.din(n8380), .dout(n8383));
    jdff dff_B_Qusatsm47_0(.din(n8383), .dout(n8386));
    jdff dff_B_xLARylk14_0(.din(n3124), .dout(n8389));
    jdff dff_B_Y78YgRbs9_0(.din(n3096), .dout(n8392));
    jdff dff_B_Szp1HVeJ0_0(.din(n8392), .dout(n8395));
    jdff dff_B_yrJTjGSX8_0(.din(n3084), .dout(n8398));
    jdff dff_A_wKweXwCq6_1(.din(n8403), .dout(n8400));
    jdff dff_A_JYNCkgNE3_1(.din(n8406), .dout(n8403));
    jdff dff_A_29vt0Iai6_1(.din(n8409), .dout(n8406));
    jdff dff_A_upaUkcFz2_1(.din(n8412), .dout(n8409));
    jdff dff_A_xwS9Vmph3_1(.din(n8415), .dout(n8412));
    jdff dff_A_QwCMM5pe6_1(.din(n8419), .dout(n8415));
    jdff dff_B_RBqfXNkC9_2(.din(n2984), .dout(n8419));
    jdff dff_B_M2eV6rMb1_0(.din(n2980), .dout(n8422));
    jdff dff_B_fECzl2j29_0(.din(n8422), .dout(n8425));
    jdff dff_B_A2vgLadr0_0(.din(n2917), .dout(n8428));
    jdff dff_A_1Do7kB6g2_0(.din(n8433), .dout(n8430));
    jdff dff_A_hFQ53zNg9_0(.din(n2910), .dout(n8433));
    jdff dff_A_TnOnyZIt6_1(.din(n2872), .dout(n8436));
    jdff dff_B_vsnB5BLX1_1(.din(n2011), .dout(n8440));
    jdff dff_B_Hlblfcs99_1(.din(n8440), .dout(n8443));
    jdff dff_B_CF1uAkos3_1(.din(n8443), .dout(n8446));
    jdff dff_B_omwt6g2n2_1(.din(n8446), .dout(n8449));
    jdff dff_B_zEB8zR890_0(.din(n2833), .dout(n8452));
    jdff dff_B_X0fm0r7M0_0(.din(n8452), .dout(n8455));
    jdff dff_A_b3Ut7UhH7_1(.din(n2383), .dout(n8457));
    jdff dff_A_op38Mzqe5_1(.din(n8463), .dout(n8460));
    jdff dff_A_uxOA9Led6_1(.din(n8466), .dout(n8463));
    jdff dff_A_TXy3bDe50_1(.din(n8469), .dout(n8466));
    jdff dff_A_u8gNdpKz3_1(.din(n2062), .dout(n8469));
    jdff dff_B_NjHQMahz2_1(.din(n2032), .dout(n8473));
    jdff dff_B_UQ2eWhvW8_0(.din(n2039), .dout(n8476));
    jdff dff_B_rz3yo8bX1_0(.din(n2003), .dout(n8479));
    jdff dff_B_pgl8Hcza8_0(.din(n8479), .dout(n8482));
    jdff dff_B_iEn66Zu24_0(.din(n8482), .dout(n8485));
    jdff dff_A_9oY2BN3F2_0(.din(n8490), .dout(n8487));
    jdff dff_A_nSYGefZu7_0(.din(n1944), .dout(n8490));
    jdff dff_A_YZHuPk2K1_1(.din(n8496), .dout(n8493));
    jdff dff_A_WfDfgt2O1_1(.din(n1909), .dout(n8496));
    jdff dff_A_F4VMf2ru8_1(.din(n8502), .dout(n8499));
    jdff dff_A_HiQIEYI01_1(.din(n8506), .dout(n8502));
    jdff dff_B_zZtQAI2w2_2(.din(n1882), .dout(n8506));
    jdff dff_A_9nUYdiC35_1(.din(n8511), .dout(n8508));
    jdff dff_A_jmBMnJRL4_1(.din(n8514), .dout(n8511));
    jdff dff_A_c7cyeEG07_1(.din(n8517), .dout(n8514));
    jdff dff_A_oja2GgdL4_1(.din(n8521), .dout(n8517));
    jdff dff_B_qex5kdE77_2(.din(n1855), .dout(n8521));
    jdff dff_B_E2BqAmmD6_1(.din(n2992), .dout(n8524));
    jdff dff_B_hlUP6DoB9_1(.din(n8524), .dout(n8527));
    jdff dff_B_gUT1FJ6E2_1(.din(n8527), .dout(n8530));
    jdff dff_B_VebpQi8Y0_1(.din(n8530), .dout(n8533));
    jdff dff_B_Iv8egv9x3_0(.din(n3020), .dout(n8536));
    jdff dff_B_QS8e2wgJ2_0(.din(n8536), .dout(n8539));
    jdff dff_B_0r9OQegj7_0(.din(n3008), .dout(n8542));
    jdff dff_B_cf8N8jNw3_1(.din(n2643), .dout(n8545));
    jdff dff_B_hzR408JK2_1(.din(n2672), .dout(n8548));
    jdff dff_B_dHwOYEWc2_1(.din(n2699), .dout(n8551));
    jdff dff_B_jbgvIvE76_1(.din(n8551), .dout(n8554));
    jdff dff_B_gUelUwAH4_1(.din(n2657), .dout(n8557));
    jdff dff_B_DjlADNOI5_1(.din(n8557), .dout(n8560));
    jdff dff_B_Jfuhpsui9_1(.din(G89), .dout(n8563));
    jdff dff_B_vti9Bbka6_1(.din(n8563), .dout(n8566));
    jdff dff_B_K6n9Gu5M3_1(.din(n8566), .dout(n8569));
    jdff dff_B_oKPFqOOM6_1(.din(n8569), .dout(n8572));
    jdff dff_B_zGP8pgHY2_1(.din(n8572), .dout(n8575));
    jdff dff_A_Dbnl3XpI9_0(.din(n2661), .dout(n8577));
    jdff dff_B_La6IPfwy8_1(.din(n2598), .dout(n8581));
    jdff dff_A_hfnE4kP47_1(.din(n2635), .dout(n8583));
    jdff dff_A_DYqfH4B18_0(.din(n8590), .dout(n8586));
    jdff dff_B_mUrVDMiY4_3(.din(n2534), .dout(n8590));
    jdff dff_B_NunZNfAB4_0(.din(n2530), .dout(n8593));
    jdff dff_B_UPaggQHO7_0(.din(n8593), .dout(n8596));
    jdff dff_A_yVSrZYYS8_0(.din(n8602), .dout(n8598));
    jdff dff_B_JyTawwKo8_2(.din(n3072), .dout(n8602));
    jdff dff_B_73b3XT5p2_0(.din(n3068), .dout(n8605));
    jdff dff_B_yYE49MnY2_0(.din(n3056), .dout(n8608));
    jdff dff_B_bSp9X1LY2_0(.din(n3048), .dout(n8611));
    jdff dff_B_Crt9Bh7Q1_0(.din(n3040), .dout(n8614));
    jdff dff_B_ipreZXo37_0(.din(n8614), .dout(n8617));
    jdff dff_B_E1vqs5So6_2(.din(n2499), .dout(n8620));
    jdff dff_A_FaUhQEIr8_1(.din(n2464), .dout(n8622));
    jdff dff_B_oyvPw3HP8_0(.din(n2449), .dout(n8626));
    jdff dff_A_uSouiXpl1_0(.din(n8631), .dout(n8628));
    jdff dff_A_kpWQCibZ0_0(.din(n2416), .dout(n8631));
    jdff dff_A_KeBEqL1b9_0(.din(n8637), .dout(n8634));
    jdff dff_A_eXNx4TLQ8_0(.din(n8640), .dout(n8637));
    jdff dff_A_7geiDjfL8_0(.din(n8643), .dout(n8640));
    jdff dff_A_x8erXmeB9_0(.din(n2379), .dout(n8643));
    jdff dff_B_olKMC4kn6_1(.din(n2276), .dout(n8647));
    jdff dff_B_BB9j9eEC6_1(.din(n2291), .dout(n8650));
    jdff dff_B_eyGmmzk53_0(.din(n2287), .dout(n8653));
    jdff dff_B_hc7iIvA21_1(.din(n2231), .dout(n8656));
    jdff dff_A_4emVkdrr4_0(.din(n8661), .dout(n8658));
    jdff dff_A_34VAu1QY2_0(.din(n8664), .dout(n8661));
    jdff dff_A_ZsIGRV5g6_0(.din(n8667), .dout(n8664));
    jdff dff_A_DxoGZ2jD9_0(.din(n8670), .dout(n8667));
    jdff dff_A_KOtvCfEw3_0(.din(n8673), .dout(n8670));
    jdff dff_A_FS4dxPOV8_0(.din(n2825), .dout(n8673));
    jdff dff_B_BaWeFQ4N1_0(.din(n2821), .dout(n8677));
    jdff dff_A_KD4wimPd0_0(.din(n2318), .dout(n8679));
    jdff dff_A_IUzccUPO8_2(.din(n2356), .dout(n8682));
    jdff dff_A_YBvaUdOP4_1(.din(n2348), .dout(n8685));
    jdff dff_A_wB9sN0yI0_0(.din(n2227), .dout(n8688));
    jdff dff_A_cZ3tvlSy3_0(.din(n8694), .dout(n8691));
    jdff dff_A_30epYld30_0(.din(n8697), .dout(n8694));
    jdff dff_A_tK5Ktzi97_0(.din(n8700), .dout(n8697));
    jdff dff_A_tNzfigGw5_0(.din(n8703), .dout(n8700));
    jdff dff_A_M6GKYzr27_0(.din(n8706), .dout(n8703));
    jdff dff_A_yE9Belt04_0(.din(n8709), .dout(n8706));
    jdff dff_A_NdAjGV575_0(.din(n8719), .dout(n8709));
    jdff dff_A_n3OppnbW5_2(.din(n8719), .dout(n8712));
    jdff dff_B_0A8unDCZ9_3(.din(n2173), .dout(n8716));
    jdff dff_B_EsG6Kwdn3_3(.din(n8716), .dout(n8719));
    jdff dff_A_BxmbYe4G3_0(.din(n8724), .dout(n8721));
    jdff dff_A_vxfEyPsa7_0(.din(n8727), .dout(n8724));
    jdff dff_A_DoJtKWku7_0(.din(n8730), .dout(n8727));
    jdff dff_A_wblS193s2_0(.din(n8733), .dout(n8730));
    jdff dff_A_ioM7agik6_0(.din(n8736), .dout(n8733));
    jdff dff_A_a30oBt2Z5_0(.din(n8739), .dout(n8736));
    jdff dff_A_olH5ydUu8_0(.din(n8743), .dout(n8739));
    jdff dff_B_BGQRYwhH0_2(.din(n2789), .dout(n8743));
    jdff dff_B_ocApAAlI3_1(.din(n2749), .dout(n8746));
    jdff dff_B_hntVSUkP1_1(.din(n2753), .dout(n8749));
    jdff dff_B_HRf6BwCS8_1(.din(n8749), .dout(n8752));
    jdff dff_A_rQDQa0fV1_0(.din(n8794), .dout(n8754));
    jdff dff_B_Qcden2jP5_2(.din(n4452), .dout(n8758));
    jdff dff_B_VOOtMusF2_2(.din(n8758), .dout(n8761));
    jdff dff_B_IblNFaSL7_2(.din(n8761), .dout(n8764));
    jdff dff_B_KxNlxfcE2_2(.din(n8764), .dout(n8767));
    jdff dff_B_x5jDJCzn2_2(.din(n8767), .dout(n8770));
    jdff dff_B_RwQl9RZp8_2(.din(n8770), .dout(n8773));
    jdff dff_B_wQV5JdOo7_2(.din(n8773), .dout(n8776));
    jdff dff_B_WKJbX2TY6_2(.din(n8776), .dout(n8779));
    jdff dff_B_YJqjLwA85_2(.din(n8779), .dout(n8782));
    jdff dff_B_UJMbps260_2(.din(n8782), .dout(n8785));
    jdff dff_B_H8qyBEwP5_2(.din(n8785), .dout(n8788));
    jdff dff_B_eQgywDC07_2(.din(n8788), .dout(n8791));
    jdff dff_B_zDz5HAab4_2(.din(n8791), .dout(n8794));
    jdff dff_A_U5A0OWvQ2_0(.din(n8833), .dout(n8796));
    jdff dff_B_8OKTv9XE9_2(.din(n4455), .dout(n8800));
    jdff dff_B_GD9uVb5h8_2(.din(n8800), .dout(n8803));
    jdff dff_B_U2Q129iN0_2(.din(n8803), .dout(n8806));
    jdff dff_B_NgjrwS3f3_2(.din(n8806), .dout(n8809));
    jdff dff_B_EM70p3Km8_2(.din(n8809), .dout(n8812));
    jdff dff_B_xayyrLPC6_2(.din(n8812), .dout(n8815));
    jdff dff_B_0gN2yr7p2_2(.din(n8815), .dout(n8818));
    jdff dff_B_Eo2L0ZQs7_2(.din(n8818), .dout(n8821));
    jdff dff_B_ps9EMUV09_2(.din(n8821), .dout(n8824));
    jdff dff_B_w6PwYQ2n3_2(.din(n8824), .dout(n8827));
    jdff dff_B_SITQzVFv6_2(.din(n8827), .dout(n8830));
    jdff dff_B_0l4IU0o40_2(.din(n8830), .dout(n8833));
    jdff dff_B_mKUwH91I0_1(.din(n4551), .dout(n8836));
    jdff dff_B_kdpLK6Ir2_1(.din(n8836), .dout(n8839));
    jdff dff_B_pKPkoAf66_1(.din(n8839), .dout(n8842));
    jdff dff_B_7X10Oy2z1_1(.din(n8842), .dout(n8845));
    jdff dff_B_YHswpmBN6_1(.din(n8845), .dout(n8848));
    jdff dff_B_hTLr99948_1(.din(n8848), .dout(n8851));
    jdff dff_B_kh0mG0oH5_1(.din(n8851), .dout(n8854));
    jdff dff_B_UXERPa0q1_1(.din(n8854), .dout(n8857));
    jdff dff_B_wiYCOpmh7_1(.din(n8857), .dout(n8860));
    jdff dff_B_YnIuCaKP6_1(.din(n8860), .dout(n8863));
    jdff dff_B_NWEmCtOZ2_1(.din(n8863), .dout(n8866));
    jdff dff_B_wCjmDPvJ6_1(.din(n8866), .dout(n8869));
    jdff dff_A_D6vLbTgQ8_0(.din(n8923), .dout(n8871));
    jdff dff_B_53fwDjvP2_2(.din(n4522), .dout(n8875));
    jdff dff_B_QOYar6qD9_2(.din(n8875), .dout(n8878));
    jdff dff_B_vleLRqDg6_2(.din(n8878), .dout(n8881));
    jdff dff_B_3bb3j1dn9_2(.din(n8881), .dout(n8884));
    jdff dff_B_IPMENRrq7_2(.din(n8884), .dout(n8887));
    jdff dff_B_o3Jo6RyQ2_2(.din(n8887), .dout(n8890));
    jdff dff_B_jhaJRz5v8_2(.din(n8890), .dout(n8893));
    jdff dff_B_LDnfabSV4_2(.din(n8893), .dout(n8896));
    jdff dff_B_LU6tQWlE5_2(.din(n8896), .dout(n8899));
    jdff dff_B_koyHqIvp9_2(.din(n8899), .dout(n8902));
    jdff dff_B_uYehnKMl7_2(.din(n8902), .dout(n8905));
    jdff dff_B_XagOhMGU8_2(.din(n8905), .dout(n8908));
    jdff dff_B_WRvEsVRJ4_2(.din(n8908), .dout(n8911));
    jdff dff_B_0DdkLjYW4_2(.din(n8911), .dout(n8914));
    jdff dff_B_KFLkPMMh7_2(.din(n8914), .dout(n8917));
    jdff dff_B_NaOW4y5v8_2(.din(n8917), .dout(n8920));
    jdff dff_B_6nDF9O8S7_2(.din(n8920), .dout(n8923));
    jdff dff_B_x5PVJcHZ1_1(.din(n4562), .dout(n8926));
    jdff dff_B_EhEJoKax5_1(.din(n8926), .dout(n8929));
    jdff dff_B_gh8Zhfvx7_1(.din(n8929), .dout(n8932));
    jdff dff_B_cZNQdkW77_1(.din(n8932), .dout(n8935));
    jdff dff_B_I7eyIFiw4_1(.din(n8935), .dout(n8938));
    jdff dff_B_zZiQPSHB6_1(.din(n8938), .dout(n8941));
    jdff dff_B_MkJ4RXvv1_1(.din(n8941), .dout(n8944));
    jdff dff_B_N3I8Jjz22_1(.din(n8944), .dout(n8947));
    jdff dff_B_f0Uny1RB5_1(.din(n8947), .dout(n8950));
    jdff dff_B_asBaZ9r35_1(.din(n8950), .dout(n8953));
    jdff dff_B_BeNWbI3f0_1(.din(n8953), .dout(n8956));
    jdff dff_B_latO3i3i6_1(.din(n8956), .dout(n8959));
    jdff dff_B_nxH7yyo68_1(.din(n8959), .dout(n8962));
    jdff dff_B_KQXKqvIk2_0(.din(n4528), .dout(n8965));
    jdff dff_B_IZwVng5o1_0(.din(n8965), .dout(n8968));
    jdff dff_B_vzpbRXCp6_0(.din(n8968), .dout(n8971));
    jdff dff_B_2Bc6UJop7_0(.din(n8971), .dout(n8974));
    jdff dff_B_sqMfXfB26_0(.din(n8974), .dout(n8977));
    jdff dff_B_okDF1nOz8_0(.din(n8977), .dout(n8980));
    jdff dff_B_3Hwed9uF8_0(.din(n8980), .dout(n8983));
    jdff dff_B_gce3rBAo9_0(.din(n8983), .dout(n8986));
    jdff dff_B_PrrVwQBD1_0(.din(n8986), .dout(n8989));
    jdff dff_B_mhxu8Eq72_0(.din(n8989), .dout(n8992));
    jdff dff_B_2ErCsl821_0(.din(n8992), .dout(n8995));
    jdff dff_B_09oTuabG4_0(.din(n8995), .dout(n8998));
    jdff dff_B_HjQBwVVw1_0(.din(n8998), .dout(n9001));
    jdff dff_B_KHPRBnxK0_0(.din(n9001), .dout(n9004));
    jdff dff_A_0Tg0GVpc8_0(.din(n9055), .dout(n9006));
    jdff dff_B_NpolJDHj7_2(.din(n4525), .dout(n9010));
    jdff dff_B_aTtyaxgO4_2(.din(n9010), .dout(n9013));
    jdff dff_B_cvk4diKq2_2(.din(n9013), .dout(n9016));
    jdff dff_B_XN4lpS7F4_2(.din(n9016), .dout(n9019));
    jdff dff_B_VzR6Q3Nw9_2(.din(n9019), .dout(n9022));
    jdff dff_B_WaMjxWFi9_2(.din(n9022), .dout(n9025));
    jdff dff_B_wzO7q3NX5_2(.din(n9025), .dout(n9028));
    jdff dff_B_EljRkBnR8_2(.din(n9028), .dout(n9031));
    jdff dff_B_FjHYRCtP3_2(.din(n9031), .dout(n9034));
    jdff dff_B_Wyodgqcx1_2(.din(n9034), .dout(n9037));
    jdff dff_B_5WyXIVz35_2(.din(n9037), .dout(n9040));
    jdff dff_B_CvXfG5r89_2(.din(n9040), .dout(n9043));
    jdff dff_B_mbFam3nO9_2(.din(n9043), .dout(n9046));
    jdff dff_B_XHdLJZGC4_2(.din(n9046), .dout(n9049));
    jdff dff_B_UQDYOXCH3_2(.din(n9049), .dout(n9052));
    jdff dff_B_Hq71TNA62_2(.din(n9052), .dout(n9055));
    jdff dff_B_mr5mYk7H5_0(.din(n4598), .dout(n9058));
    jdff dff_B_QD0a7OGU7_0(.din(n4594), .dout(n9061));
    jdff dff_B_P52bzwOL2_0(.din(n9061), .dout(n9064));
    jdff dff_B_6E67m9nk2_0(.din(n9064), .dout(n9067));
    jdff dff_B_o6C0FC1J8_0(.din(n9067), .dout(n9070));
    jdff dff_B_gmsbbxjL8_0(.din(n9070), .dout(n9073));
    jdff dff_B_pP0s51ua1_0(.din(n9073), .dout(n9076));
    jdff dff_B_173T7hMJ2_0(.din(n3729), .dout(n9079));
    jdff dff_B_Q74RQj760_0(.din(n3717), .dout(n9082));
    jdff dff_B_HWQXCFiG4_1(.din(n3705), .dout(n9085));
    jdff dff_B_NHTV8UlK1_1(.din(n3697), .dout(n9088));
    jdff dff_B_fWbOweMG4_0(.din(n3669), .dout(n9091));
    jdff dff_B_fjEFjj683_1(.din(n3641), .dout(n9094));
    jdff dff_B_EhhukHxl3_1(.din(n9094), .dout(n9097));
    jdff dff_B_uzyJlzBQ0_1(.din(n3633), .dout(n9100));
    jdff dff_B_9IECpHVC3_1(.din(n3583), .dout(n9103));
    jdff dff_B_Wv8yPjb91_1(.din(n9103), .dout(n9106));
    jdff dff_B_pSO67Ttc4_1(.din(n9106), .dout(n9109));
    jdff dff_B_Y3DHXPlw4_1(.din(n9109), .dout(n9112));
    jdff dff_B_DJ4w6L5y8_1(.din(n3587), .dout(n9115));
    jdff dff_B_OGURsFGT2_1(.din(n9115), .dout(n9118));
    jdff dff_B_W377iLEv9_1(.din(n9118), .dout(n9121));
    jdff dff_B_SyQToNJc4_1(.din(n9121), .dout(n9124));
    jdff dff_B_BdmlA7k07_1(.din(n3605), .dout(n9127));
    jdff dff_B_9gASExGS4_0(.din(n3579), .dout(n9130));
    jdff dff_B_tDGVdp7M2_0(.din(n9130), .dout(n9133));
    jdff dff_B_sVv5WnBc8_1(.din(n3499), .dout(n9136));
    jdff dff_B_rqPeaL4Q4_1(.din(n9136), .dout(n9139));
    jdff dff_B_UYU4h3RQ3_1(.din(n9139), .dout(n9142));
    jdff dff_B_oe85dSHx4_1(.din(n9142), .dout(n9145));
    jdff dff_B_Z1bZWMPx7_1(.din(n9145), .dout(n9148));
    jdff dff_B_TvFokxhq6_1(.din(n3507), .dout(n9151));
    jdff dff_B_xHL8bKfi8_1(.din(n9151), .dout(n9154));
    jdff dff_B_ORUhP1w48_1(.din(n9154), .dout(n9157));
    jdff dff_B_boMQhpJ27_0(.din(n3559), .dout(n9160));
    jdff dff_B_Mq6MvMiN9_0(.din(n9160), .dout(n9163));
    jdff dff_B_opeCNCVQ1_0(.din(n9163), .dout(n9166));
    jdff dff_B_bpWNMMEc7_0(.din(n9166), .dout(n9169));
    jdff dff_B_cRJVO95d6_0(.din(n4276), .dout(n9172));
    jdff dff_B_B2EznjiX3_0(.din(n9172), .dout(n9175));
    jdff dff_B_gjvsLsyS4_0(.din(n9175), .dout(n9178));
    jdff dff_B_WHtaxa8G1_1(.din(n4209), .dout(n9181));
    jdff dff_B_nlwoff1o3_1(.din(n9181), .dout(n9184));
    jdff dff_B_0ZQfZymY9_1(.din(n9184), .dout(n9187));
    jdff dff_B_BRbGO4Yg4_1(.din(n4213), .dout(n9190));
    jdff dff_B_cIktG6lr3_1(.din(n9190), .dout(n9193));
    jdff dff_B_LfJWX3D13_1(.din(n9193), .dout(n9196));
    jdff dff_B_MCaZvy6c3_0(.din(n4264), .dout(n9199));
    jdff dff_B_2hXY8mZJ4_0(.din(n9199), .dout(n9202));
    jdff dff_B_uQvFpwT72_0(.din(n9202), .dout(n9205));
    jdff dff_B_ZhNlUfdm8_0(.din(G174), .dout(n9208));
    jdff dff_B_OEvkFNga5_0(.din(G173), .dout(n9211));
    jdff dff_B_bRo8Z4hO6_0(.din(G176), .dout(n9214));
    jdff dff_B_kwT9n1fz3_0(.din(G175), .dout(n9217));
    jdff dff_B_jMZecd1B1_0(.din(n1952), .dout(n9220));
    jdff dff_B_xFKgSs601_0(.din(G177), .dout(n9223));
    jdff dff_B_mds2AIK08_0(.din(n1913), .dout(n9226));
    jdff dff_B_2pGwruPz1_0(.din(n1859), .dout(n9229));
    jdff dff_A_FCPrPmIm8_0(.din(n1890), .dout(n9231));
    jdff dff_B_uYOex2N95_0(.din(n1886), .dout(n9235));
    jdff dff_B_1NXFRMjk4_1(.din(n4111), .dout(n9238));
    jdff dff_B_rreQ0XYf0_1(.din(n9238), .dout(n9241));
    jdff dff_B_gICgOpXL2_1(.din(n4169), .dout(n9244));
    jdff dff_B_yLk5tBE51_1(.din(n9244), .dout(n9247));
    jdff dff_B_p3lLlLER1_1(.din(n4172), .dout(n9250));
    jdff dff_B_Ua5UgG9c8_0(.din(n4161), .dout(n9253));
    jdff dff_B_N64ZuN0W7_0(.din(n4157), .dout(n9256));
    jdff dff_B_rtQVUCQU1_0(.din(n2541), .dout(n9259));
    jdff dff_B_fPYqTgMv3_0(.din(n9259), .dout(n9262));
    jdff dff_B_83WXd5ql7_0(.din(n2679), .dout(n9265));
    jdff dff_B_ppmXzpJe8_0(.din(n9265), .dout(n9268));
    jdff dff_B_1MoapjDq3_0(.din(n2612), .dout(n9271));
    jdff dff_B_PhDfeFx85_0(.din(n9271), .dout(n9274));
    jdff dff_B_rf7vgArF7_0(.din(n2571), .dout(n9277));
    jdff dff_B_rVvKV7Bp3_0(.din(n9277), .dout(n9280));
    jdff dff_B_n43mFXus8_1(.din(n4119), .dout(n9283));
    jdff dff_B_lQ8Q3Dii3_1(.din(n9283), .dout(n9286));
    jdff dff_B_v0ffNHLM7_1(.din(n9286), .dout(n9289));
    jdff dff_B_CN1hRy5D4_0(.din(n2506), .dout(n9292));
    jdff dff_B_7XSr0N1X0_0(.din(n9292), .dout(n9295));
    jdff dff_A_xTpTo3FQ6_1(.din(n2480), .dout(n9297));
    jdff dff_B_8XEg0JBA1_0(.din(n2476), .dout(n9301));
    jdff dff_B_0p1asTaz8_0(.din(n2426), .dout(n9304));
    jdff dff_B_GHMBKMEz3_0(.din(n9304), .dout(n9307));
    jdff dff_B_3u7H70DV1_0(.din(n4115), .dout(n9310));
    jdff dff_B_ACQkRp2d8_0(.din(G44), .dout(n9313));
    jdff dff_B_ZkCoSXX81_0(.din(n4099), .dout(n9316));
    jdff dff_B_lXAUZjrw9_0(.din(n9316), .dout(n9319));
    jdff dff_B_FVEpOpmI2_0(.din(n2295), .dout(n9322));
    jdff dff_B_Cq4SEy4M3_0(.din(n2177), .dout(n9325));
    jdff dff_B_VWQRY0eh8_0(.din(n2235), .dout(n9328));
    jdff dff_B_pEGy5yFX6_0(.din(n2204), .dout(n9331));
    jdff dff_B_QcCZd2tT0_0(.din(n4077), .dout(n9334));
    jdff dff_B_lMdIjjqA3_0(.din(G115), .dout(n9337));
    jdff dff_A_jov50joB5_1(.din(n4073), .dout(n9339));
    jdff dff_B_y2mL8afH4_0(.din(n2145), .dout(n9343));
    jdff dff_B_yCOS2wms3_0(.din(n2118), .dout(n9346));
    jdff dff_B_BdF6J7Nd9_0(.din(n2090), .dout(n9349));
    jdff dff_B_UYt0YtB46_0(.din(n2066), .dout(n9352));
    jdff dff_A_VL9wH6h17_0(.din(n9357), .dout(n9354));
    jdff dff_A_XC64y0ZQ7_0(.din(n2329), .dout(n9357));
    jdff dff_B_h00Pwn007_0(.din(n2325), .dout(n9361));
    jdff dff_B_fIb3v3qv5_1(.din(n4023), .dout(n9364));
    jdff dff_B_xEb6tKc84_0(.din(n4049), .dout(n9367));
    jdff dff_B_P2YIAgvt6_0(.din(n9367), .dout(n9370));
    jdff dff_B_4Ng3MVty1_0(.din(n4045), .dout(n9373));
    jdff dff_B_mxs537I87_0(.din(n9373), .dout(n9376));
    jdff dff_A_2DeFixeh3_2(.din(n9381), .dout(n9378));
    jdff dff_A_p6fYGlLf3_2(.din(G18), .dout(n9381));
    jdff dff_A_n6hM84nC4_0(.din(n9387), .dout(n9384));
    jdff dff_A_VqC2Fu7o5_0(.din(n3271), .dout(n9387));
    jdff dff_B_7fLkiLQM3_0(.din(G168), .dout(n9391));
    jdff dff_A_c2BPqbnV3_0(.din(n9396), .dout(n9393));
    jdff dff_A_v1DXBwy66_0(.din(n3198), .dout(n9396));
    jdff dff_B_t28gJu808_0(.din(G169), .dout(n9400));
    jdff dff_A_tvyGr8hS2_0(.din(n1245), .dout(n9402));
    jdff dff_A_mwjuaXS58_1(.din(n1245), .dout(n9405));
    jdff dff_B_cmy3iLci6_1(.din(n3993), .dout(n9409));
    jdff dff_B_b19WWDy46_0(.din(G166), .dout(n9412));
    jdff dff_A_RBRzs81B1_0(.din(n3140), .dout(n9414));
    jdff dff_B_FnEjt97S5_0(.din(G167), .dout(n9418));
    jdff dff_A_L9yEVs9h8_0(.din(n9423), .dout(n9420));
    jdff dff_A_GksR6ZpJ8_0(.din(n9426), .dout(n9423));
    jdff dff_A_CfZ6Oqln4_0(.din(n3990), .dout(n9426));
    jdff dff_B_64dqJnW15_1(.din(n3788), .dout(n9430));
    jdff dff_B_W3BPbTjj3_1(.din(n9430), .dout(n9433));
    jdff dff_B_OP2RUF7k2_0(.din(n3966), .dout(n9436));
    jdff dff_B_Lcgy86XL0_0(.din(n1901), .dout(n9439));
    jdff dff_B_U1958RBQ3_0(.din(n1874), .dout(n9442));
    jdff dff_B_hfEIVdUV0_1(.din(n3954), .dout(n9445));
    jdff dff_B_ZvV1HQX72_0(.din(n1967), .dout(n9448));
    jdff dff_B_m2voZ3vE6_0(.din(n1928), .dout(n9451));
    jdff dff_A_xccNKG1p6_1(.din(G2208), .dout(n9453));
    jdff dff_B_UY3GNvtW9_0(.din(n2968), .dout(n9457));
    jdff dff_B_eCcZfGh83_0(.din(n2944), .dout(n9460));
    jdff dff_B_gbjOsGnH4_0(.din(n2891), .dout(n9463));
    jdff dff_B_l5t1Lzlf2_0(.din(n2864), .dout(n9466));
    jdff dff_A_81yKPvvS6_0(.din(n9471), .dout(n9468));
    jdff dff_A_MOHz5gvg5_0(.din(n1851), .dout(n9471));
    jdff dff_B_Ys5oJSE10_0(.din(n1847), .dout(n9475));
    jdff dff_B_NBUZtjFn9_1(.din(n3887), .dout(n9478));
    jdff dff_B_Q9WaGEmw0_0(.din(n3915), .dout(n9481));
    jdff dff_B_9hGaIqOb4_0(.din(n9481), .dout(n9484));
    jdff dff_B_R6DqXCQT1_0(.din(n3286), .dout(n9487));
    jdff dff_A_1y77Buen6_0(.din(G18), .dout(n9489));
    jdff dff_B_FkoeeYcx3_0(.din(n3182), .dout(n9493));
    jdff dff_A_Um3i6k0s2_0(.din(n3159), .dout(n9495));
    jdff dff_B_zwpHeb496_0(.din(n3155), .dout(n9499));
    jdff dff_B_hCoIS9vy3_1(.din(n3879), .dout(n9502));
    jdff dff_B_4F3mVGZg2_0(.din(n3232), .dout(n9505));
    jdff dff_B_6eM1AfF22_0(.din(n3213), .dout(n9508));
    jdff dff_A_Aax5Nc2t1_1(.din(G1459), .dout(n9510));
    jdff dff_B_AqWoWdRJ9_1(.din(n3826), .dout(n9514));
    jdff dff_B_1rCp1k1u8_1(.din(n9514), .dout(n9517));
    jdff dff_B_UT9nz9814_1(.din(n3830), .dout(n9520));
    jdff dff_B_fsMbef7P3_1(.din(n9520), .dout(n9523));
    jdff dff_B_aLTbXciP5_1(.din(n3833), .dout(n9526));
    jdff dff_A_Rjv8E4uC9_1(.din(n2522), .dout(n9528));
    jdff dff_A_DWrTK79g5_2(.din(n2522), .dout(n9531));
    jdff dff_B_IUEL5QAU1_1(.din(n2514), .dout(n9535));
    jdff dff_B_hNhDWOew7_1(.din(n2484), .dout(n9538));
    jdff dff_A_8QpsK7Yt1_1(.din(n2445), .dout(n9540));
    jdff dff_A_5CD2Eegm4_2(.din(n2445), .dout(n9543));
    jdff dff_B_PUf4qp3b3_1(.din(n2434), .dout(n9547));
    jdff dff_A_1PkpiUyh1_1(.din(n2412), .dout(n9549));
    jdff dff_A_QYNBPp378_2(.din(n2412), .dout(n9552));
    jdff dff_B_JfloGEvr0_1(.din(n2401), .dout(n9556));
    jdff dff_A_SJRSbQzT0_1(.din(n2590), .dout(n9558));
    jdff dff_A_M23IpCZd7_2(.din(n2590), .dout(n9561));
    jdff dff_B_uXICOqHD1_1(.din(n2579), .dout(n9565));
    jdff dff_A_Omj3E1au7_0(.din(n2695), .dout(n9567));
    jdff dff_A_OMALyz483_2(.din(n2695), .dout(n9570));
    jdff dff_B_tcaMqhgn1_1(.din(n2687), .dout(n9574));
    jdff dff_A_d6l7CZCQ0_1(.din(n2631), .dout(n9576));
    jdff dff_A_r5guVyE14_2(.din(n2631), .dout(n9579));
    jdff dff_B_zE8vol1i0_1(.din(n2620), .dout(n9583));
    jdff dff_A_IJjwYJTk3_0(.din(n9588), .dout(n9585));
    jdff dff_A_MeVxKv7k8_0(.din(n3823), .dout(n9588));
    jdff dff_A_ZmKoTLCU6_1(.din(G3698), .dout(n9591));
    jdff dff_B_CzetVjBx0_3(.din(n2560), .dout(n9595));
    jdff dff_B_Bh5QiV947_1(.din(n2549), .dout(n9598));
    jdff dff_B_pos8EslO2_1(.din(n3741), .dout(n9601));
    jdff dff_B_bgi1gc382_1(.din(n9601), .dout(n9604));
    jdff dff_B_DbGk8HA50_1(.din(n9604), .dout(n9607));
    jdff dff_B_SJTdq7ix4_1(.din(n3749), .dout(n9610));
    jdff dff_B_GSjpiOkW6_0(.din(n3776), .dout(n9613));
    jdff dff_B_8LCFIIXv6_0(.din(n9613), .dout(n9616));
    jdff dff_A_8eJPHOff4_1(.din(G4393), .dout(n9618));
    jdff dff_A_3iXJCCI03_1(.din(n455), .dout(n9621));
    jdff dff_B_aDgzSQ3W6_1(.din(n2153), .dout(n9625));
    jdff dff_B_sNtu3yve4_1(.din(n2126), .dout(n9628));
    jdff dff_B_XUlCmyH13_1(.din(n2098), .dout(n9631));
    jdff dff_B_B0owYQxb4_1(.din(n2074), .dout(n9634));
    jdff dff_B_F9BIbIMB5_1(.din(n2303), .dout(n9637));
    jdff dff_B_WDAEk5L34_1(.din(n2185), .dout(n9640));
    jdff dff_A_bQRHzGDs9_0(.din(n2344), .dout(n9642));
    jdff dff_B_02keszY75_1(.din(n2333), .dout(n9646));
    jdff dff_B_DAJuA5HC0_1(.din(n2243), .dout(n9649));
    jdff dff_B_P2O9N3ze6_1(.din(n2212), .dout(n9652));
    jdff dff_B_WBgQZcFf6_3(.din(n1824), .dout(n9655));
    jdff dff_B_Bcaf6cA64_3(.din(n9655), .dout(n9658));
    jdff dff_B_3eVDKZ8r3_3(.din(n9658), .dout(n9661));
    jdff dff_B_lqrthS1O3_3(.din(n9661), .dout(n9664));
    jdff dff_B_Jj3NHDP84_3(.din(n9664), .dout(n9667));
    jdff dff_B_KXnUiTzW5_3(.din(n9667), .dout(n9670));
    jdff dff_B_JD2Rz16V0_3(.din(n9670), .dout(n9673));
    jdff dff_B_aR637i0J9_3(.din(n9673), .dout(n9676));
    jdff dff_B_TJ6EZ4fW9_3(.din(n9676), .dout(n9679));
    jdff dff_B_uJQ2eOXl4_3(.din(n9679), .dout(n9682));
    jdff dff_B_0CMEndwP5_3(.din(n9682), .dout(n9685));
    jdff dff_B_V69zn5WE9_3(.din(n9685), .dout(n9688));
    jdff dff_B_SbyWKT4c1_3(.din(n9688), .dout(n9691));
    jdff dff_B_b5gDHqmV4_3(.din(n9691), .dout(n9694));
    jdff dff_B_kkRlhK8R5_3(.din(n9694), .dout(n9697));
    jdff dff_B_CXby5lLn8_3(.din(n9697), .dout(n9700));
    jdff dff_B_jh6Pz9Zb5_3(.din(n9700), .dout(n9703));
    jdff dff_B_5R7QQSBq3_3(.din(n9703), .dout(n9706));
    jdff dff_B_cB0oiWbK4_3(.din(n9706), .dout(n9709));
    jdff dff_B_ohEwP5um6_3(.din(n9709), .dout(n9712));
    jdff dff_B_fJVRGy5q8_3(.din(n9712), .dout(n9715));
    jdff dff_B_2oZZjT7X1_1(.din(n1813), .dout(n9718));
    jdff dff_B_KgojfExN2_1(.din(n4635), .dout(n9721));
    jdff dff_B_8UnFFy893_1(.din(n9721), .dout(n9724));
    jdff dff_B_tuSUn7M79_1(.din(n9724), .dout(n9727));
    jdff dff_B_bOcn9bFA5_1(.din(n9727), .dout(n9730));
    jdff dff_B_rCxV8oK94_1(.din(n9730), .dout(n9733));
    jdff dff_B_pXv33GAe6_1(.din(n9733), .dout(n9736));
    jdff dff_B_YSYV19dJ5_1(.din(n9736), .dout(n9739));
    jdff dff_B_ATGUKbGM5_1(.din(n9739), .dout(n9742));
    jdff dff_B_SzUDHR6b7_1(.din(n9742), .dout(n9745));
    jdff dff_B_LpWTZVwP6_1(.din(n9745), .dout(n9748));
    jdff dff_B_p6Dvi9i21_1(.din(n9748), .dout(n9751));
    jdff dff_B_oUEGXJvf0_1(.din(n9751), .dout(n9754));
    jdff dff_B_5FxkY6i03_1(.din(n9754), .dout(n9757));
    jdff dff_B_z5Hs1uc00_1(.din(n9757), .dout(n9760));
    jdff dff_B_yo79W8XW9_1(.din(n9760), .dout(n9763));
    jdff dff_A_X8KAt6jb7_0(.din(n1807), .dout(n9765));
    jdff dff_A_mNktjaKO5_1(.din(n1807), .dout(n9768));
    jdff dff_A_lX3g4Itf2_0(.din(n9799), .dout(n9771));
    jdff dff_B_dM42cA8C7_2(.din(n4701), .dout(n9775));
    jdff dff_B_MJTYYIxQ6_2(.din(n9775), .dout(n9778));
    jdff dff_B_GXOXjQLM0_2(.din(n9778), .dout(n9781));
    jdff dff_B_zEDiIaCw9_2(.din(n9781), .dout(n9784));
    jdff dff_B_G2n4ifS46_2(.din(n9784), .dout(n9787));
    jdff dff_B_yjrW8SYW8_2(.din(n9787), .dout(n9790));
    jdff dff_B_ldsqRPJP1_2(.din(n9790), .dout(n9793));
    jdff dff_B_AU69szzi5_2(.din(n9793), .dout(n9796));
    jdff dff_B_R8RVR4Em2_2(.din(n9796), .dout(n9799));
    jdff dff_A_ltbWdfQG3_0(.din(n9823), .dout(n9801));
    jdff dff_B_44HkEJvN5_2(.din(n4704), .dout(n9805));
    jdff dff_B_Qogw2FEU5_2(.din(n9805), .dout(n9808));
    jdff dff_B_c373aXyp3_2(.din(n9808), .dout(n9811));
    jdff dff_B_G54LPRDw9_2(.din(n9811), .dout(n9814));
    jdff dff_B_XD9VrQfq4_2(.din(n9814), .dout(n9817));
    jdff dff_B_BBr7EVxo5_2(.din(n9817), .dout(n9820));
    jdff dff_B_EsLk7yv80_2(.din(n9820), .dout(n9823));
    jdff dff_B_t0V9Cd6B6_1(.din(n4820), .dout(n9826));
    jdff dff_B_KUAIJL757_1(.din(n9826), .dout(n9829));
    jdff dff_B_oFG2qDPi6_1(.din(n9829), .dout(n9832));
    jdff dff_B_qu9AU5DH7_1(.din(n9832), .dout(n9835));
    jdff dff_B_e1LrZ9FG8_1(.din(n9835), .dout(n9838));
    jdff dff_B_Kqxsl6xq7_1(.din(n9838), .dout(n9841));
    jdff dff_B_0BdZoDHv6_1(.din(n9841), .dout(n9844));
    jdff dff_B_HtZdZ1D74_1(.din(n9844), .dout(n9847));
    jdff dff_B_iCMngwBU5_1(.din(n9847), .dout(n9850));
    jdff dff_B_d5fv3hk86_1(.din(n9850), .dout(n9853));
    jdff dff_B_SoWd5YXX4_1(.din(n9853), .dout(n9856));
    jdff dff_B_ryspUru82_1(.din(n9856), .dout(n9859));
    jdff dff_B_aYOpmNQu3_1(.din(n9859), .dout(n9862));
    jdff dff_B_9zrF3Isv5_1(.din(n9862), .dout(n9865));
    jdff dff_B_U8EmEL2h4_1(.din(n9865), .dout(n9868));
    jdff dff_B_LNzOzkYx4_0(.din(n4998), .dout(n9871));
    jdff dff_B_gnBCZDhH4_0(.din(n9871), .dout(n9874));
    jdff dff_B_J5xJEgnn2_0(.din(n4990), .dout(n9877));
    jdff dff_B_QTp7Gtxt6_0(.din(n9877), .dout(n9880));
    jdff dff_B_xR1d7E2a2_1(.din(n4948), .dout(n9883));
    jdff dff_B_u3cQHpfZ3_1(.din(n9883), .dout(n9886));
    jdff dff_B_AM7IyKHC6_1(.din(n9886), .dout(n9889));
    jdff dff_B_aI1HuN814_1(.din(n9889), .dout(n9892));
    jdff dff_B_HkRHqI9f6_1(.din(n4952), .dout(n9895));
    jdff dff_B_V4RiUXRg5_1(.din(n9895), .dout(n9898));
    jdff dff_B_AF1N2f3f8_1(.din(n9898), .dout(n9901));
    jdff dff_B_RAz5LPa67_1(.din(n9901), .dout(n9904));
    jdff dff_B_PSFf9n4w9_1(.din(n9904), .dout(n9907));
    jdff dff_B_HFTzXLQg0_1(.din(n9907), .dout(n9910));
    jdff dff_B_PYhRQtCE6_1(.din(n9910), .dout(n9913));
    jdff dff_B_X1okK80g2_1(.din(n4967), .dout(n9916));
    jdff dff_B_aeoxuii34_0(.din(n4974), .dout(n9919));
    jdff dff_B_Nh6WyFZo2_1(.din(n4970), .dout(n9922));
    jdff dff_B_xVxqDQz99_0(.din(n4956), .dout(n9925));
    jdff dff_A_189A6ZlH4_1(.din(n9930), .dout(n9927));
    jdff dff_A_eTuTsUzN9_1(.din(n9933), .dout(n9930));
    jdff dff_A_YeVLCuEd5_1(.din(n9936), .dout(n9933));
    jdff dff_A_7Sb9knEw0_1(.din(n9939), .dout(n9936));
    jdff dff_A_sBamll1V9_1(.din(n9942), .dout(n9939));
    jdff dff_A_pWlNBqqc1_1(.din(n9945), .dout(n9942));
    jdff dff_A_HTXHixWY6_1(.din(n9948), .dout(n9945));
    jdff dff_A_qm6gHRym3_1(.din(n9951), .dout(n9948));
    jdff dff_A_buTZcA207_1(.din(n9954), .dout(n9951));
    jdff dff_A_gQJETuFf1_1(.din(n4496), .dout(n9954));
    jdff dff_B_Qst8B18I0_1(.din(n4489), .dout(n9958));
    jdff dff_A_WVjGtuSH1_1(.din(n9963), .dout(n9960));
    jdff dff_A_mLbPJ5GU7_1(.din(n9966), .dout(n9963));
    jdff dff_A_OEGK5aPO0_1(.din(n9969), .dout(n9966));
    jdff dff_A_cA44UuRA4_1(.din(n9972), .dout(n9969));
    jdff dff_A_dtyJ8XnP2_1(.din(n9975), .dout(n9972));
    jdff dff_A_JTWpSgbv7_1(.din(n9978), .dout(n9975));
    jdff dff_A_TMhhQwq76_1(.din(n9981), .dout(n9978));
    jdff dff_A_sy9AdmYK5_1(.din(n9984), .dout(n9981));
    jdff dff_A_SuUZyTFP8_1(.din(n9988), .dout(n9984));
    jdff dff_B_KlXKBtaX3_2(.din(n4458), .dout(n9988));
    jdff dff_B_cUKLYI2q2_0(.din(n4936), .dout(n9991));
    jdff dff_B_LMw4H1BS8_0(.din(n9991), .dout(n9994));
    jdff dff_B_nHV2rcZB0_0(.din(n9994), .dout(n9997));
    jdff dff_B_3Z2683L62_1(.din(n4912), .dout(n10000));
    jdff dff_B_INRxn0Zf8_1(.din(n10000), .dout(n10003));
    jdff dff_B_qYyCQUq50_0(.din(n4924), .dout(n10006));
    jdff dff_B_puz4657M8_0(.din(n10006), .dout(n10009));
    jdff dff_B_h1hNkmOI9_0(.din(n10009), .dout(n10012));
    jdff dff_B_WS9Io77u8_1(.din(n4916), .dout(n10015));
    jdff dff_A_t08G5Bbe2_1(.din(n10020), .dout(n10017));
    jdff dff_A_LJD4TZIk5_1(.din(n10023), .dout(n10020));
    jdff dff_A_N9e8tcqr4_1(.din(n10026), .dout(n10023));
    jdff dff_A_F0FfSBz80_1(.din(n10029), .dout(n10026));
    jdff dff_A_B62EhZho3_1(.din(n10032), .dout(n10029));
    jdff dff_A_gKREzjCS2_1(.din(n10035), .dout(n10032));
    jdff dff_A_iasVbBSK8_1(.din(n10038), .dout(n10035));
    jdff dff_A_zCPEnLGe2_1(.din(n10041), .dout(n10038));
    jdff dff_A_HnnnsTka4_1(.din(n10060), .dout(n10041));
    jdff dff_B_kXOVzd9I2_2(.din(n4449), .dout(n10045));
    jdff dff_B_HTieYIFO7_2(.din(n10045), .dout(n10048));
    jdff dff_B_nevWWI0v8_2(.din(n10048), .dout(n10051));
    jdff dff_B_iSRBWQMZ6_2(.din(n10051), .dout(n10054));
    jdff dff_B_NIXbY9Ao0_2(.din(n10054), .dout(n10057));
    jdff dff_B_WUarIzIc6_2(.din(n10057), .dout(n10060));
    jdff dff_A_kUmEGgAQ2_1(.din(n4896), .dout(n10062));
    jdff dff_B_bKnFP9Jd3_0(.din(n4881), .dout(n10066));
    jdff dff_B_majlC20b5_0(.din(n10066), .dout(n10069));
    jdff dff_B_gLo6NdRF1_0(.din(n10069), .dout(n10072));
    jdff dff_B_Mm9GiAn24_0(.din(n10072), .dout(n10075));
    jdff dff_B_qRoOA2Qd9_0(.din(n10075), .dout(n10078));
    jdff dff_B_UMNJLbhl3_1(.din(n4854), .dout(n10081));
    jdff dff_B_4Vp9XJcD5_1(.din(n10081), .dout(n10084));
    jdff dff_B_9THo75lP0_1(.din(n10084), .dout(n10087));
    jdff dff_B_7Hmehq3E6_1(.din(n10087), .dout(n10090));
    jdff dff_B_r8AFxmE49_1(.din(n10090), .dout(n10093));
    jdff dff_B_jMIpVqyN4_1(.din(n10093), .dout(n10096));
    jdff dff_B_WfMAqJW37_0(.din(n4869), .dout(n10099));
    jdff dff_A_wXk9aqtR3_1(.din(n10104), .dout(n10101));
    jdff dff_A_C957GCgo6_1(.din(n10107), .dout(n10104));
    jdff dff_A_4vVxTJGK5_1(.din(n10110), .dout(n10107));
    jdff dff_A_fBWZPxuy6_1(.din(n10113), .dout(n10110));
    jdff dff_A_fTYnZjd86_1(.din(n10116), .dout(n10113));
    jdff dff_A_twiNsobd1_1(.din(n10119), .dout(n10116));
    jdff dff_A_Ad1WD2fp6_1(.din(n10122), .dout(n10119));
    jdff dff_A_se79etU97_1(.din(n10125), .dout(n10122));
    jdff dff_A_pOl1XUOm4_1(.din(n10128), .dout(n10125));
    jdff dff_A_JL2dJkcJ1_1(.din(n10131), .dout(n10128));
    jdff dff_A_vE50oDBr4_1(.din(n10135), .dout(n10131));
    jdff dff_B_UthSIp5O4_2(.din(n4612), .dout(n10135));
    jdff dff_B_8ozVRkdB5_0(.din(n4846), .dout(n10138));
    jdff dff_B_eAaxFN4c8_0(.din(n10138), .dout(n10141));
    jdff dff_B_GRpiWZ8t0_0(.din(n10141), .dout(n10144));
    jdff dff_B_sJXleZJV5_0(.din(n10144), .dout(n10147));
    jdff dff_B_82qNFKIF8_0(.din(n10147), .dout(n10150));
    jdff dff_B_B5qAVPdK2_0(.din(n10150), .dout(n10153));
    jdff dff_B_KoHBeDLk7_0(.din(n4830), .dout(n10156));
    jdff dff_A_xqicetMq9_0(.din(n10161), .dout(n10158));
    jdff dff_A_tj41q6wh8_0(.din(n10213), .dout(n10161));
    jdff dff_A_E6LFlpmq0_2(.din(n10167), .dout(n10164));
    jdff dff_A_k9KSXCIp0_2(.din(n10170), .dout(n10167));
    jdff dff_A_VYR4DypP3_2(.din(n10173), .dout(n10170));
    jdff dff_A_73fzXHMZ8_2(.din(n10176), .dout(n10173));
    jdff dff_A_PxD9yZqd5_2(.din(n10179), .dout(n10176));
    jdff dff_A_w0Iz6dlr5_2(.din(n10182), .dout(n10179));
    jdff dff_A_XqWRHUXo0_2(.din(n10185), .dout(n10182));
    jdff dff_A_DW5A0erl8_2(.din(n10188), .dout(n10185));
    jdff dff_A_BwmJgd5x7_2(.din(n10191), .dout(n10188));
    jdff dff_A_SLMe2BuB5_2(.din(n10194), .dout(n10191));
    jdff dff_A_uAmDQLEZ8_2(.din(n10197), .dout(n10194));
    jdff dff_A_NSIIuSUk2_2(.din(n10200), .dout(n10197));
    jdff dff_A_dlooAmvU0_2(.din(n10213), .dout(n10200));
    jdff dff_B_bRi3SU7w6_3(.din(n4609), .dout(n10204));
    jdff dff_B_Mb7QQDlE8_3(.din(n10204), .dout(n10207));
    jdff dff_B_atMmZB8Y1_3(.din(n10207), .dout(n10210));
    jdff dff_B_SI0CUn5e3_3(.din(n10210), .dout(n10213));
    jdff dff_A_BIyh4ZNm7_1(.din(n10218), .dout(n10215));
    jdff dff_A_bU0yKjex8_1(.din(n10221), .dout(n10218));
    jdff dff_A_garw6vSx8_1(.din(n10224), .dout(n10221));
    jdff dff_A_0bdyKZb81_1(.din(n10227), .dout(n10224));
    jdff dff_A_iatti9uZ2_1(.din(n4823), .dout(n10227));
    jdff dff_A_2EEXSPAA6_1(.din(n10233), .dout(n10230));
    jdff dff_A_54ofLsbF8_1(.din(n10236), .dout(n10233));
    jdff dff_A_7jKDsxoq3_1(.din(n10239), .dout(n10236));
    jdff dff_A_O2xzF8Dh2_1(.din(n10242), .dout(n10239));
    jdff dff_A_8QDMDMFw1_1(.din(n10245), .dout(n10242));
    jdff dff_A_mvDqumTc6_1(.din(n10248), .dout(n10245));
    jdff dff_A_uX2DG70z2_1(.din(n10264), .dout(n10248));
    jdff dff_B_jNmrxi3S8_2(.din(n4646), .dout(n10252));
    jdff dff_B_cZdZCxDD9_2(.din(n10252), .dout(n10255));
    jdff dff_B_Nc8LrthW4_2(.din(n10255), .dout(n10258));
    jdff dff_B_sThnjLOW4_2(.din(n10258), .dout(n10261));
    jdff dff_B_2jMqZwdh5_2(.din(n10261), .dout(n10264));
    jdff dff_B_kyfv9RBk3_0(.din(n5148), .dout(n10267));
    jdff dff_B_qMcc0HEP6_0(.din(n10267), .dout(n10270));
    jdff dff_B_YLdHd6tD0_0(.din(n10270), .dout(n10273));
    jdff dff_B_9YfKdWK08_1(.din(n5057), .dout(n10276));
    jdff dff_B_UQKYH9Ol9_1(.din(n10276), .dout(n10279));
    jdff dff_B_zccf1NQR1_1(.din(n10279), .dout(n10282));
    jdff dff_B_DsDLv6TT5_1(.din(n10282), .dout(n10285));
    jdff dff_B_Kf49E3wu8_1(.din(n10285), .dout(n10288));
    jdff dff_B_XjMt2yO34_1(.din(n10288), .dout(n10291));
    jdff dff_B_SySFhhGT3_1(.din(n10291), .dout(n10294));
    jdff dff_B_cNLpmMdh9_1(.din(n10294), .dout(n10297));
    jdff dff_B_MGzbcxmn3_1(.din(n10297), .dout(n10300));
    jdff dff_B_JUnEuirv2_1(.din(n10300), .dout(n10303));
    jdff dff_B_BhTQqvKk4_1(.din(n10303), .dout(n10306));
    jdff dff_B_OKiIDr9X6_1(.din(n10306), .dout(n10309));
    jdff dff_B_2O444AIl1_1(.din(n10309), .dout(n10312));
    jdff dff_B_EsPNKSXH3_1(.din(n10312), .dout(n10315));
    jdff dff_B_p4HONLhX2_1(.din(n10315), .dout(n10318));
    jdff dff_B_x2kVBAV96_1(.din(n10318), .dout(n10321));
    jdff dff_B_8qb9JnrM6_1(.din(n10321), .dout(n10324));
    jdff dff_B_bVCbw5jP6_0(.din(n5136), .dout(n10327));
    jdff dff_B_7FIOKbKe8_0(.din(n10327), .dout(n10330));
    jdff dff_B_9zCOOAxD2_0(.din(n5124), .dout(n10333));
    jdff dff_B_92bLwit86_0(.din(n10333), .dout(n10336));
    jdff dff_B_1nNq9ubr4_0(.din(n10336), .dout(n10339));
    jdff dff_B_WYKqQNdS8_0(.din(n10339), .dout(n10342));
    jdff dff_B_jgRtkKpr3_0(.din(n10342), .dout(n10345));
    jdff dff_B_E5nqfP4x2_0(.din(n10345), .dout(n10348));
    jdff dff_B_F2TP6eVx6_1(.din(n5101), .dout(n10351));
    jdff dff_B_cPEWPHhX5_1(.din(n10351), .dout(n10354));
    jdff dff_B_AQXSGaOY9_1(.din(n10354), .dout(n10357));
    jdff dff_B_Jdd7TguC6_0(.din(n5108), .dout(n10360));
    jdff dff_B_AsBXhVOA6_0(.din(n5093), .dout(n10363));
    jdff dff_B_gtqeDLaA1_0(.din(n10363), .dout(n10366));
    jdff dff_B_qUMsoeRw8_0(.din(n5085), .dout(n10369));
    jdff dff_B_54ePHx2p1_0(.din(n10369), .dout(n10372));
    jdff dff_B_VuDupfmp4_0(.din(n10372), .dout(n10375));
    jdff dff_B_UXMno1W47_0(.din(n10375), .dout(n10378));
    jdff dff_B_eqgWUqGr2_0(.din(n10378), .dout(n10381));
    jdff dff_B_d7qp4tb85_0(.din(n10381), .dout(n10384));
    jdff dff_B_11Q2SXGH8_0(.din(n5081), .dout(n10387));
    jdff dff_B_g6FwZoqP4_0(.din(n10387), .dout(n10390));
    jdff dff_B_oJAojJul3_0(.din(n10390), .dout(n10393));
    jdff dff_B_7T2CMOVL2_0(.din(n10393), .dout(n10396));
    jdff dff_B_qqXNUt202_0(.din(n10396), .dout(n10399));
    jdff dff_B_ESh5Qf9G8_0(.din(n5077), .dout(n10402));
    jdff dff_B_zxuyijCv3_0(.din(n10402), .dout(n10405));
    jdff dff_B_XZZm6ftf0_0(.din(n5061), .dout(n10408));
    jdff dff_A_PXGPS2LS4_1(.din(n10413), .dout(n10410));
    jdff dff_A_1W9ogM5S2_1(.din(n10416), .dout(n10413));
    jdff dff_A_YAhy02zL6_1(.din(n10419), .dout(n10416));
    jdff dff_A_hJn7yT7j7_1(.din(n10477), .dout(n10419));
    jdff dff_A_KuhxwjDN7_2(.din(n10425), .dout(n10422));
    jdff dff_A_9B3hDVd52_2(.din(n10428), .dout(n10425));
    jdff dff_A_VRs2VgW55_2(.din(n10431), .dout(n10428));
    jdff dff_A_uEyEvH4i8_2(.din(n10434), .dout(n10431));
    jdff dff_A_mTIZ4Kb78_2(.din(n10437), .dout(n10434));
    jdff dff_A_TwBweXs65_2(.din(n10440), .dout(n10437));
    jdff dff_A_yFR6T61W9_2(.din(n10443), .dout(n10440));
    jdff dff_A_LOyNwaeG2_2(.din(n10446), .dout(n10443));
    jdff dff_A_0VUNrvOx1_2(.din(n10449), .dout(n10446));
    jdff dff_A_K9bwiR2B9_2(.din(n10452), .dout(n10449));
    jdff dff_A_o0RjupcQ4_2(.din(n10455), .dout(n10452));
    jdff dff_A_5Ppzryr87_2(.din(n10458), .dout(n10455));
    jdff dff_A_D2lhm79R9_2(.din(n10461), .dout(n10458));
    jdff dff_A_whQeeJ9W9_2(.din(n10464), .dout(n10461));
    jdff dff_A_LDUmc2re1_2(.din(n10467), .dout(n10464));
    jdff dff_A_t7v2Foso9_2(.din(n10477), .dout(n10467));
    jdff dff_B_riTkMIhQ1_3(.din(n4519), .dout(n10471));
    jdff dff_B_BA6ypliL0_3(.din(n10471), .dout(n10474));
    jdff dff_B_prn8QpJd1_3(.din(n10474), .dout(n10477));
    jdff dff_B_uP0Es38F6_0(.din(n5049), .dout(n10480));
    jdff dff_B_ySHsmOrS1_0(.din(n10480), .dout(n10483));
    jdff dff_B_p8TN8DnC6_0(.din(n10483), .dout(n10486));
    jdff dff_B_PI4UAjCe7_0(.din(n10486), .dout(n10489));
    jdff dff_B_ULeS2Hdb5_0(.din(n5045), .dout(n10492));
    jdff dff_B_8MufqKta2_0(.din(n10492), .dout(n10495));
    jdff dff_B_BFXyUr5n4_0(.din(n10495), .dout(n10498));
    jdff dff_B_xS7EoXhY9_0(.din(n10498), .dout(n10501));
    jdff dff_B_M7sTA4wo4_0(.din(n5037), .dout(n10504));
    jdff dff_B_WMdstgmH6_0(.din(n5029), .dout(n10507));
    jdff dff_B_dQ2XVzZb1_0(.din(n10507), .dout(n10510));
    jdff dff_B_pBDQt7Fm1_0(.din(n10510), .dout(n10513));
    jdff dff_A_hYRC2GmT0_1(.din(n10518), .dout(n10515));
    jdff dff_A_ETdLGiEY0_1(.din(n10521), .dout(n10518));
    jdff dff_A_csLbnYY68_1(.din(n10524), .dout(n10521));
    jdff dff_A_KbhxKYfc1_1(.din(n10527), .dout(n10524));
    jdff dff_A_KIdcbo8U6_1(.din(n10530), .dout(n10527));
    jdff dff_A_cIAROaMX8_1(.din(n10533), .dout(n10530));
    jdff dff_A_ykPomkwX5_1(.din(n10570), .dout(n10533));
    jdff dff_B_wrLotaPu8_2(.din(n4683), .dout(n10537));
    jdff dff_B_qlpbRo6X8_2(.din(n10537), .dout(n10540));
    jdff dff_B_OslxSPui1_2(.din(n10540), .dout(n10543));
    jdff dff_B_LMZAH95D2_2(.din(n10543), .dout(n10546));
    jdff dff_B_W7sI2l7y4_2(.din(n10546), .dout(n10549));
    jdff dff_B_jY4d4e6v0_2(.din(n10549), .dout(n10552));
    jdff dff_B_xfjsJTi02_2(.din(n10552), .dout(n10555));
    jdff dff_B_MZyPwBM32_2(.din(n10555), .dout(n10558));
    jdff dff_B_XHc56SKP0_2(.din(n10558), .dout(n10561));
    jdff dff_B_ixzvRv4d5_2(.din(n10561), .dout(n10564));
    jdff dff_B_Ue1tB1dW8_2(.din(n10564), .dout(n10567));
    jdff dff_B_2rNbrDSn7_2(.din(n10567), .dout(n10570));
    jdff dff_B_HuXvoX1q7_0(.din(n4410), .dout(n10573));
    jdff dff_B_wIXhcqSn5_0(.din(n10573), .dout(n10576));
    jdff dff_B_AnSrUlyW8_0(.din(n10576), .dout(n10579));
    jdff dff_B_oUAMA5Bw9_0(.din(n10579), .dout(n10582));
    jdff dff_B_blBRfFA76_0(.din(n10582), .dout(n10585));
    jdff dff_B_RVNBsr5A7_0(.din(n10585), .dout(n10588));
    jdff dff_B_Feo5D2xO0_0(.din(n10588), .dout(n10591));
    jdff dff_B_vdXXe8U12_0(.din(n10591), .dout(n10594));
    jdff dff_B_mecUcKPL7_0(.din(n4399), .dout(n10597));
    jdff dff_B_6JClkLPU5_0(.din(n10597), .dout(n10600));
    jdff dff_B_iot4Zr9i4_0(.din(n10600), .dout(n10603));
    jdff dff_B_o9eZOgmS1_0(.din(n10603), .dout(n10606));
    jdff dff_B_GIOaFgy69_3(.din(n1799), .dout(n10609));
    jdff dff_B_AthcAGN26_3(.din(n10609), .dout(n10612));
    jdff dff_B_02lejIxl3_3(.din(n10612), .dout(n10615));
    jdff dff_B_Xp3YSTii9_3(.din(n10615), .dout(n10618));
    jdff dff_B_WHQ1Ggsp6_3(.din(n10618), .dout(n10621));
    jdff dff_B_CsnQHbpm0_3(.din(n10621), .dout(n10624));
    jdff dff_B_lLWNjJ9j3_3(.din(n10624), .dout(n10627));
    jdff dff_B_y3fjucnV8_3(.din(n10627), .dout(n10630));
    jdff dff_B_qJra4Pqc5_3(.din(n10630), .dout(n10633));
    jdff dff_B_l1SLN5z83_3(.din(n10633), .dout(n10636));
    jdff dff_B_vBcehRgJ4_3(.din(n10636), .dout(n10639));
    jdff dff_B_syuzaC8i3_3(.din(n10639), .dout(n10642));
    jdff dff_B_xWHdXOLP2_3(.din(n10642), .dout(n10645));
    jdff dff_B_fQZma7k94_3(.din(n10645), .dout(n10648));
    jdff dff_B_nKlIzAtF4_3(.din(n10648), .dout(n10651));
    jdff dff_B_fiaUomy91_3(.din(n10651), .dout(n10654));
    jdff dff_B_1rzDFzsj1_3(.din(n10654), .dout(n10657));
    jdff dff_B_wcNfDzhL9_3(.din(n10657), .dout(n10660));
    jdff dff_B_FivChyJd2_3(.din(n10660), .dout(n10663));
    jdff dff_A_2pLA6sGi2_0(.din(n10668), .dout(n10665));
    jdff dff_A_IScrSnDp4_0(.din(n10671), .dout(n10668));
    jdff dff_A_RIj09X6r4_0(.din(n10674), .dout(n10671));
    jdff dff_A_5miIlYs52_0(.din(n10677), .dout(n10674));
    jdff dff_A_8S2mVXtp5_0(.din(n10680), .dout(n10677));
    jdff dff_A_bVnIap0S4_0(.din(n10683), .dout(n10680));
    jdff dff_A_RUIAskX05_0(.din(n10686), .dout(n10683));
    jdff dff_A_bqr44H7R8_0(.din(n10689), .dout(n10686));
    jdff dff_A_s2bnclLQ6_0(.din(n10692), .dout(n10689));
    jdff dff_A_NKs9K9fI5_0(.din(n10695), .dout(n10692));
    jdff dff_A_rVwvjIRN8_0(.din(n10698), .dout(n10695));
    jdff dff_A_TEOTdLan2_0(.din(n10701), .dout(n10698));
    jdff dff_A_4pEt9iRe8_0(.din(n10704), .dout(n10701));
    jdff dff_A_2fsMJv6Z9_0(.din(n1796), .dout(n10704));
    jdff dff_A_rYs4GucR6_1(.din(n10710), .dout(n10707));
    jdff dff_A_DSUFAiTB4_1(.din(n10713), .dout(n10710));
    jdff dff_A_AAIVqFnq0_1(.din(n10716), .dout(n10713));
    jdff dff_A_aKdzrLD49_1(.din(n10719), .dout(n10716));
    jdff dff_A_93P75Fw56_1(.din(n1781), .dout(n10719));
    jdff dff_A_63JeO8yX5_1(.din(n10725), .dout(n10722));
    jdff dff_A_RToS7jYS6_1(.din(n10728), .dout(n10725));
    jdff dff_A_0N8FCyks1_1(.din(n10731), .dout(n10728));
    jdff dff_A_6EiRPQPw6_1(.din(n10734), .dout(n10731));
    jdff dff_A_DUwVtVMp5_1(.din(n1778), .dout(n10734));
    jdff dff_B_5GJbIelO2_1(.din(n1693), .dout(n10738));
    jdff dff_B_6QqI81sW6_1(.din(n10738), .dout(n10741));
    jdff dff_B_31axOZ779_1(.din(n10741), .dout(n10744));
    jdff dff_B_WcgBQG6L5_1(.din(n10744), .dout(n10747));
    jdff dff_B_AW24cn5E4_1(.din(n10747), .dout(n10750));
    jdff dff_B_98DFixQV3_1(.din(n10750), .dout(n10753));
    jdff dff_B_6CyJdoem4_1(.din(n10753), .dout(n10756));
    jdff dff_B_j5sFEgj30_1(.din(n10756), .dout(n10759));
    jdff dff_B_nBGwLroT7_1(.din(n10759), .dout(n10762));
    jdff dff_B_dBcfTNrF6_1(.din(n10762), .dout(n10765));
    jdff dff_B_QSBeyMPl2_1(.din(n1697), .dout(n10768));
    jdff dff_B_31TRHZrU5_1(.din(n10768), .dout(n10771));
    jdff dff_B_j117HOou5_1(.din(n10771), .dout(n10774));
    jdff dff_B_nAACLr1z2_1(.din(n10774), .dout(n10777));
    jdff dff_B_DQ1EHF7V3_1(.din(n10777), .dout(n10780));
    jdff dff_B_xJnr10EK2_1(.din(n10780), .dout(n10783));
    jdff dff_B_qnY7mpwh9_1(.din(n10783), .dout(n10786));
    jdff dff_B_CrkyE9VK5_1(.din(n10786), .dout(n10789));
    jdff dff_B_R8R1GegZ9_1(.din(n10789), .dout(n10792));
    jdff dff_A_b3NQQGGA8_0(.din(n10797), .dout(n10794));
    jdff dff_A_QP6gin3t0_0(.din(n10800), .dout(n10797));
    jdff dff_A_Cy4gb3jU5_0(.din(n10803), .dout(n10800));
    jdff dff_A_XtNZ2cwT4_0(.din(n10806), .dout(n10803));
    jdff dff_A_uztjHBXS0_0(.din(n10809), .dout(n10806));
    jdff dff_A_AFbJ8nJ87_0(.din(n10812), .dout(n10809));
    jdff dff_A_F2FgUrfK6_0(.din(n10815), .dout(n10812));
    jdff dff_A_0ehuDGa37_0(.din(n10818), .dout(n10815));
    jdff dff_A_geo1gBGY6_0(.din(n10821), .dout(n10818));
    jdff dff_A_QVllah6X5_0(.din(n10824), .dout(n10821));
    jdff dff_A_W7cqJDbd8_0(.din(n1767), .dout(n10824));
    jdff dff_B_mMspoOhi8_1(.din(n1708), .dout(n10828));
    jdff dff_B_SbXtGPCx1_1(.din(n10828), .dout(n10831));
    jdff dff_B_3RZrnDtC6_1(.din(n10831), .dout(n10834));
    jdff dff_B_k26eojcT9_1(.din(n10834), .dout(n10837));
    jdff dff_B_eirtcAzx3_1(.din(n10837), .dout(n10840));
    jdff dff_B_USI1XqZs9_1(.din(n1712), .dout(n10843));
    jdff dff_B_lbDXiSBl2_1(.din(n10843), .dout(n10846));
    jdff dff_B_c7vP74jz2_1(.din(n10846), .dout(n10849));
    jdff dff_B_fuS5g3We1_1(.din(n10849), .dout(n10852));
    jdff dff_B_ZrU08K1A0_0(.din(n1744), .dout(n10855));
    jdff dff_A_pDvDnkNp0_0(.din(n10860), .dout(n10857));
    jdff dff_A_VHmyh0658_0(.din(n10863), .dout(n10860));
    jdff dff_A_llREnJMm9_0(.din(n10866), .dout(n10863));
    jdff dff_A_5plgl53j5_0(.din(n10869), .dout(n10866));
    jdff dff_A_FUNQwxCo7_0(.din(n10872), .dout(n10869));
    jdff dff_A_rFRXfMHw8_0(.din(n10875), .dout(n10872));
    jdff dff_A_Heppkal78_0(.din(n10878), .dout(n10875));
    jdff dff_A_S98k5jCQ7_0(.din(n10881), .dout(n10878));
    jdff dff_A_yGyzPe4B2_0(.din(n10884), .dout(n10881));
    jdff dff_A_7FMjB3Vu6_0(.din(n10887), .dout(n10884));
    jdff dff_A_63wWsD236_0(.din(n10890), .dout(n10887));
    jdff dff_A_VnPbcDzP7_0(.din(n1740), .dout(n10890));
    jdff dff_A_u7F2Q8m55_1(.din(n10896), .dout(n10893));
    jdff dff_A_OXz8K64H4_1(.din(n10899), .dout(n10896));
    jdff dff_A_h6WxvGi87_1(.din(n10902), .dout(n10899));
    jdff dff_A_N1hFQIAX4_1(.din(n10905), .dout(n10902));
    jdff dff_A_kqHA7SEI9_1(.din(n10908), .dout(n10905));
    jdff dff_A_OHcH1tg02_1(.din(n10911), .dout(n10908));
    jdff dff_A_pIWS2X621_1(.din(n10914), .dout(n10911));
    jdff dff_A_Cy9aYAbq4_1(.din(n10917), .dout(n10914));
    jdff dff_A_fSmbRiGw6_1(.din(n10920), .dout(n10917));
    jdff dff_A_ntRiys6G6_1(.din(n10923), .dout(n10920));
    jdff dff_A_GtSFQ6Iu6_1(.din(n10926), .dout(n10923));
    jdff dff_A_NxWtbGzu4_1(.din(n10929), .dout(n10926));
    jdff dff_A_h48hVY0p1_1(.din(n10932), .dout(n10929));
    jdff dff_A_39wYxN6T5_1(.din(n10935), .dout(n10932));
    jdff dff_A_ywic1fHk4_1(.din(n10938), .dout(n10935));
    jdff dff_A_ohcuHZ8E6_1(.din(n10941), .dout(n10938));
    jdff dff_A_T8J0NI7b7_1(.din(n1740), .dout(n10941));
    jdff dff_A_N0r6384D1_1(.din(n1722), .dout(n10944));
    jdff dff_A_1IQtyevN2_1(.din(n10963), .dout(n10947));
    jdff dff_B_3CWIUYUh5_2(.din(n1704), .dout(n10951));
    jdff dff_B_ZSb2eyue1_2(.din(n10951), .dout(n10954));
    jdff dff_B_UEr6zIbv1_2(.din(n10954), .dout(n10957));
    jdff dff_B_JqLPROAF1_2(.din(n10957), .dout(n10960));
    jdff dff_B_FRjIx0s29_2(.din(n10960), .dout(n10963));
    jdff dff_A_0uQLXxFj7_0(.din(n10968), .dout(n10965));
    jdff dff_A_se3lgJdO6_0(.din(n10971), .dout(n10968));
    jdff dff_A_tw1W2qY31_0(.din(n10974), .dout(n10971));
    jdff dff_A_HijjC0fh7_0(.din(n10977), .dout(n10974));
    jdff dff_A_OzFdgeut2_0(.din(n1701), .dout(n10977));
    jdff dff_B_a6vI01Xa7_0(.din(n1685), .dout(n10981));
    jdff dff_B_PbVZSAaj7_0(.din(n10981), .dout(n10984));
    jdff dff_B_zoGqrCsr9_0(.din(n10984), .dout(n10987));
    jdff dff_B_8TrRRcVy0_0(.din(n10987), .dout(n10990));
    jdff dff_B_UD8zV4Fo8_0(.din(n10990), .dout(n10993));
    jdff dff_B_3vhR5FRd5_0(.din(n10993), .dout(n10996));
    jdff dff_B_egxG1bLp0_0(.din(n10996), .dout(n10999));
    jdff dff_B_wzsIbGOs3_0(.din(n10999), .dout(n11002));
    jdff dff_B_M597tXan2_0(.din(n11002), .dout(n11005));
    jdff dff_B_oSwk6T4H0_0(.din(n11005), .dout(n11008));
    jdff dff_B_lbYoKhjc4_0(.din(n11008), .dout(n11011));
    jdff dff_B_v6k1PaaS2_0(.din(n11011), .dout(n11014));
    jdff dff_A_nRk0F1yu3_0(.din(n11019), .dout(n11016));
    jdff dff_A_9F0lqJYL3_0(.din(n11022), .dout(n11019));
    jdff dff_A_ahdHbyKk0_0(.din(n11025), .dout(n11022));
    jdff dff_A_BsN9hC1e8_0(.din(n11028), .dout(n11025));
    jdff dff_A_bmHVwHPA3_0(.din(n1678), .dout(n11028));
    jdff dff_A_8v14q7Rr6_1(.din(n11034), .dout(n11031));
    jdff dff_A_bxt3cWg04_1(.din(n1674), .dout(n11034));
    jdff dff_A_ROvKrg5y1_2(.din(n1674), .dout(n11037));
    jdff dff_A_IUaQs51h2_0(.din(n11043), .dout(n11040));
    jdff dff_A_RQV5umD88_0(.din(n11046), .dout(n11043));
    jdff dff_A_DZvNQCFr8_0(.din(n11049), .dout(n11046));
    jdff dff_A_Efe0r4uT8_0(.din(n11052), .dout(n11049));
    jdff dff_A_BOeQg6d50_0(.din(n11055), .dout(n11052));
    jdff dff_A_mcxyT3IL0_0(.din(n11058), .dout(n11055));
    jdff dff_A_83idBDcV2_0(.din(n11061), .dout(n11058));
    jdff dff_A_1SOOwDKX2_0(.din(n11064), .dout(n11061));
    jdff dff_A_GfgfAQdm0_0(.din(n11067), .dout(n11064));
    jdff dff_A_qN9E9QMu1_0(.din(n11070), .dout(n11067));
    jdff dff_A_SZwoJk737_0(.din(n11073), .dout(n11070));
    jdff dff_A_FoAN2lGm2_0(.din(n11076), .dout(n11073));
    jdff dff_A_U9khHxe71_0(.din(n11079), .dout(n11076));
    jdff dff_A_LOgY3SDJ6_0(.din(n11082), .dout(n11079));
    jdff dff_A_24HZQlwX4_0(.din(n11085), .dout(n11082));
    jdff dff_A_Hk3heCbt6_0(.din(n1670), .dout(n11085));
    jdff dff_A_dy8idU0p2_1(.din(n11091), .dout(n11088));
    jdff dff_A_0k3ywTYN8_1(.din(n11094), .dout(n11091));
    jdff dff_A_FfUNx92S1_1(.din(n11097), .dout(n11094));
    jdff dff_A_xeqNNqnp7_1(.din(n11100), .dout(n11097));
    jdff dff_A_uhzyLWyT7_1(.din(n11103), .dout(n11100));
    jdff dff_A_yI1dmKmU2_1(.din(n11106), .dout(n11103));
    jdff dff_A_7ed9KzhY5_1(.din(n11109), .dout(n11106));
    jdff dff_A_g9dXKNb59_1(.din(n11112), .dout(n11109));
    jdff dff_A_fivInbil4_1(.din(n11115), .dout(n11112));
    jdff dff_A_TuC4Q1IY3_1(.din(n11118), .dout(n11115));
    jdff dff_A_zHTplkiB0_1(.din(n11121), .dout(n11118));
    jdff dff_A_HCOkP9kF2_1(.din(n11124), .dout(n11121));
    jdff dff_A_pFcKP18F0_1(.din(n11127), .dout(n11124));
    jdff dff_A_aQekNMNG6_1(.din(n11130), .dout(n11127));
    jdff dff_A_BrggSZaM2_1(.din(n11133), .dout(n11130));
    jdff dff_A_ksJ7tGhk9_1(.din(n1670), .dout(n11133));
    jdff dff_B_ntO3dZxz6_0(.din(G209), .dout(n11137));
    jdff dff_B_Eb137lpD7_3(.din(n1658), .dout(n11140));
    jdff dff_B_1b42s4Cf3_3(.din(n11140), .dout(n11143));
    jdff dff_A_FXzQTZBz9_0(.din(n11148), .dout(n11145));
    jdff dff_A_W3wYQSli9_0(.din(n11151), .dout(n11148));
    jdff dff_A_JXQWSPKi0_0(.din(n11154), .dout(n11151));
    jdff dff_A_Vtxl6EgM4_0(.din(n11157), .dout(n11154));
    jdff dff_A_IS4t9m6n0_0(.din(n11160), .dout(n11157));
    jdff dff_A_qnmJzlNA5_0(.din(n11163), .dout(n11160));
    jdff dff_A_traQn1J99_0(.din(n11166), .dout(n11163));
    jdff dff_A_0KY4L7qb6_0(.din(n11169), .dout(n11166));
    jdff dff_A_cLN2eEGx0_0(.din(n11172), .dout(n11169));
    jdff dff_A_J3qQsUsv8_0(.din(n11175), .dout(n11172));
    jdff dff_A_hpwijWbA4_0(.din(n11178), .dout(n11175));
    jdff dff_A_w8FTFYUL0_0(.din(n11181), .dout(n11178));
    jdff dff_A_6Hl9xR1E1_0(.din(n11184), .dout(n11181));
    jdff dff_A_jPop937a0_0(.din(n11187), .dout(n11184));
    jdff dff_A_csVXd10E6_0(.din(n11190), .dout(n11187));
    jdff dff_A_m1C0VH770_0(.din(n11193), .dout(n11190));
    jdff dff_A_CIVjT5VM8_0(.din(n11196), .dout(n11193));
    jdff dff_A_v7RfquDs0_0(.din(n1655), .dout(n11196));
    jdff dff_A_QUy4eyxe1_1(.din(n11202), .dout(n11199));
    jdff dff_A_phBDlMg71_1(.din(n11205), .dout(n11202));
    jdff dff_A_fIC2p0Xx1_1(.din(n11208), .dout(n11205));
    jdff dff_A_uCNOdBRd7_1(.din(n11211), .dout(n11208));
    jdff dff_A_A0vxmUpU9_1(.din(n11214), .dout(n11211));
    jdff dff_A_TxJfzI5u1_1(.din(n11217), .dout(n11214));
    jdff dff_A_9Q4iBcA39_1(.din(n11220), .dout(n11217));
    jdff dff_A_OKZphSOh1_1(.din(n11223), .dout(n11220));
    jdff dff_A_pVVPqvYX2_1(.din(n11226), .dout(n11223));
    jdff dff_A_QZfrvL4I7_1(.din(n11229), .dout(n11226));
    jdff dff_A_8O7LrDql9_1(.din(n11232), .dout(n11229));
    jdff dff_A_FhDUAYYh0_1(.din(n11235), .dout(n11232));
    jdff dff_A_mzieiADk9_1(.din(n1655), .dout(n11235));
    jdff dff_A_ohXg0I1s7_0(.din(n11241), .dout(n11238));
    jdff dff_A_1aqJqf1o2_0(.din(n1647), .dout(n11241));
    jdff dff_B_k0FUDk4O7_0(.din(G216), .dout(n11245));
    jdff dff_B_UFEOpjR45_2(.din(n1643), .dout(n11248));
    jdff dff_B_xfvM5hH19_2(.din(n11248), .dout(n11251));
    jdff dff_A_D4pDAyua3_0(.din(n11256), .dout(n11253));
    jdff dff_A_dA0aAkgi9_0(.din(n11259), .dout(n11256));
    jdff dff_A_66mRX9688_0(.din(n11262), .dout(n11259));
    jdff dff_A_6HCsU9672_0(.din(G1469), .dout(n11262));
    jdff dff_A_iVqUbNYz1_0(.din(n11268), .dout(n11265));
    jdff dff_A_Rt6Qggwj7_0(.din(n1628), .dout(n11268));
    jdff dff_B_XHcYUwEC3_0(.din(G215), .dout(n11272));
    jdff dff_B_ZdNvDYb41_2(.din(n1624), .dout(n11275));
    jdff dff_B_xceFMOFW7_2(.din(n11275), .dout(n11278));
    jdff dff_A_IuovkDfs4_0(.din(n11283), .dout(n11280));
    jdff dff_A_A3N2WasT5_0(.din(n11286), .dout(n11283));
    jdff dff_A_v0z01ZgM1_0(.din(n11289), .dout(n11286));
    jdff dff_A_pPlrvx5T9_0(.din(G106), .dout(n11289));
    jdff dff_B_n7oZ3W448_0(.din(G214), .dout(n11293));
    jdff dff_B_rNlhbg6w2_3(.din(n1609), .dout(n11296));
    jdff dff_B_pmxFTMoD6_3(.din(n11296), .dout(n11299));
    jdff dff_A_N0kDuRwy6_1(.din(n11304), .dout(n11301));
    jdff dff_A_Ivn3BrT31_1(.din(n1606), .dout(n11304));
    jdff dff_B_tR2LbQ4n4_0(.din(G213), .dout(n11308));
    jdff dff_B_z6Iml3TC6_3(.din(n1594), .dout(n11311));
    jdff dff_B_VXaHy9Hx2_3(.din(n11311), .dout(n11314));
    jdff dff_A_LhYOVxyI5_1(.din(n11319), .dout(n11316));
    jdff dff_A_Ug3mK5NG0_1(.din(n11322), .dout(n11319));
    jdff dff_A_7wd10qIo0_1(.din(n11325), .dout(n11322));
    jdff dff_A_EAb3kC1d5_1(.din(n11328), .dout(n11325));
    jdff dff_A_MAQeO5oo4_1(.din(n11331), .dout(n11328));
    jdff dff_A_B6LaQCym1_1(.din(n11334), .dout(n11331));
    jdff dff_A_mRWBJonj2_1(.din(n11337), .dout(n11334));
    jdff dff_A_15KflhwZ3_1(.din(n11340), .dout(n11337));
    jdff dff_A_HSuaGMv20_1(.din(n1587), .dout(n11340));
    jdff dff_B_fVfsT3JD2_1(.din(n1531), .dout(n11344));
    jdff dff_B_Mkxo0zjz7_1(.din(n11344), .dout(n11347));
    jdff dff_B_Z7mHQ0hz1_1(.din(n11347), .dout(n11350));
    jdff dff_B_M9KreNBI5_1(.din(n11350), .dout(n11353));
    jdff dff_B_hAhFDvod4_0(.din(n1579), .dout(n11356));
    jdff dff_B_QRx72X1R3_0(.din(n11356), .dout(n11359));
    jdff dff_A_nx74sppU0_0(.din(n11364), .dout(n11361));
    jdff dff_A_pLdcDt4v1_0(.din(n11367), .dout(n11364));
    jdff dff_A_UmgNyxXY9_0(.din(n11370), .dout(n11367));
    jdff dff_A_whLRc9xJ3_0(.din(n11373), .dout(n11370));
    jdff dff_A_mdlHZwOP4_0(.din(n11376), .dout(n11373));
    jdff dff_A_1lprh0ls4_0(.din(n11379), .dout(n11376));
    jdff dff_A_afMyLor28_0(.din(n11382), .dout(n11379));
    jdff dff_A_vQHn923G0_0(.din(n11385), .dout(n11382));
    jdff dff_A_H5ozfvEf8_0(.din(n11388), .dout(n11385));
    jdff dff_A_Bn4mYZrY0_0(.din(n11391), .dout(n11388));
    jdff dff_A_1fPSTm731_0(.din(n11394), .dout(n11391));
    jdff dff_A_hPBh4mk55_0(.din(n11397), .dout(n11394));
    jdff dff_A_LAnBHev18_0(.din(n11400), .dout(n11397));
    jdff dff_A_N85r8T5u6_0(.din(n11403), .dout(n11400));
    jdff dff_A_bYH1Yk4w1_0(.din(n1575), .dout(n11403));
    jdff dff_A_piWLtxRU3_1(.din(n11409), .dout(n11406));
    jdff dff_A_wne7cskn8_1(.din(n11412), .dout(n11409));
    jdff dff_A_sUtFUMxE0_1(.din(n1575), .dout(n11412));
    jdff dff_A_mni2gDwA4_1(.din(n11418), .dout(n11415));
    jdff dff_A_9qscZx968_1(.din(n11421), .dout(n11418));
    jdff dff_A_DOr04mro5_1(.din(n11424), .dout(n11421));
    jdff dff_A_VTSm0hsC0_1(.din(n11427), .dout(n11424));
    jdff dff_A_ZCxDpFtE6_1(.din(n11430), .dout(n11427));
    jdff dff_A_ucRnVag98_1(.din(n11433), .dout(n11430));
    jdff dff_A_0EK1odHV0_1(.din(n11436), .dout(n11433));
    jdff dff_A_PMyYqndW8_1(.din(n11439), .dout(n11436));
    jdff dff_A_DB7tKIUf7_1(.din(n11442), .dout(n11439));
    jdff dff_A_YR6YSlRF7_1(.din(n11445), .dout(n11442));
    jdff dff_A_IpbrTOhL4_1(.din(n11448), .dout(n11445));
    jdff dff_A_LnBaAuQd1_1(.din(n1557), .dout(n11448));
    jdff dff_B_C4tzDZ6m2_1(.din(n1542), .dout(n11452));
    jdff dff_A_NlXmhPtA6_0(.din(n1546), .dout(n11454));
    jdff dff_A_qb3jlVHQ1_1(.din(n11460), .dout(n11457));
    jdff dff_A_imvC1xlh9_1(.din(n11463), .dout(n11460));
    jdff dff_A_SlLxopcg6_1(.din(n11466), .dout(n11463));
    jdff dff_A_SntQfvgC6_1(.din(n11469), .dout(n11466));
    jdff dff_A_rORgkK0L6_1(.din(n11472), .dout(n11469));
    jdff dff_A_i8Ge2UoJ1_1(.din(n11475), .dout(n11472));
    jdff dff_A_xTDhwCkA7_1(.din(n11478), .dout(n11475));
    jdff dff_A_u1XntUmo6_1(.din(n11481), .dout(n11478));
    jdff dff_A_A3w1LbOh4_1(.din(n11484), .dout(n11481));
    jdff dff_A_hAcYqbdW5_1(.din(n11487), .dout(n11484));
    jdff dff_A_URvGaDG78_1(.din(n11490), .dout(n11487));
    jdff dff_A_o77milgf7_1(.din(n11493), .dout(n11490));
    jdff dff_A_UkMHL19G4_1(.din(n11496), .dout(n11493));
    jdff dff_A_TYce3fmA5_1(.din(n11499), .dout(n11496));
    jdff dff_A_xKhpYeJo3_1(.din(n1546), .dout(n11499));
    jdff dff_A_TF2dRplP6_0(.din(n11505), .dout(n11502));
    jdff dff_A_NSQ0FXRP2_0(.din(n11508), .dout(n11505));
    jdff dff_A_xjREGCon4_0(.din(n11511), .dout(n11508));
    jdff dff_A_gTFgY2Nd6_0(.din(n11514), .dout(n11511));
    jdff dff_A_YdIucaZ67_0(.din(n11517), .dout(n11514));
    jdff dff_A_WVB6Expa2_0(.din(n11520), .dout(n11517));
    jdff dff_A_b9qFrL5p4_0(.din(n11523), .dout(n11520));
    jdff dff_A_kZNUPEa16_0(.din(n11526), .dout(n11523));
    jdff dff_A_UzbzHfDK9_0(.din(n11529), .dout(n11526));
    jdff dff_A_bO5DoJI41_0(.din(n11532), .dout(n11529));
    jdff dff_A_BhdhF3A34_0(.din(n11535), .dout(n11532));
    jdff dff_A_H378nXVf0_0(.din(n11538), .dout(n11535));
    jdff dff_A_xApNFDDi8_0(.din(n11541), .dout(n11538));
    jdff dff_A_htWSNZ0U3_0(.din(n11548), .dout(n11541));
    jdff dff_B_8bzvD6Xj6_2(.din(n1538), .dout(n11545));
    jdff dff_B_64BnYiHV3_2(.din(n11545), .dout(n11548));
    jdff dff_A_kTkwB2Kb6_0(.din(n11553), .dout(n11550));
    jdff dff_A_g5E6Xoil8_0(.din(n11556), .dout(n11553));
    jdff dff_A_PxZd0RBT7_0(.din(n11559), .dout(n11556));
    jdff dff_A_e1l956lS8_0(.din(n11562), .dout(n11559));
    jdff dff_A_8nXhsAqp5_0(.din(n1535), .dout(n11562));
    jdff dff_B_ePSTFwxn2_0(.din(n1520), .dout(n11566));
    jdff dff_B_dZZlInJA2_0(.din(n11566), .dout(n11569));
    jdff dff_B_5FdAPyX25_0(.din(n11569), .dout(n11572));
    jdff dff_B_yE7AFs3X2_0(.din(n11572), .dout(n11575));
    jdff dff_B_P4AxfDd10_0(.din(n11575), .dout(n11578));
    jdff dff_B_2dTI95Ag6_0(.din(n11578), .dout(n11581));
    jdff dff_B_GJhZjZyj5_0(.din(n11581), .dout(n11584));
    jdff dff_B_GF1bxYkC6_0(.din(n11584), .dout(n11587));
    jdff dff_B_cDhyUstl7_0(.din(n11587), .dout(n11590));
    jdff dff_B_hyaXkRZh4_0(.din(n11590), .dout(n11593));
    jdff dff_B_5bVHzCoB6_0(.din(n11593), .dout(n11596));
    jdff dff_A_dI8kEoUQ0_0(.din(n11601), .dout(n11598));
    jdff dff_A_v283yLyc2_0(.din(n11604), .dout(n11601));
    jdff dff_A_9CzZbaMW0_0(.din(n11607), .dout(n11604));
    jdff dff_A_PTXyHzPb2_0(.din(n11610), .dout(n11607));
    jdff dff_A_7yrQxVyh3_0(.din(n11613), .dout(n11610));
    jdff dff_A_hXgRrwjt0_0(.din(n11616), .dout(n11613));
    jdff dff_A_mQ7JHL7A0_0(.din(n11619), .dout(n11616));
    jdff dff_A_jJWjSZLk1_0(.din(n11622), .dout(n11619));
    jdff dff_A_tGKiAFJ45_0(.din(n11625), .dout(n11622));
    jdff dff_A_OAwK0ZCv7_0(.din(n11628), .dout(n11625));
    jdff dff_A_GJ4scgZd6_0(.din(n11631), .dout(n11628));
    jdff dff_A_YBLe62Qq7_0(.din(n1517), .dout(n11631));
    jdff dff_A_U3iOSSB60_0(.din(n1509), .dout(n11634));
    jdff dff_A_BhhxFeUR3_0(.din(n11640), .dout(n11637));
    jdff dff_A_z6Z7PJLr0_0(.din(n1501), .dout(n11640));
    jdff dff_B_gmR2tVV00_0(.din(G154), .dout(n11644));
    jdff dff_B_Wun7VePb7_2(.din(n1497), .dout(n11647));
    jdff dff_B_TLKxVHrz8_2(.din(n11647), .dout(n11650));
    jdff dff_A_5KOVEoVw7_0(.din(n11655), .dout(n11652));
    jdff dff_A_ZMWNQO8U4_0(.din(n11658), .dout(n11655));
    jdff dff_A_MwA18U3m5_0(.din(n11661), .dout(n11658));
    jdff dff_A_9uuk3uJU2_0(.din(G2253), .dout(n11661));
    jdff dff_A_PlpkORAv3_0(.din(n11667), .dout(n11664));
    jdff dff_A_EX3ZzQQk9_0(.din(n1486), .dout(n11667));
    jdff dff_B_9U7qMuqH0_0(.din(G153), .dout(n11671));
    jdff dff_B_wkLN8WmT3_2(.din(n1482), .dout(n11674));
    jdff dff_B_KqGlf3EU9_2(.din(n11674), .dout(n11677));
    jdff dff_A_H4W4do6z0_0(.din(n11682), .dout(n11679));
    jdff dff_A_oif6KGoZ0_0(.din(n11685), .dout(n11682));
    jdff dff_A_8cHYjrwL0_0(.din(n11688), .dout(n11685));
    jdff dff_A_Of6m4djP1_0(.din(G2256), .dout(n11688));
    jdff dff_A_s8YrdGsc3_0(.din(n11694), .dout(n11691));
    jdff dff_A_RnCEZq7s6_0(.din(n11697), .dout(n11694));
    jdff dff_A_tjQ9oybE9_0(.din(n11700), .dout(n11697));
    jdff dff_A_CWdmyTBg6_0(.din(n11703), .dout(n11700));
    jdff dff_A_xgzkMFPV2_0(.din(n11706), .dout(n11703));
    jdff dff_A_n6EGCexi3_0(.din(n11709), .dout(n11706));
    jdff dff_A_Lyuesbap7_0(.din(n11712), .dout(n11709));
    jdff dff_A_UaKZasdC2_0(.din(n11715), .dout(n11712));
    jdff dff_A_xVfsRKwD1_0(.din(n11718), .dout(n11715));
    jdff dff_A_I12FHI8l0_0(.din(n11721), .dout(n11718));
    jdff dff_A_NRpGR77t6_0(.din(n11724), .dout(n11721));
    jdff dff_A_kOdyl9j68_0(.din(n11727), .dout(n11724));
    jdff dff_A_YcCrtlXV4_0(.din(n11730), .dout(n11727));
    jdff dff_A_DqfIZIe95_0(.din(n1475), .dout(n11730));
    jdff dff_A_OnR7F0Ov0_0(.din(n11736), .dout(n11733));
    jdff dff_A_xUWqSw9H1_0(.din(n1467), .dout(n11736));
    jdff dff_B_q90zLv3b6_0(.din(G156), .dout(n11740));
    jdff dff_A_8IlHPIpi6_1(.din(n11745), .dout(n11742));
    jdff dff_A_hhuo9bPa3_1(.din(n1463), .dout(n11745));
    jdff dff_A_jOYC5UJN4_2(.din(n11751), .dout(n11748));
    jdff dff_A_82enB9Zl4_2(.din(n1463), .dout(n11751));
    jdff dff_A_K6kRUXt23_1(.din(n11757), .dout(n11754));
    jdff dff_A_lzE1Hsi35_1(.din(n11760), .dout(n11757));
    jdff dff_A_L8NjtLMm4_1(.din(n11763), .dout(n11760));
    jdff dff_A_mBJGbxOA3_1(.din(G2239), .dout(n11763));
    jdff dff_A_Jx6Nmo0H4_2(.din(n11769), .dout(n11766));
    jdff dff_A_Inpx9wdH7_2(.din(n11772), .dout(n11769));
    jdff dff_A_1sTzqk7F1_2(.din(n11775), .dout(n11772));
    jdff dff_A_n9sFzddv8_2(.din(n11778), .dout(n11775));
    jdff dff_A_5hBpT9Dg3_2(.din(n11781), .dout(n11778));
    jdff dff_A_H9zOAFHx9_2(.din(n11784), .dout(n11781));
    jdff dff_A_DepeEy322_2(.din(n11787), .dout(n11784));
    jdff dff_A_xiHKryJN7_2(.din(n11790), .dout(n11787));
    jdff dff_A_zCrUtDH90_2(.din(n11793), .dout(n11790));
    jdff dff_A_eN39hUaF2_2(.din(n11796), .dout(n11793));
    jdff dff_A_pLg4OBT42_2(.din(n11799), .dout(n11796));
    jdff dff_A_66N60CTd1_2(.din(n11802), .dout(n11799));
    jdff dff_A_famUi9Ow7_2(.din(n11805), .dout(n11802));
    jdff dff_A_FlQ3axMt0_2(.din(n11808), .dout(n11805));
    jdff dff_A_w0z19Z6F8_2(.din(n11811), .dout(n11808));
    jdff dff_A_QOjGnQml7_2(.din(n1460), .dout(n11811));
    jdff dff_A_j7dIH2GR1_0(.din(n11817), .dout(n11814));
    jdff dff_A_Kir7Rrku2_0(.din(n1452), .dout(n11817));
    jdff dff_B_ushaR9vI3_0(.din(G155), .dout(n11821));
    jdff dff_B_g6uKnzF50_2(.din(n1448), .dout(n11824));
    jdff dff_B_an6MDwmU2_2(.din(n11824), .dout(n11827));
    jdff dff_A_7hEVAEFb8_1(.din(n11832), .dout(n11829));
    jdff dff_A_HWHE1biM3_1(.din(n11835), .dout(n11832));
    jdff dff_A_prTVDyTp7_1(.din(n11838), .dout(n11835));
    jdff dff_A_8ufHP8OR6_1(.din(n11841), .dout(n11838));
    jdff dff_A_6arFQ3iJ3_1(.din(n1441), .dout(n11841));
    jdff dff_B_7BmYyDMm7_1(.din(n1363), .dout(n11845));
    jdff dff_B_SlYEXmrL8_1(.din(n11845), .dout(n11848));
    jdff dff_B_xlCfDRVl8_1(.din(n11848), .dout(n11851));
    jdff dff_B_LHWRhSg61_1(.din(n11851), .dout(n11854));
    jdff dff_B_bOwuuzCy2_1(.din(n11854), .dout(n11857));
    jdff dff_B_9fDOTzUJ0_1(.din(n11857), .dout(n11860));
    jdff dff_B_D5Q2xOZA1_1(.din(n1370), .dout(n11863));
    jdff dff_B_yME1aZo34_1(.din(n11863), .dout(n11866));
    jdff dff_B_rpVKhQ6F6_1(.din(n11866), .dout(n11869));
    jdff dff_B_l3n405Ep5_1(.din(n11869), .dout(n11872));
    jdff dff_B_IFTfh1mX6_1(.din(n11872), .dout(n11875));
    jdff dff_A_81XBlqvm4_0(.din(n11880), .dout(n11877));
    jdff dff_A_D1phObl95_0(.din(n11883), .dout(n11880));
    jdff dff_A_uHmO9OH33_0(.din(n11886), .dout(n11883));
    jdff dff_A_h3AVsrzd6_0(.din(n11889), .dout(n11886));
    jdff dff_A_REXG7Zhp7_0(.din(n11892), .dout(n11889));
    jdff dff_A_vklsPczg5_0(.din(n11895), .dout(n11892));
    jdff dff_A_4QMJZCK65_0(.din(n11898), .dout(n11895));
    jdff dff_A_VsAIbkmZ9_0(.din(n11901), .dout(n11898));
    jdff dff_A_KrygBMp55_0(.din(n1433), .dout(n11901));
    jdff dff_B_6pPOnS6H0_1(.din(n1377), .dout(n11905));
    jdff dff_B_TlsEcBTW6_1(.din(n11905), .dout(n11908));
    jdff dff_B_iTUWS4sz1_1(.din(n11908), .dout(n11911));
    jdff dff_B_bO2tCcQc4_1(.din(n11911), .dout(n11914));
    jdff dff_B_x1Yl5yVa8_1(.din(n1384), .dout(n11917));
    jdff dff_B_wFDA0cag7_1(.din(n11917), .dout(n11920));
    jdff dff_B_PSNRXKgT4_1(.din(n11920), .dout(n11923));
    jdff dff_A_wjUihQaD1_1(.din(n11928), .dout(n11925));
    jdff dff_A_x70VSDT46_1(.din(n11931), .dout(n11928));
    jdff dff_A_KmiCco6I6_1(.din(n11934), .dout(n11931));
    jdff dff_A_JyowotkQ5_1(.din(n11937), .dout(n11934));
    jdff dff_A_5jgCpFzy0_1(.din(n11940), .dout(n11937));
    jdff dff_A_AmXvraAA1_1(.din(n11943), .dout(n11940));
    jdff dff_A_8UQcol652_1(.din(n11946), .dout(n11943));
    jdff dff_A_WbBHUvTq9_1(.din(n11949), .dout(n11946));
    jdff dff_A_9cezoIdV4_1(.din(n11952), .dout(n11949));
    jdff dff_A_AeGQcbZC4_1(.din(n1425), .dout(n11952));
    jdff dff_A_JOD0nreV1_0(.din(n11958), .dout(n11955));
    jdff dff_A_Nei84SfY4_0(.din(n1414), .dout(n11958));
    jdff dff_A_OyMjnSER3_0(.din(n11964), .dout(n11961));
    jdff dff_A_nv66cA3z1_0(.din(n1406), .dout(n11964));
    jdff dff_A_PGBKZuMi7_0(.din(n11970), .dout(n11967));
    jdff dff_A_D2YnCEkM4_0(.din(n11973), .dout(n11970));
    jdff dff_A_FuQ2lwZi3_0(.din(n11976), .dout(n11973));
    jdff dff_A_8CDfmc8z6_0(.din(n1398), .dout(n11976));
    jdff dff_A_gFW2FglF0_1(.din(n11982), .dout(n11979));
    jdff dff_A_MfH5EZsL5_1(.din(n11985), .dout(n11982));
    jdff dff_A_OgMELuPM1_1(.din(n11988), .dout(n11985));
    jdff dff_A_lI0VZls23_1(.din(n11991), .dout(n11988));
    jdff dff_A_y36RNCp36_1(.din(n11994), .dout(n11991));
    jdff dff_A_auSOT7Ez1_1(.din(n11997), .dout(n11994));
    jdff dff_A_07zLDTuy0_1(.din(n12000), .dout(n11997));
    jdff dff_A_3Gaffbtx8_1(.din(n12003), .dout(n12000));
    jdff dff_A_Legihi8a8_1(.din(n12006), .dout(n12003));
    jdff dff_A_pRiVCr5C8_1(.din(n12009), .dout(n12006));
    jdff dff_A_nQrK5SOy7_1(.din(n12012), .dout(n12009));
    jdff dff_A_90PfBetN6_1(.din(n12015), .dout(n12012));
    jdff dff_A_sIc5B8IA5_1(.din(n1398), .dout(n12015));
    jdff dff_A_bpIZOWyw1_0(.din(n12021), .dout(n12018));
    jdff dff_A_gsuy1xhg7_0(.din(n12024), .dout(n12021));
    jdff dff_A_NVkVw5Rr0_0(.din(n12027), .dout(n12024));
    jdff dff_A_9kPS5u6Z9_0(.din(n12030), .dout(n12027));
    jdff dff_A_cOrKHC8r7_0(.din(n1374), .dout(n12030));
    jdff dff_B_ALmpcn5E2_0(.din(n1352), .dout(n12034));
    jdff dff_B_8DMOOf4i3_0(.din(n12034), .dout(n12037));
    jdff dff_B_m293t9WZ8_0(.din(n12037), .dout(n12040));
    jdff dff_B_gmoTMHaR0_0(.din(n12040), .dout(n12043));
    jdff dff_B_d5sNZA4I3_0(.din(n12043), .dout(n12046));
    jdff dff_B_IDfMCid82_0(.din(n12046), .dout(n12049));
    jdff dff_B_3MDwyOK57_0(.din(n12049), .dout(n12052));
    jdff dff_B_fuApnOfa2_0(.din(n12052), .dout(n12055));
    jdff dff_A_zcwsYSNy8_0(.din(n12060), .dout(n12057));
    jdff dff_A_lLbhIJXG0_0(.din(n12063), .dout(n12060));
    jdff dff_A_pM3KtXqT8_0(.din(n12066), .dout(n12063));
    jdff dff_A_ps7QqfkW5_0(.din(n12069), .dout(n12066));
    jdff dff_A_z7tTAFy69_0(.din(n12072), .dout(n12069));
    jdff dff_A_No7cUPur3_0(.din(n12075), .dout(n12072));
    jdff dff_A_PTQffy812_0(.din(n12078), .dout(n12075));
    jdff dff_A_6lDzlWRP6_0(.din(n12081), .dout(n12078));
    jdff dff_A_LwVKvSsc3_0(.din(n1349), .dout(n12081));
    jdff dff_A_VcZ0ObV67_1(.din(n1337), .dout(n12084));
    jdff dff_B_DeBhIout9_0(.din(n1329), .dout(n12088));
    jdff dff_B_lV3ChrZN8_0(.din(G144), .dout(n12091));
    jdff dff_B_xZ08vA4y3_2(.din(n1321), .dout(n12094));
    jdff dff_B_WDEbrLem7_2(.din(n12094), .dout(n12097));
    jdff dff_A_fzbjfxrA9_0(.din(n12102), .dout(n12099));
    jdff dff_A_479Mr7cO0_0(.din(n12105), .dout(n12102));
    jdff dff_A_W3X3aebx9_0(.din(n12108), .dout(n12105));
    jdff dff_A_mm6HwVJP0_0(.din(G2224), .dout(n12108));
    jdff dff_B_D5js8nOw4_0(.din(n1310), .dout(n12112));
    jdff dff_B_1N5R0yCL3_0(.din(G135), .dout(n12115));
    jdff dff_B_0K0C5rfL1_2(.din(n1302), .dout(n12118));
    jdff dff_B_0BNgGgMg3_2(.din(n12118), .dout(n12121));
    jdff dff_A_cm1WQzw24_0(.din(n12126), .dout(n12123));
    jdff dff_A_AxAcsGCx7_0(.din(n12129), .dout(n12126));
    jdff dff_A_UmwWKvEW7_0(.din(n12132), .dout(n12129));
    jdff dff_A_1rQxkaMZ6_0(.din(G2230), .dout(n12132));
    jdff dff_A_zXQNcWHq8_0(.din(n12138), .dout(n12135));
    jdff dff_A_LZhMNDa49_0(.din(n12141), .dout(n12138));
    jdff dff_A_IYbuSqnC5_0(.din(n12144), .dout(n12141));
    jdff dff_A_hTIxALdH9_0(.din(n12147), .dout(n12144));
    jdff dff_A_MKUfhvux9_0(.din(n12150), .dout(n12147));
    jdff dff_A_2mCGjD1i9_0(.din(n12153), .dout(n12150));
    jdff dff_A_QL5ApbaD7_0(.din(n12156), .dout(n12153));
    jdff dff_A_Gz8E25yi4_0(.din(n12159), .dout(n12156));
    jdff dff_A_iuTt8jDK2_0(.din(n12162), .dout(n12159));
    jdff dff_A_4Px20A4r9_0(.din(n12165), .dout(n12162));
    jdff dff_A_iK6pO9725_0(.din(n12168), .dout(n12165));
    jdff dff_A_BLNwJD364_0(.din(n1295), .dout(n12168));
    jdff dff_A_GcFNFohd4_1(.din(n12174), .dout(n12171));
    jdff dff_A_GipSjDUt4_1(.din(n12177), .dout(n12174));
    jdff dff_A_OP4lTLMV3_1(.din(n12180), .dout(n12177));
    jdff dff_A_qtJnsGNi4_1(.din(n1295), .dout(n12180));
    jdff dff_A_q2fnkuVw8_2(.din(n12186), .dout(n12183));
    jdff dff_A_batIeYWG1_2(.din(n12189), .dout(n12186));
    jdff dff_A_OINP2Htl1_2(.din(n12192), .dout(n12189));
    jdff dff_A_f7oh9e0H0_2(.din(n12195), .dout(n12192));
    jdff dff_A_7qcirIbk1_2(.din(n12198), .dout(n12195));
    jdff dff_A_NZAOmBEF5_2(.din(n12201), .dout(n12198));
    jdff dff_A_Z41uG3Qb5_2(.din(n12204), .dout(n12201));
    jdff dff_A_dct5lZS76_2(.din(n12207), .dout(n12204));
    jdff dff_A_6B2059224_2(.din(n12210), .dout(n12207));
    jdff dff_A_kTiYQC3z8_2(.din(n12213), .dout(n12210));
    jdff dff_A_1G46lzN70_2(.din(n12216), .dout(n12213));
    jdff dff_A_AR6PB7eS3_2(.din(n1295), .dout(n12216));
    jdff dff_B_3C2QXZfv3_0(.din(n1287), .dout(n12220));
    jdff dff_B_rnocEosP8_0(.din(G147), .dout(n12223));
    jdff dff_B_77YsmIWU1_2(.din(n1279), .dout(n12226));
    jdff dff_B_sKxW7ouH5_2(.din(n12226), .dout(n12229));
    jdff dff_A_wILlbT7T3_2(.din(n12234), .dout(n12231));
    jdff dff_A_4YWfzSay5_2(.din(n12237), .dout(n12234));
    jdff dff_A_Kne2JWyF3_2(.din(n12240), .dout(n12237));
    jdff dff_A_6MKETmv02_2(.din(n12243), .dout(n12240));
    jdff dff_A_BFa9jBAm4_2(.din(n12246), .dout(n12243));
    jdff dff_A_UZhSkQ3u9_2(.din(n12249), .dout(n12246));
    jdff dff_A_QcSwRD9w2_2(.din(n12252), .dout(n12249));
    jdff dff_A_zFfFWEtR2_2(.din(n12255), .dout(n12252));
    jdff dff_A_yICARhwM9_2(.din(n12258), .dout(n12255));
    jdff dff_A_SW4xabWb7_2(.din(n12261), .dout(n12258));
    jdff dff_A_rpso9bRS2_2(.din(n12264), .dout(n12261));
    jdff dff_A_gRtxQXhT5_2(.din(n12267), .dout(n12264));
    jdff dff_A_txnbFa000_2(.din(n12270), .dout(n12267));
    jdff dff_A_xnCWaTuR7_2(.din(n1276), .dout(n12270));
    jdff dff_A_Ao79kSAN0_2(.din(n1272), .dout(n12273));
    jdff dff_B_KhfQAqlt3_0(.din(n1268), .dout(n12277));
    jdff dff_B_3uEs4dVE0_0(.din(G138), .dout(n12280));
    jdff dff_B_oNNov6Cs0_3(.din(n1260), .dout(n12283));
    jdff dff_B_syGTL4xv9_3(.din(n12283), .dout(n12286));
    jdff dff_A_iL4NUDBV5_0(.din(n12291), .dout(n12288));
    jdff dff_A_kb6YfBSF5_0(.din(n12294), .dout(n12291));
    jdff dff_A_bUkzMEKL9_0(.din(n12297), .dout(n12294));
    jdff dff_A_7k2u0Uhk4_0(.din(n1257), .dout(n12297));
    jdff dff_A_mBGChZA09_2(.din(n12303), .dout(n12300));
    jdff dff_A_KB6PSNHp2_2(.din(n1257), .dout(n12303));
    jdff dff_B_gkRoOqZ43_0(.din(G157), .dout(n12307));
    jdff dff_A_FdM5IzSU3_0(.din(n12312), .dout(n12309));
    jdff dff_A_yGaO7Vih8_0(.din(n12315), .dout(n12312));
    jdff dff_A_VMS3oj4g6_0(.din(n1242), .dout(n12315));
    jdff dff_A_d8qwEVrX0_1(.din(n1242), .dout(n12318));
    jdff dff_B_yVkI5nMr4_2(.din(n1238), .dout(n12322));
    jdff dff_B_YAXYqcGI0_2(.din(n12322), .dout(n12325));
    jdff dff_A_u6ht5Zzm1_0(.din(n12330), .dout(n12327));
    jdff dff_A_fPsIodG79_0(.din(n12333), .dout(n12330));
    jdff dff_A_soUu5tBA0_0(.din(n12336), .dout(n12333));
    jdff dff_A_j7vDye4R5_0(.din(G2236), .dout(n12336));
    jdff dff_B_6qNqKJ7I7_0(.din(n1231), .dout(n12340));
    jdff dff_B_zhQ5zoaN3_0(.din(n12340), .dout(n12343));
    jdff dff_B_oZxpILHP5_0(.din(n12343), .dout(n12346));
    jdff dff_B_eqNB2x3B1_0(.din(n12346), .dout(n12349));
    jdff dff_A_pf5blDt83_0(.din(n12354), .dout(n12351));
    jdff dff_A_GJmzwBgT8_0(.din(n12357), .dout(n12354));
    jdff dff_A_j8v0MkH30_0(.din(n12360), .dout(n12357));
    jdff dff_A_ugtOsKZg0_0(.din(n12363), .dout(n12360));
    jdff dff_A_GOtlVnN46_0(.din(n1228), .dout(n12363));
    jdff dff_B_j2k8mZZE5_1(.din(n1178), .dout(n12367));
    jdff dff_B_v4dk76pM1_1(.din(n12367), .dout(n12370));
    jdff dff_B_INxAodTD2_1(.din(n12370), .dout(n12373));
    jdff dff_B_3EeUhV7m3_1(.din(n1182), .dout(n12376));
    jdff dff_B_4KCJDPpx6_1(.din(n12376), .dout(n12379));
    jdff dff_B_YYMfaYUU9_1(.din(n12379), .dout(n12382));
    jdff dff_B_bU2JFqUT9_1(.din(n12382), .dout(n12385));
    jdff dff_B_DTSOZ4kH2_0(.din(n1164), .dout(n12388));
    jdff dff_B_HVTNJEOF6_0(.din(n12388), .dout(n12391));
    jdff dff_B_SnIFAloN7_0(.din(n12391), .dout(n12394));
    jdff dff_B_6UuhMnFy3_0(.din(n12394), .dout(n12397));
    jdff dff_B_6h0p151i4_0(.din(n12397), .dout(n12400));
    jdff dff_B_g93XN7Hd9_0(.din(n12400), .dout(n12403));
    jdff dff_B_Cd0jMb9i0_0(.din(n12403), .dout(n12406));
    jdff dff_A_0tNitACA4_0(.din(n12411), .dout(n12408));
    jdff dff_A_NqvdE97N4_0(.din(n12414), .dout(n12411));
    jdff dff_A_V0ljnoLg8_0(.din(n12417), .dout(n12414));
    jdff dff_A_ccNtsWX08_0(.din(n12420), .dout(n12417));
    jdff dff_A_FIyJsI0G3_0(.din(n12423), .dout(n12420));
    jdff dff_A_xnYzgbV02_0(.din(n12426), .dout(n12423));
    jdff dff_A_5Z8h4EPz9_0(.din(n12429), .dout(n12426));
    jdff dff_A_DjpXitUl9_0(.din(n1161), .dout(n12429));
    jdff dff_A_JovB0lwN3_0(.din(n12435), .dout(n12432));
    jdff dff_A_E5K7alzc4_0(.din(n12438), .dout(n12435));
    jdff dff_A_KJ3vDEya8_0(.din(n12441), .dout(n12438));
    jdff dff_A_eheffV112_0(.din(n12444), .dout(n12441));
    jdff dff_A_joYyMP7n7_0(.din(n12447), .dout(n12444));
    jdff dff_A_KU3rHIqv9_0(.din(n12450), .dout(n12447));
    jdff dff_A_hB3e9Lal8_0(.din(n12453), .dout(n12450));
    jdff dff_A_czRxNlFA7_0(.din(n12456), .dout(n12453));
    jdff dff_A_xfECxXcF3_0(.din(n12459), .dout(n12456));
    jdff dff_A_PJSjd5ZO0_0(.din(n12462), .dout(n12459));
    jdff dff_A_EXpZaSpZ3_0(.din(n12465), .dout(n12462));
    jdff dff_A_R5aBBOiV2_0(.din(n12468), .dout(n12465));
    jdff dff_A_1GIilQCR3_0(.din(n1134), .dout(n12468));
    jdff dff_A_px7SGiXE3_0(.din(n12474), .dout(n12471));
    jdff dff_A_m3rSiGQ31_0(.din(n12477), .dout(n12474));
    jdff dff_A_suR2No9l5_0(.din(n12480), .dout(n12477));
    jdff dff_A_0NvkXn7P2_0(.din(n12483), .dout(n12480));
    jdff dff_A_Mk4ll8HJ2_0(.din(n12486), .dout(n12483));
    jdff dff_A_G0ExnXCE7_0(.din(n12489), .dout(n12486));
    jdff dff_A_niLYAnRN9_0(.din(n12492), .dout(n12489));
    jdff dff_A_BFIbBuJj1_0(.din(n12495), .dout(n12492));
    jdff dff_A_CmHLRX2u3_0(.din(n1115), .dout(n12495));
    jdff dff_A_CJ2XfhFk2_0(.din(n12501), .dout(n12498));
    jdff dff_A_VCRb9KBz1_0(.din(n12504), .dout(n12501));
    jdff dff_A_wh4rldlH9_0(.din(n12507), .dout(n12504));
    jdff dff_A_kusIEkBs1_0(.din(n12510), .dout(n12507));
    jdff dff_A_DpbZDXwP0_0(.din(n12513), .dout(n12510));
    jdff dff_A_lPdV6RPk9_0(.din(n12516), .dout(n12513));
    jdff dff_A_dDUxUmdE1_0(.din(n12519), .dout(n12516));
    jdff dff_A_mmuEb3QL8_0(.din(n12522), .dout(n12519));
    jdff dff_A_AhamDzMV9_0(.din(n12525), .dout(n12522));
    jdff dff_A_CscisU493_0(.din(n1111), .dout(n12525));
    jdff dff_A_vO6IatWr4_0(.din(n12531), .dout(n12528));
    jdff dff_A_rJFI9lK38_0(.din(n12534), .dout(n12531));
    jdff dff_A_qKcgb3jQ7_0(.din(n12537), .dout(n12534));
    jdff dff_A_gDjcuU4m7_0(.din(n12540), .dout(n12537));
    jdff dff_A_KfEs8R6r0_0(.din(n12543), .dout(n12540));
    jdff dff_A_kRLrKGtV7_0(.din(n12546), .dout(n12543));
    jdff dff_A_HiBM4pVC7_0(.din(n12549), .dout(n12546));
    jdff dff_A_EGetv3MI1_0(.din(n12552), .dout(n12549));
    jdff dff_A_cKy94sAX5_0(.din(n12555), .dout(n12552));
    jdff dff_A_tXHQJMnv0_0(.din(n12558), .dout(n12555));
    jdff dff_A_ZxbK0vmW0_0(.din(n4680), .dout(n12558));
    jdff dff_A_gMf7R9sU2_1(.din(n12564), .dout(n12561));
    jdff dff_A_D5fs9vIB1_1(.din(n12567), .dout(n12564));
    jdff dff_A_3K7rC5Qk6_1(.din(n12570), .dout(n12567));
    jdff dff_A_WiNWTh6M3_1(.din(n12573), .dout(n12570));
    jdff dff_A_AZaIBfQd3_1(.din(n12576), .dout(n12573));
    jdff dff_A_0gFLWxzC7_1(.din(n12579), .dout(n12576));
    jdff dff_A_ranaJklK5_1(.din(n12582), .dout(n12579));
    jdff dff_A_4FRVz7XB5_1(.din(n12585), .dout(n12582));
    jdff dff_A_jEvkwzsX6_1(.din(n12588), .dout(n12585));
    jdff dff_A_t6sEAL5Z8_1(.din(n12591), .dout(n12588));
    jdff dff_A_iwIUXNDC4_1(.din(n12594), .dout(n12591));
    jdff dff_A_MbKVSPC10_1(.din(n12597), .dout(n12594));
    jdff dff_A_hfE9EebZ0_1(.din(n12600), .dout(n12597));
    jdff dff_A_2LREpPro2_1(.din(n12603), .dout(n12600));
    jdff dff_A_GAxHeVLN5_1(.din(n12606), .dout(n12603));
    jdff dff_A_bvKcreuB4_1(.din(n12609), .dout(n12606));
    jdff dff_A_hIUtR8a03_1(.din(n12612), .dout(n12609));
    jdff dff_A_PBd0LuDz8_1(.din(n12615), .dout(n12612));
    jdff dff_A_RGme1VQO3_1(.din(n4680), .dout(n12615));
    jdff dff_B_uHLU5VDr0_0(.din(n4676), .dout(n12619));
    jdff dff_A_eAUesVzk7_1(.din(n12624), .dout(n12621));
    jdff dff_A_xFztVBjF1_1(.din(n12627), .dout(n12624));
    jdff dff_A_xmevM6pX6_1(.din(n12630), .dout(n12627));
    jdff dff_A_IjN4mPtd6_1(.din(n12633), .dout(n12630));
    jdff dff_A_5KN7Waln8_1(.din(n12636), .dout(n12633));
    jdff dff_A_oeUb5HEf1_1(.din(n12639), .dout(n12636));
    jdff dff_A_WgF7CZ8P1_1(.din(n12642), .dout(n12639));
    jdff dff_A_2VlzlvdJ3_1(.din(n12645), .dout(n12642));
    jdff dff_A_aeGU1Iix2_1(.din(n12648), .dout(n12645));
    jdff dff_A_t5iGKbeR6_1(.din(n12651), .dout(n12648));
    jdff dff_A_gx9i3qNR3_1(.din(n12654), .dout(n12651));
    jdff dff_A_6aVfz3u40_1(.din(n12657), .dout(n12654));
    jdff dff_A_DrolHScC2_1(.din(n12660), .dout(n12657));
    jdff dff_A_S4OE00AN7_1(.din(n12663), .dout(n12660));
    jdff dff_A_R9H01SW31_1(.din(n12666), .dout(n12663));
    jdff dff_A_n78vXkR71_1(.din(n12669), .dout(n12666));
    jdff dff_A_eagtifbf5_1(.din(n12672), .dout(n12669));
    jdff dff_A_DInUTTPn0_1(.din(n12675), .dout(n12672));
    jdff dff_A_dzkYWVGd4_1(.din(n12678), .dout(n12675));
    jdff dff_A_EvcAKS2p6_1(.din(n12681), .dout(n12678));
    jdff dff_A_9zWEW9xr4_1(.din(n494), .dout(n12681));
    jdff dff_A_FDYHxj9q1_0(.din(n12687), .dout(n12684));
    jdff dff_A_YVjUeDoE8_0(.din(n12690), .dout(n12687));
    jdff dff_A_5gGa3kNr3_0(.din(G38), .dout(n12690));
    jdff dff_A_VmzUsI6k4_2(.din(G38), .dout(n12693));
    jdff dff_A_WJWqTm6j3_1(.din(G38), .dout(n12696));
    jdff dff_A_GrQxdQNd2_2(.din(n12702), .dout(n12699));
    jdff dff_A_DvvVmoVy6_2(.din(G38), .dout(n12702));
    jdff dff_B_H54XB8QL4_1(.din(n5160), .dout(n12706));
    jdff dff_B_kEK1mXdw5_1(.din(n12706), .dout(n12709));
    jdff dff_B_5dHBPNPx4_1(.din(n12709), .dout(n12712));
    jdff dff_B_mIULG2T30_1(.din(n12712), .dout(n12715));
    jdff dff_B_2zhiKpty8_1(.din(n12715), .dout(n12718));
    jdff dff_B_4A3Dnlax8_1(.din(n12718), .dout(n12721));
    jdff dff_B_pA6yzUWF7_1(.din(n12721), .dout(n12724));
    jdff dff_B_60QWl5sd9_1(.din(n12724), .dout(n12727));
    jdff dff_B_xqiXDl2v5_1(.din(n12727), .dout(n12730));
    jdff dff_B_ceOtUC3a3_1(.din(n12730), .dout(n12733));
    jdff dff_B_WPeyNfHw0_1(.din(n12733), .dout(n12736));
    jdff dff_B_ASHbUCWz7_1(.din(n12736), .dout(n12739));
    jdff dff_B_OKEBBw1v9_1(.din(n5233), .dout(n12742));
    jdff dff_B_xMBW8gtM9_1(.din(n12742), .dout(n12745));
    jdff dff_B_ez4oe8O89_1(.din(n5287), .dout(n12748));
    jdff dff_B_tP5QGGy90_1(.din(n12748), .dout(n12751));
    jdff dff_B_4Gm3sYUt8_1(.din(n5295), .dout(n12754));
    jdff dff_B_FUVbq3kE0_1(.din(n12754), .dout(n12757));
    jdff dff_B_82E0SqC84_1(.din(n12757), .dout(n12760));
    jdff dff_B_H0YLKs2Y6_1(.din(n12760), .dout(n12763));
    jdff dff_B_AMKVK5VG7_1(.din(n12763), .dout(n12766));
    jdff dff_B_79HMWNLb4_1(.din(n12766), .dout(n12769));
    jdff dff_B_nw132nbh3_1(.din(n5299), .dout(n12772));
    jdff dff_B_wwJVCGX44_1(.din(n12772), .dout(n12775));
    jdff dff_B_MkWhOmse4_1(.din(n12775), .dout(n12778));
    jdff dff_B_MjDQdwRa4_1(.din(n12778), .dout(n12781));
    jdff dff_B_1UGtU2pP1_1(.din(n12781), .dout(n12784));
    jdff dff_B_eYsFY6Dz2_1(.din(n12784), .dout(n12787));
    jdff dff_B_ldlJ2nWL0_1(.din(n12787), .dout(n12790));
    jdff dff_B_lxx2CanO3_1(.din(n12790), .dout(n12793));
    jdff dff_B_tmvJ6XVG7_1(.din(n5311), .dout(n12796));
    jdff dff_B_nGaZYB9h6_1(.din(n12796), .dout(n12799));
    jdff dff_B_9XJZ6PK16_0(.din(n5303), .dout(n12802));
    jdff dff_B_4stDTBS90_0(.din(n12802), .dout(n12805));
    jdff dff_A_g0sE4gYu5_1(.din(n12810), .dout(n12807));
    jdff dff_A_WG64xLY17_1(.din(n12813), .dout(n12810));
    jdff dff_A_sjwH9waE9_1(.din(n12816), .dout(n12813));
    jdff dff_A_Qzifh2BF2_1(.din(n12819), .dout(n12816));
    jdff dff_A_XyOJ4ZVF4_1(.din(n12822), .dout(n12819));
    jdff dff_A_KtsyxYg13_1(.din(n4739), .dout(n12822));
    jdff dff_A_Ed8GysSM6_1(.din(n12828), .dout(n12825));
    jdff dff_A_VkjFpfeo2_1(.din(n12831), .dout(n12828));
    jdff dff_A_L9MFRLub6_1(.din(n12834), .dout(n12831));
    jdff dff_A_t1OorFeT8_1(.din(n12837), .dout(n12834));
    jdff dff_A_pJKJ5JGS9_1(.din(n4707), .dout(n12837));
    jdff dff_B_AFVHb2Dm8_1(.din(n5245), .dout(n12841));
    jdff dff_B_VTOZJaWd5_1(.din(n12841), .dout(n12844));
    jdff dff_B_zMT5VBaP1_1(.din(n12844), .dout(n12847));
    jdff dff_B_Jmwo1Vpq5_1(.din(n12847), .dout(n12850));
    jdff dff_B_hIlveP8D7_1(.din(n12850), .dout(n12853));
    jdff dff_B_2yNwb2Rz4_1(.din(n12853), .dout(n12856));
    jdff dff_B_XKqHvp1z8_0(.din(n5267), .dout(n12859));
    jdff dff_A_KjU7AqUT0_1(.din(n12864), .dout(n12861));
    jdff dff_A_tLo5OXNk5_1(.din(n12867), .dout(n12864));
    jdff dff_A_5lvn2ewi5_1(.din(n12870), .dout(n12867));
    jdff dff_A_W1Q2ulZp0_1(.din(n12873), .dout(n12870));
    jdff dff_A_iO7mZrfs7_1(.din(n12876), .dout(n12873));
    jdff dff_A_Y5jRghTd6_1(.din(n12879), .dout(n12876));
    jdff dff_A_0WAxktpG4_1(.din(n4750), .dout(n12879));
    jdff dff_A_syDZq2026_1(.din(n12885), .dout(n12882));
    jdff dff_A_F77pSxzR3_1(.din(n12888), .dout(n12885));
    jdff dff_A_jLvMlcrl4_1(.din(n12891), .dout(n12888));
    jdff dff_A_JR4JKGp92_1(.din(n12894), .dout(n12891));
    jdff dff_A_vaUUkInl2_1(.din(n12913), .dout(n12894));
    jdff dff_B_donYkLVC3_2(.din(n4698), .dout(n12898));
    jdff dff_B_mbjCN1LT8_2(.din(n12898), .dout(n12901));
    jdff dff_B_IoS9XBZo6_2(.din(n12901), .dout(n12904));
    jdff dff_B_WdTyTBTI2_2(.din(n12904), .dout(n12907));
    jdff dff_B_p5naMZBK5_2(.din(n12907), .dout(n12910));
    jdff dff_B_jllnJNpC9_2(.din(n12910), .dout(n12913));
    jdff dff_B_2ZlPMjFp5_2(.din(n5248), .dout(n12916));
    jdff dff_B_4ORWPjYZ0_1(.din(n5237), .dout(n12919));
    jdff dff_B_IERriCYy9_0(.din(n5225), .dout(n12922));
    jdff dff_B_EjHF14WT6_0(.din(n12922), .dout(n12925));
    jdff dff_B_ornnWYyA2_1(.din(n5198), .dout(n12928));
    jdff dff_B_IDeAhHgO2_1(.din(n12928), .dout(n12931));
    jdff dff_B_86ioJiNl5_1(.din(n12931), .dout(n12934));
    jdff dff_B_DpYNnzbp2_1(.din(n12934), .dout(n12937));
    jdff dff_B_1DOt81Ad4_1(.din(n12937), .dout(n12940));
    jdff dff_B_sel0X8RR9_0(.din(n5217), .dout(n12943));
    jdff dff_A_FnpgA7eZ4_0(.din(n1220), .dout(n12945));
    jdff dff_A_Ng5qy9pI2_1(.din(n12951), .dout(n12948));
    jdff dff_A_kUyaWBU63_1(.din(n12954), .dout(n12951));
    jdff dff_A_lRVvlXKr1_1(.din(n12957), .dout(n12954));
    jdff dff_A_4BSE3NL41_1(.din(n12960), .dout(n12957));
    jdff dff_A_bHanTw4u7_1(.din(n12963), .dout(n12960));
    jdff dff_A_P3pamEE47_1(.din(n12966), .dout(n12963));
    jdff dff_A_5E4wL1zE3_1(.din(n12969), .dout(n12966));
    jdff dff_A_XixEvbBh8_1(.din(n1220), .dout(n12969));
    jdff dff_A_IynqEskC4_1(.din(n12975), .dout(n12972));
    jdff dff_A_0gA4mnx75_1(.din(n4369), .dout(n12975));
    jdff dff_B_vi9gKCrh7_0(.din(n4358), .dout(n12979));
    jdff dff_B_Pr4cRVXm5_0(.din(n5186), .dout(n12982));
    jdff dff_B_Eh2Rk16E7_0(.din(n12982), .dout(n12985));
    jdff dff_B_VkEavW1t2_0(.din(n12985), .dout(n12988));
    jdff dff_B_9ZpuAkHu2_0(.din(n5182), .dout(n12991));
    jdff dff_B_RjQZLPU06_0(.din(n12991), .dout(n12994));
    jdff dff_B_XX9PT8uf5_0(.din(n12994), .dout(n12997));
    jdff dff_A_CMDxxD1q7_2(.din(n13002), .dout(n12999));
    jdff dff_A_CCfkFeBt8_2(.din(n13005), .dout(n13002));
    jdff dff_A_4GL5I2FX7_2(.din(n13008), .dout(n13005));
    jdff dff_A_9C6nb4KK7_2(.din(n13011), .dout(n13008));
    jdff dff_A_CHLv29ha1_2(.din(n13014), .dout(n13011));
    jdff dff_A_27sUQoDV3_2(.din(n13017), .dout(n13014));
    jdff dff_A_I8542ZhQ6_2(.din(n13020), .dout(n13017));
    jdff dff_A_IGyUEtNS0_2(.din(n4796), .dout(n13020));
    jdff dff_A_opi42OKV6_1(.din(n13026), .dout(n13023));
    jdff dff_A_50Pk9rpa7_1(.din(n1092), .dout(n13026));
    jdff dff_A_h97gtSDy3_2(.din(n13032), .dout(n13029));
    jdff dff_A_KDwJqF2U7_2(.din(n13035), .dout(n13032));
    jdff dff_A_nyalX7Vu4_2(.din(n13038), .dout(n13035));
    jdff dff_A_EJWBJjO24_2(.din(n13041), .dout(n13038));
    jdff dff_A_kyC7fiAW9_2(.din(n13044), .dout(n13041));
    jdff dff_A_gSCgWGLe3_2(.din(n13047), .dout(n13044));
    jdff dff_A_UasxrxzM1_2(.din(n13050), .dout(n13047));
    jdff dff_A_3loQDpa12_2(.din(n13053), .dout(n13050));
    jdff dff_A_tJTwwsdY4_2(.din(n13056), .dout(n13053));
    jdff dff_A_RAC4MjRG2_2(.din(n13059), .dout(n13056));
    jdff dff_A_ihl4IpdQ5_2(.din(n13062), .dout(n13059));
    jdff dff_A_GMvBdxUO4_2(.din(n1092), .dout(n13062));
    jdff dff_B_OIKxCJxU6_1(.din(n5163), .dout(n13066));
    jdff dff_B_GJv8SWDd3_1(.din(n13066), .dout(n13069));
    jdff dff_B_xgc1Od2f3_1(.din(n13069), .dout(n13072));
    jdff dff_B_mm7fPUEe4_1(.din(n13072), .dout(n13075));
    jdff dff_B_2DsdV5O88_0(.din(n5170), .dout(n13078));
    jdff dff_A_x19YsS0i6_1(.din(n13087), .dout(n13080));
    jdff dff_B_SAlCeFYl0_2(.din(n1186), .dout(n13084));
    jdff dff_B_rFAGAFOx4_2(.din(n13084), .dout(n13087));
    jdff dff_A_fzKjvWig5_1(.din(n13092), .dout(n13089));
    jdff dff_A_HtvCpDy58_1(.din(n13095), .dout(n13092));
    jdff dff_A_Ns2WddQp2_1(.din(n13098), .dout(n13095));
    jdff dff_A_s7orHyME7_1(.din(n13101), .dout(n13098));
    jdff dff_A_9BI1CyFY4_1(.din(n13104), .dout(n13101));
    jdff dff_A_sKP7S97R2_1(.din(n13107), .dout(n13104));
    jdff dff_A_7MI3tEFm7_1(.din(n13110), .dout(n13107));
    jdff dff_A_lwZauxQ99_1(.din(n13113), .dout(n13110));
    jdff dff_A_W9Oe9Irk5_1(.din(n1212), .dout(n13113));
    jdff dff_A_nCU9MRR05_1(.din(n13119), .dout(n13116));
    jdff dff_A_hHJMPfl68_1(.din(n13122), .dout(n13119));
    jdff dff_A_UqO1TnTV9_1(.din(n13125), .dout(n13122));
    jdff dff_A_iGjyd2mM3_1(.din(n13128), .dout(n13125));
    jdff dff_A_fNXRIG3F4_1(.din(n13131), .dout(n13128));
    jdff dff_A_6qYis3IZ4_1(.din(n13134), .dout(n13131));
    jdff dff_A_GIqro3PQ5_1(.din(n13137), .dout(n13134));
    jdff dff_A_pvqZuXdk9_1(.din(n13140), .dout(n13137));
    jdff dff_A_TcSk9PEH7_1(.din(n13143), .dout(n13140));
    jdff dff_A_fIfmGo6g3_1(.din(n13146), .dout(n13143));
    jdff dff_A_ck0iszft9_1(.din(n1204), .dout(n13146));
    jdff dff_B_PcBIj1gP7_1(.din(n1099), .dout(n13150));
    jdff dff_B_4FoRgvuD6_0(.din(G35), .dout(n13153));
    jdff dff_A_AqZSHEOy8_1(.din(n13158), .dout(n13155));
    jdff dff_A_4E7K3r0y5_1(.din(n1095), .dout(n13158));
    jdff dff_A_EiVtXFOz7_2(.din(n13164), .dout(n13161));
    jdff dff_A_JIK2jnnq1_2(.din(n1095), .dout(n13164));
    jdff dff_A_lAvt5qLZ3_1(.din(n13170), .dout(n13167));
    jdff dff_A_KCyLF0xG5_1(.din(n13173), .dout(n13170));
    jdff dff_A_3jSymNVW0_1(.din(n13176), .dout(n13173));
    jdff dff_A_8eBzixrq7_1(.din(G4420), .dout(n13176));
    jdff dff_A_DgDAJlvf3_2(.din(n13182), .dout(n13179));
    jdff dff_A_Iuxr2gKJ8_2(.din(n1092), .dout(n13182));
    jdff dff_A_pE32UJ6Y0_0(.din(n13188), .dout(n13185));
    jdff dff_A_5dgnjyY68_0(.din(n13192), .dout(n13188));
    jdff dff_B_JGSCKHOj3_2(.din(n1200), .dout(n13192));
    jdff dff_B_fzUH6Gwg3_1(.din(n1080), .dout(n13195));
    jdff dff_B_AJSqunPQ4_0(.din(G32), .dout(n13198));
    jdff dff_A_EhA8q3zh6_1(.din(n13203), .dout(n13200));
    jdff dff_A_rPxpNk2v5_1(.din(n1076), .dout(n13203));
    jdff dff_A_6cgcbzJM4_2(.din(n13209), .dout(n13206));
    jdff dff_A_t8sJnWpR2_2(.din(n1076), .dout(n13209));
    jdff dff_A_fDzA0mv00_0(.din(n13215), .dout(n13212));
    jdff dff_A_o5zNdw3o6_0(.din(n13218), .dout(n13215));
    jdff dff_A_Q9lzvkjn7_0(.din(n13221), .dout(n13218));
    jdff dff_A_gCT6V1oP9_0(.din(n13224), .dout(n13221));
    jdff dff_A_o1KJXdOF0_0(.din(n13227), .dout(n13224));
    jdff dff_A_DSPztC9M3_0(.din(n13230), .dout(n13227));
    jdff dff_A_4Jyj9n3U1_0(.din(n13233), .dout(n13230));
    jdff dff_A_v7Y8xzsW1_0(.din(n13236), .dout(n13233));
    jdff dff_A_EZo0lXF13_0(.din(n1196), .dout(n13236));
    jdff dff_A_wUx0yTa09_0(.din(n13242), .dout(n13239));
    jdff dff_A_UzABrpJR6_0(.din(n13245), .dout(n13242));
    jdff dff_A_EYlpZPJq4_0(.din(n1193), .dout(n13245));
    jdff dff_A_egm8n0ej7_1(.din(n1134), .dout(n13248));
    jdff dff_B_yAKEZt6k3_1(.din(n1122), .dout(n13252));
    jdff dff_B_84iRtvq86_0(.din(G66), .dout(n13255));
    jdff dff_A_0iBeJp9B8_1(.din(n13260), .dout(n13257));
    jdff dff_A_T9rOa2NS6_1(.din(n1118), .dout(n13260));
    jdff dff_A_6gtT0VQr7_2(.din(n13266), .dout(n13263));
    jdff dff_A_bcAtzUew4_2(.din(n1118), .dout(n13266));
    jdff dff_A_XB3GkqvB2_1(.din(n13272), .dout(n13269));
    jdff dff_A_r1Eae4on4_1(.din(n13275), .dout(n13272));
    jdff dff_A_BKMaKKir6_1(.din(n13278), .dout(n13275));
    jdff dff_A_VgHUHFeN3_1(.din(G4437), .dout(n13278));
    jdff dff_A_5nLHnB6C4_1(.din(n1069), .dout(n13281));
    jdff dff_B_nM3yZrsY8_1(.din(n994), .dout(n13285));
    jdff dff_B_lUP2YVfW1_1(.din(n13285), .dout(n13288));
    jdff dff_B_B0NN0BAE9_1(.din(n13288), .dout(n13291));
    jdff dff_B_FX4kO5pn5_1(.din(n13291), .dout(n13294));
    jdff dff_B_G3a7yDBn7_1(.din(n13294), .dout(n13297));
    jdff dff_B_ReywKQIc6_1(.din(n13297), .dout(n13300));
    jdff dff_B_4c1rMKSY1_1(.din(n1001), .dout(n13303));
    jdff dff_B_kVQlZe7Y6_1(.din(n13303), .dout(n13306));
    jdff dff_B_VV4ipEa63_1(.din(n13306), .dout(n13309));
    jdff dff_B_NU9PT9Tc7_1(.din(n13309), .dout(n13312));
    jdff dff_B_7bPW3G278_1(.din(n13312), .dout(n13315));
    jdff dff_A_u77RTt2G0_1(.din(n13320), .dout(n13317));
    jdff dff_A_qgFMoNKm5_1(.din(n13323), .dout(n13320));
    jdff dff_A_XTAzeNi84_1(.din(n13326), .dout(n13323));
    jdff dff_A_0LzmGCC08_1(.din(n13329), .dout(n13326));
    jdff dff_A_5qzCAV2S8_1(.din(n1061), .dout(n13329));
    jdff dff_B_uW98lKMF6_1(.din(n1015), .dout(n13333));
    jdff dff_B_wJZHFkYc5_1(.din(n13333), .dout(n13336));
    jdff dff_B_RSpnqIE92_1(.din(n13336), .dout(n13339));
    jdff dff_A_GsSCDuzU2_1(.din(n13344), .dout(n13341));
    jdff dff_A_Lh6XoaEJ7_1(.din(n13347), .dout(n13344));
    jdff dff_A_vznTILIU3_1(.din(n13350), .dout(n13347));
    jdff dff_A_DMkJGa9p8_1(.din(n13353), .dout(n13350));
    jdff dff_A_xvBOGYZI5_1(.din(n13356), .dout(n13353));
    jdff dff_A_pH4My2IA7_1(.din(n1053), .dout(n13356));
    jdff dff_A_NdcOEkCb6_0(.din(n1045), .dout(n13359));
    jdff dff_A_6U1UqLW16_0(.din(n1037), .dout(n13362));
    jdff dff_A_xxOlJ3CW8_0(.din(n13368), .dout(n13365));
    jdff dff_A_U0hXA5h91_0(.din(n1034), .dout(n13368));
    jdff dff_A_JE9mLRAe8_2(.din(n13374), .dout(n13371));
    jdff dff_A_YOXyXLCP3_2(.din(n13377), .dout(n13374));
    jdff dff_A_QXQ9j92N2_2(.din(n13380), .dout(n13377));
    jdff dff_A_zIdw6yhx1_2(.din(n1026), .dout(n13380));
    jdff dff_A_L8v9zKPK0_1(.din(n13387), .dout(n13383));
    jdff dff_B_BpLrxlZp9_2(.din(n1019), .dout(n13387));
    jdff dff_A_zzibIUZP2_0(.din(n1011), .dout(n13389));
    jdff dff_A_WeQLK4OR9_0(.din(n13405), .dout(n13392));
    jdff dff_B_KV71pfwJ2_2(.din(n1008), .dout(n13396));
    jdff dff_B_pMrX8p496_2(.din(n13396), .dout(n13399));
    jdff dff_B_EYruc3vf3_2(.din(n13399), .dout(n13402));
    jdff dff_B_Kmrt3sfJ7_2(.din(n13402), .dout(n13405));
    jdff dff_B_VVfKKsny1_0(.din(n983), .dout(n13408));
    jdff dff_B_vqSnrWII8_0(.din(n13408), .dout(n13411));
    jdff dff_B_2GNWMdUI1_0(.din(n13411), .dout(n13414));
    jdff dff_A_u1xDV8Vf1_0(.din(n13419), .dout(n13416));
    jdff dff_A_iRiUx5rP2_0(.din(n13422), .dout(n13419));
    jdff dff_A_0siaQzSh6_0(.din(n13425), .dout(n13422));
    jdff dff_A_tOfU8hJU1_0(.din(n980), .dout(n13425));
    jdff dff_A_6t7b2Fct8_0(.din(n13431), .dout(n13428));
    jdff dff_A_5pYyDCjl1_0(.din(n13434), .dout(n13431));
    jdff dff_A_F5L11Xlj2_0(.din(n13437), .dout(n13434));
    jdff dff_A_ajUlbdyL5_0(.din(n976), .dout(n13437));
    jdff dff_A_ldFYse3U6_0(.din(n13443), .dout(n13440));
    jdff dff_A_8uUtDvTF5_0(.din(n13446), .dout(n13443));
    jdff dff_A_tTHkCHta4_0(.din(n13449), .dout(n13446));
    jdff dff_A_kwfy8KXb7_0(.din(n13452), .dout(n13449));
    jdff dff_A_kqH5AU9u5_0(.din(n13455), .dout(n13452));
    jdff dff_A_qEgsXavU1_0(.din(n13458), .dout(n13455));
    jdff dff_A_PXkeGuLe9_0(.din(n926), .dout(n13458));
    jdff dff_A_fdpewNTe8_1(.din(n13464), .dout(n13461));
    jdff dff_A_WvhCOYmd0_1(.din(n13467), .dout(n13464));
    jdff dff_A_tVXKqJGB9_1(.din(n926), .dout(n13467));
    jdff dff_A_EP0sGnie1_2(.din(n13473), .dout(n13470));
    jdff dff_A_hKmYyrgv9_2(.din(n13476), .dout(n13473));
    jdff dff_A_p77vMcCr0_2(.din(n13479), .dout(n13476));
    jdff dff_A_ojFg92OK0_2(.din(n13482), .dout(n13479));
    jdff dff_A_VvOpbdxn0_2(.din(n13485), .dout(n13482));
    jdff dff_A_ENMNb7XV9_2(.din(n13488), .dout(n13485));
    jdff dff_A_NwdEVlzB8_2(.din(n926), .dout(n13488));
    jdff dff_B_I7HteV6h8_1(.din(n911), .dout(n13492));
    jdff dff_B_EYX6X5V06_0(.din(G118), .dout(n13495));
    jdff dff_A_TDelmwbm7_0(.din(n13500), .dout(n13497));
    jdff dff_A_okpQ7hcA6_0(.din(n13503), .dout(n13500));
    jdff dff_A_o0jEiWOW7_0(.din(n13506), .dout(n13503));
    jdff dff_A_F6zSoCrM3_0(.din(G4394), .dout(n13506));
    jdff dff_A_UMlRGQE61_1(.din(n907), .dout(n13509));
    jdff dff_A_Ar2t3l8F8_1(.din(n907), .dout(n13512));
    jdff dff_A_ZtNUuRnv6_2(.din(n13518), .dout(n13515));
    jdff dff_A_3o7m0Os36_2(.din(n13521), .dout(n13518));
    jdff dff_A_k7JJI3cr8_2(.din(n13524), .dout(n13521));
    jdff dff_A_atQfae210_2(.din(n13527), .dout(n13524));
    jdff dff_A_1iOGvwmI5_2(.din(n13530), .dout(n13527));
    jdff dff_A_sdAdEEBW6_2(.din(n13533), .dout(n13530));
    jdff dff_A_gk9VVL3Z7_2(.din(n13536), .dout(n13533));
    jdff dff_A_CUvmDf5J0_2(.din(n13539), .dout(n13536));
    jdff dff_A_abvw01o64_2(.din(n13542), .dout(n13539));
    jdff dff_A_KGEqSJ7R2_2(.din(n907), .dout(n13542));
    jdff dff_B_QMTRnMAr5_1(.din(n895), .dout(n13546));
    jdff dff_B_Y2u8jKVw1_0(.din(G97), .dout(n13549));
    jdff dff_B_T69QBFzD0_3(.din(n891), .dout(n13552));
    jdff dff_B_QCLCXMcC4_3(.din(n13552), .dout(n13555));
    jdff dff_A_TnqZL3N03_0(.din(n13560), .dout(n13557));
    jdff dff_A_3WBdhEWs9_0(.din(n13563), .dout(n13560));
    jdff dff_A_vmr5aENK6_0(.din(n13566), .dout(n13563));
    jdff dff_A_R0cohlg94_0(.din(n888), .dout(n13566));
    jdff dff_A_azehETn11_2(.din(n13572), .dout(n13569));
    jdff dff_A_sclD5zdd4_2(.din(n13575), .dout(n13572));
    jdff dff_A_Iu8Av3AH3_2(.din(n888), .dout(n13575));
    jdff dff_B_wSeJvHvY2_1(.din(n876), .dout(n13579));
    jdff dff_B_Bzm4aaA47_0(.din(G47), .dout(n13582));
    jdff dff_B_G4bOJIy79_2(.din(n872), .dout(n13585));
    jdff dff_B_jr5IL4iN8_2(.din(n13585), .dout(n13588));
    jdff dff_A_yoOFCVWY1_0(.din(n13593), .dout(n13590));
    jdff dff_A_1ETaXjQF7_0(.din(n13596), .dout(n13593));
    jdff dff_A_70SR8ZAK3_0(.din(n13599), .dout(n13596));
    jdff dff_A_YppMUfdg6_0(.din(G4415), .dout(n13599));
    jdff dff_A_4OlQz9K68_0(.din(n13605), .dout(n13602));
    jdff dff_A_o4THdZ0n0_0(.din(n13608), .dout(n13605));
    jdff dff_A_plzDQIpw4_0(.din(n13611), .dout(n13608));
    jdff dff_A_b5VbxXny3_0(.din(n869), .dout(n13611));
    jdff dff_A_GO7S0n6C9_1(.din(n865), .dout(n13614));
    jdff dff_A_sqp9Njm17_1(.din(n13620), .dout(n13617));
    jdff dff_A_ayvScaaT2_1(.din(n818), .dout(n13620));
    jdff dff_A_dfPLcqln1_0(.din(n13626), .dout(n13623));
    jdff dff_A_kXBd5JXl6_0(.din(n13629), .dout(n13626));
    jdff dff_A_mjnJcMV75_0(.din(n13632), .dout(n13629));
    jdff dff_A_ttlRrIgr0_0(.din(n13635), .dout(n13632));
    jdff dff_A_0szJyxE99_0(.din(n13638), .dout(n13635));
    jdff dff_A_WJQMmuie9_0(.din(n13641), .dout(n13638));
    jdff dff_A_NBaBoVcZ7_0(.din(n794), .dout(n13641));
    jdff dff_A_IiN5JI5s8_0(.din(n13647), .dout(n13644));
    jdff dff_A_W5tLDX4L7_0(.din(n13650), .dout(n13647));
    jdff dff_A_7zf17ZJ46_0(.din(n13657), .dout(n13650));
    jdff dff_B_XJUEGaX61_2(.din(n761), .dout(n13654));
    jdff dff_B_cteXpGLd6_2(.din(n13654), .dout(n13657));
    jdff dff_A_rYZP6bhc0_0(.din(n13662), .dout(n13659));
    jdff dff_A_lXbV1seQ8_0(.din(n13665), .dout(n13662));
    jdff dff_A_OloIHzAR1_0(.din(n13668), .dout(n13665));
    jdff dff_A_T2HkbbHv0_0(.din(n13671), .dout(n13668));
    jdff dff_A_GTbnRU559_0(.din(n13674), .dout(n13671));
    jdff dff_A_mtPxmBZR7_0(.din(n757), .dout(n13674));
    jdff dff_A_p7UtFTKd6_1(.din(n13680), .dout(n13677));
    jdff dff_A_zUKcF8oA4_1(.din(n735), .dout(n13680));
    jdff dff_A_IxiQpLBq7_1(.din(n968), .dout(n13683));
    jdff dff_B_5hU4vHiZ8_1(.din(n953), .dout(n13687));
    jdff dff_B_0QEtDJod2_0(.din(G94), .dout(n13690));
    jdff dff_A_bIhfmbo90_0(.din(n13695), .dout(n13692));
    jdff dff_A_mdiprYfS9_0(.din(n13698), .dout(n13695));
    jdff dff_A_mb7C1QHa8_0(.din(n13701), .dout(n13698));
    jdff dff_A_J2qPaUXQ6_0(.din(G4405), .dout(n13701));
    jdff dff_A_xdlzvDjW9_0(.din(n949), .dout(n13704));
    jdff dff_A_x71sLdCq3_2(.din(n949), .dout(n13707));
    jdff dff_B_JjtPmCHB3_1(.din(n937), .dout(n13711));
    jdff dff_B_r7ZZahyA5_0(.din(G121), .dout(n13714));
    jdff dff_B_vh3Uguei7_2(.din(n933), .dout(n13717));
    jdff dff_B_2P58I5eT7_2(.din(n13717), .dout(n13720));
    jdff dff_A_vIvxKYgN7_0(.din(n13725), .dout(n13722));
    jdff dff_A_U9HEbJgo5_0(.din(n13728), .dout(n13725));
    jdff dff_A_K48xyCr10_0(.din(n13731), .dout(n13728));
    jdff dff_A_6pxG1Fq52_0(.din(G4410), .dout(n13731));
    jdff dff_A_5EbDisAo9_0(.din(n13737), .dout(n13734));
    jdff dff_A_IlnJLqiF5_0(.din(n1153), .dout(n13737));
    jdff dff_A_TzbzIG4M8_1(.din(n13743), .dout(n13740));
    jdff dff_A_9LNjiWNT4_1(.din(n13746), .dout(n13743));
    jdff dff_A_TO5rHO6z6_1(.din(n13749), .dout(n13746));
    jdff dff_A_xb40rgLK8_1(.din(n13752), .dout(n13749));
    jdff dff_A_3bsSzGkA5_1(.din(n13755), .dout(n13752));
    jdff dff_A_OL3a0SAZ9_1(.din(n13758), .dout(n13755));
    jdff dff_A_LqKGtasU1_1(.din(n13761), .dout(n13758));
    jdff dff_A_NdTm2IRH8_1(.din(n13764), .dout(n13761));
    jdff dff_A_UIODt7P69_1(.din(n13767), .dout(n13764));
    jdff dff_A_KJ01KZjo3_1(.din(n13770), .dout(n13767));
    jdff dff_A_HpI7Zu6e0_1(.din(n13773), .dout(n13770));
    jdff dff_A_nW4mItQv2_1(.din(n1153), .dout(n13773));
    jdff dff_B_Uq25joIQ0_1(.din(n1141), .dout(n13777));
    jdff dff_B_RbOHchf68_0(.din(G50), .dout(n13780));
    jdff dff_B_Th2dA3IE6_2(.din(n1137), .dout(n13783));
    jdff dff_B_clWffWiI2_2(.din(n13783), .dout(n13786));
    jdff dff_A_232Wcgk02_0(.din(n13791), .dout(n13788));
    jdff dff_A_h4ekmAyz2_0(.din(n13794), .dout(n13791));
    jdff dff_A_MAUrdrhs9_0(.din(n13797), .dout(n13794));
    jdff dff_A_vK1SaVCu5_0(.din(G4432), .dout(n13797));
    jdff dff_B_zr9TvNSk1_1(.din(n5354), .dout(n13801));
    jdff dff_B_Wfe7UT0x5_1(.din(n13801), .dout(n13804));
    jdff dff_B_KqnuhGgy5_1(.din(n13804), .dout(n13807));
    jdff dff_B_kmOdv2Jc1_1(.din(n13807), .dout(n13810));
    jdff dff_B_2iXF6qVS1_1(.din(n13810), .dout(n13813));
    jdff dff_B_VR6pvUXp8_1(.din(n13813), .dout(n13816));
    jdff dff_B_Z8lwB16C9_1(.din(n13816), .dout(n13819));
    jdff dff_B_aMHTsw7C1_1(.din(n13819), .dout(n13822));
    jdff dff_B_NpLUcPD67_1(.din(n13822), .dout(n13825));
    jdff dff_B_KBuj21bs4_1(.din(n13825), .dout(n13828));
    jdff dff_B_VzJehx210_1(.din(n13828), .dout(n13831));
    jdff dff_B_U7wBcD9C1_1(.din(n13831), .dout(n13834));
    jdff dff_B_iXzO8Qrp3_1(.din(n13834), .dout(n13837));
    jdff dff_B_KiFOFoT63_1(.din(n13837), .dout(n13840));
    jdff dff_B_3LGbg9YE5_1(.din(n13840), .dout(n13843));
    jdff dff_B_YN8G514S2_1(.din(n5461), .dout(n13846));
    jdff dff_B_Ot2uxS2b8_1(.din(n13846), .dout(n13849));
    jdff dff_B_LqYwp0DK4_1(.din(n13849), .dout(n13852));
    jdff dff_B_cC0B5eQI6_0(.din(n5609), .dout(n13855));
    jdff dff_B_mHSsPA474_1(.din(n5597), .dout(n13858));
    jdff dff_B_FqaGOYoO0_1(.din(n13858), .dout(n13861));
    jdff dff_B_29kOIiyV1_0(.din(n5583), .dout(n13864));
    jdff dff_B_AOo5QAEB4_0(.din(n13864), .dout(n13867));
    jdff dff_B_4WpU1ehT3_0(.din(n13867), .dout(n13870));
    jdff dff_B_fvd44txS3_0(.din(n13870), .dout(n13873));
    jdff dff_B_H5omkcwW9_0(.din(n13873), .dout(n13876));
    jdff dff_B_ryHRoTbl5_0(.din(n13876), .dout(n13879));
    jdff dff_B_tUAfxP7n4_0(.din(n13879), .dout(n13882));
    jdff dff_B_H0K3lUBb0_1(.din(n5552), .dout(n13885));
    jdff dff_B_xleab02x0_1(.din(n13885), .dout(n13888));
    jdff dff_B_tuMJqVnd7_1(.din(n13888), .dout(n13891));
    jdff dff_B_2bGQ9w4O4_1(.din(n13891), .dout(n13894));
    jdff dff_B_FuQFIgH88_1(.din(n13894), .dout(n13897));
    jdff dff_B_CIsA5jLb0_1(.din(n5555), .dout(n13900));
    jdff dff_B_hWdk9Lp90_1(.din(n13900), .dout(n13903));
    jdff dff_B_v2w6Y5368_1(.din(n13903), .dout(n13906));
    jdff dff_B_BaY2riKL9_1(.din(n13906), .dout(n13909));
    jdff dff_A_I1cbKSU18_1(.din(n13914), .dout(n13911));
    jdff dff_A_qiZJRdEy0_1(.din(n13917), .dout(n13914));
    jdff dff_A_riHYd6Xt7_1(.din(n13920), .dout(n13917));
    jdff dff_A_ybqhCZ7i9_1(.din(n5540), .dout(n13920));
    jdff dff_B_yaGAndz76_1(.din(n5524), .dout(n13924));
    jdff dff_A_qRjD17OP6_0(.din(n13929), .dout(n13926));
    jdff dff_A_dTfLmEGw5_0(.din(n13932), .dout(n13929));
    jdff dff_A_azqyXgUa4_0(.din(n13945), .dout(n13932));
    jdff dff_B_78qQyTrY1_2(.din(n3395), .dout(n13936));
    jdff dff_B_zFxoyLqs4_2(.din(n13936), .dout(n13939));
    jdff dff_B_yKeTjvzk6_2(.din(n13939), .dout(n13942));
    jdff dff_B_pfOlVf9R1_2(.din(n13942), .dout(n13945));
    jdff dff_A_T06DSO181_1(.din(n13950), .dout(n13947));
    jdff dff_A_bUccLvCp0_1(.din(n13953), .dout(n13950));
    jdff dff_A_4DWiGXIG0_1(.din(n5495), .dout(n13953));
    jdff dff_B_OGgUC0wS8_1(.din(n5472), .dout(n13957));
    jdff dff_B_REeW9gvT5_1(.din(n13957), .dout(n13960));
    jdff dff_B_psoXIpxT9_0(.din(n5479), .dout(n13963));
    jdff dff_B_jxRLmfFY1_0(.din(n13963), .dout(n13966));
    jdff dff_A_ZJHbP3dP6_0(.din(n13971), .dout(n13968));
    jdff dff_A_CBVuSnub1_0(.din(n13974), .dout(n13971));
    jdff dff_A_ZPEdoOs90_0(.din(n5465), .dout(n13974));
    jdff dff_A_vpVwBZGG7_1(.din(n3431), .dout(n13977));
    jdff dff_B_rjvqatEd1_1(.din(n5398), .dout(n13981));
    jdff dff_B_wHCiczz55_1(.din(n13981), .dout(n13984));
    jdff dff_B_JRcaNep85_1(.din(n13984), .dout(n13987));
    jdff dff_B_QUIsBXBh1_1(.din(n5439), .dout(n13990));
    jdff dff_B_j4SVgvbl0_1(.din(n13990), .dout(n13993));
    jdff dff_B_4Wj5yp2j5_1(.din(n5442), .dout(n13996));
    jdff dff_B_qAlmacbT0_1(.din(n13996), .dout(n13999));
    jdff dff_B_Lzk0vi2H7_1(.din(n13999), .dout(n14002));
    jdff dff_B_zd0yajDr0_1(.din(n14002), .dout(n14005));
    jdff dff_B_lbznyI1u1_1(.din(n14005), .dout(n14008));
    jdff dff_A_9qZgzsNs9_0(.din(n14013), .dout(n14010));
    jdff dff_A_TdBdHRL18_0(.din(n14016), .dout(n14013));
    jdff dff_A_9yFEB4Tk7_0(.din(n14019), .dout(n14016));
    jdff dff_A_6Yzdt3Ak2_0(.din(n4355), .dout(n14019));
    jdff dff_B_o9uY41Ac7_1(.din(n4317), .dout(n14023));
    jdff dff_A_cV1ghasb7_1(.din(n4298), .dout(n14025));
    jdff dff_A_MK79zHne4_0(.din(n14031), .dout(n14028));
    jdff dff_A_mqnS2Z4X2_0(.din(n14034), .dout(n14031));
    jdff dff_A_Pbera6bC7_0(.din(G3705), .dout(n14034));
    jdff dff_A_MV8HZdIY7_1(.din(n14040), .dout(n14037));
    jdff dff_A_wEcAMxBO0_1(.din(n14043), .dout(n14040));
    jdff dff_A_r4uRtzhq8_1(.din(G3705), .dout(n14043));
    jdff dff_A_kNbcT2hR0_0(.din(n14049), .dout(n14046));
    jdff dff_A_BXHabmH63_0(.din(n14052), .dout(n14049));
    jdff dff_A_CszolQZC5_0(.din(n14055), .dout(n14052));
    jdff dff_A_7BAqe4RH3_0(.din(n14058), .dout(n14055));
    jdff dff_A_sOHOWnrF9_0(.din(n482), .dout(n14058));
    jdff dff_B_qH8YMZAq3_0(.din(n463), .dout(n14062));
    jdff dff_A_zgO2fUiT9_1(.din(n14067), .dout(n14064));
    jdff dff_A_5wPFBUs39_1(.din(n4294), .dout(n14067));
    jdff dff_A_YU2PxwHh9_1(.din(n4291), .dout(n14070));
    jdff dff_A_u9w86PM44_2(.din(n14076), .dout(n14073));
    jdff dff_A_1fPZMeRr7_2(.din(n4291), .dout(n14076));
    jdff dff_B_P9QBsc5k9_0(.din(n4287), .dout(n14080));
    jdff dff_A_8VN8W2Jp5_0(.din(n14085), .dout(n14082));
    jdff dff_A_FFoxzIYb8_0(.din(n14088), .dout(n14085));
    jdff dff_A_fUSrVCF72_0(.din(G3717), .dout(n14088));
    jdff dff_A_UZkBPwWu9_1(.din(n14094), .dout(n14091));
    jdff dff_A_BRbsPw8B7_1(.din(n14097), .dout(n14094));
    jdff dff_A_SXnMlaJE4_1(.din(G3717), .dout(n14097));
    jdff dff_B_vA4D5r9z7_0(.din(n5431), .dout(n14101));
    jdff dff_B_wtTzXQZ68_0(.din(n14101), .dout(n14104));
    jdff dff_B_5MKJui9C7_0(.din(n14104), .dout(n14107));
    jdff dff_B_iWkXe2AJ4_0(.din(n14107), .dout(n14110));
    jdff dff_A_BxX42A2O3_1(.din(n14115), .dout(n14112));
    jdff dff_A_5gRjoGy61_1(.din(n14118), .dout(n14115));
    jdff dff_A_0WhToFMW5_1(.din(n5417), .dout(n14118));
    jdff dff_A_fDmLV9JP5_1(.din(n14124), .dout(n14121));
    jdff dff_A_wWhXJe5g4_1(.din(n14127), .dout(n14124));
    jdff dff_A_oqZruxcR8_1(.din(n14130), .dout(n14127));
    jdff dff_A_PKKRSAtR4_1(.din(n857), .dout(n14130));
    jdff dff_A_DOXs29d90_1(.din(n14136), .dout(n14133));
    jdff dff_A_X1w6X3UH9_1(.din(n14139), .dout(n14136));
    jdff dff_A_oJGc6wik0_1(.din(n14142), .dout(n14139));
    jdff dff_A_tvCdJFBR8_1(.din(n14145), .dout(n14142));
    jdff dff_A_bMRYvsgy9_1(.din(n5406), .dout(n14145));
    jdff dff_B_KeNprzu58_0(.din(n5402), .dout(n14149));
    jdff dff_A_sTYy0b9H1_1(.din(n707), .dout(n14151));
    jdff dff_A_sBgJxJKt1_1(.din(n695), .dout(n14154));
    jdff dff_B_5GHdNSKJ6_1(.din(n679), .dout(n14158));
    jdff dff_A_Oh3JpdHS7_0(.din(n14163), .dout(n14160));
    jdff dff_A_6M5Ju3np0_0(.din(n14166), .dout(n14163));
    jdff dff_A_5vS2KP6j3_0(.din(n14169), .dout(n14166));
    jdff dff_A_uuWTafWp4_0(.din(n14172), .dout(n14169));
    jdff dff_A_iqDMWr1G8_0(.din(n14175), .dout(n14172));
    jdff dff_A_2ORK7MJ96_0(.din(n14178), .dout(n14175));
    jdff dff_A_ruTERdd65_0(.din(n14181), .dout(n14178));
    jdff dff_A_PFrRtPz72_0(.din(n687), .dout(n14181));
    jdff dff_A_v76VSXqZ6_1(.din(n14187), .dout(n14184));
    jdff dff_A_JAoynUOq8_1(.din(n14190), .dout(n14187));
    jdff dff_A_rShiufyc4_1(.din(n14193), .dout(n14190));
    jdff dff_A_u95AvtUA5_1(.din(n14196), .dout(n14193));
    jdff dff_A_Mu6B6EbU7_1(.din(n687), .dout(n14196));
    jdff dff_A_8TRro6Rh2_0(.din(n14202), .dout(n14199));
    jdff dff_A_74cnW4016_0(.din(n671), .dout(n14202));
    jdff dff_A_qPeJQYRD1_0(.din(n667), .dout(n14205));
    jdff dff_A_9H4knwf08_1(.din(n667), .dout(n14208));
    jdff dff_A_AIM5S5t53_0(.din(n14214), .dout(n14211));
    jdff dff_A_5gSkhRnC7_0(.din(n14248), .dout(n14214));
    jdff dff_A_TbXBDE7v1_2(.din(n14220), .dout(n14217));
    jdff dff_A_68KSUdat4_2(.din(n14223), .dout(n14220));
    jdff dff_A_B6Cf6Acw1_2(.din(n14226), .dout(n14223));
    jdff dff_A_WFaEeLe79_2(.din(n14229), .dout(n14226));
    jdff dff_A_8oLxctnW1_2(.din(n14232), .dout(n14229));
    jdff dff_A_G9vcx2wh9_2(.din(n14235), .dout(n14232));
    jdff dff_A_36dz6SZj6_2(.din(n14238), .dout(n14235));
    jdff dff_A_PWZDMPJl4_2(.din(n14241), .dout(n14238));
    jdff dff_A_WWKtgBrA9_2(.din(n14244), .dout(n14241));
    jdff dff_A_b2eYmO4R5_2(.din(n14248), .dout(n14244));
    jdff dff_B_KidPtzUp6_3(.din(n452), .dout(n14248));
    jdff dff_A_wN9Pvajd7_2(.din(n14253), .dout(n14250));
    jdff dff_A_VW7Yj6298_2(.din(n647), .dout(n14253));
    jdff dff_A_DknvD8Cx1_1(.din(n627), .dout(n14256));
    jdff dff_A_hy19a9jk7_1(.din(n14262), .dout(n14259));
    jdff dff_A_UK6liytN6_1(.din(n14265), .dout(n14262));
    jdff dff_A_Y35dsLT03_1(.din(n14268), .dout(n14265));
    jdff dff_A_NW0XW22D6_1(.din(n14271), .dout(n14268));
    jdff dff_A_5hMSZaFC4_1(.din(n14274), .dout(n14271));
    jdff dff_A_JmylGvGX8_1(.din(n14277), .dout(n14274));
    jdff dff_A_GRIDOSq39_1(.din(n14280), .dout(n14277));
    jdff dff_A_0cOZA6cA9_1(.din(n14283), .dout(n14280));
    jdff dff_A_7gf8DVbR1_1(.din(n627), .dout(n14283));
    jdff dff_A_fn373POl2_2(.din(n14289), .dout(n14286));
    jdff dff_A_Agm25rVm7_2(.din(n14292), .dout(n14289));
    jdff dff_A_QTlFZtkZ7_2(.din(n627), .dout(n14292));
    jdff dff_B_ijgckosu9_1(.din(n605), .dout(n14296));
    jdff dff_B_sTsRkrCo0_1(.din(n14296), .dout(n14299));
    jdff dff_A_0fReXTFg6_0(.din(n14304), .dout(n14301));
    jdff dff_A_kVT3uzCz5_0(.din(n14307), .dout(n14304));
    jdff dff_A_MeHNMQtc8_0(.din(G3705), .dout(n14307));
    jdff dff_A_uSWqszjk6_0(.din(n602), .dout(n14310));
    jdff dff_A_sK9IWy2v7_0(.din(n471), .dout(n14313));
    jdff dff_A_MSVHLPQs9_1(.din(n14355), .dout(n14316));
    jdff dff_A_ZxAd4Hdj4_2(.din(n14322), .dout(n14319));
    jdff dff_A_xb6S6qui0_2(.din(n14325), .dout(n14322));
    jdff dff_A_nMiP9VN05_2(.din(n14328), .dout(n14325));
    jdff dff_A_fNiV9ITl2_2(.din(n14331), .dout(n14328));
    jdff dff_A_oaivMi756_2(.din(n14335), .dout(n14331));
    jdff dff_B_26IBZNyP1_3(.din(n583), .dout(n14335));
    jdff dff_A_5Sf6yYef6_0(.din(n459), .dout(n14337));
    jdff dff_A_DItjsZtr7_0(.din(n14343), .dout(n14340));
    jdff dff_A_aE5bhzcy6_0(.din(n14346), .dout(n14343));
    jdff dff_A_VMwgvIR75_0(.din(G41), .dout(n14346));
    jdff dff_A_1JWV0Pyl7_1(.din(G41), .dout(n14349));
    jdff dff_A_NVapzCBn3_1(.din(n579), .dout(n14352));
    jdff dff_A_iUgl4et14_0(.din(G3701), .dout(n14355));
    jdff dff_A_7xgMrx8f8_0(.din(n14361), .dout(n14358));
    jdff dff_A_L8oEP3pi9_0(.din(n14364), .dout(n14361));
    jdff dff_A_CM5uF7Q79_0(.din(n14367), .dout(n14364));
    jdff dff_A_jQm4POQd1_0(.din(n14370), .dout(n14367));
    jdff dff_A_ueMveMMH3_0(.din(n14373), .dout(n14370));
    jdff dff_A_7njmmzcU3_0(.din(n14376), .dout(n14373));
    jdff dff_A_JivydptM7_0(.din(n14379), .dout(n14376));
    jdff dff_A_FHod2HfN7_0(.din(n14382), .dout(n14379));
    jdff dff_A_n9lY1H8r0_0(.din(n14385), .dout(n14382));
    jdff dff_A_DsbOikcy1_0(.din(n14388), .dout(n14385));
    jdff dff_A_QLd0u7Pk2_0(.din(n14404), .dout(n14388));
    jdff dff_A_t2vvxLIv2_2(.din(n14404), .dout(n14391));
    jdff dff_B_P9oTzFiG0_3(.din(n576), .dout(n14395));
    jdff dff_B_pLDP2Vqt9_3(.din(n14395), .dout(n14398));
    jdff dff_B_TBNi1hV02_3(.din(n14398), .dout(n14401));
    jdff dff_B_mLOxX17m9_3(.din(n14401), .dout(n14404));
    jdff dff_A_X2hJZbNH9_1(.din(n14409), .dout(n14406));
    jdff dff_A_rTCYYuTb9_1(.din(n14412), .dout(n14409));
    jdff dff_A_MJsQ6nGm6_1(.din(n14415), .dout(n14412));
    jdff dff_A_BpQsFthV1_1(.din(n14418), .dout(n14415));
    jdff dff_A_ms5Q6tOQ7_1(.din(G4526), .dout(n14418));
    jdff dff_A_9PM9D7hK7_1(.din(n14424), .dout(n14421));
    jdff dff_A_WKlATLgI7_1(.din(n14427), .dout(n14424));
    jdff dff_A_fy6nSdI54_1(.din(n14430), .dout(n14427));
    jdff dff_A_PgvoQJuA2_1(.din(n14433), .dout(n14430));
    jdff dff_A_UdbUjPSL4_1(.din(n14436), .dout(n14433));
    jdff dff_A_VpOZSvnH0_1(.din(n14439), .dout(n14436));
    jdff dff_A_PRsLHwbW7_1(.din(n14442), .dout(n14439));
    jdff dff_A_VDwri5zt0_1(.din(n14445), .dout(n14442));
    jdff dff_A_6LaLYoZz7_1(.din(n14448), .dout(n14445));
    jdff dff_A_XDKhkYet6_1(.din(n14451), .dout(n14448));
    jdff dff_A_DLlCpuQU8_1(.din(n14454), .dout(n14451));
    jdff dff_A_Vvn0hPCn1_1(.din(n14457), .dout(n14454));
    jdff dff_A_YOC4rDdX5_1(.din(n14460), .dout(n14457));
    jdff dff_A_2bAkTEUW4_1(.din(n14463), .dout(n14460));
    jdff dff_A_d505jNZO2_1(.din(G4526), .dout(n14463));
    jdff dff_A_9M9WJaAl2_2(.din(n14469), .dout(n14466));
    jdff dff_A_vPudiIHb7_2(.din(n14472), .dout(n14469));
    jdff dff_A_nuR6vZS55_2(.din(n14475), .dout(n14472));
    jdff dff_A_u6pCXeVY1_2(.din(n14478), .dout(n14475));
    jdff dff_A_FlXCStQ04_2(.din(n14481), .dout(n14478));
    jdff dff_A_CGzIPUJQ0_2(.din(G4526), .dout(n14481));
    jdff dff_A_fptldo2Z1_1(.din(n573), .dout(n14484));
    jdff dff_A_UfqrjIig3_2(.din(n14490), .dout(n14487));
    jdff dff_A_XjEUdPLg8_2(.din(n14493), .dout(n14490));
    jdff dff_A_8zOw0JFN9_2(.din(n573), .dout(n14493));
    jdff dff_A_ujmd7dth2_1(.din(n548), .dout(n14496));
    jdff dff_A_fxhrM4H85_2(.din(n14502), .dout(n14499));
    jdff dff_A_QCnVwtnx0_2(.din(n548), .dout(n14502));
    jdff dff_A_NsVQY6dY5_0(.din(n14508), .dout(n14505));
    jdff dff_A_tlg9K5ml4_0(.din(n14511), .dout(n14508));
    jdff dff_A_uFNboZ7w4_0(.din(n544), .dout(n14511));
    jdff dff_A_KIbxWG680_1(.din(n14517), .dout(n14514));
    jdff dff_A_nsY4tZgM7_1(.din(n14520), .dout(n14517));
    jdff dff_A_T4oDNzeA1_1(.din(n14523), .dout(n14520));
    jdff dff_A_lAUA7D2V6_1(.din(n14526), .dout(n14523));
    jdff dff_A_E1HN2sYi3_1(.din(n14529), .dout(n14526));
    jdff dff_A_gi09h5j40_1(.din(n14532), .dout(n14529));
    jdff dff_A_AiXPINR31_1(.din(n14535), .dout(n14532));
    jdff dff_A_c0J9rYi81_1(.din(n14538), .dout(n14535));
    jdff dff_A_wDZaEiJY1_1(.din(n14541), .dout(n14538));
    jdff dff_A_YFnBr3dz8_1(.din(n14544), .dout(n14541));
    jdff dff_A_rLEOKtgO7_1(.din(n14547), .dout(n14544));
    jdff dff_A_Y7XVqhIw2_1(.din(n14550), .dout(n14547));
    jdff dff_A_2xgicKFQ5_1(.din(n14553), .dout(n14550));
    jdff dff_A_k9uy9nRV1_1(.din(n544), .dout(n14553));
    jdff dff_A_lxXH7riZ8_2(.din(n14559), .dout(n14556));
    jdff dff_A_isE6yyPm5_2(.din(n14562), .dout(n14559));
    jdff dff_A_yXdKgWiP7_2(.din(n14565), .dout(n14562));
    jdff dff_A_JeDlUWyh1_2(.din(n544), .dout(n14565));
    jdff dff_A_pzV3NkDf7_2(.din(n537), .dout(n14568));
    jdff dff_A_Y5zX2Jn48_1(.din(n14574), .dout(n14571));
    jdff dff_A_Awt1ZS5b6_1(.din(n14577), .dout(n14574));
    jdff dff_A_f4GZOwov5_1(.din(n14580), .dout(n14577));
    jdff dff_A_MjfUwtZn7_1(.din(G3717), .dout(n14580));
    jdff dff_A_QzaHcTNw8_1(.din(n14586), .dout(n14583));
    jdff dff_A_xNRUv05R1_1(.din(n14589), .dout(n14586));
    jdff dff_A_zfdkBFJC6_1(.din(n14592), .dout(n14589));
    jdff dff_A_qxygZq8W6_1(.din(n14595), .dout(n14592));
    jdff dff_A_viZejYLv6_1(.din(n14598), .dout(n14595));
    jdff dff_A_xBUmBKqi3_1(.din(n14601), .dout(n14598));
    jdff dff_A_aPEOWLYQ7_1(.din(n519), .dout(n14601));
    jdff dff_A_sCnlMVHi9_2(.din(n519), .dout(n14604));
    jdff dff_A_O1OWSXsT9_1(.din(n14610), .dout(n14607));
    jdff dff_A_O09Sv88N4_1(.din(n14613), .dout(n14610));
    jdff dff_A_myC7Op7m9_1(.din(n14616), .dout(n14613));
    jdff dff_A_lVTS1oef4_1(.din(n14619), .dout(n14616));
    jdff dff_A_1F408bzs9_1(.din(n14622), .dout(n14619));
    jdff dff_A_OvmsPZXt0_1(.din(n519), .dout(n14622));
    jdff dff_A_kGUs8Ygl7_2(.din(n14628), .dout(n14625));
    jdff dff_A_2PKsHjju1_2(.din(n14631), .dout(n14628));
    jdff dff_A_O3pZ11if4_2(.din(n14634), .dout(n14631));
    jdff dff_A_G4vODcwN8_2(.din(n14637), .dout(n14634));
    jdff dff_A_BfEahovQ1_2(.din(n14640), .dout(n14637));
    jdff dff_A_IPFhCnFv0_2(.din(n14643), .dout(n14640));
    jdff dff_A_bUV5ZSHt7_2(.din(n14646), .dout(n14643));
    jdff dff_A_nvfLFF5L2_2(.din(n519), .dout(n14646));
    jdff dff_A_siTTxv4V7_1(.din(G18), .dout(n14649));
    jdff dff_A_7OWMYmKc6_1(.din(n14655), .dout(n14652));
    jdff dff_A_rkwUqV5s2_1(.din(n497), .dout(n14655));
    jdff dff_A_A0c8EOMR5_0(.din(n14661), .dout(n14658));
    jdff dff_A_oT3PokxN3_0(.din(n14664), .dout(n14661));
    jdff dff_A_WhROGiIe9_0(.din(G3723), .dout(n14664));
    jdff dff_A_9SzzS9C42_2(.din(n14670), .dout(n14667));
    jdff dff_A_9IeOG2S09_2(.din(n14673), .dout(n14670));
    jdff dff_A_heDmG2sM6_2(.din(G3723), .dout(n14673));
    jdff dff_B_IDWVY7Qp0_0(.din(n5382), .dout(n14677));
    jdff dff_B_HKpF9qpd8_0(.din(n14677), .dout(n14680));
    jdff dff_B_glvbTKBU9_0(.din(n14680), .dout(n14683));
    jdff dff_B_M0X3wcWY0_0(.din(n14683), .dout(n14686));
    jdff dff_B_XYYkBOti0_0(.din(n14686), .dout(n14689));
    jdff dff_A_bxT6hRH78_0(.din(n14694), .dout(n14691));
    jdff dff_A_n78Njfyl6_0(.din(n14697), .dout(n14694));
    jdff dff_A_c3nTc5gs1_0(.din(n14700), .dout(n14697));
    jdff dff_A_J4TEJD776_0(.din(n14703), .dout(n14700));
    jdff dff_A_N99NFegW8_0(.din(n5379), .dout(n14703));
    jdff dff_A_srNQeTzb1_2(.din(n14709), .dout(n14706));
    jdff dff_A_O97I3AvY0_2(.din(n14712), .dout(n14709));
    jdff dff_A_epmZ90cf7_2(.din(n14715), .dout(n14712));
    jdff dff_A_ORIrRChN2_2(.din(n14718), .dout(n14715));
    jdff dff_A_nkNKKBf63_2(.din(n14721), .dout(n14718));
    jdff dff_A_ua17eETB6_2(.din(n3479), .dout(n14721));
    jdff dff_A_Z8dSX2lB7_2(.din(n14727), .dout(n14724));
    jdff dff_A_N77G8Ucv9_2(.din(n14730), .dout(n14727));
    jdff dff_A_7gOmAGjr3_2(.din(n14733), .dout(n14730));
    jdff dff_A_ZIz1Wk376_2(.din(n14736), .dout(n14733));
    jdff dff_A_a9jK7E3F3_2(.din(n14739), .dout(n14736));
    jdff dff_A_jj0BgXic4_2(.din(n14742), .dout(n14739));
    jdff dff_A_M2sNt5aJ0_2(.din(n14745), .dout(n14742));
    jdff dff_A_SuogiHgF1_2(.din(n732), .dout(n14745));
    jdff dff_B_8HgM9npp3_1(.din(n5357), .dout(n14749));
    jdff dff_A_WQ7rGcbR6_1(.din(n14754), .dout(n14751));
    jdff dff_A_7KKGRqGr4_1(.din(n829), .dout(n14754));
    jdff dff_A_Eo8pjj496_0(.din(n853), .dout(n14757));
    jdff dff_A_iiFUvMV99_1(.din(n14763), .dout(n14760));
    jdff dff_A_e9pqetUX0_1(.din(n14766), .dout(n14763));
    jdff dff_A_BI8gDIYZ4_1(.din(n14769), .dout(n14766));
    jdff dff_A_c1RFncXA6_1(.din(n14772), .dout(n14769));
    jdff dff_A_UFFdpIeU1_1(.din(n849), .dout(n14772));
    jdff dff_A_Ei9lQM4A3_1(.din(n14778), .dout(n14775));
    jdff dff_A_VNLWXNkb2_1(.din(n14781), .dout(n14778));
    jdff dff_A_EnvjuNp65_1(.din(n14784), .dout(n14781));
    jdff dff_A_UKT2WkAc4_1(.din(n14787), .dout(n14784));
    jdff dff_A_x11vc7E51_1(.din(n14790), .dout(n14787));
    jdff dff_A_3lQu6qF98_1(.din(n14793), .dout(n14790));
    jdff dff_A_v5z2xYqi5_1(.din(n841), .dout(n14793));
    jdff dff_A_Pa5T8Khv1_0(.din(n14799), .dout(n14796));
    jdff dff_A_8LcK8OjW1_0(.din(n14802), .dout(n14799));
    jdff dff_A_FABQIxU61_0(.din(G3729), .dout(n14802));
    jdff dff_A_oU161Ncu3_2(.din(n14808), .dout(n14805));
    jdff dff_A_PsQowceb7_2(.din(n14811), .dout(n14808));
    jdff dff_A_aF5AZzhG1_2(.din(G3729), .dout(n14811));
    jdff dff_B_h21CaGwJ6_1(.din(n710), .dout(n14815));
    jdff dff_B_l6O1nGen5_1(.din(n14815), .dout(n14818));
    jdff dff_B_aoQ4cO6G4_2(.din(n837), .dout(n14821));
    jdff dff_A_Ez3fDP7O2_0(.din(G18), .dout(n14823));
    jdff dff_A_LnfPSjCj1_2(.din(G18), .dout(n14826));
    jdff dff_A_5wOY19y38_0(.din(n14832), .dout(n14829));
    jdff dff_A_TwEkicrX2_0(.din(n14835), .dout(n14832));
    jdff dff_A_HfR9wvXH0_0(.din(G3737), .dout(n14835));
    jdff dff_A_xFFZkzla9_1(.din(n14841), .dout(n14838));
    jdff dff_A_l1nYXMXi6_1(.din(n14844), .dout(n14841));
    jdff dff_A_S887kdNf8_1(.din(n14847), .dout(n14844));
    jdff dff_A_ldZ1KY7c8_1(.din(n14850), .dout(n14847));
    jdff dff_A_YkCQntDW9_1(.din(n14853), .dout(n14850));
    jdff dff_A_41bqDbRo2_1(.din(n833), .dout(n14853));
    jdff dff_A_fSaZrFse3_2(.din(n833), .dout(n14856));
    jdff dff_A_zlrFOdIx5_2(.din(n14862), .dout(n14859));
    jdff dff_A_Oh7A8BMG5_2(.din(n14865), .dout(n14862));
    jdff dff_A_Mbxmu5IA8_2(.din(n794), .dout(n14865));
    jdff dff_A_7nHzeAQE8_0(.din(n14871), .dout(n14868));
    jdff dff_A_i8MxtEqX8_0(.din(n14874), .dout(n14871));
    jdff dff_A_gJo61eAj1_0(.din(n14877), .dout(n14874));
    jdff dff_A_jCSaDnGt3_0(.din(n14881), .dout(n14877));
    jdff dff_B_PlwNksKA7_2(.din(n790), .dout(n14881));
    jdff dff_A_UiYgcqjj0_0(.din(n14886), .dout(n14883));
    jdff dff_A_4K5YfUEq1_0(.din(n14889), .dout(n14886));
    jdff dff_A_qYFnchSb5_0(.din(n14892), .dout(n14889));
    jdff dff_A_qg2u1FFT9_0(.din(n783), .dout(n14892));
    jdff dff_A_NME46QeS8_1(.din(G18), .dout(n14895));
    jdff dff_A_hrTl2yRI2_0(.din(n14901), .dout(n14898));
    jdff dff_A_ZBdNzVag3_0(.din(n14904), .dout(n14901));
    jdff dff_A_6QumpSRY2_0(.din(G3749), .dout(n14904));
    jdff dff_A_zAZyEvqU4_1(.din(n14910), .dout(n14907));
    jdff dff_A_S2y8jGwy7_1(.din(n14913), .dout(n14910));
    jdff dff_A_eBkTexpT7_1(.din(n14916), .dout(n14913));
    jdff dff_A_1GyyuEdD3_1(.din(n14919), .dout(n14916));
    jdff dff_A_7Jc62E2n3_1(.din(n14922), .dout(n14919));
    jdff dff_A_Pgbhg1V60_1(.din(n14925), .dout(n14922));
    jdff dff_A_yGPNZGOU3_1(.din(n14932), .dout(n14925));
    jdff dff_A_DQ9xXhsI5_2(.din(n14932), .dout(n14928));
    jdff dff_B_JFMYzIFG6_3(.din(n810), .dout(n14932));
    jdff dff_B_44dd0rRk9_1(.din(n798), .dout(n14935));
    jdff dff_B_hcyQBnBz9_0(.din(G124), .dout(n14938));
    jdff dff_A_JffuGsQJ7_2(.din(G18), .dout(n14940));
    jdff dff_A_cXHyq6OK4_1(.din(G18), .dout(n14943));
    jdff dff_A_984qphLh4_2(.din(G18), .dout(n14946));
    jdff dff_A_n0yhwvps7_2(.din(G18), .dout(n14949));
    jdff dff_A_yxDm7fX93_0(.din(n14958), .dout(n14952));
    jdff dff_A_j8emn42k0_1(.din(n14958), .dout(n14955));
    jdff dff_A_Mop6iPGY8_0(.din(n14961), .dout(n14958));
    jdff dff_A_WIVPdZkN8_0(.din(n14964), .dout(n14961));
    jdff dff_A_vVahhG232_0(.din(G3743), .dout(n14964));
    jdff dff_A_hSoXGY9p8_1(.din(n4294), .dout(n14967));
    jdff dff_A_rsI4cXCp7_2(.din(n14973), .dout(n14970));
    jdff dff_A_s7ItAJyX3_2(.din(n14976), .dout(n14973));
    jdff dff_A_EagitJIb6_2(.din(n14979), .dout(n14976));
    jdff dff_A_GOOt5XX88_2(.din(n573), .dout(n14979));
    jdff dff_B_8A4vRwvi3_1(.din(n551), .dout(n14983));
    jdff dff_B_Lmpe7ff84_1(.din(n14983), .dout(n14986));
    jdff dff_A_g8Yd2so27_0(.din(G18), .dout(n14988));
    jdff dff_A_e7OVtupO2_2(.din(G18), .dout(n14991));
    jdff dff_A_DIwKuMg99_0(.din(n14997), .dout(n14994));
    jdff dff_A_7OXfBqVa7_0(.din(n15000), .dout(n14997));
    jdff dff_A_nDhm2kq96_0(.din(G3711), .dout(n15000));
    jdff dff_A_Lj9zbcUa6_1(.din(n5628), .dout(n15003));
    jdff dff_A_ywehXCUa1_0(.din(n15003), .dout(n15006));
    jdff dff_A_hpZHBmGS3_0(.din(n15006), .dout(n15009));
    jdff dff_A_sfSARdCR5_0(.din(n15009), .dout(n15012));
    jdff dff_A_nBd1YF5H6_0(.din(n15012), .dout(n15015));
    jdff dff_A_M3jxpyfz4_0(.din(n15015), .dout(n15018));
    jdff dff_A_PFYmG4hZ5_0(.din(n15018), .dout(n15021));
    jdff dff_A_eiOEw5107_0(.din(n15021), .dout(n15024));
    jdff dff_A_YXbuUOnv8_0(.din(n15024), .dout(n15027));
    jdff dff_A_XCVPSGM95_0(.din(n15027), .dout(n15030));
    jdff dff_A_ZX6fe0lf9_0(.din(n15030), .dout(n15033));
    jdff dff_A_uWzz0TLL9_0(.din(n15033), .dout(n15036));
    jdff dff_A_EfuQuOuc9_0(.din(n15036), .dout(n15039));
    jdff dff_A_hgvHOupC1_0(.din(n15039), .dout(n15042));
    jdff dff_A_wtqYKzGc1_0(.din(n15042), .dout(n15045));
    jdff dff_A_7XduDj1U7_0(.din(n15045), .dout(n15048));
    jdff dff_A_A7GNF2XS4_0(.din(n15048), .dout(n15051));
    jdff dff_A_CEmI8Lxr6_0(.din(n15051), .dout(n15054));
    jdff dff_A_5PrQnNSk7_0(.din(n15054), .dout(n15057));
    jdff dff_A_2sPFJEsh9_0(.din(n15057), .dout(n15060));
    jdff dff_A_9b6dwdyC6_0(.din(n15060), .dout(n15063));
    jdff dff_A_aZWE634o2_0(.din(n15063), .dout(n15066));
    jdff dff_A_BEWgpPnm6_0(.din(n15066), .dout(n15069));
    jdff dff_A_MNU1QNoV9_0(.din(n15069), .dout(n15072));
    jdff dff_A_LX11k00f7_0(.din(n15072), .dout(n15075));
    jdff dff_A_iNnnpCsJ0_0(.din(n15075), .dout(G2));
    jdff dff_A_bKUyBodi8_1(.din(n5631), .dout(n15081));
    jdff dff_A_v285L7xL5_0(.din(n15081), .dout(n15084));
    jdff dff_A_rUDYX13a7_0(.din(n15084), .dout(n15087));
    jdff dff_A_4tDnO5nJ5_0(.din(n15087), .dout(n15090));
    jdff dff_A_h0o3o1xr8_0(.din(n15090), .dout(n15093));
    jdff dff_A_OYeP2yOu7_0(.din(n15093), .dout(n15096));
    jdff dff_A_uKTFaQJ35_0(.din(n15096), .dout(n15099));
    jdff dff_A_eUrAMSmT5_0(.din(n15099), .dout(n15102));
    jdff dff_A_yHDXYlgH7_0(.din(n15102), .dout(n15105));
    jdff dff_A_TMxFEqwz9_0(.din(n15105), .dout(n15108));
    jdff dff_A_tVliGP8n1_0(.din(n15108), .dout(n15111));
    jdff dff_A_nt2KtYtx8_0(.din(n15111), .dout(n15114));
    jdff dff_A_8p4nqR3a8_0(.din(n15114), .dout(n15117));
    jdff dff_A_BKsLBISq9_0(.din(n15117), .dout(n15120));
    jdff dff_A_YZsBBmMq7_0(.din(n15120), .dout(n15123));
    jdff dff_A_lSdz3bWj1_0(.din(n15123), .dout(n15126));
    jdff dff_A_C3PejpNi8_0(.din(n15126), .dout(n15129));
    jdff dff_A_1tqrNl0d8_0(.din(n15129), .dout(n15132));
    jdff dff_A_7dJI4oOY1_0(.din(n15132), .dout(n15135));
    jdff dff_A_JG1vOCvW3_0(.din(n15135), .dout(n15138));
    jdff dff_A_MdcULH4j6_0(.din(n15138), .dout(n15141));
    jdff dff_A_rnzCGt0E3_0(.din(n15141), .dout(n15144));
    jdff dff_A_LpNmMvXA5_0(.din(n15144), .dout(n15147));
    jdff dff_A_8pPVXDib0_0(.din(n15147), .dout(n15150));
    jdff dff_A_wOKaWCPZ0_0(.din(n15150), .dout(n15153));
    jdff dff_A_4RoSXpPO6_0(.din(n15153), .dout(G3));
    jdff dff_A_ykkR7BTX5_1(.din(n5634), .dout(n15159));
    jdff dff_A_EpDTHM1d0_0(.din(n15159), .dout(n15162));
    jdff dff_A_brZ3xIhE2_0(.din(n15162), .dout(n15165));
    jdff dff_A_mqLJ9KNt3_0(.din(n15165), .dout(n15168));
    jdff dff_A_ToyAXf8w3_0(.din(n15168), .dout(n15171));
    jdff dff_A_LuN51aD65_0(.din(n15171), .dout(n15174));
    jdff dff_A_XH5w1yxR1_0(.din(n15174), .dout(n15177));
    jdff dff_A_3nAWI0la7_0(.din(n15177), .dout(n15180));
    jdff dff_A_ZRPZAtOX5_0(.din(n15180), .dout(n15183));
    jdff dff_A_c7HJVQT50_0(.din(n15183), .dout(n15186));
    jdff dff_A_7wrTDaOS1_0(.din(n15186), .dout(n15189));
    jdff dff_A_VAz7b4Gi5_0(.din(n15189), .dout(n15192));
    jdff dff_A_6SFwqig01_0(.din(n15192), .dout(n15195));
    jdff dff_A_IOVpHB1G7_0(.din(n15195), .dout(n15198));
    jdff dff_A_RyEOauqP4_0(.din(n15198), .dout(n15201));
    jdff dff_A_6ZTgUnNV6_0(.din(n15201), .dout(n15204));
    jdff dff_A_VThvqpi84_0(.din(n15204), .dout(n15207));
    jdff dff_A_K5pe7vPB7_0(.din(n15207), .dout(n15210));
    jdff dff_A_K3AtxB7M4_0(.din(n15210), .dout(n15213));
    jdff dff_A_A9TpM5qa7_0(.din(n15213), .dout(n15216));
    jdff dff_A_jhEdUKFC0_0(.din(n15216), .dout(n15219));
    jdff dff_A_Coq6BMl46_0(.din(n15219), .dout(n15222));
    jdff dff_A_hv1lnQ6D7_0(.din(n15222), .dout(n15225));
    jdff dff_A_AVvk53uu6_0(.din(n15225), .dout(n15228));
    jdff dff_A_zRW9CPGS3_0(.din(n15228), .dout(n15231));
    jdff dff_A_teD8M2gk8_0(.din(n15231), .dout(G450));
    jdff dff_A_5BZl4JPk1_1(.din(n5637), .dout(n15237));
    jdff dff_A_PIJL7jhG7_0(.din(n15237), .dout(n15240));
    jdff dff_A_FnQYp6ul2_0(.din(n15240), .dout(n15243));
    jdff dff_A_i4X35nkB3_0(.din(n15243), .dout(n15246));
    jdff dff_A_X1aQbOx61_0(.din(n15246), .dout(n15249));
    jdff dff_A_Tz9Ll54v1_0(.din(n15249), .dout(n15252));
    jdff dff_A_N9m2u4dY9_0(.din(n15252), .dout(n15255));
    jdff dff_A_xSNJ1BTN8_0(.din(n15255), .dout(n15258));
    jdff dff_A_4kKgQLrM4_0(.din(n15258), .dout(n15261));
    jdff dff_A_h1PCNJ8L1_0(.din(n15261), .dout(n15264));
    jdff dff_A_LWfeLkUz3_0(.din(n15264), .dout(n15267));
    jdff dff_A_XFMDUF8M2_0(.din(n15267), .dout(n15270));
    jdff dff_A_USC1GW618_0(.din(n15270), .dout(n15273));
    jdff dff_A_f0pTPOsW2_0(.din(n15273), .dout(n15276));
    jdff dff_A_6dARqQ2a3_0(.din(n15276), .dout(n15279));
    jdff dff_A_svgvGrkX3_0(.din(n15279), .dout(n15282));
    jdff dff_A_qZKJUXgl6_0(.din(n15282), .dout(n15285));
    jdff dff_A_aw2zk8MI0_0(.din(n15285), .dout(n15288));
    jdff dff_A_FnH9o1Tb4_0(.din(n15288), .dout(n15291));
    jdff dff_A_eOlFEr7z1_0(.din(n15291), .dout(n15294));
    jdff dff_A_bVOZMBm67_0(.din(n15294), .dout(n15297));
    jdff dff_A_14yrAvKb5_0(.din(n15297), .dout(n15300));
    jdff dff_A_lkSNs8He8_0(.din(n15300), .dout(n15303));
    jdff dff_A_vvfK3lCp9_0(.din(n15303), .dout(n15306));
    jdff dff_A_v2yELCdE9_0(.din(n15306), .dout(n15309));
    jdff dff_A_3PEnCtBv8_0(.din(n15309), .dout(G448));
    jdff dff_A_lpzyHoCB3_1(.din(n5640), .dout(n15315));
    jdff dff_A_oDbiegJ57_0(.din(n15315), .dout(n15318));
    jdff dff_A_Hhzsciea1_0(.din(n15318), .dout(n15321));
    jdff dff_A_YwcUCT5Z8_0(.din(n15321), .dout(n15324));
    jdff dff_A_n817RTmT7_0(.din(n15324), .dout(n15327));
    jdff dff_A_nxrsyCh59_0(.din(n15327), .dout(n15330));
    jdff dff_A_7voHvPDZ3_0(.din(n15330), .dout(n15333));
    jdff dff_A_UqJ05x1V3_0(.din(n15333), .dout(n15336));
    jdff dff_A_5n1Pyn2d8_0(.din(n15336), .dout(n15339));
    jdff dff_A_u8dNkfQO1_0(.din(n15339), .dout(n15342));
    jdff dff_A_1yUxlyNT3_0(.din(n15342), .dout(n15345));
    jdff dff_A_0N75zwGr0_0(.din(n15345), .dout(n15348));
    jdff dff_A_1rln8GPN5_0(.din(n15348), .dout(n15351));
    jdff dff_A_9yOpdUW36_0(.din(n15351), .dout(n15354));
    jdff dff_A_FdeNCbK17_0(.din(n15354), .dout(n15357));
    jdff dff_A_SWqyt6at7_0(.din(n15357), .dout(n15360));
    jdff dff_A_JZ3Vvpni9_0(.din(n15360), .dout(n15363));
    jdff dff_A_i8ZCNfUd9_0(.din(n15363), .dout(n15366));
    jdff dff_A_0lmWSpFa0_0(.din(n15366), .dout(n15369));
    jdff dff_A_3j3Lnv4x0_0(.din(n15369), .dout(n15372));
    jdff dff_A_fqLPO4jp5_0(.din(n15372), .dout(n15375));
    jdff dff_A_y7pZHwE02_0(.din(n15375), .dout(n15378));
    jdff dff_A_sUDznM3e7_0(.din(n15378), .dout(n15381));
    jdff dff_A_4KUrw3ax4_0(.din(n15381), .dout(n15384));
    jdff dff_A_9XzUPOPa3_0(.din(n15384), .dout(n15387));
    jdff dff_A_LrxXiihK5_0(.din(n15387), .dout(G444));
    jdff dff_A_rEh14yc44_1(.din(n5643), .dout(n15393));
    jdff dff_A_WHwPWy2u7_0(.din(n15393), .dout(n15396));
    jdff dff_A_u3PY3FCf3_0(.din(n15396), .dout(n15399));
    jdff dff_A_IAxjzWOd2_0(.din(n15399), .dout(n15402));
    jdff dff_A_tkmeiAQe7_0(.din(n15402), .dout(n15405));
    jdff dff_A_E7tDs0jO9_0(.din(n15405), .dout(n15408));
    jdff dff_A_PvvokCLV7_0(.din(n15408), .dout(n15411));
    jdff dff_A_UjGj5Ycc8_0(.din(n15411), .dout(n15414));
    jdff dff_A_1F61HQYx6_0(.din(n15414), .dout(n15417));
    jdff dff_A_ixNBkNpN0_0(.din(n15417), .dout(n15420));
    jdff dff_A_VrxocDes2_0(.din(n15420), .dout(n15423));
    jdff dff_A_wT6ECk2p1_0(.din(n15423), .dout(n15426));
    jdff dff_A_Oq07xbS00_0(.din(n15426), .dout(n15429));
    jdff dff_A_2CA241fZ3_0(.din(n15429), .dout(n15432));
    jdff dff_A_nDr6tM732_0(.din(n15432), .dout(n15435));
    jdff dff_A_zvMdIWmt8_0(.din(n15435), .dout(n15438));
    jdff dff_A_0BcZrKz53_0(.din(n15438), .dout(n15441));
    jdff dff_A_XcAMIdEi2_0(.din(n15441), .dout(n15444));
    jdff dff_A_EK9vnq0r5_0(.din(n15444), .dout(n15447));
    jdff dff_A_M64VN9N93_0(.din(n15447), .dout(n15450));
    jdff dff_A_PXIRguxK4_0(.din(n15450), .dout(n15453));
    jdff dff_A_1dGvCvkD2_0(.din(n15453), .dout(n15456));
    jdff dff_A_aGWXHUdU9_0(.din(n15456), .dout(n15459));
    jdff dff_A_oKOQuPsj7_0(.din(n15459), .dout(n15462));
    jdff dff_A_PMovNCDZ8_0(.din(n15462), .dout(n15465));
    jdff dff_A_RUro9E0k3_0(.din(n15465), .dout(G442));
    jdff dff_A_Qb2jOS5o0_1(.din(n5646), .dout(n15471));
    jdff dff_A_tIWBtJn27_0(.din(n15471), .dout(n15474));
    jdff dff_A_OA0wYm853_0(.din(n15474), .dout(n15477));
    jdff dff_A_G3QHnqgV6_0(.din(n15477), .dout(n15480));
    jdff dff_A_gFSGMReh4_0(.din(n15480), .dout(n15483));
    jdff dff_A_XM9QDtR27_0(.din(n15483), .dout(n15486));
    jdff dff_A_F7xGfi0s8_0(.din(n15486), .dout(n15489));
    jdff dff_A_OWvvromt7_0(.din(n15489), .dout(n15492));
    jdff dff_A_PX9v89ft9_0(.din(n15492), .dout(n15495));
    jdff dff_A_piwCPmhX3_0(.din(n15495), .dout(n15498));
    jdff dff_A_NO5XX01t3_0(.din(n15498), .dout(n15501));
    jdff dff_A_5f7o3nb18_0(.din(n15501), .dout(n15504));
    jdff dff_A_2oEv4P7U4_0(.din(n15504), .dout(n15507));
    jdff dff_A_SlzhVd5S8_0(.din(n15507), .dout(n15510));
    jdff dff_A_cSzB5Gr83_0(.din(n15510), .dout(n15513));
    jdff dff_A_t2p3AynC4_0(.din(n15513), .dout(n15516));
    jdff dff_A_fE6VYTnp9_0(.din(n15516), .dout(n15519));
    jdff dff_A_KIr9fKK00_0(.din(n15519), .dout(n15522));
    jdff dff_A_rDeUE6176_0(.din(n15522), .dout(n15525));
    jdff dff_A_HaGEhSji1_0(.din(n15525), .dout(n15528));
    jdff dff_A_Inbqn0dD7_0(.din(n15528), .dout(n15531));
    jdff dff_A_3q9vZQW89_0(.din(n15531), .dout(n15534));
    jdff dff_A_IGygduFJ1_0(.din(n15534), .dout(n15537));
    jdff dff_A_Bv5RYsxJ9_0(.din(n15537), .dout(n15540));
    jdff dff_A_zDxST4zS3_0(.din(n15540), .dout(n15543));
    jdff dff_A_bZbRI6vH5_0(.din(n15543), .dout(G440));
    jdff dff_A_lmpG2qDt1_1(.din(n5649), .dout(n15549));
    jdff dff_A_uNDxEd1U6_0(.din(n15549), .dout(n15552));
    jdff dff_A_goDTdAAp2_0(.din(n15552), .dout(n15555));
    jdff dff_A_XRqvAbIk7_0(.din(n15555), .dout(n15558));
    jdff dff_A_gsrNM9RN2_0(.din(n15558), .dout(n15561));
    jdff dff_A_guYgLIJS6_0(.din(n15561), .dout(n15564));
    jdff dff_A_9AMwW71b3_0(.din(n15564), .dout(n15567));
    jdff dff_A_ykmvIyn41_0(.din(n15567), .dout(n15570));
    jdff dff_A_xoOlKdZ24_0(.din(n15570), .dout(n15573));
    jdff dff_A_GburK90B9_0(.din(n15573), .dout(n15576));
    jdff dff_A_OeN8qLYi2_0(.din(n15576), .dout(n15579));
    jdff dff_A_EvhxFCeK1_0(.din(n15579), .dout(n15582));
    jdff dff_A_O203UWHR0_0(.din(n15582), .dout(n15585));
    jdff dff_A_FeU06reW0_0(.din(n15585), .dout(n15588));
    jdff dff_A_ZBYZw6Ck2_0(.din(n15588), .dout(n15591));
    jdff dff_A_KQ5R8WS64_0(.din(n15591), .dout(n15594));
    jdff dff_A_paOEspV96_0(.din(n15594), .dout(n15597));
    jdff dff_A_sjJDN5VP2_0(.din(n15597), .dout(n15600));
    jdff dff_A_QS5hikjm0_0(.din(n15600), .dout(n15603));
    jdff dff_A_pS4Sz9By5_0(.din(n15603), .dout(n15606));
    jdff dff_A_U3z2FtCz3_0(.din(n15606), .dout(n15609));
    jdff dff_A_FrdDRHar5_0(.din(n15609), .dout(n15612));
    jdff dff_A_r8DucLA32_0(.din(n15612), .dout(n15615));
    jdff dff_A_pX4mqxh24_0(.din(n15615), .dout(n15618));
    jdff dff_A_0BrYTy6u5_0(.din(n15618), .dout(n15621));
    jdff dff_A_6BcXm8jQ7_0(.din(n15621), .dout(G438));
    jdff dff_A_6XQh2fku4_1(.din(n5652), .dout(n15627));
    jdff dff_A_refaBZnK1_0(.din(n15627), .dout(n15630));
    jdff dff_A_v7pSivbv4_0(.din(n15630), .dout(n15633));
    jdff dff_A_5WO8c8WX3_0(.din(n15633), .dout(n15636));
    jdff dff_A_9ctrAMm45_0(.din(n15636), .dout(n15639));
    jdff dff_A_XG5Z3lUp0_0(.din(n15639), .dout(n15642));
    jdff dff_A_mIdx8PiL0_0(.din(n15642), .dout(n15645));
    jdff dff_A_s97xlK6J4_0(.din(n15645), .dout(n15648));
    jdff dff_A_MgW2xVXs6_0(.din(n15648), .dout(n15651));
    jdff dff_A_hYAfsJQT8_0(.din(n15651), .dout(n15654));
    jdff dff_A_4HD76SjN7_0(.din(n15654), .dout(n15657));
    jdff dff_A_lmRroHVc8_0(.din(n15657), .dout(n15660));
    jdff dff_A_Y5QSLk240_0(.din(n15660), .dout(n15663));
    jdff dff_A_850XsCfT5_0(.din(n15663), .dout(n15666));
    jdff dff_A_JBpYG9X07_0(.din(n15666), .dout(n15669));
    jdff dff_A_WjllqeKO9_0(.din(n15669), .dout(n15672));
    jdff dff_A_i7k7jgCg0_0(.din(n15672), .dout(n15675));
    jdff dff_A_yloCJqOE0_0(.din(n15675), .dout(n15678));
    jdff dff_A_0OnIPhgy8_0(.din(n15678), .dout(n15681));
    jdff dff_A_z8RBLO0Y4_0(.din(n15681), .dout(n15684));
    jdff dff_A_4ecQ7nfB0_0(.din(n15684), .dout(n15687));
    jdff dff_A_3C99x4QS6_0(.din(n15687), .dout(n15690));
    jdff dff_A_FP1CR0gh5_0(.din(n15690), .dout(n15693));
    jdff dff_A_xSRs55z35_0(.din(n15693), .dout(n15696));
    jdff dff_A_skyWf8pi4_0(.din(n15696), .dout(n15699));
    jdff dff_A_9kzeriYN3_0(.din(n15699), .dout(G496));
    jdff dff_A_hlgqtfXa0_1(.din(n5655), .dout(n15705));
    jdff dff_A_tbOYvf3p0_0(.din(n15705), .dout(n15708));
    jdff dff_A_hLJMW56M1_0(.din(n15708), .dout(n15711));
    jdff dff_A_dejgQg8S3_0(.din(n15711), .dout(n15714));
    jdff dff_A_ps2e0bHv0_0(.din(n15714), .dout(n15717));
    jdff dff_A_eStmDrLs9_0(.din(n15717), .dout(n15720));
    jdff dff_A_m7KfGna07_0(.din(n15720), .dout(n15723));
    jdff dff_A_3SlH0Ty24_0(.din(n15723), .dout(n15726));
    jdff dff_A_oG9KUfTy3_0(.din(n15726), .dout(n15729));
    jdff dff_A_wjNvo2rN9_0(.din(n15729), .dout(n15732));
    jdff dff_A_2TqheRFW2_0(.din(n15732), .dout(n15735));
    jdff dff_A_NoRlpiHW3_0(.din(n15735), .dout(n15738));
    jdff dff_A_YGEGc6Wu1_0(.din(n15738), .dout(n15741));
    jdff dff_A_4iv8EiES8_0(.din(n15741), .dout(n15744));
    jdff dff_A_74ndzxJd2_0(.din(n15744), .dout(n15747));
    jdff dff_A_6UgmVWUd7_0(.din(n15747), .dout(n15750));
    jdff dff_A_BrI94TK16_0(.din(n15750), .dout(n15753));
    jdff dff_A_UKYlCVZ00_0(.din(n15753), .dout(n15756));
    jdff dff_A_0CxWStX33_0(.din(n15756), .dout(n15759));
    jdff dff_A_1cE0Kbcx5_0(.din(n15759), .dout(n15762));
    jdff dff_A_Bc9wqrlK4_0(.din(n15762), .dout(n15765));
    jdff dff_A_pgItJNNg9_0(.din(n15765), .dout(n15768));
    jdff dff_A_CTE9SC373_0(.din(n15768), .dout(n15771));
    jdff dff_A_0b5GBUFN6_0(.din(n15771), .dout(n15774));
    jdff dff_A_iTnffcDf9_0(.din(n15774), .dout(n15777));
    jdff dff_A_plhMp4FJ4_0(.din(n15777), .dout(G494));
    jdff dff_A_k7VluDx66_1(.din(n5658), .dout(n15783));
    jdff dff_A_4JCyLnPT8_0(.din(n15783), .dout(n15786));
    jdff dff_A_CqQVVofU5_0(.din(n15786), .dout(n15789));
    jdff dff_A_0tGO98om5_0(.din(n15789), .dout(n15792));
    jdff dff_A_cus2wNyR3_0(.din(n15792), .dout(n15795));
    jdff dff_A_ykwg2N3S4_0(.din(n15795), .dout(n15798));
    jdff dff_A_rHEvjDg05_0(.din(n15798), .dout(n15801));
    jdff dff_A_Nr2H2tn92_0(.din(n15801), .dout(n15804));
    jdff dff_A_OWbhJzUE5_0(.din(n15804), .dout(n15807));
    jdff dff_A_SyABLrul8_0(.din(n15807), .dout(n15810));
    jdff dff_A_oAEcGWz79_0(.din(n15810), .dout(n15813));
    jdff dff_A_1JtRs0mg6_0(.din(n15813), .dout(n15816));
    jdff dff_A_QvhOosfP7_0(.din(n15816), .dout(n15819));
    jdff dff_A_cldCjiAI9_0(.din(n15819), .dout(n15822));
    jdff dff_A_2dCumnk10_0(.din(n15822), .dout(n15825));
    jdff dff_A_drQEzZcd0_0(.din(n15825), .dout(n15828));
    jdff dff_A_6m0xKfwG8_0(.din(n15828), .dout(n15831));
    jdff dff_A_EMeWYtEd7_0(.din(n15831), .dout(n15834));
    jdff dff_A_mq1eryS33_0(.din(n15834), .dout(n15837));
    jdff dff_A_vw7Fow2q3_0(.din(n15837), .dout(n15840));
    jdff dff_A_7X219nVw4_0(.din(n15840), .dout(n15843));
    jdff dff_A_zTqGXTec1_0(.din(n15843), .dout(n15846));
    jdff dff_A_SVAf83Wu1_0(.din(n15846), .dout(n15849));
    jdff dff_A_GYtMXHAg0_0(.din(n15849), .dout(n15852));
    jdff dff_A_Lg75cSrF3_0(.din(n15852), .dout(n15855));
    jdff dff_A_7Aqi7KFB9_0(.din(n15855), .dout(G492));
    jdff dff_A_f0loBwmj7_1(.din(n5661), .dout(n15861));
    jdff dff_A_UA06XAEd3_0(.din(n15861), .dout(n15864));
    jdff dff_A_KQkcnd6s5_0(.din(n15864), .dout(n15867));
    jdff dff_A_Xebfgn7k8_0(.din(n15867), .dout(n15870));
    jdff dff_A_Kb6DbJdl0_0(.din(n15870), .dout(n15873));
    jdff dff_A_oiQwF4St6_0(.din(n15873), .dout(n15876));
    jdff dff_A_7LVfNoyI8_0(.din(n15876), .dout(n15879));
    jdff dff_A_fbw2mTka4_0(.din(n15879), .dout(n15882));
    jdff dff_A_sguDky4c4_0(.din(n15882), .dout(n15885));
    jdff dff_A_6G8WXdwX6_0(.din(n15885), .dout(n15888));
    jdff dff_A_uVPYL2Fk3_0(.din(n15888), .dout(n15891));
    jdff dff_A_4VR2xzza4_0(.din(n15891), .dout(n15894));
    jdff dff_A_3c7hkXfT7_0(.din(n15894), .dout(n15897));
    jdff dff_A_PLL3p1Ae0_0(.din(n15897), .dout(n15900));
    jdff dff_A_UDPIlZY19_0(.din(n15900), .dout(n15903));
    jdff dff_A_gPGJ0XNR6_0(.din(n15903), .dout(n15906));
    jdff dff_A_VApq8idV0_0(.din(n15906), .dout(n15909));
    jdff dff_A_PCnDiEUn8_0(.din(n15909), .dout(n15912));
    jdff dff_A_QcPzhlbh9_0(.din(n15912), .dout(n15915));
    jdff dff_A_PErFiEsZ7_0(.din(n15915), .dout(n15918));
    jdff dff_A_LPQLaZXx8_0(.din(n15918), .dout(n15921));
    jdff dff_A_nU3rmj2L1_0(.din(n15921), .dout(n15924));
    jdff dff_A_K9Z7zOhI0_0(.din(n15924), .dout(n15927));
    jdff dff_A_5J3jbhlA4_0(.din(n15927), .dout(n15930));
    jdff dff_A_qfbcGDFo5_0(.din(n15930), .dout(n15933));
    jdff dff_A_W040WQg59_0(.din(n15933), .dout(G490));
    jdff dff_A_KZTb2yWC7_1(.din(n5664), .dout(n15939));
    jdff dff_A_9m7fLkwH1_0(.din(n15939), .dout(n15942));
    jdff dff_A_9o66xI0j9_0(.din(n15942), .dout(n15945));
    jdff dff_A_74RbtHo87_0(.din(n15945), .dout(n15948));
    jdff dff_A_SJrsLISZ6_0(.din(n15948), .dout(n15951));
    jdff dff_A_YDCImGTg2_0(.din(n15951), .dout(n15954));
    jdff dff_A_pKIbaLtX3_0(.din(n15954), .dout(n15957));
    jdff dff_A_8u03lCP34_0(.din(n15957), .dout(n15960));
    jdff dff_A_XAn5zpBf1_0(.din(n15960), .dout(n15963));
    jdff dff_A_ji7vzwIU7_0(.din(n15963), .dout(n15966));
    jdff dff_A_0CFrNTyK3_0(.din(n15966), .dout(n15969));
    jdff dff_A_SpUmqvJX4_0(.din(n15969), .dout(n15972));
    jdff dff_A_JFCxMApy4_0(.din(n15972), .dout(n15975));
    jdff dff_A_2o52tIzB6_0(.din(n15975), .dout(n15978));
    jdff dff_A_X0IpWm9L2_0(.din(n15978), .dout(n15981));
    jdff dff_A_67dkHOgN2_0(.din(n15981), .dout(n15984));
    jdff dff_A_gC4IHWYU7_0(.din(n15984), .dout(n15987));
    jdff dff_A_NuZIAZZe1_0(.din(n15987), .dout(n15990));
    jdff dff_A_YurapNLy8_0(.din(n15990), .dout(n15993));
    jdff dff_A_BLCgKjbE5_0(.din(n15993), .dout(n15996));
    jdff dff_A_nHtR25q09_0(.din(n15996), .dout(n15999));
    jdff dff_A_5m64xqTj3_0(.din(n15999), .dout(n16002));
    jdff dff_A_C39eLG786_0(.din(n16002), .dout(n16005));
    jdff dff_A_Z5fCVx9H0_0(.din(n16005), .dout(n16008));
    jdff dff_A_Ypbcdhpv7_0(.din(n16008), .dout(n16011));
    jdff dff_A_Qm1nj8Uz2_0(.din(n16011), .dout(G488));
    jdff dff_A_QLfkh51b8_1(.din(n5667), .dout(n16017));
    jdff dff_A_DUa9HZnC3_0(.din(n16017), .dout(n16020));
    jdff dff_A_UlCDh2JK1_0(.din(n16020), .dout(n16023));
    jdff dff_A_N2V6AKne6_0(.din(n16023), .dout(n16026));
    jdff dff_A_cG8znGBF0_0(.din(n16026), .dout(n16029));
    jdff dff_A_jU9dvUXv4_0(.din(n16029), .dout(n16032));
    jdff dff_A_6cpxOmBw2_0(.din(n16032), .dout(n16035));
    jdff dff_A_mc0wcpd06_0(.din(n16035), .dout(n16038));
    jdff dff_A_LHj9tWjm9_0(.din(n16038), .dout(n16041));
    jdff dff_A_1hts7Ibg8_0(.din(n16041), .dout(n16044));
    jdff dff_A_oB5odyPv2_0(.din(n16044), .dout(n16047));
    jdff dff_A_MKcANnJ04_0(.din(n16047), .dout(n16050));
    jdff dff_A_9CFgohJx4_0(.din(n16050), .dout(n16053));
    jdff dff_A_QwEVE3bG8_0(.din(n16053), .dout(n16056));
    jdff dff_A_vd3cvdKb9_0(.din(n16056), .dout(n16059));
    jdff dff_A_f0Zkd5IP9_0(.din(n16059), .dout(n16062));
    jdff dff_A_W3zNEd0U5_0(.din(n16062), .dout(n16065));
    jdff dff_A_z1aJ5j6L9_0(.din(n16065), .dout(n16068));
    jdff dff_A_FjTypjNG6_0(.din(n16068), .dout(n16071));
    jdff dff_A_G7vqqoYa4_0(.din(n16071), .dout(n16074));
    jdff dff_A_xw6jvl1U5_0(.din(n16074), .dout(n16077));
    jdff dff_A_SDEeN8se9_0(.din(n16077), .dout(n16080));
    jdff dff_A_bIifVykH6_0(.din(n16080), .dout(n16083));
    jdff dff_A_CtIWqBnI8_0(.din(n16083), .dout(n16086));
    jdff dff_A_5PdX3Cv19_0(.din(n16086), .dout(n16089));
    jdff dff_A_RIUIkOOA8_0(.din(n16089), .dout(G486));
    jdff dff_A_OfURwhBQ4_1(.din(n5670), .dout(n16095));
    jdff dff_A_ytSQMmZV7_0(.din(n16095), .dout(n16098));
    jdff dff_A_yINPCqiF1_0(.din(n16098), .dout(n16101));
    jdff dff_A_aX0zZrfI5_0(.din(n16101), .dout(n16104));
    jdff dff_A_Z4owilih7_0(.din(n16104), .dout(n16107));
    jdff dff_A_tA2mEIM04_0(.din(n16107), .dout(n16110));
    jdff dff_A_RNvZio891_0(.din(n16110), .dout(n16113));
    jdff dff_A_7PgBZI536_0(.din(n16113), .dout(n16116));
    jdff dff_A_ZMV5J3RQ6_0(.din(n16116), .dout(n16119));
    jdff dff_A_zDAudBa62_0(.din(n16119), .dout(n16122));
    jdff dff_A_drX3DFpO8_0(.din(n16122), .dout(n16125));
    jdff dff_A_iwCJhtCM6_0(.din(n16125), .dout(n16128));
    jdff dff_A_VnZKnpWY9_0(.din(n16128), .dout(n16131));
    jdff dff_A_uRyf39Wa0_0(.din(n16131), .dout(n16134));
    jdff dff_A_XCCaCKBf8_0(.din(n16134), .dout(n16137));
    jdff dff_A_0RZ9zW1X4_0(.din(n16137), .dout(n16140));
    jdff dff_A_WfZcjshR7_0(.din(n16140), .dout(n16143));
    jdff dff_A_B88VNbXs3_0(.din(n16143), .dout(n16146));
    jdff dff_A_YkKK2TBb4_0(.din(n16146), .dout(n16149));
    jdff dff_A_3JpGJlkj6_0(.din(n16149), .dout(n16152));
    jdff dff_A_aRnGBIFF9_0(.din(n16152), .dout(n16155));
    jdff dff_A_9LIutuJ13_0(.din(n16155), .dout(n16158));
    jdff dff_A_AagqdROk1_0(.din(n16158), .dout(n16161));
    jdff dff_A_QmDodXM35_0(.din(n16161), .dout(n16164));
    jdff dff_A_9HjBWwfe6_0(.din(n16164), .dout(n16167));
    jdff dff_A_980EDFiP5_0(.din(n16167), .dout(G484));
    jdff dff_A_fIekaECE3_1(.din(n5673), .dout(n16173));
    jdff dff_A_bk775PTy5_0(.din(n16173), .dout(n16176));
    jdff dff_A_IIfDcN731_0(.din(n16176), .dout(n16179));
    jdff dff_A_5PMu0ONu2_0(.din(n16179), .dout(n16182));
    jdff dff_A_eLol9rpd9_0(.din(n16182), .dout(n16185));
    jdff dff_A_PLHaiAic9_0(.din(n16185), .dout(n16188));
    jdff dff_A_mZTV7jyz6_0(.din(n16188), .dout(n16191));
    jdff dff_A_lcJl65Ah2_0(.din(n16191), .dout(n16194));
    jdff dff_A_6QXCIqm39_0(.din(n16194), .dout(n16197));
    jdff dff_A_dSNySXUc9_0(.din(n16197), .dout(n16200));
    jdff dff_A_7l5v8nxi4_0(.din(n16200), .dout(n16203));
    jdff dff_A_rNrrtCYT4_0(.din(n16203), .dout(n16206));
    jdff dff_A_CHI7qLaG5_0(.din(n16206), .dout(n16209));
    jdff dff_A_sELod8Nb5_0(.din(n16209), .dout(n16212));
    jdff dff_A_xf27V03z0_0(.din(n16212), .dout(n16215));
    jdff dff_A_7tmE429A8_0(.din(n16215), .dout(n16218));
    jdff dff_A_MESAuxb88_0(.din(n16218), .dout(n16221));
    jdff dff_A_vwHscXbt7_0(.din(n16221), .dout(n16224));
    jdff dff_A_PLGKFfh65_0(.din(n16224), .dout(n16227));
    jdff dff_A_d75bt1mm2_0(.din(n16227), .dout(n16230));
    jdff dff_A_etmB4GOC4_0(.din(n16230), .dout(n16233));
    jdff dff_A_sBArkJi94_0(.din(n16233), .dout(n16236));
    jdff dff_A_Z8MyH8wl9_0(.din(n16236), .dout(n16239));
    jdff dff_A_Z2kC9TQE6_0(.din(n16239), .dout(n16242));
    jdff dff_A_nLGhbYri1_0(.din(n16242), .dout(n16245));
    jdff dff_A_CCE3pTEC0_0(.din(n16245), .dout(G482));
    jdff dff_A_gOv57F6o7_1(.din(n5676), .dout(n16251));
    jdff dff_A_4ycNk5ue3_0(.din(n16251), .dout(n16254));
    jdff dff_A_kQb6alwb4_0(.din(n16254), .dout(n16257));
    jdff dff_A_750YHGfC0_0(.din(n16257), .dout(n16260));
    jdff dff_A_1jsP5YW74_0(.din(n16260), .dout(n16263));
    jdff dff_A_rQRGYg105_0(.din(n16263), .dout(n16266));
    jdff dff_A_pGGC2MO08_0(.din(n16266), .dout(n16269));
    jdff dff_A_hz0j8EbO0_0(.din(n16269), .dout(n16272));
    jdff dff_A_wvPlMp6f5_0(.din(n16272), .dout(n16275));
    jdff dff_A_te0lC6vD2_0(.din(n16275), .dout(n16278));
    jdff dff_A_lTnOwFar8_0(.din(n16278), .dout(n16281));
    jdff dff_A_axSqLTYo9_0(.din(n16281), .dout(n16284));
    jdff dff_A_vVKtUhnG0_0(.din(n16284), .dout(n16287));
    jdff dff_A_gKwZEhym9_0(.din(n16287), .dout(n16290));
    jdff dff_A_SQYHVqPZ2_0(.din(n16290), .dout(n16293));
    jdff dff_A_GszOT3Ft5_0(.din(n16293), .dout(n16296));
    jdff dff_A_1KIl7Y784_0(.din(n16296), .dout(n16299));
    jdff dff_A_HGmNnvMP1_0(.din(n16299), .dout(n16302));
    jdff dff_A_fjvhIx1R6_0(.din(n16302), .dout(n16305));
    jdff dff_A_VKCNYq9P8_0(.din(n16305), .dout(n16308));
    jdff dff_A_lM8MGmMt3_0(.din(n16308), .dout(n16311));
    jdff dff_A_N8yYnooQ6_0(.din(n16311), .dout(n16314));
    jdff dff_A_NSmpGyrU1_0(.din(n16314), .dout(n16317));
    jdff dff_A_PWWzkdMT3_0(.din(n16317), .dout(n16320));
    jdff dff_A_AcKnVu8F1_0(.din(n16320), .dout(n16323));
    jdff dff_A_1IMPCMjz6_0(.din(n16323), .dout(G480));
    jdff dff_A_11QQyRH85_1(.din(n5679), .dout(n16329));
    jdff dff_A_UjXJohJy7_0(.din(n16329), .dout(n16332));
    jdff dff_A_ShEUuRJO0_0(.din(n16332), .dout(n16335));
    jdff dff_A_tg3mlVew4_0(.din(n16335), .dout(n16338));
    jdff dff_A_4J1i6TzQ3_0(.din(n16338), .dout(n16341));
    jdff dff_A_7ZwDlCyW6_0(.din(n16341), .dout(n16344));
    jdff dff_A_VXPcrupP7_0(.din(n16344), .dout(n16347));
    jdff dff_A_Itga5flg1_0(.din(n16347), .dout(n16350));
    jdff dff_A_VwnCLoSN9_0(.din(n16350), .dout(n16353));
    jdff dff_A_91dpDgg91_0(.din(n16353), .dout(n16356));
    jdff dff_A_UpWY8KVq9_0(.din(n16356), .dout(n16359));
    jdff dff_A_bAoMvQUp4_0(.din(n16359), .dout(n16362));
    jdff dff_A_UgK6i5xj8_0(.din(n16362), .dout(n16365));
    jdff dff_A_3H0IbKDz8_0(.din(n16365), .dout(n16368));
    jdff dff_A_wbSVtmAL5_0(.din(n16368), .dout(n16371));
    jdff dff_A_83nN3jnE0_0(.din(n16371), .dout(n16374));
    jdff dff_A_52jTadLY9_0(.din(n16374), .dout(n16377));
    jdff dff_A_Bt01Oqwz6_0(.din(n16377), .dout(n16380));
    jdff dff_A_BAh45ch20_0(.din(n16380), .dout(n16383));
    jdff dff_A_lVSsa0Tp3_0(.din(n16383), .dout(n16386));
    jdff dff_A_WlWbRkXP1_0(.din(n16386), .dout(n16389));
    jdff dff_A_P2OROSa06_0(.din(n16389), .dout(n16392));
    jdff dff_A_SxaMNOeq4_0(.din(n16392), .dout(n16395));
    jdff dff_A_yA0kOM8s5_0(.din(n16395), .dout(n16398));
    jdff dff_A_2QpzgJ2M6_0(.din(n16398), .dout(n16401));
    jdff dff_A_Cnhvxw4A4_0(.din(n16401), .dout(G560));
    jdff dff_A_9okMP1UV2_1(.din(n5682), .dout(n16407));
    jdff dff_A_W0z5pZCe5_0(.din(n16407), .dout(n16410));
    jdff dff_A_tqrobSO45_0(.din(n16410), .dout(n16413));
    jdff dff_A_olNmtkdm8_0(.din(n16413), .dout(n16416));
    jdff dff_A_vckhYKQb4_0(.din(n16416), .dout(n16419));
    jdff dff_A_kBPXqeMc7_0(.din(n16419), .dout(n16422));
    jdff dff_A_g3WJ2c3N6_0(.din(n16422), .dout(n16425));
    jdff dff_A_wM3Xz4T23_0(.din(n16425), .dout(n16428));
    jdff dff_A_CCiZ0XNY6_0(.din(n16428), .dout(n16431));
    jdff dff_A_xLCoukH15_0(.din(n16431), .dout(n16434));
    jdff dff_A_XGY4ms5n3_0(.din(n16434), .dout(n16437));
    jdff dff_A_G41BNQGi2_0(.din(n16437), .dout(n16440));
    jdff dff_A_FL7zkHKh0_0(.din(n16440), .dout(n16443));
    jdff dff_A_3HXQdHjF9_0(.din(n16443), .dout(n16446));
    jdff dff_A_5gDjCqpK0_0(.din(n16446), .dout(n16449));
    jdff dff_A_nOXzo6UW1_0(.din(n16449), .dout(n16452));
    jdff dff_A_9zHsPENT5_0(.din(n16452), .dout(n16455));
    jdff dff_A_SSqTzJ4a8_0(.din(n16455), .dout(n16458));
    jdff dff_A_WC0oSFax0_0(.din(n16458), .dout(n16461));
    jdff dff_A_Nw7VJFwA3_0(.din(n16461), .dout(n16464));
    jdff dff_A_a2kMC4mj5_0(.din(n16464), .dout(n16467));
    jdff dff_A_FMGgHupn6_0(.din(n16467), .dout(n16470));
    jdff dff_A_F6impo4g7_0(.din(n16470), .dout(n16473));
    jdff dff_A_T8b8AyAx1_0(.din(n16473), .dout(n16476));
    jdff dff_A_B7P0jwiJ3_0(.din(n16476), .dout(n16479));
    jdff dff_A_QByHr7ms8_0(.din(n16479), .dout(G542));
    jdff dff_A_XMLPmksm8_1(.din(n5685), .dout(n16485));
    jdff dff_A_nXCBi7Zg4_0(.din(n16485), .dout(n16488));
    jdff dff_A_vata1kJy9_0(.din(n16488), .dout(n16491));
    jdff dff_A_X5xU5kKc2_0(.din(n16491), .dout(n16494));
    jdff dff_A_OcHyEATI4_0(.din(n16494), .dout(n16497));
    jdff dff_A_xtrwPTaF7_0(.din(n16497), .dout(n16500));
    jdff dff_A_TuikUtQJ5_0(.din(n16500), .dout(n16503));
    jdff dff_A_ScJYNUfR6_0(.din(n16503), .dout(n16506));
    jdff dff_A_EFkx2fPr0_0(.din(n16506), .dout(n16509));
    jdff dff_A_05fRovvS0_0(.din(n16509), .dout(n16512));
    jdff dff_A_gOoMGAOP1_0(.din(n16512), .dout(n16515));
    jdff dff_A_6CdV0Dx76_0(.din(n16515), .dout(n16518));
    jdff dff_A_vhsbPAM43_0(.din(n16518), .dout(n16521));
    jdff dff_A_U2PW0Nf06_0(.din(n16521), .dout(n16524));
    jdff dff_A_x6PQxXnG6_0(.din(n16524), .dout(n16527));
    jdff dff_A_g1Ki7iYn5_0(.din(n16527), .dout(n16530));
    jdff dff_A_LSN81seR6_0(.din(n16530), .dout(n16533));
    jdff dff_A_umLDc4e32_0(.din(n16533), .dout(n16536));
    jdff dff_A_D3Z8w65C0_0(.din(n16536), .dout(n16539));
    jdff dff_A_kZ0VP6MF3_0(.din(n16539), .dout(n16542));
    jdff dff_A_9MQfuMzn7_0(.din(n16542), .dout(n16545));
    jdff dff_A_Q4hBb8IV3_0(.din(n16545), .dout(n16548));
    jdff dff_A_zSXUF6JB8_0(.din(n16548), .dout(n16551));
    jdff dff_A_FxPuHxzq9_0(.din(n16551), .dout(n16554));
    jdff dff_A_fIEu4iUG2_0(.din(n16554), .dout(n16557));
    jdff dff_A_aSYzNRAE5_0(.din(n16557), .dout(G558));
    jdff dff_A_RwGKFHG76_1(.din(n5688), .dout(n16563));
    jdff dff_A_pSsJqAGi2_0(.din(n16563), .dout(n16566));
    jdff dff_A_QTQ3LRou3_0(.din(n16566), .dout(n16569));
    jdff dff_A_zHpTy2Ma4_0(.din(n16569), .dout(n16572));
    jdff dff_A_6U9Q47tX8_0(.din(n16572), .dout(n16575));
    jdff dff_A_vQSlVRYl5_0(.din(n16575), .dout(n16578));
    jdff dff_A_lqbPE6rA9_0(.din(n16578), .dout(n16581));
    jdff dff_A_DhQ8CBJN5_0(.din(n16581), .dout(n16584));
    jdff dff_A_0mmd6iAP6_0(.din(n16584), .dout(n16587));
    jdff dff_A_B4B3iqNi7_0(.din(n16587), .dout(n16590));
    jdff dff_A_6V3SgN718_0(.din(n16590), .dout(n16593));
    jdff dff_A_xPzwMw5Y4_0(.din(n16593), .dout(n16596));
    jdff dff_A_pFhm7M850_0(.din(n16596), .dout(n16599));
    jdff dff_A_DHgizohK1_0(.din(n16599), .dout(n16602));
    jdff dff_A_QoKQdfTy8_0(.din(n16602), .dout(n16605));
    jdff dff_A_xdsvHBIa9_0(.din(n16605), .dout(n16608));
    jdff dff_A_FqKVM69n1_0(.din(n16608), .dout(n16611));
    jdff dff_A_z73PWgP01_0(.din(n16611), .dout(n16614));
    jdff dff_A_KZNvMPRo8_0(.din(n16614), .dout(n16617));
    jdff dff_A_DDY7NAzT2_0(.din(n16617), .dout(n16620));
    jdff dff_A_WmMGUKcV8_0(.din(n16620), .dout(n16623));
    jdff dff_A_Eu8t7ZoD2_0(.din(n16623), .dout(n16626));
    jdff dff_A_Ui7AEILB9_0(.din(n16626), .dout(n16629));
    jdff dff_A_MXzLsN6d8_0(.din(n16629), .dout(n16632));
    jdff dff_A_uaTHpDKo8_0(.din(n16632), .dout(n16635));
    jdff dff_A_yI6apG2r3_0(.din(n16635), .dout(G556));
    jdff dff_A_o7j95bj09_1(.din(n5691), .dout(n16641));
    jdff dff_A_RCk2tpz64_0(.din(n16641), .dout(n16644));
    jdff dff_A_9iGhDWcK7_0(.din(n16644), .dout(n16647));
    jdff dff_A_dsHEauon1_0(.din(n16647), .dout(n16650));
    jdff dff_A_8AZu8qJD2_0(.din(n16650), .dout(n16653));
    jdff dff_A_7uOv7Jir4_0(.din(n16653), .dout(n16656));
    jdff dff_A_0Cliso2d7_0(.din(n16656), .dout(n16659));
    jdff dff_A_1qFCwSei7_0(.din(n16659), .dout(n16662));
    jdff dff_A_G4vSpu0G5_0(.din(n16662), .dout(n16665));
    jdff dff_A_wE2z1JIn6_0(.din(n16665), .dout(n16668));
    jdff dff_A_bcaSGDxa1_0(.din(n16668), .dout(n16671));
    jdff dff_A_JKQi14PJ0_0(.din(n16671), .dout(n16674));
    jdff dff_A_C0DiUZfg5_0(.din(n16674), .dout(n16677));
    jdff dff_A_XkoFf4qk1_0(.din(n16677), .dout(n16680));
    jdff dff_A_Sb6cXqc88_0(.din(n16680), .dout(n16683));
    jdff dff_A_HXKwbOBe7_0(.din(n16683), .dout(n16686));
    jdff dff_A_SsSbmzrP0_0(.din(n16686), .dout(n16689));
    jdff dff_A_fT3hszoY9_0(.din(n16689), .dout(n16692));
    jdff dff_A_4jYnIGsu8_0(.din(n16692), .dout(n16695));
    jdff dff_A_mSQhwvnh6_0(.din(n16695), .dout(n16698));
    jdff dff_A_R2BG7Hr51_0(.din(n16698), .dout(n16701));
    jdff dff_A_qiy3e5fv6_0(.din(n16701), .dout(n16704));
    jdff dff_A_v4Qi1qBk1_0(.din(n16704), .dout(n16707));
    jdff dff_A_DZwuPhxq7_0(.din(n16707), .dout(n16710));
    jdff dff_A_gcSvZpbq3_0(.din(n16710), .dout(n16713));
    jdff dff_A_h2PKgTfh5_0(.din(n16713), .dout(G554));
    jdff dff_A_SwcSZ5mu2_1(.din(n5694), .dout(n16719));
    jdff dff_A_I5TtFsPO3_0(.din(n16719), .dout(n16722));
    jdff dff_A_I7sBW1ym7_0(.din(n16722), .dout(n16725));
    jdff dff_A_8nuYlqo78_0(.din(n16725), .dout(n16728));
    jdff dff_A_H1pT0KGG1_0(.din(n16728), .dout(n16731));
    jdff dff_A_mTgeVoxi5_0(.din(n16731), .dout(n16734));
    jdff dff_A_r4j6ACKh3_0(.din(n16734), .dout(n16737));
    jdff dff_A_OpoqpKPM1_0(.din(n16737), .dout(n16740));
    jdff dff_A_JlLzhrCR7_0(.din(n16740), .dout(n16743));
    jdff dff_A_1NKXrdeO7_0(.din(n16743), .dout(n16746));
    jdff dff_A_FY8pf0bB7_0(.din(n16746), .dout(n16749));
    jdff dff_A_qNhI5oZQ8_0(.din(n16749), .dout(n16752));
    jdff dff_A_ex65tSP45_0(.din(n16752), .dout(n16755));
    jdff dff_A_LzjMLhai6_0(.din(n16755), .dout(n16758));
    jdff dff_A_0s70ksDY3_0(.din(n16758), .dout(n16761));
    jdff dff_A_eahvI2Tw5_0(.din(n16761), .dout(n16764));
    jdff dff_A_O5ChEaQ90_0(.din(n16764), .dout(n16767));
    jdff dff_A_xUzzNqTC1_0(.din(n16767), .dout(n16770));
    jdff dff_A_JTDcJUGE2_0(.din(n16770), .dout(n16773));
    jdff dff_A_OrQMIMW96_0(.din(n16773), .dout(n16776));
    jdff dff_A_Z0MWjToV7_0(.din(n16776), .dout(n16779));
    jdff dff_A_asxkmu0C6_0(.din(n16779), .dout(n16782));
    jdff dff_A_CnTbIlim7_0(.din(n16782), .dout(n16785));
    jdff dff_A_5eOxR1ck5_0(.din(n16785), .dout(n16788));
    jdff dff_A_YRco1Ivp7_0(.din(n16788), .dout(n16791));
    jdff dff_A_WqGolFye2_0(.din(n16791), .dout(G552));
    jdff dff_A_UOFpF7hR0_1(.din(n5697), .dout(n16797));
    jdff dff_A_DFmfw6vG3_0(.din(n16797), .dout(n16800));
    jdff dff_A_ne2TrUOm7_0(.din(n16800), .dout(n16803));
    jdff dff_A_HixFBzjI3_0(.din(n16803), .dout(n16806));
    jdff dff_A_NtJ9bVEG1_0(.din(n16806), .dout(n16809));
    jdff dff_A_QP80W6xl8_0(.din(n16809), .dout(n16812));
    jdff dff_A_sufIrqeR3_0(.din(n16812), .dout(n16815));
    jdff dff_A_QHxrtEBw3_0(.din(n16815), .dout(n16818));
    jdff dff_A_RmGhJCkc5_0(.din(n16818), .dout(n16821));
    jdff dff_A_gjMK7HsI2_0(.din(n16821), .dout(n16824));
    jdff dff_A_63XSR0MP2_0(.din(n16824), .dout(n16827));
    jdff dff_A_ldZWNcFg1_0(.din(n16827), .dout(n16830));
    jdff dff_A_sgeEwrXI0_0(.din(n16830), .dout(n16833));
    jdff dff_A_T1s58ywb7_0(.din(n16833), .dout(n16836));
    jdff dff_A_cS2UAUHB4_0(.din(n16836), .dout(n16839));
    jdff dff_A_hHRRzcPO5_0(.din(n16839), .dout(n16842));
    jdff dff_A_GMB2abC96_0(.din(n16842), .dout(n16845));
    jdff dff_A_SUMRqDyo5_0(.din(n16845), .dout(n16848));
    jdff dff_A_bdWj76Op9_0(.din(n16848), .dout(n16851));
    jdff dff_A_DqUTDiHQ6_0(.din(n16851), .dout(n16854));
    jdff dff_A_2reMXbBq1_0(.din(n16854), .dout(n16857));
    jdff dff_A_h7KHJgaO4_0(.din(n16857), .dout(n16860));
    jdff dff_A_dwLIIFPH4_0(.din(n16860), .dout(n16863));
    jdff dff_A_1Wbd86ql5_0(.din(n16863), .dout(n16866));
    jdff dff_A_E6XSqH0Y5_0(.din(n16866), .dout(n16869));
    jdff dff_A_XzveyaxA5_0(.din(n16869), .dout(G550));
    jdff dff_A_3rAom8zd6_1(.din(n5700), .dout(n16875));
    jdff dff_A_fYXRzNNc1_0(.din(n16875), .dout(n16878));
    jdff dff_A_Mtc00sxC0_0(.din(n16878), .dout(n16881));
    jdff dff_A_t5bc0efI2_0(.din(n16881), .dout(n16884));
    jdff dff_A_C3oAI2Fi4_0(.din(n16884), .dout(n16887));
    jdff dff_A_FH2lil4W1_0(.din(n16887), .dout(n16890));
    jdff dff_A_QqZeptEe5_0(.din(n16890), .dout(n16893));
    jdff dff_A_BvkR98yw1_0(.din(n16893), .dout(n16896));
    jdff dff_A_wBytA4eS0_0(.din(n16896), .dout(n16899));
    jdff dff_A_W1Nj9btQ3_0(.din(n16899), .dout(n16902));
    jdff dff_A_WIoNprCO3_0(.din(n16902), .dout(n16905));
    jdff dff_A_oTH6z8ii4_0(.din(n16905), .dout(n16908));
    jdff dff_A_iNIdyMhq9_0(.din(n16908), .dout(n16911));
    jdff dff_A_wr3GPQIf2_0(.din(n16911), .dout(n16914));
    jdff dff_A_RN5oxCKr4_0(.din(n16914), .dout(n16917));
    jdff dff_A_GBLQJdzc8_0(.din(n16917), .dout(n16920));
    jdff dff_A_6GrH231a8_0(.din(n16920), .dout(n16923));
    jdff dff_A_LzCj4MQa3_0(.din(n16923), .dout(n16926));
    jdff dff_A_YNuIQ53q7_0(.din(n16926), .dout(n16929));
    jdff dff_A_Qv19K5je0_0(.din(n16929), .dout(n16932));
    jdff dff_A_uVgXRt9m1_0(.din(n16932), .dout(n16935));
    jdff dff_A_0fqMLhtF9_0(.din(n16935), .dout(n16938));
    jdff dff_A_IxknPB2B0_0(.din(n16938), .dout(n16941));
    jdff dff_A_lDRYKVjv0_0(.din(n16941), .dout(n16944));
    jdff dff_A_rfayoZ0G4_0(.din(n16944), .dout(n16947));
    jdff dff_A_HGvALjB69_0(.din(n16947), .dout(G548));
    jdff dff_A_jC7At71Q2_1(.din(n5703), .dout(n16953));
    jdff dff_A_LxBBIU8o3_0(.din(n16953), .dout(n16956));
    jdff dff_A_r9UDQrDN1_0(.din(n16956), .dout(n16959));
    jdff dff_A_FkUvftfL8_0(.din(n16959), .dout(n16962));
    jdff dff_A_tDVD6uAd0_0(.din(n16962), .dout(n16965));
    jdff dff_A_ujznNtWB1_0(.din(n16965), .dout(n16968));
    jdff dff_A_9u2bSJuP0_0(.din(n16968), .dout(n16971));
    jdff dff_A_6A8laloR9_0(.din(n16971), .dout(n16974));
    jdff dff_A_4bnnsnk34_0(.din(n16974), .dout(n16977));
    jdff dff_A_hCILH0XJ5_0(.din(n16977), .dout(n16980));
    jdff dff_A_8E1PgMP80_0(.din(n16980), .dout(n16983));
    jdff dff_A_cOc4c2bI7_0(.din(n16983), .dout(n16986));
    jdff dff_A_it3y7hed1_0(.din(n16986), .dout(n16989));
    jdff dff_A_GhWC7yu38_0(.din(n16989), .dout(n16992));
    jdff dff_A_H5skBDB29_0(.din(n16992), .dout(n16995));
    jdff dff_A_6obFelOy3_0(.din(n16995), .dout(n16998));
    jdff dff_A_cJ7KDIQ20_0(.din(n16998), .dout(n17001));
    jdff dff_A_9qrHKiPs2_0(.din(n17001), .dout(n17004));
    jdff dff_A_yclbE7nM1_0(.din(n17004), .dout(n17007));
    jdff dff_A_WHkxj6nR7_0(.din(n17007), .dout(n17010));
    jdff dff_A_ADqu8nAL5_0(.din(n17010), .dout(n17013));
    jdff dff_A_wvVlABbh6_0(.din(n17013), .dout(n17016));
    jdff dff_A_V6m99F9k9_0(.din(n17016), .dout(n17019));
    jdff dff_A_iGzYGW3S4_0(.din(n17019), .dout(n17022));
    jdff dff_A_L4fSNyRt2_0(.din(n17022), .dout(n17025));
    jdff dff_A_Cu3qY5nH9_0(.din(n17025), .dout(G546));
    jdff dff_A_O7RMNuf06_1(.din(n5706), .dout(n17031));
    jdff dff_A_doiTLMWg7_0(.din(n17031), .dout(n17034));
    jdff dff_A_pg5VpNzU3_0(.din(n17034), .dout(n17037));
    jdff dff_A_uWjlNu2E3_0(.din(n17037), .dout(n17040));
    jdff dff_A_ljXNqORV6_0(.din(n17040), .dout(n17043));
    jdff dff_A_WqFnMp7F1_0(.din(n17043), .dout(n17046));
    jdff dff_A_yIgB1hws4_0(.din(n17046), .dout(n17049));
    jdff dff_A_3Mn7T0Mc1_0(.din(n17049), .dout(n17052));
    jdff dff_A_vKDjREg19_0(.din(n17052), .dout(n17055));
    jdff dff_A_y6BvsBzb5_0(.din(n17055), .dout(n17058));
    jdff dff_A_JefxyndS9_0(.din(n17058), .dout(n17061));
    jdff dff_A_OWHgQ3gL0_0(.din(n17061), .dout(n17064));
    jdff dff_A_w8U8XJOq5_0(.din(n17064), .dout(n17067));
    jdff dff_A_QbVkguio0_0(.din(n17067), .dout(n17070));
    jdff dff_A_NT8Dk4SR2_0(.din(n17070), .dout(n17073));
    jdff dff_A_aRnnqE9j7_0(.din(n17073), .dout(n17076));
    jdff dff_A_jkl0cphT9_0(.din(n17076), .dout(n17079));
    jdff dff_A_MIVY0kBj5_0(.din(n17079), .dout(n17082));
    jdff dff_A_I2AoVKde4_0(.din(n17082), .dout(n17085));
    jdff dff_A_4pytqjya8_0(.din(n17085), .dout(n17088));
    jdff dff_A_EP2uysYu8_0(.din(n17088), .dout(n17091));
    jdff dff_A_OylISZWJ4_0(.din(n17091), .dout(n17094));
    jdff dff_A_U3RlEzgC0_0(.din(n17094), .dout(n17097));
    jdff dff_A_SkPYBmGP8_0(.din(n17097), .dout(n17100));
    jdff dff_A_fDWQvJ6h5_0(.din(n17100), .dout(n17103));
    jdff dff_A_6MiqYO5M0_0(.din(n17103), .dout(G544));
    jdff dff_A_cykvuITa8_1(.din(n5709), .dout(n17109));
    jdff dff_A_770ukYv22_0(.din(n17109), .dout(n17112));
    jdff dff_A_aJRWQdhK0_0(.din(n17112), .dout(n17115));
    jdff dff_A_lKFzJtcr0_0(.din(n17115), .dout(n17118));
    jdff dff_A_q9bJKAqu5_0(.din(n17118), .dout(n17121));
    jdff dff_A_zVZkXWJq6_0(.din(n17121), .dout(n17124));
    jdff dff_A_xo0s4Jdx9_0(.din(n17124), .dout(n17127));
    jdff dff_A_qYZ9UaqO6_0(.din(n17127), .dout(n17130));
    jdff dff_A_zeNUlbEx4_0(.din(n17130), .dout(n17133));
    jdff dff_A_WqjG7eI77_0(.din(n17133), .dout(n17136));
    jdff dff_A_1Zn3Ue1k8_0(.din(n17136), .dout(n17139));
    jdff dff_A_u1bfDX7C2_0(.din(n17139), .dout(n17142));
    jdff dff_A_E1CkVYeH5_0(.din(n17142), .dout(n17145));
    jdff dff_A_TymXuwcy5_0(.din(n17145), .dout(n17148));
    jdff dff_A_wG4UJRUV2_0(.din(n17148), .dout(n17151));
    jdff dff_A_DMadvdJh4_0(.din(n17151), .dout(n17154));
    jdff dff_A_bM89scTp8_0(.din(n17154), .dout(n17157));
    jdff dff_A_jUY7NL5b5_0(.din(n17157), .dout(n17160));
    jdff dff_A_aMmGBlsD6_0(.din(n17160), .dout(n17163));
    jdff dff_A_s7grm0hQ4_0(.din(n17163), .dout(n17166));
    jdff dff_A_56FFMSOa8_0(.din(n17166), .dout(n17169));
    jdff dff_A_VhFAjZOL5_0(.din(n17169), .dout(n17172));
    jdff dff_A_rSbD6nUO1_0(.din(n17172), .dout(n17175));
    jdff dff_A_4S3Q3aPN4_0(.din(n17175), .dout(n17178));
    jdff dff_A_f2bmOJli8_0(.din(n17178), .dout(n17181));
    jdff dff_A_Ub6SdZnE2_0(.din(n17181), .dout(G540));
    jdff dff_A_ZmdyHmdd8_1(.din(n5712), .dout(n17187));
    jdff dff_A_mcWpOpJu8_0(.din(n17187), .dout(n17190));
    jdff dff_A_JAMipuF20_0(.din(n17190), .dout(n17193));
    jdff dff_A_lcdRUCoI8_0(.din(n17193), .dout(n17196));
    jdff dff_A_l0sFi7ci9_0(.din(n17196), .dout(n17199));
    jdff dff_A_14pZ2zFV1_0(.din(n17199), .dout(n17202));
    jdff dff_A_kM4IefWL3_0(.din(n17202), .dout(n17205));
    jdff dff_A_3SC9EuCc1_0(.din(n17205), .dout(n17208));
    jdff dff_A_p9rERASQ0_0(.din(n17208), .dout(n17211));
    jdff dff_A_w18NPP820_0(.din(n17211), .dout(n17214));
    jdff dff_A_xQNOfzUB7_0(.din(n17214), .dout(n17217));
    jdff dff_A_z1NqDnVO2_0(.din(n17217), .dout(n17220));
    jdff dff_A_Pznzn9Fh9_0(.din(n17220), .dout(n17223));
    jdff dff_A_RnIBIxir5_0(.din(n17223), .dout(n17226));
    jdff dff_A_bilz34lm8_0(.din(n17226), .dout(n17229));
    jdff dff_A_AefvOYKG9_0(.din(n17229), .dout(n17232));
    jdff dff_A_DhX6PBLq1_0(.din(n17232), .dout(n17235));
    jdff dff_A_7kpp6Y2X0_0(.din(n17235), .dout(n17238));
    jdff dff_A_il0yoA8c2_0(.din(n17238), .dout(n17241));
    jdff dff_A_VNUV6xRn4_0(.din(n17241), .dout(n17244));
    jdff dff_A_UsKiHWMT2_0(.din(n17244), .dout(n17247));
    jdff dff_A_RhI2wq0z5_0(.din(n17247), .dout(n17250));
    jdff dff_A_NTf5VPGD7_0(.din(n17250), .dout(n17253));
    jdff dff_A_bTcdFqlR5_0(.din(n17253), .dout(n17256));
    jdff dff_A_1E3cOk3U5_0(.din(n17256), .dout(n17259));
    jdff dff_A_6latRHez4_0(.din(n17259), .dout(G538));
    jdff dff_A_bVT2Wp258_1(.din(n5715), .dout(n17265));
    jdff dff_A_TWjxMiy76_0(.din(n17265), .dout(n17268));
    jdff dff_A_ZEcQB5Jl7_0(.din(n17268), .dout(n17271));
    jdff dff_A_DNfbcwZX4_0(.din(n17271), .dout(n17274));
    jdff dff_A_rt1KetpS8_0(.din(n17274), .dout(n17277));
    jdff dff_A_d83EbDdg2_0(.din(n17277), .dout(n17280));
    jdff dff_A_3bZAt0Hm5_0(.din(n17280), .dout(n17283));
    jdff dff_A_gBrCuvdu4_0(.din(n17283), .dout(n17286));
    jdff dff_A_W5yMHXz95_0(.din(n17286), .dout(n17289));
    jdff dff_A_ZZ9zmRnp3_0(.din(n17289), .dout(n17292));
    jdff dff_A_31WN9WR89_0(.din(n17292), .dout(n17295));
    jdff dff_A_dGioZHas1_0(.din(n17295), .dout(n17298));
    jdff dff_A_NP4F7CHk5_0(.din(n17298), .dout(n17301));
    jdff dff_A_txfAdmnr5_0(.din(n17301), .dout(n17304));
    jdff dff_A_dE6GOoFS8_0(.din(n17304), .dout(n17307));
    jdff dff_A_bL9jkJr21_0(.din(n17307), .dout(n17310));
    jdff dff_A_PCsnKyw47_0(.din(n17310), .dout(n17313));
    jdff dff_A_WKZ7MFIb3_0(.din(n17313), .dout(n17316));
    jdff dff_A_dehq0JxD4_0(.din(n17316), .dout(n17319));
    jdff dff_A_PRdaNg3o0_0(.din(n17319), .dout(n17322));
    jdff dff_A_73lR5fPK3_0(.din(n17322), .dout(n17325));
    jdff dff_A_BwZ9htRo1_0(.din(n17325), .dout(n17328));
    jdff dff_A_VUwT3GaX3_0(.din(n17328), .dout(n17331));
    jdff dff_A_apxQIS8p5_0(.din(n17331), .dout(n17334));
    jdff dff_A_CK0UtfAN4_0(.din(n17334), .dout(n17337));
    jdff dff_A_9vdyOd9n5_0(.din(n17337), .dout(G536));
    jdff dff_A_1ISwIh973_1(.din(n5718), .dout(n17343));
    jdff dff_A_xxcJnGPc1_0(.din(n17343), .dout(n17346));
    jdff dff_A_1f89aRfw3_0(.din(n17346), .dout(n17349));
    jdff dff_A_zaiDhMWa6_0(.din(n17349), .dout(n17352));
    jdff dff_A_xlZk6Hun3_0(.din(n17352), .dout(n17355));
    jdff dff_A_IiRPdPLX1_0(.din(n17355), .dout(n17358));
    jdff dff_A_AmsLyTTL7_0(.din(n17358), .dout(n17361));
    jdff dff_A_UYH5WbYg5_0(.din(n17361), .dout(n17364));
    jdff dff_A_xzCKYHee1_0(.din(n17364), .dout(n17367));
    jdff dff_A_F0ydn2vw7_0(.din(n17367), .dout(n17370));
    jdff dff_A_lf1zOueQ8_0(.din(n17370), .dout(n17373));
    jdff dff_A_mrDtIXis0_0(.din(n17373), .dout(n17376));
    jdff dff_A_CiyHWuyA4_0(.din(n17376), .dout(n17379));
    jdff dff_A_5yH4yel01_0(.din(n17379), .dout(n17382));
    jdff dff_A_zLGMLEYs7_0(.din(n17382), .dout(n17385));
    jdff dff_A_V1JJ2rO97_0(.din(n17385), .dout(n17388));
    jdff dff_A_4oZSJe060_0(.din(n17388), .dout(n17391));
    jdff dff_A_t118G6i42_0(.din(n17391), .dout(n17394));
    jdff dff_A_Ot5bP7Dg0_0(.din(n17394), .dout(n17397));
    jdff dff_A_Ty92eDGb9_0(.din(n17397), .dout(n17400));
    jdff dff_A_qKlU8vAu5_0(.din(n17400), .dout(n17403));
    jdff dff_A_qzBzlYFR7_0(.din(n17403), .dout(n17406));
    jdff dff_A_qOnaJgEF2_0(.din(n17406), .dout(n17409));
    jdff dff_A_rP1B7lWF8_0(.din(n17409), .dout(n17412));
    jdff dff_A_qbRmjG5t1_0(.din(n17412), .dout(n17415));
    jdff dff_A_CAN7PF2s2_0(.din(n17415), .dout(G534));
    jdff dff_A_uyVV29G02_1(.din(n5721), .dout(n17421));
    jdff dff_A_YpAS42Pd0_0(.din(n17421), .dout(n17424));
    jdff dff_A_aABiHqDV8_0(.din(n17424), .dout(n17427));
    jdff dff_A_wUqlU6bb6_0(.din(n17427), .dout(n17430));
    jdff dff_A_HpeNI6hu8_0(.din(n17430), .dout(n17433));
    jdff dff_A_31ifhgLe3_0(.din(n17433), .dout(n17436));
    jdff dff_A_20LL0kXl3_0(.din(n17436), .dout(n17439));
    jdff dff_A_5frTfrNj9_0(.din(n17439), .dout(n17442));
    jdff dff_A_MnRCGrLU2_0(.din(n17442), .dout(n17445));
    jdff dff_A_iyKzf2e81_0(.din(n17445), .dout(n17448));
    jdff dff_A_bHVODOSr4_0(.din(n17448), .dout(n17451));
    jdff dff_A_BgMe5zfd0_0(.din(n17451), .dout(n17454));
    jdff dff_A_IYQi4gKK1_0(.din(n17454), .dout(n17457));
    jdff dff_A_vyipA3Is1_0(.din(n17457), .dout(n17460));
    jdff dff_A_QQxLPPac5_0(.din(n17460), .dout(n17463));
    jdff dff_A_bYELoScb0_0(.din(n17463), .dout(n17466));
    jdff dff_A_zy7vFfa32_0(.din(n17466), .dout(n17469));
    jdff dff_A_JDIrwvVA2_0(.din(n17469), .dout(n17472));
    jdff dff_A_627Yje469_0(.din(n17472), .dout(n17475));
    jdff dff_A_TMA9OBaf5_0(.din(n17475), .dout(n17478));
    jdff dff_A_O8OwSJCu5_0(.din(n17478), .dout(n17481));
    jdff dff_A_wsyX4SW31_0(.din(n17481), .dout(n17484));
    jdff dff_A_Y70sezAz6_0(.din(n17484), .dout(n17487));
    jdff dff_A_dc3tr08t9_0(.din(n17487), .dout(n17490));
    jdff dff_A_C1dJ18Gh8_0(.din(n17490), .dout(n17493));
    jdff dff_A_XzuygA3z9_0(.din(n17493), .dout(G532));
    jdff dff_A_paBQc1dR5_1(.din(n5724), .dout(n17499));
    jdff dff_A_KrKWbOFh4_0(.din(n17499), .dout(n17502));
    jdff dff_A_owVCqCIt3_0(.din(n17502), .dout(n17505));
    jdff dff_A_8tjNKYJW7_0(.din(n17505), .dout(n17508));
    jdff dff_A_IKRWkruj3_0(.din(n17508), .dout(n17511));
    jdff dff_A_7ILXqpvi9_0(.din(n17511), .dout(n17514));
    jdff dff_A_9ssq8esx2_0(.din(n17514), .dout(n17517));
    jdff dff_A_mz5ZwWi41_0(.din(n17517), .dout(n17520));
    jdff dff_A_S3H3brTp1_0(.din(n17520), .dout(n17523));
    jdff dff_A_R3hJPeZ30_0(.din(n17523), .dout(n17526));
    jdff dff_A_M19Bz4np1_0(.din(n17526), .dout(n17529));
    jdff dff_A_1xd8j4TM9_0(.din(n17529), .dout(n17532));
    jdff dff_A_bjysYcGH5_0(.din(n17532), .dout(n17535));
    jdff dff_A_yFlYAY4Q1_0(.din(n17535), .dout(n17538));
    jdff dff_A_Itab8r2P7_0(.din(n17538), .dout(n17541));
    jdff dff_A_nxHJwfuq2_0(.din(n17541), .dout(n17544));
    jdff dff_A_qjpSuRHT0_0(.din(n17544), .dout(n17547));
    jdff dff_A_M21h6pYF5_0(.din(n17547), .dout(n17550));
    jdff dff_A_meqkVuQd2_0(.din(n17550), .dout(n17553));
    jdff dff_A_1SqBkC2z1_0(.din(n17553), .dout(n17556));
    jdff dff_A_mfmqXWB09_0(.din(n17556), .dout(n17559));
    jdff dff_A_wkbJbniV5_0(.din(n17559), .dout(n17562));
    jdff dff_A_bDCKCygv0_0(.din(n17562), .dout(n17565));
    jdff dff_A_tRoI4P0z5_0(.din(n17565), .dout(n17568));
    jdff dff_A_Ulamf9mu4_0(.din(n17568), .dout(n17571));
    jdff dff_A_DLzrrKos7_0(.din(n17571), .dout(G530));
    jdff dff_A_BhtDhst74_1(.din(n5727), .dout(n17577));
    jdff dff_A_PAVZXrKf0_0(.din(n17577), .dout(n17580));
    jdff dff_A_01cYpg8b6_0(.din(n17580), .dout(n17583));
    jdff dff_A_fajuVp6Z6_0(.din(n17583), .dout(n17586));
    jdff dff_A_DJXiWyPe2_0(.din(n17586), .dout(n17589));
    jdff dff_A_dlsyUagO4_0(.din(n17589), .dout(n17592));
    jdff dff_A_vmKx730D5_0(.din(n17592), .dout(n17595));
    jdff dff_A_0RmeoFv85_0(.din(n17595), .dout(n17598));
    jdff dff_A_IZaZ4JT98_0(.din(n17598), .dout(n17601));
    jdff dff_A_o7wAR7Kf5_0(.din(n17601), .dout(n17604));
    jdff dff_A_ZWrN8TAT6_0(.din(n17604), .dout(n17607));
    jdff dff_A_GC1pX1l39_0(.din(n17607), .dout(n17610));
    jdff dff_A_DAT3tjR14_0(.din(n17610), .dout(n17613));
    jdff dff_A_Lp3fWjAx2_0(.din(n17613), .dout(n17616));
    jdff dff_A_HhyK5uS78_0(.din(n17616), .dout(n17619));
    jdff dff_A_I6VdQDZF7_0(.din(n17619), .dout(n17622));
    jdff dff_A_sBPhlIxo5_0(.din(n17622), .dout(n17625));
    jdff dff_A_gZb17gAj1_0(.din(n17625), .dout(n17628));
    jdff dff_A_3eYdNwvV9_0(.din(n17628), .dout(n17631));
    jdff dff_A_hKabU6aP9_0(.din(n17631), .dout(n17634));
    jdff dff_A_GRmOsZCc2_0(.din(n17634), .dout(n17637));
    jdff dff_A_jOt2u3W90_0(.din(n17637), .dout(n17640));
    jdff dff_A_2nW35xZC6_0(.din(n17640), .dout(n17643));
    jdff dff_A_pEyMk4PZ2_0(.din(n17643), .dout(n17646));
    jdff dff_A_Ef2unXg22_0(.din(n17646), .dout(n17649));
    jdff dff_A_f6nhjreC0_0(.din(n17649), .dout(G528));
    jdff dff_A_xoVdo85w5_1(.din(n5730), .dout(n17655));
    jdff dff_A_5gDDdwws1_0(.din(n17655), .dout(n17658));
    jdff dff_A_tDSURJ8L5_0(.din(n17658), .dout(n17661));
    jdff dff_A_7T47Z8Ee6_0(.din(n17661), .dout(n17664));
    jdff dff_A_0qzoXbNm6_0(.din(n17664), .dout(n17667));
    jdff dff_A_emAtNjXO1_0(.din(n17667), .dout(n17670));
    jdff dff_A_Gm5iDwRD3_0(.din(n17670), .dout(n17673));
    jdff dff_A_ijIOBYxc4_0(.din(n17673), .dout(n17676));
    jdff dff_A_jFEJhcw94_0(.din(n17676), .dout(n17679));
    jdff dff_A_JVvijcYU1_0(.din(n17679), .dout(n17682));
    jdff dff_A_yGx7oG0K3_0(.din(n17682), .dout(n17685));
    jdff dff_A_FHiqnv7H8_0(.din(n17685), .dout(n17688));
    jdff dff_A_f0gM1s5W2_0(.din(n17688), .dout(n17691));
    jdff dff_A_4iHu8ezz9_0(.din(n17691), .dout(n17694));
    jdff dff_A_mJY6w7js8_0(.din(n17694), .dout(n17697));
    jdff dff_A_LD26rznv4_0(.din(n17697), .dout(n17700));
    jdff dff_A_HNHrvkNo8_0(.din(n17700), .dout(n17703));
    jdff dff_A_Qj9BCZR75_0(.din(n17703), .dout(n17706));
    jdff dff_A_5czEvGOu2_0(.din(n17706), .dout(n17709));
    jdff dff_A_nsgSRCgU3_0(.din(n17709), .dout(n17712));
    jdff dff_A_okbHxb314_0(.din(n17712), .dout(n17715));
    jdff dff_A_5ZmMUI1l1_0(.din(n17715), .dout(n17718));
    jdff dff_A_6hMGT60p9_0(.din(n17718), .dout(n17721));
    jdff dff_A_HuYc30OT2_0(.din(n17721), .dout(n17724));
    jdff dff_A_NbavnChT7_0(.din(n17724), .dout(n17727));
    jdff dff_A_xNJ98UHb0_0(.din(n17727), .dout(G526));
    jdff dff_A_7CNN2QGj1_1(.din(n5733), .dout(n17733));
    jdff dff_A_wPADSHmc3_0(.din(n17733), .dout(n17736));
    jdff dff_A_UfqHfyUg4_0(.din(n17736), .dout(n17739));
    jdff dff_A_XLoXWYXv6_0(.din(n17739), .dout(n17742));
    jdff dff_A_9CZaF95Y6_0(.din(n17742), .dout(n17745));
    jdff dff_A_fXX5esH14_0(.din(n17745), .dout(n17748));
    jdff dff_A_H6sED84P5_0(.din(n17748), .dout(n17751));
    jdff dff_A_ixSHJUKU4_0(.din(n17751), .dout(n17754));
    jdff dff_A_Ax5ViNf71_0(.din(n17754), .dout(n17757));
    jdff dff_A_xIk4ZfjZ1_0(.din(n17757), .dout(n17760));
    jdff dff_A_ww5h3tzY7_0(.din(n17760), .dout(n17763));
    jdff dff_A_T2WSgOqE8_0(.din(n17763), .dout(n17766));
    jdff dff_A_H7KwQJ684_0(.din(n17766), .dout(n17769));
    jdff dff_A_AB3GZso39_0(.din(n17769), .dout(n17772));
    jdff dff_A_tEJ9L1XR0_0(.din(n17772), .dout(n17775));
    jdff dff_A_XObD0KSJ3_0(.din(n17775), .dout(n17778));
    jdff dff_A_ftVRf9Jn2_0(.din(n17778), .dout(n17781));
    jdff dff_A_VfMZnpqv9_0(.din(n17781), .dout(n17784));
    jdff dff_A_CzQ4pz1a5_0(.din(n17784), .dout(n17787));
    jdff dff_A_OOAtbI1m4_0(.din(n17787), .dout(n17790));
    jdff dff_A_Gsx3K5yd6_0(.din(n17790), .dout(n17793));
    jdff dff_A_FESGzfjc1_0(.din(n17793), .dout(n17796));
    jdff dff_A_4E4cdKaC4_0(.din(n17796), .dout(n17799));
    jdff dff_A_gYgrfdEk4_0(.din(n17799), .dout(n17802));
    jdff dff_A_EVpZsa9A0_0(.din(n17802), .dout(n17805));
    jdff dff_A_kLXAngYK6_0(.din(n17805), .dout(G524));
    jdff dff_A_rfiYBFTn8_1(.din(n316), .dout(n17811));
    jdff dff_A_KBv17TNX9_0(.din(n17811), .dout(n17814));
    jdff dff_A_eYF8b48w9_0(.din(n17814), .dout(n17817));
    jdff dff_A_Bws8PJEh4_0(.din(n17817), .dout(n17820));
    jdff dff_A_3DAFSLe24_0(.din(n17820), .dout(n17823));
    jdff dff_A_EqiYcGl26_0(.din(n17823), .dout(n17826));
    jdff dff_A_kvlIc9Fz3_0(.din(n17826), .dout(n17829));
    jdff dff_A_6Z60N6TK4_0(.din(n17829), .dout(n17832));
    jdff dff_A_6FalZRrc5_0(.din(n17832), .dout(n17835));
    jdff dff_A_v7Zzebew6_0(.din(n17835), .dout(n17838));
    jdff dff_A_lDTvXDzZ3_0(.din(n17838), .dout(n17841));
    jdff dff_A_8yNCk5pb1_0(.din(n17841), .dout(n17844));
    jdff dff_A_HXlHmMDz8_0(.din(n17844), .dout(n17847));
    jdff dff_A_YAQm3VGj2_0(.din(n17847), .dout(n17850));
    jdff dff_A_TyTEpEEQ6_0(.din(n17850), .dout(n17853));
    jdff dff_A_GnILxcXe2_0(.din(n17853), .dout(n17856));
    jdff dff_A_BjlgeGGf3_0(.din(n17856), .dout(n17859));
    jdff dff_A_LWN4IjBz3_0(.din(n17859), .dout(n17862));
    jdff dff_A_7CQEVQDv5_0(.din(n17862), .dout(n17865));
    jdff dff_A_Svu2ui5v0_0(.din(n17865), .dout(n17868));
    jdff dff_A_5SUASKkG3_0(.din(n17868), .dout(n17871));
    jdff dff_A_vEzzzN135_0(.din(n17871), .dout(n17874));
    jdff dff_A_GvabwsAo3_0(.din(n17874), .dout(n17877));
    jdff dff_A_srrWgsu77_0(.din(n17877), .dout(n17880));
    jdff dff_A_o1tEZ4r95_0(.din(n17880), .dout(n17883));
    jdff dff_A_NhoOKTcF7_0(.din(n17883), .dout(G279));
    jdff dff_A_vzwKrL7w6_1(.din(n5736), .dout(n17889));
    jdff dff_A_6JOIMAZh5_0(.din(n17889), .dout(n17892));
    jdff dff_A_HXCK9GeG6_0(.din(n17892), .dout(n17895));
    jdff dff_A_jnAEY3hC4_0(.din(n17895), .dout(n17898));
    jdff dff_A_5T71wfnt9_0(.din(n17898), .dout(n17901));
    jdff dff_A_RSOKYoRU9_0(.din(n17901), .dout(n17904));
    jdff dff_A_kMdOAi0x2_0(.din(n17904), .dout(n17907));
    jdff dff_A_J3I9FHX88_0(.din(n17907), .dout(n17910));
    jdff dff_A_zerZj92j0_0(.din(n17910), .dout(n17913));
    jdff dff_A_pox6fFuC4_0(.din(n17913), .dout(n17916));
    jdff dff_A_Duz2K8qb1_0(.din(n17916), .dout(n17919));
    jdff dff_A_sCyRjIMc0_0(.din(n17919), .dout(n17922));
    jdff dff_A_cq5ftkKE6_0(.din(n17922), .dout(n17925));
    jdff dff_A_YLNZXz9w3_0(.din(n17925), .dout(n17928));
    jdff dff_A_iEgz1ea65_0(.din(n17928), .dout(n17931));
    jdff dff_A_cw8y85bi0_0(.din(n17931), .dout(n17934));
    jdff dff_A_Uslt2Quc2_0(.din(n17934), .dout(n17937));
    jdff dff_A_nczOkbvE2_0(.din(n17937), .dout(n17940));
    jdff dff_A_LMIHyfFj4_0(.din(n17940), .dout(n17943));
    jdff dff_A_6chGvKM88_0(.din(n17943), .dout(n17946));
    jdff dff_A_bRBAi5Lb3_0(.din(n17946), .dout(n17949));
    jdff dff_A_OW8nLXc88_0(.din(n17949), .dout(n17952));
    jdff dff_A_3TrrA0Ne9_0(.din(n17952), .dout(n17955));
    jdff dff_A_ISuiKvfN8_0(.din(n17955), .dout(n17958));
    jdff dff_A_ctXFwlbt2_0(.din(n17958), .dout(n17961));
    jdff dff_A_7eIriKKN8_0(.din(n17961), .dout(G436));
    jdff dff_A_FaNycJh43_1(.din(n5739), .dout(n17967));
    jdff dff_A_qGY3H2J69_0(.din(n17967), .dout(n17970));
    jdff dff_A_lsSkBHxA3_0(.din(n17970), .dout(n17973));
    jdff dff_A_GcliZzoZ7_0(.din(n17973), .dout(n17976));
    jdff dff_A_vV6ldDxr2_0(.din(n17976), .dout(n17979));
    jdff dff_A_YWZF2o7m3_0(.din(n17979), .dout(n17982));
    jdff dff_A_ySXUJJNC7_0(.din(n17982), .dout(n17985));
    jdff dff_A_HgFrOgpO1_0(.din(n17985), .dout(n17988));
    jdff dff_A_MCzTh2bB6_0(.din(n17988), .dout(n17991));
    jdff dff_A_KecxzNaP9_0(.din(n17991), .dout(n17994));
    jdff dff_A_BORnleMq9_0(.din(n17994), .dout(n17997));
    jdff dff_A_cssMt9s20_0(.din(n17997), .dout(n18000));
    jdff dff_A_ZnpVQHlJ1_0(.din(n18000), .dout(n18003));
    jdff dff_A_deleM0tD5_0(.din(n18003), .dout(n18006));
    jdff dff_A_ErLBn5y45_0(.din(n18006), .dout(n18009));
    jdff dff_A_55Q1owVA1_0(.din(n18009), .dout(n18012));
    jdff dff_A_LbLt0Dhv2_0(.din(n18012), .dout(n18015));
    jdff dff_A_LstWs4qX6_0(.din(n18015), .dout(n18018));
    jdff dff_A_NACdGWnd0_0(.din(n18018), .dout(n18021));
    jdff dff_A_O7Pr7R1k4_0(.din(n18021), .dout(n18024));
    jdff dff_A_GjOo3sNm4_0(.din(n18024), .dout(n18027));
    jdff dff_A_K2M5jAHP2_0(.din(n18027), .dout(n18030));
    jdff dff_A_MJuuir9n5_0(.din(n18030), .dout(n18033));
    jdff dff_A_robZoaqS9_0(.din(n18033), .dout(n18036));
    jdff dff_A_gAIBCOyk9_0(.din(n18036), .dout(n18039));
    jdff dff_A_AMKGO00a5_0(.din(n18039), .dout(G478));
    jdff dff_A_brqg9SVn2_1(.din(n5742), .dout(n18045));
    jdff dff_A_i2nClWBd8_0(.din(n18045), .dout(n18048));
    jdff dff_A_rjGy2gj30_0(.din(n18048), .dout(n18051));
    jdff dff_A_8a2xj6IU7_0(.din(n18051), .dout(n18054));
    jdff dff_A_SIGElxjj8_0(.din(n18054), .dout(n18057));
    jdff dff_A_wJTkngWn6_0(.din(n18057), .dout(n18060));
    jdff dff_A_mLbAkSGR0_0(.din(n18060), .dout(n18063));
    jdff dff_A_klxBYdW41_0(.din(n18063), .dout(n18066));
    jdff dff_A_Xbv4C9a58_0(.din(n18066), .dout(n18069));
    jdff dff_A_aoc4nmTr8_0(.din(n18069), .dout(n18072));
    jdff dff_A_ZSaE2QXU7_0(.din(n18072), .dout(n18075));
    jdff dff_A_266lQG9v2_0(.din(n18075), .dout(n18078));
    jdff dff_A_ACClf9oO2_0(.din(n18078), .dout(n18081));
    jdff dff_A_xt4hKMK18_0(.din(n18081), .dout(n18084));
    jdff dff_A_8EV2gJwp6_0(.din(n18084), .dout(n18087));
    jdff dff_A_0qYkfXI60_0(.din(n18087), .dout(n18090));
    jdff dff_A_3JpaDPRG0_0(.din(n18090), .dout(n18093));
    jdff dff_A_29vsu59F3_0(.din(n18093), .dout(n18096));
    jdff dff_A_9K2fRsf20_0(.din(n18096), .dout(n18099));
    jdff dff_A_wexf8Kp48_0(.din(n18099), .dout(n18102));
    jdff dff_A_MOslUsCL4_0(.din(n18102), .dout(n18105));
    jdff dff_A_wtQqCkoa2_0(.din(n18105), .dout(n18108));
    jdff dff_A_JpM7Yh8f2_0(.din(n18108), .dout(n18111));
    jdff dff_A_WozjK2822_0(.din(n18111), .dout(n18114));
    jdff dff_A_oR7RuUwk7_0(.din(n18114), .dout(n18117));
    jdff dff_A_UJXTa3yz1_0(.din(n18117), .dout(G522));
    jdff dff_A_ZwI2TXIA4_2(.din(n320), .dout(n18123));
    jdff dff_A_sYOBUnNc1_0(.din(n18123), .dout(n18126));
    jdff dff_A_SWDkKvin7_0(.din(n18126), .dout(n18129));
    jdff dff_A_JjIlIpCG1_0(.din(n18129), .dout(n18132));
    jdff dff_A_ABN2chsT9_0(.din(n18132), .dout(n18135));
    jdff dff_A_Btkxkv7A9_0(.din(n18135), .dout(n18138));
    jdff dff_A_cwgUJgkC7_0(.din(n18138), .dout(n18141));
    jdff dff_A_vipA9yt70_0(.din(n18141), .dout(n18144));
    jdff dff_A_OdKV93LJ2_0(.din(n18144), .dout(n18147));
    jdff dff_A_kSn5jDc07_0(.din(n18147), .dout(n18150));
    jdff dff_A_KNQPhlBV5_0(.din(n18150), .dout(n18153));
    jdff dff_A_ZrlN9XDj7_0(.din(n18153), .dout(n18156));
    jdff dff_A_qHJFyHS24_0(.din(n18156), .dout(n18159));
    jdff dff_A_8CNmKfhf2_0(.din(n18159), .dout(n18162));
    jdff dff_A_zWxyZbO43_0(.din(n18162), .dout(n18165));
    jdff dff_A_2c8CazQk6_0(.din(n18165), .dout(n18168));
    jdff dff_A_3Ah7ubNf7_0(.din(n18168), .dout(n18171));
    jdff dff_A_m0PycPBr2_0(.din(n18171), .dout(n18174));
    jdff dff_A_3errfxBV5_0(.din(n18174), .dout(n18177));
    jdff dff_A_4lcwrkSK1_0(.din(n18177), .dout(n18180));
    jdff dff_A_O2j4AT3g2_0(.din(n18180), .dout(n18183));
    jdff dff_A_Apx7J8mW7_0(.din(n18183), .dout(n18186));
    jdff dff_A_e7RAeC0K0_0(.din(n18186), .dout(n18189));
    jdff dff_A_QjToOTvY1_0(.din(n18189), .dout(n18192));
    jdff dff_A_tVxoQLMN0_0(.din(n18192), .dout(n18195));
    jdff dff_A_7lcWiGlO9_0(.din(n18195), .dout(G402));
    jdff dff_A_amYEkAj00_1(.din(n344), .dout(n18201));
    jdff dff_A_LaqWwdLI9_0(.din(n18201), .dout(n18204));
    jdff dff_A_AKECcuck3_0(.din(n18204), .dout(n18207));
    jdff dff_A_RpsUUWyQ1_0(.din(n18207), .dout(n18210));
    jdff dff_A_eROdEdx10_0(.din(n18210), .dout(n18213));
    jdff dff_A_4DHT6LpY4_0(.din(n18213), .dout(n18216));
    jdff dff_A_5mDj9NIa8_0(.din(n18216), .dout(n18219));
    jdff dff_A_bw0vr69i8_0(.din(n18219), .dout(n18222));
    jdff dff_A_dLmmBDjx3_0(.din(n18222), .dout(n18225));
    jdff dff_A_vPFBJJbJ9_0(.din(n18225), .dout(n18228));
    jdff dff_A_Twal4M3a4_0(.din(n18228), .dout(n18231));
    jdff dff_A_oqWc8lh36_0(.din(n18231), .dout(n18234));
    jdff dff_A_U6HvmVBJ8_0(.din(n18234), .dout(n18237));
    jdff dff_A_aoOGWk9v8_0(.din(n18237), .dout(n18240));
    jdff dff_A_1Jo9rpXr5_0(.din(n18240), .dout(n18243));
    jdff dff_A_xQ9nMkpX1_0(.din(n18243), .dout(n18246));
    jdff dff_A_5SbnuXRR1_0(.din(n18246), .dout(n18249));
    jdff dff_A_w3mJGjV52_0(.din(n18249), .dout(n18252));
    jdff dff_A_7gPHDzAO7_0(.din(n18252), .dout(n18255));
    jdff dff_A_fUfY2IBG8_0(.din(n18255), .dout(n18258));
    jdff dff_A_WkWstzRA6_0(.din(n18258), .dout(n18261));
    jdff dff_A_8QG85tXQ5_0(.din(n18261), .dout(n18264));
    jdff dff_A_rPwfwKyQ7_0(.din(n18264), .dout(n18267));
    jdff dff_A_GnEmrQDq6_0(.din(n18267), .dout(G404));
    jdff dff_A_t6zLtL210_1(.din(n368), .dout(n18273));
    jdff dff_A_0GahgdHp1_0(.din(n18273), .dout(n18276));
    jdff dff_A_jMA16JGn6_0(.din(n18276), .dout(n18279));
    jdff dff_A_TDTUcUn22_0(.din(n18279), .dout(n18282));
    jdff dff_A_jWjxuwBj5_0(.din(n18282), .dout(n18285));
    jdff dff_A_lkwW53Hb9_0(.din(n18285), .dout(n18288));
    jdff dff_A_WpFj8LLB2_0(.din(n18288), .dout(n18291));
    jdff dff_A_aolWF1GW7_0(.din(n18291), .dout(n18294));
    jdff dff_A_GWLXQRzp2_0(.din(n18294), .dout(n18297));
    jdff dff_A_qO5YtnWr3_0(.din(n18297), .dout(n18300));
    jdff dff_A_BSs8seSw3_0(.din(n18300), .dout(n18303));
    jdff dff_A_OWT6ucqT4_0(.din(n18303), .dout(n18306));
    jdff dff_A_z4W6vr4U3_0(.din(n18306), .dout(n18309));
    jdff dff_A_E9n4eXgP9_0(.din(n18309), .dout(n18312));
    jdff dff_A_w3jBFa2V8_0(.din(n18312), .dout(n18315));
    jdff dff_A_OYdpdVrd2_0(.din(n18315), .dout(n18318));
    jdff dff_A_7wJGjD7S5_0(.din(n18318), .dout(n18321));
    jdff dff_A_8KaPnuhh1_0(.din(n18321), .dout(n18324));
    jdff dff_A_eIuhuls23_0(.din(n18324), .dout(n18327));
    jdff dff_A_4UfwIdWz5_0(.din(n18327), .dout(n18330));
    jdff dff_A_6pgKHLx60_0(.din(n18330), .dout(n18333));
    jdff dff_A_uyafAuev0_0(.din(n18333), .dout(n18336));
    jdff dff_A_ZvUt2NIY0_0(.din(n18336), .dout(n18339));
    jdff dff_A_Chpxamw89_0(.din(n18339), .dout(G406));
    jdff dff_A_08FIgT3x3_1(.din(n392), .dout(n18345));
    jdff dff_A_DEWlQHHu2_0(.din(n18345), .dout(n18348));
    jdff dff_A_NMtfxNaz9_0(.din(n18348), .dout(n18351));
    jdff dff_A_QEoySopq9_0(.din(n18351), .dout(n18354));
    jdff dff_A_8Q0uVE093_0(.din(n18354), .dout(n18357));
    jdff dff_A_ZFv72X4T8_0(.din(n18357), .dout(n18360));
    jdff dff_A_CXac6MEm2_0(.din(n18360), .dout(n18363));
    jdff dff_A_DMK9C7R25_0(.din(n18363), .dout(n18366));
    jdff dff_A_LQkf1OU52_0(.din(n18366), .dout(n18369));
    jdff dff_A_1GojHfPY9_0(.din(n18369), .dout(n18372));
    jdff dff_A_qRdmqRbv7_0(.din(n18372), .dout(n18375));
    jdff dff_A_K6kgOyaC8_0(.din(n18375), .dout(n18378));
    jdff dff_A_z9ssNojK7_0(.din(n18378), .dout(n18381));
    jdff dff_A_D9iUZg1s9_0(.din(n18381), .dout(n18384));
    jdff dff_A_d5h4aF7y9_0(.din(n18384), .dout(n18387));
    jdff dff_A_p4SBo7ed9_0(.din(n18387), .dout(n18390));
    jdff dff_A_OUFQjWLF5_0(.din(n18390), .dout(n18393));
    jdff dff_A_GKB4SBDy1_0(.din(n18393), .dout(n18396));
    jdff dff_A_pBwVRTGm3_0(.din(n18396), .dout(n18399));
    jdff dff_A_Y2ftOXnw3_0(.din(n18399), .dout(n18402));
    jdff dff_A_rycyxBW90_0(.din(n18402), .dout(n18405));
    jdff dff_A_6Hi7eGz54_0(.din(n18405), .dout(n18408));
    jdff dff_A_cm03bSxK5_0(.din(n18408), .dout(n18411));
    jdff dff_A_HanoiqVF5_0(.din(n18411), .dout(G408));
    jdff dff_A_OYPAWhe44_1(.din(n416), .dout(n18417));
    jdff dff_A_Dp7qLDe60_0(.din(n18417), .dout(n18420));
    jdff dff_A_RQOGItHR2_0(.din(n18420), .dout(n18423));
    jdff dff_A_qsVKNdr56_0(.din(n18423), .dout(n18426));
    jdff dff_A_1VrXme1e0_0(.din(n18426), .dout(n18429));
    jdff dff_A_Z7DtqWKy9_0(.din(n18429), .dout(n18432));
    jdff dff_A_AyOK5qy39_0(.din(n18432), .dout(n18435));
    jdff dff_A_XHSITl1N6_0(.din(n18435), .dout(n18438));
    jdff dff_A_25gz9LWm6_0(.din(n18438), .dout(n18441));
    jdff dff_A_tMyhFtJO9_0(.din(n18441), .dout(n18444));
    jdff dff_A_CxaKyIIo8_0(.din(n18444), .dout(n18447));
    jdff dff_A_CnP9KI3A0_0(.din(n18447), .dout(n18450));
    jdff dff_A_zsbHjANn7_0(.din(n18450), .dout(n18453));
    jdff dff_A_8CoC8X014_0(.din(n18453), .dout(n18456));
    jdff dff_A_XhWbLnqH2_0(.din(n18456), .dout(n18459));
    jdff dff_A_T0i8zvlZ5_0(.din(n18459), .dout(n18462));
    jdff dff_A_Gqjgf0B03_0(.din(n18462), .dout(n18465));
    jdff dff_A_vMeWpli98_0(.din(n18465), .dout(n18468));
    jdff dff_A_Uz9TNndU9_0(.din(n18468), .dout(n18471));
    jdff dff_A_XvS0LSSn0_0(.din(n18471), .dout(n18474));
    jdff dff_A_PPBrGKr10_0(.din(n18474), .dout(n18477));
    jdff dff_A_rM2fcNiD2_0(.din(n18477), .dout(n18480));
    jdff dff_A_OP2oINcU6_0(.din(n18480), .dout(n18483));
    jdff dff_A_0x6LqtEa7_0(.din(n18483), .dout(G410));
    jdff dff_A_72jiinuu9_1(.din(n5745), .dout(n18489));
    jdff dff_A_9EfaEjWq2_0(.din(n18489), .dout(n18492));
    jdff dff_A_JJ9ymX5w3_0(.din(n18492), .dout(n18495));
    jdff dff_A_oIQSNchm2_0(.din(n18495), .dout(n18498));
    jdff dff_A_6GloHEU80_0(.din(n18498), .dout(n18501));
    jdff dff_A_dKoQ4bme0_0(.din(n18501), .dout(n18504));
    jdff dff_A_foZ7Xmps6_0(.din(n18504), .dout(n18507));
    jdff dff_A_hs7SzKHx5_0(.din(n18507), .dout(n18510));
    jdff dff_A_aABwAC8k3_0(.din(n18510), .dout(n18513));
    jdff dff_A_987uaKlJ6_0(.din(n18513), .dout(n18516));
    jdff dff_A_RIApDNOh1_0(.din(n18516), .dout(n18519));
    jdff dff_A_fFDtMKm58_0(.din(n18519), .dout(n18522));
endmodule

