// Benchmark "top" written by ABC on Thu May 28 22:02:41 2020

module rf_square ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \asquared[0] , \asquared[1] , \asquared[2] , \asquared[3] ,
    \asquared[4] , \asquared[5] , \asquared[6] , \asquared[7] ,
    \asquared[8] , \asquared[9] , \asquared[10] , \asquared[11] ,
    \asquared[12] , \asquared[13] , \asquared[14] , \asquared[15] ,
    \asquared[16] , \asquared[17] , \asquared[18] , \asquared[19] ,
    \asquared[20] , \asquared[21] , \asquared[22] , \asquared[23] ,
    \asquared[24] , \asquared[25] , \asquared[26] , \asquared[27] ,
    \asquared[28] , \asquared[29] , \asquared[30] , \asquared[31] ,
    \asquared[32] , \asquared[33] , \asquared[34] , \asquared[35] ,
    \asquared[36] , \asquared[37] , \asquared[38] , \asquared[39] ,
    \asquared[40] , \asquared[41] , \asquared[42] , \asquared[43] ,
    \asquared[44] , \asquared[45] , \asquared[46] , \asquared[47] ,
    \asquared[48] , \asquared[49] , \asquared[50] , \asquared[51] ,
    \asquared[52] , \asquared[53] , \asquared[54] , \asquared[55] ,
    \asquared[56] , \asquared[57] , \asquared[58] , \asquared[59] ,
    \asquared[60] , \asquared[61] , \asquared[62] , \asquared[63] ,
    \asquared[64] , \asquared[65] , \asquared[66] , \asquared[67] ,
    \asquared[68] , \asquared[69] , \asquared[70] , \asquared[71] ,
    \asquared[72] , \asquared[73] , \asquared[74] , \asquared[75] ,
    \asquared[76] , \asquared[77] , \asquared[78] , \asquared[79] ,
    \asquared[80] , \asquared[81] , \asquared[82] , \asquared[83] ,
    \asquared[84] , \asquared[85] , \asquared[86] , \asquared[87] ,
    \asquared[88] , \asquared[89] , \asquared[90] , \asquared[91] ,
    \asquared[92] , \asquared[93] , \asquared[94] , \asquared[95] ,
    \asquared[96] , \asquared[97] , \asquared[98] , \asquared[99] ,
    \asquared[100] , \asquared[101] , \asquared[102] , \asquared[103] ,
    \asquared[104] , \asquared[105] , \asquared[106] , \asquared[107] ,
    \asquared[108] , \asquared[109] , \asquared[110] , \asquared[111] ,
    \asquared[112] , \asquared[113] , \asquared[114] , \asquared[115] ,
    \asquared[116] , \asquared[117] , \asquared[118] , \asquared[119] ,
    \asquared[120] , \asquared[121] , \asquared[122] , \asquared[123] ,
    \asquared[124] , \asquared[125] , \asquared[126] , \asquared[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ;
  output \asquared[0] , \asquared[1] , \asquared[2] , \asquared[3] ,
    \asquared[4] , \asquared[5] , \asquared[6] , \asquared[7] ,
    \asquared[8] , \asquared[9] , \asquared[10] , \asquared[11] ,
    \asquared[12] , \asquared[13] , \asquared[14] , \asquared[15] ,
    \asquared[16] , \asquared[17] , \asquared[18] , \asquared[19] ,
    \asquared[20] , \asquared[21] , \asquared[22] , \asquared[23] ,
    \asquared[24] , \asquared[25] , \asquared[26] , \asquared[27] ,
    \asquared[28] , \asquared[29] , \asquared[30] , \asquared[31] ,
    \asquared[32] , \asquared[33] , \asquared[34] , \asquared[35] ,
    \asquared[36] , \asquared[37] , \asquared[38] , \asquared[39] ,
    \asquared[40] , \asquared[41] , \asquared[42] , \asquared[43] ,
    \asquared[44] , \asquared[45] , \asquared[46] , \asquared[47] ,
    \asquared[48] , \asquared[49] , \asquared[50] , \asquared[51] ,
    \asquared[52] , \asquared[53] , \asquared[54] , \asquared[55] ,
    \asquared[56] , \asquared[57] , \asquared[58] , \asquared[59] ,
    \asquared[60] , \asquared[61] , \asquared[62] , \asquared[63] ,
    \asquared[64] , \asquared[65] , \asquared[66] , \asquared[67] ,
    \asquared[68] , \asquared[69] , \asquared[70] , \asquared[71] ,
    \asquared[72] , \asquared[73] , \asquared[74] , \asquared[75] ,
    \asquared[76] , \asquared[77] , \asquared[78] , \asquared[79] ,
    \asquared[80] , \asquared[81] , \asquared[82] , \asquared[83] ,
    \asquared[84] , \asquared[85] , \asquared[86] , \asquared[87] ,
    \asquared[88] , \asquared[89] , \asquared[90] , \asquared[91] ,
    \asquared[92] , \asquared[93] , \asquared[94] , \asquared[95] ,
    \asquared[96] , \asquared[97] , \asquared[98] , \asquared[99] ,
    \asquared[100] , \asquared[101] , \asquared[102] , \asquared[103] ,
    \asquared[104] , \asquared[105] , \asquared[106] , \asquared[107] ,
    \asquared[108] , \asquared[109] , \asquared[110] , \asquared[111] ,
    \asquared[112] , \asquared[113] , \asquared[114] , \asquared[115] ,
    \asquared[116] , \asquared[117] , \asquared[118] , \asquared[119] ,
    \asquared[120] , \asquared[121] , \asquared[122] , \asquared[123] ,
    \asquared[124] , \asquared[125] , \asquared[126] , \asquared[127] ;
  wire n193, n195, n197, n198, n199, n200, n201, n202, n203, n204, n206,
    n207, n208, n209, n210, n212, n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n231, n232,
    n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n245,
    n246, n247, n248, n249, n250, n252, n253, n254, n255, n256, n257, n258,
    n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
    n271, n272, n273, n274, n275, n276, n277, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
    n296, n297, n298, n299, n300, n301, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
    n358, n359, n360, n361, n362, n363, n364, n366, n367, n368, n369, n370,
    n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
    n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
    n407, n408, n409, n410, n411, n412, n413, n414, n415, n417, n418, n419,
    n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
    n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n461, n462, n463, n464, n465, n466, n467, n468,
    n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
    n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
    n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n521, n522, n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
    n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
    n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
    n566, n567, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
    n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n618, n619, n620, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
    n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
    n676, n677, n678, n679, n680, n681, n682, n684, n685, n686, n687, n688,
    n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
    n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
    n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
    n749, n750, n751, n752, n753, n754, n755, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n815, n816, n817, n818, n819, n820, n821, n822,
    n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
    n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
    n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
    n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
    n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
    n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n900, n901, n902, n903, n904, n905, n906, n907,
    n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
    n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
    n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
    n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
    n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
    n968, n969, n970, n971, n972, n974, n975, n976, n977, n978, n979, n980,
    n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
    n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
    n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
    n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
    n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
    n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
    n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
    n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
    n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
    n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
    n1135, n1136, n1137, n1138, n1140, n1141, n1142, n1143, n1144, n1145,
    n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
    n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
    n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
    n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
    n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
    n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
    n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
    n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
    n1307, n1308, n1309, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
    n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
    n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
    n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
    n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
    n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
    n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
    n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
    n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
    n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
    n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
    n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
    n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
    n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
    n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
    n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
    n1499, n1500, n1501, n1502, n1503, n1504, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
    n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
    n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
    n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
    n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
    n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
    n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
    n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
    n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
    n1610, n1611, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
    n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
    n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
    n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
    n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
    n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
    n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
    n1711, n1712, n1713, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
    n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
    n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
    n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
    n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
    n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
    n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
    n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
    n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
    n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
    n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
    n1822, n1823, n1824, n1825, n1826, n1827, n1829, n1830, n1831, n1832,
    n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
    n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
    n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
    n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
    n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
    n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
    n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
    n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
    n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
    n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
    n1933, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
    n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
    n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
    n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
    n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
    n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
    n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
    n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
    n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
    n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
    n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
    n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2064,
    n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
    n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
    n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
    n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
    n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
    n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
    n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
    n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
    n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
    n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
    n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
    n2175, n2176, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
    n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
    n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
    n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
    n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
    n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
    n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
    n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
    n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
    n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
    n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
    n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
    n2296, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
    n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
    n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
    n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
    n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
    n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
    n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
    n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
    n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
    n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
    n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
    n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
    n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
    n2427, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
    n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
    n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
    n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
    n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
    n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
    n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
    n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
    n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
    n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
    n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
    n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
    n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
    n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2568,
    n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
    n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
    n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
    n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
    n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
    n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
    n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
    n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
    n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
    n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
    n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
    n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
    n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2697, n2698, n2699,
    n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
    n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
    n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
    n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
    n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
    n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
    n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
    n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
    n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
    n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
    n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
    n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
    n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2860,
    n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
    n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
    n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
    n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
    n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
    n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
    n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
    n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
    n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
    n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
    n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
    n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
    n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
    n2991, n2992, n2993, n2994, n2996, n2997, n2998, n2999, n3000, n3001,
    n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
    n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
    n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
    n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
    n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
    n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
    n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
    n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
    n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
    n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
    n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
    n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
    n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
    n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
    n3142, n3143, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
    n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
    n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
    n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
    n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
    n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
    n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
    n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
    n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
    n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
    n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
    n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
    n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
    n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
    n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
    n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
    n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
    n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
    n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
    n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
    n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
    n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
    n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
    n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
    n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
    n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
    n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
    n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
    n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
    n3434, n3435, n3436, n3437, n3438, n3440, n3441, n3442, n3443, n3444,
    n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
    n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
    n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
    n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
    n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
    n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
    n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
    n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
    n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
    n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
    n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
    n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
    n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
    n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
    n3585, n3586, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
    n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
    n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
    n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
    n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
    n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
    n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
    n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
    n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
    n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
    n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
    n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
    n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
    n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
    n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
    n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
    n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
    n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3764, n3765, n3766,
    n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
    n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
    n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
    n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
    n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
    n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
    n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
    n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
    n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
    n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
    n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
    n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
    n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
    n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
    n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
    n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
    n3927, n3928, n3929, n3930, n3931, n3933, n3934, n3935, n3936, n3937,
    n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
    n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
    n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
    n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
    n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
    n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
    n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
    n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
    n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
    n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
    n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
    n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
    n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
    n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
    n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
    n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
    n4098, n4099, n4100, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
    n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
    n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
    n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
    n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
    n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
    n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
    n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
    n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
    n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
    n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
    n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
    n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
    n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
    n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
    n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
    n4259, n4260, n4261, n4262, n4263, n4264, n4266, n4267, n4268, n4269,
    n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
    n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
    n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
    n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
    n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
    n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
    n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
    n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
    n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
    n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
    n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
    n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
    n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
    n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
    n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
    n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
    n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
    n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
    n4450, n4451, n4452, n4453, n4454, n4456, n4457, n4458, n4459, n4460,
    n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
    n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
    n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
    n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
    n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
    n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
    n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
    n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
    n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
    n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
    n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
    n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
    n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
    n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
    n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
    n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4620, n4621,
    n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
    n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
    n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
    n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
    n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
    n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
    n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
    n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
    n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
    n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
    n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
    n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
    n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
    n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
    n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
    n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
    n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
    n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
    n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
    n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
    n4822, n4823, n4824, n4825, n4827, n4828, n4829, n4830, n4831, n4832,
    n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
    n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
    n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
    n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
    n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
    n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
    n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
    n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
    n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
    n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
    n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
    n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
    n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
    n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
    n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
    n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
    n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
    n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5011, n5012, n5013,
    n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
    n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
    n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
    n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
    n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
    n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
    n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
    n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
    n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
    n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
    n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
    n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
    n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
    n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
    n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
    n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
    n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
    n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
    n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
    n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5212, n5213, n5214,
    n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
    n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
    n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
    n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
    n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
    n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
    n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
    n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
    n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
    n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
    n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
    n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
    n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
    n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
    n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
    n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
    n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
    n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
    n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
    n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5413, n5414, n5415,
    n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
    n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
    n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
    n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
    n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
    n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
    n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
    n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
    n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
    n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
    n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
    n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
    n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
    n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
    n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
    n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
    n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
    n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
    n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
    n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
    n5616, n5617, n5618, n5619, n5620, n5622, n5623, n5624, n5625, n5626,
    n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
    n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
    n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
    n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
    n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
    n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
    n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
    n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
    n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
    n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
    n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
    n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
    n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
    n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
    n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
    n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
    n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
    n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
    n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
    n5817, n5818, n5819, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
    n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
    n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
    n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
    n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
    n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
    n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
    n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
    n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
    n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
    n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
    n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
    n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
    n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
    n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
    n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
    n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
    n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
    n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
    n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
    n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
    n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
    n6038, n6039, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
    n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
    n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
    n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
    n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
    n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
    n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
    n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
    n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
    n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
    n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
    n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
    n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
    n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
    n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
    n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
    n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
    n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
    n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
    n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
    n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
    n6249, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
    n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
    n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
    n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
    n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
    n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
    n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
    n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
    n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
    n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
    n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
    n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
    n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
    n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
    n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
    n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
    n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
    n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
    n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
    n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
    n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
    n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
    n6470, n6471, n6472, n6473, n6475, n6476, n6477, n6478, n6479, n6480,
    n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
    n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
    n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
    n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
    n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
    n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
    n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
    n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
    n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
    n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
    n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
    n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
    n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
    n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
    n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
    n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
    n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
    n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
    n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
    n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6681,
    n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
    n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
    n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
    n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
    n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
    n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
    n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
    n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
    n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
    n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
    n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
    n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
    n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
    n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
    n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
    n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
    n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
    n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
    n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
    n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
    n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
    n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
    n6902, n6903, n6904, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
    n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
    n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
    n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
    n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
    n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
    n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
    n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
    n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
    n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
    n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
    n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
    n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
    n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
    n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
    n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
    n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
    n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
    n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
    n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
    n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
    n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7121, n7122, n7123,
    n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
    n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
    n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
    n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
    n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
    n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
    n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
    n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
    n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
    n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
    n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
    n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
    n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
    n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
    n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
    n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
    n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
    n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
    n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
    n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
    n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
    n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
    n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
    n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
    n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7373, n7374,
    n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
    n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
    n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
    n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
    n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
    n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
    n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
    n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
    n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
    n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
    n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
    n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
    n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
    n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
    n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
    n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
    n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
    n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
    n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
    n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
    n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
    n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
    n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
    n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
    n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
    n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
    n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
    n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
    n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
    n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
    n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
    n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
    n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
    n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
    n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
    n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
    n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
    n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
    n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
    n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
    n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
    n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
    n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
    n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
    n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
    n7826, n7827, n7828, n7829, n7831, n7832, n7833, n7834, n7835, n7836,
    n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
    n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
    n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
    n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
    n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
    n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
    n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
    n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
    n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
    n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
    n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
    n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
    n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
    n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
    n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
    n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
    n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
    n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
    n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
    n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
    n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
    n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
    n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8066, n8067,
    n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
    n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
    n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
    n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
    n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
    n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
    n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
    n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
    n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
    n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
    n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
    n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
    n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
    n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
    n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
    n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
    n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
    n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
    n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
    n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
    n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
    n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
    n8288, n8289, n8290, n8291, n8293, n8294, n8295, n8296, n8297, n8298,
    n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
    n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
    n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
    n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
    n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
    n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
    n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
    n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
    n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
    n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
    n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
    n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
    n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
    n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
    n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
    n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
    n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
    n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
    n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
    n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
    n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
    n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
    n8519, n8520, n8521, n8522, n8523, n8524, n8526, n8527, n8528, n8529,
    n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
    n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
    n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
    n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
    n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
    n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
    n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
    n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
    n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
    n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
    n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
    n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
    n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
    n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
    n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
    n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
    n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
    n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
    n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
    n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
    n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
    n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
    n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
    n8760, n8761, n8762, n8763, n8765, n8766, n8767, n8768, n8769, n8770,
    n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
    n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
    n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
    n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
    n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
    n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
    n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
    n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
    n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
    n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
    n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
    n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
    n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
    n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
    n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
    n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
    n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
    n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
    n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
    n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
    n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8981,
    n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
    n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
    n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
    n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
    n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
    n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
    n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
    n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
    n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
    n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
    n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
    n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
    n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
    n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
    n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
    n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
    n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
    n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
    n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
    n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
    n9182, n9183, n9184, n9185, n9186, n9187, n9189, n9190, n9191, n9192,
    n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
    n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
    n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
    n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
    n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
    n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
    n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
    n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
    n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
    n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
    n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
    n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
    n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
    n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
    n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
    n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
    n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
    n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
    n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
    n9383, n9384, n9385, n9386, n9387, n9388, n9390, n9391, n9392, n9393,
    n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
    n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
    n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
    n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
    n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
    n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
    n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
    n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
    n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
    n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
    n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
    n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
    n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
    n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
    n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
    n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
    n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
    n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
    n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
    n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
    n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
    n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
    n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
    n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
    n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
    n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
    n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
    n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
    n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
    n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
    n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
    n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
    n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
    n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
    n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
    n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
    n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
    n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
    n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
    n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
    n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9805,
    n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
    n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
    n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
    n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
    n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
    n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
    n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
    n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
    n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
    n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
    n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
    n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
    n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
    n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
    n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
    n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
    n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
    n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
    n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
    n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
    n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
    n10014, n10015, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
    n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
    n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
    n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
    n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
    n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
    n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
    n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
    n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
    n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
    n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
    n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
    n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
    n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
    n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
    n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
    n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
    n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
    n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
    n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
    n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
    n10204, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
    n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
    n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
    n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
    n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
    n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
    n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
    n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
    n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
    n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
    n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
    n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
    n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
    n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
    n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
    n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
    n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
    n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
    n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
    n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
    n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
    n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
    n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
    n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
    n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
    n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
    n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
    n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
    n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
    n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
    n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
    n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
    n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
    n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
    n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
    n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
    n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
    n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
    n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
    n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
    n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
    n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
    n10584, n10585, n10586, n10587, n10588, n10589, n10591, n10592, n10593,
    n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
    n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
    n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
    n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
    n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
    n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
    n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
    n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
    n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
    n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
    n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
    n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
    n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
    n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
    n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
    n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
    n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
    n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
    n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
    n10765, n10766, n10767, n10768, n10769, n10771, n10772, n10773, n10774,
    n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
    n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
    n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
    n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
    n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
    n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
    n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
    n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
    n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
    n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
    n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
    n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
    n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
    n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
    n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
    n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
    n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
    n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
    n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
    n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
    n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
    n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
    n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
    n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
    n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
    n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
    n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
    n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
    n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
    n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
    n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
    n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
    n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
    n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
    n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
    n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
    n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
    n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
    n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11126, n11127,
    n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
    n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
    n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
    n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
    n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
    n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
    n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
    n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
    n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
    n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
    n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
    n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
    n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
    n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
    n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
    n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
    n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
    n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
    n11290, n11291, n11292, n11293, n11294, n11296, n11297, n11298, n11299,
    n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
    n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
    n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
    n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
    n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
    n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
    n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
    n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
    n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
    n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
    n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
    n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
    n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
    n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
    n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
    n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
    n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
    n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
    n11462, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
    n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
    n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
    n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
    n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
    n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
    n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
    n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
    n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
    n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
    n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
    n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
    n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
    n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
    n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
    n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
    n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
    n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
    n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11633, n11634,
    n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
    n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
    n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
    n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
    n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
    n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
    n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
    n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
    n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
    n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
    n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
    n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
    n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
    n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
    n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
    n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
    n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
    n11788, n11789, n11790, n11791, n11792, n11793, n11795, n11796, n11797,
    n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
    n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
    n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
    n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
    n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
    n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
    n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
    n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
    n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
    n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
    n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
    n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
    n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
    n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
    n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
    n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
    n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
    n11951, n11952, n11953, n11955, n11956, n11957, n11958, n11959, n11960,
    n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
    n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
    n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
    n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
    n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
    n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
    n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
    n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
    n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
    n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
    n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
    n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
    n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
    n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
    n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
    n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
    n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
    n12114, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
    n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
    n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
    n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
    n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
    n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
    n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
    n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
    n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
    n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
    n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
    n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
    n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
    n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
    n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
    n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
    n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
    n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
    n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
    n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
    n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
    n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
    n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
    n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
    n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
    n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
    n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
    n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
    n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
    n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
    n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
    n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
    n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
    n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12422,
    n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
    n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
    n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
    n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
    n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
    n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
    n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
    n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
    n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
    n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
    n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
    n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
    n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
    n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
    n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
    n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
    n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
    n12576, n12577, n12578, n12579, n12581, n12582, n12583, n12584, n12585,
    n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
    n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
    n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
    n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
    n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
    n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
    n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
    n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
    n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
    n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
    n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
    n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
    n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
    n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
    n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12720, n12721,
    n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
    n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
    n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
    n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
    n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
    n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
    n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
    n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
    n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
    n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
    n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
    n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
    n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
    n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
    n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12857,
    n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
    n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
    n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
    n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
    n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
    n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
    n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
    n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
    n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
    n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
    n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
    n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
    n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
    n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
    n12984, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
    n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
    n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
    n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
    n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
    n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
    n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
    n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
    n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
    n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
    n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
    n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
    n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
    n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
    n13111, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
    n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
    n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
    n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
    n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
    n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
    n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
    n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
    n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
    n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
    n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
    n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
    n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
    n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
    n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
    n13247, n13248, n13249, n13250, n13252, n13253, n13254, n13255, n13256,
    n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
    n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
    n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
    n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
    n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
    n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
    n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
    n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
    n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
    n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
    n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
    n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
    n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
    n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
    n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
    n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
    n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
    n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
    n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
    n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
    n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
    n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
    n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
    n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
    n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
    n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
    n13492, n13493, n13494, n13495, n13496, n13498, n13499, n13500, n13501,
    n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
    n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
    n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
    n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
    n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
    n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
    n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
    n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
    n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
    n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
    n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
    n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
    n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
    n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
    n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
    n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
    n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
    n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
    n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
    n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
    n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
    n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
    n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
    n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
    n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
    n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
    n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
    n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
    n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
    n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
    n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
    n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
    n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
    n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
    n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
    n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
    n13828, n13829, n13830, n13831, n13833, n13834, n13835, n13836, n13837,
    n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
    n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
    n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
    n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
    n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
    n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
    n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
    n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
    n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
    n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
    n13928, n13929, n13930, n13931, n13932, n13933, n13935, n13936, n13937,
    n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
    n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
    n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
    n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
    n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
    n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
    n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
    n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
    n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
    n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
    n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
    n14037, n14038, n14039, n14040, n14042, n14043, n14044, n14045, n14046,
    n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
    n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
    n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
    n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
    n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
    n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
    n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
    n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
    n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
    n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
    n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14146,
    n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
    n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
    n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
    n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
    n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
    n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
    n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
    n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
    n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
    n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
    n14237, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
    n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
    n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
    n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
    n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
    n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
    n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
    n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
    n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
    n14319, n14320, n14321, n14322, n14323, n14324, n14326, n14327, n14328,
    n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
    n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
    n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
    n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
    n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
    n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
    n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
    n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
    n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
    n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14418, n14419,
    n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
    n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
    n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
    n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
    n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
    n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
    n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
    n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
    n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
    n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
    n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
    n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
    n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
    n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
    n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
    n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
    n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14573, n14574,
    n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
    n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
    n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
    n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
    n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
    n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
    n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
    n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14647,
    n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
    n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
    n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
    n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
    n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
    n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
    n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
    n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
    n14720, n14721, n14722, n14724, n14725, n14726, n14727, n14728, n14729,
    n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
    n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
    n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
    n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
    n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
    n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
    n14784, n14785, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
    n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
    n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
    n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
    n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
    n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
    n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
    n14848, n14849, n14850, n14852, n14853, n14854, n14855, n14856, n14857,
    n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
    n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
    n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
    n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
    n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
    n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
    n14912, n14913, n14914, n14916, n14917, n14918, n14919, n14920, n14921,
    n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
    n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
    n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
    n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
    n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
    n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14976,
    n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
    n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
    n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
    n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
    n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
    n15022, n15023, n15024, n15026, n15027, n15028, n15029, n15030, n15031,
    n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
    n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
    n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
    n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
    n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15076, n15077,
    n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
    n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
    n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
    n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
    n15114, n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
    n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
    n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
    n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
    n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15160,
    n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
    n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
    n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
    n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15197,
    n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
    n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
    n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
    n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
    n15234, n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
    n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
    n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
    n15262, n15263, n15264, n15265, n15267, n15268, n15269, n15270, n15271,
    n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
    n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
    n15290, n15291, n15292, n15293, n15295, n15296, n15297, n15298, n15299,
    n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
    n15309, n15310, n15311, n15312, n15313, n15314, n15316, n15317, n15318,
    n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
    n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
    n15337, n15338, n15339, n15341, n15342, n15343, n15344, n15345, n15346,
    n15347, n15348, n15349, n15350, n15351, n15353, n15354, n15355, n15356,
    n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
    n15366, n15368, n15369, n15370, n15371, n15373;
  zero g00000(.dout(\asquared[1] ));
  jnot g00001(.din(\a[0] ), .dout(n193));
  jand g00002(.dina(\a[1] ), .dinb(n193), .dout(\asquared[2] ));
  jxor g00003(.dina(\a[2] ), .dinb(\a[1] ), .dout(n195));
  jand g00004(.dina(n195), .dinb(\a[0] ), .dout(\asquared[3] ));
  jand g00005(.dina(\a[3] ), .dinb(\a[2] ), .dout(n197));
  jand g00006(.dina(n197), .dinb(\a[0] ), .dout(n198));
  jnot g00007(.din(n198), .dout(n199));
  jnot g00008(.din(\a[1] ), .dout(n200));
  jand g00009(.dina(\a[2] ), .dinb(n200), .dout(n201));
  jor  g00010(.dina(\a[3] ), .dinb(\a[2] ), .dout(n202));
  jand g00011(.dina(n202), .dinb(\a[0] ), .dout(n203));
  jor  g00012(.dina(n203), .dinb(n201), .dout(n204));
  jand g00013(.dina(n204), .dinb(n199), .dout(\asquared[4] ));
  jand g00014(.dina(\a[2] ), .dinb(\a[1] ), .dout(n206));
  jand g00015(.dina(\a[3] ), .dinb(\a[1] ), .dout(n207));
  jand g00016(.dina(\a[4] ), .dinb(\a[0] ), .dout(n208));
  jxor g00017(.dina(n208), .dinb(n207), .dout(n209));
  jxor g00018(.dina(n209), .dinb(n206), .dout(n210));
  jxor g00019(.dina(n210), .dinb(n198), .dout(\asquared[5] ));
  jand g00020(.dina(n208), .dinb(n207), .dout(n212));
  jand g00021(.dina(\a[4] ), .dinb(\a[1] ), .dout(n213));
  jand g00022(.dina(\a[5] ), .dinb(\a[0] ), .dout(n214));
  jor  g00023(.dina(n214), .dinb(n213), .dout(n215));
  jnot g00024(.din(\a[4] ), .dout(n216));
  jor  g00025(.dina(n216), .dinb(n193), .dout(n217));
  jnot g00026(.din(\a[5] ), .dout(n218));
  jor  g00027(.dina(n218), .dinb(n200), .dout(n219));
  jor  g00028(.dina(n219), .dinb(n217), .dout(n220));
  jand g00029(.dina(n220), .dinb(n215), .dout(n221));
  jxor g00030(.dina(n221), .dinb(n212), .dout(n222));
  jnot g00031(.din(\a[2] ), .dout(n223));
  jand g00032(.dina(\a[3] ), .dinb(n223), .dout(n224));
  jxor g00033(.dina(n224), .dinb(n222), .dout(n225));
  jor  g00034(.dina(n209), .dinb(n206), .dout(n226));
  jand g00035(.dina(n209), .dinb(n206), .dout(n227));
  jor  g00036(.dina(n227), .dinb(n198), .dout(n228));
  jand g00037(.dina(n228), .dinb(n226), .dout(n229));
  jxor g00038(.dina(n229), .dinb(n225), .dout(\asquared[6] ));
  jand g00039(.dina(\a[4] ), .dinb(\a[2] ), .dout(n231));
  jnot g00040(.din(n231), .dout(n232));
  jand g00041(.dina(n232), .dinb(n219), .dout(n233));
  jand g00042(.dina(\a[5] ), .dinb(\a[2] ), .dout(n234));
  jand g00043(.dina(n234), .dinb(n213), .dout(n235));
  jor  g00044(.dina(n235), .dinb(n233), .dout(n236));
  jand g00045(.dina(\a[6] ), .dinb(\a[0] ), .dout(n237));
  jor  g00046(.dina(n237), .dinb(n197), .dout(n238));
  jnot g00047(.din(n238), .dout(n239));
  jand g00048(.dina(n198), .dinb(\a[6] ), .dout(n240));
  jor  g00049(.dina(n240), .dinb(n239), .dout(n241));
  jxor g00050(.dina(n241), .dinb(n236), .dout(n242));
  jnot g00051(.din(n220), .dout(n243));
  jor  g00052(.dina(n212), .dinb(n243), .dout(n245));
  jxor g00053(.dina(n245), .dinb(n242), .dout(n246));
  jand g00054(.dina(n224), .dinb(n222), .dout(n247));
  jor  g00055(.dina(n224), .dinb(n222), .dout(n248));
  jand g00056(.dina(n229), .dinb(n248), .dout(n249));
  jor  g00057(.dina(n249), .dinb(n247), .dout(n250));
  jxor g00058(.dina(n250), .dinb(n246), .dout(\asquared[7] ));
  jnot g00059(.din(n240), .dout(n252));
  jor  g00060(.dina(n241), .dinb(n236), .dout(n253));
  jand g00061(.dina(n253), .dinb(n252), .dout(n254));
  jnot g00062(.din(n254), .dout(n255));
  jand g00063(.dina(\a[6] ), .dinb(\a[1] ), .dout(n256));
  jxor g00064(.dina(n256), .dinb(n216), .dout(n257));
  jnot g00065(.din(n257), .dout(n258));
  jor  g00066(.dina(n258), .dinb(n235), .dout(n259));
  jnot g00067(.din(\a[6] ), .dout(n260));
  jand g00068(.dina(n235), .dinb(n260), .dout(n261));
  jnot g00069(.din(n261), .dout(n262));
  jand g00070(.dina(n262), .dinb(n259), .dout(n263));
  jxor g00071(.dina(n263), .dinb(n255), .dout(n264));
  jand g00072(.dina(\a[7] ), .dinb(\a[0] ), .dout(n265));
  jand g00073(.dina(\a[4] ), .dinb(\a[3] ), .dout(n266));
  jor  g00074(.dina(n266), .dinb(n234), .dout(n267));
  jand g00075(.dina(\a[5] ), .dinb(\a[3] ), .dout(n268));
  jand g00076(.dina(n268), .dinb(n231), .dout(n269));
  jnot g00077(.din(n269), .dout(n270));
  jand g00078(.dina(n270), .dinb(n267), .dout(n271));
  jxor g00079(.dina(n271), .dinb(n265), .dout(n272));
  jxor g00080(.dina(n272), .dinb(n264), .dout(n273));
  jand g00081(.dina(n245), .dinb(n242), .dout(n274));
  jor  g00082(.dina(n245), .dinb(n242), .dout(n275));
  jand g00083(.dina(n250), .dinb(n275), .dout(n276));
  jor  g00084(.dina(n276), .dinb(n274), .dout(n277));
  jxor g00085(.dina(n277), .dinb(n273), .dout(\asquared[8] ));
  jand g00086(.dina(n263), .dinb(n255), .dout(n279));
  jor  g00087(.dina(n279), .dinb(n261), .dout(n280));
  jand g00088(.dina(n271), .dinb(n265), .dout(n281));
  jor  g00089(.dina(n281), .dinb(n269), .dout(n282));
  jand g00090(.dina(\a[7] ), .dinb(\a[1] ), .dout(n283));
  jxor g00091(.dina(n283), .dinb(n268), .dout(n284));
  jxor g00092(.dina(n284), .dinb(n282), .dout(n285));
  jand g00093(.dina(n256), .dinb(\a[4] ), .dout(n286));
  jand g00094(.dina(\a[8] ), .dinb(\a[0] ), .dout(n287));
  jand g00095(.dina(\a[6] ), .dinb(\a[2] ), .dout(n288));
  jor  g00096(.dina(n288), .dinb(n287), .dout(n289));
  jnot g00097(.din(n289), .dout(n290));
  jand g00098(.dina(\a[8] ), .dinb(\a[2] ), .dout(n291));
  jand g00099(.dina(n291), .dinb(n237), .dout(n292));
  jor  g00100(.dina(n292), .dinb(n290), .dout(n293));
  jxor g00101(.dina(n293), .dinb(n286), .dout(n294));
  jnot g00102(.din(n294), .dout(n295));
  jxor g00103(.dina(n295), .dinb(n285), .dout(n296));
  jxor g00104(.dina(n296), .dinb(n280), .dout(n297));
  jand g00105(.dina(n272), .dinb(n264), .dout(n298));
  jor  g00106(.dina(n272), .dinb(n264), .dout(n299));
  jand g00107(.dina(n277), .dinb(n299), .dout(n300));
  jor  g00108(.dina(n300), .dinb(n298), .dout(n301));
  jxor g00109(.dina(n301), .dinb(n297), .dout(\asquared[9] ));
  jand g00110(.dina(n284), .dinb(n282), .dout(n303));
  jand g00111(.dina(n295), .dinb(n285), .dout(n304));
  jor  g00112(.dina(n304), .dinb(n303), .dout(n305));
  jand g00113(.dina(n283), .dinb(n268), .dout(n306));
  jand g00114(.dina(\a[9] ), .dinb(\a[0] ), .dout(n307));
  jxor g00115(.dina(n307), .dinb(n306), .dout(n308));
  jand g00116(.dina(\a[8] ), .dinb(\a[5] ), .dout(n309));
  jand g00117(.dina(n309), .dinb(\a[1] ), .dout(n310));
  jnot g00118(.din(n310), .dout(n311));
  jand g00119(.dina(n311), .dinb(\a[5] ), .dout(n312));
  jand g00120(.dina(\a[8] ), .dinb(\a[1] ), .dout(n313));
  jand g00121(.dina(n313), .dinb(n218), .dout(n314));
  jor  g00122(.dina(n314), .dinb(n312), .dout(n315));
  jxor g00123(.dina(n315), .dinb(n308), .dout(n316));
  jand g00124(.dina(n289), .dinb(n286), .dout(n317));
  jor  g00125(.dina(n317), .dinb(n292), .dout(n318));
  jand g00126(.dina(\a[7] ), .dinb(\a[2] ), .dout(n319));
  jand g00127(.dina(\a[5] ), .dinb(\a[4] ), .dout(n320));
  jand g00128(.dina(\a[6] ), .dinb(\a[3] ), .dout(n321));
  jor  g00129(.dina(n321), .dinb(n320), .dout(n322));
  jand g00130(.dina(\a[6] ), .dinb(\a[4] ), .dout(n323));
  jand g00131(.dina(n323), .dinb(n268), .dout(n324));
  jnot g00132(.din(n324), .dout(n325));
  jand g00133(.dina(n325), .dinb(n322), .dout(n326));
  jxor g00134(.dina(n326), .dinb(n319), .dout(n327));
  jxor g00135(.dina(n327), .dinb(n318), .dout(n328));
  jxor g00136(.dina(n328), .dinb(n316), .dout(n329));
  jxor g00137(.dina(n329), .dinb(n305), .dout(n330));
  jand g00138(.dina(n296), .dinb(n280), .dout(n331));
  jor  g00139(.dina(n296), .dinb(n280), .dout(n332));
  jand g00140(.dina(n301), .dinb(n332), .dout(n333));
  jor  g00141(.dina(n333), .dinb(n331), .dout(n334));
  jxor g00142(.dina(n334), .dinb(n330), .dout(\asquared[10] ));
  jand g00143(.dina(n327), .dinb(n318), .dout(n336));
  jand g00144(.dina(n328), .dinb(n316), .dout(n337));
  jor  g00145(.dina(n337), .dinb(n336), .dout(n338));
  jand g00146(.dina(n326), .dinb(n319), .dout(n339));
  jor  g00147(.dina(n339), .dinb(n324), .dout(n340));
  jand g00148(.dina(\a[9] ), .dinb(\a[1] ), .dout(n341));
  jor  g00149(.dina(n341), .dinb(n323), .dout(n342));
  jand g00150(.dina(\a[9] ), .dinb(\a[4] ), .dout(n343));
  jand g00151(.dina(n343), .dinb(n256), .dout(n344));
  jnot g00152(.din(n344), .dout(n345));
  jand g00153(.dina(n345), .dinb(n342), .dout(n346));
  jxor g00154(.dina(n346), .dinb(n310), .dout(n347));
  jxor g00155(.dina(n347), .dinb(n340), .dout(n348));
  jnot g00156(.din(n291), .dout(n349));
  jand g00157(.dina(\a[7] ), .dinb(\a[3] ), .dout(n350));
  jand g00158(.dina(\a[10] ), .dinb(\a[0] ), .dout(n351));
  jxor g00159(.dina(n351), .dinb(n350), .dout(n352));
  jxor g00160(.dina(n352), .dinb(n349), .dout(n353));
  jnot g00161(.din(n353), .dout(n354));
  jand g00162(.dina(n307), .dinb(n306), .dout(n355));
  jand g00163(.dina(n315), .dinb(n308), .dout(n356));
  jor  g00164(.dina(n356), .dinb(n355), .dout(n357));
  jxor g00165(.dina(n357), .dinb(n354), .dout(n358));
  jxor g00166(.dina(n358), .dinb(n348), .dout(n359));
  jxor g00167(.dina(n359), .dinb(n338), .dout(n360));
  jand g00168(.dina(n329), .dinb(n305), .dout(n361));
  jor  g00169(.dina(n329), .dinb(n305), .dout(n362));
  jand g00170(.dina(n334), .dinb(n362), .dout(n363));
  jor  g00171(.dina(n363), .dinb(n361), .dout(n364));
  jxor g00172(.dina(n364), .dinb(n360), .dout(\asquared[11] ));
  jand g00173(.dina(n357), .dinb(n354), .dout(n366));
  jand g00174(.dina(n358), .dinb(n348), .dout(n367));
  jor  g00175(.dina(n367), .dinb(n366), .dout(n368));
  jand g00176(.dina(\a[9] ), .dinb(\a[2] ), .dout(n369));
  jand g00177(.dina(\a[8] ), .dinb(\a[3] ), .dout(n370));
  jor  g00178(.dina(n370), .dinb(n369), .dout(n371));
  jand g00179(.dina(\a[9] ), .dinb(\a[3] ), .dout(n372));
  jand g00180(.dina(n372), .dinb(n291), .dout(n373));
  jnot g00181(.din(n373), .dout(n374));
  jand g00182(.dina(n374), .dinb(n371), .dout(n375));
  jxor g00183(.dina(n375), .dinb(n345), .dout(n376));
  jnot g00184(.din(n376), .dout(n377));
  jand g00185(.dina(n256), .dinb(\a[10] ), .dout(n378));
  jnot g00186(.din(n378), .dout(n379));
  jand g00187(.dina(n379), .dinb(\a[6] ), .dout(n380));
  jand g00188(.dina(\a[10] ), .dinb(\a[1] ), .dout(n381));
  jand g00189(.dina(n381), .dinb(n260), .dout(n382));
  jor  g00190(.dina(n382), .dinb(n380), .dout(n383));
  jand g00191(.dina(n351), .dinb(n350), .dout(n384));
  jnot g00192(.din(n384), .dout(n385));
  jnot g00193(.din(n350), .dout(n386));
  jnot g00194(.din(n351), .dout(n387));
  jand g00195(.dina(n387), .dinb(n386), .dout(n388));
  jor  g00196(.dina(n388), .dinb(n349), .dout(n389));
  jand g00197(.dina(n389), .dinb(n385), .dout(n390));
  jnot g00198(.din(n390), .dout(n391));
  jxor g00199(.dina(n391), .dinb(n383), .dout(n392));
  jxor g00200(.dina(n392), .dinb(n377), .dout(n393));
  jand g00201(.dina(n346), .dinb(n310), .dout(n394));
  jand g00202(.dina(n347), .dinb(n340), .dout(n395));
  jor  g00203(.dina(n395), .dinb(n394), .dout(n396));
  jand g00204(.dina(\a[11] ), .dinb(\a[0] ), .dout(n397));
  jand g00205(.dina(\a[6] ), .dinb(\a[5] ), .dout(n398));
  jand g00206(.dina(\a[7] ), .dinb(\a[4] ), .dout(n399));
  jor  g00207(.dina(n399), .dinb(n398), .dout(n400));
  jand g00208(.dina(\a[7] ), .dinb(\a[5] ), .dout(n401));
  jand g00209(.dina(n401), .dinb(n323), .dout(n402));
  jnot g00210(.din(n402), .dout(n403));
  jand g00211(.dina(n403), .dinb(n400), .dout(n404));
  jxor g00212(.dina(n404), .dinb(n397), .dout(n405));
  jxor g00213(.dina(n405), .dinb(n396), .dout(n406));
  jxor g00214(.dina(n406), .dinb(n393), .dout(n407));
  jxor g00215(.dina(n407), .dinb(n368), .dout(n408));
  jand g00216(.dina(n359), .dinb(n338), .dout(n409));
  jnot g00217(.din(n338), .dout(n410));
  jnot g00218(.din(n359), .dout(n411));
  jand g00219(.dina(n411), .dinb(n410), .dout(n412));
  jnot g00220(.din(n412), .dout(n413));
  jand g00221(.dina(n364), .dinb(n413), .dout(n414));
  jor  g00222(.dina(n414), .dinb(n409), .dout(n415));
  jxor g00223(.dina(n415), .dinb(n408), .dout(\asquared[12] ));
  jand g00224(.dina(n405), .dinb(n396), .dout(n417));
  jand g00225(.dina(n406), .dinb(n393), .dout(n418));
  jor  g00226(.dina(n418), .dinb(n417), .dout(n419));
  jand g00227(.dina(n391), .dinb(n383), .dout(n420));
  jand g00228(.dina(n392), .dinb(n377), .dout(n421));
  jor  g00229(.dina(n421), .dinb(n420), .dout(n422));
  jand g00230(.dina(\a[11] ), .dinb(\a[1] ), .dout(n423));
  jor  g00231(.dina(n423), .dinb(n401), .dout(n424));
  jand g00232(.dina(\a[11] ), .dinb(\a[5] ), .dout(n425));
  jand g00233(.dina(n425), .dinb(n283), .dout(n426));
  jnot g00234(.din(n426), .dout(n427));
  jand g00235(.dina(n427), .dinb(n424), .dout(n428));
  jand g00236(.dina(\a[8] ), .dinb(\a[4] ), .dout(n429));
  jnot g00237(.din(n429), .dout(n430));
  jxor g00238(.dina(n430), .dinb(n378), .dout(n431));
  jxor g00239(.dina(n431), .dinb(n428), .dout(n432));
  jnot g00240(.din(n432), .dout(n433));
  jxor g00241(.dina(n433), .dinb(n422), .dout(n434));
  jand g00242(.dina(n404), .dinb(n397), .dout(n435));
  jor  g00243(.dina(n435), .dinb(n402), .dout(n436));
  jand g00244(.dina(n371), .dinb(n344), .dout(n437));
  jor  g00245(.dina(n437), .dinb(n373), .dout(n438));
  jxor g00246(.dina(n438), .dinb(n436), .dout(n439));
  jnot g00247(.din(n372), .dout(n440));
  jand g00248(.dina(\a[10] ), .dinb(\a[2] ), .dout(n441));
  jand g00249(.dina(\a[12] ), .dinb(\a[0] ), .dout(n442));
  jor  g00250(.dina(n442), .dinb(n441), .dout(n443));
  jand g00251(.dina(\a[12] ), .dinb(\a[2] ), .dout(n444));
  jand g00252(.dina(n444), .dinb(n351), .dout(n445));
  jnot g00253(.din(n445), .dout(n446));
  jand g00254(.dina(n446), .dinb(n443), .dout(n447));
  jxor g00255(.dina(n447), .dinb(n440), .dout(n448));
  jnot g00256(.din(n448), .dout(n449));
  jxor g00257(.dina(n449), .dinb(n439), .dout(n450));
  jxor g00258(.dina(n450), .dinb(n434), .dout(n451));
  jxor g00259(.dina(n451), .dinb(n419), .dout(n452));
  jand g00260(.dina(n407), .dinb(n368), .dout(n453));
  jnot g00261(.din(n368), .dout(n454));
  jnot g00262(.din(n407), .dout(n455));
  jand g00263(.dina(n455), .dinb(n454), .dout(n456));
  jnot g00264(.din(n456), .dout(n457));
  jand g00265(.dina(n415), .dinb(n457), .dout(n458));
  jor  g00266(.dina(n458), .dinb(n453), .dout(n459));
  jxor g00267(.dina(n459), .dinb(n452), .dout(\asquared[13] ));
  jand g00268(.dina(\a[11] ), .dinb(\a[2] ), .dout(n461));
  jand g00269(.dina(\a[7] ), .dinb(\a[6] ), .dout(n462));
  jor  g00270(.dina(n462), .dinb(n309), .dout(n463));
  jnot g00271(.din(n463), .dout(n464));
  jand g00272(.dina(\a[8] ), .dinb(\a[6] ), .dout(n465));
  jand g00273(.dina(n465), .dinb(n401), .dout(n466));
  jor  g00274(.dina(n466), .dinb(n464), .dout(n467));
  jxor g00275(.dina(n467), .dinb(n461), .dout(n468));
  jnot g00276(.din(n468), .dout(n469));
  jand g00277(.dina(\a[10] ), .dinb(\a[3] ), .dout(n470));
  jand g00278(.dina(\a[13] ), .dinb(\a[0] ), .dout(n471));
  jor  g00279(.dina(n471), .dinb(n343), .dout(n472));
  jnot g00280(.din(n472), .dout(n473));
  jand g00281(.dina(\a[13] ), .dinb(\a[4] ), .dout(n474));
  jand g00282(.dina(n474), .dinb(n307), .dout(n475));
  jor  g00283(.dina(n475), .dinb(n473), .dout(n476));
  jxor g00284(.dina(n476), .dinb(n470), .dout(n477));
  jnot g00285(.din(n477), .dout(n478));
  jand g00286(.dina(n430), .dinb(n379), .dout(n479));
  jnot g00287(.din(n479), .dout(n480));
  jand g00288(.dina(n429), .dinb(n378), .dout(n481));
  jor  g00289(.dina(n481), .dinb(n428), .dout(n482));
  jand g00290(.dina(n482), .dinb(n480), .dout(n483));
  jxor g00291(.dina(n483), .dinb(n478), .dout(n484));
  jxor g00292(.dina(n484), .dinb(n469), .dout(n485));
  jnot g00293(.din(\a[12] ), .dout(n486));
  jand g00294(.dina(n426), .dinb(n486), .dout(n487));
  jnot g00295(.din(n487), .dout(n488));
  jand g00296(.dina(n283), .dinb(\a[12] ), .dout(n489));
  jnot g00297(.din(n489), .dout(n490));
  jand g00298(.dina(\a[12] ), .dinb(\a[1] ), .dout(n491));
  jor  g00299(.dina(n491), .dinb(\a[7] ), .dout(n492));
  jand g00300(.dina(n492), .dinb(n490), .dout(n493));
  jor  g00301(.dina(n493), .dinb(n426), .dout(n494));
  jand g00302(.dina(n494), .dinb(n488), .dout(n495));
  jand g00303(.dina(n443), .dinb(n372), .dout(n496));
  jor  g00304(.dina(n496), .dinb(n445), .dout(n497));
  jxor g00305(.dina(n497), .dinb(n495), .dout(n498));
  jnot g00306(.din(n498), .dout(n499));
  jand g00307(.dina(n438), .dinb(n436), .dout(n500));
  jnot g00308(.din(n500), .dout(n501));
  jnot g00309(.din(n436), .dout(n502));
  jnot g00310(.din(n438), .dout(n503));
  jand g00311(.dina(n503), .dinb(n502), .dout(n504));
  jor  g00312(.dina(n448), .dinb(n504), .dout(n505));
  jand g00313(.dina(n505), .dinb(n501), .dout(n506));
  jxor g00314(.dina(n506), .dinb(n499), .dout(n507));
  jand g00315(.dina(n433), .dinb(n422), .dout(n508));
  jand g00316(.dina(n450), .dinb(n434), .dout(n509));
  jor  g00317(.dina(n509), .dinb(n508), .dout(n510));
  jxor g00318(.dina(n510), .dinb(n507), .dout(n511));
  jxor g00319(.dina(n511), .dinb(n485), .dout(n512));
  jand g00320(.dina(n451), .dinb(n419), .dout(n513));
  jnot g00321(.din(n419), .dout(n514));
  jnot g00322(.din(n451), .dout(n515));
  jand g00323(.dina(n515), .dinb(n514), .dout(n516));
  jnot g00324(.din(n516), .dout(n517));
  jand g00325(.dina(n459), .dinb(n517), .dout(n518));
  jor  g00326(.dina(n518), .dinb(n513), .dout(n519));
  jxor g00327(.dina(n519), .dinb(n512), .dout(\asquared[14] ));
  jor  g00328(.dina(n506), .dinb(n499), .dout(n521));
  jand g00329(.dina(n510), .dinb(n507), .dout(n522));
  jnot g00330(.din(n522), .dout(n523));
  jand g00331(.dina(n523), .dinb(n521), .dout(n524));
  jnot g00332(.din(n524), .dout(n525));
  jand g00333(.dina(n483), .dinb(n478), .dout(n526));
  jand g00334(.dina(n484), .dinb(n469), .dout(n527));
  jor  g00335(.dina(n527), .dinb(n526), .dout(n528));
  jand g00336(.dina(\a[13] ), .dinb(\a[1] ), .dout(n529));
  jxor g00337(.dina(n529), .dinb(n465), .dout(n530));
  jand g00338(.dina(n463), .dinb(n461), .dout(n531));
  jor  g00339(.dina(n531), .dinb(n466), .dout(n532));
  jxor g00340(.dina(n532), .dinb(n530), .dout(n533));
  jand g00341(.dina(n472), .dinb(n470), .dout(n534));
  jor  g00342(.dina(n534), .dinb(n475), .dout(n535));
  jxor g00343(.dina(n535), .dinb(n533), .dout(n536));
  jxor g00344(.dina(n536), .dinb(n528), .dout(n537));
  jand g00345(.dina(n497), .dinb(n495), .dout(n538));
  jor  g00346(.dina(n538), .dinb(n487), .dout(n539));
  jand g00347(.dina(\a[10] ), .dinb(\a[4] ), .dout(n540));
  jand g00348(.dina(\a[9] ), .dinb(\a[5] ), .dout(n541));
  jor  g00349(.dina(n541), .dinb(n540), .dout(n542));
  jand g00350(.dina(\a[10] ), .dinb(\a[5] ), .dout(n543));
  jand g00351(.dina(n543), .dinb(n343), .dout(n544));
  jnot g00352(.din(n544), .dout(n545));
  jand g00353(.dina(n545), .dinb(n542), .dout(n546));
  jxor g00354(.dina(n546), .dinb(n490), .dout(n547));
  jnot g00355(.din(n547), .dout(n548));
  jand g00356(.dina(\a[14] ), .dinb(\a[0] ), .dout(n549));
  jand g00357(.dina(\a[11] ), .dinb(\a[3] ), .dout(n550));
  jor  g00358(.dina(n550), .dinb(n444), .dout(n551));
  jand g00359(.dina(\a[12] ), .dinb(\a[3] ), .dout(n552));
  jand g00360(.dina(n552), .dinb(n461), .dout(n553));
  jnot g00361(.din(n553), .dout(n554));
  jand g00362(.dina(n554), .dinb(n551), .dout(n555));
  jxor g00363(.dina(n555), .dinb(n549), .dout(n556));
  jxor g00364(.dina(n556), .dinb(n548), .dout(n557));
  jxor g00365(.dina(n557), .dinb(n539), .dout(n558));
  jxor g00366(.dina(n558), .dinb(n537), .dout(n559));
  jxor g00367(.dina(n559), .dinb(n525), .dout(n560));
  jand g00368(.dina(n511), .dinb(n485), .dout(n561));
  jnot g00369(.din(n485), .dout(n562));
  jnot g00370(.din(n511), .dout(n563));
  jand g00371(.dina(n563), .dinb(n562), .dout(n564));
  jnot g00372(.din(n564), .dout(n565));
  jand g00373(.dina(n519), .dinb(n565), .dout(n566));
  jor  g00374(.dina(n566), .dinb(n561), .dout(n567));
  jxor g00375(.dina(n567), .dinb(n560), .dout(\asquared[15] ));
  jand g00376(.dina(n536), .dinb(n528), .dout(n569));
  jand g00377(.dina(n558), .dinb(n537), .dout(n570));
  jor  g00378(.dina(n570), .dinb(n569), .dout(n571));
  jand g00379(.dina(n532), .dinb(n530), .dout(n572));
  jand g00380(.dina(n535), .dinb(n533), .dout(n573));
  jor  g00381(.dina(n573), .dinb(n572), .dout(n574));
  jand g00382(.dina(\a[13] ), .dinb(\a[2] ), .dout(n575));
  jand g00383(.dina(\a[8] ), .dinb(\a[7] ), .dout(n576));
  jnot g00384(.din(n576), .dout(n577));
  jand g00385(.dina(\a[9] ), .dinb(\a[6] ), .dout(n578));
  jxor g00386(.dina(n578), .dinb(n577), .dout(n579));
  jxor g00387(.dina(n579), .dinb(n575), .dout(n580));
  jnot g00388(.din(n580), .dout(n581));
  jand g00389(.dina(\a[14] ), .dinb(\a[1] ), .dout(n582));
  jxor g00390(.dina(n582), .dinb(\a[8] ), .dout(n583));
  jand g00391(.dina(n529), .dinb(n465), .dout(n584));
  jand g00392(.dina(\a[11] ), .dinb(\a[4] ), .dout(n585));
  jxor g00393(.dina(n585), .dinb(n584), .dout(n586));
  jxor g00394(.dina(n586), .dinb(n583), .dout(n587));
  jxor g00395(.dina(n587), .dinb(n581), .dout(n588));
  jxor g00396(.dina(n588), .dinb(n574), .dout(n589));
  jand g00397(.dina(n556), .dinb(n548), .dout(n590));
  jand g00398(.dina(n557), .dinb(n539), .dout(n591));
  jor  g00399(.dina(n591), .dinb(n590), .dout(n592));
  jnot g00400(.din(n592), .dout(n593));
  jand g00401(.dina(n555), .dinb(n549), .dout(n594));
  jor  g00402(.dina(n594), .dinb(n553), .dout(n595));
  jand g00403(.dina(n542), .dinb(n489), .dout(n596));
  jor  g00404(.dina(n596), .dinb(n544), .dout(n597));
  jxor g00405(.dina(n597), .dinb(n595), .dout(n598));
  jand g00406(.dina(\a[15] ), .dinb(\a[10] ), .dout(n599));
  jand g00407(.dina(n599), .dinb(\a[0] ), .dout(n600));
  jand g00408(.dina(n552), .dinb(\a[10] ), .dout(n601));
  jor  g00409(.dina(n601), .dinb(n600), .dout(n602));
  jand g00410(.dina(n602), .dinb(\a[5] ), .dout(n603));
  jand g00411(.dina(\a[15] ), .dinb(\a[0] ), .dout(n604));
  jand g00412(.dina(n604), .dinb(n552), .dout(n605));
  jnot g00413(.din(n605), .dout(n606));
  jand g00414(.dina(n606), .dinb(n603), .dout(n607));
  jnot g00415(.din(n607), .dout(n608));
  jxor g00416(.dina(n604), .dinb(n552), .dout(n609));
  jor  g00417(.dina(n609), .dinb(n543), .dout(n610));
  jand g00418(.dina(n610), .dinb(n608), .dout(n611));
  jnot g00419(.din(n611), .dout(n612));
  jxor g00420(.dina(n612), .dinb(n598), .dout(n613));
  jxor g00421(.dina(n613), .dinb(n593), .dout(n614));
  jxor g00422(.dina(n614), .dinb(n589), .dout(n615));
  jxor g00423(.dina(n615), .dinb(n571), .dout(n616));
  jand g00424(.dina(n559), .dinb(n525), .dout(n617));
  jor  g00425(.dina(n559), .dinb(n525), .dout(n618));
  jand g00426(.dina(n567), .dinb(n618), .dout(n619));
  jor  g00427(.dina(n619), .dinb(n617), .dout(n620));
  jxor g00428(.dina(n620), .dinb(n616), .dout(\asquared[16] ));
  jor  g00429(.dina(n613), .dinb(n593), .dout(n622));
  jand g00430(.dina(n614), .dinb(n589), .dout(n623));
  jnot g00431(.din(n623), .dout(n624));
  jand g00432(.dina(n624), .dinb(n622), .dout(n625));
  jnot g00433(.din(n625), .dout(n626));
  jand g00434(.dina(n587), .dinb(n581), .dout(n627));
  jand g00435(.dina(n588), .dinb(n574), .dout(n628));
  jor  g00436(.dina(n628), .dinb(n627), .dout(n629));
  jand g00437(.dina(n585), .dinb(n584), .dout(n630));
  jand g00438(.dina(n586), .dinb(n583), .dout(n631));
  jor  g00439(.dina(n631), .dinb(n630), .dout(n632));
  jor  g00440(.dina(n605), .dinb(n603), .dout(n633));
  jxor g00441(.dina(n633), .dinb(n632), .dout(n634));
  jnot g00442(.din(n425), .dout(n635));
  jand g00443(.dina(\a[10] ), .dinb(\a[6] ), .dout(n636));
  jand g00444(.dina(\a[16] ), .dinb(\a[0] ), .dout(n637));
  jor  g00445(.dina(n637), .dinb(n636), .dout(n638));
  jand g00446(.dina(\a[16] ), .dinb(\a[6] ), .dout(n639));
  jand g00447(.dina(n639), .dinb(n351), .dout(n640));
  jnot g00448(.din(n640), .dout(n641));
  jand g00449(.dina(n641), .dinb(n638), .dout(n642));
  jxor g00450(.dina(n642), .dinb(n635), .dout(n643));
  jnot g00451(.din(n643), .dout(n644));
  jxor g00452(.dina(n644), .dinb(n634), .dout(n645));
  jxor g00453(.dina(n645), .dinb(n629), .dout(n646));
  jand g00454(.dina(n582), .dinb(\a[8] ), .dout(n647));
  jand g00455(.dina(\a[9] ), .dinb(\a[7] ), .dout(n648));
  jand g00456(.dina(\a[15] ), .dinb(\a[1] ), .dout(n649));
  jxor g00457(.dina(n649), .dinb(n648), .dout(n650));
  jxor g00458(.dina(n650), .dinb(n647), .dout(n651));
  jnot g00459(.din(n578), .dout(n652));
  jand g00460(.dina(n652), .dinb(n577), .dout(n653));
  jnot g00461(.din(n653), .dout(n654));
  jand g00462(.dina(n578), .dinb(n576), .dout(n655));
  jor  g00463(.dina(n655), .dinb(n575), .dout(n656));
  jand g00464(.dina(n656), .dinb(n654), .dout(n657));
  jxor g00465(.dina(n657), .dinb(n651), .dout(n658));
  jand g00466(.dina(\a[12] ), .dinb(\a[4] ), .dout(n659));
  jand g00467(.dina(\a[13] ), .dinb(\a[3] ), .dout(n660));
  jand g00468(.dina(\a[14] ), .dinb(\a[2] ), .dout(n661));
  jor  g00469(.dina(n661), .dinb(n660), .dout(n662));
  jnot g00470(.din(n662), .dout(n663));
  jand g00471(.dina(\a[14] ), .dinb(\a[3] ), .dout(n664));
  jand g00472(.dina(n664), .dinb(n575), .dout(n665));
  jor  g00473(.dina(n665), .dinb(n663), .dout(n666));
  jxor g00474(.dina(n666), .dinb(n659), .dout(n667));
  jand g00475(.dina(n597), .dinb(n595), .dout(n668));
  jnot g00476(.din(n668), .dout(n669));
  jnot g00477(.din(n595), .dout(n670));
  jnot g00478(.din(n597), .dout(n671));
  jand g00479(.dina(n671), .dinb(n670), .dout(n672));
  jor  g00480(.dina(n612), .dinb(n672), .dout(n673));
  jand g00481(.dina(n673), .dinb(n669), .dout(n674));
  jxor g00482(.dina(n674), .dinb(n667), .dout(n675));
  jxor g00483(.dina(n675), .dinb(n658), .dout(n676));
  jxor g00484(.dina(n676), .dinb(n646), .dout(n677));
  jxor g00485(.dina(n677), .dinb(n626), .dout(n678));
  jand g00486(.dina(n615), .dinb(n571), .dout(n679));
  jor  g00487(.dina(n615), .dinb(n571), .dout(n680));
  jand g00488(.dina(n620), .dinb(n680), .dout(n681));
  jor  g00489(.dina(n681), .dinb(n679), .dout(n682));
  jxor g00490(.dina(n682), .dinb(n678), .dout(\asquared[17] ));
  jand g00491(.dina(n645), .dinb(n629), .dout(n684));
  jand g00492(.dina(n676), .dinb(n646), .dout(n685));
  jor  g00493(.dina(n685), .dinb(n684), .dout(n686));
  jor  g00494(.dina(n674), .dinb(n667), .dout(n687));
  jand g00495(.dina(n675), .dinb(n658), .dout(n688));
  jnot g00496(.din(n688), .dout(n689));
  jand g00497(.dina(n689), .dinb(n687), .dout(n690));
  jnot g00498(.din(n690), .dout(n691));
  jand g00499(.dina(\a[9] ), .dinb(\a[8] ), .dout(n692));
  jand g00500(.dina(\a[10] ), .dinb(\a[7] ), .dout(n693));
  jor  g00501(.dina(n693), .dinb(n692), .dout(n694));
  jnot g00502(.din(n694), .dout(n695));
  jand g00503(.dina(\a[10] ), .dinb(\a[8] ), .dout(n696));
  jand g00504(.dina(n696), .dinb(n648), .dout(n697));
  jor  g00505(.dina(n697), .dinb(n695), .dout(n698));
  jxor g00506(.dina(n698), .dinb(n664), .dout(n699));
  jand g00507(.dina(n649), .dinb(n648), .dout(n700));
  jand g00508(.dina(\a[12] ), .dinb(\a[5] ), .dout(n701));
  jand g00509(.dina(\a[17] ), .dinb(\a[0] ), .dout(n702));
  jnot g00510(.din(n702), .dout(n703));
  jxor g00511(.dina(n703), .dinb(n701), .dout(n704));
  jxor g00512(.dina(n704), .dinb(n700), .dout(n705));
  jxor g00513(.dina(n705), .dinb(n699), .dout(n706));
  jand g00514(.dina(\a[15] ), .dinb(\a[11] ), .dout(n707));
  jand g00515(.dina(n707), .dinb(\a[2] ), .dout(n708));
  jand g00516(.dina(n474), .dinb(\a[11] ), .dout(n709));
  jor  g00517(.dina(n709), .dinb(n708), .dout(n710));
  jand g00518(.dina(n710), .dinb(\a[6] ), .dout(n711));
  jand g00519(.dina(\a[15] ), .dinb(\a[4] ), .dout(n712));
  jand g00520(.dina(n712), .dinb(n575), .dout(n713));
  jnot g00521(.din(n713), .dout(n714));
  jand g00522(.dina(n714), .dinb(n711), .dout(n715));
  jnot g00523(.din(n715), .dout(n716));
  jand g00524(.dina(\a[11] ), .dinb(\a[6] ), .dout(n717));
  jand g00525(.dina(\a[15] ), .dinb(\a[2] ), .dout(n718));
  jor  g00526(.dina(n718), .dinb(n474), .dout(n719));
  jand g00527(.dina(n719), .dinb(n714), .dout(n720));
  jor  g00528(.dina(n720), .dinb(n717), .dout(n721));
  jand g00529(.dina(n721), .dinb(n716), .dout(n722));
  jxor g00530(.dina(n722), .dinb(n706), .dout(n723));
  jxor g00531(.dina(n723), .dinb(n691), .dout(n724));
  jand g00532(.dina(n650), .dinb(n647), .dout(n725));
  jand g00533(.dina(n657), .dinb(n651), .dout(n726));
  jor  g00534(.dina(n726), .dinb(n725), .dout(n727));
  jand g00535(.dina(n633), .dinb(n632), .dout(n728));
  jnot g00536(.din(n728), .dout(n729));
  jnot g00537(.din(n632), .dout(n730));
  jnot g00538(.din(n633), .dout(n731));
  jand g00539(.dina(n731), .dinb(n730), .dout(n732));
  jor  g00540(.dina(n643), .dinb(n732), .dout(n733));
  jand g00541(.dina(n733), .dinb(n729), .dout(n734));
  jnot g00542(.din(n734), .dout(n735));
  jxor g00543(.dina(n735), .dinb(n727), .dout(n736));
  jand g00544(.dina(\a[16] ), .dinb(\a[1] ), .dout(n737));
  jor  g00545(.dina(n737), .dinb(\a[9] ), .dout(n738));
  jand g00546(.dina(\a[16] ), .dinb(\a[9] ), .dout(n739));
  jand g00547(.dina(n739), .dinb(\a[1] ), .dout(n740));
  jnot g00548(.din(n740), .dout(n741));
  jand g00549(.dina(n741), .dinb(n738), .dout(n742));
  jand g00550(.dina(n662), .dinb(n659), .dout(n743));
  jor  g00551(.dina(n743), .dinb(n665), .dout(n744));
  jxor g00552(.dina(n744), .dinb(n742), .dout(n745));
  jand g00553(.dina(n638), .dinb(n425), .dout(n746));
  jor  g00554(.dina(n746), .dinb(n640), .dout(n747));
  jxor g00555(.dina(n747), .dinb(n745), .dout(n748));
  jxor g00556(.dina(n748), .dinb(n736), .dout(n749));
  jxor g00557(.dina(n749), .dinb(n724), .dout(n750));
  jxor g00558(.dina(n750), .dinb(n686), .dout(n751));
  jand g00559(.dina(n677), .dinb(n626), .dout(n752));
  jor  g00560(.dina(n677), .dinb(n626), .dout(n753));
  jand g00561(.dina(n682), .dinb(n753), .dout(n754));
  jor  g00562(.dina(n754), .dinb(n752), .dout(n755));
  jxor g00563(.dina(n755), .dinb(n751), .dout(\asquared[18] ));
  jand g00564(.dina(n723), .dinb(n691), .dout(n757));
  jand g00565(.dina(n749), .dinb(n724), .dout(n758));
  jor  g00566(.dina(n758), .dinb(n757), .dout(n759));
  jand g00567(.dina(n694), .dinb(n664), .dout(n760));
  jor  g00568(.dina(n760), .dinb(n697), .dout(n761));
  jor  g00569(.dina(n713), .dinb(n711), .dout(n762));
  jxor g00570(.dina(n762), .dinb(n761), .dout(n763));
  jnot g00571(.din(n701), .dout(n764));
  jand g00572(.dina(n703), .dinb(n764), .dout(n765));
  jnot g00573(.din(n765), .dout(n766));
  jand g00574(.dina(n702), .dinb(n701), .dout(n767));
  jor  g00575(.dina(n767), .dinb(n700), .dout(n768));
  jand g00576(.dina(n768), .dinb(n766), .dout(n769));
  jxor g00577(.dina(n769), .dinb(n763), .dout(n770));
  jand g00578(.dina(n744), .dinb(n742), .dout(n771));
  jand g00579(.dina(n747), .dinb(n745), .dout(n772));
  jor  g00580(.dina(n772), .dinb(n771), .dout(n773));
  jnot g00581(.din(n773), .dout(n774));
  jor  g00582(.dina(n705), .dinb(n699), .dout(n775));
  jand g00583(.dina(n722), .dinb(n706), .dout(n776));
  jnot g00584(.din(n776), .dout(n777));
  jand g00585(.dina(n777), .dinb(n775), .dout(n778));
  jxor g00586(.dina(n778), .dinb(n774), .dout(n779));
  jxor g00587(.dina(n779), .dinb(n770), .dout(n780));
  jand g00588(.dina(n735), .dinb(n727), .dout(n781));
  jand g00589(.dina(n748), .dinb(n736), .dout(n782));
  jor  g00590(.dina(n782), .dinb(n781), .dout(n783));
  jand g00591(.dina(\a[12] ), .dinb(\a[6] ), .dout(n784));
  jxor g00592(.dina(n784), .dinb(n740), .dout(n785));
  jand g00593(.dina(\a[17] ), .dinb(\a[1] ), .dout(n786));
  jxor g00594(.dina(n786), .dinb(n696), .dout(n787));
  jxor g00595(.dina(n787), .dinb(n785), .dout(n788));
  jand g00596(.dina(\a[11] ), .dinb(\a[7] ), .dout(n789));
  jnot g00597(.din(n789), .dout(n790));
  jand g00598(.dina(\a[18] ), .dinb(\a[0] ), .dout(n791));
  jand g00599(.dina(\a[13] ), .dinb(\a[5] ), .dout(n792));
  jxor g00600(.dina(n792), .dinb(n791), .dout(n793));
  jxor g00601(.dina(n793), .dinb(n790), .dout(n794));
  jand g00602(.dina(\a[14] ), .dinb(\a[4] ), .dout(n795));
  jnot g00603(.din(n795), .dout(n796));
  jand g00604(.dina(\a[15] ), .dinb(\a[3] ), .dout(n797));
  jand g00605(.dina(\a[16] ), .dinb(\a[2] ), .dout(n798));
  jor  g00606(.dina(n798), .dinb(n797), .dout(n799));
  jand g00607(.dina(\a[16] ), .dinb(\a[3] ), .dout(n800));
  jand g00608(.dina(n800), .dinb(n718), .dout(n801));
  jnot g00609(.din(n801), .dout(n802));
  jand g00610(.dina(n802), .dinb(n799), .dout(n803));
  jxor g00611(.dina(n803), .dinb(n796), .dout(n804));
  jxor g00612(.dina(n804), .dinb(n794), .dout(n805));
  jxor g00613(.dina(n805), .dinb(n788), .dout(n806));
  jxor g00614(.dina(n806), .dinb(n783), .dout(n807));
  jxor g00615(.dina(n807), .dinb(n780), .dout(n808));
  jxor g00616(.dina(n808), .dinb(n759), .dout(n809));
  jand g00617(.dina(n750), .dinb(n686), .dout(n810));
  jor  g00618(.dina(n750), .dinb(n686), .dout(n811));
  jand g00619(.dina(n755), .dinb(n811), .dout(n812));
  jor  g00620(.dina(n812), .dinb(n810), .dout(n813));
  jxor g00621(.dina(n813), .dinb(n809), .dout(\asquared[19] ));
  jor  g00622(.dina(n804), .dinb(n794), .dout(n815));
  jand g00623(.dina(n805), .dinb(n788), .dout(n816));
  jnot g00624(.din(n816), .dout(n817));
  jand g00625(.dina(n817), .dinb(n815), .dout(n818));
  jnot g00626(.din(n818), .dout(n819));
  jand g00627(.dina(n786), .dinb(n696), .dout(n820));
  jand g00628(.dina(\a[18] ), .dinb(\a[1] ), .dout(n821));
  jxor g00629(.dina(n821), .dinb(\a[10] ), .dout(n822));
  jor  g00630(.dina(n822), .dinb(n820), .dout(n823));
  jnot g00631(.din(\a[18] ), .dout(n824));
  jand g00632(.dina(n820), .dinb(n824), .dout(n825));
  jnot g00633(.din(n825), .dout(n826));
  jand g00634(.dina(n826), .dinb(n823), .dout(n827));
  jand g00635(.dina(n802), .dinb(n796), .dout(n828));
  jnot g00636(.din(n828), .dout(n829));
  jand g00637(.dina(n829), .dinb(n799), .dout(n830));
  jxor g00638(.dina(n830), .dinb(n827), .dout(n831));
  jxor g00639(.dina(n831), .dinb(n819), .dout(n832));
  jand g00640(.dina(n784), .dinb(n740), .dout(n833));
  jand g00641(.dina(n787), .dinb(n785), .dout(n834));
  jor  g00642(.dina(n834), .dinb(n833), .dout(n835));
  jnot g00643(.din(n835), .dout(n836));
  jand g00644(.dina(n792), .dinb(n791), .dout(n837));
  jnot g00645(.din(n837), .dout(n838));
  jnot g00646(.din(n791), .dout(n839));
  jnot g00647(.din(n792), .dout(n840));
  jand g00648(.dina(n840), .dinb(n839), .dout(n841));
  jor  g00649(.dina(n841), .dinb(n790), .dout(n842));
  jand g00650(.dina(n842), .dinb(n838), .dout(n843));
  jxor g00651(.dina(n843), .dinb(n836), .dout(n844));
  jnot g00652(.din(n800), .dout(n845));
  jand g00653(.dina(\a[10] ), .dinb(\a[9] ), .dout(n846));
  jand g00654(.dina(\a[11] ), .dinb(\a[8] ), .dout(n847));
  jxor g00655(.dina(n847), .dinb(n846), .dout(n848));
  jxor g00656(.dina(n848), .dinb(n845), .dout(n849));
  jnot g00657(.din(n849), .dout(n850));
  jxor g00658(.dina(n850), .dinb(n844), .dout(n851));
  jxor g00659(.dina(n851), .dinb(n832), .dout(n852));
  jand g00660(.dina(n762), .dinb(n761), .dout(n853));
  jand g00661(.dina(n769), .dinb(n763), .dout(n854));
  jor  g00662(.dina(n854), .dinb(n853), .dout(n855));
  jand g00663(.dina(\a[14] ), .dinb(\a[5] ), .dout(n856));
  jand g00664(.dina(\a[13] ), .dinb(\a[6] ), .dout(n857));
  jand g00665(.dina(\a[12] ), .dinb(\a[7] ), .dout(n858));
  jor  g00666(.dina(n858), .dinb(n857), .dout(n859));
  jnot g00667(.din(n859), .dout(n860));
  jand g00668(.dina(\a[13] ), .dinb(\a[7] ), .dout(n861));
  jand g00669(.dina(n861), .dinb(n784), .dout(n862));
  jor  g00670(.dina(n862), .dinb(n860), .dout(n863));
  jxor g00671(.dina(n863), .dinb(n856), .dout(n864));
  jnot g00672(.din(n864), .dout(n865));
  jand g00673(.dina(n208), .dinb(\a[15] ), .dout(n866));
  jand g00674(.dina(\a[17] ), .dinb(\a[2] ), .dout(n867));
  jand g00675(.dina(n867), .dinb(\a[0] ), .dout(n868));
  jor  g00676(.dina(n868), .dinb(n866), .dout(n869));
  jand g00677(.dina(n869), .dinb(\a[19] ), .dout(n870));
  jnot g00678(.din(n870), .dout(n871));
  jor  g00679(.dina(n867), .dinb(n712), .dout(n872));
  jand g00680(.dina(\a[17] ), .dinb(\a[4] ), .dout(n873));
  jand g00681(.dina(n873), .dinb(n718), .dout(n874));
  jnot g00682(.din(n874), .dout(n875));
  jand g00683(.dina(n875), .dinb(n872), .dout(n876));
  jand g00684(.dina(n876), .dinb(n871), .dout(n877));
  jnot g00685(.din(n876), .dout(n878));
  jand g00686(.dina(\a[19] ), .dinb(\a[0] ), .dout(n879));
  jand g00687(.dina(n879), .dinb(n878), .dout(n880));
  jor  g00688(.dina(n880), .dinb(n877), .dout(n881));
  jxor g00689(.dina(n881), .dinb(n865), .dout(n882));
  jxor g00690(.dina(n882), .dinb(n855), .dout(n883));
  jnot g00691(.din(n883), .dout(n884));
  jor  g00692(.dina(n778), .dinb(n774), .dout(n885));
  jand g00693(.dina(n779), .dinb(n770), .dout(n886));
  jnot g00694(.din(n886), .dout(n887));
  jand g00695(.dina(n887), .dinb(n885), .dout(n888));
  jxor g00696(.dina(n888), .dinb(n884), .dout(n889));
  jxor g00697(.dina(n889), .dinb(n852), .dout(n890));
  jand g00698(.dina(n806), .dinb(n783), .dout(n891));
  jand g00699(.dina(n807), .dinb(n780), .dout(n892));
  jor  g00700(.dina(n892), .dinb(n891), .dout(n893));
  jxor g00701(.dina(n893), .dinb(n890), .dout(n894));
  jand g00702(.dina(n808), .dinb(n759), .dout(n895));
  jor  g00703(.dina(n808), .dinb(n759), .dout(n896));
  jand g00704(.dina(n813), .dinb(n896), .dout(n897));
  jor  g00705(.dina(n897), .dinb(n895), .dout(n898));
  jxor g00706(.dina(n898), .dinb(n894), .dout(\asquared[20] ));
  jor  g00707(.dina(n888), .dinb(n884), .dout(n900));
  jand g00708(.dina(n889), .dinb(n852), .dout(n901));
  jnot g00709(.din(n901), .dout(n902));
  jand g00710(.dina(n902), .dinb(n900), .dout(n903));
  jnot g00711(.din(n903), .dout(n904));
  jand g00712(.dina(n830), .dinb(n827), .dout(n905));
  jor  g00713(.dina(n905), .dinb(n825), .dout(n906));
  jnot g00714(.din(n906), .dout(n907));
  jand g00715(.dina(\a[18] ), .dinb(\a[2] ), .dout(n908));
  jand g00716(.dina(\a[17] ), .dinb(\a[3] ), .dout(n909));
  jand g00717(.dina(\a[16] ), .dinb(\a[4] ), .dout(n910));
  jor  g00718(.dina(n910), .dinb(n909), .dout(n911));
  jnot g00719(.din(n911), .dout(n912));
  jand g00720(.dina(n873), .dinb(n800), .dout(n913));
  jor  g00721(.dina(n913), .dinb(n912), .dout(n914));
  jxor g00722(.dina(n914), .dinb(n908), .dout(n915));
  jxor g00723(.dina(n915), .dinb(n907), .dout(n916));
  jand g00724(.dina(n843), .dinb(n836), .dout(n917));
  jor  g00725(.dina(n843), .dinb(n836), .dout(n918));
  jand g00726(.dina(n849), .dinb(n918), .dout(n919));
  jor  g00727(.dina(n919), .dinb(n917), .dout(n920));
  jnot g00728(.din(n920), .dout(n921));
  jxor g00729(.dina(n921), .dinb(n916), .dout(n922));
  jand g00730(.dina(n831), .dinb(n819), .dout(n923));
  jand g00731(.dina(n851), .dinb(n832), .dout(n924));
  jor  g00732(.dina(n924), .dinb(n923), .dout(n925));
  jxor g00733(.dina(n925), .dinb(n922), .dout(n926));
  jand g00734(.dina(n881), .dinb(n865), .dout(n927));
  jand g00735(.dina(n882), .dinb(n855), .dout(n928));
  jor  g00736(.dina(n928), .dinb(n927), .dout(n929));
  jand g00737(.dina(n875), .dinb(n871), .dout(n930));
  jnot g00738(.din(n930), .dout(n931));
  jand g00739(.dina(\a[11] ), .dinb(\a[9] ), .dout(n932));
  jand g00740(.dina(\a[19] ), .dinb(\a[1] ), .dout(n933));
  jxor g00741(.dina(n933), .dinb(n932), .dout(n934));
  jnot g00742(.din(n846), .dout(n935));
  jnot g00743(.din(n847), .dout(n936));
  jand g00744(.dina(n936), .dinb(n935), .dout(n937));
  jnot g00745(.din(n937), .dout(n938));
  jand g00746(.dina(n847), .dinb(n846), .dout(n939));
  jor  g00747(.dina(n939), .dinb(n800), .dout(n940));
  jand g00748(.dina(n940), .dinb(n938), .dout(n941));
  jxor g00749(.dina(n941), .dinb(n934), .dout(n942));
  jxor g00750(.dina(n942), .dinb(n931), .dout(n943));
  jxor g00751(.dina(n943), .dinb(n929), .dout(n944));
  jand g00752(.dina(n821), .dinb(\a[10] ), .dout(n945));
  jand g00753(.dina(\a[20] ), .dinb(\a[0] ), .dout(n946));
  jxor g00754(.dina(n946), .dinb(n861), .dout(n947));
  jxor g00755(.dina(n947), .dinb(n945), .dout(n948));
  jand g00756(.dina(n859), .dinb(n856), .dout(n949));
  jor  g00757(.dina(n949), .dinb(n862), .dout(n950));
  jxor g00758(.dina(n950), .dinb(n948), .dout(n951));
  jnot g00759(.din(n951), .dout(n952));
  jand g00760(.dina(\a[12] ), .dinb(\a[8] ), .dout(n953));
  jand g00761(.dina(\a[15] ), .dinb(\a[5] ), .dout(n954));
  jand g00762(.dina(\a[14] ), .dinb(\a[6] ), .dout(n955));
  jor  g00763(.dina(n955), .dinb(n954), .dout(n956));
  jnot g00764(.din(n956), .dout(n957));
  jand g00765(.dina(\a[15] ), .dinb(\a[6] ), .dout(n958));
  jand g00766(.dina(n958), .dinb(n856), .dout(n959));
  jor  g00767(.dina(n959), .dinb(n957), .dout(n960));
  jxor g00768(.dina(n960), .dinb(n953), .dout(n961));
  jxor g00769(.dina(n961), .dinb(n952), .dout(n962));
  jxor g00770(.dina(n962), .dinb(n944), .dout(n963));
  jxor g00771(.dina(n963), .dinb(n926), .dout(n964));
  jxor g00772(.dina(n964), .dinb(n904), .dout(n965));
  jand g00773(.dina(n893), .dinb(n890), .dout(n966));
  jnot g00774(.din(n890), .dout(n967));
  jnot g00775(.din(n893), .dout(n968));
  jand g00776(.dina(n968), .dinb(n967), .dout(n969));
  jnot g00777(.din(n969), .dout(n970));
  jand g00778(.dina(n898), .dinb(n970), .dout(n971));
  jor  g00779(.dina(n971), .dinb(n966), .dout(n972));
  jxor g00780(.dina(n972), .dinb(n965), .dout(\asquared[21] ));
  jand g00781(.dina(n925), .dinb(n922), .dout(n974));
  jand g00782(.dina(n963), .dinb(n926), .dout(n975));
  jor  g00783(.dina(n975), .dinb(n974), .dout(n976));
  jand g00784(.dina(n911), .dinb(n908), .dout(n977));
  jor  g00785(.dina(n977), .dinb(n913), .dout(n978));
  jand g00786(.dina(n956), .dinb(n953), .dout(n979));
  jor  g00787(.dina(n979), .dinb(n959), .dout(n980));
  jxor g00788(.dina(n980), .dinb(n978), .dout(n981));
  jand g00789(.dina(n946), .dinb(n861), .dout(n982));
  jand g00790(.dina(n947), .dinb(n945), .dout(n983));
  jor  g00791(.dina(n983), .dinb(n982), .dout(n984));
  jxor g00792(.dina(n984), .dinb(n981), .dout(n985));
  jnot g00793(.din(n985), .dout(n986));
  jor  g00794(.dina(n915), .dinb(n907), .dout(n987));
  jand g00795(.dina(n921), .dinb(n916), .dout(n988));
  jnot g00796(.din(n988), .dout(n989));
  jand g00797(.dina(n989), .dinb(n987), .dout(n990));
  jxor g00798(.dina(n990), .dinb(n986), .dout(n991));
  jnot g00799(.din(n873), .dout(n992));
  jand g00800(.dina(\a[11] ), .dinb(\a[10] ), .dout(n993));
  jand g00801(.dina(\a[12] ), .dinb(\a[9] ), .dout(n994));
  jor  g00802(.dina(n994), .dinb(n993), .dout(n995));
  jand g00803(.dina(\a[12] ), .dinb(\a[10] ), .dout(n996));
  jand g00804(.dina(n996), .dinb(n932), .dout(n997));
  jnot g00805(.din(n997), .dout(n998));
  jand g00806(.dina(n998), .dinb(n995), .dout(n999));
  jxor g00807(.dina(n999), .dinb(n992), .dout(n1000));
  jnot g00808(.din(n958), .dout(n1001));
  jand g00809(.dina(\a[13] ), .dinb(\a[8] ), .dout(n1002));
  jand g00810(.dina(\a[14] ), .dinb(\a[7] ), .dout(n1003));
  jor  g00811(.dina(n1003), .dinb(n1002), .dout(n1004));
  jand g00812(.dina(\a[14] ), .dinb(\a[8] ), .dout(n1005));
  jand g00813(.dina(n1005), .dinb(n861), .dout(n1006));
  jnot g00814(.din(n1006), .dout(n1007));
  jand g00815(.dina(n1007), .dinb(n1004), .dout(n1008));
  jxor g00816(.dina(n1008), .dinb(n1001), .dout(n1009));
  jand g00817(.dina(n798), .dinb(\a[19] ), .dout(n1010));
  jand g00818(.dina(\a[18] ), .dinb(\a[3] ), .dout(n1011));
  jand g00819(.dina(n1011), .dinb(\a[16] ), .dout(n1012));
  jor  g00820(.dina(n1012), .dinb(n1010), .dout(n1013));
  jand g00821(.dina(n1013), .dinb(\a[5] ), .dout(n1014));
  jnot g00822(.din(n1014), .dout(n1015));
  jand g00823(.dina(\a[19] ), .dinb(\a[2] ), .dout(n1016));
  jor  g00824(.dina(n1016), .dinb(n1011), .dout(n1017));
  jand g00825(.dina(\a[19] ), .dinb(\a[3] ), .dout(n1018));
  jand g00826(.dina(n1018), .dinb(n908), .dout(n1019));
  jnot g00827(.din(n1019), .dout(n1020));
  jand g00828(.dina(n1020), .dinb(n1017), .dout(n1021));
  jand g00829(.dina(n1021), .dinb(n1015), .dout(n1022));
  jnot g00830(.din(n1021), .dout(n1023));
  jand g00831(.dina(\a[16] ), .dinb(\a[5] ), .dout(n1024));
  jand g00832(.dina(n1024), .dinb(n1023), .dout(n1025));
  jor  g00833(.dina(n1025), .dinb(n1022), .dout(n1026));
  jxor g00834(.dina(n1026), .dinb(n1009), .dout(n1027));
  jxor g00835(.dina(n1027), .dinb(n1000), .dout(n1028));
  jxor g00836(.dina(n1028), .dinb(n991), .dout(n1029));
  jand g00837(.dina(n941), .dinb(n934), .dout(n1030));
  jand g00838(.dina(n942), .dinb(n931), .dout(n1031));
  jor  g00839(.dina(n1031), .dinb(n1030), .dout(n1032));
  jand g00840(.dina(n933), .dinb(n932), .dout(n1033));
  jand g00841(.dina(\a[21] ), .dinb(\a[0] ), .dout(n1034));
  jxor g00842(.dina(n1034), .dinb(n1033), .dout(n1035));
  jand g00843(.dina(\a[20] ), .dinb(\a[1] ), .dout(n1036));
  jxor g00844(.dina(n1036), .dinb(\a[11] ), .dout(n1037));
  jxor g00845(.dina(n1037), .dinb(n1035), .dout(n1038));
  jxor g00846(.dina(n1038), .dinb(n1032), .dout(n1039));
  jnot g00847(.din(n1039), .dout(n1040));
  jand g00848(.dina(n950), .dinb(n948), .dout(n1041));
  jnot g00849(.din(n1041), .dout(n1042));
  jor  g00850(.dina(n961), .dinb(n952), .dout(n1043));
  jand g00851(.dina(n1043), .dinb(n1042), .dout(n1044));
  jxor g00852(.dina(n1044), .dinb(n1040), .dout(n1045));
  jand g00853(.dina(n943), .dinb(n929), .dout(n1046));
  jand g00854(.dina(n962), .dinb(n944), .dout(n1047));
  jor  g00855(.dina(n1047), .dinb(n1046), .dout(n1048));
  jxor g00856(.dina(n1048), .dinb(n1045), .dout(n1049));
  jxor g00857(.dina(n1049), .dinb(n1029), .dout(n1050));
  jxor g00858(.dina(n1050), .dinb(n976), .dout(n1051));
  jand g00859(.dina(n964), .dinb(n904), .dout(n1052));
  jor  g00860(.dina(n964), .dinb(n904), .dout(n1053));
  jand g00861(.dina(n972), .dinb(n1053), .dout(n1054));
  jor  g00862(.dina(n1054), .dinb(n1052), .dout(n1055));
  jxor g00863(.dina(n1055), .dinb(n1051), .dout(\asquared[22] ));
  jand g00864(.dina(n1048), .dinb(n1045), .dout(n1057));
  jand g00865(.dina(n1049), .dinb(n1029), .dout(n1058));
  jor  g00866(.dina(n1058), .dinb(n1057), .dout(n1059));
  jand g00867(.dina(n1020), .dinb(n1015), .dout(n1060));
  jnot g00868(.din(n1060), .dout(n1061));
  jand g00869(.dina(n1004), .dinb(n958), .dout(n1062));
  jor  g00870(.dina(n1062), .dinb(n1006), .dout(n1063));
  jxor g00871(.dina(n1063), .dinb(n1061), .dout(n1064));
  jand g00872(.dina(n1034), .dinb(n1033), .dout(n1065));
  jand g00873(.dina(n1037), .dinb(n1035), .dout(n1066));
  jor  g00874(.dina(n1066), .dinb(n1065), .dout(n1067));
  jxor g00875(.dina(n1067), .dinb(n1064), .dout(n1068));
  jnot g00876(.din(n1068), .dout(n1069));
  jand g00877(.dina(n1038), .dinb(n1032), .dout(n1070));
  jnot g00878(.din(n1070), .dout(n1071));
  jor  g00879(.dina(n1044), .dinb(n1040), .dout(n1072));
  jand g00880(.dina(n1072), .dinb(n1071), .dout(n1073));
  jxor g00881(.dina(n1073), .dinb(n1069), .dout(n1074));
  jand g00882(.dina(\a[13] ), .dinb(\a[9] ), .dout(n1075));
  jnot g00883(.din(n639), .dout(n1076));
  jand g00884(.dina(\a[20] ), .dinb(\a[2] ), .dout(n1077));
  jxor g00885(.dina(n1077), .dinb(n1076), .dout(n1078));
  jxor g00886(.dina(n1078), .dinb(n1075), .dout(n1079));
  jnot g00887(.din(n1079), .dout(n1080));
  jand g00888(.dina(\a[22] ), .dinb(\a[0] ), .dout(n1081));
  jand g00889(.dina(\a[15] ), .dinb(\a[7] ), .dout(n1082));
  jor  g00890(.dina(n1082), .dinb(n1005), .dout(n1083));
  jand g00891(.dina(\a[15] ), .dinb(\a[8] ), .dout(n1084));
  jand g00892(.dina(n1084), .dinb(n1003), .dout(n1085));
  jnot g00893(.din(n1085), .dout(n1086));
  jand g00894(.dina(n1086), .dinb(n1083), .dout(n1087));
  jxor g00895(.dina(n1087), .dinb(n1081), .dout(n1088));
  jxor g00896(.dina(n1088), .dinb(n1080), .dout(n1089));
  jand g00897(.dina(\a[19] ), .dinb(\a[4] ), .dout(n1090));
  jand g00898(.dina(n1090), .dinb(n1011), .dout(n1091));
  jand g00899(.dina(\a[17] ), .dinb(\a[5] ), .dout(n1092));
  jand g00900(.dina(n1092), .dinb(n1018), .dout(n1093));
  jor  g00901(.dina(n1093), .dinb(n1091), .dout(n1094));
  jand g00902(.dina(\a[18] ), .dinb(\a[5] ), .dout(n1095));
  jand g00903(.dina(n1095), .dinb(n873), .dout(n1096));
  jnot g00904(.din(n1096), .dout(n1097));
  jand g00905(.dina(n1097), .dinb(n1094), .dout(n1098));
  jnot g00906(.din(n1098), .dout(n1099));
  jand g00907(.dina(\a[18] ), .dinb(\a[4] ), .dout(n1100));
  jor  g00908(.dina(n1100), .dinb(n1092), .dout(n1101));
  jand g00909(.dina(n1101), .dinb(n1097), .dout(n1102));
  jor  g00910(.dina(n1102), .dinb(n1018), .dout(n1103));
  jand g00911(.dina(n1103), .dinb(n1099), .dout(n1104));
  jxor g00912(.dina(n1104), .dinb(n1089), .dout(n1105));
  jxor g00913(.dina(n1105), .dinb(n1074), .dout(n1106));
  jor  g00914(.dina(n990), .dinb(n986), .dout(n1107));
  jand g00915(.dina(n1028), .dinb(n991), .dout(n1108));
  jnot g00916(.din(n1108), .dout(n1109));
  jand g00917(.dina(n1109), .dinb(n1107), .dout(n1110));
  jnot g00918(.din(n1110), .dout(n1111));
  jand g00919(.dina(n980), .dinb(n978), .dout(n1112));
  jand g00920(.dina(n984), .dinb(n981), .dout(n1113));
  jor  g00921(.dina(n1113), .dinb(n1112), .dout(n1114));
  jand g00922(.dina(n1036), .dinb(\a[11] ), .dout(n1115));
  jand g00923(.dina(\a[21] ), .dinb(\a[1] ), .dout(n1116));
  jxor g00924(.dina(n1116), .dinb(n996), .dout(n1117));
  jxor g00925(.dina(n1117), .dinb(n1115), .dout(n1118));
  jand g00926(.dina(n995), .dinb(n873), .dout(n1119));
  jor  g00927(.dina(n1119), .dinb(n997), .dout(n1120));
  jxor g00928(.dina(n1120), .dinb(n1118), .dout(n1121));
  jxor g00929(.dina(n1121), .dinb(n1114), .dout(n1122));
  jnot g00930(.din(n1122), .dout(n1123));
  jnot g00931(.din(n1009), .dout(n1124));
  jand g00932(.dina(n1026), .dinb(n1124), .dout(n1125));
  jnot g00933(.din(n1125), .dout(n1126));
  jnot g00934(.din(n1026), .dout(n1127));
  jand g00935(.dina(n1127), .dinb(n1009), .dout(n1128));
  jor  g00936(.dina(n1128), .dinb(n1000), .dout(n1129));
  jand g00937(.dina(n1129), .dinb(n1126), .dout(n1130));
  jxor g00938(.dina(n1130), .dinb(n1123), .dout(n1131));
  jxor g00939(.dina(n1131), .dinb(n1111), .dout(n1132));
  jxor g00940(.dina(n1132), .dinb(n1106), .dout(n1133));
  jxor g00941(.dina(n1133), .dinb(n1059), .dout(n1134));
  jand g00942(.dina(n1050), .dinb(n976), .dout(n1135));
  jor  g00943(.dina(n1050), .dinb(n976), .dout(n1136));
  jand g00944(.dina(n1055), .dinb(n1136), .dout(n1137));
  jor  g00945(.dina(n1137), .dinb(n1135), .dout(n1138));
  jxor g00946(.dina(n1138), .dinb(n1134), .dout(\asquared[23] ));
  jand g00947(.dina(n1131), .dinb(n1111), .dout(n1140));
  jand g00948(.dina(n1132), .dinb(n1106), .dout(n1141));
  jor  g00949(.dina(n1141), .dinb(n1140), .dout(n1142));
  jand g00950(.dina(n1121), .dinb(n1114), .dout(n1143));
  jnot g00951(.din(n1143), .dout(n1144));
  jor  g00952(.dina(n1130), .dinb(n1123), .dout(n1145));
  jand g00953(.dina(n1145), .dinb(n1144), .dout(n1146));
  jand g00954(.dina(n1117), .dinb(n1115), .dout(n1147));
  jand g00955(.dina(n1120), .dinb(n1118), .dout(n1148));
  jor  g00956(.dina(n1148), .dinb(n1147), .dout(n1149));
  jand g00957(.dina(\a[12] ), .dinb(\a[11] ), .dout(n1150));
  jand g00958(.dina(\a[13] ), .dinb(\a[10] ), .dout(n1151));
  jor  g00959(.dina(n1151), .dinb(n1150), .dout(n1152));
  jnot g00960(.din(n1152), .dout(n1153));
  jand g00961(.dina(\a[13] ), .dinb(\a[11] ), .dout(n1154));
  jand g00962(.dina(n1154), .dinb(n996), .dout(n1155));
  jor  g00963(.dina(n1155), .dinb(n1153), .dout(n1156));
  jxor g00964(.dina(n1156), .dinb(n1090), .dout(n1157));
  jnot g00965(.din(n1157), .dout(n1158));
  jand g00966(.dina(\a[17] ), .dinb(\a[6] ), .dout(n1159));
  jand g00967(.dina(\a[20] ), .dinb(\a[3] ), .dout(n1160));
  jor  g00968(.dina(n1160), .dinb(n1095), .dout(n1161));
  jand g00969(.dina(\a[20] ), .dinb(\a[5] ), .dout(n1162));
  jand g00970(.dina(n1162), .dinb(n1011), .dout(n1163));
  jnot g00971(.din(n1163), .dout(n1164));
  jand g00972(.dina(n1164), .dinb(n1161), .dout(n1165));
  jxor g00973(.dina(n1165), .dinb(n1159), .dout(n1166));
  jxor g00974(.dina(n1166), .dinb(n1158), .dout(n1167));
  jxor g00975(.dina(n1167), .dinb(n1149), .dout(n1168));
  jand g00976(.dina(\a[16] ), .dinb(\a[7] ), .dout(n1169));
  jand g00977(.dina(\a[14] ), .dinb(\a[9] ), .dout(n1170));
  jor  g00978(.dina(n1170), .dinb(n1084), .dout(n1171));
  jnot g00979(.din(n1171), .dout(n1172));
  jand g00980(.dina(\a[15] ), .dinb(\a[9] ), .dout(n1173));
  jand g00981(.dina(n1173), .dinb(n1005), .dout(n1174));
  jor  g00982(.dina(n1174), .dinb(n1172), .dout(n1175));
  jxor g00983(.dina(n1175), .dinb(n1169), .dout(n1176));
  jnot g00984(.din(n1176), .dout(n1177));
  jand g00985(.dina(n1087), .dinb(n1081), .dout(n1178));
  jor  g00986(.dina(n1178), .dinb(n1085), .dout(n1179));
  jnot g00987(.din(n1179), .dout(n1180));
  jand g00988(.dina(n1116), .dinb(n996), .dout(n1181));
  jand g00989(.dina(\a[23] ), .dinb(\a[0] ), .dout(n1182));
  jand g00990(.dina(\a[21] ), .dinb(\a[2] ), .dout(n1183));
  jor  g00991(.dina(n1183), .dinb(n1182), .dout(n1184));
  jnot g00992(.din(n1184), .dout(n1185));
  jand g00993(.dina(\a[23] ), .dinb(\a[2] ), .dout(n1186));
  jand g00994(.dina(n1186), .dinb(n1034), .dout(n1187));
  jor  g00995(.dina(n1187), .dinb(n1185), .dout(n1188));
  jxor g00996(.dina(n1188), .dinb(n1181), .dout(n1189));
  jxor g00997(.dina(n1189), .dinb(n1180), .dout(n1190));
  jxor g00998(.dina(n1190), .dinb(n1177), .dout(n1191));
  jxor g00999(.dina(n1191), .dinb(n1168), .dout(n1192));
  jnot g01000(.din(n1192), .dout(n1193));
  jxor g01001(.dina(n1193), .dinb(n1146), .dout(n1194));
  jor  g01002(.dina(n1073), .dinb(n1069), .dout(n1195));
  jand g01003(.dina(n1105), .dinb(n1074), .dout(n1196));
  jnot g01004(.din(n1196), .dout(n1197));
  jand g01005(.dina(n1197), .dinb(n1195), .dout(n1198));
  jnot g01006(.din(n1198), .dout(n1199));
  jand g01007(.dina(n1063), .dinb(n1061), .dout(n1200));
  jand g01008(.dina(n1067), .dinb(n1064), .dout(n1201));
  jor  g01009(.dina(n1201), .dinb(n1200), .dout(n1202));
  jand g01010(.dina(n1088), .dinb(n1080), .dout(n1203));
  jand g01011(.dina(n1104), .dinb(n1089), .dout(n1204));
  jor  g01012(.dina(n1204), .dinb(n1203), .dout(n1205));
  jxor g01013(.dina(n1205), .dinb(n1202), .dout(n1206));
  jand g01014(.dina(\a[22] ), .dinb(\a[1] ), .dout(n1207));
  jxor g01015(.dina(n1207), .dinb(\a[12] ), .dout(n1208));
  jor  g01016(.dina(n1096), .dinb(n1094), .dout(n1209));
  jxor g01017(.dina(n1209), .dinb(n1208), .dout(n1210));
  jnot g01018(.din(n1077), .dout(n1211));
  jand g01019(.dina(n1211), .dinb(n1076), .dout(n1212));
  jnot g01020(.din(n1212), .dout(n1213));
  jand g01021(.dina(n1077), .dinb(n639), .dout(n1214));
  jor  g01022(.dina(n1214), .dinb(n1075), .dout(n1215));
  jand g01023(.dina(n1215), .dinb(n1213), .dout(n1216));
  jxor g01024(.dina(n1216), .dinb(n1210), .dout(n1217));
  jxor g01025(.dina(n1217), .dinb(n1206), .dout(n1218));
  jxor g01026(.dina(n1218), .dinb(n1199), .dout(n1219));
  jxor g01027(.dina(n1219), .dinb(n1194), .dout(n1220));
  jxor g01028(.dina(n1220), .dinb(n1142), .dout(n1221));
  jand g01029(.dina(n1133), .dinb(n1059), .dout(n1222));
  jor  g01030(.dina(n1133), .dinb(n1059), .dout(n1223));
  jand g01031(.dina(n1138), .dinb(n1223), .dout(n1224));
  jor  g01032(.dina(n1224), .dinb(n1222), .dout(n1225));
  jxor g01033(.dina(n1225), .dinb(n1221), .dout(\asquared[24] ));
  jand g01034(.dina(n1218), .dinb(n1199), .dout(n1227));
  jand g01035(.dina(n1219), .dinb(n1194), .dout(n1228));
  jor  g01036(.dina(n1228), .dinb(n1227), .dout(n1229));
  jand g01037(.dina(n1209), .dinb(n1208), .dout(n1230));
  jand g01038(.dina(n1216), .dinb(n1210), .dout(n1231));
  jor  g01039(.dina(n1231), .dinb(n1230), .dout(n1232));
  jand g01040(.dina(n1207), .dinb(\a[12] ), .dout(n1233));
  jand g01041(.dina(\a[24] ), .dinb(\a[0] ), .dout(n1234));
  jxor g01042(.dina(n1234), .dinb(n1233), .dout(n1235));
  jand g01043(.dina(\a[23] ), .dinb(\a[1] ), .dout(n1236));
  jxor g01044(.dina(n1236), .dinb(n1154), .dout(n1237));
  jnot g01045(.din(n1237), .dout(n1238));
  jxor g01046(.dina(n1238), .dinb(n1235), .dout(n1239));
  jand g01047(.dina(\a[17] ), .dinb(\a[7] ), .dout(n1240));
  jand g01048(.dina(\a[22] ), .dinb(\a[2] ), .dout(n1241));
  jand g01049(.dina(\a[18] ), .dinb(\a[6] ), .dout(n1242));
  jor  g01050(.dina(n1242), .dinb(n1241), .dout(n1243));
  jnot g01051(.din(n1243), .dout(n1244));
  jand g01052(.dina(\a[22] ), .dinb(\a[6] ), .dout(n1245));
  jand g01053(.dina(n1245), .dinb(n908), .dout(n1246));
  jor  g01054(.dina(n1246), .dinb(n1244), .dout(n1247));
  jxor g01055(.dina(n1247), .dinb(n1240), .dout(n1248));
  jxor g01056(.dina(n1248), .dinb(n1239), .dout(n1249));
  jxor g01057(.dina(n1249), .dinb(n1232), .dout(n1250));
  jand g01058(.dina(\a[16] ), .dinb(\a[8] ), .dout(n1251));
  jand g01059(.dina(\a[14] ), .dinb(\a[10] ), .dout(n1252));
  jor  g01060(.dina(n1252), .dinb(n1173), .dout(n1253));
  jnot g01061(.din(n1253), .dout(n1254));
  jand g01062(.dina(n1170), .dinb(n599), .dout(n1255));
  jor  g01063(.dina(n1255), .dinb(n1254), .dout(n1256));
  jxor g01064(.dina(n1256), .dinb(n1251), .dout(n1257));
  jnot g01065(.din(n1257), .dout(n1258));
  jand g01066(.dina(\a[21] ), .dinb(\a[3] ), .dout(n1259));
  jand g01067(.dina(\a[19] ), .dinb(\a[5] ), .dout(n1260));
  jand g01068(.dina(\a[20] ), .dinb(\a[4] ), .dout(n1261));
  jor  g01069(.dina(n1261), .dinb(n1260), .dout(n1262));
  jnot g01070(.din(n1262), .dout(n1263));
  jand g01071(.dina(n1162), .dinb(n1090), .dout(n1264));
  jor  g01072(.dina(n1264), .dinb(n1263), .dout(n1265));
  jxor g01073(.dina(n1265), .dinb(n1259), .dout(n1266));
  jnot g01074(.din(n1266), .dout(n1267));
  jand g01075(.dina(n1184), .dinb(n1181), .dout(n1268));
  jor  g01076(.dina(n1268), .dinb(n1187), .dout(n1269));
  jxor g01077(.dina(n1269), .dinb(n1267), .dout(n1270));
  jxor g01078(.dina(n1270), .dinb(n1258), .dout(n1271));
  jxor g01079(.dina(n1271), .dinb(n1250), .dout(n1272));
  jand g01080(.dina(n1205), .dinb(n1202), .dout(n1273));
  jand g01081(.dina(n1217), .dinb(n1206), .dout(n1274));
  jor  g01082(.dina(n1274), .dinb(n1273), .dout(n1275));
  jxor g01083(.dina(n1275), .dinb(n1272), .dout(n1276));
  jand g01084(.dina(n1191), .dinb(n1168), .dout(n1277));
  jnot g01085(.din(n1277), .dout(n1278));
  jor  g01086(.dina(n1193), .dinb(n1146), .dout(n1279));
  jand g01087(.dina(n1279), .dinb(n1278), .dout(n1280));
  jand g01088(.dina(n1165), .dinb(n1159), .dout(n1281));
  jor  g01089(.dina(n1281), .dinb(n1163), .dout(n1282));
  jand g01090(.dina(n1152), .dinb(n1090), .dout(n1283));
  jor  g01091(.dina(n1283), .dinb(n1155), .dout(n1284));
  jxor g01092(.dina(n1284), .dinb(n1282), .dout(n1285));
  jand g01093(.dina(n1171), .dinb(n1169), .dout(n1286));
  jor  g01094(.dina(n1286), .dinb(n1174), .dout(n1287));
  jxor g01095(.dina(n1287), .dinb(n1285), .dout(n1288));
  jand g01096(.dina(n1166), .dinb(n1158), .dout(n1289));
  jand g01097(.dina(n1167), .dinb(n1149), .dout(n1290));
  jor  g01098(.dina(n1290), .dinb(n1289), .dout(n1291));
  jnot g01099(.din(n1291), .dout(n1292));
  jor  g01100(.dina(n1189), .dinb(n1180), .dout(n1293));
  jand g01101(.dina(n1190), .dinb(n1177), .dout(n1294));
  jnot g01102(.din(n1294), .dout(n1295));
  jand g01103(.dina(n1295), .dinb(n1293), .dout(n1296));
  jxor g01104(.dina(n1296), .dinb(n1292), .dout(n1297));
  jxor g01105(.dina(n1297), .dinb(n1288), .dout(n1298));
  jnot g01106(.din(n1298), .dout(n1299));
  jxor g01107(.dina(n1299), .dinb(n1280), .dout(n1300));
  jxor g01108(.dina(n1300), .dinb(n1276), .dout(n1301));
  jxor g01109(.dina(n1301), .dinb(n1229), .dout(n1302));
  jand g01110(.dina(n1220), .dinb(n1142), .dout(n1303));
  jnot g01111(.din(n1142), .dout(n1304));
  jnot g01112(.din(n1220), .dout(n1305));
  jand g01113(.dina(n1305), .dinb(n1304), .dout(n1306));
  jnot g01114(.din(n1306), .dout(n1307));
  jand g01115(.dina(n1225), .dinb(n1307), .dout(n1308));
  jor  g01116(.dina(n1308), .dinb(n1303), .dout(n1309));
  jxor g01117(.dina(n1309), .dinb(n1302), .dout(\asquared[25] ));
  jor  g01118(.dina(n1299), .dinb(n1280), .dout(n1311));
  jand g01119(.dina(n1300), .dinb(n1276), .dout(n1312));
  jnot g01120(.din(n1312), .dout(n1313));
  jand g01121(.dina(n1313), .dinb(n1311), .dout(n1314));
  jand g01122(.dina(n1243), .dinb(n1240), .dout(n1315));
  jor  g01123(.dina(n1315), .dinb(n1246), .dout(n1316));
  jand g01124(.dina(n1253), .dinb(n1251), .dout(n1317));
  jor  g01125(.dina(n1317), .dinb(n1255), .dout(n1318));
  jxor g01126(.dina(n1318), .dinb(n1316), .dout(n1319));
  jor  g01127(.dina(n1234), .dinb(n1233), .dout(n1320));
  jand g01128(.dina(n1234), .dinb(n1233), .dout(n1321));
  jor  g01129(.dina(n1237), .dinb(n1321), .dout(n1322));
  jand g01130(.dina(n1322), .dinb(n1320), .dout(n1323));
  jxor g01131(.dina(n1323), .dinb(n1319), .dout(n1324));
  jand g01132(.dina(n1269), .dinb(n1267), .dout(n1325));
  jand g01133(.dina(n1270), .dinb(n1258), .dout(n1326));
  jor  g01134(.dina(n1326), .dinb(n1325), .dout(n1327));
  jxor g01135(.dina(n1327), .dinb(n1324), .dout(n1328));
  jnot g01136(.din(n1328), .dout(n1329));
  jor  g01137(.dina(n1248), .dinb(n1239), .dout(n1330));
  jand g01138(.dina(n1249), .dinb(n1232), .dout(n1331));
  jnot g01139(.din(n1331), .dout(n1332));
  jand g01140(.dina(n1332), .dinb(n1330), .dout(n1333));
  jxor g01141(.dina(n1333), .dinb(n1329), .dout(n1334));
  jand g01142(.dina(n1271), .dinb(n1250), .dout(n1335));
  jand g01143(.dina(n1275), .dinb(n1272), .dout(n1336));
  jor  g01144(.dina(n1336), .dinb(n1335), .dout(n1337));
  jxor g01145(.dina(n1337), .dinb(n1334), .dout(n1338));
  jand g01146(.dina(n1262), .dinb(n1259), .dout(n1339));
  jor  g01147(.dina(n1339), .dinb(n1264), .dout(n1340));
  jand g01148(.dina(\a[24] ), .dinb(\a[1] ), .dout(n1341));
  jnot g01149(.din(\a[13] ), .dout(n1342));
  jand g01150(.dina(n1236), .dinb(n1154), .dout(n1343));
  jor  g01151(.dina(n1343), .dinb(n1342), .dout(n1344));
  jxor g01152(.dina(n1344), .dinb(n1341), .dout(n1345));
  jnot g01153(.din(n1345), .dout(n1346));
  jxor g01154(.dina(n1346), .dinb(n1340), .dout(n1347));
  jand g01155(.dina(n1284), .dinb(n1282), .dout(n1348));
  jand g01156(.dina(n1287), .dinb(n1285), .dout(n1349));
  jor  g01157(.dina(n1349), .dinb(n1348), .dout(n1350));
  jnot g01158(.din(n1350), .dout(n1351));
  jand g01159(.dina(\a[13] ), .dinb(\a[12] ), .dout(n1352));
  jnot g01160(.din(n1352), .dout(n1353));
  jand g01161(.dina(\a[14] ), .dinb(\a[11] ), .dout(n1354));
  jxor g01162(.dina(n1354), .dinb(n1353), .dout(n1355));
  jxor g01163(.dina(n1355), .dinb(n1162), .dout(n1356));
  jxor g01164(.dina(n1356), .dinb(n1351), .dout(n1357));
  jxor g01165(.dina(n1357), .dinb(n1347), .dout(n1358));
  jor  g01166(.dina(n1296), .dinb(n1292), .dout(n1359));
  jand g01167(.dina(n1297), .dinb(n1288), .dout(n1360));
  jnot g01168(.din(n1360), .dout(n1361));
  jand g01169(.dina(n1361), .dinb(n1359), .dout(n1362));
  jnot g01170(.din(n1362), .dout(n1363));
  jand g01171(.dina(\a[25] ), .dinb(\a[0] ), .dout(n1364));
  jor  g01172(.dina(n1364), .dinb(n1186), .dout(n1365));
  jand g01173(.dina(\a[25] ), .dinb(\a[2] ), .dout(n1366));
  jand g01174(.dina(n1366), .dinb(n1182), .dout(n1367));
  jnot g01175(.din(n1367), .dout(n1368));
  jand g01176(.dina(n1368), .dinb(n1365), .dout(n1369));
  jxor g01177(.dina(n1369), .dinb(n599), .dout(n1370));
  jnot g01178(.din(n1370), .dout(n1371));
  jand g01179(.dina(\a[18] ), .dinb(\a[7] ), .dout(n1372));
  jnot g01180(.din(n1372), .dout(n1373));
  jand g01181(.dina(\a[17] ), .dinb(\a[8] ), .dout(n1374));
  jor  g01182(.dina(n1374), .dinb(n739), .dout(n1375));
  jand g01183(.dina(\a[17] ), .dinb(\a[9] ), .dout(n1376));
  jand g01184(.dina(n1376), .dinb(n1251), .dout(n1377));
  jnot g01185(.din(n1377), .dout(n1378));
  jand g01186(.dina(n1378), .dinb(n1375), .dout(n1379));
  jxor g01187(.dina(n1379), .dinb(n1373), .dout(n1380));
  jxor g01188(.dina(n1380), .dinb(n1371), .dout(n1381));
  jand g01189(.dina(n1018), .dinb(\a[22] ), .dout(n1382));
  jand g01190(.dina(\a[21] ), .dinb(\a[4] ), .dout(n1383));
  jand g01191(.dina(n1383), .dinb(\a[19] ), .dout(n1384));
  jor  g01192(.dina(n1384), .dinb(n1382), .dout(n1385));
  jand g01193(.dina(n1385), .dinb(\a[6] ), .dout(n1386));
  jnot g01194(.din(n1386), .dout(n1387));
  jand g01195(.dina(\a[22] ), .dinb(\a[3] ), .dout(n1388));
  jor  g01196(.dina(n1388), .dinb(n1383), .dout(n1389));
  jand g01197(.dina(\a[22] ), .dinb(\a[4] ), .dout(n1390));
  jand g01198(.dina(n1390), .dinb(n1259), .dout(n1391));
  jnot g01199(.din(n1391), .dout(n1392));
  jand g01200(.dina(n1392), .dinb(n1389), .dout(n1393));
  jand g01201(.dina(n1393), .dinb(n1387), .dout(n1394));
  jnot g01202(.din(n1393), .dout(n1395));
  jand g01203(.dina(\a[19] ), .dinb(\a[6] ), .dout(n1396));
  jand g01204(.dina(n1396), .dinb(n1395), .dout(n1397));
  jor  g01205(.dina(n1397), .dinb(n1394), .dout(n1398));
  jxor g01206(.dina(n1398), .dinb(n1381), .dout(n1399));
  jxor g01207(.dina(n1399), .dinb(n1363), .dout(n1400));
  jxor g01208(.dina(n1400), .dinb(n1358), .dout(n1401));
  jxor g01209(.dina(n1401), .dinb(n1338), .dout(n1402));
  jnot g01210(.din(n1402), .dout(n1403));
  jxor g01211(.dina(n1403), .dinb(n1314), .dout(n1404));
  jand g01212(.dina(n1301), .dinb(n1229), .dout(n1405));
  jor  g01213(.dina(n1301), .dinb(n1229), .dout(n1406));
  jand g01214(.dina(n1309), .dinb(n1406), .dout(n1407));
  jor  g01215(.dina(n1407), .dinb(n1405), .dout(n1408));
  jxor g01216(.dina(n1408), .dinb(n1404), .dout(\asquared[26] ));
  jand g01217(.dina(n1337), .dinb(n1334), .dout(n1410));
  jand g01218(.dina(n1401), .dinb(n1338), .dout(n1411));
  jor  g01219(.dina(n1411), .dinb(n1410), .dout(n1412));
  jand g01220(.dina(n1399), .dinb(n1363), .dout(n1413));
  jand g01221(.dina(n1400), .dinb(n1358), .dout(n1414));
  jor  g01222(.dina(n1414), .dinb(n1413), .dout(n1415));
  jor  g01223(.dina(n1356), .dinb(n1351), .dout(n1416));
  jand g01224(.dina(n1357), .dinb(n1347), .dout(n1417));
  jnot g01225(.din(n1417), .dout(n1418));
  jand g01226(.dina(n1418), .dinb(n1416), .dout(n1419));
  jnot g01227(.din(n1419), .dout(n1420));
  jand g01228(.dina(n1392), .dinb(n1387), .dout(n1421));
  jnot g01229(.din(n1421), .dout(n1422));
  jand g01230(.dina(\a[14] ), .dinb(\a[12] ), .dout(n1423));
  jand g01231(.dina(\a[25] ), .dinb(\a[1] ), .dout(n1424));
  jxor g01232(.dina(n1424), .dinb(n1423), .dout(n1425));
  jnot g01233(.din(n1354), .dout(n1426));
  jand g01234(.dina(n1426), .dinb(n1353), .dout(n1427));
  jnot g01235(.din(n1427), .dout(n1428));
  jand g01236(.dina(n1354), .dinb(n1352), .dout(n1429));
  jor  g01237(.dina(n1429), .dinb(n1162), .dout(n1430));
  jand g01238(.dina(n1430), .dinb(n1428), .dout(n1431));
  jxor g01239(.dina(n1431), .dinb(n1425), .dout(n1432));
  jxor g01240(.dina(n1432), .dinb(n1422), .dout(n1433));
  jnot g01241(.din(n1380), .dout(n1434));
  jand g01242(.dina(n1434), .dinb(n1370), .dout(n1435));
  jand g01243(.dina(n1380), .dinb(n1371), .dout(n1436));
  jnot g01244(.din(n1436), .dout(n1437));
  jand g01245(.dina(n1398), .dinb(n1437), .dout(n1438));
  jor  g01246(.dina(n1438), .dinb(n1435), .dout(n1439));
  jxor g01247(.dina(n1439), .dinb(n1433), .dout(n1440));
  jxor g01248(.dina(n1440), .dinb(n1420), .dout(n1441));
  jxor g01249(.dina(n1441), .dinb(n1415), .dout(n1442));
  jand g01250(.dina(n1327), .dinb(n1324), .dout(n1443));
  jnot g01251(.din(n1443), .dout(n1444));
  jor  g01252(.dina(n1333), .dinb(n1329), .dout(n1445));
  jand g01253(.dina(n1445), .dinb(n1444), .dout(n1446));
  jnot g01254(.din(n1446), .dout(n1447));
  jand g01255(.dina(\a[20] ), .dinb(\a[6] ), .dout(n1448));
  jand g01256(.dina(\a[21] ), .dinb(\a[5] ), .dout(n1449));
  jor  g01257(.dina(n1449), .dinb(n1448), .dout(n1450));
  jnot g01258(.din(n1450), .dout(n1451));
  jand g01259(.dina(\a[21] ), .dinb(\a[6] ), .dout(n1452));
  jand g01260(.dina(n1452), .dinb(n1162), .dout(n1453));
  jor  g01261(.dina(n1453), .dinb(n1451), .dout(n1454));
  jxor g01262(.dina(n1454), .dinb(n1390), .dout(n1455));
  jnot g01263(.din(n1455), .dout(n1456));
  jand g01264(.dina(\a[24] ), .dinb(\a[2] ), .dout(n1457));
  jnot g01265(.din(n1457), .dout(n1458));
  jand g01266(.dina(\a[23] ), .dinb(\a[3] ), .dout(n1459));
  jand g01267(.dina(\a[19] ), .dinb(\a[7] ), .dout(n1460));
  jxor g01268(.dina(n1460), .dinb(n1459), .dout(n1461));
  jxor g01269(.dina(n1461), .dinb(n1458), .dout(n1462));
  jand g01270(.dina(\a[16] ), .dinb(\a[10] ), .dout(n1463));
  jor  g01271(.dina(n1463), .dinb(n707), .dout(n1464));
  jnot g01272(.din(n1464), .dout(n1465));
  jand g01273(.dina(\a[16] ), .dinb(\a[11] ), .dout(n1466));
  jand g01274(.dina(n1466), .dinb(n599), .dout(n1467));
  jor  g01275(.dina(n1467), .dinb(n1465), .dout(n1468));
  jxor g01276(.dina(n1468), .dinb(n1376), .dout(n1469));
  jxor g01277(.dina(n1469), .dinb(n1462), .dout(n1470));
  jxor g01278(.dina(n1470), .dinb(n1456), .dout(n1471));
  jxor g01279(.dina(n1471), .dinb(n1447), .dout(n1472));
  jand g01280(.dina(n1318), .dinb(n1316), .dout(n1473));
  jand g01281(.dina(n1323), .dinb(n1319), .dout(n1474));
  jor  g01282(.dina(n1474), .dinb(n1473), .dout(n1475));
  jand g01283(.dina(n1346), .dinb(n1340), .dout(n1476));
  jnot g01284(.din(\a[24] ), .dout(n1477));
  jand g01285(.dina(n1343), .dinb(n1477), .dout(n1478));
  jor  g01286(.dina(n1478), .dinb(n1476), .dout(n1479));
  jxor g01287(.dina(n1479), .dinb(n1475), .dout(n1480));
  jand g01288(.dina(n1369), .dinb(n599), .dout(n1481));
  jor  g01289(.dina(n1481), .dinb(n1367), .dout(n1482));
  jand g01290(.dina(n1378), .dinb(n1373), .dout(n1483));
  jnot g01291(.din(n1483), .dout(n1484));
  jand g01292(.dina(n1484), .dinb(n1375), .dout(n1485));
  jxor g01293(.dina(n1485), .dinb(n1482), .dout(n1486));
  jand g01294(.dina(n1341), .dinb(\a[13] ), .dout(n1487));
  jand g01295(.dina(\a[26] ), .dinb(\a[0] ), .dout(n1488));
  jnot g01296(.din(n1488), .dout(n1489));
  jand g01297(.dina(\a[18] ), .dinb(\a[8] ), .dout(n1490));
  jxor g01298(.dina(n1490), .dinb(n1489), .dout(n1491));
  jxor g01299(.dina(n1491), .dinb(n1487), .dout(n1492));
  jnot g01300(.din(n1492), .dout(n1493));
  jxor g01301(.dina(n1493), .dinb(n1486), .dout(n1494));
  jxor g01302(.dina(n1494), .dinb(n1480), .dout(n1495));
  jxor g01303(.dina(n1495), .dinb(n1472), .dout(n1496));
  jxor g01304(.dina(n1496), .dinb(n1442), .dout(n1497));
  jxor g01305(.dina(n1497), .dinb(n1412), .dout(n1498));
  jor  g01306(.dina(n1403), .dinb(n1314), .dout(n1499));
  jnot g01307(.din(n1499), .dout(n1500));
  jand g01308(.dina(n1403), .dinb(n1314), .dout(n1501));
  jnot g01309(.din(n1501), .dout(n1502));
  jand g01310(.dina(n1408), .dinb(n1502), .dout(n1503));
  jor  g01311(.dina(n1503), .dinb(n1500), .dout(n1504));
  jxor g01312(.dina(n1504), .dinb(n1498), .dout(\asquared[27] ));
  jand g01313(.dina(n1441), .dinb(n1415), .dout(n1506));
  jand g01314(.dina(n1496), .dinb(n1442), .dout(n1507));
  jor  g01315(.dina(n1507), .dinb(n1506), .dout(n1508));
  jand g01316(.dina(n1471), .dinb(n1447), .dout(n1509));
  jand g01317(.dina(n1495), .dinb(n1472), .dout(n1510));
  jor  g01318(.dina(n1510), .dinb(n1509), .dout(n1511));
  jand g01319(.dina(n1464), .dinb(n1376), .dout(n1512));
  jor  g01320(.dina(n1512), .dinb(n1467), .dout(n1513));
  jand g01321(.dina(n1450), .dinb(n1390), .dout(n1514));
  jor  g01322(.dina(n1514), .dinb(n1453), .dout(n1515));
  jxor g01323(.dina(n1515), .dinb(n1513), .dout(n1516));
  jand g01324(.dina(n1460), .dinb(n1459), .dout(n1517));
  jnot g01325(.din(n1517), .dout(n1518));
  jnot g01326(.din(n1459), .dout(n1519));
  jnot g01327(.din(n1460), .dout(n1520));
  jand g01328(.dina(n1520), .dinb(n1519), .dout(n1521));
  jor  g01329(.dina(n1521), .dinb(n1458), .dout(n1522));
  jand g01330(.dina(n1522), .dinb(n1518), .dout(n1523));
  jnot g01331(.din(n1523), .dout(n1524));
  jxor g01332(.dina(n1524), .dinb(n1516), .dout(n1525));
  jand g01333(.dina(n1479), .dinb(n1475), .dout(n1526));
  jand g01334(.dina(n1494), .dinb(n1480), .dout(n1527));
  jor  g01335(.dina(n1527), .dinb(n1526), .dout(n1528));
  jxor g01336(.dina(n1528), .dinb(n1525), .dout(n1529));
  jand g01337(.dina(n1424), .dinb(n1423), .dout(n1530));
  jand g01338(.dina(\a[27] ), .dinb(\a[0] ), .dout(n1531));
  jxor g01339(.dina(n1531), .dinb(n1530), .dout(n1532));
  jand g01340(.dina(n582), .dinb(\a[26] ), .dout(n1533));
  jnot g01341(.din(n1533), .dout(n1534));
  jand g01342(.dina(n1534), .dinb(\a[14] ), .dout(n1535));
  jnot g01343(.din(\a[14] ), .dout(n1536));
  jand g01344(.dina(\a[26] ), .dinb(\a[1] ), .dout(n1537));
  jand g01345(.dina(n1537), .dinb(n1536), .dout(n1538));
  jor  g01346(.dina(n1538), .dinb(n1535), .dout(n1539));
  jxor g01347(.dina(n1539), .dinb(n1532), .dout(n1540));
  jand g01348(.dina(\a[22] ), .dinb(\a[5] ), .dout(n1541));
  jand g01349(.dina(\a[14] ), .dinb(\a[13] ), .dout(n1542));
  jand g01350(.dina(\a[15] ), .dinb(\a[12] ), .dout(n1543));
  jor  g01351(.dina(n1543), .dinb(n1542), .dout(n1544));
  jnot g01352(.din(n1544), .dout(n1545));
  jand g01353(.dina(\a[15] ), .dinb(\a[13] ), .dout(n1546));
  jand g01354(.dina(n1546), .dinb(n1423), .dout(n1547));
  jor  g01355(.dina(n1547), .dinb(n1545), .dout(n1548));
  jxor g01356(.dina(n1548), .dinb(n1541), .dout(n1549));
  jand g01357(.dina(\a[24] ), .dinb(\a[3] ), .dout(n1550));
  jnot g01358(.din(n1550), .dout(n1551));
  jand g01359(.dina(\a[23] ), .dinb(\a[4] ), .dout(n1552));
  jxor g01360(.dina(n1552), .dinb(n1452), .dout(n1553));
  jxor g01361(.dina(n1553), .dinb(n1551), .dout(n1554));
  jxor g01362(.dina(n1554), .dinb(n1549), .dout(n1555));
  jxor g01363(.dina(n1555), .dinb(n1540), .dout(n1556));
  jxor g01364(.dina(n1556), .dinb(n1529), .dout(n1557));
  jxor g01365(.dina(n1557), .dinb(n1511), .dout(n1558));
  jand g01366(.dina(n1439), .dinb(n1433), .dout(n1559));
  jand g01367(.dina(n1440), .dinb(n1420), .dout(n1560));
  jor  g01368(.dina(n1560), .dinb(n1559), .dout(n1561));
  jand g01369(.dina(\a[20] ), .dinb(\a[7] ), .dout(n1562));
  jor  g01370(.dina(n1562), .dinb(n1366), .dout(n1563));
  jand g01371(.dina(\a[25] ), .dinb(\a[7] ), .dout(n1564));
  jand g01372(.dina(n1564), .dinb(n1077), .dout(n1565));
  jnot g01373(.din(n1565), .dout(n1566));
  jand g01374(.dina(n1566), .dinb(n1563), .dout(n1567));
  jxor g01375(.dina(n1567), .dinb(n1466), .dout(n1568));
  jnot g01376(.din(n1490), .dout(n1569));
  jand g01377(.dina(n1569), .dinb(n1489), .dout(n1570));
  jnot g01378(.din(n1570), .dout(n1571));
  jand g01379(.dina(n1490), .dinb(n1488), .dout(n1572));
  jor  g01380(.dina(n1572), .dinb(n1487), .dout(n1573));
  jand g01381(.dina(n1573), .dinb(n1571), .dout(n1574));
  jxor g01382(.dina(n1574), .dinb(n1568), .dout(n1575));
  jnot g01383(.din(n1575), .dout(n1576));
  jand g01384(.dina(\a[19] ), .dinb(\a[8] ), .dout(n1577));
  jand g01385(.dina(\a[18] ), .dinb(\a[9] ), .dout(n1578));
  jand g01386(.dina(\a[17] ), .dinb(\a[10] ), .dout(n1579));
  jor  g01387(.dina(n1579), .dinb(n1578), .dout(n1580));
  jnot g01388(.din(n1580), .dout(n1581));
  jand g01389(.dina(\a[18] ), .dinb(\a[10] ), .dout(n1582));
  jand g01390(.dina(n1582), .dinb(n1376), .dout(n1583));
  jor  g01391(.dina(n1583), .dinb(n1581), .dout(n1584));
  jxor g01392(.dina(n1584), .dinb(n1577), .dout(n1585));
  jxor g01393(.dina(n1585), .dinb(n1576), .dout(n1586));
  jxor g01394(.dina(n1586), .dinb(n1561), .dout(n1587));
  jand g01395(.dina(n1431), .dinb(n1425), .dout(n1588));
  jand g01396(.dina(n1432), .dinb(n1422), .dout(n1589));
  jor  g01397(.dina(n1589), .dinb(n1588), .dout(n1590));
  jnot g01398(.din(n1482), .dout(n1591));
  jnot g01399(.din(n1485), .dout(n1592));
  jand g01400(.dina(n1592), .dinb(n1591), .dout(n1593));
  jnot g01401(.din(n1593), .dout(n1594));
  jand g01402(.dina(n1485), .dinb(n1482), .dout(n1595));
  jor  g01403(.dina(n1493), .dinb(n1595), .dout(n1596));
  jand g01404(.dina(n1596), .dinb(n1594), .dout(n1597));
  jxor g01405(.dina(n1597), .dinb(n1590), .dout(n1598));
  jnot g01406(.din(n1598), .dout(n1599));
  jor  g01407(.dina(n1469), .dinb(n1462), .dout(n1600));
  jand g01408(.dina(n1470), .dinb(n1456), .dout(n1601));
  jnot g01409(.din(n1601), .dout(n1602));
  jand g01410(.dina(n1602), .dinb(n1600), .dout(n1603));
  jxor g01411(.dina(n1603), .dinb(n1599), .dout(n1604));
  jxor g01412(.dina(n1604), .dinb(n1587), .dout(n1605));
  jxor g01413(.dina(n1605), .dinb(n1558), .dout(n1606));
  jxor g01414(.dina(n1606), .dinb(n1508), .dout(n1607));
  jand g01415(.dina(n1497), .dinb(n1412), .dout(n1608));
  jor  g01416(.dina(n1497), .dinb(n1412), .dout(n1609));
  jand g01417(.dina(n1504), .dinb(n1609), .dout(n1610));
  jor  g01418(.dina(n1610), .dinb(n1608), .dout(n1611));
  jxor g01419(.dina(n1611), .dinb(n1607), .dout(\asquared[28] ));
  jand g01420(.dina(n1528), .dinb(n1525), .dout(n1613));
  jand g01421(.dina(n1556), .dinb(n1529), .dout(n1614));
  jor  g01422(.dina(n1614), .dinb(n1613), .dout(n1615));
  jand g01423(.dina(\a[21] ), .dinb(\a[7] ), .dout(n1616));
  jand g01424(.dina(\a[23] ), .dinb(\a[5] ), .dout(n1617));
  jor  g01425(.dina(n1617), .dinb(n1245), .dout(n1618));
  jnot g01426(.din(n1618), .dout(n1619));
  jand g01427(.dina(\a[23] ), .dinb(\a[6] ), .dout(n1620));
  jand g01428(.dina(n1620), .dinb(n1541), .dout(n1621));
  jor  g01429(.dina(n1621), .dinb(n1619), .dout(n1622));
  jxor g01430(.dina(n1622), .dinb(n1616), .dout(n1623));
  jnot g01431(.din(n1623), .dout(n1624));
  jand g01432(.dina(n1531), .dinb(n1530), .dout(n1625));
  jand g01433(.dina(n1539), .dinb(n1532), .dout(n1626));
  jor  g01434(.dina(n1626), .dinb(n1625), .dout(n1627));
  jand g01435(.dina(\a[20] ), .dinb(\a[8] ), .dout(n1628));
  jnot g01436(.din(n1628), .dout(n1629));
  jand g01437(.dina(\a[25] ), .dinb(\a[3] ), .dout(n1630));
  jand g01438(.dina(\a[24] ), .dinb(\a[4] ), .dout(n1631));
  jor  g01439(.dina(n1631), .dinb(n1630), .dout(n1632));
  jand g01440(.dina(\a[25] ), .dinb(\a[4] ), .dout(n1633));
  jand g01441(.dina(n1633), .dinb(n1550), .dout(n1634));
  jnot g01442(.din(n1634), .dout(n1635));
  jand g01443(.dina(n1635), .dinb(n1632), .dout(n1636));
  jxor g01444(.dina(n1636), .dinb(n1629), .dout(n1637));
  jnot g01445(.din(n1637), .dout(n1638));
  jxor g01446(.dina(n1638), .dinb(n1627), .dout(n1639));
  jxor g01447(.dina(n1639), .dinb(n1624), .dout(n1640));
  jxor g01448(.dina(n1640), .dinb(n1615), .dout(n1641));
  jor  g01449(.dina(n1554), .dinb(n1549), .dout(n1642));
  jand g01450(.dina(n1555), .dinb(n1540), .dout(n1643));
  jnot g01451(.din(n1643), .dout(n1644));
  jand g01452(.dina(n1644), .dinb(n1642), .dout(n1645));
  jnot g01453(.din(n1645), .dout(n1646));
  jand g01454(.dina(n1574), .dinb(n1568), .dout(n1647));
  jnot g01455(.din(n1647), .dout(n1648));
  jor  g01456(.dina(n1585), .dinb(n1576), .dout(n1649));
  jand g01457(.dina(n1649), .dinb(n1648), .dout(n1650));
  jnot g01458(.din(n1650), .dout(n1651));
  jand g01459(.dina(n1544), .dinb(n1541), .dout(n1652));
  jor  g01460(.dina(n1652), .dinb(n1547), .dout(n1653));
  jand g01461(.dina(\a[27] ), .dinb(\a[1] ), .dout(n1654));
  jxor g01462(.dina(n1654), .dinb(n1546), .dout(n1655));
  jxor g01463(.dina(n1655), .dinb(n1533), .dout(n1656));
  jxor g01464(.dina(n1656), .dinb(n1653), .dout(n1657));
  jxor g01465(.dina(n1657), .dinb(n1651), .dout(n1658));
  jxor g01466(.dina(n1658), .dinb(n1646), .dout(n1659));
  jxor g01467(.dina(n1659), .dinb(n1641), .dout(n1660));
  jand g01468(.dina(n1557), .dinb(n1511), .dout(n1661));
  jand g01469(.dina(n1605), .dinb(n1558), .dout(n1662));
  jor  g01470(.dina(n1662), .dinb(n1661), .dout(n1663));
  jand g01471(.dina(n1586), .dinb(n1561), .dout(n1664));
  jand g01472(.dina(n1604), .dinb(n1587), .dout(n1665));
  jor  g01473(.dina(n1665), .dinb(n1664), .dout(n1666));
  jand g01474(.dina(n1580), .dinb(n1577), .dout(n1667));
  jor  g01475(.dina(n1667), .dinb(n1583), .dout(n1668));
  jand g01476(.dina(n1552), .dinb(n1452), .dout(n1669));
  jnot g01477(.din(n1669), .dout(n1670));
  jnot g01478(.din(n1452), .dout(n1671));
  jnot g01479(.din(n1552), .dout(n1672));
  jand g01480(.dina(n1672), .dinb(n1671), .dout(n1673));
  jor  g01481(.dina(n1673), .dinb(n1551), .dout(n1674));
  jand g01482(.dina(n1674), .dinb(n1670), .dout(n1675));
  jnot g01483(.din(n1675), .dout(n1676));
  jxor g01484(.dina(n1676), .dinb(n1668), .dout(n1677));
  jand g01485(.dina(n1567), .dinb(n1466), .dout(n1678));
  jor  g01486(.dina(n1678), .dinb(n1565), .dout(n1679));
  jxor g01487(.dina(n1679), .dinb(n1677), .dout(n1680));
  jnot g01488(.din(n1680), .dout(n1681));
  jand g01489(.dina(n1597), .dinb(n1590), .dout(n1682));
  jnot g01490(.din(n1682), .dout(n1683));
  jor  g01491(.dina(n1603), .dinb(n1599), .dout(n1684));
  jand g01492(.dina(n1684), .dinb(n1683), .dout(n1685));
  jxor g01493(.dina(n1685), .dinb(n1681), .dout(n1686));
  jand g01494(.dina(n1515), .dinb(n1513), .dout(n1687));
  jand g01495(.dina(n1524), .dinb(n1516), .dout(n1688));
  jor  g01496(.dina(n1688), .dinb(n1687), .dout(n1689));
  jand g01497(.dina(\a[26] ), .dinb(\a[2] ), .dout(n1690));
  jand g01498(.dina(\a[19] ), .dinb(\a[9] ), .dout(n1691));
  jor  g01499(.dina(n1691), .dinb(n1582), .dout(n1692));
  jnot g01500(.din(n1692), .dout(n1693));
  jand g01501(.dina(\a[19] ), .dinb(\a[10] ), .dout(n1694));
  jand g01502(.dina(n1694), .dinb(n1578), .dout(n1695));
  jor  g01503(.dina(n1695), .dinb(n1693), .dout(n1696));
  jxor g01504(.dina(n1696), .dinb(n1690), .dout(n1697));
  jand g01505(.dina(\a[17] ), .dinb(\a[11] ), .dout(n1698));
  jnot g01506(.din(n1698), .dout(n1699));
  jand g01507(.dina(\a[28] ), .dinb(\a[0] ), .dout(n1700));
  jand g01508(.dina(\a[16] ), .dinb(\a[12] ), .dout(n1701));
  jxor g01509(.dina(n1701), .dinb(n1700), .dout(n1702));
  jxor g01510(.dina(n1702), .dinb(n1699), .dout(n1703));
  jxor g01511(.dina(n1703), .dinb(n1697), .dout(n1704));
  jxor g01512(.dina(n1704), .dinb(n1689), .dout(n1705));
  jxor g01513(.dina(n1705), .dinb(n1686), .dout(n1706));
  jxor g01514(.dina(n1706), .dinb(n1666), .dout(n1707));
  jxor g01515(.dina(n1707), .dinb(n1663), .dout(n1708));
  jxor g01516(.dina(n1708), .dinb(n1660), .dout(n1709));
  jand g01517(.dina(n1606), .dinb(n1508), .dout(n1710));
  jor  g01518(.dina(n1606), .dinb(n1508), .dout(n1711));
  jand g01519(.dina(n1611), .dinb(n1711), .dout(n1712));
  jor  g01520(.dina(n1712), .dinb(n1710), .dout(n1713));
  jxor g01521(.dina(n1713), .dinb(n1709), .dout(\asquared[29] ));
  jand g01522(.dina(n1706), .dinb(n1666), .dout(n1715));
  jand g01523(.dina(n1707), .dinb(n1663), .dout(n1716));
  jor  g01524(.dina(n1716), .dinb(n1715), .dout(n1717));
  jor  g01525(.dina(n1685), .dinb(n1681), .dout(n1718));
  jand g01526(.dina(n1705), .dinb(n1686), .dout(n1719));
  jnot g01527(.din(n1719), .dout(n1720));
  jand g01528(.dina(n1720), .dinb(n1718), .dout(n1721));
  jnot g01529(.din(n1721), .dout(n1722));
  jand g01530(.dina(n1657), .dinb(n1651), .dout(n1723));
  jand g01531(.dina(n1658), .dinb(n1646), .dout(n1724));
  jor  g01532(.dina(n1724), .dinb(n1723), .dout(n1725));
  jxor g01533(.dina(n1725), .dinb(n1722), .dout(n1726));
  jor  g01534(.dina(n1703), .dinb(n1697), .dout(n1727));
  jand g01535(.dina(n1704), .dinb(n1689), .dout(n1728));
  jnot g01536(.din(n1728), .dout(n1729));
  jand g01537(.dina(n1729), .dinb(n1727), .dout(n1730));
  jnot g01538(.din(n1730), .dout(n1731));
  jand g01539(.dina(n1638), .dinb(n1627), .dout(n1732));
  jand g01540(.dina(n1639), .dinb(n1624), .dout(n1733));
  jor  g01541(.dina(n1733), .dinb(n1732), .dout(n1734));
  jxor g01542(.dina(n1734), .dinb(n1731), .dout(n1735));
  jand g01543(.dina(n1692), .dinb(n1690), .dout(n1736));
  jor  g01544(.dina(n1736), .dinb(n1695), .dout(n1737));
  jnot g01545(.din(n1737), .dout(n1738));
  jand g01546(.dina(n1701), .dinb(n1700), .dout(n1739));
  jnot g01547(.din(n1739), .dout(n1740));
  jnot g01548(.din(n1700), .dout(n1741));
  jnot g01549(.din(n1701), .dout(n1742));
  jand g01550(.dina(n1742), .dinb(n1741), .dout(n1743));
  jor  g01551(.dina(n1743), .dinb(n1699), .dout(n1744));
  jand g01552(.dina(n1744), .dinb(n1740), .dout(n1745));
  jxor g01553(.dina(n1745), .dinb(n1738), .dout(n1746));
  jand g01554(.dina(n1654), .dinb(n1546), .dout(n1747));
  jand g01555(.dina(\a[29] ), .dinb(\a[0] ), .dout(n1748));
  jand g01556(.dina(\a[27] ), .dinb(\a[2] ), .dout(n1749));
  jor  g01557(.dina(n1749), .dinb(n1748), .dout(n1750));
  jnot g01558(.din(n1750), .dout(n1751));
  jand g01559(.dina(\a[29] ), .dinb(\a[2] ), .dout(n1752));
  jand g01560(.dina(n1752), .dinb(n1531), .dout(n1753));
  jor  g01561(.dina(n1753), .dinb(n1751), .dout(n1754));
  jxor g01562(.dina(n1754), .dinb(n1747), .dout(n1755));
  jnot g01563(.din(n1755), .dout(n1756));
  jxor g01564(.dina(n1756), .dinb(n1746), .dout(n1757));
  jxor g01565(.dina(n1757), .dinb(n1735), .dout(n1758));
  jxor g01566(.dina(n1758), .dinb(n1726), .dout(n1759));
  jand g01567(.dina(n1640), .dinb(n1615), .dout(n1760));
  jand g01568(.dina(n1659), .dinb(n1641), .dout(n1761));
  jor  g01569(.dina(n1761), .dinb(n1760), .dout(n1762));
  jand g01570(.dina(n1676), .dinb(n1668), .dout(n1763));
  jand g01571(.dina(n1679), .dinb(n1677), .dout(n1764));
  jor  g01572(.dina(n1764), .dinb(n1763), .dout(n1765));
  jand g01573(.dina(n1655), .dinb(n1533), .dout(n1766));
  jand g01574(.dina(n1656), .dinb(n1653), .dout(n1767));
  jor  g01575(.dina(n1767), .dinb(n1766), .dout(n1768));
  jand g01576(.dina(\a[15] ), .dinb(\a[14] ), .dout(n1769));
  jnot g01577(.din(n1769), .dout(n1770));
  jand g01578(.dina(\a[16] ), .dinb(\a[13] ), .dout(n1771));
  jxor g01579(.dina(n1771), .dinb(n1770), .dout(n1772));
  jxor g01580(.dina(n1772), .dinb(n1620), .dout(n1773));
  jnot g01581(.din(n1773), .dout(n1774));
  jxor g01582(.dina(n1774), .dinb(n1768), .dout(n1775));
  jxor g01583(.dina(n1775), .dinb(n1765), .dout(n1776));
  jand g01584(.dina(n649), .dinb(\a[28] ), .dout(n1777));
  jnot g01585(.din(n1777), .dout(n1778));
  jand g01586(.dina(\a[28] ), .dinb(\a[1] ), .dout(n1779));
  jor  g01587(.dina(n1779), .dinb(\a[15] ), .dout(n1780));
  jand g01588(.dina(n1780), .dinb(n1778), .dout(n1781));
  jand g01589(.dina(n1618), .dinb(n1616), .dout(n1782));
  jor  g01590(.dina(n1782), .dinb(n1621), .dout(n1783));
  jxor g01591(.dina(n1783), .dinb(n1781), .dout(n1784));
  jand g01592(.dina(n1635), .dinb(n1629), .dout(n1785));
  jnot g01593(.din(n1785), .dout(n1786));
  jand g01594(.dina(n1786), .dinb(n1632), .dout(n1787));
  jxor g01595(.dina(n1787), .dinb(n1784), .dout(n1788));
  jand g01596(.dina(\a[22] ), .dinb(\a[7] ), .dout(n1789));
  jand g01597(.dina(\a[24] ), .dinb(\a[5] ), .dout(n1790));
  jor  g01598(.dina(n1790), .dinb(n1789), .dout(n1791));
  jnot g01599(.din(n1791), .dout(n1792));
  jand g01600(.dina(\a[24] ), .dinb(\a[7] ), .dout(n1793));
  jand g01601(.dina(n1793), .dinb(n1541), .dout(n1794));
  jor  g01602(.dina(n1794), .dinb(n1792), .dout(n1795));
  jxor g01603(.dina(n1795), .dinb(n1633), .dout(n1796));
  jand g01604(.dina(\a[20] ), .dinb(\a[9] ), .dout(n1797));
  jand g01605(.dina(\a[18] ), .dinb(\a[11] ), .dout(n1798));
  jor  g01606(.dina(n1798), .dinb(n1694), .dout(n1799));
  jnot g01607(.din(n1799), .dout(n1800));
  jand g01608(.dina(\a[19] ), .dinb(\a[11] ), .dout(n1801));
  jand g01609(.dina(n1801), .dinb(n1582), .dout(n1802));
  jor  g01610(.dina(n1802), .dinb(n1800), .dout(n1803));
  jxor g01611(.dina(n1803), .dinb(n1797), .dout(n1804));
  jand g01612(.dina(\a[17] ), .dinb(\a[12] ), .dout(n1805));
  jand g01613(.dina(\a[26] ), .dinb(\a[3] ), .dout(n1806));
  jand g01614(.dina(\a[21] ), .dinb(\a[8] ), .dout(n1807));
  jor  g01615(.dina(n1807), .dinb(n1806), .dout(n1808));
  jand g01616(.dina(\a[26] ), .dinb(\a[8] ), .dout(n1809));
  jand g01617(.dina(n1809), .dinb(n1259), .dout(n1810));
  jnot g01618(.din(n1810), .dout(n1811));
  jand g01619(.dina(n1811), .dinb(n1808), .dout(n1812));
  jxor g01620(.dina(n1812), .dinb(n1805), .dout(n1813));
  jxor g01621(.dina(n1813), .dinb(n1804), .dout(n1814));
  jxor g01622(.dina(n1814), .dinb(n1796), .dout(n1815));
  jxor g01623(.dina(n1815), .dinb(n1788), .dout(n1816));
  jxor g01624(.dina(n1816), .dinb(n1776), .dout(n1817));
  jxor g01625(.dina(n1817), .dinb(n1762), .dout(n1818));
  jxor g01626(.dina(n1818), .dinb(n1759), .dout(n1819));
  jxor g01627(.dina(n1819), .dinb(n1717), .dout(n1820));
  jand g01628(.dina(n1708), .dinb(n1660), .dout(n1821));
  jnot g01629(.din(n1660), .dout(n1822));
  jnot g01630(.din(n1708), .dout(n1823));
  jand g01631(.dina(n1823), .dinb(n1822), .dout(n1824));
  jnot g01632(.din(n1824), .dout(n1825));
  jand g01633(.dina(n1713), .dinb(n1825), .dout(n1826));
  jor  g01634(.dina(n1826), .dinb(n1821), .dout(n1827));
  jxor g01635(.dina(n1827), .dinb(n1820), .dout(\asquared[30] ));
  jand g01636(.dina(n1817), .dinb(n1762), .dout(n1829));
  jand g01637(.dina(n1818), .dinb(n1759), .dout(n1830));
  jor  g01638(.dina(n1830), .dinb(n1829), .dout(n1831));
  jand g01639(.dina(n1783), .dinb(n1781), .dout(n1832));
  jand g01640(.dina(n1787), .dinb(n1784), .dout(n1833));
  jor  g01641(.dina(n1833), .dinb(n1832), .dout(n1834));
  jnot g01642(.din(n1834), .dout(n1835));
  jand g01643(.dina(\a[30] ), .dinb(\a[0] ), .dout(n1836));
  jxor g01644(.dina(n1836), .dinb(n1777), .dout(n1837));
  jand g01645(.dina(\a[16] ), .dinb(\a[14] ), .dout(n1838));
  jand g01646(.dina(\a[29] ), .dinb(\a[1] ), .dout(n1839));
  jxor g01647(.dina(n1839), .dinb(n1838), .dout(n1840));
  jnot g01648(.din(n1840), .dout(n1841));
  jxor g01649(.dina(n1841), .dinb(n1837), .dout(n1842));
  jxor g01650(.dina(n1842), .dinb(n1835), .dout(n1843));
  jand g01651(.dina(n1745), .dinb(n1738), .dout(n1844));
  jnot g01652(.din(n1844), .dout(n1845));
  jnot g01653(.din(n1745), .dout(n1846));
  jand g01654(.dina(n1846), .dinb(n1737), .dout(n1847));
  jor  g01655(.dina(n1756), .dinb(n1847), .dout(n1848));
  jand g01656(.dina(n1848), .dinb(n1845), .dout(n1849));
  jxor g01657(.dina(n1849), .dinb(n1843), .dout(n1850));
  jand g01658(.dina(n1815), .dinb(n1788), .dout(n1851));
  jand g01659(.dina(n1816), .dinb(n1776), .dout(n1852));
  jor  g01660(.dina(n1852), .dinb(n1851), .dout(n1853));
  jxor g01661(.dina(n1853), .dinb(n1850), .dout(n1854));
  jand g01662(.dina(n1791), .dinb(n1633), .dout(n1855));
  jor  g01663(.dina(n1855), .dinb(n1794), .dout(n1856));
  jnot g01664(.din(n1771), .dout(n1857));
  jand g01665(.dina(n1857), .dinb(n1770), .dout(n1858));
  jnot g01666(.din(n1858), .dout(n1859));
  jand g01667(.dina(n1771), .dinb(n1769), .dout(n1860));
  jor  g01668(.dina(n1860), .dinb(n1620), .dout(n1861));
  jand g01669(.dina(n1861), .dinb(n1859), .dout(n1862));
  jxor g01670(.dina(n1862), .dinb(n1856), .dout(n1863));
  jand g01671(.dina(\a[17] ), .dinb(\a[13] ), .dout(n1864));
  jand g01672(.dina(\a[28] ), .dinb(\a[2] ), .dout(n1865));
  jnot g01673(.din(n1865), .dout(n1866));
  jand g01674(.dina(\a[21] ), .dinb(\a[9] ), .dout(n1867));
  jxor g01675(.dina(n1867), .dinb(n1866), .dout(n1868));
  jxor g01676(.dina(n1868), .dinb(n1864), .dout(n1869));
  jnot g01677(.din(n1869), .dout(n1870));
  jxor g01678(.dina(n1870), .dinb(n1863), .dout(n1871));
  jnot g01679(.din(n1804), .dout(n1872));
  jor  g01680(.dina(n1813), .dinb(n1872), .dout(n1873));
  jnot g01681(.din(n1796), .dout(n1874));
  jand g01682(.dina(n1813), .dinb(n1872), .dout(n1875));
  jor  g01683(.dina(n1875), .dinb(n1874), .dout(n1876));
  jand g01684(.dina(n1876), .dinb(n1873), .dout(n1877));
  jxor g01685(.dina(n1877), .dinb(n1871), .dout(n1878));
  jand g01686(.dina(n1812), .dinb(n1805), .dout(n1879));
  jor  g01687(.dina(n1879), .dinb(n1810), .dout(n1880));
  jand g01688(.dina(n1799), .dinb(n1797), .dout(n1881));
  jor  g01689(.dina(n1881), .dinb(n1802), .dout(n1882));
  jxor g01690(.dina(n1882), .dinb(n1880), .dout(n1883));
  jand g01691(.dina(n1750), .dinb(n1747), .dout(n1884));
  jor  g01692(.dina(n1884), .dinb(n1753), .dout(n1885));
  jxor g01693(.dina(n1885), .dinb(n1883), .dout(n1886));
  jxor g01694(.dina(n1886), .dinb(n1878), .dout(n1887));
  jxor g01695(.dina(n1887), .dinb(n1854), .dout(n1888));
  jand g01696(.dina(n1725), .dinb(n1722), .dout(n1889));
  jand g01697(.dina(n1758), .dinb(n1726), .dout(n1890));
  jor  g01698(.dina(n1890), .dinb(n1889), .dout(n1891));
  jand g01699(.dina(n1774), .dinb(n1768), .dout(n1892));
  jand g01700(.dina(n1775), .dinb(n1765), .dout(n1893));
  jor  g01701(.dina(n1893), .dinb(n1892), .dout(n1894));
  jand g01702(.dina(\a[20] ), .dinb(\a[10] ), .dout(n1895));
  jnot g01703(.din(n1895), .dout(n1896));
  jand g01704(.dina(\a[18] ), .dinb(\a[12] ), .dout(n1897));
  jor  g01705(.dina(n1897), .dinb(n1801), .dout(n1898));
  jand g01706(.dina(\a[19] ), .dinb(\a[12] ), .dout(n1899));
  jand g01707(.dina(n1899), .dinb(n1798), .dout(n1900));
  jnot g01708(.din(n1900), .dout(n1901));
  jand g01709(.dina(n1901), .dinb(n1898), .dout(n1902));
  jxor g01710(.dina(n1902), .dinb(n1896), .dout(n1903));
  jand g01711(.dina(\a[25] ), .dinb(\a[5] ), .dout(n1904));
  jnot g01712(.din(n1904), .dout(n1905));
  jand g01713(.dina(\a[23] ), .dinb(\a[7] ), .dout(n1906));
  jand g01714(.dina(\a[24] ), .dinb(\a[6] ), .dout(n1907));
  jor  g01715(.dina(n1907), .dinb(n1906), .dout(n1908));
  jand g01716(.dina(n1793), .dinb(n1620), .dout(n1909));
  jnot g01717(.din(n1909), .dout(n1910));
  jand g01718(.dina(n1910), .dinb(n1908), .dout(n1911));
  jxor g01719(.dina(n1911), .dinb(n1905), .dout(n1912));
  jand g01720(.dina(\a[27] ), .dinb(\a[3] ), .dout(n1913));
  jnot g01721(.din(n1913), .dout(n1914));
  jand g01722(.dina(\a[26] ), .dinb(\a[4] ), .dout(n1915));
  jand g01723(.dina(\a[22] ), .dinb(\a[8] ), .dout(n1916));
  jxor g01724(.dina(n1916), .dinb(n1915), .dout(n1917));
  jxor g01725(.dina(n1917), .dinb(n1914), .dout(n1918));
  jnot g01726(.din(n1918), .dout(n1919));
  jxor g01727(.dina(n1919), .dinb(n1912), .dout(n1920));
  jxor g01728(.dina(n1920), .dinb(n1903), .dout(n1921));
  jxor g01729(.dina(n1921), .dinb(n1894), .dout(n1922));
  jand g01730(.dina(n1734), .dinb(n1731), .dout(n1923));
  jand g01731(.dina(n1757), .dinb(n1735), .dout(n1924));
  jor  g01732(.dina(n1924), .dinb(n1923), .dout(n1925));
  jxor g01733(.dina(n1925), .dinb(n1922), .dout(n1926));
  jxor g01734(.dina(n1926), .dinb(n1891), .dout(n1927));
  jxor g01735(.dina(n1927), .dinb(n1888), .dout(n1928));
  jxor g01736(.dina(n1928), .dinb(n1831), .dout(n1929));
  jand g01737(.dina(n1819), .dinb(n1717), .dout(n1930));
  jor  g01738(.dina(n1819), .dinb(n1717), .dout(n1931));
  jand g01739(.dina(n1827), .dinb(n1931), .dout(n1932));
  jor  g01740(.dina(n1932), .dinb(n1930), .dout(n1933));
  jxor g01741(.dina(n1933), .dinb(n1929), .dout(\asquared[31] ));
  jand g01742(.dina(n1926), .dinb(n1891), .dout(n1935));
  jand g01743(.dina(n1927), .dinb(n1888), .dout(n1936));
  jor  g01744(.dina(n1936), .dinb(n1935), .dout(n1937));
  jand g01745(.dina(n1853), .dinb(n1850), .dout(n1938));
  jand g01746(.dina(n1887), .dinb(n1854), .dout(n1939));
  jor  g01747(.dina(n1939), .dinb(n1938), .dout(n1940));
  jand g01748(.dina(n1877), .dinb(n1871), .dout(n1941));
  jand g01749(.dina(n1886), .dinb(n1878), .dout(n1942));
  jor  g01750(.dina(n1942), .dinb(n1941), .dout(n1943));
  jand g01751(.dina(\a[20] ), .dinb(\a[11] ), .dout(n1944));
  jnot g01752(.din(n1944), .dout(n1945));
  jand g01753(.dina(\a[18] ), .dinb(\a[13] ), .dout(n1946));
  jor  g01754(.dina(n1946), .dinb(n1899), .dout(n1947));
  jand g01755(.dina(\a[19] ), .dinb(\a[13] ), .dout(n1948));
  jand g01756(.dina(n1948), .dinb(n1897), .dout(n1949));
  jnot g01757(.din(n1949), .dout(n1950));
  jand g01758(.dina(n1950), .dinb(n1947), .dout(n1951));
  jxor g01759(.dina(n1951), .dinb(n1945), .dout(n1952));
  jand g01760(.dina(n1836), .dinb(n1777), .dout(n1953));
  jnot g01761(.din(n1953), .dout(n1954));
  jnot g01762(.din(n1836), .dout(n1955));
  jand g01763(.dina(n1955), .dinb(n1778), .dout(n1956));
  jor  g01764(.dina(n1841), .dinb(n1956), .dout(n1957));
  jand g01765(.dina(n1957), .dinb(n1954), .dout(n1958));
  jxor g01766(.dina(n1958), .dinb(n1952), .dout(n1959));
  jand g01767(.dina(\a[21] ), .dinb(\a[10] ), .dout(n1960));
  jand g01768(.dina(\a[31] ), .dinb(\a[0] ), .dout(n1961));
  jand g01769(.dina(\a[22] ), .dinb(\a[9] ), .dout(n1962));
  jor  g01770(.dina(n1962), .dinb(n1961), .dout(n1963));
  jand g01771(.dina(\a[31] ), .dinb(\a[9] ), .dout(n1964));
  jand g01772(.dina(n1964), .dinb(n1081), .dout(n1965));
  jnot g01773(.din(n1965), .dout(n1966));
  jand g01774(.dina(n1966), .dinb(n1963), .dout(n1967));
  jxor g01775(.dina(n1967), .dinb(n1960), .dout(n1968));
  jxor g01776(.dina(n1968), .dinb(n1959), .dout(n1969));
  jand g01777(.dina(\a[28] ), .dinb(\a[3] ), .dout(n1970));
  jand g01778(.dina(\a[27] ), .dinb(\a[4] ), .dout(n1971));
  jor  g01779(.dina(n1971), .dinb(n1970), .dout(n1972));
  jnot g01780(.din(n1972), .dout(n1973));
  jand g01781(.dina(\a[28] ), .dinb(\a[4] ), .dout(n1974));
  jand g01782(.dina(n1974), .dinb(n1913), .dout(n1975));
  jor  g01783(.dina(n1975), .dinb(n1973), .dout(n1976));
  jxor g01784(.dina(n1976), .dinb(n1752), .dout(n1977));
  jand g01785(.dina(\a[25] ), .dinb(\a[6] ), .dout(n1978));
  jand g01786(.dina(\a[16] ), .dinb(\a[15] ), .dout(n1979));
  jand g01787(.dina(\a[17] ), .dinb(\a[14] ), .dout(n1980));
  jor  g01788(.dina(n1980), .dinb(n1979), .dout(n1981));
  jnot g01789(.din(n1981), .dout(n1982));
  jand g01790(.dina(\a[17] ), .dinb(\a[15] ), .dout(n1983));
  jand g01791(.dina(n1983), .dinb(n1838), .dout(n1984));
  jor  g01792(.dina(n1984), .dinb(n1982), .dout(n1985));
  jxor g01793(.dina(n1985), .dinb(n1978), .dout(n1986));
  jand g01794(.dina(\a[23] ), .dinb(\a[8] ), .dout(n1987));
  jand g01795(.dina(\a[26] ), .dinb(\a[5] ), .dout(n1988));
  jor  g01796(.dina(n1988), .dinb(n1793), .dout(n1989));
  jand g01797(.dina(\a[26] ), .dinb(\a[7] ), .dout(n1990));
  jand g01798(.dina(n1990), .dinb(n1790), .dout(n1991));
  jnot g01799(.din(n1991), .dout(n1992));
  jand g01800(.dina(n1992), .dinb(n1989), .dout(n1993));
  jxor g01801(.dina(n1993), .dinb(n1987), .dout(n1994));
  jxor g01802(.dina(n1994), .dinb(n1986), .dout(n1995));
  jxor g01803(.dina(n1995), .dinb(n1977), .dout(n1996));
  jxor g01804(.dina(n1996), .dinb(n1969), .dout(n1997));
  jxor g01805(.dina(n1997), .dinb(n1943), .dout(n1998));
  jxor g01806(.dina(n1998), .dinb(n1940), .dout(n1999));
  jand g01807(.dina(n1921), .dinb(n1894), .dout(n2000));
  jand g01808(.dina(n1925), .dinb(n1922), .dout(n2001));
  jor  g01809(.dina(n2001), .dinb(n2000), .dout(n2002));
  jand g01810(.dina(n1882), .dinb(n1880), .dout(n2003));
  jand g01811(.dina(n1885), .dinb(n1883), .dout(n2004));
  jor  g01812(.dina(n2004), .dinb(n2003), .dout(n2005));
  jnot g01813(.din(n1856), .dout(n2006));
  jnot g01814(.din(n1862), .dout(n2007));
  jand g01815(.dina(n2007), .dinb(n2006), .dout(n2008));
  jnot g01816(.din(n2008), .dout(n2009));
  jand g01817(.dina(n1862), .dinb(n1856), .dout(n2010));
  jor  g01818(.dina(n1870), .dinb(n2010), .dout(n2011));
  jand g01819(.dina(n2011), .dinb(n2009), .dout(n2012));
  jxor g01820(.dina(n2012), .dinb(n2005), .dout(n2013));
  jand g01821(.dina(n1908), .dinb(n1904), .dout(n2014));
  jor  g01822(.dina(n2014), .dinb(n1909), .dout(n2015));
  jand g01823(.dina(\a[30] ), .dinb(\a[1] ), .dout(n2016));
  jnot g01824(.din(\a[16] ), .dout(n2017));
  jand g01825(.dina(n1839), .dinb(n1838), .dout(n2018));
  jor  g01826(.dina(n2018), .dinb(n2017), .dout(n2019));
  jxor g01827(.dina(n2019), .dinb(n2016), .dout(n2020));
  jnot g01828(.din(n2020), .dout(n2021));
  jxor g01829(.dina(n2021), .dinb(n2015), .dout(n2022));
  jxor g01830(.dina(n2022), .dinb(n2013), .dout(n2023));
  jxor g01831(.dina(n2023), .dinb(n2002), .dout(n2024));
  jnot g01832(.din(n1867), .dout(n2025));
  jand g01833(.dina(n2025), .dinb(n1866), .dout(n2026));
  jnot g01834(.din(n2026), .dout(n2027));
  jand g01835(.dina(n1867), .dinb(n1865), .dout(n2028));
  jor  g01836(.dina(n2028), .dinb(n1864), .dout(n2029));
  jand g01837(.dina(n2029), .dinb(n2027), .dout(n2030));
  jnot g01838(.din(n1915), .dout(n2031));
  jnot g01839(.din(n1916), .dout(n2032));
  jand g01840(.dina(n2032), .dinb(n2031), .dout(n2033));
  jnot g01841(.din(n2033), .dout(n2034));
  jand g01842(.dina(n1916), .dinb(n1915), .dout(n2035));
  jor  g01843(.dina(n2035), .dinb(n1913), .dout(n2036));
  jand g01844(.dina(n2036), .dinb(n2034), .dout(n2037));
  jxor g01845(.dina(n2037), .dinb(n2030), .dout(n2038));
  jand g01846(.dina(n1898), .dinb(n1895), .dout(n2039));
  jor  g01847(.dina(n2039), .dinb(n1900), .dout(n2040));
  jxor g01848(.dina(n2040), .dinb(n2038), .dout(n2041));
  jnot g01849(.din(n2041), .dout(n2042));
  jnot g01850(.din(n1912), .dout(n2043));
  jand g01851(.dina(n1919), .dinb(n2043), .dout(n2044));
  jnot g01852(.din(n2044), .dout(n2045));
  jand g01853(.dina(n1918), .dinb(n1912), .dout(n2046));
  jor  g01854(.dina(n2046), .dinb(n1903), .dout(n2047));
  jand g01855(.dina(n2047), .dinb(n2045), .dout(n2048));
  jxor g01856(.dina(n2048), .dinb(n2042), .dout(n2049));
  jnot g01857(.din(n2049), .dout(n2050));
  jor  g01858(.dina(n1842), .dinb(n1835), .dout(n2051));
  jand g01859(.dina(n1849), .dinb(n1843), .dout(n2052));
  jnot g01860(.din(n2052), .dout(n2053));
  jand g01861(.dina(n2053), .dinb(n2051), .dout(n2054));
  jxor g01862(.dina(n2054), .dinb(n2050), .dout(n2055));
  jxor g01863(.dina(n2055), .dinb(n2024), .dout(n2056));
  jxor g01864(.dina(n2056), .dinb(n1999), .dout(n2057));
  jxor g01865(.dina(n2057), .dinb(n1937), .dout(n2058));
  jand g01866(.dina(n1928), .dinb(n1831), .dout(n2059));
  jor  g01867(.dina(n1928), .dinb(n1831), .dout(n2060));
  jand g01868(.dina(n1933), .dinb(n2060), .dout(n2061));
  jor  g01869(.dina(n2061), .dinb(n2059), .dout(n2062));
  jxor g01870(.dina(n2062), .dinb(n2058), .dout(\asquared[32] ));
  jand g01871(.dina(n1998), .dinb(n1940), .dout(n2064));
  jand g01872(.dina(n2056), .dinb(n1999), .dout(n2065));
  jor  g01873(.dina(n2065), .dinb(n2064), .dout(n2066));
  jand g01874(.dina(n2023), .dinb(n2002), .dout(n2067));
  jand g01875(.dina(n2055), .dinb(n2024), .dout(n2068));
  jor  g01876(.dina(n2068), .dinb(n2067), .dout(n2069));
  jor  g01877(.dina(n2048), .dinb(n2042), .dout(n2070));
  jor  g01878(.dina(n2054), .dinb(n2050), .dout(n2071));
  jand g01879(.dina(n2071), .dinb(n2070), .dout(n2072));
  jnot g01880(.din(n2072), .dout(n2073));
  jand g01881(.dina(n2021), .dinb(n2015), .dout(n2074));
  jnot g01882(.din(\a[30] ), .dout(n2075));
  jand g01883(.dina(n2018), .dinb(n2075), .dout(n2076));
  jor  g01884(.dina(n2076), .dinb(n2074), .dout(n2077));
  jand g01885(.dina(\a[24] ), .dinb(\a[8] ), .dout(n2078));
  jand g01886(.dina(\a[26] ), .dinb(\a[6] ), .dout(n2079));
  jor  g01887(.dina(n2079), .dinb(n1564), .dout(n2080));
  jnot g01888(.din(n2080), .dout(n2081));
  jand g01889(.dina(n1990), .dinb(n1978), .dout(n2082));
  jor  g01890(.dina(n2082), .dinb(n2081), .dout(n2083));
  jxor g01891(.dina(n2083), .dinb(n2078), .dout(n2084));
  jnot g01892(.din(n2084), .dout(n2085));
  jand g01893(.dina(\a[23] ), .dinb(\a[9] ), .dout(n2086));
  jnot g01894(.din(n1974), .dout(n2087));
  jand g01895(.dina(\a[27] ), .dinb(\a[5] ), .dout(n2088));
  jnot g01896(.din(n2088), .dout(n2089));
  jand g01897(.dina(n2089), .dinb(n2087), .dout(n2090));
  jand g01898(.dina(\a[28] ), .dinb(\a[5] ), .dout(n2091));
  jand g01899(.dina(n2091), .dinb(n1971), .dout(n2092));
  jor  g01900(.dina(n2092), .dinb(n2090), .dout(n2093));
  jnot g01901(.din(n2093), .dout(n2094));
  jxor g01902(.dina(n2094), .dinb(n2086), .dout(n2095));
  jxor g01903(.dina(n2095), .dinb(n2085), .dout(n2096));
  jxor g01904(.dina(n2096), .dinb(n2077), .dout(n2097));
  jand g01905(.dina(\a[21] ), .dinb(\a[11] ), .dout(n2098));
  jnot g01906(.din(n2098), .dout(n2099));
  jand g01907(.dina(\a[20] ), .dinb(\a[12] ), .dout(n2100));
  jor  g01908(.dina(n2100), .dinb(n1948), .dout(n2101));
  jand g01909(.dina(\a[20] ), .dinb(\a[13] ), .dout(n2102));
  jand g01910(.dina(n2102), .dinb(n1899), .dout(n2103));
  jnot g01911(.din(n2103), .dout(n2104));
  jand g01912(.dina(n2104), .dinb(n2101), .dout(n2105));
  jxor g01913(.dina(n2105), .dinb(n2099), .dout(n2106));
  jand g01914(.dina(n2016), .dinb(\a[16] ), .dout(n2107));
  jnot g01915(.din(n2107), .dout(n2108));
  jand g01916(.dina(\a[32] ), .dinb(\a[0] ), .dout(n2109));
  jand g01917(.dina(\a[30] ), .dinb(\a[2] ), .dout(n2110));
  jor  g01918(.dina(n2110), .dinb(n2109), .dout(n2111));
  jand g01919(.dina(\a[32] ), .dinb(\a[2] ), .dout(n2112));
  jand g01920(.dina(n2112), .dinb(n1836), .dout(n2113));
  jnot g01921(.din(n2113), .dout(n2114));
  jand g01922(.dina(n2114), .dinb(n2111), .dout(n2115));
  jxor g01923(.dina(n2115), .dinb(n2108), .dout(n2116));
  jxor g01924(.dina(n2116), .dinb(n2106), .dout(n2117));
  jand g01925(.dina(\a[18] ), .dinb(\a[14] ), .dout(n2118));
  jand g01926(.dina(\a[29] ), .dinb(\a[3] ), .dout(n2119));
  jnot g01927(.din(n2119), .dout(n2120));
  jand g01928(.dina(\a[22] ), .dinb(\a[10] ), .dout(n2121));
  jxor g01929(.dina(n2121), .dinb(n2120), .dout(n2122));
  jxor g01930(.dina(n2122), .dinb(n2118), .dout(n2123));
  jnot g01931(.din(n2123), .dout(n2124));
  jxor g01932(.dina(n2124), .dinb(n2117), .dout(n2125));
  jxor g01933(.dina(n2125), .dinb(n2097), .dout(n2126));
  jxor g01934(.dina(n2126), .dinb(n2073), .dout(n2127));
  jxor g01935(.dina(n2127), .dinb(n2069), .dout(n2128));
  jand g01936(.dina(n2012), .dinb(n2005), .dout(n2129));
  jand g01937(.dina(n2022), .dinb(n2013), .dout(n2130));
  jor  g01938(.dina(n2130), .dinb(n2129), .dout(n2131));
  jand g01939(.dina(n1967), .dinb(n1960), .dout(n2132));
  jor  g01940(.dina(n2132), .dinb(n1965), .dout(n2133));
  jand g01941(.dina(n1947), .dinb(n1944), .dout(n2134));
  jor  g01942(.dina(n2134), .dinb(n1949), .dout(n2135));
  jxor g01943(.dina(n2135), .dinb(n2133), .dout(n2136));
  jand g01944(.dina(n1972), .dinb(n1752), .dout(n2137));
  jor  g01945(.dina(n2137), .dinb(n1975), .dout(n2138));
  jxor g01946(.dina(n2138), .dinb(n2136), .dout(n2139));
  jand g01947(.dina(n1993), .dinb(n1987), .dout(n2140));
  jor  g01948(.dina(n2140), .dinb(n1991), .dout(n2141));
  jand g01949(.dina(\a[31] ), .dinb(\a[1] ), .dout(n2142));
  jxor g01950(.dina(n2142), .dinb(n1983), .dout(n2143));
  jand g01951(.dina(n1981), .dinb(n1978), .dout(n2144));
  jor  g01952(.dina(n2144), .dinb(n1984), .dout(n2145));
  jxor g01953(.dina(n2145), .dinb(n2143), .dout(n2146));
  jxor g01954(.dina(n2146), .dinb(n2141), .dout(n2147));
  jxor g01955(.dina(n2147), .dinb(n2139), .dout(n2148));
  jxor g01956(.dina(n2148), .dinb(n2131), .dout(n2149));
  jnot g01957(.din(n1952), .dout(n2150));
  jnot g01958(.din(n1958), .dout(n2151));
  jand g01959(.dina(n2151), .dinb(n2150), .dout(n2152));
  jand g01960(.dina(n1968), .dinb(n1959), .dout(n2153));
  jor  g01961(.dina(n2153), .dinb(n2152), .dout(n2154));
  jand g01962(.dina(n2037), .dinb(n2030), .dout(n2155));
  jand g01963(.dina(n2040), .dinb(n2038), .dout(n2156));
  jor  g01964(.dina(n2156), .dinb(n2155), .dout(n2157));
  jxor g01965(.dina(n2157), .dinb(n2154), .dout(n2158));
  jnot g01966(.din(n1986), .dout(n2159));
  jor  g01967(.dina(n1994), .dinb(n2159), .dout(n2160));
  jnot g01968(.din(n1977), .dout(n2161));
  jand g01969(.dina(n1994), .dinb(n2159), .dout(n2162));
  jor  g01970(.dina(n2162), .dinb(n2161), .dout(n2163));
  jand g01971(.dina(n2163), .dinb(n2160), .dout(n2164));
  jxor g01972(.dina(n2164), .dinb(n2158), .dout(n2165));
  jand g01973(.dina(n1996), .dinb(n1969), .dout(n2166));
  jand g01974(.dina(n1997), .dinb(n1943), .dout(n2167));
  jor  g01975(.dina(n2167), .dinb(n2166), .dout(n2168));
  jxor g01976(.dina(n2168), .dinb(n2165), .dout(n2169));
  jxor g01977(.dina(n2169), .dinb(n2149), .dout(n2170));
  jxor g01978(.dina(n2170), .dinb(n2128), .dout(n2171));
  jxor g01979(.dina(n2171), .dinb(n2066), .dout(n2172));
  jand g01980(.dina(n2057), .dinb(n1937), .dout(n2173));
  jor  g01981(.dina(n2057), .dinb(n1937), .dout(n2174));
  jand g01982(.dina(n2062), .dinb(n2174), .dout(n2175));
  jor  g01983(.dina(n2175), .dinb(n2173), .dout(n2176));
  jxor g01984(.dina(n2176), .dinb(n2172), .dout(\asquared[33] ));
  jand g01985(.dina(n2135), .dinb(n2133), .dout(n2178));
  jand g01986(.dina(n2138), .dinb(n2136), .dout(n2179));
  jor  g01987(.dina(n2179), .dinb(n2178), .dout(n2180));
  jand g01988(.dina(n2116), .dinb(n2106), .dout(n2181));
  jnot g01989(.din(n2181), .dout(n2182));
  jnot g01990(.din(n2106), .dout(n2183));
  jnot g01991(.din(n2116), .dout(n2184));
  jand g01992(.dina(n2184), .dinb(n2183), .dout(n2185));
  jor  g01993(.dina(n2124), .dinb(n2185), .dout(n2186));
  jand g01994(.dina(n2186), .dinb(n2182), .dout(n2187));
  jxor g01995(.dina(n2187), .dinb(n2180), .dout(n2188));
  jand g01996(.dina(n2095), .dinb(n2085), .dout(n2189));
  jand g01997(.dina(n2096), .dinb(n2077), .dout(n2190));
  jor  g01998(.dina(n2190), .dinb(n2189), .dout(n2191));
  jxor g01999(.dina(n2191), .dinb(n2188), .dout(n2192));
  jand g02000(.dina(n2125), .dinb(n2097), .dout(n2193));
  jand g02001(.dina(n2126), .dinb(n2073), .dout(n2194));
  jor  g02002(.dina(n2194), .dinb(n2193), .dout(n2195));
  jxor g02003(.dina(n2195), .dinb(n2192), .dout(n2196));
  jand g02004(.dina(n2111), .dinb(n2107), .dout(n2197));
  jor  g02005(.dina(n2197), .dinb(n2113), .dout(n2198));
  jand g02006(.dina(n2101), .dinb(n2098), .dout(n2199));
  jor  g02007(.dina(n2199), .dinb(n2103), .dout(n2200));
  jxor g02008(.dina(n2200), .dinb(n2198), .dout(n2201));
  jnot g02009(.din(n2121), .dout(n2202));
  jand g02010(.dina(n2202), .dinb(n2120), .dout(n2203));
  jnot g02011(.din(n2203), .dout(n2204));
  jand g02012(.dina(n2121), .dinb(n2119), .dout(n2205));
  jor  g02013(.dina(n2205), .dinb(n2118), .dout(n2206));
  jand g02014(.dina(n2206), .dinb(n2204), .dout(n2207));
  jxor g02015(.dina(n2207), .dinb(n2201), .dout(n2208));
  jand g02016(.dina(n2094), .dinb(n2086), .dout(n2209));
  jor  g02017(.dina(n2209), .dinb(n2092), .dout(n2210));
  jand g02018(.dina(n2080), .dinb(n2078), .dout(n2211));
  jor  g02019(.dina(n2211), .dinb(n2082), .dout(n2212));
  jxor g02020(.dina(n2212), .dinb(n2210), .dout(n2213));
  jand g02021(.dina(\a[31] ), .dinb(\a[2] ), .dout(n2214));
  jand g02022(.dina(\a[33] ), .dinb(\a[0] ), .dout(n2215));
  jnot g02023(.din(n2215), .dout(n2216));
  jand g02024(.dina(\a[22] ), .dinb(\a[11] ), .dout(n2217));
  jnot g02025(.din(n2217), .dout(n2218));
  jand g02026(.dina(n2218), .dinb(n2216), .dout(n2219));
  jand g02027(.dina(\a[33] ), .dinb(\a[11] ), .dout(n2220));
  jand g02028(.dina(n2220), .dinb(n1081), .dout(n2221));
  jor  g02029(.dina(n2221), .dinb(n2219), .dout(n2222));
  jxor g02030(.dina(n2222), .dinb(n2214), .dout(n2223));
  jnot g02031(.din(n2223), .dout(n2224));
  jxor g02032(.dina(n2224), .dinb(n2213), .dout(n2225));
  jxor g02033(.dina(n2225), .dinb(n2208), .dout(n2226));
  jnot g02034(.din(n1990), .dout(n2227));
  jand g02035(.dina(\a[17] ), .dinb(\a[16] ), .dout(n2228));
  jand g02036(.dina(\a[18] ), .dinb(\a[15] ), .dout(n2229));
  jor  g02037(.dina(n2229), .dinb(n2228), .dout(n2230));
  jand g02038(.dina(\a[18] ), .dinb(\a[16] ), .dout(n2231));
  jand g02039(.dina(n2231), .dinb(n1983), .dout(n2232));
  jnot g02040(.din(n2232), .dout(n2233));
  jand g02041(.dina(n2233), .dinb(n2230), .dout(n2234));
  jxor g02042(.dina(n2234), .dinb(n2227), .dout(n2235));
  jnot g02043(.din(n2091), .dout(n2236));
  jand g02044(.dina(\a[25] ), .dinb(\a[8] ), .dout(n2237));
  jand g02045(.dina(\a[27] ), .dinb(\a[6] ), .dout(n2238));
  jor  g02046(.dina(n2238), .dinb(n2237), .dout(n2239));
  jand g02047(.dina(\a[27] ), .dinb(\a[8] ), .dout(n2240));
  jand g02048(.dina(n2240), .dinb(n1978), .dout(n2241));
  jnot g02049(.din(n2241), .dout(n2242));
  jand g02050(.dina(n2242), .dinb(n2239), .dout(n2243));
  jxor g02051(.dina(n2243), .dinb(n2236), .dout(n2244));
  jand g02052(.dina(\a[30] ), .dinb(\a[3] ), .dout(n2245));
  jnot g02053(.din(n2245), .dout(n2246));
  jand g02054(.dina(\a[29] ), .dinb(\a[4] ), .dout(n2247));
  jand g02055(.dina(\a[24] ), .dinb(\a[9] ), .dout(n2248));
  jxor g02056(.dina(n2248), .dinb(n2247), .dout(n2249));
  jxor g02057(.dina(n2249), .dinb(n2246), .dout(n2250));
  jnot g02058(.din(n2250), .dout(n2251));
  jxor g02059(.dina(n2251), .dinb(n2244), .dout(n2252));
  jxor g02060(.dina(n2252), .dinb(n2235), .dout(n2253));
  jxor g02061(.dina(n2253), .dinb(n2226), .dout(n2254));
  jxor g02062(.dina(n2254), .dinb(n2196), .dout(n2255));
  jand g02063(.dina(n2145), .dinb(n2143), .dout(n2256));
  jand g02064(.dina(n2146), .dinb(n2141), .dout(n2257));
  jor  g02065(.dina(n2257), .dinb(n2256), .dout(n2258));
  jand g02066(.dina(\a[21] ), .dinb(\a[12] ), .dout(n2259));
  jand g02067(.dina(\a[19] ), .dinb(\a[14] ), .dout(n2260));
  jor  g02068(.dina(n2260), .dinb(n2102), .dout(n2261));
  jnot g02069(.din(n2261), .dout(n2262));
  jand g02070(.dina(\a[20] ), .dinb(\a[14] ), .dout(n2263));
  jand g02071(.dina(n2263), .dinb(n1948), .dout(n2264));
  jor  g02072(.dina(n2264), .dinb(n2262), .dout(n2265));
  jxor g02073(.dina(n2265), .dinb(n2259), .dout(n2266));
  jnot g02074(.din(n2266), .dout(n2267));
  jand g02075(.dina(\a[32] ), .dinb(\a[1] ), .dout(n2268));
  jxor g02076(.dina(n2268), .dinb(\a[17] ), .dout(n2269));
  jand g02077(.dina(n2142), .dinb(n1983), .dout(n2270));
  jand g02078(.dina(\a[23] ), .dinb(\a[10] ), .dout(n2271));
  jxor g02079(.dina(n2271), .dinb(n2270), .dout(n2272));
  jxor g02080(.dina(n2272), .dinb(n2269), .dout(n2273));
  jxor g02081(.dina(n2273), .dinb(n2267), .dout(n2274));
  jxor g02082(.dina(n2274), .dinb(n2258), .dout(n2275));
  jand g02083(.dina(n2157), .dinb(n2154), .dout(n2276));
  jand g02084(.dina(n2164), .dinb(n2158), .dout(n2277));
  jor  g02085(.dina(n2277), .dinb(n2276), .dout(n2278));
  jxor g02086(.dina(n2278), .dinb(n2275), .dout(n2279));
  jand g02087(.dina(n2147), .dinb(n2139), .dout(n2280));
  jand g02088(.dina(n2148), .dinb(n2131), .dout(n2281));
  jor  g02089(.dina(n2281), .dinb(n2280), .dout(n2282));
  jxor g02090(.dina(n2282), .dinb(n2279), .dout(n2283));
  jand g02091(.dina(n2168), .dinb(n2165), .dout(n2284));
  jand g02092(.dina(n2169), .dinb(n2149), .dout(n2285));
  jor  g02093(.dina(n2285), .dinb(n2284), .dout(n2286));
  jxor g02094(.dina(n2286), .dinb(n2283), .dout(n2287));
  jxor g02095(.dina(n2287), .dinb(n2255), .dout(n2288));
  jand g02096(.dina(n2127), .dinb(n2069), .dout(n2289));
  jand g02097(.dina(n2170), .dinb(n2128), .dout(n2290));
  jor  g02098(.dina(n2290), .dinb(n2289), .dout(n2291));
  jxor g02099(.dina(n2291), .dinb(n2288), .dout(n2292));
  jand g02100(.dina(n2171), .dinb(n2066), .dout(n2293));
  jor  g02101(.dina(n2171), .dinb(n2066), .dout(n2294));
  jand g02102(.dina(n2176), .dinb(n2294), .dout(n2295));
  jor  g02103(.dina(n2295), .dinb(n2293), .dout(n2296));
  jxor g02104(.dina(n2296), .dinb(n2292), .dout(\asquared[34] ));
  jand g02105(.dina(n2286), .dinb(n2283), .dout(n2298));
  jand g02106(.dina(n2287), .dinb(n2255), .dout(n2299));
  jor  g02107(.dina(n2299), .dinb(n2298), .dout(n2300));
  jand g02108(.dina(n2278), .dinb(n2275), .dout(n2301));
  jand g02109(.dina(n2282), .dinb(n2279), .dout(n2302));
  jor  g02110(.dina(n2302), .dinb(n2301), .dout(n2303));
  jnot g02111(.din(n2219), .dout(n2304));
  jand g02112(.dina(n2304), .dinb(n2214), .dout(n2305));
  jor  g02113(.dina(n2305), .dinb(n2221), .dout(n2306));
  jand g02114(.dina(n2248), .dinb(n2247), .dout(n2307));
  jnot g02115(.din(n2307), .dout(n2308));
  jnot g02116(.din(n2247), .dout(n2309));
  jnot g02117(.din(n2248), .dout(n2310));
  jand g02118(.dina(n2310), .dinb(n2309), .dout(n2311));
  jor  g02119(.dina(n2311), .dinb(n2246), .dout(n2312));
  jand g02120(.dina(n2312), .dinb(n2308), .dout(n2313));
  jnot g02121(.din(n2313), .dout(n2314));
  jxor g02122(.dina(n2314), .dinb(n2306), .dout(n2315));
  jand g02123(.dina(n2239), .dinb(n2091), .dout(n2316));
  jor  g02124(.dina(n2316), .dinb(n2241), .dout(n2317));
  jxor g02125(.dina(n2317), .dinb(n2315), .dout(n2318));
  jand g02126(.dina(n2268), .dinb(\a[17] ), .dout(n2319));
  jand g02127(.dina(\a[33] ), .dinb(\a[1] ), .dout(n2320));
  jxor g02128(.dina(n2320), .dinb(n2231), .dout(n2321));
  jxor g02129(.dina(n2321), .dinb(n2319), .dout(n2322));
  jand g02130(.dina(n2230), .dinb(n1990), .dout(n2323));
  jor  g02131(.dina(n2323), .dinb(n2232), .dout(n2324));
  jxor g02132(.dina(n2324), .dinb(n2322), .dout(n2325));
  jnot g02133(.din(n2325), .dout(n2326));
  jnot g02134(.din(n2244), .dout(n2327));
  jand g02135(.dina(n2251), .dinb(n2327), .dout(n2328));
  jnot g02136(.din(n2328), .dout(n2329));
  jand g02137(.dina(n2250), .dinb(n2244), .dout(n2330));
  jor  g02138(.dina(n2330), .dinb(n2235), .dout(n2331));
  jand g02139(.dina(n2331), .dinb(n2329), .dout(n2332));
  jxor g02140(.dina(n2332), .dinb(n2326), .dout(n2333));
  jxor g02141(.dina(n2333), .dinb(n2318), .dout(n2334));
  jand g02142(.dina(n2273), .dinb(n2267), .dout(n2335));
  jand g02143(.dina(n2274), .dinb(n2258), .dout(n2336));
  jor  g02144(.dina(n2336), .dinb(n2335), .dout(n2337));
  jand g02145(.dina(n2271), .dinb(n2270), .dout(n2338));
  jand g02146(.dina(n2272), .dinb(n2269), .dout(n2339));
  jor  g02147(.dina(n2339), .dinb(n2338), .dout(n2340));
  jand g02148(.dina(n2261), .dinb(n2259), .dout(n2341));
  jor  g02149(.dina(n2341), .dinb(n2264), .dout(n2342));
  jxor g02150(.dina(n2342), .dinb(n2340), .dout(n2343));
  jand g02151(.dina(\a[23] ), .dinb(\a[11] ), .dout(n2344));
  jand g02152(.dina(\a[22] ), .dinb(\a[12] ), .dout(n2345));
  jor  g02153(.dina(n2345), .dinb(n2344), .dout(n2346));
  jnot g02154(.din(n2346), .dout(n2347));
  jand g02155(.dina(\a[23] ), .dinb(\a[12] ), .dout(n2348));
  jand g02156(.dina(n2348), .dinb(n2217), .dout(n2349));
  jor  g02157(.dina(n2349), .dinb(n2347), .dout(n2350));
  jxor g02158(.dina(n2350), .dinb(n2112), .dout(n2351));
  jnot g02159(.din(n2351), .dout(n2352));
  jxor g02160(.dina(n2352), .dinb(n2343), .dout(n2353));
  jxor g02161(.dina(n2353), .dinb(n2337), .dout(n2354));
  jand g02162(.dina(\a[28] ), .dinb(\a[6] ), .dout(n2355));
  jnot g02163(.din(n2355), .dout(n2356));
  jand g02164(.dina(\a[27] ), .dinb(\a[7] ), .dout(n2357));
  jor  g02165(.dina(n2357), .dinb(n1809), .dout(n2358));
  jand g02166(.dina(n2240), .dinb(n1990), .dout(n2359));
  jnot g02167(.din(n2359), .dout(n2360));
  jand g02168(.dina(n2360), .dinb(n2358), .dout(n2361));
  jxor g02169(.dina(n2361), .dinb(n2356), .dout(n2362));
  jand g02170(.dina(\a[21] ), .dinb(\a[13] ), .dout(n2363));
  jnot g02171(.din(n2363), .dout(n2364));
  jand g02172(.dina(\a[19] ), .dinb(\a[15] ), .dout(n2365));
  jor  g02173(.dina(n2365), .dinb(n2263), .dout(n2366));
  jand g02174(.dina(\a[20] ), .dinb(\a[15] ), .dout(n2367));
  jand g02175(.dina(n2367), .dinb(n2260), .dout(n2368));
  jnot g02176(.din(n2368), .dout(n2369));
  jand g02177(.dina(n2369), .dinb(n2366), .dout(n2370));
  jxor g02178(.dina(n2370), .dinb(n2364), .dout(n2371));
  jand g02179(.dina(\a[24] ), .dinb(\a[10] ), .dout(n2372));
  jnot g02180(.din(n2372), .dout(n2373));
  jand g02181(.dina(\a[29] ), .dinb(\a[5] ), .dout(n2374));
  jand g02182(.dina(\a[25] ), .dinb(\a[9] ), .dout(n2375));
  jxor g02183(.dina(n2375), .dinb(n2374), .dout(n2376));
  jxor g02184(.dina(n2376), .dinb(n2373), .dout(n2377));
  jnot g02185(.din(n2377), .dout(n2378));
  jxor g02186(.dina(n2378), .dinb(n2371), .dout(n2379));
  jxor g02187(.dina(n2379), .dinb(n2362), .dout(n2380));
  jxor g02188(.dina(n2380), .dinb(n2354), .dout(n2381));
  jxor g02189(.dina(n2381), .dinb(n2334), .dout(n2382));
  jxor g02190(.dina(n2382), .dinb(n2303), .dout(n2383));
  jand g02191(.dina(n2195), .dinb(n2192), .dout(n2384));
  jand g02192(.dina(n2254), .dinb(n2196), .dout(n2385));
  jor  g02193(.dina(n2385), .dinb(n2384), .dout(n2386));
  jand g02194(.dina(n2225), .dinb(n2208), .dout(n2387));
  jand g02195(.dina(n2253), .dinb(n2226), .dout(n2388));
  jor  g02196(.dina(n2388), .dinb(n2387), .dout(n2389));
  jand g02197(.dina(n2187), .dinb(n2180), .dout(n2390));
  jand g02198(.dina(n2191), .dinb(n2188), .dout(n2391));
  jor  g02199(.dina(n2391), .dinb(n2390), .dout(n2392));
  jxor g02200(.dina(n2392), .dinb(n2389), .dout(n2393));
  jand g02201(.dina(n2200), .dinb(n2198), .dout(n2394));
  jand g02202(.dina(n2207), .dinb(n2201), .dout(n2395));
  jor  g02203(.dina(n2395), .dinb(n2394), .dout(n2396));
  jand g02204(.dina(\a[31] ), .dinb(\a[3] ), .dout(n2397));
  jand g02205(.dina(\a[30] ), .dinb(\a[4] ), .dout(n2398));
  jor  g02206(.dina(n2398), .dinb(n2397), .dout(n2399));
  jand g02207(.dina(\a[31] ), .dinb(\a[4] ), .dout(n2400));
  jand g02208(.dina(n2400), .dinb(n2245), .dout(n2401));
  jnot g02209(.din(n2401), .dout(n2402));
  jand g02210(.dina(n2402), .dinb(n2399), .dout(n2403));
  jand g02211(.dina(\a[34] ), .dinb(\a[0] ), .dout(n2404));
  jnot g02212(.din(n2404), .dout(n2405));
  jxor g02213(.dina(n2405), .dinb(n2403), .dout(n2406));
  jnot g02214(.din(n2406), .dout(n2407));
  jxor g02215(.dina(n2407), .dinb(n2396), .dout(n2408));
  jnot g02216(.din(n2210), .dout(n2409));
  jnot g02217(.din(n2212), .dout(n2410));
  jand g02218(.dina(n2410), .dinb(n2409), .dout(n2411));
  jnot g02219(.din(n2411), .dout(n2412));
  jand g02220(.dina(n2212), .dinb(n2210), .dout(n2413));
  jor  g02221(.dina(n2224), .dinb(n2413), .dout(n2414));
  jand g02222(.dina(n2414), .dinb(n2412), .dout(n2415));
  jxor g02223(.dina(n2415), .dinb(n2408), .dout(n2416));
  jxor g02224(.dina(n2416), .dinb(n2393), .dout(n2417));
  jxor g02225(.dina(n2417), .dinb(n2386), .dout(n2418));
  jxor g02226(.dina(n2418), .dinb(n2383), .dout(n2419));
  jxor g02227(.dina(n2419), .dinb(n2300), .dout(n2420));
  jand g02228(.dina(n2291), .dinb(n2288), .dout(n2421));
  jnot g02229(.din(n2288), .dout(n2422));
  jnot g02230(.din(n2291), .dout(n2423));
  jand g02231(.dina(n2423), .dinb(n2422), .dout(n2424));
  jnot g02232(.din(n2424), .dout(n2425));
  jand g02233(.dina(n2296), .dinb(n2425), .dout(n2426));
  jor  g02234(.dina(n2426), .dinb(n2421), .dout(n2427));
  jxor g02235(.dina(n2427), .dinb(n2420), .dout(\asquared[35] ));
  jand g02236(.dina(n2417), .dinb(n2386), .dout(n2429));
  jand g02237(.dina(n2418), .dinb(n2383), .dout(n2430));
  jor  g02238(.dina(n2430), .dinb(n2429), .dout(n2431));
  jand g02239(.dina(n2381), .dinb(n2334), .dout(n2432));
  jand g02240(.dina(n2382), .dinb(n2303), .dout(n2433));
  jor  g02241(.dina(n2433), .dinb(n2432), .dout(n2434));
  jand g02242(.dina(n2314), .dinb(n2306), .dout(n2435));
  jand g02243(.dina(n2317), .dinb(n2315), .dout(n2436));
  jor  g02244(.dina(n2436), .dinb(n2435), .dout(n2437));
  jand g02245(.dina(n2321), .dinb(n2319), .dout(n2438));
  jand g02246(.dina(n2324), .dinb(n2322), .dout(n2439));
  jor  g02247(.dina(n2439), .dinb(n2438), .dout(n2440));
  jxor g02248(.dina(n2440), .dinb(n2437), .dout(n2441));
  jnot g02249(.din(n2340), .dout(n2442));
  jnot g02250(.din(n2342), .dout(n2443));
  jand g02251(.dina(n2443), .dinb(n2442), .dout(n2444));
  jnot g02252(.din(n2444), .dout(n2445));
  jand g02253(.dina(n2342), .dinb(n2340), .dout(n2446));
  jor  g02254(.dina(n2352), .dinb(n2446), .dout(n2447));
  jand g02255(.dina(n2447), .dinb(n2445), .dout(n2448));
  jxor g02256(.dina(n2448), .dinb(n2441), .dout(n2449));
  jnot g02257(.din(n2449), .dout(n2450));
  jor  g02258(.dina(n2332), .dinb(n2326), .dout(n2451));
  jand g02259(.dina(n2333), .dinb(n2318), .dout(n2452));
  jnot g02260(.din(n2452), .dout(n2453));
  jand g02261(.dina(n2453), .dinb(n2451), .dout(n2454));
  jxor g02262(.dina(n2454), .dinb(n2450), .dout(n2455));
  jand g02263(.dina(n2353), .dinb(n2337), .dout(n2456));
  jand g02264(.dina(n2380), .dinb(n2354), .dout(n2457));
  jor  g02265(.dina(n2457), .dinb(n2456), .dout(n2458));
  jxor g02266(.dina(n2458), .dinb(n2455), .dout(n2459));
  jxor g02267(.dina(n2459), .dinb(n2434), .dout(n2460));
  jand g02268(.dina(n2392), .dinb(n2389), .dout(n2461));
  jand g02269(.dina(n2416), .dinb(n2393), .dout(n2462));
  jor  g02270(.dina(n2462), .dinb(n2461), .dout(n2463));
  jand g02271(.dina(n2346), .dinb(n2112), .dout(n2464));
  jor  g02272(.dina(n2464), .dinb(n2349), .dout(n2465));
  jand g02273(.dina(n2366), .dinb(n2363), .dout(n2466));
  jor  g02274(.dina(n2466), .dinb(n2368), .dout(n2467));
  jxor g02275(.dina(n2467), .dinb(n2465), .dout(n2468));
  jand g02276(.dina(n2404), .dinb(n2399), .dout(n2469));
  jor  g02277(.dina(n2469), .dinb(n2401), .dout(n2470));
  jxor g02278(.dina(n2470), .dinb(n2468), .dout(n2471));
  jand g02279(.dina(n821), .dinb(\a[34] ), .dout(n2472));
  jnot g02280(.din(n2472), .dout(n2473));
  jand g02281(.dina(\a[34] ), .dinb(\a[1] ), .dout(n2474));
  jor  g02282(.dina(n2474), .dinb(\a[18] ), .dout(n2475));
  jand g02283(.dina(n2475), .dinb(n2473), .dout(n2476));
  jand g02284(.dina(n2358), .dinb(n2355), .dout(n2477));
  jor  g02285(.dina(n2477), .dinb(n2359), .dout(n2478));
  jxor g02286(.dina(n2478), .dinb(n2476), .dout(n2479));
  jnot g02287(.din(n2374), .dout(n2480));
  jnot g02288(.din(n2375), .dout(n2481));
  jand g02289(.dina(n2481), .dinb(n2480), .dout(n2482));
  jnot g02290(.din(n2482), .dout(n2483));
  jand g02291(.dina(n2375), .dinb(n2374), .dout(n2484));
  jor  g02292(.dina(n2484), .dinb(n2372), .dout(n2485));
  jand g02293(.dina(n2485), .dinb(n2483), .dout(n2486));
  jxor g02294(.dina(n2486), .dinb(n2479), .dout(n2487));
  jnot g02295(.din(n2487), .dout(n2488));
  jnot g02296(.din(n2371), .dout(n2489));
  jand g02297(.dina(n2378), .dinb(n2489), .dout(n2490));
  jnot g02298(.din(n2490), .dout(n2491));
  jand g02299(.dina(n2377), .dinb(n2371), .dout(n2492));
  jor  g02300(.dina(n2492), .dinb(n2362), .dout(n2493));
  jand g02301(.dina(n2493), .dinb(n2491), .dout(n2494));
  jxor g02302(.dina(n2494), .dinb(n2488), .dout(n2495));
  jxor g02303(.dina(n2495), .dinb(n2471), .dout(n2496));
  jxor g02304(.dina(n2496), .dinb(n2463), .dout(n2497));
  jand g02305(.dina(n2407), .dinb(n2396), .dout(n2498));
  jand g02306(.dina(n2415), .dinb(n2408), .dout(n2499));
  jor  g02307(.dina(n2499), .dinb(n2498), .dout(n2500));
  jand g02308(.dina(\a[26] ), .dinb(\a[9] ), .dout(n2501));
  jand g02309(.dina(\a[25] ), .dinb(\a[10] ), .dout(n2502));
  jor  g02310(.dina(n2502), .dinb(n2501), .dout(n2503));
  jnot g02311(.din(n2503), .dout(n2504));
  jand g02312(.dina(\a[26] ), .dinb(\a[10] ), .dout(n2505));
  jand g02313(.dina(n2505), .dinb(n2375), .dout(n2506));
  jor  g02314(.dina(n2506), .dinb(n2504), .dout(n2507));
  jxor g02315(.dina(n2507), .dinb(n2400), .dout(n2508));
  jnot g02316(.din(n2508), .dout(n2509));
  jand g02317(.dina(\a[28] ), .dinb(\a[7] ), .dout(n2510));
  jand g02318(.dina(\a[18] ), .dinb(\a[17] ), .dout(n2511));
  jnot g02319(.din(n2511), .dout(n2512));
  jand g02320(.dina(\a[19] ), .dinb(\a[16] ), .dout(n2513));
  jxor g02321(.dina(n2513), .dinb(n2512), .dout(n2514));
  jxor g02322(.dina(n2514), .dinb(n2510), .dout(n2515));
  jnot g02323(.din(n2515), .dout(n2516));
  jand g02324(.dina(\a[30] ), .dinb(\a[5] ), .dout(n2517));
  jand g02325(.dina(\a[29] ), .dinb(\a[6] ), .dout(n2518));
  jor  g02326(.dina(n2518), .dinb(n2240), .dout(n2519));
  jand g02327(.dina(\a[29] ), .dinb(\a[8] ), .dout(n2520));
  jand g02328(.dina(n2520), .dinb(n2238), .dout(n2521));
  jnot g02329(.din(n2521), .dout(n2522));
  jand g02330(.dina(n2522), .dinb(n2519), .dout(n2523));
  jxor g02331(.dina(n2523), .dinb(n2517), .dout(n2524));
  jxor g02332(.dina(n2524), .dinb(n2516), .dout(n2525));
  jxor g02333(.dina(n2525), .dinb(n2509), .dout(n2526));
  jxor g02334(.dina(n2526), .dinb(n2500), .dout(n2527));
  jand g02335(.dina(\a[22] ), .dinb(\a[13] ), .dout(n2528));
  jnot g02336(.din(n2528), .dout(n2529));
  jand g02337(.dina(\a[21] ), .dinb(\a[14] ), .dout(n2530));
  jor  g02338(.dina(n2530), .dinb(n2367), .dout(n2531));
  jand g02339(.dina(\a[21] ), .dinb(\a[15] ), .dout(n2532));
  jand g02340(.dina(n2532), .dinb(n2263), .dout(n2533));
  jnot g02341(.din(n2533), .dout(n2534));
  jand g02342(.dina(n2534), .dinb(n2531), .dout(n2535));
  jxor g02343(.dina(n2535), .dinb(n2529), .dout(n2536));
  jand g02344(.dina(\a[32] ), .dinb(\a[3] ), .dout(n2537));
  jnot g02345(.din(n2537), .dout(n2538));
  jand g02346(.dina(\a[24] ), .dinb(\a[11] ), .dout(n2539));
  jor  g02347(.dina(n2539), .dinb(n2348), .dout(n2540));
  jand g02348(.dina(\a[24] ), .dinb(\a[12] ), .dout(n2541));
  jand g02349(.dina(n2541), .dinb(n2344), .dout(n2542));
  jnot g02350(.din(n2542), .dout(n2543));
  jand g02351(.dina(n2543), .dinb(n2540), .dout(n2544));
  jxor g02352(.dina(n2544), .dinb(n2538), .dout(n2545));
  jnot g02353(.din(n2545), .dout(n2546));
  jand g02354(.dina(n2320), .dinb(n2231), .dout(n2547));
  jnot g02355(.din(n2547), .dout(n2548));
  jand g02356(.dina(\a[35] ), .dinb(\a[0] ), .dout(n2549));
  jand g02357(.dina(\a[33] ), .dinb(\a[2] ), .dout(n2550));
  jor  g02358(.dina(n2550), .dinb(n2549), .dout(n2551));
  jand g02359(.dina(\a[35] ), .dinb(\a[2] ), .dout(n2552));
  jand g02360(.dina(n2552), .dinb(n2215), .dout(n2553));
  jnot g02361(.din(n2553), .dout(n2554));
  jand g02362(.dina(n2554), .dinb(n2551), .dout(n2555));
  jxor g02363(.dina(n2555), .dinb(n2548), .dout(n2556));
  jxor g02364(.dina(n2556), .dinb(n2546), .dout(n2557));
  jxor g02365(.dina(n2557), .dinb(n2536), .dout(n2558));
  jxor g02366(.dina(n2558), .dinb(n2527), .dout(n2559));
  jxor g02367(.dina(n2559), .dinb(n2497), .dout(n2560));
  jxor g02368(.dina(n2560), .dinb(n2460), .dout(n2561));
  jxor g02369(.dina(n2561), .dinb(n2431), .dout(n2562));
  jand g02370(.dina(n2419), .dinb(n2300), .dout(n2563));
  jor  g02371(.dina(n2419), .dinb(n2300), .dout(n2564));
  jand g02372(.dina(n2427), .dinb(n2564), .dout(n2565));
  jor  g02373(.dina(n2565), .dinb(n2563), .dout(n2566));
  jxor g02374(.dina(n2566), .dinb(n2562), .dout(\asquared[36] ));
  jand g02375(.dina(n2459), .dinb(n2434), .dout(n2568));
  jand g02376(.dina(n2560), .dinb(n2460), .dout(n2569));
  jor  g02377(.dina(n2569), .dinb(n2568), .dout(n2570));
  jand g02378(.dina(n2496), .dinb(n2463), .dout(n2571));
  jand g02379(.dina(n2559), .dinb(n2497), .dout(n2572));
  jor  g02380(.dina(n2572), .dinb(n2571), .dout(n2573));
  jand g02381(.dina(n2467), .dinb(n2465), .dout(n2574));
  jand g02382(.dina(n2470), .dinb(n2468), .dout(n2575));
  jor  g02383(.dina(n2575), .dinb(n2574), .dout(n2576));
  jand g02384(.dina(n2478), .dinb(n2476), .dout(n2577));
  jand g02385(.dina(n2486), .dinb(n2479), .dout(n2578));
  jor  g02386(.dina(n2578), .dinb(n2577), .dout(n2579));
  jxor g02387(.dina(n2579), .dinb(n2576), .dout(n2580));
  jnot g02388(.din(n2580), .dout(n2581));
  jnot g02389(.din(n2556), .dout(n2582));
  jand g02390(.dina(n2582), .dinb(n2546), .dout(n2583));
  jnot g02391(.din(n2583), .dout(n2584));
  jand g02392(.dina(n2556), .dinb(n2545), .dout(n2585));
  jor  g02393(.dina(n2585), .dinb(n2536), .dout(n2586));
  jand g02394(.dina(n2586), .dinb(n2584), .dout(n2587));
  jxor g02395(.dina(n2587), .dinb(n2581), .dout(n2588));
  jnot g02396(.din(n2588), .dout(n2589));
  jor  g02397(.dina(n2494), .dinb(n2488), .dout(n2590));
  jand g02398(.dina(n2495), .dinb(n2471), .dout(n2591));
  jnot g02399(.din(n2591), .dout(n2592));
  jand g02400(.dina(n2592), .dinb(n2590), .dout(n2593));
  jxor g02401(.dina(n2593), .dinb(n2589), .dout(n2594));
  jand g02402(.dina(n2526), .dinb(n2500), .dout(n2595));
  jand g02403(.dina(n2558), .dinb(n2527), .dout(n2596));
  jor  g02404(.dina(n2596), .dinb(n2595), .dout(n2597));
  jxor g02405(.dina(n2597), .dinb(n2594), .dout(n2598));
  jxor g02406(.dina(n2598), .dinb(n2573), .dout(n2599));
  jor  g02407(.dina(n2454), .dinb(n2450), .dout(n2600));
  jand g02408(.dina(n2458), .dinb(n2455), .dout(n2601));
  jnot g02409(.din(n2601), .dout(n2602));
  jand g02410(.dina(n2602), .dinb(n2600), .dout(n2603));
  jnot g02411(.din(n2603), .dout(n2604));
  jand g02412(.dina(n2523), .dinb(n2517), .dout(n2605));
  jor  g02413(.dina(n2605), .dinb(n2521), .dout(n2606));
  jand g02414(.dina(n2503), .dinb(n2400), .dout(n2607));
  jor  g02415(.dina(n2607), .dinb(n2506), .dout(n2608));
  jxor g02416(.dina(n2608), .dinb(n2606), .dout(n2609));
  jnot g02417(.din(n2513), .dout(n2610));
  jand g02418(.dina(n2610), .dinb(n2512), .dout(n2611));
  jnot g02419(.din(n2611), .dout(n2612));
  jand g02420(.dina(n2513), .dinb(n2511), .dout(n2613));
  jor  g02421(.dina(n2613), .dinb(n2510), .dout(n2614));
  jand g02422(.dina(n2614), .dinb(n2612), .dout(n2615));
  jxor g02423(.dina(n2615), .dinb(n2609), .dout(n2616));
  jand g02424(.dina(n2540), .dinb(n2537), .dout(n2617));
  jor  g02425(.dina(n2617), .dinb(n2542), .dout(n2618));
  jand g02426(.dina(n2531), .dinb(n2528), .dout(n2619));
  jor  g02427(.dina(n2619), .dinb(n2533), .dout(n2620));
  jxor g02428(.dina(n2620), .dinb(n2618), .dout(n2621));
  jand g02429(.dina(n2551), .dinb(n2547), .dout(n2622));
  jor  g02430(.dina(n2622), .dinb(n2553), .dout(n2623));
  jxor g02431(.dina(n2623), .dinb(n2621), .dout(n2624));
  jor  g02432(.dina(n2524), .dinb(n2516), .dout(n2625));
  jand g02433(.dina(n2524), .dinb(n2516), .dout(n2626));
  jor  g02434(.dina(n2626), .dinb(n2509), .dout(n2627));
  jand g02435(.dina(n2627), .dinb(n2625), .dout(n2628));
  jxor g02436(.dina(n2628), .dinb(n2624), .dout(n2629));
  jxor g02437(.dina(n2629), .dinb(n2616), .dout(n2630));
  jxor g02438(.dina(n2630), .dinb(n2604), .dout(n2631));
  jand g02439(.dina(n2440), .dinb(n2437), .dout(n2632));
  jand g02440(.dina(n2448), .dinb(n2441), .dout(n2633));
  jor  g02441(.dina(n2633), .dinb(n2632), .dout(n2634));
  jand g02442(.dina(\a[36] ), .dinb(\a[0] ), .dout(n2635));
  jxor g02443(.dina(n2635), .dinb(n2472), .dout(n2636));
  jand g02444(.dina(\a[19] ), .dinb(\a[17] ), .dout(n2637));
  jand g02445(.dina(\a[35] ), .dinb(\a[1] ), .dout(n2638));
  jxor g02446(.dina(n2638), .dinb(n2637), .dout(n2639));
  jnot g02447(.din(n2639), .dout(n2640));
  jxor g02448(.dina(n2640), .dinb(n2636), .dout(n2641));
  jnot g02449(.din(n2641), .dout(n2642));
  jand g02450(.dina(\a[22] ), .dinb(\a[14] ), .dout(n2643));
  jand g02451(.dina(\a[20] ), .dinb(\a[16] ), .dout(n2644));
  jor  g02452(.dina(n2644), .dinb(n2532), .dout(n2645));
  jnot g02453(.din(n2645), .dout(n2646));
  jand g02454(.dina(\a[21] ), .dinb(\a[16] ), .dout(n2647));
  jand g02455(.dina(n2647), .dinb(n2367), .dout(n2648));
  jor  g02456(.dina(n2648), .dinb(n2646), .dout(n2649));
  jxor g02457(.dina(n2649), .dinb(n2643), .dout(n2650));
  jand g02458(.dina(\a[33] ), .dinb(\a[3] ), .dout(n2651));
  jand g02459(.dina(\a[32] ), .dinb(\a[4] ), .dout(n2652));
  jnot g02460(.din(n2652), .dout(n2653));
  jand g02461(.dina(\a[25] ), .dinb(\a[11] ), .dout(n2654));
  jxor g02462(.dina(n2654), .dinb(n2653), .dout(n2655));
  jxor g02463(.dina(n2655), .dinb(n2651), .dout(n2656));
  jxor g02464(.dina(n2656), .dinb(n2650), .dout(n2657));
  jxor g02465(.dina(n2657), .dinb(n2642), .dout(n2658));
  jxor g02466(.dina(n2658), .dinb(n2634), .dout(n2659));
  jand g02467(.dina(\a[30] ), .dinb(\a[6] ), .dout(n2660));
  jand g02468(.dina(\a[29] ), .dinb(\a[7] ), .dout(n2661));
  jand g02469(.dina(\a[28] ), .dinb(\a[8] ), .dout(n2662));
  jor  g02470(.dina(n2662), .dinb(n2661), .dout(n2663));
  jnot g02471(.din(n2663), .dout(n2664));
  jand g02472(.dina(n2520), .dinb(n2510), .dout(n2665));
  jor  g02473(.dina(n2665), .dinb(n2664), .dout(n2666));
  jxor g02474(.dina(n2666), .dinb(n2660), .dout(n2667));
  jand g02475(.dina(\a[31] ), .dinb(\a[5] ), .dout(n2668));
  jand g02476(.dina(\a[27] ), .dinb(\a[9] ), .dout(n2669));
  jor  g02477(.dina(n2669), .dinb(n2668), .dout(n2670));
  jnot g02478(.din(n2670), .dout(n2671));
  jand g02479(.dina(n2088), .dinb(n1964), .dout(n2672));
  jor  g02480(.dina(n2672), .dinb(n2671), .dout(n2673));
  jxor g02481(.dina(n2673), .dinb(n2505), .dout(n2674));
  jand g02482(.dina(\a[34] ), .dinb(\a[2] ), .dout(n2675));
  jand g02483(.dina(\a[23] ), .dinb(\a[13] ), .dout(n2676));
  jor  g02484(.dina(n2676), .dinb(n2541), .dout(n2677));
  jand g02485(.dina(\a[24] ), .dinb(\a[13] ), .dout(n2678));
  jand g02486(.dina(n2678), .dinb(n2348), .dout(n2679));
  jnot g02487(.din(n2679), .dout(n2680));
  jand g02488(.dina(n2680), .dinb(n2677), .dout(n2681));
  jxor g02489(.dina(n2681), .dinb(n2675), .dout(n2682));
  jxor g02490(.dina(n2682), .dinb(n2674), .dout(n2683));
  jxor g02491(.dina(n2683), .dinb(n2667), .dout(n2684));
  jxor g02492(.dina(n2684), .dinb(n2659), .dout(n2685));
  jxor g02493(.dina(n2685), .dinb(n2631), .dout(n2686));
  jxor g02494(.dina(n2686), .dinb(n2599), .dout(n2687));
  jxor g02495(.dina(n2687), .dinb(n2570), .dout(n2688));
  jand g02496(.dina(n2561), .dinb(n2431), .dout(n2689));
  jnot g02497(.din(n2431), .dout(n2690));
  jnot g02498(.din(n2561), .dout(n2691));
  jand g02499(.dina(n2691), .dinb(n2690), .dout(n2692));
  jnot g02500(.din(n2692), .dout(n2693));
  jand g02501(.dina(n2566), .dinb(n2693), .dout(n2694));
  jor  g02502(.dina(n2694), .dinb(n2689), .dout(n2695));
  jxor g02503(.dina(n2695), .dinb(n2688), .dout(\asquared[37] ));
  jand g02504(.dina(n2598), .dinb(n2573), .dout(n2697));
  jand g02505(.dina(n2686), .dinb(n2599), .dout(n2698));
  jor  g02506(.dina(n2698), .dinb(n2697), .dout(n2699));
  jor  g02507(.dina(n2593), .dinb(n2589), .dout(n2700));
  jand g02508(.dina(n2597), .dinb(n2594), .dout(n2701));
  jnot g02509(.din(n2701), .dout(n2702));
  jand g02510(.dina(n2702), .dinb(n2700), .dout(n2703));
  jnot g02511(.din(n2703), .dout(n2704));
  jand g02512(.dina(n2681), .dinb(n2675), .dout(n2705));
  jor  g02513(.dina(n2705), .dinb(n2679), .dout(n2706));
  jand g02514(.dina(n2645), .dinb(n2643), .dout(n2707));
  jor  g02515(.dina(n2707), .dinb(n2648), .dout(n2708));
  jnot g02516(.din(n2654), .dout(n2709));
  jand g02517(.dina(n2709), .dinb(n2653), .dout(n2710));
  jnot g02518(.din(n2710), .dout(n2711));
  jand g02519(.dina(n2654), .dinb(n2652), .dout(n2712));
  jor  g02520(.dina(n2712), .dinb(n2651), .dout(n2713));
  jand g02521(.dina(n2713), .dinb(n2711), .dout(n2714));
  jxor g02522(.dina(n2714), .dinb(n2708), .dout(n2715));
  jxor g02523(.dina(n2715), .dinb(n2706), .dout(n2716));
  jnot g02524(.din(n2716), .dout(n2717));
  jor  g02525(.dina(n2656), .dinb(n2650), .dout(n2718));
  jand g02526(.dina(n2657), .dinb(n2642), .dout(n2719));
  jnot g02527(.din(n2719), .dout(n2720));
  jand g02528(.dina(n2720), .dinb(n2718), .dout(n2721));
  jxor g02529(.dina(n2721), .dinb(n2717), .dout(n2722));
  jand g02530(.dina(n2670), .dinb(n2505), .dout(n2723));
  jor  g02531(.dina(n2723), .dinb(n2672), .dout(n2724));
  jnot g02532(.din(n2635), .dout(n2725));
  jand g02533(.dina(n2725), .dinb(n2473), .dout(n2726));
  jnot g02534(.din(n2726), .dout(n2727));
  jand g02535(.dina(n2635), .dinb(n2472), .dout(n2728));
  jor  g02536(.dina(n2639), .dinb(n2728), .dout(n2729));
  jand g02537(.dina(n2729), .dinb(n2727), .dout(n2730));
  jxor g02538(.dina(n2730), .dinb(n2724), .dout(n2731));
  jand g02539(.dina(\a[23] ), .dinb(\a[14] ), .dout(n2732));
  jand g02540(.dina(\a[22] ), .dinb(\a[15] ), .dout(n2733));
  jor  g02541(.dina(n2733), .dinb(n2732), .dout(n2734));
  jnot g02542(.din(n2734), .dout(n2735));
  jand g02543(.dina(\a[23] ), .dinb(\a[15] ), .dout(n2736));
  jand g02544(.dina(n2736), .dinb(n2643), .dout(n2737));
  jor  g02545(.dina(n2737), .dinb(n2735), .dout(n2738));
  jxor g02546(.dina(n2738), .dinb(n2678), .dout(n2739));
  jnot g02547(.din(n2739), .dout(n2740));
  jxor g02548(.dina(n2740), .dinb(n2731), .dout(n2741));
  jxor g02549(.dina(n2741), .dinb(n2722), .dout(n2742));
  jxor g02550(.dina(n2742), .dinb(n2704), .dout(n2743));
  jand g02551(.dina(n2620), .dinb(n2618), .dout(n2744));
  jand g02552(.dina(n2623), .dinb(n2621), .dout(n2745));
  jor  g02553(.dina(n2745), .dinb(n2744), .dout(n2746));
  jand g02554(.dina(\a[19] ), .dinb(\a[18] ), .dout(n2747));
  jand g02555(.dina(\a[20] ), .dinb(\a[17] ), .dout(n2748));
  jor  g02556(.dina(n2748), .dinb(n2747), .dout(n2749));
  jnot g02557(.din(n2749), .dout(n2750));
  jand g02558(.dina(\a[20] ), .dinb(\a[18] ), .dout(n2751));
  jand g02559(.dina(n2751), .dinb(n2637), .dout(n2752));
  jor  g02560(.dina(n2752), .dinb(n2750), .dout(n2753));
  jxor g02561(.dina(n2753), .dinb(n2520), .dout(n2754));
  jnot g02562(.din(n2754), .dout(n2755));
  jand g02563(.dina(\a[26] ), .dinb(\a[11] ), .dout(n2756));
  jand g02564(.dina(\a[32] ), .dinb(\a[5] ), .dout(n2757));
  jand g02565(.dina(\a[27] ), .dinb(\a[10] ), .dout(n2758));
  jor  g02566(.dina(n2758), .dinb(n2757), .dout(n2759));
  jand g02567(.dina(\a[32] ), .dinb(\a[10] ), .dout(n2760));
  jand g02568(.dina(n2760), .dinb(n2088), .dout(n2761));
  jnot g02569(.din(n2761), .dout(n2762));
  jand g02570(.dina(n2762), .dinb(n2759), .dout(n2763));
  jxor g02571(.dina(n2763), .dinb(n2756), .dout(n2764));
  jxor g02572(.dina(n2764), .dinb(n2755), .dout(n2765));
  jxor g02573(.dina(n2765), .dinb(n2746), .dout(n2766));
  jnot g02574(.din(n2766), .dout(n2767));
  jand g02575(.dina(n2579), .dinb(n2576), .dout(n2768));
  jnot g02576(.din(n2768), .dout(n2769));
  jor  g02577(.dina(n2587), .dinb(n2581), .dout(n2770));
  jand g02578(.dina(n2770), .dinb(n2769), .dout(n2771));
  jxor g02579(.dina(n2771), .dinb(n2767), .dout(n2772));
  jand g02580(.dina(\a[28] ), .dinb(\a[9] ), .dout(n2773));
  jnot g02581(.din(n2773), .dout(n2774));
  jand g02582(.dina(\a[31] ), .dinb(\a[6] ), .dout(n2775));
  jand g02583(.dina(\a[30] ), .dinb(\a[7] ), .dout(n2776));
  jor  g02584(.dina(n2776), .dinb(n2775), .dout(n2777));
  jand g02585(.dina(\a[31] ), .dinb(\a[7] ), .dout(n2778));
  jand g02586(.dina(n2778), .dinb(n2660), .dout(n2779));
  jnot g02587(.din(n2779), .dout(n2780));
  jand g02588(.dina(n2780), .dinb(n2777), .dout(n2781));
  jxor g02589(.dina(n2781), .dinb(n2774), .dout(n2782));
  jnot g02590(.din(n2647), .dout(n2783));
  jand g02591(.dina(\a[34] ), .dinb(\a[3] ), .dout(n2784));
  jor  g02592(.dina(n2784), .dinb(n2552), .dout(n2785));
  jand g02593(.dina(\a[35] ), .dinb(\a[3] ), .dout(n2786));
  jand g02594(.dina(n2786), .dinb(n2675), .dout(n2787));
  jnot g02595(.din(n2787), .dout(n2788));
  jand g02596(.dina(n2788), .dinb(n2785), .dout(n2789));
  jxor g02597(.dina(n2789), .dinb(n2783), .dout(n2790));
  jand g02598(.dina(n442), .dinb(\a[25] ), .dout(n2791));
  jand g02599(.dina(n208), .dinb(\a[33] ), .dout(n2792));
  jor  g02600(.dina(n2792), .dinb(n2791), .dout(n2793));
  jand g02601(.dina(n2793), .dinb(\a[37] ), .dout(n2794));
  jnot g02602(.din(n2794), .dout(n2795));
  jand g02603(.dina(\a[25] ), .dinb(\a[12] ), .dout(n2796));
  jand g02604(.dina(\a[33] ), .dinb(\a[4] ), .dout(n2797));
  jor  g02605(.dina(n2797), .dinb(n2796), .dout(n2798));
  jand g02606(.dina(\a[33] ), .dinb(\a[12] ), .dout(n2799));
  jand g02607(.dina(n2799), .dinb(n1633), .dout(n2800));
  jnot g02608(.din(n2800), .dout(n2801));
  jand g02609(.dina(n2801), .dinb(n2798), .dout(n2802));
  jand g02610(.dina(n2802), .dinb(n2795), .dout(n2803));
  jnot g02611(.din(n2802), .dout(n2804));
  jand g02612(.dina(\a[37] ), .dinb(\a[0] ), .dout(n2805));
  jand g02613(.dina(n2805), .dinb(n2804), .dout(n2806));
  jor  g02614(.dina(n2806), .dinb(n2803), .dout(n2807));
  jxor g02615(.dina(n2807), .dinb(n2790), .dout(n2808));
  jxor g02616(.dina(n2808), .dinb(n2782), .dout(n2809));
  jxor g02617(.dina(n2809), .dinb(n2772), .dout(n2810));
  jxor g02618(.dina(n2810), .dinb(n2743), .dout(n2811));
  jand g02619(.dina(n2630), .dinb(n2604), .dout(n2812));
  jand g02620(.dina(n2685), .dinb(n2631), .dout(n2813));
  jor  g02621(.dina(n2813), .dinb(n2812), .dout(n2814));
  jand g02622(.dina(n2628), .dinb(n2624), .dout(n2815));
  jand g02623(.dina(n2629), .dinb(n2616), .dout(n2816));
  jor  g02624(.dina(n2816), .dinb(n2815), .dout(n2817));
  jand g02625(.dina(n2608), .dinb(n2606), .dout(n2818));
  jand g02626(.dina(n2615), .dinb(n2609), .dout(n2819));
  jor  g02627(.dina(n2819), .dinb(n2818), .dout(n2820));
  jand g02628(.dina(n2663), .dinb(n2660), .dout(n2821));
  jor  g02629(.dina(n2821), .dinb(n2665), .dout(n2822));
  jnot g02630(.din(\a[36] ), .dout(n2823));
  jand g02631(.dina(n2638), .dinb(n2637), .dout(n2824));
  jand g02632(.dina(n2824), .dinb(n2823), .dout(n2825));
  jnot g02633(.din(n2825), .dout(n2826));
  jand g02634(.dina(n933), .dinb(\a[36] ), .dout(n2827));
  jnot g02635(.din(n2827), .dout(n2828));
  jand g02636(.dina(\a[36] ), .dinb(\a[1] ), .dout(n2829));
  jor  g02637(.dina(n2829), .dinb(\a[19] ), .dout(n2830));
  jand g02638(.dina(n2830), .dinb(n2828), .dout(n2831));
  jor  g02639(.dina(n2831), .dinb(n2824), .dout(n2832));
  jand g02640(.dina(n2832), .dinb(n2826), .dout(n2833));
  jxor g02641(.dina(n2833), .dinb(n2822), .dout(n2834));
  jxor g02642(.dina(n2834), .dinb(n2820), .dout(n2835));
  jnot g02643(.din(n2674), .dout(n2836));
  jor  g02644(.dina(n2682), .dinb(n2836), .dout(n2837));
  jnot g02645(.din(n2667), .dout(n2838));
  jand g02646(.dina(n2682), .dinb(n2836), .dout(n2839));
  jor  g02647(.dina(n2839), .dinb(n2838), .dout(n2840));
  jand g02648(.dina(n2840), .dinb(n2837), .dout(n2841));
  jxor g02649(.dina(n2841), .dinb(n2835), .dout(n2842));
  jxor g02650(.dina(n2842), .dinb(n2817), .dout(n2843));
  jor  g02651(.dina(n2658), .dinb(n2634), .dout(n2844));
  jand g02652(.dina(n2658), .dinb(n2634), .dout(n2845));
  jor  g02653(.dina(n2684), .dinb(n2845), .dout(n2846));
  jand g02654(.dina(n2846), .dinb(n2844), .dout(n2847));
  jxor g02655(.dina(n2847), .dinb(n2843), .dout(n2848));
  jxor g02656(.dina(n2848), .dinb(n2814), .dout(n2849));
  jxor g02657(.dina(n2849), .dinb(n2811), .dout(n2850));
  jxor g02658(.dina(n2850), .dinb(n2699), .dout(n2851));
  jand g02659(.dina(n2687), .dinb(n2570), .dout(n2852));
  jnot g02660(.din(n2570), .dout(n2853));
  jnot g02661(.din(n2687), .dout(n2854));
  jand g02662(.dina(n2854), .dinb(n2853), .dout(n2855));
  jnot g02663(.din(n2855), .dout(n2856));
  jand g02664(.dina(n2695), .dinb(n2856), .dout(n2857));
  jor  g02665(.dina(n2857), .dinb(n2852), .dout(n2858));
  jxor g02666(.dina(n2858), .dinb(n2851), .dout(\asquared[38] ));
  jand g02667(.dina(n2848), .dinb(n2814), .dout(n2860));
  jand g02668(.dina(n2849), .dinb(n2811), .dout(n2861));
  jor  g02669(.dina(n2861), .dinb(n2860), .dout(n2862));
  jand g02670(.dina(n2742), .dinb(n2704), .dout(n2863));
  jand g02671(.dina(n2810), .dinb(n2743), .dout(n2864));
  jor  g02672(.dina(n2864), .dinb(n2863), .dout(n2865));
  jand g02673(.dina(n2801), .dinb(n2795), .dout(n2866));
  jnot g02674(.din(n2866), .dout(n2867));
  jand g02675(.dina(n2785), .dinb(n2647), .dout(n2868));
  jor  g02676(.dina(n2868), .dinb(n2787), .dout(n2869));
  jxor g02677(.dina(n2869), .dinb(n2867), .dout(n2870));
  jand g02678(.dina(n2734), .dinb(n2678), .dout(n2871));
  jor  g02679(.dina(n2871), .dinb(n2737), .dout(n2872));
  jxor g02680(.dina(n2872), .dinb(n2870), .dout(n2873));
  jand g02681(.dina(n2764), .dinb(n2755), .dout(n2874));
  jand g02682(.dina(n2765), .dinb(n2746), .dout(n2875));
  jor  g02683(.dina(n2875), .dinb(n2874), .dout(n2876));
  jxor g02684(.dina(n2876), .dinb(n2873), .dout(n2877));
  jand g02685(.dina(\a[29] ), .dinb(\a[9] ), .dout(n2878));
  jand g02686(.dina(\a[30] ), .dinb(\a[8] ), .dout(n2879));
  jor  g02687(.dina(n2879), .dinb(n2778), .dout(n2880));
  jnot g02688(.din(n2880), .dout(n2881));
  jand g02689(.dina(\a[31] ), .dinb(\a[8] ), .dout(n2882));
  jand g02690(.dina(n2882), .dinb(n2776), .dout(n2883));
  jor  g02691(.dina(n2883), .dinb(n2881), .dout(n2884));
  jxor g02692(.dina(n2884), .dinb(n2878), .dout(n2885));
  jnot g02693(.din(n2885), .dout(n2886));
  jand g02694(.dina(\a[22] ), .dinb(\a[16] ), .dout(n2887));
  jand g02695(.dina(\a[21] ), .dinb(\a[17] ), .dout(n2888));
  jor  g02696(.dina(n2888), .dinb(n2887), .dout(n2889));
  jnot g02697(.din(n2889), .dout(n2890));
  jand g02698(.dina(\a[22] ), .dinb(\a[17] ), .dout(n2891));
  jand g02699(.dina(n2891), .dinb(n2647), .dout(n2892));
  jor  g02700(.dina(n2892), .dinb(n2890), .dout(n2893));
  jxor g02701(.dina(n2893), .dinb(n2736), .dout(n2894));
  jand g02702(.dina(\a[33] ), .dinb(\a[5] ), .dout(n2895));
  jand g02703(.dina(\a[32] ), .dinb(\a[6] ), .dout(n2896));
  jnot g02704(.din(n2896), .dout(n2897));
  jand g02705(.dina(\a[28] ), .dinb(\a[10] ), .dout(n2898));
  jxor g02706(.dina(n2898), .dinb(n2897), .dout(n2899));
  jxor g02707(.dina(n2899), .dinb(n2895), .dout(n2900));
  jxor g02708(.dina(n2900), .dinb(n2894), .dout(n2901));
  jxor g02709(.dina(n2901), .dinb(n2886), .dout(n2902));
  jxor g02710(.dina(n2902), .dinb(n2877), .dout(n2903));
  jor  g02711(.dina(n2771), .dinb(n2767), .dout(n2904));
  jand g02712(.dina(n2809), .dinb(n2772), .dout(n2905));
  jnot g02713(.din(n2905), .dout(n2906));
  jand g02714(.dina(n2906), .dinb(n2904), .dout(n2907));
  jor  g02715(.dina(n2721), .dinb(n2717), .dout(n2908));
  jand g02716(.dina(n2741), .dinb(n2722), .dout(n2909));
  jnot g02717(.din(n2909), .dout(n2910));
  jand g02718(.dina(n2910), .dinb(n2908), .dout(n2911));
  jxor g02719(.dina(n2911), .dinb(n2907), .dout(n2912));
  jxor g02720(.dina(n2912), .dinb(n2903), .dout(n2913));
  jxor g02721(.dina(n2913), .dinb(n2865), .dout(n2914));
  jand g02722(.dina(n2842), .dinb(n2817), .dout(n2915));
  jand g02723(.dina(n2847), .dinb(n2843), .dout(n2916));
  jor  g02724(.dina(n2916), .dinb(n2915), .dout(n2917));
  jnot g02725(.din(n2790), .dout(n2918));
  jand g02726(.dina(n2807), .dinb(n2918), .dout(n2919));
  jnot g02727(.din(n2919), .dout(n2920));
  jnot g02728(.din(n2807), .dout(n2921));
  jand g02729(.dina(n2921), .dinb(n2790), .dout(n2922));
  jor  g02730(.dina(n2922), .dinb(n2782), .dout(n2923));
  jand g02731(.dina(n2923), .dinb(n2920), .dout(n2924));
  jnot g02732(.din(n2724), .dout(n2925));
  jnot g02733(.din(n2730), .dout(n2926));
  jand g02734(.dina(n2926), .dinb(n2925), .dout(n2927));
  jnot g02735(.din(n2927), .dout(n2928));
  jand g02736(.dina(n2730), .dinb(n2724), .dout(n2929));
  jor  g02737(.dina(n2740), .dinb(n2929), .dout(n2930));
  jand g02738(.dina(n2930), .dinb(n2928), .dout(n2931));
  jnot g02739(.din(n2931), .dout(n2932));
  jxor g02740(.dina(n2932), .dinb(n2924), .dout(n2933));
  jand g02741(.dina(\a[37] ), .dinb(\a[1] ), .dout(n2934));
  jxor g02742(.dina(n2934), .dinb(n2751), .dout(n2935));
  jand g02743(.dina(n2749), .dinb(n2520), .dout(n2936));
  jor  g02744(.dina(n2936), .dinb(n2752), .dout(n2937));
  jxor g02745(.dina(n2937), .dinb(n2935), .dout(n2938));
  jand g02746(.dina(n2777), .dinb(n2773), .dout(n2939));
  jor  g02747(.dina(n2939), .dinb(n2779), .dout(n2940));
  jxor g02748(.dina(n2940), .dinb(n2938), .dout(n2941));
  jxor g02749(.dina(n2941), .dinb(n2933), .dout(n2942));
  jxor g02750(.dina(n2942), .dinb(n2917), .dout(n2943));
  jand g02751(.dina(n2714), .dinb(n2708), .dout(n2944));
  jand g02752(.dina(n2715), .dinb(n2706), .dout(n2945));
  jor  g02753(.dina(n2945), .dinb(n2944), .dout(n2946));
  jand g02754(.dina(n2833), .dinb(n2822), .dout(n2947));
  jor  g02755(.dina(n2947), .dinb(n2825), .dout(n2948));
  jnot g02756(.din(n2948), .dout(n2949));
  jand g02757(.dina(\a[26] ), .dinb(\a[12] ), .dout(n2950));
  jand g02758(.dina(\a[34] ), .dinb(\a[4] ), .dout(n2951));
  jand g02759(.dina(\a[27] ), .dinb(\a[11] ), .dout(n2952));
  jor  g02760(.dina(n2952), .dinb(n2951), .dout(n2953));
  jnot g02761(.din(n2953), .dout(n2954));
  jand g02762(.dina(\a[34] ), .dinb(\a[11] ), .dout(n2955));
  jand g02763(.dina(n2955), .dinb(n1971), .dout(n2956));
  jor  g02764(.dina(n2956), .dinb(n2954), .dout(n2957));
  jxor g02765(.dina(n2957), .dinb(n2950), .dout(n2958));
  jxor g02766(.dina(n2958), .dinb(n2949), .dout(n2959));
  jxor g02767(.dina(n2959), .dinb(n2946), .dout(n2960));
  jand g02768(.dina(n2834), .dinb(n2820), .dout(n2961));
  jand g02769(.dina(n2841), .dinb(n2835), .dout(n2962));
  jor  g02770(.dina(n2962), .dinb(n2961), .dout(n2963));
  jand g02771(.dina(\a[25] ), .dinb(\a[13] ), .dout(n2964));
  jand g02772(.dina(\a[24] ), .dinb(\a[14] ), .dout(n2965));
  jor  g02773(.dina(n2965), .dinb(n2964), .dout(n2966));
  jnot g02774(.din(n2966), .dout(n2967));
  jand g02775(.dina(\a[25] ), .dinb(\a[14] ), .dout(n2968));
  jand g02776(.dina(n2968), .dinb(n2678), .dout(n2969));
  jor  g02777(.dina(n2969), .dinb(n2967), .dout(n2970));
  jxor g02778(.dina(n2970), .dinb(n2786), .dout(n2971));
  jnot g02779(.din(n2971), .dout(n2972));
  jand g02780(.dina(n2763), .dinb(n2756), .dout(n2973));
  jor  g02781(.dina(n2973), .dinb(n2761), .dout(n2974));
  jnot g02782(.din(n2974), .dout(n2975));
  jand g02783(.dina(\a[38] ), .dinb(\a[0] ), .dout(n2976));
  jand g02784(.dina(\a[36] ), .dinb(\a[2] ), .dout(n2977));
  jor  g02785(.dina(n2977), .dinb(n2976), .dout(n2978));
  jand g02786(.dina(\a[38] ), .dinb(\a[2] ), .dout(n2979));
  jand g02787(.dina(n2979), .dinb(n2635), .dout(n2980));
  jnot g02788(.din(n2980), .dout(n2981));
  jand g02789(.dina(n2981), .dinb(n2978), .dout(n2982));
  jxor g02790(.dina(n2982), .dinb(n2828), .dout(n2983));
  jxor g02791(.dina(n2983), .dinb(n2975), .dout(n2984));
  jxor g02792(.dina(n2984), .dinb(n2972), .dout(n2985));
  jxor g02793(.dina(n2985), .dinb(n2963), .dout(n2986));
  jxor g02794(.dina(n2986), .dinb(n2960), .dout(n2987));
  jxor g02795(.dina(n2987), .dinb(n2943), .dout(n2988));
  jxor g02796(.dina(n2988), .dinb(n2914), .dout(n2989));
  jxor g02797(.dina(n2989), .dinb(n2862), .dout(n2990));
  jand g02798(.dina(n2850), .dinb(n2699), .dout(n2991));
  jor  g02799(.dina(n2850), .dinb(n2699), .dout(n2992));
  jand g02800(.dina(n2858), .dinb(n2992), .dout(n2993));
  jor  g02801(.dina(n2993), .dinb(n2991), .dout(n2994));
  jxor g02802(.dina(n2994), .dinb(n2990), .dout(\asquared[39] ));
  jand g02803(.dina(n2913), .dinb(n2865), .dout(n2996));
  jand g02804(.dina(n2988), .dinb(n2914), .dout(n2997));
  jor  g02805(.dina(n2997), .dinb(n2996), .dout(n2998));
  jand g02806(.dina(n2942), .dinb(n2917), .dout(n2999));
  jand g02807(.dina(n2987), .dinb(n2943), .dout(n3000));
  jor  g02808(.dina(n3000), .dinb(n2999), .dout(n3001));
  jand g02809(.dina(n2985), .dinb(n2963), .dout(n3002));
  jand g02810(.dina(n2986), .dinb(n2960), .dout(n3003));
  jor  g02811(.dina(n3003), .dinb(n3002), .dout(n3004));
  jand g02812(.dina(n2937), .dinb(n2935), .dout(n3005));
  jand g02813(.dina(n2940), .dinb(n2938), .dout(n3006));
  jor  g02814(.dina(n3006), .dinb(n3005), .dout(n3007));
  jand g02815(.dina(n2934), .dinb(n2751), .dout(n3008));
  jand g02816(.dina(\a[39] ), .dinb(\a[0] ), .dout(n3009));
  jxor g02817(.dina(n3009), .dinb(n3008), .dout(n3010));
  jand g02818(.dina(n1036), .dinb(\a[38] ), .dout(n3011));
  jnot g02819(.din(n3011), .dout(n3012));
  jand g02820(.dina(n3012), .dinb(\a[20] ), .dout(n3013));
  jnot g02821(.din(\a[20] ), .dout(n3014));
  jand g02822(.dina(\a[38] ), .dinb(\a[1] ), .dout(n3015));
  jand g02823(.dina(n3015), .dinb(n3014), .dout(n3016));
  jor  g02824(.dina(n3016), .dinb(n3013), .dout(n3017));
  jxor g02825(.dina(n3017), .dinb(n3010), .dout(n3018));
  jxor g02826(.dina(n3018), .dinb(n3007), .dout(n3019));
  jand g02827(.dina(n2869), .dinb(n2867), .dout(n3020));
  jand g02828(.dina(n2872), .dinb(n2870), .dout(n3021));
  jor  g02829(.dina(n3021), .dinb(n3020), .dout(n3022));
  jxor g02830(.dina(n3022), .dinb(n3019), .dout(n3023));
  jand g02831(.dina(n2966), .dinb(n2786), .dout(n3024));
  jor  g02832(.dina(n3024), .dinb(n2969), .dout(n3025));
  jand g02833(.dina(n2978), .dinb(n2827), .dout(n3026));
  jor  g02834(.dina(n3026), .dinb(n2980), .dout(n3027));
  jxor g02835(.dina(n3027), .dinb(n3025), .dout(n3028));
  jand g02836(.dina(n2889), .dinb(n2736), .dout(n3029));
  jor  g02837(.dina(n3029), .dinb(n2892), .dout(n3030));
  jxor g02838(.dina(n3030), .dinb(n3028), .dout(n3031));
  jor  g02839(.dina(n2900), .dinb(n2894), .dout(n3032));
  jand g02840(.dina(n2901), .dinb(n2886), .dout(n3033));
  jnot g02841(.din(n3033), .dout(n3034));
  jand g02842(.dina(n3034), .dinb(n3032), .dout(n3035));
  jor  g02843(.dina(n2983), .dinb(n2975), .dout(n3036));
  jand g02844(.dina(n2984), .dinb(n2972), .dout(n3037));
  jnot g02845(.din(n3037), .dout(n3038));
  jand g02846(.dina(n3038), .dinb(n3036), .dout(n3039));
  jxor g02847(.dina(n3039), .dinb(n3035), .dout(n3040));
  jxor g02848(.dina(n3040), .dinb(n3031), .dout(n3041));
  jxor g02849(.dina(n3041), .dinb(n3023), .dout(n3042));
  jxor g02850(.dina(n3042), .dinb(n3004), .dout(n3043));
  jxor g02851(.dina(n3043), .dinb(n3001), .dout(n3044));
  jor  g02852(.dina(n2932), .dinb(n2924), .dout(n3045));
  jand g02853(.dina(n2941), .dinb(n2933), .dout(n3046));
  jnot g02854(.din(n3046), .dout(n3047));
  jand g02855(.dina(n3047), .dinb(n3045), .dout(n3048));
  jnot g02856(.din(n3048), .dout(n3049));
  jand g02857(.dina(\a[24] ), .dinb(\a[15] ), .dout(n3050));
  jand g02858(.dina(\a[23] ), .dinb(\a[16] ), .dout(n3051));
  jor  g02859(.dina(n3051), .dinb(n3050), .dout(n3052));
  jnot g02860(.din(n3052), .dout(n3053));
  jand g02861(.dina(\a[24] ), .dinb(\a[16] ), .dout(n3054));
  jand g02862(.dina(n3054), .dinb(n2736), .dout(n3055));
  jor  g02863(.dina(n3055), .dinb(n3053), .dout(n3056));
  jxor g02864(.dina(n3056), .dinb(n2968), .dout(n3057));
  jand g02865(.dina(\a[37] ), .dinb(\a[2] ), .dout(n3058));
  jnot g02866(.din(n3058), .dout(n3059));
  jand g02867(.dina(\a[36] ), .dinb(\a[3] ), .dout(n3060));
  jand g02868(.dina(\a[26] ), .dinb(\a[13] ), .dout(n3061));
  jxor g02869(.dina(n3061), .dinb(n3060), .dout(n3062));
  jxor g02870(.dina(n3062), .dinb(n3059), .dout(n3063));
  jxor g02871(.dina(n3063), .dinb(n3057), .dout(n3064));
  jand g02872(.dina(\a[33] ), .dinb(\a[7] ), .dout(n3065));
  jand g02873(.dina(n3065), .dinb(n2896), .dout(n3066));
  jand g02874(.dina(\a[33] ), .dinb(\a[6] ), .dout(n3067));
  jand g02875(.dina(\a[30] ), .dinb(\a[9] ), .dout(n3068));
  jand g02876(.dina(n3068), .dinb(n3067), .dout(n3069));
  jor  g02877(.dina(n3069), .dinb(n3066), .dout(n3070));
  jand g02878(.dina(\a[32] ), .dinb(\a[9] ), .dout(n3071));
  jand g02879(.dina(n3071), .dinb(n2776), .dout(n3072));
  jnot g02880(.din(n3072), .dout(n3073));
  jand g02881(.dina(n3073), .dinb(n3070), .dout(n3074));
  jnot g02882(.din(n3074), .dout(n3075));
  jand g02883(.dina(\a[32] ), .dinb(\a[7] ), .dout(n3076));
  jor  g02884(.dina(n3076), .dinb(n3068), .dout(n3077));
  jand g02885(.dina(n3077), .dinb(n3073), .dout(n3078));
  jor  g02886(.dina(n3078), .dinb(n3067), .dout(n3079));
  jand g02887(.dina(n3079), .dinb(n3075), .dout(n3080));
  jxor g02888(.dina(n3080), .dinb(n3064), .dout(n3081));
  jxor g02889(.dina(n3081), .dinb(n3049), .dout(n3082));
  jand g02890(.dina(n2876), .dinb(n2873), .dout(n3083));
  jand g02891(.dina(n2902), .dinb(n2877), .dout(n3084));
  jor  g02892(.dina(n3084), .dinb(n3083), .dout(n3085));
  jxor g02893(.dina(n3085), .dinb(n3082), .dout(n3086));
  jor  g02894(.dina(n2911), .dinb(n2907), .dout(n3087));
  jand g02895(.dina(n2912), .dinb(n2903), .dout(n3088));
  jnot g02896(.din(n3088), .dout(n3089));
  jand g02897(.dina(n3089), .dinb(n3087), .dout(n3090));
  jnot g02898(.din(n3090), .dout(n3091));
  jand g02899(.dina(n2880), .dinb(n2878), .dout(n3092));
  jor  g02900(.dina(n3092), .dinb(n2883), .dout(n3093));
  jand g02901(.dina(n2953), .dinb(n2950), .dout(n3094));
  jor  g02902(.dina(n3094), .dinb(n2956), .dout(n3095));
  jxor g02903(.dina(n3095), .dinb(n3093), .dout(n3096));
  jnot g02904(.din(n2898), .dout(n3097));
  jand g02905(.dina(n3097), .dinb(n2897), .dout(n3098));
  jnot g02906(.din(n3098), .dout(n3099));
  jand g02907(.dina(n2898), .dinb(n2896), .dout(n3100));
  jor  g02908(.dina(n3100), .dinb(n2895), .dout(n3101));
  jand g02909(.dina(n3101), .dinb(n3099), .dout(n3102));
  jxor g02910(.dina(n3102), .dinb(n3096), .dout(n3103));
  jnot g02911(.din(n3103), .dout(n3104));
  jor  g02912(.dina(n2958), .dinb(n2949), .dout(n3105));
  jand g02913(.dina(n2959), .dinb(n2946), .dout(n3106));
  jnot g02914(.din(n3106), .dout(n3107));
  jand g02915(.dina(n3107), .dinb(n3105), .dout(n3108));
  jxor g02916(.dina(n3108), .dinb(n3104), .dout(n3109));
  jand g02917(.dina(\a[20] ), .dinb(\a[19] ), .dout(n3110));
  jand g02918(.dina(\a[21] ), .dinb(\a[18] ), .dout(n3111));
  jor  g02919(.dina(n3111), .dinb(n3110), .dout(n3112));
  jnot g02920(.din(n3112), .dout(n3113));
  jand g02921(.dina(\a[21] ), .dinb(\a[19] ), .dout(n3114));
  jand g02922(.dina(n3114), .dinb(n2751), .dout(n3115));
  jor  g02923(.dina(n3115), .dinb(n3113), .dout(n3116));
  jxor g02924(.dina(n3116), .dinb(n2882), .dout(n3117));
  jand g02925(.dina(\a[35] ), .dinb(\a[4] ), .dout(n3118));
  jnot g02926(.din(n3118), .dout(n3119));
  jand g02927(.dina(\a[27] ), .dinb(\a[12] ), .dout(n3120));
  jxor g02928(.dina(n3120), .dinb(n3119), .dout(n3121));
  jxor g02929(.dina(n3121), .dinb(n2891), .dout(n3122));
  jxor g02930(.dina(n3122), .dinb(n3117), .dout(n3123));
  jnot g02931(.din(n3123), .dout(n3124));
  jand g02932(.dina(\a[28] ), .dinb(\a[11] ), .dout(n3125));
  jand g02933(.dina(\a[29] ), .dinb(\a[10] ), .dout(n3126));
  jand g02934(.dina(\a[34] ), .dinb(\a[5] ), .dout(n3127));
  jor  g02935(.dina(n3127), .dinb(n3126), .dout(n3128));
  jnot g02936(.din(n3128), .dout(n3129));
  jand g02937(.dina(\a[34] ), .dinb(\a[10] ), .dout(n3130));
  jand g02938(.dina(n3130), .dinb(n2374), .dout(n3131));
  jor  g02939(.dina(n3131), .dinb(n3129), .dout(n3132));
  jxor g02940(.dina(n3132), .dinb(n3125), .dout(n3133));
  jxor g02941(.dina(n3133), .dinb(n3124), .dout(n3134));
  jxor g02942(.dina(n3134), .dinb(n3109), .dout(n3135));
  jxor g02943(.dina(n3135), .dinb(n3091), .dout(n3136));
  jxor g02944(.dina(n3136), .dinb(n3086), .dout(n3137));
  jxor g02945(.dina(n3137), .dinb(n3044), .dout(n3138));
  jxor g02946(.dina(n3138), .dinb(n2998), .dout(n3139));
  jand g02947(.dina(n2989), .dinb(n2862), .dout(n3140));
  jor  g02948(.dina(n2989), .dinb(n2862), .dout(n3141));
  jand g02949(.dina(n2994), .dinb(n3141), .dout(n3142));
  jor  g02950(.dina(n3142), .dinb(n3140), .dout(n3143));
  jxor g02951(.dina(n3143), .dinb(n3139), .dout(\asquared[40] ));
  jand g02952(.dina(n3043), .dinb(n3001), .dout(n3145));
  jand g02953(.dina(n3137), .dinb(n3044), .dout(n3146));
  jor  g02954(.dina(n3146), .dinb(n3145), .dout(n3147));
  jand g02955(.dina(n3052), .dinb(n2968), .dout(n3148));
  jor  g02956(.dina(n3148), .dinb(n3055), .dout(n3149));
  jor  g02957(.dina(n3072), .dinb(n3070), .dout(n3150));
  jxor g02958(.dina(n3150), .dinb(n3149), .dout(n3151));
  jand g02959(.dina(n3009), .dinb(n3008), .dout(n3152));
  jand g02960(.dina(n3017), .dinb(n3010), .dout(n3153));
  jor  g02961(.dina(n3153), .dinb(n3152), .dout(n3154));
  jxor g02962(.dina(n3154), .dinb(n3151), .dout(n3155));
  jand g02963(.dina(n3018), .dinb(n3007), .dout(n3156));
  jand g02964(.dina(n3022), .dinb(n3019), .dout(n3157));
  jor  g02965(.dina(n3157), .dinb(n3156), .dout(n3158));
  jxor g02966(.dina(n3158), .dinb(n3155), .dout(n3159));
  jand g02967(.dina(\a[36] ), .dinb(\a[4] ), .dout(n3160));
  jnot g02968(.din(n3160), .dout(n3161));
  jand g02969(.dina(\a[28] ), .dinb(\a[12] ), .dout(n3162));
  jand g02970(.dina(\a[35] ), .dinb(\a[5] ), .dout(n3163));
  jxor g02971(.dina(n3163), .dinb(n3162), .dout(n3164));
  jxor g02972(.dina(n3164), .dinb(n3161), .dout(n3165));
  jand g02973(.dina(\a[32] ), .dinb(\a[8] ), .dout(n3166));
  jor  g02974(.dina(n3166), .dinb(n1964), .dout(n3167));
  jnot g02975(.din(n3167), .dout(n3168));
  jand g02976(.dina(n3071), .dinb(n2882), .dout(n3169));
  jor  g02977(.dina(n3169), .dinb(n3168), .dout(n3170));
  jxor g02978(.dina(n3170), .dinb(n3065), .dout(n3171));
  jand g02979(.dina(\a[22] ), .dinb(\a[18] ), .dout(n3172));
  jand g02980(.dina(\a[40] ), .dinb(\a[0] ), .dout(n3173));
  jor  g02981(.dina(n3173), .dinb(n2979), .dout(n3174));
  jand g02982(.dina(\a[40] ), .dinb(\a[2] ), .dout(n3175));
  jand g02983(.dina(n3175), .dinb(n2976), .dout(n3176));
  jnot g02984(.din(n3176), .dout(n3177));
  jand g02985(.dina(n3177), .dinb(n3174), .dout(n3178));
  jxor g02986(.dina(n3178), .dinb(n3172), .dout(n3179));
  jxor g02987(.dina(n3179), .dinb(n3171), .dout(n3180));
  jxor g02988(.dina(n3180), .dinb(n3165), .dout(n3181));
  jxor g02989(.dina(n3181), .dinb(n3159), .dout(n3182));
  jand g02990(.dina(n3041), .dinb(n3023), .dout(n3183));
  jand g02991(.dina(n3042), .dinb(n3004), .dout(n3184));
  jor  g02992(.dina(n3184), .dinb(n3183), .dout(n3185));
  jxor g02993(.dina(n3185), .dinb(n3182), .dout(n3186));
  jor  g02994(.dina(n3039), .dinb(n3035), .dout(n3187));
  jand g02995(.dina(n3040), .dinb(n3031), .dout(n3188));
  jnot g02996(.din(n3188), .dout(n3189));
  jand g02997(.dina(n3189), .dinb(n3187), .dout(n3190));
  jnot g02998(.din(n3190), .dout(n3191));
  jand g02999(.dina(\a[25] ), .dinb(\a[15] ), .dout(n3192));
  jand g03000(.dina(\a[23] ), .dinb(\a[17] ), .dout(n3193));
  jor  g03001(.dina(n3193), .dinb(n3054), .dout(n3194));
  jnot g03002(.din(n3194), .dout(n3195));
  jand g03003(.dina(\a[24] ), .dinb(\a[17] ), .dout(n3196));
  jand g03004(.dina(n3196), .dinb(n3051), .dout(n3197));
  jor  g03005(.dina(n3197), .dinb(n3195), .dout(n3198));
  jxor g03006(.dina(n3198), .dinb(n3192), .dout(n3199));
  jnot g03007(.din(n3199), .dout(n3200));
  jand g03008(.dina(\a[37] ), .dinb(\a[3] ), .dout(n3201));
  jand g03009(.dina(\a[27] ), .dinb(\a[13] ), .dout(n3202));
  jand g03010(.dina(\a[26] ), .dinb(\a[14] ), .dout(n3203));
  jor  g03011(.dina(n3203), .dinb(n3202), .dout(n3204));
  jand g03012(.dina(\a[27] ), .dinb(\a[14] ), .dout(n3205));
  jand g03013(.dina(n3205), .dinb(n3061), .dout(n3206));
  jnot g03014(.din(n3206), .dout(n3207));
  jand g03015(.dina(n3207), .dinb(n3204), .dout(n3208));
  jxor g03016(.dina(n3208), .dinb(n3201), .dout(n3209));
  jxor g03017(.dina(n3209), .dinb(n3200), .dout(n3210));
  jand g03018(.dina(\a[29] ), .dinb(\a[11] ), .dout(n3211));
  jand g03019(.dina(\a[34] ), .dinb(\a[6] ), .dout(n3212));
  jnot g03020(.din(n3212), .dout(n3213));
  jand g03021(.dina(\a[30] ), .dinb(\a[10] ), .dout(n3214));
  jxor g03022(.dina(n3214), .dinb(n3213), .dout(n3215));
  jxor g03023(.dina(n3215), .dinb(n3211), .dout(n3216));
  jnot g03024(.din(n3216), .dout(n3217));
  jxor g03025(.dina(n3217), .dinb(n3210), .dout(n3218));
  jxor g03026(.dina(n3218), .dinb(n3191), .dout(n3219));
  jand g03027(.dina(n3095), .dinb(n3093), .dout(n3220));
  jand g03028(.dina(n3102), .dinb(n3096), .dout(n3221));
  jor  g03029(.dina(n3221), .dinb(n3220), .dout(n3222));
  jand g03030(.dina(n3027), .dinb(n3025), .dout(n3223));
  jand g03031(.dina(n3030), .dinb(n3028), .dout(n3224));
  jor  g03032(.dina(n3224), .dinb(n3223), .dout(n3225));
  jxor g03033(.dina(n3225), .dinb(n3222), .dout(n3226));
  jand g03034(.dina(\a[39] ), .dinb(\a[1] ), .dout(n3227));
  jxor g03035(.dina(n3227), .dinb(n3114), .dout(n3228));
  jxor g03036(.dina(n3228), .dinb(n3011), .dout(n3229));
  jand g03037(.dina(n3112), .dinb(n2882), .dout(n3230));
  jor  g03038(.dina(n3230), .dinb(n3115), .dout(n3231));
  jxor g03039(.dina(n3231), .dinb(n3229), .dout(n3232));
  jxor g03040(.dina(n3232), .dinb(n3226), .dout(n3233));
  jxor g03041(.dina(n3233), .dinb(n3219), .dout(n3234));
  jxor g03042(.dina(n3234), .dinb(n3186), .dout(n3235));
  jand g03043(.dina(n3081), .dinb(n3049), .dout(n3236));
  jand g03044(.dina(n3085), .dinb(n3082), .dout(n3237));
  jor  g03045(.dina(n3237), .dinb(n3236), .dout(n3238));
  jor  g03046(.dina(n3108), .dinb(n3104), .dout(n3239));
  jand g03047(.dina(n3134), .dinb(n3109), .dout(n3240));
  jnot g03048(.din(n3240), .dout(n3241));
  jand g03049(.dina(n3241), .dinb(n3239), .dout(n3242));
  jnot g03050(.din(n3242), .dout(n3243));
  jand g03051(.dina(n3128), .dinb(n3125), .dout(n3244));
  jor  g03052(.dina(n3244), .dinb(n3131), .dout(n3245));
  jand g03053(.dina(n3061), .dinb(n3060), .dout(n3246));
  jnot g03054(.din(n3246), .dout(n3247));
  jnot g03055(.din(n3060), .dout(n3248));
  jnot g03056(.din(n3061), .dout(n3249));
  jand g03057(.dina(n3249), .dinb(n3248), .dout(n3250));
  jor  g03058(.dina(n3250), .dinb(n3059), .dout(n3251));
  jand g03059(.dina(n3251), .dinb(n3247), .dout(n3252));
  jnot g03060(.din(n3252), .dout(n3253));
  jxor g03061(.dina(n3253), .dinb(n3245), .dout(n3254));
  jnot g03062(.din(n3120), .dout(n3255));
  jand g03063(.dina(n3255), .dinb(n3119), .dout(n3256));
  jnot g03064(.din(n3256), .dout(n3257));
  jand g03065(.dina(n3120), .dinb(n3118), .dout(n3258));
  jor  g03066(.dina(n3258), .dinb(n2891), .dout(n3259));
  jand g03067(.dina(n3259), .dinb(n3257), .dout(n3260));
  jxor g03068(.dina(n3260), .dinb(n3254), .dout(n3261));
  jor  g03069(.dina(n3122), .dinb(n3117), .dout(n3262));
  jor  g03070(.dina(n3133), .dinb(n3124), .dout(n3263));
  jand g03071(.dina(n3263), .dinb(n3262), .dout(n3264));
  jor  g03072(.dina(n3063), .dinb(n3057), .dout(n3265));
  jand g03073(.dina(n3080), .dinb(n3064), .dout(n3266));
  jnot g03074(.din(n3266), .dout(n3267));
  jand g03075(.dina(n3267), .dinb(n3265), .dout(n3268));
  jxor g03076(.dina(n3268), .dinb(n3264), .dout(n3269));
  jxor g03077(.dina(n3269), .dinb(n3261), .dout(n3270));
  jxor g03078(.dina(n3270), .dinb(n3243), .dout(n3271));
  jxor g03079(.dina(n3271), .dinb(n3238), .dout(n3272));
  jand g03080(.dina(n3135), .dinb(n3091), .dout(n3273));
  jand g03081(.dina(n3136), .dinb(n3086), .dout(n3274));
  jor  g03082(.dina(n3274), .dinb(n3273), .dout(n3275));
  jxor g03083(.dina(n3275), .dinb(n3272), .dout(n3276));
  jxor g03084(.dina(n3276), .dinb(n3235), .dout(n3277));
  jxor g03085(.dina(n3277), .dinb(n3147), .dout(n3278));
  jand g03086(.dina(n3138), .dinb(n2998), .dout(n3279));
  jor  g03087(.dina(n3138), .dinb(n2998), .dout(n3280));
  jand g03088(.dina(n3143), .dinb(n3280), .dout(n3281));
  jor  g03089(.dina(n3281), .dinb(n3279), .dout(n3282));
  jxor g03090(.dina(n3282), .dinb(n3278), .dout(\asquared[41] ));
  jand g03091(.dina(n3275), .dinb(n3272), .dout(n3284));
  jand g03092(.dina(n3276), .dinb(n3235), .dout(n3285));
  jor  g03093(.dina(n3285), .dinb(n3284), .dout(n3286));
  jand g03094(.dina(n3218), .dinb(n3191), .dout(n3287));
  jand g03095(.dina(n3233), .dinb(n3219), .dout(n3288));
  jor  g03096(.dina(n3288), .dinb(n3287), .dout(n3289));
  jand g03097(.dina(n3158), .dinb(n3155), .dout(n3290));
  jand g03098(.dina(n3181), .dinb(n3159), .dout(n3291));
  jor  g03099(.dina(n3291), .dinb(n3290), .dout(n3292));
  jand g03100(.dina(n3208), .dinb(n3201), .dout(n3293));
  jor  g03101(.dina(n3293), .dinb(n3206), .dout(n3294));
  jand g03102(.dina(n3178), .dinb(n3172), .dout(n3295));
  jor  g03103(.dina(n3295), .dinb(n3176), .dout(n3296));
  jand g03104(.dina(n3194), .dinb(n3192), .dout(n3297));
  jor  g03105(.dina(n3297), .dinb(n3197), .dout(n3298));
  jxor g03106(.dina(n3298), .dinb(n3296), .dout(n3299));
  jxor g03107(.dina(n3299), .dinb(n3294), .dout(n3300));
  jnot g03108(.din(n3171), .dout(n3301));
  jor  g03109(.dina(n3179), .dinb(n3301), .dout(n3302));
  jnot g03110(.din(n3165), .dout(n3303));
  jand g03111(.dina(n3179), .dinb(n3301), .dout(n3304));
  jor  g03112(.dina(n3304), .dinb(n3303), .dout(n3305));
  jand g03113(.dina(n3305), .dinb(n3302), .dout(n3306));
  jxor g03114(.dina(n3306), .dinb(n3300), .dout(n3307));
  jand g03115(.dina(n1116), .dinb(\a[40] ), .dout(n3308));
  jnot g03116(.din(n3308), .dout(n3309));
  jand g03117(.dina(\a[40] ), .dinb(\a[1] ), .dout(n3310));
  jor  g03118(.dina(n3310), .dinb(\a[21] ), .dout(n3311));
  jand g03119(.dina(n3311), .dinb(n3309), .dout(n3312));
  jand g03120(.dina(n3167), .dinb(n3065), .dout(n3313));
  jor  g03121(.dina(n3313), .dinb(n3169), .dout(n3314));
  jxor g03122(.dina(n3314), .dinb(n3312), .dout(n3315));
  jnot g03123(.din(n3214), .dout(n3316));
  jand g03124(.dina(n3316), .dinb(n3213), .dout(n3317));
  jnot g03125(.din(n3317), .dout(n3318));
  jand g03126(.dina(n3214), .dinb(n3212), .dout(n3319));
  jor  g03127(.dina(n3319), .dinb(n3211), .dout(n3320));
  jand g03128(.dina(n3320), .dinb(n3318), .dout(n3321));
  jxor g03129(.dina(n3321), .dinb(n3315), .dout(n3322));
  jxor g03130(.dina(n3322), .dinb(n3307), .dout(n3323));
  jxor g03131(.dina(n3323), .dinb(n3292), .dout(n3324));
  jxor g03132(.dina(n3324), .dinb(n3289), .dout(n3325));
  jand g03133(.dina(n3185), .dinb(n3182), .dout(n3326));
  jand g03134(.dina(n3234), .dinb(n3186), .dout(n3327));
  jor  g03135(.dina(n3327), .dinb(n3326), .dout(n3328));
  jxor g03136(.dina(n3328), .dinb(n3325), .dout(n3329));
  jand g03137(.dina(n3150), .dinb(n3149), .dout(n3330));
  jand g03138(.dina(n3154), .dinb(n3151), .dout(n3331));
  jor  g03139(.dina(n3331), .dinb(n3330), .dout(n3332));
  jand g03140(.dina(n3253), .dinb(n3245), .dout(n3333));
  jand g03141(.dina(n3260), .dinb(n3254), .dout(n3334));
  jor  g03142(.dina(n3334), .dinb(n3333), .dout(n3335));
  jxor g03143(.dina(n3335), .dinb(n3332), .dout(n3336));
  jor  g03144(.dina(n3209), .dinb(n3200), .dout(n3337));
  jand g03145(.dina(n3209), .dinb(n3200), .dout(n3338));
  jor  g03146(.dina(n3217), .dinb(n3338), .dout(n3339));
  jand g03147(.dina(n3339), .dinb(n3337), .dout(n3340));
  jxor g03148(.dina(n3340), .dinb(n3336), .dout(n3341));
  jor  g03149(.dina(n3268), .dinb(n3264), .dout(n3342));
  jand g03150(.dina(n3269), .dinb(n3261), .dout(n3343));
  jnot g03151(.din(n3343), .dout(n3344));
  jand g03152(.dina(n3344), .dinb(n3342), .dout(n3345));
  jnot g03153(.din(n3345), .dout(n3346));
  jand g03154(.dina(n3227), .dinb(n3114), .dout(n3347));
  jand g03155(.dina(\a[41] ), .dinb(\a[0] ), .dout(n3348));
  jand g03156(.dina(\a[39] ), .dinb(\a[2] ), .dout(n3349));
  jor  g03157(.dina(n3349), .dinb(n3348), .dout(n3350));
  jand g03158(.dina(\a[41] ), .dinb(\a[2] ), .dout(n3351));
  jand g03159(.dina(n3351), .dinb(n3009), .dout(n3352));
  jnot g03160(.din(n3352), .dout(n3353));
  jand g03161(.dina(n3353), .dinb(n3350), .dout(n3354));
  jxor g03162(.dina(n3354), .dinb(n3347), .dout(n3355));
  jnot g03163(.din(n3355), .dout(n3356));
  jand g03164(.dina(n3163), .dinb(n3162), .dout(n3357));
  jnot g03165(.din(n3357), .dout(n3358));
  jnot g03166(.din(n3162), .dout(n3359));
  jnot g03167(.din(n3163), .dout(n3360));
  jand g03168(.dina(n3360), .dinb(n3359), .dout(n3361));
  jor  g03169(.dina(n3361), .dinb(n3161), .dout(n3362));
  jand g03170(.dina(n3362), .dinb(n3358), .dout(n3363));
  jxor g03171(.dina(n3363), .dinb(n3356), .dout(n3364));
  jnot g03172(.din(n3364), .dout(n3365));
  jand g03173(.dina(\a[38] ), .dinb(\a[3] ), .dout(n3366));
  jand g03174(.dina(\a[28] ), .dinb(\a[13] ), .dout(n3367));
  jand g03175(.dina(\a[26] ), .dinb(\a[15] ), .dout(n3368));
  jor  g03176(.dina(n3368), .dinb(n3367), .dout(n3369));
  jnot g03177(.din(n3369), .dout(n3370));
  jand g03178(.dina(\a[28] ), .dinb(\a[15] ), .dout(n3371));
  jand g03179(.dina(n3371), .dinb(n3061), .dout(n3372));
  jor  g03180(.dina(n3372), .dinb(n3370), .dout(n3373));
  jxor g03181(.dina(n3373), .dinb(n3366), .dout(n3374));
  jxor g03182(.dina(n3374), .dinb(n3365), .dout(n3375));
  jxor g03183(.dina(n3375), .dinb(n3346), .dout(n3376));
  jxor g03184(.dina(n3376), .dinb(n3341), .dout(n3377));
  jand g03185(.dina(n3270), .dinb(n3243), .dout(n3378));
  jand g03186(.dina(n3271), .dinb(n3238), .dout(n3379));
  jor  g03187(.dina(n3379), .dinb(n3378), .dout(n3380));
  jand g03188(.dina(n3228), .dinb(n3011), .dout(n3381));
  jand g03189(.dina(n3231), .dinb(n3229), .dout(n3382));
  jor  g03190(.dina(n3382), .dinb(n3381), .dout(n3383));
  jand g03191(.dina(\a[33] ), .dinb(\a[8] ), .dout(n3384));
  jand g03192(.dina(\a[21] ), .dinb(\a[20] ), .dout(n3385));
  jnot g03193(.din(n3385), .dout(n3386));
  jand g03194(.dina(\a[22] ), .dinb(\a[19] ), .dout(n3387));
  jxor g03195(.dina(n3387), .dinb(n3386), .dout(n3388));
  jxor g03196(.dina(n3388), .dinb(n3384), .dout(n3389));
  jnot g03197(.din(n3389), .dout(n3390));
  jand g03198(.dina(\a[36] ), .dinb(\a[5] ), .dout(n3391));
  jand g03199(.dina(\a[35] ), .dinb(\a[6] ), .dout(n3392));
  jand g03200(.dina(\a[30] ), .dinb(\a[11] ), .dout(n3393));
  jor  g03201(.dina(n3393), .dinb(n3392), .dout(n3394));
  jand g03202(.dina(\a[35] ), .dinb(\a[11] ), .dout(n3395));
  jand g03203(.dina(n3395), .dinb(n2660), .dout(n3396));
  jnot g03204(.din(n3396), .dout(n3397));
  jand g03205(.dina(n3397), .dinb(n3394), .dout(n3398));
  jxor g03206(.dina(n3398), .dinb(n3391), .dout(n3399));
  jxor g03207(.dina(n3399), .dinb(n3390), .dout(n3400));
  jxor g03208(.dina(n3400), .dinb(n3383), .dout(n3401));
  jand g03209(.dina(n3225), .dinb(n3222), .dout(n3402));
  jand g03210(.dina(n3232), .dinb(n3226), .dout(n3403));
  jor  g03211(.dina(n3403), .dinb(n3402), .dout(n3404));
  jxor g03212(.dina(n3404), .dinb(n3401), .dout(n3405));
  jand g03213(.dina(\a[25] ), .dinb(\a[16] ), .dout(n3406));
  jand g03214(.dina(\a[23] ), .dinb(\a[18] ), .dout(n3407));
  jor  g03215(.dina(n3407), .dinb(n3196), .dout(n3408));
  jnot g03216(.din(n3408), .dout(n3409));
  jand g03217(.dina(\a[24] ), .dinb(\a[18] ), .dout(n3410));
  jand g03218(.dina(n3410), .dinb(n3193), .dout(n3411));
  jor  g03219(.dina(n3411), .dinb(n3409), .dout(n3412));
  jxor g03220(.dina(n3412), .dinb(n3406), .dout(n3413));
  jnot g03221(.din(n3205), .dout(n3414));
  jand g03222(.dina(\a[37] ), .dinb(\a[4] ), .dout(n3415));
  jand g03223(.dina(\a[29] ), .dinb(\a[12] ), .dout(n3416));
  jxor g03224(.dina(n3416), .dinb(n3415), .dout(n3417));
  jxor g03225(.dina(n3417), .dinb(n3414), .dout(n3418));
  jxor g03226(.dina(n3418), .dinb(n3413), .dout(n3419));
  jnot g03227(.din(n3419), .dout(n3420));
  jand g03228(.dina(\a[31] ), .dinb(\a[10] ), .dout(n3421));
  jand g03229(.dina(\a[34] ), .dinb(\a[7] ), .dout(n3422));
  jor  g03230(.dina(n3422), .dinb(n3071), .dout(n3423));
  jnot g03231(.din(n3423), .dout(n3424));
  jand g03232(.dina(\a[34] ), .dinb(\a[9] ), .dout(n3425));
  jand g03233(.dina(n3425), .dinb(n3076), .dout(n3426));
  jor  g03234(.dina(n3426), .dinb(n3424), .dout(n3427));
  jxor g03235(.dina(n3427), .dinb(n3421), .dout(n3428));
  jxor g03236(.dina(n3428), .dinb(n3420), .dout(n3429));
  jxor g03237(.dina(n3429), .dinb(n3405), .dout(n3430));
  jxor g03238(.dina(n3430), .dinb(n3380), .dout(n3431));
  jxor g03239(.dina(n3431), .dinb(n3377), .dout(n3432));
  jxor g03240(.dina(n3432), .dinb(n3329), .dout(n3433));
  jxor g03241(.dina(n3433), .dinb(n3286), .dout(n3434));
  jand g03242(.dina(n3277), .dinb(n3147), .dout(n3435));
  jor  g03243(.dina(n3277), .dinb(n3147), .dout(n3436));
  jand g03244(.dina(n3282), .dinb(n3436), .dout(n3437));
  jor  g03245(.dina(n3437), .dinb(n3435), .dout(n3438));
  jxor g03246(.dina(n3438), .dinb(n3434), .dout(\asquared[42] ));
  jand g03247(.dina(n3328), .dinb(n3325), .dout(n3440));
  jand g03248(.dina(n3432), .dinb(n3329), .dout(n3441));
  jor  g03249(.dina(n3441), .dinb(n3440), .dout(n3442));
  jand g03250(.dina(n3430), .dinb(n3380), .dout(n3443));
  jand g03251(.dina(n3431), .dinb(n3377), .dout(n3444));
  jor  g03252(.dina(n3444), .dinb(n3443), .dout(n3445));
  jand g03253(.dina(n3375), .dinb(n3346), .dout(n3446));
  jand g03254(.dina(n3376), .dinb(n3341), .dout(n3447));
  jor  g03255(.dina(n3447), .dinb(n3446), .dout(n3448));
  jand g03256(.dina(n3298), .dinb(n3296), .dout(n3449));
  jand g03257(.dina(n3299), .dinb(n3294), .dout(n3450));
  jor  g03258(.dina(n3450), .dinb(n3449), .dout(n3451));
  jnot g03259(.din(n3451), .dout(n3452));
  jor  g03260(.dina(n3363), .dinb(n3356), .dout(n3453));
  jor  g03261(.dina(n3374), .dinb(n3365), .dout(n3454));
  jand g03262(.dina(n3454), .dinb(n3453), .dout(n3455));
  jxor g03263(.dina(n3455), .dinb(n3452), .dout(n3456));
  jnot g03264(.din(n3456), .dout(n3457));
  jor  g03265(.dina(n3418), .dinb(n3413), .dout(n3458));
  jor  g03266(.dina(n3428), .dinb(n3420), .dout(n3459));
  jand g03267(.dina(n3459), .dinb(n3458), .dout(n3460));
  jxor g03268(.dina(n3460), .dinb(n3457), .dout(n3461));
  jand g03269(.dina(n3404), .dinb(n3401), .dout(n3462));
  jand g03270(.dina(n3429), .dinb(n3405), .dout(n3463));
  jor  g03271(.dina(n3463), .dinb(n3462), .dout(n3464));
  jxor g03272(.dina(n3464), .dinb(n3461), .dout(n3465));
  jxor g03273(.dina(n3465), .dinb(n3448), .dout(n3466));
  jxor g03274(.dina(n3466), .dinb(n3445), .dout(n3467));
  jand g03275(.dina(n3314), .dinb(n3312), .dout(n3468));
  jand g03276(.dina(n3321), .dinb(n3315), .dout(n3469));
  jor  g03277(.dina(n3469), .dinb(n3468), .dout(n3470));
  jand g03278(.dina(\a[29] ), .dinb(\a[13] ), .dout(n3471));
  jnot g03279(.din(n3471), .dout(n3472));
  jand g03280(.dina(\a[37] ), .dinb(\a[5] ), .dout(n3473));
  jand g03281(.dina(\a[30] ), .dinb(\a[12] ), .dout(n3474));
  jxor g03282(.dina(n3474), .dinb(n3473), .dout(n3475));
  jxor g03283(.dina(n3475), .dinb(n3472), .dout(n3476));
  jand g03284(.dina(\a[42] ), .dinb(\a[0] ), .dout(n3477));
  jxor g03285(.dina(n3477), .dinb(n3308), .dout(n3478));
  jand g03286(.dina(\a[22] ), .dinb(\a[20] ), .dout(n3479));
  jand g03287(.dina(\a[41] ), .dinb(\a[1] ), .dout(n3480));
  jxor g03288(.dina(n3480), .dinb(n3479), .dout(n3481));
  jnot g03289(.din(n3481), .dout(n3482));
  jxor g03290(.dina(n3482), .dinb(n3478), .dout(n3483));
  jxor g03291(.dina(n3483), .dinb(n3476), .dout(n3484));
  jxor g03292(.dina(n3484), .dinb(n3470), .dout(n3485));
  jand g03293(.dina(n3306), .dinb(n3300), .dout(n3486));
  jand g03294(.dina(n3322), .dinb(n3307), .dout(n3487));
  jor  g03295(.dina(n3487), .dinb(n3486), .dout(n3488));
  jxor g03296(.dina(n3488), .dinb(n3485), .dout(n3489));
  jand g03297(.dina(n3398), .dinb(n3391), .dout(n3490));
  jor  g03298(.dina(n3490), .dinb(n3396), .dout(n3491));
  jand g03299(.dina(n3416), .dinb(n3415), .dout(n3492));
  jnot g03300(.din(n3492), .dout(n3493));
  jnot g03301(.din(n3415), .dout(n3494));
  jnot g03302(.din(n3416), .dout(n3495));
  jand g03303(.dina(n3495), .dinb(n3494), .dout(n3496));
  jor  g03304(.dina(n3496), .dinb(n3414), .dout(n3497));
  jand g03305(.dina(n3497), .dinb(n3493), .dout(n3498));
  jnot g03306(.din(n3498), .dout(n3499));
  jnot g03307(.din(n3387), .dout(n3500));
  jand g03308(.dina(n3500), .dinb(n3386), .dout(n3501));
  jnot g03309(.din(n3501), .dout(n3502));
  jand g03310(.dina(n3387), .dinb(n3385), .dout(n3503));
  jor  g03311(.dina(n3503), .dinb(n3384), .dout(n3504));
  jand g03312(.dina(n3504), .dinb(n3502), .dout(n3505));
  jxor g03313(.dina(n3505), .dinb(n3499), .dout(n3506));
  jxor g03314(.dina(n3506), .dinb(n3491), .dout(n3507));
  jand g03315(.dina(n3399), .dinb(n3390), .dout(n3508));
  jand g03316(.dina(n3400), .dinb(n3383), .dout(n3509));
  jor  g03317(.dina(n3509), .dinb(n3508), .dout(n3510));
  jxor g03318(.dina(n3510), .dinb(n3507), .dout(n3511));
  jand g03319(.dina(n3369), .dinb(n3366), .dout(n3512));
  jor  g03320(.dina(n3512), .dinb(n3372), .dout(n3513));
  jand g03321(.dina(n3408), .dinb(n3406), .dout(n3514));
  jor  g03322(.dina(n3514), .dinb(n3411), .dout(n3515));
  jxor g03323(.dina(n3515), .dinb(n3513), .dout(n3516));
  jand g03324(.dina(n3354), .dinb(n3347), .dout(n3517));
  jor  g03325(.dina(n3517), .dinb(n3352), .dout(n3518));
  jxor g03326(.dina(n3518), .dinb(n3516), .dout(n3519));
  jxor g03327(.dina(n3519), .dinb(n3511), .dout(n3520));
  jxor g03328(.dina(n3520), .dinb(n3489), .dout(n3521));
  jand g03329(.dina(n3323), .dinb(n3292), .dout(n3522));
  jand g03330(.dina(n3324), .dinb(n3289), .dout(n3523));
  jor  g03331(.dina(n3523), .dinb(n3522), .dout(n3524));
  jand g03332(.dina(n3335), .dinb(n3332), .dout(n3525));
  jand g03333(.dina(n3340), .dinb(n3336), .dout(n3526));
  jor  g03334(.dina(n3526), .dinb(n3525), .dout(n3527));
  jand g03335(.dina(\a[33] ), .dinb(\a[9] ), .dout(n3528));
  jand g03336(.dina(\a[34] ), .dinb(\a[8] ), .dout(n3529));
  jor  g03337(.dina(n3529), .dinb(n3528), .dout(n3530));
  jnot g03338(.din(n3530), .dout(n3531));
  jand g03339(.dina(n3425), .dinb(n3384), .dout(n3532));
  jor  g03340(.dina(n3532), .dinb(n3531), .dout(n3533));
  jxor g03341(.dina(n3533), .dinb(n2760), .dout(n3534));
  jnot g03342(.din(n3534), .dout(n3535));
  jand g03343(.dina(\a[36] ), .dinb(\a[6] ), .dout(n3536));
  jnot g03344(.din(n3536), .dout(n3537));
  jand g03345(.dina(\a[35] ), .dinb(\a[7] ), .dout(n3538));
  jand g03346(.dina(\a[31] ), .dinb(\a[11] ), .dout(n3539));
  jxor g03347(.dina(n3539), .dinb(n3538), .dout(n3540));
  jxor g03348(.dina(n3540), .dinb(n3537), .dout(n3541));
  jnot g03349(.din(n3541), .dout(n3542));
  jand g03350(.dina(n3423), .dinb(n3421), .dout(n3543));
  jor  g03351(.dina(n3543), .dinb(n3426), .dout(n3544));
  jxor g03352(.dina(n3544), .dinb(n3542), .dout(n3545));
  jxor g03353(.dina(n3545), .dinb(n3535), .dout(n3546));
  jxor g03354(.dina(n3546), .dinb(n3527), .dout(n3547));
  jand g03355(.dina(\a[27] ), .dinb(\a[15] ), .dout(n3548));
  jnot g03356(.din(n3548), .dout(n3549));
  jand g03357(.dina(\a[38] ), .dinb(\a[4] ), .dout(n3550));
  jand g03358(.dina(\a[28] ), .dinb(\a[14] ), .dout(n3551));
  jor  g03359(.dina(n3551), .dinb(n3550), .dout(n3552));
  jand g03360(.dina(\a[38] ), .dinb(\a[14] ), .dout(n3553));
  jand g03361(.dina(n3553), .dinb(n1974), .dout(n3554));
  jnot g03362(.din(n3554), .dout(n3555));
  jand g03363(.dina(n3555), .dinb(n3552), .dout(n3556));
  jxor g03364(.dina(n3556), .dinb(n3549), .dout(n3557));
  jand g03365(.dina(\a[25] ), .dinb(\a[17] ), .dout(n3558));
  jnot g03366(.din(n3558), .dout(n3559));
  jand g03367(.dina(\a[23] ), .dinb(\a[19] ), .dout(n3560));
  jor  g03368(.dina(n3560), .dinb(n3410), .dout(n3561));
  jand g03369(.dina(\a[24] ), .dinb(\a[19] ), .dout(n3562));
  jand g03370(.dina(n3562), .dinb(n3407), .dout(n3563));
  jnot g03371(.din(n3563), .dout(n3564));
  jand g03372(.dina(n3564), .dinb(n3561), .dout(n3565));
  jxor g03373(.dina(n3565), .dinb(n3559), .dout(n3566));
  jnot g03374(.din(n3175), .dout(n3567));
  jand g03375(.dina(\a[39] ), .dinb(\a[3] ), .dout(n3568));
  jand g03376(.dina(\a[26] ), .dinb(\a[16] ), .dout(n3569));
  jxor g03377(.dina(n3569), .dinb(n3568), .dout(n3570));
  jxor g03378(.dina(n3570), .dinb(n3567), .dout(n3571));
  jnot g03379(.din(n3571), .dout(n3572));
  jxor g03380(.dina(n3572), .dinb(n3566), .dout(n3573));
  jxor g03381(.dina(n3573), .dinb(n3557), .dout(n3574));
  jxor g03382(.dina(n3574), .dinb(n3547), .dout(n3575));
  jxor g03383(.dina(n3575), .dinb(n3524), .dout(n3576));
  jxor g03384(.dina(n3576), .dinb(n3521), .dout(n3577));
  jxor g03385(.dina(n3577), .dinb(n3467), .dout(n3578));
  jxor g03386(.dina(n3578), .dinb(n3442), .dout(n3579));
  jand g03387(.dina(n3433), .dinb(n3286), .dout(n3580));
  jnot g03388(.din(n3286), .dout(n3581));
  jnot g03389(.din(n3433), .dout(n3582));
  jand g03390(.dina(n3582), .dinb(n3581), .dout(n3583));
  jnot g03391(.din(n3583), .dout(n3584));
  jand g03392(.dina(n3438), .dinb(n3584), .dout(n3585));
  jor  g03393(.dina(n3585), .dinb(n3580), .dout(n3586));
  jxor g03394(.dina(n3586), .dinb(n3579), .dout(\asquared[43] ));
  jand g03395(.dina(n3466), .dinb(n3445), .dout(n3588));
  jand g03396(.dina(n3577), .dinb(n3467), .dout(n3589));
  jor  g03397(.dina(n3589), .dinb(n3588), .dout(n3590));
  jand g03398(.dina(n3464), .dinb(n3461), .dout(n3591));
  jand g03399(.dina(n3465), .dinb(n3448), .dout(n3592));
  jor  g03400(.dina(n3592), .dinb(n3591), .dout(n3593));
  jor  g03401(.dina(n3455), .dinb(n3452), .dout(n3594));
  jor  g03402(.dina(n3460), .dinb(n3457), .dout(n3595));
  jand g03403(.dina(n3595), .dinb(n3594), .dout(n3596));
  jnot g03404(.din(n3596), .dout(n3597));
  jand g03405(.dina(\a[26] ), .dinb(\a[17] ), .dout(n3598));
  jnot g03406(.din(n3598), .dout(n3599));
  jand g03407(.dina(\a[25] ), .dinb(\a[18] ), .dout(n3600));
  jor  g03408(.dina(n3600), .dinb(n3562), .dout(n3601));
  jand g03409(.dina(\a[25] ), .dinb(\a[19] ), .dout(n3602));
  jand g03410(.dina(n3602), .dinb(n3410), .dout(n3603));
  jnot g03411(.din(n3603), .dout(n3604));
  jand g03412(.dina(n3604), .dinb(n3601), .dout(n3605));
  jxor g03413(.dina(n3605), .dinb(n3599), .dout(n3606));
  jand g03414(.dina(\a[29] ), .dinb(\a[14] ), .dout(n3607));
  jnot g03415(.din(n3607), .dout(n3608));
  jand g03416(.dina(\a[27] ), .dinb(\a[16] ), .dout(n3609));
  jor  g03417(.dina(n3609), .dinb(n3371), .dout(n3610));
  jand g03418(.dina(\a[28] ), .dinb(\a[16] ), .dout(n3611));
  jand g03419(.dina(n3611), .dinb(n3548), .dout(n3612));
  jnot g03420(.din(n3612), .dout(n3613));
  jand g03421(.dina(n3613), .dinb(n3610), .dout(n3614));
  jxor g03422(.dina(n3614), .dinb(n3608), .dout(n3615));
  jand g03423(.dina(\a[39] ), .dinb(\a[4] ), .dout(n3616));
  jnot g03424(.din(n3616), .dout(n3617));
  jand g03425(.dina(\a[43] ), .dinb(\a[0] ), .dout(n3618));
  jand g03426(.dina(\a[40] ), .dinb(\a[3] ), .dout(n3619));
  jxor g03427(.dina(n3619), .dinb(n3618), .dout(n3620));
  jxor g03428(.dina(n3620), .dinb(n3617), .dout(n3621));
  jnot g03429(.din(n3621), .dout(n3622));
  jxor g03430(.dina(n3622), .dinb(n3615), .dout(n3623));
  jxor g03431(.dina(n3623), .dinb(n3606), .dout(n3624));
  jand g03432(.dina(\a[22] ), .dinb(\a[21] ), .dout(n3625));
  jand g03433(.dina(\a[23] ), .dinb(\a[20] ), .dout(n3626));
  jor  g03434(.dina(n3626), .dinb(n3625), .dout(n3627));
  jnot g03435(.din(n3627), .dout(n3628));
  jand g03436(.dina(\a[23] ), .dinb(\a[21] ), .dout(n3629));
  jand g03437(.dina(n3629), .dinb(n3479), .dout(n3630));
  jor  g03438(.dina(n3630), .dinb(n3628), .dout(n3631));
  jxor g03439(.dina(n3631), .dinb(n3425), .dout(n3632));
  jnot g03440(.din(n3632), .dout(n3633));
  jand g03441(.dina(\a[36] ), .dinb(\a[7] ), .dout(n3634));
  jand g03442(.dina(\a[33] ), .dinb(\a[10] ), .dout(n3635));
  jand g03443(.dina(\a[35] ), .dinb(\a[8] ), .dout(n3636));
  jor  g03444(.dina(n3636), .dinb(n3635), .dout(n3637));
  jand g03445(.dina(\a[35] ), .dinb(\a[10] ), .dout(n3638));
  jand g03446(.dina(n3638), .dinb(n3384), .dout(n3639));
  jnot g03447(.din(n3639), .dout(n3640));
  jand g03448(.dina(n3640), .dinb(n3637), .dout(n3641));
  jxor g03449(.dina(n3641), .dinb(n3634), .dout(n3642));
  jxor g03450(.dina(n3642), .dinb(n3633), .dout(n3643));
  jand g03451(.dina(\a[38] ), .dinb(\a[5] ), .dout(n3644));
  jnot g03452(.din(n3644), .dout(n3645));
  jand g03453(.dina(\a[30] ), .dinb(\a[13] ), .dout(n3646));
  jxor g03454(.dina(n3646), .dinb(n3645), .dout(n3647));
  jxor g03455(.dina(n3647), .dinb(n3351), .dout(n3648));
  jnot g03456(.din(n3648), .dout(n3649));
  jxor g03457(.dina(n3649), .dinb(n3643), .dout(n3650));
  jxor g03458(.dina(n3650), .dinb(n3624), .dout(n3651));
  jxor g03459(.dina(n3651), .dinb(n3597), .dout(n3652));
  jxor g03460(.dina(n3652), .dinb(n3593), .dout(n3653));
  jor  g03461(.dina(n3483), .dinb(n3476), .dout(n3654));
  jand g03462(.dina(n3484), .dinb(n3470), .dout(n3655));
  jnot g03463(.din(n3655), .dout(n3656));
  jand g03464(.dina(n3656), .dinb(n3654), .dout(n3657));
  jnot g03465(.din(n3657), .dout(n3658));
  jand g03466(.dina(n3552), .dinb(n3548), .dout(n3659));
  jor  g03467(.dina(n3659), .dinb(n3554), .dout(n3660));
  jand g03468(.dina(n3539), .dinb(n3538), .dout(n3661));
  jnot g03469(.din(n3661), .dout(n3662));
  jnot g03470(.din(n3538), .dout(n3663));
  jnot g03471(.din(n3539), .dout(n3664));
  jand g03472(.dina(n3664), .dinb(n3663), .dout(n3665));
  jor  g03473(.dina(n3665), .dinb(n3537), .dout(n3666));
  jand g03474(.dina(n3666), .dinb(n3662), .dout(n3667));
  jnot g03475(.din(n3667), .dout(n3668));
  jxor g03476(.dina(n3668), .dinb(n3660), .dout(n3669));
  jand g03477(.dina(n3561), .dinb(n3558), .dout(n3670));
  jor  g03478(.dina(n3670), .dinb(n3563), .dout(n3671));
  jxor g03479(.dina(n3671), .dinb(n3669), .dout(n3672));
  jand g03480(.dina(n3474), .dinb(n3473), .dout(n3673));
  jnot g03481(.din(n3673), .dout(n3674));
  jnot g03482(.din(n3473), .dout(n3675));
  jnot g03483(.din(n3474), .dout(n3676));
  jand g03484(.dina(n3676), .dinb(n3675), .dout(n3677));
  jor  g03485(.dina(n3677), .dinb(n3472), .dout(n3678));
  jand g03486(.dina(n3678), .dinb(n3674), .dout(n3679));
  jand g03487(.dina(n3569), .dinb(n3568), .dout(n3680));
  jnot g03488(.din(n3680), .dout(n3681));
  jnot g03489(.din(n3568), .dout(n3682));
  jnot g03490(.din(n3569), .dout(n3683));
  jand g03491(.dina(n3683), .dinb(n3682), .dout(n3684));
  jor  g03492(.dina(n3684), .dinb(n3567), .dout(n3685));
  jand g03493(.dina(n3685), .dinb(n3681), .dout(n3686));
  jxor g03494(.dina(n3686), .dinb(n3679), .dout(n3687));
  jand g03495(.dina(n3477), .dinb(n3308), .dout(n3688));
  jnot g03496(.din(n3688), .dout(n3689));
  jnot g03497(.din(n3477), .dout(n3690));
  jand g03498(.dina(n3690), .dinb(n3309), .dout(n3691));
  jor  g03499(.dina(n3482), .dinb(n3691), .dout(n3692));
  jand g03500(.dina(n3692), .dinb(n3689), .dout(n3693));
  jnot g03501(.din(n3693), .dout(n3694));
  jxor g03502(.dina(n3694), .dinb(n3687), .dout(n3695));
  jxor g03503(.dina(n3695), .dinb(n3672), .dout(n3696));
  jxor g03504(.dina(n3696), .dinb(n3658), .dout(n3697));
  jand g03505(.dina(n3515), .dinb(n3513), .dout(n3698));
  jand g03506(.dina(n3518), .dinb(n3516), .dout(n3699));
  jor  g03507(.dina(n3699), .dinb(n3698), .dout(n3700));
  jand g03508(.dina(n3505), .dinb(n3499), .dout(n3701));
  jand g03509(.dina(n3506), .dinb(n3491), .dout(n3702));
  jor  g03510(.dina(n3702), .dinb(n3701), .dout(n3703));
  jnot g03511(.din(n3703), .dout(n3704));
  jand g03512(.dina(\a[31] ), .dinb(\a[12] ), .dout(n3705));
  jand g03513(.dina(\a[32] ), .dinb(\a[11] ), .dout(n3706));
  jand g03514(.dina(\a[37] ), .dinb(\a[6] ), .dout(n3707));
  jnot g03515(.din(n3707), .dout(n3708));
  jxor g03516(.dina(n3708), .dinb(n3706), .dout(n3709));
  jxor g03517(.dina(n3709), .dinb(n3705), .dout(n3710));
  jxor g03518(.dina(n3710), .dinb(n3704), .dout(n3711));
  jxor g03519(.dina(n3711), .dinb(n3700), .dout(n3712));
  jand g03520(.dina(n3510), .dinb(n3507), .dout(n3713));
  jand g03521(.dina(n3519), .dinb(n3511), .dout(n3714));
  jor  g03522(.dina(n3714), .dinb(n3713), .dout(n3715));
  jxor g03523(.dina(n3715), .dinb(n3712), .dout(n3716));
  jxor g03524(.dina(n3716), .dinb(n3697), .dout(n3717));
  jxor g03525(.dina(n3717), .dinb(n3653), .dout(n3718));
  jand g03526(.dina(n3575), .dinb(n3524), .dout(n3719));
  jand g03527(.dina(n3576), .dinb(n3521), .dout(n3720));
  jor  g03528(.dina(n3720), .dinb(n3719), .dout(n3721));
  jand g03529(.dina(n3488), .dinb(n3485), .dout(n3722));
  jand g03530(.dina(n3520), .dinb(n3489), .dout(n3723));
  jor  g03531(.dina(n3723), .dinb(n3722), .dout(n3724));
  jand g03532(.dina(n3546), .dinb(n3527), .dout(n3725));
  jand g03533(.dina(n3574), .dinb(n3547), .dout(n3726));
  jor  g03534(.dina(n3726), .dinb(n3725), .dout(n3727));
  jand g03535(.dina(n3544), .dinb(n3542), .dout(n3728));
  jand g03536(.dina(n3545), .dinb(n3535), .dout(n3729));
  jor  g03537(.dina(n3729), .dinb(n3728), .dout(n3730));
  jand g03538(.dina(n3480), .dinb(n3479), .dout(n3731));
  jand g03539(.dina(n1207), .dinb(\a[42] ), .dout(n3732));
  jnot g03540(.din(n3732), .dout(n3733));
  jand g03541(.dina(\a[42] ), .dinb(\a[1] ), .dout(n3734));
  jor  g03542(.dina(n3734), .dinb(\a[22] ), .dout(n3735));
  jand g03543(.dina(n3735), .dinb(n3733), .dout(n3736));
  jor  g03544(.dina(n3736), .dinb(n3731), .dout(n3737));
  jnot g03545(.din(\a[42] ), .dout(n3738));
  jand g03546(.dina(n3731), .dinb(n3738), .dout(n3739));
  jnot g03547(.din(n3739), .dout(n3740));
  jand g03548(.dina(n3740), .dinb(n3737), .dout(n3741));
  jand g03549(.dina(n3530), .dinb(n2760), .dout(n3742));
  jor  g03550(.dina(n3742), .dinb(n3532), .dout(n3743));
  jxor g03551(.dina(n3743), .dinb(n3741), .dout(n3744));
  jxor g03552(.dina(n3744), .dinb(n3730), .dout(n3745));
  jnot g03553(.din(n3745), .dout(n3746));
  jnot g03554(.din(n3566), .dout(n3747));
  jand g03555(.dina(n3572), .dinb(n3747), .dout(n3748));
  jnot g03556(.din(n3748), .dout(n3749));
  jand g03557(.dina(n3571), .dinb(n3566), .dout(n3750));
  jor  g03558(.dina(n3750), .dinb(n3557), .dout(n3751));
  jand g03559(.dina(n3751), .dinb(n3749), .dout(n3752));
  jxor g03560(.dina(n3752), .dinb(n3746), .dout(n3753));
  jxor g03561(.dina(n3753), .dinb(n3727), .dout(n3754));
  jxor g03562(.dina(n3754), .dinb(n3724), .dout(n3755));
  jxor g03563(.dina(n3755), .dinb(n3721), .dout(n3756));
  jxor g03564(.dina(n3756), .dinb(n3718), .dout(n3757));
  jxor g03565(.dina(n3757), .dinb(n3590), .dout(n3758));
  jand g03566(.dina(n3578), .dinb(n3442), .dout(n3759));
  jor  g03567(.dina(n3578), .dinb(n3442), .dout(n3760));
  jand g03568(.dina(n3586), .dinb(n3760), .dout(n3761));
  jor  g03569(.dina(n3761), .dinb(n3759), .dout(n3762));
  jxor g03570(.dina(n3762), .dinb(n3758), .dout(\asquared[44] ));
  jand g03571(.dina(n3755), .dinb(n3721), .dout(n3764));
  jand g03572(.dina(n3756), .dinb(n3718), .dout(n3765));
  jor  g03573(.dina(n3765), .dinb(n3764), .dout(n3766));
  jand g03574(.dina(n3652), .dinb(n3593), .dout(n3767));
  jand g03575(.dina(n3717), .dinb(n3653), .dout(n3768));
  jor  g03576(.dina(n3768), .dinb(n3767), .dout(n3769));
  jand g03577(.dina(n3715), .dinb(n3712), .dout(n3770));
  jand g03578(.dina(n3716), .dinb(n3697), .dout(n3771));
  jor  g03579(.dina(n3771), .dinb(n3770), .dout(n3772));
  jand g03580(.dina(n3650), .dinb(n3624), .dout(n3773));
  jand g03581(.dina(n3651), .dinb(n3597), .dout(n3774));
  jor  g03582(.dina(n3774), .dinb(n3773), .dout(n3775));
  jand g03583(.dina(n3619), .dinb(n3618), .dout(n3776));
  jnot g03584(.din(n3776), .dout(n3777));
  jnot g03585(.din(n3618), .dout(n3778));
  jnot g03586(.din(n3619), .dout(n3779));
  jand g03587(.dina(n3779), .dinb(n3778), .dout(n3780));
  jor  g03588(.dina(n3780), .dinb(n3617), .dout(n3781));
  jand g03589(.dina(n3781), .dinb(n3777), .dout(n3782));
  jnot g03590(.din(n3782), .dout(n3783));
  jnot g03591(.din(n3646), .dout(n3784));
  jand g03592(.dina(n3784), .dinb(n3645), .dout(n3785));
  jnot g03593(.din(n3785), .dout(n3786));
  jand g03594(.dina(n3646), .dinb(n3644), .dout(n3787));
  jor  g03595(.dina(n3787), .dinb(n3351), .dout(n3788));
  jand g03596(.dina(n3788), .dinb(n3786), .dout(n3789));
  jxor g03597(.dina(n3789), .dinb(n3783), .dout(n3790));
  jand g03598(.dina(n3601), .dinb(n3598), .dout(n3791));
  jor  g03599(.dina(n3791), .dinb(n3603), .dout(n3792));
  jxor g03600(.dina(n3792), .dinb(n3790), .dout(n3793));
  jnot g03601(.din(n3615), .dout(n3794));
  jand g03602(.dina(n3622), .dinb(n3794), .dout(n3795));
  jnot g03603(.din(n3795), .dout(n3796));
  jand g03604(.dina(n3621), .dinb(n3615), .dout(n3797));
  jor  g03605(.dina(n3797), .dinb(n3606), .dout(n3798));
  jand g03606(.dina(n3798), .dinb(n3796), .dout(n3799));
  jnot g03607(.din(n3799), .dout(n3800));
  jor  g03608(.dina(n3642), .dinb(n3633), .dout(n3801));
  jand g03609(.dina(n3642), .dinb(n3633), .dout(n3802));
  jor  g03610(.dina(n3649), .dinb(n3802), .dout(n3803));
  jand g03611(.dina(n3803), .dinb(n3801), .dout(n3804));
  jxor g03612(.dina(n3804), .dinb(n3800), .dout(n3805));
  jxor g03613(.dina(n3805), .dinb(n3793), .dout(n3806));
  jxor g03614(.dina(n3806), .dinb(n3775), .dout(n3807));
  jxor g03615(.dina(n3807), .dinb(n3772), .dout(n3808));
  jxor g03616(.dina(n3808), .dinb(n3769), .dout(n3809));
  jand g03617(.dina(n3753), .dinb(n3727), .dout(n3810));
  jand g03618(.dina(n3754), .dinb(n3724), .dout(n3811));
  jor  g03619(.dina(n3811), .dinb(n3810), .dout(n3812));
  jand g03620(.dina(n3744), .dinb(n3730), .dout(n3813));
  jnot g03621(.din(n3813), .dout(n3814));
  jor  g03622(.dina(n3752), .dinb(n3746), .dout(n3815));
  jand g03623(.dina(n3815), .dinb(n3814), .dout(n3816));
  jnot g03624(.din(n3816), .dout(n3817));
  jand g03625(.dina(\a[38] ), .dinb(\a[6] ), .dout(n3818));
  jand g03626(.dina(\a[37] ), .dinb(\a[7] ), .dout(n3819));
  jor  g03627(.dina(n3819), .dinb(n2220), .dout(n3820));
  jnot g03628(.din(n3820), .dout(n3821));
  jand g03629(.dina(\a[37] ), .dinb(\a[11] ), .dout(n3822));
  jand g03630(.dina(n3822), .dinb(n3065), .dout(n3823));
  jor  g03631(.dina(n3823), .dinb(n3821), .dout(n3824));
  jxor g03632(.dina(n3824), .dinb(n3818), .dout(n3825));
  jand g03633(.dina(\a[26] ), .dinb(\a[18] ), .dout(n3826));
  jand g03634(.dina(\a[24] ), .dinb(\a[20] ), .dout(n3827));
  jor  g03635(.dina(n3827), .dinb(n3602), .dout(n3828));
  jnot g03636(.din(n3828), .dout(n3829));
  jand g03637(.dina(\a[25] ), .dinb(\a[20] ), .dout(n3830));
  jand g03638(.dina(n3830), .dinb(n3562), .dout(n3831));
  jor  g03639(.dina(n3831), .dinb(n3829), .dout(n3832));
  jxor g03640(.dina(n3832), .dinb(n3826), .dout(n3833));
  jand g03641(.dina(\a[41] ), .dinb(\a[3] ), .dout(n3834));
  jand g03642(.dina(\a[29] ), .dinb(\a[15] ), .dout(n3835));
  jand g03643(.dina(\a[27] ), .dinb(\a[17] ), .dout(n3836));
  jor  g03644(.dina(n3836), .dinb(n3835), .dout(n3837));
  jand g03645(.dina(\a[29] ), .dinb(\a[17] ), .dout(n3838));
  jand g03646(.dina(n3838), .dinb(n3548), .dout(n3839));
  jnot g03647(.din(n3839), .dout(n3840));
  jand g03648(.dina(n3840), .dinb(n3837), .dout(n3841));
  jxor g03649(.dina(n3841), .dinb(n3834), .dout(n3842));
  jxor g03650(.dina(n3842), .dinb(n3833), .dout(n3843));
  jxor g03651(.dina(n3843), .dinb(n3825), .dout(n3844));
  jand g03652(.dina(\a[39] ), .dinb(\a[5] ), .dout(n3845));
  jnot g03653(.din(n3845), .dout(n3846));
  jand g03654(.dina(\a[32] ), .dinb(\a[12] ), .dout(n3847));
  jand g03655(.dina(\a[31] ), .dinb(\a[13] ), .dout(n3848));
  jor  g03656(.dina(n3848), .dinb(n3847), .dout(n3849));
  jand g03657(.dina(\a[32] ), .dinb(\a[13] ), .dout(n3850));
  jand g03658(.dina(n3850), .dinb(n3705), .dout(n3851));
  jnot g03659(.din(n3851), .dout(n3852));
  jand g03660(.dina(n3852), .dinb(n3849), .dout(n3853));
  jxor g03661(.dina(n3853), .dinb(n3846), .dout(n3854));
  jand g03662(.dina(\a[36] ), .dinb(\a[8] ), .dout(n3855));
  jnot g03663(.din(n3855), .dout(n3856));
  jand g03664(.dina(\a[35] ), .dinb(\a[9] ), .dout(n3857));
  jor  g03665(.dina(n3857), .dinb(n3130), .dout(n3858));
  jand g03666(.dina(n3638), .dinb(n3425), .dout(n3859));
  jnot g03667(.din(n3859), .dout(n3860));
  jand g03668(.dina(n3860), .dinb(n3858), .dout(n3861));
  jxor g03669(.dina(n3861), .dinb(n3856), .dout(n3862));
  jnot g03670(.din(n3611), .dout(n3863));
  jand g03671(.dina(\a[40] ), .dinb(\a[4] ), .dout(n3864));
  jand g03672(.dina(\a[30] ), .dinb(\a[14] ), .dout(n3865));
  jxor g03673(.dina(n3865), .dinb(n3864), .dout(n3866));
  jxor g03674(.dina(n3866), .dinb(n3863), .dout(n3867));
  jnot g03675(.din(n3867), .dout(n3868));
  jxor g03676(.dina(n3868), .dinb(n3862), .dout(n3869));
  jxor g03677(.dina(n3869), .dinb(n3854), .dout(n3870));
  jxor g03678(.dina(n3870), .dinb(n3844), .dout(n3871));
  jxor g03679(.dina(n3871), .dinb(n3817), .dout(n3872));
  jxor g03680(.dina(n3872), .dinb(n3812), .dout(n3873));
  jor  g03681(.dina(n3710), .dinb(n3704), .dout(n3874));
  jand g03682(.dina(n3711), .dinb(n3700), .dout(n3875));
  jnot g03683(.din(n3875), .dout(n3876));
  jand g03684(.dina(n3876), .dinb(n3874), .dout(n3877));
  jnot g03685(.din(n3877), .dout(n3878));
  jand g03686(.dina(n3641), .dinb(n3634), .dout(n3879));
  jor  g03687(.dina(n3879), .dinb(n3639), .dout(n3880));
  jand g03688(.dina(\a[43] ), .dinb(\a[1] ), .dout(n3881));
  jxor g03689(.dina(n3881), .dinb(n3629), .dout(n3882));
  jand g03690(.dina(n3627), .dinb(n3425), .dout(n3883));
  jor  g03691(.dina(n3883), .dinb(n3630), .dout(n3884));
  jxor g03692(.dina(n3884), .dinb(n3882), .dout(n3885));
  jxor g03693(.dina(n3885), .dinb(n3880), .dout(n3886));
  jand g03694(.dina(n3610), .dinb(n3607), .dout(n3887));
  jor  g03695(.dina(n3887), .dinb(n3612), .dout(n3888));
  jnot g03696(.din(n3706), .dout(n3889));
  jand g03697(.dina(n3708), .dinb(n3889), .dout(n3890));
  jnot g03698(.din(n3890), .dout(n3891));
  jand g03699(.dina(n3707), .dinb(n3706), .dout(n3892));
  jor  g03700(.dina(n3892), .dinb(n3705), .dout(n3893));
  jand g03701(.dina(n3893), .dinb(n3891), .dout(n3894));
  jxor g03702(.dina(n3894), .dinb(n3888), .dout(n3895));
  jand g03703(.dina(\a[44] ), .dinb(\a[0] ), .dout(n3896));
  jand g03704(.dina(\a[42] ), .dinb(\a[2] ), .dout(n3897));
  jor  g03705(.dina(n3897), .dinb(n3896), .dout(n3898));
  jand g03706(.dina(\a[44] ), .dinb(\a[2] ), .dout(n3899));
  jand g03707(.dina(n3899), .dinb(n3477), .dout(n3900));
  jnot g03708(.din(n3900), .dout(n3901));
  jand g03709(.dina(n3901), .dinb(n3898), .dout(n3902));
  jxor g03710(.dina(n3902), .dinb(n3733), .dout(n3903));
  jnot g03711(.din(n3903), .dout(n3904));
  jxor g03712(.dina(n3904), .dinb(n3895), .dout(n3905));
  jxor g03713(.dina(n3905), .dinb(n3886), .dout(n3906));
  jxor g03714(.dina(n3906), .dinb(n3878), .dout(n3907));
  jand g03715(.dina(n3695), .dinb(n3672), .dout(n3908));
  jand g03716(.dina(n3696), .dinb(n3658), .dout(n3909));
  jor  g03717(.dina(n3909), .dinb(n3908), .dout(n3910));
  jnot g03718(.din(n3679), .dout(n3911));
  jnot g03719(.din(n3686), .dout(n3912));
  jand g03720(.dina(n3912), .dinb(n3911), .dout(n3913));
  jand g03721(.dina(n3694), .dinb(n3687), .dout(n3914));
  jor  g03722(.dina(n3914), .dinb(n3913), .dout(n3915));
  jand g03723(.dina(n3743), .dinb(n3741), .dout(n3916));
  jor  g03724(.dina(n3916), .dinb(n3739), .dout(n3917));
  jxor g03725(.dina(n3917), .dinb(n3915), .dout(n3918));
  jand g03726(.dina(n3668), .dinb(n3660), .dout(n3919));
  jand g03727(.dina(n3671), .dinb(n3669), .dout(n3920));
  jor  g03728(.dina(n3920), .dinb(n3919), .dout(n3921));
  jxor g03729(.dina(n3921), .dinb(n3918), .dout(n3922));
  jxor g03730(.dina(n3922), .dinb(n3910), .dout(n3923));
  jxor g03731(.dina(n3923), .dinb(n3907), .dout(n3924));
  jxor g03732(.dina(n3924), .dinb(n3873), .dout(n3925));
  jxor g03733(.dina(n3925), .dinb(n3809), .dout(n3926));
  jxor g03734(.dina(n3926), .dinb(n3766), .dout(n3927));
  jand g03735(.dina(n3757), .dinb(n3590), .dout(n3928));
  jor  g03736(.dina(n3757), .dinb(n3590), .dout(n3929));
  jand g03737(.dina(n3762), .dinb(n3929), .dout(n3930));
  jor  g03738(.dina(n3930), .dinb(n3928), .dout(n3931));
  jxor g03739(.dina(n3931), .dinb(n3927), .dout(\asquared[45] ));
  jand g03740(.dina(n3808), .dinb(n3769), .dout(n3933));
  jand g03741(.dina(n3925), .dinb(n3809), .dout(n3934));
  jor  g03742(.dina(n3934), .dinb(n3933), .dout(n3935));
  jand g03743(.dina(n3872), .dinb(n3812), .dout(n3936));
  jand g03744(.dina(n3924), .dinb(n3873), .dout(n3937));
  jor  g03745(.dina(n3937), .dinb(n3936), .dout(n3938));
  jand g03746(.dina(n3841), .dinb(n3834), .dout(n3939));
  jor  g03747(.dina(n3939), .dinb(n3839), .dout(n3940));
  jand g03748(.dina(n3898), .dinb(n3732), .dout(n3941));
  jor  g03749(.dina(n3941), .dinb(n3900), .dout(n3942));
  jxor g03750(.dina(n3942), .dinb(n3940), .dout(n3943));
  jand g03751(.dina(n3828), .dinb(n3826), .dout(n3944));
  jor  g03752(.dina(n3944), .dinb(n3831), .dout(n3945));
  jxor g03753(.dina(n3945), .dinb(n3943), .dout(n3946));
  jand g03754(.dina(n3917), .dinb(n3915), .dout(n3947));
  jand g03755(.dina(n3921), .dinb(n3918), .dout(n3948));
  jor  g03756(.dina(n3948), .dinb(n3947), .dout(n3949));
  jxor g03757(.dina(n3949), .dinb(n3946), .dout(n3950));
  jand g03758(.dina(n3881), .dinb(n3629), .dout(n3951));
  jand g03759(.dina(\a[42] ), .dinb(\a[3] ), .dout(n3952));
  jxor g03760(.dina(n3952), .dinb(n3951), .dout(n3953));
  jand g03761(.dina(n1236), .dinb(\a[44] ), .dout(n3954));
  jnot g03762(.din(n3954), .dout(n3955));
  jand g03763(.dina(n3955), .dinb(\a[23] ), .dout(n3956));
  jnot g03764(.din(\a[23] ), .dout(n3957));
  jand g03765(.dina(\a[44] ), .dinb(\a[1] ), .dout(n3958));
  jand g03766(.dina(n3958), .dinb(n3957), .dout(n3959));
  jor  g03767(.dina(n3959), .dinb(n3956), .dout(n3960));
  jxor g03768(.dina(n3960), .dinb(n3953), .dout(n3961));
  jand g03769(.dina(\a[30] ), .dinb(\a[15] ), .dout(n3962));
  jand g03770(.dina(\a[29] ), .dinb(\a[16] ), .dout(n3963));
  jand g03771(.dina(\a[28] ), .dinb(\a[17] ), .dout(n3964));
  jor  g03772(.dina(n3964), .dinb(n3963), .dout(n3965));
  jnot g03773(.din(n3965), .dout(n3966));
  jand g03774(.dina(n3838), .dinb(n3611), .dout(n3967));
  jor  g03775(.dina(n3967), .dinb(n3966), .dout(n3968));
  jxor g03776(.dina(n3968), .dinb(n3962), .dout(n3969));
  jnot g03777(.din(n3969), .dout(n3970));
  jand g03778(.dina(\a[39] ), .dinb(\a[6] ), .dout(n3971));
  jor  g03779(.dina(n3971), .dinb(n2955), .dout(n3972));
  jand g03780(.dina(\a[39] ), .dinb(\a[11] ), .dout(n3973));
  jand g03781(.dina(n3973), .dinb(n3212), .dout(n3974));
  jnot g03782(.din(n3974), .dout(n3975));
  jand g03783(.dina(n3975), .dinb(n3972), .dout(n3976));
  jxor g03784(.dina(n3976), .dinb(n2799), .dout(n3977));
  jxor g03785(.dina(n3977), .dinb(n3970), .dout(n3978));
  jxor g03786(.dina(n3978), .dinb(n3961), .dout(n3979));
  jxor g03787(.dina(n3979), .dinb(n3950), .dout(n3980));
  jand g03788(.dina(n3870), .dinb(n3844), .dout(n3981));
  jand g03789(.dina(n3871), .dinb(n3817), .dout(n3982));
  jor  g03790(.dina(n3982), .dinb(n3981), .dout(n3983));
  jand g03791(.dina(n3922), .dinb(n3910), .dout(n3984));
  jand g03792(.dina(n3923), .dinb(n3907), .dout(n3985));
  jor  g03793(.dina(n3985), .dinb(n3984), .dout(n3986));
  jxor g03794(.dina(n3986), .dinb(n3983), .dout(n3987));
  jxor g03795(.dina(n3987), .dinb(n3980), .dout(n3988));
  jxor g03796(.dina(n3988), .dinb(n3938), .dout(n3989));
  jand g03797(.dina(n3806), .dinb(n3775), .dout(n3990));
  jand g03798(.dina(n3807), .dinb(n3772), .dout(n3991));
  jor  g03799(.dina(n3991), .dinb(n3990), .dout(n3992));
  jand g03800(.dina(n3804), .dinb(n3800), .dout(n3993));
  jand g03801(.dina(n3805), .dinb(n3793), .dout(n3994));
  jor  g03802(.dina(n3994), .dinb(n3993), .dout(n3995));
  jand g03803(.dina(\a[24] ), .dinb(\a[21] ), .dout(n3996));
  jand g03804(.dina(\a[23] ), .dinb(\a[22] ), .dout(n3997));
  jor  g03805(.dina(n3997), .dinb(n3996), .dout(n3998));
  jnot g03806(.din(n3998), .dout(n3999));
  jand g03807(.dina(\a[24] ), .dinb(\a[22] ), .dout(n4000));
  jand g03808(.dina(n4000), .dinb(n3629), .dout(n4001));
  jor  g03809(.dina(n4001), .dinb(n3999), .dout(n4002));
  jxor g03810(.dina(n4002), .dinb(n3638), .dout(n4003));
  jand g03811(.dina(\a[38] ), .dinb(\a[7] ), .dout(n4004));
  jand g03812(.dina(\a[37] ), .dinb(\a[8] ), .dout(n4005));
  jand g03813(.dina(\a[36] ), .dinb(\a[9] ), .dout(n4006));
  jor  g03814(.dina(n4006), .dinb(n4005), .dout(n4007));
  jnot g03815(.din(n4007), .dout(n4008));
  jand g03816(.dina(\a[37] ), .dinb(\a[9] ), .dout(n4009));
  jand g03817(.dina(n4009), .dinb(n3855), .dout(n4010));
  jor  g03818(.dina(n4010), .dinb(n4008), .dout(n4011));
  jxor g03819(.dina(n4011), .dinb(n4004), .dout(n4012));
  jand g03820(.dina(\a[45] ), .dinb(\a[0] ), .dout(n4013));
  jand g03821(.dina(\a[43] ), .dinb(\a[2] ), .dout(n4014));
  jand g03822(.dina(\a[41] ), .dinb(\a[4] ), .dout(n4015));
  jor  g03823(.dina(n4015), .dinb(n4014), .dout(n4016));
  jand g03824(.dina(\a[43] ), .dinb(\a[4] ), .dout(n4017));
  jand g03825(.dina(n4017), .dinb(n3351), .dout(n4018));
  jnot g03826(.din(n4018), .dout(n4019));
  jand g03827(.dina(n4019), .dinb(n4016), .dout(n4020));
  jxor g03828(.dina(n4020), .dinb(n4013), .dout(n4021));
  jxor g03829(.dina(n4021), .dinb(n4012), .dout(n4022));
  jxor g03830(.dina(n4022), .dinb(n4003), .dout(n4023));
  jand g03831(.dina(\a[31] ), .dinb(\a[14] ), .dout(n4024));
  jnot g03832(.din(n4024), .dout(n4025));
  jand g03833(.dina(\a[40] ), .dinb(\a[5] ), .dout(n4026));
  jxor g03834(.dina(n4026), .dinb(n3850), .dout(n4027));
  jxor g03835(.dina(n4027), .dinb(n4025), .dout(n4028));
  jand g03836(.dina(\a[27] ), .dinb(\a[18] ), .dout(n4029));
  jnot g03837(.din(n4029), .dout(n4030));
  jand g03838(.dina(\a[26] ), .dinb(\a[19] ), .dout(n4031));
  jor  g03839(.dina(n4031), .dinb(n3830), .dout(n4032));
  jand g03840(.dina(\a[26] ), .dinb(\a[20] ), .dout(n4033));
  jand g03841(.dina(n4033), .dinb(n3602), .dout(n4034));
  jnot g03842(.din(n4034), .dout(n4035));
  jand g03843(.dina(n4035), .dinb(n4032), .dout(n4036));
  jxor g03844(.dina(n4036), .dinb(n4030), .dout(n4037));
  jand g03845(.dina(n3858), .dinb(n3855), .dout(n4038));
  jor  g03846(.dina(n4038), .dinb(n3859), .dout(n4039));
  jxor g03847(.dina(n4039), .dinb(n4037), .dout(n4040));
  jxor g03848(.dina(n4040), .dinb(n4028), .dout(n4041));
  jxor g03849(.dina(n4041), .dinb(n4023), .dout(n4042));
  jxor g03850(.dina(n4042), .dinb(n3995), .dout(n4043));
  jxor g03851(.dina(n4043), .dinb(n3992), .dout(n4044));
  jand g03852(.dina(n3789), .dinb(n3783), .dout(n4045));
  jand g03853(.dina(n3792), .dinb(n3790), .dout(n4046));
  jor  g03854(.dina(n4046), .dinb(n4045), .dout(n4047));
  jnot g03855(.din(n3888), .dout(n4048));
  jnot g03856(.din(n3894), .dout(n4049));
  jand g03857(.dina(n4049), .dinb(n4048), .dout(n4050));
  jnot g03858(.din(n4050), .dout(n4051));
  jand g03859(.dina(n3894), .dinb(n3888), .dout(n4052));
  jor  g03860(.dina(n3904), .dinb(n4052), .dout(n4053));
  jand g03861(.dina(n4053), .dinb(n4051), .dout(n4054));
  jxor g03862(.dina(n4054), .dinb(n4047), .dout(n4055));
  jand g03863(.dina(n3884), .dinb(n3882), .dout(n4056));
  jand g03864(.dina(n3885), .dinb(n3880), .dout(n4057));
  jor  g03865(.dina(n4057), .dinb(n4056), .dout(n4058));
  jxor g03866(.dina(n4058), .dinb(n4055), .dout(n4059));
  jand g03867(.dina(n3905), .dinb(n3886), .dout(n4060));
  jand g03868(.dina(n3906), .dinb(n3878), .dout(n4061));
  jor  g03869(.dina(n4061), .dinb(n4060), .dout(n4062));
  jxor g03870(.dina(n4062), .dinb(n4059), .dout(n4063));
  jand g03871(.dina(n3820), .dinb(n3818), .dout(n4064));
  jor  g03872(.dina(n4064), .dinb(n3823), .dout(n4065));
  jand g03873(.dina(n3865), .dinb(n3864), .dout(n4066));
  jnot g03874(.din(n4066), .dout(n4067));
  jnot g03875(.din(n3864), .dout(n4068));
  jnot g03876(.din(n3865), .dout(n4069));
  jand g03877(.dina(n4069), .dinb(n4068), .dout(n4070));
  jor  g03878(.dina(n4070), .dinb(n3863), .dout(n4071));
  jand g03879(.dina(n4071), .dinb(n4067), .dout(n4072));
  jnot g03880(.din(n4072), .dout(n4073));
  jxor g03881(.dina(n4073), .dinb(n4065), .dout(n4074));
  jand g03882(.dina(n3849), .dinb(n3845), .dout(n4075));
  jor  g03883(.dina(n4075), .dinb(n3851), .dout(n4076));
  jxor g03884(.dina(n4076), .dinb(n4074), .dout(n4077));
  jnot g03885(.din(n3862), .dout(n4078));
  jand g03886(.dina(n3868), .dinb(n4078), .dout(n4079));
  jnot g03887(.din(n4079), .dout(n4080));
  jand g03888(.dina(n3867), .dinb(n3862), .dout(n4081));
  jor  g03889(.dina(n4081), .dinb(n3854), .dout(n4082));
  jand g03890(.dina(n4082), .dinb(n4080), .dout(n4083));
  jnot g03891(.din(n4083), .dout(n4084));
  jnot g03892(.din(n3833), .dout(n4085));
  jor  g03893(.dina(n3842), .dinb(n4085), .dout(n4086));
  jnot g03894(.din(n3825), .dout(n4087));
  jand g03895(.dina(n3842), .dinb(n4085), .dout(n4088));
  jor  g03896(.dina(n4088), .dinb(n4087), .dout(n4089));
  jand g03897(.dina(n4089), .dinb(n4086), .dout(n4090));
  jxor g03898(.dina(n4090), .dinb(n4084), .dout(n4091));
  jxor g03899(.dina(n4091), .dinb(n4077), .dout(n4092));
  jxor g03900(.dina(n4092), .dinb(n4063), .dout(n4093));
  jxor g03901(.dina(n4093), .dinb(n4044), .dout(n4094));
  jxor g03902(.dina(n4094), .dinb(n3989), .dout(n4095));
  jxor g03903(.dina(n4095), .dinb(n3935), .dout(n4096));
  jand g03904(.dina(n3926), .dinb(n3766), .dout(n4097));
  jor  g03905(.dina(n3926), .dinb(n3766), .dout(n4098));
  jand g03906(.dina(n3931), .dinb(n4098), .dout(n4099));
  jor  g03907(.dina(n4099), .dinb(n4097), .dout(n4100));
  jxor g03908(.dina(n4100), .dinb(n4096), .dout(\asquared[46] ));
  jand g03909(.dina(n3988), .dinb(n3938), .dout(n4102));
  jand g03910(.dina(n4094), .dinb(n3989), .dout(n4103));
  jor  g03911(.dina(n4103), .dinb(n4102), .dout(n4104));
  jand g03912(.dina(n4043), .dinb(n3992), .dout(n4105));
  jand g03913(.dina(n4093), .dinb(n4044), .dout(n4106));
  jor  g03914(.dina(n4106), .dinb(n4105), .dout(n4107));
  jand g03915(.dina(n4062), .dinb(n4059), .dout(n4108));
  jand g03916(.dina(n4092), .dinb(n4063), .dout(n4109));
  jor  g03917(.dina(n4109), .dinb(n4108), .dout(n4110));
  jand g03918(.dina(n4041), .dinb(n4023), .dout(n4111));
  jand g03919(.dina(n4042), .dinb(n3995), .dout(n4112));
  jor  g03920(.dina(n4112), .dinb(n4111), .dout(n4113));
  jxor g03921(.dina(n4113), .dinb(n4110), .dout(n4114));
  jand g03922(.dina(n4073), .dinb(n4065), .dout(n4115));
  jand g03923(.dina(n4076), .dinb(n4074), .dout(n4116));
  jor  g03924(.dina(n4116), .dinb(n4115), .dout(n4117));
  jand g03925(.dina(\a[32] ), .dinb(\a[14] ), .dout(n4118));
  jnot g03926(.din(n4118), .dout(n4119));
  jand g03927(.dina(\a[40] ), .dinb(\a[6] ), .dout(n4120));
  jand g03928(.dina(\a[33] ), .dinb(\a[13] ), .dout(n4121));
  jxor g03929(.dina(n4121), .dinb(n4120), .dout(n4122));
  jxor g03930(.dina(n4122), .dinb(n4119), .dout(n4123));
  jnot g03931(.din(n4123), .dout(n4124));
  jand g03932(.dina(\a[31] ), .dinb(\a[15] ), .dout(n4125));
  jand g03933(.dina(\a[41] ), .dinb(\a[5] ), .dout(n4126));
  jor  g03934(.dina(n4126), .dinb(n4125), .dout(n4127));
  jand g03935(.dina(\a[41] ), .dinb(\a[15] ), .dout(n4128));
  jand g03936(.dina(n4128), .dinb(n2668), .dout(n4129));
  jnot g03937(.din(n4129), .dout(n4130));
  jand g03938(.dina(n4130), .dinb(n4127), .dout(n4131));
  jxor g03939(.dina(n4131), .dinb(n3899), .dout(n4132));
  jxor g03940(.dina(n4132), .dinb(n4124), .dout(n4133));
  jxor g03941(.dina(n4133), .dinb(n4117), .dout(n4134));
  jand g03942(.dina(n3976), .dinb(n2799), .dout(n4135));
  jor  g03943(.dina(n4135), .dinb(n3974), .dout(n4136));
  jand g03944(.dina(n3965), .dinb(n3962), .dout(n4137));
  jor  g03945(.dina(n4137), .dinb(n3967), .dout(n4138));
  jand g03946(.dina(n4032), .dinb(n4029), .dout(n4139));
  jor  g03947(.dina(n4139), .dinb(n4034), .dout(n4140));
  jxor g03948(.dina(n4140), .dinb(n4138), .dout(n4141));
  jxor g03949(.dina(n4141), .dinb(n4136), .dout(n4142));
  jand g03950(.dina(n4054), .dinb(n4047), .dout(n4143));
  jand g03951(.dina(n4058), .dinb(n4055), .dout(n4144));
  jor  g03952(.dina(n4144), .dinb(n4143), .dout(n4145));
  jxor g03953(.dina(n4145), .dinb(n4142), .dout(n4146));
  jxor g03954(.dina(n4146), .dinb(n4134), .dout(n4147));
  jxor g03955(.dina(n4147), .dinb(n4114), .dout(n4148));
  jxor g03956(.dina(n4148), .dinb(n4107), .dout(n4149));
  jxor g03957(.dina(n4149), .dinb(n4104), .dout(n4150));
  jand g03958(.dina(n3986), .dinb(n3983), .dout(n4151));
  jand g03959(.dina(n3987), .dinb(n3980), .dout(n4152));
  jor  g03960(.dina(n4152), .dinb(n4151), .dout(n4153));
  jand g03961(.dina(n4090), .dinb(n4084), .dout(n4154));
  jand g03962(.dina(n4091), .dinb(n4077), .dout(n4155));
  jor  g03963(.dina(n4155), .dinb(n4154), .dout(n4156));
  jand g03964(.dina(\a[34] ), .dinb(\a[12] ), .dout(n4157));
  jand g03965(.dina(\a[39] ), .dinb(\a[7] ), .dout(n4158));
  jand g03966(.dina(\a[38] ), .dinb(\a[8] ), .dout(n4159));
  jor  g03967(.dina(n4159), .dinb(n4158), .dout(n4160));
  jnot g03968(.din(n4160), .dout(n4161));
  jand g03969(.dina(\a[39] ), .dinb(\a[8] ), .dout(n4162));
  jand g03970(.dina(n4162), .dinb(n4004), .dout(n4163));
  jor  g03971(.dina(n4163), .dinb(n4161), .dout(n4164));
  jxor g03972(.dina(n4164), .dinb(n4157), .dout(n4165));
  jnot g03973(.din(n4165), .dout(n4166));
  jand g03974(.dina(n3952), .dinb(n3951), .dout(n4167));
  jand g03975(.dina(n3960), .dinb(n3953), .dout(n4168));
  jor  g03976(.dina(n4168), .dinb(n4167), .dout(n4169));
  jand g03977(.dina(\a[30] ), .dinb(\a[16] ), .dout(n4170));
  jand g03978(.dina(\a[28] ), .dinb(\a[18] ), .dout(n4171));
  jor  g03979(.dina(n4171), .dinb(n3838), .dout(n4172));
  jnot g03980(.din(n4172), .dout(n4173));
  jand g03981(.dina(\a[29] ), .dinb(\a[18] ), .dout(n4174));
  jand g03982(.dina(n4174), .dinb(n3964), .dout(n4175));
  jor  g03983(.dina(n4175), .dinb(n4173), .dout(n4176));
  jxor g03984(.dina(n4176), .dinb(n4170), .dout(n4177));
  jnot g03985(.din(n4177), .dout(n4178));
  jxor g03986(.dina(n4178), .dinb(n4169), .dout(n4179));
  jxor g03987(.dina(n4179), .dinb(n4166), .dout(n4180));
  jand g03988(.dina(\a[27] ), .dinb(\a[19] ), .dout(n4181));
  jnot g03989(.din(n4181), .dout(n4182));
  jand g03990(.dina(\a[25] ), .dinb(\a[21] ), .dout(n4183));
  jor  g03991(.dina(n4183), .dinb(n4033), .dout(n4184));
  jand g03992(.dina(\a[26] ), .dinb(\a[21] ), .dout(n4185));
  jand g03993(.dina(n4185), .dinb(n3830), .dout(n4186));
  jnot g03994(.din(n4186), .dout(n4187));
  jand g03995(.dina(n4187), .dinb(n4184), .dout(n4188));
  jxor g03996(.dina(n4188), .dinb(n4182), .dout(n4189));
  jnot g03997(.din(n4009), .dout(n4190));
  jand g03998(.dina(\a[36] ), .dinb(\a[10] ), .dout(n4191));
  jor  g03999(.dina(n4191), .dinb(n3395), .dout(n4192));
  jand g04000(.dina(\a[36] ), .dinb(\a[11] ), .dout(n4193));
  jand g04001(.dina(n4193), .dinb(n3638), .dout(n4194));
  jnot g04002(.din(n4194), .dout(n4195));
  jand g04003(.dina(n4195), .dinb(n4192), .dout(n4196));
  jxor g04004(.dina(n4196), .dinb(n4190), .dout(n4197));
  jand g04005(.dina(\a[43] ), .dinb(\a[3] ), .dout(n4198));
  jnot g04006(.din(n4198), .dout(n4199));
  jand g04007(.dina(\a[46] ), .dinb(\a[0] ), .dout(n4200));
  jand g04008(.dina(\a[42] ), .dinb(\a[4] ), .dout(n4201));
  jxor g04009(.dina(n4201), .dinb(n4200), .dout(n4202));
  jxor g04010(.dina(n4202), .dinb(n4199), .dout(n4203));
  jnot g04011(.din(n4203), .dout(n4204));
  jxor g04012(.dina(n4204), .dinb(n4197), .dout(n4205));
  jxor g04013(.dina(n4205), .dinb(n4189), .dout(n4206));
  jxor g04014(.dina(n4206), .dinb(n4180), .dout(n4207));
  jxor g04015(.dina(n4207), .dinb(n4156), .dout(n4208));
  jxor g04016(.dina(n4208), .dinb(n4153), .dout(n4209));
  jnot g04017(.din(n4037), .dout(n4210));
  jand g04018(.dina(n4039), .dinb(n4210), .dout(n4211));
  jnot g04019(.din(n4211), .dout(n4212));
  jnot g04020(.din(n4039), .dout(n4213));
  jand g04021(.dina(n4213), .dinb(n4037), .dout(n4214));
  jor  g04022(.dina(n4214), .dinb(n4028), .dout(n4215));
  jand g04023(.dina(n4215), .dinb(n4212), .dout(n4216));
  jnot g04024(.din(n4216), .dout(n4217));
  jnot g04025(.din(n4012), .dout(n4218));
  jor  g04026(.dina(n4021), .dinb(n4218), .dout(n4219));
  jnot g04027(.din(n4003), .dout(n4220));
  jand g04028(.dina(n4021), .dinb(n4218), .dout(n4221));
  jor  g04029(.dina(n4221), .dinb(n4220), .dout(n4222));
  jand g04030(.dina(n4222), .dinb(n4219), .dout(n4223));
  jxor g04031(.dina(n4223), .dinb(n4217), .dout(n4224));
  jand g04032(.dina(n3977), .dinb(n3970), .dout(n4225));
  jand g04033(.dina(n3978), .dinb(n3961), .dout(n4226));
  jor  g04034(.dina(n4226), .dinb(n4225), .dout(n4227));
  jxor g04035(.dina(n4227), .dinb(n4224), .dout(n4228));
  jand g04036(.dina(n3949), .dinb(n3946), .dout(n4229));
  jand g04037(.dina(n3979), .dinb(n3950), .dout(n4230));
  jor  g04038(.dina(n4230), .dinb(n4229), .dout(n4231));
  jand g04039(.dina(n4020), .dinb(n4013), .dout(n4232));
  jor  g04040(.dina(n4232), .dinb(n4018), .dout(n4233));
  jnot g04041(.din(n4233), .dout(n4234));
  jand g04042(.dina(n4026), .dinb(n3850), .dout(n4235));
  jnot g04043(.din(n4235), .dout(n4236));
  jnot g04044(.din(n3850), .dout(n4237));
  jnot g04045(.din(n4026), .dout(n4238));
  jand g04046(.dina(n4238), .dinb(n4237), .dout(n4239));
  jor  g04047(.dina(n4239), .dinb(n4025), .dout(n4240));
  jand g04048(.dina(n4240), .dinb(n4236), .dout(n4241));
  jxor g04049(.dina(n4241), .dinb(n4234), .dout(n4242));
  jand g04050(.dina(n4007), .dinb(n4004), .dout(n4243));
  jor  g04051(.dina(n4243), .dinb(n4010), .dout(n4244));
  jxor g04052(.dina(n4244), .dinb(n4242), .dout(n4245));
  jand g04053(.dina(n3942), .dinb(n3940), .dout(n4246));
  jand g04054(.dina(n3945), .dinb(n3943), .dout(n4247));
  jor  g04055(.dina(n4247), .dinb(n4246), .dout(n4248));
  jand g04056(.dina(n3998), .dinb(n3638), .dout(n4249));
  jor  g04057(.dina(n4249), .dinb(n4001), .dout(n4250));
  jand g04058(.dina(\a[45] ), .dinb(\a[1] ), .dout(n4251));
  jxor g04059(.dina(n4251), .dinb(n4000), .dout(n4252));
  jxor g04060(.dina(n4252), .dinb(n3954), .dout(n4253));
  jxor g04061(.dina(n4253), .dinb(n4250), .dout(n4254));
  jxor g04062(.dina(n4254), .dinb(n4248), .dout(n4255));
  jxor g04063(.dina(n4255), .dinb(n4245), .dout(n4256));
  jxor g04064(.dina(n4256), .dinb(n4231), .dout(n4257));
  jxor g04065(.dina(n4257), .dinb(n4228), .dout(n4258));
  jxor g04066(.dina(n4258), .dinb(n4209), .dout(n4259));
  jxor g04067(.dina(n4259), .dinb(n4150), .dout(n4260));
  jand g04068(.dina(n4095), .dinb(n3935), .dout(n4261));
  jor  g04069(.dina(n4095), .dinb(n3935), .dout(n4262));
  jand g04070(.dina(n4100), .dinb(n4262), .dout(n4263));
  jor  g04071(.dina(n4263), .dinb(n4261), .dout(n4264));
  jxor g04072(.dina(n4264), .dinb(n4260), .dout(\asquared[47] ));
  jand g04073(.dina(n4148), .dinb(n4107), .dout(n4266));
  jand g04074(.dina(n4149), .dinb(n4104), .dout(n4267));
  jor  g04075(.dina(n4267), .dinb(n4266), .dout(n4268));
  jand g04076(.dina(n4113), .dinb(n4110), .dout(n4269));
  jand g04077(.dina(n4147), .dinb(n4114), .dout(n4270));
  jor  g04078(.dina(n4270), .dinb(n4269), .dout(n4271));
  jand g04079(.dina(n4256), .dinb(n4231), .dout(n4272));
  jand g04080(.dina(n4257), .dinb(n4228), .dout(n4273));
  jor  g04081(.dina(n4273), .dinb(n4272), .dout(n4274));
  jxor g04082(.dina(n4274), .dinb(n4271), .dout(n4275));
  jand g04083(.dina(n4131), .dinb(n3899), .dout(n4276));
  jor  g04084(.dina(n4276), .dinb(n4129), .dout(n4277));
  jand g04085(.dina(n4184), .dinb(n4181), .dout(n4278));
  jor  g04086(.dina(n4278), .dinb(n4186), .dout(n4279));
  jxor g04087(.dina(n4279), .dinb(n4277), .dout(n4280));
  jnot g04088(.din(n4280), .dout(n4281));
  jand g04089(.dina(n4201), .dinb(n4200), .dout(n4282));
  jnot g04090(.din(n4282), .dout(n4283));
  jnot g04091(.din(n4200), .dout(n4284));
  jnot g04092(.din(n4201), .dout(n4285));
  jand g04093(.dina(n4285), .dinb(n4284), .dout(n4286));
  jor  g04094(.dina(n4286), .dinb(n4199), .dout(n4287));
  jand g04095(.dina(n4287), .dinb(n4283), .dout(n4288));
  jxor g04096(.dina(n4288), .dinb(n4281), .dout(n4289));
  jnot g04097(.din(n4289), .dout(n4290));
  jnot g04098(.din(n4197), .dout(n4291));
  jand g04099(.dina(n4204), .dinb(n4291), .dout(n4292));
  jnot g04100(.din(n4292), .dout(n4293));
  jand g04101(.dina(n4203), .dinb(n4197), .dout(n4294));
  jor  g04102(.dina(n4294), .dinb(n4189), .dout(n4295));
  jand g04103(.dina(n4295), .dinb(n4293), .dout(n4296));
  jxor g04104(.dina(n4296), .dinb(n4290), .dout(n4297));
  jand g04105(.dina(n4132), .dinb(n4124), .dout(n4298));
  jand g04106(.dina(n4133), .dinb(n4117), .dout(n4299));
  jor  g04107(.dina(n4299), .dinb(n4298), .dout(n4300));
  jxor g04108(.dina(n4300), .dinb(n4297), .dout(n4301));
  jand g04109(.dina(n4206), .dinb(n4180), .dout(n4302));
  jand g04110(.dina(n4207), .dinb(n4156), .dout(n4303));
  jor  g04111(.dina(n4303), .dinb(n4302), .dout(n4304));
  jand g04112(.dina(n4145), .dinb(n4142), .dout(n4305));
  jand g04113(.dina(n4146), .dinb(n4134), .dout(n4306));
  jor  g04114(.dina(n4306), .dinb(n4305), .dout(n4307));
  jxor g04115(.dina(n4307), .dinb(n4304), .dout(n4308));
  jxor g04116(.dina(n4308), .dinb(n4301), .dout(n4309));
  jxor g04117(.dina(n4309), .dinb(n4275), .dout(n4310));
  jand g04118(.dina(n4208), .dinb(n4153), .dout(n4311));
  jand g04119(.dina(n4258), .dinb(n4209), .dout(n4312));
  jor  g04120(.dina(n4312), .dinb(n4311), .dout(n4313));
  jand g04121(.dina(n4140), .dinb(n4138), .dout(n4314));
  jand g04122(.dina(n4141), .dinb(n4136), .dout(n4315));
  jor  g04123(.dina(n4315), .dinb(n4314), .dout(n4316));
  jand g04124(.dina(n4252), .dinb(n3954), .dout(n4317));
  jand g04125(.dina(n4253), .dinb(n4250), .dout(n4318));
  jor  g04126(.dina(n4318), .dinb(n4317), .dout(n4319));
  jand g04127(.dina(\a[34] ), .dinb(\a[13] ), .dout(n4320));
  jand g04128(.dina(\a[35] ), .dinb(\a[12] ), .dout(n4321));
  jand g04129(.dina(\a[40] ), .dinb(\a[7] ), .dout(n4322));
  jor  g04130(.dina(n4322), .dinb(n4321), .dout(n4323));
  jnot g04131(.din(n4323), .dout(n4324));
  jand g04132(.dina(\a[40] ), .dinb(\a[12] ), .dout(n4325));
  jand g04133(.dina(n4325), .dinb(n3538), .dout(n4326));
  jor  g04134(.dina(n4326), .dinb(n4324), .dout(n4327));
  jxor g04135(.dina(n4327), .dinb(n4320), .dout(n4328));
  jnot g04136(.din(n4328), .dout(n4329));
  jxor g04137(.dina(n4329), .dinb(n4319), .dout(n4330));
  jxor g04138(.dina(n4330), .dinb(n4316), .dout(n4331));
  jand g04139(.dina(n4254), .dinb(n4248), .dout(n4332));
  jand g04140(.dina(n4255), .dinb(n4245), .dout(n4333));
  jor  g04141(.dina(n4333), .dinb(n4332), .dout(n4334));
  jxor g04142(.dina(n4334), .dinb(n4331), .dout(n4335));
  jand g04143(.dina(n4223), .dinb(n4217), .dout(n4336));
  jand g04144(.dina(n4227), .dinb(n4224), .dout(n4337));
  jor  g04145(.dina(n4337), .dinb(n4336), .dout(n4338));
  jxor g04146(.dina(n4338), .dinb(n4335), .dout(n4339));
  jand g04147(.dina(n4178), .dinb(n4169), .dout(n4340));
  jand g04148(.dina(n4179), .dinb(n4166), .dout(n4341));
  jor  g04149(.dina(n4341), .dinb(n4340), .dout(n4342));
  jnot g04150(.din(n4342), .dout(n4343));
  jor  g04151(.dina(n4241), .dinb(n4234), .dout(n4344));
  jand g04152(.dina(n4244), .dinb(n4242), .dout(n4345));
  jnot g04153(.din(n4345), .dout(n4346));
  jand g04154(.dina(n4346), .dinb(n4344), .dout(n4347));
  jxor g04155(.dina(n4347), .dinb(n4343), .dout(n4348));
  jand g04156(.dina(\a[46] ), .dinb(\a[1] ), .dout(n4349));
  jor  g04157(.dina(n4349), .dinb(\a[24] ), .dout(n4350));
  jand g04158(.dina(\a[46] ), .dinb(\a[24] ), .dout(n4351));
  jand g04159(.dina(n4351), .dinb(\a[1] ), .dout(n4352));
  jnot g04160(.din(n4352), .dout(n4353));
  jand g04161(.dina(n4353), .dinb(n4350), .dout(n4354));
  jand g04162(.dina(n4192), .dinb(n4009), .dout(n4355));
  jor  g04163(.dina(n4355), .dinb(n4194), .dout(n4356));
  jxor g04164(.dina(n4356), .dinb(n4354), .dout(n4357));
  jand g04165(.dina(n4160), .dinb(n4157), .dout(n4358));
  jor  g04166(.dina(n4358), .dinb(n4163), .dout(n4359));
  jxor g04167(.dina(n4359), .dinb(n4357), .dout(n4360));
  jxor g04168(.dina(n4360), .dinb(n4348), .dout(n4361));
  jand g04169(.dina(n4172), .dinb(n4170), .dout(n4362));
  jor  g04170(.dina(n4362), .dinb(n4175), .dout(n4363));
  jnot g04171(.din(n4363), .dout(n4364));
  jand g04172(.dina(n4121), .dinb(n4120), .dout(n4365));
  jnot g04173(.din(n4365), .dout(n4366));
  jnot g04174(.din(n4120), .dout(n4367));
  jnot g04175(.din(n4121), .dout(n4368));
  jand g04176(.dina(n4368), .dinb(n4367), .dout(n4369));
  jor  g04177(.dina(n4369), .dinb(n4119), .dout(n4370));
  jand g04178(.dina(n4370), .dinb(n4366), .dout(n4371));
  jxor g04179(.dina(n4371), .dinb(n4364), .dout(n4372));
  jand g04180(.dina(\a[44] ), .dinb(\a[3] ), .dout(n4373));
  jand g04181(.dina(\a[32] ), .dinb(\a[15] ), .dout(n4374));
  jor  g04182(.dina(n4374), .dinb(n4017), .dout(n4375));
  jnot g04183(.din(n4375), .dout(n4376));
  jand g04184(.dina(\a[43] ), .dinb(\a[15] ), .dout(n4377));
  jand g04185(.dina(n4377), .dinb(n2652), .dout(n4378));
  jor  g04186(.dina(n4378), .dinb(n4376), .dout(n4379));
  jxor g04187(.dina(n4379), .dinb(n4373), .dout(n4380));
  jnot g04188(.din(n4380), .dout(n4381));
  jxor g04189(.dina(n4381), .dinb(n4372), .dout(n4382));
  jand g04190(.dina(\a[42] ), .dinb(\a[5] ), .dout(n4383));
  jand g04191(.dina(\a[41] ), .dinb(\a[6] ), .dout(n4384));
  jand g04192(.dina(\a[33] ), .dinb(\a[14] ), .dout(n4385));
  jor  g04193(.dina(n4385), .dinb(n4384), .dout(n4386));
  jnot g04194(.din(n4386), .dout(n4387));
  jand g04195(.dina(\a[41] ), .dinb(\a[14] ), .dout(n4388));
  jand g04196(.dina(n4388), .dinb(n3067), .dout(n4389));
  jor  g04197(.dina(n4389), .dinb(n4387), .dout(n4390));
  jxor g04198(.dina(n4390), .dinb(n4383), .dout(n4391));
  jand g04199(.dina(\a[37] ), .dinb(\a[10] ), .dout(n4392));
  jand g04200(.dina(\a[24] ), .dinb(\a[23] ), .dout(n4393));
  jand g04201(.dina(\a[25] ), .dinb(\a[22] ), .dout(n4394));
  jor  g04202(.dina(n4394), .dinb(n4393), .dout(n4395));
  jnot g04203(.din(n4395), .dout(n4396));
  jand g04204(.dina(\a[25] ), .dinb(\a[23] ), .dout(n4397));
  jand g04205(.dina(n4397), .dinb(n4000), .dout(n4398));
  jor  g04206(.dina(n4398), .dinb(n4396), .dout(n4399));
  jxor g04207(.dina(n4399), .dinb(n4392), .dout(n4400));
  jand g04208(.dina(\a[38] ), .dinb(\a[9] ), .dout(n4401));
  jor  g04209(.dina(n4401), .dinb(n4193), .dout(n4402));
  jand g04210(.dina(\a[38] ), .dinb(\a[11] ), .dout(n4403));
  jand g04211(.dina(n4403), .dinb(n4006), .dout(n4404));
  jnot g04212(.din(n4404), .dout(n4405));
  jand g04213(.dina(n4405), .dinb(n4402), .dout(n4406));
  jxor g04214(.dina(n4406), .dinb(n4162), .dout(n4407));
  jxor g04215(.dina(n4407), .dinb(n4400), .dout(n4408));
  jxor g04216(.dina(n4408), .dinb(n4391), .dout(n4409));
  jxor g04217(.dina(n4409), .dinb(n4382), .dout(n4410));
  jand g04218(.dina(\a[28] ), .dinb(\a[19] ), .dout(n4411));
  jnot g04219(.din(n4411), .dout(n4412));
  jand g04220(.dina(\a[27] ), .dinb(\a[20] ), .dout(n4413));
  jor  g04221(.dina(n4413), .dinb(n4185), .dout(n4414));
  jand g04222(.dina(\a[27] ), .dinb(\a[21] ), .dout(n4415));
  jand g04223(.dina(n4415), .dinb(n4033), .dout(n4416));
  jnot g04224(.din(n4416), .dout(n4417));
  jand g04225(.dina(n4417), .dinb(n4414), .dout(n4418));
  jxor g04226(.dina(n4418), .dinb(n4412), .dout(n4419));
  jand g04227(.dina(\a[31] ), .dinb(\a[16] ), .dout(n4420));
  jnot g04228(.din(n4420), .dout(n4421));
  jand g04229(.dina(\a[30] ), .dinb(\a[17] ), .dout(n4422));
  jor  g04230(.dina(n4422), .dinb(n4174), .dout(n4423));
  jand g04231(.dina(\a[30] ), .dinb(\a[18] ), .dout(n4424));
  jand g04232(.dina(n4424), .dinb(n3838), .dout(n4425));
  jnot g04233(.din(n4425), .dout(n4426));
  jand g04234(.dina(n4426), .dinb(n4423), .dout(n4427));
  jxor g04235(.dina(n4427), .dinb(n4421), .dout(n4428));
  jnot g04236(.din(n4428), .dout(n4429));
  jand g04237(.dina(n4251), .dinb(n4000), .dout(n4430));
  jnot g04238(.din(n4430), .dout(n4431));
  jand g04239(.dina(\a[47] ), .dinb(\a[0] ), .dout(n4432));
  jand g04240(.dina(\a[45] ), .dinb(\a[2] ), .dout(n4433));
  jor  g04241(.dina(n4433), .dinb(n4432), .dout(n4434));
  jand g04242(.dina(\a[47] ), .dinb(\a[2] ), .dout(n4435));
  jand g04243(.dina(n4435), .dinb(n4013), .dout(n4436));
  jnot g04244(.din(n4436), .dout(n4437));
  jand g04245(.dina(n4437), .dinb(n4434), .dout(n4438));
  jxor g04246(.dina(n4438), .dinb(n4431), .dout(n4439));
  jxor g04247(.dina(n4439), .dinb(n4429), .dout(n4440));
  jxor g04248(.dina(n4440), .dinb(n4419), .dout(n4441));
  jxor g04249(.dina(n4441), .dinb(n4410), .dout(n4442));
  jxor g04250(.dina(n4442), .dinb(n4361), .dout(n4443));
  jxor g04251(.dina(n4443), .dinb(n4339), .dout(n4444));
  jxor g04252(.dina(n4444), .dinb(n4313), .dout(n4445));
  jxor g04253(.dina(n4445), .dinb(n4310), .dout(n4446));
  jxor g04254(.dina(n4446), .dinb(n4268), .dout(n4447));
  jand g04255(.dina(n4259), .dinb(n4150), .dout(n4448));
  jnot g04256(.din(n4150), .dout(n4449));
  jnot g04257(.din(n4259), .dout(n4450));
  jand g04258(.dina(n4450), .dinb(n4449), .dout(n4451));
  jnot g04259(.din(n4451), .dout(n4452));
  jand g04260(.dina(n4264), .dinb(n4452), .dout(n4453));
  jor  g04261(.dina(n4453), .dinb(n4448), .dout(n4454));
  jxor g04262(.dina(n4454), .dinb(n4447), .dout(\asquared[48] ));
  jand g04263(.dina(n4444), .dinb(n4313), .dout(n4456));
  jand g04264(.dina(n4445), .dinb(n4310), .dout(n4457));
  jor  g04265(.dina(n4457), .dinb(n4456), .dout(n4458));
  jand g04266(.dina(n4274), .dinb(n4271), .dout(n4459));
  jand g04267(.dina(n4309), .dinb(n4275), .dout(n4460));
  jor  g04268(.dina(n4460), .dinb(n4459), .dout(n4461));
  jand g04269(.dina(n4307), .dinb(n4304), .dout(n4462));
  jand g04270(.dina(n4308), .dinb(n4301), .dout(n4463));
  jor  g04271(.dina(n4463), .dinb(n4462), .dout(n4464));
  jand g04272(.dina(n4334), .dinb(n4331), .dout(n4465));
  jand g04273(.dina(n4338), .dinb(n4335), .dout(n4466));
  jor  g04274(.dina(n4466), .dinb(n4465), .dout(n4467));
  jand g04275(.dina(n4329), .dinb(n4319), .dout(n4468));
  jand g04276(.dina(n4330), .dinb(n4316), .dout(n4469));
  jor  g04277(.dina(n4469), .dinb(n4468), .dout(n4470));
  jand g04278(.dina(\a[39] ), .dinb(\a[9] ), .dout(n4471));
  jand g04279(.dina(\a[38] ), .dinb(\a[10] ), .dout(n4472));
  jor  g04280(.dina(n4472), .dinb(n3822), .dout(n4473));
  jnot g04281(.din(n4473), .dout(n4474));
  jand g04282(.dina(n4403), .dinb(n4392), .dout(n4475));
  jor  g04283(.dina(n4475), .dinb(n4474), .dout(n4476));
  jxor g04284(.dina(n4476), .dinb(n4471), .dout(n4477));
  jnot g04285(.din(n4477), .dout(n4478));
  jand g04286(.dina(\a[34] ), .dinb(\a[14] ), .dout(n4479));
  jnot g04287(.din(n4479), .dout(n4480));
  jand g04288(.dina(\a[42] ), .dinb(\a[6] ), .dout(n4481));
  jand g04289(.dina(\a[35] ), .dinb(\a[13] ), .dout(n4482));
  jxor g04290(.dina(n4482), .dinb(n4481), .dout(n4483));
  jxor g04291(.dina(n4483), .dinb(n4480), .dout(n4484));
  jand g04292(.dina(\a[41] ), .dinb(\a[7] ), .dout(n4485));
  jand g04293(.dina(\a[40] ), .dinb(\a[8] ), .dout(n4486));
  jand g04294(.dina(\a[36] ), .dinb(\a[12] ), .dout(n4487));
  jor  g04295(.dina(n4487), .dinb(n4486), .dout(n4488));
  jnot g04296(.din(n4488), .dout(n4489));
  jand g04297(.dina(n4325), .dinb(n3855), .dout(n4490));
  jor  g04298(.dina(n4490), .dinb(n4489), .dout(n4491));
  jxor g04299(.dina(n4491), .dinb(n4485), .dout(n4492));
  jxor g04300(.dina(n4492), .dinb(n4484), .dout(n4493));
  jxor g04301(.dina(n4493), .dinb(n4478), .dout(n4494));
  jxor g04302(.dina(n4494), .dinb(n4470), .dout(n4495));
  jand g04303(.dina(\a[31] ), .dinb(\a[17] ), .dout(n4496));
  jand g04304(.dina(\a[29] ), .dinb(\a[19] ), .dout(n4497));
  jor  g04305(.dina(n4497), .dinb(n4424), .dout(n4498));
  jnot g04306(.din(n4498), .dout(n4499));
  jand g04307(.dina(\a[30] ), .dinb(\a[19] ), .dout(n4500));
  jand g04308(.dina(n4500), .dinb(n4174), .dout(n4501));
  jor  g04309(.dina(n4501), .dinb(n4499), .dout(n4502));
  jxor g04310(.dina(n4502), .dinb(n4496), .dout(n4503));
  jand g04311(.dina(\a[28] ), .dinb(\a[20] ), .dout(n4504));
  jand g04312(.dina(\a[26] ), .dinb(\a[22] ), .dout(n4505));
  jor  g04313(.dina(n4505), .dinb(n4415), .dout(n4506));
  jnot g04314(.din(n4506), .dout(n4507));
  jand g04315(.dina(\a[27] ), .dinb(\a[22] ), .dout(n4508));
  jand g04316(.dina(n4508), .dinb(n4185), .dout(n4509));
  jor  g04317(.dina(n4509), .dinb(n4507), .dout(n4510));
  jxor g04318(.dina(n4510), .dinb(n4504), .dout(n4511));
  jand g04319(.dina(\a[44] ), .dinb(\a[4] ), .dout(n4512));
  jand g04320(.dina(\a[43] ), .dinb(\a[5] ), .dout(n4513));
  jand g04321(.dina(\a[33] ), .dinb(\a[15] ), .dout(n4514));
  jor  g04322(.dina(n4514), .dinb(n4513), .dout(n4515));
  jand g04323(.dina(n4377), .dinb(n2895), .dout(n4516));
  jnot g04324(.din(n4516), .dout(n4517));
  jand g04325(.dina(n4517), .dinb(n4515), .dout(n4518));
  jxor g04326(.dina(n4518), .dinb(n4512), .dout(n4519));
  jxor g04327(.dina(n4519), .dinb(n4511), .dout(n4520));
  jxor g04328(.dina(n4520), .dinb(n4503), .dout(n4521));
  jxor g04329(.dina(n4521), .dinb(n4495), .dout(n4522));
  jxor g04330(.dina(n4522), .dinb(n4467), .dout(n4523));
  jxor g04331(.dina(n4523), .dinb(n4464), .dout(n4524));
  jxor g04332(.dina(n4524), .dinb(n4461), .dout(n4525));
  jand g04333(.dina(n4406), .dinb(n4162), .dout(n4526));
  jor  g04334(.dina(n4526), .dinb(n4404), .dout(n4527));
  jand g04335(.dina(n4414), .dinb(n4411), .dout(n4528));
  jor  g04336(.dina(n4528), .dinb(n4416), .dout(n4529));
  jxor g04337(.dina(n4529), .dinb(n4527), .dout(n4530));
  jand g04338(.dina(n4386), .dinb(n4383), .dout(n4531));
  jor  g04339(.dina(n4531), .dinb(n4389), .dout(n4532));
  jxor g04340(.dina(n4532), .dinb(n4530), .dout(n4533));
  jnot g04341(.din(n4400), .dout(n4534));
  jor  g04342(.dina(n4407), .dinb(n4534), .dout(n4535));
  jnot g04343(.din(n4391), .dout(n4536));
  jand g04344(.dina(n4407), .dinb(n4534), .dout(n4537));
  jor  g04345(.dina(n4537), .dinb(n4536), .dout(n4538));
  jand g04346(.dina(n4538), .dinb(n4535), .dout(n4539));
  jxor g04347(.dina(n4539), .dinb(n4533), .dout(n4540));
  jand g04348(.dina(n4323), .dinb(n4320), .dout(n4541));
  jor  g04349(.dina(n4541), .dinb(n4326), .dout(n4542));
  jand g04350(.dina(n4395), .dinb(n4392), .dout(n4543));
  jor  g04351(.dina(n4543), .dinb(n4398), .dout(n4544));
  jxor g04352(.dina(n4544), .dinb(n4542), .dout(n4545));
  jand g04353(.dina(\a[46] ), .dinb(\a[2] ), .dout(n4546));
  jnot g04354(.din(n4546), .dout(n4547));
  jand g04355(.dina(\a[45] ), .dinb(\a[3] ), .dout(n4548));
  jand g04356(.dina(\a[32] ), .dinb(\a[16] ), .dout(n4549));
  jxor g04357(.dina(n4549), .dinb(n4548), .dout(n4550));
  jxor g04358(.dina(n4550), .dinb(n4547), .dout(n4551));
  jnot g04359(.din(n4551), .dout(n4552));
  jxor g04360(.dina(n4552), .dinb(n4545), .dout(n4553));
  jxor g04361(.dina(n4553), .dinb(n4540), .dout(n4554));
  jand g04362(.dina(n4409), .dinb(n4382), .dout(n4555));
  jand g04363(.dina(n4441), .dinb(n4410), .dout(n4556));
  jor  g04364(.dina(n4556), .dinb(n4555), .dout(n4557));
  jxor g04365(.dina(n4557), .dinb(n4554), .dout(n4558));
  jand g04366(.dina(n4423), .dinb(n4420), .dout(n4559));
  jor  g04367(.dina(n4559), .dinb(n4425), .dout(n4560));
  jand g04368(.dina(n4375), .dinb(n4373), .dout(n4561));
  jor  g04369(.dina(n4561), .dinb(n4378), .dout(n4562));
  jxor g04370(.dina(n4562), .dinb(n4560), .dout(n4563));
  jand g04371(.dina(n4434), .dinb(n4430), .dout(n4564));
  jor  g04372(.dina(n4564), .dinb(n4436), .dout(n4565));
  jxor g04373(.dina(n4565), .dinb(n4563), .dout(n4566));
  jand g04374(.dina(n4356), .dinb(n4354), .dout(n4567));
  jand g04375(.dina(n4359), .dinb(n4357), .dout(n4568));
  jor  g04376(.dina(n4568), .dinb(n4567), .dout(n4569));
  jnot g04377(.din(n4569), .dout(n4570));
  jnot g04378(.din(n4439), .dout(n4571));
  jand g04379(.dina(n4571), .dinb(n4429), .dout(n4572));
  jnot g04380(.din(n4572), .dout(n4573));
  jand g04381(.dina(n4439), .dinb(n4428), .dout(n4574));
  jor  g04382(.dina(n4574), .dinb(n4419), .dout(n4575));
  jand g04383(.dina(n4575), .dinb(n4573), .dout(n4576));
  jxor g04384(.dina(n4576), .dinb(n4570), .dout(n4577));
  jxor g04385(.dina(n4577), .dinb(n4566), .dout(n4578));
  jxor g04386(.dina(n4578), .dinb(n4558), .dout(n4579));
  jand g04387(.dina(n4442), .dinb(n4361), .dout(n4580));
  jand g04388(.dina(n4443), .dinb(n4339), .dout(n4581));
  jor  g04389(.dina(n4581), .dinb(n4580), .dout(n4582));
  jor  g04390(.dina(n4296), .dinb(n4290), .dout(n4583));
  jand g04391(.dina(n4300), .dinb(n4297), .dout(n4584));
  jnot g04392(.din(n4584), .dout(n4585));
  jand g04393(.dina(n4585), .dinb(n4583), .dout(n4586));
  jor  g04394(.dina(n4347), .dinb(n4343), .dout(n4587));
  jand g04395(.dina(n4360), .dinb(n4348), .dout(n4588));
  jnot g04396(.din(n4588), .dout(n4589));
  jand g04397(.dina(n4589), .dinb(n4587), .dout(n4590));
  jxor g04398(.dina(n4590), .dinb(n4586), .dout(n4591));
  jand g04399(.dina(n4279), .dinb(n4277), .dout(n4592));
  jnot g04400(.din(n4592), .dout(n4593));
  jor  g04401(.dina(n4288), .dinb(n4281), .dout(n4594));
  jand g04402(.dina(n4594), .dinb(n4593), .dout(n4595));
  jand g04403(.dina(\a[48] ), .dinb(\a[0] ), .dout(n4596));
  jxor g04404(.dina(n4596), .dinb(n4352), .dout(n4597));
  jand g04405(.dina(\a[47] ), .dinb(\a[1] ), .dout(n4598));
  jxor g04406(.dina(n4598), .dinb(n4397), .dout(n4599));
  jnot g04407(.din(n4599), .dout(n4600));
  jxor g04408(.dina(n4600), .dinb(n4597), .dout(n4601));
  jxor g04409(.dina(n4601), .dinb(n4595), .dout(n4602));
  jand g04410(.dina(n4371), .dinb(n4364), .dout(n4603));
  jnot g04411(.din(n4603), .dout(n4604));
  jnot g04412(.din(n4371), .dout(n4605));
  jand g04413(.dina(n4605), .dinb(n4363), .dout(n4606));
  jor  g04414(.dina(n4381), .dinb(n4606), .dout(n4607));
  jand g04415(.dina(n4607), .dinb(n4604), .dout(n4608));
  jxor g04416(.dina(n4608), .dinb(n4602), .dout(n4609));
  jxor g04417(.dina(n4609), .dinb(n4591), .dout(n4610));
  jxor g04418(.dina(n4610), .dinb(n4582), .dout(n4611));
  jxor g04419(.dina(n4611), .dinb(n4579), .dout(n4612));
  jxor g04420(.dina(n4612), .dinb(n4525), .dout(n4613));
  jxor g04421(.dina(n4613), .dinb(n4458), .dout(n4614));
  jand g04422(.dina(n4446), .dinb(n4268), .dout(n4615));
  jor  g04423(.dina(n4446), .dinb(n4268), .dout(n4616));
  jand g04424(.dina(n4454), .dinb(n4616), .dout(n4617));
  jor  g04425(.dina(n4617), .dinb(n4615), .dout(n4618));
  jxor g04426(.dina(n4618), .dinb(n4614), .dout(\asquared[49] ));
  jand g04427(.dina(n4610), .dinb(n4582), .dout(n4620));
  jand g04428(.dina(n4611), .dinb(n4579), .dout(n4621));
  jor  g04429(.dina(n4621), .dinb(n4620), .dout(n4622));
  jand g04430(.dina(n4557), .dinb(n4554), .dout(n4623));
  jand g04431(.dina(n4578), .dinb(n4558), .dout(n4624));
  jor  g04432(.dina(n4624), .dinb(n4623), .dout(n4625));
  jor  g04433(.dina(n4590), .dinb(n4586), .dout(n4626));
  jand g04434(.dina(n4609), .dinb(n4591), .dout(n4627));
  jnot g04435(.din(n4627), .dout(n4628));
  jand g04436(.dina(n4628), .dinb(n4626), .dout(n4629));
  jnot g04437(.din(n4629), .dout(n4630));
  jand g04438(.dina(\a[33] ), .dinb(\a[16] ), .dout(n4631));
  jand g04439(.dina(\a[32] ), .dinb(\a[17] ), .dout(n4632));
  jand g04440(.dina(\a[31] ), .dinb(\a[18] ), .dout(n4633));
  jor  g04441(.dina(n4633), .dinb(n4632), .dout(n4634));
  jnot g04442(.din(n4634), .dout(n4635));
  jand g04443(.dina(\a[32] ), .dinb(\a[18] ), .dout(n4636));
  jand g04444(.dina(n4636), .dinb(n4496), .dout(n4637));
  jor  g04445(.dina(n4637), .dinb(n4635), .dout(n4638));
  jxor g04446(.dina(n4638), .dinb(n4631), .dout(n4639));
  jnot g04447(.din(n4639), .dout(n4640));
  jand g04448(.dina(\a[49] ), .dinb(\a[0] ), .dout(n4641));
  jnot g04449(.din(n4641), .dout(n4642));
  jand g04450(.dina(\a[45] ), .dinb(\a[4] ), .dout(n4643));
  jand g04451(.dina(\a[44] ), .dinb(\a[5] ), .dout(n4644));
  jor  g04452(.dina(n4644), .dinb(n4643), .dout(n4645));
  jand g04453(.dina(\a[45] ), .dinb(\a[5] ), .dout(n4646));
  jand g04454(.dina(n4646), .dinb(n4512), .dout(n4647));
  jnot g04455(.din(n4647), .dout(n4648));
  jand g04456(.dina(n4648), .dinb(n4645), .dout(n4649));
  jxor g04457(.dina(n4649), .dinb(n4642), .dout(n4650));
  jand g04458(.dina(n4596), .dinb(n4352), .dout(n4651));
  jnot g04459(.din(n4651), .dout(n4652));
  jnot g04460(.din(n4596), .dout(n4653));
  jand g04461(.dina(n4653), .dinb(n4353), .dout(n4654));
  jor  g04462(.dina(n4600), .dinb(n4654), .dout(n4655));
  jand g04463(.dina(n4655), .dinb(n4652), .dout(n4656));
  jxor g04464(.dina(n4656), .dinb(n4650), .dout(n4657));
  jxor g04465(.dina(n4657), .dinb(n4640), .dout(n4658));
  jand g04466(.dina(\a[40] ), .dinb(\a[9] ), .dout(n4659));
  jand g04467(.dina(\a[37] ), .dinb(\a[12] ), .dout(n4660));
  jand g04468(.dina(\a[39] ), .dinb(\a[10] ), .dout(n4661));
  jor  g04469(.dina(n4661), .dinb(n4660), .dout(n4662));
  jnot g04470(.din(n4662), .dout(n4663));
  jand g04471(.dina(\a[39] ), .dinb(\a[12] ), .dout(n4664));
  jand g04472(.dina(n4664), .dinb(n4392), .dout(n4665));
  jor  g04473(.dina(n4665), .dinb(n4663), .dout(n4666));
  jxor g04474(.dina(n4666), .dinb(n4659), .dout(n4667));
  jand g04475(.dina(\a[29] ), .dinb(\a[20] ), .dout(n4668));
  jand g04476(.dina(\a[28] ), .dinb(\a[21] ), .dout(n4669));
  jor  g04477(.dina(n4669), .dinb(n4668), .dout(n4670));
  jnot g04478(.din(n4670), .dout(n4671));
  jand g04479(.dina(\a[29] ), .dinb(\a[21] ), .dout(n4672));
  jand g04480(.dina(n4672), .dinb(n4504), .dout(n4673));
  jor  g04481(.dina(n4673), .dinb(n4671), .dout(n4674));
  jxor g04482(.dina(n4674), .dinb(n4500), .dout(n4675));
  jand g04483(.dina(\a[46] ), .dinb(\a[3] ), .dout(n4676));
  jor  g04484(.dina(n4676), .dinb(n4435), .dout(n4677));
  jand g04485(.dina(\a[47] ), .dinb(\a[3] ), .dout(n4678));
  jand g04486(.dina(n4678), .dinb(n4546), .dout(n4679));
  jnot g04487(.din(n4679), .dout(n4680));
  jand g04488(.dina(n4680), .dinb(n4677), .dout(n4681));
  jxor g04489(.dina(n4681), .dinb(n4508), .dout(n4682));
  jxor g04490(.dina(n4682), .dinb(n4675), .dout(n4683));
  jxor g04491(.dina(n4683), .dinb(n4667), .dout(n4684));
  jxor g04492(.dina(n4684), .dinb(n4658), .dout(n4685));
  jand g04493(.dina(\a[34] ), .dinb(\a[15] ), .dout(n4686));
  jand g04494(.dina(\a[43] ), .dinb(\a[6] ), .dout(n4687));
  jand g04495(.dina(\a[35] ), .dinb(\a[14] ), .dout(n4688));
  jor  g04496(.dina(n4688), .dinb(n4687), .dout(n4689));
  jnot g04497(.din(n4689), .dout(n4690));
  jand g04498(.dina(\a[43] ), .dinb(\a[14] ), .dout(n4691));
  jand g04499(.dina(n4691), .dinb(n3392), .dout(n4692));
  jor  g04500(.dina(n4692), .dinb(n4690), .dout(n4693));
  jxor g04501(.dina(n4693), .dinb(n4686), .dout(n4694));
  jnot g04502(.din(n4694), .dout(n4695));
  jand g04503(.dina(\a[25] ), .dinb(\a[24] ), .dout(n4696));
  jnot g04504(.din(n4696), .dout(n4697));
  jand g04505(.dina(\a[26] ), .dinb(\a[23] ), .dout(n4698));
  jxor g04506(.dina(n4698), .dinb(n4697), .dout(n4699));
  jxor g04507(.dina(n4699), .dinb(n4403), .dout(n4700));
  jnot g04508(.din(n4700), .dout(n4701));
  jand g04509(.dina(\a[36] ), .dinb(\a[13] ), .dout(n4702));
  jand g04510(.dina(\a[42] ), .dinb(\a[7] ), .dout(n4703));
  jand g04511(.dina(\a[41] ), .dinb(\a[8] ), .dout(n4704));
  jor  g04512(.dina(n4704), .dinb(n4703), .dout(n4705));
  jand g04513(.dina(\a[42] ), .dinb(\a[8] ), .dout(n4706));
  jand g04514(.dina(n4706), .dinb(n4485), .dout(n4707));
  jnot g04515(.din(n4707), .dout(n4708));
  jand g04516(.dina(n4708), .dinb(n4705), .dout(n4709));
  jxor g04517(.dina(n4709), .dinb(n4702), .dout(n4710));
  jxor g04518(.dina(n4710), .dinb(n4701), .dout(n4711));
  jxor g04519(.dina(n4711), .dinb(n4695), .dout(n4712));
  jxor g04520(.dina(n4712), .dinb(n4685), .dout(n4713));
  jxor g04521(.dina(n4713), .dinb(n4630), .dout(n4714));
  jxor g04522(.dina(n4714), .dinb(n4625), .dout(n4715));
  jxor g04523(.dina(n4715), .dinb(n4622), .dout(n4716));
  jand g04524(.dina(n4498), .dinb(n4496), .dout(n4717));
  jor  g04525(.dina(n4717), .dinb(n4501), .dout(n4718));
  jand g04526(.dina(n4482), .dinb(n4481), .dout(n4719));
  jnot g04527(.din(n4719), .dout(n4720));
  jnot g04528(.din(n4481), .dout(n4721));
  jnot g04529(.din(n4482), .dout(n4722));
  jand g04530(.dina(n4722), .dinb(n4721), .dout(n4723));
  jor  g04531(.dina(n4723), .dinb(n4480), .dout(n4724));
  jand g04532(.dina(n4724), .dinb(n4720), .dout(n4725));
  jnot g04533(.din(n4725), .dout(n4726));
  jxor g04534(.dina(n4726), .dinb(n4718), .dout(n4727));
  jand g04535(.dina(n4488), .dinb(n4485), .dout(n4728));
  jor  g04536(.dina(n4728), .dinb(n4490), .dout(n4729));
  jxor g04537(.dina(n4729), .dinb(n4727), .dout(n4730));
  jnot g04538(.din(n4511), .dout(n4731));
  jor  g04539(.dina(n4519), .dinb(n4731), .dout(n4732));
  jnot g04540(.din(n4503), .dout(n4733));
  jand g04541(.dina(n4519), .dinb(n4731), .dout(n4734));
  jor  g04542(.dina(n4734), .dinb(n4733), .dout(n4735));
  jand g04543(.dina(n4735), .dinb(n4732), .dout(n4736));
  jxor g04544(.dina(n4736), .dinb(n4730), .dout(n4737));
  jnot g04545(.din(n4737), .dout(n4738));
  jor  g04546(.dina(n4601), .dinb(n4595), .dout(n4739));
  jand g04547(.dina(n4608), .dinb(n4602), .dout(n4740));
  jnot g04548(.din(n4740), .dout(n4741));
  jand g04549(.dina(n4741), .dinb(n4739), .dout(n4742));
  jxor g04550(.dina(n4742), .dinb(n4738), .dout(n4743));
  jand g04551(.dina(n4494), .dinb(n4470), .dout(n4744));
  jand g04552(.dina(n4521), .dinb(n4495), .dout(n4745));
  jor  g04553(.dina(n4745), .dinb(n4744), .dout(n4746));
  jxor g04554(.dina(n4746), .dinb(n4743), .dout(n4747));
  jand g04555(.dina(n4518), .dinb(n4512), .dout(n4748));
  jor  g04556(.dina(n4748), .dinb(n4516), .dout(n4749));
  jnot g04557(.din(n4749), .dout(n4750));
  jand g04558(.dina(n4549), .dinb(n4548), .dout(n4751));
  jnot g04559(.din(n4751), .dout(n4752));
  jnot g04560(.din(n4548), .dout(n4753));
  jnot g04561(.din(n4549), .dout(n4754));
  jand g04562(.dina(n4754), .dinb(n4753), .dout(n4755));
  jor  g04563(.dina(n4755), .dinb(n4547), .dout(n4756));
  jand g04564(.dina(n4756), .dinb(n4752), .dout(n4757));
  jxor g04565(.dina(n4757), .dinb(n4750), .dout(n4758));
  jand g04566(.dina(n4506), .dinb(n4504), .dout(n4759));
  jor  g04567(.dina(n4759), .dinb(n4509), .dout(n4760));
  jxor g04568(.dina(n4760), .dinb(n4758), .dout(n4761));
  jor  g04569(.dina(n4492), .dinb(n4484), .dout(n4762));
  jand g04570(.dina(n4493), .dinb(n4478), .dout(n4763));
  jnot g04571(.din(n4763), .dout(n4764));
  jand g04572(.dina(n4764), .dinb(n4762), .dout(n4765));
  jnot g04573(.din(n4765), .dout(n4766));
  jand g04574(.dina(n4598), .dinb(n4397), .dout(n4767));
  jand g04575(.dina(n1424), .dinb(\a[48] ), .dout(n4768));
  jnot g04576(.din(n4768), .dout(n4769));
  jand g04577(.dina(\a[48] ), .dinb(\a[1] ), .dout(n4770));
  jor  g04578(.dina(n4770), .dinb(\a[25] ), .dout(n4771));
  jand g04579(.dina(n4771), .dinb(n4769), .dout(n4772));
  jor  g04580(.dina(n4772), .dinb(n4767), .dout(n4773));
  jnot g04581(.din(\a[48] ), .dout(n4774));
  jand g04582(.dina(n4767), .dinb(n4774), .dout(n4775));
  jnot g04583(.din(n4775), .dout(n4776));
  jand g04584(.dina(n4776), .dinb(n4773), .dout(n4777));
  jand g04585(.dina(n4473), .dinb(n4471), .dout(n4778));
  jor  g04586(.dina(n4778), .dinb(n4475), .dout(n4779));
  jxor g04587(.dina(n4779), .dinb(n4777), .dout(n4780));
  jxor g04588(.dina(n4780), .dinb(n4766), .dout(n4781));
  jxor g04589(.dina(n4781), .dinb(n4761), .dout(n4782));
  jxor g04590(.dina(n4782), .dinb(n4747), .dout(n4783));
  jand g04591(.dina(n4522), .dinb(n4467), .dout(n4784));
  jand g04592(.dina(n4523), .dinb(n4464), .dout(n4785));
  jor  g04593(.dina(n4785), .dinb(n4784), .dout(n4786));
  jand g04594(.dina(n4529), .dinb(n4527), .dout(n4787));
  jand g04595(.dina(n4532), .dinb(n4530), .dout(n4788));
  jor  g04596(.dina(n4788), .dinb(n4787), .dout(n4789));
  jnot g04597(.din(n4542), .dout(n4790));
  jnot g04598(.din(n4544), .dout(n4791));
  jand g04599(.dina(n4791), .dinb(n4790), .dout(n4792));
  jnot g04600(.din(n4792), .dout(n4793));
  jand g04601(.dina(n4544), .dinb(n4542), .dout(n4794));
  jor  g04602(.dina(n4552), .dinb(n4794), .dout(n4795));
  jand g04603(.dina(n4795), .dinb(n4793), .dout(n4796));
  jxor g04604(.dina(n4796), .dinb(n4789), .dout(n4797));
  jand g04605(.dina(n4562), .dinb(n4560), .dout(n4798));
  jand g04606(.dina(n4565), .dinb(n4563), .dout(n4799));
  jor  g04607(.dina(n4799), .dinb(n4798), .dout(n4800));
  jxor g04608(.dina(n4800), .dinb(n4797), .dout(n4801));
  jand g04609(.dina(n4539), .dinb(n4533), .dout(n4802));
  jand g04610(.dina(n4553), .dinb(n4540), .dout(n4803));
  jor  g04611(.dina(n4803), .dinb(n4802), .dout(n4804));
  jnot g04612(.din(n4804), .dout(n4805));
  jor  g04613(.dina(n4576), .dinb(n4570), .dout(n4806));
  jand g04614(.dina(n4577), .dinb(n4566), .dout(n4807));
  jnot g04615(.din(n4807), .dout(n4808));
  jand g04616(.dina(n4808), .dinb(n4806), .dout(n4809));
  jxor g04617(.dina(n4809), .dinb(n4805), .dout(n4810));
  jxor g04618(.dina(n4810), .dinb(n4801), .dout(n4811));
  jxor g04619(.dina(n4811), .dinb(n4786), .dout(n4812));
  jxor g04620(.dina(n4812), .dinb(n4783), .dout(n4813));
  jxor g04621(.dina(n4813), .dinb(n4716), .dout(n4814));
  jand g04622(.dina(n4524), .dinb(n4461), .dout(n4815));
  jand g04623(.dina(n4612), .dinb(n4525), .dout(n4816));
  jor  g04624(.dina(n4816), .dinb(n4815), .dout(n4817));
  jxor g04625(.dina(n4817), .dinb(n4814), .dout(n4818));
  jand g04626(.dina(n4613), .dinb(n4458), .dout(n4819));
  jnot g04627(.din(n4458), .dout(n4820));
  jnot g04628(.din(n4613), .dout(n4821));
  jand g04629(.dina(n4821), .dinb(n4820), .dout(n4822));
  jnot g04630(.din(n4822), .dout(n4823));
  jand g04631(.dina(n4618), .dinb(n4823), .dout(n4824));
  jor  g04632(.dina(n4824), .dinb(n4819), .dout(n4825));
  jxor g04633(.dina(n4825), .dinb(n4818), .dout(\asquared[50] ));
  jand g04634(.dina(n4715), .dinb(n4622), .dout(n4827));
  jand g04635(.dina(n4813), .dinb(n4716), .dout(n4828));
  jor  g04636(.dina(n4828), .dinb(n4827), .dout(n4829));
  jand g04637(.dina(n4811), .dinb(n4786), .dout(n4830));
  jand g04638(.dina(n4812), .dinb(n4783), .dout(n4831));
  jor  g04639(.dina(n4831), .dinb(n4830), .dout(n4832));
  jand g04640(.dina(n4746), .dinb(n4743), .dout(n4833));
  jand g04641(.dina(n4782), .dinb(n4747), .dout(n4834));
  jor  g04642(.dina(n4834), .dinb(n4833), .dout(n4835));
  jor  g04643(.dina(n4809), .dinb(n4805), .dout(n4836));
  jand g04644(.dina(n4810), .dinb(n4801), .dout(n4837));
  jnot g04645(.din(n4837), .dout(n4838));
  jand g04646(.dina(n4838), .dinb(n4836), .dout(n4839));
  jnot g04647(.din(n4839), .dout(n4840));
  jand g04648(.dina(n4779), .dinb(n4777), .dout(n4841));
  jor  g04649(.dina(n4841), .dinb(n4775), .dout(n4842));
  jand g04650(.dina(\a[28] ), .dinb(\a[22] ), .dout(n4843));
  jnot g04651(.din(n4843), .dout(n4844));
  jand g04652(.dina(\a[27] ), .dinb(\a[23] ), .dout(n4845));
  jxor g04653(.dina(n4845), .dinb(n4636), .dout(n4846));
  jxor g04654(.dina(n4846), .dinb(n4844), .dout(n4847));
  jnot g04655(.din(n4847), .dout(n4848));
  jand g04656(.dina(\a[34] ), .dinb(\a[16] ), .dout(n4849));
  jand g04657(.dina(\a[35] ), .dinb(\a[15] ), .dout(n4850));
  jor  g04658(.dina(n4850), .dinb(n4646), .dout(n4851));
  jand g04659(.dina(\a[45] ), .dinb(\a[15] ), .dout(n4852));
  jand g04660(.dina(n4852), .dinb(n3163), .dout(n4853));
  jnot g04661(.din(n4853), .dout(n4854));
  jand g04662(.dina(n4854), .dinb(n4851), .dout(n4855));
  jxor g04663(.dina(n4855), .dinb(n4849), .dout(n4856));
  jxor g04664(.dina(n4856), .dinb(n4848), .dout(n4857));
  jxor g04665(.dina(n4857), .dinb(n4842), .dout(n4858));
  jand g04666(.dina(\a[31] ), .dinb(\a[19] ), .dout(n4859));
  jnot g04667(.din(n4859), .dout(n4860));
  jand g04668(.dina(\a[30] ), .dinb(\a[20] ), .dout(n4861));
  jor  g04669(.dina(n4861), .dinb(n4672), .dout(n4862));
  jand g04670(.dina(\a[30] ), .dinb(\a[21] ), .dout(n4863));
  jand g04671(.dina(n4863), .dinb(n4668), .dout(n4864));
  jnot g04672(.din(n4864), .dout(n4865));
  jand g04673(.dina(n4865), .dinb(n4862), .dout(n4866));
  jxor g04674(.dina(n4866), .dinb(n4860), .dout(n4867));
  jnot g04675(.din(n4678), .dout(n4868));
  jand g04676(.dina(\a[46] ), .dinb(\a[4] ), .dout(n4869));
  jand g04677(.dina(\a[33] ), .dinb(\a[17] ), .dout(n4870));
  jor  g04678(.dina(n4870), .dinb(n4869), .dout(n4871));
  jand g04679(.dina(\a[46] ), .dinb(\a[17] ), .dout(n4872));
  jand g04680(.dina(n4872), .dinb(n2797), .dout(n4873));
  jnot g04681(.din(n4873), .dout(n4874));
  jand g04682(.dina(n4874), .dinb(n4871), .dout(n4875));
  jxor g04683(.dina(n4875), .dinb(n4868), .dout(n4876));
  jnot g04684(.din(n4876), .dout(n4877));
  jand g04685(.dina(\a[50] ), .dinb(\a[0] ), .dout(n4878));
  jand g04686(.dina(\a[48] ), .dinb(\a[2] ), .dout(n4879));
  jor  g04687(.dina(n4879), .dinb(n4878), .dout(n4880));
  jand g04688(.dina(\a[50] ), .dinb(\a[2] ), .dout(n4881));
  jand g04689(.dina(n4881), .dinb(n4596), .dout(n4882));
  jnot g04690(.din(n4882), .dout(n4883));
  jand g04691(.dina(n4883), .dinb(n4880), .dout(n4884));
  jxor g04692(.dina(n4884), .dinb(n4769), .dout(n4885));
  jxor g04693(.dina(n4885), .dinb(n4877), .dout(n4886));
  jxor g04694(.dina(n4886), .dinb(n4867), .dout(n4887));
  jand g04695(.dina(\a[38] ), .dinb(\a[12] ), .dout(n4888));
  jnot g04696(.din(n4888), .dout(n4889));
  jand g04697(.dina(\a[40] ), .dinb(\a[10] ), .dout(n4890));
  jor  g04698(.dina(n4890), .dinb(n3973), .dout(n4891));
  jand g04699(.dina(\a[40] ), .dinb(\a[11] ), .dout(n4892));
  jand g04700(.dina(n4892), .dinb(n4661), .dout(n4893));
  jnot g04701(.din(n4893), .dout(n4894));
  jand g04702(.dina(n4894), .dinb(n4891), .dout(n4895));
  jxor g04703(.dina(n4895), .dinb(n4889), .dout(n4896));
  jnot g04704(.din(n4706), .dout(n4897));
  jand g04705(.dina(\a[37] ), .dinb(\a[13] ), .dout(n4898));
  jand g04706(.dina(\a[41] ), .dinb(\a[9] ), .dout(n4899));
  jor  g04707(.dina(n4899), .dinb(n4898), .dout(n4900));
  jand g04708(.dina(\a[41] ), .dinb(\a[13] ), .dout(n4901));
  jand g04709(.dina(n4901), .dinb(n4009), .dout(n4902));
  jnot g04710(.din(n4902), .dout(n4903));
  jand g04711(.dina(n4903), .dinb(n4900), .dout(n4904));
  jxor g04712(.dina(n4904), .dinb(n4897), .dout(n4905));
  jand g04713(.dina(\a[44] ), .dinb(\a[6] ), .dout(n4906));
  jnot g04714(.din(n4906), .dout(n4907));
  jand g04715(.dina(\a[43] ), .dinb(\a[7] ), .dout(n4908));
  jand g04716(.dina(\a[36] ), .dinb(\a[14] ), .dout(n4909));
  jxor g04717(.dina(n4909), .dinb(n4908), .dout(n4910));
  jxor g04718(.dina(n4910), .dinb(n4907), .dout(n4911));
  jnot g04719(.din(n4911), .dout(n4912));
  jxor g04720(.dina(n4912), .dinb(n4905), .dout(n4913));
  jxor g04721(.dina(n4913), .dinb(n4896), .dout(n4914));
  jxor g04722(.dina(n4914), .dinb(n4887), .dout(n4915));
  jxor g04723(.dina(n4915), .dinb(n4858), .dout(n4916));
  jxor g04724(.dina(n4916), .dinb(n4840), .dout(n4917));
  jxor g04725(.dina(n4917), .dinb(n4835), .dout(n4918));
  jxor g04726(.dina(n4918), .dinb(n4832), .dout(n4919));
  jand g04727(.dina(n4713), .dinb(n4630), .dout(n4920));
  jand g04728(.dina(n4714), .dinb(n4625), .dout(n4921));
  jor  g04729(.dina(n4921), .dinb(n4920), .dout(n4922));
  jand g04730(.dina(n4736), .dinb(n4730), .dout(n4923));
  jnot g04731(.din(n4923), .dout(n4924));
  jor  g04732(.dina(n4742), .dinb(n4738), .dout(n4925));
  jand g04733(.dina(n4925), .dinb(n4924), .dout(n4926));
  jnot g04734(.din(n4926), .dout(n4927));
  jand g04735(.dina(n4780), .dinb(n4766), .dout(n4928));
  jand g04736(.dina(n4781), .dinb(n4761), .dout(n4929));
  jor  g04737(.dina(n4929), .dinb(n4928), .dout(n4930));
  jxor g04738(.dina(n4930), .dinb(n4927), .dout(n4931));
  jand g04739(.dina(n4726), .dinb(n4718), .dout(n4932));
  jand g04740(.dina(n4729), .dinb(n4727), .dout(n4933));
  jor  g04741(.dina(n4933), .dinb(n4932), .dout(n4934));
  jnot g04742(.din(n4934), .dout(n4935));
  jor  g04743(.dina(n4757), .dinb(n4750), .dout(n4936));
  jand g04744(.dina(n4760), .dinb(n4758), .dout(n4937));
  jnot g04745(.din(n4937), .dout(n4938));
  jand g04746(.dina(n4938), .dinb(n4936), .dout(n4939));
  jxor g04747(.dina(n4939), .dinb(n4935), .dout(n4940));
  jand g04748(.dina(n4681), .dinb(n4508), .dout(n4941));
  jor  g04749(.dina(n4941), .dinb(n4679), .dout(n4942));
  jand g04750(.dina(n4645), .dinb(n4641), .dout(n4943));
  jor  g04751(.dina(n4943), .dinb(n4647), .dout(n4944));
  jxor g04752(.dina(n4944), .dinb(n4942), .dout(n4945));
  jand g04753(.dina(n4689), .dinb(n4686), .dout(n4946));
  jor  g04754(.dina(n4946), .dinb(n4692), .dout(n4947));
  jxor g04755(.dina(n4947), .dinb(n4945), .dout(n4948));
  jxor g04756(.dina(n4948), .dinb(n4940), .dout(n4949));
  jxor g04757(.dina(n4949), .dinb(n4931), .dout(n4950));
  jxor g04758(.dina(n4950), .dinb(n4922), .dout(n4951));
  jnot g04759(.din(n4650), .dout(n4952));
  jnot g04760(.din(n4656), .dout(n4953));
  jand g04761(.dina(n4953), .dinb(n4952), .dout(n4954));
  jand g04762(.dina(n4657), .dinb(n4640), .dout(n4955));
  jor  g04763(.dina(n4955), .dinb(n4954), .dout(n4956));
  jnot g04764(.din(n4675), .dout(n4957));
  jor  g04765(.dina(n4682), .dinb(n4957), .dout(n4958));
  jnot g04766(.din(n4667), .dout(n4959));
  jand g04767(.dina(n4682), .dinb(n4957), .dout(n4960));
  jor  g04768(.dina(n4960), .dinb(n4959), .dout(n4961));
  jand g04769(.dina(n4961), .dinb(n4958), .dout(n4962));
  jxor g04770(.dina(n4962), .dinb(n4956), .dout(n4963));
  jand g04771(.dina(\a[26] ), .dinb(\a[24] ), .dout(n4964));
  jand g04772(.dina(\a[49] ), .dinb(\a[1] ), .dout(n4965));
  jxor g04773(.dina(n4965), .dinb(n4964), .dout(n4966));
  jnot g04774(.din(n4698), .dout(n4967));
  jand g04775(.dina(n4967), .dinb(n4697), .dout(n4968));
  jnot g04776(.din(n4968), .dout(n4969));
  jand g04777(.dina(n4698), .dinb(n4696), .dout(n4970));
  jor  g04778(.dina(n4970), .dinb(n4403), .dout(n4971));
  jand g04779(.dina(n4971), .dinb(n4969), .dout(n4972));
  jxor g04780(.dina(n4972), .dinb(n4966), .dout(n4973));
  jand g04781(.dina(n4662), .dinb(n4659), .dout(n4974));
  jor  g04782(.dina(n4974), .dinb(n4665), .dout(n4975));
  jxor g04783(.dina(n4975), .dinb(n4973), .dout(n4976));
  jxor g04784(.dina(n4976), .dinb(n4963), .dout(n4977));
  jand g04785(.dina(n4709), .dinb(n4702), .dout(n4978));
  jor  g04786(.dina(n4978), .dinb(n4707), .dout(n4979));
  jand g04787(.dina(n4670), .dinb(n4500), .dout(n4980));
  jor  g04788(.dina(n4980), .dinb(n4673), .dout(n4981));
  jand g04789(.dina(n4634), .dinb(n4631), .dout(n4982));
  jor  g04790(.dina(n4982), .dinb(n4637), .dout(n4983));
  jxor g04791(.dina(n4983), .dinb(n4981), .dout(n4984));
  jxor g04792(.dina(n4984), .dinb(n4979), .dout(n4985));
  jor  g04793(.dina(n4710), .dinb(n4701), .dout(n4986));
  jand g04794(.dina(n4710), .dinb(n4701), .dout(n4987));
  jor  g04795(.dina(n4987), .dinb(n4695), .dout(n4988));
  jand g04796(.dina(n4988), .dinb(n4986), .dout(n4989));
  jxor g04797(.dina(n4989), .dinb(n4985), .dout(n4990));
  jand g04798(.dina(n4796), .dinb(n4789), .dout(n4991));
  jand g04799(.dina(n4800), .dinb(n4797), .dout(n4992));
  jor  g04800(.dina(n4992), .dinb(n4991), .dout(n4993));
  jxor g04801(.dina(n4993), .dinb(n4990), .dout(n4994));
  jand g04802(.dina(n4684), .dinb(n4658), .dout(n4995));
  jand g04803(.dina(n4712), .dinb(n4685), .dout(n4996));
  jor  g04804(.dina(n4996), .dinb(n4995), .dout(n4997));
  jxor g04805(.dina(n4997), .dinb(n4994), .dout(n4998));
  jxor g04806(.dina(n4998), .dinb(n4977), .dout(n4999));
  jxor g04807(.dina(n4999), .dinb(n4951), .dout(n5000));
  jxor g04808(.dina(n5000), .dinb(n4919), .dout(n5001));
  jxor g04809(.dina(n5001), .dinb(n4829), .dout(n5002));
  jand g04810(.dina(n4817), .dinb(n4814), .dout(n5003));
  jnot g04811(.din(n4814), .dout(n5004));
  jnot g04812(.din(n4817), .dout(n5005));
  jand g04813(.dina(n5005), .dinb(n5004), .dout(n5006));
  jnot g04814(.din(n5006), .dout(n5007));
  jand g04815(.dina(n4825), .dinb(n5007), .dout(n5008));
  jor  g04816(.dina(n5008), .dinb(n5003), .dout(n5009));
  jxor g04817(.dina(n5009), .dinb(n5002), .dout(\asquared[51] ));
  jand g04818(.dina(n4918), .dinb(n4832), .dout(n5011));
  jand g04819(.dina(n5000), .dinb(n4919), .dout(n5012));
  jor  g04820(.dina(n5012), .dinb(n5011), .dout(n5013));
  jand g04821(.dina(n4950), .dinb(n4922), .dout(n5014));
  jand g04822(.dina(n4999), .dinb(n4951), .dout(n5015));
  jor  g04823(.dina(n5015), .dinb(n5014), .dout(n5016));
  jand g04824(.dina(n4997), .dinb(n4994), .dout(n5017));
  jand g04825(.dina(n4998), .dinb(n4977), .dout(n5018));
  jor  g04826(.dina(n5018), .dinb(n5017), .dout(n5019));
  jand g04827(.dina(n4930), .dinb(n4927), .dout(n5020));
  jand g04828(.dina(n4949), .dinb(n4931), .dout(n5021));
  jor  g04829(.dina(n5021), .dinb(n5020), .dout(n5022));
  jand g04830(.dina(n4983), .dinb(n4981), .dout(n5023));
  jand g04831(.dina(n4984), .dinb(n4979), .dout(n5024));
  jor  g04832(.dina(n5024), .dinb(n5023), .dout(n5025));
  jand g04833(.dina(n4965), .dinb(n4964), .dout(n5026));
  jand g04834(.dina(\a[51] ), .dinb(\a[0] ), .dout(n5027));
  jxor g04835(.dina(n5027), .dinb(n5026), .dout(n5028));
  jand g04836(.dina(\a[50] ), .dinb(\a[1] ), .dout(n5029));
  jxor g04837(.dina(n5029), .dinb(\a[26] ), .dout(n5030));
  jnot g04838(.din(n5030), .dout(n5031));
  jxor g04839(.dina(n5031), .dinb(n5028), .dout(n5032));
  jand g04840(.dina(\a[34] ), .dinb(\a[17] ), .dout(n5033));
  jand g04841(.dina(\a[31] ), .dinb(\a[20] ), .dout(n5034));
  jand g04842(.dina(\a[32] ), .dinb(\a[19] ), .dout(n5035));
  jor  g04843(.dina(n5035), .dinb(n5034), .dout(n5036));
  jnot g04844(.din(n5036), .dout(n5037));
  jand g04845(.dina(\a[32] ), .dinb(\a[20] ), .dout(n5038));
  jand g04846(.dina(n5038), .dinb(n4859), .dout(n5039));
  jor  g04847(.dina(n5039), .dinb(n5037), .dout(n5040));
  jxor g04848(.dina(n5040), .dinb(n5033), .dout(n5041));
  jxor g04849(.dina(n5041), .dinb(n5032), .dout(n5042));
  jxor g04850(.dina(n5042), .dinb(n5025), .dout(n5043));
  jand g04851(.dina(\a[26] ), .dinb(\a[25] ), .dout(n5044));
  jand g04852(.dina(\a[27] ), .dinb(\a[24] ), .dout(n5045));
  jor  g04853(.dina(n5045), .dinb(n5044), .dout(n5046));
  jnot g04854(.din(n5046), .dout(n5047));
  jand g04855(.dina(\a[27] ), .dinb(\a[25] ), .dout(n5048));
  jand g04856(.dina(n5048), .dinb(n4964), .dout(n5049));
  jor  g04857(.dina(n5049), .dinb(n5047), .dout(n5050));
  jxor g04858(.dina(n5050), .dinb(n4892), .dout(n5051));
  jnot g04859(.din(n5051), .dout(n5052));
  jand g04860(.dina(\a[44] ), .dinb(\a[7] ), .dout(n5053));
  jand g04861(.dina(\a[38] ), .dinb(\a[13] ), .dout(n5054));
  jand g04862(.dina(\a[43] ), .dinb(\a[8] ), .dout(n5055));
  jor  g04863(.dina(n5055), .dinb(n5054), .dout(n5056));
  jand g04864(.dina(\a[43] ), .dinb(\a[13] ), .dout(n5057));
  jand g04865(.dina(n5057), .dinb(n4159), .dout(n5058));
  jnot g04866(.din(n5058), .dout(n5059));
  jand g04867(.dina(n5059), .dinb(n5056), .dout(n5060));
  jxor g04868(.dina(n5060), .dinb(n5053), .dout(n5061));
  jnot g04869(.din(n5061), .dout(n5062));
  jand g04870(.dina(\a[42] ), .dinb(\a[9] ), .dout(n5063));
  jand g04871(.dina(\a[41] ), .dinb(\a[10] ), .dout(n5064));
  jor  g04872(.dina(n5064), .dinb(n4664), .dout(n5065));
  jnot g04873(.din(n5065), .dout(n5066));
  jand g04874(.dina(\a[41] ), .dinb(\a[12] ), .dout(n5067));
  jand g04875(.dina(n5067), .dinb(n4661), .dout(n5068));
  jor  g04876(.dina(n5068), .dinb(n5066), .dout(n5069));
  jxor g04877(.dina(n5069), .dinb(n5063), .dout(n5070));
  jxor g04878(.dina(n5070), .dinb(n5062), .dout(n5071));
  jxor g04879(.dina(n5071), .dinb(n5052), .dout(n5072));
  jand g04880(.dina(\a[36] ), .dinb(\a[15] ), .dout(n5073));
  jnot g04881(.din(n5073), .dout(n5074));
  jand g04882(.dina(\a[45] ), .dinb(\a[6] ), .dout(n5075));
  jand g04883(.dina(\a[37] ), .dinb(\a[14] ), .dout(n5076));
  jor  g04884(.dina(n5076), .dinb(n5075), .dout(n5077));
  jand g04885(.dina(\a[45] ), .dinb(\a[14] ), .dout(n5078));
  jand g04886(.dina(n5078), .dinb(n3707), .dout(n5079));
  jnot g04887(.din(n5079), .dout(n5080));
  jand g04888(.dina(n5080), .dinb(n5077), .dout(n5081));
  jxor g04889(.dina(n5081), .dinb(n5074), .dout(n5082));
  jnot g04890(.din(n4863), .dout(n5083));
  jand g04891(.dina(\a[29] ), .dinb(\a[22] ), .dout(n5084));
  jand g04892(.dina(\a[28] ), .dinb(\a[23] ), .dout(n5085));
  jor  g04893(.dina(n5085), .dinb(n5084), .dout(n5086));
  jand g04894(.dina(\a[29] ), .dinb(\a[23] ), .dout(n5087));
  jand g04895(.dina(n5087), .dinb(n4843), .dout(n5088));
  jnot g04896(.din(n5088), .dout(n5089));
  jand g04897(.dina(n5089), .dinb(n5086), .dout(n5090));
  jxor g04898(.dina(n5090), .dinb(n5083), .dout(n5091));
  jand g04899(.dina(\a[33] ), .dinb(\a[18] ), .dout(n5092));
  jnot g04900(.din(n5092), .dout(n5093));
  jand g04901(.dina(\a[46] ), .dinb(\a[5] ), .dout(n5094));
  jand g04902(.dina(\a[35] ), .dinb(\a[16] ), .dout(n5095));
  jxor g04903(.dina(n5095), .dinb(n5094), .dout(n5096));
  jxor g04904(.dina(n5096), .dinb(n5093), .dout(n5097));
  jnot g04905(.din(n5097), .dout(n5098));
  jxor g04906(.dina(n5098), .dinb(n5091), .dout(n5099));
  jxor g04907(.dina(n5099), .dinb(n5082), .dout(n5100));
  jxor g04908(.dina(n5100), .dinb(n5072), .dout(n5101));
  jxor g04909(.dina(n5101), .dinb(n5043), .dout(n5102));
  jxor g04910(.dina(n5102), .dinb(n5022), .dout(n5103));
  jxor g04911(.dina(n5103), .dinb(n5019), .dout(n5104));
  jxor g04912(.dina(n5104), .dinb(n5016), .dout(n5105));
  jand g04913(.dina(n4916), .dinb(n4840), .dout(n5106));
  jand g04914(.dina(n4917), .dinb(n4835), .dout(n5107));
  jor  g04915(.dina(n5107), .dinb(n5106), .dout(n5108));
  jand g04916(.dina(n4989), .dinb(n4985), .dout(n5109));
  jand g04917(.dina(n4993), .dinb(n4990), .dout(n5110));
  jor  g04918(.dina(n5110), .dinb(n5109), .dout(n5111));
  jand g04919(.dina(n4962), .dinb(n4956), .dout(n5112));
  jand g04920(.dina(n4976), .dinb(n4963), .dout(n5113));
  jor  g04921(.dina(n5113), .dinb(n5112), .dout(n5114));
  jxor g04922(.dina(n5114), .dinb(n5111), .dout(n5115));
  jand g04923(.dina(n4944), .dinb(n4942), .dout(n5116));
  jand g04924(.dina(n4947), .dinb(n4945), .dout(n5117));
  jor  g04925(.dina(n5117), .dinb(n5116), .dout(n5118));
  jand g04926(.dina(n4972), .dinb(n4966), .dout(n5119));
  jand g04927(.dina(n4975), .dinb(n4973), .dout(n5120));
  jor  g04928(.dina(n5120), .dinb(n5119), .dout(n5121));
  jxor g04929(.dina(n5121), .dinb(n5118), .dout(n5122));
  jnot g04930(.din(n5122), .dout(n5123));
  jnot g04931(.din(n4885), .dout(n5124));
  jand g04932(.dina(n5124), .dinb(n4877), .dout(n5125));
  jnot g04933(.din(n5125), .dout(n5126));
  jand g04934(.dina(n4885), .dinb(n4876), .dout(n5127));
  jor  g04935(.dina(n5127), .dinb(n4867), .dout(n5128));
  jand g04936(.dina(n5128), .dinb(n5126), .dout(n5129));
  jxor g04937(.dina(n5129), .dinb(n5123), .dout(n5130));
  jxor g04938(.dina(n5130), .dinb(n5115), .dout(n5131));
  jxor g04939(.dina(n5131), .dinb(n5108), .dout(n5132));
  jand g04940(.dina(n4914), .dinb(n4887), .dout(n5133));
  jand g04941(.dina(n4915), .dinb(n4858), .dout(n5134));
  jor  g04942(.dina(n5134), .dinb(n5133), .dout(n5135));
  jand g04943(.dina(n4856), .dinb(n4848), .dout(n5136));
  jand g04944(.dina(n4857), .dinb(n4842), .dout(n5137));
  jor  g04945(.dina(n5137), .dinb(n5136), .dout(n5138));
  jand g04946(.dina(n4855), .dinb(n4849), .dout(n5139));
  jor  g04947(.dina(n5139), .dinb(n4853), .dout(n5140));
  jand g04948(.dina(n4891), .dinb(n4888), .dout(n5141));
  jor  g04949(.dina(n5141), .dinb(n4893), .dout(n5142));
  jxor g04950(.dina(n5142), .dinb(n5140), .dout(n5143));
  jand g04951(.dina(\a[49] ), .dinb(\a[2] ), .dout(n5144));
  jand g04952(.dina(\a[48] ), .dinb(\a[3] ), .dout(n5145));
  jand g04953(.dina(\a[47] ), .dinb(\a[4] ), .dout(n5146));
  jor  g04954(.dina(n5146), .dinb(n5145), .dout(n5147));
  jnot g04955(.din(n5147), .dout(n5148));
  jand g04956(.dina(\a[48] ), .dinb(\a[4] ), .dout(n5149));
  jand g04957(.dina(n5149), .dinb(n4678), .dout(n5150));
  jor  g04958(.dina(n5150), .dinb(n5148), .dout(n5151));
  jxor g04959(.dina(n5151), .dinb(n5144), .dout(n5152));
  jnot g04960(.din(n5152), .dout(n5153));
  jxor g04961(.dina(n5153), .dinb(n5143), .dout(n5154));
  jxor g04962(.dina(n5154), .dinb(n5138), .dout(n5155));
  jnot g04963(.din(n5155), .dout(n5156));
  jor  g04964(.dina(n4939), .dinb(n4935), .dout(n5157));
  jand g04965(.dina(n4948), .dinb(n4940), .dout(n5158));
  jnot g04966(.din(n5158), .dout(n5159));
  jand g04967(.dina(n5159), .dinb(n5157), .dout(n5160));
  jxor g04968(.dina(n5160), .dinb(n5156), .dout(n5161));
  jxor g04969(.dina(n5161), .dinb(n5135), .dout(n5162));
  jand g04970(.dina(n4900), .dinb(n4706), .dout(n5163));
  jor  g04971(.dina(n5163), .dinb(n4902), .dout(n5164));
  jand g04972(.dina(n4909), .dinb(n4908), .dout(n5165));
  jnot g04973(.din(n5165), .dout(n5166));
  jnot g04974(.din(n4908), .dout(n5167));
  jnot g04975(.din(n4909), .dout(n5168));
  jand g04976(.dina(n5168), .dinb(n5167), .dout(n5169));
  jor  g04977(.dina(n5169), .dinb(n4907), .dout(n5170));
  jand g04978(.dina(n5170), .dinb(n5166), .dout(n5171));
  jnot g04979(.din(n5171), .dout(n5172));
  jxor g04980(.dina(n5172), .dinb(n5164), .dout(n5173));
  jand g04981(.dina(n4845), .dinb(n4636), .dout(n5174));
  jnot g04982(.din(n5174), .dout(n5175));
  jnot g04983(.din(n4636), .dout(n5176));
  jnot g04984(.din(n4845), .dout(n5177));
  jand g04985(.dina(n5177), .dinb(n5176), .dout(n5178));
  jor  g04986(.dina(n5178), .dinb(n4844), .dout(n5179));
  jand g04987(.dina(n5179), .dinb(n5175), .dout(n5180));
  jnot g04988(.din(n5180), .dout(n5181));
  jxor g04989(.dina(n5181), .dinb(n5173), .dout(n5182));
  jnot g04990(.din(n5182), .dout(n5183));
  jnot g04991(.din(n4905), .dout(n5184));
  jand g04992(.dina(n4912), .dinb(n5184), .dout(n5185));
  jnot g04993(.din(n5185), .dout(n5186));
  jand g04994(.dina(n4911), .dinb(n4905), .dout(n5187));
  jor  g04995(.dina(n5187), .dinb(n4896), .dout(n5188));
  jand g04996(.dina(n5188), .dinb(n5186), .dout(n5189));
  jxor g04997(.dina(n5189), .dinb(n5183), .dout(n5190));
  jand g04998(.dina(n4871), .dinb(n4678), .dout(n5191));
  jor  g04999(.dina(n5191), .dinb(n4873), .dout(n5192));
  jand g05000(.dina(n4862), .dinb(n4859), .dout(n5193));
  jor  g05001(.dina(n5193), .dinb(n4864), .dout(n5194));
  jxor g05002(.dina(n5194), .dinb(n5192), .dout(n5195));
  jand g05003(.dina(n4880), .dinb(n4768), .dout(n5196));
  jor  g05004(.dina(n5196), .dinb(n4882), .dout(n5197));
  jxor g05005(.dina(n5197), .dinb(n5195), .dout(n5198));
  jxor g05006(.dina(n5198), .dinb(n5190), .dout(n5199));
  jxor g05007(.dina(n5199), .dinb(n5162), .dout(n5200));
  jxor g05008(.dina(n5200), .dinb(n5132), .dout(n5201));
  jxor g05009(.dina(n5201), .dinb(n5105), .dout(n5202));
  jxor g05010(.dina(n5202), .dinb(n5013), .dout(n5203));
  jand g05011(.dina(n5001), .dinb(n4829), .dout(n5204));
  jnot g05012(.din(n4829), .dout(n5205));
  jnot g05013(.din(n5001), .dout(n5206));
  jand g05014(.dina(n5206), .dinb(n5205), .dout(n5207));
  jnot g05015(.din(n5207), .dout(n5208));
  jand g05016(.dina(n5009), .dinb(n5208), .dout(n5209));
  jor  g05017(.dina(n5209), .dinb(n5204), .dout(n5210));
  jxor g05018(.dina(n5210), .dinb(n5203), .dout(\asquared[52] ));
  jand g05019(.dina(n5104), .dinb(n5016), .dout(n5212));
  jand g05020(.dina(n5201), .dinb(n5105), .dout(n5213));
  jor  g05021(.dina(n5213), .dinb(n5212), .dout(n5214));
  jand g05022(.dina(n5161), .dinb(n5135), .dout(n5215));
  jand g05023(.dina(n5199), .dinb(n5162), .dout(n5216));
  jor  g05024(.dina(n5216), .dinb(n5215), .dout(n5217));
  jand g05025(.dina(n5114), .dinb(n5111), .dout(n5218));
  jand g05026(.dina(n5130), .dinb(n5115), .dout(n5219));
  jor  g05027(.dina(n5219), .dinb(n5218), .dout(n5220));
  jor  g05028(.dina(n5189), .dinb(n5183), .dout(n5221));
  jand g05029(.dina(n5198), .dinb(n5190), .dout(n5222));
  jnot g05030(.din(n5222), .dout(n5223));
  jand g05031(.dina(n5223), .dinb(n5221), .dout(n5224));
  jnot g05032(.din(n5224), .dout(n5225));
  jand g05033(.dina(\a[30] ), .dinb(\a[22] ), .dout(n5226));
  jand g05034(.dina(\a[28] ), .dinb(\a[24] ), .dout(n5227));
  jor  g05035(.dina(n5227), .dinb(n5087), .dout(n5228));
  jnot g05036(.din(n5228), .dout(n5229));
  jand g05037(.dina(\a[29] ), .dinb(\a[24] ), .dout(n5230));
  jand g05038(.dina(n5230), .dinb(n5085), .dout(n5231));
  jor  g05039(.dina(n5231), .dinb(n5229), .dout(n5232));
  jxor g05040(.dina(n5232), .dinb(n5226), .dout(n5233));
  jnot g05041(.din(n5233), .dout(n5234));
  jand g05042(.dina(\a[34] ), .dinb(\a[18] ), .dout(n5235));
  jand g05043(.dina(\a[31] ), .dinb(\a[21] ), .dout(n5236));
  jor  g05044(.dina(n5236), .dinb(n5038), .dout(n5237));
  jand g05045(.dina(\a[32] ), .dinb(\a[21] ), .dout(n5238));
  jand g05046(.dina(n5238), .dinb(n5034), .dout(n5239));
  jnot g05047(.din(n5239), .dout(n5240));
  jand g05048(.dina(n5240), .dinb(n5237), .dout(n5241));
  jxor g05049(.dina(n5241), .dinb(n5235), .dout(n5242));
  jxor g05050(.dina(n5242), .dinb(n5234), .dout(n5243));
  jnot g05051(.din(n5243), .dout(n5244));
  jand g05052(.dina(\a[39] ), .dinb(\a[13] ), .dout(n5245));
  jand g05053(.dina(\a[43] ), .dinb(\a[9] ), .dout(n5246));
  jor  g05054(.dina(n5246), .dinb(n5245), .dout(n5247));
  jnot g05055(.din(n5247), .dout(n5248));
  jand g05056(.dina(n5057), .dinb(n4471), .dout(n5249));
  jor  g05057(.dina(n5249), .dinb(n5248), .dout(n5250));
  jxor g05058(.dina(n5250), .dinb(n3553), .dout(n5251));
  jxor g05059(.dina(n5251), .dinb(n5244), .dout(n5252));
  jand g05060(.dina(\a[37] ), .dinb(\a[15] ), .dout(n5253));
  jand g05061(.dina(\a[45] ), .dinb(\a[7] ), .dout(n5254));
  jand g05062(.dina(\a[44] ), .dinb(\a[8] ), .dout(n5255));
  jor  g05063(.dina(n5255), .dinb(n5254), .dout(n5256));
  jnot g05064(.din(n5256), .dout(n5257));
  jand g05065(.dina(\a[45] ), .dinb(\a[8] ), .dout(n5258));
  jand g05066(.dina(n5258), .dinb(n5053), .dout(n5259));
  jor  g05067(.dina(n5259), .dinb(n5257), .dout(n5260));
  jxor g05068(.dina(n5260), .dinb(n5253), .dout(n5261));
  jand g05069(.dina(\a[42] ), .dinb(\a[10] ), .dout(n5262));
  jand g05070(.dina(\a[41] ), .dinb(\a[11] ), .dout(n5263));
  jor  g05071(.dina(n5263), .dinb(n4325), .dout(n5264));
  jnot g05072(.din(n5264), .dout(n5265));
  jand g05073(.dina(n5067), .dinb(n4892), .dout(n5266));
  jor  g05074(.dina(n5266), .dinb(n5265), .dout(n5267));
  jxor g05075(.dina(n5267), .dinb(n5262), .dout(n5268));
  jand g05076(.dina(\a[47] ), .dinb(\a[5] ), .dout(n5269));
  jand g05077(.dina(\a[36] ), .dinb(\a[16] ), .dout(n5270));
  jand g05078(.dina(\a[46] ), .dinb(\a[6] ), .dout(n5271));
  jor  g05079(.dina(n5271), .dinb(n5270), .dout(n5272));
  jand g05080(.dina(\a[46] ), .dinb(\a[16] ), .dout(n5273));
  jand g05081(.dina(n5273), .dinb(n3536), .dout(n5274));
  jnot g05082(.din(n5274), .dout(n5275));
  jand g05083(.dina(n5275), .dinb(n5272), .dout(n5276));
  jxor g05084(.dina(n5276), .dinb(n5269), .dout(n5277));
  jxor g05085(.dina(n5277), .dinb(n5268), .dout(n5278));
  jxor g05086(.dina(n5278), .dinb(n5261), .dout(n5279));
  jxor g05087(.dina(n5279), .dinb(n5252), .dout(n5280));
  jxor g05088(.dina(n5280), .dinb(n5225), .dout(n5281));
  jxor g05089(.dina(n5281), .dinb(n5220), .dout(n5282));
  jxor g05090(.dina(n5282), .dinb(n5217), .dout(n5283));
  jand g05091(.dina(n5131), .dinb(n5108), .dout(n5284));
  jand g05092(.dina(n5200), .dinb(n5132), .dout(n5285));
  jor  g05093(.dina(n5285), .dinb(n5284), .dout(n5286));
  jxor g05094(.dina(n5286), .dinb(n5283), .dout(n5287));
  jand g05095(.dina(n5102), .dinb(n5022), .dout(n5288));
  jand g05096(.dina(n5103), .dinb(n5019), .dout(n5289));
  jor  g05097(.dina(n5289), .dinb(n5288), .dout(n5290));
  jand g05098(.dina(n5172), .dinb(n5164), .dout(n5291));
  jand g05099(.dina(n5181), .dinb(n5173), .dout(n5292));
  jor  g05100(.dina(n5292), .dinb(n5291), .dout(n5293));
  jand g05101(.dina(n5194), .dinb(n5192), .dout(n5294));
  jand g05102(.dina(n5197), .dinb(n5195), .dout(n5295));
  jor  g05103(.dina(n5295), .dinb(n5294), .dout(n5296));
  jand g05104(.dina(\a[33] ), .dinb(\a[19] ), .dout(n5297));
  jand g05105(.dina(\a[49] ), .dinb(\a[3] ), .dout(n5298));
  jor  g05106(.dina(n5298), .dinb(n4881), .dout(n5299));
  jnot g05107(.din(n5299), .dout(n5300));
  jand g05108(.dina(\a[50] ), .dinb(\a[3] ), .dout(n5301));
  jand g05109(.dina(n5301), .dinb(n5144), .dout(n5302));
  jor  g05110(.dina(n5302), .dinb(n5300), .dout(n5303));
  jxor g05111(.dina(n5303), .dinb(n5297), .dout(n5304));
  jnot g05112(.din(n5304), .dout(n5305));
  jxor g05113(.dina(n5305), .dinb(n5296), .dout(n5306));
  jxor g05114(.dina(n5306), .dinb(n5293), .dout(n5307));
  jnot g05115(.din(n5307), .dout(n5308));
  jand g05116(.dina(n5154), .dinb(n5138), .dout(n5309));
  jnot g05117(.din(n5309), .dout(n5310));
  jor  g05118(.dina(n5160), .dinb(n5156), .dout(n5311));
  jand g05119(.dina(n5311), .dinb(n5310), .dout(n5312));
  jxor g05120(.dina(n5312), .dinb(n5308), .dout(n5313));
  jor  g05121(.dina(n5070), .dinb(n5062), .dout(n5314));
  jand g05122(.dina(n5071), .dinb(n5052), .dout(n5315));
  jnot g05123(.din(n5315), .dout(n5316));
  jand g05124(.dina(n5316), .dinb(n5314), .dout(n5317));
  jnot g05125(.din(n5317), .dout(n5318));
  jand g05126(.dina(n5029), .dinb(\a[26] ), .dout(n5319));
  jand g05127(.dina(\a[51] ), .dinb(\a[1] ), .dout(n5320));
  jxor g05128(.dina(n5320), .dinb(n5048), .dout(n5321));
  jxor g05129(.dina(n5321), .dinb(n5319), .dout(n5322));
  jand g05130(.dina(n5046), .dinb(n4892), .dout(n5323));
  jor  g05131(.dina(n5323), .dinb(n5049), .dout(n5324));
  jxor g05132(.dina(n5324), .dinb(n5322), .dout(n5325));
  jnot g05133(.din(n5140), .dout(n5326));
  jnot g05134(.din(n5142), .dout(n5327));
  jand g05135(.dina(n5327), .dinb(n5326), .dout(n5328));
  jnot g05136(.din(n5328), .dout(n5329));
  jand g05137(.dina(n5142), .dinb(n5140), .dout(n5330));
  jor  g05138(.dina(n5153), .dinb(n5330), .dout(n5331));
  jand g05139(.dina(n5331), .dinb(n5329), .dout(n5332));
  jxor g05140(.dina(n5332), .dinb(n5325), .dout(n5333));
  jxor g05141(.dina(n5333), .dinb(n5318), .dout(n5334));
  jxor g05142(.dina(n5334), .dinb(n5313), .dout(n5335));
  jxor g05143(.dina(n5335), .dinb(n5290), .dout(n5336));
  jor  g05144(.dina(n5041), .dinb(n5032), .dout(n5337));
  jand g05145(.dina(n5042), .dinb(n5025), .dout(n5338));
  jnot g05146(.din(n5338), .dout(n5339));
  jand g05147(.dina(n5339), .dinb(n5337), .dout(n5340));
  jnot g05148(.din(n5340), .dout(n5341));
  jand g05149(.dina(n5065), .dinb(n5063), .dout(n5342));
  jor  g05150(.dina(n5342), .dinb(n5068), .dout(n5343));
  jor  g05151(.dina(n5027), .dinb(n5026), .dout(n5344));
  jand g05152(.dina(n5027), .dinb(n5026), .dout(n5345));
  jor  g05153(.dina(n5030), .dinb(n5345), .dout(n5346));
  jand g05154(.dina(n5346), .dinb(n5344), .dout(n5347));
  jxor g05155(.dina(n5347), .dinb(n5343), .dout(n5348));
  jand g05156(.dina(n702), .dinb(\a[35] ), .dout(n5349));
  jand g05157(.dina(n208), .dinb(\a[48] ), .dout(n5350));
  jor  g05158(.dina(n5350), .dinb(n5349), .dout(n5351));
  jand g05159(.dina(n5351), .dinb(\a[52] ), .dout(n5352));
  jnot g05160(.din(n5352), .dout(n5353));
  jand g05161(.dina(\a[35] ), .dinb(\a[17] ), .dout(n5354));
  jxor g05162(.dina(n5354), .dinb(n5149), .dout(n5355));
  jand g05163(.dina(n5355), .dinb(n5353), .dout(n5356));
  jnot g05164(.din(n5355), .dout(n5357));
  jand g05165(.dina(\a[52] ), .dinb(\a[0] ), .dout(n5358));
  jand g05166(.dina(n5358), .dinb(n5357), .dout(n5359));
  jor  g05167(.dina(n5359), .dinb(n5356), .dout(n5360));
  jxor g05168(.dina(n5360), .dinb(n5348), .dout(n5361));
  jxor g05169(.dina(n5361), .dinb(n5341), .dout(n5362));
  jnot g05170(.din(n5362), .dout(n5363));
  jand g05171(.dina(n5121), .dinb(n5118), .dout(n5364));
  jnot g05172(.din(n5364), .dout(n5365));
  jor  g05173(.dina(n5129), .dinb(n5123), .dout(n5366));
  jand g05174(.dina(n5366), .dinb(n5365), .dout(n5367));
  jxor g05175(.dina(n5367), .dinb(n5363), .dout(n5368));
  jand g05176(.dina(n5100), .dinb(n5072), .dout(n5369));
  jand g05177(.dina(n5101), .dinb(n5043), .dout(n5370));
  jor  g05178(.dina(n5370), .dinb(n5369), .dout(n5371));
  jand g05179(.dina(n5060), .dinb(n5053), .dout(n5372));
  jor  g05180(.dina(n5372), .dinb(n5058), .dout(n5373));
  jnot g05181(.din(n5373), .dout(n5374));
  jand g05182(.dina(n5095), .dinb(n5094), .dout(n5375));
  jnot g05183(.din(n5375), .dout(n5376));
  jnot g05184(.din(n5094), .dout(n5377));
  jnot g05185(.din(n5095), .dout(n5378));
  jand g05186(.dina(n5378), .dinb(n5377), .dout(n5379));
  jor  g05187(.dina(n5379), .dinb(n5093), .dout(n5380));
  jand g05188(.dina(n5380), .dinb(n5376), .dout(n5381));
  jxor g05189(.dina(n5381), .dinb(n5374), .dout(n5382));
  jand g05190(.dina(n5086), .dinb(n4863), .dout(n5383));
  jor  g05191(.dina(n5383), .dinb(n5088), .dout(n5384));
  jxor g05192(.dina(n5384), .dinb(n5382), .dout(n5385));
  jand g05193(.dina(n5036), .dinb(n5033), .dout(n5386));
  jor  g05194(.dina(n5386), .dinb(n5039), .dout(n5387));
  jand g05195(.dina(n5147), .dinb(n5144), .dout(n5388));
  jor  g05196(.dina(n5388), .dinb(n5150), .dout(n5389));
  jxor g05197(.dina(n5389), .dinb(n5387), .dout(n5390));
  jand g05198(.dina(n5077), .dinb(n5073), .dout(n5391));
  jor  g05199(.dina(n5391), .dinb(n5079), .dout(n5392));
  jxor g05200(.dina(n5392), .dinb(n5390), .dout(n5393));
  jnot g05201(.din(n5393), .dout(n5394));
  jnot g05202(.din(n5091), .dout(n5395));
  jand g05203(.dina(n5098), .dinb(n5395), .dout(n5396));
  jnot g05204(.din(n5396), .dout(n5397));
  jand g05205(.dina(n5097), .dinb(n5091), .dout(n5398));
  jor  g05206(.dina(n5398), .dinb(n5082), .dout(n5399));
  jand g05207(.dina(n5399), .dinb(n5397), .dout(n5400));
  jxor g05208(.dina(n5400), .dinb(n5394), .dout(n5401));
  jxor g05209(.dina(n5401), .dinb(n5385), .dout(n5402));
  jxor g05210(.dina(n5402), .dinb(n5371), .dout(n5403));
  jxor g05211(.dina(n5403), .dinb(n5368), .dout(n5404));
  jxor g05212(.dina(n5404), .dinb(n5336), .dout(n5405));
  jxor g05213(.dina(n5405), .dinb(n5287), .dout(n5406));
  jxor g05214(.dina(n5406), .dinb(n5214), .dout(n5407));
  jand g05215(.dina(n5202), .dinb(n5013), .dout(n5408));
  jor  g05216(.dina(n5202), .dinb(n5013), .dout(n5409));
  jand g05217(.dina(n5210), .dinb(n5409), .dout(n5410));
  jor  g05218(.dina(n5410), .dinb(n5408), .dout(n5411));
  jxor g05219(.dina(n5411), .dinb(n5407), .dout(\asquared[53] ));
  jand g05220(.dina(n5286), .dinb(n5283), .dout(n5413));
  jand g05221(.dina(n5405), .dinb(n5287), .dout(n5414));
  jor  g05222(.dina(n5414), .dinb(n5413), .dout(n5415));
  jand g05223(.dina(n5335), .dinb(n5290), .dout(n5416));
  jand g05224(.dina(n5404), .dinb(n5336), .dout(n5417));
  jor  g05225(.dina(n5417), .dinb(n5416), .dout(n5418));
  jand g05226(.dina(n5402), .dinb(n5371), .dout(n5419));
  jand g05227(.dina(n5403), .dinb(n5368), .dout(n5420));
  jor  g05228(.dina(n5420), .dinb(n5419), .dout(n5421));
  jand g05229(.dina(n5305), .dinb(n5296), .dout(n5422));
  jand g05230(.dina(n5306), .dinb(n5293), .dout(n5423));
  jor  g05231(.dina(n5423), .dinb(n5422), .dout(n5424));
  jand g05232(.dina(\a[34] ), .dinb(\a[19] ), .dout(n5425));
  jnot g05233(.din(n5425), .dout(n5426));
  jand g05234(.dina(\a[33] ), .dinb(\a[20] ), .dout(n5427));
  jor  g05235(.dina(n5427), .dinb(n5238), .dout(n5428));
  jand g05236(.dina(\a[33] ), .dinb(\a[21] ), .dout(n5429));
  jand g05237(.dina(n5429), .dinb(n5038), .dout(n5430));
  jnot g05238(.din(n5430), .dout(n5431));
  jand g05239(.dina(n5431), .dinb(n5428), .dout(n5432));
  jxor g05240(.dina(n5432), .dinb(n5426), .dout(n5433));
  jand g05241(.dina(\a[49] ), .dinb(\a[4] ), .dout(n5434));
  jnot g05242(.din(n5434), .dout(n5435));
  jand g05243(.dina(\a[36] ), .dinb(\a[17] ), .dout(n5436));
  jand g05244(.dina(\a[35] ), .dinb(\a[18] ), .dout(n5437));
  jor  g05245(.dina(n5437), .dinb(n5436), .dout(n5438));
  jand g05246(.dina(\a[36] ), .dinb(\a[18] ), .dout(n5439));
  jand g05247(.dina(n5439), .dinb(n5354), .dout(n5440));
  jnot g05248(.din(n5440), .dout(n5441));
  jand g05249(.dina(n5441), .dinb(n5438), .dout(n5442));
  jxor g05250(.dina(n5442), .dinb(n5435), .dout(n5443));
  jnot g05251(.din(n5443), .dout(n5444));
  jand g05252(.dina(n5320), .dinb(n5048), .dout(n5445));
  jnot g05253(.din(n5445), .dout(n5446));
  jnot g05254(.din(n5301), .dout(n5447));
  jand g05255(.dina(\a[51] ), .dinb(\a[2] ), .dout(n5448));
  jnot g05256(.din(n5448), .dout(n5449));
  jand g05257(.dina(n5449), .dinb(n5447), .dout(n5450));
  jnot g05258(.din(n5450), .dout(n5451));
  jand g05259(.dina(\a[51] ), .dinb(\a[3] ), .dout(n5452));
  jand g05260(.dina(n5452), .dinb(n4881), .dout(n5453));
  jnot g05261(.din(n5453), .dout(n5454));
  jand g05262(.dina(n5454), .dinb(n5451), .dout(n5455));
  jxor g05263(.dina(n5455), .dinb(n5446), .dout(n5456));
  jxor g05264(.dina(n5456), .dinb(n5444), .dout(n5457));
  jxor g05265(.dina(n5457), .dinb(n5433), .dout(n5458));
  jxor g05266(.dina(n5458), .dinb(n5424), .dout(n5459));
  jand g05267(.dina(\a[53] ), .dinb(\a[0] ), .dout(n5460));
  jand g05268(.dina(\a[48] ), .dinb(\a[5] ), .dout(n5461));
  jand g05269(.dina(\a[37] ), .dinb(\a[16] ), .dout(n5462));
  jor  g05270(.dina(n5462), .dinb(n5461), .dout(n5463));
  jnot g05271(.din(n5463), .dout(n5464));
  jand g05272(.dina(\a[48] ), .dinb(\a[16] ), .dout(n5465));
  jand g05273(.dina(n5465), .dinb(n3473), .dout(n5466));
  jor  g05274(.dina(n5466), .dinb(n5464), .dout(n5467));
  jxor g05275(.dina(n5467), .dinb(n5460), .dout(n5468));
  jnot g05276(.din(n5468), .dout(n5469));
  jand g05277(.dina(\a[39] ), .dinb(\a[14] ), .dout(n5470));
  jand g05278(.dina(\a[44] ), .dinb(\a[9] ), .dout(n5471));
  jor  g05279(.dina(n5471), .dinb(n5470), .dout(n5472));
  jand g05280(.dina(\a[44] ), .dinb(\a[14] ), .dout(n5473));
  jand g05281(.dina(n5473), .dinb(n4471), .dout(n5474));
  jnot g05282(.din(n5474), .dout(n5475));
  jand g05283(.dina(n5475), .dinb(n5472), .dout(n5476));
  jxor g05284(.dina(n5476), .dinb(n5258), .dout(n5477));
  jnot g05285(.din(n5477), .dout(n5478));
  jand g05286(.dina(\a[47] ), .dinb(\a[6] ), .dout(n5479));
  jand g05287(.dina(\a[46] ), .dinb(\a[7] ), .dout(n5480));
  jnot g05288(.din(n5480), .dout(n5481));
  jand g05289(.dina(\a[38] ), .dinb(\a[15] ), .dout(n5482));
  jxor g05290(.dina(n5482), .dinb(n5481), .dout(n5483));
  jxor g05291(.dina(n5483), .dinb(n5479), .dout(n5484));
  jxor g05292(.dina(n5484), .dinb(n5478), .dout(n5485));
  jxor g05293(.dina(n5485), .dinb(n5469), .dout(n5486));
  jxor g05294(.dina(n5486), .dinb(n5459), .dout(n5487));
  jand g05295(.dina(n5332), .dinb(n5325), .dout(n5488));
  jand g05296(.dina(n5333), .dinb(n5318), .dout(n5489));
  jor  g05297(.dina(n5489), .dinb(n5488), .dout(n5490));
  jand g05298(.dina(\a[42] ), .dinb(\a[11] ), .dout(n5491));
  jand g05299(.dina(\a[27] ), .dinb(\a[26] ), .dout(n5492));
  jand g05300(.dina(\a[28] ), .dinb(\a[25] ), .dout(n5493));
  jor  g05301(.dina(n5493), .dinb(n5492), .dout(n5494));
  jnot g05302(.din(n5494), .dout(n5495));
  jand g05303(.dina(\a[28] ), .dinb(\a[26] ), .dout(n5496));
  jand g05304(.dina(n5496), .dinb(n5048), .dout(n5497));
  jor  g05305(.dina(n5497), .dinb(n5495), .dout(n5498));
  jxor g05306(.dina(n5498), .dinb(n5491), .dout(n5499));
  jand g05307(.dina(\a[31] ), .dinb(\a[22] ), .dout(n5500));
  jand g05308(.dina(\a[30] ), .dinb(\a[23] ), .dout(n5501));
  jor  g05309(.dina(n5501), .dinb(n5230), .dout(n5502));
  jnot g05310(.din(n5502), .dout(n5503));
  jand g05311(.dina(\a[30] ), .dinb(\a[24] ), .dout(n5504));
  jand g05312(.dina(n5504), .dinb(n5087), .dout(n5505));
  jor  g05313(.dina(n5505), .dinb(n5503), .dout(n5506));
  jxor g05314(.dina(n5506), .dinb(n5500), .dout(n5507));
  jand g05315(.dina(\a[40] ), .dinb(\a[13] ), .dout(n5508));
  jand g05316(.dina(\a[43] ), .dinb(\a[10] ), .dout(n5509));
  jor  g05317(.dina(n5509), .dinb(n5067), .dout(n5510));
  jand g05318(.dina(\a[43] ), .dinb(\a[12] ), .dout(n5511));
  jand g05319(.dina(n5511), .dinb(n5064), .dout(n5512));
  jnot g05320(.din(n5512), .dout(n5513));
  jand g05321(.dina(n5513), .dinb(n5510), .dout(n5514));
  jxor g05322(.dina(n5514), .dinb(n5508), .dout(n5515));
  jxor g05323(.dina(n5515), .dinb(n5507), .dout(n5516));
  jxor g05324(.dina(n5516), .dinb(n5499), .dout(n5517));
  jxor g05325(.dina(n5517), .dinb(n5490), .dout(n5518));
  jnot g05326(.din(n5518), .dout(n5519));
  jor  g05327(.dina(n5400), .dinb(n5394), .dout(n5520));
  jand g05328(.dina(n5401), .dinb(n5385), .dout(n5521));
  jnot g05329(.din(n5521), .dout(n5522));
  jand g05330(.dina(n5522), .dinb(n5520), .dout(n5523));
  jxor g05331(.dina(n5523), .dinb(n5519), .dout(n5524));
  jxor g05332(.dina(n5524), .dinb(n5487), .dout(n5525));
  jxor g05333(.dina(n5525), .dinb(n5421), .dout(n5526));
  jxor g05334(.dina(n5526), .dinb(n5418), .dout(n5527));
  jor  g05335(.dina(n5312), .dinb(n5308), .dout(n5528));
  jand g05336(.dina(n5334), .dinb(n5313), .dout(n5529));
  jnot g05337(.din(n5529), .dout(n5530));
  jand g05338(.dina(n5530), .dinb(n5528), .dout(n5531));
  jnot g05339(.din(n5531), .dout(n5532));
  jand g05340(.dina(n5354), .dinb(n5149), .dout(n5533));
  jor  g05341(.dina(n5533), .dinb(n5352), .dout(n5534));
  jand g05342(.dina(n5299), .dinb(n5297), .dout(n5535));
  jor  g05343(.dina(n5535), .dinb(n5302), .dout(n5536));
  jxor g05344(.dina(n5536), .dinb(n5534), .dout(n5537));
  jand g05345(.dina(n5228), .dinb(n5226), .dout(n5538));
  jor  g05346(.dina(n5538), .dinb(n5231), .dout(n5539));
  jxor g05347(.dina(n5539), .dinb(n5537), .dout(n5540));
  jand g05348(.dina(n5242), .dinb(n5234), .dout(n5541));
  jnot g05349(.din(n5541), .dout(n5542));
  jor  g05350(.dina(n5251), .dinb(n5244), .dout(n5543));
  jand g05351(.dina(n5543), .dinb(n5542), .dout(n5544));
  jnot g05352(.din(n5544), .dout(n5545));
  jnot g05353(.din(n5343), .dout(n5546));
  jnot g05354(.din(n5347), .dout(n5547));
  jand g05355(.dina(n5547), .dinb(n5546), .dout(n5548));
  jnot g05356(.din(n5548), .dout(n5549));
  jand g05357(.dina(n5347), .dinb(n5343), .dout(n5550));
  jor  g05358(.dina(n5360), .dinb(n5550), .dout(n5551));
  jand g05359(.dina(n5551), .dinb(n5549), .dout(n5552));
  jxor g05360(.dina(n5552), .dinb(n5545), .dout(n5553));
  jxor g05361(.dina(n5553), .dinb(n5540), .dout(n5554));
  jand g05362(.dina(n5276), .dinb(n5269), .dout(n5555));
  jor  g05363(.dina(n5555), .dinb(n5274), .dout(n5556));
  jand g05364(.dina(n5241), .dinb(n5235), .dout(n5557));
  jor  g05365(.dina(n5557), .dinb(n5239), .dout(n5558));
  jxor g05366(.dina(n5558), .dinb(n5556), .dout(n5559));
  jand g05367(.dina(n5256), .dinb(n5253), .dout(n5560));
  jor  g05368(.dina(n5560), .dinb(n5259), .dout(n5561));
  jxor g05369(.dina(n5561), .dinb(n5559), .dout(n5562));
  jand g05370(.dina(n1654), .dinb(\a[52] ), .dout(n5563));
  jnot g05371(.din(n5563), .dout(n5564));
  jand g05372(.dina(\a[52] ), .dinb(\a[1] ), .dout(n5565));
  jor  g05373(.dina(n5565), .dinb(\a[27] ), .dout(n5566));
  jand g05374(.dina(n5566), .dinb(n5564), .dout(n5567));
  jand g05375(.dina(n5264), .dinb(n5262), .dout(n5568));
  jor  g05376(.dina(n5568), .dinb(n5266), .dout(n5569));
  jxor g05377(.dina(n5569), .dinb(n5567), .dout(n5570));
  jand g05378(.dina(n5247), .dinb(n3553), .dout(n5571));
  jor  g05379(.dina(n5571), .dinb(n5249), .dout(n5572));
  jxor g05380(.dina(n5572), .dinb(n5570), .dout(n5573));
  jnot g05381(.din(n5268), .dout(n5574));
  jor  g05382(.dina(n5277), .dinb(n5574), .dout(n5575));
  jnot g05383(.din(n5261), .dout(n5576));
  jand g05384(.dina(n5277), .dinb(n5574), .dout(n5577));
  jor  g05385(.dina(n5577), .dinb(n5576), .dout(n5578));
  jand g05386(.dina(n5578), .dinb(n5575), .dout(n5579));
  jxor g05387(.dina(n5579), .dinb(n5573), .dout(n5580));
  jxor g05388(.dina(n5580), .dinb(n5562), .dout(n5581));
  jxor g05389(.dina(n5581), .dinb(n5554), .dout(n5582));
  jxor g05390(.dina(n5582), .dinb(n5532), .dout(n5583));
  jand g05391(.dina(n5279), .dinb(n5252), .dout(n5584));
  jand g05392(.dina(n5280), .dinb(n5225), .dout(n5585));
  jor  g05393(.dina(n5585), .dinb(n5584), .dout(n5586));
  jor  g05394(.dina(n5381), .dinb(n5374), .dout(n5587));
  jand g05395(.dina(n5384), .dinb(n5382), .dout(n5588));
  jnot g05396(.din(n5588), .dout(n5589));
  jand g05397(.dina(n5589), .dinb(n5587), .dout(n5590));
  jnot g05398(.din(n5590), .dout(n5591));
  jand g05399(.dina(n5321), .dinb(n5319), .dout(n5592));
  jand g05400(.dina(n5324), .dinb(n5322), .dout(n5593));
  jor  g05401(.dina(n5593), .dinb(n5592), .dout(n5594));
  jxor g05402(.dina(n5594), .dinb(n5591), .dout(n5595));
  jand g05403(.dina(n5389), .dinb(n5387), .dout(n5596));
  jand g05404(.dina(n5392), .dinb(n5390), .dout(n5597));
  jor  g05405(.dina(n5597), .dinb(n5596), .dout(n5598));
  jxor g05406(.dina(n5598), .dinb(n5595), .dout(n5599));
  jnot g05407(.din(n5599), .dout(n5600));
  jand g05408(.dina(n5361), .dinb(n5341), .dout(n5601));
  jnot g05409(.din(n5601), .dout(n5602));
  jor  g05410(.dina(n5367), .dinb(n5363), .dout(n5603));
  jand g05411(.dina(n5603), .dinb(n5602), .dout(n5604));
  jxor g05412(.dina(n5604), .dinb(n5600), .dout(n5605));
  jxor g05413(.dina(n5605), .dinb(n5586), .dout(n5606));
  jand g05414(.dina(n5281), .dinb(n5220), .dout(n5607));
  jand g05415(.dina(n5282), .dinb(n5217), .dout(n5608));
  jor  g05416(.dina(n5608), .dinb(n5607), .dout(n5609));
  jxor g05417(.dina(n5609), .dinb(n5606), .dout(n5610));
  jxor g05418(.dina(n5610), .dinb(n5583), .dout(n5611));
  jxor g05419(.dina(n5611), .dinb(n5527), .dout(n5612));
  jxor g05420(.dina(n5612), .dinb(n5415), .dout(n5613));
  jand g05421(.dina(n5406), .dinb(n5214), .dout(n5614));
  jnot g05422(.din(n5214), .dout(n5615));
  jnot g05423(.din(n5406), .dout(n5616));
  jand g05424(.dina(n5616), .dinb(n5615), .dout(n5617));
  jnot g05425(.din(n5617), .dout(n5618));
  jand g05426(.dina(n5411), .dinb(n5618), .dout(n5619));
  jor  g05427(.dina(n5619), .dinb(n5614), .dout(n5620));
  jxor g05428(.dina(n5620), .dinb(n5613), .dout(\asquared[54] ));
  jand g05429(.dina(n5526), .dinb(n5418), .dout(n5622));
  jand g05430(.dina(n5611), .dinb(n5527), .dout(n5623));
  jor  g05431(.dina(n5623), .dinb(n5622), .dout(n5624));
  jand g05432(.dina(n5609), .dinb(n5606), .dout(n5625));
  jand g05433(.dina(n5610), .dinb(n5583), .dout(n5626));
  jor  g05434(.dina(n5626), .dinb(n5625), .dout(n5627));
  jand g05435(.dina(n5581), .dinb(n5554), .dout(n5628));
  jand g05436(.dina(n5582), .dinb(n5532), .dout(n5629));
  jor  g05437(.dina(n5629), .dinb(n5628), .dout(n5630));
  jnot g05438(.din(n5630), .dout(n5631));
  jor  g05439(.dina(n5604), .dinb(n5600), .dout(n5632));
  jand g05440(.dina(n5605), .dinb(n5586), .dout(n5633));
  jnot g05441(.din(n5633), .dout(n5634));
  jand g05442(.dina(n5634), .dinb(n5632), .dout(n5635));
  jxor g05443(.dina(n5635), .dinb(n5631), .dout(n5636));
  jand g05444(.dina(n5579), .dinb(n5573), .dout(n5637));
  jand g05445(.dina(n5580), .dinb(n5562), .dout(n5638));
  jor  g05446(.dina(n5638), .dinb(n5637), .dout(n5639));
  jand g05447(.dina(n5552), .dinb(n5545), .dout(n5640));
  jand g05448(.dina(n5553), .dinb(n5540), .dout(n5641));
  jor  g05449(.dina(n5641), .dinb(n5640), .dout(n5642));
  jand g05450(.dina(\a[31] ), .dinb(\a[23] ), .dout(n5643));
  jand g05451(.dina(\a[29] ), .dinb(\a[25] ), .dout(n5644));
  jor  g05452(.dina(n5644), .dinb(n5504), .dout(n5645));
  jnot g05453(.din(n5645), .dout(n5646));
  jand g05454(.dina(\a[30] ), .dinb(\a[25] ), .dout(n5647));
  jand g05455(.dina(n5647), .dinb(n5230), .dout(n5648));
  jor  g05456(.dina(n5648), .dinb(n5646), .dout(n5649));
  jxor g05457(.dina(n5649), .dinb(n5643), .dout(n5650));
  jnot g05458(.din(n5650), .dout(n5651));
  jand g05459(.dina(\a[35] ), .dinb(\a[19] ), .dout(n5652));
  jand g05460(.dina(\a[32] ), .dinb(\a[22] ), .dout(n5653));
  jor  g05461(.dina(n5653), .dinb(n5429), .dout(n5654));
  jand g05462(.dina(\a[33] ), .dinb(\a[22] ), .dout(n5655));
  jand g05463(.dina(n5655), .dinb(n5238), .dout(n5656));
  jnot g05464(.din(n5656), .dout(n5657));
  jand g05465(.dina(n5657), .dinb(n5654), .dout(n5658));
  jxor g05466(.dina(n5658), .dinb(n5652), .dout(n5659));
  jxor g05467(.dina(n5659), .dinb(n5651), .dout(n5660));
  jnot g05468(.din(n5660), .dout(n5661));
  jand g05469(.dina(\a[54] ), .dinb(\a[0] ), .dout(n5662));
  jxor g05470(.dina(n5662), .dinb(n5563), .dout(n5663));
  jand g05471(.dina(\a[53] ), .dinb(\a[1] ), .dout(n5664));
  jxor g05472(.dina(n5664), .dinb(n5496), .dout(n5665));
  jnot g05473(.din(n5665), .dout(n5666));
  jxor g05474(.dina(n5666), .dinb(n5663), .dout(n5667));
  jxor g05475(.dina(n5667), .dinb(n5661), .dout(n5668));
  jxor g05476(.dina(n5668), .dinb(n5642), .dout(n5669));
  jxor g05477(.dina(n5669), .dinb(n5639), .dout(n5670));
  jxor g05478(.dina(n5670), .dinb(n5636), .dout(n5671));
  jxor g05479(.dina(n5671), .dinb(n5627), .dout(n5672));
  jand g05480(.dina(n5524), .dinb(n5487), .dout(n5673));
  jand g05481(.dina(n5525), .dinb(n5421), .dout(n5674));
  jor  g05482(.dina(n5674), .dinb(n5673), .dout(n5675));
  jand g05483(.dina(n5558), .dinb(n5556), .dout(n5676));
  jand g05484(.dina(n5561), .dinb(n5559), .dout(n5677));
  jor  g05485(.dina(n5677), .dinb(n5676), .dout(n5678));
  jand g05486(.dina(n5536), .dinb(n5534), .dout(n5679));
  jand g05487(.dina(n5539), .dinb(n5537), .dout(n5680));
  jor  g05488(.dina(n5680), .dinb(n5679), .dout(n5681));
  jxor g05489(.dina(n5681), .dinb(n5678), .dout(n5682));
  jand g05490(.dina(n5569), .dinb(n5567), .dout(n5683));
  jand g05491(.dina(n5572), .dinb(n5570), .dout(n5684));
  jor  g05492(.dina(n5684), .dinb(n5683), .dout(n5685));
  jxor g05493(.dina(n5685), .dinb(n5682), .dout(n5686));
  jand g05494(.dina(n5458), .dinb(n5424), .dout(n5687));
  jand g05495(.dina(n5486), .dinb(n5459), .dout(n5688));
  jor  g05496(.dina(n5688), .dinb(n5687), .dout(n5689));
  jxor g05497(.dina(n5689), .dinb(n5686), .dout(n5690));
  jand g05498(.dina(n5463), .dinb(n5460), .dout(n5691));
  jor  g05499(.dina(n5691), .dinb(n5466), .dout(n5692));
  jnot g05500(.din(n5482), .dout(n5693));
  jand g05501(.dina(n5693), .dinb(n5481), .dout(n5694));
  jnot g05502(.din(n5694), .dout(n5695));
  jand g05503(.dina(n5482), .dinb(n5480), .dout(n5696));
  jor  g05504(.dina(n5696), .dinb(n5479), .dout(n5697));
  jand g05505(.dina(n5697), .dinb(n5695), .dout(n5698));
  jxor g05506(.dina(n5698), .dinb(n5692), .dout(n5699));
  jand g05507(.dina(n5494), .dinb(n5491), .dout(n5700));
  jor  g05508(.dina(n5700), .dinb(n5497), .dout(n5701));
  jxor g05509(.dina(n5701), .dinb(n5699), .dout(n5702));
  jand g05510(.dina(n5438), .dinb(n5434), .dout(n5703));
  jor  g05511(.dina(n5703), .dinb(n5440), .dout(n5704));
  jand g05512(.dina(n5428), .dinb(n5425), .dout(n5705));
  jor  g05513(.dina(n5705), .dinb(n5430), .dout(n5706));
  jxor g05514(.dina(n5706), .dinb(n5704), .dout(n5707));
  jand g05515(.dina(n5502), .dinb(n5500), .dout(n5708));
  jor  g05516(.dina(n5708), .dinb(n5505), .dout(n5709));
  jxor g05517(.dina(n5709), .dinb(n5707), .dout(n5710));
  jnot g05518(.din(n5710), .dout(n5711));
  jor  g05519(.dina(n5484), .dinb(n5478), .dout(n5712));
  jand g05520(.dina(n5485), .dinb(n5469), .dout(n5713));
  jnot g05521(.din(n5713), .dout(n5714));
  jand g05522(.dina(n5714), .dinb(n5712), .dout(n5715));
  jxor g05523(.dina(n5715), .dinb(n5711), .dout(n5716));
  jxor g05524(.dina(n5716), .dinb(n5702), .dout(n5717));
  jxor g05525(.dina(n5717), .dinb(n5690), .dout(n5718));
  jxor g05526(.dina(n5718), .dinb(n5675), .dout(n5719));
  jand g05527(.dina(n5594), .dinb(n5591), .dout(n5720));
  jand g05528(.dina(n5598), .dinb(n5595), .dout(n5721));
  jor  g05529(.dina(n5721), .dinb(n5720), .dout(n5722));
  jand g05530(.dina(\a[37] ), .dinb(\a[17] ), .dout(n5723));
  jnot g05531(.din(n5723), .dout(n5724));
  jand g05532(.dina(\a[48] ), .dinb(\a[6] ), .dout(n5725));
  jand g05533(.dina(\a[38] ), .dinb(\a[16] ), .dout(n5726));
  jor  g05534(.dina(n5726), .dinb(n5725), .dout(n5727));
  jand g05535(.dina(n5465), .dinb(n3818), .dout(n5728));
  jnot g05536(.din(n5728), .dout(n5729));
  jand g05537(.dina(n5729), .dinb(n5727), .dout(n5730));
  jxor g05538(.dina(n5730), .dinb(n5724), .dout(n5731));
  jnot g05539(.din(n4901), .dout(n5732));
  jand g05540(.dina(\a[42] ), .dinb(\a[12] ), .dout(n5733));
  jand g05541(.dina(\a[43] ), .dinb(\a[11] ), .dout(n5734));
  jor  g05542(.dina(n5734), .dinb(n5733), .dout(n5735));
  jand g05543(.dina(n5511), .dinb(n5491), .dout(n5736));
  jnot g05544(.din(n5736), .dout(n5737));
  jand g05545(.dina(n5737), .dinb(n5735), .dout(n5738));
  jxor g05546(.dina(n5738), .dinb(n5732), .dout(n5739));
  jand g05547(.dina(\a[34] ), .dinb(\a[20] ), .dout(n5740));
  jnot g05548(.din(n5740), .dout(n5741));
  jand g05549(.dina(\a[49] ), .dinb(\a[5] ), .dout(n5742));
  jxor g05550(.dina(n5742), .dinb(n5439), .dout(n5743));
  jxor g05551(.dina(n5743), .dinb(n5741), .dout(n5744));
  jnot g05552(.din(n5744), .dout(n5745));
  jxor g05553(.dina(n5745), .dinb(n5739), .dout(n5746));
  jxor g05554(.dina(n5746), .dinb(n5731), .dout(n5747));
  jxor g05555(.dina(n5747), .dinb(n5722), .dout(n5748));
  jand g05556(.dina(\a[47] ), .dinb(\a[7] ), .dout(n5749));
  jand g05557(.dina(\a[39] ), .dinb(\a[15] ), .dout(n5750));
  jand g05558(.dina(n5750), .dinb(n5749), .dout(n5751));
  jand g05559(.dina(\a[47] ), .dinb(\a[8] ), .dout(n5752));
  jand g05560(.dina(n5752), .dinb(n5480), .dout(n5753));
  jor  g05561(.dina(n5753), .dinb(n5751), .dout(n5754));
  jand g05562(.dina(\a[46] ), .dinb(\a[8] ), .dout(n5755));
  jand g05563(.dina(n5755), .dinb(n5750), .dout(n5756));
  jnot g05564(.din(n5756), .dout(n5757));
  jand g05565(.dina(n5757), .dinb(n5754), .dout(n5758));
  jnot g05566(.din(n5758), .dout(n5759));
  jxor g05567(.dina(n5755), .dinb(n5750), .dout(n5760));
  jor  g05568(.dina(n5760), .dinb(n5749), .dout(n5761));
  jand g05569(.dina(n5761), .dinb(n5759), .dout(n5762));
  jand g05570(.dina(\a[52] ), .dinb(\a[2] ), .dout(n5763));
  jand g05571(.dina(\a[50] ), .dinb(\a[4] ), .dout(n5764));
  jor  g05572(.dina(n5764), .dinb(n5452), .dout(n5765));
  jand g05573(.dina(\a[51] ), .dinb(\a[4] ), .dout(n5766));
  jand g05574(.dina(n5766), .dinb(n5301), .dout(n5767));
  jnot g05575(.din(n5767), .dout(n5768));
  jand g05576(.dina(n5768), .dinb(n5765), .dout(n5769));
  jxor g05577(.dina(n5769), .dinb(n5763), .dout(n5770));
  jxor g05578(.dina(n5770), .dinb(n5762), .dout(n5771));
  jnot g05579(.din(n5771), .dout(n5772));
  jand g05580(.dina(\a[45] ), .dinb(\a[9] ), .dout(n5773));
  jand g05581(.dina(\a[40] ), .dinb(\a[14] ), .dout(n5774));
  jand g05582(.dina(\a[44] ), .dinb(\a[10] ), .dout(n5775));
  jor  g05583(.dina(n5775), .dinb(n5774), .dout(n5776));
  jnot g05584(.din(n5776), .dout(n5777));
  jand g05585(.dina(n5473), .dinb(n4890), .dout(n5778));
  jor  g05586(.dina(n5778), .dinb(n5777), .dout(n5779));
  jxor g05587(.dina(n5779), .dinb(n5773), .dout(n5780));
  jxor g05588(.dina(n5780), .dinb(n5772), .dout(n5781));
  jxor g05589(.dina(n5781), .dinb(n5748), .dout(n5782));
  jand g05590(.dina(n5517), .dinb(n5490), .dout(n5783));
  jnot g05591(.din(n5783), .dout(n5784));
  jor  g05592(.dina(n5523), .dinb(n5519), .dout(n5785));
  jand g05593(.dina(n5785), .dinb(n5784), .dout(n5786));
  jnot g05594(.din(n5786), .dout(n5787));
  jand g05595(.dina(n5514), .dinb(n5508), .dout(n5788));
  jor  g05596(.dina(n5788), .dinb(n5512), .dout(n5789));
  jand g05597(.dina(n5476), .dinb(n5258), .dout(n5790));
  jor  g05598(.dina(n5790), .dinb(n5474), .dout(n5791));
  jand g05599(.dina(n5451), .dinb(n5445), .dout(n5792));
  jor  g05600(.dina(n5792), .dinb(n5453), .dout(n5793));
  jxor g05601(.dina(n5793), .dinb(n5791), .dout(n5794));
  jxor g05602(.dina(n5794), .dinb(n5789), .dout(n5795));
  jnot g05603(.din(n5456), .dout(n5796));
  jand g05604(.dina(n5796), .dinb(n5444), .dout(n5797));
  jnot g05605(.din(n5797), .dout(n5798));
  jand g05606(.dina(n5456), .dinb(n5443), .dout(n5799));
  jor  g05607(.dina(n5799), .dinb(n5433), .dout(n5800));
  jand g05608(.dina(n5800), .dinb(n5798), .dout(n5801));
  jnot g05609(.din(n5801), .dout(n5802));
  jnot g05610(.din(n5507), .dout(n5803));
  jor  g05611(.dina(n5515), .dinb(n5803), .dout(n5804));
  jnot g05612(.din(n5499), .dout(n5805));
  jand g05613(.dina(n5515), .dinb(n5803), .dout(n5806));
  jor  g05614(.dina(n5806), .dinb(n5805), .dout(n5807));
  jand g05615(.dina(n5807), .dinb(n5804), .dout(n5808));
  jxor g05616(.dina(n5808), .dinb(n5802), .dout(n5809));
  jxor g05617(.dina(n5809), .dinb(n5795), .dout(n5810));
  jxor g05618(.dina(n5810), .dinb(n5787), .dout(n5811));
  jxor g05619(.dina(n5811), .dinb(n5782), .dout(n5812));
  jxor g05620(.dina(n5812), .dinb(n5719), .dout(n5813));
  jxor g05621(.dina(n5813), .dinb(n5672), .dout(n5814));
  jxor g05622(.dina(n5814), .dinb(n5624), .dout(n5815));
  jand g05623(.dina(n5612), .dinb(n5415), .dout(n5816));
  jor  g05624(.dina(n5612), .dinb(n5415), .dout(n5817));
  jand g05625(.dina(n5620), .dinb(n5817), .dout(n5818));
  jor  g05626(.dina(n5818), .dinb(n5816), .dout(n5819));
  jxor g05627(.dina(n5819), .dinb(n5815), .dout(\asquared[55] ));
  jand g05628(.dina(n5671), .dinb(n5627), .dout(n5821));
  jand g05629(.dina(n5813), .dinb(n5672), .dout(n5822));
  jor  g05630(.dina(n5822), .dinb(n5821), .dout(n5823));
  jor  g05631(.dina(n5635), .dinb(n5631), .dout(n5824));
  jand g05632(.dina(n5670), .dinb(n5636), .dout(n5825));
  jnot g05633(.din(n5825), .dout(n5826));
  jand g05634(.dina(n5826), .dinb(n5824), .dout(n5827));
  jnot g05635(.din(n5827), .dout(n5828));
  jand g05636(.dina(n5747), .dinb(n5722), .dout(n5829));
  jand g05637(.dina(n5781), .dinb(n5748), .dout(n5830));
  jor  g05638(.dina(n5830), .dinb(n5829), .dout(n5831));
  jand g05639(.dina(n5698), .dinb(n5692), .dout(n5832));
  jand g05640(.dina(n5701), .dinb(n5699), .dout(n5833));
  jor  g05641(.dina(n5833), .dinb(n5832), .dout(n5834));
  jand g05642(.dina(n5793), .dinb(n5791), .dout(n5835));
  jand g05643(.dina(n5794), .dinb(n5789), .dout(n5836));
  jor  g05644(.dina(n5836), .dinb(n5835), .dout(n5837));
  jxor g05645(.dina(n5837), .dinb(n5834), .dout(n5838));
  jand g05646(.dina(n5735), .dinb(n4901), .dout(n5839));
  jor  g05647(.dina(n5839), .dinb(n5736), .dout(n5840));
  jnot g05648(.din(\a[54] ), .dout(n5841));
  jand g05649(.dina(n5664), .dinb(n5496), .dout(n5842));
  jand g05650(.dina(n5842), .dinb(n5841), .dout(n5843));
  jnot g05651(.din(n5843), .dout(n5844));
  jand g05652(.dina(\a[54] ), .dinb(\a[28] ), .dout(n5845));
  jand g05653(.dina(n5845), .dinb(\a[1] ), .dout(n5846));
  jnot g05654(.din(n5846), .dout(n5847));
  jand g05655(.dina(\a[54] ), .dinb(\a[1] ), .dout(n5848));
  jor  g05656(.dina(n5848), .dinb(\a[28] ), .dout(n5849));
  jand g05657(.dina(n5849), .dinb(n5847), .dout(n5850));
  jor  g05658(.dina(n5850), .dinb(n5842), .dout(n5851));
  jand g05659(.dina(n5851), .dinb(n5844), .dout(n5852));
  jxor g05660(.dina(n5852), .dinb(n5840), .dout(n5853));
  jxor g05661(.dina(n5853), .dinb(n5838), .dout(n5854));
  jxor g05662(.dina(n5854), .dinb(n5831), .dout(n5855));
  jand g05663(.dina(n5769), .dinb(n5763), .dout(n5856));
  jor  g05664(.dina(n5856), .dinb(n5767), .dout(n5857));
  jand g05665(.dina(n5776), .dinb(n5773), .dout(n5858));
  jor  g05666(.dina(n5858), .dinb(n5778), .dout(n5859));
  jxor g05667(.dina(n5859), .dinb(n5857), .dout(n5860));
  jnot g05668(.din(n5860), .dout(n5861));
  jand g05669(.dina(n5742), .dinb(n5439), .dout(n5862));
  jnot g05670(.din(n5862), .dout(n5863));
  jnot g05671(.din(n5439), .dout(n5864));
  jnot g05672(.din(n5742), .dout(n5865));
  jand g05673(.dina(n5865), .dinb(n5864), .dout(n5866));
  jor  g05674(.dina(n5866), .dinb(n5741), .dout(n5867));
  jand g05675(.dina(n5867), .dinb(n5863), .dout(n5868));
  jxor g05676(.dina(n5868), .dinb(n5861), .dout(n5869));
  jnot g05677(.din(n5869), .dout(n5870));
  jand g05678(.dina(n5659), .dinb(n5651), .dout(n5871));
  jnot g05679(.din(n5871), .dout(n5872));
  jor  g05680(.dina(n5667), .dinb(n5661), .dout(n5873));
  jand g05681(.dina(n5873), .dinb(n5872), .dout(n5874));
  jxor g05682(.dina(n5874), .dinb(n5870), .dout(n5875));
  jor  g05683(.dina(n5756), .dinb(n5754), .dout(n5876));
  jnot g05684(.din(n5876), .dout(n5877));
  jand g05685(.dina(n5662), .dinb(n5563), .dout(n5878));
  jnot g05686(.din(n5878), .dout(n5879));
  jnot g05687(.din(n5662), .dout(n5880));
  jand g05688(.dina(n5880), .dinb(n5564), .dout(n5881));
  jor  g05689(.dina(n5666), .dinb(n5881), .dout(n5882));
  jand g05690(.dina(n5882), .dinb(n5879), .dout(n5883));
  jxor g05691(.dina(n5883), .dinb(n5877), .dout(n5884));
  jand g05692(.dina(\a[50] ), .dinb(\a[5] ), .dout(n5885));
  jand g05693(.dina(\a[37] ), .dinb(\a[18] ), .dout(n5886));
  jand g05694(.dina(\a[36] ), .dinb(\a[19] ), .dout(n5887));
  jor  g05695(.dina(n5887), .dinb(n5886), .dout(n5888));
  jnot g05696(.din(n5888), .dout(n5889));
  jand g05697(.dina(\a[37] ), .dinb(\a[19] ), .dout(n5890));
  jand g05698(.dina(n5890), .dinb(n5439), .dout(n5891));
  jor  g05699(.dina(n5891), .dinb(n5889), .dout(n5892));
  jxor g05700(.dina(n5892), .dinb(n5885), .dout(n5893));
  jnot g05701(.din(n5893), .dout(n5894));
  jxor g05702(.dina(n5894), .dinb(n5884), .dout(n5895));
  jxor g05703(.dina(n5895), .dinb(n5875), .dout(n5896));
  jxor g05704(.dina(n5896), .dinb(n5855), .dout(n5897));
  jxor g05705(.dina(n5897), .dinb(n5828), .dout(n5898));
  jand g05706(.dina(n5668), .dinb(n5642), .dout(n5899));
  jand g05707(.dina(n5669), .dinb(n5639), .dout(n5900));
  jor  g05708(.dina(n5900), .dinb(n5899), .dout(n5901));
  jand g05709(.dina(n5658), .dinb(n5652), .dout(n5902));
  jor  g05710(.dina(n5902), .dinb(n5656), .dout(n5903));
  jand g05711(.dina(n5645), .dinb(n5643), .dout(n5904));
  jor  g05712(.dina(n5904), .dinb(n5648), .dout(n5905));
  jxor g05713(.dina(n5905), .dinb(n5903), .dout(n5906));
  jand g05714(.dina(n5727), .dinb(n5723), .dout(n5907));
  jor  g05715(.dina(n5907), .dinb(n5728), .dout(n5908));
  jxor g05716(.dina(n5908), .dinb(n5906), .dout(n5909));
  jand g05717(.dina(n5770), .dinb(n5762), .dout(n5910));
  jnot g05718(.din(n5910), .dout(n5911));
  jor  g05719(.dina(n5780), .dinb(n5772), .dout(n5912));
  jand g05720(.dina(n5912), .dinb(n5911), .dout(n5913));
  jnot g05721(.din(n5739), .dout(n5914));
  jand g05722(.dina(n5745), .dinb(n5914), .dout(n5915));
  jnot g05723(.din(n5915), .dout(n5916));
  jand g05724(.dina(n5744), .dinb(n5739), .dout(n5917));
  jor  g05725(.dina(n5917), .dinb(n5731), .dout(n5918));
  jand g05726(.dina(n5918), .dinb(n5916), .dout(n5919));
  jxor g05727(.dina(n5919), .dinb(n5913), .dout(n5920));
  jxor g05728(.dina(n5920), .dinb(n5909), .dout(n5921));
  jxor g05729(.dina(n5921), .dinb(n5901), .dout(n5922));
  jand g05730(.dina(n5681), .dinb(n5678), .dout(n5923));
  jand g05731(.dina(n5685), .dinb(n5682), .dout(n5924));
  jor  g05732(.dina(n5924), .dinb(n5923), .dout(n5925));
  jand g05733(.dina(\a[39] ), .dinb(\a[16] ), .dout(n5926));
  jand g05734(.dina(\a[48] ), .dinb(\a[7] ), .dout(n5927));
  jor  g05735(.dina(n5927), .dinb(n5752), .dout(n5928));
  jnot g05736(.din(n5928), .dout(n5929));
  jand g05737(.dina(\a[48] ), .dinb(\a[8] ), .dout(n5930));
  jand g05738(.dina(n5930), .dinb(n5749), .dout(n5931));
  jor  g05739(.dina(n5931), .dinb(n5929), .dout(n5932));
  jxor g05740(.dina(n5932), .dinb(n5926), .dout(n5933));
  jnot g05741(.din(n5933), .dout(n5934));
  jand g05742(.dina(\a[28] ), .dinb(\a[27] ), .dout(n5935));
  jnot g05743(.din(n5935), .dout(n5936));
  jand g05744(.dina(\a[29] ), .dinb(\a[26] ), .dout(n5937));
  jxor g05745(.dina(n5937), .dinb(n5936), .dout(n5938));
  jxor g05746(.dina(n5938), .dinb(n5511), .dout(n5939));
  jnot g05747(.din(n5939), .dout(n5940));
  jand g05748(.dina(\a[45] ), .dinb(\a[10] ), .dout(n5941));
  jand g05749(.dina(\a[42] ), .dinb(\a[13] ), .dout(n5942));
  jand g05750(.dina(\a[44] ), .dinb(\a[11] ), .dout(n5943));
  jor  g05751(.dina(n5943), .dinb(n5942), .dout(n5944));
  jand g05752(.dina(\a[44] ), .dinb(\a[13] ), .dout(n5945));
  jand g05753(.dina(n5945), .dinb(n5491), .dout(n5946));
  jnot g05754(.din(n5946), .dout(n5947));
  jand g05755(.dina(n5947), .dinb(n5944), .dout(n5948));
  jxor g05756(.dina(n5948), .dinb(n5941), .dout(n5949));
  jxor g05757(.dina(n5949), .dinb(n5940), .dout(n5950));
  jxor g05758(.dina(n5950), .dinb(n5934), .dout(n5951));
  jxor g05759(.dina(n5951), .dinb(n5925), .dout(n5952));
  jand g05760(.dina(\a[32] ), .dinb(\a[23] ), .dout(n5953));
  jnot g05761(.din(n5953), .dout(n5954));
  jand g05762(.dina(\a[31] ), .dinb(\a[24] ), .dout(n5955));
  jor  g05763(.dina(n5955), .dinb(n5647), .dout(n5956));
  jand g05764(.dina(\a[31] ), .dinb(\a[25] ), .dout(n5957));
  jand g05765(.dina(n5957), .dinb(n5504), .dout(n5958));
  jnot g05766(.din(n5958), .dout(n5959));
  jand g05767(.dina(n5959), .dinb(n5956), .dout(n5960));
  jxor g05768(.dina(n5960), .dinb(n5954), .dout(n5961));
  jand g05769(.dina(\a[35] ), .dinb(\a[20] ), .dout(n5962));
  jnot g05770(.din(n5962), .dout(n5963));
  jand g05771(.dina(\a[34] ), .dinb(\a[21] ), .dout(n5964));
  jor  g05772(.dina(n5964), .dinb(n5655), .dout(n5965));
  jand g05773(.dina(\a[34] ), .dinb(\a[22] ), .dout(n5966));
  jand g05774(.dina(n5966), .dinb(n5429), .dout(n5967));
  jnot g05775(.din(n5967), .dout(n5968));
  jand g05776(.dina(n5968), .dinb(n5965), .dout(n5969));
  jxor g05777(.dina(n5969), .dinb(n5963), .dout(n5970));
  jand g05778(.dina(n208), .dinb(\a[51] ), .dout(n5971));
  jand g05779(.dina(\a[53] ), .dinb(\a[2] ), .dout(n5972));
  jand g05780(.dina(n5972), .dinb(\a[0] ), .dout(n5973));
  jor  g05781(.dina(n5973), .dinb(n5971), .dout(n5974));
  jand g05782(.dina(n5974), .dinb(\a[55] ), .dout(n5975));
  jnot g05783(.din(n5975), .dout(n5976));
  jor  g05784(.dina(n5972), .dinb(n5766), .dout(n5977));
  jand g05785(.dina(\a[53] ), .dinb(\a[4] ), .dout(n5978));
  jand g05786(.dina(n5978), .dinb(n5448), .dout(n5979));
  jnot g05787(.din(n5979), .dout(n5980));
  jand g05788(.dina(n5980), .dinb(n5977), .dout(n5981));
  jand g05789(.dina(n5981), .dinb(n5976), .dout(n5982));
  jnot g05790(.din(n5981), .dout(n5983));
  jand g05791(.dina(\a[55] ), .dinb(\a[0] ), .dout(n5984));
  jand g05792(.dina(n5984), .dinb(n5983), .dout(n5985));
  jor  g05793(.dina(n5985), .dinb(n5982), .dout(n5986));
  jxor g05794(.dina(n5986), .dinb(n5970), .dout(n5987));
  jxor g05795(.dina(n5987), .dinb(n5961), .dout(n5988));
  jxor g05796(.dina(n5988), .dinb(n5952), .dout(n5989));
  jxor g05797(.dina(n5989), .dinb(n5922), .dout(n5990));
  jxor g05798(.dina(n5990), .dinb(n5898), .dout(n5991));
  jand g05799(.dina(n5718), .dinb(n5675), .dout(n5992));
  jand g05800(.dina(n5812), .dinb(n5719), .dout(n5993));
  jor  g05801(.dina(n5993), .dinb(n5992), .dout(n5994));
  jand g05802(.dina(n5810), .dinb(n5787), .dout(n5995));
  jand g05803(.dina(n5811), .dinb(n5782), .dout(n5996));
  jor  g05804(.dina(n5996), .dinb(n5995), .dout(n5997));
  jand g05805(.dina(n5689), .dinb(n5686), .dout(n5998));
  jand g05806(.dina(n5717), .dinb(n5690), .dout(n5999));
  jor  g05807(.dina(n5999), .dinb(n5998), .dout(n6000));
  jor  g05808(.dina(n5715), .dinb(n5711), .dout(n6001));
  jand g05809(.dina(n5716), .dinb(n5702), .dout(n6002));
  jnot g05810(.din(n6002), .dout(n6003));
  jand g05811(.dina(n6003), .dinb(n6001), .dout(n6004));
  jnot g05812(.din(n6004), .dout(n6005));
  jand g05813(.dina(n5706), .dinb(n5704), .dout(n6006));
  jand g05814(.dina(n5709), .dinb(n5707), .dout(n6007));
  jor  g05815(.dina(n6007), .dinb(n6006), .dout(n6008));
  jand g05816(.dina(\a[40] ), .dinb(\a[15] ), .dout(n6009));
  jnot g05817(.din(n6009), .dout(n6010));
  jand g05818(.dina(\a[46] ), .dinb(\a[9] ), .dout(n6011));
  jxor g05819(.dina(n6011), .dinb(n4388), .dout(n6012));
  jxor g05820(.dina(n6012), .dinb(n6010), .dout(n6013));
  jnot g05821(.din(n6013), .dout(n6014));
  jand g05822(.dina(\a[52] ), .dinb(\a[3] ), .dout(n6015));
  jand g05823(.dina(\a[49] ), .dinb(\a[6] ), .dout(n6016));
  jand g05824(.dina(\a[38] ), .dinb(\a[17] ), .dout(n6017));
  jor  g05825(.dina(n6017), .dinb(n6016), .dout(n6018));
  jand g05826(.dina(\a[49] ), .dinb(\a[17] ), .dout(n6019));
  jand g05827(.dina(n6019), .dinb(n3818), .dout(n6020));
  jnot g05828(.din(n6020), .dout(n6021));
  jand g05829(.dina(n6021), .dinb(n6018), .dout(n6022));
  jxor g05830(.dina(n6022), .dinb(n6015), .dout(n6023));
  jxor g05831(.dina(n6023), .dinb(n6014), .dout(n6024));
  jxor g05832(.dina(n6024), .dinb(n6008), .dout(n6025));
  jand g05833(.dina(n5808), .dinb(n5802), .dout(n6026));
  jand g05834(.dina(n5809), .dinb(n5795), .dout(n6027));
  jor  g05835(.dina(n6027), .dinb(n6026), .dout(n6028));
  jxor g05836(.dina(n6028), .dinb(n6025), .dout(n6029));
  jxor g05837(.dina(n6029), .dinb(n6005), .dout(n6030));
  jxor g05838(.dina(n6030), .dinb(n6000), .dout(n6031));
  jxor g05839(.dina(n6031), .dinb(n5997), .dout(n6032));
  jxor g05840(.dina(n6032), .dinb(n5994), .dout(n6033));
  jxor g05841(.dina(n6033), .dinb(n5991), .dout(n6034));
  jxor g05842(.dina(n6034), .dinb(n5823), .dout(n6035));
  jand g05843(.dina(n5814), .dinb(n5624), .dout(n6036));
  jor  g05844(.dina(n5814), .dinb(n5624), .dout(n6037));
  jand g05845(.dina(n5819), .dinb(n6037), .dout(n6038));
  jor  g05846(.dina(n6038), .dinb(n6036), .dout(n6039));
  jxor g05847(.dina(n6039), .dinb(n6035), .dout(\asquared[56] ));
  jand g05848(.dina(n6032), .dinb(n5994), .dout(n6041));
  jand g05849(.dina(n6033), .dinb(n5991), .dout(n6042));
  jor  g05850(.dina(n6042), .dinb(n6041), .dout(n6043));
  jand g05851(.dina(\a[40] ), .dinb(\a[16] ), .dout(n6044));
  jnot g05852(.din(n6044), .dout(n6045));
  jor  g05853(.dina(n5930), .dinb(n4128), .dout(n6046));
  jand g05854(.dina(\a[48] ), .dinb(\a[15] ), .dout(n6047));
  jand g05855(.dina(n6047), .dinb(n4704), .dout(n6048));
  jnot g05856(.din(n6048), .dout(n6049));
  jand g05857(.dina(n6049), .dinb(n6046), .dout(n6050));
  jxor g05858(.dina(n6050), .dinb(n6045), .dout(n6051));
  jand g05859(.dina(\a[45] ), .dinb(\a[11] ), .dout(n6052));
  jnot g05860(.din(n6052), .dout(n6053));
  jand g05861(.dina(\a[44] ), .dinb(\a[12] ), .dout(n6054));
  jor  g05862(.dina(n6054), .dinb(n5057), .dout(n6055));
  jand g05863(.dina(n5945), .dinb(n5511), .dout(n6056));
  jnot g05864(.din(n6056), .dout(n6057));
  jand g05865(.dina(n6057), .dinb(n6055), .dout(n6058));
  jxor g05866(.dina(n6058), .dinb(n6053), .dout(n6059));
  jand g05867(.dina(\a[50] ), .dinb(\a[6] ), .dout(n6060));
  jnot g05868(.din(n6060), .dout(n6061));
  jand g05869(.dina(\a[49] ), .dinb(\a[7] ), .dout(n6062));
  jand g05870(.dina(\a[39] ), .dinb(\a[17] ), .dout(n6063));
  jxor g05871(.dina(n6063), .dinb(n6062), .dout(n6064));
  jxor g05872(.dina(n6064), .dinb(n6061), .dout(n6065));
  jnot g05873(.din(n6065), .dout(n6066));
  jxor g05874(.dina(n6066), .dinb(n6059), .dout(n6067));
  jxor g05875(.dina(n6067), .dinb(n6051), .dout(n6068));
  jand g05876(.dina(\a[47] ), .dinb(\a[9] ), .dout(n6069));
  jand g05877(.dina(\a[42] ), .dinb(\a[14] ), .dout(n6070));
  jand g05878(.dina(\a[46] ), .dinb(\a[10] ), .dout(n6071));
  jor  g05879(.dina(n6071), .dinb(n6070), .dout(n6072));
  jnot g05880(.din(n6072), .dout(n6073));
  jand g05881(.dina(\a[46] ), .dinb(\a[14] ), .dout(n6074));
  jand g05882(.dina(n6074), .dinb(n5262), .dout(n6075));
  jor  g05883(.dina(n6075), .dinb(n6073), .dout(n6076));
  jxor g05884(.dina(n6076), .dinb(n6069), .dout(n6077));
  jand g05885(.dina(\a[32] ), .dinb(\a[24] ), .dout(n6078));
  jand g05886(.dina(\a[30] ), .dinb(\a[26] ), .dout(n6079));
  jor  g05887(.dina(n6079), .dinb(n5957), .dout(n6080));
  jnot g05888(.din(n6080), .dout(n6081));
  jand g05889(.dina(\a[31] ), .dinb(\a[26] ), .dout(n6082));
  jand g05890(.dina(n6082), .dinb(n5647), .dout(n6083));
  jor  g05891(.dina(n6083), .dinb(n6081), .dout(n6084));
  jxor g05892(.dina(n6084), .dinb(n6078), .dout(n6085));
  jand g05893(.dina(\a[36] ), .dinb(\a[20] ), .dout(n6086));
  jand g05894(.dina(\a[33] ), .dinb(\a[23] ), .dout(n6087));
  jor  g05895(.dina(n6087), .dinb(n5966), .dout(n6088));
  jand g05896(.dina(\a[34] ), .dinb(\a[23] ), .dout(n6089));
  jand g05897(.dina(n6089), .dinb(n5655), .dout(n6090));
  jnot g05898(.din(n6090), .dout(n6091));
  jand g05899(.dina(n6091), .dinb(n6088), .dout(n6092));
  jxor g05900(.dina(n6092), .dinb(n6086), .dout(n6093));
  jxor g05901(.dina(n6093), .dinb(n6085), .dout(n6094));
  jxor g05902(.dina(n6094), .dinb(n6077), .dout(n6095));
  jxor g05903(.dina(n6095), .dinb(n6068), .dout(n6096));
  jand g05904(.dina(\a[56] ), .dinb(\a[0] ), .dout(n6097));
  jand g05905(.dina(\a[54] ), .dinb(\a[2] ), .dout(n6098));
  jor  g05906(.dina(n6098), .dinb(n6097), .dout(n6099));
  jand g05907(.dina(\a[56] ), .dinb(\a[2] ), .dout(n6100));
  jand g05908(.dina(n6100), .dinb(n5662), .dout(n6101));
  jnot g05909(.din(n6101), .dout(n6102));
  jand g05910(.dina(n6102), .dinb(n6099), .dout(n6103));
  jxor g05911(.dina(n6103), .dinb(n5846), .dout(n6104));
  jand g05912(.dina(n5928), .dinb(n5926), .dout(n6105));
  jor  g05913(.dina(n6105), .dinb(n5931), .dout(n6106));
  jxor g05914(.dina(n6106), .dinb(n6104), .dout(n6107));
  jand g05915(.dina(\a[53] ), .dinb(\a[3] ), .dout(n6108));
  jnot g05916(.din(n6108), .dout(n6109));
  jand g05917(.dina(\a[52] ), .dinb(\a[4] ), .dout(n6110));
  jxor g05918(.dina(n6110), .dinb(n5890), .dout(n6111));
  jxor g05919(.dina(n6111), .dinb(n6109), .dout(n6112));
  jnot g05920(.din(n6112), .dout(n6113));
  jxor g05921(.dina(n6113), .dinb(n6107), .dout(n6114));
  jxor g05922(.dina(n6114), .dinb(n6096), .dout(n6115));
  jand g05923(.dina(n6028), .dinb(n6025), .dout(n6116));
  jand g05924(.dina(n6029), .dinb(n6005), .dout(n6117));
  jor  g05925(.dina(n6117), .dinb(n6116), .dout(n6118));
  jand g05926(.dina(n6022), .dinb(n6015), .dout(n6119));
  jor  g05927(.dina(n6119), .dinb(n6020), .dout(n6120));
  jand g05928(.dina(n5965), .dinb(n5962), .dout(n6121));
  jor  g05929(.dina(n6121), .dinb(n5967), .dout(n6122));
  jand g05930(.dina(n5956), .dinb(n5953), .dout(n6123));
  jor  g05931(.dina(n6123), .dinb(n5958), .dout(n6124));
  jxor g05932(.dina(n6124), .dinb(n6122), .dout(n6125));
  jxor g05933(.dina(n6125), .dinb(n6120), .dout(n6126));
  jand g05934(.dina(n5948), .dinb(n5941), .dout(n6127));
  jor  g05935(.dina(n6127), .dinb(n5946), .dout(n6128));
  jand g05936(.dina(\a[29] ), .dinb(\a[27] ), .dout(n6129));
  jand g05937(.dina(\a[55] ), .dinb(\a[1] ), .dout(n6130));
  jxor g05938(.dina(n6130), .dinb(n6129), .dout(n6131));
  jnot g05939(.din(n5937), .dout(n6132));
  jand g05940(.dina(n6132), .dinb(n5936), .dout(n6133));
  jnot g05941(.din(n6133), .dout(n6134));
  jand g05942(.dina(n5937), .dinb(n5935), .dout(n6135));
  jor  g05943(.dina(n6135), .dinb(n5511), .dout(n6136));
  jand g05944(.dina(n6136), .dinb(n6134), .dout(n6137));
  jxor g05945(.dina(n6137), .dinb(n6131), .dout(n6138));
  jxor g05946(.dina(n6138), .dinb(n6128), .dout(n6139));
  jor  g05947(.dina(n5949), .dinb(n5940), .dout(n6140));
  jand g05948(.dina(n5949), .dinb(n5940), .dout(n6141));
  jor  g05949(.dina(n6141), .dinb(n5934), .dout(n6142));
  jand g05950(.dina(n6142), .dinb(n6140), .dout(n6143));
  jxor g05951(.dina(n6143), .dinb(n6139), .dout(n6144));
  jxor g05952(.dina(n6144), .dinb(n6126), .dout(n6145));
  jxor g05953(.dina(n6145), .dinb(n6118), .dout(n6146));
  jxor g05954(.dina(n6146), .dinb(n6115), .dout(n6147));
  jand g05955(.dina(n6030), .dinb(n6000), .dout(n6148));
  jand g05956(.dina(n6031), .dinb(n5997), .dout(n6149));
  jor  g05957(.dina(n6149), .dinb(n6148), .dout(n6150));
  jand g05958(.dina(n5980), .dinb(n5976), .dout(n6151));
  jnot g05959(.din(n6151), .dout(n6152));
  jand g05960(.dina(n5888), .dinb(n5885), .dout(n6153));
  jor  g05961(.dina(n6153), .dinb(n5891), .dout(n6154));
  jxor g05962(.dina(n6154), .dinb(n6152), .dout(n6155));
  jnot g05963(.din(n6155), .dout(n6156));
  jand g05964(.dina(n6011), .dinb(n4388), .dout(n6157));
  jnot g05965(.din(n6157), .dout(n6158));
  jnot g05966(.din(n4388), .dout(n6159));
  jnot g05967(.din(n6011), .dout(n6160));
  jand g05968(.dina(n6160), .dinb(n6159), .dout(n6161));
  jor  g05969(.dina(n6161), .dinb(n6010), .dout(n6162));
  jand g05970(.dina(n6162), .dinb(n6158), .dout(n6163));
  jxor g05971(.dina(n6163), .dinb(n6156), .dout(n6164));
  jand g05972(.dina(n6023), .dinb(n6014), .dout(n6165));
  jand g05973(.dina(n6024), .dinb(n6008), .dout(n6166));
  jor  g05974(.dina(n6166), .dinb(n6165), .dout(n6167));
  jxor g05975(.dina(n6167), .dinb(n6164), .dout(n6168));
  jand g05976(.dina(n5837), .dinb(n5834), .dout(n6169));
  jand g05977(.dina(n5853), .dinb(n5838), .dout(n6170));
  jor  g05978(.dina(n6170), .dinb(n6169), .dout(n6171));
  jxor g05979(.dina(n6171), .dinb(n6168), .dout(n6172));
  jand g05980(.dina(n5905), .dinb(n5903), .dout(n6173));
  jand g05981(.dina(n5908), .dinb(n5906), .dout(n6174));
  jor  g05982(.dina(n6174), .dinb(n6173), .dout(n6175));
  jand g05983(.dina(n5883), .dinb(n5877), .dout(n6176));
  jnot g05984(.din(n6176), .dout(n6177));
  jnot g05985(.din(n5883), .dout(n6178));
  jand g05986(.dina(n6178), .dinb(n5876), .dout(n6179));
  jor  g05987(.dina(n5894), .dinb(n6179), .dout(n6180));
  jand g05988(.dina(n6180), .dinb(n6177), .dout(n6181));
  jxor g05989(.dina(n6181), .dinb(n6175), .dout(n6182));
  jnot g05990(.din(n6182), .dout(n6183));
  jnot g05991(.din(n5970), .dout(n6184));
  jand g05992(.dina(n5986), .dinb(n6184), .dout(n6185));
  jnot g05993(.din(n6185), .dout(n6186));
  jnot g05994(.din(n5986), .dout(n6187));
  jand g05995(.dina(n6187), .dinb(n5970), .dout(n6188));
  jor  g05996(.dina(n6188), .dinb(n5961), .dout(n6189));
  jand g05997(.dina(n6189), .dinb(n6186), .dout(n6190));
  jxor g05998(.dina(n6190), .dinb(n6183), .dout(n6191));
  jand g05999(.dina(n5951), .dinb(n5925), .dout(n6192));
  jand g06000(.dina(n5988), .dinb(n5952), .dout(n6193));
  jor  g06001(.dina(n6193), .dinb(n6192), .dout(n6194));
  jxor g06002(.dina(n6194), .dinb(n6191), .dout(n6195));
  jxor g06003(.dina(n6195), .dinb(n6172), .dout(n6196));
  jxor g06004(.dina(n6196), .dinb(n6150), .dout(n6197));
  jxor g06005(.dina(n6197), .dinb(n6147), .dout(n6198));
  jand g06006(.dina(n5859), .dinb(n5857), .dout(n6199));
  jnot g06007(.din(n6199), .dout(n6200));
  jor  g06008(.dina(n5868), .dinb(n5861), .dout(n6201));
  jand g06009(.dina(n6201), .dinb(n6200), .dout(n6202));
  jnot g06010(.din(n6202), .dout(n6203));
  jand g06011(.dina(n5852), .dinb(n5840), .dout(n6204));
  jor  g06012(.dina(n6204), .dinb(n5843), .dout(n6205));
  jnot g06013(.din(n6205), .dout(n6206));
  jand g06014(.dina(\a[35] ), .dinb(\a[21] ), .dout(n6207));
  jand g06015(.dina(\a[51] ), .dinb(\a[5] ), .dout(n6208));
  jand g06016(.dina(\a[38] ), .dinb(\a[18] ), .dout(n6209));
  jor  g06017(.dina(n6209), .dinb(n6208), .dout(n6210));
  jnot g06018(.din(n6210), .dout(n6211));
  jand g06019(.dina(\a[51] ), .dinb(\a[18] ), .dout(n6212));
  jand g06020(.dina(n6212), .dinb(n3644), .dout(n6213));
  jor  g06021(.dina(n6213), .dinb(n6211), .dout(n6214));
  jxor g06022(.dina(n6214), .dinb(n6207), .dout(n6215));
  jxor g06023(.dina(n6215), .dinb(n6206), .dout(n6216));
  jxor g06024(.dina(n6216), .dinb(n6203), .dout(n6217));
  jnot g06025(.din(n6217), .dout(n6218));
  jor  g06026(.dina(n5919), .dinb(n5913), .dout(n6219));
  jand g06027(.dina(n5920), .dinb(n5909), .dout(n6220));
  jnot g06028(.din(n6220), .dout(n6221));
  jand g06029(.dina(n6221), .dinb(n6219), .dout(n6222));
  jxor g06030(.dina(n6222), .dinb(n6218), .dout(n6223));
  jand g06031(.dina(n5874), .dinb(n5870), .dout(n6224));
  jnot g06032(.din(n6224), .dout(n6225));
  jnot g06033(.din(n5874), .dout(n6226));
  jand g06034(.dina(n6226), .dinb(n5869), .dout(n6227));
  jor  g06035(.dina(n5895), .dinb(n6227), .dout(n6228));
  jand g06036(.dina(n6228), .dinb(n6225), .dout(n6229));
  jxor g06037(.dina(n6229), .dinb(n6223), .dout(n6230));
  jor  g06038(.dina(n5854), .dinb(n5831), .dout(n6231));
  jand g06039(.dina(n5854), .dinb(n5831), .dout(n6232));
  jor  g06040(.dina(n5896), .dinb(n6232), .dout(n6233));
  jand g06041(.dina(n6233), .dinb(n6231), .dout(n6234));
  jxor g06042(.dina(n6234), .dinb(n6230), .dout(n6235));
  jand g06043(.dina(n5921), .dinb(n5901), .dout(n6236));
  jand g06044(.dina(n5989), .dinb(n5922), .dout(n6237));
  jor  g06045(.dina(n6237), .dinb(n6236), .dout(n6238));
  jxor g06046(.dina(n6238), .dinb(n6235), .dout(n6239));
  jand g06047(.dina(n5897), .dinb(n5828), .dout(n6240));
  jand g06048(.dina(n5990), .dinb(n5898), .dout(n6241));
  jor  g06049(.dina(n6241), .dinb(n6240), .dout(n6242));
  jxor g06050(.dina(n6242), .dinb(n6239), .dout(n6243));
  jxor g06051(.dina(n6243), .dinb(n6198), .dout(n6244));
  jxor g06052(.dina(n6244), .dinb(n6043), .dout(n6245));
  jand g06053(.dina(n6034), .dinb(n5823), .dout(n6246));
  jor  g06054(.dina(n6034), .dinb(n5823), .dout(n6247));
  jand g06055(.dina(n6039), .dinb(n6247), .dout(n6248));
  jor  g06056(.dina(n6248), .dinb(n6246), .dout(n6249));
  jxor g06057(.dina(n6249), .dinb(n6245), .dout(\asquared[57] ));
  jand g06058(.dina(n6242), .dinb(n6239), .dout(n6251));
  jand g06059(.dina(n6243), .dinb(n6198), .dout(n6252));
  jor  g06060(.dina(n6252), .dinb(n6251), .dout(n6253));
  jand g06061(.dina(n6234), .dinb(n6230), .dout(n6254));
  jand g06062(.dina(n6238), .dinb(n6235), .dout(n6255));
  jor  g06063(.dina(n6255), .dinb(n6254), .dout(n6256));
  jand g06064(.dina(n6137), .dinb(n6131), .dout(n6257));
  jand g06065(.dina(n6138), .dinb(n6128), .dout(n6258));
  jor  g06066(.dina(n6258), .dinb(n6257), .dout(n6259));
  jnot g06067(.din(n6104), .dout(n6260));
  jnot g06068(.din(n6106), .dout(n6261));
  jand g06069(.dina(n6261), .dinb(n6260), .dout(n6262));
  jnot g06070(.din(n6262), .dout(n6263));
  jand g06071(.dina(n6106), .dinb(n6104), .dout(n6264));
  jor  g06072(.dina(n6113), .dinb(n6264), .dout(n6265));
  jand g06073(.dina(n6265), .dinb(n6263), .dout(n6266));
  jxor g06074(.dina(n6266), .dinb(n6259), .dout(n6267));
  jnot g06075(.din(n6085), .dout(n6268));
  jor  g06076(.dina(n6093), .dinb(n6268), .dout(n6269));
  jnot g06077(.din(n6077), .dout(n6270));
  jand g06078(.dina(n6093), .dinb(n6268), .dout(n6271));
  jor  g06079(.dina(n6271), .dinb(n6270), .dout(n6272));
  jand g06080(.dina(n6272), .dinb(n6269), .dout(n6273));
  jxor g06081(.dina(n6273), .dinb(n6267), .dout(n6274));
  jand g06082(.dina(n6095), .dinb(n6068), .dout(n6275));
  jand g06083(.dina(n6114), .dinb(n6096), .dout(n6276));
  jor  g06084(.dina(n6276), .dinb(n6275), .dout(n6277));
  jxor g06085(.dina(n6277), .dinb(n6274), .dout(n6278));
  jand g06086(.dina(n6046), .dinb(n6044), .dout(n6279));
  jor  g06087(.dina(n6279), .dinb(n6048), .dout(n6280));
  jand g06088(.dina(n6080), .dinb(n6078), .dout(n6281));
  jor  g06089(.dina(n6281), .dinb(n6083), .dout(n6282));
  jxor g06090(.dina(n6282), .dinb(n6280), .dout(n6283));
  jand g06091(.dina(n6063), .dinb(n6062), .dout(n6284));
  jnot g06092(.din(n6284), .dout(n6285));
  jnot g06093(.din(n6062), .dout(n6286));
  jnot g06094(.din(n6063), .dout(n6287));
  jand g06095(.dina(n6287), .dinb(n6286), .dout(n6288));
  jor  g06096(.dina(n6288), .dinb(n6061), .dout(n6289));
  jand g06097(.dina(n6289), .dinb(n6285), .dout(n6290));
  jnot g06098(.din(n6290), .dout(n6291));
  jxor g06099(.dina(n6291), .dinb(n6283), .dout(n6292));
  jand g06100(.dina(n6092), .dinb(n6086), .dout(n6293));
  jor  g06101(.dina(n6293), .dinb(n6090), .dout(n6294));
  jnot g06102(.din(n6294), .dout(n6295));
  jand g06103(.dina(n6110), .dinb(n5890), .dout(n6296));
  jnot g06104(.din(n6296), .dout(n6297));
  jnot g06105(.din(n5890), .dout(n6298));
  jnot g06106(.din(n6110), .dout(n6299));
  jand g06107(.dina(n6299), .dinb(n6298), .dout(n6300));
  jor  g06108(.dina(n6300), .dinb(n6109), .dout(n6301));
  jand g06109(.dina(n6301), .dinb(n6297), .dout(n6302));
  jxor g06110(.dina(n6302), .dinb(n6295), .dout(n6303));
  jand g06111(.dina(n6103), .dinb(n5846), .dout(n6304));
  jor  g06112(.dina(n6304), .dinb(n6101), .dout(n6305));
  jxor g06113(.dina(n6305), .dinb(n6303), .dout(n6306));
  jxor g06114(.dina(n6306), .dinb(n6292), .dout(n6307));
  jnot g06115(.din(n6307), .dout(n6308));
  jnot g06116(.din(n6059), .dout(n6309));
  jand g06117(.dina(n6066), .dinb(n6309), .dout(n6310));
  jnot g06118(.din(n6310), .dout(n6311));
  jand g06119(.dina(n6065), .dinb(n6059), .dout(n6312));
  jor  g06120(.dina(n6312), .dinb(n6051), .dout(n6313));
  jand g06121(.dina(n6313), .dinb(n6311), .dout(n6314));
  jxor g06122(.dina(n6314), .dinb(n6308), .dout(n6315));
  jxor g06123(.dina(n6315), .dinb(n6278), .dout(n6316));
  jxor g06124(.dina(n6316), .dinb(n6256), .dout(n6317));
  jand g06125(.dina(n6181), .dinb(n6175), .dout(n6318));
  jnot g06126(.din(n6318), .dout(n6319));
  jor  g06127(.dina(n6190), .dinb(n6183), .dout(n6320));
  jand g06128(.dina(n6320), .dinb(n6319), .dout(n6321));
  jnot g06129(.din(n6321), .dout(n6322));
  jand g06130(.dina(\a[42] ), .dinb(\a[15] ), .dout(n6323));
  jand g06131(.dina(\a[48] ), .dinb(\a[9] ), .dout(n6324));
  jand g06132(.dina(\a[47] ), .dinb(\a[10] ), .dout(n6325));
  jor  g06133(.dina(n6325), .dinb(n6324), .dout(n6326));
  jnot g06134(.din(n6326), .dout(n6327));
  jand g06135(.dina(\a[48] ), .dinb(\a[10] ), .dout(n6328));
  jand g06136(.dina(n6328), .dinb(n6069), .dout(n6329));
  jor  g06137(.dina(n6329), .dinb(n6327), .dout(n6330));
  jxor g06138(.dina(n6330), .dinb(n6323), .dout(n6331));
  jand g06139(.dina(\a[52] ), .dinb(\a[5] ), .dout(n6332));
  jand g06140(.dina(\a[38] ), .dinb(\a[19] ), .dout(n6333));
  jand g06141(.dina(\a[37] ), .dinb(\a[20] ), .dout(n6334));
  jor  g06142(.dina(n6334), .dinb(n6333), .dout(n6335));
  jnot g06143(.din(n6335), .dout(n6336));
  jand g06144(.dina(\a[38] ), .dinb(\a[20] ), .dout(n6337));
  jand g06145(.dina(n6337), .dinb(n5890), .dout(n6338));
  jor  g06146(.dina(n6338), .dinb(n6336), .dout(n6339));
  jxor g06147(.dina(n6339), .dinb(n6332), .dout(n6340));
  jand g06148(.dina(\a[54] ), .dinb(\a[3] ), .dout(n6341));
  jand g06149(.dina(\a[55] ), .dinb(\a[2] ), .dout(n6342));
  jor  g06150(.dina(n6342), .dinb(n5978), .dout(n6343));
  jand g06151(.dina(\a[55] ), .dinb(\a[4] ), .dout(n6344));
  jand g06152(.dina(n6344), .dinb(n5972), .dout(n6345));
  jnot g06153(.din(n6345), .dout(n6346));
  jand g06154(.dina(n6346), .dinb(n6343), .dout(n6347));
  jxor g06155(.dina(n6347), .dinb(n6341), .dout(n6348));
  jxor g06156(.dina(n6348), .dinb(n6340), .dout(n6349));
  jxor g06157(.dina(n6349), .dinb(n6331), .dout(n6350));
  jand g06158(.dina(\a[39] ), .dinb(\a[18] ), .dout(n6351));
  jand g06159(.dina(\a[51] ), .dinb(\a[6] ), .dout(n6352));
  jand g06160(.dina(\a[40] ), .dinb(\a[17] ), .dout(n6353));
  jor  g06161(.dina(n6353), .dinb(n6352), .dout(n6354));
  jnot g06162(.din(n6354), .dout(n6355));
  jand g06163(.dina(\a[51] ), .dinb(\a[17] ), .dout(n6356));
  jand g06164(.dina(n6356), .dinb(n4120), .dout(n6357));
  jor  g06165(.dina(n6357), .dinb(n6355), .dout(n6358));
  jxor g06166(.dina(n6358), .dinb(n6351), .dout(n6359));
  jand g06167(.dina(\a[45] ), .dinb(\a[12] ), .dout(n6360));
  jand g06168(.dina(\a[29] ), .dinb(\a[28] ), .dout(n6361));
  jand g06169(.dina(\a[30] ), .dinb(\a[27] ), .dout(n6362));
  jor  g06170(.dina(n6362), .dinb(n6361), .dout(n6363));
  jnot g06171(.din(n6363), .dout(n6364));
  jand g06172(.dina(\a[30] ), .dinb(\a[28] ), .dout(n6365));
  jand g06173(.dina(n6365), .dinb(n6129), .dout(n6366));
  jor  g06174(.dina(n6366), .dinb(n6364), .dout(n6367));
  jxor g06175(.dina(n6367), .dinb(n6360), .dout(n6368));
  jand g06176(.dina(\a[46] ), .dinb(\a[11] ), .dout(n6369));
  jor  g06177(.dina(n6369), .dinb(n5945), .dout(n6370));
  jand g06178(.dina(\a[46] ), .dinb(\a[13] ), .dout(n6371));
  jand g06179(.dina(n6371), .dinb(n5943), .dout(n6372));
  jnot g06180(.din(n6372), .dout(n6373));
  jand g06181(.dina(n6373), .dinb(n6370), .dout(n6374));
  jxor g06182(.dina(n6374), .dinb(n4691), .dout(n6375));
  jxor g06183(.dina(n6375), .dinb(n6368), .dout(n6376));
  jxor g06184(.dina(n6376), .dinb(n6359), .dout(n6377));
  jxor g06185(.dina(n6377), .dinb(n6350), .dout(n6378));
  jxor g06186(.dina(n6378), .dinb(n6322), .dout(n6379));
  jor  g06187(.dina(n6222), .dinb(n6218), .dout(n6380));
  jand g06188(.dina(n6229), .dinb(n6223), .dout(n6381));
  jnot g06189(.din(n6381), .dout(n6382));
  jand g06190(.dina(n6382), .dinb(n6380), .dout(n6383));
  jnot g06191(.din(n6383), .dout(n6384));
  jand g06192(.dina(n6072), .dinb(n6069), .dout(n6385));
  jor  g06193(.dina(n6385), .dinb(n6075), .dout(n6386));
  jand g06194(.dina(n6210), .dinb(n6207), .dout(n6387));
  jor  g06195(.dina(n6387), .dinb(n6213), .dout(n6388));
  jxor g06196(.dina(n6388), .dinb(n6386), .dout(n6389));
  jand g06197(.dina(n6055), .dinb(n6052), .dout(n6390));
  jor  g06198(.dina(n6390), .dinb(n6056), .dout(n6391));
  jxor g06199(.dina(n6391), .dinb(n6389), .dout(n6392));
  jnot g06200(.din(n6392), .dout(n6393));
  jor  g06201(.dina(n6215), .dinb(n6206), .dout(n6394));
  jand g06202(.dina(n6216), .dinb(n6203), .dout(n6395));
  jnot g06203(.din(n6395), .dout(n6396));
  jand g06204(.dina(n6396), .dinb(n6394), .dout(n6397));
  jxor g06205(.dina(n6397), .dinb(n6393), .dout(n6398));
  jand g06206(.dina(\a[33] ), .dinb(\a[24] ), .dout(n6399));
  jand g06207(.dina(\a[32] ), .dinb(\a[25] ), .dout(n6400));
  jor  g06208(.dina(n6400), .dinb(n6082), .dout(n6401));
  jnot g06209(.din(n6401), .dout(n6402));
  jand g06210(.dina(\a[32] ), .dinb(\a[26] ), .dout(n6403));
  jand g06211(.dina(n6403), .dinb(n5957), .dout(n6404));
  jor  g06212(.dina(n6404), .dinb(n6402), .dout(n6405));
  jxor g06213(.dina(n6405), .dinb(n6399), .dout(n6406));
  jand g06214(.dina(\a[36] ), .dinb(\a[21] ), .dout(n6407));
  jand g06215(.dina(\a[35] ), .dinb(\a[22] ), .dout(n6408));
  jor  g06216(.dina(n6408), .dinb(n6089), .dout(n6409));
  jnot g06217(.din(n6409), .dout(n6410));
  jand g06218(.dina(\a[35] ), .dinb(\a[23] ), .dout(n6411));
  jand g06219(.dina(n6411), .dinb(n5966), .dout(n6412));
  jor  g06220(.dina(n6412), .dinb(n6410), .dout(n6413));
  jxor g06221(.dina(n6413), .dinb(n6407), .dout(n6414));
  jand g06222(.dina(\a[50] ), .dinb(\a[7] ), .dout(n6415));
  jand g06223(.dina(\a[49] ), .dinb(\a[8] ), .dout(n6416));
  jand g06224(.dina(\a[41] ), .dinb(\a[16] ), .dout(n6417));
  jor  g06225(.dina(n6417), .dinb(n6416), .dout(n6418));
  jand g06226(.dina(\a[49] ), .dinb(\a[16] ), .dout(n6419));
  jand g06227(.dina(n6419), .dinb(n4704), .dout(n6420));
  jnot g06228(.din(n6420), .dout(n6421));
  jand g06229(.dina(n6421), .dinb(n6418), .dout(n6422));
  jxor g06230(.dina(n6422), .dinb(n6415), .dout(n6423));
  jxor g06231(.dina(n6423), .dinb(n6414), .dout(n6424));
  jxor g06232(.dina(n6424), .dinb(n6406), .dout(n6425));
  jxor g06233(.dina(n6425), .dinb(n6398), .dout(n6426));
  jxor g06234(.dina(n6426), .dinb(n6384), .dout(n6427));
  jxor g06235(.dina(n6427), .dinb(n6379), .dout(n6428));
  jxor g06236(.dina(n6428), .dinb(n6317), .dout(n6429));
  jand g06237(.dina(n6196), .dinb(n6150), .dout(n6430));
  jand g06238(.dina(n6197), .dinb(n6147), .dout(n6431));
  jor  g06239(.dina(n6431), .dinb(n6430), .dout(n6432));
  jand g06240(.dina(n6145), .dinb(n6118), .dout(n6433));
  jand g06241(.dina(n6146), .dinb(n6115), .dout(n6434));
  jor  g06242(.dina(n6434), .dinb(n6433), .dout(n6435));
  jand g06243(.dina(n6194), .dinb(n6191), .dout(n6436));
  jand g06244(.dina(n6195), .dinb(n6172), .dout(n6437));
  jor  g06245(.dina(n6437), .dinb(n6436), .dout(n6438));
  jand g06246(.dina(n6167), .dinb(n6164), .dout(n6439));
  jand g06247(.dina(n6171), .dinb(n6168), .dout(n6440));
  jor  g06248(.dina(n6440), .dinb(n6439), .dout(n6441));
  jand g06249(.dina(n6143), .dinb(n6139), .dout(n6442));
  jand g06250(.dina(n6144), .dinb(n6126), .dout(n6443));
  jor  g06251(.dina(n6443), .dinb(n6442), .dout(n6444));
  jxor g06252(.dina(n6444), .dinb(n6441), .dout(n6445));
  jand g06253(.dina(n6130), .dinb(n6129), .dout(n6446));
  jand g06254(.dina(\a[57] ), .dinb(\a[0] ), .dout(n6447));
  jxor g06255(.dina(n6447), .dinb(n6446), .dout(n6448));
  jand g06256(.dina(\a[56] ), .dinb(\a[1] ), .dout(n6449));
  jxor g06257(.dina(n6449), .dinb(\a[29] ), .dout(n6450));
  jnot g06258(.din(n6450), .dout(n6451));
  jxor g06259(.dina(n6451), .dinb(n6448), .dout(n6452));
  jnot g06260(.din(n6452), .dout(n6453));
  jand g06261(.dina(n6124), .dinb(n6122), .dout(n6454));
  jand g06262(.dina(n6125), .dinb(n6120), .dout(n6455));
  jor  g06263(.dina(n6455), .dinb(n6454), .dout(n6456));
  jxor g06264(.dina(n6456), .dinb(n6453), .dout(n6457));
  jnot g06265(.din(n6457), .dout(n6458));
  jand g06266(.dina(n6154), .dinb(n6152), .dout(n6459));
  jnot g06267(.din(n6459), .dout(n6460));
  jor  g06268(.dina(n6163), .dinb(n6156), .dout(n6461));
  jand g06269(.dina(n6461), .dinb(n6460), .dout(n6462));
  jxor g06270(.dina(n6462), .dinb(n6458), .dout(n6463));
  jxor g06271(.dina(n6463), .dinb(n6445), .dout(n6464));
  jxor g06272(.dina(n6464), .dinb(n6438), .dout(n6465));
  jxor g06273(.dina(n6465), .dinb(n6435), .dout(n6466));
  jxor g06274(.dina(n6466), .dinb(n6432), .dout(n6467));
  jxor g06275(.dina(n6467), .dinb(n6429), .dout(n6468));
  jxor g06276(.dina(n6468), .dinb(n6253), .dout(n6469));
  jand g06277(.dina(n6244), .dinb(n6043), .dout(n6470));
  jor  g06278(.dina(n6244), .dinb(n6043), .dout(n6471));
  jand g06279(.dina(n6249), .dinb(n6471), .dout(n6472));
  jor  g06280(.dina(n6472), .dinb(n6470), .dout(n6473));
  jxor g06281(.dina(n6473), .dinb(n6469), .dout(\asquared[58] ));
  jand g06282(.dina(n6466), .dinb(n6432), .dout(n6475));
  jand g06283(.dina(n6467), .dinb(n6429), .dout(n6476));
  jor  g06284(.dina(n6476), .dinb(n6475), .dout(n6477));
  jand g06285(.dina(n6316), .dinb(n6256), .dout(n6478));
  jand g06286(.dina(n6428), .dinb(n6317), .dout(n6479));
  jor  g06287(.dina(n6479), .dinb(n6478), .dout(n6480));
  jand g06288(.dina(n6277), .dinb(n6274), .dout(n6481));
  jand g06289(.dina(n6315), .dinb(n6278), .dout(n6482));
  jor  g06290(.dina(n6482), .dinb(n6481), .dout(n6483));
  jor  g06291(.dina(n6397), .dinb(n6393), .dout(n6484));
  jand g06292(.dina(n6425), .dinb(n6398), .dout(n6485));
  jnot g06293(.din(n6485), .dout(n6486));
  jand g06294(.dina(n6486), .dinb(n6484), .dout(n6487));
  jnot g06295(.din(n6487), .dout(n6488));
  jand g06296(.dina(n6388), .dinb(n6386), .dout(n6489));
  jand g06297(.dina(n6391), .dinb(n6389), .dout(n6490));
  jor  g06298(.dina(n6490), .dinb(n6489), .dout(n6491));
  jnot g06299(.din(n6491), .dout(n6492));
  jor  g06300(.dina(n6302), .dinb(n6295), .dout(n6493));
  jand g06301(.dina(n6305), .dinb(n6303), .dout(n6494));
  jnot g06302(.din(n6494), .dout(n6495));
  jand g06303(.dina(n6495), .dinb(n6493), .dout(n6496));
  jxor g06304(.dina(n6496), .dinb(n6492), .dout(n6497));
  jand g06305(.dina(n6282), .dinb(n6280), .dout(n6498));
  jand g06306(.dina(n6291), .dinb(n6283), .dout(n6499));
  jor  g06307(.dina(n6499), .dinb(n6498), .dout(n6500));
  jxor g06308(.dina(n6500), .dinb(n6497), .dout(n6501));
  jnot g06309(.din(n6501), .dout(n6502));
  jand g06310(.dina(n6306), .dinb(n6292), .dout(n6503));
  jnot g06311(.din(n6503), .dout(n6504));
  jor  g06312(.dina(n6314), .dinb(n6308), .dout(n6505));
  jand g06313(.dina(n6505), .dinb(n6504), .dout(n6506));
  jxor g06314(.dina(n6506), .dinb(n6502), .dout(n6507));
  jxor g06315(.dina(n6507), .dinb(n6488), .dout(n6508));
  jxor g06316(.dina(n6508), .dinb(n6483), .dout(n6509));
  jand g06317(.dina(n6426), .dinb(n6384), .dout(n6510));
  jand g06318(.dina(n6427), .dinb(n6379), .dout(n6511));
  jor  g06319(.dina(n6511), .dinb(n6510), .dout(n6512));
  jxor g06320(.dina(n6512), .dinb(n6509), .dout(n6513));
  jxor g06321(.dina(n6513), .dinb(n6480), .dout(n6514));
  jand g06322(.dina(n6464), .dinb(n6438), .dout(n6515));
  jand g06323(.dina(n6465), .dinb(n6435), .dout(n6516));
  jor  g06324(.dina(n6516), .dinb(n6515), .dout(n6517));
  jand g06325(.dina(n6377), .dinb(n6350), .dout(n6518));
  jand g06326(.dina(n6378), .dinb(n6322), .dout(n6519));
  jor  g06327(.dina(n6519), .dinb(n6518), .dout(n6520));
  jand g06328(.dina(n6449), .dinb(\a[29] ), .dout(n6521));
  jand g06329(.dina(\a[57] ), .dinb(\a[1] ), .dout(n6522));
  jxor g06330(.dina(n6522), .dinb(n6365), .dout(n6523));
  jxor g06331(.dina(n6523), .dinb(n6521), .dout(n6524));
  jand g06332(.dina(n6363), .dinb(n6360), .dout(n6525));
  jor  g06333(.dina(n6525), .dinb(n6366), .dout(n6526));
  jxor g06334(.dina(n6526), .dinb(n6524), .dout(n6527));
  jnot g06335(.din(n6340), .dout(n6528));
  jor  g06336(.dina(n6348), .dinb(n6528), .dout(n6529));
  jnot g06337(.din(n6331), .dout(n6530));
  jand g06338(.dina(n6348), .dinb(n6528), .dout(n6531));
  jor  g06339(.dina(n6531), .dinb(n6530), .dout(n6532));
  jand g06340(.dina(n6532), .dinb(n6529), .dout(n6533));
  jxor g06341(.dina(n6533), .dinb(n6527), .dout(n6534));
  jnot g06342(.din(n6368), .dout(n6535));
  jor  g06343(.dina(n6375), .dinb(n6535), .dout(n6536));
  jnot g06344(.din(n6359), .dout(n6537));
  jand g06345(.dina(n6375), .dinb(n6535), .dout(n6538));
  jor  g06346(.dina(n6538), .dinb(n6537), .dout(n6539));
  jand g06347(.dina(n6539), .dinb(n6536), .dout(n6540));
  jxor g06348(.dina(n6540), .dinb(n6534), .dout(n6541));
  jxor g06349(.dina(n6541), .dinb(n6520), .dout(n6542));
  jand g06350(.dina(n6326), .dinb(n6323), .dout(n6543));
  jor  g06351(.dina(n6543), .dinb(n6329), .dout(n6544));
  jand g06352(.dina(n6401), .dinb(n6399), .dout(n6545));
  jor  g06353(.dina(n6545), .dinb(n6404), .dout(n6546));
  jxor g06354(.dina(n6546), .dinb(n6544), .dout(n6547));
  jand g06355(.dina(n6409), .dinb(n6407), .dout(n6548));
  jor  g06356(.dina(n6548), .dinb(n6412), .dout(n6549));
  jxor g06357(.dina(n6549), .dinb(n6547), .dout(n6550));
  jand g06358(.dina(n6374), .dinb(n4691), .dout(n6551));
  jor  g06359(.dina(n6551), .dinb(n6372), .dout(n6552));
  jand g06360(.dina(n6347), .dinb(n6341), .dout(n6553));
  jor  g06361(.dina(n6553), .dinb(n6345), .dout(n6554));
  jand g06362(.dina(n6335), .dinb(n6332), .dout(n6555));
  jor  g06363(.dina(n6555), .dinb(n6338), .dout(n6556));
  jxor g06364(.dina(n6556), .dinb(n6554), .dout(n6557));
  jxor g06365(.dina(n6557), .dinb(n6552), .dout(n6558));
  jxor g06366(.dina(n6558), .dinb(n6550), .dout(n6559));
  jnot g06367(.din(n6414), .dout(n6560));
  jor  g06368(.dina(n6423), .dinb(n6560), .dout(n6561));
  jnot g06369(.din(n6406), .dout(n6562));
  jand g06370(.dina(n6423), .dinb(n6560), .dout(n6563));
  jor  g06371(.dina(n6563), .dinb(n6562), .dout(n6564));
  jand g06372(.dina(n6564), .dinb(n6561), .dout(n6565));
  jxor g06373(.dina(n6565), .dinb(n6559), .dout(n6566));
  jxor g06374(.dina(n6566), .dinb(n6542), .dout(n6567));
  jxor g06375(.dina(n6567), .dinb(n6517), .dout(n6568));
  jand g06376(.dina(n6266), .dinb(n6259), .dout(n6569));
  jand g06377(.dina(n6273), .dinb(n6267), .dout(n6570));
  jor  g06378(.dina(n6570), .dinb(n6569), .dout(n6571));
  jand g06379(.dina(\a[41] ), .dinb(\a[17] ), .dout(n6572));
  jnot g06380(.din(n6572), .dout(n6573));
  jand g06381(.dina(\a[49] ), .dinb(\a[9] ), .dout(n6574));
  jand g06382(.dina(\a[42] ), .dinb(\a[16] ), .dout(n6575));
  jor  g06383(.dina(n6575), .dinb(n6574), .dout(n6576));
  jand g06384(.dina(n6419), .dinb(n5063), .dout(n6577));
  jnot g06385(.din(n6577), .dout(n6578));
  jand g06386(.dina(n6578), .dinb(n6576), .dout(n6579));
  jxor g06387(.dina(n6579), .dinb(n6573), .dout(n6580));
  jand g06388(.dina(\a[53] ), .dinb(\a[5] ), .dout(n6581));
  jnot g06389(.din(n6581), .dout(n6582));
  jand g06390(.dina(\a[37] ), .dinb(\a[21] ), .dout(n6583));
  jor  g06391(.dina(n6583), .dinb(n6337), .dout(n6584));
  jand g06392(.dina(\a[38] ), .dinb(\a[21] ), .dout(n6585));
  jand g06393(.dina(n6585), .dinb(n6334), .dout(n6586));
  jnot g06394(.din(n6586), .dout(n6587));
  jand g06395(.dina(n6587), .dinb(n6584), .dout(n6588));
  jxor g06396(.dina(n6588), .dinb(n6582), .dout(n6589));
  jnot g06397(.din(n6100), .dout(n6590));
  jand g06398(.dina(\a[58] ), .dinb(\a[0] ), .dout(n6591));
  jand g06399(.dina(\a[54] ), .dinb(\a[4] ), .dout(n6592));
  jxor g06400(.dina(n6592), .dinb(n6591), .dout(n6593));
  jxor g06401(.dina(n6593), .dinb(n6590), .dout(n6594));
  jnot g06402(.din(n6594), .dout(n6595));
  jxor g06403(.dina(n6595), .dinb(n6589), .dout(n6596));
  jxor g06404(.dina(n6596), .dinb(n6580), .dout(n6597));
  jand g06405(.dina(\a[33] ), .dinb(\a[25] ), .dout(n6598));
  jand g06406(.dina(\a[31] ), .dinb(\a[27] ), .dout(n6599));
  jor  g06407(.dina(n6599), .dinb(n6403), .dout(n6600));
  jnot g06408(.din(n6600), .dout(n6601));
  jand g06409(.dina(\a[32] ), .dinb(\a[27] ), .dout(n6602));
  jand g06410(.dina(n6602), .dinb(n6082), .dout(n6603));
  jor  g06411(.dina(n6603), .dinb(n6601), .dout(n6604));
  jxor g06412(.dina(n6604), .dinb(n6598), .dout(n6605));
  jand g06413(.dina(\a[36] ), .dinb(\a[22] ), .dout(n6606));
  jand g06414(.dina(\a[34] ), .dinb(\a[24] ), .dout(n6607));
  jor  g06415(.dina(n6607), .dinb(n6411), .dout(n6608));
  jnot g06416(.din(n6608), .dout(n6609));
  jand g06417(.dina(\a[35] ), .dinb(\a[24] ), .dout(n6610));
  jand g06418(.dina(n6610), .dinb(n6089), .dout(n6611));
  jor  g06419(.dina(n6611), .dinb(n6609), .dout(n6612));
  jxor g06420(.dina(n6612), .dinb(n6606), .dout(n6613));
  jand g06421(.dina(\a[40] ), .dinb(\a[18] ), .dout(n6614));
  jand g06422(.dina(\a[51] ), .dinb(\a[7] ), .dout(n6615));
  jand g06423(.dina(\a[50] ), .dinb(\a[8] ), .dout(n6616));
  jor  g06424(.dina(n6616), .dinb(n6615), .dout(n6617));
  jand g06425(.dina(\a[51] ), .dinb(\a[8] ), .dout(n6618));
  jand g06426(.dina(n6618), .dinb(n6415), .dout(n6619));
  jnot g06427(.din(n6619), .dout(n6620));
  jand g06428(.dina(n6620), .dinb(n6617), .dout(n6621));
  jxor g06429(.dina(n6621), .dinb(n6614), .dout(n6622));
  jxor g06430(.dina(n6622), .dinb(n6613), .dout(n6623));
  jxor g06431(.dina(n6623), .dinb(n6605), .dout(n6624));
  jxor g06432(.dina(n6624), .dinb(n6597), .dout(n6625));
  jxor g06433(.dina(n6625), .dinb(n6571), .dout(n6626));
  jand g06434(.dina(n6444), .dinb(n6441), .dout(n6627));
  jand g06435(.dina(n6463), .dinb(n6445), .dout(n6628));
  jor  g06436(.dina(n6628), .dinb(n6627), .dout(n6629));
  jand g06437(.dina(n6422), .dinb(n6415), .dout(n6630));
  jor  g06438(.dina(n6630), .dinb(n6420), .dout(n6631));
  jand g06439(.dina(n6354), .dinb(n6351), .dout(n6632));
  jor  g06440(.dina(n6632), .dinb(n6357), .dout(n6633));
  jxor g06441(.dina(n6633), .dinb(n6631), .dout(n6634));
  jor  g06442(.dina(n6447), .dinb(n6446), .dout(n6635));
  jand g06443(.dina(n6447), .dinb(n6446), .dout(n6636));
  jor  g06444(.dina(n6450), .dinb(n6636), .dout(n6637));
  jand g06445(.dina(n6637), .dinb(n6635), .dout(n6638));
  jxor g06446(.dina(n6638), .dinb(n6634), .dout(n6639));
  jnot g06447(.din(n6639), .dout(n6640));
  jand g06448(.dina(n6456), .dinb(n6453), .dout(n6641));
  jnot g06449(.din(n6641), .dout(n6642));
  jor  g06450(.dina(n6462), .dinb(n6458), .dout(n6643));
  jand g06451(.dina(n6643), .dinb(n6642), .dout(n6644));
  jxor g06452(.dina(n6644), .dinb(n6640), .dout(n6645));
  jand g06453(.dina(\a[45] ), .dinb(\a[13] ), .dout(n6646));
  jand g06454(.dina(\a[46] ), .dinb(\a[12] ), .dout(n6647));
  jor  g06455(.dina(n6647), .dinb(n6646), .dout(n6648));
  jnot g06456(.din(n6648), .dout(n6649));
  jand g06457(.dina(n6371), .dinb(n6360), .dout(n6650));
  jor  g06458(.dina(n6650), .dinb(n6649), .dout(n6651));
  jxor g06459(.dina(n6651), .dinb(n5473), .dout(n6652));
  jnot g06460(.din(n6652), .dout(n6653));
  jand g06461(.dina(\a[47] ), .dinb(\a[11] ), .dout(n6654));
  jor  g06462(.dina(n6654), .dinb(n4377), .dout(n6655));
  jand g06463(.dina(\a[47] ), .dinb(\a[15] ), .dout(n6656));
  jand g06464(.dina(n6656), .dinb(n5734), .dout(n6657));
  jnot g06465(.din(n6657), .dout(n6658));
  jand g06466(.dina(n6658), .dinb(n6655), .dout(n6659));
  jxor g06467(.dina(n6659), .dinb(n6328), .dout(n6660));
  jxor g06468(.dina(n6660), .dinb(n6653), .dout(n6661));
  jand g06469(.dina(\a[55] ), .dinb(\a[3] ), .dout(n6662));
  jand g06470(.dina(\a[39] ), .dinb(\a[19] ), .dout(n6663));
  jnot g06471(.din(n6663), .dout(n6664));
  jand g06472(.dina(\a[52] ), .dinb(\a[6] ), .dout(n6665));
  jxor g06473(.dina(n6665), .dinb(n6664), .dout(n6666));
  jxor g06474(.dina(n6666), .dinb(n6662), .dout(n6667));
  jnot g06475(.din(n6667), .dout(n6668));
  jxor g06476(.dina(n6668), .dinb(n6661), .dout(n6669));
  jxor g06477(.dina(n6669), .dinb(n6645), .dout(n6670));
  jxor g06478(.dina(n6670), .dinb(n6629), .dout(n6671));
  jxor g06479(.dina(n6671), .dinb(n6626), .dout(n6672));
  jxor g06480(.dina(n6672), .dinb(n6568), .dout(n6673));
  jxor g06481(.dina(n6673), .dinb(n6514), .dout(n6674));
  jxor g06482(.dina(n6674), .dinb(n6477), .dout(n6675));
  jand g06483(.dina(n6468), .dinb(n6253), .dout(n6676));
  jor  g06484(.dina(n6468), .dinb(n6253), .dout(n6677));
  jand g06485(.dina(n6473), .dinb(n6677), .dout(n6678));
  jor  g06486(.dina(n6678), .dinb(n6676), .dout(n6679));
  jxor g06487(.dina(n6679), .dinb(n6675), .dout(\asquared[59] ));
  jand g06488(.dina(n6567), .dinb(n6517), .dout(n6681));
  jand g06489(.dina(n6672), .dinb(n6568), .dout(n6682));
  jor  g06490(.dina(n6682), .dinb(n6681), .dout(n6683));
  jand g06491(.dina(n6670), .dinb(n6629), .dout(n6684));
  jand g06492(.dina(n6671), .dinb(n6626), .dout(n6685));
  jor  g06493(.dina(n6685), .dinb(n6684), .dout(n6686));
  jand g06494(.dina(n6541), .dinb(n6520), .dout(n6687));
  jand g06495(.dina(n6566), .dinb(n6542), .dout(n6688));
  jor  g06496(.dina(n6688), .dinb(n6687), .dout(n6689));
  jor  g06497(.dina(n6644), .dinb(n6640), .dout(n6690));
  jand g06498(.dina(n6669), .dinb(n6645), .dout(n6691));
  jnot g06499(.din(n6691), .dout(n6692));
  jand g06500(.dina(n6692), .dinb(n6690), .dout(n6693));
  jnot g06501(.din(n6693), .dout(n6694));
  jand g06502(.dina(n6633), .dinb(n6631), .dout(n6695));
  jand g06503(.dina(n6638), .dinb(n6634), .dout(n6696));
  jor  g06504(.dina(n6696), .dinb(n6695), .dout(n6697));
  jand g06505(.dina(n6556), .dinb(n6554), .dout(n6698));
  jand g06506(.dina(n6557), .dinb(n6552), .dout(n6699));
  jor  g06507(.dina(n6699), .dinb(n6698), .dout(n6700));
  jxor g06508(.dina(n6700), .dinb(n6697), .dout(n6701));
  jand g06509(.dina(n6546), .dinb(n6544), .dout(n6702));
  jand g06510(.dina(n6549), .dinb(n6547), .dout(n6703));
  jor  g06511(.dina(n6703), .dinb(n6702), .dout(n6704));
  jxor g06512(.dina(n6704), .dinb(n6701), .dout(n6705));
  jand g06513(.dina(n6558), .dinb(n6550), .dout(n6706));
  jand g06514(.dina(n6565), .dinb(n6559), .dout(n6707));
  jor  g06515(.dina(n6707), .dinb(n6706), .dout(n6708));
  jxor g06516(.dina(n6708), .dinb(n6705), .dout(n6709));
  jxor g06517(.dina(n6709), .dinb(n6694), .dout(n6710));
  jxor g06518(.dina(n6710), .dinb(n6689), .dout(n6711));
  jxor g06519(.dina(n6711), .dinb(n6686), .dout(n6712));
  jxor g06520(.dina(n6712), .dinb(n6683), .dout(n6713));
  jand g06521(.dina(n6508), .dinb(n6483), .dout(n6714));
  jand g06522(.dina(n6512), .dinb(n6509), .dout(n6715));
  jor  g06523(.dina(n6715), .dinb(n6714), .dout(n6716));
  jor  g06524(.dina(n6660), .dinb(n6653), .dout(n6717));
  jand g06525(.dina(n6660), .dinb(n6653), .dout(n6718));
  jor  g06526(.dina(n6668), .dinb(n6718), .dout(n6719));
  jand g06527(.dina(n6719), .dinb(n6717), .dout(n6720));
  jnot g06528(.din(n6613), .dout(n6721));
  jor  g06529(.dina(n6622), .dinb(n6721), .dout(n6722));
  jnot g06530(.din(n6605), .dout(n6723));
  jand g06531(.dina(n6622), .dinb(n6721), .dout(n6724));
  jor  g06532(.dina(n6724), .dinb(n6723), .dout(n6725));
  jand g06533(.dina(n6725), .dinb(n6722), .dout(n6726));
  jxor g06534(.dina(n6726), .dinb(n6720), .dout(n6727));
  jnot g06535(.din(n6727), .dout(n6728));
  jnot g06536(.din(n6589), .dout(n6729));
  jand g06537(.dina(n6595), .dinb(n6729), .dout(n6730));
  jnot g06538(.din(n6730), .dout(n6731));
  jand g06539(.dina(n6594), .dinb(n6589), .dout(n6732));
  jor  g06540(.dina(n6732), .dinb(n6580), .dout(n6733));
  jand g06541(.dina(n6733), .dinb(n6731), .dout(n6734));
  jxor g06542(.dina(n6734), .dinb(n6728), .dout(n6735));
  jand g06543(.dina(n6624), .dinb(n6597), .dout(n6736));
  jand g06544(.dina(n6625), .dinb(n6571), .dout(n6737));
  jor  g06545(.dina(n6737), .dinb(n6736), .dout(n6738));
  jand g06546(.dina(n6592), .dinb(n6591), .dout(n6739));
  jnot g06547(.din(n6739), .dout(n6740));
  jnot g06548(.din(n6591), .dout(n6741));
  jnot g06549(.din(n6592), .dout(n6742));
  jand g06550(.dina(n6742), .dinb(n6741), .dout(n6743));
  jor  g06551(.dina(n6743), .dinb(n6590), .dout(n6744));
  jand g06552(.dina(n6744), .dinb(n6740), .dout(n6745));
  jnot g06553(.din(n6745), .dout(n6746));
  jnot g06554(.din(n6665), .dout(n6747));
  jand g06555(.dina(n6747), .dinb(n6664), .dout(n6748));
  jnot g06556(.din(n6748), .dout(n6749));
  jand g06557(.dina(n6665), .dinb(n6663), .dout(n6750));
  jor  g06558(.dina(n6750), .dinb(n6662), .dout(n6751));
  jand g06559(.dina(n6751), .dinb(n6749), .dout(n6752));
  jxor g06560(.dina(n6752), .dinb(n6746), .dout(n6753));
  jand g06561(.dina(n6576), .dinb(n6572), .dout(n6754));
  jor  g06562(.dina(n6754), .dinb(n6577), .dout(n6755));
  jxor g06563(.dina(n6755), .dinb(n6753), .dout(n6756));
  jand g06564(.dina(n6621), .dinb(n6614), .dout(n6757));
  jor  g06565(.dina(n6757), .dinb(n6619), .dout(n6758));
  jand g06566(.dina(n6584), .dinb(n6581), .dout(n6759));
  jor  g06567(.dina(n6759), .dinb(n6586), .dout(n6760));
  jand g06568(.dina(n6608), .dinb(n6606), .dout(n6761));
  jor  g06569(.dina(n6761), .dinb(n6611), .dout(n6762));
  jxor g06570(.dina(n6762), .dinb(n6760), .dout(n6763));
  jxor g06571(.dina(n6763), .dinb(n6758), .dout(n6764));
  jand g06572(.dina(n6659), .dinb(n6328), .dout(n6765));
  jor  g06573(.dina(n6765), .dinb(n6657), .dout(n6766));
  jand g06574(.dina(n2016), .dinb(\a[58] ), .dout(n6767));
  jnot g06575(.din(n6767), .dout(n6768));
  jand g06576(.dina(\a[58] ), .dinb(\a[1] ), .dout(n6769));
  jor  g06577(.dina(n6769), .dinb(\a[30] ), .dout(n6770));
  jand g06578(.dina(n6770), .dinb(n6768), .dout(n6771));
  jand g06579(.dina(n6648), .dinb(n5473), .dout(n6772));
  jor  g06580(.dina(n6772), .dinb(n6650), .dout(n6773));
  jxor g06581(.dina(n6773), .dinb(n6771), .dout(n6774));
  jxor g06582(.dina(n6774), .dinb(n6766), .dout(n6775));
  jxor g06583(.dina(n6775), .dinb(n6764), .dout(n6776));
  jxor g06584(.dina(n6776), .dinb(n6756), .dout(n6777));
  jxor g06585(.dina(n6777), .dinb(n6738), .dout(n6778));
  jxor g06586(.dina(n6778), .dinb(n6735), .dout(n6779));
  jxor g06587(.dina(n6779), .dinb(n6716), .dout(n6780));
  jor  g06588(.dina(n6506), .dinb(n6502), .dout(n6781));
  jand g06589(.dina(n6507), .dinb(n6488), .dout(n6782));
  jnot g06590(.din(n6782), .dout(n6783));
  jand g06591(.dina(n6783), .dinb(n6781), .dout(n6784));
  jnot g06592(.din(n6784), .dout(n6785));
  jand g06593(.dina(n6533), .dinb(n6527), .dout(n6786));
  jand g06594(.dina(n6540), .dinb(n6534), .dout(n6787));
  jor  g06595(.dina(n6787), .dinb(n6786), .dout(n6788));
  jnot g06596(.din(n6344), .dout(n6789));
  jand g06597(.dina(\a[54] ), .dinb(\a[5] ), .dout(n6790));
  jand g06598(.dina(\a[40] ), .dinb(\a[19] ), .dout(n6791));
  jxor g06599(.dina(n6791), .dinb(n6790), .dout(n6792));
  jxor g06600(.dina(n6792), .dinb(n6789), .dout(n6793));
  jnot g06601(.din(n6793), .dout(n6794));
  jand g06602(.dina(n6600), .dinb(n6598), .dout(n6795));
  jor  g06603(.dina(n6795), .dinb(n6603), .dout(n6796));
  jnot g06604(.din(n6796), .dout(n6797));
  jand g06605(.dina(n6522), .dinb(n6365), .dout(n6798));
  jand g06606(.dina(\a[57] ), .dinb(\a[2] ), .dout(n6799));
  jand g06607(.dina(\a[56] ), .dinb(\a[3] ), .dout(n6800));
  jor  g06608(.dina(n6800), .dinb(n6799), .dout(n6801));
  jnot g06609(.din(n6801), .dout(n6802));
  jand g06610(.dina(\a[57] ), .dinb(\a[3] ), .dout(n6803));
  jand g06611(.dina(n6803), .dinb(n6100), .dout(n6804));
  jor  g06612(.dina(n6804), .dinb(n6802), .dout(n6805));
  jxor g06613(.dina(n6805), .dinb(n6798), .dout(n6806));
  jxor g06614(.dina(n6806), .dinb(n6797), .dout(n6807));
  jxor g06615(.dina(n6807), .dinb(n6794), .dout(n6808));
  jand g06616(.dina(\a[43] ), .dinb(\a[16] ), .dout(n6809));
  jand g06617(.dina(\a[42] ), .dinb(\a[17] ), .dout(n6810));
  jor  g06618(.dina(n6810), .dinb(n6809), .dout(n6811));
  jnot g06619(.din(n6811), .dout(n6812));
  jand g06620(.dina(\a[43] ), .dinb(\a[17] ), .dout(n6813));
  jand g06621(.dina(n6813), .dinb(n6575), .dout(n6814));
  jor  g06622(.dina(n6814), .dinb(n6812), .dout(n6815));
  jxor g06623(.dina(n6815), .dinb(n6618), .dout(n6816));
  jnot g06624(.din(n6816), .dout(n6817));
  jand g06625(.dina(\a[30] ), .dinb(\a[29] ), .dout(n6818));
  jnot g06626(.din(n6818), .dout(n6819));
  jand g06627(.dina(\a[31] ), .dinb(\a[28] ), .dout(n6820));
  jxor g06628(.dina(n6820), .dinb(n6819), .dout(n6821));
  jxor g06629(.dina(n6821), .dinb(n6371), .dout(n6822));
  jnot g06630(.din(n6822), .dout(n6823));
  jand g06631(.dina(\a[48] ), .dinb(\a[11] ), .dout(n6824));
  jand g06632(.dina(\a[47] ), .dinb(\a[12] ), .dout(n6825));
  jor  g06633(.dina(n6825), .dinb(n5078), .dout(n6826));
  jand g06634(.dina(\a[47] ), .dinb(\a[14] ), .dout(n6827));
  jand g06635(.dina(n6827), .dinb(n6360), .dout(n6828));
  jnot g06636(.din(n6828), .dout(n6829));
  jand g06637(.dina(n6829), .dinb(n6826), .dout(n6830));
  jxor g06638(.dina(n6830), .dinb(n6824), .dout(n6831));
  jxor g06639(.dina(n6831), .dinb(n6823), .dout(n6832));
  jxor g06640(.dina(n6832), .dinb(n6817), .dout(n6833));
  jxor g06641(.dina(n6833), .dinb(n6808), .dout(n6834));
  jxor g06642(.dina(n6834), .dinb(n6788), .dout(n6835));
  jxor g06643(.dina(n6835), .dinb(n6785), .dout(n6836));
  jand g06644(.dina(n6523), .dinb(n6521), .dout(n6837));
  jand g06645(.dina(n6526), .dinb(n6524), .dout(n6838));
  jor  g06646(.dina(n6838), .dinb(n6837), .dout(n6839));
  jand g06647(.dina(\a[50] ), .dinb(\a[9] ), .dout(n6840));
  jand g06648(.dina(\a[44] ), .dinb(\a[15] ), .dout(n6841));
  jand g06649(.dina(\a[49] ), .dinb(\a[10] ), .dout(n6842));
  jor  g06650(.dina(n6842), .dinb(n6841), .dout(n6843));
  jnot g06651(.din(n6843), .dout(n6844));
  jand g06652(.dina(\a[49] ), .dinb(\a[15] ), .dout(n6845));
  jand g06653(.dina(n6845), .dinb(n5775), .dout(n6846));
  jor  g06654(.dina(n6846), .dinb(n6844), .dout(n6847));
  jxor g06655(.dina(n6847), .dinb(n6840), .dout(n6848));
  jnot g06656(.din(n6848), .dout(n6849));
  jand g06657(.dina(\a[53] ), .dinb(\a[6] ), .dout(n6850));
  jand g06658(.dina(\a[52] ), .dinb(\a[7] ), .dout(n6851));
  jand g06659(.dina(\a[41] ), .dinb(\a[18] ), .dout(n6852));
  jor  g06660(.dina(n6852), .dinb(n6851), .dout(n6853));
  jand g06661(.dina(\a[52] ), .dinb(\a[18] ), .dout(n6854));
  jand g06662(.dina(n6854), .dinb(n4485), .dout(n6855));
  jnot g06663(.din(n6855), .dout(n6856));
  jand g06664(.dina(n6856), .dinb(n6853), .dout(n6857));
  jxor g06665(.dina(n6857), .dinb(n6850), .dout(n6858));
  jxor g06666(.dina(n6858), .dinb(n6849), .dout(n6859));
  jxor g06667(.dina(n6859), .dinb(n6839), .dout(n6860));
  jnot g06668(.din(n6860), .dout(n6861));
  jor  g06669(.dina(n6496), .dinb(n6492), .dout(n6862));
  jand g06670(.dina(n6500), .dinb(n6497), .dout(n6863));
  jnot g06671(.din(n6863), .dout(n6864));
  jand g06672(.dina(n6864), .dinb(n6862), .dout(n6865));
  jxor g06673(.dina(n6865), .dinb(n6861), .dout(n6866));
  jand g06674(.dina(\a[33] ), .dinb(\a[26] ), .dout(n6867));
  jand g06675(.dina(\a[59] ), .dinb(\a[0] ), .dout(n6868));
  jor  g06676(.dina(n6868), .dinb(n6602), .dout(n6869));
  jnot g06677(.din(n6869), .dout(n6870));
  jand g06678(.dina(\a[59] ), .dinb(\a[27] ), .dout(n6871));
  jand g06679(.dina(n6871), .dinb(n2109), .dout(n6872));
  jor  g06680(.dina(n6872), .dinb(n6870), .dout(n6873));
  jxor g06681(.dina(n6873), .dinb(n6867), .dout(n6874));
  jand g06682(.dina(\a[36] ), .dinb(\a[23] ), .dout(n6875));
  jand g06683(.dina(\a[34] ), .dinb(\a[25] ), .dout(n6876));
  jor  g06684(.dina(n6876), .dinb(n6610), .dout(n6877));
  jnot g06685(.din(n6877), .dout(n6878));
  jand g06686(.dina(\a[35] ), .dinb(\a[25] ), .dout(n6879));
  jand g06687(.dina(n6879), .dinb(n6607), .dout(n6880));
  jor  g06688(.dina(n6880), .dinb(n6878), .dout(n6881));
  jxor g06689(.dina(n6881), .dinb(n6875), .dout(n6882));
  jand g06690(.dina(\a[39] ), .dinb(\a[20] ), .dout(n6883));
  jand g06691(.dina(\a[37] ), .dinb(\a[22] ), .dout(n6884));
  jor  g06692(.dina(n6884), .dinb(n6585), .dout(n6885));
  jand g06693(.dina(\a[38] ), .dinb(\a[22] ), .dout(n6886));
  jand g06694(.dina(n6886), .dinb(n6583), .dout(n6887));
  jnot g06695(.din(n6887), .dout(n6888));
  jand g06696(.dina(n6888), .dinb(n6885), .dout(n6889));
  jxor g06697(.dina(n6889), .dinb(n6883), .dout(n6890));
  jxor g06698(.dina(n6890), .dinb(n6882), .dout(n6891));
  jxor g06699(.dina(n6891), .dinb(n6874), .dout(n6892));
  jxor g06700(.dina(n6892), .dinb(n6866), .dout(n6893));
  jxor g06701(.dina(n6893), .dinb(n6836), .dout(n6894));
  jxor g06702(.dina(n6894), .dinb(n6780), .dout(n6895));
  jxor g06703(.dina(n6895), .dinb(n6713), .dout(n6896));
  jand g06704(.dina(n6513), .dinb(n6480), .dout(n6897));
  jand g06705(.dina(n6673), .dinb(n6514), .dout(n6898));
  jor  g06706(.dina(n6898), .dinb(n6897), .dout(n6899));
  jxor g06707(.dina(n6899), .dinb(n6896), .dout(n6900));
  jand g06708(.dina(n6674), .dinb(n6477), .dout(n6901));
  jor  g06709(.dina(n6674), .dinb(n6477), .dout(n6902));
  jand g06710(.dina(n6679), .dinb(n6902), .dout(n6903));
  jor  g06711(.dina(n6903), .dinb(n6901), .dout(n6904));
  jxor g06712(.dina(n6904), .dinb(n6900), .dout(\asquared[60] ));
  jand g06713(.dina(n6712), .dinb(n6683), .dout(n6906));
  jand g06714(.dina(n6895), .dinb(n6713), .dout(n6907));
  jor  g06715(.dina(n6907), .dinb(n6906), .dout(n6908));
  jand g06716(.dina(n6779), .dinb(n6716), .dout(n6909));
  jand g06717(.dina(n6894), .dinb(n6780), .dout(n6910));
  jor  g06718(.dina(n6910), .dinb(n6909), .dout(n6911));
  jand g06719(.dina(n6835), .dinb(n6785), .dout(n6912));
  jand g06720(.dina(n6893), .dinb(n6836), .dout(n6913));
  jor  g06721(.dina(n6913), .dinb(n6912), .dout(n6914));
  jand g06722(.dina(n6777), .dinb(n6738), .dout(n6915));
  jand g06723(.dina(n6778), .dinb(n6735), .dout(n6916));
  jor  g06724(.dina(n6916), .dinb(n6915), .dout(n6917));
  jand g06725(.dina(n6762), .dinb(n6760), .dout(n6918));
  jand g06726(.dina(n6763), .dinb(n6758), .dout(n6919));
  jor  g06727(.dina(n6919), .dinb(n6918), .dout(n6920));
  jand g06728(.dina(n6752), .dinb(n6746), .dout(n6921));
  jand g06729(.dina(n6755), .dinb(n6753), .dout(n6922));
  jor  g06730(.dina(n6922), .dinb(n6921), .dout(n6923));
  jxor g06731(.dina(n6923), .dinb(n6920), .dout(n6924));
  jnot g06732(.din(n6924), .dout(n6925));
  jor  g06733(.dina(n6806), .dinb(n6797), .dout(n6926));
  jand g06734(.dina(n6807), .dinb(n6794), .dout(n6927));
  jnot g06735(.din(n6927), .dout(n6928));
  jand g06736(.dina(n6928), .dinb(n6926), .dout(n6929));
  jxor g06737(.dina(n6929), .dinb(n6925), .dout(n6930));
  jnot g06738(.din(n6930), .dout(n6931));
  jand g06739(.dina(n6726), .dinb(n6720), .dout(n6932));
  jnot g06740(.din(n6932), .dout(n6933));
  jor  g06741(.dina(n6734), .dinb(n6728), .dout(n6934));
  jand g06742(.dina(n6934), .dinb(n6933), .dout(n6935));
  jxor g06743(.dina(n6935), .dinb(n6931), .dout(n6936));
  jnot g06744(.din(n6936), .dout(n6937));
  jor  g06745(.dina(n6865), .dinb(n6861), .dout(n6938));
  jand g06746(.dina(n6892), .dinb(n6866), .dout(n6939));
  jnot g06747(.din(n6939), .dout(n6940));
  jand g06748(.dina(n6940), .dinb(n6938), .dout(n6941));
  jxor g06749(.dina(n6941), .dinb(n6937), .dout(n6942));
  jxor g06750(.dina(n6942), .dinb(n6917), .dout(n6943));
  jxor g06751(.dina(n6943), .dinb(n6914), .dout(n6944));
  jxor g06752(.dina(n6944), .dinb(n6911), .dout(n6945));
  jand g06753(.dina(n6775), .dinb(n6764), .dout(n6946));
  jand g06754(.dina(n6776), .dinb(n6756), .dout(n6947));
  jor  g06755(.dina(n6947), .dinb(n6946), .dout(n6948));
  jand g06756(.dina(n6773), .dinb(n6771), .dout(n6949));
  jand g06757(.dina(n6774), .dinb(n6766), .dout(n6950));
  jor  g06758(.dina(n6950), .dinb(n6949), .dout(n6951));
  jand g06759(.dina(\a[60] ), .dinb(\a[0] ), .dout(n6952));
  jxor g06760(.dina(n6952), .dinb(n6767), .dout(n6953));
  jand g06761(.dina(\a[31] ), .dinb(\a[29] ), .dout(n6954));
  jand g06762(.dina(\a[59] ), .dinb(\a[1] ), .dout(n6955));
  jxor g06763(.dina(n6955), .dinb(n6954), .dout(n6956));
  jnot g06764(.din(n6956), .dout(n6957));
  jxor g06765(.dina(n6957), .dinb(n6953), .dout(n6958));
  jand g06766(.dina(\a[33] ), .dinb(\a[27] ), .dout(n6959));
  jnot g06767(.din(n6959), .dout(n6960));
  jand g06768(.dina(\a[32] ), .dinb(\a[28] ), .dout(n6961));
  jand g06769(.dina(\a[37] ), .dinb(\a[23] ), .dout(n6962));
  jxor g06770(.dina(n6962), .dinb(n6961), .dout(n6963));
  jxor g06771(.dina(n6963), .dinb(n6960), .dout(n6964));
  jxor g06772(.dina(n6964), .dinb(n6958), .dout(n6965));
  jxor g06773(.dina(n6965), .dinb(n6951), .dout(n6966));
  jand g06774(.dina(\a[55] ), .dinb(\a[5] ), .dout(n6967));
  jnot g06775(.din(n6967), .dout(n6968));
  jand g06776(.dina(\a[54] ), .dinb(\a[6] ), .dout(n6969));
  jand g06777(.dina(\a[41] ), .dinb(\a[19] ), .dout(n6970));
  jxor g06778(.dina(n6970), .dinb(n6969), .dout(n6971));
  jxor g06779(.dina(n6971), .dinb(n6968), .dout(n6972));
  jnot g06780(.din(n6972), .dout(n6973));
  jand g06781(.dina(\a[53] ), .dinb(\a[7] ), .dout(n6974));
  jnot g06782(.din(n6974), .dout(n6975));
  jand g06783(.dina(\a[52] ), .dinb(\a[8] ), .dout(n6976));
  jand g06784(.dina(\a[42] ), .dinb(\a[18] ), .dout(n6977));
  jxor g06785(.dina(n6977), .dinb(n6976), .dout(n6978));
  jxor g06786(.dina(n6978), .dinb(n6975), .dout(n6979));
  jnot g06787(.din(n6074), .dout(n6980));
  jand g06788(.dina(\a[48] ), .dinb(\a[12] ), .dout(n6981));
  jand g06789(.dina(\a[47] ), .dinb(\a[13] ), .dout(n6982));
  jor  g06790(.dina(n6982), .dinb(n6981), .dout(n6983));
  jand g06791(.dina(\a[48] ), .dinb(\a[13] ), .dout(n6984));
  jand g06792(.dina(n6984), .dinb(n6825), .dout(n6985));
  jnot g06793(.din(n6985), .dout(n6986));
  jand g06794(.dina(n6986), .dinb(n6983), .dout(n6987));
  jxor g06795(.dina(n6987), .dinb(n6980), .dout(n6988));
  jxor g06796(.dina(n6988), .dinb(n6979), .dout(n6989));
  jxor g06797(.dina(n6989), .dinb(n6973), .dout(n6990));
  jxor g06798(.dina(n6990), .dinb(n6966), .dout(n6991));
  jxor g06799(.dina(n6991), .dinb(n6948), .dout(n6992));
  jand g06800(.dina(n6708), .dinb(n6705), .dout(n6993));
  jand g06801(.dina(n6709), .dinb(n6694), .dout(n6994));
  jor  g06802(.dina(n6994), .dinb(n6993), .dout(n6995));
  jand g06803(.dina(n6700), .dinb(n6697), .dout(n6996));
  jand g06804(.dina(n6704), .dinb(n6701), .dout(n6997));
  jor  g06805(.dina(n6997), .dinb(n6996), .dout(n6998));
  jand g06806(.dina(\a[36] ), .dinb(\a[24] ), .dout(n6999));
  jand g06807(.dina(\a[34] ), .dinb(\a[26] ), .dout(n7000));
  jor  g06808(.dina(n7000), .dinb(n6879), .dout(n7001));
  jnot g06809(.din(n7001), .dout(n7002));
  jand g06810(.dina(\a[35] ), .dinb(\a[26] ), .dout(n7003));
  jand g06811(.dina(n7003), .dinb(n6876), .dout(n7004));
  jor  g06812(.dina(n7004), .dinb(n7002), .dout(n7005));
  jxor g06813(.dina(n7005), .dinb(n6999), .dout(n7006));
  jand g06814(.dina(\a[40] ), .dinb(\a[20] ), .dout(n7007));
  jand g06815(.dina(\a[39] ), .dinb(\a[21] ), .dout(n7008));
  jor  g06816(.dina(n7008), .dinb(n6886), .dout(n7009));
  jnot g06817(.din(n7009), .dout(n7010));
  jand g06818(.dina(\a[39] ), .dinb(\a[22] ), .dout(n7011));
  jand g06819(.dina(n7011), .dinb(n6585), .dout(n7012));
  jor  g06820(.dina(n7012), .dinb(n7010), .dout(n7013));
  jxor g06821(.dina(n7013), .dinb(n7007), .dout(n7014));
  jand g06822(.dina(\a[58] ), .dinb(\a[2] ), .dout(n7015));
  jand g06823(.dina(\a[56] ), .dinb(\a[4] ), .dout(n7016));
  jor  g06824(.dina(n7016), .dinb(n6803), .dout(n7017));
  jand g06825(.dina(\a[57] ), .dinb(\a[4] ), .dout(n7018));
  jand g06826(.dina(n7018), .dinb(n6800), .dout(n7019));
  jnot g06827(.din(n7019), .dout(n7020));
  jand g06828(.dina(n7020), .dinb(n7017), .dout(n7021));
  jxor g06829(.dina(n7021), .dinb(n7015), .dout(n7022));
  jxor g06830(.dina(n7022), .dinb(n7014), .dout(n7023));
  jxor g06831(.dina(n7023), .dinb(n7006), .dout(n7024));
  jxor g06832(.dina(n7024), .dinb(n6998), .dout(n7025));
  jand g06833(.dina(\a[50] ), .dinb(\a[10] ), .dout(n7026));
  jand g06834(.dina(\a[49] ), .dinb(\a[11] ), .dout(n7027));
  jor  g06835(.dina(n7027), .dinb(n4852), .dout(n7028));
  jnot g06836(.din(n7028), .dout(n7029));
  jand g06837(.dina(n6845), .dinb(n6052), .dout(n7030));
  jor  g06838(.dina(n7030), .dinb(n7029), .dout(n7031));
  jxor g06839(.dina(n7031), .dinb(n7026), .dout(n7032));
  jnot g06840(.din(n7032), .dout(n7033));
  jand g06841(.dina(n6830), .dinb(n6824), .dout(n7034));
  jor  g06842(.dina(n7034), .dinb(n6828), .dout(n7035));
  jnot g06843(.din(n7035), .dout(n7036));
  jand g06844(.dina(\a[51] ), .dinb(\a[9] ), .dout(n7037));
  jand g06845(.dina(\a[44] ), .dinb(\a[16] ), .dout(n7038));
  jor  g06846(.dina(n7038), .dinb(n7037), .dout(n7039));
  jnot g06847(.din(n7039), .dout(n7040));
  jand g06848(.dina(\a[51] ), .dinb(\a[16] ), .dout(n7041));
  jand g06849(.dina(n7041), .dinb(n5471), .dout(n7042));
  jor  g06850(.dina(n7042), .dinb(n7040), .dout(n7043));
  jxor g06851(.dina(n7043), .dinb(n6813), .dout(n7044));
  jxor g06852(.dina(n7044), .dinb(n7036), .dout(n7045));
  jxor g06853(.dina(n7045), .dinb(n7033), .dout(n7046));
  jxor g06854(.dina(n7046), .dinb(n7025), .dout(n7047));
  jxor g06855(.dina(n7047), .dinb(n6995), .dout(n7048));
  jxor g06856(.dina(n7048), .dinb(n6992), .dout(n7049));
  jand g06857(.dina(n6710), .dinb(n6689), .dout(n7050));
  jand g06858(.dina(n6711), .dinb(n6686), .dout(n7051));
  jor  g06859(.dina(n7051), .dinb(n7050), .dout(n7052));
  jand g06860(.dina(n6857), .dinb(n6850), .dout(n7053));
  jor  g06861(.dina(n7053), .dinb(n6855), .dout(n7054));
  jand g06862(.dina(n6811), .dinb(n6618), .dout(n7055));
  jor  g06863(.dina(n7055), .dinb(n6814), .dout(n7056));
  jxor g06864(.dina(n7056), .dinb(n7054), .dout(n7057));
  jnot g06865(.din(n6820), .dout(n7058));
  jand g06866(.dina(n7058), .dinb(n6819), .dout(n7059));
  jnot g06867(.din(n7059), .dout(n7060));
  jand g06868(.dina(n6820), .dinb(n6818), .dout(n7061));
  jor  g06869(.dina(n7061), .dinb(n6371), .dout(n7062));
  jand g06870(.dina(n7062), .dinb(n7060), .dout(n7063));
  jxor g06871(.dina(n7063), .dinb(n7057), .dout(n7064));
  jnot g06872(.din(n6882), .dout(n7065));
  jor  g06873(.dina(n6890), .dinb(n7065), .dout(n7066));
  jnot g06874(.din(n6874), .dout(n7067));
  jand g06875(.dina(n6890), .dinb(n7065), .dout(n7068));
  jor  g06876(.dina(n7068), .dinb(n7067), .dout(n7069));
  jand g06877(.dina(n7069), .dinb(n7066), .dout(n7070));
  jxor g06878(.dina(n7070), .dinb(n7064), .dout(n7071));
  jor  g06879(.dina(n6831), .dinb(n6823), .dout(n7072));
  jand g06880(.dina(n6831), .dinb(n6823), .dout(n7073));
  jor  g06881(.dina(n7073), .dinb(n6817), .dout(n7074));
  jand g06882(.dina(n7074), .dinb(n7072), .dout(n7075));
  jxor g06883(.dina(n7075), .dinb(n7071), .dout(n7076));
  jand g06884(.dina(n6833), .dinb(n6808), .dout(n7077));
  jand g06885(.dina(n6834), .dinb(n6788), .dout(n7078));
  jor  g06886(.dina(n7078), .dinb(n7077), .dout(n7079));
  jand g06887(.dina(n6858), .dinb(n6849), .dout(n7080));
  jand g06888(.dina(n6859), .dinb(n6839), .dout(n7081));
  jor  g06889(.dina(n7081), .dinb(n7080), .dout(n7082));
  jand g06890(.dina(n6889), .dinb(n6883), .dout(n7083));
  jor  g06891(.dina(n7083), .dinb(n6887), .dout(n7084));
  jnot g06892(.din(n7084), .dout(n7085));
  jand g06893(.dina(n6791), .dinb(n6790), .dout(n7086));
  jnot g06894(.din(n7086), .dout(n7087));
  jnot g06895(.din(n6790), .dout(n7088));
  jnot g06896(.din(n6791), .dout(n7089));
  jand g06897(.dina(n7089), .dinb(n7088), .dout(n7090));
  jor  g06898(.dina(n7090), .dinb(n6789), .dout(n7091));
  jand g06899(.dina(n7091), .dinb(n7087), .dout(n7092));
  jxor g06900(.dina(n7092), .dinb(n7085), .dout(n7093));
  jand g06901(.dina(n6877), .dinb(n6875), .dout(n7094));
  jor  g06902(.dina(n7094), .dinb(n6880), .dout(n7095));
  jxor g06903(.dina(n7095), .dinb(n7093), .dout(n7096));
  jand g06904(.dina(n6801), .dinb(n6798), .dout(n7097));
  jor  g06905(.dina(n7097), .dinb(n6804), .dout(n7098));
  jand g06906(.dina(n6869), .dinb(n6867), .dout(n7099));
  jor  g06907(.dina(n7099), .dinb(n6872), .dout(n7100));
  jxor g06908(.dina(n7100), .dinb(n7098), .dout(n7101));
  jand g06909(.dina(n6843), .dinb(n6840), .dout(n7102));
  jor  g06910(.dina(n7102), .dinb(n6846), .dout(n7103));
  jxor g06911(.dina(n7103), .dinb(n7101), .dout(n7104));
  jxor g06912(.dina(n7104), .dinb(n7096), .dout(n7105));
  jxor g06913(.dina(n7105), .dinb(n7082), .dout(n7106));
  jxor g06914(.dina(n7106), .dinb(n7079), .dout(n7107));
  jxor g06915(.dina(n7107), .dinb(n7076), .dout(n7108));
  jxor g06916(.dina(n7108), .dinb(n7052), .dout(n7109));
  jxor g06917(.dina(n7109), .dinb(n7049), .dout(n7110));
  jxor g06918(.dina(n7110), .dinb(n6945), .dout(n7111));
  jxor g06919(.dina(n7111), .dinb(n6908), .dout(n7112));
  jand g06920(.dina(n6899), .dinb(n6896), .dout(n7113));
  jnot g06921(.din(n6896), .dout(n7114));
  jnot g06922(.din(n6899), .dout(n7115));
  jand g06923(.dina(n7115), .dinb(n7114), .dout(n7116));
  jnot g06924(.din(n7116), .dout(n7117));
  jand g06925(.dina(n6904), .dinb(n7117), .dout(n7118));
  jor  g06926(.dina(n7118), .dinb(n7113), .dout(n7119));
  jxor g06927(.dina(n7119), .dinb(n7112), .dout(\asquared[61] ));
  jand g06928(.dina(n6944), .dinb(n6911), .dout(n7121));
  jand g06929(.dina(n7110), .dinb(n6945), .dout(n7122));
  jor  g06930(.dina(n7122), .dinb(n7121), .dout(n7123));
  jand g06931(.dina(n6942), .dinb(n6917), .dout(n7124));
  jand g06932(.dina(n6943), .dinb(n6914), .dout(n7125));
  jor  g06933(.dina(n7125), .dinb(n7124), .dout(n7126));
  jand g06934(.dina(n6990), .dinb(n6966), .dout(n7127));
  jand g06935(.dina(n6991), .dinb(n6948), .dout(n7128));
  jor  g06936(.dina(n7128), .dinb(n7127), .dout(n7129));
  jand g06937(.dina(n7039), .dinb(n6813), .dout(n7130));
  jor  g06938(.dina(n7130), .dinb(n7042), .dout(n7131));
  jand g06939(.dina(n6977), .dinb(n6976), .dout(n7132));
  jnot g06940(.din(n7132), .dout(n7133));
  jnot g06941(.din(n6976), .dout(n7134));
  jnot g06942(.din(n6977), .dout(n7135));
  jand g06943(.dina(n7135), .dinb(n7134), .dout(n7136));
  jor  g06944(.dina(n7136), .dinb(n6975), .dout(n7137));
  jand g06945(.dina(n7137), .dinb(n7133), .dout(n7138));
  jnot g06946(.din(n7138), .dout(n7139));
  jxor g06947(.dina(n7139), .dinb(n7131), .dout(n7140));
  jnot g06948(.din(n6952), .dout(n7141));
  jand g06949(.dina(n7141), .dinb(n6768), .dout(n7142));
  jnot g06950(.din(n7142), .dout(n7143));
  jand g06951(.dina(n6952), .dinb(n6767), .dout(n7144));
  jor  g06952(.dina(n6956), .dinb(n7144), .dout(n7145));
  jand g06953(.dina(n7145), .dinb(n7143), .dout(n7146));
  jxor g06954(.dina(n7146), .dinb(n7140), .dout(n7147));
  jand g06955(.dina(n6988), .dinb(n6979), .dout(n7148));
  jnot g06956(.din(n7148), .dout(n7149));
  jnot g06957(.din(n6979), .dout(n7150));
  jnot g06958(.din(n6988), .dout(n7151));
  jand g06959(.dina(n7151), .dinb(n7150), .dout(n7152));
  jor  g06960(.dina(n7152), .dinb(n6973), .dout(n7153));
  jand g06961(.dina(n7153), .dinb(n7149), .dout(n7154));
  jxor g06962(.dina(n7154), .dinb(n7147), .dout(n7155));
  jnot g06963(.din(n7155), .dout(n7156));
  jor  g06964(.dina(n6964), .dinb(n6958), .dout(n7157));
  jand g06965(.dina(n6965), .dinb(n6951), .dout(n7158));
  jnot g06966(.din(n7158), .dout(n7159));
  jand g06967(.dina(n7159), .dinb(n7157), .dout(n7160));
  jxor g06968(.dina(n7160), .dinb(n7156), .dout(n7161));
  jand g06969(.dina(n7001), .dinb(n6999), .dout(n7162));
  jor  g06970(.dina(n7162), .dinb(n7004), .dout(n7163));
  jand g06971(.dina(n6962), .dinb(n6961), .dout(n7164));
  jnot g06972(.din(n7164), .dout(n7165));
  jnot g06973(.din(n6961), .dout(n7166));
  jnot g06974(.din(n6962), .dout(n7167));
  jand g06975(.dina(n7167), .dinb(n7166), .dout(n7168));
  jor  g06976(.dina(n7168), .dinb(n6960), .dout(n7169));
  jand g06977(.dina(n7169), .dinb(n7165), .dout(n7170));
  jnot g06978(.din(n7170), .dout(n7171));
  jxor g06979(.dina(n7171), .dinb(n7163), .dout(n7172));
  jand g06980(.dina(n7009), .dinb(n7007), .dout(n7173));
  jor  g06981(.dina(n7173), .dinb(n7012), .dout(n7174));
  jxor g06982(.dina(n7174), .dinb(n7172), .dout(n7175));
  jand g06983(.dina(n7021), .dinb(n7015), .dout(n7176));
  jor  g06984(.dina(n7176), .dinb(n7019), .dout(n7177));
  jnot g06985(.din(n7177), .dout(n7178));
  jand g06986(.dina(n6970), .dinb(n6969), .dout(n7179));
  jnot g06987(.din(n7179), .dout(n7180));
  jnot g06988(.din(n6969), .dout(n7181));
  jnot g06989(.din(n6970), .dout(n7182));
  jand g06990(.dina(n7182), .dinb(n7181), .dout(n7183));
  jor  g06991(.dina(n7183), .dinb(n6968), .dout(n7184));
  jand g06992(.dina(n7184), .dinb(n7180), .dout(n7185));
  jxor g06993(.dina(n7185), .dinb(n7178), .dout(n7186));
  jand g06994(.dina(n7028), .dinb(n7026), .dout(n7187));
  jor  g06995(.dina(n7187), .dinb(n7030), .dout(n7188));
  jxor g06996(.dina(n7188), .dinb(n7186), .dout(n7189));
  jxor g06997(.dina(n7189), .dinb(n7175), .dout(n7190));
  jnot g06998(.din(n7014), .dout(n7191));
  jor  g06999(.dina(n7022), .dinb(n7191), .dout(n7192));
  jnot g07000(.din(n7006), .dout(n7193));
  jand g07001(.dina(n7022), .dinb(n7191), .dout(n7194));
  jor  g07002(.dina(n7194), .dinb(n7193), .dout(n7195));
  jand g07003(.dina(n7195), .dinb(n7192), .dout(n7196));
  jxor g07004(.dina(n7196), .dinb(n7190), .dout(n7197));
  jxor g07005(.dina(n7197), .dinb(n7161), .dout(n7198));
  jxor g07006(.dina(n7198), .dinb(n7129), .dout(n7199));
  jxor g07007(.dina(n7199), .dinb(n7126), .dout(n7200));
  jand g07008(.dina(n7106), .dinb(n7079), .dout(n7201));
  jand g07009(.dina(n7107), .dinb(n7076), .dout(n7202));
  jor  g07010(.dina(n7202), .dinb(n7201), .dout(n7203));
  jor  g07011(.dina(n6935), .dinb(n6931), .dout(n7204));
  jor  g07012(.dina(n6941), .dinb(n6937), .dout(n7205));
  jand g07013(.dina(n7205), .dinb(n7204), .dout(n7206));
  jnot g07014(.din(n7206), .dout(n7207));
  jand g07015(.dina(n6923), .dinb(n6920), .dout(n7208));
  jnot g07016(.din(n7208), .dout(n7209));
  jor  g07017(.dina(n6929), .dinb(n6925), .dout(n7210));
  jand g07018(.dina(n7210), .dinb(n7209), .dout(n7211));
  jnot g07019(.din(n7211), .dout(n7212));
  jand g07020(.dina(\a[31] ), .dinb(\a[30] ), .dout(n7213));
  jand g07021(.dina(\a[32] ), .dinb(\a[29] ), .dout(n7214));
  jor  g07022(.dina(n7214), .dinb(n7213), .dout(n7215));
  jnot g07023(.din(n7215), .dout(n7216));
  jand g07024(.dina(\a[32] ), .dinb(\a[30] ), .dout(n7217));
  jand g07025(.dina(n7217), .dinb(n6954), .dout(n7218));
  jor  g07026(.dina(n7218), .dinb(n7216), .dout(n7219));
  jxor g07027(.dina(n7219), .dinb(n6984), .dout(n7220));
  jnot g07028(.din(n7220), .dout(n7221));
  jand g07029(.dina(\a[50] ), .dinb(\a[11] ), .dout(n7222));
  jand g07030(.dina(\a[49] ), .dinb(\a[12] ), .dout(n7223));
  jor  g07031(.dina(n7223), .dinb(n6827), .dout(n7224));
  jnot g07032(.din(n7224), .dout(n7225));
  jand g07033(.dina(\a[49] ), .dinb(\a[14] ), .dout(n7226));
  jand g07034(.dina(n7226), .dinb(n6825), .dout(n7227));
  jor  g07035(.dina(n7227), .dinb(n7225), .dout(n7228));
  jxor g07036(.dina(n7228), .dinb(n7222), .dout(n7229));
  jand g07037(.dina(\a[45] ), .dinb(\a[16] ), .dout(n7230));
  jand g07038(.dina(\a[46] ), .dinb(\a[15] ), .dout(n7231));
  jand g07039(.dina(\a[51] ), .dinb(\a[10] ), .dout(n7232));
  jor  g07040(.dina(n7232), .dinb(n7231), .dout(n7233));
  jnot g07041(.din(n7233), .dout(n7234));
  jand g07042(.dina(\a[51] ), .dinb(\a[15] ), .dout(n7235));
  jand g07043(.dina(n7235), .dinb(n6071), .dout(n7236));
  jor  g07044(.dina(n7236), .dinb(n7234), .dout(n7237));
  jxor g07045(.dina(n7237), .dinb(n7230), .dout(n7238));
  jxor g07046(.dina(n7238), .dinb(n7229), .dout(n7239));
  jxor g07047(.dina(n7239), .dinb(n7221), .dout(n7240));
  jxor g07048(.dina(n7240), .dinb(n7212), .dout(n7241));
  jand g07049(.dina(\a[37] ), .dinb(\a[24] ), .dout(n7242));
  jand g07050(.dina(\a[36] ), .dinb(\a[25] ), .dout(n7243));
  jor  g07051(.dina(n7243), .dinb(n7242), .dout(n7244));
  jnot g07052(.din(n7244), .dout(n7245));
  jand g07053(.dina(\a[37] ), .dinb(\a[25] ), .dout(n7246));
  jand g07054(.dina(n7246), .dinb(n6999), .dout(n7247));
  jor  g07055(.dina(n7247), .dinb(n7245), .dout(n7248));
  jxor g07056(.dina(n7248), .dinb(n7011), .dout(n7249));
  jand g07057(.dina(\a[55] ), .dinb(\a[6] ), .dout(n7250));
  jand g07058(.dina(\a[41] ), .dinb(\a[20] ), .dout(n7251));
  jand g07059(.dina(\a[40] ), .dinb(\a[21] ), .dout(n7252));
  jor  g07060(.dina(n7252), .dinb(n7251), .dout(n7253));
  jnot g07061(.din(n7253), .dout(n7254));
  jand g07062(.dina(\a[41] ), .dinb(\a[21] ), .dout(n7255));
  jand g07063(.dina(n7255), .dinb(n7007), .dout(n7256));
  jor  g07064(.dina(n7256), .dinb(n7254), .dout(n7257));
  jxor g07065(.dina(n7257), .dinb(n7250), .dout(n7258));
  jand g07066(.dina(\a[61] ), .dinb(\a[0] ), .dout(n7259));
  jand g07067(.dina(\a[59] ), .dinb(\a[2] ), .dout(n7260));
  jand g07068(.dina(\a[56] ), .dinb(\a[5] ), .dout(n7261));
  jor  g07069(.dina(n7261), .dinb(n7260), .dout(n7262));
  jand g07070(.dina(\a[59] ), .dinb(\a[5] ), .dout(n7263));
  jand g07071(.dina(n7263), .dinb(n6100), .dout(n7264));
  jnot g07072(.din(n7264), .dout(n7265));
  jand g07073(.dina(n7265), .dinb(n7262), .dout(n7266));
  jxor g07074(.dina(n7266), .dinb(n7259), .dout(n7267));
  jxor g07075(.dina(n7267), .dinb(n7258), .dout(n7268));
  jxor g07076(.dina(n7268), .dinb(n7249), .dout(n7269));
  jxor g07077(.dina(n7269), .dinb(n7241), .dout(n7270));
  jxor g07078(.dina(n7270), .dinb(n7207), .dout(n7271));
  jxor g07079(.dina(n7271), .dinb(n7203), .dout(n7272));
  jxor g07080(.dina(n7272), .dinb(n7200), .dout(n7273));
  jand g07081(.dina(n7108), .dinb(n7052), .dout(n7274));
  jand g07082(.dina(n7109), .dinb(n7049), .dout(n7275));
  jor  g07083(.dina(n7275), .dinb(n7274), .dout(n7276));
  jand g07084(.dina(n7047), .dinb(n6995), .dout(n7277));
  jand g07085(.dina(n7048), .dinb(n6992), .dout(n7278));
  jor  g07086(.dina(n7278), .dinb(n7277), .dout(n7279));
  jand g07087(.dina(n7024), .dinb(n6998), .dout(n7280));
  jand g07088(.dina(n7046), .dinb(n7025), .dout(n7281));
  jor  g07089(.dina(n7281), .dinb(n7280), .dout(n7282));
  jor  g07090(.dina(n7044), .dinb(n7036), .dout(n7283));
  jand g07091(.dina(n7045), .dinb(n7033), .dout(n7284));
  jnot g07092(.din(n7284), .dout(n7285));
  jand g07093(.dina(n7285), .dinb(n7283), .dout(n7286));
  jnot g07094(.din(n7286), .dout(n7287));
  jor  g07095(.dina(n7092), .dinb(n7085), .dout(n7288));
  jand g07096(.dina(n7095), .dinb(n7093), .dout(n7289));
  jnot g07097(.din(n7289), .dout(n7290));
  jand g07098(.dina(n7290), .dinb(n7288), .dout(n7291));
  jnot g07099(.din(n7291), .dout(n7292));
  jand g07100(.dina(\a[60] ), .dinb(\a[1] ), .dout(n7293));
  jnot g07101(.din(\a[31] ), .dout(n7294));
  jand g07102(.dina(n6955), .dinb(n6954), .dout(n7295));
  jor  g07103(.dina(n7295), .dinb(n7294), .dout(n7296));
  jxor g07104(.dina(n7296), .dinb(n7293), .dout(n7297));
  jnot g07105(.din(n7297), .dout(n7298));
  jand g07106(.dina(n6986), .dinb(n6980), .dout(n7299));
  jnot g07107(.din(n7299), .dout(n7300));
  jand g07108(.dina(n7300), .dinb(n6983), .dout(n7301));
  jxor g07109(.dina(n7301), .dinb(n7298), .dout(n7302));
  jxor g07110(.dina(n7302), .dinb(n7292), .dout(n7303));
  jxor g07111(.dina(n7303), .dinb(n7287), .dout(n7304));
  jand g07112(.dina(n7100), .dinb(n7098), .dout(n7305));
  jand g07113(.dina(n7103), .dinb(n7101), .dout(n7306));
  jor  g07114(.dina(n7306), .dinb(n7305), .dout(n7307));
  jand g07115(.dina(n7056), .dinb(n7054), .dout(n7308));
  jand g07116(.dina(n7063), .dinb(n7057), .dout(n7309));
  jor  g07117(.dina(n7309), .dinb(n7308), .dout(n7310));
  jnot g07118(.din(n7310), .dout(n7311));
  jand g07119(.dina(\a[38] ), .dinb(\a[23] ), .dout(n7312));
  jand g07120(.dina(\a[58] ), .dinb(\a[3] ), .dout(n7313));
  jor  g07121(.dina(n7313), .dinb(n7018), .dout(n7314));
  jnot g07122(.din(n7314), .dout(n7315));
  jand g07123(.dina(\a[58] ), .dinb(\a[4] ), .dout(n7316));
  jand g07124(.dina(n7316), .dinb(n6803), .dout(n7317));
  jor  g07125(.dina(n7317), .dinb(n7315), .dout(n7318));
  jxor g07126(.dina(n7318), .dinb(n7312), .dout(n7319));
  jxor g07127(.dina(n7319), .dinb(n7311), .dout(n7320));
  jxor g07128(.dina(n7320), .dinb(n7307), .dout(n7321));
  jxor g07129(.dina(n7321), .dinb(n7304), .dout(n7322));
  jxor g07130(.dina(n7322), .dinb(n7282), .dout(n7323));
  jand g07131(.dina(n7070), .dinb(n7064), .dout(n7324));
  jand g07132(.dina(n7075), .dinb(n7071), .dout(n7325));
  jor  g07133(.dina(n7325), .dinb(n7324), .dout(n7326));
  jand g07134(.dina(n7104), .dinb(n7096), .dout(n7327));
  jand g07135(.dina(n7105), .dinb(n7082), .dout(n7328));
  jor  g07136(.dina(n7328), .dinb(n7327), .dout(n7329));
  jand g07137(.dina(\a[34] ), .dinb(\a[27] ), .dout(n7330));
  jand g07138(.dina(\a[33] ), .dinb(\a[28] ), .dout(n7331));
  jor  g07139(.dina(n7331), .dinb(n7330), .dout(n7332));
  jnot g07140(.din(n7332), .dout(n7333));
  jand g07141(.dina(\a[34] ), .dinb(\a[28] ), .dout(n7334));
  jand g07142(.dina(n7334), .dinb(n6959), .dout(n7335));
  jor  g07143(.dina(n7335), .dinb(n7333), .dout(n7336));
  jxor g07144(.dina(n7336), .dinb(n7003), .dout(n7337));
  jand g07145(.dina(\a[43] ), .dinb(\a[18] ), .dout(n7338));
  jand g07146(.dina(\a[52] ), .dinb(\a[9] ), .dout(n7339));
  jand g07147(.dina(\a[44] ), .dinb(\a[17] ), .dout(n7340));
  jor  g07148(.dina(n7340), .dinb(n7339), .dout(n7341));
  jnot g07149(.din(n7341), .dout(n7342));
  jand g07150(.dina(\a[52] ), .dinb(\a[17] ), .dout(n7343));
  jand g07151(.dina(n7343), .dinb(n5471), .dout(n7344));
  jor  g07152(.dina(n7344), .dinb(n7342), .dout(n7345));
  jxor g07153(.dina(n7345), .dinb(n7338), .dout(n7346));
  jand g07154(.dina(\a[42] ), .dinb(\a[19] ), .dout(n7347));
  jand g07155(.dina(\a[54] ), .dinb(\a[7] ), .dout(n7348));
  jand g07156(.dina(\a[53] ), .dinb(\a[8] ), .dout(n7349));
  jor  g07157(.dina(n7349), .dinb(n7348), .dout(n7350));
  jand g07158(.dina(\a[54] ), .dinb(\a[8] ), .dout(n7351));
  jand g07159(.dina(n7351), .dinb(n6974), .dout(n7352));
  jnot g07160(.din(n7352), .dout(n7353));
  jand g07161(.dina(n7353), .dinb(n7350), .dout(n7354));
  jxor g07162(.dina(n7354), .dinb(n7347), .dout(n7355));
  jxor g07163(.dina(n7355), .dinb(n7346), .dout(n7356));
  jxor g07164(.dina(n7356), .dinb(n7337), .dout(n7357));
  jxor g07165(.dina(n7357), .dinb(n7329), .dout(n7358));
  jxor g07166(.dina(n7358), .dinb(n7326), .dout(n7359));
  jxor g07167(.dina(n7359), .dinb(n7323), .dout(n7360));
  jxor g07168(.dina(n7360), .dinb(n7279), .dout(n7361));
  jxor g07169(.dina(n7361), .dinb(n7276), .dout(n7362));
  jxor g07170(.dina(n7362), .dinb(n7273), .dout(n7363));
  jxor g07171(.dina(n7363), .dinb(n7123), .dout(n7364));
  jand g07172(.dina(n7111), .dinb(n6908), .dout(n7365));
  jnot g07173(.din(n6908), .dout(n7366));
  jnot g07174(.din(n7111), .dout(n7367));
  jand g07175(.dina(n7367), .dinb(n7366), .dout(n7368));
  jnot g07176(.din(n7368), .dout(n7369));
  jand g07177(.dina(n7119), .dinb(n7369), .dout(n7370));
  jor  g07178(.dina(n7370), .dinb(n7365), .dout(n7371));
  jxor g07179(.dina(n7371), .dinb(n7364), .dout(\asquared[62] ));
  jand g07180(.dina(n7361), .dinb(n7276), .dout(n7373));
  jand g07181(.dina(n7362), .dinb(n7273), .dout(n7374));
  jor  g07182(.dina(n7374), .dinb(n7373), .dout(n7375));
  jand g07183(.dina(n7359), .dinb(n7323), .dout(n7376));
  jand g07184(.dina(n7360), .dinb(n7279), .dout(n7377));
  jor  g07185(.dina(n7377), .dinb(n7376), .dout(n7378));
  jand g07186(.dina(n7233), .dinb(n7230), .dout(n7379));
  jor  g07187(.dina(n7379), .dinb(n7236), .dout(n7380));
  jand g07188(.dina(n7341), .dinb(n7338), .dout(n7381));
  jor  g07189(.dina(n7381), .dinb(n7344), .dout(n7382));
  jxor g07190(.dina(n7382), .dinb(n7380), .dout(n7383));
  jand g07191(.dina(\a[59] ), .dinb(\a[3] ), .dout(n7384));
  jand g07192(.dina(\a[57] ), .dinb(\a[5] ), .dout(n7385));
  jor  g07193(.dina(n7385), .dinb(n7316), .dout(n7386));
  jnot g07194(.din(n7386), .dout(n7387));
  jand g07195(.dina(\a[58] ), .dinb(\a[5] ), .dout(n7388));
  jand g07196(.dina(n7388), .dinb(n7018), .dout(n7389));
  jor  g07197(.dina(n7389), .dinb(n7387), .dout(n7390));
  jxor g07198(.dina(n7390), .dinb(n7384), .dout(n7391));
  jnot g07199(.din(n7391), .dout(n7392));
  jxor g07200(.dina(n7392), .dinb(n7383), .dout(n7393));
  jnot g07201(.din(n7346), .dout(n7394));
  jor  g07202(.dina(n7355), .dinb(n7394), .dout(n7395));
  jnot g07203(.din(n7337), .dout(n7396));
  jand g07204(.dina(n7355), .dinb(n7394), .dout(n7397));
  jor  g07205(.dina(n7397), .dinb(n7396), .dout(n7398));
  jand g07206(.dina(n7398), .dinb(n7395), .dout(n7399));
  jxor g07207(.dina(n7399), .dinb(n7393), .dout(n7400));
  jnot g07208(.din(n7400), .dout(n7401));
  jor  g07209(.dina(n7319), .dinb(n7311), .dout(n7402));
  jand g07210(.dina(n7320), .dinb(n7307), .dout(n7403));
  jnot g07211(.din(n7403), .dout(n7404));
  jand g07212(.dina(n7404), .dinb(n7402), .dout(n7405));
  jxor g07213(.dina(n7405), .dinb(n7401), .dout(n7406));
  jand g07214(.dina(n7139), .dinb(n7131), .dout(n7407));
  jand g07215(.dina(n7146), .dinb(n7140), .dout(n7408));
  jor  g07216(.dina(n7408), .dinb(n7407), .dout(n7409));
  jand g07217(.dina(n7301), .dinb(n7298), .dout(n7410));
  jnot g07218(.din(\a[60] ), .dout(n7411));
  jand g07219(.dina(n7295), .dinb(n7411), .dout(n7412));
  jor  g07220(.dina(n7412), .dinb(n7410), .dout(n7413));
  jxor g07221(.dina(n7413), .dinb(n7409), .dout(n7414));
  jand g07222(.dina(n7171), .dinb(n7163), .dout(n7415));
  jand g07223(.dina(n7174), .dinb(n7172), .dout(n7416));
  jor  g07224(.dina(n7416), .dinb(n7415), .dout(n7417));
  jxor g07225(.dina(n7417), .dinb(n7414), .dout(n7418));
  jand g07226(.dina(n7240), .dinb(n7212), .dout(n7419));
  jand g07227(.dina(n7269), .dinb(n7241), .dout(n7420));
  jor  g07228(.dina(n7420), .dinb(n7419), .dout(n7421));
  jxor g07229(.dina(n7421), .dinb(n7418), .dout(n7422));
  jxor g07230(.dina(n7422), .dinb(n7406), .dout(n7423));
  jxor g07231(.dina(n7423), .dinb(n7378), .dout(n7424));
  jand g07232(.dina(n7197), .dinb(n7161), .dout(n7425));
  jand g07233(.dina(n7198), .dinb(n7129), .dout(n7426));
  jor  g07234(.dina(n7426), .dinb(n7425), .dout(n7427));
  jand g07235(.dina(n7321), .dinb(n7304), .dout(n7428));
  jand g07236(.dina(n7322), .dinb(n7282), .dout(n7429));
  jor  g07237(.dina(n7429), .dinb(n7428), .dout(n7430));
  jand g07238(.dina(\a[53] ), .dinb(\a[9] ), .dout(n7431));
  jnot g07239(.din(n7431), .dout(n7432));
  jand g07240(.dina(\a[52] ), .dinb(\a[10] ), .dout(n7433));
  jand g07241(.dina(\a[45] ), .dinb(\a[17] ), .dout(n7434));
  jor  g07242(.dina(n7434), .dinb(n7433), .dout(n7435));
  jand g07243(.dina(n7343), .dinb(n5941), .dout(n7436));
  jnot g07244(.din(n7436), .dout(n7437));
  jand g07245(.dina(n7437), .dinb(n7435), .dout(n7438));
  jxor g07246(.dina(n7438), .dinb(n7432), .dout(n7439));
  jnot g07247(.din(n7255), .dout(n7440));
  jand g07248(.dina(\a[36] ), .dinb(\a[26] ), .dout(n7441));
  jor  g07249(.dina(n7441), .dinb(n7246), .dout(n7442));
  jand g07250(.dina(\a[37] ), .dinb(\a[26] ), .dout(n7443));
  jand g07251(.dina(n7443), .dinb(n7243), .dout(n7444));
  jnot g07252(.din(n7444), .dout(n7445));
  jand g07253(.dina(n7445), .dinb(n7442), .dout(n7446));
  jxor g07254(.dina(n7446), .dinb(n7440), .dout(n7447));
  jnot g07255(.din(n7447), .dout(n7448));
  jand g07256(.dina(n7293), .dinb(\a[31] ), .dout(n7449));
  jnot g07257(.din(n7449), .dout(n7450));
  jand g07258(.dina(\a[62] ), .dinb(\a[0] ), .dout(n7451));
  jand g07259(.dina(\a[60] ), .dinb(\a[2] ), .dout(n7452));
  jor  g07260(.dina(n7452), .dinb(n7451), .dout(n7453));
  jand g07261(.dina(\a[62] ), .dinb(\a[2] ), .dout(n7454));
  jand g07262(.dina(n7454), .dinb(n6952), .dout(n7455));
  jnot g07263(.din(n7455), .dout(n7456));
  jand g07264(.dina(n7456), .dinb(n7453), .dout(n7457));
  jxor g07265(.dina(n7457), .dinb(n7450), .dout(n7458));
  jxor g07266(.dina(n7458), .dinb(n7448), .dout(n7459));
  jxor g07267(.dina(n7459), .dinb(n7439), .dout(n7460));
  jand g07268(.dina(\a[42] ), .dinb(\a[20] ), .dout(n7461));
  jand g07269(.dina(\a[56] ), .dinb(\a[6] ), .dout(n7462));
  jand g07270(.dina(\a[55] ), .dinb(\a[7] ), .dout(n7463));
  jor  g07271(.dina(n7463), .dinb(n7462), .dout(n7464));
  jnot g07272(.din(n7464), .dout(n7465));
  jand g07273(.dina(\a[56] ), .dinb(\a[7] ), .dout(n7466));
  jand g07274(.dina(n7466), .dinb(n7250), .dout(n7467));
  jor  g07275(.dina(n7467), .dinb(n7465), .dout(n7468));
  jxor g07276(.dina(n7468), .dinb(n7461), .dout(n7469));
  jand g07277(.dina(\a[50] ), .dinb(\a[12] ), .dout(n7470));
  jand g07278(.dina(\a[49] ), .dinb(\a[13] ), .dout(n7471));
  jand g07279(.dina(\a[48] ), .dinb(\a[14] ), .dout(n7472));
  jor  g07280(.dina(n7472), .dinb(n7471), .dout(n7473));
  jnot g07281(.din(n7473), .dout(n7474));
  jand g07282(.dina(n7226), .dinb(n6984), .dout(n7475));
  jor  g07283(.dina(n7475), .dinb(n7474), .dout(n7476));
  jxor g07284(.dina(n7476), .dinb(n7470), .dout(n7477));
  jand g07285(.dina(\a[51] ), .dinb(\a[11] ), .dout(n7478));
  jor  g07286(.dina(n7478), .dinb(n6656), .dout(n7479));
  jand g07287(.dina(n7235), .dinb(n6654), .dout(n7480));
  jnot g07288(.din(n7480), .dout(n7481));
  jand g07289(.dina(n7481), .dinb(n7479), .dout(n7482));
  jxor g07290(.dina(n7482), .dinb(n5273), .dout(n7483));
  jxor g07291(.dina(n7483), .dinb(n7477), .dout(n7484));
  jxor g07292(.dina(n7484), .dinb(n7469), .dout(n7485));
  jxor g07293(.dina(n7485), .dinb(n7460), .dout(n7486));
  jand g07294(.dina(\a[40] ), .dinb(\a[22] ), .dout(n7487));
  jand g07295(.dina(\a[39] ), .dinb(\a[23] ), .dout(n7488));
  jand g07296(.dina(\a[38] ), .dinb(\a[24] ), .dout(n7489));
  jor  g07297(.dina(n7489), .dinb(n7488), .dout(n7490));
  jnot g07298(.din(n7490), .dout(n7491));
  jand g07299(.dina(\a[39] ), .dinb(\a[24] ), .dout(n7492));
  jand g07300(.dina(n7492), .dinb(n7312), .dout(n7493));
  jor  g07301(.dina(n7493), .dinb(n7491), .dout(n7494));
  jxor g07302(.dina(n7494), .dinb(n7487), .dout(n7495));
  jand g07303(.dina(\a[35] ), .dinb(\a[27] ), .dout(n7496));
  jand g07304(.dina(\a[33] ), .dinb(\a[29] ), .dout(n7497));
  jor  g07305(.dina(n7497), .dinb(n7334), .dout(n7498));
  jnot g07306(.din(n7498), .dout(n7499));
  jand g07307(.dina(\a[34] ), .dinb(\a[29] ), .dout(n7500));
  jand g07308(.dina(n7500), .dinb(n7331), .dout(n7501));
  jor  g07309(.dina(n7501), .dinb(n7499), .dout(n7502));
  jxor g07310(.dina(n7502), .dinb(n7496), .dout(n7503));
  jand g07311(.dina(\a[43] ), .dinb(\a[19] ), .dout(n7504));
  jand g07312(.dina(\a[44] ), .dinb(\a[18] ), .dout(n7505));
  jor  g07313(.dina(n7505), .dinb(n7351), .dout(n7506));
  jand g07314(.dina(\a[54] ), .dinb(\a[18] ), .dout(n7507));
  jand g07315(.dina(n7507), .dinb(n5255), .dout(n7508));
  jnot g07316(.din(n7508), .dout(n7509));
  jand g07317(.dina(n7509), .dinb(n7506), .dout(n7510));
  jxor g07318(.dina(n7510), .dinb(n7504), .dout(n7511));
  jxor g07319(.dina(n7511), .dinb(n7503), .dout(n7512));
  jxor g07320(.dina(n7512), .dinb(n7495), .dout(n7513));
  jxor g07321(.dina(n7513), .dinb(n7486), .dout(n7514));
  jxor g07322(.dina(n7514), .dinb(n7430), .dout(n7515));
  jxor g07323(.dina(n7515), .dinb(n7427), .dout(n7516));
  jxor g07324(.dina(n7516), .dinb(n7424), .dout(n7517));
  jand g07325(.dina(n7199), .dinb(n7126), .dout(n7518));
  jand g07326(.dina(n7272), .dinb(n7200), .dout(n7519));
  jor  g07327(.dina(n7519), .dinb(n7518), .dout(n7520));
  jand g07328(.dina(n7357), .dinb(n7329), .dout(n7521));
  jand g07329(.dina(n7358), .dinb(n7326), .dout(n7522));
  jor  g07330(.dina(n7522), .dinb(n7521), .dout(n7523));
  jor  g07331(.dina(n7185), .dinb(n7178), .dout(n7524));
  jand g07332(.dina(n7188), .dinb(n7186), .dout(n7525));
  jnot g07333(.din(n7525), .dout(n7526));
  jand g07334(.dina(n7526), .dinb(n7524), .dout(n7527));
  jnot g07335(.din(n7527), .dout(n7528));
  jnot g07336(.din(n7258), .dout(n7529));
  jor  g07337(.dina(n7267), .dinb(n7529), .dout(n7530));
  jnot g07338(.din(n7249), .dout(n7531));
  jand g07339(.dina(n7267), .dinb(n7529), .dout(n7532));
  jor  g07340(.dina(n7532), .dinb(n7531), .dout(n7533));
  jand g07341(.dina(n7533), .dinb(n7530), .dout(n7534));
  jxor g07342(.dina(n7534), .dinb(n7528), .dout(n7535));
  jnot g07343(.din(n7535), .dout(n7536));
  jor  g07344(.dina(n7238), .dinb(n7229), .dout(n7537));
  jand g07345(.dina(n7239), .dinb(n7221), .dout(n7538));
  jnot g07346(.din(n7538), .dout(n7539));
  jand g07347(.dina(n7539), .dinb(n7537), .dout(n7540));
  jxor g07348(.dina(n7540), .dinb(n7536), .dout(n7541));
  jand g07349(.dina(n7354), .dinb(n7347), .dout(n7542));
  jor  g07350(.dina(n7542), .dinb(n7352), .dout(n7543));
  jand g07351(.dina(n7266), .dinb(n7259), .dout(n7544));
  jor  g07352(.dina(n7544), .dinb(n7264), .dout(n7545));
  jand g07353(.dina(n7253), .dinb(n7250), .dout(n7546));
  jor  g07354(.dina(n7546), .dinb(n7256), .dout(n7547));
  jxor g07355(.dina(n7547), .dinb(n7545), .dout(n7548));
  jxor g07356(.dina(n7548), .dinb(n7543), .dout(n7549));
  jand g07357(.dina(n7332), .dinb(n7003), .dout(n7550));
  jor  g07358(.dina(n7550), .dinb(n7335), .dout(n7551));
  jand g07359(.dina(n7314), .dinb(n7312), .dout(n7552));
  jor  g07360(.dina(n7552), .dinb(n7317), .dout(n7553));
  jxor g07361(.dina(n7553), .dinb(n7551), .dout(n7554));
  jand g07362(.dina(n7244), .dinb(n7011), .dout(n7555));
  jor  g07363(.dina(n7555), .dinb(n7247), .dout(n7556));
  jxor g07364(.dina(n7556), .dinb(n7554), .dout(n7557));
  jand g07365(.dina(\a[61] ), .dinb(\a[1] ), .dout(n7558));
  jxor g07366(.dina(n7558), .dinb(n7217), .dout(n7559));
  jand g07367(.dina(n7215), .dinb(n6984), .dout(n7560));
  jor  g07368(.dina(n7560), .dinb(n7218), .dout(n7561));
  jxor g07369(.dina(n7561), .dinb(n7559), .dout(n7562));
  jand g07370(.dina(n7224), .dinb(n7222), .dout(n7563));
  jor  g07371(.dina(n7563), .dinb(n7227), .dout(n7564));
  jxor g07372(.dina(n7564), .dinb(n7562), .dout(n7565));
  jxor g07373(.dina(n7565), .dinb(n7557), .dout(n7566));
  jxor g07374(.dina(n7566), .dinb(n7549), .dout(n7567));
  jxor g07375(.dina(n7567), .dinb(n7541), .dout(n7568));
  jxor g07376(.dina(n7568), .dinb(n7523), .dout(n7569));
  jand g07377(.dina(n7189), .dinb(n7175), .dout(n7570));
  jand g07378(.dina(n7196), .dinb(n7190), .dout(n7571));
  jor  g07379(.dina(n7571), .dinb(n7570), .dout(n7572));
  jand g07380(.dina(n7302), .dinb(n7292), .dout(n7573));
  jand g07381(.dina(n7303), .dinb(n7287), .dout(n7574));
  jor  g07382(.dina(n7574), .dinb(n7573), .dout(n7575));
  jxor g07383(.dina(n7575), .dinb(n7572), .dout(n7576));
  jnot g07384(.din(n7576), .dout(n7577));
  jand g07385(.dina(n7154), .dinb(n7147), .dout(n7578));
  jnot g07386(.din(n7578), .dout(n7579));
  jor  g07387(.dina(n7160), .dinb(n7156), .dout(n7580));
  jand g07388(.dina(n7580), .dinb(n7579), .dout(n7581));
  jxor g07389(.dina(n7581), .dinb(n7577), .dout(n7582));
  jand g07390(.dina(n7270), .dinb(n7207), .dout(n7583));
  jand g07391(.dina(n7271), .dinb(n7203), .dout(n7584));
  jor  g07392(.dina(n7584), .dinb(n7583), .dout(n7585));
  jxor g07393(.dina(n7585), .dinb(n7582), .dout(n7586));
  jxor g07394(.dina(n7586), .dinb(n7569), .dout(n7587));
  jxor g07395(.dina(n7587), .dinb(n7520), .dout(n7588));
  jxor g07396(.dina(n7588), .dinb(n7517), .dout(n7589));
  jxor g07397(.dina(n7589), .dinb(n7375), .dout(n7590));
  jand g07398(.dina(n7363), .dinb(n7123), .dout(n7591));
  jor  g07399(.dina(n7363), .dinb(n7123), .dout(n7592));
  jand g07400(.dina(n7371), .dinb(n7592), .dout(n7593));
  jor  g07401(.dina(n7593), .dinb(n7591), .dout(n7594));
  jxor g07402(.dina(n7594), .dinb(n7590), .dout(\asquared[63] ));
  jand g07403(.dina(n7587), .dinb(n7520), .dout(n7596));
  jand g07404(.dina(n7588), .dinb(n7517), .dout(n7597));
  jor  g07405(.dina(n7597), .dinb(n7596), .dout(n7598));
  jand g07406(.dina(n7423), .dinb(n7378), .dout(n7599));
  jand g07407(.dina(n7516), .dinb(n7424), .dout(n7600));
  jor  g07408(.dina(n7600), .dinb(n7599), .dout(n7601));
  jand g07409(.dina(n7514), .dinb(n7430), .dout(n7602));
  jand g07410(.dina(n7515), .dinb(n7427), .dout(n7603));
  jor  g07411(.dina(n7603), .dinb(n7602), .dout(n7604));
  jand g07412(.dina(n7565), .dinb(n7557), .dout(n7605));
  jand g07413(.dina(n7566), .dinb(n7549), .dout(n7606));
  jor  g07414(.dina(n7606), .dinb(n7605), .dout(n7607));
  jnot g07415(.din(n7607), .dout(n7608));
  jand g07416(.dina(n7534), .dinb(n7528), .dout(n7609));
  jnot g07417(.din(n7609), .dout(n7610));
  jor  g07418(.dina(n7540), .dinb(n7536), .dout(n7611));
  jand g07419(.dina(n7611), .dinb(n7610), .dout(n7612));
  jxor g07420(.dina(n7612), .dinb(n7608), .dout(n7613));
  jnot g07421(.din(n7613), .dout(n7614));
  jand g07422(.dina(n7399), .dinb(n7393), .dout(n7615));
  jnot g07423(.din(n7615), .dout(n7616));
  jor  g07424(.dina(n7405), .dinb(n7401), .dout(n7617));
  jand g07425(.dina(n7617), .dinb(n7616), .dout(n7618));
  jxor g07426(.dina(n7618), .dinb(n7614), .dout(n7619));
  jand g07427(.dina(n7553), .dinb(n7551), .dout(n7620));
  jand g07428(.dina(n7556), .dinb(n7554), .dout(n7621));
  jor  g07429(.dina(n7621), .dinb(n7620), .dout(n7622));
  jnot g07430(.din(n7380), .dout(n7623));
  jnot g07431(.din(n7382), .dout(n7624));
  jand g07432(.dina(n7624), .dinb(n7623), .dout(n7625));
  jnot g07433(.din(n7625), .dout(n7626));
  jand g07434(.dina(n7382), .dinb(n7380), .dout(n7627));
  jor  g07435(.dina(n7392), .dinb(n7627), .dout(n7628));
  jand g07436(.dina(n7628), .dinb(n7626), .dout(n7629));
  jxor g07437(.dina(n7629), .dinb(n7622), .dout(n7630));
  jand g07438(.dina(n7561), .dinb(n7559), .dout(n7631));
  jand g07439(.dina(n7564), .dinb(n7562), .dout(n7632));
  jor  g07440(.dina(n7632), .dinb(n7631), .dout(n7633));
  jxor g07441(.dina(n7633), .dinb(n7630), .dout(n7634));
  jand g07442(.dina(n7485), .dinb(n7460), .dout(n7635));
  jand g07443(.dina(n7513), .dinb(n7486), .dout(n7636));
  jor  g07444(.dina(n7636), .dinb(n7635), .dout(n7637));
  jxor g07445(.dina(n7637), .dinb(n7634), .dout(n7638));
  jand g07446(.dina(n7490), .dinb(n7487), .dout(n7639));
  jor  g07447(.dina(n7639), .dinb(n7493), .dout(n7640));
  jand g07448(.dina(n7464), .dinb(n7461), .dout(n7641));
  jor  g07449(.dina(n7641), .dinb(n7467), .dout(n7642));
  jxor g07450(.dina(n7642), .dinb(n7640), .dout(n7643));
  jand g07451(.dina(n7473), .dinb(n7470), .dout(n7644));
  jor  g07452(.dina(n7644), .dinb(n7475), .dout(n7645));
  jxor g07453(.dina(n7645), .dinb(n7643), .dout(n7646));
  jand g07454(.dina(n7386), .dinb(n7384), .dout(n7647));
  jor  g07455(.dina(n7647), .dinb(n7389), .dout(n7648));
  jand g07456(.dina(n7442), .dinb(n7255), .dout(n7649));
  jor  g07457(.dina(n7649), .dinb(n7444), .dout(n7650));
  jxor g07458(.dina(n7650), .dinb(n7648), .dout(n7651));
  jand g07459(.dina(n7453), .dinb(n7449), .dout(n7652));
  jor  g07460(.dina(n7652), .dinb(n7455), .dout(n7653));
  jxor g07461(.dina(n7653), .dinb(n7651), .dout(n7654));
  jand g07462(.dina(n7547), .dinb(n7545), .dout(n7655));
  jand g07463(.dina(n7548), .dinb(n7543), .dout(n7656));
  jor  g07464(.dina(n7656), .dinb(n7655), .dout(n7657));
  jxor g07465(.dina(n7657), .dinb(n7654), .dout(n7658));
  jxor g07466(.dina(n7658), .dinb(n7646), .dout(n7659));
  jxor g07467(.dina(n7659), .dinb(n7638), .dout(n7660));
  jxor g07468(.dina(n7660), .dinb(n7619), .dout(n7661));
  jxor g07469(.dina(n7661), .dinb(n7604), .dout(n7662));
  jxor g07470(.dina(n7662), .dinb(n7601), .dout(n7663));
  jand g07471(.dina(n7585), .dinb(n7582), .dout(n7664));
  jand g07472(.dina(n7586), .dinb(n7569), .dout(n7665));
  jor  g07473(.dina(n7665), .dinb(n7664), .dout(n7666));
  jand g07474(.dina(n7575), .dinb(n7572), .dout(n7667));
  jnot g07475(.din(n7667), .dout(n7668));
  jor  g07476(.dina(n7581), .dinb(n7577), .dout(n7669));
  jand g07477(.dina(n7669), .dinb(n7668), .dout(n7670));
  jnot g07478(.din(n7670), .dout(n7671));
  jand g07479(.dina(n7510), .dinb(n7504), .dout(n7672));
  jor  g07480(.dina(n7672), .dinb(n7508), .dout(n7673));
  jand g07481(.dina(n7498), .dinb(n7496), .dout(n7674));
  jor  g07482(.dina(n7674), .dinb(n7501), .dout(n7675));
  jand g07483(.dina(n7435), .dinb(n7431), .dout(n7676));
  jor  g07484(.dina(n7676), .dinb(n7436), .dout(n7677));
  jxor g07485(.dina(n7677), .dinb(n7675), .dout(n7678));
  jxor g07486(.dina(n7678), .dinb(n7673), .dout(n7679));
  jnot g07487(.din(n7503), .dout(n7680));
  jor  g07488(.dina(n7511), .dinb(n7680), .dout(n7681));
  jnot g07489(.din(n7495), .dout(n7682));
  jand g07490(.dina(n7511), .dinb(n7680), .dout(n7683));
  jor  g07491(.dina(n7683), .dinb(n7682), .dout(n7684));
  jand g07492(.dina(n7684), .dinb(n7681), .dout(n7685));
  jxor g07493(.dina(n7685), .dinb(n7679), .dout(n7686));
  jnot g07494(.din(n7477), .dout(n7687));
  jor  g07495(.dina(n7483), .dinb(n7687), .dout(n7688));
  jnot g07496(.din(n7469), .dout(n7689));
  jand g07497(.dina(n7483), .dinb(n7687), .dout(n7690));
  jor  g07498(.dina(n7690), .dinb(n7689), .dout(n7691));
  jand g07499(.dina(n7691), .dinb(n7688), .dout(n7692));
  jxor g07500(.dina(n7692), .dinb(n7686), .dout(n7693));
  jand g07501(.dina(n7413), .dinb(n7409), .dout(n7694));
  jand g07502(.dina(n7417), .dinb(n7414), .dout(n7695));
  jor  g07503(.dina(n7695), .dinb(n7694), .dout(n7696));
  jnot g07504(.din(n7696), .dout(n7697));
  jnot g07505(.din(n7458), .dout(n7698));
  jand g07506(.dina(n7698), .dinb(n7448), .dout(n7699));
  jnot g07507(.din(n7699), .dout(n7700));
  jand g07508(.dina(n7458), .dinb(n7447), .dout(n7701));
  jor  g07509(.dina(n7701), .dinb(n7439), .dout(n7702));
  jand g07510(.dina(n7702), .dinb(n7700), .dout(n7703));
  jxor g07511(.dina(n7703), .dinb(n7697), .dout(n7704));
  jand g07512(.dina(n7558), .dinb(n7217), .dout(n7705));
  jand g07513(.dina(\a[63] ), .dinb(\a[0] ), .dout(n7706));
  jxor g07514(.dina(n7706), .dinb(n7705), .dout(n7707));
  jnot g07515(.din(n7707), .dout(n7708));
  jand g07516(.dina(n2268), .dinb(\a[62] ), .dout(n7709));
  jnot g07517(.din(n7709), .dout(n7710));
  jand g07518(.dina(\a[62] ), .dinb(\a[1] ), .dout(n7711));
  jor  g07519(.dina(n7711), .dinb(\a[32] ), .dout(n7712));
  jand g07520(.dina(n7712), .dinb(n7710), .dout(n7713));
  jxor g07521(.dina(n7713), .dinb(n7708), .dout(n7714));
  jnot g07522(.din(n7714), .dout(n7715));
  jand g07523(.dina(\a[36] ), .dinb(\a[27] ), .dout(n7716));
  jand g07524(.dina(\a[35] ), .dinb(\a[28] ), .dout(n7717));
  jor  g07525(.dina(n7717), .dinb(n7500), .dout(n7718));
  jnot g07526(.din(n7718), .dout(n7719));
  jand g07527(.dina(\a[35] ), .dinb(\a[29] ), .dout(n7720));
  jand g07528(.dina(n7720), .dinb(n7334), .dout(n7721));
  jor  g07529(.dina(n7721), .dinb(n7719), .dout(n7722));
  jxor g07530(.dina(n7722), .dinb(n7716), .dout(n7723));
  jnot g07531(.din(n7723), .dout(n7724));
  jand g07532(.dina(\a[38] ), .dinb(\a[25] ), .dout(n7725));
  jor  g07533(.dina(n7725), .dinb(n7443), .dout(n7726));
  jand g07534(.dina(\a[38] ), .dinb(\a[26] ), .dout(n7727));
  jand g07535(.dina(n7727), .dinb(n7246), .dout(n7728));
  jnot g07536(.din(n7728), .dout(n7729));
  jand g07537(.dina(n7729), .dinb(n7726), .dout(n7730));
  jxor g07538(.dina(n7730), .dinb(n7492), .dout(n7731));
  jxor g07539(.dina(n7731), .dinb(n7724), .dout(n7732));
  jxor g07540(.dina(n7732), .dinb(n7715), .dout(n7733));
  jxor g07541(.dina(n7733), .dinb(n7704), .dout(n7734));
  jxor g07542(.dina(n7734), .dinb(n7693), .dout(n7735));
  jxor g07543(.dina(n7735), .dinb(n7671), .dout(n7736));
  jxor g07544(.dina(n7736), .dinb(n7666), .dout(n7737));
  jand g07545(.dina(n7567), .dinb(n7541), .dout(n7738));
  jand g07546(.dina(n7568), .dinb(n7523), .dout(n7739));
  jor  g07547(.dina(n7739), .dinb(n7738), .dout(n7740));
  jand g07548(.dina(n7421), .dinb(n7418), .dout(n7741));
  jand g07549(.dina(n7422), .dinb(n7406), .dout(n7742));
  jor  g07550(.dina(n7742), .dinb(n7741), .dout(n7743));
  jand g07551(.dina(\a[42] ), .dinb(\a[21] ), .dout(n7744));
  jand g07552(.dina(\a[41] ), .dinb(\a[22] ), .dout(n7745));
  jor  g07553(.dina(n7745), .dinb(n7744), .dout(n7746));
  jnot g07554(.din(n7746), .dout(n7747));
  jand g07555(.dina(\a[42] ), .dinb(\a[22] ), .dout(n7748));
  jand g07556(.dina(n7748), .dinb(n7255), .dout(n7749));
  jor  g07557(.dina(n7749), .dinb(n7747), .dout(n7750));
  jxor g07558(.dina(n7750), .dinb(n7388), .dout(n7751));
  jnot g07559(.din(n7751), .dout(n7752));
  jand g07560(.dina(n7482), .dinb(n5273), .dout(n7753));
  jor  g07561(.dina(n7753), .dinb(n7480), .dout(n7754));
  jnot g07562(.din(n7754), .dout(n7755));
  jand g07563(.dina(\a[61] ), .dinb(\a[2] ), .dout(n7756));
  jand g07564(.dina(\a[60] ), .dinb(\a[3] ), .dout(n7757));
  jand g07565(.dina(\a[59] ), .dinb(\a[4] ), .dout(n7758));
  jor  g07566(.dina(n7758), .dinb(n7757), .dout(n7759));
  jnot g07567(.din(n7759), .dout(n7760));
  jand g07568(.dina(\a[60] ), .dinb(\a[4] ), .dout(n7761));
  jand g07569(.dina(n7761), .dinb(n7384), .dout(n7762));
  jor  g07570(.dina(n7762), .dinb(n7760), .dout(n7763));
  jxor g07571(.dina(n7763), .dinb(n7756), .dout(n7764));
  jxor g07572(.dina(n7764), .dinb(n7755), .dout(n7765));
  jxor g07573(.dina(n7765), .dinb(n7752), .dout(n7766));
  jnot g07574(.din(n7466), .dout(n7767));
  jand g07575(.dina(\a[55] ), .dinb(\a[8] ), .dout(n7768));
  jand g07576(.dina(\a[44] ), .dinb(\a[19] ), .dout(n7769));
  jor  g07577(.dina(n7769), .dinb(n7768), .dout(n7770));
  jand g07578(.dina(\a[55] ), .dinb(\a[19] ), .dout(n7771));
  jand g07579(.dina(n7771), .dinb(n5255), .dout(n7772));
  jnot g07580(.din(n7772), .dout(n7773));
  jand g07581(.dina(n7773), .dinb(n7770), .dout(n7774));
  jxor g07582(.dina(n7774), .dinb(n7767), .dout(n7775));
  jand g07583(.dina(\a[40] ), .dinb(\a[23] ), .dout(n7776));
  jnot g07584(.din(n7776), .dout(n7777));
  jand g07585(.dina(\a[57] ), .dinb(\a[6] ), .dout(n7778));
  jand g07586(.dina(\a[43] ), .dinb(\a[20] ), .dout(n7779));
  jxor g07587(.dina(n7779), .dinb(n7778), .dout(n7780));
  jxor g07588(.dina(n7780), .dinb(n7777), .dout(n7781));
  jnot g07589(.din(n7226), .dout(n7782));
  jand g07590(.dina(\a[32] ), .dinb(\a[31] ), .dout(n7783));
  jand g07591(.dina(\a[33] ), .dinb(\a[30] ), .dout(n7784));
  jxor g07592(.dina(n7784), .dinb(n7783), .dout(n7785));
  jxor g07593(.dina(n7785), .dinb(n7782), .dout(n7786));
  jnot g07594(.din(n7786), .dout(n7787));
  jxor g07595(.dina(n7787), .dinb(n7781), .dout(n7788));
  jxor g07596(.dina(n7788), .dinb(n7775), .dout(n7789));
  jxor g07597(.dina(n7789), .dinb(n7766), .dout(n7790));
  jand g07598(.dina(\a[53] ), .dinb(\a[10] ), .dout(n7791));
  jand g07599(.dina(\a[52] ), .dinb(\a[11] ), .dout(n7792));
  jand g07600(.dina(\a[47] ), .dinb(\a[16] ), .dout(n7793));
  jor  g07601(.dina(n7793), .dinb(n7792), .dout(n7794));
  jnot g07602(.din(n7794), .dout(n7795));
  jand g07603(.dina(\a[52] ), .dinb(\a[16] ), .dout(n7796));
  jand g07604(.dina(n7796), .dinb(n6654), .dout(n7797));
  jor  g07605(.dina(n7797), .dinb(n7795), .dout(n7798));
  jxor g07606(.dina(n7798), .dinb(n7791), .dout(n7799));
  jnot g07607(.din(n7799), .dout(n7800));
  jand g07608(.dina(\a[45] ), .dinb(\a[18] ), .dout(n7801));
  jand g07609(.dina(\a[54] ), .dinb(\a[9] ), .dout(n7802));
  jor  g07610(.dina(n7802), .dinb(n4872), .dout(n7803));
  jand g07611(.dina(\a[54] ), .dinb(\a[17] ), .dout(n7804));
  jand g07612(.dina(n7804), .dinb(n6011), .dout(n7805));
  jnot g07613(.din(n7805), .dout(n7806));
  jand g07614(.dina(n7806), .dinb(n7803), .dout(n7807));
  jxor g07615(.dina(n7807), .dinb(n7801), .dout(n7808));
  jxor g07616(.dina(n7808), .dinb(n7800), .dout(n7809));
  jnot g07617(.din(n7809), .dout(n7810));
  jand g07618(.dina(\a[50] ), .dinb(\a[13] ), .dout(n7811));
  jand g07619(.dina(\a[51] ), .dinb(\a[12] ), .dout(n7812));
  jor  g07620(.dina(n7812), .dinb(n7811), .dout(n7813));
  jnot g07621(.din(n7813), .dout(n7814));
  jand g07622(.dina(\a[51] ), .dinb(\a[13] ), .dout(n7815));
  jand g07623(.dina(n7815), .dinb(n7470), .dout(n7816));
  jor  g07624(.dina(n7816), .dinb(n7814), .dout(n7817));
  jxor g07625(.dina(n7817), .dinb(n6047), .dout(n7818));
  jxor g07626(.dina(n7818), .dinb(n7810), .dout(n7819));
  jxor g07627(.dina(n7819), .dinb(n7790), .dout(n7820));
  jxor g07628(.dina(n7820), .dinb(n7743), .dout(n7821));
  jxor g07629(.dina(n7821), .dinb(n7740), .dout(n7822));
  jxor g07630(.dina(n7822), .dinb(n7737), .dout(n7823));
  jxor g07631(.dina(n7823), .dinb(n7663), .dout(n7824));
  jxor g07632(.dina(n7824), .dinb(n7598), .dout(n7825));
  jand g07633(.dina(n7589), .dinb(n7375), .dout(n7826));
  jor  g07634(.dina(n7589), .dinb(n7375), .dout(n7827));
  jand g07635(.dina(n7594), .dinb(n7827), .dout(n7828));
  jor  g07636(.dina(n7828), .dinb(n7826), .dout(n7829));
  jxor g07637(.dina(n7829), .dinb(n7825), .dout(\asquared[64] ));
  jand g07638(.dina(n7660), .dinb(n7619), .dout(n7831));
  jand g07639(.dina(n7661), .dinb(n7604), .dout(n7832));
  jor  g07640(.dina(n7832), .dinb(n7831), .dout(n7833));
  jand g07641(.dina(n7730), .dinb(n7492), .dout(n7834));
  jor  g07642(.dina(n7834), .dinb(n7728), .dout(n7835));
  jand g07643(.dina(n7813), .dinb(n6047), .dout(n7836));
  jor  g07644(.dina(n7836), .dinb(n7816), .dout(n7837));
  jxor g07645(.dina(n7837), .dinb(n7835), .dout(n7838));
  jand g07646(.dina(n7794), .dinb(n7791), .dout(n7839));
  jor  g07647(.dina(n7839), .dinb(n7797), .dout(n7840));
  jxor g07648(.dina(n7840), .dinb(n7838), .dout(n7841));
  jnot g07649(.din(n7841), .dout(n7842));
  jnot g07650(.din(n7781), .dout(n7843));
  jand g07651(.dina(n7787), .dinb(n7843), .dout(n7844));
  jnot g07652(.din(n7844), .dout(n7845));
  jand g07653(.dina(n7786), .dinb(n7781), .dout(n7846));
  jor  g07654(.dina(n7846), .dinb(n7775), .dout(n7847));
  jand g07655(.dina(n7847), .dinb(n7845), .dout(n7848));
  jxor g07656(.dina(n7848), .dinb(n7842), .dout(n7849));
  jnot g07657(.din(n7849), .dout(n7850));
  jand g07658(.dina(n7808), .dinb(n7800), .dout(n7851));
  jnot g07659(.din(n7851), .dout(n7852));
  jor  g07660(.dina(n7818), .dinb(n7810), .dout(n7853));
  jand g07661(.dina(n7853), .dinb(n7852), .dout(n7854));
  jxor g07662(.dina(n7854), .dinb(n7850), .dout(n7855));
  jnot g07663(.din(n7855), .dout(n7856));
  jor  g07664(.dina(n7612), .dinb(n7608), .dout(n7857));
  jor  g07665(.dina(n7618), .dinb(n7614), .dout(n7858));
  jand g07666(.dina(n7858), .dinb(n7857), .dout(n7859));
  jxor g07667(.dina(n7859), .dinb(n7856), .dout(n7860));
  jand g07668(.dina(n7629), .dinb(n7622), .dout(n7861));
  jand g07669(.dina(n7633), .dinb(n7630), .dout(n7862));
  jor  g07670(.dina(n7862), .dinb(n7861), .dout(n7863));
  jor  g07671(.dina(n7764), .dinb(n7755), .dout(n7864));
  jand g07672(.dina(n7765), .dinb(n7752), .dout(n7865));
  jnot g07673(.din(n7865), .dout(n7866));
  jand g07674(.dina(n7866), .dinb(n7864), .dout(n7867));
  jnot g07675(.din(n7867), .dout(n7868));
  jxor g07676(.dina(n7868), .dinb(n7863), .dout(n7869));
  jnot g07677(.din(n7783), .dout(n7870));
  jnot g07678(.din(n7784), .dout(n7871));
  jand g07679(.dina(n7871), .dinb(n7870), .dout(n7872));
  jnot g07680(.din(n7872), .dout(n7873));
  jand g07681(.dina(n7784), .dinb(n7783), .dout(n7874));
  jor  g07682(.dina(n7874), .dinb(n7226), .dout(n7875));
  jand g07683(.dina(n7875), .dinb(n7873), .dout(n7876));
  jand g07684(.dina(\a[63] ), .dinb(\a[1] ), .dout(n7877));
  jor  g07685(.dina(n7877), .dinb(n7709), .dout(n7878));
  jand g07686(.dina(n7709), .dinb(\a[63] ), .dout(n7879));
  jnot g07687(.din(n7879), .dout(n7880));
  jand g07688(.dina(n7880), .dinb(n7878), .dout(n7881));
  jxor g07689(.dina(n7881), .dinb(n7876), .dout(n7882));
  jand g07690(.dina(\a[53] ), .dinb(\a[11] ), .dout(n7883));
  jand g07691(.dina(\a[52] ), .dinb(\a[12] ), .dout(n7884));
  jor  g07692(.dina(n7884), .dinb(n7883), .dout(n7885));
  jnot g07693(.din(n7885), .dout(n7886));
  jand g07694(.dina(\a[53] ), .dinb(\a[12] ), .dout(n7887));
  jand g07695(.dina(n7887), .dinb(n7792), .dout(n7888));
  jor  g07696(.dina(n7888), .dinb(n7886), .dout(n7889));
  jxor g07697(.dina(n7889), .dinb(n7815), .dout(n7890));
  jand g07698(.dina(\a[55] ), .dinb(\a[9] ), .dout(n7891));
  jnot g07699(.din(n7891), .dout(n7892));
  jand g07700(.dina(\a[54] ), .dinb(\a[10] ), .dout(n7893));
  jxor g07701(.dina(n7893), .dinb(n6845), .dout(n7894));
  jxor g07702(.dina(n7894), .dinb(n7892), .dout(n7895));
  jxor g07703(.dina(n7895), .dinb(n7890), .dout(n7896));
  jxor g07704(.dina(n7896), .dinb(n7882), .dout(n7897));
  jxor g07705(.dina(n7897), .dinb(n7869), .dout(n7898));
  jxor g07706(.dina(n7898), .dinb(n7860), .dout(n7899));
  jxor g07707(.dina(n7899), .dinb(n7833), .dout(n7900));
  jand g07708(.dina(n7637), .dinb(n7634), .dout(n7901));
  jand g07709(.dina(n7659), .dinb(n7638), .dout(n7902));
  jor  g07710(.dina(n7902), .dinb(n7901), .dout(n7903));
  jand g07711(.dina(\a[61] ), .dinb(\a[3] ), .dout(n7904));
  jor  g07712(.dina(n7904), .dinb(n7761), .dout(n7905));
  jnot g07713(.din(n7905), .dout(n7906));
  jand g07714(.dina(\a[61] ), .dinb(\a[4] ), .dout(n7907));
  jand g07715(.dina(n7907), .dinb(n7757), .dout(n7908));
  jor  g07716(.dina(n7908), .dinb(n7906), .dout(n7909));
  jxor g07717(.dina(n7909), .dinb(n7454), .dout(n7910));
  jnot g07718(.din(n7910), .dout(n7911));
  jand g07719(.dina(\a[46] ), .dinb(\a[18] ), .dout(n7912));
  jand g07720(.dina(\a[45] ), .dinb(\a[19] ), .dout(n7913));
  jor  g07721(.dina(n7913), .dinb(n7912), .dout(n7914));
  jnot g07722(.din(n7914), .dout(n7915));
  jand g07723(.dina(\a[46] ), .dinb(\a[19] ), .dout(n7916));
  jand g07724(.dina(n7916), .dinb(n7801), .dout(n7917));
  jor  g07725(.dina(n7917), .dinb(n7915), .dout(n7918));
  jxor g07726(.dina(n7918), .dinb(n7263), .dout(n7919));
  jnot g07727(.din(n7919), .dout(n7920));
  jor  g07728(.dina(n7706), .dinb(n7705), .dout(n7921));
  jand g07729(.dina(n7706), .dinb(n7705), .dout(n7922));
  jor  g07730(.dina(n7713), .dinb(n7922), .dout(n7923));
  jand g07731(.dina(n7923), .dinb(n7921), .dout(n7924));
  jxor g07732(.dina(n7924), .dinb(n7920), .dout(n7925));
  jxor g07733(.dina(n7925), .dinb(n7911), .dout(n7926));
  jand g07734(.dina(\a[50] ), .dinb(\a[14] ), .dout(n7927));
  jand g07735(.dina(\a[33] ), .dinb(\a[31] ), .dout(n7928));
  jand g07736(.dina(\a[34] ), .dinb(\a[30] ), .dout(n7929));
  jor  g07737(.dina(n7929), .dinb(n7928), .dout(n7930));
  jnot g07738(.din(n7930), .dout(n7931));
  jand g07739(.dina(\a[34] ), .dinb(\a[31] ), .dout(n7932));
  jand g07740(.dina(n7932), .dinb(n7784), .dout(n7933));
  jor  g07741(.dina(n7933), .dinb(n7931), .dout(n7934));
  jxor g07742(.dina(n7934), .dinb(n7927), .dout(n7935));
  jand g07743(.dina(\a[37] ), .dinb(\a[27] ), .dout(n7936));
  jand g07744(.dina(\a[36] ), .dinb(\a[28] ), .dout(n7937));
  jor  g07745(.dina(n7937), .dinb(n7720), .dout(n7938));
  jnot g07746(.din(n7938), .dout(n7939));
  jand g07747(.dina(\a[36] ), .dinb(\a[29] ), .dout(n7940));
  jand g07748(.dina(n7940), .dinb(n7717), .dout(n7941));
  jor  g07749(.dina(n7941), .dinb(n7939), .dout(n7942));
  jxor g07750(.dina(n7942), .dinb(n7936), .dout(n7943));
  jand g07751(.dina(\a[56] ), .dinb(\a[8] ), .dout(n7944));
  jor  g07752(.dina(n7944), .dinb(n5465), .dout(n7945));
  jand g07753(.dina(\a[56] ), .dinb(\a[16] ), .dout(n7946));
  jand g07754(.dina(n7946), .dinb(n5930), .dout(n7947));
  jnot g07755(.din(n7947), .dout(n7948));
  jand g07756(.dina(n7948), .dinb(n7945), .dout(n7949));
  jxor g07757(.dina(n7949), .dinb(n7727), .dout(n7950));
  jxor g07758(.dina(n7950), .dinb(n7943), .dout(n7951));
  jxor g07759(.dina(n7951), .dinb(n7935), .dout(n7952));
  jxor g07760(.dina(n7952), .dinb(n7926), .dout(n7953));
  jand g07761(.dina(\a[41] ), .dinb(\a[23] ), .dout(n7954));
  jand g07762(.dina(\a[40] ), .dinb(\a[24] ), .dout(n7955));
  jand g07763(.dina(\a[39] ), .dinb(\a[25] ), .dout(n7956));
  jor  g07764(.dina(n7956), .dinb(n7955), .dout(n7957));
  jnot g07765(.din(n7957), .dout(n7958));
  jand g07766(.dina(\a[40] ), .dinb(\a[25] ), .dout(n7959));
  jand g07767(.dina(n7959), .dinb(n7492), .dout(n7960));
  jor  g07768(.dina(n7960), .dinb(n7958), .dout(n7961));
  jxor g07769(.dina(n7961), .dinb(n7954), .dout(n7962));
  jand g07770(.dina(\a[44] ), .dinb(\a[20] ), .dout(n7963));
  jand g07771(.dina(\a[43] ), .dinb(\a[21] ), .dout(n7964));
  jor  g07772(.dina(n7964), .dinb(n7748), .dout(n7965));
  jnot g07773(.din(n7965), .dout(n7966));
  jand g07774(.dina(\a[43] ), .dinb(\a[22] ), .dout(n7967));
  jand g07775(.dina(n7967), .dinb(n7744), .dout(n7968));
  jor  g07776(.dina(n7968), .dinb(n7966), .dout(n7969));
  jxor g07777(.dina(n7969), .dinb(n7963), .dout(n7970));
  jand g07778(.dina(\a[58] ), .dinb(\a[6] ), .dout(n7971));
  jand g07779(.dina(\a[47] ), .dinb(\a[17] ), .dout(n7972));
  jand g07780(.dina(\a[57] ), .dinb(\a[7] ), .dout(n7973));
  jor  g07781(.dina(n7973), .dinb(n7972), .dout(n7974));
  jand g07782(.dina(\a[57] ), .dinb(\a[17] ), .dout(n7975));
  jand g07783(.dina(n7975), .dinb(n5749), .dout(n7976));
  jnot g07784(.din(n7976), .dout(n7977));
  jand g07785(.dina(n7977), .dinb(n7974), .dout(n7978));
  jxor g07786(.dina(n7978), .dinb(n7971), .dout(n7979));
  jxor g07787(.dina(n7979), .dinb(n7970), .dout(n7980));
  jxor g07788(.dina(n7980), .dinb(n7962), .dout(n7981));
  jxor g07789(.dina(n7981), .dinb(n7953), .dout(n7982));
  jxor g07790(.dina(n7982), .dinb(n7903), .dout(n7983));
  jand g07791(.dina(n7642), .dinb(n7640), .dout(n7984));
  jand g07792(.dina(n7645), .dinb(n7643), .dout(n7985));
  jor  g07793(.dina(n7985), .dinb(n7984), .dout(n7986));
  jand g07794(.dina(n7677), .dinb(n7675), .dout(n7987));
  jand g07795(.dina(n7678), .dinb(n7673), .dout(n7988));
  jor  g07796(.dina(n7988), .dinb(n7987), .dout(n7989));
  jxor g07797(.dina(n7989), .dinb(n7986), .dout(n7990));
  jand g07798(.dina(n7650), .dinb(n7648), .dout(n7991));
  jand g07799(.dina(n7653), .dinb(n7651), .dout(n7992));
  jor  g07800(.dina(n7992), .dinb(n7991), .dout(n7993));
  jxor g07801(.dina(n7993), .dinb(n7990), .dout(n7994));
  jand g07802(.dina(n7685), .dinb(n7679), .dout(n7995));
  jand g07803(.dina(n7692), .dinb(n7686), .dout(n7996));
  jor  g07804(.dina(n7996), .dinb(n7995), .dout(n7997));
  jand g07805(.dina(n7657), .dinb(n7654), .dout(n7998));
  jand g07806(.dina(n7658), .dinb(n7646), .dout(n7999));
  jor  g07807(.dina(n7999), .dinb(n7998), .dout(n8000));
  jxor g07808(.dina(n8000), .dinb(n7997), .dout(n8001));
  jxor g07809(.dina(n8001), .dinb(n7994), .dout(n8002));
  jxor g07810(.dina(n8002), .dinb(n7983), .dout(n8003));
  jxor g07811(.dina(n8003), .dinb(n7900), .dout(n8004));
  jand g07812(.dina(n7736), .dinb(n7666), .dout(n8005));
  jand g07813(.dina(n7822), .dinb(n7737), .dout(n8006));
  jor  g07814(.dina(n8006), .dinb(n8005), .dout(n8007));
  jand g07815(.dina(n7820), .dinb(n7743), .dout(n8008));
  jand g07816(.dina(n7821), .dinb(n7740), .dout(n8009));
  jor  g07817(.dina(n8009), .dinb(n8008), .dout(n8010));
  jand g07818(.dina(n7734), .dinb(n7693), .dout(n8011));
  jand g07819(.dina(n7735), .dinb(n7671), .dout(n8012));
  jor  g07820(.dina(n8012), .dinb(n8011), .dout(n8013));
  jand g07821(.dina(n7789), .dinb(n7766), .dout(n8014));
  jand g07822(.dina(n7819), .dinb(n7790), .dout(n8015));
  jor  g07823(.dina(n8015), .dinb(n8014), .dout(n8016));
  jnot g07824(.din(n8016), .dout(n8017));
  jor  g07825(.dina(n7703), .dinb(n7697), .dout(n8018));
  jand g07826(.dina(n7733), .dinb(n7704), .dout(n8019));
  jnot g07827(.din(n8019), .dout(n8020));
  jand g07828(.dina(n8020), .dinb(n8018), .dout(n8021));
  jxor g07829(.dina(n8021), .dinb(n8017), .dout(n8022));
  jand g07830(.dina(n7731), .dinb(n7724), .dout(n8023));
  jand g07831(.dina(n7732), .dinb(n7715), .dout(n8024));
  jor  g07832(.dina(n8024), .dinb(n8023), .dout(n8025));
  jand g07833(.dina(n7807), .dinb(n7801), .dout(n8026));
  jor  g07834(.dina(n8026), .dinb(n7805), .dout(n8027));
  jnot g07835(.din(n7778), .dout(n8028));
  jnot g07836(.din(n7779), .dout(n8029));
  jand g07837(.dina(n8029), .dinb(n8028), .dout(n8030));
  jnot g07838(.din(n8030), .dout(n8031));
  jand g07839(.dina(n7779), .dinb(n7778), .dout(n8032));
  jor  g07840(.dina(n8032), .dinb(n7776), .dout(n8033));
  jand g07841(.dina(n8033), .dinb(n8031), .dout(n8034));
  jxor g07842(.dina(n8034), .dinb(n8027), .dout(n8035));
  jand g07843(.dina(n7718), .dinb(n7716), .dout(n8036));
  jor  g07844(.dina(n8036), .dinb(n7721), .dout(n8037));
  jxor g07845(.dina(n8037), .dinb(n8035), .dout(n8038));
  jand g07846(.dina(n7746), .dinb(n7388), .dout(n8039));
  jor  g07847(.dina(n8039), .dinb(n7749), .dout(n8040));
  jand g07848(.dina(n7759), .dinb(n7756), .dout(n8041));
  jor  g07849(.dina(n8041), .dinb(n7762), .dout(n8042));
  jxor g07850(.dina(n8042), .dinb(n8040), .dout(n8043));
  jand g07851(.dina(n7770), .dinb(n7466), .dout(n8044));
  jor  g07852(.dina(n8044), .dinb(n7772), .dout(n8045));
  jxor g07853(.dina(n8045), .dinb(n8043), .dout(n8046));
  jxor g07854(.dina(n8046), .dinb(n8038), .dout(n8047));
  jxor g07855(.dina(n8047), .dinb(n8025), .dout(n8048));
  jxor g07856(.dina(n8048), .dinb(n8022), .dout(n8049));
  jxor g07857(.dina(n8049), .dinb(n8013), .dout(n8050));
  jxor g07858(.dina(n8050), .dinb(n8010), .dout(n8051));
  jxor g07859(.dina(n8051), .dinb(n8007), .dout(n8052));
  jxor g07860(.dina(n8052), .dinb(n8004), .dout(n8053));
  jand g07861(.dina(n7662), .dinb(n7601), .dout(n8054));
  jand g07862(.dina(n7823), .dinb(n7663), .dout(n8055));
  jor  g07863(.dina(n8055), .dinb(n8054), .dout(n8056));
  jxor g07864(.dina(n8056), .dinb(n8053), .dout(n8057));
  jand g07865(.dina(n7824), .dinb(n7598), .dout(n8058));
  jnot g07866(.din(n7598), .dout(n8059));
  jnot g07867(.din(n7824), .dout(n8060));
  jand g07868(.dina(n8060), .dinb(n8059), .dout(n8061));
  jnot g07869(.din(n8061), .dout(n8062));
  jand g07870(.dina(n7829), .dinb(n8062), .dout(n8063));
  jor  g07871(.dina(n8063), .dinb(n8058), .dout(n8064));
  jxor g07872(.dina(n8064), .dinb(n8057), .dout(\asquared[65] ));
  jand g07873(.dina(n8051), .dinb(n8007), .dout(n8066));
  jand g07874(.dina(n8052), .dinb(n8004), .dout(n8067));
  jor  g07875(.dina(n8067), .dinb(n8066), .dout(n8068));
  jand g07876(.dina(n7899), .dinb(n7833), .dout(n8069));
  jand g07877(.dina(n8003), .dinb(n7900), .dout(n8070));
  jor  g07878(.dina(n8070), .dinb(n8069), .dout(n8071));
  jand g07879(.dina(n7982), .dinb(n7903), .dout(n8072));
  jand g07880(.dina(n8002), .dinb(n7983), .dout(n8073));
  jor  g07881(.dina(n8073), .dinb(n8072), .dout(n8074));
  jor  g07882(.dina(n7859), .dinb(n7856), .dout(n8075));
  jand g07883(.dina(n7898), .dinb(n7860), .dout(n8076));
  jnot g07884(.din(n8076), .dout(n8077));
  jand g07885(.dina(n8077), .dinb(n8075), .dout(n8078));
  jnot g07886(.din(n8078), .dout(n8079));
  jand g07887(.dina(n7952), .dinb(n7926), .dout(n8080));
  jand g07888(.dina(n7981), .dinb(n7953), .dout(n8081));
  jor  g07889(.dina(n8081), .dinb(n8080), .dout(n8082));
  jand g07890(.dina(n7868), .dinb(n7863), .dout(n8083));
  jand g07891(.dina(n7897), .dinb(n7869), .dout(n8084));
  jor  g07892(.dina(n8084), .dinb(n8083), .dout(n8085));
  jxor g07893(.dina(n8085), .dinb(n8082), .dout(n8086));
  jor  g07894(.dina(n7895), .dinb(n7890), .dout(n8087));
  jand g07895(.dina(n7896), .dinb(n7882), .dout(n8088));
  jnot g07896(.din(n8088), .dout(n8089));
  jand g07897(.dina(n8089), .dinb(n8087), .dout(n8090));
  jnot g07898(.din(n8090), .dout(n8091));
  jand g07899(.dina(n7978), .dinb(n7971), .dout(n8092));
  jor  g07900(.dina(n8092), .dinb(n7976), .dout(n8093));
  jand g07901(.dina(n7957), .dinb(n7954), .dout(n8094));
  jor  g07902(.dina(n8094), .dinb(n7960), .dout(n8095));
  jand g07903(.dina(n7893), .dinb(n6845), .dout(n8096));
  jnot g07904(.din(n8096), .dout(n8097));
  jnot g07905(.din(n6845), .dout(n8098));
  jnot g07906(.din(n7893), .dout(n8099));
  jand g07907(.dina(n8099), .dinb(n8098), .dout(n8100));
  jor  g07908(.dina(n8100), .dinb(n7892), .dout(n8101));
  jand g07909(.dina(n8101), .dinb(n8097), .dout(n8102));
  jnot g07910(.din(n8102), .dout(n8103));
  jxor g07911(.dina(n8103), .dinb(n8095), .dout(n8104));
  jxor g07912(.dina(n8104), .dinb(n8093), .dout(n8105));
  jand g07913(.dina(n7949), .dinb(n7727), .dout(n8106));
  jor  g07914(.dina(n8106), .dinb(n7947), .dout(n8107));
  jand g07915(.dina(n7905), .dinb(n7454), .dout(n8108));
  jor  g07916(.dina(n8108), .dinb(n7908), .dout(n8109));
  jand g07917(.dina(n7914), .dinb(n7263), .dout(n8110));
  jor  g07918(.dina(n8110), .dinb(n7917), .dout(n8111));
  jxor g07919(.dina(n8111), .dinb(n8109), .dout(n8112));
  jxor g07920(.dina(n8112), .dinb(n8107), .dout(n8113));
  jxor g07921(.dina(n8113), .dinb(n8105), .dout(n8114));
  jxor g07922(.dina(n8114), .dinb(n8091), .dout(n8115));
  jxor g07923(.dina(n8115), .dinb(n8086), .dout(n8116));
  jxor g07924(.dina(n8116), .dinb(n8079), .dout(n8117));
  jxor g07925(.dina(n8117), .dinb(n8074), .dout(n8118));
  jxor g07926(.dina(n8118), .dinb(n8071), .dout(n8119));
  jand g07927(.dina(n8049), .dinb(n8013), .dout(n8120));
  jand g07928(.dina(n8050), .dinb(n8010), .dout(n8121));
  jor  g07929(.dina(n8121), .dinb(n8120), .dout(n8122));
  jand g07930(.dina(n7965), .dinb(n7963), .dout(n8123));
  jor  g07931(.dina(n8123), .dinb(n7968), .dout(n8124));
  jand g07932(.dina(n7938), .dinb(n7936), .dout(n8125));
  jor  g07933(.dina(n8125), .dinb(n7941), .dout(n8126));
  jxor g07934(.dina(n8126), .dinb(n8124), .dout(n8127));
  jand g07935(.dina(n7885), .dinb(n7815), .dout(n8128));
  jor  g07936(.dina(n8128), .dinb(n7888), .dout(n8129));
  jxor g07937(.dina(n8129), .dinb(n8127), .dout(n8130));
  jnot g07938(.din(n7943), .dout(n8131));
  jor  g07939(.dina(n7950), .dinb(n8131), .dout(n8132));
  jnot g07940(.din(n7935), .dout(n8133));
  jand g07941(.dina(n7950), .dinb(n8131), .dout(n8134));
  jor  g07942(.dina(n8134), .dinb(n8133), .dout(n8135));
  jand g07943(.dina(n8135), .dinb(n8132), .dout(n8136));
  jxor g07944(.dina(n8136), .dinb(n8130), .dout(n8137));
  jnot g07945(.din(n7970), .dout(n8138));
  jor  g07946(.dina(n7979), .dinb(n8138), .dout(n8139));
  jnot g07947(.din(n7962), .dout(n8140));
  jand g07948(.dina(n7979), .dinb(n8138), .dout(n8141));
  jor  g07949(.dina(n8141), .dinb(n8140), .dout(n8142));
  jand g07950(.dina(n8142), .dinb(n8139), .dout(n8143));
  jxor g07951(.dina(n8143), .dinb(n8137), .dout(n8144));
  jand g07952(.dina(n8000), .dinb(n7997), .dout(n8145));
  jand g07953(.dina(n8001), .dinb(n7994), .dout(n8146));
  jor  g07954(.dina(n8146), .dinb(n8145), .dout(n8147));
  jxor g07955(.dina(n8147), .dinb(n8144), .dout(n8148));
  jand g07956(.dina(n7989), .dinb(n7986), .dout(n8149));
  jand g07957(.dina(n7993), .dinb(n7990), .dout(n8150));
  jor  g07958(.dina(n8150), .dinb(n8149), .dout(n8151));
  jand g07959(.dina(n7924), .dinb(n7920), .dout(n8152));
  jand g07960(.dina(n7925), .dinb(n7911), .dout(n8153));
  jor  g07961(.dina(n8153), .dinb(n8152), .dout(n8154));
  jxor g07962(.dina(n8154), .dinb(n8151), .dout(n8155));
  jand g07963(.dina(\a[63] ), .dinb(\a[2] ), .dout(n8156));
  jor  g07964(.dina(n8156), .dinb(n7907), .dout(n8157));
  jand g07965(.dina(\a[63] ), .dinb(\a[4] ), .dout(n8158));
  jand g07966(.dina(n8158), .dinb(n7756), .dout(n8159));
  jnot g07967(.din(n8159), .dout(n8160));
  jand g07968(.dina(n8160), .dinb(n8157), .dout(n8161));
  jand g07969(.dina(n7930), .dinb(n7927), .dout(n8162));
  jor  g07970(.dina(n8162), .dinb(n7933), .dout(n8163));
  jxor g07971(.dina(n8163), .dinb(n8161), .dout(n8164));
  jand g07972(.dina(\a[51] ), .dinb(\a[14] ), .dout(n8165));
  jand g07973(.dina(\a[50] ), .dinb(\a[15] ), .dout(n8166));
  jor  g07974(.dina(n8166), .dinb(n8165), .dout(n8167));
  jnot g07975(.din(n8167), .dout(n8168));
  jand g07976(.dina(n7927), .dinb(n7235), .dout(n8169));
  jor  g07977(.dina(n8169), .dinb(n8168), .dout(n8170));
  jxor g07978(.dina(n8170), .dinb(n6419), .dout(n8171));
  jnot g07979(.din(n7887), .dout(n8172));
  jand g07980(.dina(\a[52] ), .dinb(\a[13] ), .dout(n8173));
  jand g07981(.dina(\a[47] ), .dinb(\a[18] ), .dout(n8174));
  jxor g07982(.dina(n8174), .dinb(n8173), .dout(n8175));
  jxor g07983(.dina(n8175), .dinb(n8172), .dout(n8176));
  jxor g07984(.dina(n8176), .dinb(n8171), .dout(n8177));
  jxor g07985(.dina(n8177), .dinb(n8164), .dout(n8178));
  jxor g07986(.dina(n8178), .dinb(n8155), .dout(n8179));
  jxor g07987(.dina(n8179), .dinb(n8148), .dout(n8180));
  jxor g07988(.dina(n8180), .dinb(n8122), .dout(n8181));
  jand g07989(.dina(n7837), .dinb(n7835), .dout(n8182));
  jand g07990(.dina(n7840), .dinb(n7838), .dout(n8183));
  jor  g07991(.dina(n8183), .dinb(n8182), .dout(n8184));
  jand g07992(.dina(n8034), .dinb(n8027), .dout(n8185));
  jand g07993(.dina(n8037), .dinb(n8035), .dout(n8186));
  jor  g07994(.dina(n8186), .dinb(n8185), .dout(n8187));
  jxor g07995(.dina(n8187), .dinb(n8184), .dout(n8188));
  jand g07996(.dina(n8042), .dinb(n8040), .dout(n8189));
  jand g07997(.dina(n8045), .dinb(n8043), .dout(n8190));
  jor  g07998(.dina(n8190), .dinb(n8189), .dout(n8191));
  jxor g07999(.dina(n8191), .dinb(n8188), .dout(n8192));
  jand g08000(.dina(n8046), .dinb(n8038), .dout(n8193));
  jand g08001(.dina(n8047), .dinb(n8025), .dout(n8194));
  jor  g08002(.dina(n8194), .dinb(n8193), .dout(n8195));
  jnot g08003(.din(n8195), .dout(n8196));
  jor  g08004(.dina(n7848), .dinb(n7842), .dout(n8197));
  jor  g08005(.dina(n7854), .dinb(n7850), .dout(n8198));
  jand g08006(.dina(n8198), .dinb(n8197), .dout(n8199));
  jxor g08007(.dina(n8199), .dinb(n8196), .dout(n8200));
  jxor g08008(.dina(n8200), .dinb(n8192), .dout(n8201));
  jor  g08009(.dina(n8021), .dinb(n8017), .dout(n8202));
  jand g08010(.dina(n8048), .dinb(n8022), .dout(n8203));
  jnot g08011(.din(n8203), .dout(n8204));
  jand g08012(.dina(n8204), .dinb(n8202), .dout(n8205));
  jnot g08013(.din(n8205), .dout(n8206));
  jand g08014(.dina(\a[60] ), .dinb(\a[5] ), .dout(n8207));
  jand g08015(.dina(\a[59] ), .dinb(\a[6] ), .dout(n8208));
  jand g08016(.dina(\a[58] ), .dinb(\a[7] ), .dout(n8209));
  jor  g08017(.dina(n8209), .dinb(n8208), .dout(n8210));
  jnot g08018(.din(n8210), .dout(n8211));
  jand g08019(.dina(\a[59] ), .dinb(\a[7] ), .dout(n8212));
  jand g08020(.dina(n8212), .dinb(n7971), .dout(n8213));
  jor  g08021(.dina(n8213), .dinb(n8211), .dout(n8214));
  jxor g08022(.dina(n8214), .dinb(n8207), .dout(n8215));
  jnot g08023(.din(n8215), .dout(n8216));
  jand g08024(.dina(\a[57] ), .dinb(\a[8] ), .dout(n8217));
  jand g08025(.dina(\a[44] ), .dinb(\a[21] ), .dout(n8218));
  jor  g08026(.dina(n8218), .dinb(n7967), .dout(n8219));
  jnot g08027(.din(n8219), .dout(n8220));
  jand g08028(.dina(\a[44] ), .dinb(\a[22] ), .dout(n8221));
  jand g08029(.dina(n8221), .dinb(n7964), .dout(n8222));
  jor  g08030(.dina(n8222), .dinb(n8220), .dout(n8223));
  jxor g08031(.dina(n8223), .dinb(n8217), .dout(n8224));
  jnot g08032(.din(n8224), .dout(n8225));
  jand g08033(.dina(n7881), .dinb(n7876), .dout(n8226));
  jor  g08034(.dina(n8226), .dinb(n7879), .dout(n8227));
  jxor g08035(.dina(n8227), .dinb(n8225), .dout(n8228));
  jxor g08036(.dina(n8228), .dinb(n8216), .dout(n8229));
  jand g08037(.dina(\a[48] ), .dinb(\a[17] ), .dout(n8230));
  jnot g08038(.din(\a[33] ), .dout(n8231));
  jand g08039(.dina(\a[62] ), .dinb(\a[3] ), .dout(n8232));
  jxor g08040(.dina(n8232), .dinb(n8231), .dout(n8233));
  jxor g08041(.dina(n8233), .dinb(n8230), .dout(n8234));
  jnot g08042(.din(n8234), .dout(n8235));
  jnot g08043(.din(n7916), .dout(n8236));
  jand g08044(.dina(\a[54] ), .dinb(\a[11] ), .dout(n8237));
  jxor g08045(.dina(n8237), .dinb(n8236), .dout(n8238));
  jxor g08046(.dina(n8238), .dinb(n7940), .dout(n8239));
  jand g08047(.dina(\a[35] ), .dinb(\a[30] ), .dout(n8240));
  jand g08048(.dina(\a[33] ), .dinb(\a[32] ), .dout(n8241));
  jor  g08049(.dina(n8241), .dinb(n7932), .dout(n8242));
  jnot g08050(.din(n8242), .dout(n8243));
  jand g08051(.dina(\a[34] ), .dinb(\a[32] ), .dout(n8244));
  jand g08052(.dina(n8244), .dinb(n7928), .dout(n8245));
  jor  g08053(.dina(n8245), .dinb(n8243), .dout(n8246));
  jxor g08054(.dina(n8246), .dinb(n8240), .dout(n8247));
  jxor g08055(.dina(n8247), .dinb(n8239), .dout(n8248));
  jxor g08056(.dina(n8248), .dinb(n8235), .dout(n8249));
  jxor g08057(.dina(n8249), .dinb(n8229), .dout(n8250));
  jand g08058(.dina(\a[39] ), .dinb(\a[26] ), .dout(n8251));
  jnot g08059(.din(n8251), .dout(n8252));
  jand g08060(.dina(\a[37] ), .dinb(\a[28] ), .dout(n8253));
  jand g08061(.dina(\a[38] ), .dinb(\a[27] ), .dout(n8254));
  jor  g08062(.dina(n8254), .dinb(n8253), .dout(n8255));
  jand g08063(.dina(\a[38] ), .dinb(\a[28] ), .dout(n8256));
  jand g08064(.dina(n8256), .dinb(n7936), .dout(n8257));
  jnot g08065(.din(n8257), .dout(n8258));
  jand g08066(.dina(n8258), .dinb(n8255), .dout(n8259));
  jxor g08067(.dina(n8259), .dinb(n8252), .dout(n8260));
  jand g08068(.dina(\a[42] ), .dinb(\a[23] ), .dout(n8261));
  jnot g08069(.din(n8261), .dout(n8262));
  jand g08070(.dina(\a[41] ), .dinb(\a[24] ), .dout(n8263));
  jor  g08071(.dina(n8263), .dinb(n7959), .dout(n8264));
  jand g08072(.dina(\a[41] ), .dinb(\a[25] ), .dout(n8265));
  jand g08073(.dina(n8265), .dinb(n7955), .dout(n8266));
  jnot g08074(.din(n8266), .dout(n8267));
  jand g08075(.dina(n8267), .dinb(n8264), .dout(n8268));
  jxor g08076(.dina(n8268), .dinb(n8262), .dout(n8269));
  jand g08077(.dina(\a[56] ), .dinb(\a[9] ), .dout(n8270));
  jnot g08078(.din(n8270), .dout(n8271));
  jand g08079(.dina(\a[55] ), .dinb(\a[10] ), .dout(n8272));
  jand g08080(.dina(\a[45] ), .dinb(\a[20] ), .dout(n8273));
  jxor g08081(.dina(n8273), .dinb(n8272), .dout(n8274));
  jxor g08082(.dina(n8274), .dinb(n8271), .dout(n8275));
  jnot g08083(.din(n8275), .dout(n8276));
  jxor g08084(.dina(n8276), .dinb(n8269), .dout(n8277));
  jxor g08085(.dina(n8277), .dinb(n8260), .dout(n8278));
  jxor g08086(.dina(n8278), .dinb(n8250), .dout(n8279));
  jxor g08087(.dina(n8279), .dinb(n8206), .dout(n8280));
  jxor g08088(.dina(n8280), .dinb(n8201), .dout(n8281));
  jxor g08089(.dina(n8281), .dinb(n8181), .dout(n8282));
  jxor g08090(.dina(n8282), .dinb(n8119), .dout(n8283));
  jxor g08091(.dina(n8283), .dinb(n8068), .dout(n8284));
  jand g08092(.dina(n8056), .dinb(n8053), .dout(n8285));
  jnot g08093(.din(n8053), .dout(n8286));
  jnot g08094(.din(n8056), .dout(n8287));
  jand g08095(.dina(n8287), .dinb(n8286), .dout(n8288));
  jnot g08096(.din(n8288), .dout(n8289));
  jand g08097(.dina(n8064), .dinb(n8289), .dout(n8290));
  jor  g08098(.dina(n8290), .dinb(n8285), .dout(n8291));
  jxor g08099(.dina(n8291), .dinb(n8284), .dout(\asquared[66] ));
  jand g08100(.dina(n8118), .dinb(n8071), .dout(n8293));
  jand g08101(.dina(n8282), .dinb(n8119), .dout(n8294));
  jor  g08102(.dina(n8294), .dinb(n8293), .dout(n8295));
  jand g08103(.dina(n8116), .dinb(n8079), .dout(n8296));
  jand g08104(.dina(n8117), .dinb(n8074), .dout(n8297));
  jor  g08105(.dina(n8297), .dinb(n8296), .dout(n8298));
  jand g08106(.dina(n8279), .dinb(n8206), .dout(n8299));
  jand g08107(.dina(n8280), .dinb(n8201), .dout(n8300));
  jor  g08108(.dina(n8300), .dinb(n8299), .dout(n8301));
  jxor g08109(.dina(n8301), .dinb(n8298), .dout(n8302));
  jand g08110(.dina(n8085), .dinb(n8082), .dout(n8303));
  jand g08111(.dina(n8115), .dinb(n8086), .dout(n8304));
  jor  g08112(.dina(n8304), .dinb(n8303), .dout(n8305));
  jand g08113(.dina(\a[56] ), .dinb(\a[10] ), .dout(n8306));
  jand g08114(.dina(\a[40] ), .dinb(\a[26] ), .dout(n8307));
  jor  g08115(.dina(n8307), .dinb(n8265), .dout(n8308));
  jnot g08116(.din(n8308), .dout(n8309));
  jand g08117(.dina(\a[41] ), .dinb(\a[26] ), .dout(n8310));
  jand g08118(.dina(n8310), .dinb(n7959), .dout(n8311));
  jor  g08119(.dina(n8311), .dinb(n8309), .dout(n8312));
  jxor g08120(.dina(n8312), .dinb(n8306), .dout(n8313));
  jand g08121(.dina(\a[46] ), .dinb(\a[20] ), .dout(n8314));
  jand g08122(.dina(\a[45] ), .dinb(\a[21] ), .dout(n8315));
  jor  g08123(.dina(n8315), .dinb(n8221), .dout(n8316));
  jnot g08124(.din(n8316), .dout(n8317));
  jand g08125(.dina(\a[45] ), .dinb(\a[22] ), .dout(n8318));
  jand g08126(.dina(n8318), .dinb(n8218), .dout(n8319));
  jor  g08127(.dina(n8319), .dinb(n8317), .dout(n8320));
  jxor g08128(.dina(n8320), .dinb(n8314), .dout(n8321));
  jand g08129(.dina(\a[43] ), .dinb(\a[23] ), .dout(n8322));
  jand g08130(.dina(\a[57] ), .dinb(\a[9] ), .dout(n8323));
  jand g08131(.dina(\a[42] ), .dinb(\a[24] ), .dout(n8324));
  jor  g08132(.dina(n8324), .dinb(n8323), .dout(n8325));
  jand g08133(.dina(\a[57] ), .dinb(\a[24] ), .dout(n8326));
  jand g08134(.dina(n8326), .dinb(n5063), .dout(n8327));
  jnot g08135(.din(n8327), .dout(n8328));
  jand g08136(.dina(n8328), .dinb(n8325), .dout(n8329));
  jxor g08137(.dina(n8329), .dinb(n8322), .dout(n8330));
  jxor g08138(.dina(n8330), .dinb(n8321), .dout(n8331));
  jxor g08139(.dina(n8331), .dinb(n8313), .dout(n8332));
  jand g08140(.dina(\a[50] ), .dinb(\a[16] ), .dout(n8333));
  jor  g08141(.dina(n8333), .dinb(n6019), .dout(n8334));
  jnot g08142(.din(n8334), .dout(n8335));
  jand g08143(.dina(\a[50] ), .dinb(\a[17] ), .dout(n8336));
  jand g08144(.dina(n8336), .dinb(n6419), .dout(n8337));
  jor  g08145(.dina(n8337), .dinb(n8335), .dout(n8338));
  jxor g08146(.dina(n8338), .dinb(n8244), .dout(n8339));
  jand g08147(.dina(\a[52] ), .dinb(\a[14] ), .dout(n8340));
  jand g08148(.dina(\a[36] ), .dinb(\a[30] ), .dout(n8341));
  jand g08149(.dina(\a[35] ), .dinb(\a[31] ), .dout(n8342));
  jor  g08150(.dina(n8342), .dinb(n8341), .dout(n8343));
  jnot g08151(.din(n8343), .dout(n8344));
  jand g08152(.dina(\a[36] ), .dinb(\a[31] ), .dout(n8345));
  jand g08153(.dina(n8345), .dinb(n8240), .dout(n8346));
  jor  g08154(.dina(n8346), .dinb(n8344), .dout(n8347));
  jxor g08155(.dina(n8347), .dinb(n8340), .dout(n8348));
  jand g08156(.dina(\a[48] ), .dinb(\a[18] ), .dout(n8349));
  jand g08157(.dina(\a[53] ), .dinb(\a[13] ), .dout(n8350));
  jor  g08158(.dina(n8350), .dinb(n7235), .dout(n8351));
  jand g08159(.dina(\a[53] ), .dinb(\a[15] ), .dout(n8352));
  jand g08160(.dina(n8352), .dinb(n7815), .dout(n8353));
  jnot g08161(.din(n8353), .dout(n8354));
  jand g08162(.dina(n8354), .dinb(n8351), .dout(n8355));
  jxor g08163(.dina(n8355), .dinb(n8349), .dout(n8356));
  jxor g08164(.dina(n8356), .dinb(n8348), .dout(n8357));
  jxor g08165(.dina(n8357), .dinb(n8339), .dout(n8358));
  jxor g08166(.dina(n8358), .dinb(n8332), .dout(n8359));
  jand g08167(.dina(\a[55] ), .dinb(\a[11] ), .dout(n8360));
  jnot g08168(.din(n8360), .dout(n8361));
  jand g08169(.dina(\a[47] ), .dinb(\a[19] ), .dout(n8362));
  jand g08170(.dina(\a[54] ), .dinb(\a[12] ), .dout(n8363));
  jxor g08171(.dina(n8363), .dinb(n8362), .dout(n8364));
  jxor g08172(.dina(n8364), .dinb(n8361), .dout(n8365));
  jand g08173(.dina(\a[39] ), .dinb(\a[27] ), .dout(n8366));
  jand g08174(.dina(\a[37] ), .dinb(\a[29] ), .dout(n8367));
  jor  g08175(.dina(n8367), .dinb(n8256), .dout(n8368));
  jnot g08176(.din(n8368), .dout(n8369));
  jand g08177(.dina(\a[38] ), .dinb(\a[29] ), .dout(n8370));
  jand g08178(.dina(n8370), .dinb(n8253), .dout(n8371));
  jor  g08179(.dina(n8371), .dinb(n8369), .dout(n8372));
  jxor g08180(.dina(n8372), .dinb(n8366), .dout(n8373));
  jand g08181(.dina(\a[63] ), .dinb(\a[3] ), .dout(n8374));
  jand g08182(.dina(\a[61] ), .dinb(\a[5] ), .dout(n8375));
  jand g08183(.dina(\a[62] ), .dinb(\a[4] ), .dout(n8376));
  jor  g08184(.dina(n8376), .dinb(n8375), .dout(n8377));
  jand g08185(.dina(\a[62] ), .dinb(\a[5] ), .dout(n8378));
  jand g08186(.dina(n8378), .dinb(n7907), .dout(n8379));
  jnot g08187(.din(n8379), .dout(n8380));
  jand g08188(.dina(n8380), .dinb(n8377), .dout(n8381));
  jxor g08189(.dina(n8381), .dinb(n8374), .dout(n8382));
  jxor g08190(.dina(n8382), .dinb(n8373), .dout(n8383));
  jxor g08191(.dina(n8383), .dinb(n8365), .dout(n8384));
  jxor g08192(.dina(n8384), .dinb(n8359), .dout(n8385));
  jxor g08193(.dina(n8385), .dinb(n8305), .dout(n8386));
  jand g08194(.dina(n8103), .dinb(n8095), .dout(n8387));
  jand g08195(.dina(n8104), .dinb(n8093), .dout(n8388));
  jor  g08196(.dina(n8388), .dinb(n8387), .dout(n8389));
  jand g08197(.dina(n8111), .dinb(n8109), .dout(n8390));
  jand g08198(.dina(n8112), .dinb(n8107), .dout(n8391));
  jor  g08199(.dina(n8391), .dinb(n8390), .dout(n8392));
  jxor g08200(.dina(n8392), .dinb(n8389), .dout(n8393));
  jand g08201(.dina(n8126), .dinb(n8124), .dout(n8394));
  jand g08202(.dina(n8129), .dinb(n8127), .dout(n8395));
  jor  g08203(.dina(n8395), .dinb(n8394), .dout(n8396));
  jxor g08204(.dina(n8396), .dinb(n8393), .dout(n8397));
  jand g08205(.dina(n8113), .dinb(n8105), .dout(n8398));
  jand g08206(.dina(n8114), .dinb(n8091), .dout(n8399));
  jor  g08207(.dina(n8399), .dinb(n8398), .dout(n8400));
  jand g08208(.dina(n8136), .dinb(n8130), .dout(n8401));
  jand g08209(.dina(n8143), .dinb(n8137), .dout(n8402));
  jor  g08210(.dina(n8402), .dinb(n8401), .dout(n8403));
  jxor g08211(.dina(n8403), .dinb(n8400), .dout(n8404));
  jxor g08212(.dina(n8404), .dinb(n8397), .dout(n8405));
  jxor g08213(.dina(n8405), .dinb(n8386), .dout(n8406));
  jxor g08214(.dina(n8406), .dinb(n8302), .dout(n8407));
  jand g08215(.dina(n8180), .dinb(n8122), .dout(n8408));
  jand g08216(.dina(n8281), .dinb(n8181), .dout(n8409));
  jor  g08217(.dina(n8409), .dinb(n8408), .dout(n8410));
  jor  g08218(.dina(n8199), .dinb(n8196), .dout(n8411));
  jand g08219(.dina(n8200), .dinb(n8192), .dout(n8412));
  jnot g08220(.din(n8412), .dout(n8413));
  jand g08221(.dina(n8413), .dinb(n8411), .dout(n8414));
  jnot g08222(.din(n8414), .dout(n8415));
  jand g08223(.dina(n8187), .dinb(n8184), .dout(n8416));
  jand g08224(.dina(n8191), .dinb(n8188), .dout(n8417));
  jor  g08225(.dina(n8417), .dinb(n8416), .dout(n8418));
  jor  g08226(.dina(n8176), .dinb(n8171), .dout(n8419));
  jand g08227(.dina(n8177), .dinb(n8164), .dout(n8420));
  jnot g08228(.din(n8420), .dout(n8421));
  jand g08229(.dina(n8421), .dinb(n8419), .dout(n8422));
  jnot g08230(.din(n8422), .dout(n8423));
  jand g08231(.dina(n8163), .dinb(n8161), .dout(n8424));
  jor  g08232(.dina(n8424), .dinb(n8159), .dout(n8425));
  jand g08233(.dina(n8255), .dinb(n8251), .dout(n8426));
  jor  g08234(.dina(n8426), .dinb(n8257), .dout(n8427));
  jxor g08235(.dina(n8427), .dinb(n8425), .dout(n8428));
  jand g08236(.dina(\a[60] ), .dinb(\a[6] ), .dout(n8429));
  jand g08237(.dina(\a[58] ), .dinb(\a[8] ), .dout(n8430));
  jor  g08238(.dina(n8430), .dinb(n8212), .dout(n8431));
  jnot g08239(.din(n8431), .dout(n8432));
  jand g08240(.dina(\a[59] ), .dinb(\a[8] ), .dout(n8433));
  jand g08241(.dina(n8433), .dinb(n8209), .dout(n8434));
  jor  g08242(.dina(n8434), .dinb(n8432), .dout(n8435));
  jxor g08243(.dina(n8435), .dinb(n8429), .dout(n8436));
  jnot g08244(.din(n8436), .dout(n8437));
  jxor g08245(.dina(n8437), .dinb(n8428), .dout(n8438));
  jxor g08246(.dina(n8438), .dinb(n8423), .dout(n8439));
  jxor g08247(.dina(n8439), .dinb(n8418), .dout(n8440));
  jand g08248(.dina(n8242), .dinb(n8240), .dout(n8441));
  jor  g08249(.dina(n8441), .dinb(n8245), .dout(n8442));
  jnot g08250(.din(n8232), .dout(n8443));
  jand g08251(.dina(n8443), .dinb(n8231), .dout(n8444));
  jnot g08252(.din(n8444), .dout(n8445));
  jand g08253(.dina(n8232), .dinb(\a[33] ), .dout(n8446));
  jor  g08254(.dina(n8446), .dinb(n8230), .dout(n8447));
  jand g08255(.dina(n8447), .dinb(n8445), .dout(n8448));
  jxor g08256(.dina(n8448), .dinb(n8442), .dout(n8449));
  jand g08257(.dina(n8167), .dinb(n6419), .dout(n8450));
  jor  g08258(.dina(n8450), .dinb(n8169), .dout(n8451));
  jxor g08259(.dina(n8451), .dinb(n8449), .dout(n8452));
  jand g08260(.dina(n8210), .dinb(n8207), .dout(n8453));
  jor  g08261(.dina(n8453), .dinb(n8213), .dout(n8454));
  jand g08262(.dina(n8219), .dinb(n8217), .dout(n8455));
  jor  g08263(.dina(n8455), .dinb(n8222), .dout(n8456));
  jxor g08264(.dina(n8456), .dinb(n8454), .dout(n8457));
  jnot g08265(.din(n8237), .dout(n8458));
  jand g08266(.dina(n8458), .dinb(n8236), .dout(n8459));
  jnot g08267(.din(n8459), .dout(n8460));
  jand g08268(.dina(n8237), .dinb(n7916), .dout(n8461));
  jor  g08269(.dina(n8461), .dinb(n7940), .dout(n8462));
  jand g08270(.dina(n8462), .dinb(n8460), .dout(n8463));
  jxor g08271(.dina(n8463), .dinb(n8457), .dout(n8464));
  jnot g08272(.din(n8464), .dout(n8465));
  jor  g08273(.dina(n8247), .dinb(n8239), .dout(n8466));
  jand g08274(.dina(n8248), .dinb(n8235), .dout(n8467));
  jnot g08275(.din(n8467), .dout(n8468));
  jand g08276(.dina(n8468), .dinb(n8466), .dout(n8469));
  jxor g08277(.dina(n8469), .dinb(n8465), .dout(n8470));
  jxor g08278(.dina(n8470), .dinb(n8452), .dout(n8471));
  jxor g08279(.dina(n8471), .dinb(n8440), .dout(n8472));
  jxor g08280(.dina(n8472), .dinb(n8415), .dout(n8473));
  jand g08281(.dina(n8147), .dinb(n8144), .dout(n8474));
  jand g08282(.dina(n8179), .dinb(n8148), .dout(n8475));
  jor  g08283(.dina(n8475), .dinb(n8474), .dout(n8476));
  jand g08284(.dina(n8174), .dinb(n8173), .dout(n8477));
  jnot g08285(.din(n8477), .dout(n8478));
  jnot g08286(.din(n8173), .dout(n8479));
  jnot g08287(.din(n8174), .dout(n8480));
  jand g08288(.dina(n8480), .dinb(n8479), .dout(n8481));
  jor  g08289(.dina(n8481), .dinb(n8172), .dout(n8482));
  jand g08290(.dina(n8482), .dinb(n8478), .dout(n8483));
  jand g08291(.dina(n8273), .dinb(n8272), .dout(n8484));
  jnot g08292(.din(n8484), .dout(n8485));
  jnot g08293(.din(n8272), .dout(n8486));
  jnot g08294(.din(n8273), .dout(n8487));
  jand g08295(.dina(n8487), .dinb(n8486), .dout(n8488));
  jor  g08296(.dina(n8488), .dinb(n8271), .dout(n8489));
  jand g08297(.dina(n8489), .dinb(n8485), .dout(n8490));
  jxor g08298(.dina(n8490), .dinb(n8483), .dout(n8491));
  jand g08299(.dina(n8264), .dinb(n8261), .dout(n8492));
  jor  g08300(.dina(n8492), .dinb(n8266), .dout(n8493));
  jxor g08301(.dina(n8493), .dinb(n8491), .dout(n8494));
  jand g08302(.dina(n8227), .dinb(n8225), .dout(n8495));
  jand g08303(.dina(n8228), .dinb(n8216), .dout(n8496));
  jor  g08304(.dina(n8496), .dinb(n8495), .dout(n8497));
  jxor g08305(.dina(n8497), .dinb(n8494), .dout(n8498));
  jnot g08306(.din(n8498), .dout(n8499));
  jnot g08307(.din(n8269), .dout(n8500));
  jand g08308(.dina(n8276), .dinb(n8500), .dout(n8501));
  jnot g08309(.din(n8501), .dout(n8502));
  jand g08310(.dina(n8275), .dinb(n8269), .dout(n8503));
  jor  g08311(.dina(n8503), .dinb(n8260), .dout(n8504));
  jand g08312(.dina(n8504), .dinb(n8502), .dout(n8505));
  jxor g08313(.dina(n8505), .dinb(n8499), .dout(n8506));
  jand g08314(.dina(n8154), .dinb(n8151), .dout(n8507));
  jand g08315(.dina(n8178), .dinb(n8155), .dout(n8508));
  jor  g08316(.dina(n8508), .dinb(n8507), .dout(n8509));
  jor  g08317(.dina(n8249), .dinb(n8229), .dout(n8510));
  jand g08318(.dina(n8249), .dinb(n8229), .dout(n8511));
  jor  g08319(.dina(n8278), .dinb(n8511), .dout(n8512));
  jand g08320(.dina(n8512), .dinb(n8510), .dout(n8513));
  jxor g08321(.dina(n8513), .dinb(n8509), .dout(n8514));
  jxor g08322(.dina(n8514), .dinb(n8506), .dout(n8515));
  jxor g08323(.dina(n8515), .dinb(n8476), .dout(n8516));
  jxor g08324(.dina(n8516), .dinb(n8473), .dout(n8517));
  jxor g08325(.dina(n8517), .dinb(n8410), .dout(n8518));
  jxor g08326(.dina(n8518), .dinb(n8407), .dout(n8519));
  jxor g08327(.dina(n8519), .dinb(n8295), .dout(n8520));
  jand g08328(.dina(n8283), .dinb(n8068), .dout(n8521));
  jor  g08329(.dina(n8283), .dinb(n8068), .dout(n8522));
  jand g08330(.dina(n8291), .dinb(n8522), .dout(n8523));
  jor  g08331(.dina(n8523), .dinb(n8521), .dout(n8524));
  jxor g08332(.dina(n8524), .dinb(n8520), .dout(\asquared[67] ));
  jand g08333(.dina(n8517), .dinb(n8410), .dout(n8526));
  jand g08334(.dina(n8518), .dinb(n8407), .dout(n8527));
  jor  g08335(.dina(n8527), .dinb(n8526), .dout(n8528));
  jand g08336(.dina(n8301), .dinb(n8298), .dout(n8529));
  jand g08337(.dina(n8406), .dinb(n8302), .dout(n8530));
  jor  g08338(.dina(n8530), .dinb(n8529), .dout(n8531));
  jand g08339(.dina(n8471), .dinb(n8440), .dout(n8532));
  jand g08340(.dina(n8472), .dinb(n8415), .dout(n8533));
  jor  g08341(.dina(n8533), .dinb(n8532), .dout(n8534));
  jand g08342(.dina(n8403), .dinb(n8400), .dout(n8535));
  jand g08343(.dina(n8404), .dinb(n8397), .dout(n8536));
  jor  g08344(.dina(n8536), .dinb(n8535), .dout(n8537));
  jnot g08345(.din(n8321), .dout(n8538));
  jor  g08346(.dina(n8330), .dinb(n8538), .dout(n8539));
  jnot g08347(.din(n8313), .dout(n8540));
  jand g08348(.dina(n8330), .dinb(n8538), .dout(n8541));
  jor  g08349(.dina(n8541), .dinb(n8540), .dout(n8542));
  jand g08350(.dina(n8542), .dinb(n8539), .dout(n8543));
  jnot g08351(.din(n8425), .dout(n8544));
  jnot g08352(.din(n8427), .dout(n8545));
  jand g08353(.dina(n8545), .dinb(n8544), .dout(n8546));
  jnot g08354(.din(n8546), .dout(n8547));
  jand g08355(.dina(n8427), .dinb(n8425), .dout(n8548));
  jor  g08356(.dina(n8437), .dinb(n8548), .dout(n8549));
  jand g08357(.dina(n8549), .dinb(n8547), .dout(n8550));
  jxor g08358(.dina(n8550), .dinb(n8543), .dout(n8551));
  jnot g08359(.din(n8373), .dout(n8552));
  jor  g08360(.dina(n8382), .dinb(n8552), .dout(n8553));
  jnot g08361(.din(n8365), .dout(n8554));
  jand g08362(.dina(n8382), .dinb(n8552), .dout(n8555));
  jor  g08363(.dina(n8555), .dinb(n8554), .dout(n8556));
  jand g08364(.dina(n8556), .dinb(n8553), .dout(n8557));
  jxor g08365(.dina(n8557), .dinb(n8551), .dout(n8558));
  jand g08366(.dina(n8381), .dinb(n8374), .dout(n8559));
  jor  g08367(.dina(n8559), .dinb(n8379), .dout(n8560));
  jand g08368(.dina(n8431), .dinb(n8429), .dout(n8561));
  jor  g08369(.dina(n8561), .dinb(n8434), .dout(n8562));
  jxor g08370(.dina(n8562), .dinb(n8560), .dout(n8563));
  jand g08371(.dina(n8368), .dinb(n8366), .dout(n8564));
  jor  g08372(.dina(n8564), .dinb(n8371), .dout(n8565));
  jxor g08373(.dina(n8565), .dinb(n8563), .dout(n8566));
  jand g08374(.dina(n8329), .dinb(n8322), .dout(n8567));
  jor  g08375(.dina(n8567), .dinb(n8327), .dout(n8568));
  jand g08376(.dina(n8308), .dinb(n8306), .dout(n8569));
  jor  g08377(.dina(n8569), .dinb(n8311), .dout(n8570));
  jxor g08378(.dina(n8570), .dinb(n8568), .dout(n8571));
  jand g08379(.dina(n8316), .dinb(n8314), .dout(n8572));
  jor  g08380(.dina(n8572), .dinb(n8319), .dout(n8573));
  jxor g08381(.dina(n8573), .dinb(n8571), .dout(n8574));
  jand g08382(.dina(\a[61] ), .dinb(\a[6] ), .dout(n8575));
  jand g08383(.dina(n8334), .dinb(n8244), .dout(n8576));
  jor  g08384(.dina(n8576), .dinb(n8337), .dout(n8577));
  jxor g08385(.dina(n8577), .dinb(n8575), .dout(n8578));
  jand g08386(.dina(n8343), .dinb(n8340), .dout(n8579));
  jor  g08387(.dina(n8579), .dinb(n8346), .dout(n8580));
  jxor g08388(.dina(n8580), .dinb(n8578), .dout(n8581));
  jxor g08389(.dina(n8581), .dinb(n8574), .dout(n8582));
  jxor g08390(.dina(n8582), .dinb(n8566), .dout(n8583));
  jxor g08391(.dina(n8583), .dinb(n8558), .dout(n8584));
  jxor g08392(.dina(n8584), .dinb(n8537), .dout(n8585));
  jxor g08393(.dina(n8585), .dinb(n8534), .dout(n8586));
  jand g08394(.dina(n8355), .dinb(n8349), .dout(n8587));
  jor  g08395(.dina(n8587), .dinb(n8353), .dout(n8588));
  jnot g08396(.din(n8588), .dout(n8589));
  jand g08397(.dina(n8363), .dinb(n8362), .dout(n8590));
  jnot g08398(.din(n8590), .dout(n8591));
  jnot g08399(.din(n8362), .dout(n8592));
  jnot g08400(.din(n8363), .dout(n8593));
  jand g08401(.dina(n8593), .dinb(n8592), .dout(n8594));
  jor  g08402(.dina(n8594), .dinb(n8361), .dout(n8595));
  jand g08403(.dina(n8595), .dinb(n8591), .dout(n8596));
  jxor g08404(.dina(n8596), .dinb(n8589), .dout(n8597));
  jand g08405(.dina(\a[57] ), .dinb(\a[10] ), .dout(n8598));
  jnot g08406(.din(n8598), .dout(n8599));
  jand g08407(.dina(\a[56] ), .dinb(\a[11] ), .dout(n8600));
  jand g08408(.dina(\a[47] ), .dinb(\a[20] ), .dout(n8601));
  jor  g08409(.dina(n8601), .dinb(n8600), .dout(n8602));
  jand g08410(.dina(\a[56] ), .dinb(\a[20] ), .dout(n8603));
  jand g08411(.dina(n8603), .dinb(n6654), .dout(n8604));
  jnot g08412(.din(n8604), .dout(n8605));
  jand g08413(.dina(n8605), .dinb(n8602), .dout(n8606));
  jxor g08414(.dina(n8606), .dinb(n8599), .dout(n8607));
  jnot g08415(.din(n8607), .dout(n8608));
  jxor g08416(.dina(n8608), .dinb(n8597), .dout(n8609));
  jnot g08417(.din(n8348), .dout(n8610));
  jor  g08418(.dina(n8356), .dinb(n8610), .dout(n8611));
  jnot g08419(.din(n8339), .dout(n8612));
  jand g08420(.dina(n8356), .dinb(n8610), .dout(n8613));
  jor  g08421(.dina(n8613), .dinb(n8612), .dout(n8614));
  jand g08422(.dina(n8614), .dinb(n8611), .dout(n8615));
  jxor g08423(.dina(n8615), .dinb(n8609), .dout(n8616));
  jand g08424(.dina(n8392), .dinb(n8389), .dout(n8617));
  jand g08425(.dina(n8396), .dinb(n8393), .dout(n8618));
  jor  g08426(.dina(n8618), .dinb(n8617), .dout(n8619));
  jxor g08427(.dina(n8619), .dinb(n8616), .dout(n8620));
  jand g08428(.dina(n8358), .dinb(n8332), .dout(n8621));
  jand g08429(.dina(n8384), .dinb(n8359), .dout(n8622));
  jor  g08430(.dina(n8622), .dinb(n8621), .dout(n8623));
  jand g08431(.dina(n8438), .dinb(n8423), .dout(n8624));
  jand g08432(.dina(n8439), .dinb(n8418), .dout(n8625));
  jor  g08433(.dina(n8625), .dinb(n8624), .dout(n8626));
  jxor g08434(.dina(n8626), .dinb(n8623), .dout(n8627));
  jxor g08435(.dina(n8627), .dinb(n8620), .dout(n8628));
  jxor g08436(.dina(n8628), .dinb(n8586), .dout(n8629));
  jxor g08437(.dina(n8629), .dinb(n8531), .dout(n8630));
  jand g08438(.dina(n8515), .dinb(n8476), .dout(n8631));
  jand g08439(.dina(n8516), .dinb(n8473), .dout(n8632));
  jor  g08440(.dina(n8632), .dinb(n8631), .dout(n8633));
  jand g08441(.dina(n8385), .dinb(n8305), .dout(n8634));
  jand g08442(.dina(n8405), .dinb(n8386), .dout(n8635));
  jor  g08443(.dina(n8635), .dinb(n8634), .dout(n8636));
  jxor g08444(.dina(n8636), .dinb(n8633), .dout(n8637));
  jand g08445(.dina(n8513), .dinb(n8509), .dout(n8638));
  jand g08446(.dina(n8514), .dinb(n8506), .dout(n8639));
  jor  g08447(.dina(n8639), .dinb(n8638), .dout(n8640));
  jand g08448(.dina(\a[55] ), .dinb(\a[12] ), .dout(n8641));
  jand g08449(.dina(\a[54] ), .dinb(\a[13] ), .dout(n8642));
  jor  g08450(.dina(n8642), .dinb(n8641), .dout(n8643));
  jnot g08451(.din(n8643), .dout(n8644));
  jand g08452(.dina(\a[55] ), .dinb(\a[13] ), .dout(n8645));
  jand g08453(.dina(n8645), .dinb(n8363), .dout(n8646));
  jor  g08454(.dina(n8646), .dinb(n8644), .dout(n8647));
  jxor g08455(.dina(n8647), .dinb(n8370), .dout(n8648));
  jnot g08456(.din(n8648), .dout(n8649));
  jand g08457(.dina(\a[49] ), .dinb(\a[18] ), .dout(n8650));
  jnot g08458(.din(n8650), .dout(n8651));
  jnot g08459(.din(\a[34] ), .dout(n8652));
  jnot g08460(.din(n8378), .dout(n8653));
  jand g08461(.dina(n8653), .dinb(n8652), .dout(n8654));
  jnot g08462(.din(n8654), .dout(n8655));
  jand g08463(.dina(n3127), .dinb(\a[62] ), .dout(n8656));
  jnot g08464(.din(n8656), .dout(n8657));
  jand g08465(.dina(n8657), .dinb(n8655), .dout(n8658));
  jor  g08466(.dina(n8658), .dinb(n8651), .dout(n8659));
  jand g08467(.dina(n8655), .dinb(n8650), .dout(n8660));
  jor  g08468(.dina(n8660), .dinb(n8656), .dout(n8661));
  jnot g08469(.din(n8661), .dout(n8662));
  jand g08470(.dina(n8662), .dinb(n8655), .dout(n8663));
  jnot g08471(.din(n8663), .dout(n8664));
  jand g08472(.dina(n8664), .dinb(n8659), .dout(n8665));
  jand g08473(.dina(\a[35] ), .dinb(\a[32] ), .dout(n8666));
  jand g08474(.dina(\a[34] ), .dinb(\a[33] ), .dout(n8667));
  jor  g08475(.dina(n8667), .dinb(n8666), .dout(n8668));
  jnot g08476(.din(n8668), .dout(n8669));
  jand g08477(.dina(\a[35] ), .dinb(\a[33] ), .dout(n8670));
  jand g08478(.dina(n8670), .dinb(n8244), .dout(n8671));
  jor  g08479(.dina(n8671), .dinb(n8669), .dout(n8672));
  jxor g08480(.dina(n8672), .dinb(n8345), .dout(n8673));
  jxor g08481(.dina(n8673), .dinb(n8665), .dout(n8674));
  jxor g08482(.dina(n8674), .dinb(n8649), .dout(n8675));
  jand g08483(.dina(\a[44] ), .dinb(\a[23] ), .dout(n8676));
  jand g08484(.dina(\a[43] ), .dinb(\a[24] ), .dout(n8677));
  jor  g08485(.dina(n8677), .dinb(n8676), .dout(n8678));
  jnot g08486(.din(n8678), .dout(n8679));
  jand g08487(.dina(\a[44] ), .dinb(\a[24] ), .dout(n8680));
  jand g08488(.dina(n8680), .dinb(n8322), .dout(n8681));
  jor  g08489(.dina(n8681), .dinb(n8679), .dout(n8682));
  jxor g08490(.dina(n8682), .dinb(n8318), .dout(n8683));
  jnot g08491(.din(n8683), .dout(n8684));
  jand g08492(.dina(\a[60] ), .dinb(\a[7] ), .dout(n8685));
  jand g08493(.dina(\a[58] ), .dinb(\a[9] ), .dout(n8686));
  jor  g08494(.dina(n8686), .dinb(n8433), .dout(n8687));
  jand g08495(.dina(\a[59] ), .dinb(\a[9] ), .dout(n8688));
  jand g08496(.dina(n8688), .dinb(n8430), .dout(n8689));
  jnot g08497(.din(n8689), .dout(n8690));
  jand g08498(.dina(n8690), .dinb(n8687), .dout(n8691));
  jxor g08499(.dina(n8691), .dinb(n8685), .dout(n8692));
  jxor g08500(.dina(n8692), .dinb(n8684), .dout(n8693));
  jand g08501(.dina(\a[52] ), .dinb(\a[15] ), .dout(n8694));
  jnot g08502(.din(n7041), .dout(n8695));
  jand g08503(.dina(\a[37] ), .dinb(\a[30] ), .dout(n8696));
  jxor g08504(.dina(n8696), .dinb(n8695), .dout(n8697));
  jxor g08505(.dina(n8697), .dinb(n8694), .dout(n8698));
  jnot g08506(.din(n8698), .dout(n8699));
  jxor g08507(.dina(n8699), .dinb(n8693), .dout(n8700));
  jxor g08508(.dina(n8700), .dinb(n8675), .dout(n8701));
  jnot g08509(.din(n8158), .dout(n8702));
  jand g08510(.dina(\a[40] ), .dinb(\a[27] ), .dout(n8703));
  jand g08511(.dina(\a[39] ), .dinb(\a[28] ), .dout(n8704));
  jor  g08512(.dina(n8704), .dinb(n8703), .dout(n8705));
  jand g08513(.dina(\a[40] ), .dinb(\a[28] ), .dout(n8706));
  jand g08514(.dina(n8706), .dinb(n8366), .dout(n8707));
  jnot g08515(.din(n8707), .dout(n8708));
  jand g08516(.dina(n8708), .dinb(n8705), .dout(n8709));
  jxor g08517(.dina(n8709), .dinb(n8702), .dout(n8710));
  jand g08518(.dina(\a[42] ), .dinb(\a[25] ), .dout(n8711));
  jnot g08519(.din(n8711), .dout(n8712));
  jand g08520(.dina(\a[46] ), .dinb(\a[21] ), .dout(n8713));
  jxor g08521(.dina(n8713), .dinb(n8310), .dout(n8714));
  jxor g08522(.dina(n8714), .dinb(n8712), .dout(n8715));
  jand g08523(.dina(\a[53] ), .dinb(\a[48] ), .dout(n8716));
  jand g08524(.dina(n8716), .dinb(\a[14] ), .dout(n8717));
  jand g08525(.dina(n8336), .dinb(\a[48] ), .dout(n8718));
  jor  g08526(.dina(n8718), .dinb(n8717), .dout(n8719));
  jand g08527(.dina(n8719), .dinb(\a[19] ), .dout(n8720));
  jnot g08528(.din(n8720), .dout(n8721));
  jand g08529(.dina(\a[53] ), .dinb(\a[14] ), .dout(n8722));
  jxor g08530(.dina(n8722), .dinb(n8336), .dout(n8723));
  jand g08531(.dina(n8723), .dinb(n8721), .dout(n8724));
  jnot g08532(.din(n8723), .dout(n8725));
  jand g08533(.dina(\a[48] ), .dinb(\a[19] ), .dout(n8726));
  jand g08534(.dina(n8726), .dinb(n8725), .dout(n8727));
  jor  g08535(.dina(n8727), .dinb(n8724), .dout(n8728));
  jxor g08536(.dina(n8728), .dinb(n8715), .dout(n8729));
  jxor g08537(.dina(n8729), .dinb(n8710), .dout(n8730));
  jxor g08538(.dina(n8730), .dinb(n8701), .dout(n8731));
  jxor g08539(.dina(n8731), .dinb(n8640), .dout(n8732));
  jand g08540(.dina(n8456), .dinb(n8454), .dout(n8733));
  jand g08541(.dina(n8463), .dinb(n8457), .dout(n8734));
  jor  g08542(.dina(n8734), .dinb(n8733), .dout(n8735));
  jnot g08543(.din(n8483), .dout(n8736));
  jnot g08544(.din(n8490), .dout(n8737));
  jand g08545(.dina(n8737), .dinb(n8736), .dout(n8738));
  jand g08546(.dina(n8493), .dinb(n8491), .dout(n8739));
  jor  g08547(.dina(n8739), .dinb(n8738), .dout(n8740));
  jxor g08548(.dina(n8740), .dinb(n8735), .dout(n8741));
  jand g08549(.dina(n8448), .dinb(n8442), .dout(n8742));
  jand g08550(.dina(n8451), .dinb(n8449), .dout(n8743));
  jor  g08551(.dina(n8743), .dinb(n8742), .dout(n8744));
  jxor g08552(.dina(n8744), .dinb(n8741), .dout(n8745));
  jor  g08553(.dina(n8469), .dinb(n8465), .dout(n8746));
  jand g08554(.dina(n8470), .dinb(n8452), .dout(n8747));
  jnot g08555(.din(n8747), .dout(n8748));
  jand g08556(.dina(n8748), .dinb(n8746), .dout(n8749));
  jand g08557(.dina(n8497), .dinb(n8494), .dout(n8750));
  jnot g08558(.din(n8750), .dout(n8751));
  jor  g08559(.dina(n8505), .dinb(n8499), .dout(n8752));
  jand g08560(.dina(n8752), .dinb(n8751), .dout(n8753));
  jxor g08561(.dina(n8753), .dinb(n8749), .dout(n8754));
  jxor g08562(.dina(n8754), .dinb(n8745), .dout(n8755));
  jxor g08563(.dina(n8755), .dinb(n8732), .dout(n8756));
  jxor g08564(.dina(n8756), .dinb(n8637), .dout(n8757));
  jxor g08565(.dina(n8757), .dinb(n8630), .dout(n8758));
  jxor g08566(.dina(n8758), .dinb(n8528), .dout(n8759));
  jand g08567(.dina(n8519), .dinb(n8295), .dout(n8760));
  jor  g08568(.dina(n8519), .dinb(n8295), .dout(n8761));
  jand g08569(.dina(n8524), .dinb(n8761), .dout(n8762));
  jor  g08570(.dina(n8762), .dinb(n8760), .dout(n8763));
  jxor g08571(.dina(n8763), .dinb(n8759), .dout(\asquared[68] ));
  jand g08572(.dina(n8629), .dinb(n8531), .dout(n8765));
  jand g08573(.dina(n8757), .dinb(n8630), .dout(n8766));
  jor  g08574(.dina(n8766), .dinb(n8765), .dout(n8767));
  jand g08575(.dina(n8585), .dinb(n8534), .dout(n8768));
  jand g08576(.dina(n8628), .dinb(n8586), .dout(n8769));
  jor  g08577(.dina(n8769), .dinb(n8768), .dout(n8770));
  jand g08578(.dina(n8731), .dinb(n8640), .dout(n8771));
  jand g08579(.dina(n8755), .dinb(n8732), .dout(n8772));
  jor  g08580(.dina(n8772), .dinb(n8771), .dout(n8773));
  jand g08581(.dina(n8626), .dinb(n8623), .dout(n8774));
  jand g08582(.dina(n8627), .dinb(n8620), .dout(n8775));
  jor  g08583(.dina(n8775), .dinb(n8774), .dout(n8776));
  jand g08584(.dina(n8581), .dinb(n8574), .dout(n8777));
  jand g08585(.dina(n8582), .dinb(n8566), .dout(n8778));
  jor  g08586(.dina(n8778), .dinb(n8777), .dout(n8779));
  jand g08587(.dina(n8550), .dinb(n8543), .dout(n8780));
  jand g08588(.dina(n8557), .dinb(n8551), .dout(n8781));
  jor  g08589(.dina(n8781), .dinb(n8780), .dout(n8782));
  jxor g08590(.dina(n8782), .dinb(n8779), .dout(n8783));
  jand g08591(.dina(n8615), .dinb(n8609), .dout(n8784));
  jand g08592(.dina(n8619), .dinb(n8616), .dout(n8785));
  jor  g08593(.dina(n8785), .dinb(n8784), .dout(n8786));
  jxor g08594(.dina(n8786), .dinb(n8783), .dout(n8787));
  jand g08595(.dina(\a[38] ), .dinb(\a[30] ), .dout(n8788));
  jand g08596(.dina(\a[37] ), .dinb(\a[31] ), .dout(n8789));
  jand g08597(.dina(\a[36] ), .dinb(\a[32] ), .dout(n8790));
  jor  g08598(.dina(n8790), .dinb(n8789), .dout(n8791));
  jnot g08599(.din(n8791), .dout(n8792));
  jand g08600(.dina(\a[37] ), .dinb(\a[32] ), .dout(n8793));
  jand g08601(.dina(n8793), .dinb(n8345), .dout(n8794));
  jor  g08602(.dina(n8794), .dinb(n8792), .dout(n8795));
  jxor g08603(.dina(n8795), .dinb(n8788), .dout(n8796));
  jnot g08604(.din(n8796), .dout(n8797));
  jand g08605(.dina(\a[50] ), .dinb(\a[18] ), .dout(n8798));
  jand g08606(.dina(\a[49] ), .dinb(\a[19] ), .dout(n8799));
  jor  g08607(.dina(n8799), .dinb(n8798), .dout(n8800));
  jand g08608(.dina(\a[50] ), .dinb(\a[19] ), .dout(n8801));
  jand g08609(.dina(n8801), .dinb(n8650), .dout(n8802));
  jnot g08610(.din(n8802), .dout(n8803));
  jand g08611(.dina(n8803), .dinb(n8800), .dout(n8804));
  jxor g08612(.dina(n8804), .dinb(n8670), .dout(n8805));
  jxor g08613(.dina(n8805), .dinb(n8797), .dout(n8806));
  jnot g08614(.din(n8806), .dout(n8807));
  jand g08615(.dina(\a[56] ), .dinb(\a[12] ), .dout(n8808));
  jnot g08616(.din(n6356), .dout(n8809));
  jxor g08617(.dina(n8645), .dinb(n8809), .dout(n8810));
  jxor g08618(.dina(n8810), .dinb(n8808), .dout(n8811));
  jxor g08619(.dina(n8811), .dinb(n8807), .dout(n8812));
  jand g08620(.dina(\a[43] ), .dinb(\a[25] ), .dout(n8813));
  jand g08621(.dina(\a[42] ), .dinb(\a[26] ), .dout(n8814));
  jor  g08622(.dina(n8814), .dinb(n8813), .dout(n8815));
  jnot g08623(.din(n8815), .dout(n8816));
  jand g08624(.dina(\a[43] ), .dinb(\a[26] ), .dout(n8817));
  jand g08625(.dina(n8817), .dinb(n8711), .dout(n8818));
  jor  g08626(.dina(n8818), .dinb(n8816), .dout(n8819));
  jxor g08627(.dina(n8819), .dinb(n8680), .dout(n8820));
  jand g08628(.dina(\a[48] ), .dinb(\a[20] ), .dout(n8821));
  jand g08629(.dina(\a[45] ), .dinb(\a[23] ), .dout(n8822));
  jand g08630(.dina(\a[46] ), .dinb(\a[22] ), .dout(n8823));
  jor  g08631(.dina(n8823), .dinb(n8822), .dout(n8824));
  jnot g08632(.din(n8824), .dout(n8825));
  jand g08633(.dina(\a[46] ), .dinb(\a[23] ), .dout(n8826));
  jand g08634(.dina(n8826), .dinb(n8318), .dout(n8827));
  jor  g08635(.dina(n8827), .dinb(n8825), .dout(n8828));
  jxor g08636(.dina(n8828), .dinb(n8821), .dout(n8829));
  jand g08637(.dina(\a[54] ), .dinb(\a[14] ), .dout(n8830));
  jor  g08638(.dina(n8352), .dinb(n7796), .dout(n8831));
  jand g08639(.dina(\a[53] ), .dinb(\a[16] ), .dout(n8832));
  jand g08640(.dina(n8832), .dinb(n8694), .dout(n8833));
  jnot g08641(.din(n8833), .dout(n8834));
  jand g08642(.dina(n8834), .dinb(n8831), .dout(n8835));
  jxor g08643(.dina(n8835), .dinb(n8830), .dout(n8836));
  jxor g08644(.dina(n8836), .dinb(n8829), .dout(n8837));
  jxor g08645(.dina(n8837), .dinb(n8820), .dout(n8838));
  jxor g08646(.dina(n8838), .dinb(n8812), .dout(n8839));
  jand g08647(.dina(\a[47] ), .dinb(\a[21] ), .dout(n8840));
  jand g08648(.dina(\a[63] ), .dinb(\a[5] ), .dout(n8841));
  jand g08649(.dina(\a[62] ), .dinb(\a[6] ), .dout(n8842));
  jor  g08650(.dina(n8842), .dinb(n8841), .dout(n8843));
  jnot g08651(.din(n8843), .dout(n8844));
  jand g08652(.dina(\a[63] ), .dinb(\a[6] ), .dout(n8845));
  jand g08653(.dina(n8845), .dinb(n8378), .dout(n8846));
  jor  g08654(.dina(n8846), .dinb(n8844), .dout(n8847));
  jxor g08655(.dina(n8847), .dinb(n8840), .dout(n8848));
  jand g08656(.dina(\a[41] ), .dinb(\a[27] ), .dout(n8849));
  jand g08657(.dina(\a[39] ), .dinb(\a[29] ), .dout(n8850));
  jor  g08658(.dina(n8850), .dinb(n8706), .dout(n8851));
  jnot g08659(.din(n8851), .dout(n8852));
  jand g08660(.dina(\a[40] ), .dinb(\a[29] ), .dout(n8853));
  jand g08661(.dina(n8853), .dinb(n8704), .dout(n8854));
  jor  g08662(.dina(n8854), .dinb(n8852), .dout(n8855));
  jxor g08663(.dina(n8855), .dinb(n8849), .dout(n8856));
  jand g08664(.dina(\a[58] ), .dinb(\a[10] ), .dout(n8857));
  jand g08665(.dina(\a[57] ), .dinb(\a[11] ), .dout(n8858));
  jor  g08666(.dina(n8858), .dinb(n8857), .dout(n8859));
  jand g08667(.dina(\a[58] ), .dinb(\a[11] ), .dout(n8860));
  jand g08668(.dina(n8860), .dinb(n8598), .dout(n8861));
  jnot g08669(.din(n8861), .dout(n8862));
  jand g08670(.dina(n8862), .dinb(n8859), .dout(n8863));
  jxor g08671(.dina(n8863), .dinb(n8688), .dout(n8864));
  jxor g08672(.dina(n8864), .dinb(n8856), .dout(n8865));
  jxor g08673(.dina(n8865), .dinb(n8848), .dout(n8866));
  jxor g08674(.dina(n8866), .dinb(n8839), .dout(n8867));
  jxor g08675(.dina(n8867), .dinb(n8787), .dout(n8868));
  jxor g08676(.dina(n8868), .dinb(n8776), .dout(n8869));
  jxor g08677(.dina(n8869), .dinb(n8773), .dout(n8870));
  jxor g08678(.dina(n8870), .dinb(n8770), .dout(n8871));
  jand g08679(.dina(n8636), .dinb(n8633), .dout(n8872));
  jand g08680(.dina(n8756), .dinb(n8637), .dout(n8873));
  jor  g08681(.dina(n8873), .dinb(n8872), .dout(n8874));
  jor  g08682(.dina(n8753), .dinb(n8749), .dout(n8875));
  jand g08683(.dina(n8754), .dinb(n8745), .dout(n8876));
  jnot g08684(.din(n8876), .dout(n8877));
  jand g08685(.dina(n8877), .dinb(n8875), .dout(n8878));
  jnot g08686(.din(n8878), .dout(n8879));
  jand g08687(.dina(n8722), .dinb(n8336), .dout(n8880));
  jor  g08688(.dina(n8880), .dinb(n8720), .dout(n8881));
  jnot g08689(.din(n8310), .dout(n8882));
  jnot g08690(.din(n8713), .dout(n8883));
  jand g08691(.dina(n8883), .dinb(n8882), .dout(n8884));
  jnot g08692(.din(n8884), .dout(n8885));
  jand g08693(.dina(n8713), .dinb(n8310), .dout(n8886));
  jor  g08694(.dina(n8886), .dinb(n8711), .dout(n8887));
  jand g08695(.dina(n8887), .dinb(n8885), .dout(n8888));
  jxor g08696(.dina(n8888), .dinb(n8881), .dout(n8889));
  jand g08697(.dina(n8643), .dinb(n8370), .dout(n8890));
  jor  g08698(.dina(n8890), .dinb(n8646), .dout(n8891));
  jxor g08699(.dina(n8891), .dinb(n8889), .dout(n8892));
  jor  g08700(.dina(n8673), .dinb(n8665), .dout(n8893));
  jand g08701(.dina(n8674), .dinb(n8649), .dout(n8894));
  jnot g08702(.din(n8894), .dout(n8895));
  jand g08703(.dina(n8895), .dinb(n8893), .dout(n8896));
  jnot g08704(.din(n8715), .dout(n8897));
  jand g08705(.dina(n8728), .dinb(n8897), .dout(n8898));
  jnot g08706(.din(n8898), .dout(n8899));
  jnot g08707(.din(n8728), .dout(n8900));
  jand g08708(.dina(n8900), .dinb(n8715), .dout(n8901));
  jor  g08709(.dina(n8901), .dinb(n8710), .dout(n8902));
  jand g08710(.dina(n8902), .dinb(n8899), .dout(n8903));
  jxor g08711(.dina(n8903), .dinb(n8896), .dout(n8904));
  jxor g08712(.dina(n8904), .dinb(n8892), .dout(n8905));
  jand g08713(.dina(n8740), .dinb(n8735), .dout(n8906));
  jand g08714(.dina(n8744), .dinb(n8741), .dout(n8907));
  jor  g08715(.dina(n8907), .dinb(n8906), .dout(n8908));
  jand g08716(.dina(n8691), .dinb(n8685), .dout(n8909));
  jor  g08717(.dina(n8909), .dinb(n8689), .dout(n8910));
  jand g08718(.dina(n8602), .dinb(n8598), .dout(n8911));
  jor  g08719(.dina(n8911), .dinb(n8604), .dout(n8912));
  jand g08720(.dina(n8678), .dinb(n8318), .dout(n8913));
  jor  g08721(.dina(n8913), .dinb(n8681), .dout(n8914));
  jxor g08722(.dina(n8914), .dinb(n8912), .dout(n8915));
  jxor g08723(.dina(n8915), .dinb(n8910), .dout(n8916));
  jand g08724(.dina(n8705), .dinb(n8158), .dout(n8917));
  jor  g08725(.dina(n8917), .dinb(n8707), .dout(n8918));
  jand g08726(.dina(n8668), .dinb(n8345), .dout(n8919));
  jor  g08727(.dina(n8919), .dinb(n8671), .dout(n8920));
  jxor g08728(.dina(n8920), .dinb(n8918), .dout(n8921));
  jnot g08729(.din(n8696), .dout(n8922));
  jand g08730(.dina(n8922), .dinb(n8695), .dout(n8923));
  jnot g08731(.din(n8923), .dout(n8924));
  jand g08732(.dina(n8696), .dinb(n7041), .dout(n8925));
  jor  g08733(.dina(n8925), .dinb(n8694), .dout(n8926));
  jand g08734(.dina(n8926), .dinb(n8924), .dout(n8927));
  jxor g08735(.dina(n8927), .dinb(n8921), .dout(n8928));
  jxor g08736(.dina(n8928), .dinb(n8916), .dout(n8929));
  jxor g08737(.dina(n8929), .dinb(n8908), .dout(n8930));
  jxor g08738(.dina(n8930), .dinb(n8905), .dout(n8931));
  jxor g08739(.dina(n8931), .dinb(n8879), .dout(n8932));
  jand g08740(.dina(n8583), .dinb(n8558), .dout(n8933));
  jand g08741(.dina(n8584), .dinb(n8537), .dout(n8934));
  jor  g08742(.dina(n8934), .dinb(n8933), .dout(n8935));
  jand g08743(.dina(n8700), .dinb(n8675), .dout(n8936));
  jand g08744(.dina(n8730), .dinb(n8701), .dout(n8937));
  jor  g08745(.dina(n8937), .dinb(n8936), .dout(n8938));
  jand g08746(.dina(n8570), .dinb(n8568), .dout(n8939));
  jand g08747(.dina(n8573), .dinb(n8571), .dout(n8940));
  jor  g08748(.dina(n8940), .dinb(n8939), .dout(n8941));
  jand g08749(.dina(n8596), .dinb(n8589), .dout(n8942));
  jor  g08750(.dina(n8596), .dinb(n8589), .dout(n8943));
  jand g08751(.dina(n8607), .dinb(n8943), .dout(n8944));
  jor  g08752(.dina(n8944), .dinb(n8942), .dout(n8945));
  jnot g08753(.din(n8945), .dout(n8946));
  jxor g08754(.dina(n8946), .dinb(n8941), .dout(n8947));
  jor  g08755(.dina(n8692), .dinb(n8684), .dout(n8948));
  jand g08756(.dina(n8692), .dinb(n8684), .dout(n8949));
  jor  g08757(.dina(n8699), .dinb(n8949), .dout(n8950));
  jand g08758(.dina(n8950), .dinb(n8948), .dout(n8951));
  jxor g08759(.dina(n8951), .dinb(n8947), .dout(n8952));
  jand g08760(.dina(n8577), .dinb(n8575), .dout(n8953));
  jand g08761(.dina(n8580), .dinb(n8578), .dout(n8954));
  jor  g08762(.dina(n8954), .dinb(n8953), .dout(n8955));
  jand g08763(.dina(\a[60] ), .dinb(\a[8] ), .dout(n8956));
  jand g08764(.dina(\a[61] ), .dinb(\a[7] ), .dout(n8957));
  jor  g08765(.dina(n8957), .dinb(n8956), .dout(n8958));
  jand g08766(.dina(\a[61] ), .dinb(\a[8] ), .dout(n8959));
  jand g08767(.dina(n8959), .dinb(n8685), .dout(n8960));
  jnot g08768(.din(n8960), .dout(n8961));
  jand g08769(.dina(n8961), .dinb(n8958), .dout(n8962));
  jxor g08770(.dina(n8962), .dinb(n8661), .dout(n8963));
  jxor g08771(.dina(n8963), .dinb(n8955), .dout(n8964));
  jand g08772(.dina(n8562), .dinb(n8560), .dout(n8965));
  jand g08773(.dina(n8565), .dinb(n8563), .dout(n8966));
  jor  g08774(.dina(n8966), .dinb(n8965), .dout(n8967));
  jxor g08775(.dina(n8967), .dinb(n8964), .dout(n8968));
  jxor g08776(.dina(n8968), .dinb(n8952), .dout(n8969));
  jxor g08777(.dina(n8969), .dinb(n8938), .dout(n8970));
  jxor g08778(.dina(n8970), .dinb(n8935), .dout(n8971));
  jxor g08779(.dina(n8971), .dinb(n8932), .dout(n8972));
  jxor g08780(.dina(n8972), .dinb(n8874), .dout(n8973));
  jxor g08781(.dina(n8973), .dinb(n8871), .dout(n8974));
  jxor g08782(.dina(n8974), .dinb(n8767), .dout(n8975));
  jand g08783(.dina(n8758), .dinb(n8528), .dout(n8976));
  jor  g08784(.dina(n8758), .dinb(n8528), .dout(n8977));
  jand g08785(.dina(n8763), .dinb(n8977), .dout(n8978));
  jor  g08786(.dina(n8978), .dinb(n8976), .dout(n8979));
  jxor g08787(.dina(n8979), .dinb(n8975), .dout(\asquared[69] ));
  jand g08788(.dina(n8972), .dinb(n8874), .dout(n8981));
  jand g08789(.dina(n8973), .dinb(n8871), .dout(n8982));
  jor  g08790(.dina(n8982), .dinb(n8981), .dout(n8983));
  jand g08791(.dina(n8869), .dinb(n8773), .dout(n8984));
  jand g08792(.dina(n8870), .dinb(n8770), .dout(n8985));
  jor  g08793(.dina(n8985), .dinb(n8984), .dout(n8986));
  jand g08794(.dina(n8930), .dinb(n8905), .dout(n8987));
  jand g08795(.dina(n8931), .dinb(n8879), .dout(n8988));
  jor  g08796(.dina(n8988), .dinb(n8987), .dout(n8989));
  jand g08797(.dina(n8838), .dinb(n8812), .dout(n8990));
  jand g08798(.dina(n8866), .dinb(n8839), .dout(n8991));
  jor  g08799(.dina(n8991), .dinb(n8990), .dout(n8992));
  jand g08800(.dina(n8928), .dinb(n8916), .dout(n8993));
  jand g08801(.dina(n8929), .dinb(n8908), .dout(n8994));
  jor  g08802(.dina(n8994), .dinb(n8993), .dout(n8995));
  jand g08803(.dina(n8815), .dinb(n8680), .dout(n8996));
  jor  g08804(.dina(n8996), .dinb(n8818), .dout(n8997));
  jnot g08805(.din(n8645), .dout(n8998));
  jand g08806(.dina(n8998), .dinb(n8809), .dout(n8999));
  jnot g08807(.din(n8999), .dout(n9000));
  jand g08808(.dina(n8645), .dinb(n6356), .dout(n9001));
  jor  g08809(.dina(n9001), .dinb(n8808), .dout(n9002));
  jand g08810(.dina(n9002), .dinb(n9000), .dout(n9003));
  jxor g08811(.dina(n9003), .dinb(n8997), .dout(n9004));
  jand g08812(.dina(n8851), .dinb(n8849), .dout(n9005));
  jor  g08813(.dina(n9005), .dinb(n8854), .dout(n9006));
  jxor g08814(.dina(n9006), .dinb(n9004), .dout(n9007));
  jand g08815(.dina(n8920), .dinb(n8918), .dout(n9008));
  jand g08816(.dina(n8927), .dinb(n8921), .dout(n9009));
  jor  g08817(.dina(n9009), .dinb(n9008), .dout(n9010));
  jand g08818(.dina(n8888), .dinb(n8881), .dout(n9011));
  jand g08819(.dina(n8891), .dinb(n8889), .dout(n9012));
  jor  g08820(.dina(n9012), .dinb(n9011), .dout(n9013));
  jxor g08821(.dina(n9013), .dinb(n9010), .dout(n9014));
  jxor g08822(.dina(n9014), .dinb(n9007), .dout(n9015));
  jxor g08823(.dina(n9015), .dinb(n8995), .dout(n9016));
  jxor g08824(.dina(n9016), .dinb(n8992), .dout(n9017));
  jxor g08825(.dina(n9017), .dinb(n8989), .dout(n9018));
  jand g08826(.dina(n8782), .dinb(n8779), .dout(n9019));
  jand g08827(.dina(n8786), .dinb(n8783), .dout(n9020));
  jor  g08828(.dina(n9020), .dinb(n9019), .dout(n9021));
  jand g08829(.dina(n8805), .dinb(n8797), .dout(n9022));
  jnot g08830(.din(n9022), .dout(n9023));
  jor  g08831(.dina(n8811), .dinb(n8807), .dout(n9024));
  jand g08832(.dina(n9024), .dinb(n9023), .dout(n9025));
  jnot g08833(.din(n9025), .dout(n9026));
  jnot g08834(.din(n8829), .dout(n9027));
  jor  g08835(.dina(n8836), .dinb(n9027), .dout(n9028));
  jnot g08836(.din(n8820), .dout(n9029));
  jand g08837(.dina(n8836), .dinb(n9027), .dout(n9030));
  jor  g08838(.dina(n9030), .dinb(n9029), .dout(n9031));
  jand g08839(.dina(n9031), .dinb(n9028), .dout(n9032));
  jxor g08840(.dina(n9032), .dinb(n9026), .dout(n9033));
  jand g08841(.dina(n8963), .dinb(n8955), .dout(n9034));
  jand g08842(.dina(n8967), .dinb(n8964), .dout(n9035));
  jor  g08843(.dina(n9035), .dinb(n9034), .dout(n9036));
  jxor g08844(.dina(n9036), .dinb(n9033), .dout(n9037));
  jand g08845(.dina(n8863), .dinb(n8688), .dout(n9038));
  jor  g08846(.dina(n9038), .dinb(n8861), .dout(n9039));
  jand g08847(.dina(n8843), .dinb(n8840), .dout(n9040));
  jor  g08848(.dina(n9040), .dinb(n8846), .dout(n9041));
  jxor g08849(.dina(n9041), .dinb(n9039), .dout(n9042));
  jand g08850(.dina(n8824), .dinb(n8821), .dout(n9043));
  jor  g08851(.dina(n9043), .dinb(n8827), .dout(n9044));
  jxor g08852(.dina(n9044), .dinb(n9042), .dout(n9045));
  jand g08853(.dina(n8835), .dinb(n8830), .dout(n9046));
  jor  g08854(.dina(n9046), .dinb(n8833), .dout(n9047));
  jand g08855(.dina(n8804), .dinb(n8670), .dout(n9048));
  jor  g08856(.dina(n9048), .dinb(n8802), .dout(n9049));
  jand g08857(.dina(n8791), .dinb(n8788), .dout(n9050));
  jor  g08858(.dina(n9050), .dinb(n8794), .dout(n9051));
  jxor g08859(.dina(n9051), .dinb(n9049), .dout(n9052));
  jxor g08860(.dina(n9052), .dinb(n9047), .dout(n9053));
  jnot g08861(.din(n8856), .dout(n9054));
  jor  g08862(.dina(n8864), .dinb(n9054), .dout(n9055));
  jnot g08863(.din(n8848), .dout(n9056));
  jand g08864(.dina(n8864), .dinb(n9054), .dout(n9057));
  jor  g08865(.dina(n9057), .dinb(n9056), .dout(n9058));
  jand g08866(.dina(n9058), .dinb(n9055), .dout(n9059));
  jxor g08867(.dina(n9059), .dinb(n9053), .dout(n9060));
  jxor g08868(.dina(n9060), .dinb(n9045), .dout(n9061));
  jxor g08869(.dina(n9061), .dinb(n9037), .dout(n9062));
  jxor g08870(.dina(n9062), .dinb(n9021), .dout(n9063));
  jxor g08871(.dina(n9063), .dinb(n9018), .dout(n9064));
  jxor g08872(.dina(n9064), .dinb(n8986), .dout(n9065));
  jand g08873(.dina(n8970), .dinb(n8935), .dout(n9066));
  jand g08874(.dina(n8971), .dinb(n8932), .dout(n9067));
  jor  g08875(.dina(n9067), .dinb(n9066), .dout(n9068));
  jand g08876(.dina(n8867), .dinb(n8787), .dout(n9069));
  jand g08877(.dina(n8868), .dinb(n8776), .dout(n9070));
  jor  g08878(.dina(n9070), .dinb(n9069), .dout(n9071));
  jxor g08879(.dina(n9071), .dinb(n9068), .dout(n9072));
  jand g08880(.dina(n8946), .dinb(n8941), .dout(n9073));
  jand g08881(.dina(n8951), .dinb(n8947), .dout(n9074));
  jor  g08882(.dina(n9074), .dinb(n9073), .dout(n9075));
  jand g08883(.dina(\a[42] ), .dinb(\a[27] ), .dout(n9076));
  jor  g08884(.dina(n9076), .dinb(n8817), .dout(n9077));
  jnot g08885(.din(n9077), .dout(n9078));
  jand g08886(.dina(\a[43] ), .dinb(\a[27] ), .dout(n9079));
  jand g08887(.dina(n9079), .dinb(n8814), .dout(n9080));
  jor  g08888(.dina(n9080), .dinb(n9078), .dout(n9081));
  jxor g08889(.dina(n9081), .dinb(n8845), .dout(n9082));
  jand g08890(.dina(\a[45] ), .dinb(\a[24] ), .dout(n9083));
  jand g08891(.dina(\a[44] ), .dinb(\a[25] ), .dout(n9084));
  jor  g08892(.dina(n9084), .dinb(n9083), .dout(n9085));
  jnot g08893(.din(n9085), .dout(n9086));
  jand g08894(.dina(\a[45] ), .dinb(\a[25] ), .dout(n9087));
  jand g08895(.dina(n9087), .dinb(n8680), .dout(n9088));
  jor  g08896(.dina(n9088), .dinb(n9086), .dout(n9089));
  jxor g08897(.dina(n9089), .dinb(n8826), .dout(n9090));
  jand g08898(.dina(\a[60] ), .dinb(\a[9] ), .dout(n9091));
  jand g08899(.dina(\a[59] ), .dinb(\a[10] ), .dout(n9092));
  jor  g08900(.dina(n9092), .dinb(n9091), .dout(n9093));
  jand g08901(.dina(\a[60] ), .dinb(\a[10] ), .dout(n9094));
  jand g08902(.dina(n9094), .dinb(n8688), .dout(n9095));
  jnot g08903(.din(n9095), .dout(n9096));
  jand g08904(.dina(n9096), .dinb(n9093), .dout(n9097));
  jxor g08905(.dina(n9097), .dinb(n8959), .dout(n9098));
  jxor g08906(.dina(n9098), .dinb(n9090), .dout(n9099));
  jxor g08907(.dina(n9099), .dinb(n9082), .dout(n9100));
  jxor g08908(.dina(n9100), .dinb(n9075), .dout(n9101));
  jand g08909(.dina(\a[55] ), .dinb(\a[14] ), .dout(n9102));
  jand g08910(.dina(\a[48] ), .dinb(\a[21] ), .dout(n9103));
  jand g08911(.dina(\a[47] ), .dinb(\a[22] ), .dout(n9104));
  jor  g08912(.dina(n9104), .dinb(n9103), .dout(n9105));
  jnot g08913(.din(n9105), .dout(n9106));
  jand g08914(.dina(\a[48] ), .dinb(\a[22] ), .dout(n9107));
  jand g08915(.dina(n9107), .dinb(n8840), .dout(n9108));
  jor  g08916(.dina(n9108), .dinb(n9106), .dout(n9109));
  jxor g08917(.dina(n9109), .dinb(n9102), .dout(n9110));
  jnot g08918(.din(n9110), .dout(n9111));
  jand g08919(.dina(\a[57] ), .dinb(\a[12] ), .dout(n9112));
  jand g08920(.dina(\a[56] ), .dinb(\a[13] ), .dout(n9113));
  jor  g08921(.dina(n9113), .dinb(n9112), .dout(n9114));
  jnot g08922(.din(n9114), .dout(n9115));
  jand g08923(.dina(\a[57] ), .dinb(\a[13] ), .dout(n9116));
  jand g08924(.dina(n9116), .dinb(n8808), .dout(n9117));
  jor  g08925(.dina(n9117), .dinb(n9115), .dout(n9118));
  jxor g08926(.dina(n9118), .dinb(n8860), .dout(n9119));
  jnot g08927(.din(n9119), .dout(n9120));
  jand g08928(.dina(n8962), .dinb(n8661), .dout(n9121));
  jor  g08929(.dina(n9121), .dinb(n8960), .dout(n9122));
  jxor g08930(.dina(n9122), .dinb(n9120), .dout(n9123));
  jxor g08931(.dina(n9123), .dinb(n9111), .dout(n9124));
  jxor g08932(.dina(n9124), .dinb(n9101), .dout(n9125));
  jand g08933(.dina(n8968), .dinb(n8952), .dout(n9126));
  jand g08934(.dina(n8969), .dinb(n8938), .dout(n9127));
  jor  g08935(.dina(n9127), .dinb(n9126), .dout(n9128));
  jor  g08936(.dina(n8903), .dinb(n8896), .dout(n9129));
  jand g08937(.dina(n8904), .dinb(n8892), .dout(n9130));
  jnot g08938(.din(n9130), .dout(n9131));
  jand g08939(.dina(n9131), .dinb(n9129), .dout(n9132));
  jnot g08940(.din(n9132), .dout(n9133));
  jand g08941(.dina(n8914), .dinb(n8912), .dout(n9134));
  jand g08942(.dina(n8915), .dinb(n8910), .dout(n9135));
  jor  g08943(.dina(n9135), .dinb(n9134), .dout(n9136));
  jand g08944(.dina(\a[41] ), .dinb(\a[28] ), .dout(n9137));
  jand g08945(.dina(\a[39] ), .dinb(\a[30] ), .dout(n9138));
  jor  g08946(.dina(n9138), .dinb(n8853), .dout(n9139));
  jnot g08947(.din(n9139), .dout(n9140));
  jand g08948(.dina(\a[40] ), .dinb(\a[30] ), .dout(n9141));
  jand g08949(.dina(n9141), .dinb(n8850), .dout(n9142));
  jor  g08950(.dina(n9142), .dinb(n9140), .dout(n9143));
  jxor g08951(.dina(n9143), .dinb(n9137), .dout(n9144));
  jnot g08952(.din(n9144), .dout(n9145));
  jor  g08953(.dina(n7343), .dinb(n6212), .dout(n9146));
  jand g08954(.dina(n6854), .dinb(n6356), .dout(n9147));
  jnot g08955(.din(n9147), .dout(n9148));
  jand g08956(.dina(n9148), .dinb(n9146), .dout(n9149));
  jxor g08957(.dina(n9149), .dinb(n8801), .dout(n9150));
  jxor g08958(.dina(n9150), .dinb(n9145), .dout(n9151));
  jxor g08959(.dina(n9151), .dinb(n9136), .dout(n9152));
  jand g08960(.dina(\a[54] ), .dinb(\a[15] ), .dout(n9153));
  jnot g08961(.din(n9153), .dout(n9154));
  jand g08962(.dina(\a[49] ), .dinb(\a[20] ), .dout(n9155));
  jxor g08963(.dina(n9155), .dinb(n8832), .dout(n9156));
  jxor g08964(.dina(n9156), .dinb(n9154), .dout(n9157));
  jnot g08965(.din(n9157), .dout(n9158));
  jand g08966(.dina(\a[38] ), .dinb(\a[31] ), .dout(n9159));
  jnot g08967(.din(n9159), .dout(n9160));
  jand g08968(.dina(\a[36] ), .dinb(\a[33] ), .dout(n9161));
  jor  g08969(.dina(n9161), .dinb(n8793), .dout(n9162));
  jand g08970(.dina(\a[37] ), .dinb(\a[33] ), .dout(n9163));
  jand g08971(.dina(n9163), .dinb(n8790), .dout(n9164));
  jnot g08972(.din(n9164), .dout(n9165));
  jand g08973(.dina(n9165), .dinb(n9162), .dout(n9166));
  jxor g08974(.dina(n9166), .dinb(n9160), .dout(n9167));
  jand g08975(.dina(\a[62] ), .dinb(\a[7] ), .dout(n9168));
  jnot g08976(.din(n9168), .dout(n9169));
  jand g08977(.dina(\a[35] ), .dinb(n8652), .dout(n9170));
  jxor g08978(.dina(n9170), .dinb(n9169), .dout(n9171));
  jxor g08979(.dina(n9171), .dinb(n9167), .dout(n9172));
  jxor g08980(.dina(n9172), .dinb(n9158), .dout(n9173));
  jxor g08981(.dina(n9173), .dinb(n9152), .dout(n9174));
  jxor g08982(.dina(n9174), .dinb(n9133), .dout(n9175));
  jxor g08983(.dina(n9175), .dinb(n9128), .dout(n9176));
  jxor g08984(.dina(n9176), .dinb(n9125), .dout(n9177));
  jxor g08985(.dina(n9177), .dinb(n9072), .dout(n9178));
  jxor g08986(.dina(n9178), .dinb(n9065), .dout(n9179));
  jxor g08987(.dina(n9179), .dinb(n8983), .dout(n9180));
  jand g08988(.dina(n8974), .dinb(n8767), .dout(n9181));
  jnot g08989(.din(n8767), .dout(n9182));
  jnot g08990(.din(n8974), .dout(n9183));
  jand g08991(.dina(n9183), .dinb(n9182), .dout(n9184));
  jnot g08992(.din(n9184), .dout(n9185));
  jand g08993(.dina(n8979), .dinb(n9185), .dout(n9186));
  jor  g08994(.dina(n9186), .dinb(n9181), .dout(n9187));
  jxor g08995(.dina(n9187), .dinb(n9180), .dout(\asquared[70] ));
  jand g08996(.dina(n9064), .dinb(n8986), .dout(n9189));
  jand g08997(.dina(n9178), .dinb(n9065), .dout(n9190));
  jor  g08998(.dina(n9190), .dinb(n9189), .dout(n9191));
  jand g08999(.dina(n9017), .dinb(n8989), .dout(n9192));
  jand g09000(.dina(n9063), .dinb(n9018), .dout(n9193));
  jor  g09001(.dina(n9193), .dinb(n9192), .dout(n9194));
  jand g09002(.dina(n9150), .dinb(n9145), .dout(n9195));
  jand g09003(.dina(n9151), .dinb(n9136), .dout(n9196));
  jor  g09004(.dina(n9196), .dinb(n9195), .dout(n9197));
  jand g09005(.dina(n9077), .dinb(n8845), .dout(n9198));
  jor  g09006(.dina(n9198), .dinb(n9080), .dout(n9199));
  jand g09007(.dina(n9139), .dinb(n9137), .dout(n9200));
  jor  g09008(.dina(n9200), .dinb(n9142), .dout(n9201));
  jxor g09009(.dina(n9201), .dinb(n9199), .dout(n9202));
  jand g09010(.dina(n9085), .dinb(n8826), .dout(n9203));
  jor  g09011(.dina(n9203), .dinb(n9088), .dout(n9204));
  jxor g09012(.dina(n9204), .dinb(n9202), .dout(n9205));
  jand g09013(.dina(\a[62] ), .dinb(\a[8] ), .dout(n9206));
  jnot g09014(.din(\a[35] ), .dout(n9207));
  jand g09015(.dina(n9169), .dinb(n8652), .dout(n9208));
  jor  g09016(.dina(n9208), .dinb(n9207), .dout(n9209));
  jnot g09017(.din(n9209), .dout(n9210));
  jxor g09018(.dina(n9210), .dinb(n9206), .dout(n9211));
  jand g09019(.dina(n9162), .dinb(n9159), .dout(n9212));
  jor  g09020(.dina(n9212), .dinb(n9164), .dout(n9213));
  jxor g09021(.dina(n9213), .dinb(n9211), .dout(n9214));
  jxor g09022(.dina(n9214), .dinb(n9205), .dout(n9215));
  jxor g09023(.dina(n9215), .dinb(n9197), .dout(n9216));
  jand g09024(.dina(n9173), .dinb(n9152), .dout(n9217));
  jand g09025(.dina(n9174), .dinb(n9133), .dout(n9218));
  jor  g09026(.dina(n9218), .dinb(n9217), .dout(n9219));
  jand g09027(.dina(n9122), .dinb(n9120), .dout(n9220));
  jand g09028(.dina(n9123), .dinb(n9111), .dout(n9221));
  jor  g09029(.dina(n9221), .dinb(n9220), .dout(n9222));
  jnot g09030(.din(n9090), .dout(n9223));
  jor  g09031(.dina(n9098), .dinb(n9223), .dout(n9224));
  jnot g09032(.din(n9082), .dout(n9225));
  jand g09033(.dina(n9098), .dinb(n9223), .dout(n9226));
  jor  g09034(.dina(n9226), .dinb(n9225), .dout(n9227));
  jand g09035(.dina(n9227), .dinb(n9224), .dout(n9228));
  jxor g09036(.dina(n9228), .dinb(n9222), .dout(n9229));
  jand g09037(.dina(n9171), .dinb(n9167), .dout(n9230));
  jnot g09038(.din(n9230), .dout(n9231));
  jnot g09039(.din(n9167), .dout(n9232));
  jnot g09040(.din(n9171), .dout(n9233));
  jand g09041(.dina(n9233), .dinb(n9232), .dout(n9234));
  jor  g09042(.dina(n9234), .dinb(n9158), .dout(n9235));
  jand g09043(.dina(n9235), .dinb(n9231), .dout(n9236));
  jxor g09044(.dina(n9236), .dinb(n9229), .dout(n9237));
  jxor g09045(.dina(n9237), .dinb(n9219), .dout(n9238));
  jxor g09046(.dina(n9238), .dinb(n9216), .dout(n9239));
  jxor g09047(.dina(n9239), .dinb(n9194), .dout(n9240));
  jand g09048(.dina(n9015), .dinb(n8995), .dout(n9241));
  jand g09049(.dina(n9016), .dinb(n8992), .dout(n9242));
  jor  g09050(.dina(n9242), .dinb(n9241), .dout(n9243));
  jand g09051(.dina(n9013), .dinb(n9010), .dout(n9244));
  jand g09052(.dina(n9014), .dinb(n9007), .dout(n9245));
  jor  g09053(.dina(n9245), .dinb(n9244), .dout(n9246));
  jand g09054(.dina(n9149), .dinb(n8801), .dout(n9247));
  jor  g09055(.dina(n9247), .dinb(n9147), .dout(n9248));
  jnot g09056(.din(n9248), .dout(n9249));
  jand g09057(.dina(n9155), .dinb(n8832), .dout(n9250));
  jnot g09058(.din(n9250), .dout(n9251));
  jnot g09059(.din(n8832), .dout(n9252));
  jnot g09060(.din(n9155), .dout(n9253));
  jand g09061(.dina(n9253), .dinb(n9252), .dout(n9254));
  jor  g09062(.dina(n9254), .dinb(n9154), .dout(n9255));
  jand g09063(.dina(n9255), .dinb(n9251), .dout(n9256));
  jxor g09064(.dina(n9256), .dinb(n9249), .dout(n9257));
  jand g09065(.dina(\a[38] ), .dinb(\a[32] ), .dout(n9258));
  jnot g09066(.din(n9258), .dout(n9259));
  jand g09067(.dina(\a[36] ), .dinb(\a[34] ), .dout(n9260));
  jor  g09068(.dina(n9260), .dinb(n9163), .dout(n9261));
  jand g09069(.dina(\a[37] ), .dinb(\a[34] ), .dout(n9262));
  jand g09070(.dina(n9262), .dinb(n9161), .dout(n9263));
  jnot g09071(.din(n9263), .dout(n9264));
  jand g09072(.dina(n9264), .dinb(n9261), .dout(n9265));
  jxor g09073(.dina(n9265), .dinb(n9259), .dout(n9266));
  jnot g09074(.din(n9266), .dout(n9267));
  jxor g09075(.dina(n9267), .dinb(n9257), .dout(n9268));
  jxor g09076(.dina(n9268), .dinb(n9246), .dout(n9269));
  jand g09077(.dina(\a[58] ), .dinb(\a[12] ), .dout(n9270));
  jor  g09078(.dina(n9116), .dinb(n4351), .dout(n9271));
  jnot g09079(.din(n9271), .dout(n9272));
  jand g09080(.dina(n8326), .dinb(n6371), .dout(n9273));
  jor  g09081(.dina(n9273), .dinb(n9272), .dout(n9274));
  jxor g09082(.dina(n9274), .dinb(n9270), .dout(n9275));
  jand g09083(.dina(\a[53] ), .dinb(\a[17] ), .dout(n9276));
  jand g09084(.dina(\a[54] ), .dinb(\a[16] ), .dout(n9277));
  jor  g09085(.dina(n9277), .dinb(n9276), .dout(n9278));
  jnot g09086(.din(n9278), .dout(n9279));
  jand g09087(.dina(n8832), .dinb(n7804), .dout(n9280));
  jor  g09088(.dina(n9280), .dinb(n9279), .dout(n9281));
  jxor g09089(.dina(n9281), .dinb(n6854), .dout(n9282));
  jand g09090(.dina(\a[61] ), .dinb(\a[9] ), .dout(n9283));
  jand g09091(.dina(\a[59] ), .dinb(\a[11] ), .dout(n9284));
  jor  g09092(.dina(n9284), .dinb(n9094), .dout(n9285));
  jand g09093(.dina(\a[60] ), .dinb(\a[11] ), .dout(n9286));
  jand g09094(.dina(n9286), .dinb(n9092), .dout(n9287));
  jnot g09095(.din(n9287), .dout(n9288));
  jand g09096(.dina(n9288), .dinb(n9285), .dout(n9289));
  jxor g09097(.dina(n9289), .dinb(n9283), .dout(n9290));
  jxor g09098(.dina(n9290), .dinb(n9282), .dout(n9291));
  jxor g09099(.dina(n9291), .dinb(n9275), .dout(n9292));
  jxor g09100(.dina(n9292), .dinb(n9269), .dout(n9293));
  jxor g09101(.dina(n9293), .dinb(n9243), .dout(n9294));
  jand g09102(.dina(n9059), .dinb(n9053), .dout(n9295));
  jand g09103(.dina(n9060), .dinb(n9045), .dout(n9296));
  jor  g09104(.dina(n9296), .dinb(n9295), .dout(n9297));
  jand g09105(.dina(n9051), .dinb(n9049), .dout(n9298));
  jand g09106(.dina(n9052), .dinb(n9047), .dout(n9299));
  jor  g09107(.dina(n9299), .dinb(n9298), .dout(n9300));
  jand g09108(.dina(\a[41] ), .dinb(\a[29] ), .dout(n9301));
  jand g09109(.dina(\a[39] ), .dinb(\a[31] ), .dout(n9302));
  jor  g09110(.dina(n9302), .dinb(n9141), .dout(n9303));
  jnot g09111(.din(n9303), .dout(n9304));
  jand g09112(.dina(\a[40] ), .dinb(\a[31] ), .dout(n9305));
  jand g09113(.dina(n9305), .dinb(n9138), .dout(n9306));
  jor  g09114(.dina(n9306), .dinb(n9304), .dout(n9307));
  jxor g09115(.dina(n9307), .dinb(n9301), .dout(n9308));
  jand g09116(.dina(\a[42] ), .dinb(\a[28] ), .dout(n9309));
  jand g09117(.dina(\a[47] ), .dinb(\a[23] ), .dout(n9310));
  jnot g09118(.din(n9310), .dout(n9311));
  jand g09119(.dina(\a[63] ), .dinb(\a[7] ), .dout(n9312));
  jxor g09120(.dina(n9312), .dinb(n9311), .dout(n9313));
  jxor g09121(.dina(n9313), .dinb(n9309), .dout(n9314));
  jxor g09122(.dina(n9314), .dinb(n9308), .dout(n9315));
  jxor g09123(.dina(n9315), .dinb(n9300), .dout(n9316));
  jand g09124(.dina(\a[49] ), .dinb(\a[21] ), .dout(n9317));
  jand g09125(.dina(\a[51] ), .dinb(\a[19] ), .dout(n9318));
  jand g09126(.dina(\a[50] ), .dinb(\a[20] ), .dout(n9319));
  jor  g09127(.dina(n9319), .dinb(n9318), .dout(n9320));
  jnot g09128(.din(n9320), .dout(n9321));
  jand g09129(.dina(\a[51] ), .dinb(\a[20] ), .dout(n9322));
  jand g09130(.dina(n9322), .dinb(n8801), .dout(n9323));
  jor  g09131(.dina(n9323), .dinb(n9321), .dout(n9324));
  jxor g09132(.dina(n9324), .dinb(n9317), .dout(n9325));
  jand g09133(.dina(\a[44] ), .dinb(\a[26] ), .dout(n9326));
  jor  g09134(.dina(n9326), .dinb(n9079), .dout(n9327));
  jnot g09135(.din(n9327), .dout(n9328));
  jand g09136(.dina(\a[44] ), .dinb(\a[27] ), .dout(n9329));
  jand g09137(.dina(n9329), .dinb(n8817), .dout(n9330));
  jor  g09138(.dina(n9330), .dinb(n9328), .dout(n9331));
  jxor g09139(.dina(n9331), .dinb(n9087), .dout(n9332));
  jand g09140(.dina(\a[56] ), .dinb(\a[14] ), .dout(n9333));
  jand g09141(.dina(\a[55] ), .dinb(\a[15] ), .dout(n9334));
  jor  g09142(.dina(n9334), .dinb(n9333), .dout(n9335));
  jand g09143(.dina(\a[56] ), .dinb(\a[15] ), .dout(n9336));
  jand g09144(.dina(n9336), .dinb(n9102), .dout(n9337));
  jnot g09145(.din(n9337), .dout(n9338));
  jand g09146(.dina(n9338), .dinb(n9335), .dout(n9339));
  jxor g09147(.dina(n9339), .dinb(n9107), .dout(n9340));
  jxor g09148(.dina(n9340), .dinb(n9332), .dout(n9341));
  jxor g09149(.dina(n9341), .dinb(n9325), .dout(n9342));
  jxor g09150(.dina(n9342), .dinb(n9316), .dout(n9343));
  jxor g09151(.dina(n9343), .dinb(n9297), .dout(n9344));
  jxor g09152(.dina(n9344), .dinb(n9294), .dout(n9345));
  jxor g09153(.dina(n9345), .dinb(n9240), .dout(n9346));
  jand g09154(.dina(n9175), .dinb(n9128), .dout(n9347));
  jand g09155(.dina(n9176), .dinb(n9125), .dout(n9348));
  jor  g09156(.dina(n9348), .dinb(n9347), .dout(n9349));
  jand g09157(.dina(n9061), .dinb(n9037), .dout(n9350));
  jand g09158(.dina(n9062), .dinb(n9021), .dout(n9351));
  jor  g09159(.dina(n9351), .dinb(n9350), .dout(n9352));
  jand g09160(.dina(n9100), .dinb(n9075), .dout(n9353));
  jand g09161(.dina(n9124), .dinb(n9101), .dout(n9354));
  jor  g09162(.dina(n9354), .dinb(n9353), .dout(n9355));
  jand g09163(.dina(n9032), .dinb(n9026), .dout(n9356));
  jand g09164(.dina(n9036), .dinb(n9033), .dout(n9357));
  jor  g09165(.dina(n9357), .dinb(n9356), .dout(n9358));
  jand g09166(.dina(n9097), .dinb(n8959), .dout(n9359));
  jor  g09167(.dina(n9359), .dinb(n9095), .dout(n9360));
  jand g09168(.dina(n9114), .dinb(n8860), .dout(n9361));
  jor  g09169(.dina(n9361), .dinb(n9117), .dout(n9362));
  jxor g09170(.dina(n9362), .dinb(n9360), .dout(n9363));
  jand g09171(.dina(n9105), .dinb(n9102), .dout(n9364));
  jor  g09172(.dina(n9364), .dinb(n9108), .dout(n9365));
  jxor g09173(.dina(n9365), .dinb(n9363), .dout(n9366));
  jand g09174(.dina(n9041), .dinb(n9039), .dout(n9367));
  jand g09175(.dina(n9044), .dinb(n9042), .dout(n9368));
  jor  g09176(.dina(n9368), .dinb(n9367), .dout(n9369));
  jand g09177(.dina(n9003), .dinb(n8997), .dout(n9370));
  jand g09178(.dina(n9006), .dinb(n9004), .dout(n9371));
  jor  g09179(.dina(n9371), .dinb(n9370), .dout(n9372));
  jxor g09180(.dina(n9372), .dinb(n9369), .dout(n9373));
  jxor g09181(.dina(n9373), .dinb(n9366), .dout(n9374));
  jxor g09182(.dina(n9374), .dinb(n9358), .dout(n9375));
  jxor g09183(.dina(n9375), .dinb(n9355), .dout(n9376));
  jxor g09184(.dina(n9376), .dinb(n9352), .dout(n9377));
  jxor g09185(.dina(n9377), .dinb(n9349), .dout(n9378));
  jand g09186(.dina(n9071), .dinb(n9068), .dout(n9379));
  jand g09187(.dina(n9177), .dinb(n9072), .dout(n9380));
  jor  g09188(.dina(n9380), .dinb(n9379), .dout(n9381));
  jxor g09189(.dina(n9381), .dinb(n9378), .dout(n9382));
  jxor g09190(.dina(n9382), .dinb(n9346), .dout(n9383));
  jxor g09191(.dina(n9383), .dinb(n9191), .dout(n9384));
  jand g09192(.dina(n9179), .dinb(n8983), .dout(n9385));
  jor  g09193(.dina(n9179), .dinb(n8983), .dout(n9386));
  jand g09194(.dina(n9187), .dinb(n9386), .dout(n9387));
  jor  g09195(.dina(n9387), .dinb(n9385), .dout(n9388));
  jxor g09196(.dina(n9388), .dinb(n9384), .dout(\asquared[71] ));
  jand g09197(.dina(n9381), .dinb(n9378), .dout(n9390));
  jand g09198(.dina(n9382), .dinb(n9346), .dout(n9391));
  jor  g09199(.dina(n9391), .dinb(n9390), .dout(n9392));
  jand g09200(.dina(n9293), .dinb(n9243), .dout(n9393));
  jand g09201(.dina(n9344), .dinb(n9294), .dout(n9394));
  jor  g09202(.dina(n9394), .dinb(n9393), .dout(n9395));
  jand g09203(.dina(n9210), .dinb(n9206), .dout(n9396));
  jand g09204(.dina(n9213), .dinb(n9211), .dout(n9397));
  jor  g09205(.dina(n9397), .dinb(n9396), .dout(n9398));
  jand g09206(.dina(n9256), .dinb(n9249), .dout(n9399));
  jor  g09207(.dina(n9256), .dinb(n9249), .dout(n9400));
  jand g09208(.dina(n9266), .dinb(n9400), .dout(n9401));
  jor  g09209(.dina(n9401), .dinb(n9399), .dout(n9402));
  jnot g09210(.din(n9402), .dout(n9403));
  jxor g09211(.dina(n9403), .dinb(n9398), .dout(n9404));
  jand g09212(.dina(n9201), .dinb(n9199), .dout(n9405));
  jand g09213(.dina(n9204), .dinb(n9202), .dout(n9406));
  jor  g09214(.dina(n9406), .dinb(n9405), .dout(n9407));
  jxor g09215(.dina(n9407), .dinb(n9404), .dout(n9408));
  jand g09216(.dina(n9214), .dinb(n9205), .dout(n9409));
  jand g09217(.dina(n9215), .dinb(n9197), .dout(n9410));
  jor  g09218(.dina(n9410), .dinb(n9409), .dout(n9411));
  jxor g09219(.dina(n9411), .dinb(n9408), .dout(n9412));
  jand g09220(.dina(n9268), .dinb(n9246), .dout(n9413));
  jand g09221(.dina(n9292), .dinb(n9269), .dout(n9414));
  jor  g09222(.dina(n9414), .dinb(n9413), .dout(n9415));
  jxor g09223(.dina(n9415), .dinb(n9412), .dout(n9416));
  jand g09224(.dina(n9237), .dinb(n9219), .dout(n9417));
  jand g09225(.dina(n9238), .dinb(n9216), .dout(n9418));
  jor  g09226(.dina(n9418), .dinb(n9417), .dout(n9419));
  jxor g09227(.dina(n9419), .dinb(n9416), .dout(n9420));
  jxor g09228(.dina(n9420), .dinb(n9395), .dout(n9421));
  jand g09229(.dina(n9239), .dinb(n9194), .dout(n9422));
  jand g09230(.dina(n9345), .dinb(n9240), .dout(n9423));
  jor  g09231(.dina(n9423), .dinb(n9422), .dout(n9424));
  jxor g09232(.dina(n9424), .dinb(n9421), .dout(n9425));
  jand g09233(.dina(n9376), .dinb(n9352), .dout(n9426));
  jand g09234(.dina(n9377), .dinb(n9349), .dout(n9427));
  jor  g09235(.dina(n9427), .dinb(n9426), .dout(n9428));
  jand g09236(.dina(n9342), .dinb(n9316), .dout(n9429));
  jand g09237(.dina(n9343), .dinb(n9297), .dout(n9430));
  jor  g09238(.dina(n9430), .dinb(n9429), .dout(n9431));
  jand g09239(.dina(n9362), .dinb(n9360), .dout(n9432));
  jand g09240(.dina(n9365), .dinb(n9363), .dout(n9433));
  jor  g09241(.dina(n9433), .dinb(n9432), .dout(n9434));
  jnot g09242(.din(n9282), .dout(n9435));
  jor  g09243(.dina(n9290), .dinb(n9435), .dout(n9436));
  jnot g09244(.din(n9275), .dout(n9437));
  jand g09245(.dina(n9290), .dinb(n9435), .dout(n9438));
  jor  g09246(.dina(n9438), .dinb(n9437), .dout(n9439));
  jand g09247(.dina(n9439), .dinb(n9436), .dout(n9440));
  jxor g09248(.dina(n9440), .dinb(n9434), .dout(n9441));
  jnot g09249(.din(n9332), .dout(n9442));
  jor  g09250(.dina(n9340), .dinb(n9442), .dout(n9443));
  jnot g09251(.din(n9325), .dout(n9444));
  jand g09252(.dina(n9340), .dinb(n9442), .dout(n9445));
  jor  g09253(.dina(n9445), .dinb(n9444), .dout(n9446));
  jand g09254(.dina(n9446), .dinb(n9443), .dout(n9447));
  jxor g09255(.dina(n9447), .dinb(n9441), .dout(n9448));
  jxor g09256(.dina(n9448), .dinb(n9431), .dout(n9449));
  jor  g09257(.dina(n9314), .dinb(n9308), .dout(n9450));
  jand g09258(.dina(n9315), .dinb(n9300), .dout(n9451));
  jnot g09259(.din(n9451), .dout(n9452));
  jand g09260(.dina(n9452), .dinb(n9450), .dout(n9453));
  jnot g09261(.din(n9453), .dout(n9454));
  jand g09262(.dina(n9289), .dinb(n9283), .dout(n9455));
  jor  g09263(.dina(n9455), .dinb(n9287), .dout(n9456));
  jand g09264(.dina(n9271), .dinb(n9270), .dout(n9457));
  jor  g09265(.dina(n9457), .dinb(n9273), .dout(n9458));
  jxor g09266(.dina(n9458), .dinb(n9456), .dout(n9459));
  jand g09267(.dina(n9327), .dinb(n9087), .dout(n9460));
  jor  g09268(.dina(n9460), .dinb(n9330), .dout(n9461));
  jxor g09269(.dina(n9461), .dinb(n9459), .dout(n9462));
  jand g09270(.dina(n9339), .dinb(n9107), .dout(n9463));
  jor  g09271(.dina(n9463), .dinb(n9337), .dout(n9464));
  jand g09272(.dina(n9303), .dinb(n9301), .dout(n9465));
  jor  g09273(.dina(n9465), .dinb(n9306), .dout(n9466));
  jxor g09274(.dina(n9466), .dinb(n9464), .dout(n9467));
  jnot g09275(.din(n9312), .dout(n9468));
  jand g09276(.dina(n9468), .dinb(n9311), .dout(n9469));
  jnot g09277(.din(n9469), .dout(n9470));
  jand g09278(.dina(n9312), .dinb(n9310), .dout(n9471));
  jor  g09279(.dina(n9471), .dinb(n9309), .dout(n9472));
  jand g09280(.dina(n9472), .dinb(n9470), .dout(n9473));
  jxor g09281(.dina(n9473), .dinb(n9467), .dout(n9474));
  jxor g09282(.dina(n9474), .dinb(n9462), .dout(n9475));
  jxor g09283(.dina(n9475), .dinb(n9454), .dout(n9476));
  jxor g09284(.dina(n9476), .dinb(n9449), .dout(n9477));
  jxor g09285(.dina(n9477), .dinb(n9428), .dout(n9478));
  jand g09286(.dina(n9374), .dinb(n9358), .dout(n9479));
  jand g09287(.dina(n9375), .dinb(n9355), .dout(n9480));
  jor  g09288(.dina(n9480), .dinb(n9479), .dout(n9481));
  jand g09289(.dina(n9372), .dinb(n9369), .dout(n9482));
  jand g09290(.dina(n9373), .dinb(n9366), .dout(n9483));
  jor  g09291(.dina(n9483), .dinb(n9482), .dout(n9484));
  jand g09292(.dina(n9278), .dinb(n6854), .dout(n9485));
  jor  g09293(.dina(n9485), .dinb(n9280), .dout(n9486));
  jand g09294(.dina(n9261), .dinb(n9258), .dout(n9487));
  jor  g09295(.dina(n9487), .dinb(n9263), .dout(n9488));
  jxor g09296(.dina(n9488), .dinb(n9486), .dout(n9489));
  jand g09297(.dina(\a[63] ), .dinb(\a[8] ), .dout(n9490));
  jand g09298(.dina(\a[61] ), .dinb(\a[10] ), .dout(n9491));
  jor  g09299(.dina(n9491), .dinb(n9490), .dout(n9492));
  jnot g09300(.din(n9492), .dout(n9493));
  jand g09301(.dina(\a[63] ), .dinb(\a[10] ), .dout(n9494));
  jand g09302(.dina(n9494), .dinb(n8959), .dout(n9495));
  jor  g09303(.dina(n9495), .dinb(n9493), .dout(n9496));
  jxor g09304(.dina(n9496), .dinb(n9286), .dout(n9497));
  jnot g09305(.din(n9497), .dout(n9498));
  jxor g09306(.dina(n9498), .dinb(n9489), .dout(n9499));
  jxor g09307(.dina(n9499), .dinb(n9484), .dout(n9500));
  jand g09308(.dina(\a[50] ), .dinb(\a[21] ), .dout(n9501));
  jand g09309(.dina(\a[52] ), .dinb(\a[19] ), .dout(n9502));
  jor  g09310(.dina(n9502), .dinb(n9322), .dout(n9503));
  jnot g09311(.din(n9503), .dout(n9504));
  jand g09312(.dina(\a[52] ), .dinb(\a[20] ), .dout(n9505));
  jand g09313(.dina(n9505), .dinb(n9318), .dout(n9506));
  jor  g09314(.dina(n9506), .dinb(n9504), .dout(n9507));
  jxor g09315(.dina(n9507), .dinb(n9501), .dout(n9508));
  jand g09316(.dina(\a[49] ), .dinb(\a[22] ), .dout(n9509));
  jnot g09317(.din(n9509), .dout(n9510));
  jand g09318(.dina(\a[62] ), .dinb(\a[9] ), .dout(n9511));
  jor  g09319(.dina(n9511), .dinb(\a[36] ), .dout(n9512));
  jand g09320(.dina(\a[62] ), .dinb(\a[36] ), .dout(n9513));
  jand g09321(.dina(n9513), .dinb(\a[9] ), .dout(n9514));
  jnot g09322(.din(n9514), .dout(n9515));
  jand g09323(.dina(n9515), .dinb(n9512), .dout(n9516));
  jor  g09324(.dina(n9516), .dinb(n9510), .dout(n9517));
  jand g09325(.dina(n9512), .dinb(n9509), .dout(n9518));
  jor  g09326(.dina(n9518), .dinb(n9514), .dout(n9519));
  jnot g09327(.din(n9519), .dout(n9520));
  jand g09328(.dina(n9520), .dinb(n9512), .dout(n9521));
  jnot g09329(.din(n9521), .dout(n9522));
  jand g09330(.dina(n9522), .dinb(n9517), .dout(n9523));
  jxor g09331(.dina(n9523), .dinb(n9508), .dout(n9524));
  jnot g09332(.din(n9524), .dout(n9525));
  jand g09333(.dina(\a[38] ), .dinb(\a[33] ), .dout(n9526));
  jnot g09334(.din(n9262), .dout(n9527));
  jand g09335(.dina(\a[36] ), .dinb(\a[35] ), .dout(n9528));
  jxor g09336(.dina(n9528), .dinb(n9527), .dout(n9529));
  jxor g09337(.dina(n9529), .dinb(n9526), .dout(n9530));
  jxor g09338(.dina(n9530), .dinb(n9525), .dout(n9531));
  jxor g09339(.dina(n9531), .dinb(n9500), .dout(n9532));
  jxor g09340(.dina(n9532), .dinb(n9481), .dout(n9533));
  jand g09341(.dina(n9228), .dinb(n9222), .dout(n9534));
  jand g09342(.dina(n9236), .dinb(n9229), .dout(n9535));
  jor  g09343(.dina(n9535), .dinb(n9534), .dout(n9536));
  jand g09344(.dina(\a[58] ), .dinb(\a[13] ), .dout(n9537));
  jand g09345(.dina(\a[59] ), .dinb(\a[12] ), .dout(n9538));
  jor  g09346(.dina(n9538), .dinb(n9537), .dout(n9539));
  jand g09347(.dina(\a[59] ), .dinb(\a[13] ), .dout(n9540));
  jand g09348(.dina(n9540), .dinb(n9270), .dout(n9541));
  jnot g09349(.din(n9541), .dout(n9542));
  jand g09350(.dina(n9542), .dinb(n9539), .dout(n9543));
  jand g09351(.dina(n9320), .dinb(n9317), .dout(n9544));
  jor  g09352(.dina(n9544), .dinb(n9323), .dout(n9545));
  jxor g09353(.dina(n9545), .dinb(n9543), .dout(n9546));
  jand g09354(.dina(\a[47] ), .dinb(\a[24] ), .dout(n9547));
  jand g09355(.dina(\a[46] ), .dinb(\a[25] ), .dout(n9548));
  jand g09356(.dina(\a[45] ), .dinb(\a[26] ), .dout(n9549));
  jor  g09357(.dina(n9549), .dinb(n9548), .dout(n9550));
  jnot g09358(.din(n9550), .dout(n9551));
  jand g09359(.dina(\a[46] ), .dinb(\a[26] ), .dout(n9552));
  jand g09360(.dina(n9552), .dinb(n9087), .dout(n9553));
  jor  g09361(.dina(n9553), .dinb(n9551), .dout(n9554));
  jxor g09362(.dina(n9554), .dinb(n9547), .dout(n9555));
  jnot g09363(.din(n9555), .dout(n9556));
  jand g09364(.dina(\a[57] ), .dinb(\a[14] ), .dout(n9557));
  jand g09365(.dina(\a[55] ), .dinb(\a[16] ), .dout(n9558));
  jor  g09366(.dina(n9558), .dinb(n9336), .dout(n9559));
  jand g09367(.dina(n9334), .dinb(n7946), .dout(n9560));
  jnot g09368(.din(n9560), .dout(n9561));
  jand g09369(.dina(n9561), .dinb(n9559), .dout(n9562));
  jxor g09370(.dina(n9562), .dinb(n9557), .dout(n9563));
  jxor g09371(.dina(n9563), .dinb(n9556), .dout(n9564));
  jxor g09372(.dina(n9564), .dinb(n9546), .dout(n9565));
  jand g09373(.dina(\a[48] ), .dinb(\a[23] ), .dout(n9566));
  jand g09374(.dina(\a[53] ), .dinb(\a[18] ), .dout(n9567));
  jor  g09375(.dina(n9567), .dinb(n7804), .dout(n9568));
  jnot g09376(.din(n9568), .dout(n9569));
  jand g09377(.dina(n9276), .dinb(n7507), .dout(n9570));
  jor  g09378(.dina(n9570), .dinb(n9569), .dout(n9571));
  jxor g09379(.dina(n9571), .dinb(n9566), .dout(n9572));
  jand g09380(.dina(\a[41] ), .dinb(\a[30] ), .dout(n9573));
  jand g09381(.dina(\a[39] ), .dinb(\a[32] ), .dout(n9574));
  jor  g09382(.dina(n9574), .dinb(n9305), .dout(n9575));
  jnot g09383(.din(n9575), .dout(n9576));
  jand g09384(.dina(\a[40] ), .dinb(\a[32] ), .dout(n9577));
  jand g09385(.dina(n9577), .dinb(n9302), .dout(n9578));
  jor  g09386(.dina(n9578), .dinb(n9576), .dout(n9579));
  jxor g09387(.dina(n9579), .dinb(n9573), .dout(n9580));
  jand g09388(.dina(\a[43] ), .dinb(\a[28] ), .dout(n9581));
  jand g09389(.dina(\a[42] ), .dinb(\a[29] ), .dout(n9582));
  jor  g09390(.dina(n9582), .dinb(n9581), .dout(n9583));
  jand g09391(.dina(\a[43] ), .dinb(\a[29] ), .dout(n9584));
  jand g09392(.dina(n9584), .dinb(n9309), .dout(n9585));
  jnot g09393(.din(n9585), .dout(n9586));
  jand g09394(.dina(n9586), .dinb(n9583), .dout(n9587));
  jxor g09395(.dina(n9587), .dinb(n9329), .dout(n9588));
  jxor g09396(.dina(n9588), .dinb(n9580), .dout(n9589));
  jxor g09397(.dina(n9589), .dinb(n9572), .dout(n9590));
  jxor g09398(.dina(n9590), .dinb(n9565), .dout(n9591));
  jxor g09399(.dina(n9591), .dinb(n9536), .dout(n9592));
  jxor g09400(.dina(n9592), .dinb(n9533), .dout(n9593));
  jxor g09401(.dina(n9593), .dinb(n9478), .dout(n9594));
  jxor g09402(.dina(n9594), .dinb(n9425), .dout(n9595));
  jxor g09403(.dina(n9595), .dinb(n9392), .dout(n9596));
  jand g09404(.dina(n9383), .dinb(n9191), .dout(n9597));
  jnot g09405(.din(n9191), .dout(n9598));
  jnot g09406(.din(n9383), .dout(n9599));
  jand g09407(.dina(n9599), .dinb(n9598), .dout(n9600));
  jnot g09408(.din(n9600), .dout(n9601));
  jand g09409(.dina(n9388), .dinb(n9601), .dout(n9602));
  jor  g09410(.dina(n9602), .dinb(n9597), .dout(n9603));
  jxor g09411(.dina(n9603), .dinb(n9596), .dout(\asquared[72] ));
  jand g09412(.dina(n9532), .dinb(n9481), .dout(n9605));
  jand g09413(.dina(n9592), .dinb(n9533), .dout(n9606));
  jor  g09414(.dina(n9606), .dinb(n9605), .dout(n9607));
  jand g09415(.dina(n9474), .dinb(n9462), .dout(n9608));
  jand g09416(.dina(n9475), .dinb(n9454), .dout(n9609));
  jor  g09417(.dina(n9609), .dinb(n9608), .dout(n9610));
  jand g09418(.dina(n9466), .dinb(n9464), .dout(n9611));
  jand g09419(.dina(n9473), .dinb(n9467), .dout(n9612));
  jor  g09420(.dina(n9612), .dinb(n9611), .dout(n9613));
  jand g09421(.dina(\a[41] ), .dinb(\a[31] ), .dout(n9614));
  jand g09422(.dina(\a[42] ), .dinb(\a[30] ), .dout(n9615));
  jor  g09423(.dina(n9615), .dinb(n9614), .dout(n9616));
  jnot g09424(.din(n9616), .dout(n9617));
  jand g09425(.dina(\a[42] ), .dinb(\a[31] ), .dout(n9618));
  jand g09426(.dina(n9618), .dinb(n9573), .dout(n9619));
  jor  g09427(.dina(n9619), .dinb(n9617), .dout(n9620));
  jxor g09428(.dina(n9620), .dinb(n9584), .dout(n9621));
  jnot g09429(.din(n9621), .dout(n9622));
  jnot g09430(.din(n9486), .dout(n9623));
  jnot g09431(.din(n9488), .dout(n9624));
  jand g09432(.dina(n9624), .dinb(n9623), .dout(n9625));
  jnot g09433(.din(n9625), .dout(n9626));
  jand g09434(.dina(n9488), .dinb(n9486), .dout(n9627));
  jor  g09435(.dina(n9498), .dinb(n9627), .dout(n9628));
  jand g09436(.dina(n9628), .dinb(n9626), .dout(n9629));
  jxor g09437(.dina(n9629), .dinb(n9622), .dout(n9630));
  jxor g09438(.dina(n9630), .dinb(n9613), .dout(n9631));
  jxor g09439(.dina(n9631), .dinb(n9610), .dout(n9632));
  jand g09440(.dina(n9499), .dinb(n9484), .dout(n9633));
  jand g09441(.dina(n9531), .dinb(n9500), .dout(n9634));
  jor  g09442(.dina(n9634), .dinb(n9633), .dout(n9635));
  jxor g09443(.dina(n9635), .dinb(n9632), .dout(n9636));
  jand g09444(.dina(n9448), .dinb(n9431), .dout(n9637));
  jand g09445(.dina(n9476), .dinb(n9449), .dout(n9638));
  jor  g09446(.dina(n9638), .dinb(n9637), .dout(n9639));
  jxor g09447(.dina(n9639), .dinb(n9636), .dout(n9640));
  jxor g09448(.dina(n9640), .dinb(n9607), .dout(n9641));
  jand g09449(.dina(n9477), .dinb(n9428), .dout(n9642));
  jand g09450(.dina(n9593), .dinb(n9478), .dout(n9643));
  jor  g09451(.dina(n9643), .dinb(n9642), .dout(n9644));
  jxor g09452(.dina(n9644), .dinb(n9641), .dout(n9645));
  jand g09453(.dina(n9419), .dinb(n9416), .dout(n9646));
  jand g09454(.dina(n9420), .dinb(n9395), .dout(n9647));
  jor  g09455(.dina(n9647), .dinb(n9646), .dout(n9648));
  jand g09456(.dina(n9458), .dinb(n9456), .dout(n9649));
  jand g09457(.dina(n9461), .dinb(n9459), .dout(n9650));
  jor  g09458(.dina(n9650), .dinb(n9649), .dout(n9651));
  jnot g09459(.din(n9580), .dout(n9652));
  jor  g09460(.dina(n9588), .dinb(n9652), .dout(n9653));
  jnot g09461(.din(n9572), .dout(n9654));
  jand g09462(.dina(n9588), .dinb(n9652), .dout(n9655));
  jor  g09463(.dina(n9655), .dinb(n9654), .dout(n9656));
  jand g09464(.dina(n9656), .dinb(n9653), .dout(n9657));
  jxor g09465(.dina(n9657), .dinb(n9651), .dout(n9658));
  jnot g09466(.din(n9658), .dout(n9659));
  jor  g09467(.dina(n9523), .dinb(n9508), .dout(n9660));
  jor  g09468(.dina(n9530), .dinb(n9525), .dout(n9661));
  jand g09469(.dina(n9661), .dinb(n9660), .dout(n9662));
  jxor g09470(.dina(n9662), .dinb(n9659), .dout(n9663));
  jand g09471(.dina(n9590), .dinb(n9565), .dout(n9664));
  jand g09472(.dina(n9591), .dinb(n9536), .dout(n9665));
  jor  g09473(.dina(n9665), .dinb(n9664), .dout(n9666));
  jxor g09474(.dina(n9666), .dinb(n9663), .dout(n9667));
  jand g09475(.dina(n9563), .dinb(n9556), .dout(n9668));
  jand g09476(.dina(n9564), .dinb(n9546), .dout(n9669));
  jor  g09477(.dina(n9669), .dinb(n9668), .dout(n9670));
  jand g09478(.dina(n9587), .dinb(n9329), .dout(n9671));
  jor  g09479(.dina(n9671), .dinb(n9585), .dout(n9672));
  jand g09480(.dina(n9568), .dinb(n9566), .dout(n9673));
  jor  g09481(.dina(n9673), .dinb(n9570), .dout(n9674));
  jxor g09482(.dina(n9674), .dinb(n9672), .dout(n9675));
  jand g09483(.dina(n9575), .dinb(n9573), .dout(n9676));
  jor  g09484(.dina(n9676), .dinb(n9578), .dout(n9677));
  jxor g09485(.dina(n9677), .dinb(n9675), .dout(n9678));
  jnot g09486(.din(n9528), .dout(n9679));
  jand g09487(.dina(n9679), .dinb(n9527), .dout(n9680));
  jnot g09488(.din(n9680), .dout(n9681));
  jand g09489(.dina(n9528), .dinb(n9262), .dout(n9682));
  jor  g09490(.dina(n9682), .dinb(n9526), .dout(n9683));
  jand g09491(.dina(n9683), .dinb(n9681), .dout(n9684));
  jxor g09492(.dina(n9684), .dinb(n9519), .dout(n9685));
  jand g09493(.dina(n9503), .dinb(n9501), .dout(n9686));
  jor  g09494(.dina(n9686), .dinb(n9506), .dout(n9687));
  jxor g09495(.dina(n9687), .dinb(n9685), .dout(n9688));
  jxor g09496(.dina(n9688), .dinb(n9678), .dout(n9689));
  jxor g09497(.dina(n9689), .dinb(n9670), .dout(n9690));
  jxor g09498(.dina(n9690), .dinb(n9667), .dout(n9691));
  jxor g09499(.dina(n9691), .dinb(n9648), .dout(n9692));
  jand g09500(.dina(n9440), .dinb(n9434), .dout(n9693));
  jand g09501(.dina(n9447), .dinb(n9441), .dout(n9694));
  jor  g09502(.dina(n9694), .dinb(n9693), .dout(n9695));
  jand g09503(.dina(n9545), .dinb(n9543), .dout(n9696));
  jor  g09504(.dina(n9696), .dinb(n9541), .dout(n9697));
  jand g09505(.dina(\a[60] ), .dinb(\a[12] ), .dout(n9698));
  jand g09506(.dina(\a[48] ), .dinb(\a[24] ), .dout(n9699));
  jand g09507(.dina(\a[47] ), .dinb(\a[25] ), .dout(n9700));
  jor  g09508(.dina(n9700), .dinb(n9699), .dout(n9701));
  jnot g09509(.din(n9701), .dout(n9702));
  jand g09510(.dina(\a[48] ), .dinb(\a[25] ), .dout(n9703));
  jand g09511(.dina(n9703), .dinb(n9547), .dout(n9704));
  jor  g09512(.dina(n9704), .dinb(n9702), .dout(n9705));
  jxor g09513(.dina(n9705), .dinb(n9698), .dout(n9706));
  jnot g09514(.din(n9706), .dout(n9707));
  jxor g09515(.dina(n9707), .dinb(n9697), .dout(n9708));
  jand g09516(.dina(\a[63] ), .dinb(\a[9] ), .dout(n9709));
  jand g09517(.dina(\a[62] ), .dinb(\a[10] ), .dout(n9710));
  jand g09518(.dina(\a[61] ), .dinb(\a[11] ), .dout(n9711));
  jor  g09519(.dina(n9711), .dinb(n9710), .dout(n9712));
  jand g09520(.dina(\a[62] ), .dinb(\a[11] ), .dout(n9713));
  jand g09521(.dina(n9713), .dinb(n9491), .dout(n9714));
  jnot g09522(.din(n9714), .dout(n9715));
  jand g09523(.dina(n9715), .dinb(n9712), .dout(n9716));
  jxor g09524(.dina(n9716), .dinb(n9709), .dout(n9717));
  jxor g09525(.dina(n9717), .dinb(n9708), .dout(n9718));
  jand g09526(.dina(\a[55] ), .dinb(\a[17] ), .dout(n9719));
  jnot g09527(.din(n9719), .dout(n9720));
  jor  g09528(.dina(n9505), .dinb(n7507), .dout(n9721));
  jand g09529(.dina(\a[54] ), .dinb(\a[20] ), .dout(n9722));
  jand g09530(.dina(n9722), .dinb(n6854), .dout(n9723));
  jnot g09531(.din(n9723), .dout(n9724));
  jand g09532(.dina(n9724), .dinb(n9721), .dout(n9725));
  jxor g09533(.dina(n9725), .dinb(n9720), .dout(n9726));
  jand g09534(.dina(\a[37] ), .dinb(\a[35] ), .dout(n9727));
  jnot g09535(.din(n9727), .dout(n9728));
  jand g09536(.dina(\a[51] ), .dinb(\a[21] ), .dout(n9729));
  jand g09537(.dina(\a[50] ), .dinb(\a[22] ), .dout(n9730));
  jor  g09538(.dina(n9730), .dinb(n9729), .dout(n9731));
  jand g09539(.dina(\a[51] ), .dinb(\a[22] ), .dout(n9732));
  jand g09540(.dina(n9732), .dinb(n9501), .dout(n9733));
  jnot g09541(.din(n9733), .dout(n9734));
  jand g09542(.dina(n9734), .dinb(n9731), .dout(n9735));
  jxor g09543(.dina(n9735), .dinb(n9728), .dout(n9736));
  jnot g09544(.din(n9577), .dout(n9737));
  jand g09545(.dina(\a[49] ), .dinb(\a[23] ), .dout(n9738));
  jxor g09546(.dina(n9738), .dinb(n7946), .dout(n9739));
  jxor g09547(.dina(n9739), .dinb(n9737), .dout(n9740));
  jnot g09548(.din(n9740), .dout(n9741));
  jxor g09549(.dina(n9741), .dinb(n9736), .dout(n9742));
  jxor g09550(.dina(n9742), .dinb(n9726), .dout(n9743));
  jxor g09551(.dina(n9743), .dinb(n9718), .dout(n9744));
  jxor g09552(.dina(n9744), .dinb(n9695), .dout(n9745));
  jand g09553(.dina(n9411), .dinb(n9408), .dout(n9746));
  jand g09554(.dina(n9415), .dinb(n9412), .dout(n9747));
  jor  g09555(.dina(n9747), .dinb(n9746), .dout(n9748));
  jand g09556(.dina(n9562), .dinb(n9557), .dout(n9749));
  jor  g09557(.dina(n9749), .dinb(n9560), .dout(n9750));
  jand g09558(.dina(n9550), .dinb(n9547), .dout(n9751));
  jor  g09559(.dina(n9751), .dinb(n9553), .dout(n9752));
  jxor g09560(.dina(n9752), .dinb(n9750), .dout(n9753));
  jand g09561(.dina(n9492), .dinb(n9286), .dout(n9754));
  jor  g09562(.dina(n9754), .dinb(n9495), .dout(n9755));
  jxor g09563(.dina(n9755), .dinb(n9753), .dout(n9756));
  jand g09564(.dina(n9403), .dinb(n9398), .dout(n9757));
  jand g09565(.dina(n9407), .dinb(n9404), .dout(n9758));
  jor  g09566(.dina(n9758), .dinb(n9757), .dout(n9759));
  jxor g09567(.dina(n9759), .dinb(n9756), .dout(n9760));
  jand g09568(.dina(\a[53] ), .dinb(\a[19] ), .dout(n9761));
  jand g09569(.dina(\a[38] ), .dinb(\a[34] ), .dout(n9762));
  jand g09570(.dina(\a[39] ), .dinb(\a[33] ), .dout(n9763));
  jor  g09571(.dina(n9763), .dinb(n9762), .dout(n9764));
  jnot g09572(.din(n9764), .dout(n9765));
  jand g09573(.dina(\a[39] ), .dinb(\a[34] ), .dout(n9766));
  jand g09574(.dina(n9766), .dinb(n9526), .dout(n9767));
  jor  g09575(.dina(n9767), .dinb(n9765), .dout(n9768));
  jxor g09576(.dina(n9768), .dinb(n9761), .dout(n9769));
  jand g09577(.dina(\a[45] ), .dinb(\a[27] ), .dout(n9770));
  jand g09578(.dina(\a[44] ), .dinb(\a[28] ), .dout(n9771));
  jor  g09579(.dina(n9771), .dinb(n9770), .dout(n9772));
  jnot g09580(.din(n9772), .dout(n9773));
  jand g09581(.dina(\a[45] ), .dinb(\a[28] ), .dout(n9774));
  jand g09582(.dina(n9774), .dinb(n9329), .dout(n9775));
  jor  g09583(.dina(n9775), .dinb(n9773), .dout(n9776));
  jxor g09584(.dina(n9776), .dinb(n9552), .dout(n9777));
  jand g09585(.dina(\a[58] ), .dinb(\a[14] ), .dout(n9778));
  jand g09586(.dina(\a[57] ), .dinb(\a[15] ), .dout(n9779));
  jor  g09587(.dina(n9779), .dinb(n9778), .dout(n9780));
  jand g09588(.dina(\a[58] ), .dinb(\a[15] ), .dout(n9781));
  jand g09589(.dina(n9781), .dinb(n9557), .dout(n9782));
  jnot g09590(.din(n9782), .dout(n9783));
  jand g09591(.dina(n9783), .dinb(n9780), .dout(n9784));
  jxor g09592(.dina(n9784), .dinb(n9540), .dout(n9785));
  jxor g09593(.dina(n9785), .dinb(n9777), .dout(n9786));
  jxor g09594(.dina(n9786), .dinb(n9769), .dout(n9787));
  jxor g09595(.dina(n9787), .dinb(n9760), .dout(n9788));
  jxor g09596(.dina(n9788), .dinb(n9748), .dout(n9789));
  jxor g09597(.dina(n9789), .dinb(n9745), .dout(n9790));
  jxor g09598(.dina(n9790), .dinb(n9692), .dout(n9791));
  jxor g09599(.dina(n9791), .dinb(n9645), .dout(n9792));
  jand g09600(.dina(n9424), .dinb(n9421), .dout(n9793));
  jand g09601(.dina(n9594), .dinb(n9425), .dout(n9794));
  jor  g09602(.dina(n9794), .dinb(n9793), .dout(n9795));
  jxor g09603(.dina(n9795), .dinb(n9792), .dout(n9796));
  jand g09604(.dina(n9595), .dinb(n9392), .dout(n9797));
  jnot g09605(.din(n9392), .dout(n9798));
  jnot g09606(.din(n9595), .dout(n9799));
  jand g09607(.dina(n9799), .dinb(n9798), .dout(n9800));
  jnot g09608(.din(n9800), .dout(n9801));
  jand g09609(.dina(n9603), .dinb(n9801), .dout(n9802));
  jor  g09610(.dina(n9802), .dinb(n9797), .dout(n9803));
  jxor g09611(.dina(n9803), .dinb(n9796), .dout(\asquared[73] ));
  jand g09612(.dina(n9644), .dinb(n9641), .dout(n9805));
  jand g09613(.dina(n9791), .dinb(n9645), .dout(n9806));
  jor  g09614(.dina(n9806), .dinb(n9805), .dout(n9807));
  jand g09615(.dina(n9691), .dinb(n9648), .dout(n9808));
  jand g09616(.dina(n9790), .dinb(n9692), .dout(n9809));
  jor  g09617(.dina(n9809), .dinb(n9808), .dout(n9810));
  jand g09618(.dina(n9788), .dinb(n9748), .dout(n9811));
  jand g09619(.dina(n9789), .dinb(n9745), .dout(n9812));
  jor  g09620(.dina(n9812), .dinb(n9811), .dout(n9813));
  jand g09621(.dina(n9666), .dinb(n9663), .dout(n9814));
  jand g09622(.dina(n9690), .dinb(n9667), .dout(n9815));
  jor  g09623(.dina(n9815), .dinb(n9814), .dout(n9816));
  jand g09624(.dina(n9759), .dinb(n9756), .dout(n9817));
  jand g09625(.dina(n9787), .dinb(n9760), .dout(n9818));
  jor  g09626(.dina(n9818), .dinb(n9817), .dout(n9819));
  jand g09627(.dina(n9674), .dinb(n9672), .dout(n9820));
  jand g09628(.dina(n9677), .dinb(n9675), .dout(n9821));
  jor  g09629(.dina(n9821), .dinb(n9820), .dout(n9822));
  jand g09630(.dina(n9752), .dinb(n9750), .dout(n9823));
  jand g09631(.dina(n9755), .dinb(n9753), .dout(n9824));
  jor  g09632(.dina(n9824), .dinb(n9823), .dout(n9825));
  jnot g09633(.din(n9825), .dout(n9826));
  jand g09634(.dina(\a[41] ), .dinb(\a[32] ), .dout(n9827));
  jand g09635(.dina(\a[40] ), .dinb(\a[33] ), .dout(n9828));
  jor  g09636(.dina(n9828), .dinb(n9827), .dout(n9829));
  jnot g09637(.din(n9829), .dout(n9830));
  jand g09638(.dina(\a[41] ), .dinb(\a[33] ), .dout(n9831));
  jand g09639(.dina(n9831), .dinb(n9577), .dout(n9832));
  jor  g09640(.dina(n9832), .dinb(n9830), .dout(n9833));
  jxor g09641(.dina(n9833), .dinb(n9618), .dout(n9834));
  jxor g09642(.dina(n9834), .dinb(n9826), .dout(n9835));
  jxor g09643(.dina(n9835), .dinb(n9822), .dout(n9836));
  jand g09644(.dina(n9688), .dinb(n9678), .dout(n9837));
  jand g09645(.dina(n9689), .dinb(n9670), .dout(n9838));
  jor  g09646(.dina(n9838), .dinb(n9837), .dout(n9839));
  jxor g09647(.dina(n9839), .dinb(n9836), .dout(n9840));
  jxor g09648(.dina(n9840), .dinb(n9819), .dout(n9841));
  jxor g09649(.dina(n9841), .dinb(n9816), .dout(n9842));
  jxor g09650(.dina(n9842), .dinb(n9813), .dout(n9843));
  jxor g09651(.dina(n9843), .dinb(n9810), .dout(n9844));
  jand g09652(.dina(n9639), .dinb(n9636), .dout(n9845));
  jand g09653(.dina(n9640), .dinb(n9607), .dout(n9846));
  jor  g09654(.dina(n9846), .dinb(n9845), .dout(n9847));
  jand g09655(.dina(n9707), .dinb(n9697), .dout(n9848));
  jand g09656(.dina(n9717), .dinb(n9708), .dout(n9849));
  jor  g09657(.dina(n9849), .dinb(n9848), .dout(n9850));
  jand g09658(.dina(n9684), .dinb(n9519), .dout(n9851));
  jand g09659(.dina(n9687), .dinb(n9685), .dout(n9852));
  jor  g09660(.dina(n9852), .dinb(n9851), .dout(n9853));
  jxor g09661(.dina(n9853), .dinb(n9850), .dout(n9854));
  jnot g09662(.din(n9777), .dout(n9855));
  jor  g09663(.dina(n9785), .dinb(n9855), .dout(n9856));
  jnot g09664(.din(n9769), .dout(n9857));
  jand g09665(.dina(n9785), .dinb(n9855), .dout(n9858));
  jor  g09666(.dina(n9858), .dinb(n9857), .dout(n9859));
  jand g09667(.dina(n9859), .dinb(n9856), .dout(n9860));
  jxor g09668(.dina(n9860), .dinb(n9854), .dout(n9861));
  jand g09669(.dina(n9743), .dinb(n9718), .dout(n9862));
  jand g09670(.dina(n9744), .dinb(n9695), .dout(n9863));
  jor  g09671(.dina(n9863), .dinb(n9862), .dout(n9864));
  jxor g09672(.dina(n9864), .dinb(n9861), .dout(n9865));
  jand g09673(.dina(\a[60] ), .dinb(\a[13] ), .dout(n9866));
  jand g09674(.dina(n9731), .dinb(n9727), .dout(n9867));
  jor  g09675(.dina(n9867), .dinb(n9733), .dout(n9868));
  jxor g09676(.dina(n9868), .dinb(n9866), .dout(n9869));
  jand g09677(.dina(n9764), .dinb(n9761), .dout(n9870));
  jor  g09678(.dina(n9870), .dinb(n9767), .dout(n9871));
  jxor g09679(.dina(n9871), .dinb(n9869), .dout(n9872));
  jand g09680(.dina(n9716), .dinb(n9709), .dout(n9873));
  jor  g09681(.dina(n9873), .dinb(n9714), .dout(n9874));
  jand g09682(.dina(n9701), .dinb(n9698), .dout(n9875));
  jor  g09683(.dina(n9875), .dinb(n9704), .dout(n9876));
  jxor g09684(.dina(n9876), .dinb(n9874), .dout(n9877));
  jand g09685(.dina(n9721), .dinb(n9719), .dout(n9878));
  jor  g09686(.dina(n9878), .dinb(n9723), .dout(n9879));
  jxor g09687(.dina(n9879), .dinb(n9877), .dout(n9880));
  jxor g09688(.dina(n9880), .dinb(n9872), .dout(n9881));
  jnot g09689(.din(n9881), .dout(n9882));
  jnot g09690(.din(n9736), .dout(n9883));
  jand g09691(.dina(n9741), .dinb(n9883), .dout(n9884));
  jnot g09692(.din(n9884), .dout(n9885));
  jand g09693(.dina(n9740), .dinb(n9736), .dout(n9886));
  jor  g09694(.dina(n9886), .dinb(n9726), .dout(n9887));
  jand g09695(.dina(n9887), .dinb(n9885), .dout(n9888));
  jxor g09696(.dina(n9888), .dinb(n9882), .dout(n9889));
  jxor g09697(.dina(n9889), .dinb(n9865), .dout(n9890));
  jxor g09698(.dina(n9890), .dinb(n9847), .dout(n9891));
  jand g09699(.dina(n9657), .dinb(n9651), .dout(n9892));
  jnot g09700(.din(n9892), .dout(n9893));
  jor  g09701(.dina(n9662), .dinb(n9659), .dout(n9894));
  jand g09702(.dina(n9894), .dinb(n9893), .dout(n9895));
  jnot g09703(.din(n9895), .dout(n9896));
  jnot g09704(.din(n9732), .dout(n9897));
  jand g09705(.dina(\a[53] ), .dinb(\a[20] ), .dout(n9898));
  jand g09706(.dina(\a[52] ), .dinb(\a[21] ), .dout(n9899));
  jor  g09707(.dina(n9899), .dinb(n9898), .dout(n9900));
  jand g09708(.dina(\a[53] ), .dinb(\a[21] ), .dout(n9901));
  jand g09709(.dina(n9901), .dinb(n9505), .dout(n9902));
  jnot g09710(.din(n9902), .dout(n9903));
  jand g09711(.dina(n9903), .dinb(n9900), .dout(n9904));
  jxor g09712(.dina(n9904), .dinb(n9897), .dout(n9905));
  jand g09713(.dina(\a[55] ), .dinb(\a[18] ), .dout(n9906));
  jnot g09714(.din(n9906), .dout(n9907));
  jand g09715(.dina(\a[54] ), .dinb(\a[19] ), .dout(n9908));
  jand g09716(.dina(\a[49] ), .dinb(\a[24] ), .dout(n9909));
  jor  g09717(.dina(n9909), .dinb(n9908), .dout(n9910));
  jand g09718(.dina(\a[54] ), .dinb(\a[24] ), .dout(n9911));
  jand g09719(.dina(n9911), .dinb(n8799), .dout(n9912));
  jnot g09720(.din(n9912), .dout(n9913));
  jand g09721(.dina(n9913), .dinb(n9910), .dout(n9914));
  jxor g09722(.dina(n9914), .dinb(n9907), .dout(n9915));
  jnot g09723(.din(n9915), .dout(n9916));
  jand g09724(.dina(\a[50] ), .dinb(\a[23] ), .dout(n9917));
  jnot g09725(.din(n9917), .dout(n9918));
  jor  g09726(.dina(n9713), .dinb(\a[37] ), .dout(n9919));
  jand g09727(.dina(n3822), .dinb(\a[62] ), .dout(n9920));
  jnot g09728(.din(n9920), .dout(n9921));
  jand g09729(.dina(n9921), .dinb(n9919), .dout(n9922));
  jor  g09730(.dina(n9922), .dinb(n9918), .dout(n9923));
  jand g09731(.dina(n9919), .dinb(n9917), .dout(n9924));
  jor  g09732(.dina(n9924), .dinb(n9920), .dout(n9925));
  jnot g09733(.din(n9925), .dout(n9926));
  jand g09734(.dina(n9926), .dinb(n9919), .dout(n9927));
  jnot g09735(.din(n9927), .dout(n9928));
  jand g09736(.dina(n9928), .dinb(n9923), .dout(n9929));
  jxor g09737(.dina(n9929), .dinb(n9916), .dout(n9930));
  jxor g09738(.dina(n9930), .dinb(n9905), .dout(n9931));
  jand g09739(.dina(\a[56] ), .dinb(\a[17] ), .dout(n9932));
  jand g09740(.dina(\a[47] ), .dinb(\a[26] ), .dout(n9933));
  jand g09741(.dina(\a[46] ), .dinb(\a[27] ), .dout(n9934));
  jor  g09742(.dina(n9934), .dinb(n9933), .dout(n9935));
  jnot g09743(.din(n9935), .dout(n9936));
  jand g09744(.dina(\a[47] ), .dinb(\a[27] ), .dout(n9937));
  jand g09745(.dina(n9937), .dinb(n9552), .dout(n9938));
  jor  g09746(.dina(n9938), .dinb(n9936), .dout(n9939));
  jxor g09747(.dina(n9939), .dinb(n9932), .dout(n9940));
  jnot g09748(.din(n9940), .dout(n9941));
  jnot g09749(.din(n7946), .dout(n9942));
  jnot g09750(.din(n9738), .dout(n9943));
  jand g09751(.dina(n9943), .dinb(n9942), .dout(n9944));
  jnot g09752(.din(n9944), .dout(n9945));
  jand g09753(.dina(n9738), .dinb(n7946), .dout(n9946));
  jor  g09754(.dina(n9946), .dinb(n9577), .dout(n9947));
  jand g09755(.dina(n9947), .dinb(n9945), .dout(n9948));
  jxor g09756(.dina(n9948), .dinb(n9941), .dout(n9949));
  jand g09757(.dina(\a[59] ), .dinb(\a[14] ), .dout(n9950));
  jand g09758(.dina(\a[57] ), .dinb(\a[16] ), .dout(n9951));
  jor  g09759(.dina(n9951), .dinb(n9781), .dout(n9952));
  jand g09760(.dina(\a[58] ), .dinb(\a[16] ), .dout(n9953));
  jand g09761(.dina(n9953), .dinb(n9779), .dout(n9954));
  jnot g09762(.din(n9954), .dout(n9955));
  jand g09763(.dina(n9955), .dinb(n9952), .dout(n9956));
  jxor g09764(.dina(n9956), .dinb(n9950), .dout(n9957));
  jxor g09765(.dina(n9957), .dinb(n9949), .dout(n9958));
  jxor g09766(.dina(n9958), .dinb(n9931), .dout(n9959));
  jxor g09767(.dina(n9959), .dinb(n9896), .dout(n9960));
  jand g09768(.dina(n9631), .dinb(n9610), .dout(n9961));
  jand g09769(.dina(n9635), .dinb(n9632), .dout(n9962));
  jor  g09770(.dina(n9962), .dinb(n9961), .dout(n9963));
  jand g09771(.dina(n9784), .dinb(n9540), .dout(n9964));
  jor  g09772(.dina(n9964), .dinb(n9782), .dout(n9965));
  jand g09773(.dina(n9772), .dinb(n9552), .dout(n9966));
  jor  g09774(.dina(n9966), .dinb(n9775), .dout(n9967));
  jxor g09775(.dina(n9967), .dinb(n9965), .dout(n9968));
  jand g09776(.dina(n9616), .dinb(n9584), .dout(n9969));
  jor  g09777(.dina(n9969), .dinb(n9619), .dout(n9970));
  jxor g09778(.dina(n9970), .dinb(n9968), .dout(n9971));
  jand g09779(.dina(n9629), .dinb(n9622), .dout(n9972));
  jand g09780(.dina(n9630), .dinb(n9613), .dout(n9973));
  jor  g09781(.dina(n9973), .dinb(n9972), .dout(n9974));
  jxor g09782(.dina(n9974), .dinb(n9971), .dout(n9975));
  jand g09783(.dina(\a[44] ), .dinb(\a[29] ), .dout(n9976));
  jand g09784(.dina(\a[43] ), .dinb(\a[30] ), .dout(n9977));
  jor  g09785(.dina(n9977), .dinb(n9976), .dout(n9978));
  jnot g09786(.din(n9978), .dout(n9979));
  jand g09787(.dina(\a[44] ), .dinb(\a[30] ), .dout(n9980));
  jand g09788(.dina(n9980), .dinb(n9584), .dout(n9981));
  jor  g09789(.dina(n9981), .dinb(n9979), .dout(n9982));
  jxor g09790(.dina(n9982), .dinb(n9774), .dout(n9983));
  jnot g09791(.din(n9983), .dout(n9984));
  jand g09792(.dina(\a[61] ), .dinb(\a[12] ), .dout(n9985));
  jor  g09793(.dina(n9985), .dinb(n9494), .dout(n9986));
  jand g09794(.dina(\a[63] ), .dinb(\a[12] ), .dout(n9987));
  jand g09795(.dina(n9987), .dinb(n9491), .dout(n9988));
  jnot g09796(.din(n9988), .dout(n9989));
  jand g09797(.dina(n9989), .dinb(n9986), .dout(n9990));
  jxor g09798(.dina(n9990), .dinb(n9703), .dout(n9991));
  jxor g09799(.dina(n9991), .dinb(n9984), .dout(n9992));
  jnot g09800(.din(n9992), .dout(n9993));
  jand g09801(.dina(\a[38] ), .dinb(\a[35] ), .dout(n9994));
  jand g09802(.dina(\a[37] ), .dinb(\a[36] ), .dout(n9995));
  jor  g09803(.dina(n9995), .dinb(n9994), .dout(n9996));
  jnot g09804(.din(n9996), .dout(n9997));
  jand g09805(.dina(\a[38] ), .dinb(\a[36] ), .dout(n9998));
  jand g09806(.dina(n9998), .dinb(n9727), .dout(n9999));
  jor  g09807(.dina(n9999), .dinb(n9997), .dout(n10000));
  jxor g09808(.dina(n10000), .dinb(n9766), .dout(n10001));
  jxor g09809(.dina(n10001), .dinb(n9993), .dout(n10002));
  jxor g09810(.dina(n10002), .dinb(n9975), .dout(n10003));
  jxor g09811(.dina(n10003), .dinb(n9963), .dout(n10004));
  jxor g09812(.dina(n10004), .dinb(n9960), .dout(n10005));
  jxor g09813(.dina(n10005), .dinb(n9891), .dout(n10006));
  jxor g09814(.dina(n10006), .dinb(n9844), .dout(n10007));
  jxor g09815(.dina(n10007), .dinb(n9807), .dout(n10008));
  jand g09816(.dina(n9795), .dinb(n9792), .dout(n10009));
  jnot g09817(.din(n9792), .dout(n10010));
  jnot g09818(.din(n9795), .dout(n10011));
  jand g09819(.dina(n10011), .dinb(n10010), .dout(n10012));
  jnot g09820(.din(n10012), .dout(n10013));
  jand g09821(.dina(n9803), .dinb(n10013), .dout(n10014));
  jor  g09822(.dina(n10014), .dinb(n10009), .dout(n10015));
  jxor g09823(.dina(n10015), .dinb(n10008), .dout(\asquared[74] ));
  jand g09824(.dina(n9843), .dinb(n9810), .dout(n10017));
  jand g09825(.dina(n10006), .dinb(n9844), .dout(n10018));
  jor  g09826(.dina(n10018), .dinb(n10017), .dout(n10019));
  jand g09827(.dina(n9890), .dinb(n9847), .dout(n10020));
  jand g09828(.dina(n10005), .dinb(n9891), .dout(n10021));
  jor  g09829(.dina(n10021), .dinb(n10020), .dout(n10022));
  jand g09830(.dina(n10003), .dinb(n9963), .dout(n10023));
  jand g09831(.dina(n10004), .dinb(n9960), .dout(n10024));
  jor  g09832(.dina(n10024), .dinb(n10023), .dout(n10025));
  jand g09833(.dina(n9864), .dinb(n9861), .dout(n10026));
  jand g09834(.dina(n9889), .dinb(n9865), .dout(n10027));
  jor  g09835(.dina(n10027), .dinb(n10026), .dout(n10028));
  jand g09836(.dina(n9876), .dinb(n9874), .dout(n10029));
  jand g09837(.dina(n9879), .dinb(n9877), .dout(n10030));
  jor  g09838(.dina(n10030), .dinb(n10029), .dout(n10031));
  jand g09839(.dina(n9868), .dinb(n9866), .dout(n10032));
  jand g09840(.dina(n9871), .dinb(n9869), .dout(n10033));
  jor  g09841(.dina(n10033), .dinb(n10032), .dout(n10034));
  jxor g09842(.dina(n10034), .dinb(n10031), .dout(n10035));
  jor  g09843(.dina(n9948), .dinb(n9941), .dout(n10036));
  jand g09844(.dina(n9948), .dinb(n9941), .dout(n10037));
  jor  g09845(.dina(n9957), .dinb(n10037), .dout(n10038));
  jand g09846(.dina(n10038), .dinb(n10036), .dout(n10039));
  jxor g09847(.dina(n10039), .dinb(n10035), .dout(n10040));
  jand g09848(.dina(n9880), .dinb(n9872), .dout(n10041));
  jnot g09849(.din(n10041), .dout(n10042));
  jor  g09850(.dina(n9888), .dinb(n9882), .dout(n10043));
  jand g09851(.dina(n10043), .dinb(n10042), .dout(n10044));
  jnot g09852(.din(n10044), .dout(n10045));
  jand g09853(.dina(n9853), .dinb(n9850), .dout(n10046));
  jand g09854(.dina(n9860), .dinb(n9854), .dout(n10047));
  jor  g09855(.dina(n10047), .dinb(n10046), .dout(n10048));
  jxor g09856(.dina(n10048), .dinb(n10045), .dout(n10049));
  jxor g09857(.dina(n10049), .dinb(n10040), .dout(n10050));
  jxor g09858(.dina(n10050), .dinb(n10028), .dout(n10051));
  jxor g09859(.dina(n10051), .dinb(n10025), .dout(n10052));
  jxor g09860(.dina(n10052), .dinb(n10022), .dout(n10053));
  jand g09861(.dina(n9841), .dinb(n9816), .dout(n10054));
  jand g09862(.dina(n9842), .dinb(n9813), .dout(n10055));
  jor  g09863(.dina(n10055), .dinb(n10054), .dout(n10056));
  jnot g09864(.din(n9929), .dout(n10057));
  jand g09865(.dina(n10057), .dinb(n9916), .dout(n10058));
  jnot g09866(.din(n10058), .dout(n10059));
  jand g09867(.dina(n9929), .dinb(n9915), .dout(n10060));
  jor  g09868(.dina(n10060), .dinb(n9905), .dout(n10061));
  jand g09869(.dina(n10061), .dinb(n10059), .dout(n10062));
  jand g09870(.dina(n9829), .dinb(n9618), .dout(n10063));
  jor  g09871(.dina(n10063), .dinb(n9832), .dout(n10064));
  jand g09872(.dina(n9996), .dinb(n9766), .dout(n10065));
  jor  g09873(.dina(n10065), .dinb(n9999), .dout(n10066));
  jxor g09874(.dina(n10066), .dinb(n10064), .dout(n10067));
  jand g09875(.dina(\a[60] ), .dinb(\a[14] ), .dout(n10068));
  jand g09876(.dina(\a[59] ), .dinb(\a[15] ), .dout(n10069));
  jor  g09877(.dina(n10069), .dinb(n9953), .dout(n10070));
  jnot g09878(.din(n10070), .dout(n10071));
  jand g09879(.dina(\a[59] ), .dinb(\a[16] ), .dout(n10072));
  jand g09880(.dina(n10072), .dinb(n9781), .dout(n10073));
  jor  g09881(.dina(n10073), .dinb(n10071), .dout(n10074));
  jxor g09882(.dina(n10074), .dinb(n10068), .dout(n10075));
  jnot g09883(.din(n10075), .dout(n10076));
  jxor g09884(.dina(n10076), .dinb(n10067), .dout(n10077));
  jnot g09885(.din(n10077), .dout(n10078));
  jxor g09886(.dina(n10078), .dinb(n10062), .dout(n10079));
  jnot g09887(.din(n10079), .dout(n10080));
  jor  g09888(.dina(n9834), .dinb(n9826), .dout(n10081));
  jand g09889(.dina(n9835), .dinb(n9822), .dout(n10082));
  jnot g09890(.din(n10082), .dout(n10083));
  jand g09891(.dina(n10083), .dinb(n10081), .dout(n10084));
  jxor g09892(.dina(n10084), .dinb(n10080), .dout(n10085));
  jand g09893(.dina(n9958), .dinb(n9931), .dout(n10086));
  jand g09894(.dina(n9959), .dinb(n9896), .dout(n10087));
  jor  g09895(.dina(n10087), .dinb(n10086), .dout(n10088));
  jand g09896(.dina(n9974), .dinb(n9971), .dout(n10089));
  jand g09897(.dina(n10002), .dinb(n9975), .dout(n10090));
  jor  g09898(.dina(n10090), .dinb(n10089), .dout(n10091));
  jxor g09899(.dina(n10091), .dinb(n10088), .dout(n10092));
  jxor g09900(.dina(n10092), .dinb(n10085), .dout(n10093));
  jxor g09901(.dina(n10093), .dinb(n10056), .dout(n10094));
  jand g09902(.dina(n9839), .dinb(n9836), .dout(n10095));
  jand g09903(.dina(n9840), .dinb(n9819), .dout(n10096));
  jor  g09904(.dina(n10096), .dinb(n10095), .dout(n10097));
  jand g09905(.dina(n9956), .dinb(n9950), .dout(n10098));
  jor  g09906(.dina(n10098), .dinb(n9954), .dout(n10099));
  jand g09907(.dina(n9935), .dinb(n9932), .dout(n10100));
  jor  g09908(.dina(n10100), .dinb(n9938), .dout(n10101));
  jand g09909(.dina(n9978), .dinb(n9774), .dout(n10102));
  jor  g09910(.dina(n10102), .dinb(n9981), .dout(n10103));
  jxor g09911(.dina(n10103), .dinb(n10101), .dout(n10104));
  jxor g09912(.dina(n10104), .dinb(n10099), .dout(n10105));
  jand g09913(.dina(n9990), .dinb(n9703), .dout(n10106));
  jor  g09914(.dina(n10106), .dinb(n9988), .dout(n10107));
  jand g09915(.dina(n9910), .dinb(n9906), .dout(n10108));
  jor  g09916(.dina(n10108), .dinb(n9912), .dout(n10109));
  jand g09917(.dina(n9900), .dinb(n9732), .dout(n10110));
  jor  g09918(.dina(n10110), .dinb(n9902), .dout(n10111));
  jxor g09919(.dina(n10111), .dinb(n10109), .dout(n10112));
  jxor g09920(.dina(n10112), .dinb(n10107), .dout(n10113));
  jnot g09921(.din(n10113), .dout(n10114));
  jand g09922(.dina(n9991), .dinb(n9984), .dout(n10115));
  jnot g09923(.din(n10115), .dout(n10116));
  jor  g09924(.dina(n10001), .dinb(n9993), .dout(n10117));
  jand g09925(.dina(n10117), .dinb(n10116), .dout(n10118));
  jxor g09926(.dina(n10118), .dinb(n10114), .dout(n10119));
  jxor g09927(.dina(n10119), .dinb(n10105), .dout(n10120));
  jxor g09928(.dina(n10120), .dinb(n10097), .dout(n10121));
  jand g09929(.dina(n9967), .dinb(n9965), .dout(n10122));
  jand g09930(.dina(n9970), .dinb(n9968), .dout(n10123));
  jor  g09931(.dina(n10123), .dinb(n10122), .dout(n10124));
  jand g09932(.dina(\a[61] ), .dinb(\a[13] ), .dout(n10125));
  jand g09933(.dina(\a[62] ), .dinb(\a[12] ), .dout(n10126));
  jor  g09934(.dina(n10126), .dinb(n10125), .dout(n10127));
  jand g09935(.dina(\a[62] ), .dinb(\a[13] ), .dout(n10128));
  jand g09936(.dina(n10128), .dinb(n9985), .dout(n10129));
  jnot g09937(.din(n10129), .dout(n10130));
  jand g09938(.dina(n10130), .dinb(n10127), .dout(n10131));
  jxor g09939(.dina(n10131), .dinb(n9925), .dout(n10132));
  jnot g09940(.din(n10132), .dout(n10133));
  jand g09941(.dina(\a[45] ), .dinb(\a[29] ), .dout(n10134));
  jnot g09942(.din(n7975), .dout(n10135));
  jxor g09943(.dina(n9980), .dinb(n10135), .dout(n10136));
  jxor g09944(.dina(n10136), .dinb(n10134), .dout(n10137));
  jxor g09945(.dina(n10137), .dinb(n10133), .dout(n10138));
  jxor g09946(.dina(n10138), .dinb(n10124), .dout(n10139));
  jand g09947(.dina(\a[48] ), .dinb(\a[26] ), .dout(n10140));
  jand g09948(.dina(\a[46] ), .dinb(\a[28] ), .dout(n10141));
  jor  g09949(.dina(n10141), .dinb(n9937), .dout(n10142));
  jnot g09950(.din(n10142), .dout(n10143));
  jand g09951(.dina(\a[47] ), .dinb(\a[28] ), .dout(n10144));
  jand g09952(.dina(n10144), .dinb(n9934), .dout(n10145));
  jor  g09953(.dina(n10145), .dinb(n10143), .dout(n10146));
  jxor g09954(.dina(n10146), .dinb(n10140), .dout(n10147));
  jand g09955(.dina(\a[56] ), .dinb(\a[18] ), .dout(n10148));
  jand g09956(.dina(\a[49] ), .dinb(\a[25] ), .dout(n10149));
  jor  g09957(.dina(n10149), .dinb(n10148), .dout(n10150));
  jnot g09958(.din(n10150), .dout(n10151));
  jand g09959(.dina(\a[56] ), .dinb(\a[25] ), .dout(n10152));
  jand g09960(.dina(n10152), .dinb(n8650), .dout(n10153));
  jor  g09961(.dina(n10153), .dinb(n10151), .dout(n10154));
  jxor g09962(.dina(n10154), .dinb(n9831), .dout(n10155));
  jand g09963(.dina(\a[63] ), .dinb(\a[11] ), .dout(n10156));
  jand g09964(.dina(\a[43] ), .dinb(\a[31] ), .dout(n10157));
  jand g09965(.dina(\a[42] ), .dinb(\a[32] ), .dout(n10158));
  jor  g09966(.dina(n10158), .dinb(n10157), .dout(n10159));
  jand g09967(.dina(\a[43] ), .dinb(\a[32] ), .dout(n10160));
  jand g09968(.dina(n10160), .dinb(n9618), .dout(n10161));
  jnot g09969(.din(n10161), .dout(n10162));
  jand g09970(.dina(n10162), .dinb(n10159), .dout(n10163));
  jxor g09971(.dina(n10163), .dinb(n10156), .dout(n10164));
  jxor g09972(.dina(n10164), .dinb(n10155), .dout(n10165));
  jxor g09973(.dina(n10165), .dinb(n10147), .dout(n10166));
  jand g09974(.dina(\a[51] ), .dinb(\a[23] ), .dout(n10167));
  jand g09975(.dina(\a[50] ), .dinb(\a[24] ), .dout(n10168));
  jor  g09976(.dina(n10168), .dinb(n10167), .dout(n10169));
  jnot g09977(.din(n10169), .dout(n10170));
  jand g09978(.dina(\a[51] ), .dinb(\a[24] ), .dout(n10171));
  jand g09979(.dina(n10171), .dinb(n9917), .dout(n10172));
  jor  g09980(.dina(n10172), .dinb(n10170), .dout(n10173));
  jxor g09981(.dina(n10173), .dinb(n9998), .dout(n10174));
  jand g09982(.dina(\a[40] ), .dinb(\a[34] ), .dout(n10175));
  jand g09983(.dina(\a[39] ), .dinb(\a[35] ), .dout(n10176));
  jor  g09984(.dina(n10176), .dinb(n10175), .dout(n10177));
  jnot g09985(.din(n10177), .dout(n10178));
  jand g09986(.dina(\a[40] ), .dinb(\a[35] ), .dout(n10179));
  jand g09987(.dina(n10179), .dinb(n9766), .dout(n10180));
  jor  g09988(.dina(n10180), .dinb(n10178), .dout(n10181));
  jxor g09989(.dina(n10181), .dinb(n9722), .dout(n10182));
  jand g09990(.dina(\a[52] ), .dinb(\a[22] ), .dout(n10183));
  jor  g09991(.dina(n9901), .dinb(n7771), .dout(n10184));
  jand g09992(.dina(\a[55] ), .dinb(\a[21] ), .dout(n10185));
  jand g09993(.dina(n10185), .dinb(n9761), .dout(n10186));
  jnot g09994(.din(n10186), .dout(n10187));
  jand g09995(.dina(n10187), .dinb(n10184), .dout(n10188));
  jxor g09996(.dina(n10188), .dinb(n10183), .dout(n10189));
  jxor g09997(.dina(n10189), .dinb(n10182), .dout(n10190));
  jxor g09998(.dina(n10190), .dinb(n10174), .dout(n10191));
  jxor g09999(.dina(n10191), .dinb(n10166), .dout(n10192));
  jxor g10000(.dina(n10192), .dinb(n10139), .dout(n10193));
  jxor g10001(.dina(n10193), .dinb(n10121), .dout(n10194));
  jxor g10002(.dina(n10194), .dinb(n10094), .dout(n10195));
  jxor g10003(.dina(n10195), .dinb(n10053), .dout(n10196));
  jxor g10004(.dina(n10196), .dinb(n10019), .dout(n10197));
  jand g10005(.dina(n10007), .dinb(n9807), .dout(n10198));
  jnot g10006(.din(n9807), .dout(n10199));
  jnot g10007(.din(n10007), .dout(n10200));
  jand g10008(.dina(n10200), .dinb(n10199), .dout(n10201));
  jnot g10009(.din(n10201), .dout(n10202));
  jand g10010(.dina(n10015), .dinb(n10202), .dout(n10203));
  jor  g10011(.dina(n10203), .dinb(n10198), .dout(n10204));
  jxor g10012(.dina(n10204), .dinb(n10197), .dout(\asquared[75] ));
  jand g10013(.dina(n10052), .dinb(n10022), .dout(n10206));
  jand g10014(.dina(n10195), .dinb(n10053), .dout(n10207));
  jor  g10015(.dina(n10207), .dinb(n10206), .dout(n10208));
  jand g10016(.dina(n10050), .dinb(n10028), .dout(n10209));
  jand g10017(.dina(n10051), .dinb(n10025), .dout(n10210));
  jor  g10018(.dina(n10210), .dinb(n10209), .dout(n10211));
  jand g10019(.dina(n10111), .dinb(n10109), .dout(n10212));
  jand g10020(.dina(n10112), .dinb(n10107), .dout(n10213));
  jor  g10021(.dina(n10213), .dinb(n10212), .dout(n10214));
  jnot g10022(.din(n10064), .dout(n10215));
  jnot g10023(.din(n10066), .dout(n10216));
  jand g10024(.dina(n10216), .dinb(n10215), .dout(n10217));
  jnot g10025(.din(n10217), .dout(n10218));
  jand g10026(.dina(n10066), .dinb(n10064), .dout(n10219));
  jor  g10027(.dina(n10076), .dinb(n10219), .dout(n10220));
  jand g10028(.dina(n10220), .dinb(n10218), .dout(n10221));
  jxor g10029(.dina(n10221), .dinb(n10214), .dout(n10222));
  jand g10030(.dina(n10103), .dinb(n10101), .dout(n10223));
  jand g10031(.dina(n10104), .dinb(n10099), .dout(n10224));
  jor  g10032(.dina(n10224), .dinb(n10223), .dout(n10225));
  jxor g10033(.dina(n10225), .dinb(n10222), .dout(n10226));
  jand g10034(.dina(n10191), .dinb(n10166), .dout(n10227));
  jand g10035(.dina(n10192), .dinb(n10139), .dout(n10228));
  jor  g10036(.dina(n10228), .dinb(n10227), .dout(n10229));
  jxor g10037(.dina(n10229), .dinb(n10226), .dout(n10230));
  jor  g10038(.dina(n10137), .dinb(n10133), .dout(n10231));
  jand g10039(.dina(n10138), .dinb(n10124), .dout(n10232));
  jnot g10040(.din(n10232), .dout(n10233));
  jand g10041(.dina(n10233), .dinb(n10231), .dout(n10234));
  jnot g10042(.din(n10234), .dout(n10235));
  jand g10043(.dina(n10188), .dinb(n10183), .dout(n10236));
  jor  g10044(.dina(n10236), .dinb(n10186), .dout(n10237));
  jand g10045(.dina(n10177), .dinb(n9722), .dout(n10238));
  jor  g10046(.dina(n10238), .dinb(n10180), .dout(n10239));
  jand g10047(.dina(n10169), .dinb(n9998), .dout(n10240));
  jor  g10048(.dina(n10240), .dinb(n10172), .dout(n10241));
  jxor g10049(.dina(n10241), .dinb(n10239), .dout(n10242));
  jxor g10050(.dina(n10242), .dinb(n10237), .dout(n10243));
  jand g10051(.dina(n10163), .dinb(n10156), .dout(n10244));
  jor  g10052(.dina(n10244), .dinb(n10161), .dout(n10245));
  jand g10053(.dina(n10150), .dinb(n9831), .dout(n10246));
  jor  g10054(.dina(n10246), .dinb(n10153), .dout(n10247));
  jxor g10055(.dina(n10247), .dinb(n10245), .dout(n10248));
  jand g10056(.dina(n10131), .dinb(n9925), .dout(n10249));
  jor  g10057(.dina(n10249), .dinb(n10129), .dout(n10250));
  jxor g10058(.dina(n10250), .dinb(n10248), .dout(n10251));
  jxor g10059(.dina(n10251), .dinb(n10243), .dout(n10252));
  jxor g10060(.dina(n10252), .dinb(n10235), .dout(n10253));
  jxor g10061(.dina(n10253), .dinb(n10230), .dout(n10254));
  jxor g10062(.dina(n10254), .dinb(n10211), .dout(n10255));
  jand g10063(.dina(n10048), .dinb(n10045), .dout(n10256));
  jand g10064(.dina(n10049), .dinb(n10040), .dout(n10257));
  jor  g10065(.dina(n10257), .dinb(n10256), .dout(n10258));
  jand g10066(.dina(n10142), .dinb(n10140), .dout(n10259));
  jor  g10067(.dina(n10259), .dinb(n10145), .dout(n10260));
  jnot g10068(.din(n9980), .dout(n10261));
  jand g10069(.dina(n10261), .dinb(n10135), .dout(n10262));
  jnot g10070(.din(n10262), .dout(n10263));
  jand g10071(.dina(n9980), .dinb(n7975), .dout(n10264));
  jor  g10072(.dina(n10264), .dinb(n10134), .dout(n10265));
  jand g10073(.dina(n10265), .dinb(n10263), .dout(n10266));
  jxor g10074(.dina(n10266), .dinb(n10260), .dout(n10267));
  jand g10075(.dina(n10070), .dinb(n10068), .dout(n10268));
  jor  g10076(.dina(n10268), .dinb(n10073), .dout(n10269));
  jxor g10077(.dina(n10269), .dinb(n10267), .dout(n10270));
  jnot g10078(.din(n10182), .dout(n10271));
  jor  g10079(.dina(n10189), .dinb(n10271), .dout(n10272));
  jnot g10080(.din(n10174), .dout(n10273));
  jand g10081(.dina(n10189), .dinb(n10271), .dout(n10274));
  jor  g10082(.dina(n10274), .dinb(n10273), .dout(n10275));
  jand g10083(.dina(n10275), .dinb(n10272), .dout(n10276));
  jnot g10084(.din(n10155), .dout(n10277));
  jor  g10085(.dina(n10164), .dinb(n10277), .dout(n10278));
  jnot g10086(.din(n10147), .dout(n10279));
  jand g10087(.dina(n10164), .dinb(n10277), .dout(n10280));
  jor  g10088(.dina(n10280), .dinb(n10279), .dout(n10281));
  jand g10089(.dina(n10281), .dinb(n10278), .dout(n10282));
  jxor g10090(.dina(n10282), .dinb(n10276), .dout(n10283));
  jxor g10091(.dina(n10283), .dinb(n10270), .dout(n10284));
  jxor g10092(.dina(n10284), .dinb(n10258), .dout(n10285));
  jand g10093(.dina(n10034), .dinb(n10031), .dout(n10286));
  jand g10094(.dina(n10039), .dinb(n10035), .dout(n10287));
  jor  g10095(.dina(n10287), .dinb(n10286), .dout(n10288));
  jand g10096(.dina(\a[52] ), .dinb(\a[23] ), .dout(n10289));
  jand g10097(.dina(\a[39] ), .dinb(\a[36] ), .dout(n10290));
  jor  g10098(.dina(n10290), .dinb(n10179), .dout(n10291));
  jnot g10099(.din(n10291), .dout(n10292));
  jand g10100(.dina(\a[40] ), .dinb(\a[36] ), .dout(n10293));
  jand g10101(.dina(n10293), .dinb(n10176), .dout(n10294));
  jor  g10102(.dina(n10294), .dinb(n10292), .dout(n10295));
  jxor g10103(.dina(n10295), .dinb(n10289), .dout(n10296));
  jnot g10104(.din(n10296), .dout(n10297));
  jand g10105(.dina(\a[45] ), .dinb(\a[30] ), .dout(n10298));
  jand g10106(.dina(\a[56] ), .dinb(\a[19] ), .dout(n10299));
  jor  g10107(.dina(n10299), .dinb(n9987), .dout(n10300));
  jand g10108(.dina(\a[63] ), .dinb(\a[19] ), .dout(n10301));
  jand g10109(.dina(n10301), .dinb(n8808), .dout(n10302));
  jnot g10110(.din(n10302), .dout(n10303));
  jand g10111(.dina(n10303), .dinb(n10300), .dout(n10304));
  jxor g10112(.dina(n10304), .dinb(n10298), .dout(n10305));
  jxor g10113(.dina(n10305), .dinb(n10297), .dout(n10306));
  jnot g10114(.din(n10128), .dout(n10307));
  jnot g10115(.din(\a[37] ), .dout(n10308));
  jand g10116(.dina(\a[38] ), .dinb(n10308), .dout(n10309));
  jxor g10117(.dina(n10309), .dinb(n10307), .dout(n10310));
  jnot g10118(.din(n10310), .dout(n10311));
  jxor g10119(.dina(n10311), .dinb(n10306), .dout(n10312));
  jxor g10120(.dina(n10312), .dinb(n10288), .dout(n10313));
  jand g10121(.dina(\a[48] ), .dinb(\a[27] ), .dout(n10314));
  jand g10122(.dina(\a[46] ), .dinb(\a[29] ), .dout(n10315));
  jor  g10123(.dina(n10315), .dinb(n10144), .dout(n10316));
  jnot g10124(.din(n10316), .dout(n10317));
  jand g10125(.dina(\a[47] ), .dinb(\a[29] ), .dout(n10318));
  jand g10126(.dina(n10318), .dinb(n10141), .dout(n10319));
  jor  g10127(.dina(n10319), .dinb(n10317), .dout(n10320));
  jxor g10128(.dina(n10320), .dinb(n10314), .dout(n10321));
  jand g10129(.dina(\a[58] ), .dinb(\a[17] ), .dout(n10322));
  jand g10130(.dina(\a[49] ), .dinb(\a[26] ), .dout(n10323));
  jand g10131(.dina(\a[57] ), .dinb(\a[18] ), .dout(n10324));
  jor  g10132(.dina(n10324), .dinb(n10323), .dout(n10325));
  jnot g10133(.din(n10325), .dout(n10326));
  jand g10134(.dina(\a[57] ), .dinb(\a[26] ), .dout(n10327));
  jand g10135(.dina(n10327), .dinb(n8650), .dout(n10328));
  jor  g10136(.dina(n10328), .dinb(n10326), .dout(n10329));
  jxor g10137(.dina(n10329), .dinb(n10322), .dout(n10330));
  jand g10138(.dina(\a[61] ), .dinb(\a[14] ), .dout(n10331));
  jand g10139(.dina(\a[60] ), .dinb(\a[15] ), .dout(n10332));
  jor  g10140(.dina(n10332), .dinb(n10072), .dout(n10333));
  jand g10141(.dina(\a[60] ), .dinb(\a[16] ), .dout(n10334));
  jand g10142(.dina(n10334), .dinb(n10069), .dout(n10335));
  jnot g10143(.din(n10335), .dout(n10336));
  jand g10144(.dina(n10336), .dinb(n10333), .dout(n10337));
  jxor g10145(.dina(n10337), .dinb(n10331), .dout(n10338));
  jxor g10146(.dina(n10338), .dinb(n10330), .dout(n10339));
  jxor g10147(.dina(n10339), .dinb(n10321), .dout(n10340));
  jxor g10148(.dina(n10340), .dinb(n10313), .dout(n10341));
  jxor g10149(.dina(n10341), .dinb(n10285), .dout(n10342));
  jxor g10150(.dina(n10342), .dinb(n10255), .dout(n10343));
  jand g10151(.dina(n10120), .dinb(n10097), .dout(n10344));
  jand g10152(.dina(n10193), .dinb(n10121), .dout(n10345));
  jor  g10153(.dina(n10345), .dinb(n10344), .dout(n10346));
  jand g10154(.dina(n10091), .dinb(n10088), .dout(n10347));
  jand g10155(.dina(n10092), .dinb(n10085), .dout(n10348));
  jor  g10156(.dina(n10348), .dinb(n10347), .dout(n10349));
  jor  g10157(.dina(n10078), .dinb(n10062), .dout(n10350));
  jor  g10158(.dina(n10084), .dinb(n10080), .dout(n10351));
  jand g10159(.dina(n10351), .dinb(n10350), .dout(n10352));
  jnot g10160(.din(n10352), .dout(n10353));
  jor  g10161(.dina(n10118), .dinb(n10114), .dout(n10354));
  jand g10162(.dina(n10119), .dinb(n10105), .dout(n10355));
  jnot g10163(.din(n10355), .dout(n10356));
  jand g10164(.dina(n10356), .dinb(n10354), .dout(n10357));
  jnot g10165(.din(n10357), .dout(n10358));
  jand g10166(.dina(\a[54] ), .dinb(\a[21] ), .dout(n10359));
  jnot g10167(.din(n10359), .dout(n10360));
  jand g10168(.dina(\a[53] ), .dinb(\a[22] ), .dout(n10361));
  jor  g10169(.dina(n10361), .dinb(n10171), .dout(n10362));
  jand g10170(.dina(\a[53] ), .dinb(\a[24] ), .dout(n10363));
  jand g10171(.dina(n10363), .dinb(n9732), .dout(n10364));
  jnot g10172(.din(n10364), .dout(n10365));
  jand g10173(.dina(n10365), .dinb(n10362), .dout(n10366));
  jxor g10174(.dina(n10366), .dinb(n10360), .dout(n10367));
  jand g10175(.dina(\a[44] ), .dinb(\a[31] ), .dout(n10368));
  jnot g10176(.din(n10368), .dout(n10369));
  jand g10177(.dina(\a[42] ), .dinb(\a[33] ), .dout(n10370));
  jor  g10178(.dina(n10370), .dinb(n10160), .dout(n10371));
  jand g10179(.dina(\a[43] ), .dinb(\a[33] ), .dout(n10372));
  jand g10180(.dina(n10372), .dinb(n10158), .dout(n10373));
  jnot g10181(.din(n10373), .dout(n10374));
  jand g10182(.dina(n10374), .dinb(n10371), .dout(n10375));
  jxor g10183(.dina(n10375), .dinb(n10369), .dout(n10376));
  jand g10184(.dina(\a[41] ), .dinb(\a[34] ), .dout(n10377));
  jnot g10185(.din(n10377), .dout(n10378));
  jand g10186(.dina(\a[55] ), .dinb(\a[20] ), .dout(n10379));
  jand g10187(.dina(\a[50] ), .dinb(\a[25] ), .dout(n10380));
  jxor g10188(.dina(n10380), .dinb(n10379), .dout(n10381));
  jxor g10189(.dina(n10381), .dinb(n10378), .dout(n10382));
  jnot g10190(.din(n10382), .dout(n10383));
  jxor g10191(.dina(n10383), .dinb(n10376), .dout(n10384));
  jxor g10192(.dina(n10384), .dinb(n10367), .dout(n10385));
  jxor g10193(.dina(n10385), .dinb(n10358), .dout(n10386));
  jxor g10194(.dina(n10386), .dinb(n10353), .dout(n10387));
  jxor g10195(.dina(n10387), .dinb(n10349), .dout(n10388));
  jxor g10196(.dina(n10388), .dinb(n10346), .dout(n10389));
  jand g10197(.dina(n10093), .dinb(n10056), .dout(n10390));
  jand g10198(.dina(n10194), .dinb(n10094), .dout(n10391));
  jor  g10199(.dina(n10391), .dinb(n10390), .dout(n10392));
  jxor g10200(.dina(n10392), .dinb(n10389), .dout(n10393));
  jxor g10201(.dina(n10393), .dinb(n10343), .dout(n10394));
  jxor g10202(.dina(n10394), .dinb(n10208), .dout(n10395));
  jand g10203(.dina(n10196), .dinb(n10019), .dout(n10396));
  jnot g10204(.din(n10019), .dout(n10397));
  jnot g10205(.din(n10196), .dout(n10398));
  jand g10206(.dina(n10398), .dinb(n10397), .dout(n10399));
  jnot g10207(.din(n10399), .dout(n10400));
  jand g10208(.dina(n10204), .dinb(n10400), .dout(n10401));
  jor  g10209(.dina(n10401), .dinb(n10396), .dout(n10402));
  jxor g10210(.dina(n10402), .dinb(n10395), .dout(\asquared[76] ));
  jand g10211(.dina(n10392), .dinb(n10389), .dout(n10404));
  jand g10212(.dina(n10393), .dinb(n10343), .dout(n10405));
  jor  g10213(.dina(n10405), .dinb(n10404), .dout(n10406));
  jand g10214(.dina(n10254), .dinb(n10211), .dout(n10407));
  jand g10215(.dina(n10342), .dinb(n10255), .dout(n10408));
  jor  g10216(.dina(n10408), .dinb(n10407), .dout(n10409));
  jand g10217(.dina(n10284), .dinb(n10258), .dout(n10410));
  jand g10218(.dina(n10341), .dinb(n10285), .dout(n10411));
  jor  g10219(.dina(n10411), .dinb(n10410), .dout(n10412));
  jand g10220(.dina(n10229), .dinb(n10226), .dout(n10413));
  jand g10221(.dina(n10253), .dinb(n10230), .dout(n10414));
  jor  g10222(.dina(n10414), .dinb(n10413), .dout(n10415));
  jand g10223(.dina(n10251), .dinb(n10243), .dout(n10416));
  jand g10224(.dina(n10252), .dinb(n10235), .dout(n10417));
  jor  g10225(.dina(n10417), .dinb(n10416), .dout(n10418));
  jand g10226(.dina(n10282), .dinb(n10276), .dout(n10419));
  jand g10227(.dina(n10283), .dinb(n10270), .dout(n10420));
  jor  g10228(.dina(n10420), .dinb(n10419), .dout(n10421));
  jand g10229(.dina(\a[54] ), .dinb(\a[22] ), .dout(n10422));
  jor  g10230(.dina(n10422), .dinb(n10185), .dout(n10423));
  jnot g10231(.din(n10423), .dout(n10424));
  jand g10232(.dina(\a[55] ), .dinb(\a[22] ), .dout(n10425));
  jand g10233(.dina(n10425), .dinb(n10359), .dout(n10426));
  jor  g10234(.dina(n10426), .dinb(n10424), .dout(n10427));
  jxor g10235(.dina(n10427), .dinb(n8603), .dout(n10428));
  jnot g10236(.din(n10428), .dout(n10429));
  jand g10237(.dina(\a[57] ), .dinb(\a[19] ), .dout(n10430));
  jnot g10238(.din(n10430), .dout(n10431));
  jand g10239(.dina(\a[53] ), .dinb(\a[23] ), .dout(n10432));
  jxor g10240(.dina(n10432), .dinb(n10431), .dout(n10433));
  jxor g10241(.dina(n10433), .dinb(n10372), .dout(n10434));
  jnot g10242(.din(n10434), .dout(n10435));
  jand g10243(.dina(\a[63] ), .dinb(\a[13] ), .dout(n10436));
  jand g10244(.dina(\a[45] ), .dinb(\a[31] ), .dout(n10437));
  jand g10245(.dina(\a[44] ), .dinb(\a[32] ), .dout(n10438));
  jor  g10246(.dina(n10438), .dinb(n10437), .dout(n10439));
  jand g10247(.dina(\a[45] ), .dinb(\a[32] ), .dout(n10440));
  jand g10248(.dina(n10440), .dinb(n10368), .dout(n10441));
  jnot g10249(.din(n10441), .dout(n10442));
  jand g10250(.dina(n10442), .dinb(n10439), .dout(n10443));
  jxor g10251(.dina(n10443), .dinb(n10436), .dout(n10444));
  jxor g10252(.dina(n10444), .dinb(n10435), .dout(n10445));
  jxor g10253(.dina(n10445), .dinb(n10429), .dout(n10446));
  jxor g10254(.dina(n10446), .dinb(n10421), .dout(n10447));
  jxor g10255(.dina(n10447), .dinb(n10418), .dout(n10448));
  jxor g10256(.dina(n10448), .dinb(n10415), .dout(n10449));
  jxor g10257(.dina(n10449), .dinb(n10412), .dout(n10450));
  jxor g10258(.dina(n10450), .dinb(n10409), .dout(n10451));
  jand g10259(.dina(n10387), .dinb(n10349), .dout(n10452));
  jand g10260(.dina(n10388), .dinb(n10346), .dout(n10453));
  jor  g10261(.dina(n10453), .dinb(n10452), .dout(n10454));
  jand g10262(.dina(n10247), .dinb(n10245), .dout(n10455));
  jand g10263(.dina(n10250), .dinb(n10248), .dout(n10456));
  jor  g10264(.dina(n10456), .dinb(n10455), .dout(n10457));
  jand g10265(.dina(n10266), .dinb(n10260), .dout(n10458));
  jand g10266(.dina(n10269), .dinb(n10267), .dout(n10459));
  jor  g10267(.dina(n10459), .dinb(n10458), .dout(n10460));
  jxor g10268(.dina(n10460), .dinb(n10457), .dout(n10461));
  jand g10269(.dina(n10241), .dinb(n10239), .dout(n10462));
  jand g10270(.dina(n10242), .dinb(n10237), .dout(n10463));
  jor  g10271(.dina(n10463), .dinb(n10462), .dout(n10464));
  jxor g10272(.dina(n10464), .dinb(n10461), .dout(n10465));
  jand g10273(.dina(n10312), .dinb(n10288), .dout(n10466));
  jand g10274(.dina(n10340), .dinb(n10313), .dout(n10467));
  jor  g10275(.dina(n10467), .dinb(n10466), .dout(n10468));
  jxor g10276(.dina(n10468), .dinb(n10465), .dout(n10469));
  jand g10277(.dina(n10304), .dinb(n10298), .dout(n10470));
  jor  g10278(.dina(n10470), .dinb(n10302), .dout(n10471));
  jand g10279(.dina(n10316), .dinb(n10314), .dout(n10472));
  jor  g10280(.dina(n10472), .dinb(n10319), .dout(n10473));
  jnot g10281(.din(n10379), .dout(n10474));
  jnot g10282(.din(n10380), .dout(n10475));
  jand g10283(.dina(n10475), .dinb(n10474), .dout(n10476));
  jnot g10284(.din(n10476), .dout(n10477));
  jand g10285(.dina(n10380), .dinb(n10379), .dout(n10478));
  jor  g10286(.dina(n10478), .dinb(n10377), .dout(n10479));
  jand g10287(.dina(n10479), .dinb(n10477), .dout(n10480));
  jxor g10288(.dina(n10480), .dinb(n10473), .dout(n10481));
  jxor g10289(.dina(n10481), .dinb(n10471), .dout(n10482));
  jnot g10290(.din(\a[38] ), .dout(n10483));
  jand g10291(.dina(n10307), .dinb(n10308), .dout(n10484));
  jor  g10292(.dina(n10484), .dinb(n10483), .dout(n10485));
  jnot g10293(.din(n10485), .dout(n10486));
  jand g10294(.dina(\a[62] ), .dinb(\a[14] ), .dout(n10487));
  jxor g10295(.dina(n10487), .dinb(n10486), .dout(n10488));
  jand g10296(.dina(n10291), .dinb(n10289), .dout(n10489));
  jor  g10297(.dina(n10489), .dinb(n10294), .dout(n10490));
  jxor g10298(.dina(n10490), .dinb(n10488), .dout(n10491));
  jnot g10299(.din(n10491), .dout(n10492));
  jnot g10300(.din(n10376), .dout(n10493));
  jand g10301(.dina(n10383), .dinb(n10493), .dout(n10494));
  jnot g10302(.din(n10494), .dout(n10495));
  jand g10303(.dina(n10382), .dinb(n10376), .dout(n10496));
  jor  g10304(.dina(n10496), .dinb(n10367), .dout(n10497));
  jand g10305(.dina(n10497), .dinb(n10495), .dout(n10498));
  jxor g10306(.dina(n10498), .dinb(n10492), .dout(n10499));
  jxor g10307(.dina(n10499), .dinb(n10482), .dout(n10500));
  jxor g10308(.dina(n10500), .dinb(n10469), .dout(n10501));
  jxor g10309(.dina(n10501), .dinb(n10454), .dout(n10502));
  jand g10310(.dina(n10385), .dinb(n10358), .dout(n10503));
  jand g10311(.dina(n10386), .dinb(n10353), .dout(n10504));
  jor  g10312(.dina(n10504), .dinb(n10503), .dout(n10505));
  jand g10313(.dina(n10337), .dinb(n10331), .dout(n10506));
  jor  g10314(.dina(n10506), .dinb(n10335), .dout(n10507));
  jand g10315(.dina(n10325), .dinb(n10322), .dout(n10508));
  jor  g10316(.dina(n10508), .dinb(n10328), .dout(n10509));
  jxor g10317(.dina(n10509), .dinb(n10507), .dout(n10510));
  jand g10318(.dina(n10371), .dinb(n10368), .dout(n10511));
  jor  g10319(.dina(n10511), .dinb(n10373), .dout(n10512));
  jxor g10320(.dina(n10512), .dinb(n10510), .dout(n10513));
  jnot g10321(.din(n10330), .dout(n10514));
  jor  g10322(.dina(n10338), .dinb(n10514), .dout(n10515));
  jnot g10323(.din(n10321), .dout(n10516));
  jand g10324(.dina(n10338), .dinb(n10514), .dout(n10517));
  jor  g10325(.dina(n10517), .dinb(n10516), .dout(n10518));
  jand g10326(.dina(n10518), .dinb(n10515), .dout(n10519));
  jor  g10327(.dina(n10305), .dinb(n10297), .dout(n10520));
  jand g10328(.dina(n10305), .dinb(n10297), .dout(n10521));
  jor  g10329(.dina(n10311), .dinb(n10521), .dout(n10522));
  jand g10330(.dina(n10522), .dinb(n10520), .dout(n10523));
  jxor g10331(.dina(n10523), .dinb(n10519), .dout(n10524));
  jxor g10332(.dina(n10524), .dinb(n10513), .dout(n10525));
  jxor g10333(.dina(n10525), .dinb(n10505), .dout(n10526));
  jand g10334(.dina(n10221), .dinb(n10214), .dout(n10527));
  jand g10335(.dina(n10225), .dinb(n10222), .dout(n10528));
  jor  g10336(.dina(n10528), .dinb(n10527), .dout(n10529));
  jand g10337(.dina(\a[39] ), .dinb(\a[37] ), .dout(n10530));
  jand g10338(.dina(\a[51] ), .dinb(\a[25] ), .dout(n10531));
  jand g10339(.dina(\a[52] ), .dinb(\a[24] ), .dout(n10532));
  jor  g10340(.dina(n10532), .dinb(n10531), .dout(n10533));
  jnot g10341(.din(n10533), .dout(n10534));
  jand g10342(.dina(\a[52] ), .dinb(\a[25] ), .dout(n10535));
  jand g10343(.dina(n10535), .dinb(n10171), .dout(n10536));
  jor  g10344(.dina(n10536), .dinb(n10534), .dout(n10537));
  jxor g10345(.dina(n10537), .dinb(n10530), .dout(n10538));
  jand g10346(.dina(\a[42] ), .dinb(\a[34] ), .dout(n10539));
  jand g10347(.dina(\a[41] ), .dinb(\a[35] ), .dout(n10540));
  jor  g10348(.dina(n10540), .dinb(n10293), .dout(n10541));
  jnot g10349(.din(n10541), .dout(n10542));
  jand g10350(.dina(\a[41] ), .dinb(\a[36] ), .dout(n10543));
  jand g10351(.dina(n10543), .dinb(n10179), .dout(n10544));
  jor  g10352(.dina(n10544), .dinb(n10542), .dout(n10545));
  jxor g10353(.dina(n10545), .dinb(n10539), .dout(n10546));
  jand g10354(.dina(\a[48] ), .dinb(\a[28] ), .dout(n10547));
  jand g10355(.dina(\a[46] ), .dinb(\a[30] ), .dout(n10548));
  jor  g10356(.dina(n10548), .dinb(n10318), .dout(n10549));
  jand g10357(.dina(\a[47] ), .dinb(\a[30] ), .dout(n10550));
  jand g10358(.dina(n10550), .dinb(n10315), .dout(n10551));
  jnot g10359(.din(n10551), .dout(n10552));
  jand g10360(.dina(n10552), .dinb(n10549), .dout(n10553));
  jxor g10361(.dina(n10553), .dinb(n10547), .dout(n10554));
  jxor g10362(.dina(n10554), .dinb(n10546), .dout(n10555));
  jxor g10363(.dina(n10555), .dinb(n10538), .dout(n10556));
  jxor g10364(.dina(n10556), .dinb(n10529), .dout(n10557));
  jand g10365(.dina(\a[58] ), .dinb(\a[18] ), .dout(n10558));
  jand g10366(.dina(\a[50] ), .dinb(\a[26] ), .dout(n10559));
  jand g10367(.dina(\a[49] ), .dinb(\a[27] ), .dout(n10560));
  jor  g10368(.dina(n10560), .dinb(n10559), .dout(n10561));
  jnot g10369(.din(n10561), .dout(n10562));
  jand g10370(.dina(\a[50] ), .dinb(\a[27] ), .dout(n10563));
  jand g10371(.dina(n10563), .dinb(n10323), .dout(n10564));
  jor  g10372(.dina(n10564), .dinb(n10562), .dout(n10565));
  jxor g10373(.dina(n10565), .dinb(n10558), .dout(n10566));
  jnot g10374(.din(n10566), .dout(n10567));
  jand g10375(.dina(\a[61] ), .dinb(\a[15] ), .dout(n10568));
  jand g10376(.dina(\a[59] ), .dinb(\a[17] ), .dout(n10569));
  jor  g10377(.dina(n10569), .dinb(n10334), .dout(n10570));
  jnot g10378(.din(n10570), .dout(n10571));
  jand g10379(.dina(\a[60] ), .dinb(\a[17] ), .dout(n10572));
  jand g10380(.dina(n10572), .dinb(n10072), .dout(n10573));
  jor  g10381(.dina(n10573), .dinb(n10571), .dout(n10574));
  jxor g10382(.dina(n10574), .dinb(n10568), .dout(n10575));
  jnot g10383(.din(n10575), .dout(n10576));
  jand g10384(.dina(n10362), .dinb(n10359), .dout(n10577));
  jor  g10385(.dina(n10577), .dinb(n10364), .dout(n10578));
  jxor g10386(.dina(n10578), .dinb(n10576), .dout(n10579));
  jxor g10387(.dina(n10579), .dinb(n10567), .dout(n10580));
  jxor g10388(.dina(n10580), .dinb(n10557), .dout(n10581));
  jxor g10389(.dina(n10581), .dinb(n10526), .dout(n10582));
  jxor g10390(.dina(n10582), .dinb(n10502), .dout(n10583));
  jxor g10391(.dina(n10583), .dinb(n10451), .dout(n10584));
  jxor g10392(.dina(n10584), .dinb(n10406), .dout(n10585));
  jand g10393(.dina(n10394), .dinb(n10208), .dout(n10586));
  jor  g10394(.dina(n10394), .dinb(n10208), .dout(n10587));
  jand g10395(.dina(n10402), .dinb(n10587), .dout(n10588));
  jor  g10396(.dina(n10588), .dinb(n10586), .dout(n10589));
  jxor g10397(.dina(n10589), .dinb(n10585), .dout(\asquared[77] ));
  jand g10398(.dina(n10450), .dinb(n10409), .dout(n10591));
  jand g10399(.dina(n10583), .dinb(n10451), .dout(n10592));
  jor  g10400(.dina(n10592), .dinb(n10591), .dout(n10593));
  jand g10401(.dina(n10501), .dinb(n10454), .dout(n10594));
  jand g10402(.dina(n10582), .dinb(n10502), .dout(n10595));
  jor  g10403(.dina(n10595), .dinb(n10594), .dout(n10596));
  jand g10404(.dina(n10525), .dinb(n10505), .dout(n10597));
  jand g10405(.dina(n10581), .dinb(n10526), .dout(n10598));
  jor  g10406(.dina(n10598), .dinb(n10597), .dout(n10599));
  jand g10407(.dina(n10468), .dinb(n10465), .dout(n10600));
  jand g10408(.dina(n10500), .dinb(n10469), .dout(n10601));
  jor  g10409(.dina(n10601), .dinb(n10600), .dout(n10602));
  jor  g10410(.dina(n10498), .dinb(n10492), .dout(n10603));
  jand g10411(.dina(n10499), .dinb(n10482), .dout(n10604));
  jnot g10412(.din(n10604), .dout(n10605));
  jand g10413(.dina(n10605), .dinb(n10603), .dout(n10606));
  jnot g10414(.din(n10606), .dout(n10607));
  jand g10415(.dina(n10523), .dinb(n10519), .dout(n10608));
  jand g10416(.dina(n10524), .dinb(n10513), .dout(n10609));
  jor  g10417(.dina(n10609), .dinb(n10608), .dout(n10610));
  jand g10418(.dina(\a[61] ), .dinb(\a[16] ), .dout(n10611));
  jnot g10419(.din(n10611), .dout(n10612));
  jand g10420(.dina(\a[44] ), .dinb(\a[33] ), .dout(n10613));
  jor  g10421(.dina(n10613), .dinb(n10440), .dout(n10614));
  jand g10422(.dina(\a[45] ), .dinb(\a[33] ), .dout(n10615));
  jand g10423(.dina(n10615), .dinb(n10438), .dout(n10616));
  jnot g10424(.din(n10616), .dout(n10617));
  jand g10425(.dina(n10617), .dinb(n10614), .dout(n10618));
  jxor g10426(.dina(n10618), .dinb(n10612), .dout(n10619));
  jnot g10427(.din(n10535), .dout(n10620));
  jand g10428(.dina(\a[54] ), .dinb(\a[23] ), .dout(n10621));
  jor  g10429(.dina(n10621), .dinb(n10363), .dout(n10622));
  jand g10430(.dina(n10432), .dinb(n9911), .dout(n10623));
  jnot g10431(.din(n10623), .dout(n10624));
  jand g10432(.dina(n10624), .dinb(n10622), .dout(n10625));
  jxor g10433(.dina(n10625), .dinb(n10620), .dout(n10626));
  jand g10434(.dina(\a[43] ), .dinb(\a[34] ), .dout(n10627));
  jnot g10435(.din(n10627), .dout(n10628));
  jand g10436(.dina(\a[51] ), .dinb(\a[26] ), .dout(n10629));
  jxor g10437(.dina(n10629), .dinb(n10425), .dout(n10630));
  jxor g10438(.dina(n10630), .dinb(n10628), .dout(n10631));
  jnot g10439(.din(n10631), .dout(n10632));
  jxor g10440(.dina(n10632), .dinb(n10626), .dout(n10633));
  jxor g10441(.dina(n10633), .dinb(n10619), .dout(n10634));
  jxor g10442(.dina(n10634), .dinb(n10610), .dout(n10635));
  jxor g10443(.dina(n10635), .dinb(n10607), .dout(n10636));
  jxor g10444(.dina(n10636), .dinb(n10602), .dout(n10637));
  jxor g10445(.dina(n10637), .dinb(n10599), .dout(n10638));
  jxor g10446(.dina(n10638), .dinb(n10596), .dout(n10639));
  jand g10447(.dina(n10448), .dinb(n10415), .dout(n10640));
  jand g10448(.dina(n10449), .dinb(n10412), .dout(n10641));
  jor  g10449(.dina(n10641), .dinb(n10640), .dout(n10642));
  jand g10450(.dina(n10509), .dinb(n10507), .dout(n10643));
  jand g10451(.dina(n10512), .dinb(n10510), .dout(n10644));
  jor  g10452(.dina(n10644), .dinb(n10643), .dout(n10645));
  jand g10453(.dina(\a[59] ), .dinb(\a[18] ), .dout(n10646));
  jor  g10454(.dina(n10646), .dinb(n10572), .dout(n10647));
  jand g10455(.dina(\a[60] ), .dinb(\a[18] ), .dout(n10648));
  jand g10456(.dina(n10648), .dinb(n10569), .dout(n10649));
  jnot g10457(.din(n10649), .dout(n10650));
  jand g10458(.dina(n10650), .dinb(n10647), .dout(n10651));
  jand g10459(.dina(n10533), .dinb(n10530), .dout(n10652));
  jor  g10460(.dina(n10652), .dinb(n10536), .dout(n10653));
  jxor g10461(.dina(n10653), .dinb(n10651), .dout(n10654));
  jxor g10462(.dina(n10654), .dinb(n10645), .dout(n10655));
  jand g10463(.dina(n10480), .dinb(n10473), .dout(n10656));
  jand g10464(.dina(n10481), .dinb(n10471), .dout(n10657));
  jor  g10465(.dina(n10657), .dinb(n10656), .dout(n10658));
  jxor g10466(.dina(n10658), .dinb(n10655), .dout(n10659));
  jand g10467(.dina(n10556), .dinb(n10529), .dout(n10660));
  jand g10468(.dina(n10580), .dinb(n10557), .dout(n10661));
  jor  g10469(.dina(n10661), .dinb(n10660), .dout(n10662));
  jxor g10470(.dina(n10662), .dinb(n10659), .dout(n10663));
  jand g10471(.dina(n10443), .dinb(n10436), .dout(n10664));
  jor  g10472(.dina(n10664), .dinb(n10441), .dout(n10665));
  jand g10473(.dina(n10553), .dinb(n10547), .dout(n10666));
  jor  g10474(.dina(n10666), .dinb(n10551), .dout(n10667));
  jand g10475(.dina(n10423), .dinb(n8603), .dout(n10668));
  jor  g10476(.dina(n10668), .dinb(n10426), .dout(n10669));
  jxor g10477(.dina(n10669), .dinb(n10667), .dout(n10670));
  jxor g10478(.dina(n10670), .dinb(n10665), .dout(n10671));
  jand g10479(.dina(n10561), .dinb(n10558), .dout(n10672));
  jor  g10480(.dina(n10672), .dinb(n10564), .dout(n10673));
  jand g10481(.dina(n10570), .dinb(n10568), .dout(n10674));
  jor  g10482(.dina(n10674), .dinb(n10573), .dout(n10675));
  jxor g10483(.dina(n10675), .dinb(n10673), .dout(n10676));
  jnot g10484(.din(n10432), .dout(n10677));
  jand g10485(.dina(n10677), .dinb(n10431), .dout(n10678));
  jnot g10486(.din(n10678), .dout(n10679));
  jand g10487(.dina(n10432), .dinb(n10430), .dout(n10680));
  jor  g10488(.dina(n10680), .dinb(n10372), .dout(n10681));
  jand g10489(.dina(n10681), .dinb(n10679), .dout(n10682));
  jxor g10490(.dina(n10682), .dinb(n10676), .dout(n10683));
  jor  g10491(.dina(n10444), .dinb(n10435), .dout(n10684));
  jand g10492(.dina(n10444), .dinb(n10435), .dout(n10685));
  jor  g10493(.dina(n10685), .dinb(n10429), .dout(n10686));
  jand g10494(.dina(n10686), .dinb(n10684), .dout(n10687));
  jxor g10495(.dina(n10687), .dinb(n10683), .dout(n10688));
  jxor g10496(.dina(n10688), .dinb(n10671), .dout(n10689));
  jxor g10497(.dina(n10689), .dinb(n10663), .dout(n10690));
  jxor g10498(.dina(n10690), .dinb(n10642), .dout(n10691));
  jand g10499(.dina(n10487), .dinb(n10486), .dout(n10692));
  jand g10500(.dina(n10490), .dinb(n10488), .dout(n10693));
  jor  g10501(.dina(n10693), .dinb(n10692), .dout(n10694));
  jand g10502(.dina(n10578), .dinb(n10576), .dout(n10695));
  jand g10503(.dina(n10579), .dinb(n10567), .dout(n10696));
  jor  g10504(.dina(n10696), .dinb(n10695), .dout(n10697));
  jxor g10505(.dina(n10697), .dinb(n10694), .dout(n10698));
  jnot g10506(.din(n10546), .dout(n10699));
  jor  g10507(.dina(n10554), .dinb(n10699), .dout(n10700));
  jnot g10508(.din(n10538), .dout(n10701));
  jand g10509(.dina(n10554), .dinb(n10699), .dout(n10702));
  jor  g10510(.dina(n10702), .dinb(n10701), .dout(n10703));
  jand g10511(.dina(n10703), .dinb(n10700), .dout(n10704));
  jxor g10512(.dina(n10704), .dinb(n10698), .dout(n10705));
  jand g10513(.dina(n10446), .dinb(n10421), .dout(n10706));
  jand g10514(.dina(n10447), .dinb(n10418), .dout(n10707));
  jor  g10515(.dina(n10707), .dinb(n10706), .dout(n10708));
  jxor g10516(.dina(n10708), .dinb(n10705), .dout(n10709));
  jand g10517(.dina(n10460), .dinb(n10457), .dout(n10710));
  jand g10518(.dina(n10464), .dinb(n10461), .dout(n10711));
  jor  g10519(.dina(n10711), .dinb(n10710), .dout(n10712));
  jand g10520(.dina(\a[42] ), .dinb(\a[35] ), .dout(n10713));
  jand g10521(.dina(\a[40] ), .dinb(\a[37] ), .dout(n10714));
  jor  g10522(.dina(n10714), .dinb(n10543), .dout(n10715));
  jnot g10523(.din(n10715), .dout(n10716));
  jand g10524(.dina(\a[41] ), .dinb(\a[37] ), .dout(n10717));
  jand g10525(.dina(n10717), .dinb(n10293), .dout(n10718));
  jor  g10526(.dina(n10718), .dinb(n10716), .dout(n10719));
  jxor g10527(.dina(n10719), .dinb(n10713), .dout(n10720));
  jnot g10528(.din(n10720), .dout(n10721));
  jand g10529(.dina(\a[63] ), .dinb(\a[14] ), .dout(n10722));
  jand g10530(.dina(\a[46] ), .dinb(\a[31] ), .dout(n10723));
  jor  g10531(.dina(n10723), .dinb(n10722), .dout(n10724));
  jand g10532(.dina(\a[63] ), .dinb(\a[31] ), .dout(n10725));
  jand g10533(.dina(n10725), .dinb(n6074), .dout(n10726));
  jnot g10534(.din(n10726), .dout(n10727));
  jand g10535(.dina(n10727), .dinb(n10724), .dout(n10728));
  jxor g10536(.dina(n10728), .dinb(n10550), .dout(n10729));
  jxor g10537(.dina(n10729), .dinb(n10721), .dout(n10730));
  jand g10538(.dina(\a[62] ), .dinb(\a[15] ), .dout(n10731));
  jnot g10539(.din(n10731), .dout(n10732));
  jand g10540(.dina(\a[39] ), .dinb(n10483), .dout(n10733));
  jxor g10541(.dina(n10733), .dinb(n10732), .dout(n10734));
  jnot g10542(.din(n10734), .dout(n10735));
  jxor g10543(.dina(n10735), .dinb(n10730), .dout(n10736));
  jxor g10544(.dina(n10736), .dinb(n10712), .dout(n10737));
  jand g10545(.dina(\a[49] ), .dinb(\a[28] ), .dout(n10738));
  jand g10546(.dina(\a[48] ), .dinb(\a[29] ), .dout(n10739));
  jor  g10547(.dina(n10739), .dinb(n10738), .dout(n10740));
  jnot g10548(.din(n10740), .dout(n10741));
  jand g10549(.dina(\a[49] ), .dinb(\a[29] ), .dout(n10742));
  jand g10550(.dina(n10742), .dinb(n10547), .dout(n10743));
  jor  g10551(.dina(n10743), .dinb(n10741), .dout(n10744));
  jxor g10552(.dina(n10744), .dinb(n10563), .dout(n10745));
  jnot g10553(.din(n10745), .dout(n10746));
  jand g10554(.dina(\a[58] ), .dinb(\a[19] ), .dout(n10747));
  jand g10555(.dina(\a[57] ), .dinb(\a[20] ), .dout(n10748));
  jand g10556(.dina(\a[56] ), .dinb(\a[21] ), .dout(n10749));
  jor  g10557(.dina(n10749), .dinb(n10748), .dout(n10750));
  jnot g10558(.din(n10750), .dout(n10751));
  jand g10559(.dina(\a[57] ), .dinb(\a[21] ), .dout(n10752));
  jand g10560(.dina(n10752), .dinb(n8603), .dout(n10753));
  jor  g10561(.dina(n10753), .dinb(n10751), .dout(n10754));
  jxor g10562(.dina(n10754), .dinb(n10747), .dout(n10755));
  jnot g10563(.din(n10755), .dout(n10756));
  jand g10564(.dina(n10541), .dinb(n10539), .dout(n10757));
  jor  g10565(.dina(n10757), .dinb(n10544), .dout(n10758));
  jxor g10566(.dina(n10758), .dinb(n10756), .dout(n10759));
  jxor g10567(.dina(n10759), .dinb(n10746), .dout(n10760));
  jxor g10568(.dina(n10760), .dinb(n10737), .dout(n10761));
  jxor g10569(.dina(n10761), .dinb(n10709), .dout(n10762));
  jxor g10570(.dina(n10762), .dinb(n10691), .dout(n10763));
  jxor g10571(.dina(n10763), .dinb(n10639), .dout(n10764));
  jxor g10572(.dina(n10764), .dinb(n10593), .dout(n10765));
  jand g10573(.dina(n10584), .dinb(n10406), .dout(n10766));
  jor  g10574(.dina(n10584), .dinb(n10406), .dout(n10767));
  jand g10575(.dina(n10589), .dinb(n10767), .dout(n10768));
  jor  g10576(.dina(n10768), .dinb(n10766), .dout(n10769));
  jxor g10577(.dina(n10769), .dinb(n10765), .dout(\asquared[78] ));
  jand g10578(.dina(n10638), .dinb(n10596), .dout(n10771));
  jand g10579(.dina(n10763), .dinb(n10639), .dout(n10772));
  jor  g10580(.dina(n10772), .dinb(n10771), .dout(n10773));
  jand g10581(.dina(n10708), .dinb(n10705), .dout(n10774));
  jand g10582(.dina(n10761), .dinb(n10709), .dout(n10775));
  jor  g10583(.dina(n10775), .dinb(n10774), .dout(n10776));
  jand g10584(.dina(n10662), .dinb(n10659), .dout(n10777));
  jand g10585(.dina(n10689), .dinb(n10663), .dout(n10778));
  jor  g10586(.dina(n10778), .dinb(n10777), .dout(n10779));
  jand g10587(.dina(n10697), .dinb(n10694), .dout(n10780));
  jand g10588(.dina(n10704), .dinb(n10698), .dout(n10781));
  jor  g10589(.dina(n10781), .dinb(n10780), .dout(n10782));
  jand g10590(.dina(\a[63] ), .dinb(\a[15] ), .dout(n10783));
  jand g10591(.dina(\a[62] ), .dinb(\a[16] ), .dout(n10784));
  jand g10592(.dina(\a[61] ), .dinb(\a[17] ), .dout(n10785));
  jor  g10593(.dina(n10785), .dinb(n10784), .dout(n10786));
  jnot g10594(.din(n10786), .dout(n10787));
  jand g10595(.dina(\a[62] ), .dinb(\a[17] ), .dout(n10788));
  jand g10596(.dina(n10788), .dinb(n10611), .dout(n10789));
  jor  g10597(.dina(n10789), .dinb(n10787), .dout(n10790));
  jxor g10598(.dina(n10790), .dinb(n10783), .dout(n10791));
  jand g10599(.dina(\a[51] ), .dinb(\a[27] ), .dout(n10792));
  jand g10600(.dina(\a[50] ), .dinb(\a[28] ), .dout(n10793));
  jor  g10601(.dina(n10793), .dinb(n10742), .dout(n10794));
  jnot g10602(.din(n10794), .dout(n10795));
  jand g10603(.dina(\a[50] ), .dinb(\a[29] ), .dout(n10796));
  jand g10604(.dina(n10796), .dinb(n10738), .dout(n10797));
  jor  g10605(.dina(n10797), .dinb(n10795), .dout(n10798));
  jxor g10606(.dina(n10798), .dinb(n10792), .dout(n10799));
  jand g10607(.dina(\a[59] ), .dinb(\a[19] ), .dout(n10800));
  jor  g10608(.dina(n10800), .dinb(n10752), .dout(n10801));
  jand g10609(.dina(\a[59] ), .dinb(\a[21] ), .dout(n10802));
  jand g10610(.dina(n10802), .dinb(n10430), .dout(n10803));
  jnot g10611(.din(n10803), .dout(n10804));
  jand g10612(.dina(n10804), .dinb(n10801), .dout(n10805));
  jxor g10613(.dina(n10805), .dinb(n10648), .dout(n10806));
  jxor g10614(.dina(n10806), .dinb(n10799), .dout(n10807));
  jxor g10615(.dina(n10807), .dinb(n10791), .dout(n10808));
  jand g10616(.dina(\a[53] ), .dinb(\a[25] ), .dout(n10809));
  jand g10617(.dina(\a[56] ), .dinb(\a[22] ), .dout(n10810));
  jor  g10618(.dina(n10810), .dinb(n9911), .dout(n10811));
  jnot g10619(.din(n10811), .dout(n10812));
  jand g10620(.dina(\a[56] ), .dinb(\a[24] ), .dout(n10813));
  jand g10621(.dina(n10813), .dinb(n10422), .dout(n10814));
  jor  g10622(.dina(n10814), .dinb(n10812), .dout(n10815));
  jxor g10623(.dina(n10815), .dinb(n10809), .dout(n10816));
  jnot g10624(.din(n10816), .dout(n10817));
  jand g10625(.dina(\a[58] ), .dinb(\a[20] ), .dout(n10818));
  jand g10626(.dina(\a[48] ), .dinb(\a[30] ), .dout(n10819));
  jand g10627(.dina(\a[47] ), .dinb(\a[31] ), .dout(n10820));
  jor  g10628(.dina(n10820), .dinb(n10819), .dout(n10821));
  jand g10629(.dina(\a[48] ), .dinb(\a[31] ), .dout(n10822));
  jand g10630(.dina(n10822), .dinb(n10550), .dout(n10823));
  jnot g10631(.din(n10823), .dout(n10824));
  jand g10632(.dina(n10824), .dinb(n10821), .dout(n10825));
  jxor g10633(.dina(n10825), .dinb(n10818), .dout(n10826));
  jand g10634(.dina(\a[46] ), .dinb(\a[32] ), .dout(n10827));
  jand g10635(.dina(\a[44] ), .dinb(\a[34] ), .dout(n10828));
  jor  g10636(.dina(n10828), .dinb(n10615), .dout(n10829));
  jand g10637(.dina(\a[45] ), .dinb(\a[34] ), .dout(n10830));
  jand g10638(.dina(n10830), .dinb(n10613), .dout(n10831));
  jnot g10639(.din(n10831), .dout(n10832));
  jand g10640(.dina(n10832), .dinb(n10829), .dout(n10833));
  jxor g10641(.dina(n10833), .dinb(n10827), .dout(n10834));
  jxor g10642(.dina(n10834), .dinb(n10826), .dout(n10835));
  jxor g10643(.dina(n10835), .dinb(n10817), .dout(n10836));
  jxor g10644(.dina(n10836), .dinb(n10808), .dout(n10837));
  jxor g10645(.dina(n10837), .dinb(n10782), .dout(n10838));
  jxor g10646(.dina(n10838), .dinb(n10779), .dout(n10839));
  jxor g10647(.dina(n10839), .dinb(n10776), .dout(n10840));
  jand g10648(.dina(n10690), .dinb(n10642), .dout(n10841));
  jand g10649(.dina(n10762), .dinb(n10691), .dout(n10842));
  jor  g10650(.dina(n10842), .dinb(n10841), .dout(n10843));
  jxor g10651(.dina(n10843), .dinb(n10840), .dout(n10844));
  jand g10652(.dina(n10636), .dinb(n10602), .dout(n10845));
  jand g10653(.dina(n10637), .dinb(n10599), .dout(n10846));
  jor  g10654(.dina(n10846), .dinb(n10845), .dout(n10847));
  jand g10655(.dina(n10758), .dinb(n10756), .dout(n10848));
  jand g10656(.dina(n10759), .dinb(n10746), .dout(n10849));
  jor  g10657(.dina(n10849), .dinb(n10848), .dout(n10850));
  jor  g10658(.dina(n10729), .dinb(n10721), .dout(n10851));
  jand g10659(.dina(n10729), .dinb(n10721), .dout(n10852));
  jor  g10660(.dina(n10735), .dinb(n10852), .dout(n10853));
  jand g10661(.dina(n10853), .dinb(n10851), .dout(n10854));
  jxor g10662(.dina(n10854), .dinb(n10850), .dout(n10855));
  jnot g10663(.din(n10855), .dout(n10856));
  jnot g10664(.din(n10626), .dout(n10857));
  jand g10665(.dina(n10632), .dinb(n10857), .dout(n10858));
  jnot g10666(.din(n10858), .dout(n10859));
  jand g10667(.dina(n10631), .dinb(n10626), .dout(n10860));
  jor  g10668(.dina(n10860), .dinb(n10619), .dout(n10861));
  jand g10669(.dina(n10861), .dinb(n10859), .dout(n10862));
  jxor g10670(.dina(n10862), .dinb(n10856), .dout(n10863));
  jand g10671(.dina(n10687), .dinb(n10683), .dout(n10864));
  jand g10672(.dina(n10688), .dinb(n10671), .dout(n10865));
  jor  g10673(.dina(n10865), .dinb(n10864), .dout(n10866));
  jxor g10674(.dina(n10866), .dinb(n10863), .dout(n10867));
  jnot g10675(.din(\a[39] ), .dout(n10868));
  jand g10676(.dina(n10732), .dinb(n10483), .dout(n10869));
  jor  g10677(.dina(n10869), .dinb(n10868), .dout(n10870));
  jnot g10678(.din(n10870), .dout(n10871));
  jand g10679(.dina(n10715), .dinb(n10713), .dout(n10872));
  jor  g10680(.dina(n10872), .dinb(n10718), .dout(n10873));
  jxor g10681(.dina(n10873), .dinb(n10871), .dout(n10874));
  jand g10682(.dina(n10622), .dinb(n10535), .dout(n10875));
  jor  g10683(.dina(n10875), .dinb(n10623), .dout(n10876));
  jxor g10684(.dina(n10876), .dinb(n10874), .dout(n10877));
  jand g10685(.dina(n10728), .dinb(n10550), .dout(n10878));
  jor  g10686(.dina(n10878), .dinb(n10726), .dout(n10879));
  jand g10687(.dina(n10740), .dinb(n10563), .dout(n10880));
  jor  g10688(.dina(n10880), .dinb(n10743), .dout(n10881));
  jxor g10689(.dina(n10881), .dinb(n10879), .dout(n10882));
  jand g10690(.dina(n10614), .dinb(n10611), .dout(n10883));
  jor  g10691(.dina(n10883), .dinb(n10616), .dout(n10884));
  jxor g10692(.dina(n10884), .dinb(n10882), .dout(n10885));
  jand g10693(.dina(n10675), .dinb(n10673), .dout(n10886));
  jand g10694(.dina(n10682), .dinb(n10676), .dout(n10887));
  jor  g10695(.dina(n10887), .dinb(n10886), .dout(n10888));
  jxor g10696(.dina(n10888), .dinb(n10885), .dout(n10889));
  jxor g10697(.dina(n10889), .dinb(n10877), .dout(n10890));
  jxor g10698(.dina(n10890), .dinb(n10867), .dout(n10891));
  jxor g10699(.dina(n10891), .dinb(n10847), .dout(n10892));
  jand g10700(.dina(n10669), .dinb(n10667), .dout(n10893));
  jand g10701(.dina(n10670), .dinb(n10665), .dout(n10894));
  jor  g10702(.dina(n10894), .dinb(n10893), .dout(n10895));
  jand g10703(.dina(\a[55] ), .dinb(\a[23] ), .dout(n10896));
  jand g10704(.dina(\a[43] ), .dinb(\a[35] ), .dout(n10897));
  jand g10705(.dina(\a[42] ), .dinb(\a[36] ), .dout(n10898));
  jor  g10706(.dina(n10898), .dinb(n10897), .dout(n10899));
  jand g10707(.dina(\a[43] ), .dinb(\a[36] ), .dout(n10900));
  jand g10708(.dina(n10900), .dinb(n10713), .dout(n10901));
  jnot g10709(.din(n10901), .dout(n10902));
  jand g10710(.dina(n10902), .dinb(n10899), .dout(n10903));
  jxor g10711(.dina(n10903), .dinb(n10896), .dout(n10904));
  jnot g10712(.din(n10904), .dout(n10905));
  jand g10713(.dina(\a[40] ), .dinb(\a[38] ), .dout(n10906));
  jnot g10714(.din(n10906), .dout(n10907));
  jand g10715(.dina(\a[52] ), .dinb(\a[26] ), .dout(n10908));
  jxor g10716(.dina(n10908), .dinb(n10907), .dout(n10909));
  jxor g10717(.dina(n10909), .dinb(n10717), .dout(n10910));
  jxor g10718(.dina(n10910), .dinb(n10905), .dout(n10911));
  jxor g10719(.dina(n10911), .dinb(n10895), .dout(n10912));
  jand g10720(.dina(n10750), .dinb(n10747), .dout(n10913));
  jor  g10721(.dina(n10913), .dinb(n10753), .dout(n10914));
  jnot g10722(.din(n10425), .dout(n10915));
  jnot g10723(.din(n10629), .dout(n10916));
  jand g10724(.dina(n10916), .dinb(n10915), .dout(n10917));
  jnot g10725(.din(n10917), .dout(n10918));
  jand g10726(.dina(n10629), .dinb(n10425), .dout(n10919));
  jor  g10727(.dina(n10919), .dinb(n10627), .dout(n10920));
  jand g10728(.dina(n10920), .dinb(n10918), .dout(n10921));
  jxor g10729(.dina(n10921), .dinb(n10914), .dout(n10922));
  jand g10730(.dina(n10653), .dinb(n10651), .dout(n10923));
  jor  g10731(.dina(n10923), .dinb(n10649), .dout(n10924));
  jxor g10732(.dina(n10924), .dinb(n10922), .dout(n10925));
  jand g10733(.dina(n10654), .dinb(n10645), .dout(n10926));
  jand g10734(.dina(n10658), .dinb(n10655), .dout(n10927));
  jor  g10735(.dina(n10927), .dinb(n10926), .dout(n10928));
  jxor g10736(.dina(n10928), .dinb(n10925), .dout(n10929));
  jxor g10737(.dina(n10929), .dinb(n10912), .dout(n10930));
  jand g10738(.dina(n10634), .dinb(n10610), .dout(n10931));
  jand g10739(.dina(n10635), .dinb(n10607), .dout(n10932));
  jor  g10740(.dina(n10932), .dinb(n10931), .dout(n10933));
  jand g10741(.dina(n10736), .dinb(n10712), .dout(n10934));
  jand g10742(.dina(n10760), .dinb(n10737), .dout(n10935));
  jor  g10743(.dina(n10935), .dinb(n10934), .dout(n10936));
  jxor g10744(.dina(n10936), .dinb(n10933), .dout(n10937));
  jxor g10745(.dina(n10937), .dinb(n10930), .dout(n10938));
  jxor g10746(.dina(n10938), .dinb(n10892), .dout(n10939));
  jxor g10747(.dina(n10939), .dinb(n10844), .dout(n10940));
  jxor g10748(.dina(n10940), .dinb(n10773), .dout(n10941));
  jand g10749(.dina(n10764), .dinb(n10593), .dout(n10942));
  jor  g10750(.dina(n10764), .dinb(n10593), .dout(n10943));
  jand g10751(.dina(n10769), .dinb(n10943), .dout(n10944));
  jor  g10752(.dina(n10944), .dinb(n10942), .dout(n10945));
  jxor g10753(.dina(n10945), .dinb(n10941), .dout(\asquared[79] ));
  jand g10754(.dina(n10843), .dinb(n10840), .dout(n10947));
  jand g10755(.dina(n10939), .dinb(n10844), .dout(n10948));
  jor  g10756(.dina(n10948), .dinb(n10947), .dout(n10949));
  jand g10757(.dina(n10936), .dinb(n10933), .dout(n10950));
  jand g10758(.dina(n10937), .dinb(n10930), .dout(n10951));
  jor  g10759(.dina(n10951), .dinb(n10950), .dout(n10952));
  jand g10760(.dina(n10836), .dinb(n10808), .dout(n10953));
  jand g10761(.dina(n10837), .dinb(n10782), .dout(n10954));
  jor  g10762(.dina(n10954), .dinb(n10953), .dout(n10955));
  jand g10763(.dina(n10805), .dinb(n10648), .dout(n10956));
  jor  g10764(.dina(n10956), .dinb(n10803), .dout(n10957));
  jand g10765(.dina(n10794), .dinb(n10792), .dout(n10958));
  jor  g10766(.dina(n10958), .dinb(n10797), .dout(n10959));
  jxor g10767(.dina(n10959), .dinb(n10957), .dout(n10960));
  jand g10768(.dina(n10811), .dinb(n10809), .dout(n10961));
  jor  g10769(.dina(n10961), .dinb(n10814), .dout(n10962));
  jxor g10770(.dina(n10962), .dinb(n10960), .dout(n10963));
  jnot g10771(.din(n10963), .dout(n10964));
  jor  g10772(.dina(n10910), .dinb(n10905), .dout(n10965));
  jand g10773(.dina(n10911), .dinb(n10895), .dout(n10966));
  jnot g10774(.din(n10966), .dout(n10967));
  jand g10775(.dina(n10967), .dinb(n10965), .dout(n10968));
  jxor g10776(.dina(n10968), .dinb(n10964), .dout(n10969));
  jand g10777(.dina(n10921), .dinb(n10914), .dout(n10970));
  jand g10778(.dina(n10924), .dinb(n10922), .dout(n10971));
  jor  g10779(.dina(n10971), .dinb(n10970), .dout(n10972));
  jand g10780(.dina(\a[56] ), .dinb(\a[23] ), .dout(n10973));
  jnot g10781(.din(n10973), .dout(n10974));
  jand g10782(.dina(\a[52] ), .dinb(\a[27] ), .dout(n10975));
  jnot g10783(.din(n10975), .dout(n10976));
  jand g10784(.dina(n10976), .dinb(n10974), .dout(n10977));
  jand g10785(.dina(\a[56] ), .dinb(\a[27] ), .dout(n10978));
  jand g10786(.dina(n10978), .dinb(n10289), .dout(n10979));
  jor  g10787(.dina(n10979), .dinb(n10977), .dout(n10980));
  jxor g10788(.dina(n10980), .dinb(n10900), .dout(n10981));
  jnot g10789(.din(n10981), .dout(n10982));
  jand g10790(.dina(\a[63] ), .dinb(\a[16] ), .dout(n10983));
  jand g10791(.dina(\a[44] ), .dinb(\a[35] ), .dout(n10984));
  jor  g10792(.dina(n10984), .dinb(n10830), .dout(n10985));
  jand g10793(.dina(\a[45] ), .dinb(\a[35] ), .dout(n10986));
  jand g10794(.dina(n10986), .dinb(n10828), .dout(n10987));
  jnot g10795(.din(n10987), .dout(n10988));
  jand g10796(.dina(n10988), .dinb(n10985), .dout(n10989));
  jxor g10797(.dina(n10989), .dinb(n10983), .dout(n10990));
  jxor g10798(.dina(n10990), .dinb(n10982), .dout(n10991));
  jxor g10799(.dina(n10991), .dinb(n10972), .dout(n10992));
  jxor g10800(.dina(n10992), .dinb(n10969), .dout(n10993));
  jxor g10801(.dina(n10993), .dinb(n10955), .dout(n10994));
  jand g10802(.dina(n10903), .dinb(n10896), .dout(n10995));
  jor  g10803(.dina(n10995), .dinb(n10901), .dout(n10996));
  jand g10804(.dina(\a[61] ), .dinb(\a[18] ), .dout(n10997));
  jnot g10805(.din(n10908), .dout(n10998));
  jand g10806(.dina(n10998), .dinb(n10907), .dout(n10999));
  jnot g10807(.din(n10999), .dout(n11000));
  jand g10808(.dina(n10908), .dinb(n10906), .dout(n11001));
  jor  g10809(.dina(n11001), .dinb(n10717), .dout(n11002));
  jand g10810(.dina(n11002), .dinb(n11000), .dout(n11003));
  jxor g10811(.dina(n11003), .dinb(n10997), .dout(n11004));
  jxor g10812(.dina(n11004), .dinb(n10996), .dout(n11005));
  jand g10813(.dina(n10833), .dinb(n10827), .dout(n11006));
  jor  g10814(.dina(n11006), .dinb(n10831), .dout(n11007));
  jand g10815(.dina(n10825), .dinb(n10818), .dout(n11008));
  jor  g10816(.dina(n11008), .dinb(n10823), .dout(n11009));
  jand g10817(.dina(n10786), .dinb(n10783), .dout(n11010));
  jor  g10818(.dina(n11010), .dinb(n10789), .dout(n11011));
  jxor g10819(.dina(n11011), .dinb(n11009), .dout(n11012));
  jxor g10820(.dina(n11012), .dinb(n11007), .dout(n11013));
  jxor g10821(.dina(n11013), .dinb(n11005), .dout(n11014));
  jor  g10822(.dina(n10834), .dinb(n10826), .dout(n11015));
  jand g10823(.dina(n10834), .dinb(n10826), .dout(n11016));
  jor  g10824(.dina(n11016), .dinb(n10817), .dout(n11017));
  jand g10825(.dina(n11017), .dinb(n11015), .dout(n11018));
  jxor g10826(.dina(n11018), .dinb(n11014), .dout(n11019));
  jxor g10827(.dina(n11019), .dinb(n10994), .dout(n11020));
  jxor g10828(.dina(n11020), .dinb(n10952), .dout(n11021));
  jand g10829(.dina(n10838), .dinb(n10779), .dout(n11022));
  jand g10830(.dina(n10839), .dinb(n10776), .dout(n11023));
  jor  g10831(.dina(n11023), .dinb(n11022), .dout(n11024));
  jxor g10832(.dina(n11024), .dinb(n11021), .dout(n11025));
  jand g10833(.dina(n10866), .dinb(n10863), .dout(n11026));
  jand g10834(.dina(n10890), .dinb(n10867), .dout(n11027));
  jor  g10835(.dina(n11027), .dinb(n11026), .dout(n11028));
  jand g10836(.dina(n10888), .dinb(n10885), .dout(n11029));
  jand g10837(.dina(n10889), .dinb(n10877), .dout(n11030));
  jor  g10838(.dina(n11030), .dinb(n11029), .dout(n11031));
  jand g10839(.dina(\a[42] ), .dinb(\a[37] ), .dout(n11032));
  jand g10840(.dina(\a[40] ), .dinb(\a[39] ), .dout(n11033));
  jand g10841(.dina(\a[41] ), .dinb(\a[38] ), .dout(n11034));
  jor  g10842(.dina(n11034), .dinb(n11033), .dout(n11035));
  jnot g10843(.din(n11035), .dout(n11036));
  jand g10844(.dina(\a[41] ), .dinb(\a[39] ), .dout(n11037));
  jand g10845(.dina(n11037), .dinb(n10906), .dout(n11038));
  jor  g10846(.dina(n11038), .dinb(n11036), .dout(n11039));
  jxor g10847(.dina(n11039), .dinb(n11032), .dout(n11040));
  jnot g10848(.din(n11040), .dout(n11041));
  jand g10849(.dina(\a[55] ), .dinb(\a[24] ), .dout(n11042));
  jand g10850(.dina(\a[53] ), .dinb(\a[26] ), .dout(n11043));
  jand g10851(.dina(\a[54] ), .dinb(\a[25] ), .dout(n11044));
  jor  g10852(.dina(n11044), .dinb(n11043), .dout(n11045));
  jand g10853(.dina(\a[54] ), .dinb(\a[26] ), .dout(n11046));
  jand g10854(.dina(n11046), .dinb(n10809), .dout(n11047));
  jnot g10855(.din(n11047), .dout(n11048));
  jand g10856(.dina(n11048), .dinb(n11045), .dout(n11049));
  jxor g10857(.dina(n11049), .dinb(n11042), .dout(n11050));
  jxor g10858(.dina(n11050), .dinb(n11041), .dout(n11051));
  jand g10859(.dina(\a[51] ), .dinb(\a[28] ), .dout(n11052));
  jor  g10860(.dina(n10788), .dinb(\a[40] ), .dout(n11053));
  jnot g10861(.din(n11053), .dout(n11054));
  jand g10862(.dina(\a[62] ), .dinb(\a[40] ), .dout(n11055));
  jand g10863(.dina(n11055), .dinb(\a[17] ), .dout(n11056));
  jor  g10864(.dina(n11056), .dinb(n11054), .dout(n11057));
  jxor g10865(.dina(n11057), .dinb(n11052), .dout(n11058));
  jnot g10866(.din(n11058), .dout(n11059));
  jxor g10867(.dina(n11059), .dinb(n11051), .dout(n11060));
  jand g10868(.dina(\a[46] ), .dinb(\a[33] ), .dout(n11061));
  jand g10869(.dina(\a[47] ), .dinb(\a[32] ), .dout(n11062));
  jor  g10870(.dina(n11062), .dinb(n11061), .dout(n11063));
  jnot g10871(.din(n11063), .dout(n11064));
  jand g10872(.dina(\a[47] ), .dinb(\a[33] ), .dout(n11065));
  jand g10873(.dina(n11065), .dinb(n10827), .dout(n11066));
  jor  g10874(.dina(n11066), .dinb(n11064), .dout(n11067));
  jxor g10875(.dina(n11067), .dinb(n10822), .dout(n11068));
  jand g10876(.dina(\a[57] ), .dinb(\a[22] ), .dout(n11069));
  jand g10877(.dina(\a[49] ), .dinb(\a[30] ), .dout(n11070));
  jor  g10878(.dina(n11070), .dinb(n10796), .dout(n11071));
  jnot g10879(.din(n11071), .dout(n11072));
  jand g10880(.dina(\a[50] ), .dinb(\a[30] ), .dout(n11073));
  jand g10881(.dina(n11073), .dinb(n10742), .dout(n11074));
  jor  g10882(.dina(n11074), .dinb(n11072), .dout(n11075));
  jxor g10883(.dina(n11075), .dinb(n11069), .dout(n11076));
  jand g10884(.dina(\a[60] ), .dinb(\a[19] ), .dout(n11077));
  jand g10885(.dina(\a[59] ), .dinb(\a[20] ), .dout(n11078));
  jand g10886(.dina(\a[58] ), .dinb(\a[21] ), .dout(n11079));
  jor  g10887(.dina(n11079), .dinb(n11078), .dout(n11080));
  jand g10888(.dina(n10818), .dinb(n10802), .dout(n11081));
  jnot g10889(.din(n11081), .dout(n11082));
  jand g10890(.dina(n11082), .dinb(n11080), .dout(n11083));
  jxor g10891(.dina(n11083), .dinb(n11077), .dout(n11084));
  jxor g10892(.dina(n11084), .dinb(n11076), .dout(n11085));
  jxor g10893(.dina(n11085), .dinb(n11068), .dout(n11086));
  jxor g10894(.dina(n11086), .dinb(n11060), .dout(n11087));
  jxor g10895(.dina(n11087), .dinb(n11031), .dout(n11088));
  jxor g10896(.dina(n11088), .dinb(n11028), .dout(n11089));
  jand g10897(.dina(n10881), .dinb(n10879), .dout(n11090));
  jand g10898(.dina(n10884), .dinb(n10882), .dout(n11091));
  jor  g10899(.dina(n11091), .dinb(n11090), .dout(n11092));
  jand g10900(.dina(n10873), .dinb(n10871), .dout(n11093));
  jand g10901(.dina(n10876), .dinb(n10874), .dout(n11094));
  jor  g10902(.dina(n11094), .dinb(n11093), .dout(n11095));
  jxor g10903(.dina(n11095), .dinb(n11092), .dout(n11096));
  jnot g10904(.din(n10799), .dout(n11097));
  jor  g10905(.dina(n10806), .dinb(n11097), .dout(n11098));
  jnot g10906(.din(n10791), .dout(n11099));
  jand g10907(.dina(n10806), .dinb(n11097), .dout(n11100));
  jor  g10908(.dina(n11100), .dinb(n11099), .dout(n11101));
  jand g10909(.dina(n11101), .dinb(n11098), .dout(n11102));
  jxor g10910(.dina(n11102), .dinb(n11096), .dout(n11103));
  jnot g10911(.din(n11103), .dout(n11104));
  jand g10912(.dina(n10854), .dinb(n10850), .dout(n11105));
  jnot g10913(.din(n11105), .dout(n11106));
  jor  g10914(.dina(n10862), .dinb(n10856), .dout(n11107));
  jand g10915(.dina(n11107), .dinb(n11106), .dout(n11108));
  jxor g10916(.dina(n11108), .dinb(n11104), .dout(n11109));
  jand g10917(.dina(n10928), .dinb(n10925), .dout(n11110));
  jand g10918(.dina(n10929), .dinb(n10912), .dout(n11111));
  jor  g10919(.dina(n11111), .dinb(n11110), .dout(n11112));
  jxor g10920(.dina(n11112), .dinb(n11109), .dout(n11113));
  jxor g10921(.dina(n11113), .dinb(n11089), .dout(n11114));
  jand g10922(.dina(n10891), .dinb(n10847), .dout(n11115));
  jand g10923(.dina(n10938), .dinb(n10892), .dout(n11116));
  jor  g10924(.dina(n11116), .dinb(n11115), .dout(n11117));
  jxor g10925(.dina(n11117), .dinb(n11114), .dout(n11118));
  jxor g10926(.dina(n11118), .dinb(n11025), .dout(n11119));
  jxor g10927(.dina(n11119), .dinb(n10949), .dout(n11120));
  jand g10928(.dina(n10940), .dinb(n10773), .dout(n11121));
  jor  g10929(.dina(n10940), .dinb(n10773), .dout(n11122));
  jand g10930(.dina(n10945), .dinb(n11122), .dout(n11123));
  jor  g10931(.dina(n11123), .dinb(n11121), .dout(n11124));
  jxor g10932(.dina(n11124), .dinb(n11120), .dout(\asquared[80] ));
  jand g10933(.dina(n11117), .dinb(n11114), .dout(n11126));
  jand g10934(.dina(n11118), .dinb(n11025), .dout(n11127));
  jor  g10935(.dina(n11127), .dinb(n11126), .dout(n11128));
  jand g10936(.dina(n11020), .dinb(n10952), .dout(n11129));
  jand g10937(.dina(n11024), .dinb(n11021), .dout(n11130));
  jor  g10938(.dina(n11130), .dinb(n11129), .dout(n11131));
  jand g10939(.dina(n10993), .dinb(n10955), .dout(n11132));
  jand g10940(.dina(n11019), .dinb(n10994), .dout(n11133));
  jor  g10941(.dina(n11133), .dinb(n11132), .dout(n11134));
  jor  g10942(.dina(n11108), .dinb(n11104), .dout(n11135));
  jand g10943(.dina(n11112), .dinb(n11109), .dout(n11136));
  jnot g10944(.din(n11136), .dout(n11137));
  jand g10945(.dina(n11137), .dinb(n11135), .dout(n11138));
  jnot g10946(.din(n11138), .dout(n11139));
  jand g10947(.dina(\a[61] ), .dinb(\a[19] ), .dout(n11140));
  jand g10948(.dina(\a[62] ), .dinb(\a[18] ), .dout(n11141));
  jor  g10949(.dina(n11141), .dinb(n11140), .dout(n11142));
  jand g10950(.dina(\a[62] ), .dinb(\a[19] ), .dout(n11143));
  jand g10951(.dina(n11143), .dinb(n10997), .dout(n11144));
  jnot g10952(.din(n11144), .dout(n11145));
  jand g10953(.dina(n11145), .dinb(n11142), .dout(n11146));
  jand g10954(.dina(n11053), .dinb(n11052), .dout(n11147));
  jor  g10955(.dina(n11147), .dinb(n11056), .dout(n11148));
  jxor g10956(.dina(n11148), .dinb(n11146), .dout(n11149));
  jand g10957(.dina(\a[46] ), .dinb(\a[34] ), .dout(n11150));
  jand g10958(.dina(\a[44] ), .dinb(\a[36] ), .dout(n11151));
  jor  g10959(.dina(n11151), .dinb(n10986), .dout(n11152));
  jnot g10960(.din(n11152), .dout(n11153));
  jand g10961(.dina(\a[45] ), .dinb(\a[36] ), .dout(n11154));
  jand g10962(.dina(n11154), .dinb(n10984), .dout(n11155));
  jor  g10963(.dina(n11155), .dinb(n11153), .dout(n11156));
  jxor g10964(.dina(n11156), .dinb(n11150), .dout(n11157));
  jnot g10965(.din(n11157), .dout(n11158));
  jand g10966(.dina(\a[63] ), .dinb(\a[17] ), .dout(n11159));
  jand g10967(.dina(\a[51] ), .dinb(\a[29] ), .dout(n11160));
  jor  g10968(.dina(n11160), .dinb(n11159), .dout(n11161));
  jand g10969(.dina(\a[63] ), .dinb(\a[29] ), .dout(n11162));
  jand g10970(.dina(n11162), .dinb(n6356), .dout(n11163));
  jnot g10971(.din(n11163), .dout(n11164));
  jand g10972(.dina(n11164), .dinb(n11161), .dout(n11165));
  jxor g10973(.dina(n11165), .dinb(n11065), .dout(n11166));
  jxor g10974(.dina(n11166), .dinb(n11158), .dout(n11167));
  jxor g10975(.dina(n11167), .dinb(n11149), .dout(n11168));
  jand g10976(.dina(\a[58] ), .dinb(\a[22] ), .dout(n11169));
  jor  g10977(.dina(n11169), .dinb(n10802), .dout(n11170));
  jand g10978(.dina(\a[59] ), .dinb(\a[22] ), .dout(n11171));
  jand g10979(.dina(n11171), .dinb(n11079), .dout(n11172));
  jnot g10980(.din(n11172), .dout(n11173));
  jand g10981(.dina(n11173), .dinb(n11170), .dout(n11174));
  jand g10982(.dina(\a[60] ), .dinb(\a[20] ), .dout(n11175));
  jxor g10983(.dina(n11175), .dinb(n11174), .dout(n11176));
  jand g10984(.dina(n11035), .dinb(n11032), .dout(n11177));
  jor  g10985(.dina(n11177), .dinb(n11038), .dout(n11178));
  jxor g10986(.dina(n11178), .dinb(n11176), .dout(n11179));
  jnot g10987(.din(n11179), .dout(n11180));
  jand g10988(.dina(\a[49] ), .dinb(\a[31] ), .dout(n11181));
  jand g10989(.dina(\a[48] ), .dinb(\a[32] ), .dout(n11182));
  jor  g10990(.dina(n11182), .dinb(n11181), .dout(n11183));
  jnot g10991(.din(n11183), .dout(n11184));
  jand g10992(.dina(\a[49] ), .dinb(\a[32] ), .dout(n11185));
  jand g10993(.dina(n11185), .dinb(n10822), .dout(n11186));
  jor  g10994(.dina(n11186), .dinb(n11184), .dout(n11187));
  jxor g10995(.dina(n11187), .dinb(n11073), .dout(n11188));
  jxor g10996(.dina(n11188), .dinb(n11180), .dout(n11189));
  jand g10997(.dina(\a[53] ), .dinb(\a[27] ), .dout(n11190));
  jand g10998(.dina(\a[52] ), .dinb(\a[28] ), .dout(n11191));
  jor  g10999(.dina(n11191), .dinb(n11190), .dout(n11192));
  jnot g11000(.din(n11192), .dout(n11193));
  jand g11001(.dina(\a[53] ), .dinb(\a[28] ), .dout(n11194));
  jand g11002(.dina(n11194), .dinb(n10975), .dout(n11195));
  jor  g11003(.dina(n11195), .dinb(n11193), .dout(n11196));
  jxor g11004(.dina(n11196), .dinb(n11037), .dout(n11197));
  jand g11005(.dina(\a[55] ), .dinb(\a[25] ), .dout(n11198));
  jand g11006(.dina(\a[43] ), .dinb(\a[37] ), .dout(n11199));
  jand g11007(.dina(\a[42] ), .dinb(\a[38] ), .dout(n11200));
  jor  g11008(.dina(n11200), .dinb(n11199), .dout(n11201));
  jnot g11009(.din(n11201), .dout(n11202));
  jand g11010(.dina(\a[43] ), .dinb(\a[38] ), .dout(n11203));
  jand g11011(.dina(n11203), .dinb(n11032), .dout(n11204));
  jor  g11012(.dina(n11204), .dinb(n11202), .dout(n11205));
  jxor g11013(.dina(n11205), .dinb(n11198), .dout(n11206));
  jand g11014(.dina(\a[57] ), .dinb(\a[23] ), .dout(n11207));
  jor  g11015(.dina(n11046), .dinb(n10813), .dout(n11208));
  jand g11016(.dina(\a[56] ), .dinb(\a[26] ), .dout(n11209));
  jand g11017(.dina(n11209), .dinb(n9911), .dout(n11210));
  jnot g11018(.din(n11210), .dout(n11211));
  jand g11019(.dina(n11211), .dinb(n11208), .dout(n11212));
  jxor g11020(.dina(n11212), .dinb(n11207), .dout(n11213));
  jxor g11021(.dina(n11213), .dinb(n11206), .dout(n11214));
  jxor g11022(.dina(n11214), .dinb(n11197), .dout(n11215));
  jxor g11023(.dina(n11215), .dinb(n11189), .dout(n11216));
  jxor g11024(.dina(n11216), .dinb(n11168), .dout(n11217));
  jxor g11025(.dina(n11217), .dinb(n11139), .dout(n11218));
  jxor g11026(.dina(n11218), .dinb(n11134), .dout(n11219));
  jxor g11027(.dina(n11219), .dinb(n11131), .dout(n11220));
  jand g11028(.dina(n11088), .dinb(n11028), .dout(n11221));
  jand g11029(.dina(n11113), .dinb(n11089), .dout(n11222));
  jor  g11030(.dina(n11222), .dinb(n11221), .dout(n11223));
  jand g11031(.dina(n11086), .dinb(n11060), .dout(n11224));
  jand g11032(.dina(n11087), .dinb(n11031), .dout(n11225));
  jor  g11033(.dina(n11225), .dinb(n11224), .dout(n11226));
  jand g11034(.dina(n10989), .dinb(n10983), .dout(n11227));
  jor  g11035(.dina(n11227), .dinb(n10987), .dout(n11228));
  jand g11036(.dina(n11049), .dinb(n11042), .dout(n11229));
  jor  g11037(.dina(n11229), .dinb(n11047), .dout(n11230));
  jxor g11038(.dina(n11230), .dinb(n11228), .dout(n11231));
  jnot g11039(.din(n10977), .dout(n11232));
  jand g11040(.dina(n11232), .dinb(n10900), .dout(n11233));
  jor  g11041(.dina(n11233), .dinb(n10979), .dout(n11234));
  jxor g11042(.dina(n11234), .dinb(n11231), .dout(n11235));
  jand g11043(.dina(n10990), .dinb(n10982), .dout(n11236));
  jand g11044(.dina(n10991), .dinb(n10972), .dout(n11237));
  jor  g11045(.dina(n11237), .dinb(n11236), .dout(n11238));
  jxor g11046(.dina(n11238), .dinb(n11235), .dout(n11239));
  jand g11047(.dina(n11095), .dinb(n11092), .dout(n11240));
  jand g11048(.dina(n11102), .dinb(n11096), .dout(n11241));
  jor  g11049(.dina(n11241), .dinb(n11240), .dout(n11242));
  jxor g11050(.dina(n11242), .dinb(n11239), .dout(n11243));
  jxor g11051(.dina(n11243), .dinb(n11226), .dout(n11244));
  jand g11052(.dina(n11083), .dinb(n11077), .dout(n11245));
  jor  g11053(.dina(n11245), .dinb(n11081), .dout(n11246));
  jand g11054(.dina(n11071), .dinb(n11069), .dout(n11247));
  jor  g11055(.dina(n11247), .dinb(n11074), .dout(n11248));
  jxor g11056(.dina(n11248), .dinb(n11246), .dout(n11249));
  jand g11057(.dina(n11063), .dinb(n10822), .dout(n11250));
  jor  g11058(.dina(n11250), .dinb(n11066), .dout(n11251));
  jxor g11059(.dina(n11251), .dinb(n11249), .dout(n11252));
  jor  g11060(.dina(n11050), .dinb(n11041), .dout(n11253));
  jand g11061(.dina(n11050), .dinb(n11041), .dout(n11254));
  jor  g11062(.dina(n11059), .dinb(n11254), .dout(n11255));
  jand g11063(.dina(n11255), .dinb(n11253), .dout(n11256));
  jnot g11064(.din(n11076), .dout(n11257));
  jor  g11065(.dina(n11084), .dinb(n11257), .dout(n11258));
  jnot g11066(.din(n11068), .dout(n11259));
  jand g11067(.dina(n11084), .dinb(n11257), .dout(n11260));
  jor  g11068(.dina(n11260), .dinb(n11259), .dout(n11261));
  jand g11069(.dina(n11261), .dinb(n11258), .dout(n11262));
  jxor g11070(.dina(n11262), .dinb(n11256), .dout(n11263));
  jxor g11071(.dina(n11263), .dinb(n11252), .dout(n11264));
  jxor g11072(.dina(n11264), .dinb(n11244), .dout(n11265));
  jand g11073(.dina(n10959), .dinb(n10957), .dout(n11266));
  jand g11074(.dina(n10962), .dinb(n10960), .dout(n11267));
  jor  g11075(.dina(n11267), .dinb(n11266), .dout(n11268));
  jand g11076(.dina(n11011), .dinb(n11009), .dout(n11269));
  jand g11077(.dina(n11012), .dinb(n11007), .dout(n11270));
  jor  g11078(.dina(n11270), .dinb(n11269), .dout(n11271));
  jxor g11079(.dina(n11271), .dinb(n11268), .dout(n11272));
  jand g11080(.dina(n11003), .dinb(n10997), .dout(n11273));
  jand g11081(.dina(n11004), .dinb(n10996), .dout(n11274));
  jor  g11082(.dina(n11274), .dinb(n11273), .dout(n11275));
  jxor g11083(.dina(n11275), .dinb(n11272), .dout(n11276));
  jor  g11084(.dina(n10968), .dinb(n10964), .dout(n11277));
  jand g11085(.dina(n10992), .dinb(n10969), .dout(n11278));
  jnot g11086(.din(n11278), .dout(n11279));
  jand g11087(.dina(n11279), .dinb(n11277), .dout(n11280));
  jnot g11088(.din(n11280), .dout(n11281));
  jand g11089(.dina(n11013), .dinb(n11005), .dout(n11282));
  jand g11090(.dina(n11018), .dinb(n11014), .dout(n11283));
  jor  g11091(.dina(n11283), .dinb(n11282), .dout(n11284));
  jxor g11092(.dina(n11284), .dinb(n11281), .dout(n11285));
  jxor g11093(.dina(n11285), .dinb(n11276), .dout(n11286));
  jxor g11094(.dina(n11286), .dinb(n11265), .dout(n11287));
  jxor g11095(.dina(n11287), .dinb(n11223), .dout(n11288));
  jxor g11096(.dina(n11288), .dinb(n11220), .dout(n11289));
  jxor g11097(.dina(n11289), .dinb(n11128), .dout(n11290));
  jand g11098(.dina(n11119), .dinb(n10949), .dout(n11291));
  jor  g11099(.dina(n11119), .dinb(n10949), .dout(n11292));
  jand g11100(.dina(n11124), .dinb(n11292), .dout(n11293));
  jor  g11101(.dina(n11293), .dinb(n11291), .dout(n11294));
  jxor g11102(.dina(n11294), .dinb(n11290), .dout(\asquared[81] ));
  jand g11103(.dina(n11219), .dinb(n11131), .dout(n11296));
  jand g11104(.dina(n11288), .dinb(n11220), .dout(n11297));
  jor  g11105(.dina(n11297), .dinb(n11296), .dout(n11298));
  jand g11106(.dina(n11286), .dinb(n11265), .dout(n11299));
  jand g11107(.dina(n11287), .dinb(n11223), .dout(n11300));
  jor  g11108(.dina(n11300), .dinb(n11299), .dout(n11301));
  jand g11109(.dina(n11243), .dinb(n11226), .dout(n11302));
  jand g11110(.dina(n11264), .dinb(n11244), .dout(n11303));
  jor  g11111(.dina(n11303), .dinb(n11302), .dout(n11304));
  jand g11112(.dina(n11284), .dinb(n11281), .dout(n11305));
  jand g11113(.dina(n11285), .dinb(n11276), .dout(n11306));
  jor  g11114(.dina(n11306), .dinb(n11305), .dout(n11307));
  jand g11115(.dina(n11271), .dinb(n11268), .dout(n11308));
  jand g11116(.dina(n11275), .dinb(n11272), .dout(n11309));
  jor  g11117(.dina(n11309), .dinb(n11308), .dout(n11310));
  jnot g11118(.din(n8326), .dout(n11311));
  jand g11119(.dina(\a[48] ), .dinb(\a[33] ), .dout(n11312));
  jand g11120(.dina(\a[47] ), .dinb(\a[34] ), .dout(n11313));
  jor  g11121(.dina(n11313), .dinb(n11312), .dout(n11314));
  jand g11122(.dina(\a[48] ), .dinb(\a[34] ), .dout(n11315));
  jand g11123(.dina(n11315), .dinb(n11065), .dout(n11316));
  jnot g11124(.din(n11316), .dout(n11317));
  jand g11125(.dina(n11317), .dinb(n11314), .dout(n11318));
  jxor g11126(.dina(n11318), .dinb(n11311), .dout(n11319));
  jnot g11127(.din(n11171), .dout(n11320));
  jand g11128(.dina(\a[58] ), .dinb(\a[23] ), .dout(n11321));
  jor  g11129(.dina(n11321), .dinb(n10152), .dout(n11322));
  jand g11130(.dina(\a[58] ), .dinb(\a[25] ), .dout(n11323));
  jand g11131(.dina(n11323), .dinb(n10973), .dout(n11324));
  jnot g11132(.din(n11324), .dout(n11325));
  jand g11133(.dina(n11325), .dinb(n11322), .dout(n11326));
  jxor g11134(.dina(n11326), .dinb(n11320), .dout(n11327));
  jnot g11135(.din(n11143), .dout(n11328));
  jnot g11136(.din(\a[40] ), .dout(n11329));
  jand g11137(.dina(\a[41] ), .dinb(n11329), .dout(n11330));
  jxor g11138(.dina(n11330), .dinb(n11328), .dout(n11331));
  jnot g11139(.din(n11331), .dout(n11332));
  jxor g11140(.dina(n11332), .dinb(n11327), .dout(n11333));
  jxor g11141(.dina(n11333), .dinb(n11319), .dout(n11334));
  jxor g11142(.dina(n11334), .dinb(n11310), .dout(n11335));
  jand g11143(.dina(\a[46] ), .dinb(\a[35] ), .dout(n11336));
  jand g11144(.dina(\a[44] ), .dinb(\a[37] ), .dout(n11337));
  jor  g11145(.dina(n11337), .dinb(n11154), .dout(n11338));
  jnot g11146(.din(n11338), .dout(n11339));
  jand g11147(.dina(\a[45] ), .dinb(\a[37] ), .dout(n11340));
  jand g11148(.dina(n11340), .dinb(n11151), .dout(n11341));
  jor  g11149(.dina(n11341), .dinb(n11339), .dout(n11342));
  jxor g11150(.dina(n11342), .dinb(n11336), .dout(n11343));
  jnot g11151(.din(n11343), .dout(n11344));
  jand g11152(.dina(\a[63] ), .dinb(\a[18] ), .dout(n11345));
  jand g11153(.dina(\a[61] ), .dinb(\a[20] ), .dout(n11346));
  jand g11154(.dina(\a[60] ), .dinb(\a[21] ), .dout(n11347));
  jor  g11155(.dina(n11347), .dinb(n11346), .dout(n11348));
  jand g11156(.dina(\a[61] ), .dinb(\a[21] ), .dout(n11349));
  jand g11157(.dina(n11349), .dinb(n11175), .dout(n11350));
  jnot g11158(.din(n11350), .dout(n11351));
  jand g11159(.dina(n11351), .dinb(n11348), .dout(n11352));
  jxor g11160(.dina(n11352), .dinb(n11345), .dout(n11353));
  jxor g11161(.dina(n11353), .dinb(n11344), .dout(n11354));
  jnot g11162(.din(n11354), .dout(n11355));
  jand g11163(.dina(\a[55] ), .dinb(\a[26] ), .dout(n11356));
  jnot g11164(.din(n11194), .dout(n11357));
  jand g11165(.dina(\a[52] ), .dinb(\a[29] ), .dout(n11358));
  jnot g11166(.din(n11358), .dout(n11359));
  jand g11167(.dina(n11359), .dinb(n11357), .dout(n11360));
  jand g11168(.dina(\a[53] ), .dinb(\a[29] ), .dout(n11361));
  jand g11169(.dina(n11361), .dinb(n11191), .dout(n11362));
  jor  g11170(.dina(n11362), .dinb(n11360), .dout(n11363));
  jxor g11171(.dina(n11363), .dinb(n11356), .dout(n11364));
  jxor g11172(.dina(n11364), .dinb(n11355), .dout(n11365));
  jxor g11173(.dina(n11365), .dinb(n11335), .dout(n11366));
  jxor g11174(.dina(n11366), .dinb(n11307), .dout(n11367));
  jxor g11175(.dina(n11367), .dinb(n11304), .dout(n11368));
  jxor g11176(.dina(n11368), .dinb(n11301), .dout(n11369));
  jand g11177(.dina(n11215), .dinb(n11189), .dout(n11370));
  jand g11178(.dina(n11216), .dinb(n11168), .dout(n11371));
  jor  g11179(.dina(n11371), .dinb(n11370), .dout(n11372));
  jand g11180(.dina(n11165), .dinb(n11065), .dout(n11373));
  jor  g11181(.dina(n11373), .dinb(n11163), .dout(n11374));
  jand g11182(.dina(n11183), .dinb(n11073), .dout(n11375));
  jor  g11183(.dina(n11375), .dinb(n11186), .dout(n11376));
  jxor g11184(.dina(n11376), .dinb(n11374), .dout(n11377));
  jand g11185(.dina(n11175), .dinb(n11174), .dout(n11378));
  jor  g11186(.dina(n11378), .dinb(n11172), .dout(n11379));
  jxor g11187(.dina(n11379), .dinb(n11377), .dout(n11380));
  jand g11188(.dina(n11166), .dinb(n11158), .dout(n11381));
  jand g11189(.dina(n11167), .dinb(n11149), .dout(n11382));
  jor  g11190(.dina(n11382), .dinb(n11381), .dout(n11383));
  jxor g11191(.dina(n11383), .dinb(n11380), .dout(n11384));
  jand g11192(.dina(n11148), .dinb(n11146), .dout(n11385));
  jor  g11193(.dina(n11385), .dinb(n11144), .dout(n11386));
  jand g11194(.dina(n11152), .dinb(n11150), .dout(n11387));
  jor  g11195(.dina(n11387), .dinb(n11155), .dout(n11388));
  jxor g11196(.dina(n11388), .dinb(n11386), .dout(n11389));
  jand g11197(.dina(\a[51] ), .dinb(\a[30] ), .dout(n11390));
  jand g11198(.dina(\a[50] ), .dinb(\a[31] ), .dout(n11391));
  jor  g11199(.dina(n11391), .dinb(n11185), .dout(n11392));
  jnot g11200(.din(n11392), .dout(n11393));
  jand g11201(.dina(\a[50] ), .dinb(\a[32] ), .dout(n11394));
  jand g11202(.dina(n11394), .dinb(n11181), .dout(n11395));
  jor  g11203(.dina(n11395), .dinb(n11393), .dout(n11396));
  jxor g11204(.dina(n11396), .dinb(n11390), .dout(n11397));
  jnot g11205(.din(n11397), .dout(n11398));
  jxor g11206(.dina(n11398), .dinb(n11389), .dout(n11399));
  jxor g11207(.dina(n11399), .dinb(n11384), .dout(n11400));
  jxor g11208(.dina(n11400), .dinb(n11372), .dout(n11401));
  jand g11209(.dina(n11212), .dinb(n11207), .dout(n11402));
  jor  g11210(.dina(n11402), .dinb(n11210), .dout(n11403));
  jand g11211(.dina(n11201), .dinb(n11198), .dout(n11404));
  jor  g11212(.dina(n11404), .dinb(n11204), .dout(n11405));
  jand g11213(.dina(n11192), .dinb(n11037), .dout(n11406));
  jor  g11214(.dina(n11406), .dinb(n11195), .dout(n11407));
  jxor g11215(.dina(n11407), .dinb(n11405), .dout(n11408));
  jxor g11216(.dina(n11408), .dinb(n11403), .dout(n11409));
  jand g11217(.dina(n11178), .dinb(n11176), .dout(n11410));
  jnot g11218(.din(n11410), .dout(n11411));
  jor  g11219(.dina(n11188), .dinb(n11180), .dout(n11412));
  jand g11220(.dina(n11412), .dinb(n11411), .dout(n11413));
  jnot g11221(.din(n11413), .dout(n11414));
  jnot g11222(.din(n11206), .dout(n11415));
  jor  g11223(.dina(n11213), .dinb(n11415), .dout(n11416));
  jnot g11224(.din(n11197), .dout(n11417));
  jand g11225(.dina(n11213), .dinb(n11415), .dout(n11418));
  jor  g11226(.dina(n11418), .dinb(n11417), .dout(n11419));
  jand g11227(.dina(n11419), .dinb(n11416), .dout(n11420));
  jxor g11228(.dina(n11420), .dinb(n11414), .dout(n11421));
  jxor g11229(.dina(n11421), .dinb(n11409), .dout(n11422));
  jxor g11230(.dina(n11422), .dinb(n11401), .dout(n11423));
  jand g11231(.dina(n11217), .dinb(n11139), .dout(n11424));
  jand g11232(.dina(n11218), .dinb(n11134), .dout(n11425));
  jor  g11233(.dina(n11425), .dinb(n11424), .dout(n11426));
  jand g11234(.dina(n11230), .dinb(n11228), .dout(n11427));
  jand g11235(.dina(n11234), .dinb(n11231), .dout(n11428));
  jor  g11236(.dina(n11428), .dinb(n11427), .dout(n11429));
  jand g11237(.dina(n11248), .dinb(n11246), .dout(n11430));
  jand g11238(.dina(n11251), .dinb(n11249), .dout(n11431));
  jor  g11239(.dina(n11431), .dinb(n11430), .dout(n11432));
  jnot g11240(.din(n11432), .dout(n11433));
  jand g11241(.dina(\a[54] ), .dinb(\a[27] ), .dout(n11434));
  jand g11242(.dina(\a[42] ), .dinb(\a[39] ), .dout(n11435));
  jor  g11243(.dina(n11435), .dinb(n11203), .dout(n11436));
  jnot g11244(.din(n11436), .dout(n11437));
  jand g11245(.dina(\a[43] ), .dinb(\a[39] ), .dout(n11438));
  jand g11246(.dina(n11438), .dinb(n11200), .dout(n11439));
  jor  g11247(.dina(n11439), .dinb(n11437), .dout(n11440));
  jxor g11248(.dina(n11440), .dinb(n11434), .dout(n11441));
  jxor g11249(.dina(n11441), .dinb(n11433), .dout(n11442));
  jxor g11250(.dina(n11442), .dinb(n11429), .dout(n11443));
  jand g11251(.dina(n11238), .dinb(n11235), .dout(n11444));
  jand g11252(.dina(n11242), .dinb(n11239), .dout(n11445));
  jor  g11253(.dina(n11445), .dinb(n11444), .dout(n11446));
  jand g11254(.dina(n11262), .dinb(n11256), .dout(n11447));
  jand g11255(.dina(n11263), .dinb(n11252), .dout(n11448));
  jor  g11256(.dina(n11448), .dinb(n11447), .dout(n11449));
  jxor g11257(.dina(n11449), .dinb(n11446), .dout(n11450));
  jxor g11258(.dina(n11450), .dinb(n11443), .dout(n11451));
  jxor g11259(.dina(n11451), .dinb(n11426), .dout(n11452));
  jxor g11260(.dina(n11452), .dinb(n11423), .dout(n11453));
  jxor g11261(.dina(n11453), .dinb(n11369), .dout(n11454));
  jxor g11262(.dina(n11454), .dinb(n11298), .dout(n11455));
  jand g11263(.dina(n11289), .dinb(n11128), .dout(n11456));
  jnot g11264(.din(n11128), .dout(n11457));
  jnot g11265(.din(n11289), .dout(n11458));
  jand g11266(.dina(n11458), .dinb(n11457), .dout(n11459));
  jnot g11267(.din(n11459), .dout(n11460));
  jand g11268(.dina(n11294), .dinb(n11460), .dout(n11461));
  jor  g11269(.dina(n11461), .dinb(n11456), .dout(n11462));
  jxor g11270(.dina(n11462), .dinb(n11455), .dout(\asquared[82] ));
  jand g11271(.dina(n11368), .dinb(n11301), .dout(n11464));
  jand g11272(.dina(n11453), .dinb(n11369), .dout(n11465));
  jor  g11273(.dina(n11465), .dinb(n11464), .dout(n11466));
  jand g11274(.dina(n11451), .dinb(n11426), .dout(n11467));
  jand g11275(.dina(n11452), .dinb(n11423), .dout(n11468));
  jor  g11276(.dina(n11468), .dinb(n11467), .dout(n11469));
  jand g11277(.dina(n11400), .dinb(n11372), .dout(n11470));
  jand g11278(.dina(n11422), .dinb(n11401), .dout(n11471));
  jor  g11279(.dina(n11471), .dinb(n11470), .dout(n11472));
  jand g11280(.dina(n11449), .dinb(n11446), .dout(n11473));
  jand g11281(.dina(n11450), .dinb(n11443), .dout(n11474));
  jor  g11282(.dina(n11474), .dinb(n11473), .dout(n11475));
  jor  g11283(.dina(n11441), .dinb(n11433), .dout(n11476));
  jand g11284(.dina(n11442), .dinb(n11429), .dout(n11477));
  jnot g11285(.din(n11477), .dout(n11478));
  jand g11286(.dina(n11478), .dinb(n11476), .dout(n11479));
  jnot g11287(.din(n11479), .dout(n11480));
  jand g11288(.dina(\a[60] ), .dinb(\a[22] ), .dout(n11481));
  jnot g11289(.din(n11481), .dout(n11482));
  jand g11290(.dina(\a[58] ), .dinb(\a[24] ), .dout(n11483));
  jand g11291(.dina(\a[59] ), .dinb(\a[23] ), .dout(n11484));
  jor  g11292(.dina(n11484), .dinb(n11483), .dout(n11485));
  jand g11293(.dina(\a[59] ), .dinb(\a[24] ), .dout(n11486));
  jand g11294(.dina(n11486), .dinb(n11321), .dout(n11487));
  jnot g11295(.din(n11487), .dout(n11488));
  jand g11296(.dina(n11488), .dinb(n11485), .dout(n11489));
  jxor g11297(.dina(n11489), .dinb(n11482), .dout(n11490));
  jnot g11298(.din(n11394), .dout(n11491));
  jand g11299(.dina(\a[49] ), .dinb(\a[33] ), .dout(n11492));
  jor  g11300(.dina(n11492), .dinb(n11315), .dout(n11493));
  jand g11301(.dina(\a[49] ), .dinb(\a[34] ), .dout(n11494));
  jand g11302(.dina(n11494), .dinb(n11312), .dout(n11495));
  jnot g11303(.din(n11495), .dout(n11496));
  jand g11304(.dina(n11496), .dinb(n11493), .dout(n11497));
  jxor g11305(.dina(n11497), .dinb(n11491), .dout(n11498));
  jand g11306(.dina(\a[62] ), .dinb(\a[20] ), .dout(n11499));
  jnot g11307(.din(n11499), .dout(n11500));
  jand g11308(.dina(\a[51] ), .dinb(\a[31] ), .dout(n11501));
  jxor g11309(.dina(n11501), .dinb(n11349), .dout(n11502));
  jxor g11310(.dina(n11502), .dinb(n11500), .dout(n11503));
  jnot g11311(.din(n11503), .dout(n11504));
  jxor g11312(.dina(n11504), .dinb(n11498), .dout(n11505));
  jxor g11313(.dina(n11505), .dinb(n11490), .dout(n11506));
  jxor g11314(.dina(n11506), .dinb(n11480), .dout(n11507));
  jand g11315(.dina(\a[47] ), .dinb(\a[35] ), .dout(n11508));
  jand g11316(.dina(\a[46] ), .dinb(\a[36] ), .dout(n11509));
  jor  g11317(.dina(n11509), .dinb(n11340), .dout(n11510));
  jnot g11318(.din(n11510), .dout(n11511));
  jand g11319(.dina(\a[46] ), .dinb(\a[37] ), .dout(n11512));
  jand g11320(.dina(n11512), .dinb(n11154), .dout(n11513));
  jor  g11321(.dina(n11513), .dinb(n11511), .dout(n11514));
  jxor g11322(.dina(n11514), .dinb(n11508), .dout(n11515));
  jand g11323(.dina(\a[42] ), .dinb(\a[40] ), .dout(n11516));
  jand g11324(.dina(\a[52] ), .dinb(\a[30] ), .dout(n11517));
  jor  g11325(.dina(n11517), .dinb(n11361), .dout(n11518));
  jnot g11326(.din(n11518), .dout(n11519));
  jand g11327(.dina(\a[53] ), .dinb(\a[30] ), .dout(n11520));
  jand g11328(.dina(n11520), .dinb(n11358), .dout(n11521));
  jor  g11329(.dina(n11521), .dinb(n11519), .dout(n11522));
  jxor g11330(.dina(n11522), .dinb(n11516), .dout(n11523));
  jand g11331(.dina(\a[44] ), .dinb(\a[38] ), .dout(n11524));
  jor  g11332(.dina(n11524), .dinb(n11438), .dout(n11525));
  jand g11333(.dina(\a[44] ), .dinb(\a[39] ), .dout(n11526));
  jand g11334(.dina(n11526), .dinb(n11203), .dout(n11527));
  jnot g11335(.din(n11527), .dout(n11528));
  jand g11336(.dina(n11528), .dinb(n11525), .dout(n11529));
  jxor g11337(.dina(n11529), .dinb(n11209), .dout(n11530));
  jxor g11338(.dina(n11530), .dinb(n11523), .dout(n11531));
  jxor g11339(.dina(n11531), .dinb(n11515), .dout(n11532));
  jxor g11340(.dina(n11532), .dinb(n11507), .dout(n11533));
  jxor g11341(.dina(n11533), .dinb(n11475), .dout(n11534));
  jxor g11342(.dina(n11534), .dinb(n11472), .dout(n11535));
  jxor g11343(.dina(n11535), .dinb(n11469), .dout(n11536));
  jand g11344(.dina(n11334), .dinb(n11310), .dout(n11537));
  jand g11345(.dina(n11365), .dinb(n11335), .dout(n11538));
  jor  g11346(.dina(n11538), .dinb(n11537), .dout(n11539));
  jand g11347(.dina(n11314), .dinb(n8326), .dout(n11540));
  jor  g11348(.dina(n11540), .dinb(n11316), .dout(n11541));
  jand g11349(.dina(n11392), .dinb(n11390), .dout(n11542));
  jor  g11350(.dina(n11542), .dinb(n11395), .dout(n11543));
  jxor g11351(.dina(n11543), .dinb(n11541), .dout(n11544));
  jnot g11352(.din(n11360), .dout(n11545));
  jand g11353(.dina(n11545), .dinb(n11356), .dout(n11546));
  jor  g11354(.dina(n11546), .dinb(n11362), .dout(n11547));
  jxor g11355(.dina(n11547), .dinb(n11544), .dout(n11548));
  jand g11356(.dina(n11352), .dinb(n11345), .dout(n11549));
  jor  g11357(.dina(n11549), .dinb(n11350), .dout(n11550));
  jand g11358(.dina(n11322), .dinb(n11171), .dout(n11551));
  jor  g11359(.dina(n11551), .dinb(n11324), .dout(n11552));
  jxor g11360(.dina(n11552), .dinb(n11550), .dout(n11553));
  jand g11361(.dina(n11338), .dinb(n11336), .dout(n11554));
  jor  g11362(.dina(n11554), .dinb(n11341), .dout(n11555));
  jxor g11363(.dina(n11555), .dinb(n11553), .dout(n11556));
  jnot g11364(.din(n11556), .dout(n11557));
  jand g11365(.dina(n11353), .dinb(n11344), .dout(n11558));
  jnot g11366(.din(n11558), .dout(n11559));
  jor  g11367(.dina(n11364), .dinb(n11355), .dout(n11560));
  jand g11368(.dina(n11560), .dinb(n11559), .dout(n11561));
  jxor g11369(.dina(n11561), .dinb(n11557), .dout(n11562));
  jxor g11370(.dina(n11562), .dinb(n11548), .dout(n11563));
  jxor g11371(.dina(n11563), .dinb(n11539), .dout(n11564));
  jnot g11372(.din(n11327), .dout(n11565));
  jand g11373(.dina(n11332), .dinb(n11565), .dout(n11566));
  jnot g11374(.din(n11566), .dout(n11567));
  jand g11375(.dina(n11331), .dinb(n11327), .dout(n11568));
  jor  g11376(.dina(n11568), .dinb(n11319), .dout(n11569));
  jand g11377(.dina(n11569), .dinb(n11567), .dout(n11570));
  jnot g11378(.din(n11570), .dout(n11571));
  jnot g11379(.din(n11386), .dout(n11572));
  jnot g11380(.din(n11388), .dout(n11573));
  jand g11381(.dina(n11573), .dinb(n11572), .dout(n11574));
  jnot g11382(.din(n11574), .dout(n11575));
  jand g11383(.dina(n11388), .dinb(n11386), .dout(n11576));
  jor  g11384(.dina(n11398), .dinb(n11576), .dout(n11577));
  jand g11385(.dina(n11577), .dinb(n11575), .dout(n11578));
  jxor g11386(.dina(n11578), .dinb(n11571), .dout(n11579));
  jnot g11387(.din(\a[41] ), .dout(n11580));
  jand g11388(.dina(n11328), .dinb(n11329), .dout(n11581));
  jor  g11389(.dina(n11581), .dinb(n11580), .dout(n11582));
  jnot g11390(.din(n11582), .dout(n11583));
  jxor g11391(.dina(n11583), .dinb(n10301), .dout(n11584));
  jand g11392(.dina(n11436), .dinb(n11434), .dout(n11585));
  jor  g11393(.dina(n11585), .dinb(n11439), .dout(n11586));
  jxor g11394(.dina(n11586), .dinb(n11584), .dout(n11587));
  jxor g11395(.dina(n11587), .dinb(n11579), .dout(n11588));
  jxor g11396(.dina(n11588), .dinb(n11564), .dout(n11589));
  jand g11397(.dina(n11366), .dinb(n11307), .dout(n11590));
  jand g11398(.dina(n11367), .dinb(n11304), .dout(n11591));
  jor  g11399(.dina(n11591), .dinb(n11590), .dout(n11592));
  jand g11400(.dina(n11407), .dinb(n11405), .dout(n11593));
  jand g11401(.dina(n11408), .dinb(n11403), .dout(n11594));
  jor  g11402(.dina(n11594), .dinb(n11593), .dout(n11595));
  jand g11403(.dina(n11376), .dinb(n11374), .dout(n11596));
  jand g11404(.dina(n11379), .dinb(n11377), .dout(n11597));
  jor  g11405(.dina(n11597), .dinb(n11596), .dout(n11598));
  jand g11406(.dina(\a[55] ), .dinb(\a[28] ), .dout(n11599));
  jand g11407(.dina(n11599), .dinb(n11434), .dout(n11600));
  jand g11408(.dina(\a[57] ), .dinb(\a[25] ), .dout(n11601));
  jand g11409(.dina(n11601), .dinb(n5845), .dout(n11602));
  jor  g11410(.dina(n11602), .dinb(n11600), .dout(n11603));
  jand g11411(.dina(\a[57] ), .dinb(\a[27] ), .dout(n11604));
  jand g11412(.dina(n11604), .dinb(n11198), .dout(n11605));
  jnot g11413(.din(n11605), .dout(n11606));
  jand g11414(.dina(n11606), .dinb(n11603), .dout(n11607));
  jnot g11415(.din(n11607), .dout(n11608));
  jand g11416(.dina(\a[55] ), .dinb(\a[27] ), .dout(n11609));
  jor  g11417(.dina(n11609), .dinb(n11601), .dout(n11610));
  jand g11418(.dina(n11610), .dinb(n11606), .dout(n11611));
  jor  g11419(.dina(n11611), .dinb(n5845), .dout(n11612));
  jand g11420(.dina(n11612), .dinb(n11608), .dout(n11613));
  jxor g11421(.dina(n11613), .dinb(n11598), .dout(n11614));
  jxor g11422(.dina(n11614), .dinb(n11595), .dout(n11615));
  jand g11423(.dina(n11383), .dinb(n11380), .dout(n11616));
  jand g11424(.dina(n11399), .dinb(n11384), .dout(n11617));
  jor  g11425(.dina(n11617), .dinb(n11616), .dout(n11618));
  jand g11426(.dina(n11420), .dinb(n11414), .dout(n11619));
  jand g11427(.dina(n11421), .dinb(n11409), .dout(n11620));
  jor  g11428(.dina(n11620), .dinb(n11619), .dout(n11621));
  jxor g11429(.dina(n11621), .dinb(n11618), .dout(n11622));
  jxor g11430(.dina(n11622), .dinb(n11615), .dout(n11623));
  jxor g11431(.dina(n11623), .dinb(n11592), .dout(n11624));
  jxor g11432(.dina(n11624), .dinb(n11589), .dout(n11625));
  jxor g11433(.dina(n11625), .dinb(n11536), .dout(n11626));
  jxor g11434(.dina(n11626), .dinb(n11466), .dout(n11627));
  jand g11435(.dina(n11454), .dinb(n11298), .dout(n11628));
  jor  g11436(.dina(n11454), .dinb(n11298), .dout(n11629));
  jand g11437(.dina(n11462), .dinb(n11629), .dout(n11630));
  jor  g11438(.dina(n11630), .dinb(n11628), .dout(n11631));
  jxor g11439(.dina(n11631), .dinb(n11627), .dout(\asquared[83] ));
  jand g11440(.dina(n11535), .dinb(n11469), .dout(n11633));
  jand g11441(.dina(n11625), .dinb(n11536), .dout(n11634));
  jor  g11442(.dina(n11634), .dinb(n11633), .dout(n11635));
  jand g11443(.dina(n11623), .dinb(n11592), .dout(n11636));
  jand g11444(.dina(n11624), .dinb(n11589), .dout(n11637));
  jor  g11445(.dina(n11637), .dinb(n11636), .dout(n11638));
  jand g11446(.dina(n11563), .dinb(n11539), .dout(n11639));
  jand g11447(.dina(n11588), .dinb(n11564), .dout(n11640));
  jor  g11448(.dina(n11640), .dinb(n11639), .dout(n11641));
  jand g11449(.dina(n11621), .dinb(n11618), .dout(n11642));
  jand g11450(.dina(n11622), .dinb(n11615), .dout(n11643));
  jor  g11451(.dina(n11643), .dinb(n11642), .dout(n11644));
  jand g11452(.dina(n11613), .dinb(n11598), .dout(n11645));
  jand g11453(.dina(n11614), .dinb(n11595), .dout(n11646));
  jor  g11454(.dina(n11646), .dinb(n11645), .dout(n11647));
  jand g11455(.dina(\a[50] ), .dinb(\a[33] ), .dout(n11648));
  jnot g11456(.din(n11648), .dout(n11649));
  jand g11457(.dina(\a[48] ), .dinb(\a[35] ), .dout(n11650));
  jor  g11458(.dina(n11650), .dinb(n11494), .dout(n11651));
  jand g11459(.dina(\a[49] ), .dinb(\a[35] ), .dout(n11652));
  jand g11460(.dina(n11652), .dinb(n11315), .dout(n11653));
  jnot g11461(.din(n11653), .dout(n11654));
  jand g11462(.dina(n11654), .dinb(n11651), .dout(n11655));
  jxor g11463(.dina(n11655), .dinb(n11649), .dout(n11656));
  jand g11464(.dina(\a[54] ), .dinb(\a[29] ), .dout(n11657));
  jnot g11465(.din(n11657), .dout(n11658));
  jand g11466(.dina(\a[43] ), .dinb(\a[40] ), .dout(n11659));
  jor  g11467(.dina(n11659), .dinb(n11526), .dout(n11660));
  jand g11468(.dina(\a[44] ), .dinb(\a[40] ), .dout(n11661));
  jand g11469(.dina(n11661), .dinb(n11438), .dout(n11662));
  jnot g11470(.din(n11662), .dout(n11663));
  jand g11471(.dina(n11663), .dinb(n11660), .dout(n11664));
  jxor g11472(.dina(n11664), .dinb(n11658), .dout(n11665));
  jand g11473(.dina(\a[62] ), .dinb(\a[21] ), .dout(n11666));
  jnot g11474(.din(n11666), .dout(n11667));
  jand g11475(.dina(\a[42] ), .dinb(n11580), .dout(n11668));
  jxor g11476(.dina(n11668), .dinb(n11667), .dout(n11669));
  jnot g11477(.din(n11669), .dout(n11670));
  jxor g11478(.dina(n11670), .dinb(n11665), .dout(n11671));
  jxor g11479(.dina(n11671), .dinb(n11656), .dout(n11672));
  jxor g11480(.dina(n11672), .dinb(n11647), .dout(n11673));
  jand g11481(.dina(\a[63] ), .dinb(\a[20] ), .dout(n11674));
  jand g11482(.dina(\a[61] ), .dinb(\a[22] ), .dout(n11675));
  jor  g11483(.dina(n11675), .dinb(n11674), .dout(n11676));
  jnot g11484(.din(n11676), .dout(n11677));
  jand g11485(.dina(\a[63] ), .dinb(\a[22] ), .dout(n11678));
  jand g11486(.dina(n11678), .dinb(n11346), .dout(n11679));
  jor  g11487(.dina(n11679), .dinb(n11677), .dout(n11680));
  jxor g11488(.dina(n11680), .dinb(n10978), .dout(n11681));
  jand g11489(.dina(\a[47] ), .dinb(\a[36] ), .dout(n11682));
  jand g11490(.dina(\a[45] ), .dinb(\a[38] ), .dout(n11683));
  jor  g11491(.dina(n11683), .dinb(n11512), .dout(n11684));
  jnot g11492(.din(n11684), .dout(n11685));
  jand g11493(.dina(\a[46] ), .dinb(\a[38] ), .dout(n11686));
  jand g11494(.dina(n11686), .dinb(n11340), .dout(n11687));
  jor  g11495(.dina(n11687), .dinb(n11685), .dout(n11688));
  jxor g11496(.dina(n11688), .dinb(n11682), .dout(n11689));
  jand g11497(.dina(\a[51] ), .dinb(\a[32] ), .dout(n11690));
  jor  g11498(.dina(n11690), .dinb(n10327), .dout(n11691));
  jand g11499(.dina(\a[57] ), .dinb(\a[32] ), .dout(n11692));
  jand g11500(.dina(n11692), .dinb(n10629), .dout(n11693));
  jnot g11501(.din(n11693), .dout(n11694));
  jand g11502(.dina(n11694), .dinb(n11691), .dout(n11695));
  jxor g11503(.dina(n11695), .dinb(n11323), .dout(n11696));
  jxor g11504(.dina(n11696), .dinb(n11689), .dout(n11697));
  jxor g11505(.dina(n11697), .dinb(n11681), .dout(n11698));
  jxor g11506(.dina(n11698), .dinb(n11673), .dout(n11699));
  jxor g11507(.dina(n11699), .dinb(n11644), .dout(n11700));
  jxor g11508(.dina(n11700), .dinb(n11641), .dout(n11701));
  jxor g11509(.dina(n11701), .dinb(n11638), .dout(n11702));
  jand g11510(.dina(n11533), .dinb(n11475), .dout(n11703));
  jand g11511(.dina(n11534), .dinb(n11472), .dout(n11704));
  jor  g11512(.dina(n11704), .dinb(n11703), .dout(n11705));
  jand g11513(.dina(n11543), .dinb(n11541), .dout(n11706));
  jand g11514(.dina(n11547), .dinb(n11544), .dout(n11707));
  jor  g11515(.dina(n11707), .dinb(n11706), .dout(n11708));
  jand g11516(.dina(n11552), .dinb(n11550), .dout(n11709));
  jand g11517(.dina(n11555), .dinb(n11553), .dout(n11710));
  jor  g11518(.dina(n11710), .dinb(n11709), .dout(n11711));
  jxor g11519(.dina(n11711), .dinb(n11708), .dout(n11712));
  jnot g11520(.din(n11712), .dout(n11713));
  jnot g11521(.din(n11498), .dout(n11714));
  jand g11522(.dina(n11504), .dinb(n11714), .dout(n11715));
  jnot g11523(.din(n11715), .dout(n11716));
  jand g11524(.dina(n11503), .dinb(n11498), .dout(n11717));
  jor  g11525(.dina(n11717), .dinb(n11490), .dout(n11718));
  jand g11526(.dina(n11718), .dinb(n11716), .dout(n11719));
  jxor g11527(.dina(n11719), .dinb(n11713), .dout(n11720));
  jand g11528(.dina(n11583), .dinb(n10301), .dout(n11721));
  jand g11529(.dina(n11586), .dinb(n11584), .dout(n11722));
  jor  g11530(.dina(n11722), .dinb(n11721), .dout(n11723));
  jand g11531(.dina(\a[60] ), .dinb(\a[23] ), .dout(n11724));
  jor  g11532(.dina(n11724), .dinb(n11486), .dout(n11725));
  jand g11533(.dina(\a[60] ), .dinb(\a[24] ), .dout(n11726));
  jand g11534(.dina(n11726), .dinb(n11484), .dout(n11727));
  jnot g11535(.din(n11727), .dout(n11728));
  jand g11536(.dina(n11728), .dinb(n11725), .dout(n11729));
  jand g11537(.dina(n11518), .dinb(n11516), .dout(n11730));
  jor  g11538(.dina(n11730), .dinb(n11521), .dout(n11731));
  jxor g11539(.dina(n11731), .dinb(n11729), .dout(n11732));
  jnot g11540(.din(n11732), .dout(n11733));
  jand g11541(.dina(\a[52] ), .dinb(\a[31] ), .dout(n11734));
  jor  g11542(.dina(n11599), .dinb(n11520), .dout(n11735));
  jnot g11543(.din(n11735), .dout(n11736));
  jand g11544(.dina(\a[55] ), .dinb(\a[30] ), .dout(n11737));
  jand g11545(.dina(n11737), .dinb(n11194), .dout(n11738));
  jor  g11546(.dina(n11738), .dinb(n11736), .dout(n11739));
  jxor g11547(.dina(n11739), .dinb(n11734), .dout(n11740));
  jxor g11548(.dina(n11740), .dinb(n11733), .dout(n11741));
  jxor g11549(.dina(n11741), .dinb(n11723), .dout(n11742));
  jand g11550(.dina(n11578), .dinb(n11571), .dout(n11743));
  jand g11551(.dina(n11587), .dinb(n11579), .dout(n11744));
  jor  g11552(.dina(n11744), .dinb(n11743), .dout(n11745));
  jxor g11553(.dina(n11745), .dinb(n11742), .dout(n11746));
  jxor g11554(.dina(n11746), .dinb(n11720), .dout(n11747));
  jxor g11555(.dina(n11747), .dinb(n11705), .dout(n11748));
  jand g11556(.dina(n11529), .dinb(n11209), .dout(n11749));
  jor  g11557(.dina(n11749), .dinb(n11527), .dout(n11750));
  jand g11558(.dina(n11485), .dinb(n11481), .dout(n11751));
  jor  g11559(.dina(n11751), .dinb(n11487), .dout(n11752));
  jand g11560(.dina(n11510), .dinb(n11508), .dout(n11753));
  jor  g11561(.dina(n11753), .dinb(n11513), .dout(n11754));
  jxor g11562(.dina(n11754), .dinb(n11752), .dout(n11755));
  jxor g11563(.dina(n11755), .dinb(n11750), .dout(n11756));
  jand g11564(.dina(n11493), .dinb(n11394), .dout(n11757));
  jor  g11565(.dina(n11757), .dinb(n11495), .dout(n11758));
  jnot g11566(.din(n11349), .dout(n11759));
  jnot g11567(.din(n11501), .dout(n11760));
  jand g11568(.dina(n11760), .dinb(n11759), .dout(n11761));
  jnot g11569(.din(n11761), .dout(n11762));
  jand g11570(.dina(n11501), .dinb(n11349), .dout(n11763));
  jor  g11571(.dina(n11763), .dinb(n11499), .dout(n11764));
  jand g11572(.dina(n11764), .dinb(n11762), .dout(n11765));
  jxor g11573(.dina(n11765), .dinb(n11758), .dout(n11766));
  jor  g11574(.dina(n11605), .dinb(n11603), .dout(n11767));
  jxor g11575(.dina(n11767), .dinb(n11766), .dout(n11768));
  jnot g11576(.din(n11523), .dout(n11769));
  jor  g11577(.dina(n11530), .dinb(n11769), .dout(n11770));
  jnot g11578(.din(n11515), .dout(n11771));
  jand g11579(.dina(n11530), .dinb(n11769), .dout(n11772));
  jor  g11580(.dina(n11772), .dinb(n11771), .dout(n11773));
  jand g11581(.dina(n11773), .dinb(n11770), .dout(n11774));
  jxor g11582(.dina(n11774), .dinb(n11768), .dout(n11775));
  jxor g11583(.dina(n11775), .dinb(n11756), .dout(n11776));
  jand g11584(.dina(n11506), .dinb(n11480), .dout(n11777));
  jand g11585(.dina(n11532), .dinb(n11507), .dout(n11778));
  jor  g11586(.dina(n11778), .dinb(n11777), .dout(n11779));
  jnot g11587(.din(n11779), .dout(n11780));
  jor  g11588(.dina(n11561), .dinb(n11557), .dout(n11781));
  jand g11589(.dina(n11562), .dinb(n11548), .dout(n11782));
  jnot g11590(.din(n11782), .dout(n11783));
  jand g11591(.dina(n11783), .dinb(n11781), .dout(n11784));
  jxor g11592(.dina(n11784), .dinb(n11780), .dout(n11785));
  jxor g11593(.dina(n11785), .dinb(n11776), .dout(n11786));
  jxor g11594(.dina(n11786), .dinb(n11748), .dout(n11787));
  jxor g11595(.dina(n11787), .dinb(n11702), .dout(n11788));
  jxor g11596(.dina(n11788), .dinb(n11635), .dout(n11789));
  jand g11597(.dina(n11626), .dinb(n11466), .dout(n11790));
  jor  g11598(.dina(n11626), .dinb(n11466), .dout(n11791));
  jand g11599(.dina(n11631), .dinb(n11791), .dout(n11792));
  jor  g11600(.dina(n11792), .dinb(n11790), .dout(n11793));
  jxor g11601(.dina(n11793), .dinb(n11789), .dout(\asquared[84] ));
  jand g11602(.dina(n11701), .dinb(n11638), .dout(n11795));
  jand g11603(.dina(n11787), .dinb(n11702), .dout(n11796));
  jor  g11604(.dina(n11796), .dinb(n11795), .dout(n11797));
  jand g11605(.dina(n11699), .dinb(n11644), .dout(n11798));
  jand g11606(.dina(n11700), .dinb(n11641), .dout(n11799));
  jor  g11607(.dina(n11799), .dinb(n11798), .dout(n11800));
  jnot g11608(.din(n11800), .dout(n11801));
  jor  g11609(.dina(n11784), .dinb(n11780), .dout(n11802));
  jand g11610(.dina(n11785), .dinb(n11776), .dout(n11803));
  jnot g11611(.din(n11803), .dout(n11804));
  jand g11612(.dina(n11804), .dinb(n11802), .dout(n11805));
  jxor g11613(.dina(n11805), .dinb(n11801), .dout(n11806));
  jand g11614(.dina(n11660), .dinb(n11657), .dout(n11807));
  jor  g11615(.dina(n11807), .dinb(n11662), .dout(n11808));
  jand g11616(.dina(n11667), .dinb(n11580), .dout(n11809));
  jor  g11617(.dina(n11809), .dinb(n3738), .dout(n11810));
  jnot g11618(.din(n11810), .dout(n11811));
  jxor g11619(.dina(n11811), .dinb(n11808), .dout(n11812));
  jand g11620(.dina(n11735), .dinb(n11734), .dout(n11813));
  jor  g11621(.dina(n11813), .dinb(n11738), .dout(n11814));
  jxor g11622(.dina(n11814), .dinb(n11812), .dout(n11815));
  jnot g11623(.din(n11665), .dout(n11816));
  jand g11624(.dina(n11670), .dinb(n11816), .dout(n11817));
  jnot g11625(.din(n11817), .dout(n11818));
  jand g11626(.dina(n11669), .dinb(n11665), .dout(n11819));
  jor  g11627(.dina(n11819), .dinb(n11656), .dout(n11820));
  jand g11628(.dina(n11820), .dinb(n11818), .dout(n11821));
  jnot g11629(.din(n11821), .dout(n11822));
  jnot g11630(.din(n11689), .dout(n11823));
  jor  g11631(.dina(n11696), .dinb(n11823), .dout(n11824));
  jnot g11632(.din(n11681), .dout(n11825));
  jand g11633(.dina(n11696), .dinb(n11823), .dout(n11826));
  jor  g11634(.dina(n11826), .dinb(n11825), .dout(n11827));
  jand g11635(.dina(n11827), .dinb(n11824), .dout(n11828));
  jxor g11636(.dina(n11828), .dinb(n11822), .dout(n11829));
  jxor g11637(.dina(n11829), .dinb(n11815), .dout(n11830));
  jand g11638(.dina(n11672), .dinb(n11647), .dout(n11831));
  jand g11639(.dina(n11698), .dinb(n11673), .dout(n11832));
  jor  g11640(.dina(n11832), .dinb(n11831), .dout(n11833));
  jand g11641(.dina(n11774), .dinb(n11768), .dout(n11834));
  jand g11642(.dina(n11775), .dinb(n11756), .dout(n11835));
  jor  g11643(.dina(n11835), .dinb(n11834), .dout(n11836));
  jxor g11644(.dina(n11836), .dinb(n11833), .dout(n11837));
  jxor g11645(.dina(n11837), .dinb(n11830), .dout(n11838));
  jxor g11646(.dina(n11838), .dinb(n11806), .dout(n11839));
  jand g11647(.dina(n11747), .dinb(n11705), .dout(n11840));
  jand g11648(.dina(n11786), .dinb(n11748), .dout(n11841));
  jor  g11649(.dina(n11841), .dinb(n11840), .dout(n11842));
  jor  g11650(.dina(n11740), .dinb(n11733), .dout(n11843));
  jand g11651(.dina(n11741), .dinb(n11723), .dout(n11844));
  jnot g11652(.din(n11844), .dout(n11845));
  jand g11653(.dina(n11845), .dinb(n11843), .dout(n11846));
  jnot g11654(.din(n11846), .dout(n11847));
  jand g11655(.dina(n11731), .dinb(n11729), .dout(n11848));
  jor  g11656(.dina(n11848), .dinb(n11727), .dout(n11849));
  jand g11657(.dina(n11676), .dinb(n10978), .dout(n11850));
  jor  g11658(.dina(n11850), .dinb(n11679), .dout(n11851));
  jxor g11659(.dina(n11851), .dinb(n11849), .dout(n11852));
  jand g11660(.dina(\a[58] ), .dinb(\a[26] ), .dout(n11853));
  jand g11661(.dina(\a[53] ), .dinb(\a[31] ), .dout(n11854));
  jand g11662(.dina(\a[52] ), .dinb(\a[32] ), .dout(n11855));
  jor  g11663(.dina(n11855), .dinb(n11854), .dout(n11856));
  jnot g11664(.din(n11856), .dout(n11857));
  jand g11665(.dina(\a[53] ), .dinb(\a[32] ), .dout(n11858));
  jand g11666(.dina(n11858), .dinb(n11734), .dout(n11859));
  jor  g11667(.dina(n11859), .dinb(n11857), .dout(n11860));
  jxor g11668(.dina(n11860), .dinb(n11853), .dout(n11861));
  jnot g11669(.din(n11861), .dout(n11862));
  jxor g11670(.dina(n11862), .dinb(n11852), .dout(n11863));
  jxor g11671(.dina(n11863), .dinb(n11847), .dout(n11864));
  jnot g11672(.din(n11864), .dout(n11865));
  jand g11673(.dina(n11711), .dinb(n11708), .dout(n11866));
  jnot g11674(.din(n11866), .dout(n11867));
  jor  g11675(.dina(n11719), .dinb(n11713), .dout(n11868));
  jand g11676(.dina(n11868), .dinb(n11867), .dout(n11869));
  jxor g11677(.dina(n11869), .dinb(n11865), .dout(n11870));
  jand g11678(.dina(n11745), .dinb(n11742), .dout(n11871));
  jand g11679(.dina(n11746), .dinb(n11720), .dout(n11872));
  jor  g11680(.dina(n11872), .dinb(n11871), .dout(n11873));
  jxor g11681(.dina(n11873), .dinb(n11870), .dout(n11874));
  jand g11682(.dina(\a[50] ), .dinb(\a[34] ), .dout(n11875));
  jand g11683(.dina(\a[48] ), .dinb(\a[36] ), .dout(n11876));
  jor  g11684(.dina(n11876), .dinb(n11652), .dout(n11877));
  jnot g11685(.din(n11877), .dout(n11878));
  jand g11686(.dina(\a[49] ), .dinb(\a[36] ), .dout(n11879));
  jand g11687(.dina(n11879), .dinb(n11650), .dout(n11880));
  jor  g11688(.dina(n11880), .dinb(n11878), .dout(n11881));
  jxor g11689(.dina(n11881), .dinb(n11875), .dout(n11882));
  jand g11690(.dina(\a[51] ), .dinb(\a[33] ), .dout(n11883));
  jand g11691(.dina(\a[59] ), .dinb(\a[25] ), .dout(n11884));
  jor  g11692(.dina(n11884), .dinb(n11726), .dout(n11885));
  jnot g11693(.din(n11885), .dout(n11886));
  jand g11694(.dina(\a[60] ), .dinb(\a[25] ), .dout(n11887));
  jand g11695(.dina(n11887), .dinb(n11486), .dout(n11888));
  jor  g11696(.dina(n11888), .dinb(n11886), .dout(n11889));
  jxor g11697(.dina(n11889), .dinb(n11883), .dout(n11890));
  jand g11698(.dina(\a[63] ), .dinb(\a[21] ), .dout(n11891));
  jand g11699(.dina(\a[62] ), .dinb(\a[22] ), .dout(n11892));
  jand g11700(.dina(\a[61] ), .dinb(\a[23] ), .dout(n11893));
  jor  g11701(.dina(n11893), .dinb(n11892), .dout(n11894));
  jand g11702(.dina(\a[62] ), .dinb(\a[23] ), .dout(n11895));
  jand g11703(.dina(n11895), .dinb(n11675), .dout(n11896));
  jnot g11704(.din(n11896), .dout(n11897));
  jand g11705(.dina(n11897), .dinb(n11894), .dout(n11898));
  jxor g11706(.dina(n11898), .dinb(n11891), .dout(n11899));
  jxor g11707(.dina(n11899), .dinb(n11890), .dout(n11900));
  jxor g11708(.dina(n11900), .dinb(n11882), .dout(n11901));
  jand g11709(.dina(\a[47] ), .dinb(\a[37] ), .dout(n11902));
  jnot g11710(.din(n11902), .dout(n11903));
  jand g11711(.dina(\a[54] ), .dinb(\a[30] ), .dout(n11904));
  jor  g11712(.dina(n11904), .dinb(n11604), .dout(n11905));
  jand g11713(.dina(\a[57] ), .dinb(\a[30] ), .dout(n11906));
  jand g11714(.dina(n11906), .dinb(n11434), .dout(n11907));
  jnot g11715(.din(n11907), .dout(n11908));
  jand g11716(.dina(n11908), .dinb(n11905), .dout(n11909));
  jxor g11717(.dina(n11909), .dinb(n11903), .dout(n11910));
  jand g11718(.dina(\a[45] ), .dinb(\a[39] ), .dout(n11911));
  jnot g11719(.din(n11911), .dout(n11912));
  jand g11720(.dina(\a[43] ), .dinb(\a[41] ), .dout(n11913));
  jor  g11721(.dina(n11913), .dinb(n11661), .dout(n11914));
  jand g11722(.dina(\a[44] ), .dinb(\a[41] ), .dout(n11915));
  jand g11723(.dina(n11915), .dinb(n11659), .dout(n11916));
  jnot g11724(.din(n11916), .dout(n11917));
  jand g11725(.dina(n11917), .dinb(n11914), .dout(n11918));
  jxor g11726(.dina(n11918), .dinb(n11912), .dout(n11919));
  jand g11727(.dina(\a[56] ), .dinb(\a[28] ), .dout(n11920));
  jnot g11728(.din(n11920), .dout(n11921));
  jand g11729(.dina(\a[55] ), .dinb(\a[29] ), .dout(n11922));
  jxor g11730(.dina(n11922), .dinb(n11686), .dout(n11923));
  jxor g11731(.dina(n11923), .dinb(n11921), .dout(n11924));
  jnot g11732(.din(n11924), .dout(n11925));
  jxor g11733(.dina(n11925), .dinb(n11919), .dout(n11926));
  jxor g11734(.dina(n11926), .dinb(n11910), .dout(n11927));
  jxor g11735(.dina(n11927), .dinb(n11901), .dout(n11928));
  jand g11736(.dina(n11695), .dinb(n11323), .dout(n11929));
  jor  g11737(.dina(n11929), .dinb(n11693), .dout(n11930));
  jand g11738(.dina(n11651), .dinb(n11648), .dout(n11931));
  jor  g11739(.dina(n11931), .dinb(n11653), .dout(n11932));
  jand g11740(.dina(n11684), .dinb(n11682), .dout(n11933));
  jor  g11741(.dina(n11933), .dinb(n11687), .dout(n11934));
  jxor g11742(.dina(n11934), .dinb(n11932), .dout(n11935));
  jxor g11743(.dina(n11935), .dinb(n11930), .dout(n11936));
  jand g11744(.dina(n11754), .dinb(n11752), .dout(n11937));
  jand g11745(.dina(n11755), .dinb(n11750), .dout(n11938));
  jor  g11746(.dina(n11938), .dinb(n11937), .dout(n11939));
  jand g11747(.dina(n11765), .dinb(n11758), .dout(n11940));
  jand g11748(.dina(n11767), .dinb(n11766), .dout(n11941));
  jor  g11749(.dina(n11941), .dinb(n11940), .dout(n11942));
  jxor g11750(.dina(n11942), .dinb(n11939), .dout(n11943));
  jxor g11751(.dina(n11943), .dinb(n11936), .dout(n11944));
  jxor g11752(.dina(n11944), .dinb(n11928), .dout(n11945));
  jxor g11753(.dina(n11945), .dinb(n11874), .dout(n11946));
  jxor g11754(.dina(n11946), .dinb(n11842), .dout(n11947));
  jxor g11755(.dina(n11947), .dinb(n11839), .dout(n11948));
  jxor g11756(.dina(n11948), .dinb(n11797), .dout(n11949));
  jand g11757(.dina(n11788), .dinb(n11635), .dout(n11950));
  jor  g11758(.dina(n11788), .dinb(n11635), .dout(n11951));
  jand g11759(.dina(n11793), .dinb(n11951), .dout(n11952));
  jor  g11760(.dina(n11952), .dinb(n11950), .dout(n11953));
  jxor g11761(.dina(n11953), .dinb(n11949), .dout(\asquared[85] ));
  jand g11762(.dina(n11946), .dinb(n11842), .dout(n11955));
  jand g11763(.dina(n11947), .dinb(n11839), .dout(n11956));
  jor  g11764(.dina(n11956), .dinb(n11955), .dout(n11957));
  jand g11765(.dina(n11836), .dinb(n11833), .dout(n11958));
  jand g11766(.dina(n11837), .dinb(n11830), .dout(n11959));
  jor  g11767(.dina(n11959), .dinb(n11958), .dout(n11960));
  jand g11768(.dina(n11934), .dinb(n11932), .dout(n11961));
  jand g11769(.dina(n11935), .dinb(n11930), .dout(n11962));
  jor  g11770(.dina(n11962), .dinb(n11961), .dout(n11963));
  jand g11771(.dina(n11811), .dinb(n11808), .dout(n11964));
  jand g11772(.dina(n11814), .dinb(n11812), .dout(n11965));
  jor  g11773(.dina(n11965), .dinb(n11964), .dout(n11966));
  jxor g11774(.dina(n11966), .dinb(n11963), .dout(n11967));
  jnot g11775(.din(n11849), .dout(n11968));
  jnot g11776(.din(n11851), .dout(n11969));
  jand g11777(.dina(n11969), .dinb(n11968), .dout(n11970));
  jnot g11778(.din(n11970), .dout(n11971));
  jand g11779(.dina(n11851), .dinb(n11849), .dout(n11972));
  jor  g11780(.dina(n11862), .dinb(n11972), .dout(n11973));
  jand g11781(.dina(n11973), .dinb(n11971), .dout(n11974));
  jxor g11782(.dina(n11974), .dinb(n11967), .dout(n11975));
  jnot g11783(.din(n11975), .dout(n11976));
  jand g11784(.dina(n11863), .dinb(n11847), .dout(n11977));
  jnot g11785(.din(n11977), .dout(n11978));
  jor  g11786(.dina(n11869), .dinb(n11865), .dout(n11979));
  jand g11787(.dina(n11979), .dinb(n11978), .dout(n11980));
  jxor g11788(.dina(n11980), .dinb(n11976), .dout(n11981));
  jand g11789(.dina(n11927), .dinb(n11901), .dout(n11982));
  jand g11790(.dina(n11944), .dinb(n11928), .dout(n11983));
  jor  g11791(.dina(n11983), .dinb(n11982), .dout(n11984));
  jxor g11792(.dina(n11984), .dinb(n11981), .dout(n11985));
  jxor g11793(.dina(n11985), .dinb(n11960), .dout(n11986));
  jand g11794(.dina(n11873), .dinb(n11870), .dout(n11987));
  jand g11795(.dina(n11945), .dinb(n11874), .dout(n11988));
  jor  g11796(.dina(n11988), .dinb(n11987), .dout(n11989));
  jxor g11797(.dina(n11989), .dinb(n11986), .dout(n11990));
  jor  g11798(.dina(n11805), .dinb(n11801), .dout(n11991));
  jand g11799(.dina(n11838), .dinb(n11806), .dout(n11992));
  jnot g11800(.din(n11992), .dout(n11993));
  jand g11801(.dina(n11993), .dinb(n11991), .dout(n11994));
  jnot g11802(.din(n11994), .dout(n11995));
  jand g11803(.dina(n11828), .dinb(n11822), .dout(n11996));
  jand g11804(.dina(n11829), .dinb(n11815), .dout(n11997));
  jor  g11805(.dina(n11997), .dinb(n11996), .dout(n11998));
  jand g11806(.dina(\a[46] ), .dinb(\a[39] ), .dout(n11999));
  jnot g11807(.din(n11999), .dout(n12000));
  jand g11808(.dina(\a[45] ), .dinb(\a[40] ), .dout(n12001));
  jor  g11809(.dina(n12001), .dinb(n11915), .dout(n12002));
  jand g11810(.dina(\a[45] ), .dinb(\a[41] ), .dout(n12003));
  jand g11811(.dina(n12003), .dinb(n11661), .dout(n12004));
  jnot g11812(.din(n12004), .dout(n12005));
  jand g11813(.dina(n12005), .dinb(n12002), .dout(n12006));
  jxor g11814(.dina(n12006), .dinb(n12000), .dout(n12007));
  jnot g11815(.din(n11858), .dout(n12008));
  jand g11816(.dina(\a[52] ), .dinb(\a[33] ), .dout(n12009));
  jand g11817(.dina(\a[51] ), .dinb(\a[34] ), .dout(n12010));
  jor  g11818(.dina(n12010), .dinb(n12009), .dout(n12011));
  jand g11819(.dina(\a[52] ), .dinb(\a[34] ), .dout(n12012));
  jand g11820(.dina(n12012), .dinb(n11883), .dout(n12013));
  jnot g11821(.din(n12013), .dout(n12014));
  jand g11822(.dina(n12014), .dinb(n12011), .dout(n12015));
  jxor g11823(.dina(n12015), .dinb(n12008), .dout(n12016));
  jand g11824(.dina(\a[50] ), .dinb(\a[35] ), .dout(n12017));
  jnot g11825(.din(n12017), .dout(n12018));
  jand g11826(.dina(\a[57] ), .dinb(\a[28] ), .dout(n12019));
  jxor g11827(.dina(n12019), .dinb(n11678), .dout(n12020));
  jxor g11828(.dina(n12020), .dinb(n12018), .dout(n12021));
  jnot g11829(.din(n12021), .dout(n12022));
  jxor g11830(.dina(n12022), .dinb(n12016), .dout(n12023));
  jxor g11831(.dina(n12023), .dinb(n12007), .dout(n12024));
  jand g11832(.dina(\a[56] ), .dinb(\a[29] ), .dout(n12025));
  jnot g11833(.din(n12025), .dout(n12026));
  jand g11834(.dina(\a[54] ), .dinb(\a[31] ), .dout(n12027));
  jor  g11835(.dina(n12027), .dinb(n11737), .dout(n12028));
  jand g11836(.dina(\a[55] ), .dinb(\a[31] ), .dout(n12029));
  jand g11837(.dina(n12029), .dinb(n11904), .dout(n12030));
  jnot g11838(.din(n12030), .dout(n12031));
  jand g11839(.dina(n12031), .dinb(n12028), .dout(n12032));
  jxor g11840(.dina(n12032), .dinb(n12026), .dout(n12033));
  jnot g11841(.din(n11879), .dout(n12034));
  jand g11842(.dina(\a[48] ), .dinb(\a[37] ), .dout(n12035));
  jand g11843(.dina(\a[47] ), .dinb(\a[38] ), .dout(n12036));
  jor  g11844(.dina(n12036), .dinb(n12035), .dout(n12037));
  jand g11845(.dina(\a[48] ), .dinb(\a[38] ), .dout(n12038));
  jand g11846(.dina(n12038), .dinb(n11902), .dout(n12039));
  jnot g11847(.din(n12039), .dout(n12040));
  jand g11848(.dina(n12040), .dinb(n12037), .dout(n12041));
  jxor g11849(.dina(n12041), .dinb(n12034), .dout(n12042));
  jnot g11850(.din(n11895), .dout(n12043));
  jand g11851(.dina(\a[43] ), .dinb(n3738), .dout(n12044));
  jxor g11852(.dina(n12044), .dinb(n12043), .dout(n12045));
  jnot g11853(.din(n12045), .dout(n12046));
  jxor g11854(.dina(n12046), .dinb(n12042), .dout(n12047));
  jxor g11855(.dina(n12047), .dinb(n12033), .dout(n12048));
  jxor g11856(.dina(n12048), .dinb(n12024), .dout(n12049));
  jxor g11857(.dina(n12049), .dinb(n11998), .dout(n12050));
  jand g11858(.dina(n11898), .dinb(n11891), .dout(n12051));
  jor  g11859(.dina(n12051), .dinb(n11896), .dout(n12052));
  jand g11860(.dina(n11877), .dinb(n11875), .dout(n12053));
  jor  g11861(.dina(n12053), .dinb(n11880), .dout(n12054));
  jxor g11862(.dina(n12054), .dinb(n12052), .dout(n12055));
  jand g11863(.dina(n11885), .dinb(n11883), .dout(n12056));
  jor  g11864(.dina(n12056), .dinb(n11888), .dout(n12057));
  jxor g11865(.dina(n12057), .dinb(n12055), .dout(n12058));
  jnot g11866(.din(n11919), .dout(n12059));
  jand g11867(.dina(n11925), .dinb(n12059), .dout(n12060));
  jnot g11868(.din(n12060), .dout(n12061));
  jand g11869(.dina(n11924), .dinb(n11919), .dout(n12062));
  jor  g11870(.dina(n12062), .dinb(n11910), .dout(n12063));
  jand g11871(.dina(n12063), .dinb(n12061), .dout(n12064));
  jnot g11872(.din(n12064), .dout(n12065));
  jnot g11873(.din(n11890), .dout(n12066));
  jor  g11874(.dina(n11899), .dinb(n12066), .dout(n12067));
  jnot g11875(.din(n11882), .dout(n12068));
  jand g11876(.dina(n11899), .dinb(n12066), .dout(n12069));
  jor  g11877(.dina(n12069), .dinb(n12068), .dout(n12070));
  jand g11878(.dina(n12070), .dinb(n12067), .dout(n12071));
  jxor g11879(.dina(n12071), .dinb(n12065), .dout(n12072));
  jxor g11880(.dina(n12072), .dinb(n12058), .dout(n12073));
  jand g11881(.dina(n11942), .dinb(n11939), .dout(n12074));
  jand g11882(.dina(n11943), .dinb(n11936), .dout(n12075));
  jor  g11883(.dina(n12075), .dinb(n12074), .dout(n12076));
  jand g11884(.dina(\a[61] ), .dinb(\a[24] ), .dout(n12077));
  jand g11885(.dina(n11914), .dinb(n11911), .dout(n12078));
  jor  g11886(.dina(n12078), .dinb(n11916), .dout(n12079));
  jxor g11887(.dina(n12079), .dinb(n12077), .dout(n12080));
  jnot g11888(.din(n12080), .dout(n12081));
  jand g11889(.dina(n11922), .dinb(n11686), .dout(n12082));
  jnot g11890(.din(n12082), .dout(n12083));
  jnot g11891(.din(n11686), .dout(n12084));
  jnot g11892(.din(n11922), .dout(n12085));
  jand g11893(.dina(n12085), .dinb(n12084), .dout(n12086));
  jor  g11894(.dina(n12086), .dinb(n11921), .dout(n12087));
  jand g11895(.dina(n12087), .dinb(n12083), .dout(n12088));
  jxor g11896(.dina(n12088), .dinb(n12081), .dout(n12089));
  jand g11897(.dina(n11856), .dinb(n11853), .dout(n12090));
  jor  g11898(.dina(n12090), .dinb(n11859), .dout(n12091));
  jand g11899(.dina(n11905), .dinb(n11902), .dout(n12092));
  jor  g11900(.dina(n12092), .dinb(n11907), .dout(n12093));
  jxor g11901(.dina(n12093), .dinb(n12091), .dout(n12094));
  jand g11902(.dina(\a[59] ), .dinb(\a[26] ), .dout(n12095));
  jand g11903(.dina(\a[58] ), .dinb(\a[27] ), .dout(n12096));
  jor  g11904(.dina(n12096), .dinb(n12095), .dout(n12097));
  jnot g11905(.din(n12097), .dout(n12098));
  jand g11906(.dina(n11853), .dinb(n6871), .dout(n12099));
  jor  g11907(.dina(n12099), .dinb(n12098), .dout(n12100));
  jxor g11908(.dina(n12100), .dinb(n11887), .dout(n12101));
  jnot g11909(.din(n12101), .dout(n12102));
  jxor g11910(.dina(n12102), .dinb(n12094), .dout(n12103));
  jxor g11911(.dina(n12103), .dinb(n12089), .dout(n12104));
  jxor g11912(.dina(n12104), .dinb(n12076), .dout(n12105));
  jxor g11913(.dina(n12105), .dinb(n12073), .dout(n12106));
  jxor g11914(.dina(n12106), .dinb(n12050), .dout(n12107));
  jxor g11915(.dina(n12107), .dinb(n11995), .dout(n12108));
  jxor g11916(.dina(n12108), .dinb(n11990), .dout(n12109));
  jxor g11917(.dina(n12109), .dinb(n11957), .dout(n12110));
  jand g11918(.dina(n11948), .dinb(n11797), .dout(n12111));
  jor  g11919(.dina(n11948), .dinb(n11797), .dout(n12112));
  jand g11920(.dina(n11953), .dinb(n12112), .dout(n12113));
  jor  g11921(.dina(n12113), .dinb(n12111), .dout(n12114));
  jxor g11922(.dina(n12114), .dinb(n12110), .dout(\asquared[86] ));
  jand g11923(.dina(n12107), .dinb(n11995), .dout(n12116));
  jand g11924(.dina(n12108), .dinb(n11990), .dout(n12117));
  jor  g11925(.dina(n12117), .dinb(n12116), .dout(n12118));
  jand g11926(.dina(n12105), .dinb(n12073), .dout(n12119));
  jand g11927(.dina(n12106), .dinb(n12050), .dout(n12120));
  jor  g11928(.dina(n12120), .dinb(n12119), .dout(n12121));
  jnot g11929(.din(n12121), .dout(n12122));
  jor  g11930(.dina(n11980), .dinb(n11976), .dout(n12123));
  jand g11931(.dina(n11984), .dinb(n11981), .dout(n12124));
  jnot g11932(.din(n12124), .dout(n12125));
  jand g11933(.dina(n12125), .dinb(n12123), .dout(n12126));
  jxor g11934(.dina(n12126), .dinb(n12122), .dout(n12127));
  jand g11935(.dina(n12103), .dinb(n12089), .dout(n12128));
  jand g11936(.dina(n12104), .dinb(n12076), .dout(n12129));
  jor  g11937(.dina(n12129), .dinb(n12128), .dout(n12130));
  jand g11938(.dina(n12079), .dinb(n12077), .dout(n12131));
  jnot g11939(.din(n12131), .dout(n12132));
  jor  g11940(.dina(n12088), .dinb(n12081), .dout(n12133));
  jand g11941(.dina(n12133), .dinb(n12132), .dout(n12134));
  jnot g11942(.din(n12134), .dout(n12135));
  jand g11943(.dina(\a[61] ), .dinb(\a[25] ), .dout(n12136));
  jand g11944(.dina(\a[62] ), .dinb(\a[24] ), .dout(n12137));
  jor  g11945(.dina(n12137), .dinb(n12136), .dout(n12138));
  jand g11946(.dina(\a[62] ), .dinb(\a[25] ), .dout(n12139));
  jand g11947(.dina(n12139), .dinb(n12077), .dout(n12140));
  jnot g11948(.din(n12140), .dout(n12141));
  jand g11949(.dina(n12141), .dinb(n12138), .dout(n12142));
  jnot g11950(.din(\a[43] ), .dout(n12143));
  jand g11951(.dina(n12043), .dinb(n3738), .dout(n12144));
  jor  g11952(.dina(n12144), .dinb(n12143), .dout(n12145));
  jnot g11953(.din(n12145), .dout(n12146));
  jxor g11954(.dina(n12146), .dinb(n12142), .dout(n12147));
  jxor g11955(.dina(n12147), .dinb(n12135), .dout(n12148));
  jand g11956(.dina(n12054), .dinb(n12052), .dout(n12149));
  jand g11957(.dina(n12057), .dinb(n12055), .dout(n12150));
  jor  g11958(.dina(n12150), .dinb(n12149), .dout(n12151));
  jxor g11959(.dina(n12151), .dinb(n12148), .dout(n12152));
  jxor g11960(.dina(n12152), .dinb(n12130), .dout(n12153));
  jand g11961(.dina(n12048), .dinb(n12024), .dout(n12154));
  jand g11962(.dina(n12049), .dinb(n11998), .dout(n12155));
  jor  g11963(.dina(n12155), .dinb(n12154), .dout(n12156));
  jxor g11964(.dina(n12156), .dinb(n12153), .dout(n12157));
  jxor g11965(.dina(n12157), .dinb(n12127), .dout(n12158));
  jand g11966(.dina(n11985), .dinb(n11960), .dout(n12159));
  jand g11967(.dina(n11989), .dinb(n11986), .dout(n12160));
  jor  g11968(.dina(n12160), .dinb(n12159), .dout(n12161));
  jnot g11969(.din(n12016), .dout(n12162));
  jand g11970(.dina(n12022), .dinb(n12162), .dout(n12163));
  jnot g11971(.din(n12163), .dout(n12164));
  jand g11972(.dina(n12021), .dinb(n12016), .dout(n12165));
  jor  g11973(.dina(n12165), .dinb(n12007), .dout(n12166));
  jand g11974(.dina(n12166), .dinb(n12164), .dout(n12167));
  jnot g11975(.din(n12167), .dout(n12168));
  jnot g11976(.din(n12091), .dout(n12169));
  jnot g11977(.din(n12093), .dout(n12170));
  jand g11978(.dina(n12170), .dinb(n12169), .dout(n12171));
  jnot g11979(.din(n12171), .dout(n12172));
  jand g11980(.dina(n12093), .dinb(n12091), .dout(n12173));
  jor  g11981(.dina(n12102), .dinb(n12173), .dout(n12174));
  jand g11982(.dina(n12174), .dinb(n12172), .dout(n12175));
  jxor g11983(.dina(n12175), .dinb(n12168), .dout(n12176));
  jnot g11984(.din(n12176), .dout(n12177));
  jnot g11985(.din(n12042), .dout(n12178));
  jand g11986(.dina(n12046), .dinb(n12178), .dout(n12179));
  jnot g11987(.din(n12179), .dout(n12180));
  jand g11988(.dina(n12045), .dinb(n12042), .dout(n12181));
  jor  g11989(.dina(n12181), .dinb(n12033), .dout(n12182));
  jand g11990(.dina(n12182), .dinb(n12180), .dout(n12183));
  jxor g11991(.dina(n12183), .dinb(n12177), .dout(n12184));
  jand g11992(.dina(n11966), .dinb(n11963), .dout(n12185));
  jand g11993(.dina(n11974), .dinb(n11967), .dout(n12186));
  jor  g11994(.dina(n12186), .dinb(n12185), .dout(n12187));
  jand g11995(.dina(n12002), .dinb(n11999), .dout(n12188));
  jor  g11996(.dina(n12188), .dinb(n12004), .dout(n12189));
  jand g11997(.dina(n12028), .dinb(n12025), .dout(n12190));
  jor  g11998(.dina(n12190), .dinb(n12030), .dout(n12191));
  jxor g11999(.dina(n12191), .dinb(n12189), .dout(n12192));
  jand g12000(.dina(n12037), .dinb(n11879), .dout(n12193));
  jor  g12001(.dina(n12193), .dinb(n12039), .dout(n12194));
  jxor g12002(.dina(n12194), .dinb(n12192), .dout(n12195));
  jand g12003(.dina(n12011), .dinb(n11858), .dout(n12196));
  jor  g12004(.dina(n12196), .dinb(n12013), .dout(n12197));
  jand g12005(.dina(n12097), .dinb(n11887), .dout(n12198));
  jor  g12006(.dina(n12198), .dinb(n12099), .dout(n12199));
  jxor g12007(.dina(n12199), .dinb(n12197), .dout(n12200));
  jnot g12008(.din(n11678), .dout(n12201));
  jnot g12009(.din(n12019), .dout(n12202));
  jand g12010(.dina(n12202), .dinb(n12201), .dout(n12203));
  jnot g12011(.din(n12203), .dout(n12204));
  jand g12012(.dina(n12019), .dinb(n11678), .dout(n12205));
  jor  g12013(.dina(n12205), .dinb(n12017), .dout(n12206));
  jand g12014(.dina(n12206), .dinb(n12204), .dout(n12207));
  jxor g12015(.dina(n12207), .dinb(n12200), .dout(n12208));
  jxor g12016(.dina(n12208), .dinb(n12195), .dout(n12209));
  jxor g12017(.dina(n12209), .dinb(n12187), .dout(n12210));
  jxor g12018(.dina(n12210), .dinb(n12184), .dout(n12211));
  jand g12019(.dina(n12071), .dinb(n12065), .dout(n12212));
  jand g12020(.dina(n12072), .dinb(n12058), .dout(n12213));
  jor  g12021(.dina(n12213), .dinb(n12212), .dout(n12214));
  jand g12022(.dina(\a[56] ), .dinb(\a[30] ), .dout(n12215));
  jand g12023(.dina(\a[46] ), .dinb(\a[40] ), .dout(n12216));
  jand g12024(.dina(\a[47] ), .dinb(\a[39] ), .dout(n12217));
  jor  g12025(.dina(n12217), .dinb(n12216), .dout(n12218));
  jnot g12026(.din(n12218), .dout(n12219));
  jand g12027(.dina(\a[47] ), .dinb(\a[40] ), .dout(n12220));
  jand g12028(.dina(n12220), .dinb(n11999), .dout(n12221));
  jor  g12029(.dina(n12221), .dinb(n12219), .dout(n12222));
  jxor g12030(.dina(n12222), .dinb(n12215), .dout(n12223));
  jnot g12031(.din(n12223), .dout(n12224));
  jand g12032(.dina(\a[60] ), .dinb(\a[26] ), .dout(n12225));
  jand g12033(.dina(\a[58] ), .dinb(\a[28] ), .dout(n12226));
  jor  g12034(.dina(n12226), .dinb(n6871), .dout(n12227));
  jand g12035(.dina(\a[59] ), .dinb(\a[28] ), .dout(n12228));
  jand g12036(.dina(n12228), .dinb(n12096), .dout(n12229));
  jnot g12037(.din(n12229), .dout(n12230));
  jand g12038(.dina(n12230), .dinb(n12227), .dout(n12231));
  jxor g12039(.dina(n12231), .dinb(n12225), .dout(n12232));
  jnot g12040(.din(n12232), .dout(n12233));
  jand g12041(.dina(\a[44] ), .dinb(\a[42] ), .dout(n12234));
  jnot g12042(.din(n12234), .dout(n12235));
  jand g12043(.dina(\a[54] ), .dinb(\a[32] ), .dout(n12236));
  jxor g12044(.dina(n12236), .dinb(n12235), .dout(n12237));
  jxor g12045(.dina(n12237), .dinb(n12003), .dout(n12238));
  jxor g12046(.dina(n12238), .dinb(n12233), .dout(n12239));
  jxor g12047(.dina(n12239), .dinb(n12224), .dout(n12240));
  jand g12048(.dina(\a[57] ), .dinb(\a[29] ), .dout(n12241));
  jor  g12049(.dina(n12241), .dinb(n12029), .dout(n12242));
  jnot g12050(.din(n12242), .dout(n12243));
  jand g12051(.dina(\a[57] ), .dinb(\a[31] ), .dout(n12244));
  jand g12052(.dina(n12244), .dinb(n11922), .dout(n12245));
  jor  g12053(.dina(n12245), .dinb(n12243), .dout(n12246));
  jxor g12054(.dina(n12246), .dinb(n12038), .dout(n12247));
  jand g12055(.dina(\a[53] ), .dinb(\a[33] ), .dout(n12248));
  jand g12056(.dina(\a[51] ), .dinb(\a[35] ), .dout(n12249));
  jor  g12057(.dina(n12249), .dinb(n12012), .dout(n12250));
  jnot g12058(.din(n12250), .dout(n12251));
  jand g12059(.dina(\a[52] ), .dinb(\a[35] ), .dout(n12252));
  jand g12060(.dina(n12252), .dinb(n12010), .dout(n12253));
  jor  g12061(.dina(n12253), .dinb(n12251), .dout(n12254));
  jxor g12062(.dina(n12254), .dinb(n12248), .dout(n12255));
  jand g12063(.dina(\a[63] ), .dinb(\a[23] ), .dout(n12256));
  jand g12064(.dina(\a[50] ), .dinb(\a[36] ), .dout(n12257));
  jand g12065(.dina(\a[49] ), .dinb(\a[37] ), .dout(n12258));
  jor  g12066(.dina(n12258), .dinb(n12257), .dout(n12259));
  jand g12067(.dina(\a[50] ), .dinb(\a[37] ), .dout(n12260));
  jand g12068(.dina(n12260), .dinb(n11879), .dout(n12261));
  jnot g12069(.din(n12261), .dout(n12262));
  jand g12070(.dina(n12262), .dinb(n12259), .dout(n12263));
  jxor g12071(.dina(n12263), .dinb(n12256), .dout(n12264));
  jxor g12072(.dina(n12264), .dinb(n12255), .dout(n12265));
  jxor g12073(.dina(n12265), .dinb(n12247), .dout(n12266));
  jxor g12074(.dina(n12266), .dinb(n12240), .dout(n12267));
  jxor g12075(.dina(n12267), .dinb(n12214), .dout(n12268));
  jxor g12076(.dina(n12268), .dinb(n12211), .dout(n12269));
  jxor g12077(.dina(n12269), .dinb(n12161), .dout(n12270));
  jxor g12078(.dina(n12270), .dinb(n12158), .dout(n12271));
  jxor g12079(.dina(n12271), .dinb(n12118), .dout(n12272));
  jand g12080(.dina(n12109), .dinb(n11957), .dout(n12273));
  jor  g12081(.dina(n12109), .dinb(n11957), .dout(n12274));
  jand g12082(.dina(n12114), .dinb(n12274), .dout(n12275));
  jor  g12083(.dina(n12275), .dinb(n12273), .dout(n12276));
  jxor g12084(.dina(n12276), .dinb(n12272), .dout(\asquared[87] ));
  jand g12085(.dina(n12269), .dinb(n12161), .dout(n12278));
  jand g12086(.dina(n12270), .dinb(n12158), .dout(n12279));
  jor  g12087(.dina(n12279), .dinb(n12278), .dout(n12280));
  jand g12088(.dina(n12266), .dinb(n12240), .dout(n12281));
  jand g12089(.dina(n12267), .dinb(n12214), .dout(n12282));
  jor  g12090(.dina(n12282), .dinb(n12281), .dout(n12283));
  jand g12091(.dina(n12191), .dinb(n12189), .dout(n12284));
  jand g12092(.dina(n12194), .dinb(n12192), .dout(n12285));
  jor  g12093(.dina(n12285), .dinb(n12284), .dout(n12286));
  jnot g12094(.din(n12255), .dout(n12287));
  jor  g12095(.dina(n12264), .dinb(n12287), .dout(n12288));
  jnot g12096(.din(n12247), .dout(n12289));
  jand g12097(.dina(n12264), .dinb(n12287), .dout(n12290));
  jor  g12098(.dina(n12290), .dinb(n12289), .dout(n12291));
  jand g12099(.dina(n12291), .dinb(n12288), .dout(n12292));
  jxor g12100(.dina(n12292), .dinb(n12286), .dout(n12293));
  jnot g12101(.din(n12293), .dout(n12294));
  jor  g12102(.dina(n12238), .dinb(n12233), .dout(n12295));
  jand g12103(.dina(n12239), .dinb(n12224), .dout(n12296));
  jnot g12104(.din(n12296), .dout(n12297));
  jand g12105(.dina(n12297), .dinb(n12295), .dout(n12298));
  jxor g12106(.dina(n12298), .dinb(n12294), .dout(n12299));
  jxor g12107(.dina(n12299), .dinb(n12283), .dout(n12300));
  jand g12108(.dina(n12152), .dinb(n12130), .dout(n12301));
  jand g12109(.dina(n12156), .dinb(n12153), .dout(n12302));
  jor  g12110(.dina(n12302), .dinb(n12301), .dout(n12303));
  jxor g12111(.dina(n12303), .dinb(n12300), .dout(n12304));
  jnot g12112(.din(n12304), .dout(n12305));
  jor  g12113(.dina(n12126), .dinb(n12122), .dout(n12306));
  jand g12114(.dina(n12157), .dinb(n12127), .dout(n12307));
  jnot g12115(.din(n12307), .dout(n12308));
  jand g12116(.dina(n12308), .dinb(n12306), .dout(n12309));
  jxor g12117(.dina(n12309), .dinb(n12305), .dout(n12310));
  jand g12118(.dina(n12210), .dinb(n12184), .dout(n12311));
  jand g12119(.dina(n12268), .dinb(n12211), .dout(n12312));
  jor  g12120(.dina(n12312), .dinb(n12311), .dout(n12313));
  jand g12121(.dina(n12199), .dinb(n12197), .dout(n12314));
  jand g12122(.dina(n12207), .dinb(n12200), .dout(n12315));
  jor  g12123(.dina(n12315), .dinb(n12314), .dout(n12316));
  jand g12124(.dina(\a[56] ), .dinb(\a[31] ), .dout(n12317));
  jand g12125(.dina(\a[54] ), .dinb(\a[33] ), .dout(n12318));
  jor  g12126(.dina(n12318), .dinb(n12317), .dout(n12319));
  jnot g12127(.din(n12319), .dout(n12320));
  jand g12128(.dina(\a[56] ), .dinb(\a[33] ), .dout(n12321));
  jand g12129(.dina(n12321), .dinb(n12027), .dout(n12322));
  jor  g12130(.dina(n12322), .dinb(n12320), .dout(n12323));
  jxor g12131(.dina(n12323), .dinb(n12220), .dout(n12324));
  jnot g12132(.din(n12139), .dout(n12325));
  jand g12133(.dina(\a[44] ), .dinb(n12143), .dout(n12326));
  jxor g12134(.dina(n12326), .dinb(n12325), .dout(n12327));
  jxor g12135(.dina(n12327), .dinb(n12324), .dout(n12328));
  jxor g12136(.dina(n12328), .dinb(n12316), .dout(n12329));
  jand g12137(.dina(\a[55] ), .dinb(\a[32] ), .dout(n12330));
  jand g12138(.dina(\a[46] ), .dinb(\a[41] ), .dout(n12331));
  jand g12139(.dina(\a[45] ), .dinb(\a[42] ), .dout(n12332));
  jor  g12140(.dina(n12332), .dinb(n12331), .dout(n12333));
  jnot g12141(.din(n12333), .dout(n12334));
  jand g12142(.dina(\a[46] ), .dinb(\a[42] ), .dout(n12335));
  jand g12143(.dina(n12335), .dinb(n12003), .dout(n12336));
  jor  g12144(.dina(n12336), .dinb(n12334), .dout(n12337));
  jxor g12145(.dina(n12337), .dinb(n12330), .dout(n12338));
  jand g12146(.dina(\a[49] ), .dinb(\a[38] ), .dout(n12339));
  jand g12147(.dina(\a[48] ), .dinb(\a[39] ), .dout(n12340));
  jor  g12148(.dina(n12340), .dinb(n12339), .dout(n12341));
  jnot g12149(.din(n12341), .dout(n12342));
  jand g12150(.dina(\a[49] ), .dinb(\a[39] ), .dout(n12343));
  jand g12151(.dina(n12343), .dinb(n12038), .dout(n12344));
  jor  g12152(.dina(n12344), .dinb(n12342), .dout(n12345));
  jxor g12153(.dina(n12345), .dinb(n12260), .dout(n12346));
  jand g12154(.dina(\a[63] ), .dinb(\a[24] ), .dout(n12347));
  jand g12155(.dina(\a[61] ), .dinb(\a[26] ), .dout(n12348));
  jand g12156(.dina(\a[60] ), .dinb(\a[27] ), .dout(n12349));
  jor  g12157(.dina(n12349), .dinb(n12348), .dout(n12350));
  jand g12158(.dina(\a[61] ), .dinb(\a[27] ), .dout(n12351));
  jand g12159(.dina(n12351), .dinb(n12225), .dout(n12352));
  jnot g12160(.din(n12352), .dout(n12353));
  jand g12161(.dina(n12353), .dinb(n12350), .dout(n12354));
  jxor g12162(.dina(n12354), .dinb(n12347), .dout(n12355));
  jxor g12163(.dina(n12355), .dinb(n12346), .dout(n12356));
  jxor g12164(.dina(n12356), .dinb(n12338), .dout(n12357));
  jxor g12165(.dina(n12357), .dinb(n12329), .dout(n12358));
  jnot g12166(.din(n12252), .dout(n12359));
  jand g12167(.dina(\a[58] ), .dinb(\a[29] ), .dout(n12360));
  jand g12168(.dina(\a[51] ), .dinb(\a[36] ), .dout(n12361));
  jxor g12169(.dina(n12361), .dinb(n12360), .dout(n12362));
  jxor g12170(.dina(n12362), .dinb(n12359), .dout(n12363));
  jnot g12171(.din(n12363), .dout(n12364));
  jnot g12172(.din(n12228), .dout(n12365));
  jand g12173(.dina(\a[53] ), .dinb(\a[34] ), .dout(n12366));
  jxor g12174(.dina(n12366), .dinb(n11906), .dout(n12367));
  jxor g12175(.dina(n12367), .dinb(n12365), .dout(n12368));
  jnot g12176(.din(n12368), .dout(n12369));
  jand g12177(.dina(n12146), .dinb(n12142), .dout(n12370));
  jor  g12178(.dina(n12370), .dinb(n12140), .dout(n12371));
  jxor g12179(.dina(n12371), .dinb(n12369), .dout(n12372));
  jxor g12180(.dina(n12372), .dinb(n12364), .dout(n12373));
  jxor g12181(.dina(n12373), .dinb(n12358), .dout(n12374));
  jxor g12182(.dina(n12374), .dinb(n12313), .dout(n12375));
  jand g12183(.dina(n12208), .dinb(n12195), .dout(n12376));
  jand g12184(.dina(n12209), .dinb(n12187), .dout(n12377));
  jor  g12185(.dina(n12377), .dinb(n12376), .dout(n12378));
  jand g12186(.dina(n12175), .dinb(n12168), .dout(n12379));
  jnot g12187(.din(n12379), .dout(n12380));
  jor  g12188(.dina(n12183), .dinb(n12177), .dout(n12381));
  jand g12189(.dina(n12381), .dinb(n12380), .dout(n12382));
  jnot g12190(.din(n12382), .dout(n12383));
  jxor g12191(.dina(n12383), .dinb(n12378), .dout(n12384));
  jand g12192(.dina(n12147), .dinb(n12135), .dout(n12385));
  jand g12193(.dina(n12151), .dinb(n12148), .dout(n12386));
  jor  g12194(.dina(n12386), .dinb(n12385), .dout(n12387));
  jand g12195(.dina(n12218), .dinb(n12215), .dout(n12388));
  jor  g12196(.dina(n12388), .dinb(n12221), .dout(n12389));
  jnot g12197(.din(n12236), .dout(n12390));
  jand g12198(.dina(n12390), .dinb(n12235), .dout(n12391));
  jnot g12199(.din(n12391), .dout(n12392));
  jand g12200(.dina(n12236), .dinb(n12234), .dout(n12393));
  jor  g12201(.dina(n12393), .dinb(n12003), .dout(n12394));
  jand g12202(.dina(n12394), .dinb(n12392), .dout(n12395));
  jxor g12203(.dina(n12395), .dinb(n12389), .dout(n12396));
  jand g12204(.dina(n12242), .dinb(n12038), .dout(n12397));
  jor  g12205(.dina(n12397), .dinb(n12245), .dout(n12398));
  jxor g12206(.dina(n12398), .dinb(n12396), .dout(n12399));
  jand g12207(.dina(n12263), .dinb(n12256), .dout(n12400));
  jor  g12208(.dina(n12400), .dinb(n12261), .dout(n12401));
  jand g12209(.dina(n12231), .dinb(n12225), .dout(n12402));
  jor  g12210(.dina(n12402), .dinb(n12229), .dout(n12403));
  jand g12211(.dina(n12250), .dinb(n12248), .dout(n12404));
  jor  g12212(.dina(n12404), .dinb(n12253), .dout(n12405));
  jxor g12213(.dina(n12405), .dinb(n12403), .dout(n12406));
  jxor g12214(.dina(n12406), .dinb(n12401), .dout(n12407));
  jxor g12215(.dina(n12407), .dinb(n12399), .dout(n12408));
  jxor g12216(.dina(n12408), .dinb(n12387), .dout(n12409));
  jxor g12217(.dina(n12409), .dinb(n12384), .dout(n12410));
  jxor g12218(.dina(n12410), .dinb(n12375), .dout(n12411));
  jxor g12219(.dina(n12411), .dinb(n12310), .dout(n12412));
  jxor g12220(.dina(n12412), .dinb(n12280), .dout(n12413));
  jand g12221(.dina(n12271), .dinb(n12118), .dout(n12414));
  jnot g12222(.din(n12118), .dout(n12415));
  jnot g12223(.din(n12271), .dout(n12416));
  jand g12224(.dina(n12416), .dinb(n12415), .dout(n12417));
  jnot g12225(.din(n12417), .dout(n12418));
  jand g12226(.dina(n12276), .dinb(n12418), .dout(n12419));
  jor  g12227(.dina(n12419), .dinb(n12414), .dout(n12420));
  jxor g12228(.dina(n12420), .dinb(n12413), .dout(\asquared[88] ));
  jor  g12229(.dina(n12309), .dinb(n12305), .dout(n12422));
  jand g12230(.dina(n12411), .dinb(n12310), .dout(n12423));
  jnot g12231(.din(n12423), .dout(n12424));
  jand g12232(.dina(n12424), .dinb(n12422), .dout(n12425));
  jand g12233(.dina(n12374), .dinb(n12313), .dout(n12426));
  jand g12234(.dina(n12410), .dinb(n12375), .dout(n12427));
  jor  g12235(.dina(n12427), .dinb(n12426), .dout(n12428));
  jand g12236(.dina(n12383), .dinb(n12378), .dout(n12429));
  jand g12237(.dina(n12409), .dinb(n12384), .dout(n12430));
  jor  g12238(.dina(n12430), .dinb(n12429), .dout(n12431));
  jand g12239(.dina(n12405), .dinb(n12403), .dout(n12432));
  jand g12240(.dina(n12406), .dinb(n12401), .dout(n12433));
  jor  g12241(.dina(n12433), .dinb(n12432), .dout(n12434));
  jand g12242(.dina(n12371), .dinb(n12369), .dout(n12435));
  jand g12243(.dina(n12372), .dinb(n12364), .dout(n12436));
  jor  g12244(.dina(n12436), .dinb(n12435), .dout(n12437));
  jxor g12245(.dina(n12437), .dinb(n12434), .dout(n12438));
  jnot g12246(.din(n12346), .dout(n12439));
  jor  g12247(.dina(n12355), .dinb(n12439), .dout(n12440));
  jnot g12248(.din(n12338), .dout(n12441));
  jand g12249(.dina(n12355), .dinb(n12439), .dout(n12442));
  jor  g12250(.dina(n12442), .dinb(n12441), .dout(n12443));
  jand g12251(.dina(n12443), .dinb(n12440), .dout(n12444));
  jxor g12252(.dina(n12444), .dinb(n12438), .dout(n12445));
  jand g12253(.dina(n12357), .dinb(n12329), .dout(n12446));
  jand g12254(.dina(n12373), .dinb(n12358), .dout(n12447));
  jor  g12255(.dina(n12447), .dinb(n12446), .dout(n12448));
  jxor g12256(.dina(n12448), .dinb(n12445), .dout(n12449));
  jxor g12257(.dina(n12449), .dinb(n12431), .dout(n12450));
  jxor g12258(.dina(n12450), .dinb(n12428), .dout(n12451));
  jand g12259(.dina(n12407), .dinb(n12399), .dout(n12452));
  jand g12260(.dina(n12408), .dinb(n12387), .dout(n12453));
  jor  g12261(.dina(n12453), .dinb(n12452), .dout(n12454));
  jnot g12262(.din(n12454), .dout(n12455));
  jand g12263(.dina(n12292), .dinb(n12286), .dout(n12456));
  jnot g12264(.din(n12456), .dout(n12457));
  jor  g12265(.dina(n12298), .dinb(n12294), .dout(n12458));
  jand g12266(.dina(n12458), .dinb(n12457), .dout(n12459));
  jxor g12267(.dina(n12459), .dinb(n12455), .dout(n12460));
  jand g12268(.dina(n12354), .dinb(n12347), .dout(n12461));
  jor  g12269(.dina(n12461), .dinb(n12352), .dout(n12462));
  jnot g12270(.din(n12462), .dout(n12463));
  jand g12271(.dina(n12366), .dinb(n11906), .dout(n12464));
  jnot g12272(.din(n12464), .dout(n12465));
  jnot g12273(.din(n11906), .dout(n12466));
  jnot g12274(.din(n12366), .dout(n12467));
  jand g12275(.dina(n12467), .dinb(n12466), .dout(n12468));
  jor  g12276(.dina(n12468), .dinb(n12365), .dout(n12469));
  jand g12277(.dina(n12469), .dinb(n12465), .dout(n12470));
  jxor g12278(.dina(n12470), .dinb(n12463), .dout(n12471));
  jand g12279(.dina(n12341), .dinb(n12260), .dout(n12472));
  jor  g12280(.dina(n12472), .dinb(n12344), .dout(n12473));
  jxor g12281(.dina(n12473), .dinb(n12471), .dout(n12474));
  jor  g12282(.dina(n12327), .dinb(n12324), .dout(n12475));
  jand g12283(.dina(n12328), .dinb(n12316), .dout(n12476));
  jnot g12284(.din(n12476), .dout(n12477));
  jand g12285(.dina(n12477), .dinb(n12475), .dout(n12478));
  jnot g12286(.din(n12478), .dout(n12479));
  jand g12287(.dina(n12319), .dinb(n12220), .dout(n12480));
  jor  g12288(.dina(n12480), .dinb(n12322), .dout(n12481));
  jnot g12289(.din(n12481), .dout(n12482));
  jand g12290(.dina(n12361), .dinb(n12360), .dout(n12483));
  jnot g12291(.din(n12483), .dout(n12484));
  jnot g12292(.din(n12360), .dout(n12485));
  jnot g12293(.din(n12361), .dout(n12486));
  jand g12294(.dina(n12486), .dinb(n12485), .dout(n12487));
  jor  g12295(.dina(n12487), .dinb(n12359), .dout(n12488));
  jand g12296(.dina(n12488), .dinb(n12484), .dout(n12489));
  jxor g12297(.dina(n12489), .dinb(n12482), .dout(n12490));
  jand g12298(.dina(\a[45] ), .dinb(\a[43] ), .dout(n12491));
  jand g12299(.dina(\a[55] ), .dinb(\a[33] ), .dout(n12492));
  jand g12300(.dina(\a[54] ), .dinb(\a[34] ), .dout(n12493));
  jor  g12301(.dina(n12493), .dinb(n12492), .dout(n12494));
  jnot g12302(.din(n12494), .dout(n12495));
  jand g12303(.dina(\a[55] ), .dinb(\a[34] ), .dout(n12496));
  jand g12304(.dina(n12496), .dinb(n12318), .dout(n12497));
  jor  g12305(.dina(n12497), .dinb(n12495), .dout(n12498));
  jxor g12306(.dina(n12498), .dinb(n12491), .dout(n12499));
  jnot g12307(.din(n12499), .dout(n12500));
  jxor g12308(.dina(n12500), .dinb(n12490), .dout(n12501));
  jxor g12309(.dina(n12501), .dinb(n12479), .dout(n12502));
  jxor g12310(.dina(n12502), .dinb(n12474), .dout(n12503));
  jxor g12311(.dina(n12503), .dinb(n12460), .dout(n12504));
  jand g12312(.dina(n12299), .dinb(n12283), .dout(n12505));
  jand g12313(.dina(n12303), .dinb(n12300), .dout(n12506));
  jor  g12314(.dina(n12506), .dinb(n12505), .dout(n12507));
  jand g12315(.dina(n12395), .dinb(n12389), .dout(n12508));
  jand g12316(.dina(n12398), .dinb(n12396), .dout(n12509));
  jor  g12317(.dina(n12509), .dinb(n12508), .dout(n12510));
  jand g12318(.dina(\a[48] ), .dinb(\a[40] ), .dout(n12511));
  jand g12319(.dina(\a[58] ), .dinb(\a[30] ), .dout(n12512));
  jand g12320(.dina(\a[56] ), .dinb(\a[32] ), .dout(n12513));
  jor  g12321(.dina(n12513), .dinb(n12512), .dout(n12514));
  jnot g12322(.din(n12514), .dout(n12515));
  jand g12323(.dina(\a[58] ), .dinb(\a[32] ), .dout(n12516));
  jand g12324(.dina(n12516), .dinb(n12215), .dout(n12517));
  jor  g12325(.dina(n12517), .dinb(n12515), .dout(n12518));
  jxor g12326(.dina(n12518), .dinb(n12511), .dout(n12519));
  jnot g12327(.din(n12519), .dout(n12520));
  jand g12328(.dina(\a[59] ), .dinb(\a[29] ), .dout(n12521));
  jand g12329(.dina(\a[50] ), .dinb(\a[38] ), .dout(n12522));
  jor  g12330(.dina(n12522), .dinb(n12343), .dout(n12523));
  jand g12331(.dina(\a[50] ), .dinb(\a[39] ), .dout(n12524));
  jand g12332(.dina(n12524), .dinb(n12339), .dout(n12525));
  jnot g12333(.din(n12525), .dout(n12526));
  jand g12334(.dina(n12526), .dinb(n12523), .dout(n12527));
  jxor g12335(.dina(n12527), .dinb(n12521), .dout(n12528));
  jxor g12336(.dina(n12528), .dinb(n12520), .dout(n12529));
  jxor g12337(.dina(n12529), .dinb(n12510), .dout(n12530));
  jand g12338(.dina(\a[63] ), .dinb(\a[25] ), .dout(n12531));
  jnot g12339(.din(\a[44] ), .dout(n12532));
  jand g12340(.dina(n12325), .dinb(n12143), .dout(n12533));
  jor  g12341(.dina(n12533), .dinb(n12532), .dout(n12534));
  jnot g12342(.din(n12534), .dout(n12535));
  jxor g12343(.dina(n12535), .dinb(n12531), .dout(n12536));
  jand g12344(.dina(n12333), .dinb(n12330), .dout(n12537));
  jor  g12345(.dina(n12537), .dinb(n12336), .dout(n12538));
  jxor g12346(.dina(n12538), .dinb(n12536), .dout(n12539));
  jxor g12347(.dina(n12539), .dinb(n12530), .dout(n12540));
  jand g12348(.dina(\a[53] ), .dinb(\a[35] ), .dout(n12541));
  jand g12349(.dina(\a[51] ), .dinb(\a[37] ), .dout(n12542));
  jand g12350(.dina(\a[52] ), .dinb(\a[36] ), .dout(n12543));
  jor  g12351(.dina(n12543), .dinb(n12542), .dout(n12544));
  jnot g12352(.din(n12544), .dout(n12545));
  jand g12353(.dina(\a[52] ), .dinb(\a[37] ), .dout(n12546));
  jand g12354(.dina(n12546), .dinb(n12361), .dout(n12547));
  jor  g12355(.dina(n12547), .dinb(n12545), .dout(n12548));
  jxor g12356(.dina(n12548), .dinb(n12541), .dout(n12549));
  jand g12357(.dina(\a[47] ), .dinb(\a[41] ), .dout(n12550));
  jor  g12358(.dina(n12550), .dinb(n12335), .dout(n12551));
  jnot g12359(.din(n12551), .dout(n12552));
  jand g12360(.dina(\a[47] ), .dinb(\a[42] ), .dout(n12553));
  jand g12361(.dina(n12553), .dinb(n12331), .dout(n12554));
  jor  g12362(.dina(n12554), .dinb(n12552), .dout(n12555));
  jxor g12363(.dina(n12555), .dinb(n12244), .dout(n12556));
  jand g12364(.dina(\a[62] ), .dinb(\a[26] ), .dout(n12557));
  jand g12365(.dina(\a[60] ), .dinb(\a[28] ), .dout(n12558));
  jor  g12366(.dina(n12558), .dinb(n12351), .dout(n12559));
  jand g12367(.dina(\a[61] ), .dinb(\a[28] ), .dout(n12560));
  jand g12368(.dina(n12560), .dinb(n12349), .dout(n12561));
  jnot g12369(.din(n12561), .dout(n12562));
  jand g12370(.dina(n12562), .dinb(n12559), .dout(n12563));
  jxor g12371(.dina(n12563), .dinb(n12557), .dout(n12564));
  jxor g12372(.dina(n12564), .dinb(n12556), .dout(n12565));
  jxor g12373(.dina(n12565), .dinb(n12549), .dout(n12566));
  jxor g12374(.dina(n12566), .dinb(n12540), .dout(n12567));
  jxor g12375(.dina(n12567), .dinb(n12507), .dout(n12568));
  jxor g12376(.dina(n12568), .dinb(n12504), .dout(n12569));
  jxor g12377(.dina(n12569), .dinb(n12451), .dout(n12570));
  jnot g12378(.din(n12570), .dout(n12571));
  jxor g12379(.dina(n12571), .dinb(n12425), .dout(n12572));
  jand g12380(.dina(n12412), .dinb(n12280), .dout(n12573));
  jnot g12381(.din(n12280), .dout(n12574));
  jnot g12382(.din(n12412), .dout(n12575));
  jand g12383(.dina(n12575), .dinb(n12574), .dout(n12576));
  jnot g12384(.din(n12576), .dout(n12577));
  jand g12385(.dina(n12420), .dinb(n12577), .dout(n12578));
  jor  g12386(.dina(n12578), .dinb(n12573), .dout(n12579));
  jxor g12387(.dina(n12579), .dinb(n12572), .dout(\asquared[89] ));
  jand g12388(.dina(n12450), .dinb(n12428), .dout(n12581));
  jand g12389(.dina(n12569), .dinb(n12451), .dout(n12582));
  jor  g12390(.dina(n12582), .dinb(n12581), .dout(n12583));
  jor  g12391(.dina(n12459), .dinb(n12455), .dout(n12584));
  jand g12392(.dina(n12503), .dinb(n12460), .dout(n12585));
  jnot g12393(.din(n12585), .dout(n12586));
  jand g12394(.dina(n12586), .dinb(n12584), .dout(n12587));
  jnot g12395(.din(n12587), .dout(n12588));
  jand g12396(.dina(n12528), .dinb(n12520), .dout(n12589));
  jand g12397(.dina(n12529), .dinb(n12510), .dout(n12590));
  jor  g12398(.dina(n12590), .dinb(n12589), .dout(n12591));
  jnot g12399(.din(n12556), .dout(n12592));
  jor  g12400(.dina(n12564), .dinb(n12592), .dout(n12593));
  jnot g12401(.din(n12549), .dout(n12594));
  jand g12402(.dina(n12564), .dinb(n12592), .dout(n12595));
  jor  g12403(.dina(n12595), .dinb(n12594), .dout(n12596));
  jand g12404(.dina(n12596), .dinb(n12593), .dout(n12597));
  jxor g12405(.dina(n12597), .dinb(n12591), .dout(n12598));
  jand g12406(.dina(n12527), .dinb(n12521), .dout(n12599));
  jor  g12407(.dina(n12599), .dinb(n12525), .dout(n12600));
  jand g12408(.dina(n12551), .dinb(n12244), .dout(n12601));
  jor  g12409(.dina(n12601), .dinb(n12554), .dout(n12602));
  jxor g12410(.dina(n12602), .dinb(n12600), .dout(n12603));
  jand g12411(.dina(\a[63] ), .dinb(\a[26] ), .dout(n12604));
  jand g12412(.dina(\a[49] ), .dinb(\a[40] ), .dout(n12605));
  jor  g12413(.dina(n12605), .dinb(n12524), .dout(n12606));
  jnot g12414(.din(n12606), .dout(n12607));
  jand g12415(.dina(\a[50] ), .dinb(\a[40] ), .dout(n12608));
  jand g12416(.dina(n12608), .dinb(n12343), .dout(n12609));
  jor  g12417(.dina(n12609), .dinb(n12607), .dout(n12610));
  jxor g12418(.dina(n12610), .dinb(n12604), .dout(n12611));
  jnot g12419(.din(n12611), .dout(n12612));
  jxor g12420(.dina(n12612), .dinb(n12603), .dout(n12613));
  jxor g12421(.dina(n12613), .dinb(n12598), .dout(n12614));
  jor  g12422(.dina(n12539), .dinb(n12530), .dout(n12615));
  jand g12423(.dina(n12539), .dinb(n12530), .dout(n12616));
  jor  g12424(.dina(n12566), .dinb(n12616), .dout(n12617));
  jand g12425(.dina(n12617), .dinb(n12615), .dout(n12618));
  jxor g12426(.dina(n12618), .dinb(n12614), .dout(n12619));
  jxor g12427(.dina(n12619), .dinb(n12588), .dout(n12620));
  jand g12428(.dina(n12567), .dinb(n12507), .dout(n12621));
  jand g12429(.dina(n12568), .dinb(n12504), .dout(n12622));
  jor  g12430(.dina(n12622), .dinb(n12621), .dout(n12623));
  jxor g12431(.dina(n12623), .dinb(n12620), .dout(n12624));
  jor  g12432(.dina(n12470), .dinb(n12463), .dout(n12625));
  jand g12433(.dina(n12473), .dinb(n12471), .dout(n12626));
  jnot g12434(.din(n12626), .dout(n12627));
  jand g12435(.dina(n12627), .dinb(n12625), .dout(n12628));
  jnot g12436(.din(n12628), .dout(n12629));
  jand g12437(.dina(n12535), .dinb(n12531), .dout(n12630));
  jand g12438(.dina(n12538), .dinb(n12536), .dout(n12631));
  jor  g12439(.dina(n12631), .dinb(n12630), .dout(n12632));
  jxor g12440(.dina(n12632), .dinb(n12629), .dout(n12633));
  jand g12441(.dina(n12489), .dinb(n12482), .dout(n12634));
  jnot g12442(.din(n12634), .dout(n12635));
  jnot g12443(.din(n12489), .dout(n12636));
  jand g12444(.dina(n12636), .dinb(n12481), .dout(n12637));
  jor  g12445(.dina(n12500), .dinb(n12637), .dout(n12638));
  jand g12446(.dina(n12638), .dinb(n12635), .dout(n12639));
  jxor g12447(.dina(n12639), .dinb(n12633), .dout(n12640));
  jand g12448(.dina(n12437), .dinb(n12434), .dout(n12641));
  jand g12449(.dina(n12444), .dinb(n12438), .dout(n12642));
  jor  g12450(.dina(n12642), .dinb(n12641), .dout(n12643));
  jxor g12451(.dina(n12643), .dinb(n12640), .dout(n12644));
  jand g12452(.dina(n12501), .dinb(n12479), .dout(n12645));
  jand g12453(.dina(n12502), .dinb(n12474), .dout(n12646));
  jor  g12454(.dina(n12646), .dinb(n12645), .dout(n12647));
  jxor g12455(.dina(n12647), .dinb(n12644), .dout(n12648));
  jand g12456(.dina(n12448), .dinb(n12445), .dout(n12649));
  jand g12457(.dina(n12449), .dinb(n12431), .dout(n12650));
  jor  g12458(.dina(n12650), .dinb(n12649), .dout(n12651));
  jand g12459(.dina(n12563), .dinb(n12557), .dout(n12652));
  jor  g12460(.dina(n12652), .dinb(n12561), .dout(n12653));
  jand g12461(.dina(n12544), .dinb(n12541), .dout(n12654));
  jor  g12462(.dina(n12654), .dinb(n12547), .dout(n12655));
  jxor g12463(.dina(n12655), .dinb(n12653), .dout(n12656));
  jand g12464(.dina(n12514), .dinb(n12511), .dout(n12657));
  jor  g12465(.dina(n12657), .dinb(n12517), .dout(n12658));
  jxor g12466(.dina(n12658), .dinb(n12656), .dout(n12659));
  jand g12467(.dina(\a[60] ), .dinb(\a[29] ), .dout(n12660));
  jor  g12468(.dina(n12660), .dinb(n12560), .dout(n12661));
  jand g12469(.dina(\a[61] ), .dinb(\a[29] ), .dout(n12662));
  jand g12470(.dina(n12662), .dinb(n12558), .dout(n12663));
  jnot g12471(.din(n12663), .dout(n12664));
  jand g12472(.dina(n12664), .dinb(n12661), .dout(n12665));
  jand g12473(.dina(n12494), .dinb(n12491), .dout(n12666));
  jor  g12474(.dina(n12666), .dinb(n12497), .dout(n12667));
  jxor g12475(.dina(n12667), .dinb(n12665), .dout(n12668));
  jand g12476(.dina(\a[46] ), .dinb(\a[43] ), .dout(n12669));
  jor  g12477(.dina(n12669), .dinb(n12553), .dout(n12670));
  jnot g12478(.din(n12670), .dout(n12671));
  jand g12479(.dina(\a[47] ), .dinb(\a[43] ), .dout(n12672));
  jand g12480(.dina(n12672), .dinb(n12335), .dout(n12673));
  jor  g12481(.dina(n12673), .dinb(n12671), .dout(n12674));
  jxor g12482(.dina(n12674), .dinb(n12496), .dout(n12675));
  jand g12483(.dina(\a[62] ), .dinb(\a[27] ), .dout(n12676));
  jnot g12484(.din(n12676), .dout(n12677));
  jand g12485(.dina(\a[45] ), .dinb(n12532), .dout(n12678));
  jxor g12486(.dina(n12678), .dinb(n12677), .dout(n12679));
  jxor g12487(.dina(n12679), .dinb(n12675), .dout(n12680));
  jxor g12488(.dina(n12680), .dinb(n12668), .dout(n12681));
  jxor g12489(.dina(n12681), .dinb(n12659), .dout(n12682));
  jand g12490(.dina(\a[59] ), .dinb(\a[30] ), .dout(n12683));
  jand g12491(.dina(\a[58] ), .dinb(\a[31] ), .dout(n12684));
  jor  g12492(.dina(n12684), .dinb(n11692), .dout(n12685));
  jnot g12493(.din(n12685), .dout(n12686));
  jand g12494(.dina(n12516), .dinb(n12244), .dout(n12687));
  jor  g12495(.dina(n12687), .dinb(n12686), .dout(n12688));
  jxor g12496(.dina(n12688), .dinb(n12683), .dout(n12689));
  jand g12497(.dina(\a[53] ), .dinb(\a[36] ), .dout(n12690));
  jand g12498(.dina(\a[51] ), .dinb(\a[38] ), .dout(n12691));
  jor  g12499(.dina(n12691), .dinb(n12546), .dout(n12692));
  jnot g12500(.din(n12692), .dout(n12693));
  jand g12501(.dina(\a[52] ), .dinb(\a[38] ), .dout(n12694));
  jand g12502(.dina(n12694), .dinb(n12542), .dout(n12695));
  jor  g12503(.dina(n12695), .dinb(n12693), .dout(n12696));
  jxor g12504(.dina(n12696), .dinb(n12690), .dout(n12697));
  jand g12505(.dina(\a[48] ), .dinb(\a[41] ), .dout(n12698));
  jand g12506(.dina(\a[54] ), .dinb(\a[35] ), .dout(n12699));
  jor  g12507(.dina(n12699), .dinb(n12321), .dout(n12700));
  jand g12508(.dina(\a[56] ), .dinb(\a[35] ), .dout(n12701));
  jand g12509(.dina(n12701), .dinb(n12318), .dout(n12702));
  jnot g12510(.din(n12702), .dout(n12703));
  jand g12511(.dina(n12703), .dinb(n12700), .dout(n12704));
  jxor g12512(.dina(n12704), .dinb(n12698), .dout(n12705));
  jxor g12513(.dina(n12705), .dinb(n12697), .dout(n12706));
  jxor g12514(.dina(n12706), .dinb(n12689), .dout(n12707));
  jxor g12515(.dina(n12707), .dinb(n12682), .dout(n12708));
  jxor g12516(.dina(n12708), .dinb(n12651), .dout(n12709));
  jxor g12517(.dina(n12709), .dinb(n12648), .dout(n12710));
  jxor g12518(.dina(n12710), .dinb(n12624), .dout(n12711));
  jxor g12519(.dina(n12711), .dinb(n12583), .dout(n12712));
  jor  g12520(.dina(n12571), .dinb(n12425), .dout(n12713));
  jnot g12521(.din(n12713), .dout(n12714));
  jand g12522(.dina(n12571), .dinb(n12425), .dout(n12715));
  jnot g12523(.din(n12715), .dout(n12716));
  jand g12524(.dina(n12579), .dinb(n12716), .dout(n12717));
  jor  g12525(.dina(n12717), .dinb(n12714), .dout(n12718));
  jxor g12526(.dina(n12718), .dinb(n12712), .dout(\asquared[90] ));
  jand g12527(.dina(n12623), .dinb(n12620), .dout(n12720));
  jand g12528(.dina(n12710), .dinb(n12624), .dout(n12721));
  jor  g12529(.dina(n12721), .dinb(n12720), .dout(n12722));
  jand g12530(.dina(n12643), .dinb(n12640), .dout(n12723));
  jand g12531(.dina(n12647), .dinb(n12644), .dout(n12724));
  jor  g12532(.dina(n12724), .dinb(n12723), .dout(n12725));
  jand g12533(.dina(n12704), .dinb(n12698), .dout(n12726));
  jor  g12534(.dina(n12726), .dinb(n12702), .dout(n12727));
  jand g12535(.dina(n12670), .dinb(n12496), .dout(n12728));
  jor  g12536(.dina(n12728), .dinb(n12673), .dout(n12729));
  jnot g12537(.din(\a[45] ), .dout(n12730));
  jand g12538(.dina(n12677), .dinb(n12532), .dout(n12731));
  jor  g12539(.dina(n12731), .dinb(n12730), .dout(n12732));
  jnot g12540(.din(n12732), .dout(n12733));
  jxor g12541(.dina(n12733), .dinb(n12729), .dout(n12734));
  jxor g12542(.dina(n12734), .dinb(n12727), .dout(n12735));
  jor  g12543(.dina(n12679), .dinb(n12675), .dout(n12736));
  jand g12544(.dina(n12680), .dinb(n12668), .dout(n12737));
  jnot g12545(.din(n12737), .dout(n12738));
  jand g12546(.dina(n12738), .dinb(n12736), .dout(n12739));
  jnot g12547(.din(n12739), .dout(n12740));
  jnot g12548(.din(n12697), .dout(n12741));
  jor  g12549(.dina(n12705), .dinb(n12741), .dout(n12742));
  jnot g12550(.din(n12689), .dout(n12743));
  jand g12551(.dina(n12705), .dinb(n12741), .dout(n12744));
  jor  g12552(.dina(n12744), .dinb(n12743), .dout(n12745));
  jand g12553(.dina(n12745), .dinb(n12742), .dout(n12746));
  jxor g12554(.dina(n12746), .dinb(n12740), .dout(n12747));
  jxor g12555(.dina(n12747), .dinb(n12735), .dout(n12748));
  jor  g12556(.dina(n12681), .dinb(n12659), .dout(n12749));
  jand g12557(.dina(n12681), .dinb(n12659), .dout(n12750));
  jor  g12558(.dina(n12707), .dinb(n12750), .dout(n12751));
  jand g12559(.dina(n12751), .dinb(n12749), .dout(n12752));
  jxor g12560(.dina(n12752), .dinb(n12748), .dout(n12753));
  jxor g12561(.dina(n12753), .dinb(n12725), .dout(n12754));
  jand g12562(.dina(n12708), .dinb(n12651), .dout(n12755));
  jand g12563(.dina(n12709), .dinb(n12648), .dout(n12756));
  jor  g12564(.dina(n12756), .dinb(n12755), .dout(n12757));
  jxor g12565(.dina(n12757), .dinb(n12754), .dout(n12758));
  jand g12566(.dina(n12618), .dinb(n12614), .dout(n12759));
  jand g12567(.dina(n12619), .dinb(n12588), .dout(n12760));
  jor  g12568(.dina(n12760), .dinb(n12759), .dout(n12761));
  jand g12569(.dina(n12692), .dinb(n12690), .dout(n12762));
  jor  g12570(.dina(n12762), .dinb(n12695), .dout(n12763));
  jand g12571(.dina(n12685), .dinb(n12683), .dout(n12764));
  jor  g12572(.dina(n12764), .dinb(n12687), .dout(n12765));
  jxor g12573(.dina(n12765), .dinb(n12763), .dout(n12766));
  jand g12574(.dina(n12606), .dinb(n12604), .dout(n12767));
  jor  g12575(.dina(n12767), .dinb(n12609), .dout(n12768));
  jxor g12576(.dina(n12768), .dinb(n12766), .dout(n12769));
  jand g12577(.dina(n12632), .dinb(n12629), .dout(n12770));
  jand g12578(.dina(n12639), .dinb(n12633), .dout(n12771));
  jor  g12579(.dina(n12771), .dinb(n12770), .dout(n12772));
  jxor g12580(.dina(n12772), .dinb(n12769), .dout(n12773));
  jand g12581(.dina(\a[48] ), .dinb(\a[42] ), .dout(n12774));
  jand g12582(.dina(\a[46] ), .dinb(\a[44] ), .dout(n12775));
  jor  g12583(.dina(n12775), .dinb(n12672), .dout(n12776));
  jnot g12584(.din(n12776), .dout(n12777));
  jand g12585(.dina(\a[47] ), .dinb(\a[44] ), .dout(n12778));
  jand g12586(.dina(n12778), .dinb(n12669), .dout(n12779));
  jor  g12587(.dina(n12779), .dinb(n12777), .dout(n12780));
  jxor g12588(.dina(n12780), .dinb(n12774), .dout(n12781));
  jand g12589(.dina(\a[54] ), .dinb(\a[36] ), .dout(n12782));
  jand g12590(.dina(\a[53] ), .dinb(\a[37] ), .dout(n12783));
  jor  g12591(.dina(n12783), .dinb(n12694), .dout(n12784));
  jnot g12592(.din(n12784), .dout(n12785));
  jand g12593(.dina(\a[53] ), .dinb(\a[38] ), .dout(n12786));
  jand g12594(.dina(n12786), .dinb(n12546), .dout(n12787));
  jor  g12595(.dina(n12787), .dinb(n12785), .dout(n12788));
  jxor g12596(.dina(n12788), .dinb(n12782), .dout(n12789));
  jand g12597(.dina(\a[55] ), .dinb(\a[35] ), .dout(n12790));
  jand g12598(.dina(\a[57] ), .dinb(\a[33] ), .dout(n12791));
  jand g12599(.dina(\a[56] ), .dinb(\a[34] ), .dout(n12792));
  jor  g12600(.dina(n12792), .dinb(n12791), .dout(n12793));
  jand g12601(.dina(\a[57] ), .dinb(\a[34] ), .dout(n12794));
  jand g12602(.dina(n12794), .dinb(n12321), .dout(n12795));
  jnot g12603(.din(n12795), .dout(n12796));
  jand g12604(.dina(n12796), .dinb(n12793), .dout(n12797));
  jxor g12605(.dina(n12797), .dinb(n12790), .dout(n12798));
  jxor g12606(.dina(n12798), .dinb(n12789), .dout(n12799));
  jxor g12607(.dina(n12799), .dinb(n12781), .dout(n12800));
  jxor g12608(.dina(n12800), .dinb(n12773), .dout(n12801));
  jxor g12609(.dina(n12801), .dinb(n12761), .dout(n12802));
  jand g12610(.dina(n12597), .dinb(n12591), .dout(n12803));
  jand g12611(.dina(n12613), .dinb(n12598), .dout(n12804));
  jor  g12612(.dina(n12804), .dinb(n12803), .dout(n12805));
  jand g12613(.dina(n12655), .dinb(n12653), .dout(n12806));
  jand g12614(.dina(n12658), .dinb(n12656), .dout(n12807));
  jor  g12615(.dina(n12807), .dinb(n12806), .dout(n12808));
  jnot g12616(.din(n12808), .dout(n12809));
  jand g12617(.dina(\a[51] ), .dinb(\a[39] ), .dout(n12810));
  jand g12618(.dina(\a[49] ), .dinb(\a[41] ), .dout(n12811));
  jor  g12619(.dina(n12811), .dinb(n12608), .dout(n12812));
  jnot g12620(.din(n12812), .dout(n12813));
  jand g12621(.dina(\a[50] ), .dinb(\a[41] ), .dout(n12814));
  jand g12622(.dina(n12814), .dinb(n12605), .dout(n12815));
  jor  g12623(.dina(n12815), .dinb(n12813), .dout(n12816));
  jxor g12624(.dina(n12816), .dinb(n12810), .dout(n12817));
  jxor g12625(.dina(n12817), .dinb(n12809), .dout(n12818));
  jnot g12626(.din(n12600), .dout(n12819));
  jnot g12627(.din(n12602), .dout(n12820));
  jand g12628(.dina(n12820), .dinb(n12819), .dout(n12821));
  jnot g12629(.din(n12821), .dout(n12822));
  jand g12630(.dina(n12602), .dinb(n12600), .dout(n12823));
  jor  g12631(.dina(n12612), .dinb(n12823), .dout(n12824));
  jand g12632(.dina(n12824), .dinb(n12822), .dout(n12825));
  jxor g12633(.dina(n12825), .dinb(n12818), .dout(n12826));
  jand g12634(.dina(n12667), .dinb(n12665), .dout(n12827));
  jor  g12635(.dina(n12827), .dinb(n12663), .dout(n12828));
  jand g12636(.dina(\a[59] ), .dinb(\a[31] ), .dout(n12829));
  jor  g12637(.dina(n12829), .dinb(n12516), .dout(n12830));
  jand g12638(.dina(\a[59] ), .dinb(\a[32] ), .dout(n12831));
  jand g12639(.dina(n12831), .dinb(n12684), .dout(n12832));
  jnot g12640(.din(n12832), .dout(n12833));
  jand g12641(.dina(n12833), .dinb(n12830), .dout(n12834));
  jand g12642(.dina(\a[60] ), .dinb(\a[30] ), .dout(n12835));
  jxor g12643(.dina(n12835), .dinb(n12834), .dout(n12836));
  jxor g12644(.dina(n12836), .dinb(n12828), .dout(n12837));
  jand g12645(.dina(\a[63] ), .dinb(\a[27] ), .dout(n12838));
  jand g12646(.dina(\a[62] ), .dinb(\a[28] ), .dout(n12839));
  jor  g12647(.dina(n12839), .dinb(n12662), .dout(n12840));
  jand g12648(.dina(\a[62] ), .dinb(\a[29] ), .dout(n12841));
  jand g12649(.dina(n12841), .dinb(n12560), .dout(n12842));
  jnot g12650(.din(n12842), .dout(n12843));
  jand g12651(.dina(n12843), .dinb(n12840), .dout(n12844));
  jxor g12652(.dina(n12844), .dinb(n12838), .dout(n12845));
  jxor g12653(.dina(n12845), .dinb(n12837), .dout(n12846));
  jxor g12654(.dina(n12846), .dinb(n12826), .dout(n12847));
  jxor g12655(.dina(n12847), .dinb(n12805), .dout(n12848));
  jxor g12656(.dina(n12848), .dinb(n12802), .dout(n12849));
  jxor g12657(.dina(n12849), .dinb(n12758), .dout(n12850));
  jxor g12658(.dina(n12850), .dinb(n12722), .dout(n12851));
  jand g12659(.dina(n12711), .dinb(n12583), .dout(n12852));
  jor  g12660(.dina(n12711), .dinb(n12583), .dout(n12853));
  jand g12661(.dina(n12718), .dinb(n12853), .dout(n12854));
  jor  g12662(.dina(n12854), .dinb(n12852), .dout(n12855));
  jxor g12663(.dina(n12855), .dinb(n12851), .dout(\asquared[91] ));
  jand g12664(.dina(n12757), .dinb(n12754), .dout(n12857));
  jand g12665(.dina(n12849), .dinb(n12758), .dout(n12858));
  jor  g12666(.dina(n12858), .dinb(n12857), .dout(n12859));
  jand g12667(.dina(n12844), .dinb(n12838), .dout(n12860));
  jor  g12668(.dina(n12860), .dinb(n12842), .dout(n12861));
  jand g12669(.dina(n12784), .dinb(n12782), .dout(n12862));
  jor  g12670(.dina(n12862), .dinb(n12787), .dout(n12863));
  jxor g12671(.dina(n12863), .dinb(n12861), .dout(n12864));
  jand g12672(.dina(n12835), .dinb(n12834), .dout(n12865));
  jor  g12673(.dina(n12865), .dinb(n12832), .dout(n12866));
  jxor g12674(.dina(n12866), .dinb(n12864), .dout(n12867));
  jnot g12675(.din(n12867), .dout(n12868));
  jor  g12676(.dina(n12817), .dinb(n12809), .dout(n12869));
  jand g12677(.dina(n12825), .dinb(n12818), .dout(n12870));
  jnot g12678(.din(n12870), .dout(n12871));
  jand g12679(.dina(n12871), .dinb(n12869), .dout(n12872));
  jxor g12680(.dina(n12872), .dinb(n12868), .dout(n12873));
  jand g12681(.dina(\a[48] ), .dinb(\a[43] ), .dout(n12874));
  jor  g12682(.dina(n12874), .dinb(n12778), .dout(n12875));
  jnot g12683(.din(n12875), .dout(n12876));
  jand g12684(.dina(\a[48] ), .dinb(\a[44] ), .dout(n12877));
  jand g12685(.dina(n12877), .dinb(n12672), .dout(n12878));
  jor  g12686(.dina(n12878), .dinb(n12876), .dout(n12879));
  jxor g12687(.dina(n12879), .dinb(n12701), .dout(n12880));
  jnot g12688(.din(n12880), .dout(n12881));
  jand g12689(.dina(\a[63] ), .dinb(\a[28] ), .dout(n12882));
  jand g12690(.dina(\a[51] ), .dinb(\a[40] ), .dout(n12883));
  jor  g12691(.dina(n12883), .dinb(n12814), .dout(n12884));
  jand g12692(.dina(\a[51] ), .dinb(\a[41] ), .dout(n12885));
  jand g12693(.dina(n12885), .dinb(n12608), .dout(n12886));
  jnot g12694(.din(n12886), .dout(n12887));
  jand g12695(.dina(n12887), .dinb(n12884), .dout(n12888));
  jxor g12696(.dina(n12888), .dinb(n12882), .dout(n12889));
  jxor g12697(.dina(n12889), .dinb(n12881), .dout(n12890));
  jnot g12698(.din(n12841), .dout(n12891));
  jand g12699(.dina(\a[46] ), .dinb(n12730), .dout(n12892));
  jxor g12700(.dina(n12892), .dinb(n12891), .dout(n12893));
  jnot g12701(.din(n12893), .dout(n12894));
  jxor g12702(.dina(n12894), .dinb(n12890), .dout(n12895));
  jxor g12703(.dina(n12895), .dinb(n12873), .dout(n12896));
  jand g12704(.dina(n12752), .dinb(n12748), .dout(n12897));
  jand g12705(.dina(n12753), .dinb(n12725), .dout(n12898));
  jor  g12706(.dina(n12898), .dinb(n12897), .dout(n12899));
  jxor g12707(.dina(n12899), .dinb(n12896), .dout(n12900));
  jand g12708(.dina(n12765), .dinb(n12763), .dout(n12901));
  jand g12709(.dina(n12768), .dinb(n12766), .dout(n12902));
  jor  g12710(.dina(n12902), .dinb(n12901), .dout(n12903));
  jand g12711(.dina(n12733), .dinb(n12729), .dout(n12904));
  jand g12712(.dina(n12734), .dinb(n12727), .dout(n12905));
  jor  g12713(.dina(n12905), .dinb(n12904), .dout(n12906));
  jnot g12714(.din(n12906), .dout(n12907));
  jand g12715(.dina(\a[49] ), .dinb(\a[42] ), .dout(n12908));
  jand g12716(.dina(\a[55] ), .dinb(\a[36] ), .dout(n12909));
  jor  g12717(.dina(n12909), .dinb(n12794), .dout(n12910));
  jnot g12718(.din(n12910), .dout(n12911));
  jand g12719(.dina(\a[57] ), .dinb(\a[36] ), .dout(n12912));
  jand g12720(.dina(n12912), .dinb(n12496), .dout(n12913));
  jor  g12721(.dina(n12913), .dinb(n12911), .dout(n12914));
  jxor g12722(.dina(n12914), .dinb(n12908), .dout(n12915));
  jxor g12723(.dina(n12915), .dinb(n12907), .dout(n12916));
  jxor g12724(.dina(n12916), .dinb(n12903), .dout(n12917));
  jand g12725(.dina(n12746), .dinb(n12740), .dout(n12918));
  jand g12726(.dina(n12747), .dinb(n12735), .dout(n12919));
  jor  g12727(.dina(n12919), .dinb(n12918), .dout(n12920));
  jand g12728(.dina(\a[54] ), .dinb(\a[37] ), .dout(n12921));
  jnot g12729(.din(n12921), .dout(n12922));
  jand g12730(.dina(\a[52] ), .dinb(\a[39] ), .dout(n12923));
  jor  g12731(.dina(n12923), .dinb(n12786), .dout(n12924));
  jand g12732(.dina(\a[53] ), .dinb(\a[39] ), .dout(n12925));
  jand g12733(.dina(n12925), .dinb(n12694), .dout(n12926));
  jnot g12734(.din(n12926), .dout(n12927));
  jand g12735(.dina(n12927), .dinb(n12924), .dout(n12928));
  jxor g12736(.dina(n12928), .dinb(n12922), .dout(n12929));
  jand g12737(.dina(n12812), .dinb(n12810), .dout(n12930));
  jor  g12738(.dina(n12930), .dinb(n12815), .dout(n12931));
  jnot g12739(.din(n12931), .dout(n12932));
  jxor g12740(.dina(n12932), .dinb(n12929), .dout(n12933));
  jand g12741(.dina(\a[60] ), .dinb(\a[31] ), .dout(n12934));
  jand g12742(.dina(\a[58] ), .dinb(\a[33] ), .dout(n12935));
  jor  g12743(.dina(n12935), .dinb(n12831), .dout(n12936));
  jand g12744(.dina(\a[59] ), .dinb(\a[33] ), .dout(n12937));
  jand g12745(.dina(n12937), .dinb(n12516), .dout(n12938));
  jnot g12746(.din(n12938), .dout(n12939));
  jand g12747(.dina(n12939), .dinb(n12936), .dout(n12940));
  jxor g12748(.dina(n12940), .dinb(n12934), .dout(n12941));
  jxor g12749(.dina(n12941), .dinb(n12933), .dout(n12942));
  jxor g12750(.dina(n12942), .dinb(n12920), .dout(n12943));
  jxor g12751(.dina(n12943), .dinb(n12917), .dout(n12944));
  jxor g12752(.dina(n12944), .dinb(n12900), .dout(n12945));
  jand g12753(.dina(n12801), .dinb(n12761), .dout(n12946));
  jand g12754(.dina(n12848), .dinb(n12802), .dout(n12947));
  jor  g12755(.dina(n12947), .dinb(n12946), .dout(n12948));
  jand g12756(.dina(n12846), .dinb(n12826), .dout(n12949));
  jand g12757(.dina(n12847), .dinb(n12805), .dout(n12950));
  jor  g12758(.dina(n12950), .dinb(n12949), .dout(n12951));
  jand g12759(.dina(n12772), .dinb(n12769), .dout(n12952));
  jand g12760(.dina(n12800), .dinb(n12773), .dout(n12953));
  jor  g12761(.dina(n12953), .dinb(n12952), .dout(n12954));
  jand g12762(.dina(n12797), .dinb(n12790), .dout(n12955));
  jor  g12763(.dina(n12955), .dinb(n12795), .dout(n12956));
  jand g12764(.dina(\a[61] ), .dinb(\a[30] ), .dout(n12957));
  jand g12765(.dina(n12776), .dinb(n12774), .dout(n12958));
  jor  g12766(.dina(n12958), .dinb(n12779), .dout(n12959));
  jxor g12767(.dina(n12959), .dinb(n12957), .dout(n12960));
  jxor g12768(.dina(n12960), .dinb(n12956), .dout(n12961));
  jand g12769(.dina(n12836), .dinb(n12828), .dout(n12962));
  jand g12770(.dina(n12845), .dinb(n12837), .dout(n12963));
  jor  g12771(.dina(n12963), .dinb(n12962), .dout(n12964));
  jnot g12772(.din(n12789), .dout(n12965));
  jor  g12773(.dina(n12798), .dinb(n12965), .dout(n12966));
  jnot g12774(.din(n12781), .dout(n12967));
  jand g12775(.dina(n12798), .dinb(n12965), .dout(n12968));
  jor  g12776(.dina(n12968), .dinb(n12967), .dout(n12969));
  jand g12777(.dina(n12969), .dinb(n12966), .dout(n12970));
  jxor g12778(.dina(n12970), .dinb(n12964), .dout(n12971));
  jxor g12779(.dina(n12971), .dinb(n12961), .dout(n12972));
  jxor g12780(.dina(n12972), .dinb(n12954), .dout(n12973));
  jxor g12781(.dina(n12973), .dinb(n12951), .dout(n12974));
  jxor g12782(.dina(n12974), .dinb(n12948), .dout(n12975));
  jxor g12783(.dina(n12975), .dinb(n12945), .dout(n12976));
  jxor g12784(.dina(n12976), .dinb(n12859), .dout(n12977));
  jand g12785(.dina(n12850), .dinb(n12722), .dout(n12978));
  jnot g12786(.din(n12722), .dout(n12979));
  jnot g12787(.din(n12850), .dout(n12980));
  jand g12788(.dina(n12980), .dinb(n12979), .dout(n12981));
  jnot g12789(.din(n12981), .dout(n12982));
  jand g12790(.dina(n12855), .dinb(n12982), .dout(n12983));
  jor  g12791(.dina(n12983), .dinb(n12978), .dout(n12984));
  jxor g12792(.dina(n12984), .dinb(n12977), .dout(\asquared[92] ));
  jand g12793(.dina(n12972), .dinb(n12954), .dout(n12986));
  jand g12794(.dina(n12973), .dinb(n12951), .dout(n12987));
  jor  g12795(.dina(n12987), .dinb(n12986), .dout(n12988));
  jand g12796(.dina(n12942), .dinb(n12920), .dout(n12989));
  jand g12797(.dina(n12943), .dinb(n12917), .dout(n12990));
  jor  g12798(.dina(n12990), .dinb(n12989), .dout(n12991));
  jand g12799(.dina(n12970), .dinb(n12964), .dout(n12992));
  jand g12800(.dina(n12971), .dinb(n12961), .dout(n12993));
  jor  g12801(.dina(n12993), .dinb(n12992), .dout(n12994));
  jand g12802(.dina(n12959), .dinb(n12957), .dout(n12995));
  jand g12803(.dina(n12960), .dinb(n12956), .dout(n12996));
  jor  g12804(.dina(n12996), .dinb(n12995), .dout(n12997));
  jnot g12805(.din(\a[46] ), .dout(n12998));
  jand g12806(.dina(n12891), .dinb(n12730), .dout(n12999));
  jor  g12807(.dina(n12999), .dinb(n12998), .dout(n13000));
  jnot g12808(.din(n13000), .dout(n13001));
  jand g12809(.dina(\a[61] ), .dinb(\a[31] ), .dout(n13002));
  jand g12810(.dina(\a[62] ), .dinb(\a[30] ), .dout(n13003));
  jor  g12811(.dina(n13003), .dinb(n13002), .dout(n13004));
  jand g12812(.dina(\a[62] ), .dinb(\a[31] ), .dout(n13005));
  jand g12813(.dina(n13005), .dinb(n12957), .dout(n13006));
  jnot g12814(.din(n13006), .dout(n13007));
  jand g12815(.dina(n13007), .dinb(n13004), .dout(n13008));
  jxor g12816(.dina(n13008), .dinb(n13001), .dout(n13009));
  jnot g12817(.din(n13009), .dout(n13010));
  jand g12818(.dina(\a[52] ), .dinb(\a[40] ), .dout(n13011));
  jor  g12819(.dina(n13011), .dinb(n12885), .dout(n13012));
  jnot g12820(.din(n13012), .dout(n13013));
  jand g12821(.dina(\a[52] ), .dinb(\a[41] ), .dout(n13014));
  jand g12822(.dina(n13014), .dinb(n12883), .dout(n13015));
  jor  g12823(.dina(n13015), .dinb(n13013), .dout(n13016));
  jxor g12824(.dina(n13016), .dinb(n12925), .dout(n13017));
  jxor g12825(.dina(n13017), .dinb(n13010), .dout(n13018));
  jxor g12826(.dina(n13018), .dinb(n12997), .dout(n13019));
  jand g12827(.dina(\a[49] ), .dinb(\a[43] ), .dout(n13020));
  jnot g12828(.din(n13020), .dout(n13021));
  jand g12829(.dina(\a[47] ), .dinb(\a[45] ), .dout(n13022));
  jor  g12830(.dina(n13022), .dinb(n12877), .dout(n13023));
  jand g12831(.dina(\a[48] ), .dinb(\a[45] ), .dout(n13024));
  jand g12832(.dina(n13024), .dinb(n12778), .dout(n13025));
  jnot g12833(.din(n13025), .dout(n13026));
  jand g12834(.dina(n13026), .dinb(n13023), .dout(n13027));
  jxor g12835(.dina(n13027), .dinb(n13021), .dout(n13028));
  jand g12836(.dina(\a[58] ), .dinb(\a[34] ), .dout(n13029));
  jnot g12837(.din(n13029), .dout(n13030));
  jand g12838(.dina(\a[50] ), .dinb(\a[42] ), .dout(n13031));
  jand g12839(.dina(\a[57] ), .dinb(\a[35] ), .dout(n13032));
  jxor g12840(.dina(n13032), .dinb(n13031), .dout(n13033));
  jxor g12841(.dina(n13033), .dinb(n13030), .dout(n13034));
  jxor g12842(.dina(n13034), .dinb(n13028), .dout(n13035));
  jand g12843(.dina(\a[56] ), .dinb(\a[36] ), .dout(n13036));
  jnot g12844(.din(n12937), .dout(n13037));
  jxor g12845(.dina(n13037), .dinb(n11162), .dout(n13038));
  jxor g12846(.dina(n13038), .dinb(n13036), .dout(n13039));
  jnot g12847(.din(n13039), .dout(n13040));
  jxor g12848(.dina(n13040), .dinb(n13035), .dout(n13041));
  jxor g12849(.dina(n13041), .dinb(n13019), .dout(n13042));
  jxor g12850(.dina(n13042), .dinb(n12994), .dout(n13043));
  jxor g12851(.dina(n13043), .dinb(n12991), .dout(n13044));
  jxor g12852(.dina(n13044), .dinb(n12988), .dout(n13045));
  jand g12853(.dina(n12899), .dinb(n12896), .dout(n13046));
  jand g12854(.dina(n12944), .dinb(n12900), .dout(n13047));
  jor  g12855(.dina(n13047), .dinb(n13046), .dout(n13048));
  jand g12856(.dina(n12863), .dinb(n12861), .dout(n13049));
  jand g12857(.dina(n12866), .dinb(n12864), .dout(n13050));
  jor  g12858(.dina(n13050), .dinb(n13049), .dout(n13051));
  jand g12859(.dina(n12932), .dinb(n12929), .dout(n13052));
  jnot g12860(.din(n13052), .dout(n13053));
  jnot g12861(.din(n12929), .dout(n13054));
  jand g12862(.dina(n12931), .dinb(n13054), .dout(n13055));
  jor  g12863(.dina(n12941), .dinb(n13055), .dout(n13056));
  jand g12864(.dina(n13056), .dinb(n13053), .dout(n13057));
  jxor g12865(.dina(n13057), .dinb(n13051), .dout(n13058));
  jor  g12866(.dina(n12889), .dinb(n12881), .dout(n13059));
  jand g12867(.dina(n12889), .dinb(n12881), .dout(n13060));
  jor  g12868(.dina(n12894), .dinb(n13060), .dout(n13061));
  jand g12869(.dina(n13061), .dinb(n13059), .dout(n13062));
  jxor g12870(.dina(n13062), .dinb(n13058), .dout(n13063));
  jor  g12871(.dina(n12872), .dinb(n12868), .dout(n13064));
  jand g12872(.dina(n12895), .dinb(n12873), .dout(n13065));
  jnot g12873(.din(n13065), .dout(n13066));
  jand g12874(.dina(n13066), .dinb(n13064), .dout(n13067));
  jnot g12875(.din(n13067), .dout(n13068));
  jor  g12876(.dina(n12915), .dinb(n12907), .dout(n13069));
  jand g12877(.dina(n12916), .dinb(n12903), .dout(n13070));
  jnot g12878(.din(n13070), .dout(n13071));
  jand g12879(.dina(n13071), .dinb(n13069), .dout(n13072));
  jnot g12880(.din(n13072), .dout(n13073));
  jand g12881(.dina(n12888), .dinb(n12882), .dout(n13074));
  jor  g12882(.dina(n13074), .dinb(n12886), .dout(n13075));
  jand g12883(.dina(n12940), .dinb(n12934), .dout(n13076));
  jor  g12884(.dina(n13076), .dinb(n12938), .dout(n13077));
  jand g12885(.dina(n12924), .dinb(n12921), .dout(n13078));
  jor  g12886(.dina(n13078), .dinb(n12926), .dout(n13079));
  jxor g12887(.dina(n13079), .dinb(n13077), .dout(n13080));
  jxor g12888(.dina(n13080), .dinb(n13075), .dout(n13081));
  jand g12889(.dina(n12875), .dinb(n12701), .dout(n13082));
  jor  g12890(.dina(n13082), .dinb(n12878), .dout(n13083));
  jand g12891(.dina(n12910), .dinb(n12908), .dout(n13084));
  jor  g12892(.dina(n13084), .dinb(n12913), .dout(n13085));
  jxor g12893(.dina(n13085), .dinb(n13083), .dout(n13086));
  jand g12894(.dina(\a[60] ), .dinb(\a[32] ), .dout(n13087));
  jand g12895(.dina(\a[55] ), .dinb(\a[37] ), .dout(n13088));
  jand g12896(.dina(\a[54] ), .dinb(\a[38] ), .dout(n13089));
  jor  g12897(.dina(n13089), .dinb(n13088), .dout(n13090));
  jnot g12898(.din(n13090), .dout(n13091));
  jand g12899(.dina(\a[55] ), .dinb(\a[38] ), .dout(n13092));
  jand g12900(.dina(n13092), .dinb(n12921), .dout(n13093));
  jor  g12901(.dina(n13093), .dinb(n13091), .dout(n13094));
  jxor g12902(.dina(n13094), .dinb(n13087), .dout(n13095));
  jnot g12903(.din(n13095), .dout(n13096));
  jxor g12904(.dina(n13096), .dinb(n13086), .dout(n13097));
  jxor g12905(.dina(n13097), .dinb(n13081), .dout(n13098));
  jxor g12906(.dina(n13098), .dinb(n13073), .dout(n13099));
  jxor g12907(.dina(n13099), .dinb(n13068), .dout(n13100));
  jxor g12908(.dina(n13100), .dinb(n13063), .dout(n13101));
  jxor g12909(.dina(n13101), .dinb(n13048), .dout(n13102));
  jxor g12910(.dina(n13102), .dinb(n13045), .dout(n13103));
  jand g12911(.dina(n12974), .dinb(n12948), .dout(n13104));
  jand g12912(.dina(n12975), .dinb(n12945), .dout(n13105));
  jor  g12913(.dina(n13105), .dinb(n13104), .dout(n13106));
  jxor g12914(.dina(n13106), .dinb(n13103), .dout(n13107));
  jand g12915(.dina(n12976), .dinb(n12859), .dout(n13108));
  jor  g12916(.dina(n12976), .dinb(n12859), .dout(n13109));
  jand g12917(.dina(n12984), .dinb(n13109), .dout(n13110));
  jor  g12918(.dina(n13110), .dinb(n13108), .dout(n13111));
  jxor g12919(.dina(n13111), .dinb(n13107), .dout(\asquared[93] ));
  jand g12920(.dina(n13101), .dinb(n13048), .dout(n13113));
  jand g12921(.dina(n13102), .dinb(n13045), .dout(n13114));
  jor  g12922(.dina(n13114), .dinb(n13113), .dout(n13115));
  jand g12923(.dina(n13043), .dinb(n12991), .dout(n13116));
  jand g12924(.dina(n13044), .dinb(n12988), .dout(n13117));
  jor  g12925(.dina(n13117), .dinb(n13116), .dout(n13118));
  jand g12926(.dina(n13079), .dinb(n13077), .dout(n13119));
  jand g12927(.dina(n13080), .dinb(n13075), .dout(n13120));
  jor  g12928(.dina(n13120), .dinb(n13119), .dout(n13121));
  jnot g12929(.din(n13083), .dout(n13122));
  jnot g12930(.din(n13085), .dout(n13123));
  jand g12931(.dina(n13123), .dinb(n13122), .dout(n13124));
  jnot g12932(.din(n13124), .dout(n13125));
  jand g12933(.dina(n13085), .dinb(n13083), .dout(n13126));
  jor  g12934(.dina(n13096), .dinb(n13126), .dout(n13127));
  jand g12935(.dina(n13127), .dinb(n13125), .dout(n13128));
  jxor g12936(.dina(n13128), .dinb(n13121), .dout(n13129));
  jand g12937(.dina(n13034), .dinb(n13028), .dout(n13130));
  jnot g12938(.din(n13130), .dout(n13131));
  jnot g12939(.din(n13028), .dout(n13132));
  jnot g12940(.din(n13034), .dout(n13133));
  jand g12941(.dina(n13133), .dinb(n13132), .dout(n13134));
  jor  g12942(.dina(n13040), .dinb(n13134), .dout(n13135));
  jand g12943(.dina(n13135), .dinb(n13131), .dout(n13136));
  jxor g12944(.dina(n13136), .dinb(n13129), .dout(n13137));
  jand g12945(.dina(n13097), .dinb(n13081), .dout(n13138));
  jand g12946(.dina(n13098), .dinb(n13073), .dout(n13139));
  jor  g12947(.dina(n13139), .dinb(n13138), .dout(n13140));
  jxor g12948(.dina(n13140), .dinb(n13137), .dout(n13141));
  jor  g12949(.dina(n13017), .dinb(n13010), .dout(n13142));
  jand g12950(.dina(n13018), .dinb(n12997), .dout(n13143));
  jnot g12951(.din(n13143), .dout(n13144));
  jand g12952(.dina(n13144), .dinb(n13142), .dout(n13145));
  jnot g12953(.din(n13145), .dout(n13146));
  jand g12954(.dina(n13023), .dinb(n13020), .dout(n13147));
  jor  g12955(.dina(n13147), .dinb(n13025), .dout(n13148));
  jnot g12956(.din(n13031), .dout(n13149));
  jnot g12957(.din(n13032), .dout(n13150));
  jand g12958(.dina(n13150), .dinb(n13149), .dout(n13151));
  jnot g12959(.din(n13151), .dout(n13152));
  jand g12960(.dina(n13032), .dinb(n13031), .dout(n13153));
  jor  g12961(.dina(n13153), .dinb(n13029), .dout(n13154));
  jand g12962(.dina(n13154), .dinb(n13152), .dout(n13155));
  jxor g12963(.dina(n13155), .dinb(n13148), .dout(n13156));
  jand g12964(.dina(n13012), .dinb(n12925), .dout(n13157));
  jor  g12965(.dina(n13157), .dinb(n13015), .dout(n13158));
  jxor g12966(.dina(n13158), .dinb(n13156), .dout(n13159));
  jand g12967(.dina(n13090), .dinb(n13087), .dout(n13160));
  jor  g12968(.dina(n13160), .dinb(n13093), .dout(n13161));
  jnot g12969(.din(n11162), .dout(n13162));
  jand g12970(.dina(n13037), .dinb(n13162), .dout(n13163));
  jnot g12971(.din(n13163), .dout(n13164));
  jand g12972(.dina(n12937), .dinb(n11162), .dout(n13165));
  jor  g12973(.dina(n13165), .dinb(n13036), .dout(n13166));
  jand g12974(.dina(n13166), .dinb(n13164), .dout(n13167));
  jxor g12975(.dina(n13167), .dinb(n13161), .dout(n13168));
  jand g12976(.dina(n13008), .dinb(n13001), .dout(n13169));
  jor  g12977(.dina(n13169), .dinb(n13006), .dout(n13170));
  jxor g12978(.dina(n13170), .dinb(n13168), .dout(n13171));
  jxor g12979(.dina(n13171), .dinb(n13159), .dout(n13172));
  jxor g12980(.dina(n13172), .dinb(n13146), .dout(n13173));
  jxor g12981(.dina(n13173), .dinb(n13141), .dout(n13174));
  jxor g12982(.dina(n13174), .dinb(n13118), .dout(n13175));
  jand g12983(.dina(n13099), .dinb(n13068), .dout(n13176));
  jand g12984(.dina(n13100), .dinb(n13063), .dout(n13177));
  jor  g12985(.dina(n13177), .dinb(n13176), .dout(n13178));
  jand g12986(.dina(n13041), .dinb(n13019), .dout(n13179));
  jand g12987(.dina(n13042), .dinb(n12994), .dout(n13180));
  jor  g12988(.dina(n13180), .dinb(n13179), .dout(n13181));
  jand g12989(.dina(n13057), .dinb(n13051), .dout(n13182));
  jand g12990(.dina(n13062), .dinb(n13058), .dout(n13183));
  jor  g12991(.dina(n13183), .dinb(n13182), .dout(n13184));
  jand g12992(.dina(\a[59] ), .dinb(\a[34] ), .dout(n13185));
  jand g12993(.dina(\a[53] ), .dinb(\a[40] ), .dout(n13186));
  jor  g12994(.dina(n13186), .dinb(n13014), .dout(n13187));
  jnot g12995(.din(n13187), .dout(n13188));
  jand g12996(.dina(\a[53] ), .dinb(\a[41] ), .dout(n13189));
  jand g12997(.dina(n13189), .dinb(n13011), .dout(n13190));
  jor  g12998(.dina(n13190), .dinb(n13188), .dout(n13191));
  jxor g12999(.dina(n13191), .dinb(n13185), .dout(n13192));
  jnot g13000(.din(n13192), .dout(n13193));
  jand g13001(.dina(\a[63] ), .dinb(\a[30] ), .dout(n13194));
  jand g13002(.dina(\a[61] ), .dinb(\a[32] ), .dout(n13195));
  jand g13003(.dina(\a[60] ), .dinb(\a[33] ), .dout(n13196));
  jor  g13004(.dina(n13196), .dinb(n13195), .dout(n13197));
  jand g13005(.dina(\a[61] ), .dinb(\a[33] ), .dout(n13198));
  jand g13006(.dina(n13198), .dinb(n13087), .dout(n13199));
  jnot g13007(.din(n13199), .dout(n13200));
  jand g13008(.dina(n13200), .dinb(n13197), .dout(n13201));
  jxor g13009(.dina(n13201), .dinb(n13194), .dout(n13202));
  jnot g13010(.din(n13202), .dout(n13203));
  jand g13011(.dina(\a[58] ), .dinb(\a[35] ), .dout(n13204));
  jand g13012(.dina(\a[54] ), .dinb(\a[39] ), .dout(n13205));
  jor  g13013(.dina(n13205), .dinb(n12912), .dout(n13206));
  jnot g13014(.din(n13206), .dout(n13207));
  jand g13015(.dina(\a[57] ), .dinb(\a[39] ), .dout(n13208));
  jand g13016(.dina(n13208), .dinb(n12782), .dout(n13209));
  jor  g13017(.dina(n13209), .dinb(n13207), .dout(n13210));
  jxor g13018(.dina(n13210), .dinb(n13204), .dout(n13211));
  jxor g13019(.dina(n13211), .dinb(n13203), .dout(n13212));
  jxor g13020(.dina(n13212), .dinb(n13193), .dout(n13213));
  jand g13021(.dina(\a[51] ), .dinb(\a[42] ), .dout(n13214));
  jand g13022(.dina(\a[49] ), .dinb(\a[44] ), .dout(n13215));
  jnot g13023(.din(n13215), .dout(n13216));
  jand g13024(.dina(\a[50] ), .dinb(\a[43] ), .dout(n13217));
  jnot g13025(.din(n13217), .dout(n13218));
  jand g13026(.dina(n13218), .dinb(n13216), .dout(n13219));
  jand g13027(.dina(\a[50] ), .dinb(\a[44] ), .dout(n13220));
  jand g13028(.dina(n13220), .dinb(n13020), .dout(n13221));
  jor  g13029(.dina(n13221), .dinb(n13219), .dout(n13222));
  jxor g13030(.dina(n13222), .dinb(n13214), .dout(n13223));
  jnot g13031(.din(n13223), .dout(n13224));
  jand g13032(.dina(\a[56] ), .dinb(\a[37] ), .dout(n13225));
  jor  g13033(.dina(n13092), .dinb(n13024), .dout(n13226));
  jand g13034(.dina(\a[55] ), .dinb(\a[45] ), .dout(n13227));
  jand g13035(.dina(n13227), .dinb(n12038), .dout(n13228));
  jnot g13036(.din(n13228), .dout(n13229));
  jand g13037(.dina(n13229), .dinb(n13226), .dout(n13230));
  jxor g13038(.dina(n13230), .dinb(n13225), .dout(n13231));
  jxor g13039(.dina(n13231), .dinb(n13224), .dout(n13232));
  jnot g13040(.din(n13005), .dout(n13233));
  jand g13041(.dina(\a[47] ), .dinb(n12998), .dout(n13234));
  jxor g13042(.dina(n13234), .dinb(n13233), .dout(n13235));
  jnot g13043(.din(n13235), .dout(n13236));
  jxor g13044(.dina(n13236), .dinb(n13232), .dout(n13237));
  jxor g13045(.dina(n13237), .dinb(n13213), .dout(n13238));
  jxor g13046(.dina(n13238), .dinb(n13184), .dout(n13239));
  jxor g13047(.dina(n13239), .dinb(n13181), .dout(n13240));
  jxor g13048(.dina(n13240), .dinb(n13178), .dout(n13241));
  jxor g13049(.dina(n13241), .dinb(n13175), .dout(n13242));
  jxor g13050(.dina(n13242), .dinb(n13115), .dout(n13243));
  jand g13051(.dina(n13106), .dinb(n13103), .dout(n13244));
  jnot g13052(.din(n13103), .dout(n13245));
  jnot g13053(.din(n13106), .dout(n13246));
  jand g13054(.dina(n13246), .dinb(n13245), .dout(n13247));
  jnot g13055(.din(n13247), .dout(n13248));
  jand g13056(.dina(n13111), .dinb(n13248), .dout(n13249));
  jor  g13057(.dina(n13249), .dinb(n13244), .dout(n13250));
  jxor g13058(.dina(n13250), .dinb(n13243), .dout(\asquared[94] ));
  jand g13059(.dina(n13239), .dinb(n13181), .dout(n13252));
  jand g13060(.dina(n13240), .dinb(n13178), .dout(n13253));
  jor  g13061(.dina(n13253), .dinb(n13252), .dout(n13254));
  jand g13062(.dina(n13237), .dinb(n13213), .dout(n13255));
  jand g13063(.dina(n13238), .dinb(n13184), .dout(n13256));
  jor  g13064(.dina(n13256), .dinb(n13255), .dout(n13257));
  jand g13065(.dina(n13167), .dinb(n13161), .dout(n13258));
  jand g13066(.dina(n13170), .dinb(n13168), .dout(n13259));
  jor  g13067(.dina(n13259), .dinb(n13258), .dout(n13260));
  jand g13068(.dina(n13155), .dinb(n13148), .dout(n13261));
  jand g13069(.dina(n13158), .dinb(n13156), .dout(n13262));
  jor  g13070(.dina(n13262), .dinb(n13261), .dout(n13263));
  jxor g13071(.dina(n13263), .dinb(n13260), .dout(n13264));
  jnot g13072(.din(n13264), .dout(n13265));
  jor  g13073(.dina(n13211), .dinb(n13203), .dout(n13266));
  jand g13074(.dina(n13212), .dinb(n13193), .dout(n13267));
  jnot g13075(.din(n13267), .dout(n13268));
  jand g13076(.dina(n13268), .dinb(n13266), .dout(n13269));
  jxor g13077(.dina(n13269), .dinb(n13265), .dout(n13270));
  jand g13078(.dina(n13171), .dinb(n13159), .dout(n13271));
  jand g13079(.dina(n13172), .dinb(n13146), .dout(n13272));
  jor  g13080(.dina(n13272), .dinb(n13271), .dout(n13273));
  jxor g13081(.dina(n13273), .dinb(n13270), .dout(n13274));
  jxor g13082(.dina(n13274), .dinb(n13257), .dout(n13275));
  jxor g13083(.dina(n13275), .dinb(n13254), .dout(n13276));
  jand g13084(.dina(n13140), .dinb(n13137), .dout(n13277));
  jand g13085(.dina(n13173), .dinb(n13141), .dout(n13278));
  jor  g13086(.dina(n13278), .dinb(n13277), .dout(n13279));
  jand g13087(.dina(n13230), .dinb(n13225), .dout(n13280));
  jor  g13088(.dina(n13280), .dinb(n13228), .dout(n13281));
  jnot g13089(.din(\a[47] ), .dout(n13282));
  jand g13090(.dina(n13233), .dinb(n12998), .dout(n13283));
  jor  g13091(.dina(n13283), .dinb(n13282), .dout(n13284));
  jnot g13092(.din(n13284), .dout(n13285));
  jxor g13093(.dina(n13285), .dinb(n10725), .dout(n13286));
  jxor g13094(.dina(n13286), .dinb(n13281), .dout(n13287));
  jor  g13095(.dina(n13231), .dinb(n13224), .dout(n13288));
  jand g13096(.dina(n13231), .dinb(n13224), .dout(n13289));
  jor  g13097(.dina(n13236), .dinb(n13289), .dout(n13290));
  jand g13098(.dina(n13290), .dinb(n13288), .dout(n13291));
  jxor g13099(.dina(n13291), .dinb(n13287), .dout(n13292));
  jand g13100(.dina(n13201), .dinb(n13194), .dout(n13293));
  jor  g13101(.dina(n13293), .dinb(n13199), .dout(n13294));
  jand g13102(.dina(n13206), .dinb(n13204), .dout(n13295));
  jor  g13103(.dina(n13295), .dinb(n13209), .dout(n13296));
  jxor g13104(.dina(n13296), .dinb(n13294), .dout(n13297));
  jand g13105(.dina(n13187), .dinb(n13185), .dout(n13298));
  jor  g13106(.dina(n13298), .dinb(n13190), .dout(n13299));
  jxor g13107(.dina(n13299), .dinb(n13297), .dout(n13300));
  jxor g13108(.dina(n13300), .dinb(n13292), .dout(n13301));
  jxor g13109(.dina(n13301), .dinb(n13279), .dout(n13302));
  jand g13110(.dina(n13128), .dinb(n13121), .dout(n13303));
  jand g13111(.dina(n13136), .dinb(n13129), .dout(n13304));
  jor  g13112(.dina(n13304), .dinb(n13303), .dout(n13305));
  jand g13113(.dina(\a[54] ), .dinb(\a[40] ), .dout(n13306));
  jand g13114(.dina(\a[52] ), .dinb(\a[42] ), .dout(n13307));
  jor  g13115(.dina(n13307), .dinb(n13189), .dout(n13308));
  jnot g13116(.din(n13308), .dout(n13309));
  jand g13117(.dina(\a[53] ), .dinb(\a[42] ), .dout(n13310));
  jand g13118(.dina(n13310), .dinb(n13014), .dout(n13311));
  jor  g13119(.dina(n13311), .dinb(n13309), .dout(n13312));
  jxor g13120(.dina(n13312), .dinb(n13306), .dout(n13313));
  jnot g13121(.din(n13313), .dout(n13314));
  jand g13122(.dina(\a[58] ), .dinb(\a[36] ), .dout(n13315));
  jand g13123(.dina(\a[51] ), .dinb(\a[43] ), .dout(n13316));
  jor  g13124(.dina(n13316), .dinb(n13220), .dout(n13317));
  jand g13125(.dina(\a[51] ), .dinb(\a[44] ), .dout(n13318));
  jand g13126(.dina(n13318), .dinb(n13217), .dout(n13319));
  jnot g13127(.din(n13319), .dout(n13320));
  jand g13128(.dina(n13320), .dinb(n13317), .dout(n13321));
  jxor g13129(.dina(n13321), .dinb(n13315), .dout(n13322));
  jxor g13130(.dina(n13322), .dinb(n13314), .dout(n13323));
  jnot g13131(.din(n13323), .dout(n13324));
  jand g13132(.dina(\a[49] ), .dinb(\a[45] ), .dout(n13325));
  jand g13133(.dina(\a[48] ), .dinb(\a[46] ), .dout(n13326));
  jnot g13134(.din(n13326), .dout(n13327));
  jand g13135(.dina(\a[56] ), .dinb(\a[38] ), .dout(n13328));
  jxor g13136(.dina(n13328), .dinb(n13327), .dout(n13329));
  jxor g13137(.dina(n13329), .dinb(n13325), .dout(n13330));
  jxor g13138(.dina(n13330), .dinb(n13324), .dout(n13331));
  jxor g13139(.dina(n13331), .dinb(n13305), .dout(n13332));
  jand g13140(.dina(\a[57] ), .dinb(\a[37] ), .dout(n13333));
  jnot g13141(.din(n13333), .dout(n13334));
  jand g13142(.dina(\a[60] ), .dinb(\a[34] ), .dout(n13335));
  jand g13143(.dina(\a[55] ), .dinb(\a[39] ), .dout(n13336));
  jxor g13144(.dina(n13336), .dinb(n13335), .dout(n13337));
  jxor g13145(.dina(n13337), .dinb(n13334), .dout(n13338));
  jnot g13146(.din(n13338), .dout(n13339));
  jand g13147(.dina(\a[62] ), .dinb(\a[32] ), .dout(n13340));
  jand g13148(.dina(\a[59] ), .dinb(\a[35] ), .dout(n13341));
  jor  g13149(.dina(n13341), .dinb(n13198), .dout(n13342));
  jnot g13150(.din(n13342), .dout(n13343));
  jand g13151(.dina(\a[61] ), .dinb(\a[35] ), .dout(n13344));
  jand g13152(.dina(n13344), .dinb(n12937), .dout(n13345));
  jor  g13153(.dina(n13345), .dinb(n13343), .dout(n13346));
  jxor g13154(.dina(n13346), .dinb(n13340), .dout(n13347));
  jnot g13155(.din(n13347), .dout(n13348));
  jnot g13156(.din(n13219), .dout(n13349));
  jand g13157(.dina(n13349), .dinb(n13214), .dout(n13350));
  jor  g13158(.dina(n13350), .dinb(n13221), .dout(n13351));
  jxor g13159(.dina(n13351), .dinb(n13348), .dout(n13352));
  jxor g13160(.dina(n13352), .dinb(n13339), .dout(n13353));
  jxor g13161(.dina(n13353), .dinb(n13332), .dout(n13354));
  jxor g13162(.dina(n13354), .dinb(n13302), .dout(n13355));
  jxor g13163(.dina(n13355), .dinb(n13276), .dout(n13356));
  jand g13164(.dina(n13174), .dinb(n13118), .dout(n13357));
  jand g13165(.dina(n13241), .dinb(n13175), .dout(n13358));
  jor  g13166(.dina(n13358), .dinb(n13357), .dout(n13359));
  jxor g13167(.dina(n13359), .dinb(n13356), .dout(n13360));
  jand g13168(.dina(n13242), .dinb(n13115), .dout(n13361));
  jor  g13169(.dina(n13242), .dinb(n13115), .dout(n13362));
  jand g13170(.dina(n13250), .dinb(n13362), .dout(n13363));
  jor  g13171(.dina(n13363), .dinb(n13361), .dout(n13364));
  jxor g13172(.dina(n13364), .dinb(n13360), .dout(\asquared[95] ));
  jand g13173(.dina(n13275), .dinb(n13254), .dout(n13366));
  jand g13174(.dina(n13355), .dinb(n13276), .dout(n13367));
  jor  g13175(.dina(n13367), .dinb(n13366), .dout(n13368));
  jand g13176(.dina(n13301), .dinb(n13279), .dout(n13369));
  jand g13177(.dina(n13354), .dinb(n13302), .dout(n13370));
  jor  g13178(.dina(n13370), .dinb(n13369), .dout(n13371));
  jand g13179(.dina(n13331), .dinb(n13305), .dout(n13372));
  jand g13180(.dina(n13353), .dinb(n13332), .dout(n13373));
  jor  g13181(.dina(n13373), .dinb(n13372), .dout(n13374));
  jand g13182(.dina(n13285), .dinb(n10725), .dout(n13375));
  jand g13183(.dina(n13286), .dinb(n13281), .dout(n13376));
  jor  g13184(.dina(n13376), .dinb(n13375), .dout(n13377));
  jand g13185(.dina(\a[59] ), .dinb(\a[36] ), .dout(n13378));
  jand g13186(.dina(\a[60] ), .dinb(\a[35] ), .dout(n13379));
  jor  g13187(.dina(n13379), .dinb(n13378), .dout(n13380));
  jand g13188(.dina(\a[60] ), .dinb(\a[36] ), .dout(n13381));
  jand g13189(.dina(n13381), .dinb(n13341), .dout(n13382));
  jnot g13190(.din(n13382), .dout(n13383));
  jand g13191(.dina(n13383), .dinb(n13380), .dout(n13384));
  jnot g13192(.din(n13328), .dout(n13385));
  jand g13193(.dina(n13385), .dinb(n13327), .dout(n13386));
  jnot g13194(.din(n13386), .dout(n13387));
  jand g13195(.dina(n13328), .dinb(n13326), .dout(n13388));
  jor  g13196(.dina(n13388), .dinb(n13325), .dout(n13389));
  jand g13197(.dina(n13389), .dinb(n13387), .dout(n13390));
  jxor g13198(.dina(n13390), .dinb(n13384), .dout(n13391));
  jxor g13199(.dina(n13391), .dinb(n13377), .dout(n13392));
  jand g13200(.dina(n13296), .dinb(n13294), .dout(n13393));
  jand g13201(.dina(n13299), .dinb(n13297), .dout(n13394));
  jor  g13202(.dina(n13394), .dinb(n13393), .dout(n13395));
  jxor g13203(.dina(n13395), .dinb(n13392), .dout(n13396));
  jand g13204(.dina(n13291), .dinb(n13287), .dout(n13397));
  jand g13205(.dina(n13300), .dinb(n13292), .dout(n13398));
  jor  g13206(.dina(n13398), .dinb(n13397), .dout(n13399));
  jxor g13207(.dina(n13399), .dinb(n13396), .dout(n13400));
  jxor g13208(.dina(n13400), .dinb(n13374), .dout(n13401));
  jxor g13209(.dina(n13401), .dinb(n13371), .dout(n13402));
  jand g13210(.dina(n13273), .dinb(n13270), .dout(n13403));
  jand g13211(.dina(n13274), .dinb(n13257), .dout(n13404));
  jor  g13212(.dina(n13404), .dinb(n13403), .dout(n13405));
  jand g13213(.dina(n13342), .dinb(n13340), .dout(n13406));
  jor  g13214(.dina(n13406), .dinb(n13345), .dout(n13407));
  jand g13215(.dina(n13336), .dinb(n13335), .dout(n13408));
  jnot g13216(.din(n13408), .dout(n13409));
  jnot g13217(.din(n13335), .dout(n13410));
  jnot g13218(.din(n13336), .dout(n13411));
  jand g13219(.dina(n13411), .dinb(n13410), .dout(n13412));
  jor  g13220(.dina(n13412), .dinb(n13334), .dout(n13413));
  jand g13221(.dina(n13413), .dinb(n13409), .dout(n13414));
  jnot g13222(.din(n13414), .dout(n13415));
  jxor g13223(.dina(n13415), .dinb(n13407), .dout(n13416));
  jand g13224(.dina(n13308), .dinb(n13306), .dout(n13417));
  jor  g13225(.dina(n13417), .dinb(n13311), .dout(n13418));
  jxor g13226(.dina(n13418), .dinb(n13416), .dout(n13419));
  jand g13227(.dina(n13322), .dinb(n13314), .dout(n13420));
  jnot g13228(.din(n13420), .dout(n13421));
  jor  g13229(.dina(n13330), .dinb(n13324), .dout(n13422));
  jand g13230(.dina(n13422), .dinb(n13421), .dout(n13423));
  jnot g13231(.din(n13423), .dout(n13424));
  jand g13232(.dina(n13351), .dinb(n13348), .dout(n13425));
  jand g13233(.dina(n13352), .dinb(n13339), .dout(n13426));
  jor  g13234(.dina(n13426), .dinb(n13425), .dout(n13427));
  jxor g13235(.dina(n13427), .dinb(n13424), .dout(n13428));
  jxor g13236(.dina(n13428), .dinb(n13419), .dout(n13429));
  jxor g13237(.dina(n13429), .dinb(n13405), .dout(n13430));
  jand g13238(.dina(n13263), .dinb(n13260), .dout(n13431));
  jnot g13239(.din(n13431), .dout(n13432));
  jor  g13240(.dina(n13269), .dinb(n13265), .dout(n13433));
  jand g13241(.dina(n13433), .dinb(n13432), .dout(n13434));
  jnot g13242(.din(n13310), .dout(n13435));
  jand g13243(.dina(\a[52] ), .dinb(\a[43] ), .dout(n13436));
  jor  g13244(.dina(n13436), .dinb(n13318), .dout(n13437));
  jand g13245(.dina(\a[52] ), .dinb(\a[44] ), .dout(n13438));
  jand g13246(.dina(n13438), .dinb(n13316), .dout(n13439));
  jnot g13247(.din(n13439), .dout(n13440));
  jand g13248(.dina(n13440), .dinb(n13437), .dout(n13441));
  jxor g13249(.dina(n13441), .dinb(n13435), .dout(n13442));
  jnot g13250(.din(n13442), .dout(n13443));
  jand g13251(.dina(\a[56] ), .dinb(\a[39] ), .dout(n13444));
  jnot g13252(.din(n13444), .dout(n13445));
  jand g13253(.dina(\a[50] ), .dinb(\a[45] ), .dout(n13446));
  jand g13254(.dina(\a[49] ), .dinb(\a[46] ), .dout(n13447));
  jor  g13255(.dina(n13447), .dinb(n13446), .dout(n13448));
  jand g13256(.dina(\a[50] ), .dinb(\a[46] ), .dout(n13449));
  jand g13257(.dina(n13449), .dinb(n13325), .dout(n13450));
  jnot g13258(.din(n13450), .dout(n13451));
  jand g13259(.dina(n13451), .dinb(n13448), .dout(n13452));
  jxor g13260(.dina(n13452), .dinb(n13445), .dout(n13453));
  jand g13261(.dina(\a[62] ), .dinb(\a[33] ), .dout(n13454));
  jnot g13262(.din(n13454), .dout(n13455));
  jand g13263(.dina(\a[48] ), .dinb(n13282), .dout(n13456));
  jxor g13264(.dina(n13456), .dinb(n13455), .dout(n13457));
  jxor g13265(.dina(n13457), .dinb(n13453), .dout(n13458));
  jxor g13266(.dina(n13458), .dinb(n13443), .dout(n13459));
  jnot g13267(.din(n13459), .dout(n13460));
  jxor g13268(.dina(n13460), .dinb(n13434), .dout(n13461));
  jand g13269(.dina(n13321), .dinb(n13315), .dout(n13462));
  jor  g13270(.dina(n13462), .dinb(n13319), .dout(n13463));
  jand g13271(.dina(\a[58] ), .dinb(\a[37] ), .dout(n13464));
  jnot g13272(.din(n13464), .dout(n13465));
  jand g13273(.dina(\a[57] ), .dinb(\a[38] ), .dout(n13466));
  jand g13274(.dina(\a[55] ), .dinb(\a[40] ), .dout(n13467));
  jor  g13275(.dina(n13467), .dinb(n13466), .dout(n13468));
  jand g13276(.dina(\a[57] ), .dinb(\a[40] ), .dout(n13469));
  jand g13277(.dina(n13469), .dinb(n13092), .dout(n13470));
  jnot g13278(.din(n13470), .dout(n13471));
  jand g13279(.dina(n13471), .dinb(n13468), .dout(n13472));
  jxor g13280(.dina(n13472), .dinb(n13465), .dout(n13473));
  jnot g13281(.din(n13473), .dout(n13474));
  jxor g13282(.dina(n13474), .dinb(n13463), .dout(n13475));
  jand g13283(.dina(\a[54] ), .dinb(\a[41] ), .dout(n13476));
  jand g13284(.dina(\a[63] ), .dinb(\a[32] ), .dout(n13477));
  jand g13285(.dina(\a[61] ), .dinb(\a[34] ), .dout(n13478));
  jor  g13286(.dina(n13478), .dinb(n13477), .dout(n13479));
  jand g13287(.dina(\a[63] ), .dinb(\a[34] ), .dout(n13480));
  jand g13288(.dina(n13480), .dinb(n13195), .dout(n13481));
  jnot g13289(.din(n13481), .dout(n13482));
  jand g13290(.dina(n13482), .dinb(n13479), .dout(n13483));
  jxor g13291(.dina(n13483), .dinb(n13476), .dout(n13484));
  jxor g13292(.dina(n13484), .dinb(n13475), .dout(n13485));
  jxor g13293(.dina(n13485), .dinb(n13461), .dout(n13486));
  jxor g13294(.dina(n13486), .dinb(n13430), .dout(n13487));
  jxor g13295(.dina(n13487), .dinb(n13402), .dout(n13488));
  jxor g13296(.dina(n13488), .dinb(n13368), .dout(n13489));
  jand g13297(.dina(n13359), .dinb(n13356), .dout(n13490));
  jnot g13298(.din(n13356), .dout(n13491));
  jnot g13299(.din(n13359), .dout(n13492));
  jand g13300(.dina(n13492), .dinb(n13491), .dout(n13493));
  jnot g13301(.din(n13493), .dout(n13494));
  jand g13302(.dina(n13364), .dinb(n13494), .dout(n13495));
  jor  g13303(.dina(n13495), .dinb(n13490), .dout(n13496));
  jxor g13304(.dina(n13496), .dinb(n13489), .dout(\asquared[96] ));
  jand g13305(.dina(n13401), .dinb(n13371), .dout(n13498));
  jand g13306(.dina(n13487), .dinb(n13402), .dout(n13499));
  jor  g13307(.dina(n13499), .dinb(n13498), .dout(n13500));
  jand g13308(.dina(n13399), .dinb(n13396), .dout(n13501));
  jand g13309(.dina(n13400), .dinb(n13374), .dout(n13502));
  jor  g13310(.dina(n13502), .dinb(n13501), .dout(n13503));
  jand g13311(.dina(n13448), .dinb(n13444), .dout(n13504));
  jor  g13312(.dina(n13504), .dinb(n13450), .dout(n13505));
  jand g13313(.dina(n13455), .dinb(n13282), .dout(n13506));
  jor  g13314(.dina(n13506), .dinb(n4774), .dout(n13507));
  jnot g13315(.din(n13507), .dout(n13508));
  jxor g13316(.dina(n13508), .dinb(n13505), .dout(n13509));
  jand g13317(.dina(n13437), .dinb(n13310), .dout(n13510));
  jor  g13318(.dina(n13510), .dinb(n13439), .dout(n13511));
  jxor g13319(.dina(n13511), .dinb(n13509), .dout(n13512));
  jnot g13320(.din(n13453), .dout(n13513));
  jnot g13321(.din(n13457), .dout(n13514));
  jand g13322(.dina(n13514), .dinb(n13513), .dout(n13515));
  jnot g13323(.din(n13515), .dout(n13516));
  jand g13324(.dina(n13457), .dinb(n13453), .dout(n13517));
  jor  g13325(.dina(n13517), .dinb(n13442), .dout(n13518));
  jand g13326(.dina(n13518), .dinb(n13516), .dout(n13519));
  jnot g13327(.din(n13519), .dout(n13520));
  jnot g13328(.din(n13463), .dout(n13521));
  jand g13329(.dina(n13473), .dinb(n13521), .dout(n13522));
  jnot g13330(.din(n13522), .dout(n13523));
  jand g13331(.dina(n13474), .dinb(n13463), .dout(n13524));
  jor  g13332(.dina(n13484), .dinb(n13524), .dout(n13525));
  jand g13333(.dina(n13525), .dinb(n13523), .dout(n13526));
  jxor g13334(.dina(n13526), .dinb(n13520), .dout(n13527));
  jxor g13335(.dina(n13527), .dinb(n13512), .dout(n13528));
  jxor g13336(.dina(n13528), .dinb(n13503), .dout(n13529));
  jand g13337(.dina(n13415), .dinb(n13407), .dout(n13530));
  jand g13338(.dina(n13418), .dinb(n13416), .dout(n13531));
  jor  g13339(.dina(n13531), .dinb(n13530), .dout(n13532));
  jand g13340(.dina(\a[55] ), .dinb(\a[41] ), .dout(n13533));
  jand g13341(.dina(\a[53] ), .dinb(\a[43] ), .dout(n13534));
  jand g13342(.dina(n13534), .dinb(n13533), .dout(n13535));
  jand g13343(.dina(\a[55] ), .dinb(\a[42] ), .dout(n13536));
  jand g13344(.dina(n13536), .dinb(n13476), .dout(n13537));
  jor  g13345(.dina(n13537), .dinb(n13535), .dout(n13538));
  jand g13346(.dina(\a[54] ), .dinb(\a[43] ), .dout(n13539));
  jand g13347(.dina(n13539), .dinb(n13310), .dout(n13540));
  jnot g13348(.din(n13540), .dout(n13541));
  jand g13349(.dina(n13541), .dinb(n13538), .dout(n13542));
  jnot g13350(.din(n13542), .dout(n13543));
  jand g13351(.dina(\a[54] ), .dinb(\a[42] ), .dout(n13544));
  jor  g13352(.dina(n13544), .dinb(n13534), .dout(n13545));
  jand g13353(.dina(n13545), .dinb(n13541), .dout(n13546));
  jor  g13354(.dina(n13546), .dinb(n13533), .dout(n13547));
  jand g13355(.dina(n13547), .dinb(n13543), .dout(n13548));
  jand g13356(.dina(\a[63] ), .dinb(\a[33] ), .dout(n13549));
  jand g13357(.dina(\a[62] ), .dinb(\a[34] ), .dout(n13550));
  jor  g13358(.dina(n13550), .dinb(n13344), .dout(n13551));
  jand g13359(.dina(\a[62] ), .dinb(\a[35] ), .dout(n13552));
  jand g13360(.dina(n13552), .dinb(n13478), .dout(n13553));
  jnot g13361(.din(n13553), .dout(n13554));
  jand g13362(.dina(n13554), .dinb(n13551), .dout(n13555));
  jxor g13363(.dina(n13555), .dinb(n13549), .dout(n13556));
  jxor g13364(.dina(n13556), .dinb(n13548), .dout(n13557));
  jxor g13365(.dina(n13557), .dinb(n13532), .dout(n13558));
  jand g13366(.dina(n13483), .dinb(n13476), .dout(n13559));
  jor  g13367(.dina(n13559), .dinb(n13481), .dout(n13560));
  jand g13368(.dina(n13468), .dinb(n13464), .dout(n13561));
  jor  g13369(.dina(n13561), .dinb(n13470), .dout(n13562));
  jxor g13370(.dina(n13562), .dinb(n13560), .dout(n13563));
  jand g13371(.dina(n13390), .dinb(n13384), .dout(n13564));
  jor  g13372(.dina(n13564), .dinb(n13382), .dout(n13565));
  jxor g13373(.dina(n13565), .dinb(n13563), .dout(n13566));
  jand g13374(.dina(n13391), .dinb(n13377), .dout(n13567));
  jand g13375(.dina(n13395), .dinb(n13392), .dout(n13568));
  jor  g13376(.dina(n13568), .dinb(n13567), .dout(n13569));
  jxor g13377(.dina(n13569), .dinb(n13566), .dout(n13570));
  jxor g13378(.dina(n13570), .dinb(n13558), .dout(n13571));
  jxor g13379(.dina(n13571), .dinb(n13529), .dout(n13572));
  jand g13380(.dina(n13429), .dinb(n13405), .dout(n13573));
  jand g13381(.dina(n13486), .dinb(n13430), .dout(n13574));
  jor  g13382(.dina(n13574), .dinb(n13573), .dout(n13575));
  jand g13383(.dina(n13427), .dinb(n13424), .dout(n13576));
  jand g13384(.dina(n13428), .dinb(n13419), .dout(n13577));
  jor  g13385(.dina(n13577), .dinb(n13576), .dout(n13578));
  jand g13386(.dina(\a[51] ), .dinb(\a[45] ), .dout(n13579));
  jand g13387(.dina(\a[49] ), .dinb(\a[47] ), .dout(n13580));
  jor  g13388(.dina(n13580), .dinb(n13449), .dout(n13581));
  jnot g13389(.din(n13581), .dout(n13582));
  jand g13390(.dina(\a[50] ), .dinb(\a[47] ), .dout(n13583));
  jand g13391(.dina(n13583), .dinb(n13447), .dout(n13584));
  jor  g13392(.dina(n13584), .dinb(n13582), .dout(n13585));
  jxor g13393(.dina(n13585), .dinb(n13579), .dout(n13586));
  jand g13394(.dina(\a[58] ), .dinb(\a[38] ), .dout(n13587));
  jor  g13395(.dina(n13587), .dinb(n13208), .dout(n13588));
  jnot g13396(.din(n13588), .dout(n13589));
  jand g13397(.dina(\a[58] ), .dinb(\a[39] ), .dout(n13590));
  jand g13398(.dina(n13590), .dinb(n13466), .dout(n13591));
  jor  g13399(.dina(n13591), .dinb(n13589), .dout(n13592));
  jxor g13400(.dina(n13592), .dinb(n13438), .dout(n13593));
  jand g13401(.dina(\a[59] ), .dinb(\a[37] ), .dout(n13594));
  jand g13402(.dina(\a[56] ), .dinb(\a[40] ), .dout(n13595));
  jor  g13403(.dina(n13595), .dinb(n13594), .dout(n13596));
  jand g13404(.dina(\a[59] ), .dinb(\a[40] ), .dout(n13597));
  jand g13405(.dina(n13597), .dinb(n13225), .dout(n13598));
  jnot g13406(.din(n13598), .dout(n13599));
  jand g13407(.dina(n13599), .dinb(n13596), .dout(n13600));
  jxor g13408(.dina(n13600), .dinb(n13381), .dout(n13601));
  jxor g13409(.dina(n13601), .dinb(n13593), .dout(n13602));
  jxor g13410(.dina(n13602), .dinb(n13586), .dout(n13603));
  jxor g13411(.dina(n13603), .dinb(n13578), .dout(n13604));
  jand g13412(.dina(n13460), .dinb(n13434), .dout(n13605));
  jnot g13413(.din(n13605), .dout(n13606));
  jnot g13414(.din(n13434), .dout(n13607));
  jand g13415(.dina(n13459), .dinb(n13607), .dout(n13608));
  jor  g13416(.dina(n13485), .dinb(n13608), .dout(n13609));
  jand g13417(.dina(n13609), .dinb(n13606), .dout(n13610));
  jxor g13418(.dina(n13610), .dinb(n13604), .dout(n13611));
  jxor g13419(.dina(n13611), .dinb(n13575), .dout(n13612));
  jxor g13420(.dina(n13612), .dinb(n13572), .dout(n13613));
  jxor g13421(.dina(n13613), .dinb(n13500), .dout(n13614));
  jand g13422(.dina(n13488), .dinb(n13368), .dout(n13615));
  jor  g13423(.dina(n13488), .dinb(n13368), .dout(n13616));
  jand g13424(.dina(n13496), .dinb(n13616), .dout(n13617));
  jor  g13425(.dina(n13617), .dinb(n13615), .dout(n13618));
  jxor g13426(.dina(n13618), .dinb(n13614), .dout(\asquared[97] ));
  jand g13427(.dina(n13611), .dinb(n13575), .dout(n13620));
  jand g13428(.dina(n13612), .dinb(n13572), .dout(n13621));
  jor  g13429(.dina(n13621), .dinb(n13620), .dout(n13622));
  jand g13430(.dina(n13603), .dinb(n13578), .dout(n13623));
  jand g13431(.dina(n13610), .dinb(n13604), .dout(n13624));
  jor  g13432(.dina(n13624), .dinb(n13623), .dout(n13625));
  jand g13433(.dina(\a[61] ), .dinb(\a[36] ), .dout(n13626));
  jand g13434(.dina(n13581), .dinb(n13579), .dout(n13627));
  jor  g13435(.dina(n13627), .dinb(n13584), .dout(n13628));
  jxor g13436(.dina(n13628), .dinb(n13626), .dout(n13629));
  jand g13437(.dina(n13588), .dinb(n13438), .dout(n13630));
  jor  g13438(.dina(n13630), .dinb(n13591), .dout(n13631));
  jxor g13439(.dina(n13631), .dinb(n13629), .dout(n13632));
  jand g13440(.dina(n13562), .dinb(n13560), .dout(n13633));
  jand g13441(.dina(n13565), .dinb(n13563), .dout(n13634));
  jor  g13442(.dina(n13634), .dinb(n13633), .dout(n13635));
  jnot g13443(.din(n13593), .dout(n13636));
  jor  g13444(.dina(n13601), .dinb(n13636), .dout(n13637));
  jnot g13445(.din(n13586), .dout(n13638));
  jand g13446(.dina(n13601), .dinb(n13636), .dout(n13639));
  jor  g13447(.dina(n13639), .dinb(n13638), .dout(n13640));
  jand g13448(.dina(n13640), .dinb(n13637), .dout(n13641));
  jxor g13449(.dina(n13641), .dinb(n13635), .dout(n13642));
  jxor g13450(.dina(n13642), .dinb(n13632), .dout(n13643));
  jand g13451(.dina(n13508), .dinb(n13505), .dout(n13644));
  jand g13452(.dina(n13511), .dinb(n13509), .dout(n13645));
  jor  g13453(.dina(n13645), .dinb(n13644), .dout(n13646));
  jand g13454(.dina(\a[51] ), .dinb(\a[46] ), .dout(n13647));
  jor  g13455(.dina(n13647), .dinb(n13583), .dout(n13648));
  jnot g13456(.din(n13648), .dout(n13649));
  jand g13457(.dina(\a[51] ), .dinb(\a[47] ), .dout(n13650));
  jand g13458(.dina(n13650), .dinb(n13449), .dout(n13651));
  jor  g13459(.dina(n13651), .dinb(n13649), .dout(n13652));
  jxor g13460(.dina(n13652), .dinb(n13469), .dout(n13653));
  jnot g13461(.din(n13552), .dout(n13654));
  jand g13462(.dina(\a[49] ), .dinb(n4774), .dout(n13655));
  jxor g13463(.dina(n13655), .dinb(n13654), .dout(n13656));
  jxor g13464(.dina(n13656), .dinb(n13653), .dout(n13657));
  jxor g13465(.dina(n13657), .dinb(n13646), .dout(n13658));
  jand g13466(.dina(n13600), .dinb(n13381), .dout(n13659));
  jor  g13467(.dina(n13659), .dinb(n13598), .dout(n13660));
  jand g13468(.dina(n13555), .dinb(n13549), .dout(n13661));
  jor  g13469(.dina(n13661), .dinb(n13553), .dout(n13662));
  jxor g13470(.dina(n13662), .dinb(n13660), .dout(n13663));
  jor  g13471(.dina(n13540), .dinb(n13538), .dout(n13664));
  jxor g13472(.dina(n13664), .dinb(n13663), .dout(n13665));
  jand g13473(.dina(n13556), .dinb(n13548), .dout(n13666));
  jand g13474(.dina(n13557), .dinb(n13532), .dout(n13667));
  jor  g13475(.dina(n13667), .dinb(n13666), .dout(n13668));
  jxor g13476(.dina(n13668), .dinb(n13665), .dout(n13669));
  jxor g13477(.dina(n13669), .dinb(n13658), .dout(n13670));
  jxor g13478(.dina(n13670), .dinb(n13643), .dout(n13671));
  jxor g13479(.dina(n13671), .dinb(n13625), .dout(n13672));
  jand g13480(.dina(n13528), .dinb(n13503), .dout(n13673));
  jand g13481(.dina(n13571), .dinb(n13529), .dout(n13674));
  jor  g13482(.dina(n13674), .dinb(n13673), .dout(n13675));
  jand g13483(.dina(n13569), .dinb(n13566), .dout(n13676));
  jand g13484(.dina(n13570), .dinb(n13558), .dout(n13677));
  jor  g13485(.dina(n13677), .dinb(n13676), .dout(n13678));
  jand g13486(.dina(n13526), .dinb(n13520), .dout(n13679));
  jand g13487(.dina(n13527), .dinb(n13512), .dout(n13680));
  jor  g13488(.dina(n13680), .dinb(n13679), .dout(n13681));
  jnot g13489(.din(n13539), .dout(n13682));
  jand g13490(.dina(\a[52] ), .dinb(\a[45] ), .dout(n13683));
  jand g13491(.dina(\a[53] ), .dinb(\a[44] ), .dout(n13684));
  jor  g13492(.dina(n13684), .dinb(n13683), .dout(n13685));
  jand g13493(.dina(\a[53] ), .dinb(\a[45] ), .dout(n13686));
  jand g13494(.dina(n13686), .dinb(n13438), .dout(n13687));
  jnot g13495(.din(n13687), .dout(n13688));
  jand g13496(.dina(n13688), .dinb(n13685), .dout(n13689));
  jxor g13497(.dina(n13689), .dinb(n13682), .dout(n13690));
  jand g13498(.dina(\a[60] ), .dinb(\a[37] ), .dout(n13691));
  jnot g13499(.din(n13691), .dout(n13692));
  jand g13500(.dina(\a[59] ), .dinb(\a[38] ), .dout(n13693));
  jor  g13501(.dina(n13693), .dinb(n13590), .dout(n13694));
  jand g13502(.dina(\a[59] ), .dinb(\a[39] ), .dout(n13695));
  jand g13503(.dina(n13695), .dinb(n13587), .dout(n13696));
  jnot g13504(.din(n13696), .dout(n13697));
  jand g13505(.dina(n13697), .dinb(n13694), .dout(n13698));
  jxor g13506(.dina(n13698), .dinb(n13692), .dout(n13699));
  jand g13507(.dina(\a[56] ), .dinb(\a[41] ), .dout(n13700));
  jnot g13508(.din(n13700), .dout(n13701));
  jxor g13509(.dina(n13536), .dinb(n13480), .dout(n13702));
  jxor g13510(.dina(n13702), .dinb(n13701), .dout(n13703));
  jnot g13511(.din(n13703), .dout(n13704));
  jxor g13512(.dina(n13704), .dinb(n13699), .dout(n13705));
  jxor g13513(.dina(n13705), .dinb(n13690), .dout(n13706));
  jxor g13514(.dina(n13706), .dinb(n13681), .dout(n13707));
  jxor g13515(.dina(n13707), .dinb(n13678), .dout(n13708));
  jxor g13516(.dina(n13708), .dinb(n13675), .dout(n13709));
  jxor g13517(.dina(n13709), .dinb(n13672), .dout(n13710));
  jxor g13518(.dina(n13710), .dinb(n13622), .dout(n13711));
  jand g13519(.dina(n13613), .dinb(n13500), .dout(n13712));
  jnot g13520(.din(n13500), .dout(n13713));
  jnot g13521(.din(n13613), .dout(n13714));
  jand g13522(.dina(n13714), .dinb(n13713), .dout(n13715));
  jnot g13523(.din(n13715), .dout(n13716));
  jand g13524(.dina(n13618), .dinb(n13716), .dout(n13717));
  jor  g13525(.dina(n13717), .dinb(n13712), .dout(n13718));
  jxor g13526(.dina(n13718), .dinb(n13711), .dout(\asquared[98] ));
  jand g13527(.dina(n13708), .dinb(n13675), .dout(n13720));
  jand g13528(.dina(n13709), .dinb(n13672), .dout(n13721));
  jor  g13529(.dina(n13721), .dinb(n13720), .dout(n13722));
  jand g13530(.dina(n13706), .dinb(n13681), .dout(n13723));
  jand g13531(.dina(n13707), .dinb(n13678), .dout(n13724));
  jor  g13532(.dina(n13724), .dinb(n13723), .dout(n13725));
  jand g13533(.dina(n13662), .dinb(n13660), .dout(n13726));
  jand g13534(.dina(n13664), .dinb(n13663), .dout(n13727));
  jor  g13535(.dina(n13727), .dinb(n13726), .dout(n13728));
  jand g13536(.dina(n13628), .dinb(n13626), .dout(n13729));
  jand g13537(.dina(n13631), .dinb(n13629), .dout(n13730));
  jor  g13538(.dina(n13730), .dinb(n13729), .dout(n13731));
  jxor g13539(.dina(n13731), .dinb(n13728), .dout(n13732));
  jnot g13540(.din(n13732), .dout(n13733));
  jnot g13541(.din(n13699), .dout(n13734));
  jand g13542(.dina(n13704), .dinb(n13734), .dout(n13735));
  jnot g13543(.din(n13735), .dout(n13736));
  jand g13544(.dina(n13703), .dinb(n13699), .dout(n13737));
  jor  g13545(.dina(n13737), .dinb(n13690), .dout(n13738));
  jand g13546(.dina(n13738), .dinb(n13736), .dout(n13739));
  jxor g13547(.dina(n13739), .dinb(n13733), .dout(n13740));
  jand g13548(.dina(n13694), .dinb(n13691), .dout(n13741));
  jor  g13549(.dina(n13741), .dinb(n13696), .dout(n13742));
  jnot g13550(.din(n13480), .dout(n13743));
  jnot g13551(.din(n13536), .dout(n13744));
  jand g13552(.dina(n13744), .dinb(n13743), .dout(n13745));
  jnot g13553(.din(n13745), .dout(n13746));
  jand g13554(.dina(n13536), .dinb(n13480), .dout(n13747));
  jor  g13555(.dina(n13747), .dinb(n13700), .dout(n13748));
  jand g13556(.dina(n13748), .dinb(n13746), .dout(n13749));
  jxor g13557(.dina(n13749), .dinb(n13742), .dout(n13750));
  jand g13558(.dina(n13685), .dinb(n13539), .dout(n13751));
  jor  g13559(.dina(n13751), .dinb(n13687), .dout(n13752));
  jxor g13560(.dina(n13752), .dinb(n13750), .dout(n13753));
  jnot g13561(.din(n13753), .dout(n13754));
  jor  g13562(.dina(n13656), .dinb(n13653), .dout(n13755));
  jand g13563(.dina(n13657), .dinb(n13646), .dout(n13756));
  jnot g13564(.din(n13756), .dout(n13757));
  jand g13565(.dina(n13757), .dinb(n13755), .dout(n13758));
  jxor g13566(.dina(n13758), .dinb(n13754), .dout(n13759));
  jand g13567(.dina(\a[61] ), .dinb(\a[37] ), .dout(n13760));
  jor  g13568(.dina(n13760), .dinb(n9513), .dout(n13761));
  jand g13569(.dina(\a[62] ), .dinb(\a[37] ), .dout(n13762));
  jand g13570(.dina(n13762), .dinb(n13626), .dout(n13763));
  jnot g13571(.din(n13763), .dout(n13764));
  jand g13572(.dina(n13764), .dinb(n13761), .dout(n13765));
  jnot g13573(.din(\a[49] ), .dout(n13766));
  jand g13574(.dina(n13654), .dinb(n4774), .dout(n13767));
  jor  g13575(.dina(n13767), .dinb(n13766), .dout(n13768));
  jnot g13576(.din(n13768), .dout(n13769));
  jxor g13577(.dina(n13769), .dinb(n13765), .dout(n13770));
  jand g13578(.dina(\a[52] ), .dinb(\a[46] ), .dout(n13771));
  jand g13579(.dina(\a[50] ), .dinb(\a[48] ), .dout(n13772));
  jor  g13580(.dina(n13772), .dinb(n13650), .dout(n13773));
  jnot g13581(.din(n13773), .dout(n13774));
  jand g13582(.dina(\a[51] ), .dinb(\a[48] ), .dout(n13775));
  jand g13583(.dina(n13775), .dinb(n13583), .dout(n13776));
  jor  g13584(.dina(n13776), .dinb(n13774), .dout(n13777));
  jxor g13585(.dina(n13777), .dinb(n13771), .dout(n13778));
  jnot g13586(.din(n13778), .dout(n13779));
  jand g13587(.dina(\a[58] ), .dinb(\a[40] ), .dout(n13780));
  jor  g13588(.dina(n13780), .dinb(n13695), .dout(n13781));
  jand g13589(.dina(n13597), .dinb(n13590), .dout(n13782));
  jnot g13590(.din(n13782), .dout(n13783));
  jand g13591(.dina(n13783), .dinb(n13781), .dout(n13784));
  jxor g13592(.dina(n13784), .dinb(n13686), .dout(n13785));
  jxor g13593(.dina(n13785), .dinb(n13779), .dout(n13786));
  jxor g13594(.dina(n13786), .dinb(n13770), .dout(n13787));
  jxor g13595(.dina(n13787), .dinb(n13759), .dout(n13788));
  jxor g13596(.dina(n13788), .dinb(n13740), .dout(n13789));
  jxor g13597(.dina(n13789), .dinb(n13725), .dout(n13790));
  jand g13598(.dina(n13670), .dinb(n13643), .dout(n13791));
  jand g13599(.dina(n13671), .dinb(n13625), .dout(n13792));
  jor  g13600(.dina(n13792), .dinb(n13791), .dout(n13793));
  jand g13601(.dina(n13668), .dinb(n13665), .dout(n13794));
  jand g13602(.dina(n13669), .dinb(n13658), .dout(n13795));
  jor  g13603(.dina(n13795), .dinb(n13794), .dout(n13796));
  jand g13604(.dina(n13641), .dinb(n13635), .dout(n13797));
  jand g13605(.dina(n13642), .dinb(n13632), .dout(n13798));
  jor  g13606(.dina(n13798), .dinb(n13797), .dout(n13799));
  jand g13607(.dina(\a[55] ), .dinb(\a[43] ), .dout(n13800));
  jand g13608(.dina(\a[54] ), .dinb(\a[44] ), .dout(n13801));
  jor  g13609(.dina(n13801), .dinb(n13800), .dout(n13802));
  jand g13610(.dina(\a[55] ), .dinb(\a[44] ), .dout(n13803));
  jand g13611(.dina(n13803), .dinb(n13539), .dout(n13804));
  jnot g13612(.din(n13804), .dout(n13805));
  jand g13613(.dina(n13805), .dinb(n13802), .dout(n13806));
  jand g13614(.dina(\a[63] ), .dinb(\a[35] ), .dout(n13807));
  jxor g13615(.dina(n13807), .dinb(n13806), .dout(n13808));
  jand g13616(.dina(n13648), .dinb(n13469), .dout(n13809));
  jor  g13617(.dina(n13809), .dinb(n13651), .dout(n13810));
  jxor g13618(.dina(n13810), .dinb(n13808), .dout(n13811));
  jnot g13619(.din(n13811), .dout(n13812));
  jand g13620(.dina(\a[60] ), .dinb(\a[38] ), .dout(n13813));
  jand g13621(.dina(\a[57] ), .dinb(\a[41] ), .dout(n13814));
  jand g13622(.dina(\a[56] ), .dinb(\a[42] ), .dout(n13815));
  jor  g13623(.dina(n13815), .dinb(n13814), .dout(n13816));
  jnot g13624(.din(n13816), .dout(n13817));
  jand g13625(.dina(\a[57] ), .dinb(\a[42] ), .dout(n13818));
  jand g13626(.dina(n13818), .dinb(n13700), .dout(n13819));
  jor  g13627(.dina(n13819), .dinb(n13817), .dout(n13820));
  jxor g13628(.dina(n13820), .dinb(n13813), .dout(n13821));
  jxor g13629(.dina(n13821), .dinb(n13812), .dout(n13822));
  jxor g13630(.dina(n13822), .dinb(n13799), .dout(n13823));
  jxor g13631(.dina(n13823), .dinb(n13796), .dout(n13824));
  jxor g13632(.dina(n13824), .dinb(n13793), .dout(n13825));
  jxor g13633(.dina(n13825), .dinb(n13790), .dout(n13826));
  jxor g13634(.dina(n13826), .dinb(n13722), .dout(n13827));
  jand g13635(.dina(n13710), .dinb(n13622), .dout(n13828));
  jor  g13636(.dina(n13710), .dinb(n13622), .dout(n13829));
  jand g13637(.dina(n13718), .dinb(n13829), .dout(n13830));
  jor  g13638(.dina(n13830), .dinb(n13828), .dout(n13831));
  jxor g13639(.dina(n13831), .dinb(n13827), .dout(\asquared[99] ));
  jand g13640(.dina(n13824), .dinb(n13793), .dout(n13833));
  jand g13641(.dina(n13825), .dinb(n13790), .dout(n13834));
  jor  g13642(.dina(n13834), .dinb(n13833), .dout(n13835));
  jand g13643(.dina(n13822), .dinb(n13799), .dout(n13836));
  jand g13644(.dina(n13823), .dinb(n13796), .dout(n13837));
  jor  g13645(.dina(n13837), .dinb(n13836), .dout(n13838));
  jand g13646(.dina(n13810), .dinb(n13808), .dout(n13839));
  jnot g13647(.din(n13839), .dout(n13840));
  jor  g13648(.dina(n13821), .dinb(n13812), .dout(n13841));
  jand g13649(.dina(n13841), .dinb(n13840), .dout(n13842));
  jnot g13650(.din(n13842), .dout(n13843));
  jand g13651(.dina(n13749), .dinb(n13742), .dout(n13844));
  jand g13652(.dina(n13752), .dinb(n13750), .dout(n13845));
  jor  g13653(.dina(n13845), .dinb(n13844), .dout(n13846));
  jnot g13654(.din(n13762), .dout(n13847));
  jand g13655(.dina(\a[50] ), .dinb(n13766), .dout(n13848));
  jxor g13656(.dina(n13848), .dinb(n13847), .dout(n13849));
  jnot g13657(.din(n13849), .dout(n13850));
  jxor g13658(.dina(n13850), .dinb(n13846), .dout(n13851));
  jxor g13659(.dina(n13851), .dinb(n13843), .dout(n13852));
  jand g13660(.dina(n13784), .dinb(n13686), .dout(n13853));
  jor  g13661(.dina(n13853), .dinb(n13782), .dout(n13854));
  jand g13662(.dina(n13773), .dinb(n13771), .dout(n13855));
  jor  g13663(.dina(n13855), .dinb(n13776), .dout(n13856));
  jxor g13664(.dina(n13856), .dinb(n13854), .dout(n13857));
  jand g13665(.dina(n13807), .dinb(n13806), .dout(n13858));
  jor  g13666(.dina(n13858), .dinb(n13804), .dout(n13859));
  jxor g13667(.dina(n13859), .dinb(n13857), .dout(n13860));
  jand g13668(.dina(n13785), .dinb(n13779), .dout(n13861));
  jand g13669(.dina(n13786), .dinb(n13770), .dout(n13862));
  jor  g13670(.dina(n13862), .dinb(n13861), .dout(n13863));
  jxor g13671(.dina(n13863), .dinb(n13860), .dout(n13864));
  jand g13672(.dina(n13769), .dinb(n13765), .dout(n13865));
  jor  g13673(.dina(n13865), .dinb(n13763), .dout(n13866));
  jand g13674(.dina(n13816), .dinb(n13813), .dout(n13867));
  jor  g13675(.dina(n13867), .dinb(n13819), .dout(n13868));
  jxor g13676(.dina(n13868), .dinb(n13866), .dout(n13869));
  jand g13677(.dina(\a[63] ), .dinb(\a[36] ), .dout(n13870));
  jand g13678(.dina(\a[60] ), .dinb(\a[39] ), .dout(n13871));
  jand g13679(.dina(\a[61] ), .dinb(\a[38] ), .dout(n13872));
  jor  g13680(.dina(n13872), .dinb(n13871), .dout(n13873));
  jnot g13681(.din(n13873), .dout(n13874));
  jand g13682(.dina(\a[61] ), .dinb(\a[39] ), .dout(n13875));
  jand g13683(.dina(n13875), .dinb(n13813), .dout(n13876));
  jor  g13684(.dina(n13876), .dinb(n13874), .dout(n13877));
  jxor g13685(.dina(n13877), .dinb(n13870), .dout(n13878));
  jnot g13686(.din(n13878), .dout(n13879));
  jxor g13687(.dina(n13879), .dinb(n13869), .dout(n13880));
  jxor g13688(.dina(n13880), .dinb(n13864), .dout(n13881));
  jxor g13689(.dina(n13881), .dinb(n13852), .dout(n13882));
  jxor g13690(.dina(n13882), .dinb(n13838), .dout(n13883));
  jand g13691(.dina(n13731), .dinb(n13728), .dout(n13884));
  jnot g13692(.din(n13884), .dout(n13885));
  jor  g13693(.dina(n13739), .dinb(n13733), .dout(n13886));
  jand g13694(.dina(n13886), .dinb(n13885), .dout(n13887));
  jnot g13695(.din(n13887), .dout(n13888));
  jnot g13696(.din(n13775), .dout(n13889));
  jand g13697(.dina(\a[56] ), .dinb(\a[43] ), .dout(n13890));
  jor  g13698(.dina(n13890), .dinb(n13818), .dout(n13891));
  jand g13699(.dina(\a[57] ), .dinb(\a[43] ), .dout(n13892));
  jand g13700(.dina(n13892), .dinb(n13815), .dout(n13893));
  jnot g13701(.din(n13893), .dout(n13894));
  jand g13702(.dina(n13894), .dinb(n13891), .dout(n13895));
  jxor g13703(.dina(n13895), .dinb(n13889), .dout(n13896));
  jand g13704(.dina(\a[54] ), .dinb(\a[45] ), .dout(n13897));
  jnot g13705(.din(n13897), .dout(n13898));
  jand g13706(.dina(\a[52] ), .dinb(\a[47] ), .dout(n13899));
  jand g13707(.dina(\a[53] ), .dinb(\a[46] ), .dout(n13900));
  jor  g13708(.dina(n13900), .dinb(n13899), .dout(n13901));
  jand g13709(.dina(\a[53] ), .dinb(\a[47] ), .dout(n13902));
  jand g13710(.dina(n13902), .dinb(n13771), .dout(n13903));
  jnot g13711(.din(n13903), .dout(n13904));
  jand g13712(.dina(n13904), .dinb(n13901), .dout(n13905));
  jxor g13713(.dina(n13905), .dinb(n13898), .dout(n13906));
  jnot g13714(.din(n13597), .dout(n13907));
  jand g13715(.dina(\a[58] ), .dinb(\a[41] ), .dout(n13908));
  jxor g13716(.dina(n13908), .dinb(n13803), .dout(n13909));
  jxor g13717(.dina(n13909), .dinb(n13907), .dout(n13910));
  jnot g13718(.din(n13910), .dout(n13911));
  jxor g13719(.dina(n13911), .dinb(n13906), .dout(n13912));
  jxor g13720(.dina(n13912), .dinb(n13896), .dout(n13913));
  jxor g13721(.dina(n13913), .dinb(n13888), .dout(n13914));
  jnot g13722(.din(n13914), .dout(n13915));
  jor  g13723(.dina(n13758), .dinb(n13754), .dout(n13916));
  jand g13724(.dina(n13787), .dinb(n13759), .dout(n13917));
  jnot g13725(.din(n13917), .dout(n13918));
  jand g13726(.dina(n13918), .dinb(n13916), .dout(n13919));
  jxor g13727(.dina(n13919), .dinb(n13915), .dout(n13920));
  jand g13728(.dina(n13788), .dinb(n13740), .dout(n13921));
  jand g13729(.dina(n13789), .dinb(n13725), .dout(n13922));
  jor  g13730(.dina(n13922), .dinb(n13921), .dout(n13923));
  jxor g13731(.dina(n13923), .dinb(n13920), .dout(n13924));
  jxor g13732(.dina(n13924), .dinb(n13883), .dout(n13925));
  jxor g13733(.dina(n13925), .dinb(n13835), .dout(n13926));
  jand g13734(.dina(n13826), .dinb(n13722), .dout(n13927));
  jnot g13735(.din(n13722), .dout(n13928));
  jnot g13736(.din(n13826), .dout(n13929));
  jand g13737(.dina(n13929), .dinb(n13928), .dout(n13930));
  jnot g13738(.din(n13930), .dout(n13931));
  jand g13739(.dina(n13831), .dinb(n13931), .dout(n13932));
  jor  g13740(.dina(n13932), .dinb(n13927), .dout(n13933));
  jxor g13741(.dina(n13933), .dinb(n13926), .dout(\asquared[100] ));
  jand g13742(.dina(n13923), .dinb(n13920), .dout(n13935));
  jand g13743(.dina(n13924), .dinb(n13883), .dout(n13936));
  jor  g13744(.dina(n13936), .dinb(n13935), .dout(n13937));
  jand g13745(.dina(n13856), .dinb(n13854), .dout(n13938));
  jand g13746(.dina(n13859), .dinb(n13857), .dout(n13939));
  jor  g13747(.dina(n13939), .dinb(n13938), .dout(n13940));
  jnot g13748(.din(n13940), .dout(n13941));
  jand g13749(.dina(\a[51] ), .dinb(\a[49] ), .dout(n13942));
  jand g13750(.dina(\a[52] ), .dinb(\a[48] ), .dout(n13943));
  jor  g13751(.dina(n13943), .dinb(n13942), .dout(n13944));
  jnot g13752(.din(n13944), .dout(n13945));
  jand g13753(.dina(\a[52] ), .dinb(\a[49] ), .dout(n13946));
  jand g13754(.dina(n13946), .dinb(n13775), .dout(n13947));
  jor  g13755(.dina(n13947), .dinb(n13945), .dout(n13948));
  jxor g13756(.dina(n13948), .dinb(n13902), .dout(n13949));
  jxor g13757(.dina(n13949), .dinb(n13941), .dout(n13950));
  jnot g13758(.din(n13866), .dout(n13951));
  jnot g13759(.din(n13868), .dout(n13952));
  jand g13760(.dina(n13952), .dinb(n13951), .dout(n13953));
  jnot g13761(.din(n13953), .dout(n13954));
  jand g13762(.dina(n13868), .dinb(n13866), .dout(n13955));
  jor  g13763(.dina(n13879), .dinb(n13955), .dout(n13956));
  jand g13764(.dina(n13956), .dinb(n13954), .dout(n13957));
  jxor g13765(.dina(n13957), .dinb(n13950), .dout(n13958));
  jnot g13766(.din(n13958), .dout(n13959));
  jand g13767(.dina(n13913), .dinb(n13888), .dout(n13960));
  jnot g13768(.din(n13960), .dout(n13961));
  jor  g13769(.dina(n13919), .dinb(n13915), .dout(n13962));
  jand g13770(.dina(n13962), .dinb(n13961), .dout(n13963));
  jxor g13771(.dina(n13963), .dinb(n13959), .dout(n13964));
  jand g13772(.dina(n13873), .dinb(n13870), .dout(n13965));
  jor  g13773(.dina(n13965), .dinb(n13876), .dout(n13966));
  jand g13774(.dina(n13901), .dinb(n13897), .dout(n13967));
  jor  g13775(.dina(n13967), .dinb(n13903), .dout(n13968));
  jxor g13776(.dina(n13968), .dinb(n13966), .dout(n13969));
  jnot g13777(.din(n13803), .dout(n13970));
  jnot g13778(.din(n13908), .dout(n13971));
  jand g13779(.dina(n13971), .dinb(n13970), .dout(n13972));
  jnot g13780(.din(n13972), .dout(n13973));
  jand g13781(.dina(n13908), .dinb(n13803), .dout(n13974));
  jor  g13782(.dina(n13974), .dinb(n13597), .dout(n13975));
  jand g13783(.dina(n13975), .dinb(n13973), .dout(n13976));
  jxor g13784(.dina(n13976), .dinb(n13969), .dout(n13977));
  jnot g13785(.din(n13977), .dout(n13978));
  jnot g13786(.din(n13906), .dout(n13979));
  jand g13787(.dina(n13911), .dinb(n13979), .dout(n13980));
  jnot g13788(.din(n13980), .dout(n13981));
  jand g13789(.dina(n13910), .dinb(n13906), .dout(n13982));
  jor  g13790(.dina(n13982), .dinb(n13896), .dout(n13983));
  jand g13791(.dina(n13983), .dinb(n13981), .dout(n13984));
  jxor g13792(.dina(n13984), .dinb(n13978), .dout(n13985));
  jnot g13793(.din(\a[50] ), .dout(n13986));
  jand g13794(.dina(n13847), .dinb(n13766), .dout(n13987));
  jor  g13795(.dina(n13987), .dinb(n13986), .dout(n13988));
  jnot g13796(.din(n13988), .dout(n13989));
  jand g13797(.dina(\a[63] ), .dinb(\a[37] ), .dout(n13990));
  jxor g13798(.dina(n13990), .dinb(n13989), .dout(n13991));
  jand g13799(.dina(n13891), .dinb(n13775), .dout(n13992));
  jor  g13800(.dina(n13992), .dinb(n13893), .dout(n13993));
  jxor g13801(.dina(n13993), .dinb(n13991), .dout(n13994));
  jxor g13802(.dina(n13994), .dinb(n13985), .dout(n13995));
  jxor g13803(.dina(n13995), .dinb(n13964), .dout(n13996));
  jand g13804(.dina(n13881), .dinb(n13852), .dout(n13997));
  jand g13805(.dina(n13882), .dinb(n13838), .dout(n13998));
  jor  g13806(.dina(n13998), .dinb(n13997), .dout(n13999));
  jand g13807(.dina(n13850), .dinb(n13846), .dout(n14000));
  jand g13808(.dina(n13851), .dinb(n13843), .dout(n14001));
  jor  g13809(.dina(n14001), .dinb(n14000), .dout(n14002));
  jand g13810(.dina(\a[54] ), .dinb(\a[46] ), .dout(n14003));
  jand g13811(.dina(\a[59] ), .dinb(\a[41] ), .dout(n14004));
  jand g13812(.dina(\a[58] ), .dinb(\a[42] ), .dout(n14005));
  jor  g13813(.dina(n14005), .dinb(n14004), .dout(n14006));
  jnot g13814(.din(n14006), .dout(n14007));
  jand g13815(.dina(\a[59] ), .dinb(\a[42] ), .dout(n14008));
  jand g13816(.dina(n14008), .dinb(n13908), .dout(n14009));
  jor  g13817(.dina(n14009), .dinb(n14007), .dout(n14010));
  jxor g13818(.dina(n14010), .dinb(n14003), .dout(n14011));
  jand g13819(.dina(\a[56] ), .dinb(\a[44] ), .dout(n14012));
  jor  g13820(.dina(n14012), .dinb(n13227), .dout(n14013));
  jnot g13821(.din(n14013), .dout(n14014));
  jand g13822(.dina(\a[56] ), .dinb(\a[45] ), .dout(n14015));
  jand g13823(.dina(n14015), .dinb(n13803), .dout(n14016));
  jor  g13824(.dina(n14016), .dinb(n14014), .dout(n14017));
  jxor g13825(.dina(n14017), .dinb(n13892), .dout(n14018));
  jand g13826(.dina(\a[62] ), .dinb(\a[38] ), .dout(n14019));
  jand g13827(.dina(\a[60] ), .dinb(\a[40] ), .dout(n14020));
  jor  g13828(.dina(n14020), .dinb(n13875), .dout(n14021));
  jand g13829(.dina(\a[61] ), .dinb(\a[40] ), .dout(n14022));
  jand g13830(.dina(n14022), .dinb(n13871), .dout(n14023));
  jnot g13831(.din(n14023), .dout(n14024));
  jand g13832(.dina(n14024), .dinb(n14021), .dout(n14025));
  jxor g13833(.dina(n14025), .dinb(n14019), .dout(n14026));
  jxor g13834(.dina(n14026), .dinb(n14018), .dout(n14027));
  jxor g13835(.dina(n14027), .dinb(n14011), .dout(n14028));
  jxor g13836(.dina(n14028), .dinb(n14002), .dout(n14029));
  jand g13837(.dina(n13863), .dinb(n13860), .dout(n14030));
  jand g13838(.dina(n13880), .dinb(n13864), .dout(n14031));
  jor  g13839(.dina(n14031), .dinb(n14030), .dout(n14032));
  jxor g13840(.dina(n14032), .dinb(n14029), .dout(n14033));
  jxor g13841(.dina(n14033), .dinb(n13999), .dout(n14034));
  jxor g13842(.dina(n14034), .dinb(n13996), .dout(n14035));
  jxor g13843(.dina(n14035), .dinb(n13937), .dout(n14036));
  jand g13844(.dina(n13925), .dinb(n13835), .dout(n14037));
  jor  g13845(.dina(n13925), .dinb(n13835), .dout(n14038));
  jand g13846(.dina(n13933), .dinb(n14038), .dout(n14039));
  jor  g13847(.dina(n14039), .dinb(n14037), .dout(n14040));
  jxor g13848(.dina(n14040), .dinb(n14036), .dout(\asquared[101] ));
  jand g13849(.dina(n14033), .dinb(n13999), .dout(n14042));
  jand g13850(.dina(n14034), .dinb(n13996), .dout(n14043));
  jor  g13851(.dina(n14043), .dinb(n14042), .dout(n14044));
  jor  g13852(.dina(n13963), .dinb(n13959), .dout(n14045));
  jand g13853(.dina(n13995), .dinb(n13964), .dout(n14046));
  jnot g13854(.din(n14046), .dout(n14047));
  jand g13855(.dina(n14047), .dinb(n14045), .dout(n14048));
  jnot g13856(.din(n14048), .dout(n14049));
  jor  g13857(.dina(n13949), .dinb(n13941), .dout(n14050));
  jand g13858(.dina(n13957), .dinb(n13950), .dout(n14051));
  jnot g13859(.din(n14051), .dout(n14052));
  jand g13860(.dina(n14052), .dinb(n14050), .dout(n14053));
  jnot g13861(.din(n14053), .dout(n14054));
  jand g13862(.dina(\a[58] ), .dinb(\a[43] ), .dout(n14055));
  jor  g13863(.dina(n14055), .dinb(n14015), .dout(n14056));
  jnot g13864(.din(n14056), .dout(n14057));
  jand g13865(.dina(\a[58] ), .dinb(\a[45] ), .dout(n14058));
  jand g13866(.dina(n14058), .dinb(n13890), .dout(n14059));
  jor  g13867(.dina(n14059), .dinb(n14057), .dout(n14060));
  jxor g13868(.dina(n14060), .dinb(n14008), .dout(n14061));
  jnot g13869(.din(n14061), .dout(n14062));
  jand g13870(.dina(\a[63] ), .dinb(\a[38] ), .dout(n14063));
  jand g13871(.dina(\a[55] ), .dinb(\a[46] ), .dout(n14064));
  jand g13872(.dina(\a[54] ), .dinb(\a[47] ), .dout(n14065));
  jor  g13873(.dina(n14065), .dinb(n14064), .dout(n14066));
  jand g13874(.dina(\a[55] ), .dinb(\a[47] ), .dout(n14067));
  jand g13875(.dina(n14067), .dinb(n14003), .dout(n14068));
  jnot g13876(.din(n14068), .dout(n14069));
  jand g13877(.dina(n14069), .dinb(n14066), .dout(n14070));
  jxor g13878(.dina(n14070), .dinb(n14063), .dout(n14071));
  jxor g13879(.dina(n14071), .dinb(n14062), .dout(n14072));
  jand g13880(.dina(\a[53] ), .dinb(\a[49] ), .dout(n14073));
  jand g13881(.dina(n14073), .dinb(n13943), .dout(n14074));
  jand g13882(.dina(\a[57] ), .dinb(\a[44] ), .dout(n14075));
  jand g13883(.dina(n14075), .dinb(n8716), .dout(n14076));
  jor  g13884(.dina(n14076), .dinb(n14074), .dout(n14077));
  jand g13885(.dina(\a[57] ), .dinb(\a[49] ), .dout(n14078));
  jand g13886(.dina(n14078), .dinb(n13438), .dout(n14079));
  jnot g13887(.din(n14079), .dout(n14080));
  jand g13888(.dina(n14080), .dinb(n14077), .dout(n14081));
  jnot g13889(.din(n14081), .dout(n14082));
  jor  g13890(.dina(n14075), .dinb(n13946), .dout(n14083));
  jand g13891(.dina(n14083), .dinb(n14080), .dout(n14084));
  jor  g13892(.dina(n14084), .dinb(n8716), .dout(n14085));
  jand g13893(.dina(n14085), .dinb(n14082), .dout(n14086));
  jxor g13894(.dina(n14086), .dinb(n14072), .dout(n14087));
  jxor g13895(.dina(n14087), .dinb(n14054), .dout(n14088));
  jand g13896(.dina(n13990), .dinb(n13989), .dout(n14089));
  jand g13897(.dina(n13993), .dinb(n13991), .dout(n14090));
  jor  g13898(.dina(n14090), .dinb(n14089), .dout(n14091));
  jand g13899(.dina(\a[60] ), .dinb(\a[41] ), .dout(n14092));
  jor  g13900(.dina(n14092), .dinb(n14022), .dout(n14093));
  jand g13901(.dina(\a[61] ), .dinb(\a[41] ), .dout(n14094));
  jand g13902(.dina(n14094), .dinb(n14020), .dout(n14095));
  jnot g13903(.din(n14095), .dout(n14096));
  jand g13904(.dina(n14096), .dinb(n14093), .dout(n14097));
  jand g13905(.dina(n13944), .dinb(n13902), .dout(n14098));
  jor  g13906(.dina(n14098), .dinb(n13947), .dout(n14099));
  jxor g13907(.dina(n14099), .dinb(n14097), .dout(n14100));
  jnot g13908(.din(n14100), .dout(n14101));
  jand g13909(.dina(\a[62] ), .dinb(\a[39] ), .dout(n14102));
  jnot g13910(.din(n14102), .dout(n14103));
  jand g13911(.dina(\a[51] ), .dinb(n13986), .dout(n14104));
  jxor g13912(.dina(n14104), .dinb(n14103), .dout(n14105));
  jxor g13913(.dina(n14105), .dinb(n14101), .dout(n14106));
  jxor g13914(.dina(n14106), .dinb(n14091), .dout(n14107));
  jxor g13915(.dina(n14107), .dinb(n14088), .dout(n14108));
  jxor g13916(.dina(n14108), .dinb(n14049), .dout(n14109));
  jand g13917(.dina(n14025), .dinb(n14019), .dout(n14110));
  jor  g13918(.dina(n14110), .dinb(n14023), .dout(n14111));
  jand g13919(.dina(n14006), .dinb(n14003), .dout(n14112));
  jor  g13920(.dina(n14112), .dinb(n14009), .dout(n14113));
  jxor g13921(.dina(n14113), .dinb(n14111), .dout(n14114));
  jand g13922(.dina(n14013), .dinb(n13892), .dout(n14115));
  jor  g13923(.dina(n14115), .dinb(n14016), .dout(n14116));
  jxor g13924(.dina(n14116), .dinb(n14114), .dout(n14117));
  jand g13925(.dina(n13968), .dinb(n13966), .dout(n14118));
  jand g13926(.dina(n13976), .dinb(n13969), .dout(n14119));
  jor  g13927(.dina(n14119), .dinb(n14118), .dout(n14120));
  jnot g13928(.din(n14018), .dout(n14121));
  jor  g13929(.dina(n14026), .dinb(n14121), .dout(n14122));
  jnot g13930(.din(n14011), .dout(n14123));
  jand g13931(.dina(n14026), .dinb(n14121), .dout(n14124));
  jor  g13932(.dina(n14124), .dinb(n14123), .dout(n14125));
  jand g13933(.dina(n14125), .dinb(n14122), .dout(n14126));
  jxor g13934(.dina(n14126), .dinb(n14120), .dout(n14127));
  jxor g13935(.dina(n14127), .dinb(n14117), .dout(n14128));
  jand g13936(.dina(n14028), .dinb(n14002), .dout(n14129));
  jand g13937(.dina(n14032), .dinb(n14029), .dout(n14130));
  jor  g13938(.dina(n14130), .dinb(n14129), .dout(n14131));
  jnot g13939(.din(n14131), .dout(n14132));
  jor  g13940(.dina(n13984), .dinb(n13978), .dout(n14133));
  jand g13941(.dina(n13994), .dinb(n13985), .dout(n14134));
  jnot g13942(.din(n14134), .dout(n14135));
  jand g13943(.dina(n14135), .dinb(n14133), .dout(n14136));
  jxor g13944(.dina(n14136), .dinb(n14132), .dout(n14137));
  jxor g13945(.dina(n14137), .dinb(n14128), .dout(n14138));
  jxor g13946(.dina(n14138), .dinb(n14109), .dout(n14139));
  jxor g13947(.dina(n14139), .dinb(n14044), .dout(n14140));
  jand g13948(.dina(n14035), .dinb(n13937), .dout(n14141));
  jor  g13949(.dina(n14035), .dinb(n13937), .dout(n14142));
  jand g13950(.dina(n14040), .dinb(n14142), .dout(n14143));
  jor  g13951(.dina(n14143), .dinb(n14141), .dout(n14144));
  jxor g13952(.dina(n14144), .dinb(n14140), .dout(\asquared[102] ));
  jand g13953(.dina(n14108), .dinb(n14049), .dout(n14146));
  jand g13954(.dina(n14138), .dinb(n14109), .dout(n14147));
  jor  g13955(.dina(n14147), .dinb(n14146), .dout(n14148));
  jand g13956(.dina(n14070), .dinb(n14063), .dout(n14149));
  jor  g13957(.dina(n14149), .dinb(n14068), .dout(n14150));
  jor  g13958(.dina(n14079), .dinb(n14077), .dout(n14151));
  jnot g13959(.din(\a[51] ), .dout(n14152));
  jand g13960(.dina(n14103), .dinb(n13986), .dout(n14153));
  jor  g13961(.dina(n14153), .dinb(n14152), .dout(n14154));
  jnot g13962(.din(n14154), .dout(n14155));
  jxor g13963(.dina(n14155), .dinb(n14151), .dout(n14156));
  jxor g13964(.dina(n14156), .dinb(n14150), .dout(n14157));
  jand g13965(.dina(n14113), .dinb(n14111), .dout(n14158));
  jand g13966(.dina(n14116), .dinb(n14114), .dout(n14159));
  jor  g13967(.dina(n14159), .dinb(n14158), .dout(n14160));
  jxor g13968(.dina(n14160), .dinb(n14157), .dout(n14161));
  jand g13969(.dina(n14071), .dinb(n14062), .dout(n14162));
  jand g13970(.dina(n14086), .dinb(n14072), .dout(n14163));
  jor  g13971(.dina(n14163), .dinb(n14162), .dout(n14164));
  jxor g13972(.dina(n14164), .dinb(n14161), .dout(n14165));
  jand g13973(.dina(n14087), .dinb(n14054), .dout(n14166));
  jand g13974(.dina(n14107), .dinb(n14088), .dout(n14167));
  jor  g13975(.dina(n14167), .dinb(n14166), .dout(n14168));
  jand g13976(.dina(n14126), .dinb(n14120), .dout(n14169));
  jand g13977(.dina(n14127), .dinb(n14117), .dout(n14170));
  jor  g13978(.dina(n14170), .dinb(n14169), .dout(n14171));
  jxor g13979(.dina(n14171), .dinb(n14168), .dout(n14172));
  jxor g13980(.dina(n14172), .dinb(n14165), .dout(n14173));
  jor  g13981(.dina(n14136), .dinb(n14132), .dout(n14174));
  jand g13982(.dina(n14137), .dinb(n14128), .dout(n14175));
  jnot g13983(.din(n14175), .dout(n14176));
  jand g13984(.dina(n14176), .dinb(n14174), .dout(n14177));
  jnot g13985(.din(n14177), .dout(n14178));
  jor  g13986(.dina(n14105), .dinb(n14101), .dout(n14179));
  jand g13987(.dina(n14106), .dinb(n14091), .dout(n14180));
  jnot g13988(.din(n14180), .dout(n14181));
  jand g13989(.dina(n14181), .dinb(n14179), .dout(n14182));
  jnot g13990(.din(n14182), .dout(n14183));
  jand g13991(.dina(n14099), .dinb(n14097), .dout(n14184));
  jor  g13992(.dina(n14184), .dinb(n14095), .dout(n14185));
  jand g13993(.dina(n14056), .dinb(n14008), .dout(n14186));
  jor  g13994(.dina(n14186), .dinb(n14059), .dout(n14187));
  jxor g13995(.dina(n14187), .dinb(n14185), .dout(n14188));
  jand g13996(.dina(\a[63] ), .dinb(\a[39] ), .dout(n14189));
  jand g13997(.dina(\a[60] ), .dinb(\a[42] ), .dout(n14190));
  jor  g13998(.dina(n14190), .dinb(n14094), .dout(n14191));
  jnot g13999(.din(n14191), .dout(n14192));
  jand g14000(.dina(\a[61] ), .dinb(\a[42] ), .dout(n14193));
  jand g14001(.dina(n14193), .dinb(n14092), .dout(n14194));
  jor  g14002(.dina(n14194), .dinb(n14192), .dout(n14195));
  jxor g14003(.dina(n14195), .dinb(n14189), .dout(n14196));
  jnot g14004(.din(n14196), .dout(n14197));
  jxor g14005(.dina(n14197), .dinb(n14188), .dout(n14198));
  jxor g14006(.dina(n14198), .dinb(n14183), .dout(n14199));
  jand g14007(.dina(\a[54] ), .dinb(\a[48] ), .dout(n14200));
  jand g14008(.dina(\a[52] ), .dinb(\a[50] ), .dout(n14201));
  jor  g14009(.dina(n14201), .dinb(n14073), .dout(n14202));
  jnot g14010(.din(n14202), .dout(n14203));
  jand g14011(.dina(\a[53] ), .dinb(\a[50] ), .dout(n14204));
  jand g14012(.dina(n14204), .dinb(n13946), .dout(n14205));
  jor  g14013(.dina(n14205), .dinb(n14203), .dout(n14206));
  jxor g14014(.dina(n14206), .dinb(n14200), .dout(n14207));
  jnot g14015(.din(n14207), .dout(n14208));
  jand g14016(.dina(\a[57] ), .dinb(\a[45] ), .dout(n14209));
  jand g14017(.dina(\a[56] ), .dinb(\a[46] ), .dout(n14210));
  jor  g14018(.dina(n14210), .dinb(n14067), .dout(n14211));
  jnot g14019(.din(n14211), .dout(n14212));
  jand g14020(.dina(\a[56] ), .dinb(\a[47] ), .dout(n14213));
  jand g14021(.dina(n14213), .dinb(n14064), .dout(n14214));
  jor  g14022(.dina(n14214), .dinb(n14212), .dout(n14215));
  jxor g14023(.dina(n14215), .dinb(n14209), .dout(n14216));
  jnot g14024(.din(n14216), .dout(n14217));
  jand g14025(.dina(\a[58] ), .dinb(\a[44] ), .dout(n14218));
  jnot g14026(.din(n14218), .dout(n14219));
  jand g14027(.dina(\a[59] ), .dinb(\a[43] ), .dout(n14220));
  jnot g14028(.din(n14220), .dout(n14221));
  jand g14029(.dina(n14221), .dinb(n14219), .dout(n14222));
  jand g14030(.dina(\a[59] ), .dinb(\a[44] ), .dout(n14223));
  jand g14031(.dina(n14223), .dinb(n14055), .dout(n14224));
  jor  g14032(.dina(n14224), .dinb(n14222), .dout(n14225));
  jnot g14033(.din(n14225), .dout(n14226));
  jxor g14034(.dina(n14226), .dinb(n11055), .dout(n14227));
  jxor g14035(.dina(n14227), .dinb(n14217), .dout(n14228));
  jxor g14036(.dina(n14228), .dinb(n14208), .dout(n14229));
  jxor g14037(.dina(n14229), .dinb(n14199), .dout(n14230));
  jxor g14038(.dina(n14230), .dinb(n14178), .dout(n14231));
  jxor g14039(.dina(n14231), .dinb(n14173), .dout(n14232));
  jxor g14040(.dina(n14232), .dinb(n14148), .dout(n14233));
  jand g14041(.dina(n14139), .dinb(n14044), .dout(n14234));
  jor  g14042(.dina(n14139), .dinb(n14044), .dout(n14235));
  jand g14043(.dina(n14144), .dinb(n14235), .dout(n14236));
  jor  g14044(.dina(n14236), .dinb(n14234), .dout(n14237));
  jxor g14045(.dina(n14237), .dinb(n14233), .dout(\asquared[103] ));
  jand g14046(.dina(n14230), .dinb(n14178), .dout(n14239));
  jand g14047(.dina(n14231), .dinb(n14173), .dout(n14240));
  jor  g14048(.dina(n14240), .dinb(n14239), .dout(n14241));
  jand g14049(.dina(n14155), .dinb(n14151), .dout(n14242));
  jand g14050(.dina(n14156), .dinb(n14150), .dout(n14243));
  jor  g14051(.dina(n14243), .dinb(n14242), .dout(n14244));
  jnot g14052(.din(n14185), .dout(n14245));
  jnot g14053(.din(n14187), .dout(n14246));
  jand g14054(.dina(n14246), .dinb(n14245), .dout(n14247));
  jnot g14055(.din(n14247), .dout(n14248));
  jand g14056(.dina(n14187), .dinb(n14185), .dout(n14249));
  jor  g14057(.dina(n14197), .dinb(n14249), .dout(n14250));
  jand g14058(.dina(n14250), .dinb(n14248), .dout(n14251));
  jxor g14059(.dina(n14251), .dinb(n14244), .dout(n14252));
  jor  g14060(.dina(n14227), .dinb(n14217), .dout(n14253));
  jand g14061(.dina(n14227), .dinb(n14217), .dout(n14254));
  jor  g14062(.dina(n14254), .dinb(n14208), .dout(n14255));
  jand g14063(.dina(n14255), .dinb(n14253), .dout(n14256));
  jxor g14064(.dina(n14256), .dinb(n14252), .dout(n14257));
  jand g14065(.dina(n14198), .dinb(n14183), .dout(n14258));
  jand g14066(.dina(n14229), .dinb(n14199), .dout(n14259));
  jor  g14067(.dina(n14259), .dinb(n14258), .dout(n14260));
  jand g14068(.dina(n14160), .dinb(n14157), .dout(n14261));
  jand g14069(.dina(n14164), .dinb(n14161), .dout(n14262));
  jor  g14070(.dina(n14262), .dinb(n14261), .dout(n14263));
  jxor g14071(.dina(n14263), .dinb(n14260), .dout(n14264));
  jxor g14072(.dina(n14264), .dinb(n14257), .dout(n14265));
  jand g14073(.dina(n14171), .dinb(n14168), .dout(n14266));
  jand g14074(.dina(n14172), .dinb(n14165), .dout(n14267));
  jor  g14075(.dina(n14267), .dinb(n14266), .dout(n14268));
  jand g14076(.dina(\a[63] ), .dinb(\a[40] ), .dout(n14269));
  jand g14077(.dina(n14202), .dinb(n14200), .dout(n14270));
  jor  g14078(.dina(n14270), .dinb(n14205), .dout(n14271));
  jxor g14079(.dina(n14271), .dinb(n14269), .dout(n14272));
  jand g14080(.dina(n14211), .dinb(n14209), .dout(n14273));
  jor  g14081(.dina(n14273), .dinb(n14214), .dout(n14274));
  jxor g14082(.dina(n14274), .dinb(n14272), .dout(n14275));
  jand g14083(.dina(n14226), .dinb(n11055), .dout(n14276));
  jor  g14084(.dina(n14276), .dinb(n14224), .dout(n14277));
  jand g14085(.dina(n14191), .dinb(n14189), .dout(n14278));
  jor  g14086(.dina(n14278), .dinb(n14194), .dout(n14279));
  jxor g14087(.dina(n14279), .dinb(n14277), .dout(n14280));
  jor  g14088(.dina(n14223), .dinb(n14058), .dout(n14281));
  jnot g14089(.din(n14281), .dout(n14282));
  jand g14090(.dina(\a[59] ), .dinb(\a[45] ), .dout(n14283));
  jand g14091(.dina(n14283), .dinb(n14218), .dout(n14284));
  jor  g14092(.dina(n14284), .dinb(n14282), .dout(n14285));
  jxor g14093(.dina(n14285), .dinb(n14193), .dout(n14286));
  jnot g14094(.din(n14286), .dout(n14287));
  jxor g14095(.dina(n14287), .dinb(n14280), .dout(n14288));
  jxor g14096(.dina(n14288), .dinb(n14275), .dout(n14289));
  jand g14097(.dina(\a[55] ), .dinb(\a[48] ), .dout(n14290));
  jand g14098(.dina(\a[54] ), .dinb(\a[49] ), .dout(n14291));
  jor  g14099(.dina(n14291), .dinb(n14204), .dout(n14292));
  jnot g14100(.din(n14292), .dout(n14293));
  jand g14101(.dina(\a[54] ), .dinb(\a[50] ), .dout(n14294));
  jand g14102(.dina(n14294), .dinb(n14073), .dout(n14295));
  jor  g14103(.dina(n14295), .dinb(n14293), .dout(n14296));
  jxor g14104(.dina(n14296), .dinb(n14290), .dout(n14297));
  jnot g14105(.din(n14297), .dout(n14298));
  jand g14106(.dina(\a[60] ), .dinb(\a[43] ), .dout(n14299));
  jand g14107(.dina(\a[57] ), .dinb(\a[46] ), .dout(n14300));
  jor  g14108(.dina(n14300), .dinb(n14213), .dout(n14301));
  jand g14109(.dina(\a[57] ), .dinb(\a[47] ), .dout(n14302));
  jand g14110(.dina(n14302), .dinb(n14210), .dout(n14303));
  jnot g14111(.din(n14303), .dout(n14304));
  jand g14112(.dina(n14304), .dinb(n14301), .dout(n14305));
  jxor g14113(.dina(n14305), .dinb(n14299), .dout(n14306));
  jxor g14114(.dina(n14306), .dinb(n14298), .dout(n14307));
  jand g14115(.dina(\a[62] ), .dinb(\a[41] ), .dout(n14308));
  jnot g14116(.din(n14308), .dout(n14309));
  jand g14117(.dina(\a[52] ), .dinb(n14152), .dout(n14310));
  jxor g14118(.dina(n14310), .dinb(n14309), .dout(n14311));
  jnot g14119(.din(n14311), .dout(n14312));
  jxor g14120(.dina(n14312), .dinb(n14307), .dout(n14313));
  jxor g14121(.dina(n14313), .dinb(n14289), .dout(n14314));
  jxor g14122(.dina(n14314), .dinb(n14268), .dout(n14315));
  jxor g14123(.dina(n14315), .dinb(n14265), .dout(n14316));
  jxor g14124(.dina(n14316), .dinb(n14241), .dout(n14317));
  jand g14125(.dina(n14232), .dinb(n14148), .dout(n14318));
  jnot g14126(.din(n14148), .dout(n14319));
  jnot g14127(.din(n14232), .dout(n14320));
  jand g14128(.dina(n14320), .dinb(n14319), .dout(n14321));
  jnot g14129(.din(n14321), .dout(n14322));
  jand g14130(.dina(n14237), .dinb(n14322), .dout(n14323));
  jor  g14131(.dina(n14323), .dinb(n14318), .dout(n14324));
  jxor g14132(.dina(n14324), .dinb(n14317), .dout(\asquared[104] ));
  jand g14133(.dina(n14314), .dinb(n14268), .dout(n14326));
  jand g14134(.dina(n14315), .dinb(n14265), .dout(n14327));
  jor  g14135(.dina(n14327), .dinb(n14326), .dout(n14328));
  jand g14136(.dina(n14251), .dinb(n14244), .dout(n14329));
  jand g14137(.dina(n14256), .dinb(n14252), .dout(n14330));
  jor  g14138(.dina(n14330), .dinb(n14329), .dout(n14331));
  jnot g14139(.din(n14275), .dout(n14332));
  jnot g14140(.din(n14288), .dout(n14333));
  jand g14141(.dina(n14333), .dinb(n14332), .dout(n14334));
  jnot g14142(.din(n14334), .dout(n14335));
  jand g14143(.dina(n14288), .dinb(n14275), .dout(n14336));
  jor  g14144(.dina(n14313), .dinb(n14336), .dout(n14337));
  jand g14145(.dina(n14337), .dinb(n14335), .dout(n14338));
  jxor g14146(.dina(n14338), .dinb(n14331), .dout(n14339));
  jand g14147(.dina(n14271), .dinb(n14269), .dout(n14340));
  jand g14148(.dina(n14274), .dinb(n14272), .dout(n14341));
  jor  g14149(.dina(n14341), .dinb(n14340), .dout(n14342));
  jnot g14150(.din(\a[52] ), .dout(n14343));
  jand g14151(.dina(n14309), .dinb(n14152), .dout(n14344));
  jor  g14152(.dina(n14344), .dinb(n14343), .dout(n14345));
  jnot g14153(.din(n14345), .dout(n14346));
  jand g14154(.dina(\a[62] ), .dinb(\a[42] ), .dout(n14347));
  jand g14155(.dina(\a[63] ), .dinb(\a[41] ), .dout(n14348));
  jor  g14156(.dina(n14348), .dinb(n14347), .dout(n14349));
  jand g14157(.dina(\a[63] ), .dinb(\a[42] ), .dout(n14350));
  jand g14158(.dina(n14350), .dinb(n14308), .dout(n14351));
  jnot g14159(.din(n14351), .dout(n14352));
  jand g14160(.dina(n14352), .dinb(n14349), .dout(n14353));
  jxor g14161(.dina(n14353), .dinb(n14346), .dout(n14354));
  jxor g14162(.dina(n14354), .dinb(n14342), .dout(n14355));
  jnot g14163(.din(n14277), .dout(n14356));
  jnot g14164(.din(n14279), .dout(n14357));
  jand g14165(.dina(n14357), .dinb(n14356), .dout(n14358));
  jnot g14166(.din(n14358), .dout(n14359));
  jand g14167(.dina(n14279), .dinb(n14277), .dout(n14360));
  jor  g14168(.dina(n14287), .dinb(n14360), .dout(n14361));
  jand g14169(.dina(n14361), .dinb(n14359), .dout(n14362));
  jxor g14170(.dina(n14362), .dinb(n14355), .dout(n14363));
  jxor g14171(.dina(n14363), .dinb(n14339), .dout(n14364));
  jand g14172(.dina(n14263), .dinb(n14260), .dout(n14365));
  jand g14173(.dina(n14264), .dinb(n14257), .dout(n14366));
  jor  g14174(.dina(n14366), .dinb(n14365), .dout(n14367));
  jand g14175(.dina(n14305), .dinb(n14299), .dout(n14368));
  jor  g14176(.dina(n14368), .dinb(n14303), .dout(n14369));
  jand g14177(.dina(n14292), .dinb(n14290), .dout(n14370));
  jor  g14178(.dina(n14370), .dinb(n14295), .dout(n14371));
  jxor g14179(.dina(n14371), .dinb(n14369), .dout(n14372));
  jand g14180(.dina(n14281), .dinb(n14193), .dout(n14373));
  jor  g14181(.dina(n14373), .dinb(n14284), .dout(n14374));
  jxor g14182(.dina(n14374), .dinb(n14372), .dout(n14375));
  jor  g14183(.dina(n14306), .dinb(n14298), .dout(n14376));
  jand g14184(.dina(n14306), .dinb(n14298), .dout(n14377));
  jor  g14185(.dina(n14312), .dinb(n14377), .dout(n14378));
  jand g14186(.dina(n14378), .dinb(n14376), .dout(n14379));
  jxor g14187(.dina(n14379), .dinb(n14375), .dout(n14380));
  jand g14188(.dina(\a[58] ), .dinb(\a[46] ), .dout(n14381));
  jand g14189(.dina(\a[56] ), .dinb(\a[48] ), .dout(n14382));
  jor  g14190(.dina(n14382), .dinb(n14302), .dout(n14383));
  jnot g14191(.din(n14383), .dout(n14384));
  jand g14192(.dina(\a[57] ), .dinb(\a[48] ), .dout(n14385));
  jand g14193(.dina(n14385), .dinb(n14213), .dout(n14386));
  jor  g14194(.dina(n14386), .dinb(n14384), .dout(n14387));
  jxor g14195(.dina(n14387), .dinb(n14381), .dout(n14388));
  jnot g14196(.din(n14388), .dout(n14389));
  jand g14197(.dina(\a[60] ), .dinb(\a[44] ), .dout(n14390));
  jand g14198(.dina(\a[61] ), .dinb(\a[43] ), .dout(n14391));
  jor  g14199(.dina(n14391), .dinb(n14283), .dout(n14392));
  jand g14200(.dina(\a[61] ), .dinb(\a[45] ), .dout(n14393));
  jand g14201(.dina(n14393), .dinb(n14220), .dout(n14394));
  jnot g14202(.din(n14394), .dout(n14395));
  jand g14203(.dina(n14395), .dinb(n14392), .dout(n14396));
  jxor g14204(.dina(n14396), .dinb(n14390), .dout(n14397));
  jxor g14205(.dina(n14397), .dinb(n14389), .dout(n14398));
  jnot g14206(.din(n14398), .dout(n14399));
  jand g14207(.dina(\a[55] ), .dinb(\a[49] ), .dout(n14400));
  jand g14208(.dina(\a[53] ), .dinb(\a[51] ), .dout(n14401));
  jor  g14209(.dina(n14401), .dinb(n14294), .dout(n14402));
  jnot g14210(.din(n14402), .dout(n14403));
  jand g14211(.dina(\a[54] ), .dinb(\a[51] ), .dout(n14404));
  jand g14212(.dina(n14404), .dinb(n14204), .dout(n14405));
  jor  g14213(.dina(n14405), .dinb(n14403), .dout(n14406));
  jxor g14214(.dina(n14406), .dinb(n14400), .dout(n14407));
  jxor g14215(.dina(n14407), .dinb(n14399), .dout(n14408));
  jxor g14216(.dina(n14408), .dinb(n14380), .dout(n14409));
  jxor g14217(.dina(n14409), .dinb(n14367), .dout(n14410));
  jxor g14218(.dina(n14410), .dinb(n14364), .dout(n14411));
  jxor g14219(.dina(n14411), .dinb(n14328), .dout(n14412));
  jand g14220(.dina(n14316), .dinb(n14241), .dout(n14413));
  jor  g14221(.dina(n14316), .dinb(n14241), .dout(n14414));
  jand g14222(.dina(n14324), .dinb(n14414), .dout(n14415));
  jor  g14223(.dina(n14415), .dinb(n14413), .dout(n14416));
  jxor g14224(.dina(n14416), .dinb(n14412), .dout(\asquared[105] ));
  jand g14225(.dina(n14396), .dinb(n14390), .dout(n14418));
  jor  g14226(.dina(n14418), .dinb(n14394), .dout(n14419));
  jand g14227(.dina(n14383), .dinb(n14381), .dout(n14420));
  jor  g14228(.dina(n14420), .dinb(n14386), .dout(n14421));
  jand g14229(.dina(n14402), .dinb(n14400), .dout(n14422));
  jor  g14230(.dina(n14422), .dinb(n14405), .dout(n14423));
  jxor g14231(.dina(n14423), .dinb(n14421), .dout(n14424));
  jxor g14232(.dina(n14424), .dinb(n14419), .dout(n14425));
  jnot g14233(.din(n14425), .dout(n14426));
  jand g14234(.dina(n14397), .dinb(n14389), .dout(n14427));
  jnot g14235(.din(n14427), .dout(n14428));
  jor  g14236(.dina(n14407), .dinb(n14399), .dout(n14429));
  jand g14237(.dina(n14429), .dinb(n14428), .dout(n14430));
  jxor g14238(.dina(n14430), .dinb(n14426), .dout(n14431));
  jand g14239(.dina(n14354), .dinb(n14342), .dout(n14432));
  jand g14240(.dina(n14362), .dinb(n14355), .dout(n14433));
  jor  g14241(.dina(n14433), .dinb(n14432), .dout(n14434));
  jxor g14242(.dina(n14434), .dinb(n14431), .dout(n14435));
  jand g14243(.dina(n14338), .dinb(n14331), .dout(n14436));
  jand g14244(.dina(n14363), .dinb(n14339), .dout(n14437));
  jor  g14245(.dina(n14437), .dinb(n14436), .dout(n14438));
  jxor g14246(.dina(n14438), .dinb(n14435), .dout(n14439));
  jand g14247(.dina(n14379), .dinb(n14375), .dout(n14440));
  jand g14248(.dina(n14408), .dinb(n14380), .dout(n14441));
  jor  g14249(.dina(n14441), .dinb(n14440), .dout(n14442));
  jand g14250(.dina(n14371), .dinb(n14369), .dout(n14443));
  jand g14251(.dina(n14374), .dinb(n14372), .dout(n14444));
  jor  g14252(.dina(n14444), .dinb(n14443), .dout(n14445));
  jand g14253(.dina(\a[56] ), .dinb(\a[49] ), .dout(n14446));
  jand g14254(.dina(\a[55] ), .dinb(\a[50] ), .dout(n14447));
  jor  g14255(.dina(n14447), .dinb(n14404), .dout(n14448));
  jnot g14256(.din(n14448), .dout(n14449));
  jand g14257(.dina(\a[55] ), .dinb(\a[51] ), .dout(n14450));
  jand g14258(.dina(n14450), .dinb(n14294), .dout(n14451));
  jor  g14259(.dina(n14451), .dinb(n14449), .dout(n14452));
  jxor g14260(.dina(n14452), .dinb(n14446), .dout(n14453));
  jand g14261(.dina(\a[62] ), .dinb(\a[43] ), .dout(n14454));
  jnot g14262(.din(n14454), .dout(n14455));
  jand g14263(.dina(\a[53] ), .dinb(n14343), .dout(n14456));
  jxor g14264(.dina(n14456), .dinb(n14455), .dout(n14457));
  jxor g14265(.dina(n14457), .dinb(n14453), .dout(n14458));
  jxor g14266(.dina(n14458), .dinb(n14445), .dout(n14459));
  jand g14267(.dina(\a[59] ), .dinb(\a[46] ), .dout(n14460));
  jand g14268(.dina(\a[58] ), .dinb(\a[47] ), .dout(n14461));
  jor  g14269(.dina(n14461), .dinb(n14385), .dout(n14462));
  jnot g14270(.din(n14462), .dout(n14463));
  jand g14271(.dina(\a[58] ), .dinb(\a[48] ), .dout(n14464));
  jand g14272(.dina(n14464), .dinb(n14302), .dout(n14465));
  jor  g14273(.dina(n14465), .dinb(n14463), .dout(n14466));
  jxor g14274(.dina(n14466), .dinb(n14460), .dout(n14467));
  jnot g14275(.din(n14467), .dout(n14468));
  jand g14276(.dina(\a[61] ), .dinb(\a[44] ), .dout(n14469));
  jand g14277(.dina(\a[60] ), .dinb(\a[45] ), .dout(n14470));
  jor  g14278(.dina(n14470), .dinb(n14469), .dout(n14471));
  jnot g14279(.din(n14471), .dout(n14472));
  jand g14280(.dina(n14393), .dinb(n14390), .dout(n14473));
  jor  g14281(.dina(n14473), .dinb(n14472), .dout(n14474));
  jxor g14282(.dina(n14474), .dinb(n14350), .dout(n14475));
  jnot g14283(.din(n14475), .dout(n14476));
  jand g14284(.dina(n14353), .dinb(n14346), .dout(n14477));
  jor  g14285(.dina(n14477), .dinb(n14351), .dout(n14478));
  jxor g14286(.dina(n14478), .dinb(n14476), .dout(n14479));
  jxor g14287(.dina(n14479), .dinb(n14468), .dout(n14480));
  jxor g14288(.dina(n14480), .dinb(n14459), .dout(n14481));
  jxor g14289(.dina(n14481), .dinb(n14442), .dout(n14482));
  jxor g14290(.dina(n14482), .dinb(n14439), .dout(n14483));
  jand g14291(.dina(n14409), .dinb(n14367), .dout(n14484));
  jand g14292(.dina(n14410), .dinb(n14364), .dout(n14485));
  jor  g14293(.dina(n14485), .dinb(n14484), .dout(n14486));
  jxor g14294(.dina(n14486), .dinb(n14483), .dout(n14487));
  jand g14295(.dina(n14411), .dinb(n14328), .dout(n14488));
  jor  g14296(.dina(n14411), .dinb(n14328), .dout(n14489));
  jand g14297(.dina(n14416), .dinb(n14489), .dout(n14490));
  jor  g14298(.dina(n14490), .dinb(n14488), .dout(n14491));
  jxor g14299(.dina(n14491), .dinb(n14487), .dout(\asquared[106] ));
  jand g14300(.dina(n14438), .dinb(n14435), .dout(n14493));
  jand g14301(.dina(n14482), .dinb(n14439), .dout(n14494));
  jor  g14302(.dina(n14494), .dinb(n14493), .dout(n14495));
  jand g14303(.dina(\a[63] ), .dinb(\a[43] ), .dout(n14496));
  jnot g14304(.din(\a[53] ), .dout(n14497));
  jand g14305(.dina(n14455), .dinb(n14343), .dout(n14498));
  jor  g14306(.dina(n14498), .dinb(n14497), .dout(n14499));
  jnot g14307(.din(n14499), .dout(n14500));
  jxor g14308(.dina(n14500), .dinb(n14496), .dout(n14501));
  jand g14309(.dina(n14448), .dinb(n14446), .dout(n14502));
  jor  g14310(.dina(n14502), .dinb(n14451), .dout(n14503));
  jxor g14311(.dina(n14503), .dinb(n14501), .dout(n14504));
  jand g14312(.dina(n14478), .dinb(n14476), .dout(n14505));
  jand g14313(.dina(n14479), .dinb(n14468), .dout(n14506));
  jor  g14314(.dina(n14506), .dinb(n14505), .dout(n14507));
  jxor g14315(.dina(n14507), .dinb(n14504), .dout(n14508));
  jnot g14316(.din(n14508), .dout(n14509));
  jor  g14317(.dina(n14457), .dinb(n14453), .dout(n14510));
  jand g14318(.dina(n14458), .dinb(n14445), .dout(n14511));
  jnot g14319(.din(n14511), .dout(n14512));
  jand g14320(.dina(n14512), .dinb(n14510), .dout(n14513));
  jxor g14321(.dina(n14513), .dinb(n14509), .dout(n14514));
  jand g14322(.dina(n14480), .dinb(n14459), .dout(n14515));
  jand g14323(.dina(n14481), .dinb(n14442), .dout(n14516));
  jor  g14324(.dina(n14516), .dinb(n14515), .dout(n14517));
  jxor g14325(.dina(n14517), .dinb(n14514), .dout(n14518));
  jor  g14326(.dina(n14430), .dinb(n14426), .dout(n14519));
  jand g14327(.dina(n14434), .dinb(n14431), .dout(n14520));
  jnot g14328(.din(n14520), .dout(n14521));
  jand g14329(.dina(n14521), .dinb(n14519), .dout(n14522));
  jnot g14330(.din(n14522), .dout(n14523));
  jand g14331(.dina(n14423), .dinb(n14421), .dout(n14524));
  jand g14332(.dina(n14424), .dinb(n14419), .dout(n14525));
  jor  g14333(.dina(n14525), .dinb(n14524), .dout(n14526));
  jand g14334(.dina(\a[56] ), .dinb(\a[50] ), .dout(n14527));
  jand g14335(.dina(\a[54] ), .dinb(\a[52] ), .dout(n14528));
  jor  g14336(.dina(n14528), .dinb(n14450), .dout(n14529));
  jnot g14337(.din(n14529), .dout(n14530));
  jand g14338(.dina(\a[55] ), .dinb(\a[52] ), .dout(n14531));
  jand g14339(.dina(n14531), .dinb(n14404), .dout(n14532));
  jor  g14340(.dina(n14532), .dinb(n14530), .dout(n14533));
  jxor g14341(.dina(n14533), .dinb(n14527), .dout(n14534));
  jnot g14342(.din(n14534), .dout(n14535));
  jand g14343(.dina(\a[59] ), .dinb(\a[47] ), .dout(n14536));
  jor  g14344(.dina(n14464), .dinb(n14078), .dout(n14537));
  jand g14345(.dina(\a[58] ), .dinb(\a[49] ), .dout(n14538));
  jand g14346(.dina(n14538), .dinb(n14385), .dout(n14539));
  jnot g14347(.din(n14539), .dout(n14540));
  jand g14348(.dina(n14540), .dinb(n14537), .dout(n14541));
  jxor g14349(.dina(n14541), .dinb(n14536), .dout(n14542));
  jxor g14350(.dina(n14542), .dinb(n14535), .dout(n14543));
  jxor g14351(.dina(n14543), .dinb(n14526), .dout(n14544));
  jand g14352(.dina(n14462), .dinb(n14460), .dout(n14545));
  jor  g14353(.dina(n14545), .dinb(n14465), .dout(n14546));
  jand g14354(.dina(n14471), .dinb(n14350), .dout(n14547));
  jor  g14355(.dina(n14547), .dinb(n14473), .dout(n14548));
  jnot g14356(.din(n14548), .dout(n14549));
  jxor g14357(.dina(n14549), .dinb(n14546), .dout(n14550));
  jand g14358(.dina(\a[62] ), .dinb(\a[44] ), .dout(n14551));
  jnot g14359(.din(n14551), .dout(n14552));
  jand g14360(.dina(\a[60] ), .dinb(\a[46] ), .dout(n14553));
  jor  g14361(.dina(n14553), .dinb(n14393), .dout(n14554));
  jand g14362(.dina(\a[61] ), .dinb(\a[46] ), .dout(n14555));
  jand g14363(.dina(n14555), .dinb(n14470), .dout(n14556));
  jnot g14364(.din(n14556), .dout(n14557));
  jand g14365(.dina(n14557), .dinb(n14554), .dout(n14558));
  jxor g14366(.dina(n14558), .dinb(n14552), .dout(n14559));
  jxor g14367(.dina(n14559), .dinb(n14550), .dout(n14560));
  jxor g14368(.dina(n14560), .dinb(n14544), .dout(n14561));
  jxor g14369(.dina(n14561), .dinb(n14523), .dout(n14562));
  jxor g14370(.dina(n14562), .dinb(n14518), .dout(n14563));
  jxor g14371(.dina(n14563), .dinb(n14495), .dout(n14564));
  jand g14372(.dina(n14486), .dinb(n14483), .dout(n14565));
  jnot g14373(.din(n14483), .dout(n14566));
  jnot g14374(.din(n14486), .dout(n14567));
  jand g14375(.dina(n14567), .dinb(n14566), .dout(n14568));
  jnot g14376(.din(n14568), .dout(n14569));
  jand g14377(.dina(n14491), .dinb(n14569), .dout(n14570));
  jor  g14378(.dina(n14570), .dinb(n14565), .dout(n14571));
  jxor g14379(.dina(n14571), .dinb(n14564), .dout(\asquared[107] ));
  jand g14380(.dina(n14517), .dinb(n14514), .dout(n14573));
  jand g14381(.dina(n14562), .dinb(n14518), .dout(n14574));
  jor  g14382(.dina(n14574), .dinb(n14573), .dout(n14575));
  jand g14383(.dina(n14507), .dinb(n14504), .dout(n14576));
  jnot g14384(.din(n14576), .dout(n14577));
  jor  g14385(.dina(n14513), .dinb(n14509), .dout(n14578));
  jand g14386(.dina(n14578), .dinb(n14577), .dout(n14579));
  jnot g14387(.din(n14579), .dout(n14580));
  jand g14388(.dina(\a[60] ), .dinb(\a[47] ), .dout(n14581));
  jor  g14389(.dina(n14581), .dinb(n14555), .dout(n14582));
  jand g14390(.dina(\a[61] ), .dinb(\a[47] ), .dout(n14583));
  jand g14391(.dina(n14583), .dinb(n14553), .dout(n14584));
  jnot g14392(.din(n14584), .dout(n14585));
  jand g14393(.dina(n14585), .dinb(n14582), .dout(n14586));
  jand g14394(.dina(n14529), .dinb(n14527), .dout(n14587));
  jor  g14395(.dina(n14587), .dinb(n14532), .dout(n14588));
  jxor g14396(.dina(n14588), .dinb(n14586), .dout(n14589));
  jand g14397(.dina(\a[57] ), .dinb(\a[50] ), .dout(n14590));
  jand g14398(.dina(\a[56] ), .dinb(\a[51] ), .dout(n14591));
  jor  g14399(.dina(n14591), .dinb(n14531), .dout(n14592));
  jnot g14400(.din(n14592), .dout(n14593));
  jand g14401(.dina(\a[56] ), .dinb(\a[52] ), .dout(n14594));
  jand g14402(.dina(n14594), .dinb(n14450), .dout(n14595));
  jor  g14403(.dina(n14595), .dinb(n14593), .dout(n14596));
  jxor g14404(.dina(n14596), .dinb(n14590), .dout(n14597));
  jand g14405(.dina(\a[62] ), .dinb(\a[45] ), .dout(n14598));
  jnot g14406(.din(n14598), .dout(n14599));
  jand g14407(.dina(\a[54] ), .dinb(n14497), .dout(n14600));
  jxor g14408(.dina(n14600), .dinb(n14599), .dout(n14601));
  jxor g14409(.dina(n14601), .dinb(n14597), .dout(n14602));
  jxor g14410(.dina(n14602), .dinb(n14589), .dout(n14603));
  jand g14411(.dina(n14541), .dinb(n14536), .dout(n14604));
  jor  g14412(.dina(n14604), .dinb(n14539), .dout(n14605));
  jand g14413(.dina(n14554), .dinb(n14551), .dout(n14606));
  jor  g14414(.dina(n14606), .dinb(n14556), .dout(n14607));
  jxor g14415(.dina(n14607), .dinb(n14605), .dout(n14608));
  jand g14416(.dina(\a[59] ), .dinb(\a[48] ), .dout(n14609));
  jand g14417(.dina(\a[63] ), .dinb(\a[44] ), .dout(n14610));
  jor  g14418(.dina(n14610), .dinb(n14538), .dout(n14611));
  jnot g14419(.din(n14611), .dout(n14612));
  jand g14420(.dina(\a[63] ), .dinb(\a[58] ), .dout(n14613));
  jand g14421(.dina(n14613), .dinb(n13215), .dout(n14614));
  jor  g14422(.dina(n14614), .dinb(n14612), .dout(n14615));
  jxor g14423(.dina(n14615), .dinb(n14609), .dout(n14616));
  jnot g14424(.din(n14616), .dout(n14617));
  jxor g14425(.dina(n14617), .dinb(n14608), .dout(n14618));
  jxor g14426(.dina(n14618), .dinb(n14603), .dout(n14619));
  jxor g14427(.dina(n14619), .dinb(n14580), .dout(n14620));
  jand g14428(.dina(n14560), .dinb(n14544), .dout(n14621));
  jand g14429(.dina(n14561), .dinb(n14523), .dout(n14622));
  jor  g14430(.dina(n14622), .dinb(n14621), .dout(n14623));
  jand g14431(.dina(n14500), .dinb(n14496), .dout(n14624));
  jand g14432(.dina(n14503), .dinb(n14501), .dout(n14625));
  jor  g14433(.dina(n14625), .dinb(n14624), .dout(n14626));
  jand g14434(.dina(n14548), .dinb(n14546), .dout(n14627));
  jnot g14435(.din(n14627), .dout(n14628));
  jnot g14436(.din(n14546), .dout(n14629));
  jand g14437(.dina(n14549), .dinb(n14629), .dout(n14630));
  jor  g14438(.dina(n14559), .dinb(n14630), .dout(n14631));
  jand g14439(.dina(n14631), .dinb(n14628), .dout(n14632));
  jnot g14440(.din(n14632), .dout(n14633));
  jxor g14441(.dina(n14633), .dinb(n14626), .dout(n14634));
  jand g14442(.dina(n14542), .dinb(n14535), .dout(n14635));
  jand g14443(.dina(n14543), .dinb(n14526), .dout(n14636));
  jor  g14444(.dina(n14636), .dinb(n14635), .dout(n14637));
  jxor g14445(.dina(n14637), .dinb(n14634), .dout(n14638));
  jxor g14446(.dina(n14638), .dinb(n14623), .dout(n14639));
  jxor g14447(.dina(n14639), .dinb(n14620), .dout(n14640));
  jxor g14448(.dina(n14640), .dinb(n14575), .dout(n14641));
  jand g14449(.dina(n14563), .dinb(n14495), .dout(n14642));
  jor  g14450(.dina(n14563), .dinb(n14495), .dout(n14643));
  jand g14451(.dina(n14571), .dinb(n14643), .dout(n14644));
  jor  g14452(.dina(n14644), .dinb(n14642), .dout(n14645));
  jxor g14453(.dina(n14645), .dinb(n14641), .dout(\asquared[108] ));
  jand g14454(.dina(n14638), .dinb(n14623), .dout(n14647));
  jand g14455(.dina(n14639), .dinb(n14620), .dout(n14648));
  jor  g14456(.dina(n14648), .dinb(n14647), .dout(n14649));
  jand g14457(.dina(n14618), .dinb(n14603), .dout(n14650));
  jand g14458(.dina(n14619), .dinb(n14580), .dout(n14651));
  jor  g14459(.dina(n14651), .dinb(n14650), .dout(n14652));
  jor  g14460(.dina(n14601), .dinb(n14597), .dout(n14653));
  jand g14461(.dina(n14602), .dinb(n14589), .dout(n14654));
  jnot g14462(.din(n14654), .dout(n14655));
  jand g14463(.dina(n14655), .dinb(n14653), .dout(n14656));
  jnot g14464(.din(n14656), .dout(n14657));
  jand g14465(.dina(\a[57] ), .dinb(\a[51] ), .dout(n14658));
  jand g14466(.dina(\a[55] ), .dinb(\a[53] ), .dout(n14659));
  jor  g14467(.dina(n14659), .dinb(n14594), .dout(n14660));
  jnot g14468(.din(n14660), .dout(n14661));
  jand g14469(.dina(\a[56] ), .dinb(\a[53] ), .dout(n14662));
  jand g14470(.dina(n14662), .dinb(n14531), .dout(n14663));
  jor  g14471(.dina(n14663), .dinb(n14661), .dout(n14664));
  jxor g14472(.dina(n14664), .dinb(n14658), .dout(n14665));
  jnot g14473(.din(n14665), .dout(n14666));
  jnot g14474(.din(n14605), .dout(n14667));
  jnot g14475(.din(n14607), .dout(n14668));
  jand g14476(.dina(n14668), .dinb(n14667), .dout(n14669));
  jnot g14477(.din(n14669), .dout(n14670));
  jand g14478(.dina(n14607), .dinb(n14605), .dout(n14671));
  jor  g14479(.dina(n14617), .dinb(n14671), .dout(n14672));
  jand g14480(.dina(n14672), .dinb(n14670), .dout(n14673));
  jxor g14481(.dina(n14673), .dinb(n14666), .dout(n14674));
  jxor g14482(.dina(n14674), .dinb(n14657), .dout(n14675));
  jxor g14483(.dina(n14675), .dinb(n14652), .dout(n14676));
  jand g14484(.dina(n14592), .dinb(n14590), .dout(n14677));
  jor  g14485(.dina(n14677), .dinb(n14595), .dout(n14678));
  jand g14486(.dina(n14599), .dinb(n14497), .dout(n14679));
  jor  g14487(.dina(n14679), .dinb(n5841), .dout(n14680));
  jnot g14488(.din(n14680), .dout(n14681));
  jxor g14489(.dina(n14681), .dinb(n14678), .dout(n14682));
  jand g14490(.dina(n14611), .dinb(n14609), .dout(n14683));
  jor  g14491(.dina(n14683), .dinb(n14614), .dout(n14684));
  jxor g14492(.dina(n14684), .dinb(n14682), .dout(n14685));
  jand g14493(.dina(n14633), .dinb(n14626), .dout(n14686));
  jand g14494(.dina(n14637), .dinb(n14634), .dout(n14687));
  jor  g14495(.dina(n14687), .dinb(n14686), .dout(n14688));
  jxor g14496(.dina(n14688), .dinb(n14685), .dout(n14689));
  jand g14497(.dina(\a[60] ), .dinb(\a[48] ), .dout(n14690));
  jand g14498(.dina(\a[59] ), .dinb(\a[49] ), .dout(n14691));
  jand g14499(.dina(\a[58] ), .dinb(\a[50] ), .dout(n14692));
  jor  g14500(.dina(n14692), .dinb(n14691), .dout(n14693));
  jnot g14501(.din(n14693), .dout(n14694));
  jand g14502(.dina(\a[59] ), .dinb(\a[50] ), .dout(n14695));
  jand g14503(.dina(n14695), .dinb(n14538), .dout(n14696));
  jor  g14504(.dina(n14696), .dinb(n14694), .dout(n14697));
  jxor g14505(.dina(n14697), .dinb(n14690), .dout(n14698));
  jnot g14506(.din(n14698), .dout(n14699));
  jand g14507(.dina(\a[63] ), .dinb(\a[45] ), .dout(n14700));
  jand g14508(.dina(\a[62] ), .dinb(\a[46] ), .dout(n14701));
  jor  g14509(.dina(n14701), .dinb(n14583), .dout(n14702));
  jnot g14510(.din(n14702), .dout(n14703));
  jand g14511(.dina(\a[62] ), .dinb(\a[47] ), .dout(n14704));
  jand g14512(.dina(n14704), .dinb(n14555), .dout(n14705));
  jor  g14513(.dina(n14705), .dinb(n14703), .dout(n14706));
  jxor g14514(.dina(n14706), .dinb(n14700), .dout(n14707));
  jnot g14515(.din(n14707), .dout(n14708));
  jand g14516(.dina(n14588), .dinb(n14586), .dout(n14709));
  jor  g14517(.dina(n14709), .dinb(n14584), .dout(n14710));
  jxor g14518(.dina(n14710), .dinb(n14708), .dout(n14711));
  jxor g14519(.dina(n14711), .dinb(n14699), .dout(n14712));
  jxor g14520(.dina(n14712), .dinb(n14689), .dout(n14713));
  jxor g14521(.dina(n14713), .dinb(n14676), .dout(n14714));
  jxor g14522(.dina(n14714), .dinb(n14649), .dout(n14715));
  jand g14523(.dina(n14640), .dinb(n14575), .dout(n14716));
  jnot g14524(.din(n14575), .dout(n14717));
  jnot g14525(.din(n14640), .dout(n14718));
  jand g14526(.dina(n14718), .dinb(n14717), .dout(n14719));
  jnot g14527(.din(n14719), .dout(n14720));
  jand g14528(.dina(n14645), .dinb(n14720), .dout(n14721));
  jor  g14529(.dina(n14721), .dinb(n14716), .dout(n14722));
  jxor g14530(.dina(n14722), .dinb(n14715), .dout(\asquared[109] ));
  jand g14531(.dina(n14675), .dinb(n14652), .dout(n14724));
  jand g14532(.dina(n14713), .dinb(n14676), .dout(n14725));
  jor  g14533(.dina(n14725), .dinb(n14724), .dout(n14726));
  jand g14534(.dina(n14710), .dinb(n14708), .dout(n14727));
  jand g14535(.dina(n14711), .dinb(n14699), .dout(n14728));
  jor  g14536(.dina(n14728), .dinb(n14727), .dout(n14729));
  jand g14537(.dina(n14681), .dinb(n14678), .dout(n14730));
  jand g14538(.dina(n14684), .dinb(n14682), .dout(n14731));
  jor  g14539(.dina(n14731), .dinb(n14730), .dout(n14732));
  jnot g14540(.din(n14732), .dout(n14733));
  jnot g14541(.din(n14704), .dout(n14734));
  jand g14542(.dina(\a[55] ), .dinb(n5841), .dout(n14735));
  jxor g14543(.dina(n14735), .dinb(n14734), .dout(n14736));
  jxor g14544(.dina(n14736), .dinb(n14733), .dout(n14737));
  jxor g14545(.dina(n14737), .dinb(n14729), .dout(n14738));
  jand g14546(.dina(n14688), .dinb(n14685), .dout(n14739));
  jand g14547(.dina(n14712), .dinb(n14689), .dout(n14740));
  jor  g14548(.dina(n14740), .dinb(n14739), .dout(n14741));
  jxor g14549(.dina(n14741), .dinb(n14738), .dout(n14742));
  jand g14550(.dina(\a[63] ), .dinb(\a[46] ), .dout(n14743));
  jand g14551(.dina(n14660), .dinb(n14658), .dout(n14744));
  jor  g14552(.dina(n14744), .dinb(n14663), .dout(n14745));
  jxor g14553(.dina(n14745), .dinb(n14743), .dout(n14746));
  jand g14554(.dina(n14693), .dinb(n14690), .dout(n14747));
  jor  g14555(.dina(n14747), .dinb(n14696), .dout(n14748));
  jxor g14556(.dina(n14748), .dinb(n14746), .dout(n14749));
  jand g14557(.dina(n14673), .dinb(n14666), .dout(n14750));
  jand g14558(.dina(n14674), .dinb(n14657), .dout(n14751));
  jor  g14559(.dina(n14751), .dinb(n14750), .dout(n14752));
  jxor g14560(.dina(n14752), .dinb(n14749), .dout(n14753));
  jand g14561(.dina(\a[58] ), .dinb(\a[51] ), .dout(n14754));
  jand g14562(.dina(\a[57] ), .dinb(\a[52] ), .dout(n14755));
  jor  g14563(.dina(n14755), .dinb(n14662), .dout(n14756));
  jnot g14564(.din(n14756), .dout(n14757));
  jand g14565(.dina(\a[57] ), .dinb(\a[53] ), .dout(n14758));
  jand g14566(.dina(n14758), .dinb(n14594), .dout(n14759));
  jor  g14567(.dina(n14759), .dinb(n14757), .dout(n14760));
  jxor g14568(.dina(n14760), .dinb(n14754), .dout(n14761));
  jnot g14569(.din(n14761), .dout(n14762));
  jand g14570(.dina(\a[61] ), .dinb(\a[48] ), .dout(n14763));
  jand g14571(.dina(\a[60] ), .dinb(\a[49] ), .dout(n14764));
  jor  g14572(.dina(n14764), .dinb(n14695), .dout(n14765));
  jnot g14573(.din(n14765), .dout(n14766));
  jand g14574(.dina(\a[60] ), .dinb(\a[50] ), .dout(n14767));
  jand g14575(.dina(n14767), .dinb(n14691), .dout(n14768));
  jor  g14576(.dina(n14768), .dinb(n14766), .dout(n14769));
  jxor g14577(.dina(n14769), .dinb(n14763), .dout(n14770));
  jnot g14578(.din(n14770), .dout(n14771));
  jand g14579(.dina(n14702), .dinb(n14700), .dout(n14772));
  jor  g14580(.dina(n14772), .dinb(n14705), .dout(n14773));
  jxor g14581(.dina(n14773), .dinb(n14771), .dout(n14774));
  jxor g14582(.dina(n14774), .dinb(n14762), .dout(n14775));
  jxor g14583(.dina(n14775), .dinb(n14753), .dout(n14776));
  jxor g14584(.dina(n14776), .dinb(n14742), .dout(n14777));
  jxor g14585(.dina(n14777), .dinb(n14726), .dout(n14778));
  jand g14586(.dina(n14714), .dinb(n14649), .dout(n14779));
  jnot g14587(.din(n14649), .dout(n14780));
  jnot g14588(.din(n14714), .dout(n14781));
  jand g14589(.dina(n14781), .dinb(n14780), .dout(n14782));
  jnot g14590(.din(n14782), .dout(n14783));
  jand g14591(.dina(n14722), .dinb(n14783), .dout(n14784));
  jor  g14592(.dina(n14784), .dinb(n14779), .dout(n14785));
  jxor g14593(.dina(n14785), .dinb(n14778), .dout(\asquared[110] ));
  jand g14594(.dina(n14741), .dinb(n14738), .dout(n14787));
  jand g14595(.dina(n14776), .dinb(n14742), .dout(n14788));
  jor  g14596(.dina(n14788), .dinb(n14787), .dout(n14789));
  jand g14597(.dina(n14773), .dinb(n14771), .dout(n14790));
  jand g14598(.dina(n14774), .dinb(n14762), .dout(n14791));
  jor  g14599(.dina(n14791), .dinb(n14790), .dout(n14792));
  jand g14600(.dina(n14756), .dinb(n14754), .dout(n14793));
  jor  g14601(.dina(n14793), .dinb(n14759), .dout(n14794));
  jand g14602(.dina(n14765), .dinb(n14763), .dout(n14795));
  jor  g14603(.dina(n14795), .dinb(n14768), .dout(n14796));
  jxor g14604(.dina(n14796), .dinb(n14794), .dout(n14797));
  jand g14605(.dina(\a[61] ), .dinb(\a[49] ), .dout(n14798));
  jand g14606(.dina(\a[59] ), .dinb(\a[51] ), .dout(n14799));
  jor  g14607(.dina(n14799), .dinb(n14767), .dout(n14800));
  jnot g14608(.din(n14800), .dout(n14801));
  jand g14609(.dina(\a[60] ), .dinb(\a[51] ), .dout(n14802));
  jand g14610(.dina(n14802), .dinb(n14695), .dout(n14803));
  jor  g14611(.dina(n14803), .dinb(n14801), .dout(n14804));
  jxor g14612(.dina(n14804), .dinb(n14798), .dout(n14805));
  jnot g14613(.din(n14805), .dout(n14806));
  jxor g14614(.dina(n14806), .dinb(n14797), .dout(n14807));
  jxor g14615(.dina(n14807), .dinb(n14792), .dout(n14808));
  jnot g14616(.din(n14808), .dout(n14809));
  jor  g14617(.dina(n14736), .dinb(n14733), .dout(n14810));
  jand g14618(.dina(n14737), .dinb(n14729), .dout(n14811));
  jnot g14619(.din(n14811), .dout(n14812));
  jand g14620(.dina(n14812), .dinb(n14810), .dout(n14813));
  jxor g14621(.dina(n14813), .dinb(n14809), .dout(n14814));
  jand g14622(.dina(n14745), .dinb(n14743), .dout(n14815));
  jand g14623(.dina(n14748), .dinb(n14746), .dout(n14816));
  jor  g14624(.dina(n14816), .dinb(n14815), .dout(n14817));
  jnot g14625(.din(\a[55] ), .dout(n14818));
  jand g14626(.dina(n14734), .dinb(n5841), .dout(n14819));
  jor  g14627(.dina(n14819), .dinb(n14818), .dout(n14820));
  jnot g14628(.din(n14820), .dout(n14821));
  jand g14629(.dina(\a[62] ), .dinb(\a[48] ), .dout(n14822));
  jand g14630(.dina(\a[63] ), .dinb(\a[47] ), .dout(n14823));
  jor  g14631(.dina(n14823), .dinb(n14822), .dout(n14824));
  jand g14632(.dina(\a[63] ), .dinb(\a[48] ), .dout(n14825));
  jand g14633(.dina(n14825), .dinb(n14704), .dout(n14826));
  jnot g14634(.din(n14826), .dout(n14827));
  jand g14635(.dina(n14827), .dinb(n14824), .dout(n14828));
  jxor g14636(.dina(n14828), .dinb(n14821), .dout(n14829));
  jnot g14637(.din(n14829), .dout(n14830));
  jand g14638(.dina(\a[58] ), .dinb(\a[52] ), .dout(n14831));
  jand g14639(.dina(\a[56] ), .dinb(\a[54] ), .dout(n14832));
  jor  g14640(.dina(n14832), .dinb(n14758), .dout(n14833));
  jnot g14641(.din(n14833), .dout(n14834));
  jand g14642(.dina(\a[57] ), .dinb(\a[54] ), .dout(n14835));
  jand g14643(.dina(n14835), .dinb(n14662), .dout(n14836));
  jor  g14644(.dina(n14836), .dinb(n14834), .dout(n14837));
  jxor g14645(.dina(n14837), .dinb(n14831), .dout(n14838));
  jxor g14646(.dina(n14838), .dinb(n14830), .dout(n14839));
  jxor g14647(.dina(n14839), .dinb(n14817), .dout(n14840));
  jand g14648(.dina(n14752), .dinb(n14749), .dout(n14841));
  jand g14649(.dina(n14775), .dinb(n14753), .dout(n14842));
  jor  g14650(.dina(n14842), .dinb(n14841), .dout(n14843));
  jxor g14651(.dina(n14843), .dinb(n14840), .dout(n14844));
  jxor g14652(.dina(n14844), .dinb(n14814), .dout(n14845));
  jxor g14653(.dina(n14845), .dinb(n14789), .dout(n14846));
  jand g14654(.dina(n14777), .dinb(n14726), .dout(n14847));
  jor  g14655(.dina(n14777), .dinb(n14726), .dout(n14848));
  jand g14656(.dina(n14785), .dinb(n14848), .dout(n14849));
  jor  g14657(.dina(n14849), .dinb(n14847), .dout(n14850));
  jxor g14658(.dina(n14850), .dinb(n14846), .dout(\asquared[111] ));
  jand g14659(.dina(n14843), .dinb(n14840), .dout(n14852));
  jand g14660(.dina(n14844), .dinb(n14814), .dout(n14853));
  jor  g14661(.dina(n14853), .dinb(n14852), .dout(n14854));
  jand g14662(.dina(n14800), .dinb(n14798), .dout(n14855));
  jor  g14663(.dina(n14855), .dinb(n14803), .dout(n14856));
  jand g14664(.dina(n14833), .dinb(n14831), .dout(n14857));
  jor  g14665(.dina(n14857), .dinb(n14836), .dout(n14858));
  jxor g14666(.dina(n14858), .dinb(n14856), .dout(n14859));
  jand g14667(.dina(n14828), .dinb(n14821), .dout(n14860));
  jor  g14668(.dina(n14860), .dinb(n14826), .dout(n14861));
  jxor g14669(.dina(n14861), .dinb(n14859), .dout(n14862));
  jnot g14670(.din(n14794), .dout(n14863));
  jnot g14671(.din(n14796), .dout(n14864));
  jand g14672(.dina(n14864), .dinb(n14863), .dout(n14865));
  jnot g14673(.din(n14865), .dout(n14866));
  jand g14674(.dina(n14796), .dinb(n14794), .dout(n14867));
  jor  g14675(.dina(n14806), .dinb(n14867), .dout(n14868));
  jand g14676(.dina(n14868), .dinb(n14866), .dout(n14869));
  jxor g14677(.dina(n14869), .dinb(n14862), .dout(n14870));
  jnot g14678(.din(n14870), .dout(n14871));
  jor  g14679(.dina(n14838), .dinb(n14830), .dout(n14872));
  jand g14680(.dina(n14839), .dinb(n14817), .dout(n14873));
  jnot g14681(.din(n14873), .dout(n14874));
  jand g14682(.dina(n14874), .dinb(n14872), .dout(n14875));
  jxor g14683(.dina(n14875), .dinb(n14871), .dout(n14876));
  jand g14684(.dina(n14807), .dinb(n14792), .dout(n14877));
  jnot g14685(.din(n14877), .dout(n14878));
  jor  g14686(.dina(n14813), .dinb(n14809), .dout(n14879));
  jand g14687(.dina(n14879), .dinb(n14878), .dout(n14880));
  jnot g14688(.din(n14880), .dout(n14881));
  jand g14689(.dina(\a[59] ), .dinb(\a[52] ), .dout(n14882));
  jand g14690(.dina(\a[58] ), .dinb(\a[53] ), .dout(n14883));
  jor  g14691(.dina(n14883), .dinb(n14835), .dout(n14884));
  jnot g14692(.din(n14884), .dout(n14885));
  jand g14693(.dina(\a[58] ), .dinb(\a[54] ), .dout(n14886));
  jand g14694(.dina(n14886), .dinb(n14758), .dout(n14887));
  jor  g14695(.dina(n14887), .dinb(n14885), .dout(n14888));
  jxor g14696(.dina(n14888), .dinb(n14882), .dout(n14889));
  jnot g14697(.din(n14889), .dout(n14890));
  jand g14698(.dina(\a[62] ), .dinb(\a[49] ), .dout(n14891));
  jnot g14699(.din(n14891), .dout(n14892));
  jand g14700(.dina(\a[56] ), .dinb(n14818), .dout(n14893));
  jxor g14701(.dina(n14893), .dinb(n14892), .dout(n14894));
  jnot g14702(.din(n14894), .dout(n14895));
  jand g14703(.dina(\a[61] ), .dinb(\a[50] ), .dout(n14896));
  jor  g14704(.dina(n14896), .dinb(n14802), .dout(n14897));
  jand g14705(.dina(\a[61] ), .dinb(\a[51] ), .dout(n14898));
  jand g14706(.dina(n14898), .dinb(n14767), .dout(n14899));
  jnot g14707(.din(n14899), .dout(n14900));
  jand g14708(.dina(n14900), .dinb(n14897), .dout(n14901));
  jxor g14709(.dina(n14901), .dinb(n14825), .dout(n14902));
  jxor g14710(.dina(n14902), .dinb(n14895), .dout(n14903));
  jxor g14711(.dina(n14903), .dinb(n14890), .dout(n14904));
  jxor g14712(.dina(n14904), .dinb(n14881), .dout(n14905));
  jxor g14713(.dina(n14905), .dinb(n14876), .dout(n14906));
  jxor g14714(.dina(n14906), .dinb(n14854), .dout(n14907));
  jand g14715(.dina(n14845), .dinb(n14789), .dout(n14908));
  jnot g14716(.din(n14789), .dout(n14909));
  jnot g14717(.din(n14845), .dout(n14910));
  jand g14718(.dina(n14910), .dinb(n14909), .dout(n14911));
  jnot g14719(.din(n14911), .dout(n14912));
  jand g14720(.dina(n14850), .dinb(n14912), .dout(n14913));
  jor  g14721(.dina(n14913), .dinb(n14908), .dout(n14914));
  jxor g14722(.dina(n14914), .dinb(n14907), .dout(\asquared[112] ));
  jand g14723(.dina(n14904), .dinb(n14881), .dout(n14916));
  jand g14724(.dina(n14905), .dinb(n14876), .dout(n14917));
  jor  g14725(.dina(n14917), .dinb(n14916), .dout(n14918));
  jand g14726(.dina(n14869), .dinb(n14862), .dout(n14919));
  jnot g14727(.din(n14919), .dout(n14920));
  jor  g14728(.dina(n14875), .dinb(n14871), .dout(n14921));
  jand g14729(.dina(n14921), .dinb(n14920), .dout(n14922));
  jnot g14730(.din(n14922), .dout(n14923));
  jand g14731(.dina(\a[59] ), .dinb(\a[53] ), .dout(n14924));
  jand g14732(.dina(\a[57] ), .dinb(\a[55] ), .dout(n14925));
  jor  g14733(.dina(n14925), .dinb(n14886), .dout(n14926));
  jnot g14734(.din(n14926), .dout(n14927));
  jand g14735(.dina(\a[58] ), .dinb(\a[55] ), .dout(n14928));
  jand g14736(.dina(n14928), .dinb(n14835), .dout(n14929));
  jor  g14737(.dina(n14929), .dinb(n14927), .dout(n14930));
  jxor g14738(.dina(n14930), .dinb(n14924), .dout(n14931));
  jnot g14739(.din(n14931), .dout(n14932));
  jand g14740(.dina(n14901), .dinb(n14825), .dout(n14933));
  jor  g14741(.dina(n14933), .dinb(n14899), .dout(n14934));
  jand g14742(.dina(\a[60] ), .dinb(\a[52] ), .dout(n14935));
  jor  g14743(.dina(n14935), .dinb(n14898), .dout(n14936));
  jand g14744(.dina(\a[61] ), .dinb(\a[52] ), .dout(n14937));
  jand g14745(.dina(n14937), .dinb(n14802), .dout(n14938));
  jnot g14746(.din(n14938), .dout(n14939));
  jand g14747(.dina(n14939), .dinb(n14936), .dout(n14940));
  jand g14748(.dina(\a[63] ), .dinb(\a[49] ), .dout(n14941));
  jand g14749(.dina(n14941), .dinb(n14936), .dout(n14942));
  jnot g14750(.din(n14942), .dout(n14943));
  jand g14751(.dina(n14943), .dinb(n14940), .dout(n14944));
  jnot g14752(.din(n14940), .dout(n14945));
  jand g14753(.dina(n14941), .dinb(n14945), .dout(n14946));
  jor  g14754(.dina(n14946), .dinb(n14944), .dout(n14947));
  jxor g14755(.dina(n14947), .dinb(n14934), .dout(n14948));
  jxor g14756(.dina(n14948), .dinb(n14932), .dout(n14949));
  jxor g14757(.dina(n14949), .dinb(n14923), .dout(n14950));
  jnot g14758(.din(\a[56] ), .dout(n14951));
  jand g14759(.dina(n14892), .dinb(n14818), .dout(n14952));
  jor  g14760(.dina(n14952), .dinb(n14951), .dout(n14953));
  jnot g14761(.din(n14953), .dout(n14954));
  jand g14762(.dina(\a[62] ), .dinb(\a[50] ), .dout(n14955));
  jxor g14763(.dina(n14955), .dinb(n14954), .dout(n14956));
  jand g14764(.dina(n14884), .dinb(n14882), .dout(n14957));
  jor  g14765(.dina(n14957), .dinb(n14887), .dout(n14958));
  jxor g14766(.dina(n14958), .dinb(n14956), .dout(n14959));
  jand g14767(.dina(n14858), .dinb(n14856), .dout(n14960));
  jand g14768(.dina(n14861), .dinb(n14859), .dout(n14961));
  jor  g14769(.dina(n14961), .dinb(n14960), .dout(n14962));
  jor  g14770(.dina(n14902), .dinb(n14895), .dout(n14963));
  jand g14771(.dina(n14902), .dinb(n14895), .dout(n14964));
  jor  g14772(.dina(n14964), .dinb(n14890), .dout(n14965));
  jand g14773(.dina(n14965), .dinb(n14963), .dout(n14966));
  jxor g14774(.dina(n14966), .dinb(n14962), .dout(n14967));
  jxor g14775(.dina(n14967), .dinb(n14959), .dout(n14968));
  jxor g14776(.dina(n14968), .dinb(n14950), .dout(n14969));
  jxor g14777(.dina(n14969), .dinb(n14918), .dout(n14970));
  jand g14778(.dina(n14906), .dinb(n14854), .dout(n14971));
  jor  g14779(.dina(n14906), .dinb(n14854), .dout(n14972));
  jand g14780(.dina(n14914), .dinb(n14972), .dout(n14973));
  jor  g14781(.dina(n14973), .dinb(n14971), .dout(n14974));
  jxor g14782(.dina(n14974), .dinb(n14970), .dout(\asquared[113] ));
  jand g14783(.dina(n14949), .dinb(n14923), .dout(n14976));
  jand g14784(.dina(n14968), .dinb(n14950), .dout(n14977));
  jor  g14785(.dina(n14977), .dinb(n14976), .dout(n14978));
  jand g14786(.dina(n14955), .dinb(n14954), .dout(n14979));
  jand g14787(.dina(n14958), .dinb(n14956), .dout(n14980));
  jor  g14788(.dina(n14980), .dinb(n14979), .dout(n14981));
  jand g14789(.dina(\a[60] ), .dinb(\a[53] ), .dout(n14982));
  jor  g14790(.dina(n14982), .dinb(n14937), .dout(n14983));
  jand g14791(.dina(\a[61] ), .dinb(\a[53] ), .dout(n14984));
  jand g14792(.dina(n14984), .dinb(n14935), .dout(n14985));
  jnot g14793(.din(n14985), .dout(n14986));
  jand g14794(.dina(n14986), .dinb(n14983), .dout(n14987));
  jand g14795(.dina(n14926), .dinb(n14924), .dout(n14988));
  jor  g14796(.dina(n14988), .dinb(n14929), .dout(n14989));
  jxor g14797(.dina(n14989), .dinb(n14987), .dout(n14990));
  jxor g14798(.dina(n14990), .dinb(n14981), .dout(n14991));
  jand g14799(.dina(n14947), .dinb(n14934), .dout(n14992));
  jand g14800(.dina(n14948), .dinb(n14932), .dout(n14993));
  jor  g14801(.dina(n14993), .dinb(n14992), .dout(n14994));
  jxor g14802(.dina(n14994), .dinb(n14991), .dout(n14995));
  jand g14803(.dina(n14966), .dinb(n14962), .dout(n14996));
  jand g14804(.dina(n14967), .dinb(n14959), .dout(n14997));
  jor  g14805(.dina(n14997), .dinb(n14996), .dout(n14998));
  jand g14806(.dina(\a[63] ), .dinb(\a[50] ), .dout(n14999));
  jand g14807(.dina(\a[59] ), .dinb(\a[54] ), .dout(n15000));
  jor  g14808(.dina(n15000), .dinb(n14928), .dout(n15001));
  jnot g14809(.din(n15001), .dout(n15002));
  jand g14810(.dina(\a[59] ), .dinb(\a[55] ), .dout(n15003));
  jand g14811(.dina(n15003), .dinb(n14886), .dout(n15004));
  jor  g14812(.dina(n15004), .dinb(n15002), .dout(n15005));
  jxor g14813(.dina(n15005), .dinb(n14999), .dout(n15006));
  jand g14814(.dina(n14943), .dinb(n14939), .dout(n15007));
  jxor g14815(.dina(n15007), .dinb(n15006), .dout(n15008));
  jnot g14816(.din(n15008), .dout(n15009));
  jand g14817(.dina(\a[62] ), .dinb(\a[51] ), .dout(n15010));
  jnot g14818(.din(n15010), .dout(n15011));
  jand g14819(.dina(\a[57] ), .dinb(n14951), .dout(n15012));
  jxor g14820(.dina(n15012), .dinb(n15011), .dout(n15013));
  jxor g14821(.dina(n15013), .dinb(n15009), .dout(n15014));
  jxor g14822(.dina(n15014), .dinb(n14998), .dout(n15015));
  jxor g14823(.dina(n15015), .dinb(n14995), .dout(n15016));
  jxor g14824(.dina(n15016), .dinb(n14978), .dout(n15017));
  jand g14825(.dina(n14969), .dinb(n14918), .dout(n15018));
  jnot g14826(.din(n14918), .dout(n15019));
  jnot g14827(.din(n14969), .dout(n15020));
  jand g14828(.dina(n15020), .dinb(n15019), .dout(n15021));
  jnot g14829(.din(n15021), .dout(n15022));
  jand g14830(.dina(n14974), .dinb(n15022), .dout(n15023));
  jor  g14831(.dina(n15023), .dinb(n15018), .dout(n15024));
  jxor g14832(.dina(n15024), .dinb(n15017), .dout(\asquared[114] ));
  jand g14833(.dina(n15014), .dinb(n14998), .dout(n15026));
  jand g14834(.dina(n15015), .dinb(n14995), .dout(n15027));
  jor  g14835(.dina(n15027), .dinb(n15026), .dout(n15028));
  jnot g14836(.din(\a[57] ), .dout(n15029));
  jand g14837(.dina(n15011), .dinb(n14951), .dout(n15030));
  jor  g14838(.dina(n15030), .dinb(n15029), .dout(n15031));
  jnot g14839(.din(n15031), .dout(n15032));
  jand g14840(.dina(n15001), .dinb(n14999), .dout(n15033));
  jor  g14841(.dina(n15033), .dinb(n15004), .dout(n15034));
  jxor g14842(.dina(n15034), .dinb(n15032), .dout(n15035));
  jand g14843(.dina(n14989), .dinb(n14987), .dout(n15036));
  jor  g14844(.dina(n15036), .dinb(n14985), .dout(n15037));
  jxor g14845(.dina(n15037), .dinb(n15035), .dout(n15038));
  jand g14846(.dina(n14990), .dinb(n14981), .dout(n15039));
  jand g14847(.dina(n14994), .dinb(n14991), .dout(n15040));
  jor  g14848(.dina(n15040), .dinb(n15039), .dout(n15041));
  jxor g14849(.dina(n15041), .dinb(n15038), .dout(n15042));
  jor  g14850(.dina(n15007), .dinb(n15006), .dout(n15043));
  jor  g14851(.dina(n15013), .dinb(n15009), .dout(n15044));
  jand g14852(.dina(n15044), .dinb(n15043), .dout(n15045));
  jnot g14853(.din(n15045), .dout(n15046));
  jand g14854(.dina(\a[60] ), .dinb(\a[54] ), .dout(n15047));
  jand g14855(.dina(\a[58] ), .dinb(\a[56] ), .dout(n15048));
  jor  g14856(.dina(n15048), .dinb(n15003), .dout(n15049));
  jnot g14857(.din(n15049), .dout(n15050));
  jand g14858(.dina(\a[59] ), .dinb(\a[56] ), .dout(n15051));
  jand g14859(.dina(n15051), .dinb(n14928), .dout(n15052));
  jor  g14860(.dina(n15052), .dinb(n15050), .dout(n15053));
  jxor g14861(.dina(n15053), .dinb(n15047), .dout(n15054));
  jnot g14862(.din(n15054), .dout(n15055));
  jand g14863(.dina(\a[63] ), .dinb(\a[51] ), .dout(n15056));
  jand g14864(.dina(\a[62] ), .dinb(\a[52] ), .dout(n15057));
  jor  g14865(.dina(n15057), .dinb(n14984), .dout(n15058));
  jand g14866(.dina(\a[62] ), .dinb(\a[53] ), .dout(n15059));
  jand g14867(.dina(n15059), .dinb(n14937), .dout(n15060));
  jnot g14868(.din(n15060), .dout(n15061));
  jand g14869(.dina(n15061), .dinb(n15058), .dout(n15062));
  jxor g14870(.dina(n15062), .dinb(n15056), .dout(n15063));
  jxor g14871(.dina(n15063), .dinb(n15055), .dout(n15064));
  jxor g14872(.dina(n15064), .dinb(n15046), .dout(n15065));
  jxor g14873(.dina(n15065), .dinb(n15042), .dout(n15066));
  jxor g14874(.dina(n15066), .dinb(n15028), .dout(n15067));
  jand g14875(.dina(n15016), .dinb(n14978), .dout(n15068));
  jnot g14876(.din(n14978), .dout(n15069));
  jnot g14877(.din(n15016), .dout(n15070));
  jand g14878(.dina(n15070), .dinb(n15069), .dout(n15071));
  jnot g14879(.din(n15071), .dout(n15072));
  jand g14880(.dina(n15024), .dinb(n15072), .dout(n15073));
  jor  g14881(.dina(n15073), .dinb(n15068), .dout(n15074));
  jxor g14882(.dina(n15074), .dinb(n15067), .dout(\asquared[115] ));
  jand g14883(.dina(n15041), .dinb(n15038), .dout(n15076));
  jand g14884(.dina(n15065), .dinb(n15042), .dout(n15077));
  jor  g14885(.dina(n15077), .dinb(n15076), .dout(n15078));
  jand g14886(.dina(n15034), .dinb(n15032), .dout(n15079));
  jand g14887(.dina(n15037), .dinb(n15035), .dout(n15080));
  jor  g14888(.dina(n15080), .dinb(n15079), .dout(n15081));
  jand g14889(.dina(\a[61] ), .dinb(\a[54] ), .dout(n15082));
  jand g14890(.dina(\a[60] ), .dinb(\a[55] ), .dout(n15083));
  jor  g14891(.dina(n15083), .dinb(n15051), .dout(n15084));
  jnot g14892(.din(n15084), .dout(n15085));
  jand g14893(.dina(\a[60] ), .dinb(\a[56] ), .dout(n15086));
  jand g14894(.dina(n15086), .dinb(n15003), .dout(n15087));
  jor  g14895(.dina(n15087), .dinb(n15085), .dout(n15088));
  jxor g14896(.dina(n15088), .dinb(n15082), .dout(n15089));
  jnot g14897(.din(n15059), .dout(n15090));
  jand g14898(.dina(\a[58] ), .dinb(n15029), .dout(n15091));
  jxor g14899(.dina(n15091), .dinb(n15090), .dout(n15092));
  jxor g14900(.dina(n15092), .dinb(n15089), .dout(n15093));
  jxor g14901(.dina(n15093), .dinb(n15081), .dout(n15094));
  jand g14902(.dina(n15062), .dinb(n15056), .dout(n15095));
  jor  g14903(.dina(n15095), .dinb(n15060), .dout(n15096));
  jand g14904(.dina(\a[63] ), .dinb(\a[52] ), .dout(n15097));
  jand g14905(.dina(n15049), .dinb(n15047), .dout(n15098));
  jor  g14906(.dina(n15098), .dinb(n15052), .dout(n15099));
  jxor g14907(.dina(n15099), .dinb(n15097), .dout(n15100));
  jxor g14908(.dina(n15100), .dinb(n15096), .dout(n15101));
  jand g14909(.dina(n15063), .dinb(n15055), .dout(n15102));
  jand g14910(.dina(n15064), .dinb(n15046), .dout(n15103));
  jor  g14911(.dina(n15103), .dinb(n15102), .dout(n15104));
  jxor g14912(.dina(n15104), .dinb(n15101), .dout(n15105));
  jxor g14913(.dina(n15105), .dinb(n15094), .dout(n15106));
  jxor g14914(.dina(n15106), .dinb(n15078), .dout(n15107));
  jand g14915(.dina(n15066), .dinb(n15028), .dout(n15108));
  jnot g14916(.din(n15028), .dout(n15109));
  jnot g14917(.din(n15066), .dout(n15110));
  jand g14918(.dina(n15110), .dinb(n15109), .dout(n15111));
  jnot g14919(.din(n15111), .dout(n15112));
  jand g14920(.dina(n15074), .dinb(n15112), .dout(n15113));
  jor  g14921(.dina(n15113), .dinb(n15108), .dout(n15114));
  jxor g14922(.dina(n15114), .dinb(n15107), .dout(\asquared[116] ));
  jor  g14923(.dina(n15092), .dinb(n15089), .dout(n15116));
  jand g14924(.dina(n15093), .dinb(n15081), .dout(n15117));
  jnot g14925(.din(n15117), .dout(n15118));
  jand g14926(.dina(n15118), .dinb(n15116), .dout(n15119));
  jnot g14927(.din(n15119), .dout(n15120));
  jand g14928(.dina(n15099), .dinb(n15097), .dout(n15121));
  jand g14929(.dina(n15100), .dinb(n15096), .dout(n15122));
  jor  g14930(.dina(n15122), .dinb(n15121), .dout(n15123));
  jxor g14931(.dina(n15123), .dinb(n15120), .dout(n15124));
  jand g14932(.dina(\a[62] ), .dinb(\a[54] ), .dout(n15125));
  jand g14933(.dina(\a[63] ), .dinb(\a[53] ), .dout(n15126));
  jor  g14934(.dina(n15126), .dinb(n15125), .dout(n15127));
  jand g14935(.dina(\a[63] ), .dinb(\a[54] ), .dout(n15128));
  jand g14936(.dina(n15128), .dinb(n15059), .dout(n15129));
  jnot g14937(.din(n15129), .dout(n15130));
  jand g14938(.dina(n15130), .dinb(n15127), .dout(n15131));
  jnot g14939(.din(\a[58] ), .dout(n15132));
  jand g14940(.dina(n15090), .dinb(n15029), .dout(n15133));
  jor  g14941(.dina(n15133), .dinb(n15132), .dout(n15134));
  jnot g14942(.din(n15134), .dout(n15135));
  jxor g14943(.dina(n15135), .dinb(n15131), .dout(n15136));
  jand g14944(.dina(\a[61] ), .dinb(\a[55] ), .dout(n15137));
  jand g14945(.dina(\a[59] ), .dinb(\a[57] ), .dout(n15138));
  jor  g14946(.dina(n15138), .dinb(n15086), .dout(n15139));
  jnot g14947(.din(n15139), .dout(n15140));
  jand g14948(.dina(\a[60] ), .dinb(\a[57] ), .dout(n15141));
  jand g14949(.dina(n15141), .dinb(n15051), .dout(n15142));
  jor  g14950(.dina(n15142), .dinb(n15140), .dout(n15143));
  jxor g14951(.dina(n15143), .dinb(n15137), .dout(n15144));
  jnot g14952(.din(n15144), .dout(n15145));
  jand g14953(.dina(n15084), .dinb(n15082), .dout(n15146));
  jor  g14954(.dina(n15146), .dinb(n15087), .dout(n15147));
  jxor g14955(.dina(n15147), .dinb(n15145), .dout(n15148));
  jxor g14956(.dina(n15148), .dinb(n15136), .dout(n15149));
  jxor g14957(.dina(n15149), .dinb(n15124), .dout(n15150));
  jand g14958(.dina(n15104), .dinb(n15101), .dout(n15151));
  jand g14959(.dina(n15105), .dinb(n15094), .dout(n15152));
  jor  g14960(.dina(n15152), .dinb(n15151), .dout(n15153));
  jxor g14961(.dina(n15153), .dinb(n15150), .dout(n15154));
  jand g14962(.dina(n15106), .dinb(n15078), .dout(n15155));
  jor  g14963(.dina(n15106), .dinb(n15078), .dout(n15156));
  jand g14964(.dina(n15114), .dinb(n15156), .dout(n15157));
  jor  g14965(.dina(n15157), .dinb(n15155), .dout(n15158));
  jxor g14966(.dina(n15158), .dinb(n15154), .dout(\asquared[117] ));
  jand g14967(.dina(n15123), .dinb(n15120), .dout(n15160));
  jand g14968(.dina(n15149), .dinb(n15124), .dout(n15161));
  jor  g14969(.dina(n15161), .dinb(n15160), .dout(n15162));
  jand g14970(.dina(n15147), .dinb(n15145), .dout(n15163));
  jand g14971(.dina(n15148), .dinb(n15136), .dout(n15164));
  jor  g14972(.dina(n15164), .dinb(n15163), .dout(n15165));
  jnot g14973(.din(n15165), .dout(n15166));
  jand g14974(.dina(\a[62] ), .dinb(\a[55] ), .dout(n15167));
  jnot g14975(.din(n15167), .dout(n15168));
  jand g14976(.dina(\a[59] ), .dinb(n15132), .dout(n15169));
  jxor g14977(.dina(n15169), .dinb(n15168), .dout(n15170));
  jxor g14978(.dina(n15170), .dinb(n15166), .dout(n15171));
  jand g14979(.dina(n15135), .dinb(n15131), .dout(n15172));
  jor  g14980(.dina(n15172), .dinb(n15129), .dout(n15173));
  jand g14981(.dina(n15139), .dinb(n15137), .dout(n15174));
  jor  g14982(.dina(n15174), .dinb(n15142), .dout(n15175));
  jxor g14983(.dina(n15175), .dinb(n15173), .dout(n15176));
  jnot g14984(.din(n15141), .dout(n15177));
  jand g14985(.dina(\a[61] ), .dinb(\a[56] ), .dout(n15178));
  jnot g14986(.din(n15178), .dout(n15179));
  jand g14987(.dina(n15179), .dinb(n15177), .dout(n15180));
  jand g14988(.dina(\a[61] ), .dinb(\a[57] ), .dout(n15181));
  jand g14989(.dina(n15181), .dinb(n15086), .dout(n15182));
  jor  g14990(.dina(n15182), .dinb(n15180), .dout(n15183));
  jxor g14991(.dina(n15183), .dinb(n15128), .dout(n15184));
  jnot g14992(.din(n15184), .dout(n15185));
  jxor g14993(.dina(n15185), .dinb(n15176), .dout(n15186));
  jxor g14994(.dina(n15186), .dinb(n15171), .dout(n15187));
  jxor g14995(.dina(n15187), .dinb(n15162), .dout(n15188));
  jand g14996(.dina(n15153), .dinb(n15150), .dout(n15189));
  jnot g14997(.din(n15150), .dout(n15190));
  jnot g14998(.din(n15153), .dout(n15191));
  jand g14999(.dina(n15191), .dinb(n15190), .dout(n15192));
  jnot g15000(.din(n15192), .dout(n15193));
  jand g15001(.dina(n15158), .dinb(n15193), .dout(n15194));
  jor  g15002(.dina(n15194), .dinb(n15189), .dout(n15195));
  jxor g15003(.dina(n15195), .dinb(n15188), .dout(\asquared[118] ));
  jnot g15004(.din(\a[59] ), .dout(n15197));
  jand g15005(.dina(n15168), .dinb(n15132), .dout(n15198));
  jor  g15006(.dina(n15198), .dinb(n15197), .dout(n15199));
  jnot g15007(.din(n15199), .dout(n15200));
  jand g15008(.dina(\a[63] ), .dinb(\a[55] ), .dout(n15201));
  jxor g15009(.dina(n15201), .dinb(n15200), .dout(n15202));
  jnot g15010(.din(n15180), .dout(n15203));
  jand g15011(.dina(n15203), .dinb(n15128), .dout(n15204));
  jor  g15012(.dina(n15204), .dinb(n15182), .dout(n15205));
  jxor g15013(.dina(n15205), .dinb(n15202), .dout(n15206));
  jnot g15014(.din(n15173), .dout(n15207));
  jnot g15015(.din(n15175), .dout(n15208));
  jand g15016(.dina(n15208), .dinb(n15207), .dout(n15209));
  jnot g15017(.din(n15209), .dout(n15210));
  jand g15018(.dina(n15175), .dinb(n15173), .dout(n15211));
  jor  g15019(.dina(n15185), .dinb(n15211), .dout(n15212));
  jand g15020(.dina(n15212), .dinb(n15210), .dout(n15213));
  jnot g15021(.din(n15213), .dout(n15214));
  jand g15022(.dina(\a[62] ), .dinb(\a[56] ), .dout(n15215));
  jand g15023(.dina(\a[60] ), .dinb(\a[58] ), .dout(n15216));
  jor  g15024(.dina(n15216), .dinb(n15181), .dout(n15217));
  jnot g15025(.din(n15217), .dout(n15218));
  jand g15026(.dina(\a[61] ), .dinb(\a[58] ), .dout(n15219));
  jand g15027(.dina(n15219), .dinb(n15141), .dout(n15220));
  jor  g15028(.dina(n15220), .dinb(n15218), .dout(n15221));
  jxor g15029(.dina(n15221), .dinb(n15215), .dout(n15222));
  jxor g15030(.dina(n15222), .dinb(n15214), .dout(n15223));
  jxor g15031(.dina(n15223), .dinb(n15206), .dout(n15224));
  jnot g15032(.din(n15224), .dout(n15225));
  jor  g15033(.dina(n15170), .dinb(n15166), .dout(n15226));
  jand g15034(.dina(n15186), .dinb(n15171), .dout(n15227));
  jnot g15035(.din(n15227), .dout(n15228));
  jand g15036(.dina(n15228), .dinb(n15226), .dout(n15229));
  jxor g15037(.dina(n15229), .dinb(n15225), .dout(n15230));
  jand g15038(.dina(n15187), .dinb(n15162), .dout(n15231));
  jor  g15039(.dina(n15187), .dinb(n15162), .dout(n15232));
  jand g15040(.dina(n15195), .dinb(n15232), .dout(n15233));
  jor  g15041(.dina(n15233), .dinb(n15231), .dout(n15234));
  jxor g15042(.dina(n15234), .dinb(n15230), .dout(\asquared[119] ));
  jand g15043(.dina(n15201), .dinb(n15200), .dout(n15236));
  jand g15044(.dina(n15205), .dinb(n15202), .dout(n15237));
  jor  g15045(.dina(n15237), .dinb(n15236), .dout(n15238));
  jand g15046(.dina(\a[63] ), .dinb(\a[56] ), .dout(n15239));
  jor  g15047(.dina(n15239), .dinb(n15219), .dout(n15240));
  jand g15048(.dina(n15178), .dinb(n14613), .dout(n15241));
  jnot g15049(.din(n15241), .dout(n15242));
  jand g15050(.dina(n15242), .dinb(n15240), .dout(n15243));
  jand g15051(.dina(n15217), .dinb(n15215), .dout(n15244));
  jor  g15052(.dina(n15244), .dinb(n15220), .dout(n15245));
  jxor g15053(.dina(n15245), .dinb(n15243), .dout(n15246));
  jnot g15054(.din(n15246), .dout(n15247));
  jand g15055(.dina(\a[62] ), .dinb(\a[57] ), .dout(n15248));
  jnot g15056(.din(n15248), .dout(n15249));
  jand g15057(.dina(\a[60] ), .dinb(n15197), .dout(n15250));
  jxor g15058(.dina(n15250), .dinb(n15249), .dout(n15251));
  jxor g15059(.dina(n15251), .dinb(n15247), .dout(n15252));
  jxor g15060(.dina(n15252), .dinb(n15238), .dout(n15253));
  jor  g15061(.dina(n15222), .dinb(n15214), .dout(n15254));
  jand g15062(.dina(n15223), .dinb(n15206), .dout(n15255));
  jnot g15063(.din(n15255), .dout(n15256));
  jand g15064(.dina(n15256), .dinb(n15254), .dout(n15257));
  jnot g15065(.din(n15257), .dout(n15258));
  jxor g15066(.dina(n15258), .dinb(n15253), .dout(n15259));
  jor  g15067(.dina(n15229), .dinb(n15225), .dout(n15260));
  jnot g15068(.din(n15260), .dout(n15261));
  jand g15069(.dina(n15229), .dinb(n15225), .dout(n15262));
  jnot g15070(.din(n15262), .dout(n15263));
  jand g15071(.dina(n15234), .dinb(n15263), .dout(n15264));
  jor  g15072(.dina(n15264), .dinb(n15261), .dout(n15265));
  jxor g15073(.dina(n15265), .dinb(n15259), .dout(\asquared[120] ));
  jor  g15074(.dina(n15251), .dinb(n15247), .dout(n15267));
  jand g15075(.dina(n15252), .dinb(n15238), .dout(n15268));
  jnot g15076(.din(n15268), .dout(n15269));
  jand g15077(.dina(n15269), .dinb(n15267), .dout(n15270));
  jand g15078(.dina(n15249), .dinb(n15197), .dout(n15271));
  jor  g15079(.dina(n15271), .dinb(n7411), .dout(n15272));
  jnot g15080(.din(n15272), .dout(n15273));
  jand g15081(.dina(n15245), .dinb(n15243), .dout(n15274));
  jor  g15082(.dina(n15274), .dinb(n15241), .dout(n15275));
  jxor g15083(.dina(n15275), .dinb(n15273), .dout(n15276));
  jnot g15084(.din(n15276), .dout(n15277));
  jand g15085(.dina(\a[63] ), .dinb(\a[57] ), .dout(n15278));
  jand g15086(.dina(\a[62] ), .dinb(\a[58] ), .dout(n15279));
  jand g15087(.dina(\a[61] ), .dinb(\a[59] ), .dout(n15280));
  jor  g15088(.dina(n15280), .dinb(n15279), .dout(n15281));
  jnot g15089(.din(n15281), .dout(n15282));
  jand g15090(.dina(\a[62] ), .dinb(\a[59] ), .dout(n15283));
  jand g15091(.dina(n15283), .dinb(n15219), .dout(n15284));
  jor  g15092(.dina(n15284), .dinb(n15282), .dout(n15285));
  jxor g15093(.dina(n15285), .dinb(n15278), .dout(n15286));
  jxor g15094(.dina(n15286), .dinb(n15277), .dout(n15287));
  jnot g15095(.din(n15287), .dout(n15288));
  jxor g15096(.dina(n15288), .dinb(n15270), .dout(n15289));
  jand g15097(.dina(n15258), .dinb(n15253), .dout(n15290));
  jor  g15098(.dina(n15258), .dinb(n15253), .dout(n15291));
  jand g15099(.dina(n15265), .dinb(n15291), .dout(n15292));
  jor  g15100(.dina(n15292), .dinb(n15290), .dout(n15293));
  jxor g15101(.dina(n15293), .dinb(n15289), .dout(\asquared[121] ));
  jand g15102(.dina(n15281), .dinb(n15278), .dout(n15295));
  jor  g15103(.dina(n15295), .dinb(n15284), .dout(n15296));
  jxor g15104(.dina(n15296), .dinb(n14613), .dout(n15297));
  jnot g15105(.din(n15297), .dout(n15298));
  jnot g15106(.din(n15283), .dout(n15299));
  jand g15107(.dina(\a[61] ), .dinb(n7411), .dout(n15300));
  jxor g15108(.dina(n15300), .dinb(n15299), .dout(n15301));
  jxor g15109(.dina(n15301), .dinb(n15298), .dout(n15302));
  jnot g15110(.din(n15302), .dout(n15303));
  jand g15111(.dina(n15275), .dinb(n15273), .dout(n15304));
  jnot g15112(.din(n15304), .dout(n15305));
  jor  g15113(.dina(n15286), .dinb(n15277), .dout(n15306));
  jand g15114(.dina(n15306), .dinb(n15305), .dout(n15307));
  jxor g15115(.dina(n15307), .dinb(n15303), .dout(n15308));
  jnot g15116(.din(n15270), .dout(n15309));
  jand g15117(.dina(n15287), .dinb(n15309), .dout(n15310));
  jand g15118(.dina(n15288), .dinb(n15270), .dout(n15311));
  jnot g15119(.din(n15311), .dout(n15312));
  jand g15120(.dina(n15293), .dinb(n15312), .dout(n15313));
  jor  g15121(.dina(n15313), .dinb(n15310), .dout(n15314));
  jxor g15122(.dina(n15314), .dinb(n15308), .dout(\asquared[122] ));
  jand g15123(.dina(n15296), .dinb(n14613), .dout(n15316));
  jnot g15124(.din(n15316), .dout(n15317));
  jor  g15125(.dina(n15301), .dinb(n15298), .dout(n15318));
  jand g15126(.dina(n15318), .dinb(n15317), .dout(n15319));
  jand g15127(.dina(\a[62] ), .dinb(\a[60] ), .dout(n15320));
  jand g15128(.dina(\a[63] ), .dinb(\a[59] ), .dout(n15321));
  jor  g15129(.dina(n15321), .dinb(n15320), .dout(n15322));
  jand g15130(.dina(\a[63] ), .dinb(\a[60] ), .dout(n15323));
  jand g15131(.dina(n15323), .dinb(n15283), .dout(n15324));
  jnot g15132(.din(n15324), .dout(n15325));
  jand g15133(.dina(n15325), .dinb(n15322), .dout(n15326));
  jnot g15134(.din(\a[61] ), .dout(n15327));
  jand g15135(.dina(n15299), .dinb(n7411), .dout(n15328));
  jor  g15136(.dina(n15328), .dinb(n15327), .dout(n15329));
  jnot g15137(.din(n15329), .dout(n15330));
  jxor g15138(.dina(n15330), .dinb(n15326), .dout(n15331));
  jnot g15139(.din(n15331), .dout(n15332));
  jxor g15140(.dina(n15332), .dinb(n15319), .dout(n15333));
  jor  g15141(.dina(n15307), .dinb(n15303), .dout(n15334));
  jnot g15142(.din(n15334), .dout(n15335));
  jand g15143(.dina(n15307), .dinb(n15303), .dout(n15336));
  jnot g15144(.din(n15336), .dout(n15337));
  jand g15145(.dina(n15314), .dinb(n15337), .dout(n15338));
  jor  g15146(.dina(n15338), .dinb(n15335), .dout(n15339));
  jxor g15147(.dina(n15339), .dinb(n15333), .dout(\asquared[123] ));
  jand g15148(.dina(n15330), .dinb(n15326), .dout(n15341));
  jor  g15149(.dina(n15341), .dinb(n15324), .dout(n15342));
  jand g15150(.dina(\a[62] ), .dinb(n15327), .dout(n15343));
  jxor g15151(.dina(n15343), .dinb(n15323), .dout(n15344));
  jxor g15152(.dina(n15344), .dinb(n15342), .dout(n15345));
  jor  g15153(.dina(n15332), .dinb(n15319), .dout(n15346));
  jnot g15154(.din(n15346), .dout(n15347));
  jand g15155(.dina(n15332), .dinb(n15319), .dout(n15348));
  jnot g15156(.din(n15348), .dout(n15349));
  jand g15157(.dina(n15339), .dinb(n15349), .dout(n15350));
  jor  g15158(.dina(n15350), .dinb(n15347), .dout(n15351));
  jxor g15159(.dina(n15351), .dinb(n15345), .dout(\asquared[124] ));
  jand g15160(.dina(\a[63] ), .dinb(\a[61] ), .dout(n15353));
  jand g15161(.dina(n15353), .dinb(\a[62] ), .dout(n15354));
  jnot g15162(.din(n15354), .dout(n15355));
  jor  g15163(.dina(n15323), .dinb(\a[61] ), .dout(n15356));
  jand g15164(.dina(n15356), .dinb(\a[62] ), .dout(n15357));
  jor  g15165(.dina(n15357), .dinb(n15353), .dout(n15358));
  jand g15166(.dina(n15358), .dinb(n15355), .dout(n15359));
  jand g15167(.dina(n15344), .dinb(n15342), .dout(n15360));
  jnot g15168(.din(n15342), .dout(n15361));
  jnot g15169(.din(n15344), .dout(n15362));
  jand g15170(.dina(n15362), .dinb(n15361), .dout(n15363));
  jnot g15171(.din(n15363), .dout(n15364));
  jand g15172(.dina(n15351), .dinb(n15364), .dout(n15365));
  jor  g15173(.dina(n15365), .dinb(n15360), .dout(n15366));
  jxor g15174(.dina(n15366), .dinb(n15359), .dout(\asquared[125] ));
  jnot g15175(.din(\a[62] ), .dout(n15368));
  jand g15176(.dina(\a[63] ), .dinb(n15368), .dout(n15369));
  jor  g15177(.dina(n15366), .dinb(n15354), .dout(n15370));
  jand g15178(.dina(n15370), .dinb(n15358), .dout(n15371));
  jxor g15179(.dina(n15371), .dinb(n15369), .dout(\asquared[126] ));
  jor  g15180(.dina(n15371), .dinb(\a[62] ), .dout(n15373));
  jand g15181(.dina(n15373), .dinb(\a[63] ), .dout(\asquared[127] ));
  buf  g15182(.din(\a[0] ), .dout(\asquared[0] ));
endmodule


