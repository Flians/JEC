// Benchmark "top" written by ABC on Wed May 27 23:34:13 2020

module rf_adder ( 
    a0 , a1 , a2 , a3 , a4 , a5 , a6 , a7 , a8 ,
    a9 , a10 , a11 , a12 , a13 , a14 , a15 , a16 ,
    a17 , a18 , a19 , a20 , a21 , a22 , a23 , a24 ,
    a25 , a26 , a27 , a28 , a29 , a30 , a31 , a32 ,
    a33 , a34 , a35 , a36 , a37 , a38 , a39 , a40 ,
    a41 , a42 , a43 , a44 , a45 , a46 , a47 , a48 ,
    a49 , a50 , a51 , a52 , a53 , a54 , a55 , a56 ,
    a57 , a58 , a59 , a60 , a61 , a62 , a63 , a64 ,
    a65 , a66 , a67 , a68 , a69 , a70 , a71 , a72 ,
    a73 , a74 , a75 , a76 , a77 , a78 , a79 , a80 ,
    a81 , a82 , a83 , a84 , a85 , a86 , a87 , a88 ,
    a89 , a90 , a91 , a92 , a93 , a94 , a95 , a96 ,
    a97 , a98 , a99 , a100 , a101 , a102 , a103 ,
    a104 , a105 , a106 , a107 , a108 , a109 , a110 ,
    a111 , a112 , a113 , a114 , a115 , a116 , a117 ,
    a118 , a119 , a120 , a121 , a122 , a123 , a124 ,
    a125 , a126 , a127 , b0 , b1 , b2 , b3 , b4 ,
    b5 , b6 , b7 , b8 , b9 , b10 , b11 , b12 ,
    b13 , b14 , b15 , b16 , b17 , b18 , b19 , b20 ,
    b21 , b22 , b23 , b24 , b25 , b26 , b27 , b28 ,
    b29 , b30 , b31 , b32 , b33 , b34 , b35 , b36 ,
    b37 , b38 , b39 , b40 , b41 , b42 , b43 , b44 ,
    b45 , b46 , b47 , b48 , b49 , b50 , b51 , b52 ,
    b53 , b54 , b55 , b56 , b57 , b58 , b59 , b60 ,
    b61 , b62 , b63 , b64 , b65 , b66 , b67 , b68 ,
    b69 , b70 , b71 , b72 , b73 , b74 , b75 , b76 ,
    b77 , b78 , b79 , b80 , b81 , b82 , b83 , b84 ,
    b85 , b86 , b87 , b88 , b89 , b90 , b91 , b92 ,
    b93 , b94 , b95 , b96 , b97 , b98 , b99 ,
    b100 , b101 , b102 , b103 , b104 , b105 , b106 ,
    b107 , b108 , b109 , b110 , b111 , b112 , b113 ,
    b114 , b115 , b116 , b117 , b118 , b119 , b120 ,
    b121 , b122 , b123 , b124 , b125 , b126 , b127 ,
    f0 , f1 , f2 , f3 , f4 , f5 , f6 , f7 , f8 ,
    f9 , f10 , f11 , f12 , f13 , f14 , f15 , f16 ,
    f17 , f18 , f19 , f20 , f21 , f22 , f23 , f24 ,
    f25 , f26 , f27 , f28 , f29 , f30 , f31 , f32 ,
    f33 , f34 , f35 , f36 , f37 , f38 , f39 , f40 ,
    f41 , f42 , f43 , f44 , f45 , f46 , f47 , f48 ,
    f49 , f50 , f51 , f52 , f53 , f54 , f55 , f56 ,
    f57 , f58 , f59 , f60 , f61 , f62 , f63 , f64 ,
    f65 , f66 , f67 , f68 , f69 , f70 , f71 , f72 ,
    f73 , f74 , f75 , f76 , f77 , f78 , f79 , f80 ,
    f81 , f82 , f83 , f84 , f85 , f86 , f87 , f88 ,
    f89 , f90 , f91 , f92 , f93 , f94 , f95 , f96 ,
    f97 , f98 , f99 , f100 , f101 , f102 , f103 ,
    f104 , f105 , f106 , f107 , f108 , f109 , f110 ,
    f111 , f112 , f113 , f114 , f115 , f116 , f117 ,
    f118 , f119 , f120 , f121 , f122 , f123 , f124 ,
    f125 , f126 , f127 , cOut  );
  input  a0 , a1 , a2 , a3 , a4 , a5 , a6 , a7 ,
    a8 , a9 , a10 , a11 , a12 , a13 , a14 , a15 ,
    a16 , a17 , a18 , a19 , a20 , a21 , a22 , a23 ,
    a24 , a25 , a26 , a27 , a28 , a29 , a30 , a31 ,
    a32 , a33 , a34 , a35 , a36 , a37 , a38 , a39 ,
    a40 , a41 , a42 , a43 , a44 , a45 , a46 , a47 ,
    a48 , a49 , a50 , a51 , a52 , a53 , a54 , a55 ,
    a56 , a57 , a58 , a59 , a60 , a61 , a62 , a63 ,
    a64 , a65 , a66 , a67 , a68 , a69 , a70 , a71 ,
    a72 , a73 , a74 , a75 , a76 , a77 , a78 , a79 ,
    a80 , a81 , a82 , a83 , a84 , a85 , a86 , a87 ,
    a88 , a89 , a90 , a91 , a92 , a93 , a94 , a95 ,
    a96 , a97 , a98 , a99 , a100 , a101 , a102 ,
    a103 , a104 , a105 , a106 , a107 , a108 , a109 ,
    a110 , a111 , a112 , a113 , a114 , a115 , a116 ,
    a117 , a118 , a119 , a120 , a121 , a122 , a123 ,
    a124 , a125 , a126 , a127 , b0 , b1 , b2 , b3 ,
    b4 , b5 , b6 , b7 , b8 , b9 , b10 , b11 ,
    b12 , b13 , b14 , b15 , b16 , b17 , b18 , b19 ,
    b20 , b21 , b22 , b23 , b24 , b25 , b26 , b27 ,
    b28 , b29 , b30 , b31 , b32 , b33 , b34 , b35 ,
    b36 , b37 , b38 , b39 , b40 , b41 , b42 , b43 ,
    b44 , b45 , b46 , b47 , b48 , b49 , b50 , b51 ,
    b52 , b53 , b54 , b55 , b56 , b57 , b58 , b59 ,
    b60 , b61 , b62 , b63 , b64 , b65 , b66 , b67 ,
    b68 , b69 , b70 , b71 , b72 , b73 , b74 , b75 ,
    b76 , b77 , b78 , b79 , b80 , b81 , b82 , b83 ,
    b84 , b85 , b86 , b87 , b88 , b89 , b90 , b91 ,
    b92 , b93 , b94 , b95 , b96 , b97 , b98 , b99 ,
    b100 , b101 , b102 , b103 , b104 , b105 , b106 ,
    b107 , b108 , b109 , b110 , b111 , b112 , b113 ,
    b114 , b115 , b116 , b117 , b118 , b119 , b120 ,
    b121 , b122 , b123 , b124 , b125 , b126 , b127 ;
  output f0 , f1 , f2 , f3 , f4 , f5 , f6 , f7 ,
    f8 , f9 , f10 , f11 , f12 , f13 , f14 , f15 ,
    f16 , f17 , f18 , f19 , f20 , f21 , f22 , f23 ,
    f24 , f25 , f26 , f27 , f28 , f29 , f30 , f31 ,
    f32 , f33 , f34 , f35 , f36 , f37 , f38 , f39 ,
    f40 , f41 , f42 , f43 , f44 , f45 , f46 , f47 ,
    f48 , f49 , f50 , f51 , f52 , f53 , f54 , f55 ,
    f56 , f57 , f58 , f59 , f60 , f61 , f62 , f63 ,
    f64 , f65 , f66 , f67 , f68 , f69 , f70 , f71 ,
    f72 , f73 , f74 , f75 , f76 , f77 , f78 , f79 ,
    f80 , f81 , f82 , f83 , f84 , f85 , f86 , f87 ,
    f88 , f89 , f90 , f91 , f92 , f93 , f94 , f95 ,
    f96 , f97 , f98 , f99 , f100 , f101 , f102 ,
    f103 , f104 , f105 , f106 , f107 , f108 , f109 ,
    f110 , f111 , f112 , f113 , f114 , f115 , f116 ,
    f117 , f118 , f119 , f120 , f121 , f122 , f123 ,
    f124 , f125 , f126 , f127 , cOut;
  wire n386, n387, n389, n390, n391, n392, n393, n395, n396, n397, n398,
    n399, n401, n402, n403, n404, n405, n407, n408, n409, n410, n411, n413,
    n414, n415, n416, n417, n419, n420, n421, n422, n423, n425, n426, n427,
    n428, n429, n431, n432, n433, n434, n435, n437, n438, n439, n440, n441,
    n443, n444, n445, n446, n447, n449, n450, n451, n452, n453, n455, n456,
    n457, n458, n459, n461, n462, n463, n464, n465, n467, n468, n469, n470,
    n471, n473, n474, n475, n476, n477, n479, n480, n481, n482, n483, n485,
    n486, n487, n488, n489, n491, n492, n493, n494, n495, n497, n498, n499,
    n500, n501, n503, n504, n505, n506, n507, n509, n510, n511, n512, n513,
    n515, n516, n517, n518, n519, n521, n522, n523, n524, n525, n527, n528,
    n529, n530, n531, n533, n534, n535, n536, n537, n539, n540, n541, n542,
    n543, n545, n546, n547, n548, n549, n551, n552, n553, n554, n555, n557,
    n558, n559, n560, n561, n563, n564, n565, n566, n567, n569, n570, n571,
    n572, n573, n575, n576, n577, n578, n579, n581, n582, n583, n584, n585,
    n587, n588, n589, n590, n591, n593, n594, n595, n596, n597, n599, n600,
    n601, n602, n603, n605, n606, n607, n608, n609, n611, n612, n613, n614,
    n615, n617, n618, n619, n620, n621, n623, n624, n625, n626, n627, n629,
    n630, n631, n632, n633, n635, n636, n637, n638, n639, n641, n642, n643,
    n644, n645, n647, n648, n649, n650, n651, n653, n654, n655, n656, n657,
    n659, n660, n661, n662, n663, n665, n666, n667, n668, n669, n671, n672,
    n673, n674, n675, n677, n678, n679, n680, n681, n683, n684, n685, n686,
    n687, n689, n690, n691, n692, n693, n695, n696, n697, n698, n699, n701,
    n702, n703, n704, n705, n707, n708, n709, n710, n711, n713, n714, n715,
    n716, n717, n719, n720, n721, n722, n723, n725, n726, n727, n728, n729,
    n731, n732, n733, n734, n735, n737, n738, n739, n740, n741, n743, n744,
    n745, n746, n747, n749, n750, n751, n752, n753, n755, n756, n757, n758,
    n759, n761, n762, n763, n764, n765, n767, n768, n769, n770, n771, n773,
    n774, n775, n776, n777, n779, n780, n781, n782, n783, n785, n786, n787,
    n788, n789, n791, n792, n793, n794, n795, n797, n798, n799, n800, n801,
    n803, n804, n805, n806, n807, n809, n810, n811, n812, n813, n815, n816,
    n817, n818, n819, n821, n822, n823, n824, n825, n827, n828, n829, n830,
    n831, n833, n834, n835, n836, n837, n839, n840, n841, n842, n843, n845,
    n846, n847, n848, n849, n851, n852, n853, n854, n855, n857, n858, n859,
    n860, n861, n863, n864, n865, n866, n867, n869, n870, n871, n872, n873,
    n875, n876, n877, n878, n879, n881, n882, n883, n884, n885, n887, n888,
    n889, n890, n891, n893, n894, n895, n896, n897, n899, n900, n901, n902,
    n903, n905, n906, n907, n908, n909, n911, n912, n913, n914, n915, n917,
    n918, n919, n920, n921, n923, n924, n925, n926, n927, n929, n930, n931,
    n932, n933, n935, n936, n937, n938, n939, n941, n942, n943, n944, n945,
    n947, n948, n949, n950, n951, n953, n954, n955, n956, n957, n959, n960,
    n961, n962, n963, n965, n966, n967, n968, n969, n971, n972, n973, n974,
    n975, n977, n978, n979, n980, n981, n983, n984, n985, n986, n987, n989,
    n990, n991, n992, n993, n995, n996, n997, n998, n999, n1001, n1002,
    n1003, n1004, n1005, n1007, n1008, n1009, n1010, n1011, n1013, n1014,
    n1015, n1016, n1017, n1019, n1020, n1021, n1022, n1023, n1025, n1026,
    n1027, n1028, n1029, n1031, n1032, n1033, n1034, n1035, n1037, n1038,
    n1039, n1040, n1041, n1043, n1044, n1045, n1046, n1047, n1049, n1050,
    n1051, n1052, n1053, n1055, n1056, n1057, n1058, n1059, n1061, n1062,
    n1063, n1064, n1065, n1067, n1068, n1069, n1070, n1071, n1073, n1074,
    n1075, n1076, n1077, n1079, n1080, n1081, n1082, n1083, n1085, n1086,
    n1087, n1088, n1089, n1091, n1092, n1093, n1094, n1095, n1097, n1098,
    n1099, n1100, n1101, n1103, n1104, n1105, n1106, n1107, n1109, n1110,
    n1111, n1112, n1113, n1115, n1116, n1117, n1118, n1119, n1121, n1122,
    n1123, n1124, n1125, n1127, n1128, n1129, n1130, n1131, n1133, n1134,
    n1135, n1136, n1137, n1139, n1140, n1141, n1142, n1143, n1145, n1146,
    n1147;
  jxor g000(.dina(b0 ), .dinb(a0 ), .dout(f0 ));
  jand g001(.dina(b0 ), .dinb(a0 ), .dout(n386));
  jxor g002(.dina(b1 ), .dinb(a1 ), .dout(n387));
  jxor g003(.dina(n387), .dinb(n386), .dout(f1 ));
  jxor g004(.dina(b2 ), .dinb(a2 ), .dout(n389));
  jor  g005(.dina(b1 ), .dinb(a1 ), .dout(n390));
  jand g006(.dina(b1 ), .dinb(a1 ), .dout(n391));
  jor  g007(.dina(n391), .dinb(n386), .dout(n392));
  jand g008(.dina(n392), .dinb(n390), .dout(n393));
  jxor g009(.dina(n393), .dinb(n389), .dout(f2 ));
  jxor g010(.dina(b3 ), .dinb(a3 ), .dout(n395));
  jor  g011(.dina(b2 ), .dinb(a2 ), .dout(n396));
  jand g012(.dina(b2 ), .dinb(a2 ), .dout(n397));
  jor  g013(.dina(n393), .dinb(n397), .dout(n398));
  jand g014(.dina(n398), .dinb(n396), .dout(n399));
  jxor g015(.dina(n399), .dinb(n395), .dout(f3 ));
  jxor g016(.dina(b4 ), .dinb(a4 ), .dout(n401));
  jor  g017(.dina(b3 ), .dinb(a3 ), .dout(n402));
  jand g018(.dina(b3 ), .dinb(a3 ), .dout(n403));
  jor  g019(.dina(n399), .dinb(n403), .dout(n404));
  jand g020(.dina(n404), .dinb(n402), .dout(n405));
  jxor g021(.dina(n405), .dinb(n401), .dout(f4 ));
  jxor g022(.dina(b5 ), .dinb(a5 ), .dout(n407));
  jor  g023(.dina(b4 ), .dinb(a4 ), .dout(n408));
  jand g024(.dina(b4 ), .dinb(a4 ), .dout(n409));
  jor  g025(.dina(n405), .dinb(n409), .dout(n410));
  jand g026(.dina(n410), .dinb(n408), .dout(n411));
  jxor g027(.dina(n411), .dinb(n407), .dout(f5 ));
  jxor g028(.dina(b6 ), .dinb(a6 ), .dout(n413));
  jor  g029(.dina(b5 ), .dinb(a5 ), .dout(n414));
  jand g030(.dina(b5 ), .dinb(a5 ), .dout(n415));
  jor  g031(.dina(n411), .dinb(n415), .dout(n416));
  jand g032(.dina(n416), .dinb(n414), .dout(n417));
  jxor g033(.dina(n417), .dinb(n413), .dout(f6 ));
  jxor g034(.dina(b7 ), .dinb(a7 ), .dout(n419));
  jor  g035(.dina(b6 ), .dinb(a6 ), .dout(n420));
  jand g036(.dina(b6 ), .dinb(a6 ), .dout(n421));
  jor  g037(.dina(n417), .dinb(n421), .dout(n422));
  jand g038(.dina(n422), .dinb(n420), .dout(n423));
  jxor g039(.dina(n423), .dinb(n419), .dout(f7 ));
  jxor g040(.dina(b8 ), .dinb(a8 ), .dout(n425));
  jor  g041(.dina(b7 ), .dinb(a7 ), .dout(n426));
  jand g042(.dina(b7 ), .dinb(a7 ), .dout(n427));
  jor  g043(.dina(n423), .dinb(n427), .dout(n428));
  jand g044(.dina(n428), .dinb(n426), .dout(n429));
  jxor g045(.dina(n429), .dinb(n425), .dout(f8 ));
  jxor g046(.dina(b9 ), .dinb(a9 ), .dout(n431));
  jor  g047(.dina(b8 ), .dinb(a8 ), .dout(n432));
  jand g048(.dina(b8 ), .dinb(a8 ), .dout(n433));
  jor  g049(.dina(n429), .dinb(n433), .dout(n434));
  jand g050(.dina(n434), .dinb(n432), .dout(n435));
  jxor g051(.dina(n435), .dinb(n431), .dout(f9 ));
  jxor g052(.dina(b10 ), .dinb(a10 ), .dout(n437));
  jor  g053(.dina(b9 ), .dinb(a9 ), .dout(n438));
  jand g054(.dina(b9 ), .dinb(a9 ), .dout(n439));
  jor  g055(.dina(n435), .dinb(n439), .dout(n440));
  jand g056(.dina(n440), .dinb(n438), .dout(n441));
  jxor g057(.dina(n441), .dinb(n437), .dout(f10 ));
  jxor g058(.dina(b11 ), .dinb(a11 ), .dout(n443));
  jor  g059(.dina(b10 ), .dinb(a10 ), .dout(n444));
  jand g060(.dina(b10 ), .dinb(a10 ), .dout(n445));
  jor  g061(.dina(n441), .dinb(n445), .dout(n446));
  jand g062(.dina(n446), .dinb(n444), .dout(n447));
  jxor g063(.dina(n447), .dinb(n443), .dout(f11 ));
  jxor g064(.dina(b12 ), .dinb(a12 ), .dout(n449));
  jor  g065(.dina(b11 ), .dinb(a11 ), .dout(n450));
  jand g066(.dina(b11 ), .dinb(a11 ), .dout(n451));
  jor  g067(.dina(n447), .dinb(n451), .dout(n452));
  jand g068(.dina(n452), .dinb(n450), .dout(n453));
  jxor g069(.dina(n453), .dinb(n449), .dout(f12 ));
  jxor g070(.dina(b13 ), .dinb(a13 ), .dout(n455));
  jor  g071(.dina(b12 ), .dinb(a12 ), .dout(n456));
  jand g072(.dina(b12 ), .dinb(a12 ), .dout(n457));
  jor  g073(.dina(n453), .dinb(n457), .dout(n458));
  jand g074(.dina(n458), .dinb(n456), .dout(n459));
  jxor g075(.dina(n459), .dinb(n455), .dout(f13 ));
  jxor g076(.dina(b14 ), .dinb(a14 ), .dout(n461));
  jor  g077(.dina(b13 ), .dinb(a13 ), .dout(n462));
  jand g078(.dina(b13 ), .dinb(a13 ), .dout(n463));
  jor  g079(.dina(n459), .dinb(n463), .dout(n464));
  jand g080(.dina(n464), .dinb(n462), .dout(n465));
  jxor g081(.dina(n465), .dinb(n461), .dout(f14 ));
  jxor g082(.dina(b15 ), .dinb(a15 ), .dout(n467));
  jor  g083(.dina(b14 ), .dinb(a14 ), .dout(n468));
  jand g084(.dina(b14 ), .dinb(a14 ), .dout(n469));
  jor  g085(.dina(n465), .dinb(n469), .dout(n470));
  jand g086(.dina(n470), .dinb(n468), .dout(n471));
  jxor g087(.dina(n471), .dinb(n467), .dout(f15 ));
  jxor g088(.dina(b16 ), .dinb(a16 ), .dout(n473));
  jor  g089(.dina(b15 ), .dinb(a15 ), .dout(n474));
  jand g090(.dina(b15 ), .dinb(a15 ), .dout(n475));
  jor  g091(.dina(n471), .dinb(n475), .dout(n476));
  jand g092(.dina(n476), .dinb(n474), .dout(n477));
  jxor g093(.dina(n477), .dinb(n473), .dout(f16 ));
  jxor g094(.dina(b17 ), .dinb(a17 ), .dout(n479));
  jor  g095(.dina(b16 ), .dinb(a16 ), .dout(n480));
  jand g096(.dina(b16 ), .dinb(a16 ), .dout(n481));
  jor  g097(.dina(n477), .dinb(n481), .dout(n482));
  jand g098(.dina(n482), .dinb(n480), .dout(n483));
  jxor g099(.dina(n483), .dinb(n479), .dout(f17 ));
  jxor g100(.dina(b18 ), .dinb(a18 ), .dout(n485));
  jor  g101(.dina(b17 ), .dinb(a17 ), .dout(n486));
  jand g102(.dina(b17 ), .dinb(a17 ), .dout(n487));
  jor  g103(.dina(n483), .dinb(n487), .dout(n488));
  jand g104(.dina(n488), .dinb(n486), .dout(n489));
  jxor g105(.dina(n489), .dinb(n485), .dout(f18 ));
  jxor g106(.dina(b19 ), .dinb(a19 ), .dout(n491));
  jor  g107(.dina(b18 ), .dinb(a18 ), .dout(n492));
  jand g108(.dina(b18 ), .dinb(a18 ), .dout(n493));
  jor  g109(.dina(n489), .dinb(n493), .dout(n494));
  jand g110(.dina(n494), .dinb(n492), .dout(n495));
  jxor g111(.dina(n495), .dinb(n491), .dout(f19 ));
  jxor g112(.dina(b20 ), .dinb(a20 ), .dout(n497));
  jor  g113(.dina(b19 ), .dinb(a19 ), .dout(n498));
  jand g114(.dina(b19 ), .dinb(a19 ), .dout(n499));
  jor  g115(.dina(n495), .dinb(n499), .dout(n500));
  jand g116(.dina(n500), .dinb(n498), .dout(n501));
  jxor g117(.dina(n501), .dinb(n497), .dout(f20 ));
  jxor g118(.dina(b21 ), .dinb(a21 ), .dout(n503));
  jor  g119(.dina(b20 ), .dinb(a20 ), .dout(n504));
  jand g120(.dina(b20 ), .dinb(a20 ), .dout(n505));
  jor  g121(.dina(n501), .dinb(n505), .dout(n506));
  jand g122(.dina(n506), .dinb(n504), .dout(n507));
  jxor g123(.dina(n507), .dinb(n503), .dout(f21 ));
  jxor g124(.dina(b22 ), .dinb(a22 ), .dout(n509));
  jor  g125(.dina(b21 ), .dinb(a21 ), .dout(n510));
  jand g126(.dina(b21 ), .dinb(a21 ), .dout(n511));
  jor  g127(.dina(n507), .dinb(n511), .dout(n512));
  jand g128(.dina(n512), .dinb(n510), .dout(n513));
  jxor g129(.dina(n513), .dinb(n509), .dout(f22 ));
  jxor g130(.dina(b23 ), .dinb(a23 ), .dout(n515));
  jor  g131(.dina(b22 ), .dinb(a22 ), .dout(n516));
  jand g132(.dina(b22 ), .dinb(a22 ), .dout(n517));
  jor  g133(.dina(n513), .dinb(n517), .dout(n518));
  jand g134(.dina(n518), .dinb(n516), .dout(n519));
  jxor g135(.dina(n519), .dinb(n515), .dout(f23 ));
  jxor g136(.dina(b24 ), .dinb(a24 ), .dout(n521));
  jor  g137(.dina(b23 ), .dinb(a23 ), .dout(n522));
  jand g138(.dina(b23 ), .dinb(a23 ), .dout(n523));
  jor  g139(.dina(n519), .dinb(n523), .dout(n524));
  jand g140(.dina(n524), .dinb(n522), .dout(n525));
  jxor g141(.dina(n525), .dinb(n521), .dout(f24 ));
  jxor g142(.dina(b25 ), .dinb(a25 ), .dout(n527));
  jor  g143(.dina(b24 ), .dinb(a24 ), .dout(n528));
  jand g144(.dina(b24 ), .dinb(a24 ), .dout(n529));
  jor  g145(.dina(n525), .dinb(n529), .dout(n530));
  jand g146(.dina(n530), .dinb(n528), .dout(n531));
  jxor g147(.dina(n531), .dinb(n527), .dout(f25 ));
  jxor g148(.dina(b26 ), .dinb(a26 ), .dout(n533));
  jor  g149(.dina(b25 ), .dinb(a25 ), .dout(n534));
  jand g150(.dina(b25 ), .dinb(a25 ), .dout(n535));
  jor  g151(.dina(n531), .dinb(n535), .dout(n536));
  jand g152(.dina(n536), .dinb(n534), .dout(n537));
  jxor g153(.dina(n537), .dinb(n533), .dout(f26 ));
  jxor g154(.dina(b27 ), .dinb(a27 ), .dout(n539));
  jor  g155(.dina(b26 ), .dinb(a26 ), .dout(n540));
  jand g156(.dina(b26 ), .dinb(a26 ), .dout(n541));
  jor  g157(.dina(n537), .dinb(n541), .dout(n542));
  jand g158(.dina(n542), .dinb(n540), .dout(n543));
  jxor g159(.dina(n543), .dinb(n539), .dout(f27 ));
  jxor g160(.dina(b28 ), .dinb(a28 ), .dout(n545));
  jor  g161(.dina(b27 ), .dinb(a27 ), .dout(n546));
  jand g162(.dina(b27 ), .dinb(a27 ), .dout(n547));
  jor  g163(.dina(n543), .dinb(n547), .dout(n548));
  jand g164(.dina(n548), .dinb(n546), .dout(n549));
  jxor g165(.dina(n549), .dinb(n545), .dout(f28 ));
  jxor g166(.dina(b29 ), .dinb(a29 ), .dout(n551));
  jor  g167(.dina(b28 ), .dinb(a28 ), .dout(n552));
  jand g168(.dina(b28 ), .dinb(a28 ), .dout(n553));
  jor  g169(.dina(n549), .dinb(n553), .dout(n554));
  jand g170(.dina(n554), .dinb(n552), .dout(n555));
  jxor g171(.dina(n555), .dinb(n551), .dout(f29 ));
  jxor g172(.dina(b30 ), .dinb(a30 ), .dout(n557));
  jor  g173(.dina(b29 ), .dinb(a29 ), .dout(n558));
  jand g174(.dina(b29 ), .dinb(a29 ), .dout(n559));
  jor  g175(.dina(n555), .dinb(n559), .dout(n560));
  jand g176(.dina(n560), .dinb(n558), .dout(n561));
  jxor g177(.dina(n561), .dinb(n557), .dout(f30 ));
  jxor g178(.dina(b31 ), .dinb(a31 ), .dout(n563));
  jor  g179(.dina(b30 ), .dinb(a30 ), .dout(n564));
  jand g180(.dina(b30 ), .dinb(a30 ), .dout(n565));
  jor  g181(.dina(n561), .dinb(n565), .dout(n566));
  jand g182(.dina(n566), .dinb(n564), .dout(n567));
  jxor g183(.dina(n567), .dinb(n563), .dout(f31 ));
  jxor g184(.dina(b32 ), .dinb(a32 ), .dout(n569));
  jor  g185(.dina(b31 ), .dinb(a31 ), .dout(n570));
  jand g186(.dina(b31 ), .dinb(a31 ), .dout(n571));
  jor  g187(.dina(n567), .dinb(n571), .dout(n572));
  jand g188(.dina(n572), .dinb(n570), .dout(n573));
  jxor g189(.dina(n573), .dinb(n569), .dout(f32 ));
  jxor g190(.dina(b33 ), .dinb(a33 ), .dout(n575));
  jor  g191(.dina(b32 ), .dinb(a32 ), .dout(n576));
  jand g192(.dina(b32 ), .dinb(a32 ), .dout(n577));
  jor  g193(.dina(n573), .dinb(n577), .dout(n578));
  jand g194(.dina(n578), .dinb(n576), .dout(n579));
  jxor g195(.dina(n579), .dinb(n575), .dout(f33 ));
  jxor g196(.dina(b34 ), .dinb(a34 ), .dout(n581));
  jor  g197(.dina(b33 ), .dinb(a33 ), .dout(n582));
  jand g198(.dina(b33 ), .dinb(a33 ), .dout(n583));
  jor  g199(.dina(n579), .dinb(n583), .dout(n584));
  jand g200(.dina(n584), .dinb(n582), .dout(n585));
  jxor g201(.dina(n585), .dinb(n581), .dout(f34 ));
  jxor g202(.dina(b35 ), .dinb(a35 ), .dout(n587));
  jor  g203(.dina(b34 ), .dinb(a34 ), .dout(n588));
  jand g204(.dina(b34 ), .dinb(a34 ), .dout(n589));
  jor  g205(.dina(n585), .dinb(n589), .dout(n590));
  jand g206(.dina(n590), .dinb(n588), .dout(n591));
  jxor g207(.dina(n591), .dinb(n587), .dout(f35 ));
  jxor g208(.dina(b36 ), .dinb(a36 ), .dout(n593));
  jor  g209(.dina(b35 ), .dinb(a35 ), .dout(n594));
  jand g210(.dina(b35 ), .dinb(a35 ), .dout(n595));
  jor  g211(.dina(n591), .dinb(n595), .dout(n596));
  jand g212(.dina(n596), .dinb(n594), .dout(n597));
  jxor g213(.dina(n597), .dinb(n593), .dout(f36 ));
  jxor g214(.dina(b37 ), .dinb(a37 ), .dout(n599));
  jor  g215(.dina(b36 ), .dinb(a36 ), .dout(n600));
  jand g216(.dina(b36 ), .dinb(a36 ), .dout(n601));
  jor  g217(.dina(n597), .dinb(n601), .dout(n602));
  jand g218(.dina(n602), .dinb(n600), .dout(n603));
  jxor g219(.dina(n603), .dinb(n599), .dout(f37 ));
  jxor g220(.dina(b38 ), .dinb(a38 ), .dout(n605));
  jor  g221(.dina(b37 ), .dinb(a37 ), .dout(n606));
  jand g222(.dina(b37 ), .dinb(a37 ), .dout(n607));
  jor  g223(.dina(n603), .dinb(n607), .dout(n608));
  jand g224(.dina(n608), .dinb(n606), .dout(n609));
  jxor g225(.dina(n609), .dinb(n605), .dout(f38 ));
  jxor g226(.dina(b39 ), .dinb(a39 ), .dout(n611));
  jor  g227(.dina(b38 ), .dinb(a38 ), .dout(n612));
  jand g228(.dina(b38 ), .dinb(a38 ), .dout(n613));
  jor  g229(.dina(n609), .dinb(n613), .dout(n614));
  jand g230(.dina(n614), .dinb(n612), .dout(n615));
  jxor g231(.dina(n615), .dinb(n611), .dout(f39 ));
  jxor g232(.dina(b40 ), .dinb(a40 ), .dout(n617));
  jor  g233(.dina(b39 ), .dinb(a39 ), .dout(n618));
  jand g234(.dina(b39 ), .dinb(a39 ), .dout(n619));
  jor  g235(.dina(n615), .dinb(n619), .dout(n620));
  jand g236(.dina(n620), .dinb(n618), .dout(n621));
  jxor g237(.dina(n621), .dinb(n617), .dout(f40 ));
  jxor g238(.dina(b41 ), .dinb(a41 ), .dout(n623));
  jor  g239(.dina(b40 ), .dinb(a40 ), .dout(n624));
  jand g240(.dina(b40 ), .dinb(a40 ), .dout(n625));
  jor  g241(.dina(n621), .dinb(n625), .dout(n626));
  jand g242(.dina(n626), .dinb(n624), .dout(n627));
  jxor g243(.dina(n627), .dinb(n623), .dout(f41 ));
  jxor g244(.dina(b42 ), .dinb(a42 ), .dout(n629));
  jor  g245(.dina(b41 ), .dinb(a41 ), .dout(n630));
  jand g246(.dina(b41 ), .dinb(a41 ), .dout(n631));
  jor  g247(.dina(n627), .dinb(n631), .dout(n632));
  jand g248(.dina(n632), .dinb(n630), .dout(n633));
  jxor g249(.dina(n633), .dinb(n629), .dout(f42 ));
  jxor g250(.dina(b43 ), .dinb(a43 ), .dout(n635));
  jor  g251(.dina(b42 ), .dinb(a42 ), .dout(n636));
  jand g252(.dina(b42 ), .dinb(a42 ), .dout(n637));
  jor  g253(.dina(n633), .dinb(n637), .dout(n638));
  jand g254(.dina(n638), .dinb(n636), .dout(n639));
  jxor g255(.dina(n639), .dinb(n635), .dout(f43 ));
  jxor g256(.dina(b44 ), .dinb(a44 ), .dout(n641));
  jor  g257(.dina(b43 ), .dinb(a43 ), .dout(n642));
  jand g258(.dina(b43 ), .dinb(a43 ), .dout(n643));
  jor  g259(.dina(n639), .dinb(n643), .dout(n644));
  jand g260(.dina(n644), .dinb(n642), .dout(n645));
  jxor g261(.dina(n645), .dinb(n641), .dout(f44 ));
  jxor g262(.dina(b45 ), .dinb(a45 ), .dout(n647));
  jor  g263(.dina(b44 ), .dinb(a44 ), .dout(n648));
  jand g264(.dina(b44 ), .dinb(a44 ), .dout(n649));
  jor  g265(.dina(n645), .dinb(n649), .dout(n650));
  jand g266(.dina(n650), .dinb(n648), .dout(n651));
  jxor g267(.dina(n651), .dinb(n647), .dout(f45 ));
  jxor g268(.dina(b46 ), .dinb(a46 ), .dout(n653));
  jor  g269(.dina(b45 ), .dinb(a45 ), .dout(n654));
  jand g270(.dina(b45 ), .dinb(a45 ), .dout(n655));
  jor  g271(.dina(n651), .dinb(n655), .dout(n656));
  jand g272(.dina(n656), .dinb(n654), .dout(n657));
  jxor g273(.dina(n657), .dinb(n653), .dout(f46 ));
  jxor g274(.dina(b47 ), .dinb(a47 ), .dout(n659));
  jor  g275(.dina(b46 ), .dinb(a46 ), .dout(n660));
  jand g276(.dina(b46 ), .dinb(a46 ), .dout(n661));
  jor  g277(.dina(n657), .dinb(n661), .dout(n662));
  jand g278(.dina(n662), .dinb(n660), .dout(n663));
  jxor g279(.dina(n663), .dinb(n659), .dout(f47 ));
  jxor g280(.dina(b48 ), .dinb(a48 ), .dout(n665));
  jor  g281(.dina(b47 ), .dinb(a47 ), .dout(n666));
  jand g282(.dina(b47 ), .dinb(a47 ), .dout(n667));
  jor  g283(.dina(n663), .dinb(n667), .dout(n668));
  jand g284(.dina(n668), .dinb(n666), .dout(n669));
  jxor g285(.dina(n669), .dinb(n665), .dout(f48 ));
  jxor g286(.dina(b49 ), .dinb(a49 ), .dout(n671));
  jor  g287(.dina(b48 ), .dinb(a48 ), .dout(n672));
  jand g288(.dina(b48 ), .dinb(a48 ), .dout(n673));
  jor  g289(.dina(n669), .dinb(n673), .dout(n674));
  jand g290(.dina(n674), .dinb(n672), .dout(n675));
  jxor g291(.dina(n675), .dinb(n671), .dout(f49 ));
  jxor g292(.dina(b50 ), .dinb(a50 ), .dout(n677));
  jor  g293(.dina(b49 ), .dinb(a49 ), .dout(n678));
  jand g294(.dina(b49 ), .dinb(a49 ), .dout(n679));
  jor  g295(.dina(n675), .dinb(n679), .dout(n680));
  jand g296(.dina(n680), .dinb(n678), .dout(n681));
  jxor g297(.dina(n681), .dinb(n677), .dout(f50 ));
  jxor g298(.dina(b51 ), .dinb(a51 ), .dout(n683));
  jor  g299(.dina(b50 ), .dinb(a50 ), .dout(n684));
  jand g300(.dina(b50 ), .dinb(a50 ), .dout(n685));
  jor  g301(.dina(n681), .dinb(n685), .dout(n686));
  jand g302(.dina(n686), .dinb(n684), .dout(n687));
  jxor g303(.dina(n687), .dinb(n683), .dout(f51 ));
  jxor g304(.dina(b52 ), .dinb(a52 ), .dout(n689));
  jor  g305(.dina(b51 ), .dinb(a51 ), .dout(n690));
  jand g306(.dina(b51 ), .dinb(a51 ), .dout(n691));
  jor  g307(.dina(n687), .dinb(n691), .dout(n692));
  jand g308(.dina(n692), .dinb(n690), .dout(n693));
  jxor g309(.dina(n693), .dinb(n689), .dout(f52 ));
  jxor g310(.dina(b53 ), .dinb(a53 ), .dout(n695));
  jor  g311(.dina(b52 ), .dinb(a52 ), .dout(n696));
  jand g312(.dina(b52 ), .dinb(a52 ), .dout(n697));
  jor  g313(.dina(n693), .dinb(n697), .dout(n698));
  jand g314(.dina(n698), .dinb(n696), .dout(n699));
  jxor g315(.dina(n699), .dinb(n695), .dout(f53 ));
  jxor g316(.dina(b54 ), .dinb(a54 ), .dout(n701));
  jor  g317(.dina(b53 ), .dinb(a53 ), .dout(n702));
  jand g318(.dina(b53 ), .dinb(a53 ), .dout(n703));
  jor  g319(.dina(n699), .dinb(n703), .dout(n704));
  jand g320(.dina(n704), .dinb(n702), .dout(n705));
  jxor g321(.dina(n705), .dinb(n701), .dout(f54 ));
  jxor g322(.dina(b55 ), .dinb(a55 ), .dout(n707));
  jor  g323(.dina(b54 ), .dinb(a54 ), .dout(n708));
  jand g324(.dina(b54 ), .dinb(a54 ), .dout(n709));
  jor  g325(.dina(n705), .dinb(n709), .dout(n710));
  jand g326(.dina(n710), .dinb(n708), .dout(n711));
  jxor g327(.dina(n711), .dinb(n707), .dout(f55 ));
  jxor g328(.dina(b56 ), .dinb(a56 ), .dout(n713));
  jor  g329(.dina(b55 ), .dinb(a55 ), .dout(n714));
  jand g330(.dina(b55 ), .dinb(a55 ), .dout(n715));
  jor  g331(.dina(n711), .dinb(n715), .dout(n716));
  jand g332(.dina(n716), .dinb(n714), .dout(n717));
  jxor g333(.dina(n717), .dinb(n713), .dout(f56 ));
  jxor g334(.dina(b57 ), .dinb(a57 ), .dout(n719));
  jor  g335(.dina(b56 ), .dinb(a56 ), .dout(n720));
  jand g336(.dina(b56 ), .dinb(a56 ), .dout(n721));
  jor  g337(.dina(n717), .dinb(n721), .dout(n722));
  jand g338(.dina(n722), .dinb(n720), .dout(n723));
  jxor g339(.dina(n723), .dinb(n719), .dout(f57 ));
  jxor g340(.dina(b58 ), .dinb(a58 ), .dout(n725));
  jor  g341(.dina(b57 ), .dinb(a57 ), .dout(n726));
  jand g342(.dina(b57 ), .dinb(a57 ), .dout(n727));
  jor  g343(.dina(n723), .dinb(n727), .dout(n728));
  jand g344(.dina(n728), .dinb(n726), .dout(n729));
  jxor g345(.dina(n729), .dinb(n725), .dout(f58 ));
  jxor g346(.dina(b59 ), .dinb(a59 ), .dout(n731));
  jor  g347(.dina(b58 ), .dinb(a58 ), .dout(n732));
  jand g348(.dina(b58 ), .dinb(a58 ), .dout(n733));
  jor  g349(.dina(n729), .dinb(n733), .dout(n734));
  jand g350(.dina(n734), .dinb(n732), .dout(n735));
  jxor g351(.dina(n735), .dinb(n731), .dout(f59 ));
  jxor g352(.dina(b60 ), .dinb(a60 ), .dout(n737));
  jor  g353(.dina(b59 ), .dinb(a59 ), .dout(n738));
  jand g354(.dina(b59 ), .dinb(a59 ), .dout(n739));
  jor  g355(.dina(n735), .dinb(n739), .dout(n740));
  jand g356(.dina(n740), .dinb(n738), .dout(n741));
  jxor g357(.dina(n741), .dinb(n737), .dout(f60 ));
  jxor g358(.dina(b61 ), .dinb(a61 ), .dout(n743));
  jor  g359(.dina(b60 ), .dinb(a60 ), .dout(n744));
  jand g360(.dina(b60 ), .dinb(a60 ), .dout(n745));
  jor  g361(.dina(n741), .dinb(n745), .dout(n746));
  jand g362(.dina(n746), .dinb(n744), .dout(n747));
  jxor g363(.dina(n747), .dinb(n743), .dout(f61 ));
  jxor g364(.dina(b62 ), .dinb(a62 ), .dout(n749));
  jor  g365(.dina(b61 ), .dinb(a61 ), .dout(n750));
  jand g366(.dina(b61 ), .dinb(a61 ), .dout(n751));
  jor  g367(.dina(n747), .dinb(n751), .dout(n752));
  jand g368(.dina(n752), .dinb(n750), .dout(n753));
  jxor g369(.dina(n753), .dinb(n749), .dout(f62 ));
  jxor g370(.dina(b63 ), .dinb(a63 ), .dout(n755));
  jor  g371(.dina(b62 ), .dinb(a62 ), .dout(n756));
  jand g372(.dina(b62 ), .dinb(a62 ), .dout(n757));
  jor  g373(.dina(n753), .dinb(n757), .dout(n758));
  jand g374(.dina(n758), .dinb(n756), .dout(n759));
  jxor g375(.dina(n759), .dinb(n755), .dout(f63 ));
  jxor g376(.dina(b64 ), .dinb(a64 ), .dout(n761));
  jor  g377(.dina(b63 ), .dinb(a63 ), .dout(n762));
  jand g378(.dina(b63 ), .dinb(a63 ), .dout(n763));
  jor  g379(.dina(n759), .dinb(n763), .dout(n764));
  jand g380(.dina(n764), .dinb(n762), .dout(n765));
  jxor g381(.dina(n765), .dinb(n761), .dout(f64 ));
  jxor g382(.dina(b65 ), .dinb(a65 ), .dout(n767));
  jor  g383(.dina(b64 ), .dinb(a64 ), .dout(n768));
  jand g384(.dina(b64 ), .dinb(a64 ), .dout(n769));
  jor  g385(.dina(n765), .dinb(n769), .dout(n770));
  jand g386(.dina(n770), .dinb(n768), .dout(n771));
  jxor g387(.dina(n771), .dinb(n767), .dout(f65 ));
  jxor g388(.dina(b66 ), .dinb(a66 ), .dout(n773));
  jor  g389(.dina(b65 ), .dinb(a65 ), .dout(n774));
  jand g390(.dina(b65 ), .dinb(a65 ), .dout(n775));
  jor  g391(.dina(n771), .dinb(n775), .dout(n776));
  jand g392(.dina(n776), .dinb(n774), .dout(n777));
  jxor g393(.dina(n777), .dinb(n773), .dout(f66 ));
  jxor g394(.dina(b67 ), .dinb(a67 ), .dout(n779));
  jor  g395(.dina(b66 ), .dinb(a66 ), .dout(n780));
  jand g396(.dina(b66 ), .dinb(a66 ), .dout(n781));
  jor  g397(.dina(n777), .dinb(n781), .dout(n782));
  jand g398(.dina(n782), .dinb(n780), .dout(n783));
  jxor g399(.dina(n783), .dinb(n779), .dout(f67 ));
  jxor g400(.dina(b68 ), .dinb(a68 ), .dout(n785));
  jor  g401(.dina(b67 ), .dinb(a67 ), .dout(n786));
  jand g402(.dina(b67 ), .dinb(a67 ), .dout(n787));
  jor  g403(.dina(n783), .dinb(n787), .dout(n788));
  jand g404(.dina(n788), .dinb(n786), .dout(n789));
  jxor g405(.dina(n789), .dinb(n785), .dout(f68 ));
  jxor g406(.dina(b69 ), .dinb(a69 ), .dout(n791));
  jor  g407(.dina(b68 ), .dinb(a68 ), .dout(n792));
  jand g408(.dina(b68 ), .dinb(a68 ), .dout(n793));
  jor  g409(.dina(n789), .dinb(n793), .dout(n794));
  jand g410(.dina(n794), .dinb(n792), .dout(n795));
  jxor g411(.dina(n795), .dinb(n791), .dout(f69 ));
  jxor g412(.dina(b70 ), .dinb(a70 ), .dout(n797));
  jor  g413(.dina(b69 ), .dinb(a69 ), .dout(n798));
  jand g414(.dina(b69 ), .dinb(a69 ), .dout(n799));
  jor  g415(.dina(n795), .dinb(n799), .dout(n800));
  jand g416(.dina(n800), .dinb(n798), .dout(n801));
  jxor g417(.dina(n801), .dinb(n797), .dout(f70 ));
  jxor g418(.dina(b71 ), .dinb(a71 ), .dout(n803));
  jor  g419(.dina(b70 ), .dinb(a70 ), .dout(n804));
  jand g420(.dina(b70 ), .dinb(a70 ), .dout(n805));
  jor  g421(.dina(n801), .dinb(n805), .dout(n806));
  jand g422(.dina(n806), .dinb(n804), .dout(n807));
  jxor g423(.dina(n807), .dinb(n803), .dout(f71 ));
  jxor g424(.dina(b72 ), .dinb(a72 ), .dout(n809));
  jor  g425(.dina(b71 ), .dinb(a71 ), .dout(n810));
  jand g426(.dina(b71 ), .dinb(a71 ), .dout(n811));
  jor  g427(.dina(n807), .dinb(n811), .dout(n812));
  jand g428(.dina(n812), .dinb(n810), .dout(n813));
  jxor g429(.dina(n813), .dinb(n809), .dout(f72 ));
  jxor g430(.dina(b73 ), .dinb(a73 ), .dout(n815));
  jor  g431(.dina(b72 ), .dinb(a72 ), .dout(n816));
  jand g432(.dina(b72 ), .dinb(a72 ), .dout(n817));
  jor  g433(.dina(n813), .dinb(n817), .dout(n818));
  jand g434(.dina(n818), .dinb(n816), .dout(n819));
  jxor g435(.dina(n819), .dinb(n815), .dout(f73 ));
  jxor g436(.dina(b74 ), .dinb(a74 ), .dout(n821));
  jor  g437(.dina(b73 ), .dinb(a73 ), .dout(n822));
  jand g438(.dina(b73 ), .dinb(a73 ), .dout(n823));
  jor  g439(.dina(n819), .dinb(n823), .dout(n824));
  jand g440(.dina(n824), .dinb(n822), .dout(n825));
  jxor g441(.dina(n825), .dinb(n821), .dout(f74 ));
  jxor g442(.dina(b75 ), .dinb(a75 ), .dout(n827));
  jor  g443(.dina(b74 ), .dinb(a74 ), .dout(n828));
  jand g444(.dina(b74 ), .dinb(a74 ), .dout(n829));
  jor  g445(.dina(n825), .dinb(n829), .dout(n830));
  jand g446(.dina(n830), .dinb(n828), .dout(n831));
  jxor g447(.dina(n831), .dinb(n827), .dout(f75 ));
  jxor g448(.dina(b76 ), .dinb(a76 ), .dout(n833));
  jor  g449(.dina(b75 ), .dinb(a75 ), .dout(n834));
  jand g450(.dina(b75 ), .dinb(a75 ), .dout(n835));
  jor  g451(.dina(n831), .dinb(n835), .dout(n836));
  jand g452(.dina(n836), .dinb(n834), .dout(n837));
  jxor g453(.dina(n837), .dinb(n833), .dout(f76 ));
  jxor g454(.dina(b77 ), .dinb(a77 ), .dout(n839));
  jor  g455(.dina(b76 ), .dinb(a76 ), .dout(n840));
  jand g456(.dina(b76 ), .dinb(a76 ), .dout(n841));
  jor  g457(.dina(n837), .dinb(n841), .dout(n842));
  jand g458(.dina(n842), .dinb(n840), .dout(n843));
  jxor g459(.dina(n843), .dinb(n839), .dout(f77 ));
  jxor g460(.dina(b78 ), .dinb(a78 ), .dout(n845));
  jor  g461(.dina(b77 ), .dinb(a77 ), .dout(n846));
  jand g462(.dina(b77 ), .dinb(a77 ), .dout(n847));
  jor  g463(.dina(n843), .dinb(n847), .dout(n848));
  jand g464(.dina(n848), .dinb(n846), .dout(n849));
  jxor g465(.dina(n849), .dinb(n845), .dout(f78 ));
  jxor g466(.dina(b79 ), .dinb(a79 ), .dout(n851));
  jor  g467(.dina(b78 ), .dinb(a78 ), .dout(n852));
  jand g468(.dina(b78 ), .dinb(a78 ), .dout(n853));
  jor  g469(.dina(n849), .dinb(n853), .dout(n854));
  jand g470(.dina(n854), .dinb(n852), .dout(n855));
  jxor g471(.dina(n855), .dinb(n851), .dout(f79 ));
  jxor g472(.dina(b80 ), .dinb(a80 ), .dout(n857));
  jor  g473(.dina(b79 ), .dinb(a79 ), .dout(n858));
  jand g474(.dina(b79 ), .dinb(a79 ), .dout(n859));
  jor  g475(.dina(n855), .dinb(n859), .dout(n860));
  jand g476(.dina(n860), .dinb(n858), .dout(n861));
  jxor g477(.dina(n861), .dinb(n857), .dout(f80 ));
  jxor g478(.dina(b81 ), .dinb(a81 ), .dout(n863));
  jor  g479(.dina(b80 ), .dinb(a80 ), .dout(n864));
  jand g480(.dina(b80 ), .dinb(a80 ), .dout(n865));
  jor  g481(.dina(n861), .dinb(n865), .dout(n866));
  jand g482(.dina(n866), .dinb(n864), .dout(n867));
  jxor g483(.dina(n867), .dinb(n863), .dout(f81 ));
  jxor g484(.dina(b82 ), .dinb(a82 ), .dout(n869));
  jor  g485(.dina(b81 ), .dinb(a81 ), .dout(n870));
  jand g486(.dina(b81 ), .dinb(a81 ), .dout(n871));
  jor  g487(.dina(n867), .dinb(n871), .dout(n872));
  jand g488(.dina(n872), .dinb(n870), .dout(n873));
  jxor g489(.dina(n873), .dinb(n869), .dout(f82 ));
  jxor g490(.dina(b83 ), .dinb(a83 ), .dout(n875));
  jor  g491(.dina(b82 ), .dinb(a82 ), .dout(n876));
  jand g492(.dina(b82 ), .dinb(a82 ), .dout(n877));
  jor  g493(.dina(n873), .dinb(n877), .dout(n878));
  jand g494(.dina(n878), .dinb(n876), .dout(n879));
  jxor g495(.dina(n879), .dinb(n875), .dout(f83 ));
  jxor g496(.dina(b84 ), .dinb(a84 ), .dout(n881));
  jor  g497(.dina(b83 ), .dinb(a83 ), .dout(n882));
  jand g498(.dina(b83 ), .dinb(a83 ), .dout(n883));
  jor  g499(.dina(n879), .dinb(n883), .dout(n884));
  jand g500(.dina(n884), .dinb(n882), .dout(n885));
  jxor g501(.dina(n885), .dinb(n881), .dout(f84 ));
  jxor g502(.dina(b85 ), .dinb(a85 ), .dout(n887));
  jor  g503(.dina(b84 ), .dinb(a84 ), .dout(n888));
  jand g504(.dina(b84 ), .dinb(a84 ), .dout(n889));
  jor  g505(.dina(n885), .dinb(n889), .dout(n890));
  jand g506(.dina(n890), .dinb(n888), .dout(n891));
  jxor g507(.dina(n891), .dinb(n887), .dout(f85 ));
  jxor g508(.dina(b86 ), .dinb(a86 ), .dout(n893));
  jor  g509(.dina(b85 ), .dinb(a85 ), .dout(n894));
  jand g510(.dina(b85 ), .dinb(a85 ), .dout(n895));
  jor  g511(.dina(n891), .dinb(n895), .dout(n896));
  jand g512(.dina(n896), .dinb(n894), .dout(n897));
  jxor g513(.dina(n897), .dinb(n893), .dout(f86 ));
  jxor g514(.dina(b87 ), .dinb(a87 ), .dout(n899));
  jor  g515(.dina(b86 ), .dinb(a86 ), .dout(n900));
  jand g516(.dina(b86 ), .dinb(a86 ), .dout(n901));
  jor  g517(.dina(n897), .dinb(n901), .dout(n902));
  jand g518(.dina(n902), .dinb(n900), .dout(n903));
  jxor g519(.dina(n903), .dinb(n899), .dout(f87 ));
  jxor g520(.dina(b88 ), .dinb(a88 ), .dout(n905));
  jor  g521(.dina(b87 ), .dinb(a87 ), .dout(n906));
  jand g522(.dina(b87 ), .dinb(a87 ), .dout(n907));
  jor  g523(.dina(n903), .dinb(n907), .dout(n908));
  jand g524(.dina(n908), .dinb(n906), .dout(n909));
  jxor g525(.dina(n909), .dinb(n905), .dout(f88 ));
  jxor g526(.dina(b89 ), .dinb(a89 ), .dout(n911));
  jor  g527(.dina(b88 ), .dinb(a88 ), .dout(n912));
  jand g528(.dina(b88 ), .dinb(a88 ), .dout(n913));
  jor  g529(.dina(n909), .dinb(n913), .dout(n914));
  jand g530(.dina(n914), .dinb(n912), .dout(n915));
  jxor g531(.dina(n915), .dinb(n911), .dout(f89 ));
  jxor g532(.dina(b90 ), .dinb(a90 ), .dout(n917));
  jor  g533(.dina(b89 ), .dinb(a89 ), .dout(n918));
  jand g534(.dina(b89 ), .dinb(a89 ), .dout(n919));
  jor  g535(.dina(n915), .dinb(n919), .dout(n920));
  jand g536(.dina(n920), .dinb(n918), .dout(n921));
  jxor g537(.dina(n921), .dinb(n917), .dout(f90 ));
  jxor g538(.dina(b91 ), .dinb(a91 ), .dout(n923));
  jor  g539(.dina(b90 ), .dinb(a90 ), .dout(n924));
  jand g540(.dina(b90 ), .dinb(a90 ), .dout(n925));
  jor  g541(.dina(n921), .dinb(n925), .dout(n926));
  jand g542(.dina(n926), .dinb(n924), .dout(n927));
  jxor g543(.dina(n927), .dinb(n923), .dout(f91 ));
  jxor g544(.dina(b92 ), .dinb(a92 ), .dout(n929));
  jor  g545(.dina(b91 ), .dinb(a91 ), .dout(n930));
  jand g546(.dina(b91 ), .dinb(a91 ), .dout(n931));
  jor  g547(.dina(n927), .dinb(n931), .dout(n932));
  jand g548(.dina(n932), .dinb(n930), .dout(n933));
  jxor g549(.dina(n933), .dinb(n929), .dout(f92 ));
  jxor g550(.dina(b93 ), .dinb(a93 ), .dout(n935));
  jor  g551(.dina(b92 ), .dinb(a92 ), .dout(n936));
  jand g552(.dina(b92 ), .dinb(a92 ), .dout(n937));
  jor  g553(.dina(n933), .dinb(n937), .dout(n938));
  jand g554(.dina(n938), .dinb(n936), .dout(n939));
  jxor g555(.dina(n939), .dinb(n935), .dout(f93 ));
  jxor g556(.dina(b94 ), .dinb(a94 ), .dout(n941));
  jor  g557(.dina(b93 ), .dinb(a93 ), .dout(n942));
  jand g558(.dina(b93 ), .dinb(a93 ), .dout(n943));
  jor  g559(.dina(n939), .dinb(n943), .dout(n944));
  jand g560(.dina(n944), .dinb(n942), .dout(n945));
  jxor g561(.dina(n945), .dinb(n941), .dout(f94 ));
  jxor g562(.dina(b95 ), .dinb(a95 ), .dout(n947));
  jor  g563(.dina(b94 ), .dinb(a94 ), .dout(n948));
  jand g564(.dina(b94 ), .dinb(a94 ), .dout(n949));
  jor  g565(.dina(n945), .dinb(n949), .dout(n950));
  jand g566(.dina(n950), .dinb(n948), .dout(n951));
  jxor g567(.dina(n951), .dinb(n947), .dout(f95 ));
  jxor g568(.dina(b96 ), .dinb(a96 ), .dout(n953));
  jor  g569(.dina(b95 ), .dinb(a95 ), .dout(n954));
  jand g570(.dina(b95 ), .dinb(a95 ), .dout(n955));
  jor  g571(.dina(n951), .dinb(n955), .dout(n956));
  jand g572(.dina(n956), .dinb(n954), .dout(n957));
  jxor g573(.dina(n957), .dinb(n953), .dout(f96 ));
  jxor g574(.dina(b97 ), .dinb(a97 ), .dout(n959));
  jor  g575(.dina(b96 ), .dinb(a96 ), .dout(n960));
  jand g576(.dina(b96 ), .dinb(a96 ), .dout(n961));
  jor  g577(.dina(n957), .dinb(n961), .dout(n962));
  jand g578(.dina(n962), .dinb(n960), .dout(n963));
  jxor g579(.dina(n963), .dinb(n959), .dout(f97 ));
  jxor g580(.dina(b98 ), .dinb(a98 ), .dout(n965));
  jor  g581(.dina(b97 ), .dinb(a97 ), .dout(n966));
  jand g582(.dina(b97 ), .dinb(a97 ), .dout(n967));
  jor  g583(.dina(n963), .dinb(n967), .dout(n968));
  jand g584(.dina(n968), .dinb(n966), .dout(n969));
  jxor g585(.dina(n969), .dinb(n965), .dout(f98 ));
  jxor g586(.dina(b99 ), .dinb(a99 ), .dout(n971));
  jor  g587(.dina(b98 ), .dinb(a98 ), .dout(n972));
  jand g588(.dina(b98 ), .dinb(a98 ), .dout(n973));
  jor  g589(.dina(n969), .dinb(n973), .dout(n974));
  jand g590(.dina(n974), .dinb(n972), .dout(n975));
  jxor g591(.dina(n975), .dinb(n971), .dout(f99 ));
  jxor g592(.dina(b100 ), .dinb(a100 ), .dout(n977));
  jor  g593(.dina(b99 ), .dinb(a99 ), .dout(n978));
  jand g594(.dina(b99 ), .dinb(a99 ), .dout(n979));
  jor  g595(.dina(n975), .dinb(n979), .dout(n980));
  jand g596(.dina(n980), .dinb(n978), .dout(n981));
  jxor g597(.dina(n981), .dinb(n977), .dout(f100 ));
  jxor g598(.dina(b101 ), .dinb(a101 ), .dout(n983));
  jor  g599(.dina(b100 ), .dinb(a100 ), .dout(n984));
  jand g600(.dina(b100 ), .dinb(a100 ), .dout(n985));
  jor  g601(.dina(n981), .dinb(n985), .dout(n986));
  jand g602(.dina(n986), .dinb(n984), .dout(n987));
  jxor g603(.dina(n987), .dinb(n983), .dout(f101 ));
  jxor g604(.dina(b102 ), .dinb(a102 ), .dout(n989));
  jor  g605(.dina(b101 ), .dinb(a101 ), .dout(n990));
  jand g606(.dina(b101 ), .dinb(a101 ), .dout(n991));
  jor  g607(.dina(n987), .dinb(n991), .dout(n992));
  jand g608(.dina(n992), .dinb(n990), .dout(n993));
  jxor g609(.dina(n993), .dinb(n989), .dout(f102 ));
  jxor g610(.dina(b103 ), .dinb(a103 ), .dout(n995));
  jor  g611(.dina(b102 ), .dinb(a102 ), .dout(n996));
  jand g612(.dina(b102 ), .dinb(a102 ), .dout(n997));
  jor  g613(.dina(n993), .dinb(n997), .dout(n998));
  jand g614(.dina(n998), .dinb(n996), .dout(n999));
  jxor g615(.dina(n999), .dinb(n995), .dout(f103 ));
  jxor g616(.dina(b104 ), .dinb(a104 ), .dout(n1001));
  jor  g617(.dina(b103 ), .dinb(a103 ), .dout(n1002));
  jand g618(.dina(b103 ), .dinb(a103 ), .dout(n1003));
  jor  g619(.dina(n999), .dinb(n1003), .dout(n1004));
  jand g620(.dina(n1004), .dinb(n1002), .dout(n1005));
  jxor g621(.dina(n1005), .dinb(n1001), .dout(f104 ));
  jxor g622(.dina(b105 ), .dinb(a105 ), .dout(n1007));
  jor  g623(.dina(b104 ), .dinb(a104 ), .dout(n1008));
  jand g624(.dina(b104 ), .dinb(a104 ), .dout(n1009));
  jor  g625(.dina(n1005), .dinb(n1009), .dout(n1010));
  jand g626(.dina(n1010), .dinb(n1008), .dout(n1011));
  jxor g627(.dina(n1011), .dinb(n1007), .dout(f105 ));
  jxor g628(.dina(b106 ), .dinb(a106 ), .dout(n1013));
  jor  g629(.dina(b105 ), .dinb(a105 ), .dout(n1014));
  jand g630(.dina(b105 ), .dinb(a105 ), .dout(n1015));
  jor  g631(.dina(n1011), .dinb(n1015), .dout(n1016));
  jand g632(.dina(n1016), .dinb(n1014), .dout(n1017));
  jxor g633(.dina(n1017), .dinb(n1013), .dout(f106 ));
  jxor g634(.dina(b107 ), .dinb(a107 ), .dout(n1019));
  jor  g635(.dina(b106 ), .dinb(a106 ), .dout(n1020));
  jand g636(.dina(b106 ), .dinb(a106 ), .dout(n1021));
  jor  g637(.dina(n1017), .dinb(n1021), .dout(n1022));
  jand g638(.dina(n1022), .dinb(n1020), .dout(n1023));
  jxor g639(.dina(n1023), .dinb(n1019), .dout(f107 ));
  jxor g640(.dina(b108 ), .dinb(a108 ), .dout(n1025));
  jor  g641(.dina(b107 ), .dinb(a107 ), .dout(n1026));
  jand g642(.dina(b107 ), .dinb(a107 ), .dout(n1027));
  jor  g643(.dina(n1023), .dinb(n1027), .dout(n1028));
  jand g644(.dina(n1028), .dinb(n1026), .dout(n1029));
  jxor g645(.dina(n1029), .dinb(n1025), .dout(f108 ));
  jxor g646(.dina(b109 ), .dinb(a109 ), .dout(n1031));
  jor  g647(.dina(b108 ), .dinb(a108 ), .dout(n1032));
  jand g648(.dina(b108 ), .dinb(a108 ), .dout(n1033));
  jor  g649(.dina(n1029), .dinb(n1033), .dout(n1034));
  jand g650(.dina(n1034), .dinb(n1032), .dout(n1035));
  jxor g651(.dina(n1035), .dinb(n1031), .dout(f109 ));
  jxor g652(.dina(b110 ), .dinb(a110 ), .dout(n1037));
  jor  g653(.dina(b109 ), .dinb(a109 ), .dout(n1038));
  jand g654(.dina(b109 ), .dinb(a109 ), .dout(n1039));
  jor  g655(.dina(n1035), .dinb(n1039), .dout(n1040));
  jand g656(.dina(n1040), .dinb(n1038), .dout(n1041));
  jxor g657(.dina(n1041), .dinb(n1037), .dout(f110 ));
  jxor g658(.dina(b111 ), .dinb(a111 ), .dout(n1043));
  jor  g659(.dina(b110 ), .dinb(a110 ), .dout(n1044));
  jand g660(.dina(b110 ), .dinb(a110 ), .dout(n1045));
  jor  g661(.dina(n1041), .dinb(n1045), .dout(n1046));
  jand g662(.dina(n1046), .dinb(n1044), .dout(n1047));
  jxor g663(.dina(n1047), .dinb(n1043), .dout(f111 ));
  jxor g664(.dina(b112 ), .dinb(a112 ), .dout(n1049));
  jor  g665(.dina(b111 ), .dinb(a111 ), .dout(n1050));
  jand g666(.dina(b111 ), .dinb(a111 ), .dout(n1051));
  jor  g667(.dina(n1047), .dinb(n1051), .dout(n1052));
  jand g668(.dina(n1052), .dinb(n1050), .dout(n1053));
  jxor g669(.dina(n1053), .dinb(n1049), .dout(f112 ));
  jxor g670(.dina(b113 ), .dinb(a113 ), .dout(n1055));
  jor  g671(.dina(b112 ), .dinb(a112 ), .dout(n1056));
  jand g672(.dina(b112 ), .dinb(a112 ), .dout(n1057));
  jor  g673(.dina(n1053), .dinb(n1057), .dout(n1058));
  jand g674(.dina(n1058), .dinb(n1056), .dout(n1059));
  jxor g675(.dina(n1059), .dinb(n1055), .dout(f113 ));
  jxor g676(.dina(b114 ), .dinb(a114 ), .dout(n1061));
  jor  g677(.dina(b113 ), .dinb(a113 ), .dout(n1062));
  jand g678(.dina(b113 ), .dinb(a113 ), .dout(n1063));
  jor  g679(.dina(n1059), .dinb(n1063), .dout(n1064));
  jand g680(.dina(n1064), .dinb(n1062), .dout(n1065));
  jxor g681(.dina(n1065), .dinb(n1061), .dout(f114 ));
  jxor g682(.dina(b115 ), .dinb(a115 ), .dout(n1067));
  jor  g683(.dina(b114 ), .dinb(a114 ), .dout(n1068));
  jand g684(.dina(b114 ), .dinb(a114 ), .dout(n1069));
  jor  g685(.dina(n1065), .dinb(n1069), .dout(n1070));
  jand g686(.dina(n1070), .dinb(n1068), .dout(n1071));
  jxor g687(.dina(n1071), .dinb(n1067), .dout(f115 ));
  jxor g688(.dina(b116 ), .dinb(a116 ), .dout(n1073));
  jor  g689(.dina(b115 ), .dinb(a115 ), .dout(n1074));
  jand g690(.dina(b115 ), .dinb(a115 ), .dout(n1075));
  jor  g691(.dina(n1071), .dinb(n1075), .dout(n1076));
  jand g692(.dina(n1076), .dinb(n1074), .dout(n1077));
  jxor g693(.dina(n1077), .dinb(n1073), .dout(f116 ));
  jxor g694(.dina(b117 ), .dinb(a117 ), .dout(n1079));
  jor  g695(.dina(b116 ), .dinb(a116 ), .dout(n1080));
  jand g696(.dina(b116 ), .dinb(a116 ), .dout(n1081));
  jor  g697(.dina(n1077), .dinb(n1081), .dout(n1082));
  jand g698(.dina(n1082), .dinb(n1080), .dout(n1083));
  jxor g699(.dina(n1083), .dinb(n1079), .dout(f117 ));
  jxor g700(.dina(b118 ), .dinb(a118 ), .dout(n1085));
  jor  g701(.dina(b117 ), .dinb(a117 ), .dout(n1086));
  jand g702(.dina(b117 ), .dinb(a117 ), .dout(n1087));
  jor  g703(.dina(n1083), .dinb(n1087), .dout(n1088));
  jand g704(.dina(n1088), .dinb(n1086), .dout(n1089));
  jxor g705(.dina(n1089), .dinb(n1085), .dout(f118 ));
  jxor g706(.dina(b119 ), .dinb(a119 ), .dout(n1091));
  jor  g707(.dina(b118 ), .dinb(a118 ), .dout(n1092));
  jand g708(.dina(b118 ), .dinb(a118 ), .dout(n1093));
  jor  g709(.dina(n1089), .dinb(n1093), .dout(n1094));
  jand g710(.dina(n1094), .dinb(n1092), .dout(n1095));
  jxor g711(.dina(n1095), .dinb(n1091), .dout(f119 ));
  jxor g712(.dina(b120 ), .dinb(a120 ), .dout(n1097));
  jor  g713(.dina(b119 ), .dinb(a119 ), .dout(n1098));
  jand g714(.dina(b119 ), .dinb(a119 ), .dout(n1099));
  jor  g715(.dina(n1095), .dinb(n1099), .dout(n1100));
  jand g716(.dina(n1100), .dinb(n1098), .dout(n1101));
  jxor g717(.dina(n1101), .dinb(n1097), .dout(f120 ));
  jxor g718(.dina(b121 ), .dinb(a121 ), .dout(n1103));
  jor  g719(.dina(b120 ), .dinb(a120 ), .dout(n1104));
  jand g720(.dina(b120 ), .dinb(a120 ), .dout(n1105));
  jor  g721(.dina(n1101), .dinb(n1105), .dout(n1106));
  jand g722(.dina(n1106), .dinb(n1104), .dout(n1107));
  jxor g723(.dina(n1107), .dinb(n1103), .dout(f121 ));
  jxor g724(.dina(b122 ), .dinb(a122 ), .dout(n1109));
  jor  g725(.dina(b121 ), .dinb(a121 ), .dout(n1110));
  jand g726(.dina(b121 ), .dinb(a121 ), .dout(n1111));
  jor  g727(.dina(n1107), .dinb(n1111), .dout(n1112));
  jand g728(.dina(n1112), .dinb(n1110), .dout(n1113));
  jxor g729(.dina(n1113), .dinb(n1109), .dout(f122 ));
  jxor g730(.dina(b123 ), .dinb(a123 ), .dout(n1115));
  jor  g731(.dina(b122 ), .dinb(a122 ), .dout(n1116));
  jand g732(.dina(b122 ), .dinb(a122 ), .dout(n1117));
  jor  g733(.dina(n1113), .dinb(n1117), .dout(n1118));
  jand g734(.dina(n1118), .dinb(n1116), .dout(n1119));
  jxor g735(.dina(n1119), .dinb(n1115), .dout(f123 ));
  jxor g736(.dina(b124 ), .dinb(a124 ), .dout(n1121));
  jor  g737(.dina(b123 ), .dinb(a123 ), .dout(n1122));
  jand g738(.dina(b123 ), .dinb(a123 ), .dout(n1123));
  jor  g739(.dina(n1119), .dinb(n1123), .dout(n1124));
  jand g740(.dina(n1124), .dinb(n1122), .dout(n1125));
  jxor g741(.dina(n1125), .dinb(n1121), .dout(f124 ));
  jxor g742(.dina(b125 ), .dinb(a125 ), .dout(n1127));
  jor  g743(.dina(b124 ), .dinb(a124 ), .dout(n1128));
  jand g744(.dina(b124 ), .dinb(a124 ), .dout(n1129));
  jor  g745(.dina(n1125), .dinb(n1129), .dout(n1130));
  jand g746(.dina(n1130), .dinb(n1128), .dout(n1131));
  jxor g747(.dina(n1131), .dinb(n1127), .dout(f125 ));
  jxor g748(.dina(b126 ), .dinb(a126 ), .dout(n1133));
  jor  g749(.dina(b125 ), .dinb(a125 ), .dout(n1134));
  jand g750(.dina(b125 ), .dinb(a125 ), .dout(n1135));
  jor  g751(.dina(n1131), .dinb(n1135), .dout(n1136));
  jand g752(.dina(n1136), .dinb(n1134), .dout(n1137));
  jxor g753(.dina(n1137), .dinb(n1133), .dout(f126 ));
  jxor g754(.dina(b127 ), .dinb(a127 ), .dout(n1139));
  jor  g755(.dina(b126 ), .dinb(a126 ), .dout(n1140));
  jand g756(.dina(b126 ), .dinb(a126 ), .dout(n1141));
  jor  g757(.dina(n1137), .dinb(n1141), .dout(n1142));
  jand g758(.dina(n1142), .dinb(n1140), .dout(n1143));
  jxor g759(.dina(n1143), .dinb(n1139), .dout(f127 ));
  jor  g760(.dina(b127 ), .dinb(a127 ), .dout(n1145));
  jand g761(.dina(b127 ), .dinb(a127 ), .dout(n1146));
  jor  g762(.dina(n1143), .dinb(n1146), .dout(n1147));
  jand g763(.dina(n1147), .dinb(n1145), .dout(cOut));
endmodule


