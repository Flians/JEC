/*
rf_c6288:
	jxor: 446
	jspl: 940
	jspl3: 260
	jnot: 330
	jdff: 8448
	jand: 683
	jor: 331

Summary:
	jxor: 446
	jspl: 940
	jspl3: 260
	jnot: 330
	jdff: 8448
	jand: 683
	jor: 331

The maximum logic level gap of any gate:
	rf_c6288: 60
*/

module rf_c6288(gclk, G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat, G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat, G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat, G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat, G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat, G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat, G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat, G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat, G6270gat, G6280gat, G6287gat, G6288gat);
	input gclk;
	input G1gat;
	input G18gat;
	input G35gat;
	input G52gat;
	input G69gat;
	input G86gat;
	input G103gat;
	input G120gat;
	input G137gat;
	input G154gat;
	input G171gat;
	input G188gat;
	input G205gat;
	input G222gat;
	input G239gat;
	input G256gat;
	input G273gat;
	input G290gat;
	input G307gat;
	input G324gat;
	input G341gat;
	input G358gat;
	input G375gat;
	input G392gat;
	input G409gat;
	input G426gat;
	input G443gat;
	input G460gat;
	input G477gat;
	input G494gat;
	input G511gat;
	input G528gat;
	output G545gat;
	output G1581gat;
	output G1901gat;
	output G2223gat;
	output G2548gat;
	output G2877gat;
	output G3211gat;
	output G3552gat;
	output G3895gat;
	output G4241gat;
	output G4591gat;
	output G4946gat;
	output G5308gat;
	output G5672gat;
	output G5971gat;
	output G6123gat;
	output G6150gat;
	output G6160gat;
	output G6170gat;
	output G6180gat;
	output G6190gat;
	output G6200gat;
	output G6210gat;
	output G6220gat;
	output G6230gat;
	output G6240gat;
	output G6250gat;
	output G6260gat;
	output G6270gat;
	output G6280gat;
	output G6287gat;
	output G6288gat;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n69;
	wire n70;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1667;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1684;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1690;
	wire n1691;
	wire n1692;
	wire n1693;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1707;
	wire n1708;
	wire n1709;
	wire n1710;
	wire n1711;
	wire n1712;
	wire n1713;
	wire n1714;
	wire n1715;
	wire n1716;
	wire n1717;
	wire n1718;
	wire n1719;
	wire n1720;
	wire n1722;
	wire n1723;
	wire n1724;
	wire n1725;
	wire n1726;
	wire n1727;
	wire n1728;
	wire n1729;
	wire n1730;
	wire n1731;
	wire n1732;
	wire n1733;
	wire n1734;
	wire n1735;
	wire n1736;
	wire n1737;
	wire n1738;
	wire n1739;
	wire n1740;
	wire n1741;
	wire n1742;
	wire n1743;
	wire n1744;
	wire n1745;
	wire n1746;
	wire n1747;
	wire n1748;
	wire n1749;
	wire n1750;
	wire n1751;
	wire n1752;
	wire n1753;
	wire n1754;
	wire n1755;
	wire n1756;
	wire n1757;
	wire n1758;
	wire n1760;
	wire n1761;
	wire n1762;
	wire n1763;
	wire n1764;
	wire n1765;
	wire n1766;
	wire n1767;
	wire n1768;
	wire n1769;
	wire n1770;
	wire n1771;
	wire n1772;
	wire n1773;
	wire n1774;
	wire n1775;
	wire n1776;
	wire n1777;
	wire n1778;
	wire n1779;
	wire n1780;
	wire n1781;
	wire n1782;
	wire n1783;
	wire n1784;
	wire n1785;
	wire n1786;
	wire n1787;
	wire n1788;
	wire n1789;
	wire n1790;
	wire n1791;
	wire n1793;
	wire n1794;
	wire n1795;
	wire n1796;
	wire n1797;
	wire n1798;
	wire n1799;
	wire n1800;
	wire n1801;
	wire n1802;
	wire n1803;
	wire n1804;
	wire n1805;
	wire n1806;
	wire n1807;
	wire n1808;
	wire n1809;
	wire n1810;
	wire n1811;
	wire n1812;
	wire n1813;
	wire n1814;
	wire n1815;
	wire n1816;
	wire n1817;
	wire n1819;
	wire n1820;
	wire n1821;
	wire n1822;
	wire n1823;
	wire n1824;
	wire n1825;
	wire n1826;
	wire n1827;
	wire n1828;
	wire n1829;
	wire n1830;
	wire n1831;
	wire n1832;
	wire n1833;
	wire n1834;
	wire n1835;
	wire n1836;
	wire n1838;
	wire n1839;
	wire n1840;
	wire n1841;
	wire n1842;
	wire n1843;
	wire n1844;
	wire n1845;
	wire n1846;
	wire n1847;
	wire n1848;
	wire n1849;
	wire n1850;
	wire n1851;
	wire [2:0] w_G1gat_0;
	wire [2:0] w_G1gat_1;
	wire [2:0] w_G1gat_2;
	wire [2:0] w_G1gat_3;
	wire [2:0] w_G1gat_4;
	wire [2:0] w_G1gat_5;
	wire [2:0] w_G1gat_6;
	wire [1:0] w_G1gat_7;
	wire [2:0] w_G18gat_0;
	wire [2:0] w_G18gat_1;
	wire [2:0] w_G18gat_2;
	wire [2:0] w_G18gat_3;
	wire [2:0] w_G18gat_4;
	wire [2:0] w_G18gat_5;
	wire [2:0] w_G18gat_6;
	wire [2:0] w_G18gat_7;
	wire [2:0] w_G35gat_0;
	wire [2:0] w_G35gat_1;
	wire [2:0] w_G35gat_2;
	wire [2:0] w_G35gat_3;
	wire [2:0] w_G35gat_4;
	wire [2:0] w_G35gat_5;
	wire [2:0] w_G35gat_6;
	wire [2:0] w_G35gat_7;
	wire [2:0] w_G52gat_0;
	wire [2:0] w_G52gat_1;
	wire [2:0] w_G52gat_2;
	wire [2:0] w_G52gat_3;
	wire [2:0] w_G52gat_4;
	wire [2:0] w_G52gat_5;
	wire [2:0] w_G52gat_6;
	wire [2:0] w_G52gat_7;
	wire [2:0] w_G69gat_0;
	wire [2:0] w_G69gat_1;
	wire [2:0] w_G69gat_2;
	wire [2:0] w_G69gat_3;
	wire [2:0] w_G69gat_4;
	wire [2:0] w_G69gat_5;
	wire [2:0] w_G69gat_6;
	wire [1:0] w_G69gat_7;
	wire [2:0] w_G86gat_0;
	wire [2:0] w_G86gat_1;
	wire [2:0] w_G86gat_2;
	wire [2:0] w_G86gat_3;
	wire [2:0] w_G86gat_4;
	wire [2:0] w_G86gat_5;
	wire [2:0] w_G86gat_6;
	wire [1:0] w_G86gat_7;
	wire [2:0] w_G103gat_0;
	wire [2:0] w_G103gat_1;
	wire [2:0] w_G103gat_2;
	wire [2:0] w_G103gat_3;
	wire [2:0] w_G103gat_4;
	wire [2:0] w_G103gat_5;
	wire [2:0] w_G103gat_6;
	wire [1:0] w_G103gat_7;
	wire [2:0] w_G120gat_0;
	wire [2:0] w_G120gat_1;
	wire [2:0] w_G120gat_2;
	wire [2:0] w_G120gat_3;
	wire [2:0] w_G120gat_4;
	wire [2:0] w_G120gat_5;
	wire [2:0] w_G120gat_6;
	wire [1:0] w_G120gat_7;
	wire [2:0] w_G137gat_0;
	wire [2:0] w_G137gat_1;
	wire [2:0] w_G137gat_2;
	wire [2:0] w_G137gat_3;
	wire [2:0] w_G137gat_4;
	wire [2:0] w_G137gat_5;
	wire [2:0] w_G137gat_6;
	wire [1:0] w_G137gat_7;
	wire [2:0] w_G154gat_0;
	wire [2:0] w_G154gat_1;
	wire [2:0] w_G154gat_2;
	wire [2:0] w_G154gat_3;
	wire [2:0] w_G154gat_4;
	wire [2:0] w_G154gat_5;
	wire [2:0] w_G154gat_6;
	wire [1:0] w_G154gat_7;
	wire [2:0] w_G171gat_0;
	wire [2:0] w_G171gat_1;
	wire [2:0] w_G171gat_2;
	wire [2:0] w_G171gat_3;
	wire [2:0] w_G171gat_4;
	wire [2:0] w_G171gat_5;
	wire [2:0] w_G171gat_6;
	wire [1:0] w_G171gat_7;
	wire [2:0] w_G188gat_0;
	wire [2:0] w_G188gat_1;
	wire [2:0] w_G188gat_2;
	wire [2:0] w_G188gat_3;
	wire [2:0] w_G188gat_4;
	wire [2:0] w_G188gat_5;
	wire [2:0] w_G188gat_6;
	wire [1:0] w_G188gat_7;
	wire [2:0] w_G205gat_0;
	wire [2:0] w_G205gat_1;
	wire [2:0] w_G205gat_2;
	wire [2:0] w_G205gat_3;
	wire [2:0] w_G205gat_4;
	wire [2:0] w_G205gat_5;
	wire [2:0] w_G205gat_6;
	wire [1:0] w_G205gat_7;
	wire [2:0] w_G222gat_0;
	wire [2:0] w_G222gat_1;
	wire [2:0] w_G222gat_2;
	wire [2:0] w_G222gat_3;
	wire [2:0] w_G222gat_4;
	wire [2:0] w_G222gat_5;
	wire [2:0] w_G222gat_6;
	wire [1:0] w_G222gat_7;
	wire [2:0] w_G239gat_0;
	wire [2:0] w_G239gat_1;
	wire [2:0] w_G239gat_2;
	wire [2:0] w_G239gat_3;
	wire [2:0] w_G239gat_4;
	wire [2:0] w_G239gat_5;
	wire [2:0] w_G239gat_6;
	wire [1:0] w_G239gat_7;
	wire [2:0] w_G256gat_0;
	wire [2:0] w_G256gat_1;
	wire [2:0] w_G256gat_2;
	wire [2:0] w_G256gat_3;
	wire [2:0] w_G256gat_4;
	wire [2:0] w_G256gat_5;
	wire [2:0] w_G256gat_6;
	wire [1:0] w_G256gat_7;
	wire [2:0] w_G273gat_0;
	wire [2:0] w_G273gat_1;
	wire [2:0] w_G273gat_2;
	wire [2:0] w_G273gat_3;
	wire [2:0] w_G273gat_4;
	wire [2:0] w_G273gat_5;
	wire [2:0] w_G273gat_6;
	wire [2:0] w_G273gat_7;
	wire [2:0] w_G290gat_0;
	wire [2:0] w_G290gat_1;
	wire [2:0] w_G290gat_2;
	wire [2:0] w_G290gat_3;
	wire [2:0] w_G290gat_4;
	wire [2:0] w_G290gat_5;
	wire [2:0] w_G290gat_6;
	wire [2:0] w_G290gat_7;
	wire [2:0] w_G307gat_0;
	wire [2:0] w_G307gat_1;
	wire [2:0] w_G307gat_2;
	wire [2:0] w_G307gat_3;
	wire [2:0] w_G307gat_4;
	wire [2:0] w_G307gat_5;
	wire [2:0] w_G307gat_6;
	wire [2:0] w_G307gat_7;
	wire [2:0] w_G324gat_0;
	wire [2:0] w_G324gat_1;
	wire [2:0] w_G324gat_2;
	wire [2:0] w_G324gat_3;
	wire [2:0] w_G324gat_4;
	wire [2:0] w_G324gat_5;
	wire [2:0] w_G324gat_6;
	wire [1:0] w_G324gat_7;
	wire [2:0] w_G341gat_0;
	wire [2:0] w_G341gat_1;
	wire [2:0] w_G341gat_2;
	wire [2:0] w_G341gat_3;
	wire [2:0] w_G341gat_4;
	wire [2:0] w_G341gat_5;
	wire [2:0] w_G341gat_6;
	wire [1:0] w_G341gat_7;
	wire [2:0] w_G358gat_0;
	wire [2:0] w_G358gat_1;
	wire [2:0] w_G358gat_2;
	wire [2:0] w_G358gat_3;
	wire [2:0] w_G358gat_4;
	wire [2:0] w_G358gat_5;
	wire [2:0] w_G358gat_6;
	wire [1:0] w_G358gat_7;
	wire [2:0] w_G375gat_0;
	wire [2:0] w_G375gat_1;
	wire [2:0] w_G375gat_2;
	wire [2:0] w_G375gat_3;
	wire [2:0] w_G375gat_4;
	wire [2:0] w_G375gat_5;
	wire [2:0] w_G375gat_6;
	wire [1:0] w_G375gat_7;
	wire [2:0] w_G392gat_0;
	wire [2:0] w_G392gat_1;
	wire [2:0] w_G392gat_2;
	wire [2:0] w_G392gat_3;
	wire [2:0] w_G392gat_4;
	wire [2:0] w_G392gat_5;
	wire [2:0] w_G392gat_6;
	wire [1:0] w_G392gat_7;
	wire [2:0] w_G409gat_0;
	wire [2:0] w_G409gat_1;
	wire [2:0] w_G409gat_2;
	wire [2:0] w_G409gat_3;
	wire [2:0] w_G409gat_4;
	wire [2:0] w_G409gat_5;
	wire [2:0] w_G409gat_6;
	wire [1:0] w_G409gat_7;
	wire [2:0] w_G426gat_0;
	wire [2:0] w_G426gat_1;
	wire [2:0] w_G426gat_2;
	wire [2:0] w_G426gat_3;
	wire [2:0] w_G426gat_4;
	wire [2:0] w_G426gat_5;
	wire [2:0] w_G426gat_6;
	wire [1:0] w_G426gat_7;
	wire [2:0] w_G443gat_0;
	wire [2:0] w_G443gat_1;
	wire [2:0] w_G443gat_2;
	wire [2:0] w_G443gat_3;
	wire [2:0] w_G443gat_4;
	wire [2:0] w_G443gat_5;
	wire [2:0] w_G443gat_6;
	wire [1:0] w_G443gat_7;
	wire [2:0] w_G460gat_0;
	wire [2:0] w_G460gat_1;
	wire [2:0] w_G460gat_2;
	wire [2:0] w_G460gat_3;
	wire [2:0] w_G460gat_4;
	wire [2:0] w_G460gat_5;
	wire [2:0] w_G460gat_6;
	wire [1:0] w_G460gat_7;
	wire [2:0] w_G477gat_0;
	wire [2:0] w_G477gat_1;
	wire [2:0] w_G477gat_2;
	wire [2:0] w_G477gat_3;
	wire [2:0] w_G477gat_4;
	wire [2:0] w_G477gat_5;
	wire [2:0] w_G477gat_6;
	wire [1:0] w_G477gat_7;
	wire [2:0] w_G494gat_0;
	wire [2:0] w_G494gat_1;
	wire [2:0] w_G494gat_2;
	wire [2:0] w_G494gat_3;
	wire [2:0] w_G494gat_4;
	wire [2:0] w_G494gat_5;
	wire [2:0] w_G494gat_6;
	wire [1:0] w_G494gat_7;
	wire [2:0] w_G511gat_0;
	wire [2:0] w_G511gat_1;
	wire [2:0] w_G511gat_2;
	wire [2:0] w_G511gat_3;
	wire [2:0] w_G511gat_4;
	wire [2:0] w_G511gat_5;
	wire [2:0] w_G511gat_6;
	wire [1:0] w_G511gat_7;
	wire [2:0] w_G528gat_0;
	wire [2:0] w_G528gat_1;
	wire [2:0] w_G528gat_2;
	wire [2:0] w_G528gat_3;
	wire [2:0] w_G528gat_4;
	wire [2:0] w_G528gat_5;
	wire [2:0] w_G528gat_6;
	wire [1:0] w_G528gat_7;
	wire w_G545gat_0;
	wire G545gat_fa_;
	wire [1:0] w_n65_0;
	wire [1:0] w_n69_0;
	wire [1:0] w_n70_0;
	wire [1:0] w_n72_0;
	wire [1:0] w_n75_0;
	wire [1:0] w_n77_0;
	wire [1:0] w_n78_0;
	wire [1:0] w_n81_0;
	wire [2:0] w_n82_0;
	wire [1:0] w_n82_1;
	wire [1:0] w_n84_0;
	wire [1:0] w_n85_0;
	wire [1:0] w_n87_0;
	wire [1:0] w_n89_0;
	wire [1:0] w_n93_0;
	wire [1:0] w_n94_0;
	wire [1:0] w_n96_0;
	wire [1:0] w_n99_0;
	wire [2:0] w_n100_0;
	wire [1:0] w_n100_1;
	wire [2:0] w_n101_0;
	wire [1:0] w_n103_0;
	wire [1:0] w_n104_0;
	wire [1:0] w_n107_0;
	wire [1:0] w_n108_0;
	wire [1:0] w_n110_0;
	wire [1:0] w_n115_0;
	wire [1:0] w_n116_0;
	wire [2:0] w_n126_0;
	wire [1:0] w_n128_0;
	wire [1:0] w_n129_0;
	wire [1:0] w_n130_0;
	wire [1:0] w_n131_0;
	wire [2:0] w_n132_0;
	wire [2:0] w_n133_0;
	wire [1:0] w_n138_0;
	wire [1:0] w_n139_0;
	wire [1:0] w_n140_0;
	wire [1:0] w_n142_0;
	wire [1:0] w_n143_0;
	wire [1:0] w_n145_0;
	wire [1:0] w_n150_0;
	wire [1:0] w_n151_0;
	wire [2:0] w_n156_0;
	wire [1:0] w_n158_0;
	wire [1:0] w_n163_0;
	wire [1:0] w_n165_0;
	wire [1:0] w_n166_0;
	wire [1:0] w_n168_0;
	wire [2:0] w_n169_0;
	wire [1:0] w_n170_0;
	wire [1:0] w_n172_0;
	wire [1:0] w_n174_0;
	wire [1:0] w_n175_0;
	wire [1:0] w_n176_0;
	wire [1:0] w_n177_0;
	wire [1:0] w_n178_0;
	wire [1:0] w_n180_0;
	wire [1:0] w_n181_0;
	wire [1:0] w_n183_0;
	wire [1:0] w_n188_0;
	wire [1:0] w_n189_0;
	wire [2:0] w_n194_0;
	wire [1:0] w_n196_0;
	wire [1:0] w_n199_0;
	wire [1:0] w_n201_0;
	wire [1:0] w_n204_0;
	wire [1:0] w_n206_0;
	wire [1:0] w_n207_0;
	wire [1:0] w_n209_0;
	wire [2:0] w_n210_0;
	wire [1:0] w_n210_1;
	wire [1:0] w_n213_0;
	wire [1:0] w_n215_0;
	wire [1:0] w_n216_0;
	wire [1:0] w_n217_0;
	wire [1:0] w_n218_0;
	wire [1:0] w_n219_0;
	wire [1:0] w_n220_0;
	wire [1:0] w_n221_0;
	wire [1:0] w_n223_0;
	wire [1:0] w_n224_0;
	wire [1:0] w_n226_0;
	wire [1:0] w_n231_0;
	wire [1:0] w_n232_0;
	wire [2:0] w_n237_0;
	wire [1:0] w_n239_0;
	wire [1:0] w_n242_0;
	wire [1:0] w_n244_0;
	wire [1:0] w_n247_0;
	wire [1:0] w_n249_0;
	wire [1:0] w_n252_0;
	wire [1:0] w_n254_0;
	wire [1:0] w_n255_0;
	wire [1:0] w_n257_0;
	wire [2:0] w_n258_0;
	wire [1:0] w_n259_0;
	wire [1:0] w_n261_0;
	wire [1:0] w_n264_0;
	wire [1:0] w_n265_0;
	wire [1:0] w_n266_0;
	wire [1:0] w_n267_0;
	wire [1:0] w_n268_0;
	wire [1:0] w_n269_0;
	wire [1:0] w_n270_0;
	wire [1:0] w_n271_0;
	wire [1:0] w_n272_0;
	wire [1:0] w_n274_0;
	wire [1:0] w_n275_0;
	wire [1:0] w_n277_0;
	wire [1:0] w_n282_0;
	wire [1:0] w_n283_0;
	wire [2:0] w_n288_0;
	wire [1:0] w_n290_0;
	wire [1:0] w_n293_0;
	wire [1:0] w_n295_0;
	wire [1:0] w_n298_0;
	wire [1:0] w_n300_0;
	wire [1:0] w_n303_0;
	wire [1:0] w_n305_0;
	wire [1:0] w_n308_0;
	wire [1:0] w_n310_0;
	wire [1:0] w_n311_0;
	wire [1:0] w_n313_0;
	wire [2:0] w_n314_0;
	wire [1:0] w_n315_0;
	wire [1:0] w_n317_0;
	wire [1:0] w_n320_0;
	wire [1:0] w_n321_0;
	wire [1:0] w_n322_0;
	wire [1:0] w_n323_0;
	wire [1:0] w_n324_0;
	wire [1:0] w_n325_0;
	wire [1:0] w_n326_0;
	wire [1:0] w_n327_0;
	wire [1:0] w_n328_0;
	wire [1:0] w_n329_0;
	wire [1:0] w_n330_0;
	wire [1:0] w_n332_0;
	wire [1:0] w_n333_0;
	wire [1:0] w_n335_0;
	wire [1:0] w_n340_0;
	wire [1:0] w_n341_0;
	wire [2:0] w_n346_0;
	wire [1:0] w_n348_0;
	wire [1:0] w_n351_0;
	wire [1:0] w_n353_0;
	wire [1:0] w_n356_0;
	wire [1:0] w_n358_0;
	wire [1:0] w_n361_0;
	wire [1:0] w_n363_0;
	wire [1:0] w_n366_0;
	wire [1:0] w_n368_0;
	wire [1:0] w_n371_0;
	wire [1:0] w_n372_0;
	wire [1:0] w_n373_0;
	wire [1:0] w_n375_0;
	wire [2:0] w_n376_0;
	wire [1:0] w_n377_0;
	wire [1:0] w_n380_0;
	wire [1:0] w_n382_0;
	wire [1:0] w_n383_0;
	wire [1:0] w_n384_0;
	wire [1:0] w_n385_0;
	wire [1:0] w_n386_0;
	wire [1:0] w_n387_0;
	wire [1:0] w_n388_0;
	wire [1:0] w_n389_0;
	wire [1:0] w_n390_0;
	wire [1:0] w_n391_0;
	wire [1:0] w_n392_0;
	wire [1:0] w_n393_0;
	wire [1:0] w_n394_0;
	wire [1:0] w_n396_0;
	wire [1:0] w_n397_0;
	wire [1:0] w_n399_0;
	wire [1:0] w_n404_0;
	wire [1:0] w_n405_0;
	wire [2:0] w_n410_0;
	wire [1:0] w_n412_0;
	wire [1:0] w_n415_0;
	wire [1:0] w_n417_0;
	wire [1:0] w_n420_0;
	wire [1:0] w_n422_0;
	wire [1:0] w_n425_0;
	wire [1:0] w_n427_0;
	wire [1:0] w_n430_0;
	wire [1:0] w_n432_0;
	wire [1:0] w_n435_0;
	wire [1:0] w_n437_0;
	wire [1:0] w_n441_0;
	wire [1:0] w_n442_0;
	wire [1:0] w_n443_0;
	wire [1:0] w_n445_0;
	wire [2:0] w_n446_0;
	wire [1:0] w_n447_0;
	wire [1:0] w_n450_0;
	wire [1:0] w_n452_0;
	wire [1:0] w_n453_0;
	wire [1:0] w_n454_0;
	wire [1:0] w_n455_0;
	wire [1:0] w_n456_0;
	wire [1:0] w_n457_0;
	wire [1:0] w_n458_0;
	wire [1:0] w_n459_0;
	wire [1:0] w_n460_0;
	wire [1:0] w_n461_0;
	wire [1:0] w_n462_0;
	wire [1:0] w_n463_0;
	wire [1:0] w_n464_0;
	wire [1:0] w_n465_0;
	wire [1:0] w_n466_0;
	wire [1:0] w_n468_0;
	wire [1:0] w_n469_0;
	wire [1:0] w_n471_0;
	wire [1:0] w_n476_0;
	wire [1:0] w_n477_0;
	wire [2:0] w_n482_0;
	wire [1:0] w_n484_0;
	wire [1:0] w_n487_0;
	wire [1:0] w_n489_0;
	wire [1:0] w_n492_0;
	wire [1:0] w_n494_0;
	wire [1:0] w_n497_0;
	wire [1:0] w_n499_0;
	wire [1:0] w_n502_0;
	wire [1:0] w_n504_0;
	wire [1:0] w_n507_0;
	wire [1:0] w_n509_0;
	wire [1:0] w_n512_0;
	wire [1:0] w_n514_0;
	wire [1:0] w_n518_0;
	wire [1:0] w_n519_0;
	wire [1:0] w_n520_0;
	wire [1:0] w_n522_0;
	wire [2:0] w_n523_0;
	wire [1:0] w_n524_0;
	wire [1:0] w_n527_0;
	wire [1:0] w_n529_0;
	wire [1:0] w_n530_0;
	wire [1:0] w_n531_0;
	wire [1:0] w_n532_0;
	wire [1:0] w_n533_0;
	wire [1:0] w_n534_0;
	wire [1:0] w_n535_0;
	wire [1:0] w_n536_0;
	wire [1:0] w_n537_0;
	wire [1:0] w_n538_0;
	wire [1:0] w_n539_0;
	wire [1:0] w_n540_0;
	wire [1:0] w_n541_0;
	wire [1:0] w_n542_0;
	wire [1:0] w_n543_0;
	wire [1:0] w_n544_0;
	wire [1:0] w_n545_0;
	wire [1:0] w_n547_0;
	wire [1:0] w_n548_0;
	wire [1:0] w_n550_0;
	wire [1:0] w_n555_0;
	wire [1:0] w_n556_0;
	wire [2:0] w_n561_0;
	wire [1:0] w_n563_0;
	wire [1:0] w_n566_0;
	wire [1:0] w_n568_0;
	wire [1:0] w_n571_0;
	wire [1:0] w_n573_0;
	wire [1:0] w_n576_0;
	wire [1:0] w_n578_0;
	wire [1:0] w_n581_0;
	wire [1:0] w_n583_0;
	wire [1:0] w_n586_0;
	wire [1:0] w_n588_0;
	wire [1:0] w_n591_0;
	wire [1:0] w_n593_0;
	wire [1:0] w_n596_0;
	wire [1:0] w_n598_0;
	wire [1:0] w_n602_0;
	wire [1:0] w_n603_0;
	wire [1:0] w_n604_0;
	wire [1:0] w_n606_0;
	wire [2:0] w_n607_0;
	wire [1:0] w_n608_0;
	wire [1:0] w_n611_0;
	wire [1:0] w_n613_0;
	wire [1:0] w_n614_0;
	wire [1:0] w_n615_0;
	wire [1:0] w_n616_0;
	wire [1:0] w_n617_0;
	wire [1:0] w_n618_0;
	wire [1:0] w_n619_0;
	wire [1:0] w_n620_0;
	wire [1:0] w_n621_0;
	wire [1:0] w_n622_0;
	wire [1:0] w_n623_0;
	wire [1:0] w_n624_0;
	wire [1:0] w_n625_0;
	wire [1:0] w_n626_0;
	wire [1:0] w_n627_0;
	wire [1:0] w_n628_0;
	wire [1:0] w_n629_0;
	wire [1:0] w_n630_0;
	wire [1:0] w_n631_0;
	wire [1:0] w_n633_0;
	wire [1:0] w_n634_0;
	wire [1:0] w_n636_0;
	wire [1:0] w_n641_0;
	wire [1:0] w_n642_0;
	wire [2:0] w_n647_0;
	wire [1:0] w_n649_0;
	wire [1:0] w_n652_0;
	wire [1:0] w_n654_0;
	wire [1:0] w_n657_0;
	wire [1:0] w_n659_0;
	wire [1:0] w_n662_0;
	wire [1:0] w_n664_0;
	wire [1:0] w_n667_0;
	wire [1:0] w_n669_0;
	wire [1:0] w_n672_0;
	wire [1:0] w_n674_0;
	wire [1:0] w_n677_0;
	wire [1:0] w_n679_0;
	wire [1:0] w_n682_0;
	wire [1:0] w_n684_0;
	wire [1:0] w_n687_0;
	wire [1:0] w_n689_0;
	wire [1:0] w_n693_0;
	wire [1:0] w_n694_0;
	wire [2:0] w_n695_0;
	wire [1:0] w_n697_0;
	wire [2:0] w_n698_0;
	wire [1:0] w_n699_0;
	wire [1:0] w_n702_0;
	wire [1:0] w_n704_0;
	wire [1:0] w_n705_0;
	wire [1:0] w_n706_0;
	wire [1:0] w_n707_0;
	wire [1:0] w_n708_0;
	wire [1:0] w_n709_0;
	wire [1:0] w_n710_0;
	wire [1:0] w_n711_0;
	wire [1:0] w_n712_0;
	wire [1:0] w_n713_0;
	wire [1:0] w_n714_0;
	wire [1:0] w_n715_0;
	wire [1:0] w_n716_0;
	wire [1:0] w_n717_0;
	wire [1:0] w_n718_0;
	wire [1:0] w_n719_0;
	wire [1:0] w_n720_0;
	wire [1:0] w_n721_0;
	wire [1:0] w_n722_0;
	wire [1:0] w_n723_0;
	wire [1:0] w_n724_0;
	wire [1:0] w_n726_0;
	wire [1:0] w_n727_0;
	wire [1:0] w_n729_0;
	wire [1:0] w_n734_0;
	wire [1:0] w_n735_0;
	wire [2:0] w_n740_0;
	wire [1:0] w_n742_0;
	wire [1:0] w_n745_0;
	wire [1:0] w_n747_0;
	wire [1:0] w_n750_0;
	wire [1:0] w_n752_0;
	wire [1:0] w_n755_0;
	wire [1:0] w_n757_0;
	wire [1:0] w_n760_0;
	wire [1:0] w_n762_0;
	wire [1:0] w_n765_0;
	wire [1:0] w_n767_0;
	wire [1:0] w_n770_0;
	wire [1:0] w_n772_0;
	wire [1:0] w_n775_0;
	wire [1:0] w_n777_0;
	wire [1:0] w_n780_0;
	wire [1:0] w_n782_0;
	wire [1:0] w_n785_0;
	wire [1:0] w_n787_0;
	wire [1:0] w_n791_0;
	wire [1:0] w_n792_0;
	wire [1:0] w_n793_0;
	wire [1:0] w_n795_0;
	wire [2:0] w_n797_0;
	wire [1:0] w_n800_0;
	wire [1:0] w_n802_0;
	wire [1:0] w_n803_0;
	wire [1:0] w_n804_0;
	wire [1:0] w_n805_0;
	wire [1:0] w_n806_0;
	wire [1:0] w_n807_0;
	wire [1:0] w_n808_0;
	wire [1:0] w_n809_0;
	wire [1:0] w_n810_0;
	wire [1:0] w_n811_0;
	wire [1:0] w_n812_0;
	wire [1:0] w_n813_0;
	wire [1:0] w_n814_0;
	wire [1:0] w_n815_0;
	wire [1:0] w_n816_0;
	wire [1:0] w_n817_0;
	wire [1:0] w_n818_0;
	wire [1:0] w_n819_0;
	wire [1:0] w_n820_0;
	wire [1:0] w_n821_0;
	wire [1:0] w_n822_0;
	wire [1:0] w_n823_0;
	wire [1:0] w_n824_0;
	wire [1:0] w_n826_0;
	wire [1:0] w_n827_0;
	wire [1:0] w_n829_0;
	wire [1:0] w_n834_0;
	wire [1:0] w_n835_0;
	wire [1:0] w_n839_0;
	wire [1:0] w_n840_0;
	wire [2:0] w_n844_0;
	wire [1:0] w_n846_0;
	wire [1:0] w_n849_0;
	wire [1:0] w_n851_0;
	wire [1:0] w_n854_0;
	wire [1:0] w_n856_0;
	wire [1:0] w_n859_0;
	wire [1:0] w_n861_0;
	wire [1:0] w_n864_0;
	wire [1:0] w_n866_0;
	wire [1:0] w_n869_0;
	wire [1:0] w_n871_0;
	wire [1:0] w_n874_0;
	wire [1:0] w_n876_0;
	wire [1:0] w_n879_0;
	wire [1:0] w_n881_0;
	wire [1:0] w_n884_0;
	wire [1:0] w_n886_0;
	wire [1:0] w_n889_0;
	wire [1:0] w_n891_0;
	wire [1:0] w_n895_0;
	wire [1:0] w_n896_0;
	wire [1:0] w_n897_0;
	wire [1:0] w_n898_0;
	wire [1:0] w_n901_0;
	wire [1:0] w_n903_0;
	wire [1:0] w_n906_0;
	wire [1:0] w_n907_0;
	wire [1:0] w_n908_0;
	wire [1:0] w_n909_0;
	wire [1:0] w_n910_0;
	wire [1:0] w_n911_0;
	wire [1:0] w_n912_0;
	wire [1:0] w_n913_0;
	wire [1:0] w_n914_0;
	wire [1:0] w_n915_0;
	wire [1:0] w_n916_0;
	wire [1:0] w_n917_0;
	wire [1:0] w_n918_0;
	wire [1:0] w_n919_0;
	wire [1:0] w_n920_0;
	wire [1:0] w_n921_0;
	wire [1:0] w_n922_0;
	wire [1:0] w_n923_0;
	wire [1:0] w_n924_0;
	wire [1:0] w_n925_0;
	wire [1:0] w_n926_0;
	wire [2:0] w_n927_0;
	wire [1:0] w_n929_0;
	wire [1:0] w_n930_0;
	wire [1:0] w_n931_0;
	wire [1:0] w_n932_0;
	wire [1:0] w_n937_0;
	wire [1:0] w_n938_0;
	wire [2:0] w_n942_0;
	wire [1:0] w_n943_0;
	wire [1:0] w_n949_0;
	wire [1:0] w_n951_0;
	wire [1:0] w_n954_0;
	wire [1:0] w_n956_0;
	wire [1:0] w_n959_0;
	wire [1:0] w_n961_0;
	wire [1:0] w_n964_0;
	wire [1:0] w_n966_0;
	wire [1:0] w_n969_0;
	wire [1:0] w_n971_0;
	wire [1:0] w_n974_0;
	wire [1:0] w_n976_0;
	wire [1:0] w_n979_0;
	wire [1:0] w_n981_0;
	wire [1:0] w_n984_0;
	wire [1:0] w_n986_0;
	wire [1:0] w_n989_0;
	wire [1:0] w_n991_0;
	wire [1:0] w_n994_0;
	wire [1:0] w_n996_0;
	wire [1:0] w_n999_0;
	wire [1:0] w_n1001_0;
	wire [1:0] w_n1005_0;
	wire [1:0] w_n1006_0;
	wire [1:0] w_n1008_0;
	wire [1:0] w_n1009_0;
	wire [1:0] w_n1010_0;
	wire [1:0] w_n1011_0;
	wire [1:0] w_n1012_0;
	wire [1:0] w_n1013_0;
	wire [1:0] w_n1014_0;
	wire [1:0] w_n1015_0;
	wire [1:0] w_n1016_0;
	wire [1:0] w_n1017_0;
	wire [1:0] w_n1018_0;
	wire [1:0] w_n1019_0;
	wire [1:0] w_n1020_0;
	wire [1:0] w_n1021_0;
	wire [1:0] w_n1022_0;
	wire [1:0] w_n1023_0;
	wire [1:0] w_n1024_0;
	wire [1:0] w_n1025_0;
	wire [1:0] w_n1026_0;
	wire [1:0] w_n1027_0;
	wire [1:0] w_n1028_0;
	wire [1:0] w_n1029_0;
	wire [1:0] w_n1030_0;
	wire [1:0] w_n1031_0;
	wire [1:0] w_n1032_0;
	wire [1:0] w_n1033_0;
	wire [1:0] w_n1034_0;
	wire [1:0] w_n1035_0;
	wire [1:0] w_n1037_0;
	wire [1:0] w_n1039_0;
	wire [1:0] w_n1043_0;
	wire [1:0] w_n1044_0;
	wire [1:0] w_n1048_0;
	wire [1:0] w_n1049_0;
	wire [1:0] w_n1052_0;
	wire [1:0] w_n1054_0;
	wire [1:0] w_n1057_0;
	wire [1:0] w_n1059_0;
	wire [1:0] w_n1062_0;
	wire [1:0] w_n1064_0;
	wire [1:0] w_n1067_0;
	wire [1:0] w_n1069_0;
	wire [1:0] w_n1072_0;
	wire [1:0] w_n1074_0;
	wire [1:0] w_n1077_0;
	wire [1:0] w_n1079_0;
	wire [1:0] w_n1082_0;
	wire [1:0] w_n1084_0;
	wire [1:0] w_n1087_0;
	wire [1:0] w_n1089_0;
	wire [1:0] w_n1092_0;
	wire [1:0] w_n1094_0;
	wire [1:0] w_n1097_0;
	wire [1:0] w_n1099_0;
	wire [1:0] w_n1102_0;
	wire [1:0] w_n1103_0;
	wire [1:0] w_n1109_0;
	wire [1:0] w_n1110_0;
	wire [1:0] w_n1114_0;
	wire [1:0] w_n1115_0;
	wire [1:0] w_n1116_0;
	wire [1:0] w_n1117_0;
	wire [1:0] w_n1118_0;
	wire [1:0] w_n1119_0;
	wire [1:0] w_n1120_0;
	wire [1:0] w_n1121_0;
	wire [1:0] w_n1122_0;
	wire [1:0] w_n1123_0;
	wire [1:0] w_n1124_0;
	wire [1:0] w_n1125_0;
	wire [1:0] w_n1126_0;
	wire [1:0] w_n1127_0;
	wire [1:0] w_n1128_0;
	wire [1:0] w_n1129_0;
	wire [1:0] w_n1130_0;
	wire [1:0] w_n1131_0;
	wire [1:0] w_n1132_0;
	wire [1:0] w_n1133_0;
	wire [1:0] w_n1134_0;
	wire [1:0] w_n1135_0;
	wire [1:0] w_n1137_0;
	wire [1:0] w_n1138_0;
	wire [1:0] w_n1139_0;
	wire [1:0] w_n1140_0;
	wire [1:0] w_n1141_0;
	wire [1:0] w_n1147_0;
	wire [1:0] w_n1151_0;
	wire [1:0] w_n1152_0;
	wire [1:0] w_n1156_0;
	wire [1:0] w_n1158_0;
	wire [1:0] w_n1161_0;
	wire [1:0] w_n1163_0;
	wire [1:0] w_n1166_0;
	wire [1:0] w_n1168_0;
	wire [1:0] w_n1171_0;
	wire [1:0] w_n1173_0;
	wire [1:0] w_n1176_0;
	wire [1:0] w_n1178_0;
	wire [1:0] w_n1181_0;
	wire [1:0] w_n1183_0;
	wire [1:0] w_n1186_0;
	wire [1:0] w_n1188_0;
	wire [1:0] w_n1191_0;
	wire [1:0] w_n1193_0;
	wire [1:0] w_n1196_0;
	wire [1:0] w_n1198_0;
	wire [1:0] w_n1201_0;
	wire [1:0] w_n1203_0;
	wire [1:0] w_n1206_0;
	wire [1:0] w_n1207_0;
	wire [1:0] w_n1208_0;
	wire [1:0] w_n1210_0;
	wire [1:0] w_n1212_0;
	wire [1:0] w_n1213_0;
	wire [1:0] w_n1214_0;
	wire [1:0] w_n1215_0;
	wire [1:0] w_n1216_0;
	wire [1:0] w_n1217_0;
	wire [1:0] w_n1218_0;
	wire [1:0] w_n1219_0;
	wire [1:0] w_n1220_0;
	wire [1:0] w_n1221_0;
	wire [1:0] w_n1222_0;
	wire [1:0] w_n1223_0;
	wire [1:0] w_n1224_0;
	wire [1:0] w_n1225_0;
	wire [1:0] w_n1226_0;
	wire [1:0] w_n1227_0;
	wire [1:0] w_n1228_0;
	wire [1:0] w_n1229_0;
	wire [1:0] w_n1230_0;
	wire [1:0] w_n1231_0;
	wire [1:0] w_n1232_0;
	wire [1:0] w_n1234_0;
	wire [1:0] w_n1236_0;
	wire [1:0] w_n1237_0;
	wire [1:0] w_n1238_0;
	wire [1:0] w_n1244_0;
	wire [1:0] w_n1247_0;
	wire [1:0] w_n1248_0;
	wire [1:0] w_n1251_0;
	wire [1:0] w_n1253_0;
	wire [1:0] w_n1256_0;
	wire [1:0] w_n1258_0;
	wire [1:0] w_n1261_0;
	wire [1:0] w_n1263_0;
	wire [1:0] w_n1266_0;
	wire [1:0] w_n1268_0;
	wire [1:0] w_n1271_0;
	wire [1:0] w_n1273_0;
	wire [1:0] w_n1276_0;
	wire [1:0] w_n1278_0;
	wire [1:0] w_n1281_0;
	wire [1:0] w_n1283_0;
	wire [1:0] w_n1286_0;
	wire [1:0] w_n1288_0;
	wire [1:0] w_n1291_0;
	wire [1:0] w_n1293_0;
	wire [1:0] w_n1296_0;
	wire [1:0] w_n1297_0;
	wire [1:0] w_n1298_0;
	wire [1:0] w_n1301_0;
	wire [1:0] w_n1303_0;
	wire [1:0] w_n1304_0;
	wire [1:0] w_n1305_0;
	wire [1:0] w_n1306_0;
	wire [1:0] w_n1307_0;
	wire [1:0] w_n1308_0;
	wire [1:0] w_n1309_0;
	wire [1:0] w_n1310_0;
	wire [1:0] w_n1311_0;
	wire [1:0] w_n1312_0;
	wire [1:0] w_n1313_0;
	wire [1:0] w_n1314_0;
	wire [1:0] w_n1315_0;
	wire [1:0] w_n1316_0;
	wire [1:0] w_n1317_0;
	wire [1:0] w_n1318_0;
	wire [1:0] w_n1319_0;
	wire [1:0] w_n1320_0;
	wire [1:0] w_n1321_0;
	wire [1:0] w_n1322_0;
	wire [1:0] w_n1324_0;
	wire [1:0] w_n1325_0;
	wire [1:0] w_n1326_0;
	wire [1:0] w_n1332_0;
	wire [1:0] w_n1337_0;
	wire [1:0] w_n1338_0;
	wire [1:0] w_n1341_0;
	wire [1:0] w_n1343_0;
	wire [1:0] w_n1346_0;
	wire [1:0] w_n1348_0;
	wire [1:0] w_n1351_0;
	wire [1:0] w_n1353_0;
	wire [1:0] w_n1356_0;
	wire [1:0] w_n1358_0;
	wire [1:0] w_n1361_0;
	wire [1:0] w_n1363_0;
	wire [1:0] w_n1366_0;
	wire [1:0] w_n1368_0;
	wire [1:0] w_n1371_0;
	wire [1:0] w_n1373_0;
	wire [1:0] w_n1376_0;
	wire [1:0] w_n1378_0;
	wire [1:0] w_n1381_0;
	wire [1:0] w_n1382_0;
	wire [1:0] w_n1383_0;
	wire [1:0] w_n1386_0;
	wire [1:0] w_n1388_0;
	wire [1:0] w_n1389_0;
	wire [1:0] w_n1390_0;
	wire [1:0] w_n1391_0;
	wire [1:0] w_n1392_0;
	wire [1:0] w_n1393_0;
	wire [1:0] w_n1394_0;
	wire [1:0] w_n1395_0;
	wire [1:0] w_n1396_0;
	wire [1:0] w_n1397_0;
	wire [1:0] w_n1398_0;
	wire [1:0] w_n1399_0;
	wire [1:0] w_n1400_0;
	wire [1:0] w_n1401_0;
	wire [1:0] w_n1402_0;
	wire [1:0] w_n1403_0;
	wire [1:0] w_n1404_0;
	wire [1:0] w_n1405_0;
	wire [1:0] w_n1407_0;
	wire [1:0] w_n1409_0;
	wire [1:0] w_n1410_0;
	wire [1:0] w_n1415_0;
	wire [1:0] w_n1420_0;
	wire [1:0] w_n1421_0;
	wire [1:0] w_n1424_0;
	wire [1:0] w_n1426_0;
	wire [1:0] w_n1429_0;
	wire [1:0] w_n1431_0;
	wire [1:0] w_n1434_0;
	wire [1:0] w_n1436_0;
	wire [1:0] w_n1439_0;
	wire [1:0] w_n1441_0;
	wire [1:0] w_n1444_0;
	wire [1:0] w_n1446_0;
	wire [1:0] w_n1449_0;
	wire [1:0] w_n1451_0;
	wire [1:0] w_n1454_0;
	wire [1:0] w_n1456_0;
	wire [1:0] w_n1459_0;
	wire [1:0] w_n1460_0;
	wire [1:0] w_n1461_0;
	wire [1:0] w_n1464_0;
	wire [1:0] w_n1466_0;
	wire [1:0] w_n1467_0;
	wire [1:0] w_n1468_0;
	wire [1:0] w_n1469_0;
	wire [1:0] w_n1470_0;
	wire [1:0] w_n1471_0;
	wire [1:0] w_n1472_0;
	wire [1:0] w_n1473_0;
	wire [1:0] w_n1474_0;
	wire [1:0] w_n1475_0;
	wire [1:0] w_n1476_0;
	wire [1:0] w_n1477_0;
	wire [1:0] w_n1478_0;
	wire [1:0] w_n1479_0;
	wire [1:0] w_n1480_0;
	wire [1:0] w_n1481_0;
	wire [1:0] w_n1483_0;
	wire [1:0] w_n1485_0;
	wire [1:0] w_n1486_0;
	wire [1:0] w_n1491_0;
	wire [1:0] w_n1496_0;
	wire [1:0] w_n1497_0;
	wire [1:0] w_n1500_0;
	wire [1:0] w_n1502_0;
	wire [1:0] w_n1505_0;
	wire [1:0] w_n1507_0;
	wire [1:0] w_n1510_0;
	wire [1:0] w_n1512_0;
	wire [1:0] w_n1515_0;
	wire [1:0] w_n1517_0;
	wire [1:0] w_n1520_0;
	wire [1:0] w_n1522_0;
	wire [1:0] w_n1525_0;
	wire [1:0] w_n1527_0;
	wire [1:0] w_n1530_0;
	wire [1:0] w_n1531_0;
	wire [1:0] w_n1532_0;
	wire [1:0] w_n1535_0;
	wire [1:0] w_n1537_0;
	wire [1:0] w_n1538_0;
	wire [1:0] w_n1539_0;
	wire [1:0] w_n1540_0;
	wire [1:0] w_n1541_0;
	wire [1:0] w_n1542_0;
	wire [1:0] w_n1543_0;
	wire [1:0] w_n1544_0;
	wire [1:0] w_n1545_0;
	wire [1:0] w_n1546_0;
	wire [1:0] w_n1547_0;
	wire [1:0] w_n1548_0;
	wire [1:0] w_n1549_0;
	wire [1:0] w_n1550_0;
	wire [1:0] w_n1552_0;
	wire [1:0] w_n1554_0;
	wire [1:0] w_n1555_0;
	wire [1:0] w_n1560_0;
	wire [1:0] w_n1565_0;
	wire [1:0] w_n1566_0;
	wire [1:0] w_n1569_0;
	wire [1:0] w_n1571_0;
	wire [1:0] w_n1574_0;
	wire [1:0] w_n1576_0;
	wire [1:0] w_n1579_0;
	wire [1:0] w_n1581_0;
	wire [1:0] w_n1584_0;
	wire [1:0] w_n1586_0;
	wire [1:0] w_n1589_0;
	wire [1:0] w_n1591_0;
	wire [1:0] w_n1594_0;
	wire [1:0] w_n1595_0;
	wire [1:0] w_n1596_0;
	wire [1:0] w_n1599_0;
	wire [1:0] w_n1601_0;
	wire [1:0] w_n1602_0;
	wire [1:0] w_n1603_0;
	wire [1:0] w_n1604_0;
	wire [1:0] w_n1605_0;
	wire [1:0] w_n1606_0;
	wire [1:0] w_n1607_0;
	wire [1:0] w_n1608_0;
	wire [1:0] w_n1609_0;
	wire [1:0] w_n1610_0;
	wire [1:0] w_n1611_0;
	wire [1:0] w_n1612_0;
	wire [1:0] w_n1614_0;
	wire [1:0] w_n1616_0;
	wire [1:0] w_n1617_0;
	wire [1:0] w_n1622_0;
	wire [1:0] w_n1627_0;
	wire [1:0] w_n1628_0;
	wire [1:0] w_n1631_0;
	wire [1:0] w_n1633_0;
	wire [1:0] w_n1636_0;
	wire [1:0] w_n1638_0;
	wire [1:0] w_n1641_0;
	wire [1:0] w_n1643_0;
	wire [1:0] w_n1646_0;
	wire [1:0] w_n1648_0;
	wire [1:0] w_n1651_0;
	wire [1:0] w_n1652_0;
	wire [1:0] w_n1653_0;
	wire [1:0] w_n1656_0;
	wire [1:0] w_n1658_0;
	wire [1:0] w_n1659_0;
	wire [1:0] w_n1660_0;
	wire [1:0] w_n1661_0;
	wire [1:0] w_n1662_0;
	wire [1:0] w_n1663_0;
	wire [1:0] w_n1664_0;
	wire [1:0] w_n1665_0;
	wire [1:0] w_n1666_0;
	wire [1:0] w_n1667_0;
	wire [1:0] w_n1669_0;
	wire [1:0] w_n1671_0;
	wire [1:0] w_n1672_0;
	wire [1:0] w_n1677_0;
	wire [1:0] w_n1682_0;
	wire [1:0] w_n1684_0;
	wire [1:0] w_n1687_0;
	wire [1:0] w_n1689_0;
	wire [1:0] w_n1692_0;
	wire [1:0] w_n1694_0;
	wire [1:0] w_n1697_0;
	wire [1:0] w_n1699_0;
	wire [1:0] w_n1702_0;
	wire [1:0] w_n1703_0;
	wire [1:0] w_n1704_0;
	wire [1:0] w_n1707_0;
	wire [1:0] w_n1709_0;
	wire [1:0] w_n1710_0;
	wire [1:0] w_n1711_0;
	wire [1:0] w_n1712_0;
	wire [1:0] w_n1713_0;
	wire [1:0] w_n1714_0;
	wire [1:0] w_n1715_0;
	wire [1:0] w_n1716_0;
	wire [1:0] w_n1717_0;
	wire [1:0] w_n1719_0;
	wire [1:0] w_n1720_0;
	wire [1:0] w_n1725_0;
	wire [1:0] w_n1728_0;
	wire [1:0] w_n1730_0;
	wire [1:0] w_n1733_0;
	wire [1:0] w_n1735_0;
	wire [1:0] w_n1738_0;
	wire [1:0] w_n1740_0;
	wire [1:0] w_n1743_0;
	wire [1:0] w_n1744_0;
	wire [1:0] w_n1745_0;
	wire [1:0] w_n1748_0;
	wire [1:0] w_n1750_0;
	wire [1:0] w_n1751_0;
	wire [1:0] w_n1752_0;
	wire [1:0] w_n1753_0;
	wire [1:0] w_n1754_0;
	wire [1:0] w_n1755_0;
	wire [1:0] w_n1756_0;
	wire [1:0] w_n1757_0;
	wire [1:0] w_n1758_0;
	wire [1:0] w_n1765_0;
	wire [1:0] w_n1768_0;
	wire [1:0] w_n1770_0;
	wire [1:0] w_n1773_0;
	wire [1:0] w_n1775_0;
	wire [1:0] w_n1778_0;
	wire [1:0] w_n1779_0;
	wire [1:0] w_n1780_0;
	wire [1:0] w_n1783_0;
	wire [1:0] w_n1785_0;
	wire [1:0] w_n1786_0;
	wire [1:0] w_n1787_0;
	wire [1:0] w_n1788_0;
	wire [1:0] w_n1789_0;
	wire [1:0] w_n1790_0;
	wire [1:0] w_n1791_0;
	wire [1:0] w_n1798_0;
	wire [1:0] w_n1801_0;
	wire [1:0] w_n1803_0;
	wire [1:0] w_n1806_0;
	wire [1:0] w_n1807_0;
	wire [1:0] w_n1808_0;
	wire [1:0] w_n1811_0;
	wire [1:0] w_n1813_0;
	wire [1:0] w_n1814_0;
	wire [1:0] w_n1815_0;
	wire [1:0] w_n1816_0;
	wire [1:0] w_n1817_0;
	wire [1:0] w_n1824_0;
	wire [1:0] w_n1827_0;
	wire [1:0] w_n1828_0;
	wire [1:0] w_n1829_0;
	wire [1:0] w_n1832_0;
	wire [1:0] w_n1834_0;
	wire [1:0] w_n1835_0;
	wire [1:0] w_n1836_0;
	wire [1:0] w_n1838_0;
	wire [1:0] w_n1841_0;
	wire [1:0] w_n1848_0;
	wire [1:0] w_n1849_0;
	wire w_dff_B_ORLY9DPs0_1;
	wire w_dff_B_oZHNDDvI5_1;
	wire w_dff_B_Ij8bIAet5_1;
	wire w_dff_B_LNzalzae9_1;
	wire w_dff_B_G2992b235_1;
	wire w_dff_B_Y9xjsZpf4_1;
	wire w_dff_B_cB49q0lG3_1;
	wire w_dff_B_w7BFs5Bb5_1;
	wire w_dff_B_gK2wT7JT1_1;
	wire w_dff_B_eri50NwL8_1;
	wire w_dff_B_sHtfu03p8_1;
	wire w_dff_B_YgdLPBYN7_1;
	wire w_dff_B_7odUktbF4_1;
	wire w_dff_B_AIe7hqhN6_1;
	wire w_dff_B_LtMhjqtt0_1;
	wire w_dff_B_E8jnQa4e2_1;
	wire w_dff_B_k0vSFOZe6_1;
	wire w_dff_B_KTFb8unQ6_1;
	wire w_dff_B_JaqLzDzK5_1;
	wire w_dff_B_UaZUS7uq1_1;
	wire w_dff_B_Gw3gHxAU9_1;
	wire w_dff_B_M40SSfNW0_1;
	wire w_dff_B_k9xHOgEo2_1;
	wire w_dff_B_EBqLY7Wb5_1;
	wire w_dff_B_r2MimJxL5_1;
	wire w_dff_B_IuaNMIbD0_1;
	wire w_dff_B_IX9gG3S53_1;
	wire w_dff_B_LRtb1ykq6_1;
	wire w_dff_B_JDdX9bxa1_1;
	wire w_dff_B_g2lSI0ru0_1;
	wire w_dff_B_QBhLXg9E7_1;
	wire w_dff_B_6ndOoDWP9_1;
	wire w_dff_B_xCeUiCs86_1;
	wire w_dff_B_oAZrojAF4_1;
	wire w_dff_B_Blu890lS8_1;
	wire w_dff_B_XmDg2Ir85_1;
	wire w_dff_B_sWBqXna13_1;
	wire w_dff_B_eH6mOT2k8_1;
	wire w_dff_B_h6aemqzt4_1;
	wire w_dff_B_zCAitGh83_1;
	wire w_dff_B_yFASLsDr1_1;
	wire w_dff_B_IJSxLSEe1_1;
	wire w_dff_B_PFVS4DSZ5_1;
	wire w_dff_B_n6Xnw4qU0_1;
	wire w_dff_B_0AmiNKMU8_1;
	wire w_dff_B_dopvKpGm6_1;
	wire w_dff_B_rkGExKL76_1;
	wire w_dff_B_vaHARmQP2_1;
	wire w_dff_B_EOhZpgfC5_1;
	wire w_dff_B_1N97qTn32_1;
	wire w_dff_B_tADF5loM5_1;
	wire w_dff_B_oz165xF91_1;
	wire w_dff_B_7xNgGFpp8_1;
	wire w_dff_B_tRx9jQr35_1;
	wire w_dff_B_Ryqjbisa9_1;
	wire w_dff_B_Y3zQrAZz4_1;
	wire w_dff_B_FqB3WI4q8_1;
	wire w_dff_B_to8w4a7x0_1;
	wire w_dff_B_OU0FYghf6_1;
	wire w_dff_B_H5DkQQS58_1;
	wire w_dff_B_0lzxZQvI1_1;
	wire w_dff_B_sGY503si0_1;
	wire w_dff_B_N40UKXNQ2_1;
	wire w_dff_B_hNRrtrSy6_1;
	wire w_dff_B_kCq1Pjjp4_1;
	wire w_dff_B_5hSiQmj88_1;
	wire w_dff_B_53B8NZmX8_1;
	wire w_dff_B_sVGJtqzn0_1;
	wire w_dff_B_R1c7Z2Ac4_1;
	wire w_dff_B_Rstyn61Z1_1;
	wire w_dff_B_VB1NPt8j4_1;
	wire w_dff_B_ZXGd2pai9_1;
	wire w_dff_B_HpRRLtSh1_1;
	wire w_dff_B_BP6dCCub8_1;
	wire w_dff_B_7EYqV7Xu1_1;
	wire w_dff_B_W4LGGPQG0_1;
	wire w_dff_B_9mt1mbrt9_1;
	wire w_dff_B_MeN2bBFT2_1;
	wire w_dff_B_MNcptmay2_1;
	wire w_dff_B_80TRIpfk9_1;
	wire w_dff_B_YMAcT9ym8_1;
	wire w_dff_B_dnK0GQsU2_1;
	wire w_dff_B_Tpuf8Jvi6_1;
	wire w_dff_B_piRrKy2c2_1;
	wire w_dff_B_r4gZneIh8_1;
	wire w_dff_B_ZDLBo6Uh5_1;
	wire w_dff_B_WzugrBuw6_1;
	wire w_dff_B_vQoBen6M1_1;
	wire w_dff_B_ZqgtYdFw3_1;
	wire w_dff_B_Cq3OTBLI9_1;
	wire w_dff_B_By0i8jzb1_1;
	wire w_dff_B_sWvwVGJZ8_1;
	wire w_dff_B_VoQ6TS7b0_1;
	wire w_dff_B_Wle8A4Yf0_1;
	wire w_dff_B_UQQW8iTz5_1;
	wire w_dff_B_itdCWixZ0_1;
	wire w_dff_B_V5JRKZ0E7_1;
	wire w_dff_B_nuTxSf3V6_1;
	wire w_dff_B_NsCMPFEu6_1;
	wire w_dff_B_VTRLNAiW9_1;
	wire w_dff_B_MKOKdvzz0_1;
	wire w_dff_B_rLdClAAR1_1;
	wire w_dff_B_tjssuTd70_1;
	wire w_dff_B_OLX31m4k8_1;
	wire w_dff_B_aIeLOVwR2_1;
	wire w_dff_B_uC8AU9eC6_1;
	wire w_dff_B_IQ226zB29_1;
	wire w_dff_B_G9jovtSI4_1;
	wire w_dff_B_mmDSTvj04_1;
	wire w_dff_B_mDnqxGGm3_1;
	wire w_dff_B_BPQLcRlU0_1;
	wire w_dff_B_aiGt8Dic1_1;
	wire w_dff_B_s52Nu9LV3_1;
	wire w_dff_B_bSVOMIX40_1;
	wire w_dff_B_BJLX2naj7_1;
	wire w_dff_B_vcPR8CNy8_1;
	wire w_dff_B_EdoSg5X52_1;
	wire w_dff_B_4gsK11Xq9_1;
	wire w_dff_B_RiXaZqSO7_1;
	wire w_dff_B_YEdKv2G26_1;
	wire w_dff_B_MqDQFoRb5_1;
	wire w_dff_B_XAk9Ie3e6_1;
	wire w_dff_B_ZcCR1UC79_1;
	wire w_dff_B_RYAcUgtn8_1;
	wire w_dff_B_6U4SpEKA3_1;
	wire w_dff_B_1W6La1mW7_1;
	wire w_dff_B_U3NVz7Gm3_1;
	wire w_dff_B_uqQY5foB5_1;
	wire w_dff_B_f8Wxk0BQ4_1;
	wire w_dff_B_FdNtK8LV3_1;
	wire w_dff_B_nk4NLpLZ7_1;
	wire w_dff_B_uwf0iG056_1;
	wire w_dff_B_NfkAaFSp9_1;
	wire w_dff_B_FzXvi16b5_1;
	wire w_dff_B_ssy4zHjc9_1;
	wire w_dff_B_M4pUayoG1_1;
	wire w_dff_B_Cr8Iu6sw6_1;
	wire w_dff_B_y9oGrr659_1;
	wire w_dff_B_leFj1xjK8_1;
	wire w_dff_B_1SPpOoKH7_1;
	wire w_dff_B_yxOTRkff3_1;
	wire w_dff_B_NXBs2v549_1;
	wire w_dff_B_QxvYgTXT7_1;
	wire w_dff_B_7nDGrMEn4_1;
	wire w_dff_B_wgsWXVkt3_1;
	wire w_dff_B_Ng7TGNCt8_1;
	wire w_dff_B_eBBkXGyg4_1;
	wire w_dff_B_5oeXDePC1_1;
	wire w_dff_B_WNVXoER12_1;
	wire w_dff_B_Uh2Azmw13_1;
	wire w_dff_B_LB5rLVW66_1;
	wire w_dff_B_Q251MPaq6_1;
	wire w_dff_B_FxOmnJYt7_1;
	wire w_dff_B_b4tasGne0_1;
	wire w_dff_B_RQpEWAFG6_1;
	wire w_dff_B_udbH2LjQ4_1;
	wire w_dff_B_e6tXLClc7_1;
	wire w_dff_B_k5wDjoX28_1;
	wire w_dff_B_7n3OBNNV4_1;
	wire w_dff_B_AlWaHE5r6_1;
	wire w_dff_B_MuIFzA4v1_1;
	wire w_dff_B_xpKQQ4mf8_1;
	wire w_dff_B_TSMfxi0V4_1;
	wire w_dff_B_3Tyoumh72_1;
	wire w_dff_B_l8S7gwAd0_1;
	wire w_dff_B_teFzx1jm2_1;
	wire w_dff_B_Mb96YJlx9_1;
	wire w_dff_B_8r7Z6t1f5_1;
	wire w_dff_B_7Cm8J7323_1;
	wire w_dff_B_YO0GtC4U2_1;
	wire w_dff_B_L1iFFo4V1_1;
	wire w_dff_B_DPvSa2gd6_1;
	wire w_dff_B_NsC6prcU0_1;
	wire w_dff_B_7ROqNocH2_1;
	wire w_dff_B_QHokTbzR1_1;
	wire w_dff_B_g6Pg8PGz3_1;
	wire w_dff_B_o02MqCH97_1;
	wire w_dff_B_rzPZ16kv6_1;
	wire w_dff_B_MKEs9oF78_1;
	wire w_dff_B_NeRT2TyM7_1;
	wire w_dff_B_vjBECOxd6_1;
	wire w_dff_B_1i8tbPKA3_1;
	wire w_dff_B_843t3xRY4_1;
	wire w_dff_B_bdqLC7vo9_1;
	wire w_dff_B_TNcI5eRw5_1;
	wire w_dff_B_LwTHwz5h1_1;
	wire w_dff_B_ogKjg4TT7_1;
	wire w_dff_B_1tnGRLsd5_1;
	wire w_dff_B_VX77IbmL3_1;
	wire w_dff_B_OYPlSZWi4_1;
	wire w_dff_B_ZyFnTC5A9_1;
	wire w_dff_B_Bq9AfCGp8_1;
	wire w_dff_B_FBymBW7n1_1;
	wire w_dff_B_MBqbtgjv8_1;
	wire w_dff_B_atvdlYe82_1;
	wire w_dff_B_wuJiLk3f0_1;
	wire w_dff_B_f8wiba432_1;
	wire w_dff_B_iarYdNOs8_1;
	wire w_dff_B_SUNnvvs75_1;
	wire w_dff_B_p8pivOpx2_1;
	wire w_dff_B_WrnvBMAh0_1;
	wire w_dff_B_OMVFAJ2a6_1;
	wire w_dff_B_YElUZzDf9_1;
	wire w_dff_B_U1mmLwCZ0_1;
	wire w_dff_B_4oTRfwQr8_1;
	wire w_dff_B_dKRgVAHZ8_1;
	wire w_dff_B_UrxQXydp3_1;
	wire w_dff_B_5wtEYjLL2_1;
	wire w_dff_B_4lb9XoRh5_1;
	wire w_dff_B_I9nJ9Bc26_1;
	wire w_dff_B_ba7yHDor7_1;
	wire w_dff_B_1v9PejCt4_1;
	wire w_dff_B_E6K7aPBy9_1;
	wire w_dff_B_kjU0WIxU8_1;
	wire w_dff_B_m5VZ61L67_1;
	wire w_dff_B_hoJsCj2k7_1;
	wire w_dff_B_YNt5KqTj9_1;
	wire w_dff_B_KrtjcLqM4_1;
	wire w_dff_B_cjyca7w44_1;
	wire w_dff_B_LMGnYrWV7_1;
	wire w_dff_B_D0n8gG373_1;
	wire w_dff_B_xustH9JN0_1;
	wire w_dff_B_AdciMGAg0_1;
	wire w_dff_B_YgVZMix71_1;
	wire w_dff_B_2x8z9CsQ3_1;
	wire w_dff_B_3R5MpDEX5_1;
	wire w_dff_B_MAphkkXz6_1;
	wire w_dff_B_tBGD9mXy0_1;
	wire w_dff_B_nxywcEQT7_1;
	wire w_dff_B_43c16sot3_1;
	wire w_dff_B_YOI6Kdlw6_1;
	wire w_dff_B_4vog6DFp5_1;
	wire w_dff_B_HLRyeS8Z6_1;
	wire w_dff_B_YPLgVBAv6_1;
	wire w_dff_B_EnAH4Js65_1;
	wire w_dff_B_xvFx4mJ55_1;
	wire w_dff_B_TTSwfGcV1_1;
	wire w_dff_B_5a35RJUv5_1;
	wire w_dff_B_IkHbgszW1_1;
	wire w_dff_B_OHLiR9ce0_1;
	wire w_dff_B_aQJSDXwv1_1;
	wire w_dff_B_KEclRy8v4_1;
	wire w_dff_B_J6hTIKWU6_1;
	wire w_dff_B_1xGOBdgR8_1;
	wire w_dff_B_4I22MR9j5_1;
	wire w_dff_B_l9Znp2i90_1;
	wire w_dff_B_fX6XFwfv2_1;
	wire w_dff_B_bhERwpZM9_1;
	wire w_dff_B_vounQEKF0_1;
	wire w_dff_B_iEe7ZKqG0_1;
	wire w_dff_B_E0LBWgmp0_1;
	wire w_dff_B_fckmYLXb9_1;
	wire w_dff_B_ojD4jv0Q0_1;
	wire w_dff_B_0lII4XEZ5_1;
	wire w_dff_B_1yEjaGtF8_1;
	wire w_dff_B_16CiTP473_1;
	wire w_dff_B_GPpO06U95_1;
	wire w_dff_B_ywCLCs4H4_1;
	wire w_dff_B_cd6ipKFb5_1;
	wire w_dff_B_zxKrJ2Hg1_1;
	wire w_dff_B_4yU7EuX57_1;
	wire w_dff_B_TP0usAbO3_1;
	wire w_dff_B_sAXTRqGj2_1;
	wire w_dff_B_5ZVIeCy01_1;
	wire w_dff_B_gKeN94ss9_1;
	wire w_dff_B_mYQ91xFU0_1;
	wire w_dff_B_dqyaHDPz6_1;
	wire w_dff_B_83rQTowt2_1;
	wire w_dff_B_gGVYeCIU3_1;
	wire w_dff_B_qegBv0gk7_1;
	wire w_dff_B_ljCYe4Mi5_1;
	wire w_dff_B_eERNXww16_1;
	wire w_dff_B_1j0PqywI6_1;
	wire w_dff_B_Fp4hZQj24_1;
	wire w_dff_B_Bzd4Gd4G7_1;
	wire w_dff_B_IOkKtf9i2_1;
	wire w_dff_B_I0WggfyD7_1;
	wire w_dff_B_fonbVM4p5_1;
	wire w_dff_B_vaq0t36y3_1;
	wire w_dff_B_gorOyYwL1_1;
	wire w_dff_B_9aONanXf9_1;
	wire w_dff_B_VfrXnsV62_1;
	wire w_dff_B_Qvl9bDzk3_1;
	wire w_dff_B_A2DRuLiV4_1;
	wire w_dff_B_pjxF3ZmG0_1;
	wire w_dff_B_pCPX82E15_1;
	wire w_dff_B_P2cfAhMG6_1;
	wire w_dff_B_EcYzZ6w71_1;
	wire w_dff_B_wIr2XIFU7_1;
	wire w_dff_B_furpVV9k1_1;
	wire w_dff_B_QvHf1xwY0_1;
	wire w_dff_B_o4u3vI5k6_1;
	wire w_dff_B_kHPkxqTA9_1;
	wire w_dff_B_obd657vg8_1;
	wire w_dff_B_33mIoTbk8_1;
	wire w_dff_B_yxBmnghK9_1;
	wire w_dff_B_eXX13Pqf2_1;
	wire w_dff_B_0ueVHSbU3_1;
	wire w_dff_B_k8P4wljZ5_1;
	wire w_dff_B_xLEamzwr9_1;
	wire w_dff_B_zURI3Hdu6_1;
	wire w_dff_B_kYeKGal02_1;
	wire w_dff_B_wnEDff3J9_1;
	wire w_dff_B_vU0e0Ijl7_1;
	wire w_dff_B_TjK5C9pn3_1;
	wire w_dff_B_leCVotMu8_1;
	wire w_dff_B_Ocyxqbgr9_1;
	wire w_dff_B_3u7UaqNw8_1;
	wire w_dff_B_2SKH4sBb5_1;
	wire w_dff_B_xPcaFZLU2_1;
	wire w_dff_B_8S3jPgSq7_1;
	wire w_dff_B_vGd5woqt0_1;
	wire w_dff_B_ZTvQ8cOR8_1;
	wire w_dff_B_PirkwQWd4_1;
	wire w_dff_B_jpzYNZOM2_1;
	wire w_dff_B_Lg15YytX8_1;
	wire w_dff_B_C37td1dx7_1;
	wire w_dff_B_L6WtZiIo4_1;
	wire w_dff_B_n3S53RUV4_1;
	wire w_dff_B_hupLYL7c3_1;
	wire w_dff_B_gmBAj38L4_1;
	wire w_dff_B_qLJbvFUF3_1;
	wire w_dff_B_lMpFMA492_1;
	wire w_dff_B_DMuZ9GNp9_1;
	wire w_dff_B_eN08a2vV8_1;
	wire w_dff_B_TZVngQF69_1;
	wire w_dff_B_5aFT5H7H8_1;
	wire w_dff_B_AH6MrSp94_1;
	wire w_dff_B_fxHsrPUf6_1;
	wire w_dff_B_vYOXfILh7_1;
	wire w_dff_B_fMoeLlFX7_0;
	wire w_dff_B_sbFeo1EI5_1;
	wire w_dff_B_2INyUXAH4_1;
	wire w_dff_B_zTW8EAQk9_1;
	wire w_dff_B_kcolGlWG7_1;
	wire w_dff_B_bmKLUEvh2_1;
	wire w_dff_B_RwqUbpFi6_1;
	wire w_dff_B_ReuhXnQ20_1;
	wire w_dff_B_pAVLRkq43_1;
	wire w_dff_B_pihkHoxr6_1;
	wire w_dff_B_6xtnLTau1_1;
	wire w_dff_B_bna7xfMG2_1;
	wire w_dff_B_qeId6v1Q8_1;
	wire w_dff_B_tEIzL6Si8_1;
	wire w_dff_B_hQicRh9g9_0;
	wire w_dff_B_Zsh8d9J27_0;
	wire w_dff_B_EJ1uPLOd7_0;
	wire w_dff_B_49lDF8be5_0;
	wire w_dff_B_oubJSXAn0_0;
	wire w_dff_B_AgpVtZNU5_0;
	wire w_dff_B_aqxE7IaL6_0;
	wire w_dff_B_z2OGlrf04_0;
	wire w_dff_B_gMnJwXhg9_0;
	wire w_dff_B_MHn6vCaL1_0;
	wire w_dff_B_lO57ET7m6_0;
	wire w_dff_A_m0JjNuvI8_0;
	wire w_dff_A_XyLHhIko8_0;
	wire w_dff_A_YZyxKGH84_0;
	wire w_dff_A_zNE32iKI2_0;
	wire w_dff_A_J6oD1eTw0_0;
	wire w_dff_A_RzBZ9N197_0;
	wire w_dff_A_PbKFL8IP9_0;
	wire w_dff_A_w5ljE4UP8_0;
	wire w_dff_A_ldpsVJv72_0;
	wire w_dff_A_BIR0T2Er1_0;
	wire w_dff_A_UOZBiI5q7_0;
	wire w_dff_A_AfYw5laX3_0;
	wire w_dff_B_tWoZIzdD1_1;
	wire w_dff_B_l8E1hQ3o8_1;
	wire w_dff_B_iz9aTgB08_2;
	wire w_dff_B_bV3ZWcCp4_2;
	wire w_dff_B_qTkMv25N4_2;
	wire w_dff_B_qYKJNjHM8_2;
	wire w_dff_B_ZE0PLiXw4_2;
	wire w_dff_B_e7JmlJml1_2;
	wire w_dff_B_pSibLW3N1_2;
	wire w_dff_B_Xb5OxJb10_2;
	wire w_dff_B_2fv4WZuu7_2;
	wire w_dff_B_aU7SC2Mt6_2;
	wire w_dff_B_AMl8UHIt8_2;
	wire w_dff_B_zqxapdLY1_2;
	wire w_dff_B_r1kE9BxB6_2;
	wire w_dff_B_QatLuJBO0_2;
	wire w_dff_B_xgMpC9re1_2;
	wire w_dff_B_4XrfGHGV8_2;
	wire w_dff_B_tBJTXV7x1_2;
	wire w_dff_B_MR6tEHgC4_2;
	wire w_dff_B_e34WTH2O3_2;
	wire w_dff_B_hUnFkNs61_2;
	wire w_dff_B_RnZXvcQH5_2;
	wire w_dff_B_7ADFwLpP0_2;
	wire w_dff_B_wXScGgMg6_2;
	wire w_dff_B_A3sTDcJI9_2;
	wire w_dff_B_AUuzRjLB8_2;
	wire w_dff_B_3LPsbA4d6_2;
	wire w_dff_B_m28lmXxm5_2;
	wire w_dff_B_vGvo1yPu8_2;
	wire w_dff_B_orcXzQlX1_2;
	wire w_dff_B_TW4Lygyl1_2;
	wire w_dff_B_NehRVWgf9_2;
	wire w_dff_B_k6lnXCH26_2;
	wire w_dff_B_mtTvTe6Y9_2;
	wire w_dff_B_1Qyk3WNZ6_2;
	wire w_dff_B_CtmDnbP80_2;
	wire w_dff_B_3t6dei1P1_2;
	wire w_dff_B_7uNCo4D26_2;
	wire w_dff_B_T8ejGtNS7_2;
	wire w_dff_B_Yak9Udtk2_2;
	wire w_dff_B_R0LIlpBN7_2;
	wire w_dff_B_5SzAzHYS9_2;
	wire w_dff_B_ICHowvGj6_2;
	wire w_dff_B_J7UtQFDH1_2;
	wire w_dff_B_D6Ik5QjN1_2;
	wire w_dff_B_PMAbDxLz8_2;
	wire w_dff_B_ImRoXffv4_2;
	wire w_dff_B_Pftahw966_2;
	wire w_dff_B_lG50ej0b4_2;
	wire w_dff_B_r4AF2vQW2_2;
	wire w_dff_B_uBLBvLJo3_2;
	wire w_dff_B_fOJhEY0Y2_2;
	wire w_dff_B_ktcPXAgr7_2;
	wire w_dff_B_4OKefqFS1_2;
	wire w_dff_B_mF1Ktk8h2_2;
	wire w_dff_B_FhwPWVkg5_2;
	wire w_dff_B_ZRuRRZd25_2;
	wire w_dff_B_IgwhY4ht2_2;
	wire w_dff_B_rgzkUHGt0_2;
	wire w_dff_B_jAPfrKB49_2;
	wire w_dff_B_g4xoyXVp5_2;
	wire w_dff_B_YAyryhwi7_1;
	wire w_dff_B_n8wgVtZu5_1;
	wire w_dff_B_CEZXvmhg5_1;
	wire w_dff_B_iE86Ry8q4_1;
	wire w_dff_B_5Gr5F1uv0_1;
	wire w_dff_B_AjkQlkJc1_1;
	wire w_dff_B_lVVVOTHN7_1;
	wire w_dff_B_YjTJqmDs0_1;
	wire w_dff_B_OztWx61B7_1;
	wire w_dff_B_GCPIvll60_1;
	wire w_dff_B_wJhP7oj49_1;
	wire w_dff_B_EMOiCLTU2_0;
	wire w_dff_B_VZTT7cji8_0;
	wire w_dff_B_DC8U9q976_0;
	wire w_dff_B_3YqqsRiB0_0;
	wire w_dff_B_t7nv8bQi1_0;
	wire w_dff_B_I0yUCq319_0;
	wire w_dff_B_7Uv01WtP1_0;
	wire w_dff_B_LzStQ3BC8_0;
	wire w_dff_B_WmBNDTAf5_0;
	wire w_dff_B_4MdSaJGN5_0;
	wire w_dff_A_fmIwcrek3_1;
	wire w_dff_A_IdGKqR6F6_1;
	wire w_dff_A_xkn4FbBm7_1;
	wire w_dff_A_sJ43ChCR0_1;
	wire w_dff_A_Jnu1htZZ2_1;
	wire w_dff_A_2yfFXLks2_1;
	wire w_dff_A_ewtxhN3X2_1;
	wire w_dff_A_FQo0tz0n9_1;
	wire w_dff_A_TaYisTDI2_1;
	wire w_dff_A_JC7YBa092_1;
	wire w_dff_A_TxFnIYqv4_1;
	wire w_dff_B_q6Qq8Sg23_1;
	wire w_dff_B_Ay8glTj51_1;
	wire w_dff_B_b8Ma6md70_1;
	wire w_dff_B_aQi1gvLr0_1;
	wire w_dff_B_Ldv37RNC9_1;
	wire w_dff_B_4Nq2UBo37_1;
	wire w_dff_B_7vTiqso71_1;
	wire w_dff_B_gnm77Bmi3_1;
	wire w_dff_B_fO3h4D8N1_1;
	wire w_dff_B_OClDH2tm0_1;
	wire w_dff_B_V4tVImYF3_1;
	wire w_dff_B_m15yRGzY6_0;
	wire w_dff_B_UBlVmbjq0_0;
	wire w_dff_B_uNkVxzEa5_0;
	wire w_dff_B_KJL4lO9v3_0;
	wire w_dff_B_aPw0MuTd1_0;
	wire w_dff_B_rcNnLJ2S1_0;
	wire w_dff_B_j4djZjDh0_0;
	wire w_dff_B_82Yeytqs9_0;
	wire w_dff_B_qkz65yQF3_0;
	wire w_dff_B_k03xV37X7_0;
	wire w_dff_A_Yy2ZexX11_1;
	wire w_dff_A_6sBrAL3t7_1;
	wire w_dff_A_9BRfZH5s0_1;
	wire w_dff_A_L9cWyI3p3_1;
	wire w_dff_A_nIyoYqLH8_1;
	wire w_dff_A_dQdlcR7G4_1;
	wire w_dff_A_etzBS0ph8_1;
	wire w_dff_A_b1nMr4uH3_1;
	wire w_dff_A_LTxjtvaL4_1;
	wire w_dff_A_PfRSPYNF2_1;
	wire w_dff_A_axlC0KEc6_1;
	wire w_dff_B_kVPEUSYw5_1;
	wire w_dff_B_5l0iSaGZ3_1;
	wire w_dff_B_IIk8IVHM1_1;
	wire w_dff_B_OrVwB2EW5_1;
	wire w_dff_B_jC1WHUIe7_1;
	wire w_dff_B_JynPFKln8_1;
	wire w_dff_B_KvA4F5B44_1;
	wire w_dff_B_aYfYaXIp1_1;
	wire w_dff_B_1bzdDDi43_1;
	wire w_dff_B_IuZmrOTp9_1;
	wire w_dff_B_2lTowDer4_1;
	wire w_dff_B_C8qvizap8_0;
	wire w_dff_B_lBnjesKo5_0;
	wire w_dff_B_jz1RhArz6_0;
	wire w_dff_B_CuB6WOtN4_0;
	wire w_dff_B_zjvUSenK3_0;
	wire w_dff_B_23I54xxa7_0;
	wire w_dff_B_LPvYyFpm3_0;
	wire w_dff_B_C3nCA6dU3_0;
	wire w_dff_B_Y22ZQXVl8_0;
	wire w_dff_B_uo9daJrs0_0;
	wire w_dff_A_1wWc61pi3_1;
	wire w_dff_A_yQ3s8HxE3_1;
	wire w_dff_A_bZZlQ63Z6_1;
	wire w_dff_A_sJz3lPCI2_1;
	wire w_dff_A_AeVnl6g52_1;
	wire w_dff_A_ujEWTp711_1;
	wire w_dff_A_CjsMYCwH0_1;
	wire w_dff_A_3I90hbjW0_1;
	wire w_dff_A_P6IelWAb2_1;
	wire w_dff_A_6NepZbbQ7_1;
	wire w_dff_A_DbyttkQU3_1;
	wire w_dff_B_5IpxAz8Z3_1;
	wire w_dff_B_vmnqg6ss9_1;
	wire w_dff_B_a0HmcnQt4_1;
	wire w_dff_B_GDNd8PaH0_1;
	wire w_dff_B_Dx47z0606_1;
	wire w_dff_B_7y7VD2tk1_1;
	wire w_dff_B_RhgaHpNV8_1;
	wire w_dff_B_2eVIsDYU4_1;
	wire w_dff_B_LpGSaLql7_1;
	wire w_dff_B_B6zPzUqH3_1;
	wire w_dff_B_wn5H5gc59_1;
	wire w_dff_B_SNWo6Qzh0_0;
	wire w_dff_B_JCohFOdw7_0;
	wire w_dff_B_dBnURjkZ9_0;
	wire w_dff_B_KKfS702Q7_0;
	wire w_dff_B_SLl5u2BT3_0;
	wire w_dff_B_HcmqYFwf9_0;
	wire w_dff_B_6ZEM32JD3_0;
	wire w_dff_B_2mWIb39J0_0;
	wire w_dff_B_nnnlgVky2_0;
	wire w_dff_B_pS6Cq4dI7_0;
	wire w_dff_A_BL7JtSMX2_1;
	wire w_dff_A_gVAvQkw08_1;
	wire w_dff_A_OA5pJVT69_1;
	wire w_dff_A_19h8PTCo1_1;
	wire w_dff_A_L7S2zJkL2_1;
	wire w_dff_A_0knXNdyO8_1;
	wire w_dff_A_XLhx0YIo9_1;
	wire w_dff_A_DjUE5ZZc0_1;
	wire w_dff_A_8xz9VRPK9_1;
	wire w_dff_A_mHSJJKXo5_1;
	wire w_dff_A_RlkqRC6Q9_1;
	wire w_dff_B_v6IhuskW6_1;
	wire w_dff_B_63Mcjvni8_1;
	wire w_dff_B_wWKuo2wb4_1;
	wire w_dff_B_Bdhejcms1_1;
	wire w_dff_B_E5cBadYg7_1;
	wire w_dff_B_kvA1IVVx7_1;
	wire w_dff_B_KTiaSrYS3_1;
	wire w_dff_B_gdbnzCQD1_1;
	wire w_dff_B_YncGPHfT1_1;
	wire w_dff_B_g1SETCA08_1;
	wire w_dff_B_j8qeHvjW3_1;
	wire w_dff_B_NMCqCl6C4_0;
	wire w_dff_B_6NwIBqkQ4_0;
	wire w_dff_B_C65pYUIX2_0;
	wire w_dff_B_VrInQc6Q7_0;
	wire w_dff_B_qAXq7WAD6_0;
	wire w_dff_B_T8MwLudp5_0;
	wire w_dff_B_dDKNL7hr7_0;
	wire w_dff_B_NYILoQxo0_0;
	wire w_dff_B_plAUKf9m5_0;
	wire w_dff_A_JDqsIVPy3_1;
	wire w_dff_A_9Rl5Nb2Z0_1;
	wire w_dff_A_3yhR6Yn71_1;
	wire w_dff_A_FZKJHNdz8_1;
	wire w_dff_A_pe6LVOie1_1;
	wire w_dff_A_PRTjnTu04_1;
	wire w_dff_A_mwh0BfB78_1;
	wire w_dff_A_ho26mdp31_1;
	wire w_dff_A_G9YDQs7A9_1;
	wire w_dff_A_mHhCd8B79_1;
	wire w_dff_B_wn7ZCnbN9_1;
	wire w_dff_B_dn4JiUK64_1;
	wire w_dff_B_VUJCs6ZS0_1;
	wire w_dff_B_OrD85vZy6_1;
	wire w_dff_B_zEJMwPul2_1;
	wire w_dff_B_OWdu6gAX7_1;
	wire w_dff_B_w5AIDrQX9_1;
	wire w_dff_B_4mhNrqrI1_1;
	wire w_dff_B_OK4ySXev2_1;
	wire w_dff_B_J3ei1HvP0_1;
	wire w_dff_B_zqYyVafT0_0;
	wire w_dff_B_yFBrxJni0_0;
	wire w_dff_B_UQIfRW0B4_0;
	wire w_dff_B_73QqV5xQ9_0;
	wire w_dff_B_U7IAGtya2_0;
	wire w_dff_B_T6fUOHGE2_0;
	wire w_dff_B_Qh64Slzd2_0;
	wire w_dff_B_hwj8yCsY3_0;
	wire w_dff_A_PEMtf3vg5_1;
	wire w_dff_A_Cdu3USMO5_1;
	wire w_dff_A_zhX2MfbU8_1;
	wire w_dff_A_LFvGuECz9_1;
	wire w_dff_A_niCj6BqO6_1;
	wire w_dff_A_jxK1qrBp5_1;
	wire w_dff_A_eQCJCu5d0_1;
	wire w_dff_A_uuOsS5Nl6_1;
	wire w_dff_A_alqW54nR6_1;
	wire w_dff_B_hDIJRorC0_1;
	wire w_dff_B_XYhI3q5R6_1;
	wire w_dff_B_IT6zoV182_1;
	wire w_dff_B_91PgArA15_1;
	wire w_dff_B_hREdb58u6_1;
	wire w_dff_B_MWc4OmHJ5_1;
	wire w_dff_B_rK8WkAaj8_1;
	wire w_dff_B_BN5B8V2h3_1;
	wire w_dff_B_QPdpzU6K2_1;
	wire w_dff_B_LL8oMdvo3_1;
	wire w_dff_B_IYlB5aSd1_0;
	wire w_dff_B_ZTaSJ6TW1_0;
	wire w_dff_B_jdmB6ANR4_0;
	wire w_dff_B_3PQFhNu23_0;
	wire w_dff_B_Y0oZyQIu9_0;
	wire w_dff_B_N3LBxeXa8_0;
	wire w_dff_B_YGbr3H580_0;
	wire w_dff_B_UtgNrEWs9_0;
	wire w_dff_A_vqWjPbkR0_1;
	wire w_dff_A_fQ4eruGN5_1;
	wire w_dff_A_5M2X4v0J2_1;
	wire w_dff_A_2OamhUUX4_1;
	wire w_dff_A_iwFPN9Lb6_1;
	wire w_dff_A_OHdBHNXF9_1;
	wire w_dff_A_l60AQmtu6_1;
	wire w_dff_A_kro1kpmS6_1;
	wire w_dff_A_1K1g5fbW6_1;
	wire w_dff_B_qThZXVAS5_1;
	wire w_dff_B_4KsNT68r4_1;
	wire w_dff_B_m0321h2C0_1;
	wire w_dff_B_AtHV9SqQ6_1;
	wire w_dff_B_1taZFBdh8_1;
	wire w_dff_B_ZuRuUN8X6_1;
	wire w_dff_B_RNNhOt3S1_1;
	wire w_dff_B_PaiXs0mt7_1;
	wire w_dff_B_tH6DKS5D0_0;
	wire w_dff_B_wAzPyPXZ1_0;
	wire w_dff_B_453u6ucA1_0;
	wire w_dff_B_KBA9Z8uR9_0;
	wire w_dff_B_eK1Ui84y8_0;
	wire w_dff_B_qqrw33Vf4_0;
	wire w_dff_A_sBMcs55T8_1;
	wire w_dff_A_fyj4QY1o3_1;
	wire w_dff_A_oxyUvhSv3_1;
	wire w_dff_A_aaetnem01_1;
	wire w_dff_A_Bw5tnDwG9_1;
	wire w_dff_A_vFKT07tG1_1;
	wire w_dff_A_0GFTuX1r9_1;
	wire w_dff_B_89zGTgIV5_1;
	wire w_dff_B_tbNkuEda9_1;
	wire w_dff_B_Lf1hSQTd4_1;
	wire w_dff_B_B7Y8Xqzg5_1;
	wire w_dff_B_sipoZOv55_1;
	wire w_dff_B_I6yWBDMP5_1;
	wire w_dff_B_uM7kyvMl1_1;
	wire w_dff_B_BOAjz2Gm4_0;
	wire w_dff_B_NlqWlu6X0_0;
	wire w_dff_B_NBYt3pqa5_0;
	wire w_dff_B_WfTwraRJ8_0;
	wire w_dff_B_fW2lPW9w3_0;
	wire w_dff_A_YyE8LCpd2_1;
	wire w_dff_A_kyqDLJ360_1;
	wire w_dff_A_yVVeluAA9_1;
	wire w_dff_A_BK3FG69W3_1;
	wire w_dff_A_bd6lX0Qc8_1;
	wire w_dff_A_aEBeq1PX8_1;
	wire w_dff_B_7YPz0EEJ5_1;
	wire w_dff_B_vSqMAagr0_1;
	wire w_dff_B_g1EjlE8T9_1;
	wire w_dff_B_UukhTS6B9_1;
	wire w_dff_B_TnCH5q7Z6_1;
	wire w_dff_B_WWr6rpmz9_1;
	wire w_dff_B_fwtVPQSN3_0;
	wire w_dff_B_od5UusqG5_0;
	wire w_dff_B_L58Alc1U3_0;
	wire w_dff_B_RMHEEMGh8_0;
	wire w_dff_A_icapOvkN0_1;
	wire w_dff_A_Dh0iTn9n1_1;
	wire w_dff_A_00RSsezR6_1;
	wire w_dff_A_adH5Mp8P7_1;
	wire w_dff_A_VznJHwpx9_1;
	wire w_dff_B_EaACql833_1;
	wire w_dff_B_CNq2ygGW5_1;
	wire w_dff_B_3s0PRdKJ2_1;
	wire w_dff_A_MOiX7ir23_0;
	wire w_dff_A_K4ToNhLz9_0;
	wire w_dff_B_BFNl21zT8_1;
	wire w_dff_A_8LRjp0fZ3_0;
	wire w_dff_B_YxY9L11J6_1;
	wire w_dff_A_BLchi0CF4_1;
	wire w_dff_B_6NEy3HGz2_2;
	wire w_dff_B_uKVEnDbQ2_1;
	wire w_dff_A_6V7hrwzn6_0;
	wire w_dff_A_fNxtcm6l6_0;
	wire w_dff_A_6F0XgFpA4_0;
	wire w_dff_A_J44bVdcI7_0;
	wire w_dff_A_psvP85Nc8_0;
	wire w_dff_A_svKF7qMX4_0;
	wire w_dff_A_ceoaJjlg4_0;
	wire w_dff_A_uMh3wmh43_0;
	wire w_dff_A_W9TbWtlx1_0;
	wire w_dff_A_56uq5eD56_0;
	wire w_dff_A_pk7oJCgU3_0;
	wire w_dff_A_OWeYt4PU1_0;
	wire w_dff_A_BRlYgQwf5_0;
	wire w_dff_A_lXeA3x2S5_0;
	wire w_dff_A_izlyF6sL0_0;
	wire w_dff_A_8v87OChG1_0;
	wire w_dff_A_Q37cT2OV6_0;
	wire w_dff_A_8lR8qIBP6_0;
	wire w_dff_A_f2ymBBmN9_0;
	wire w_dff_A_uwxDyZH07_0;
	wire w_dff_A_TaJiwgA97_0;
	wire w_dff_A_JsTOEFvp2_0;
	wire w_dff_A_5XoUr31V9_0;
	wire w_dff_A_s2FCC40a3_0;
	wire w_dff_A_rCDjsYt57_0;
	wire w_dff_A_6XcoHjrL7_0;
	wire w_dff_A_plIe5c5R0_0;
	wire w_dff_A_lXIm4D0B8_0;
	wire w_dff_A_cjOmuz7j2_0;
	wire w_dff_A_MQJ1NTqI4_0;
	wire w_dff_A_6pA4xgLf6_0;
	wire w_dff_A_AVj3Kxvt1_0;
	wire w_dff_A_riwt5X847_0;
	wire w_dff_A_hQVe51HY8_0;
	wire w_dff_A_CT7W2dHd3_0;
	wire w_dff_A_lHUiqZYq7_0;
	wire w_dff_A_0DwLaxM29_0;
	wire w_dff_A_cvpYQpNF5_0;
	wire w_dff_A_K5Az5ea85_0;
	wire w_dff_A_9jw0b8U63_0;
	wire w_dff_A_UJ9I5hKy2_0;
	wire w_dff_A_0ZD60s2I6_0;
	wire w_dff_A_6Qm3LNbZ2_0;
	wire w_dff_A_4Cy19Jzl6_0;
	wire w_dff_A_nNe7f8Xx0_1;
	wire w_dff_B_cm5qEtPD6_1;
	wire w_dff_A_hpkQO7MK5_0;
	wire w_dff_A_S0gkK6by2_0;
	wire w_dff_A_wv30d5M87_0;
	wire w_dff_A_l5LiC6On9_0;
	wire w_dff_A_x8gfXW7k9_0;
	wire w_dff_A_sZ1guD3X8_0;
	wire w_dff_A_AMEnIHwt7_0;
	wire w_dff_A_XOlSkgMJ2_0;
	wire w_dff_A_BYrGcG2S3_0;
	wire w_dff_A_QEu5ft5c4_0;
	wire w_dff_A_4dHJ5FnO9_0;
	wire w_dff_A_0qZAWYTK7_0;
	wire w_dff_A_uF596t8g2_0;
	wire w_dff_A_ijqfPpKd9_0;
	wire w_dff_A_Ug3QQrpa5_0;
	wire w_dff_A_ZR61NCGG8_0;
	wire w_dff_A_v4Ozbc4b5_0;
	wire w_dff_A_WwPIPAVl7_0;
	wire w_dff_A_gb66Bs6G0_0;
	wire w_dff_A_uFyblmZr5_0;
	wire w_dff_A_jzHJH7ng6_0;
	wire w_dff_A_kvrYy2i36_0;
	wire w_dff_A_5bfFOKNy9_0;
	wire w_dff_A_YTXbspCj6_0;
	wire w_dff_A_QbgmQ9GR0_0;
	wire w_dff_A_DWtzE9Lg9_0;
	wire w_dff_A_rD2ES1qK5_0;
	wire w_dff_A_M8jWDMan9_0;
	wire w_dff_A_D9l9qJ8J3_0;
	wire w_dff_A_hd2BDvex8_0;
	wire w_dff_A_pQIeJ1yR6_0;
	wire w_dff_A_3nxdof6H0_0;
	wire w_dff_A_j3UuPga36_0;
	wire w_dff_A_jnYUxKz76_0;
	wire w_dff_A_s9qkdFRi6_0;
	wire w_dff_A_0Qx3SRCO8_0;
	wire w_dff_A_uknZAKxN2_0;
	wire w_dff_A_jIWh811E7_0;
	wire w_dff_A_CDbqx1dQ0_0;
	wire w_dff_A_zTPZjg254_0;
	wire w_dff_A_O44AF8rm8_0;
	wire w_dff_A_ve3QpJuC3_1;
	wire w_dff_B_L99dMJIv6_1;
	wire w_dff_B_KKp1gkxY3_1;
	wire w_dff_B_OprdLYLo0_1;
	wire w_dff_B_76Lwyahd0_1;
	wire w_dff_B_bwVhD8xL5_1;
	wire w_dff_B_c9FhlcRE6_1;
	wire w_dff_B_db3vdHwX2_1;
	wire w_dff_B_TzrojeaV2_1;
	wire w_dff_B_OdyuZ8aR4_1;
	wire w_dff_B_OtluU48w3_1;
	wire w_dff_B_1rwJXIys4_1;
	wire w_dff_B_yNTuvNMC9_1;
	wire w_dff_B_O7B3LFZ33_1;
	wire w_dff_B_Dt2BYe0z8_1;
	wire w_dff_B_bph5RScJ6_1;
	wire w_dff_B_srYuAKkj3_1;
	wire w_dff_B_22bIZSn63_1;
	wire w_dff_B_lYRTQzSs5_1;
	wire w_dff_B_hcq8z5Yw5_1;
	wire w_dff_B_5PdSpXBM8_1;
	wire w_dff_B_o3oBp1mo1_1;
	wire w_dff_B_eEfCfQXT7_1;
	wire w_dff_B_HTVDmjNe4_1;
	wire w_dff_B_bA9Iry2k2_1;
	wire w_dff_B_xcpF8nml9_1;
	wire w_dff_B_OyxFWTsp4_1;
	wire w_dff_B_qoWgq2Zp2_1;
	wire w_dff_B_u6EardZn0_1;
	wire w_dff_B_of8g8xc52_1;
	wire w_dff_B_Qasj3y822_1;
	wire w_dff_B_g0HV2ilx8_1;
	wire w_dff_B_A5sm3Avt5_1;
	wire w_dff_B_xuTN1zfU2_1;
	wire w_dff_B_0NtVP1NK5_1;
	wire w_dff_B_gZlEn6vm6_1;
	wire w_dff_B_VyAkWJzf9_1;
	wire w_dff_B_6piPLQWx6_1;
	wire w_dff_B_XehIwMva3_1;
	wire w_dff_A_dkFBMNyd3_0;
	wire w_dff_A_IYbI70kl3_0;
	wire w_dff_A_RV4KjewY1_0;
	wire w_dff_A_AD3xpUNw8_0;
	wire w_dff_A_pZk4GdOh0_0;
	wire w_dff_A_T0CF8oMq8_0;
	wire w_dff_A_eUxaKqhA6_0;
	wire w_dff_A_FHxmToAu5_0;
	wire w_dff_A_QsmErd6W4_0;
	wire w_dff_A_MnpNT35V7_0;
	wire w_dff_A_aQIKJJWY2_0;
	wire w_dff_A_51EP7Rqb8_0;
	wire w_dff_A_DPrAYKxd9_0;
	wire w_dff_A_BJjSs7Ka8_0;
	wire w_dff_A_6lMKKesw8_0;
	wire w_dff_A_oII8ASb93_0;
	wire w_dff_A_5vYfnKTv1_0;
	wire w_dff_A_TObYhCgW7_0;
	wire w_dff_A_0DYMsleC5_0;
	wire w_dff_A_fhKsflu15_0;
	wire w_dff_A_6DrtfXqu5_0;
	wire w_dff_A_yL4F9Vsb6_0;
	wire w_dff_A_waY3hmgA8_0;
	wire w_dff_A_KBExpihi0_0;
	wire w_dff_A_YskG4wLk4_0;
	wire w_dff_A_qpxTXPI91_0;
	wire w_dff_A_QwLV5MNt0_0;
	wire w_dff_A_xzuvi9cr1_0;
	wire w_dff_A_deE9DqQJ7_0;
	wire w_dff_A_KaBZbPk31_0;
	wire w_dff_A_OkqWzp1N0_0;
	wire w_dff_A_Ofu4lpNa4_0;
	wire w_dff_A_MQKVLyyw0_0;
	wire w_dff_A_I2smT1Jo3_0;
	wire w_dff_A_W7hnBpyI7_0;
	wire w_dff_A_bLF0rPgD2_0;
	wire w_dff_A_4iRi0tfL7_0;
	wire w_dff_A_MyPZGV0G3_0;
	wire w_dff_A_hATT4C2w2_1;
	wire w_dff_B_YKDZx7fy4_1;
	wire w_dff_B_30CAmLrj8_1;
	wire w_dff_B_0YaJDvfN2_1;
	wire w_dff_B_xYO3EXLV4_1;
	wire w_dff_B_YRhavu0M3_1;
	wire w_dff_B_gWiVubG23_1;
	wire w_dff_B_h6IxwEcD2_1;
	wire w_dff_B_o8F9vjcx2_1;
	wire w_dff_B_rd95D0NW5_1;
	wire w_dff_B_f2dDuNHD4_1;
	wire w_dff_B_6UVGXx0J7_1;
	wire w_dff_B_zzhPxBZM3_1;
	wire w_dff_B_Le6VQwOB4_1;
	wire w_dff_B_ViuBbaOd0_1;
	wire w_dff_B_8AZluf0v6_1;
	wire w_dff_B_JUi4qjU18_1;
	wire w_dff_B_JtZdrjT47_1;
	wire w_dff_B_B4lfhRrp4_1;
	wire w_dff_B_ebo5fi4h9_1;
	wire w_dff_B_Zr7omRJh7_1;
	wire w_dff_B_2K1G3JGf0_1;
	wire w_dff_B_UuRafueM8_1;
	wire w_dff_B_jkTLqjWb8_1;
	wire w_dff_B_hMUURlBV9_1;
	wire w_dff_B_WbWycBrW8_1;
	wire w_dff_B_ItSywzld8_1;
	wire w_dff_B_ItYAKeDP6_1;
	wire w_dff_B_ogltcAiF7_1;
	wire w_dff_B_sz1Trnej1_1;
	wire w_dff_B_Tqtrvtr68_1;
	wire w_dff_B_5KlUi48L2_1;
	wire w_dff_B_mFQJulWB4_1;
	wire w_dff_B_MA7cwNGm2_1;
	wire w_dff_B_gR0O5Ao48_1;
	wire w_dff_B_ycRlJSps1_1;
	wire w_dff_A_p7GUuktE2_0;
	wire w_dff_A_WHpTdWff5_0;
	wire w_dff_A_XCfgdy1a4_0;
	wire w_dff_A_DRj5AaGN2_0;
	wire w_dff_A_94I3XL4l4_0;
	wire w_dff_A_yy9zWcg31_0;
	wire w_dff_A_JeXyUzJI4_0;
	wire w_dff_A_p4iV8HMX0_0;
	wire w_dff_A_fPsliYym6_0;
	wire w_dff_A_ZKMmuNkq9_0;
	wire w_dff_A_gwudE4ZE6_0;
	wire w_dff_A_9io5mtJi6_0;
	wire w_dff_A_yYey6hKF0_0;
	wire w_dff_A_ZC2toaYY2_0;
	wire w_dff_A_I5CCOEl28_0;
	wire w_dff_A_Q1PIakiP2_0;
	wire w_dff_A_HoZCIjjc0_0;
	wire w_dff_A_gBioCk720_0;
	wire w_dff_A_fiU2mHFd9_0;
	wire w_dff_A_Gb6RctpV2_0;
	wire w_dff_A_A3rKjPti5_0;
	wire w_dff_A_8ueIGBPZ8_0;
	wire w_dff_A_MhypBxVz4_0;
	wire w_dff_A_PXkaP1gN3_0;
	wire w_dff_A_lTvnh4hg6_0;
	wire w_dff_A_401zNE1z2_0;
	wire w_dff_A_HiI0Rbrh6_0;
	wire w_dff_A_yB0SWjtR4_0;
	wire w_dff_A_BtnbUn9A9_0;
	wire w_dff_A_wYQVAkQO0_0;
	wire w_dff_A_CyWGjM0H9_0;
	wire w_dff_A_KQhmwlZn2_0;
	wire w_dff_A_3WzrqVap0_0;
	wire w_dff_A_AS5QDOLL6_0;
	wire w_dff_A_U6tTMT4n6_0;
	wire w_dff_A_aPxlJXc64_1;
	wire w_dff_B_iy31NKBE3_1;
	wire w_dff_B_RTB9HEF04_1;
	wire w_dff_B_I7c2d6g67_1;
	wire w_dff_B_gBizV6y55_1;
	wire w_dff_B_a2aYoDrQ9_1;
	wire w_dff_B_TBDvLm7N3_1;
	wire w_dff_B_IqOAo8VR3_1;
	wire w_dff_B_OSVZOmad4_1;
	wire w_dff_B_zCNee9JC4_1;
	wire w_dff_B_4ver7lNm3_1;
	wire w_dff_B_uiigXH6p4_1;
	wire w_dff_B_8VcGRPQe1_1;
	wire w_dff_B_Vxa46z4X8_1;
	wire w_dff_B_nnl1cWl62_1;
	wire w_dff_B_SEmewUDT4_1;
	wire w_dff_B_T4XHIcec4_1;
	wire w_dff_B_sKOzv35U8_1;
	wire w_dff_B_yEvHS9qk0_1;
	wire w_dff_B_Ips5b0QF2_1;
	wire w_dff_B_UWKtcUi81_1;
	wire w_dff_B_L4HA2sbK5_1;
	wire w_dff_B_YydlJqw35_1;
	wire w_dff_B_bZESkjES9_1;
	wire w_dff_B_5Uifv4636_1;
	wire w_dff_B_nyAcTbUx9_1;
	wire w_dff_B_quG33DA47_1;
	wire w_dff_B_DagU8vkE8_1;
	wire w_dff_B_NdnLBpy36_1;
	wire w_dff_B_qzLi7wxI0_1;
	wire w_dff_B_vFSrm8xK7_1;
	wire w_dff_B_fSmRDmHs5_1;
	wire w_dff_B_qOHS1r4z9_1;
	wire w_dff_A_25J1ABlK1_0;
	wire w_dff_A_dN3XHPRR1_0;
	wire w_dff_A_xhb7EiLO9_0;
	wire w_dff_A_fiM37NNF6_0;
	wire w_dff_A_Vt79zmtK1_0;
	wire w_dff_A_X86iegjD5_0;
	wire w_dff_A_1GqdSVGj9_0;
	wire w_dff_A_vNkKSNx74_0;
	wire w_dff_A_At5yY3qr4_0;
	wire w_dff_A_GGZLjlkr5_0;
	wire w_dff_A_JQnaDncF0_0;
	wire w_dff_A_gHGlTTdY7_0;
	wire w_dff_A_jEfy5eT24_0;
	wire w_dff_A_6IQDB7TZ7_0;
	wire w_dff_A_E7tr3AmN3_0;
	wire w_dff_A_hleiiF2t2_0;
	wire w_dff_A_eqLjgLOn4_0;
	wire w_dff_A_91W6l9NE5_0;
	wire w_dff_A_9e2Mw5bp3_0;
	wire w_dff_A_Bulf4hA77_0;
	wire w_dff_A_7HAxMaP98_0;
	wire w_dff_A_53WWlr557_0;
	wire w_dff_A_VJ9VPnRZ1_0;
	wire w_dff_A_1mR2f2WZ5_0;
	wire w_dff_A_pAYbq8Wm4_0;
	wire w_dff_A_vpfnu7Zo2_0;
	wire w_dff_A_8QmlS4kl5_0;
	wire w_dff_A_YVshM2O80_0;
	wire w_dff_A_BbvnutCV7_0;
	wire w_dff_A_9bNkaOUZ7_0;
	wire w_dff_A_3Z9gBS8J2_0;
	wire w_dff_A_QyYqNGcL2_0;
	wire w_dff_A_y52OnWIm4_1;
	wire w_dff_B_03OhajKk6_1;
	wire w_dff_B_78yyYrFy9_1;
	wire w_dff_B_gP9qIGun5_1;
	wire w_dff_B_a0D0ATka5_1;
	wire w_dff_B_r5GjRDuH9_1;
	wire w_dff_B_uyfJ7Mt46_1;
	wire w_dff_B_vEwSBPt70_1;
	wire w_dff_B_shnxaGXY8_1;
	wire w_dff_B_sjrSdDmm3_1;
	wire w_dff_B_WpSDGyFr8_1;
	wire w_dff_B_YSayJaUO7_1;
	wire w_dff_B_L1y1wUmA7_1;
	wire w_dff_B_DhnnIlKP4_1;
	wire w_dff_B_aPPAH2Ah1_1;
	wire w_dff_B_CbCL1So65_1;
	wire w_dff_B_tF0PQgSd6_1;
	wire w_dff_B_W1EZMm6m4_1;
	wire w_dff_B_HBH1vVDM0_1;
	wire w_dff_B_GobGod4P7_1;
	wire w_dff_B_lg1clGu56_1;
	wire w_dff_B_VGX2ImSY9_1;
	wire w_dff_B_old76uYA3_1;
	wire w_dff_B_WLCDqwmH1_1;
	wire w_dff_B_OiiVPp338_1;
	wire w_dff_B_TzjhTPpi6_1;
	wire w_dff_B_SMsTbFdw7_1;
	wire w_dff_B_rrKbl2Oz7_1;
	wire w_dff_B_9nDqJSLu7_1;
	wire w_dff_B_DQfbDQM90_1;
	wire w_dff_A_koecHf197_0;
	wire w_dff_A_88of4Y3H2_0;
	wire w_dff_A_zUKI2ipk6_0;
	wire w_dff_A_Mg1QMq1y0_0;
	wire w_dff_A_KO8gUpMt8_0;
	wire w_dff_A_bZyjf5QM0_0;
	wire w_dff_A_Jp87AN728_0;
	wire w_dff_A_Vw0XLAzK7_0;
	wire w_dff_A_j1sNWFGB9_0;
	wire w_dff_A_nX2OLA8t1_0;
	wire w_dff_A_3bBkmYjL4_0;
	wire w_dff_A_GeiHwEMD0_0;
	wire w_dff_A_WZnIHl6l9_0;
	wire w_dff_A_p5kFz4gF7_0;
	wire w_dff_A_sx8ig0DO6_0;
	wire w_dff_A_mYZKCLuz6_0;
	wire w_dff_A_1oFOzSW69_0;
	wire w_dff_A_uGPvtTVX7_0;
	wire w_dff_A_zZu1xyvL2_0;
	wire w_dff_A_VybmS4eT2_0;
	wire w_dff_A_j5yhgpTH9_0;
	wire w_dff_A_VW0iDvQY7_0;
	wire w_dff_A_lVUI89H38_0;
	wire w_dff_A_vcBEXZuq6_0;
	wire w_dff_A_QF69uTUZ8_0;
	wire w_dff_A_iaD0Ui6t2_0;
	wire w_dff_A_E4NDaTF07_0;
	wire w_dff_A_3CQsH5Ge1_0;
	wire w_dff_A_Bh1ZRL9E6_0;
	wire w_dff_A_CjzJvrro2_1;
	wire w_dff_B_jPf9d1437_1;
	wire w_dff_B_PMZhOHfG5_1;
	wire w_dff_B_7m5Ljs6L5_1;
	wire w_dff_B_91Eq0bsZ1_1;
	wire w_dff_B_caNJuHBv3_1;
	wire w_dff_B_uq5XLDR71_1;
	wire w_dff_B_7sdbKtDC6_1;
	wire w_dff_B_Hhdpf7DE2_1;
	wire w_dff_B_6UqegZxt9_1;
	wire w_dff_B_sU8svXl31_1;
	wire w_dff_B_Stgp5cb35_1;
	wire w_dff_B_qngqHhWW7_1;
	wire w_dff_B_tZVYjBeh0_1;
	wire w_dff_B_Ar81sFvH3_1;
	wire w_dff_B_3P3blIMd6_1;
	wire w_dff_B_tGnemvza7_1;
	wire w_dff_B_TSPrvUGD6_1;
	wire w_dff_B_FdpkVCvy7_1;
	wire w_dff_B_cLibVtUJ7_1;
	wire w_dff_B_hra5wWkj4_1;
	wire w_dff_B_L4Z2YD5P5_1;
	wire w_dff_B_zBbDLL0r2_1;
	wire w_dff_B_V8cBGbxW4_1;
	wire w_dff_B_cUpVF8kC7_1;
	wire w_dff_B_wop3Ppbk9_1;
	wire w_dff_B_ZBjdgUM75_1;
	wire w_dff_A_4yTvoOGG4_0;
	wire w_dff_A_f4aJ6Dam8_0;
	wire w_dff_A_lH0gg2iX6_0;
	wire w_dff_A_zUAKggiq6_0;
	wire w_dff_A_vNUFrGXP7_0;
	wire w_dff_A_UfxBdeRD1_0;
	wire w_dff_A_VdQzMsFY8_0;
	wire w_dff_A_GhDlmh643_0;
	wire w_dff_A_6B1Ba9kp1_0;
	wire w_dff_A_Orz0hikz5_0;
	wire w_dff_A_t472kEWT1_0;
	wire w_dff_A_r2bAcMBp7_0;
	wire w_dff_A_kuDJKgVV6_0;
	wire w_dff_A_4EAKvhJF0_0;
	wire w_dff_A_ScwgxVOV1_0;
	wire w_dff_A_xDNSVloW3_0;
	wire w_dff_A_mJ4UpHWR6_0;
	wire w_dff_A_FQBlAXKf7_0;
	wire w_dff_A_2rVn07hh8_0;
	wire w_dff_A_xaaj5BxM3_0;
	wire w_dff_A_ApncF34F8_0;
	wire w_dff_A_HfF4ygvD2_0;
	wire w_dff_A_TwrHOL4N2_0;
	wire w_dff_A_WBeW4mnR4_0;
	wire w_dff_A_f5dVDaYY7_0;
	wire w_dff_A_t8tAzgMp1_0;
	wire w_dff_A_CHZGfPAc5_1;
	wire w_dff_B_uPooh4ko2_1;
	wire w_dff_B_jB9bx6RJ4_1;
	wire w_dff_B_rEj5h7iN0_1;
	wire w_dff_B_y2Bpli1n5_1;
	wire w_dff_B_z1Cb8xDh4_1;
	wire w_dff_B_fg0i13d87_1;
	wire w_dff_B_KXGIOptQ6_1;
	wire w_dff_B_jcuzs3am8_1;
	wire w_dff_B_mSXkN6kp4_1;
	wire w_dff_B_noNM6B8J1_1;
	wire w_dff_B_O0RoGiIr8_1;
	wire w_dff_B_VDCUgvIi3_1;
	wire w_dff_B_GnCt8pN18_1;
	wire w_dff_B_V9ew3Jy92_1;
	wire w_dff_B_i0ViKzR78_1;
	wire w_dff_B_6ylNFGro7_1;
	wire w_dff_B_ACRkX0KM3_1;
	wire w_dff_B_LZbVOwwh8_1;
	wire w_dff_B_IH4X7iGM9_1;
	wire w_dff_B_yu6bXgS87_1;
	wire w_dff_B_k6SXAJtP2_1;
	wire w_dff_B_v1w7e7PW8_1;
	wire w_dff_B_AjWbN0rr3_1;
	wire w_dff_A_6PiLb6KC4_0;
	wire w_dff_A_Bb9UfAdB0_0;
	wire w_dff_A_HPwUAGCC3_0;
	wire w_dff_A_dFCAAs831_0;
	wire w_dff_A_Iy9sInHu9_0;
	wire w_dff_A_VclKgW8m9_0;
	wire w_dff_A_qI9EW8fy2_0;
	wire w_dff_A_xyJySTWb1_0;
	wire w_dff_A_JSmQBqyU7_0;
	wire w_dff_A_TtAhHQGa5_0;
	wire w_dff_A_RSrEA1wc2_0;
	wire w_dff_A_2eu7Rc9D6_0;
	wire w_dff_A_ke2CuF9w4_0;
	wire w_dff_A_DmWln3eR4_0;
	wire w_dff_A_JLIO5ySW8_0;
	wire w_dff_A_QR3vwlDf0_0;
	wire w_dff_A_lYlufg023_0;
	wire w_dff_A_k4nutc9v4_0;
	wire w_dff_A_vpDUgNWM4_0;
	wire w_dff_A_xMXRsrhP8_0;
	wire w_dff_A_naWIhevA7_0;
	wire w_dff_A_V1cu7Egm0_0;
	wire w_dff_A_eUbJdN5F3_0;
	wire w_dff_A_peHk2qng5_1;
	wire w_dff_B_3jm1LoUs7_1;
	wire w_dff_B_5OHO6uYD6_1;
	wire w_dff_B_YdpCmWmt5_1;
	wire w_dff_B_d2BgRoeI9_1;
	wire w_dff_B_XfRatf0y3_1;
	wire w_dff_B_zgYCR2wc2_1;
	wire w_dff_B_3nhwhcBJ4_1;
	wire w_dff_B_6ETBEvVU5_1;
	wire w_dff_B_JKJeDhBx4_1;
	wire w_dff_B_z2UOf6LZ5_1;
	wire w_dff_B_3Tk7LKh01_1;
	wire w_dff_B_5MH3Oeh13_1;
	wire w_dff_B_t99yLnjP3_1;
	wire w_dff_B_ECHD0jid6_1;
	wire w_dff_B_lksvYya75_1;
	wire w_dff_B_jqsJEwL29_1;
	wire w_dff_B_g0eg8jXV5_1;
	wire w_dff_B_umj1hFfn6_1;
	wire w_dff_B_U0LQCSR08_1;
	wire w_dff_B_pRSP3AEO9_1;
	wire w_dff_A_9DNkYF7O1_0;
	wire w_dff_A_MTW7eLSF3_0;
	wire w_dff_A_XOaFlA969_0;
	wire w_dff_A_vW6bK1cy4_0;
	wire w_dff_A_Db1PgHsM6_0;
	wire w_dff_A_wXTeGHmP5_0;
	wire w_dff_A_57S724kv0_0;
	wire w_dff_A_cHuF6PXi2_0;
	wire w_dff_A_lIFHSSwv1_0;
	wire w_dff_A_UW6i24ke9_0;
	wire w_dff_A_hz9fPhRz7_0;
	wire w_dff_A_7RfluJ9C7_0;
	wire w_dff_A_2CBO0o5u6_0;
	wire w_dff_A_wPxwHqT10_0;
	wire w_dff_A_TQfBR9oN4_0;
	wire w_dff_A_WyQ6RYTx7_0;
	wire w_dff_A_eCWI2sTG8_0;
	wire w_dff_A_S0RWZkCc7_0;
	wire w_dff_A_5eQzsYTy1_0;
	wire w_dff_A_edGf9AFJ6_0;
	wire w_dff_A_tZxpkrLk3_1;
	wire w_dff_B_h6JbXv9q1_1;
	wire w_dff_B_5pF6I5F77_1;
	wire w_dff_B_vVA7RSmo9_1;
	wire w_dff_B_mARE0DzF5_1;
	wire w_dff_B_jZnpDUjS2_1;
	wire w_dff_B_MBIWsY8n5_1;
	wire w_dff_B_JebC4doU8_1;
	wire w_dff_B_0k6QPpgW6_1;
	wire w_dff_B_0K1i2wLI0_1;
	wire w_dff_B_8ETZk4Mc5_1;
	wire w_dff_B_DqYHRLOG4_1;
	wire w_dff_B_VOnfjZ3w1_1;
	wire w_dff_B_k9OxSITD3_1;
	wire w_dff_B_CjOzhyUA6_1;
	wire w_dff_B_wpjKZvYm1_1;
	wire w_dff_B_txgUulhx8_1;
	wire w_dff_B_rd8mdpko9_1;
	wire w_dff_A_jFTrrHOP4_0;
	wire w_dff_A_HnMp1a7O1_0;
	wire w_dff_A_QOFFq5fX4_0;
	wire w_dff_A_YsTdaKn61_0;
	wire w_dff_A_55FDEM2a4_0;
	wire w_dff_A_0MrTwIOG1_0;
	wire w_dff_A_wLDUqIBe9_0;
	wire w_dff_A_GCZtswWN6_0;
	wire w_dff_A_0h0x7GFn7_0;
	wire w_dff_A_kXcckj9G0_0;
	wire w_dff_A_qLW1G1338_0;
	wire w_dff_A_a3wbc89U7_0;
	wire w_dff_A_UoZYWiHc9_0;
	wire w_dff_A_HDQ0hPqB8_0;
	wire w_dff_A_SJPEAaCf7_0;
	wire w_dff_A_OV18yayR5_0;
	wire w_dff_A_Ond58uNP5_0;
	wire w_dff_A_iWmMC9ts3_1;
	wire w_dff_B_bbmCodpv9_1;
	wire w_dff_B_T3DLMfQa1_1;
	wire w_dff_B_ZGze8S695_1;
	wire w_dff_B_KelZoE8Z9_1;
	wire w_dff_B_WZqPo0yc3_1;
	wire w_dff_B_u1qfyp3f0_1;
	wire w_dff_B_VZCzrF6J2_1;
	wire w_dff_B_ld2M7Io84_1;
	wire w_dff_B_ej3hterM9_1;
	wire w_dff_B_BNA27gul1_1;
	wire w_dff_B_1dBIy7716_1;
	wire w_dff_B_9B6EDUzt7_1;
	wire w_dff_B_AmcbYULr1_1;
	wire w_dff_B_AwKqnTL31_1;
	wire w_dff_A_DJjqOhdm7_0;
	wire w_dff_A_YvHKOKcx4_0;
	wire w_dff_A_eVvSIuyt5_0;
	wire w_dff_A_TroSCxah7_0;
	wire w_dff_A_9WzLxNoc4_0;
	wire w_dff_A_0DsPOaC91_0;
	wire w_dff_A_SUaqs6Qk8_0;
	wire w_dff_A_vedmNpOY1_0;
	wire w_dff_A_hzU4Gapk7_0;
	wire w_dff_A_DU3UOxV42_0;
	wire w_dff_A_9hV77ayo2_0;
	wire w_dff_A_T6AGU7rH3_0;
	wire w_dff_A_CCzX6Ho66_0;
	wire w_dff_A_0h3CobnG1_0;
	wire w_dff_A_kqbN4kqC7_1;
	wire w_dff_B_WDHxITla2_1;
	wire w_dff_B_YHInVKxR8_1;
	wire w_dff_B_zeOKIsAd7_1;
	wire w_dff_B_fdAkYsbd6_1;
	wire w_dff_B_rndcK6l50_1;
	wire w_dff_B_5Mq1T8Oi4_1;
	wire w_dff_B_nBl7lXVE3_1;
	wire w_dff_B_EdRrC5GC0_1;
	wire w_dff_B_0vCdFfoY2_1;
	wire w_dff_B_Y7QU2Ebk7_1;
	wire w_dff_B_TKqaCuwG8_1;
	wire w_dff_A_8kpIdcK42_0;
	wire w_dff_A_8D7AhApE5_0;
	wire w_dff_A_h55Xr0L76_0;
	wire w_dff_A_BcyEWGfB6_0;
	wire w_dff_A_uo5N9op78_0;
	wire w_dff_A_22USeGXd2_0;
	wire w_dff_A_HducLP3S1_0;
	wire w_dff_A_NOebkhnB5_0;
	wire w_dff_A_zww6rqlG3_0;
	wire w_dff_A_r6DPxvsI5_0;
	wire w_dff_A_Tooep5n49_0;
	wire w_dff_A_VpV1Wt6x7_1;
	wire w_dff_B_FxJTXI7R9_1;
	wire w_dff_B_y8vDRHA60_1;
	wire w_dff_B_63Slu4xQ8_1;
	wire w_dff_B_Rf2K9rdr8_1;
	wire w_dff_B_42yb08Af2_1;
	wire w_dff_B_19nrQdrO5_1;
	wire w_dff_B_tBHNWRrm0_1;
	wire w_dff_B_1qvD8ff13_1;
	wire w_dff_A_dTyP0f7L8_0;
	wire w_dff_A_bV00JtyD4_0;
	wire w_dff_A_U1trpJOS5_0;
	wire w_dff_A_ePo85IVu4_0;
	wire w_dff_A_ruNAtg1E0_0;
	wire w_dff_A_aYd37mFd2_0;
	wire w_dff_A_BE4QZEcY8_0;
	wire w_dff_A_JUvwpQwb8_0;
	wire w_dff_A_YXMU8p9c8_1;
	wire w_dff_B_6LZmB3Gn3_1;
	wire w_dff_B_012J1un06_1;
	wire w_dff_B_OxwRlb8w7_1;
	wire w_dff_B_jffWmVSl8_1;
	wire w_dff_B_GUp30YFz8_1;
	wire w_dff_B_CNllXBTv4_0;
	wire w_dff_A_gix6zsfO9_0;
	wire w_dff_A_IN8XLFiq7_0;
	wire w_dff_A_OgaaY1J50_0;
	wire w_dff_A_FLj6H75i3_0;
	wire w_dff_A_MuhjVLNl5_0;
	wire w_dff_A_nYOTDYLC5_0;
	wire w_dff_A_uhOhIG0A7_0;
	wire w_dff_A_HyISg1en7_1;
	wire w_dff_B_oFoXuBJi1_1;
	wire w_dff_B_uu5s7mxV8_2;
	wire w_dff_B_RrcJzKsF4_2;
	wire w_dff_B_RM9G0PvZ0_2;
	wire w_dff_B_s4PasYeV7_2;
	wire w_dff_B_vxw4WpAf9_2;
	wire w_dff_B_CIWvcv9n0_2;
	wire w_dff_B_zrqvvdgs2_2;
	wire w_dff_B_ibP34pDL5_2;
	wire w_dff_B_KvdxSQg76_2;
	wire w_dff_B_qS1V03CX0_2;
	wire w_dff_B_Z0CElkhq4_2;
	wire w_dff_B_Z4oX2eZC2_2;
	wire w_dff_B_mmnzgVYX2_2;
	wire w_dff_B_nIFa6QTK4_2;
	wire w_dff_B_jmxhQi6B0_2;
	wire w_dff_B_TCn8qOCJ0_2;
	wire w_dff_B_5LFSMMoA6_2;
	wire w_dff_B_VltZJW6A5_2;
	wire w_dff_B_N1Y9uENj0_2;
	wire w_dff_B_sYSfSS3X1_2;
	wire w_dff_B_GgAsFdPT7_2;
	wire w_dff_B_wFhOb4C65_2;
	wire w_dff_B_ESdU0vGh2_2;
	wire w_dff_B_3V9cVasK4_2;
	wire w_dff_B_0cHK6SdN2_2;
	wire w_dff_B_5mXlmx2L3_2;
	wire w_dff_B_wGCg2bAy6_2;
	wire w_dff_B_RVQJ6Jm35_2;
	wire w_dff_B_ja9cWSXL8_2;
	wire w_dff_B_Se2B2VG83_2;
	wire w_dff_B_IiGk1jLN6_2;
	wire w_dff_B_4VFrOGka8_2;
	wire w_dff_B_zSN1oP7s0_2;
	wire w_dff_B_SzOasAmJ6_2;
	wire w_dff_B_Sn72WNp93_2;
	wire w_dff_B_aUPtDaFI0_2;
	wire w_dff_B_DJwCsm9G0_2;
	wire w_dff_B_iBTf6qWn7_2;
	wire w_dff_B_LSnm5eJl7_2;
	wire w_dff_B_pBlO0dTg7_2;
	wire w_dff_B_mtHqs9xD2_2;
	wire w_dff_B_bvKCUuvs3_2;
	wire w_dff_B_QGnr771I8_2;
	wire w_dff_B_OUTFygTT9_2;
	wire w_dff_A_8FZFsssn1_0;
	wire w_dff_B_YU9Fs9yY9_1;
	wire w_dff_B_Cmju4XkZ6_2;
	wire w_dff_B_XKJLECiX2_2;
	wire w_dff_B_9iJPZpOG0_2;
	wire w_dff_B_riD7Hhbp0_2;
	wire w_dff_B_MUBFnhlV8_2;
	wire w_dff_B_oWvVhCi61_2;
	wire w_dff_B_244JvJfI4_2;
	wire w_dff_B_smPeRvbF6_2;
	wire w_dff_B_144CYuEf9_2;
	wire w_dff_B_VUKIUUqr1_2;
	wire w_dff_B_89P51siD4_2;
	wire w_dff_B_53acqq0B2_2;
	wire w_dff_B_QZyI493c2_2;
	wire w_dff_B_ieQuILvB7_2;
	wire w_dff_B_9XVzMyIm3_2;
	wire w_dff_B_CBSWQztz5_2;
	wire w_dff_B_rLPlqZ4P8_2;
	wire w_dff_B_V0N7pwgU0_2;
	wire w_dff_B_mJkgIjw38_2;
	wire w_dff_B_7JTOvEP82_2;
	wire w_dff_B_PexFvD751_2;
	wire w_dff_B_cONiCm715_2;
	wire w_dff_B_1rjeMho76_2;
	wire w_dff_B_53CgxPdn7_2;
	wire w_dff_B_HFO9JKgM9_2;
	wire w_dff_B_gNeO94Sq5_2;
	wire w_dff_B_8ZKoRUde3_2;
	wire w_dff_B_Kce3qLiA4_2;
	wire w_dff_B_N0iyvKSp3_2;
	wire w_dff_B_7hRlI4ES7_2;
	wire w_dff_B_KpSFj8zI0_2;
	wire w_dff_B_hFDt0Kgj7_2;
	wire w_dff_B_uIG9bSch6_2;
	wire w_dff_B_MO1mBpfc0_2;
	wire w_dff_B_PpjVTIOw8_2;
	wire w_dff_B_5MoCXwDb0_2;
	wire w_dff_B_wR1jJcqr2_2;
	wire w_dff_B_exRrguur1_2;
	wire w_dff_B_wcFWD4uh4_2;
	wire w_dff_B_RRR1lM4Q7_2;
	wire w_dff_B_N6d7RHoj3_2;
	wire w_dff_A_hHU6UceV1_1;
	wire w_dff_B_fzzOmr8J1_1;
	wire w_dff_B_yIf3oAeV5_1;
	wire w_dff_B_n1ODXD237_1;
	wire w_dff_B_wsJVEs0y7_1;
	wire w_dff_B_E0fa8WJR7_1;
	wire w_dff_B_4P9o2Dp96_1;
	wire w_dff_B_xnWLgX6V4_1;
	wire w_dff_B_UY0riLX37_1;
	wire w_dff_B_3BS2JmOQ3_1;
	wire w_dff_B_GSLimxgR9_1;
	wire w_dff_B_xlxmilYB6_1;
	wire w_dff_B_g0smN5WD2_1;
	wire w_dff_B_pZCtFNNp6_1;
	wire w_dff_B_YwwKu8VX9_1;
	wire w_dff_B_reuRlGSb4_1;
	wire w_dff_B_LDMW8fnj0_1;
	wire w_dff_B_ldAQpglH3_1;
	wire w_dff_B_U8ofqQwm2_1;
	wire w_dff_B_rsk4C2hf8_1;
	wire w_dff_B_0kIq5otZ5_1;
	wire w_dff_B_KghDC9zd6_1;
	wire w_dff_B_mcbKVaae7_1;
	wire w_dff_B_3jhVv5In6_1;
	wire w_dff_B_b8eEDtjU1_1;
	wire w_dff_B_iqDhQZyc2_1;
	wire w_dff_B_8xbn7ygX3_1;
	wire w_dff_B_SOSxbKXV8_1;
	wire w_dff_B_FGd2q3r20_1;
	wire w_dff_B_MAUVOqBM6_1;
	wire w_dff_B_hzdiH5tC3_1;
	wire w_dff_B_wQDkuLSQ2_1;
	wire w_dff_B_gnZ80UEL4_1;
	wire w_dff_B_6RSExyqG0_1;
	wire w_dff_B_TEwbDJuc7_1;
	wire w_dff_B_xxvzGOjw8_1;
	wire w_dff_B_k2Occ9hC0_1;
	wire w_dff_B_VV2MIwFT6_1;
	wire w_dff_B_KpqY4Roc0_1;
	wire w_dff_A_0x7sXd5j0_0;
	wire w_dff_A_1t0KfLDD4_0;
	wire w_dff_A_c1C5p1y66_0;
	wire w_dff_A_OEpCSvpc2_0;
	wire w_dff_A_HboQAD2X9_0;
	wire w_dff_A_VSaBkZhR9_0;
	wire w_dff_A_tx41zBWz7_0;
	wire w_dff_A_ar4OMavj3_0;
	wire w_dff_A_3kyOvU4F9_0;
	wire w_dff_A_QqCw3m452_0;
	wire w_dff_A_2TVhhPhf6_0;
	wire w_dff_A_eQ9CyBdA7_0;
	wire w_dff_A_Q6Bpm4h13_0;
	wire w_dff_A_zz8k9yHb4_0;
	wire w_dff_A_itMEMbUa8_0;
	wire w_dff_A_gP9gCfzn7_0;
	wire w_dff_A_EPexjiHt3_0;
	wire w_dff_A_gpcO4scG3_0;
	wire w_dff_A_hISEMg0b2_0;
	wire w_dff_A_AErJsgPT6_0;
	wire w_dff_A_XnsgTuen7_0;
	wire w_dff_A_gSUsSpUM9_0;
	wire w_dff_A_xJh2KpoY8_0;
	wire w_dff_A_aqHw9f9o2_0;
	wire w_dff_A_Z1OQV4rR3_0;
	wire w_dff_A_aW88qQaB0_0;
	wire w_dff_A_dBKO5jgt7_0;
	wire w_dff_A_tvTL01T53_0;
	wire w_dff_A_0NIWXbRw4_0;
	wire w_dff_A_RF6jJ1qM4_0;
	wire w_dff_A_wpKf0Pax1_0;
	wire w_dff_A_cSGwaseN9_0;
	wire w_dff_A_IqWGRieV0_0;
	wire w_dff_A_MquVKvAs7_0;
	wire w_dff_A_iK6EvYbl7_0;
	wire w_dff_A_ojtGVxro0_0;
	wire w_dff_A_VdfbowkM1_0;
	wire w_dff_A_7YxzHdl95_0;
	wire w_dff_A_CZ2jEFdf6_0;
	wire w_dff_B_n1qofQ7N6_1;
	wire w_dff_A_To4CQYwR5_0;
	wire w_dff_A_ggh7op5Z7_0;
	wire w_dff_A_yxOIQ4lR2_0;
	wire w_dff_A_FrkpCw5a8_0;
	wire w_dff_A_JElZmtGa1_0;
	wire w_dff_A_3mFIzyLZ1_0;
	wire w_dff_A_3HmzR6yy1_0;
	wire w_dff_A_RlOVBzJF3_0;
	wire w_dff_A_eCWTqBit2_0;
	wire w_dff_A_smlIJURR8_0;
	wire w_dff_A_Aeraraba3_0;
	wire w_dff_A_WbXmNPCy1_0;
	wire w_dff_A_fzBGNR4C0_0;
	wire w_dff_A_pDscmNUD6_0;
	wire w_dff_A_1rabCNHB7_0;
	wire w_dff_A_tEb8e0M24_0;
	wire w_dff_A_EWJSBKE89_0;
	wire w_dff_A_GMdCjHzv1_0;
	wire w_dff_A_8DzFQCZx0_0;
	wire w_dff_A_5gg0W96i4_0;
	wire w_dff_A_mF2BH9hX5_0;
	wire w_dff_A_6qLITpxo1_0;
	wire w_dff_A_gvQuIHqD6_0;
	wire w_dff_A_np2AACK71_0;
	wire w_dff_A_dSSqv5el9_0;
	wire w_dff_A_6ZcnzBpi8_0;
	wire w_dff_A_9TJo8J1h8_0;
	wire w_dff_A_A3svwYQ96_0;
	wire w_dff_A_wgUbjRhB2_0;
	wire w_dff_A_7HSPdK1j0_0;
	wire w_dff_A_htXIfznG4_0;
	wire w_dff_A_WKGGiWb44_0;
	wire w_dff_A_XareqLXt0_0;
	wire w_dff_A_gM7V1X5D8_0;
	wire w_dff_A_1KDVfjr33_0;
	wire w_dff_A_OgeeSzwv6_0;
	wire w_dff_B_T0JlXUcf3_1;
	wire w_dff_A_1FBtlnJd4_0;
	wire w_dff_A_YRhvihQA6_0;
	wire w_dff_A_2u9NoB241_0;
	wire w_dff_A_qw0GAhjs9_0;
	wire w_dff_A_QDn77CaY5_0;
	wire w_dff_A_voPjoagP0_0;
	wire w_dff_A_FJAaoLIb1_0;
	wire w_dff_A_GLoNUQPe4_0;
	wire w_dff_A_hvLyiykL5_0;
	wire w_dff_A_6E27U3Vr7_0;
	wire w_dff_A_kZyClB2W3_0;
	wire w_dff_A_szql5YIY2_0;
	wire w_dff_A_dhUrHtm81_0;
	wire w_dff_A_uVzSUWcq3_0;
	wire w_dff_A_6OhY4Zcq0_0;
	wire w_dff_A_jlwv0Zhf6_0;
	wire w_dff_A_9AwAA0PN1_0;
	wire w_dff_A_jMPHnMES8_0;
	wire w_dff_A_STtMjR668_0;
	wire w_dff_A_i4fnA0FW5_0;
	wire w_dff_A_9ca1J4kT0_0;
	wire w_dff_A_4KZVR7Fb3_0;
	wire w_dff_A_OY8XUwl90_0;
	wire w_dff_A_qWRvH4Bx0_0;
	wire w_dff_A_Vp8wa24D0_0;
	wire w_dff_A_wVfnTa6n8_0;
	wire w_dff_A_ZVuLWI3g9_0;
	wire w_dff_A_ctXthAzv4_0;
	wire w_dff_A_iQzNwUYQ3_0;
	wire w_dff_A_pB3OO0pO7_0;
	wire w_dff_A_w2rvrd2E6_0;
	wire w_dff_A_4Sqb3nNa1_0;
	wire w_dff_A_5WYeOW9D8_0;
	wire w_dff_B_SpoUZEwd0_1;
	wire w_dff_A_BonLGtCS7_0;
	wire w_dff_A_qXCCAQEi7_0;
	wire w_dff_A_hvhrF0bn2_0;
	wire w_dff_A_hZ6uZVYi5_0;
	wire w_dff_A_FpERn6Cd7_0;
	wire w_dff_A_KEBm57gp9_0;
	wire w_dff_A_Ff4uTXqb2_0;
	wire w_dff_A_4KQt9KZB9_0;
	wire w_dff_A_aSzd3V5y7_0;
	wire w_dff_A_eQBooRoZ2_0;
	wire w_dff_A_9EjCucF43_0;
	wire w_dff_A_rnB0gZ014_0;
	wire w_dff_A_D8avDmqJ8_0;
	wire w_dff_A_zjAVnxuZ6_0;
	wire w_dff_A_QgM4FMme2_0;
	wire w_dff_A_6jVIJBg65_0;
	wire w_dff_A_iSLGsF3h3_0;
	wire w_dff_A_FHou2Rh10_0;
	wire w_dff_A_GQCklcge3_0;
	wire w_dff_A_oSYctBLT9_0;
	wire w_dff_A_jFsyfJ843_0;
	wire w_dff_A_eAmjjxs99_0;
	wire w_dff_A_Oa5q03m06_0;
	wire w_dff_A_slspMlqY1_0;
	wire w_dff_A_cSBYrpul6_0;
	wire w_dff_A_lzmXifd79_0;
	wire w_dff_A_InnUBaSo2_0;
	wire w_dff_A_E2J9lZA42_0;
	wire w_dff_A_UZ7DrGWN9_0;
	wire w_dff_A_8tiOknIL2_0;
	wire w_dff_B_wkFc1ith2_1;
	wire w_dff_A_Z0qkaj588_0;
	wire w_dff_A_Mgna3mO74_0;
	wire w_dff_A_0K0H1mcN6_0;
	wire w_dff_A_U8uKCunH7_0;
	wire w_dff_A_ZCcxNhSW5_0;
	wire w_dff_A_Vq4Igk4k9_0;
	wire w_dff_A_leSBSrue9_0;
	wire w_dff_A_a1D3WmsL1_0;
	wire w_dff_A_97FYEoeL1_0;
	wire w_dff_A_NeaUB9Zu6_0;
	wire w_dff_A_wLEdSDoS0_0;
	wire w_dff_A_AZ733hQx0_0;
	wire w_dff_A_owYA2bLA9_0;
	wire w_dff_A_h1BVIcgu9_0;
	wire w_dff_A_OKGD1lo05_0;
	wire w_dff_A_L2wyClKZ6_0;
	wire w_dff_A_1pTA4NV72_0;
	wire w_dff_A_sulAL0da8_0;
	wire w_dff_A_jKqVXPEE7_0;
	wire w_dff_A_5ZzBjgKr7_0;
	wire w_dff_A_fh5MXxQN3_0;
	wire w_dff_A_kCwfeBfB8_0;
	wire w_dff_A_Se7yCc9P7_0;
	wire w_dff_A_alDo3FBj1_0;
	wire w_dff_A_jw9LVS7v8_0;
	wire w_dff_A_pPk0ZHij9_0;
	wire w_dff_A_w7T9nth90_0;
	wire w_dff_B_cNZdpEw14_1;
	wire w_dff_A_dDbcnEjY4_0;
	wire w_dff_A_JIpFM2TJ9_0;
	wire w_dff_A_UivY7Xvx2_0;
	wire w_dff_A_66jSKIFW0_0;
	wire w_dff_A_c7SNGAbI1_0;
	wire w_dff_A_Qn1WG3OA6_0;
	wire w_dff_A_UX79hV7d6_0;
	wire w_dff_A_3QMeQRYx4_0;
	wire w_dff_A_AkiNZV2m3_0;
	wire w_dff_A_4GLBo9I30_0;
	wire w_dff_A_C6znERXG9_0;
	wire w_dff_A_OTrDjAso9_0;
	wire w_dff_A_M9TN7u1o8_0;
	wire w_dff_A_SpNUAerN7_0;
	wire w_dff_A_Li1BxMt35_0;
	wire w_dff_A_hVARLdF90_0;
	wire w_dff_A_KOyFnJ6P3_0;
	wire w_dff_A_heyaKFTt6_0;
	wire w_dff_A_IfoL8a475_0;
	wire w_dff_A_qzKxelDI9_0;
	wire w_dff_A_wrjPjiGi8_0;
	wire w_dff_A_U06rrlK61_0;
	wire w_dff_A_F7GGot049_0;
	wire w_dff_A_H5a6kMnc7_0;
	wire w_dff_B_YN9xniCe7_1;
	wire w_dff_A_B3WQpwTl4_0;
	wire w_dff_A_0YemFUP72_0;
	wire w_dff_A_KRiL7IEK0_0;
	wire w_dff_A_GBy94EUE8_0;
	wire w_dff_A_zaQIbnIG7_0;
	wire w_dff_A_TRKK8lrZ0_0;
	wire w_dff_A_fHLYcBzl5_0;
	wire w_dff_A_jeGCbEct3_0;
	wire w_dff_A_xwjJ8Hl73_0;
	wire w_dff_A_l0S9gEMM7_0;
	wire w_dff_A_4eGXOV3D3_0;
	wire w_dff_A_A5zXeENM3_0;
	wire w_dff_A_pH1V3gBq1_0;
	wire w_dff_A_O5YybVCM4_0;
	wire w_dff_A_AYkCkQii3_0;
	wire w_dff_A_E8GAXqDH7_0;
	wire w_dff_A_6XWz6aFm8_0;
	wire w_dff_A_cC0z3G040_0;
	wire w_dff_A_5pWPVmoE9_0;
	wire w_dff_A_bWWMFQmV5_0;
	wire w_dff_A_vOuZa3lL8_0;
	wire w_dff_B_t7zGmDAA3_1;
	wire w_dff_A_2UkcZ4Vf5_0;
	wire w_dff_A_3tkynaLc6_0;
	wire w_dff_A_Bn60p0gt6_0;
	wire w_dff_A_LBSeKYrW7_0;
	wire w_dff_A_ktP54q1O9_0;
	wire w_dff_A_oKlHnjZ98_0;
	wire w_dff_A_5fnwKwEV0_0;
	wire w_dff_A_28cwp9BN3_0;
	wire w_dff_A_TZyYsELy1_0;
	wire w_dff_A_PdIZnOZs0_0;
	wire w_dff_A_qu5JsAQ68_0;
	wire w_dff_A_iIdUagJN7_0;
	wire w_dff_A_7DmEP9vG1_0;
	wire w_dff_A_QHMsashP2_0;
	wire w_dff_A_Z335YrJW3_0;
	wire w_dff_A_YzF7m0cY7_0;
	wire w_dff_A_Q4WRj3c35_0;
	wire w_dff_A_AoFzQpzy8_0;
	wire w_dff_B_0Uuq0fZ45_1;
	wire w_dff_A_2QI3qJVS2_0;
	wire w_dff_A_4TwJTyUU2_0;
	wire w_dff_A_zxDsxLGi9_0;
	wire w_dff_A_lCKEQrTs5_0;
	wire w_dff_A_D7FM4cfR4_0;
	wire w_dff_A_bh17kYxA5_0;
	wire w_dff_A_Y0CCq4A94_0;
	wire w_dff_A_NK5EfVlx2_0;
	wire w_dff_A_dLqodMmE1_0;
	wire w_dff_A_sagg0vuS4_0;
	wire w_dff_A_0LFcPuXD3_0;
	wire w_dff_A_cKBBEiH61_0;
	wire w_dff_A_NB7t1PsP8_0;
	wire w_dff_A_E3uuICfZ1_0;
	wire w_dff_A_AGyhUYPC7_0;
	wire w_dff_B_5lD7qqqs3_1;
	wire w_dff_A_AeuZPtDG8_0;
	wire w_dff_A_vrALIgrq6_0;
	wire w_dff_A_qH8KSHAO7_0;
	wire w_dff_A_ilmxlb7E5_0;
	wire w_dff_A_ke8BPedF2_0;
	wire w_dff_A_inHWBLTv5_0;
	wire w_dff_A_pccu4gh62_0;
	wire w_dff_A_IbKovbYn7_0;
	wire w_dff_A_fu6aqHvG5_0;
	wire w_dff_A_0EY2T5k61_0;
	wire w_dff_A_VWcmwtMh6_0;
	wire w_dff_A_m59HVWWN7_0;
	wire w_dff_B_Mhfr6fth5_1;
	wire w_dff_A_hyLvjgaq0_0;
	wire w_dff_A_fBk1XXtD8_0;
	wire w_dff_A_zOV19tar9_0;
	wire w_dff_A_cxfpP6D50_0;
	wire w_dff_A_e9mREQgc5_0;
	wire w_dff_A_dDUC5QbX1_0;
	wire w_dff_A_HeV4VCqy0_0;
	wire w_dff_A_lF7GCaFH7_0;
	wire w_dff_A_SZD2cvwN7_0;
	wire w_dff_A_ykQi1sID8_0;
	wire w_dff_A_bcA037ij8_0;
	wire w_dff_A_3cslWXqh6_1;
	wire w_dff_A_FWT5Eskw0_0;
	wire w_dff_A_100ztZiO3_0;
	wire w_dff_A_rKcGLXn78_0;
	wire w_dff_A_zmkCMecj4_0;
	wire w_dff_A_K0SsOrCV3_0;
	wire w_dff_A_dpwNAxEi6_0;
	wire w_dff_A_QvvnFDEe2_0;
	wire w_dff_B_GTzGY71r8_1;
	wire w_dff_A_JJnjh7cr5_1;
	wire w_dff_A_O3sEcoDA0_2;
	wire w_dff_A_129vUXF14_2;
	wire w_dff_A_58oNjSm74_0;
	wire w_dff_B_Xfkd7YaU7_2;
	wire w_dff_B_XYCnbEGk1_2;
	wire w_dff_B_ALEJVILM3_2;
	wire w_dff_B_hfXJN78t0_2;
	wire w_dff_B_IzVQw3Tg1_2;
	wire w_dff_B_86eJopzj1_2;
	wire w_dff_B_z0CKpGcV5_2;
	wire w_dff_B_VQGFMzn25_2;
	wire w_dff_B_pMLI55rQ1_2;
	wire w_dff_B_W07sIFpL5_2;
	wire w_dff_B_b4GITiFx9_2;
	wire w_dff_B_7vqDzFke6_2;
	wire w_dff_B_AFOV77Yp9_2;
	wire w_dff_B_LLMZEDco8_2;
	wire w_dff_B_IHcIAwtU1_2;
	wire w_dff_B_SX5AH0VY9_2;
	wire w_dff_B_skJe9Cz49_2;
	wire w_dff_B_GJkn4qjp1_2;
	wire w_dff_B_klc7ieDe0_2;
	wire w_dff_B_wwrrlaah7_2;
	wire w_dff_B_8JFqXxNQ4_2;
	wire w_dff_B_GXl8i9xh2_2;
	wire w_dff_B_1XnU7mGy5_2;
	wire w_dff_B_7yYzIjPa6_2;
	wire w_dff_B_E2v58dEj9_2;
	wire w_dff_B_GGvRfait7_2;
	wire w_dff_B_8421x3Dt3_2;
	wire w_dff_B_rIQAlWVs4_2;
	wire w_dff_B_FV3ApBIe9_2;
	wire w_dff_B_9QeiNDJJ8_2;
	wire w_dff_B_3Jm3eYIe2_2;
	wire w_dff_B_JaCMRJUa7_2;
	wire w_dff_B_7gh0oi4N6_2;
	wire w_dff_B_YrVzFK9A7_2;
	wire w_dff_B_LseRDJ8k7_2;
	wire w_dff_B_aYL9nx0e2_2;
	wire w_dff_B_77BJru3w1_2;
	wire w_dff_B_210xLPz89_2;
	wire w_dff_B_ai8Za3sR0_2;
	wire w_dff_B_7stG2Ylw7_2;
	wire w_dff_B_rD4XypI92_2;
	wire w_dff_B_9k8wHymZ8_2;
	wire w_dff_B_si7ZQzf03_2;
	wire w_dff_B_4MuhyZz56_2;
	wire w_dff_B_A3hoYYku9_2;
	wire w_dff_A_0WP8bNhx8_0;
	wire w_dff_B_ixj7yUiC0_1;
	wire w_dff_B_RdEFjcEE0_2;
	wire w_dff_B_MV4bqQJz9_2;
	wire w_dff_B_ClRaOHsw9_2;
	wire w_dff_B_UHV0fyxY3_2;
	wire w_dff_B_dygcDZ8r6_2;
	wire w_dff_B_6TgLpY779_2;
	wire w_dff_B_ir36mJq39_2;
	wire w_dff_B_8JZxrxqd7_2;
	wire w_dff_B_qmho1tvv5_2;
	wire w_dff_B_eA36qhs15_2;
	wire w_dff_B_vKHAUT8B3_2;
	wire w_dff_B_NHDgziGL8_2;
	wire w_dff_B_U12dkmG22_2;
	wire w_dff_B_qYCAoU1x6_2;
	wire w_dff_B_P1FziXA14_2;
	wire w_dff_B_KtVatRyz5_2;
	wire w_dff_B_manjh1NZ5_2;
	wire w_dff_B_QTwQ1JIM6_2;
	wire w_dff_B_9F3Cheqa6_2;
	wire w_dff_B_wYumgaWL6_2;
	wire w_dff_B_pCSDMmHc2_2;
	wire w_dff_B_WLlRa5yB2_2;
	wire w_dff_B_RlF98wIe1_2;
	wire w_dff_B_gSOEA2j56_2;
	wire w_dff_B_VXDqMmki5_2;
	wire w_dff_B_n8gUi5QA1_2;
	wire w_dff_B_PX2sR0uv3_2;
	wire w_dff_B_ZQyEPytw4_2;
	wire w_dff_B_9bhBoudj2_2;
	wire w_dff_B_CEJjXlkA2_2;
	wire w_dff_B_irtCtgqt4_2;
	wire w_dff_B_NtCTb9NO3_2;
	wire w_dff_B_QAMRhUhQ1_2;
	wire w_dff_B_L3KJJBar3_2;
	wire w_dff_B_X3hmDc9U0_2;
	wire w_dff_B_t8a7mpJc1_2;
	wire w_dff_B_eakJ78K88_2;
	wire w_dff_B_7Stnel8r1_2;
	wire w_dff_B_qFncmWYE3_2;
	wire w_dff_B_NK1cGy002_2;
	wire w_dff_B_0RTT3rWU7_2;
	wire w_dff_A_LiLLaKQ70_1;
	wire w_dff_A_JVFZYS5k2_0;
	wire w_dff_A_ThE4032i7_0;
	wire w_dff_A_b8dyL3Gc7_0;
	wire w_dff_A_MFmMa0Sk5_0;
	wire w_dff_A_hNVLQOt59_0;
	wire w_dff_A_aNJzPPnh5_0;
	wire w_dff_A_sTza9uYR8_0;
	wire w_dff_A_ucZrvFil5_0;
	wire w_dff_A_rujyZHXO7_0;
	wire w_dff_A_BTuUOtKP4_0;
	wire w_dff_A_oicvysoX1_0;
	wire w_dff_A_tmZXjUZJ1_0;
	wire w_dff_A_OP2JCiGM7_0;
	wire w_dff_A_X51ycMFW3_0;
	wire w_dff_A_ulWJkAd52_0;
	wire w_dff_A_wBkthbbs3_0;
	wire w_dff_A_efQbvt229_0;
	wire w_dff_A_QeXAeT9f6_0;
	wire w_dff_A_s7D7sebC2_0;
	wire w_dff_A_x885c7Ue6_0;
	wire w_dff_A_wiavjYbC8_0;
	wire w_dff_A_qLhJBFLE0_0;
	wire w_dff_A_1kIhnF6k7_0;
	wire w_dff_A_Z84DsC3x1_0;
	wire w_dff_A_O8e5PD9S4_0;
	wire w_dff_A_mxB2yEn90_0;
	wire w_dff_A_VLDufczS1_0;
	wire w_dff_A_tyScGpDV5_0;
	wire w_dff_A_CrJ0yvYZ5_0;
	wire w_dff_A_RrkunfDu4_0;
	wire w_dff_A_BZnmWBMG8_0;
	wire w_dff_A_JpAY9JLX4_0;
	wire w_dff_A_NN1WPiiH7_0;
	wire w_dff_A_ElRliAgJ8_0;
	wire w_dff_A_DqnCeYFm4_0;
	wire w_dff_A_Zrw86vAk2_0;
	wire w_dff_A_dfoK9Vu36_0;
	wire w_dff_A_PXYu4tFF2_0;
	wire w_dff_A_rNhfqppf1_1;
	wire w_dff_A_ERUtKZw50_2;
	wire w_dff_B_pFzgrlqQ6_1;
	wire w_dff_B_aqLqSVbb5_2;
	wire w_dff_B_8TtlUCFZ6_2;
	wire w_dff_B_fGoWAijM3_2;
	wire w_dff_B_LX6g5d3q0_2;
	wire w_dff_B_OxgyoqTX1_2;
	wire w_dff_B_ePUgQZSz9_2;
	wire w_dff_B_855WPIpP8_2;
	wire w_dff_B_1SLzG1sJ8_2;
	wire w_dff_B_ZONFmFUc2_2;
	wire w_dff_B_zgrMX4vu2_2;
	wire w_dff_B_CWoryAm58_2;
	wire w_dff_B_8PI4HxTW1_2;
	wire w_dff_B_W565hlja3_2;
	wire w_dff_B_goC2GtdM8_2;
	wire w_dff_B_zglewjTh2_2;
	wire w_dff_B_NCfsaHxY3_2;
	wire w_dff_B_izzFwD9P7_2;
	wire w_dff_B_jcVvnAzP3_2;
	wire w_dff_B_V8ljW9QM2_2;
	wire w_dff_B_RiDZEjDY7_2;
	wire w_dff_B_PiUefMaQ9_2;
	wire w_dff_B_l17r3wle0_2;
	wire w_dff_B_pjpfPEhq9_2;
	wire w_dff_B_DVx2s3wq5_2;
	wire w_dff_B_73GQfmpV4_2;
	wire w_dff_B_iiZJ8oQK7_2;
	wire w_dff_B_ETLGqHFC0_2;
	wire w_dff_B_wuc06J5x0_2;
	wire w_dff_B_2mWbSJ3u6_2;
	wire w_dff_B_UVLb67d54_2;
	wire w_dff_B_dXYrXhlm3_2;
	wire w_dff_B_sNZ6qBcz6_2;
	wire w_dff_B_GSt3l0oj2_2;
	wire w_dff_B_CGzaqclw9_2;
	wire w_dff_B_lsaBQh7J8_2;
	wire w_dff_B_YFGLmNff5_1;
	wire w_dff_B_qjeV4zON2_2;
	wire w_dff_B_8R7Ti3qY2_2;
	wire w_dff_B_84YqnIUj2_2;
	wire w_dff_B_IJnCaoWh3_2;
	wire w_dff_B_0OEM80xx5_2;
	wire w_dff_B_uV6ZS0iu8_2;
	wire w_dff_B_6Y0S37xe5_2;
	wire w_dff_B_lHV9p9xl7_2;
	wire w_dff_B_8REZEnvQ1_2;
	wire w_dff_B_VqROLeH34_2;
	wire w_dff_B_ogbzXqZ74_2;
	wire w_dff_B_t8uPvq429_2;
	wire w_dff_B_JaALiz3y5_2;
	wire w_dff_B_nRCTL3CB6_2;
	wire w_dff_B_rZWLath03_2;
	wire w_dff_B_8235HZRe8_2;
	wire w_dff_B_vj6GeHQl1_2;
	wire w_dff_B_wWrx1rJ38_2;
	wire w_dff_B_fYft93dk1_2;
	wire w_dff_B_3JYrxhaL4_2;
	wire w_dff_B_wNm6FKIX1_2;
	wire w_dff_B_2itOObFF4_2;
	wire w_dff_B_Rzkg6iNm6_2;
	wire w_dff_B_MkZbSH8v5_2;
	wire w_dff_B_LwCJR8VV8_2;
	wire w_dff_B_oPY21CCQ4_2;
	wire w_dff_B_vMqCSAr18_2;
	wire w_dff_B_vkit0yNc5_2;
	wire w_dff_B_LoFVokDw9_2;
	wire w_dff_B_JaDhI1AO8_2;
	wire w_dff_B_ZYWG448Y6_2;
	wire w_dff_B_XMyO4VcL9_2;
	wire w_dff_B_p7A5tY8K4_1;
	wire w_dff_B_SWE7pXwo9_2;
	wire w_dff_B_lOav3PfN0_2;
	wire w_dff_B_wFYf2lav8_2;
	wire w_dff_B_HZIKFsvb9_2;
	wire w_dff_B_R488Rsjb9_2;
	wire w_dff_B_098UAozT5_2;
	wire w_dff_B_iFUaAVA13_2;
	wire w_dff_B_IWrhjz9Z0_2;
	wire w_dff_B_4J5QOlcx4_2;
	wire w_dff_B_xfOBvoTR5_2;
	wire w_dff_B_03J3pO6K2_2;
	wire w_dff_B_aZn31KFm0_2;
	wire w_dff_B_226Xofee5_2;
	wire w_dff_B_lhKvZDVA2_2;
	wire w_dff_B_itQyYcEO2_2;
	wire w_dff_B_v2OoYA8f8_2;
	wire w_dff_B_w06hzSZz7_2;
	wire w_dff_B_TVmd71Bt5_2;
	wire w_dff_B_gAUP2gyM6_2;
	wire w_dff_B_pGZDE7MI4_2;
	wire w_dff_B_FF3Y9FHH8_2;
	wire w_dff_B_TlxNAIKP7_2;
	wire w_dff_B_uSV59Dl34_2;
	wire w_dff_B_r445SAU90_2;
	wire w_dff_B_pWXeHk9R5_2;
	wire w_dff_B_sVujVXx70_2;
	wire w_dff_B_IvwcZuZ52_2;
	wire w_dff_B_IqjvnNs23_2;
	wire w_dff_B_A0EP2u038_2;
	wire w_dff_B_LdbHXJz70_1;
	wire w_dff_B_remLdU3W7_2;
	wire w_dff_B_nSCTjnSp5_2;
	wire w_dff_B_EmZUjoei5_2;
	wire w_dff_B_kzvdLuxQ4_2;
	wire w_dff_B_j0nqz0qI3_2;
	wire w_dff_B_UF4stipx1_2;
	wire w_dff_B_Ong0mR9n3_2;
	wire w_dff_B_BoG9dJsj3_2;
	wire w_dff_B_4l8CMNvt4_2;
	wire w_dff_B_0AtmG2Cn7_2;
	wire w_dff_B_vaaTdudL8_2;
	wire w_dff_B_fJqk2wzJ0_2;
	wire w_dff_B_FPlSDfho2_2;
	wire w_dff_B_FukND1Vq8_2;
	wire w_dff_B_g0Om3uaU4_2;
	wire w_dff_B_Pj0dZwwN3_2;
	wire w_dff_B_Bh7jb3Mx6_2;
	wire w_dff_B_ffTQWIFS5_2;
	wire w_dff_B_wLMNGDU23_2;
	wire w_dff_B_A3BrkMmV3_2;
	wire w_dff_B_gSujsVYH1_2;
	wire w_dff_B_qErqbt8q0_2;
	wire w_dff_B_fOtmj0Vl2_2;
	wire w_dff_B_G3PK9Dmz9_2;
	wire w_dff_B_YZsqRtp03_2;
	wire w_dff_B_ahnDQaUE2_2;
	wire w_dff_B_VdB4vGKp5_1;
	wire w_dff_B_2VwStOel9_2;
	wire w_dff_B_kLxdcguU7_2;
	wire w_dff_B_7jOyGxjd9_2;
	wire w_dff_B_iAYneITv0_2;
	wire w_dff_B_7W1gMF8E6_2;
	wire w_dff_B_4heQCxFT6_2;
	wire w_dff_B_BmKSXrJd4_2;
	wire w_dff_B_YIhP0J3W2_2;
	wire w_dff_B_DxH8y57k0_2;
	wire w_dff_B_DxkGXL4K2_2;
	wire w_dff_B_LG1DRUM75_2;
	wire w_dff_B_gwkAKuOX3_2;
	wire w_dff_B_HZIXzl9R1_2;
	wire w_dff_B_t0YiUaOj3_2;
	wire w_dff_B_XaEkSQOJ5_2;
	wire w_dff_B_Ieuytx2k1_2;
	wire w_dff_B_rVH2xRnM3_2;
	wire w_dff_B_MNSiRIMK9_2;
	wire w_dff_B_gIFGXc919_2;
	wire w_dff_B_CrCxR1cm2_2;
	wire w_dff_B_gQ6syMS02_2;
	wire w_dff_B_B1MHIwkE4_2;
	wire w_dff_B_oai99Er00_2;
	wire w_dff_B_Ha01Stdo7_1;
	wire w_dff_B_kPzXdT731_2;
	wire w_dff_B_rtyGdkVm1_2;
	wire w_dff_B_vhAZV4Tc4_2;
	wire w_dff_B_gWd43pn36_2;
	wire w_dff_B_ZdFhonGr4_2;
	wire w_dff_B_Rtwqnh0h5_2;
	wire w_dff_B_HNe5PlZm0_2;
	wire w_dff_B_3SxQLx4g3_2;
	wire w_dff_B_okHSrSDq9_2;
	wire w_dff_B_3B9sHaTO1_2;
	wire w_dff_B_jpsQrg4H5_2;
	wire w_dff_B_DsHnBPqt4_2;
	wire w_dff_B_jZdjHIib2_2;
	wire w_dff_B_DBAuNXme7_2;
	wire w_dff_B_Z1xPljwx3_2;
	wire w_dff_B_a779KKf65_2;
	wire w_dff_B_t1I5GBDE3_2;
	wire w_dff_B_pLjYX2P31_2;
	wire w_dff_B_Jv3A2qaZ9_2;
	wire w_dff_B_rbZL3TVO2_2;
	wire w_dff_B_QhBkAYhP6_1;
	wire w_dff_B_3yKfvuf39_2;
	wire w_dff_B_QAyCvtyq7_2;
	wire w_dff_B_Ob3yL81s1_2;
	wire w_dff_B_SW0GfjWC1_2;
	wire w_dff_B_pdfeUBWc5_2;
	wire w_dff_B_bzFlRNgb6_2;
	wire w_dff_B_reD8dfdd1_2;
	wire w_dff_B_HlnvGXCL2_2;
	wire w_dff_B_9R9D6Qrj3_2;
	wire w_dff_B_685BWqiP9_2;
	wire w_dff_B_OjdGeNKJ3_2;
	wire w_dff_B_ryEQoQyp0_2;
	wire w_dff_B_snitgZz50_2;
	wire w_dff_B_2EI7hVaw4_2;
	wire w_dff_B_1Huhmroh3_2;
	wire w_dff_B_OnVhSGaU0_2;
	wire w_dff_B_Flxa6Eko8_2;
	wire w_dff_B_6Fhf9Eju8_1;
	wire w_dff_B_7OpAxnXt7_2;
	wire w_dff_B_j0cy7ffD7_2;
	wire w_dff_B_Peeqc6VE0_2;
	wire w_dff_B_3ekBNrqu2_2;
	wire w_dff_B_Tvh1sZvk8_2;
	wire w_dff_B_iKrspdTh0_2;
	wire w_dff_B_NT2WauMy1_2;
	wire w_dff_B_OW93GX1A8_2;
	wire w_dff_B_wPlQyK8K5_2;
	wire w_dff_B_3gwdVvUv7_2;
	wire w_dff_B_QcrKqKi74_2;
	wire w_dff_B_7XhZKsfy9_2;
	wire w_dff_B_7t7VuDNg2_2;
	wire w_dff_B_5WzUuFtq7_2;
	wire w_dff_B_ncfFgBcp6_1;
	wire w_dff_B_1SQv2chZ3_2;
	wire w_dff_B_kaNBOWuF6_2;
	wire w_dff_B_pMy8k2Y10_2;
	wire w_dff_B_CPnvODoO8_2;
	wire w_dff_B_BsS1fQvf8_2;
	wire w_dff_B_4KO8A3aG2_2;
	wire w_dff_B_WoJonN7K9_2;
	wire w_dff_B_cFRAFIlK7_2;
	wire w_dff_B_sE7s3cCi0_2;
	wire w_dff_B_2BHgDr6f3_2;
	wire w_dff_B_Hwp7sJGy6_2;
	wire w_dff_B_Rn758qRw2_1;
	wire w_dff_B_245dB2Vj1_2;
	wire w_dff_B_GxmnUU2i9_2;
	wire w_dff_B_qMjk9fbg4_2;
	wire w_dff_B_HfWphmhP3_2;
	wire w_dff_B_QZE1CIaw1_2;
	wire w_dff_B_ht3rygSr0_2;
	wire w_dff_B_E9bULjDw7_2;
	wire w_dff_B_U2AtfufT8_2;
	wire w_dff_B_6BySlTG00_1;
	wire w_dff_B_jyMdLAoA5_1;
	wire w_dff_B_55AhhSfT5_2;
	wire w_dff_B_AR0OBn1x1_2;
	wire w_dff_B_SKN6sspX6_2;
	wire w_dff_B_uXlhIgzZ4_2;
	wire w_dff_A_bcg8oVQH4_1;
	wire w_dff_A_1G0AuNFk3_0;
	wire w_dff_A_avonoj9j1_0;
	wire w_dff_A_ixNCcfTv9_1;
	wire w_dff_A_ir0jkoTy5_2;
	wire w_dff_A_srC73IwU0_2;
	wire w_dff_B_iWR1jGX20_0;
	wire w_dff_A_vNJLJ28L9_1;
	wire w_dff_A_nsNq7sN28_1;
	wire w_dff_B_YGmA32BL2_1;
	wire w_dff_B_Xe2jUCZn7_1;
	wire w_dff_B_VrfINGLF2_2;
	wire w_dff_B_XRfA1XNS1_2;
	wire w_dff_B_OcDoaZCJ1_2;
	wire w_dff_B_TgjGHPTz1_2;
	wire w_dff_B_uirphLHQ6_2;
	wire w_dff_B_pXrGjQ6a9_2;
	wire w_dff_B_z75aXurF5_2;
	wire w_dff_B_gMdAcu1U7_2;
	wire w_dff_B_SAinsTPC1_2;
	wire w_dff_B_Vz6fifrE0_2;
	wire w_dff_B_G7rr8G725_2;
	wire w_dff_B_I2mQM6LX9_2;
	wire w_dff_B_QUJcTRdT2_2;
	wire w_dff_B_2BGDN8B65_2;
	wire w_dff_B_hBQWltrx1_2;
	wire w_dff_B_TdXrTcUA7_2;
	wire w_dff_B_IpKsEiml0_2;
	wire w_dff_B_VgYxqRs84_2;
	wire w_dff_B_Jr4pzSBm6_2;
	wire w_dff_B_9v4AewAA1_2;
	wire w_dff_B_sUyJAQLP2_2;
	wire w_dff_B_iIaN59k97_2;
	wire w_dff_B_7STjTvPY6_2;
	wire w_dff_B_SrNRAmR12_2;
	wire w_dff_B_O8jpz1An2_2;
	wire w_dff_B_7T1mB0cm9_2;
	wire w_dff_B_DmaFqNAH0_2;
	wire w_dff_B_WobrmUQu2_2;
	wire w_dff_B_D2JmnkdL1_2;
	wire w_dff_B_tpgvJ9CA8_2;
	wire w_dff_B_BSOTueR98_2;
	wire w_dff_B_VQH5x6mD1_2;
	wire w_dff_B_EbjNuSer1_2;
	wire w_dff_B_ka8jStj19_2;
	wire w_dff_B_kNTlWiqX7_2;
	wire w_dff_B_afMCcITk5_2;
	wire w_dff_B_bpOdG4iR4_2;
	wire w_dff_B_EH4SD5so8_2;
	wire w_dff_B_ebJun9CI7_2;
	wire w_dff_B_Rk1dtwek0_2;
	wire w_dff_B_71HUwSnK0_2;
	wire w_dff_B_dZZyLqHf4_2;
	wire w_dff_B_QSRCM4is5_2;
	wire w_dff_B_yiuIGVGX8_2;
	wire w_dff_B_fZaMNZMF5_2;
	wire w_dff_B_la2T5edW5_2;
	wire w_dff_B_GIJup5jm6_2;
	wire w_dff_B_KiUGehzL6_1;
	wire w_dff_B_rewq4jsN8_2;
	wire w_dff_B_FsJAHL7T8_2;
	wire w_dff_B_DxbEk9Do7_2;
	wire w_dff_B_qk9p5GUp6_2;
	wire w_dff_B_HZN6197g9_2;
	wire w_dff_B_ItHsGKyE2_2;
	wire w_dff_B_hRMkurKu0_2;
	wire w_dff_B_10g616Fd4_2;
	wire w_dff_B_AjD8ZvoK2_2;
	wire w_dff_B_EsPpHUED9_2;
	wire w_dff_B_z4QvrVIP4_2;
	wire w_dff_B_EdUwjeuf8_2;
	wire w_dff_B_nYnp5rFQ8_2;
	wire w_dff_B_aRSQi7JQ7_2;
	wire w_dff_B_5C1Bkj3z8_2;
	wire w_dff_B_FNBeGY117_2;
	wire w_dff_B_TQGFwaNc2_2;
	wire w_dff_B_nMaRYxcD2_2;
	wire w_dff_B_EqTgjE9Q8_2;
	wire w_dff_B_wSvHJhfE2_2;
	wire w_dff_B_Cm294iTF6_2;
	wire w_dff_B_xmhdO6RH9_2;
	wire w_dff_B_xtH2xk4b5_2;
	wire w_dff_B_9c9MD8zi2_2;
	wire w_dff_B_yRBYk8Oe2_2;
	wire w_dff_B_MGHYPV087_2;
	wire w_dff_B_yE4eQ1Uh3_2;
	wire w_dff_B_TqRH4DC72_2;
	wire w_dff_B_QTy9EYpY8_2;
	wire w_dff_B_LR2IAJHR2_2;
	wire w_dff_B_u2lXHmpz3_2;
	wire w_dff_B_9sNQnnWr0_2;
	wire w_dff_B_JvxBIJkd5_2;
	wire w_dff_B_bdNK3aFA1_2;
	wire w_dff_B_OXb66QLL0_2;
	wire w_dff_B_ui7AadZK3_2;
	wire w_dff_B_acAocIjr2_2;
	wire w_dff_B_uObjiOEf1_2;
	wire w_dff_B_RP3MClyb5_2;
	wire w_dff_B_6ZcaJYfa8_2;
	wire w_dff_B_hSsYxRe46_2;
	wire w_dff_B_LLAZKhDn3_2;
	wire w_dff_B_4OqqlQj08_2;
	wire w_dff_B_877gKBVH1_1;
	wire w_dff_B_5jft2Vwy6_2;
	wire w_dff_B_ZN8TJwuQ8_2;
	wire w_dff_B_zTZjp51P1_2;
	wire w_dff_B_hUvwZgQR1_2;
	wire w_dff_B_FVNmkt943_2;
	wire w_dff_B_sXLylmgx7_2;
	wire w_dff_B_WANgA7vs3_2;
	wire w_dff_B_fCC3zs2y6_2;
	wire w_dff_B_x2qKhbFB6_2;
	wire w_dff_B_GUNSKsCY0_2;
	wire w_dff_B_iQmc28Lc0_2;
	wire w_dff_B_uY4a52hs4_2;
	wire w_dff_B_3iCrlnnm9_2;
	wire w_dff_B_LJLGwmyK7_2;
	wire w_dff_B_NV4ochvg1_2;
	wire w_dff_B_cTAZdZuN9_2;
	wire w_dff_B_PrHX0WOD4_2;
	wire w_dff_B_rxkKwHsc1_2;
	wire w_dff_B_8rmTXVCC1_2;
	wire w_dff_B_6nCHpHQ83_2;
	wire w_dff_B_v9bxAY7j3_2;
	wire w_dff_B_dkFlagy72_2;
	wire w_dff_B_aXPHQdB68_2;
	wire w_dff_B_dnoxVV8M8_2;
	wire w_dff_B_siVuMN1S1_2;
	wire w_dff_B_OvKBIR2v5_2;
	wire w_dff_B_VGwR5a5V8_2;
	wire w_dff_B_PfZATf5Z7_2;
	wire w_dff_B_JO5e3owO8_2;
	wire w_dff_B_QOIGMBCv0_2;
	wire w_dff_B_cOEeJdOO5_2;
	wire w_dff_B_bLVjfL3e5_2;
	wire w_dff_B_RaWgKTIy8_2;
	wire w_dff_B_l22DOOKi2_2;
	wire w_dff_B_0GbXCiTa4_2;
	wire w_dff_B_ET3KHaJ89_2;
	wire w_dff_B_zFBisT5P4_2;
	wire w_dff_B_lwCdysTz7_2;
	wire w_dff_B_vxmO1t5E1_1;
	wire w_dff_B_KgNEIDdg7_2;
	wire w_dff_B_DyOciAqY6_2;
	wire w_dff_B_AO610JJm0_2;
	wire w_dff_B_4Bx7eUcR0_2;
	wire w_dff_B_Dce8WUZR6_2;
	wire w_dff_B_NTm7gPf28_2;
	wire w_dff_B_fU6SomYh0_2;
	wire w_dff_B_OdaSii8Z4_2;
	wire w_dff_B_1niVhtcy2_2;
	wire w_dff_B_GstPYLjk1_2;
	wire w_dff_B_T8Spe6jd9_2;
	wire w_dff_B_lPRBVp1C3_2;
	wire w_dff_B_pwA5AzaO2_2;
	wire w_dff_B_BI5zecxF9_2;
	wire w_dff_B_Rf3UPpIJ2_2;
	wire w_dff_B_NJz4azqW1_2;
	wire w_dff_B_NfQ241217_2;
	wire w_dff_B_awfMdEK42_2;
	wire w_dff_B_0PeRm2hj5_2;
	wire w_dff_B_Qmg3mdtc5_2;
	wire w_dff_B_wG7tUDtG6_2;
	wire w_dff_B_oB2hDlLM6_2;
	wire w_dff_B_P7fByLw52_2;
	wire w_dff_B_4lr70A8b7_2;
	wire w_dff_B_dhwmhWxF1_2;
	wire w_dff_B_jl7oPzYT6_2;
	wire w_dff_B_2extvQgJ6_2;
	wire w_dff_B_AuJWx6rf1_2;
	wire w_dff_B_tLaxWX5T1_2;
	wire w_dff_B_bBV8Rk6E4_2;
	wire w_dff_B_HpW7zvZH0_2;
	wire w_dff_B_EipvCePu1_2;
	wire w_dff_B_l7FlFbyc1_2;
	wire w_dff_B_X2kT5Udq3_2;
	wire w_dff_B_6Gtr6lbk5_2;
	wire w_dff_B_pkXP9ILj6_1;
	wire w_dff_B_7T2LisQI8_2;
	wire w_dff_B_83iD7Qxu4_2;
	wire w_dff_B_4jDij4Gy4_2;
	wire w_dff_B_7JujXeVW3_2;
	wire w_dff_B_Y591g1cA7_2;
	wire w_dff_B_OPsknhG53_2;
	wire w_dff_B_Oet3mOMN6_2;
	wire w_dff_B_dzqTfCik5_2;
	wire w_dff_B_5eDO5SmG6_2;
	wire w_dff_B_jPoroVdG8_2;
	wire w_dff_B_iIynPmaY5_2;
	wire w_dff_B_4aihdRmi2_2;
	wire w_dff_B_O3vtcIue1_2;
	wire w_dff_B_GinTlZ4E5_2;
	wire w_dff_B_8hOLKX822_2;
	wire w_dff_B_D4wy2Okt0_2;
	wire w_dff_B_zogtRBeB2_2;
	wire w_dff_B_kcYT7JJE9_2;
	wire w_dff_B_h74PmwWU9_2;
	wire w_dff_B_fxamom8A5_2;
	wire w_dff_B_7plIDstX4_2;
	wire w_dff_B_zwt3KlqH6_2;
	wire w_dff_B_F0e8ypID5_2;
	wire w_dff_B_INyCAKn87_2;
	wire w_dff_B_bG8EAJce6_2;
	wire w_dff_B_zqeQsN1F0_2;
	wire w_dff_B_vGlcpdYO4_2;
	wire w_dff_B_EGrDx8bY8_2;
	wire w_dff_B_M3k35jO77_2;
	wire w_dff_B_V8sBfmYO8_2;
	wire w_dff_B_HMm1T04d9_2;
	wire w_dff_B_pf4x7cqt6_2;
	wire w_dff_B_BJRhwV3R5_1;
	wire w_dff_B_BQnm9l3F7_2;
	wire w_dff_B_0fs6jalb2_2;
	wire w_dff_B_tWegmQyn5_2;
	wire w_dff_B_c8BeTa936_2;
	wire w_dff_B_UT333E6g5_2;
	wire w_dff_B_7aK2YLmc4_2;
	wire w_dff_B_YSRAgxvZ2_2;
	wire w_dff_B_hZO859T94_2;
	wire w_dff_B_Rjud5mMf3_2;
	wire w_dff_B_jKvJFixD2_2;
	wire w_dff_B_o2SywZtH9_2;
	wire w_dff_B_3K0e5WII4_2;
	wire w_dff_B_FM3HVfhi8_2;
	wire w_dff_B_zWDUI0Me3_2;
	wire w_dff_B_avZ27p1p6_2;
	wire w_dff_B_NEm5x4Wc3_2;
	wire w_dff_B_C5PNdhBg2_2;
	wire w_dff_B_VKCtOqN43_2;
	wire w_dff_B_lUwmlAeX7_2;
	wire w_dff_B_Fbiezlze8_2;
	wire w_dff_B_nufP5pcR3_2;
	wire w_dff_B_uakW9DrU9_2;
	wire w_dff_B_p9UZvedm1_2;
	wire w_dff_B_eucCY8Co8_2;
	wire w_dff_B_HTzDBLQN1_2;
	wire w_dff_B_LJb31AHq0_2;
	wire w_dff_B_DzISyPcN3_2;
	wire w_dff_B_ovFfKiA53_2;
	wire w_dff_B_LjFoFNip1_2;
	wire w_dff_B_yk77LfyS1_1;
	wire w_dff_B_vX247xk67_2;
	wire w_dff_B_sokSTcOG0_2;
	wire w_dff_B_Au02DbKr4_2;
	wire w_dff_B_xAKdDGgk1_2;
	wire w_dff_B_CKOuBb2H3_2;
	wire w_dff_B_J4gbxKKz7_2;
	wire w_dff_B_HmJft7fe1_2;
	wire w_dff_B_0o4AMnh69_2;
	wire w_dff_B_uotRdzng1_2;
	wire w_dff_B_7k9pINyR9_2;
	wire w_dff_B_yzGc4yFe4_2;
	wire w_dff_B_nNtGhztX6_2;
	wire w_dff_B_C3pVjf5o5_2;
	wire w_dff_B_SiadrbWM7_2;
	wire w_dff_B_VByJf3059_2;
	wire w_dff_B_yH2hGQCi7_2;
	wire w_dff_B_PHYtLVdL3_2;
	wire w_dff_B_aWFLV4zV8_2;
	wire w_dff_B_VreCK2Zn9_2;
	wire w_dff_B_vhbocJP33_2;
	wire w_dff_B_b36eqfI50_2;
	wire w_dff_B_tsznxY1O7_2;
	wire w_dff_B_cqMgiee46_2;
	wire w_dff_B_euIm4nAl6_2;
	wire w_dff_B_tVGUx8Nc5_2;
	wire w_dff_B_KPzLWWr84_2;
	wire w_dff_B_sfAyzdid9_1;
	wire w_dff_B_tBziSE9s9_2;
	wire w_dff_B_E3WiGHgg3_2;
	wire w_dff_B_3odx0bRh1_2;
	wire w_dff_B_5xvwF1AJ0_2;
	wire w_dff_B_PXwsmNAp1_2;
	wire w_dff_B_EPR7Gnig5_2;
	wire w_dff_B_BdDlnazm5_2;
	wire w_dff_B_MNrxvM1N4_2;
	wire w_dff_B_FktG2pVH6_2;
	wire w_dff_B_QO1tV3ur3_2;
	wire w_dff_B_cHrW7Fv70_2;
	wire w_dff_B_WpCoG4pw2_2;
	wire w_dff_B_hRKP4OTP6_2;
	wire w_dff_B_aMKpDt5s2_2;
	wire w_dff_B_SBAQuFqy8_2;
	wire w_dff_B_KfWZey4c7_2;
	wire w_dff_B_1sSUDwjL5_2;
	wire w_dff_B_kRM71OWs1_2;
	wire w_dff_B_L7Re6p556_2;
	wire w_dff_B_RLZ1sl8P5_2;
	wire w_dff_B_j7Hhtgq99_2;
	wire w_dff_B_fS3wTcsS6_2;
	wire w_dff_B_SXqyNsLN2_2;
	wire w_dff_B_P8KsRJix4_1;
	wire w_dff_B_ivtSATeg6_2;
	wire w_dff_B_bSck8pg16_2;
	wire w_dff_B_PPlnoxLt1_2;
	wire w_dff_B_gVRRjAkj5_2;
	wire w_dff_B_yXvRq2zm9_2;
	wire w_dff_B_udWu3Xpw1_2;
	wire w_dff_B_HPD2iSFG7_2;
	wire w_dff_B_3wR3YO3U4_2;
	wire w_dff_B_tjZYPU2Z4_2;
	wire w_dff_B_WQXKZcJ65_2;
	wire w_dff_B_cbevVVP57_2;
	wire w_dff_B_q1NKHPOc8_2;
	wire w_dff_B_DAKdFrKw1_2;
	wire w_dff_B_kSqrz5ax3_2;
	wire w_dff_B_jT95uDpE4_2;
	wire w_dff_B_tWTx0CE57_2;
	wire w_dff_B_OTXhif4F3_2;
	wire w_dff_B_2CSl2zK59_2;
	wire w_dff_B_OMGyWvRk1_2;
	wire w_dff_B_oiv1Ej0a7_2;
	wire w_dff_B_dq2zZtCe8_1;
	wire w_dff_B_xM74ADJ29_2;
	wire w_dff_B_3eiP6WyV9_2;
	wire w_dff_B_wwcWKxWg0_2;
	wire w_dff_B_6JXvXZL78_2;
	wire w_dff_B_nhQwA36v6_2;
	wire w_dff_B_tKbfhqnV1_2;
	wire w_dff_B_u3mx4Fm42_2;
	wire w_dff_B_AHTXeoLm0_2;
	wire w_dff_B_AC2GPz4U2_2;
	wire w_dff_B_1m42DFdN0_2;
	wire w_dff_B_M8rU20jP3_2;
	wire w_dff_B_D2qZE4Ho3_2;
	wire w_dff_B_0hHmznac2_2;
	wire w_dff_B_qIOTDY6n4_2;
	wire w_dff_B_EBfLEmbc8_2;
	wire w_dff_B_VzlPzLz94_2;
	wire w_dff_B_eVcoFSmM5_2;
	wire w_dff_B_YZOkLI4o6_1;
	wire w_dff_B_xuWjU0ax0_2;
	wire w_dff_B_udVe7QZu4_2;
	wire w_dff_B_Klc1olYN9_2;
	wire w_dff_B_7yt3SJo93_2;
	wire w_dff_B_X0RUb1Vg3_2;
	wire w_dff_B_khSBdDmA2_2;
	wire w_dff_B_gmVkOzqQ9_2;
	wire w_dff_B_PJFu1ViR8_2;
	wire w_dff_B_HwKhKumH7_2;
	wire w_dff_B_OVKJk7MB5_2;
	wire w_dff_B_kFgG7cQJ0_2;
	wire w_dff_B_CgvGs1og2_2;
	wire w_dff_B_ZT1o73KG3_2;
	wire w_dff_B_Pwl0RWjL6_2;
	wire w_dff_B_emUlAaqO8_1;
	wire w_dff_B_VhQFQa4L7_2;
	wire w_dff_B_mI8afoDC6_2;
	wire w_dff_B_lD2EsLUg4_2;
	wire w_dff_B_hAofEnzJ7_2;
	wire w_dff_B_2jUyhUpQ3_2;
	wire w_dff_B_mEOz2IDu0_2;
	wire w_dff_B_21cavMbj0_2;
	wire w_dff_B_tOik5Oue3_2;
	wire w_dff_B_lfRjL2Zh3_2;
	wire w_dff_B_Eevn5yIO0_2;
	wire w_dff_B_HK1uxouA2_2;
	wire w_dff_B_CzRkLVTi9_1;
	wire w_dff_B_7w8WipcE5_2;
	wire w_dff_B_dyrzvjCK6_2;
	wire w_dff_B_c4k9w88Y8_2;
	wire w_dff_B_KUDyAe7b5_2;
	wire w_dff_B_edYnSJi39_2;
	wire w_dff_B_Z1h68yYY9_2;
	wire w_dff_B_1YazrMbv9_2;
	wire w_dff_B_eHQGTVDo8_2;
	wire w_dff_B_7gwb7JRl2_1;
	wire w_dff_B_CraBrRg64_0;
	wire w_dff_B_BzYavjYu2_2;
	wire w_dff_B_uynEtcs31_2;
	wire w_dff_B_VjiOsel71_2;
	wire w_dff_B_LYuZZ2cD3_2;
	wire w_dff_B_owZoKCNi7_1;
	wire w_dff_A_HULXV26v8_0;
	wire w_dff_A_g6UKxOzF8_0;
	wire w_dff_A_5rzIXust7_1;
	wire w_dff_B_xI4KtHss7_1;
	wire w_dff_B_UZHohOxC7_2;
	wire w_dff_B_TPMAldQH1_2;
	wire w_dff_B_5umnd9nw4_2;
	wire w_dff_B_0BLSgGkg2_2;
	wire w_dff_B_OXUIaxMq9_2;
	wire w_dff_B_S9W9NEpu2_2;
	wire w_dff_B_5LMjWyT50_2;
	wire w_dff_B_UEMTtNBy1_2;
	wire w_dff_B_eD72nMjZ9_2;
	wire w_dff_B_oNjwemyX7_2;
	wire w_dff_B_Bd2jz3141_2;
	wire w_dff_B_h9VDgHHg6_2;
	wire w_dff_B_hunrCV1g8_2;
	wire w_dff_B_Oip8vEve4_2;
	wire w_dff_B_CGb7fR6C3_2;
	wire w_dff_B_lhU3fi1G5_2;
	wire w_dff_B_LMRqX8TV9_2;
	wire w_dff_B_gbUfhRb91_2;
	wire w_dff_B_gTW28RTb5_2;
	wire w_dff_B_JzFV2ONK0_2;
	wire w_dff_B_wZ2WsLoG4_2;
	wire w_dff_B_32evhavQ6_2;
	wire w_dff_B_zRNwHgyq7_2;
	wire w_dff_B_CSIE9nZD5_2;
	wire w_dff_B_Hw8v52VP5_2;
	wire w_dff_B_Z0XSY5sY1_2;
	wire w_dff_B_hr8K6DLV8_2;
	wire w_dff_B_CpslQAyj1_2;
	wire w_dff_B_RY8Tk1dv4_2;
	wire w_dff_B_GBUU6KTQ5_2;
	wire w_dff_B_DjKzZ8ih2_2;
	wire w_dff_B_Novj0s5f8_2;
	wire w_dff_B_xk6Kvhft1_2;
	wire w_dff_B_OAoSmCH78_2;
	wire w_dff_B_apBZy1Lr3_2;
	wire w_dff_B_6vvQA9U62_2;
	wire w_dff_B_MZft0Rpa3_2;
	wire w_dff_B_Mlm0szhn8_2;
	wire w_dff_B_WmvtQHks0_2;
	wire w_dff_B_Hyy1Rhgv9_2;
	wire w_dff_B_vRqrLQ890_2;
	wire w_dff_B_4nmjdSV93_2;
	wire w_dff_B_GfL5xMsK7_2;
	wire w_dff_B_ZCZqkJND0_2;
	wire w_dff_B_aULq1Jt46_2;
	wire w_dff_B_RhxBNb8P7_0;
	wire w_dff_A_LfO3RIHK7_1;
	wire w_dff_B_JQvbpp403_1;
	wire w_dff_B_U90uMvAa1_2;
	wire w_dff_B_NoiBQRiJ2_2;
	wire w_dff_B_tL1mZXxV9_2;
	wire w_dff_B_enHzjiiw8_2;
	wire w_dff_B_rZPNWW4h8_2;
	wire w_dff_B_5d4oZ88T3_2;
	wire w_dff_B_LF8NBnL16_2;
	wire w_dff_B_aZ6ugA3w1_2;
	wire w_dff_B_6tSuWOSC7_2;
	wire w_dff_B_7VPh3tWa7_2;
	wire w_dff_B_IYxYnHIB6_2;
	wire w_dff_B_ZfUC2LkC6_2;
	wire w_dff_B_bJUgQ1XH8_2;
	wire w_dff_B_1nfqEaHb5_2;
	wire w_dff_B_HHn9aFlQ1_2;
	wire w_dff_B_GGXcCVo58_2;
	wire w_dff_B_Uuexpj197_2;
	wire w_dff_B_qmZSuspL3_2;
	wire w_dff_B_ujEsUb5c8_2;
	wire w_dff_B_WaY0OldU3_2;
	wire w_dff_B_8gIcdXQJ8_2;
	wire w_dff_B_XAq5HCEW5_2;
	wire w_dff_B_b152A6lN0_2;
	wire w_dff_B_k5sYsebK4_2;
	wire w_dff_B_p5e0Aezl2_2;
	wire w_dff_B_mIXScm0Q0_2;
	wire w_dff_B_pkiogah55_2;
	wire w_dff_B_y6dWHmgG4_2;
	wire w_dff_B_m9hCgzYF4_2;
	wire w_dff_B_QPQHOcDJ8_2;
	wire w_dff_B_Dm8NMg9V0_2;
	wire w_dff_B_5NYVmpA13_2;
	wire w_dff_B_QteqSDU96_2;
	wire w_dff_B_t2oKy07e8_2;
	wire w_dff_B_2a6sqRoH9_2;
	wire w_dff_B_AFtX9sIe1_2;
	wire w_dff_B_mv30Dwhi6_2;
	wire w_dff_B_YQa0O84W7_2;
	wire w_dff_B_Ot77QrI62_2;
	wire w_dff_B_Iuv5wbIc7_2;
	wire w_dff_B_O1NHPjoB7_2;
	wire w_dff_B_lOSBJ7tE3_1;
	wire w_dff_B_9RJNcfrF2_2;
	wire w_dff_B_aEoizBxe3_2;
	wire w_dff_B_HUhjX3n13_2;
	wire w_dff_B_FAnE5Wis5_2;
	wire w_dff_B_inS0zxTF9_2;
	wire w_dff_B_ocxw3Y8Y4_2;
	wire w_dff_B_jKQ9Slxc5_2;
	wire w_dff_B_K6n4O5zN0_2;
	wire w_dff_B_qOSioDeL5_2;
	wire w_dff_B_sqONaICq0_2;
	wire w_dff_B_Sn6e1hcZ3_2;
	wire w_dff_B_SeW8fSQC5_2;
	wire w_dff_B_HBLe2pbK5_2;
	wire w_dff_B_LW4q84Ob7_2;
	wire w_dff_B_SZByWkeP9_2;
	wire w_dff_B_efFwplAt5_2;
	wire w_dff_B_b34dtNXc7_2;
	wire w_dff_B_hUPtkb717_2;
	wire w_dff_B_iagk97iy3_2;
	wire w_dff_B_eEyigFEQ2_2;
	wire w_dff_B_Y2XLB0bw4_2;
	wire w_dff_B_upcuLzjl5_2;
	wire w_dff_B_Es71zjQl3_2;
	wire w_dff_B_CDVgHeAy7_2;
	wire w_dff_B_duaNfMR90_2;
	wire w_dff_B_PK063A7o8_2;
	wire w_dff_B_cavtLJ0J7_2;
	wire w_dff_B_Ta4lBXkR2_2;
	wire w_dff_B_nys8lKOj7_2;
	wire w_dff_B_K8vOuI1A7_2;
	wire w_dff_B_kcgKCWXT9_2;
	wire w_dff_B_w3iLftcQ4_2;
	wire w_dff_B_wyRUFoPh9_2;
	wire w_dff_B_XNdGnwWX0_2;
	wire w_dff_B_skBhd1sh3_2;
	wire w_dff_B_3azMdPCw2_2;
	wire w_dff_B_SzYlsXIl7_2;
	wire w_dff_B_dQDJWevx9_2;
	wire w_dff_B_eCtGb53e0_1;
	wire w_dff_B_TJ0XPJ058_2;
	wire w_dff_B_LFISirk68_2;
	wire w_dff_B_jKk0oP377_2;
	wire w_dff_B_42TnxQTR1_2;
	wire w_dff_B_eBVbqtvU6_2;
	wire w_dff_B_fmejP46P8_2;
	wire w_dff_B_P5Q0hKUW1_2;
	wire w_dff_B_tFj8JxWy3_2;
	wire w_dff_B_8kmoOYdH1_2;
	wire w_dff_B_xpmmf9ZZ5_2;
	wire w_dff_B_vVzBuWer4_2;
	wire w_dff_B_ia0jNExX5_2;
	wire w_dff_B_OxSmDrYf1_2;
	wire w_dff_B_yjNFD4bk2_2;
	wire w_dff_B_iN8QNmSG1_2;
	wire w_dff_B_DuOCbTw32_2;
	wire w_dff_B_v2omJpgm9_2;
	wire w_dff_B_9sJXtV8b3_2;
	wire w_dff_B_HyIdw98L7_2;
	wire w_dff_B_EmupylG62_2;
	wire w_dff_B_QFbOzZc40_2;
	wire w_dff_B_ECWOHVdg0_2;
	wire w_dff_B_Rw1BSHKQ9_2;
	wire w_dff_B_O5WmV9b73_2;
	wire w_dff_B_GxUPNd4x8_2;
	wire w_dff_B_vtbgzxZ13_2;
	wire w_dff_B_zpW5bKD34_2;
	wire w_dff_B_IJr7b9Kn5_2;
	wire w_dff_B_jpvW04FO2_2;
	wire w_dff_B_zcdynVVv1_2;
	wire w_dff_B_SOxiC8ch5_2;
	wire w_dff_B_yfTvDbjC5_2;
	wire w_dff_B_r9psN4dq6_2;
	wire w_dff_B_vZdHmVoe7_2;
	wire w_dff_B_pV0mhRZL3_2;
	wire w_dff_B_Rb5srVo57_1;
	wire w_dff_B_lZn9UF0Q4_2;
	wire w_dff_B_15z3pBvV7_2;
	wire w_dff_B_v8TT3key1_2;
	wire w_dff_B_3WxeF3as2_2;
	wire w_dff_B_cW4lRg5Y5_2;
	wire w_dff_B_on5C6lik6_2;
	wire w_dff_B_poWIt2H63_2;
	wire w_dff_B_keKaoNRj2_2;
	wire w_dff_B_YPAGzvB34_2;
	wire w_dff_B_sKfDDsa15_2;
	wire w_dff_B_145WmUMG5_2;
	wire w_dff_B_IDhYC0Mq0_2;
	wire w_dff_B_ltG2fnaH3_2;
	wire w_dff_B_fcwqtJuG0_2;
	wire w_dff_B_3iixEj0N7_2;
	wire w_dff_B_WrM8pzZb8_2;
	wire w_dff_B_4tTfQJlb0_2;
	wire w_dff_B_olsGP0uP6_2;
	wire w_dff_B_HoZJEgBU2_2;
	wire w_dff_B_26PZ9btN9_2;
	wire w_dff_B_wn9pbkMV8_2;
	wire w_dff_B_IKMYJJjS8_2;
	wire w_dff_B_0d4yX2xg0_2;
	wire w_dff_B_3XdOFMFu8_2;
	wire w_dff_B_WPiWKbN28_2;
	wire w_dff_B_3L6vqFYl4_2;
	wire w_dff_B_OtpxpA1G4_2;
	wire w_dff_B_5o0b8ZpA8_2;
	wire w_dff_B_pyChaReD3_2;
	wire w_dff_B_djIcuisx9_2;
	wire w_dff_B_E2Lm7Htj4_2;
	wire w_dff_B_eZBfBava6_2;
	wire w_dff_B_fWUgkO5b0_1;
	wire w_dff_B_6iUBDZHj4_2;
	wire w_dff_B_Fd0MyKka5_2;
	wire w_dff_B_ND8OBbwC0_2;
	wire w_dff_B_nErpmHl18_2;
	wire w_dff_B_2tEclMAK1_2;
	wire w_dff_B_lA9v8wsM5_2;
	wire w_dff_B_KnaG4l6K5_2;
	wire w_dff_B_m0I4GfXp4_2;
	wire w_dff_B_dwd3x7Ia6_2;
	wire w_dff_B_klRcr3bk7_2;
	wire w_dff_B_rl1m2nHq1_2;
	wire w_dff_B_gO1gN7Ik5_2;
	wire w_dff_B_GHym1I754_2;
	wire w_dff_B_jl9Ge0LM5_2;
	wire w_dff_B_x0QUaPVo7_2;
	wire w_dff_B_4qNuKCMZ4_2;
	wire w_dff_B_wWjawONr7_2;
	wire w_dff_B_YrfYcJyl0_2;
	wire w_dff_B_ALQWyxbg3_2;
	wire w_dff_B_VxcZ4zR37_2;
	wire w_dff_B_3SSxB3xy1_2;
	wire w_dff_B_r00RNczI8_2;
	wire w_dff_B_6TmPeOpD3_2;
	wire w_dff_B_QQGQvHcR2_2;
	wire w_dff_B_uwyEBFDM8_2;
	wire w_dff_B_PWGYKLKY5_2;
	wire w_dff_B_e6K5chWS2_2;
	wire w_dff_B_fj8Vgs8k0_2;
	wire w_dff_B_c0w64E9o7_2;
	wire w_dff_B_mxcrFEy75_1;
	wire w_dff_B_4OMtVokv1_2;
	wire w_dff_B_acoRmwt28_2;
	wire w_dff_B_9KkUNVVI6_2;
	wire w_dff_B_G1Bo0LPI7_2;
	wire w_dff_B_JICtEKpQ8_2;
	wire w_dff_B_pEUGoxrz8_2;
	wire w_dff_B_N306hy2O3_2;
	wire w_dff_B_lceEbzHj3_2;
	wire w_dff_B_gFD0s3mq0_2;
	wire w_dff_B_2lffssTC4_2;
	wire w_dff_B_Yxr7O1Uj6_2;
	wire w_dff_B_5YMx5so30_2;
	wire w_dff_B_oexpnFcj0_2;
	wire w_dff_B_AQJqsCTT4_2;
	wire w_dff_B_4psAA1UQ1_2;
	wire w_dff_B_0eo6v2GS3_2;
	wire w_dff_B_297USJ0g9_2;
	wire w_dff_B_mAYcP06y0_2;
	wire w_dff_B_NGHXSi535_2;
	wire w_dff_B_lU1WgcM25_2;
	wire w_dff_B_phJ4JOgn2_2;
	wire w_dff_B_6Lz8YEo09_2;
	wire w_dff_B_q7GzRp9T7_2;
	wire w_dff_B_43Y1xxIr5_2;
	wire w_dff_B_UDGVpLg17_2;
	wire w_dff_B_ycB40T2b3_2;
	wire w_dff_B_ygjs60Th7_1;
	wire w_dff_B_Z0Duo9dV0_2;
	wire w_dff_B_VRnX6mHH9_2;
	wire w_dff_B_hXfiWR3P6_2;
	wire w_dff_B_3jIfXF6T0_2;
	wire w_dff_B_vdyx2JQE5_2;
	wire w_dff_B_lOPKwDuT8_2;
	wire w_dff_B_l3MrveyU8_2;
	wire w_dff_B_4NWA4bwp0_2;
	wire w_dff_B_eOjGzMjl3_2;
	wire w_dff_B_x5te0b223_2;
	wire w_dff_B_ynbAoZOU9_2;
	wire w_dff_B_oaA6cAh42_2;
	wire w_dff_B_yBxAq33v3_2;
	wire w_dff_B_5faZdRXQ3_2;
	wire w_dff_B_DyBzSxvy7_2;
	wire w_dff_B_b2UQyiTc7_2;
	wire w_dff_B_EjFXhMjI9_2;
	wire w_dff_B_O4ZLzo7Q7_2;
	wire w_dff_B_OEPcdrkb7_2;
	wire w_dff_B_arWQVsp99_2;
	wire w_dff_B_xctT5K701_2;
	wire w_dff_B_DGBVxjsn9_2;
	wire w_dff_B_vZ6KDoV16_2;
	wire w_dff_B_WMEeveX70_1;
	wire w_dff_B_8xYkexNR0_2;
	wire w_dff_B_XchKCJZz6_2;
	wire w_dff_B_BcqWLi289_2;
	wire w_dff_B_7Ixca6yZ6_2;
	wire w_dff_B_GfjppUmw8_2;
	wire w_dff_B_TL87T78e5_2;
	wire w_dff_B_c6ACRB5u9_2;
	wire w_dff_B_7NIqPGV22_2;
	wire w_dff_B_648NKTum2_2;
	wire w_dff_B_uf0MxER77_2;
	wire w_dff_B_zrLxTw9F9_2;
	wire w_dff_B_8H5kqOg08_2;
	wire w_dff_B_lCivCT015_2;
	wire w_dff_B_qMyG07dM2_2;
	wire w_dff_B_TGb8nIso0_2;
	wire w_dff_B_HDWsRIIj2_2;
	wire w_dff_B_DsXCdJIH8_2;
	wire w_dff_B_sKSNMA531_2;
	wire w_dff_B_A3MxRWOn7_2;
	wire w_dff_B_DFyyoA0N0_2;
	wire w_dff_B_VvhQZ0NB6_1;
	wire w_dff_B_pgbrNAnr1_2;
	wire w_dff_B_bEdYUBvI7_2;
	wire w_dff_B_zugL85Ye3_2;
	wire w_dff_B_i48PGo582_2;
	wire w_dff_B_te4HLu1p9_2;
	wire w_dff_B_hwMFpPo93_2;
	wire w_dff_B_A60vuWWt2_2;
	wire w_dff_B_EQBRvvYW5_2;
	wire w_dff_B_QIrZ9R2b6_2;
	wire w_dff_B_aDMKBFu62_2;
	wire w_dff_B_HTRPVf4C5_2;
	wire w_dff_B_ziCjGJz67_2;
	wire w_dff_B_eIRFFKhB0_2;
	wire w_dff_B_txtJm3rF6_2;
	wire w_dff_B_k4XIAjuc1_2;
	wire w_dff_B_RNkWNosq9_2;
	wire w_dff_B_J6QBkd1c4_2;
	wire w_dff_B_UaNQnCtd9_1;
	wire w_dff_B_dighet794_2;
	wire w_dff_B_XMXdOW4Z5_2;
	wire w_dff_B_vKmnixM04_2;
	wire w_dff_B_MoWautym2_2;
	wire w_dff_B_758aSQuj9_2;
	wire w_dff_B_dFY0FqmX0_2;
	wire w_dff_B_ht9z6Nlz5_2;
	wire w_dff_B_6LLvWaqw6_2;
	wire w_dff_B_neqTqmG74_2;
	wire w_dff_B_NsYz8Tbc1_2;
	wire w_dff_B_0bhSfjpg3_2;
	wire w_dff_B_WSbE96bQ3_2;
	wire w_dff_B_TCa8Nxe60_2;
	wire w_dff_B_nnVOysn11_2;
	wire w_dff_B_ztAH3VDi4_1;
	wire w_dff_B_mwJc1BeS3_2;
	wire w_dff_B_3sxCiYtf9_2;
	wire w_dff_B_RLpQhle37_2;
	wire w_dff_B_b01OVPTv4_2;
	wire w_dff_B_YVIsgybR5_2;
	wire w_dff_B_B7qquJtX8_2;
	wire w_dff_B_Ea8Tq7lI1_2;
	wire w_dff_B_qcWevvG74_2;
	wire w_dff_B_5s5oyIZD3_2;
	wire w_dff_B_BMfrFhAf7_2;
	wire w_dff_B_cFedhM6m6_2;
	wire w_dff_B_lIUTpAE80_1;
	wire w_dff_B_uL5pjgHx5_2;
	wire w_dff_B_tHoIgdej0_2;
	wire w_dff_B_VQfOBjtP3_2;
	wire w_dff_B_xiJINwsA5_2;
	wire w_dff_B_3ZyEqvnH6_2;
	wire w_dff_B_BG0lSzJ73_2;
	wire w_dff_B_9cmf9K3G9_2;
	wire w_dff_B_nalj3afZ5_2;
	wire w_dff_B_BmR3h8NF0_1;
	wire w_dff_B_fEsB0Ljq9_0;
	wire w_dff_B_Su4WFigI8_2;
	wire w_dff_B_jnLnM26k1_2;
	wire w_dff_B_nHW52yND5_2;
	wire w_dff_B_psp5KmyI1_2;
	wire w_dff_B_74u3CizV5_1;
	wire w_dff_A_lY35Gf6q5_0;
	wire w_dff_A_4KBjmpb35_0;
	wire w_dff_A_g6U8xrxE7_0;
	wire w_dff_A_IX8YLItY8_1;
	wire w_dff_B_5P4pp9zh5_2;
	wire w_dff_B_2YkkQ9rd3_1;
	wire w_dff_B_JuqYWJY15_2;
	wire w_dff_B_MFOTu59Z4_2;
	wire w_dff_B_pUrciEDZ6_2;
	wire w_dff_B_ae0rn1Vl9_2;
	wire w_dff_B_QQMrrVrk5_2;
	wire w_dff_B_4kSfgJ1w5_2;
	wire w_dff_B_lm8Xe7PB3_2;
	wire w_dff_B_oohCaw863_2;
	wire w_dff_B_ZKqaoZ7F4_2;
	wire w_dff_B_9n80JxzK0_2;
	wire w_dff_B_9GOdYVMe1_2;
	wire w_dff_B_W0HuBbm93_2;
	wire w_dff_B_2WXWACs30_2;
	wire w_dff_B_ItzjVcsw5_2;
	wire w_dff_B_jSscDheQ5_2;
	wire w_dff_B_IFADsWC58_2;
	wire w_dff_B_X2amMj6X1_2;
	wire w_dff_B_hz0cZMFW7_2;
	wire w_dff_B_R3E6d6yl4_2;
	wire w_dff_B_Jtl4fyGM1_2;
	wire w_dff_B_0iPHElpd8_2;
	wire w_dff_B_sCXxBtso0_2;
	wire w_dff_B_hgajkR5L3_2;
	wire w_dff_B_MflVSr1N3_2;
	wire w_dff_B_uFbs19s49_2;
	wire w_dff_B_JdRzqbq86_2;
	wire w_dff_B_uEbBayz01_2;
	wire w_dff_B_966hOrhk2_2;
	wire w_dff_B_TG4B0ySn7_2;
	wire w_dff_B_vUJgjzdo4_2;
	wire w_dff_B_1Zqukoio1_2;
	wire w_dff_B_QgioRiTJ3_2;
	wire w_dff_B_m8IPSO2E5_2;
	wire w_dff_B_z0uyovCq3_2;
	wire w_dff_B_6P9Ru5e75_2;
	wire w_dff_B_Mf8FdXk30_2;
	wire w_dff_B_2vxJTD2u6_2;
	wire w_dff_B_zKVWfg8V0_2;
	wire w_dff_B_tzpUw0ad2_2;
	wire w_dff_B_SicE7c7A6_2;
	wire w_dff_B_uumtACLN2_2;
	wire w_dff_B_FZ6IXBKU5_2;
	wire w_dff_B_cSvpNLU87_2;
	wire w_dff_B_GjTXKUHD5_2;
	wire w_dff_B_mJ9wVZH48_2;
	wire w_dff_B_Y7cEae5U1_1;
	wire w_dff_B_R0URrd2P3_2;
	wire w_dff_B_hwqMBUsx1_2;
	wire w_dff_B_YErTvJtL1_2;
	wire w_dff_B_zut8PZZn6_2;
	wire w_dff_B_UbOtM6RN0_2;
	wire w_dff_B_wieL0KOK9_2;
	wire w_dff_B_pej1ijAG6_2;
	wire w_dff_B_8IfK4BbJ0_2;
	wire w_dff_B_wzqxTmUW5_2;
	wire w_dff_B_3zUfbgfe6_2;
	wire w_dff_B_9u2PPMPm8_2;
	wire w_dff_B_somNHLV52_2;
	wire w_dff_B_wL41hHxW5_2;
	wire w_dff_B_j9GT010h3_2;
	wire w_dff_B_cX1W1JIx9_2;
	wire w_dff_B_8jhoHevL2_2;
	wire w_dff_B_uC7tnTzC1_2;
	wire w_dff_B_EbtojuWS9_2;
	wire w_dff_B_ev9XnmBM8_2;
	wire w_dff_B_wOC6kAbp3_2;
	wire w_dff_B_rgSopqSd3_2;
	wire w_dff_B_4LkbpIWS1_2;
	wire w_dff_B_Cd3jsIgJ2_2;
	wire w_dff_B_Jzi6yvEP6_2;
	wire w_dff_B_fF6d4owR2_2;
	wire w_dff_B_CBEP8Hgy4_2;
	wire w_dff_B_eEsFpIIl4_2;
	wire w_dff_B_b2m5Bg1A5_2;
	wire w_dff_B_h6bXhJra1_2;
	wire w_dff_B_PAMu7WGB0_2;
	wire w_dff_B_2Bnc9tCI2_2;
	wire w_dff_B_NyIK2i0x2_2;
	wire w_dff_B_KJkA6zte2_2;
	wire w_dff_B_DCwdtyls8_2;
	wire w_dff_B_nYNWCZCP3_2;
	wire w_dff_B_3jzPG3fB9_2;
	wire w_dff_B_fzmUEzNP9_2;
	wire w_dff_B_Krivrsg29_2;
	wire w_dff_B_MIEuH8hx6_2;
	wire w_dff_B_zS3qZF2g9_2;
	wire w_dff_B_veZHBUJv1_1;
	wire w_dff_B_lLeaJOqU6_2;
	wire w_dff_B_Gpc8TddJ5_2;
	wire w_dff_B_3dtFcCsZ5_2;
	wire w_dff_B_NgCwOr0u0_2;
	wire w_dff_B_4oDTmw7D5_2;
	wire w_dff_B_HJtdDzz43_2;
	wire w_dff_B_VEuFlud65_2;
	wire w_dff_B_JW6v6wyL5_2;
	wire w_dff_B_r83ELxry2_2;
	wire w_dff_B_LOIXOIv78_2;
	wire w_dff_B_F6yoJNjV6_2;
	wire w_dff_B_zLLd9rv06_2;
	wire w_dff_B_2BhHRQih1_2;
	wire w_dff_B_JB3k6geG3_2;
	wire w_dff_B_5q3NxEkH7_2;
	wire w_dff_B_eSBQStM02_2;
	wire w_dff_B_Y8TEAzYS5_2;
	wire w_dff_B_p9w5r6di2_2;
	wire w_dff_B_o7hHWP8Z2_2;
	wire w_dff_B_Nn3vFM4n8_2;
	wire w_dff_B_tSw5WrnD2_2;
	wire w_dff_B_61w3WLDm2_2;
	wire w_dff_B_P17ohZkU7_2;
	wire w_dff_B_RjHV7ITZ0_2;
	wire w_dff_B_9Tz4lley7_2;
	wire w_dff_B_QkGmoXMf7_2;
	wire w_dff_B_6sVUDqCe5_2;
	wire w_dff_B_VwWx60VY1_2;
	wire w_dff_B_czw2cOJi9_2;
	wire w_dff_B_NZD7xLZ20_2;
	wire w_dff_B_bXjCGVl78_2;
	wire w_dff_B_ViKNaZDL6_2;
	wire w_dff_B_xm6oSMuN9_2;
	wire w_dff_B_w1Q7IhUT5_2;
	wire w_dff_B_g0wfKieS7_2;
	wire w_dff_B_yb8ttNkF6_2;
	wire w_dff_B_WFUfie7T9_2;
	wire w_dff_B_uOEOZObL3_1;
	wire w_dff_B_1ojTqbuu5_2;
	wire w_dff_B_Mu1h62B41_2;
	wire w_dff_B_h48RORwK8_2;
	wire w_dff_B_M8KCaOh65_2;
	wire w_dff_B_id2XqKqF6_2;
	wire w_dff_B_477vbMIP6_2;
	wire w_dff_B_YARh4HJy9_2;
	wire w_dff_B_iaZlrNcx3_2;
	wire w_dff_B_cXwSHk198_2;
	wire w_dff_B_RUWyyqcD6_2;
	wire w_dff_B_Z0uOcxay9_2;
	wire w_dff_B_iYnFwR0M6_2;
	wire w_dff_B_kyLjDg9w9_2;
	wire w_dff_B_pVeZ9JKP0_2;
	wire w_dff_B_LMlpdPGc4_2;
	wire w_dff_B_0pEm2brJ7_2;
	wire w_dff_B_caSTd6PM9_2;
	wire w_dff_B_PePFdTAP5_2;
	wire w_dff_B_jsD4HgHt8_2;
	wire w_dff_B_Sg1wUg0H2_2;
	wire w_dff_B_yF28aubg9_2;
	wire w_dff_B_tvAuubX99_2;
	wire w_dff_B_4BqsZZHS4_2;
	wire w_dff_B_A81Y95J23_2;
	wire w_dff_B_kPfcUBLB3_2;
	wire w_dff_B_g2enGmPe7_2;
	wire w_dff_B_fZHCOcL76_2;
	wire w_dff_B_53SXnkVu4_2;
	wire w_dff_B_kCbt8Nyg5_2;
	wire w_dff_B_fJoq84PA2_2;
	wire w_dff_B_cRtX1KIi2_2;
	wire w_dff_B_TMcWbaYf7_2;
	wire w_dff_B_GOyUKeLb9_2;
	wire w_dff_B_4P83CbSp6_2;
	wire w_dff_B_UhIogdie1_1;
	wire w_dff_B_ar28uOhU3_2;
	wire w_dff_B_Mbxc45If8_2;
	wire w_dff_B_IRIz1hRJ5_2;
	wire w_dff_B_sAwZzgXI3_2;
	wire w_dff_B_Su7aprlm6_2;
	wire w_dff_B_0uBCu5Mm2_2;
	wire w_dff_B_zevdaLSW5_2;
	wire w_dff_B_Q7unzoo97_2;
	wire w_dff_B_mjsYeI5S9_2;
	wire w_dff_B_3un0WgMB5_2;
	wire w_dff_B_J0Da3LgN1_2;
	wire w_dff_B_u054pjDB7_2;
	wire w_dff_B_k3aJothM2_2;
	wire w_dff_B_C2ncuhDq0_2;
	wire w_dff_B_U3SgzjHC2_2;
	wire w_dff_B_Fuqn5Uxb5_2;
	wire w_dff_B_4jyMa10R5_2;
	wire w_dff_B_coKJHB6e8_2;
	wire w_dff_B_rmaE43Yd5_2;
	wire w_dff_B_j4sQzHwf7_2;
	wire w_dff_B_dN0cZSOu0_2;
	wire w_dff_B_UaO0raDX3_2;
	wire w_dff_B_zAux4gZk5_2;
	wire w_dff_B_lKn1YUqf5_2;
	wire w_dff_B_386CQtn60_2;
	wire w_dff_B_rpCfMSGh8_2;
	wire w_dff_B_Sivw5WCI8_2;
	wire w_dff_B_h1mTn8qL8_2;
	wire w_dff_B_zQTzwlJ39_2;
	wire w_dff_B_wHbRWiRb4_2;
	wire w_dff_B_eSqY2FEm1_2;
	wire w_dff_B_Ty6trjOr3_1;
	wire w_dff_B_zyptDpkY2_2;
	wire w_dff_B_y4Ube5an2_2;
	wire w_dff_B_I4zNbDoI3_2;
	wire w_dff_B_iC6EmDSr4_2;
	wire w_dff_B_MrZ7h7iX8_2;
	wire w_dff_B_9C48Tz4M7_2;
	wire w_dff_B_eY43w6qp7_2;
	wire w_dff_B_94bRS6Zc3_2;
	wire w_dff_B_MnxwYbbG6_2;
	wire w_dff_B_FcPa4WaH5_2;
	wire w_dff_B_yTvnrMGf7_2;
	wire w_dff_B_tmnxWpXx3_2;
	wire w_dff_B_mP67yWkI7_2;
	wire w_dff_B_ZVEW2Wgg7_2;
	wire w_dff_B_jEqc3vX75_2;
	wire w_dff_B_meSBabrK2_2;
	wire w_dff_B_js3dBYcS8_2;
	wire w_dff_B_BNKNvkt61_2;
	wire w_dff_B_0xtg43hz4_2;
	wire w_dff_B_lgd5mQvA2_2;
	wire w_dff_B_sCW2FjgQ1_2;
	wire w_dff_B_hMKtJyxY7_2;
	wire w_dff_B_SgOIII2a1_2;
	wire w_dff_B_LwYy6BIU8_2;
	wire w_dff_B_NdHpaAPw4_2;
	wire w_dff_B_na7o3CWK8_2;
	wire w_dff_B_o4fmtzml8_2;
	wire w_dff_B_j1yGSPFY8_2;
	wire w_dff_B_aOKnKsbI5_1;
	wire w_dff_B_t8WFISp08_2;
	wire w_dff_B_44nP9i2V4_2;
	wire w_dff_B_5bAK6Yg66_2;
	wire w_dff_B_wihg9dZv6_2;
	wire w_dff_B_y7sptAQY7_2;
	wire w_dff_B_r347IwI28_2;
	wire w_dff_B_OyhCjVUy9_2;
	wire w_dff_B_Ab5EYeQs5_2;
	wire w_dff_B_5E4cWV1U8_2;
	wire w_dff_B_usSTADm85_2;
	wire w_dff_B_C9OMeGqX5_2;
	wire w_dff_B_EVQJ2NAe5_2;
	wire w_dff_B_zaFgKXCb5_2;
	wire w_dff_B_B9iZeQ1Q6_2;
	wire w_dff_B_76jpFiPs1_2;
	wire w_dff_B_GMAX2RNd1_2;
	wire w_dff_B_oYUp9omq1_2;
	wire w_dff_B_qFhHMkon7_2;
	wire w_dff_B_o3ablrzL1_2;
	wire w_dff_B_UQv29VuB1_2;
	wire w_dff_B_M7jLzGgz1_2;
	wire w_dff_B_PwLVjtrM8_2;
	wire w_dff_B_KYXnVwUT0_2;
	wire w_dff_B_kmKD18UZ3_2;
	wire w_dff_B_zR9qlZKD4_2;
	wire w_dff_B_F4vP9F4i6_1;
	wire w_dff_B_1p18hD567_2;
	wire w_dff_B_MLapcce12_2;
	wire w_dff_B_EBSLFvWC5_2;
	wire w_dff_B_APz24RGh2_2;
	wire w_dff_B_6mYl2Ci25_2;
	wire w_dff_B_AKhJBG480_2;
	wire w_dff_B_5i0imjQS0_2;
	wire w_dff_B_NUXUo0vc7_2;
	wire w_dff_B_spQShVNE1_2;
	wire w_dff_B_EQeg9lbJ2_2;
	wire w_dff_B_tLQFADPr9_2;
	wire w_dff_B_EP7XPJMF7_2;
	wire w_dff_B_l5VjWV6J7_2;
	wire w_dff_B_EhiQJxor2_2;
	wire w_dff_B_HoUupqzo8_2;
	wire w_dff_B_8xTQIdKM1_2;
	wire w_dff_B_eXlfqz2o1_2;
	wire w_dff_B_FRfXUKr84_2;
	wire w_dff_B_9KiotzSZ4_2;
	wire w_dff_B_W62zzIzD4_2;
	wire w_dff_B_3KK4QQkq5_2;
	wire w_dff_B_QpjVlIc90_2;
	wire w_dff_B_9M5pmyQ40_1;
	wire w_dff_B_3Oy4zAc83_2;
	wire w_dff_B_RbVCnQe98_2;
	wire w_dff_B_1pczOuZR7_2;
	wire w_dff_B_6yB0xafJ0_2;
	wire w_dff_B_SuSjQcXD1_2;
	wire w_dff_B_DxiDnaAc5_2;
	wire w_dff_B_qiywJnVB2_2;
	wire w_dff_B_WVtFyks58_2;
	wire w_dff_B_16hPDcOk3_2;
	wire w_dff_B_GIDQdYSE8_2;
	wire w_dff_B_hjY8zbRe0_2;
	wire w_dff_B_flV9nWky7_2;
	wire w_dff_B_f6MA30B28_2;
	wire w_dff_B_rtRNaiLF9_2;
	wire w_dff_B_Weew9LTl7_2;
	wire w_dff_B_sPbCZpbO2_2;
	wire w_dff_B_UX0a4oAJ7_2;
	wire w_dff_B_ifbYKzyJ1_2;
	wire w_dff_B_qqduDE2g4_2;
	wire w_dff_B_s9Cd84hT8_1;
	wire w_dff_B_ZSz19q7P4_2;
	wire w_dff_B_Lq2hAwIk1_2;
	wire w_dff_B_R58AkyAS8_2;
	wire w_dff_B_2bS28fJ98_2;
	wire w_dff_B_X2Svo9sr2_2;
	wire w_dff_B_JEo17NHy5_2;
	wire w_dff_B_SgkybFcA6_2;
	wire w_dff_B_LY8odb8R5_2;
	wire w_dff_B_rVpjdAN79_2;
	wire w_dff_B_lyJmV2WD3_2;
	wire w_dff_B_yUNS7d8j9_2;
	wire w_dff_B_So8gVGsf1_2;
	wire w_dff_B_E31YnTJc1_2;
	wire w_dff_B_SeWOF00b6_2;
	wire w_dff_B_1g9pyNQd0_2;
	wire w_dff_B_1WJwsVqu8_2;
	wire w_dff_B_qAkQqxEW1_1;
	wire w_dff_B_DRRdmiDW3_2;
	wire w_dff_B_urIvva7L5_2;
	wire w_dff_B_MuWDCOfI2_2;
	wire w_dff_B_IKxz5faF8_2;
	wire w_dff_B_MUQ3CgdL6_2;
	wire w_dff_B_atjKpGNi7_2;
	wire w_dff_B_OXNf1yG70_2;
	wire w_dff_B_1UWUrrwO9_2;
	wire w_dff_B_qce8hfQB1_2;
	wire w_dff_B_mGHPOroW1_2;
	wire w_dff_B_mHDzVxhK5_2;
	wire w_dff_B_Vu6i6Fll3_2;
	wire w_dff_B_WVEh5NPZ2_2;
	wire w_dff_B_BnZj7UBm8_1;
	wire w_dff_B_4QyvSVSR8_2;
	wire w_dff_B_IIx56gXe0_2;
	wire w_dff_B_6wZH7Ok81_2;
	wire w_dff_B_gkNvJvQH7_2;
	wire w_dff_B_PUvLPEbX8_2;
	wire w_dff_B_613AM2O79_2;
	wire w_dff_B_xrCZWvcG0_2;
	wire w_dff_B_ly6g3P1U1_2;
	wire w_dff_B_QaJT2DOY0_2;
	wire w_dff_B_wVO3rB1a0_2;
	wire w_dff_B_OOIwGHPY4_2;
	wire w_dff_B_TK43nvRb3_1;
	wire w_dff_B_L7G2pKg59_2;
	wire w_dff_B_0KwACUyX9_2;
	wire w_dff_B_kIK5WVBH9_2;
	wire w_dff_B_8YKbz1RU8_2;
	wire w_dff_B_F5ySW75Y5_2;
	wire w_dff_B_ffnSJ3H53_2;
	wire w_dff_B_JqLKAmu29_2;
	wire w_dff_B_NxEO5AfJ9_2;
	wire w_dff_B_p983pDwu3_1;
	wire w_dff_B_Lj5YMUYh5_2;
	wire w_dff_B_xBmmamQh7_2;
	wire w_dff_B_JlmFxbUl8_2;
	wire w_dff_B_Cjc6iVEW9_2;
	wire w_dff_B_9IuVKnvE7_1;
	wire w_dff_A_pnxRAwe47_1;
	wire w_dff_A_bReyMFdL4_2;
	wire w_dff_A_MHJ6KRGP1_2;
	wire w_dff_B_1PbYWcAW4_2;
	wire w_dff_B_RRuD0sth9_1;
	wire w_dff_B_phbo0j6D0_2;
	wire w_dff_B_8YVilGzq5_2;
	wire w_dff_B_BmzU59om7_2;
	wire w_dff_B_YVIktdGg6_2;
	wire w_dff_B_8ydDYcP81_2;
	wire w_dff_B_OQgfeYhR3_2;
	wire w_dff_B_G11Lskv29_2;
	wire w_dff_B_CQCWSLBS8_2;
	wire w_dff_B_sUEr4TXq0_2;
	wire w_dff_B_7MbSH3721_2;
	wire w_dff_B_SePz8io24_2;
	wire w_dff_B_NGQ8Tdl15_2;
	wire w_dff_B_lt75ed062_2;
	wire w_dff_B_VWqlhZly4_2;
	wire w_dff_B_ntIG5aVD8_2;
	wire w_dff_B_W8LSHsh81_2;
	wire w_dff_B_tSTUgfPQ8_2;
	wire w_dff_B_upkqrRwu6_2;
	wire w_dff_B_jy1WydnB1_2;
	wire w_dff_B_ohhgsH8T8_2;
	wire w_dff_B_stsMYuIm9_2;
	wire w_dff_B_U1tVEron5_2;
	wire w_dff_B_ZiUT98Jd3_2;
	wire w_dff_B_LaBPyo2r3_2;
	wire w_dff_B_GkAN6Om21_2;
	wire w_dff_B_tejtAvzC6_2;
	wire w_dff_B_cVencumn7_2;
	wire w_dff_B_IpnrKMFN1_2;
	wire w_dff_B_LjnXAPnO4_2;
	wire w_dff_B_INSiJQO72_2;
	wire w_dff_B_hKsAMLUP0_2;
	wire w_dff_B_oEVqmzXk3_2;
	wire w_dff_B_684SEqpv1_2;
	wire w_dff_B_SZaKRMyP0_2;
	wire w_dff_B_b7TOsfdU2_2;
	wire w_dff_B_GRC7YGEg7_2;
	wire w_dff_B_wBGrFOu90_2;
	wire w_dff_B_2ld1AzU40_2;
	wire w_dff_B_inHNCpSI0_2;
	wire w_dff_B_Q5QfrRvA9_2;
	wire w_dff_B_4HYX0Wkp9_2;
	wire w_dff_B_Z7CtsIPD6_2;
	wire w_dff_B_VF1cx7eZ3_2;
	wire w_dff_B_fExNCCvN4_2;
	wire w_dff_B_QRalWrY44_2;
	wire w_dff_B_wthlQ4w61_2;
	wire w_dff_B_sIuJ0ldn2_1;
	wire w_dff_B_6KJiEFqY2_2;
	wire w_dff_B_mw3p6vg57_2;
	wire w_dff_B_g5ipnwXZ8_2;
	wire w_dff_B_B7gmGxNR2_2;
	wire w_dff_B_Ti3DIU192_2;
	wire w_dff_B_lXKsN52i6_2;
	wire w_dff_B_1W4sHzwi9_2;
	wire w_dff_B_RAn4t7HL8_2;
	wire w_dff_B_ELJ6mODA6_2;
	wire w_dff_B_dwQbV2VH6_2;
	wire w_dff_B_O7zE7Wi63_2;
	wire w_dff_B_FtPLZGxp7_2;
	wire w_dff_B_649zuP3T6_2;
	wire w_dff_B_cFneH57W6_2;
	wire w_dff_B_DqeffqpD8_2;
	wire w_dff_B_bvBe0FNz4_2;
	wire w_dff_B_tywvN8aH2_2;
	wire w_dff_B_gLWEqJuP2_2;
	wire w_dff_B_6gYaM4J94_2;
	wire w_dff_B_RT9Hkvei7_2;
	wire w_dff_B_Zxgv8LjW3_2;
	wire w_dff_B_ZFv2T1Bh8_2;
	wire w_dff_B_DeWHq8RW5_2;
	wire w_dff_B_Fn2Kytrg2_2;
	wire w_dff_B_fOcOOTkF3_2;
	wire w_dff_B_wqZknIfA0_2;
	wire w_dff_B_XqwC3bhT1_2;
	wire w_dff_B_jiJk4psO8_2;
	wire w_dff_B_i43SwWRs6_2;
	wire w_dff_B_dXh13j5K4_2;
	wire w_dff_B_Kc0wYyDf7_2;
	wire w_dff_B_EvRJKgDR7_2;
	wire w_dff_B_NjoHizA18_2;
	wire w_dff_B_lotqe8Oh9_2;
	wire w_dff_B_AXmoDAIb4_2;
	wire w_dff_B_eLZ0OLec7_2;
	wire w_dff_B_wAglXE6F0_2;
	wire w_dff_B_UrBfy7n78_2;
	wire w_dff_B_odXcaD7i8_2;
	wire w_dff_B_M0LYrLI80_2;
	wire w_dff_B_Cg2CwX5J4_2;
	wire w_dff_B_1csLnxFv0_1;
	wire w_dff_B_b4kl91Zv3_2;
	wire w_dff_B_QsZYzkpk1_2;
	wire w_dff_B_tNrblsGQ5_2;
	wire w_dff_B_XxOCstFK5_2;
	wire w_dff_B_5ws6GyMH6_2;
	wire w_dff_B_XiBkvPrz0_2;
	wire w_dff_B_ANZU9JIL9_2;
	wire w_dff_B_S7iFtZF05_2;
	wire w_dff_B_G8OgqTJ99_2;
	wire w_dff_B_nNTVIRhW9_2;
	wire w_dff_B_Fq3mlY0W3_2;
	wire w_dff_B_42xAzjpx3_2;
	wire w_dff_B_PBaV0l5S1_2;
	wire w_dff_B_uNJs50bg3_2;
	wire w_dff_B_nJdHJFwc2_2;
	wire w_dff_B_UTjvwtPY6_2;
	wire w_dff_B_IjWk86Bp9_2;
	wire w_dff_B_pnuPGRxD0_2;
	wire w_dff_B_x8cpswUn2_2;
	wire w_dff_B_fGzF0AhU7_2;
	wire w_dff_B_bFI6WgSD4_2;
	wire w_dff_B_095JIYNe4_2;
	wire w_dff_B_EiJlTDHF4_2;
	wire w_dff_B_bQNSlO170_2;
	wire w_dff_B_NB2NLA2v6_2;
	wire w_dff_B_MGxVDMPn2_2;
	wire w_dff_B_ZXh3Z5mH3_2;
	wire w_dff_B_lqvgRkIg5_2;
	wire w_dff_B_Ec17dfrk4_2;
	wire w_dff_B_ASikrecF2_2;
	wire w_dff_B_oUB0YSab3_2;
	wire w_dff_B_rR8EqmPP1_2;
	wire w_dff_B_zjR6gQcK8_2;
	wire w_dff_B_OwcYP0uH8_2;
	wire w_dff_B_3d7wCdrG2_2;
	wire w_dff_B_mahCikNx5_2;
	wire w_dff_B_si4xxSjr1_2;
	wire w_dff_B_qyzV3BIc3_2;
	wire w_dff_B_9SfuAkYY9_1;
	wire w_dff_B_FsMcM0tO7_2;
	wire w_dff_B_2ED1pqdD9_2;
	wire w_dff_B_jzNsQ8RR5_2;
	wire w_dff_B_PRx9EmQN4_2;
	wire w_dff_B_GtqUXrql6_2;
	wire w_dff_B_JnZ8EYwP5_2;
	wire w_dff_B_5tNGFGjg9_2;
	wire w_dff_B_ddYVAcUU7_2;
	wire w_dff_B_5YFqgaWt4_2;
	wire w_dff_B_oUbmb7iS9_2;
	wire w_dff_B_Kqs9sEQy3_2;
	wire w_dff_B_o7EUY3su9_2;
	wire w_dff_B_mFHopx8k7_2;
	wire w_dff_B_vPeapwCx7_2;
	wire w_dff_B_LntdU5Z96_2;
	wire w_dff_B_LlkzF4AE4_2;
	wire w_dff_B_UoDF4jVm3_2;
	wire w_dff_B_mlborhS82_2;
	wire w_dff_B_kv6fnce34_2;
	wire w_dff_B_F5EZnrfI6_2;
	wire w_dff_B_hg5VPneE7_2;
	wire w_dff_B_Zc12SvIE2_2;
	wire w_dff_B_9JW8665k2_2;
	wire w_dff_B_GC3jK5Dl2_2;
	wire w_dff_B_g7K8x2lD0_2;
	wire w_dff_B_9zfFNM3v5_2;
	wire w_dff_B_vfkppYBB0_2;
	wire w_dff_B_JWG6VLI99_2;
	wire w_dff_B_xwEi4aM58_2;
	wire w_dff_B_m2V0cs3H6_2;
	wire w_dff_B_uhzNH2U43_2;
	wire w_dff_B_y8yadeKv2_2;
	wire w_dff_B_J8TzKbhy6_2;
	wire w_dff_B_v8I2cg8R8_2;
	wire w_dff_B_22AifnwD9_2;
	wire w_dff_B_Ow6XnM5z2_1;
	wire w_dff_B_fXdVR7Yh4_2;
	wire w_dff_B_P4h4V8Nh2_2;
	wire w_dff_B_HxI3PnX11_2;
	wire w_dff_B_KWBjY2yn2_2;
	wire w_dff_B_mKkk714A4_2;
	wire w_dff_B_qJJthC0G1_2;
	wire w_dff_B_mxh4hOpr8_2;
	wire w_dff_B_M77jESMV4_2;
	wire w_dff_B_mW368jgu3_2;
	wire w_dff_B_3CodNuHe9_2;
	wire w_dff_B_qmSuJsmC7_2;
	wire w_dff_B_cOYrjpoi4_2;
	wire w_dff_B_Z18h3vrZ8_2;
	wire w_dff_B_lYFzWjRi4_2;
	wire w_dff_B_qvJ3F9DW2_2;
	wire w_dff_B_Hf6gstuf4_2;
	wire w_dff_B_C5NwgdrA5_2;
	wire w_dff_B_YvHI9ZI63_2;
	wire w_dff_B_P5xYgdSi5_2;
	wire w_dff_B_W5nzsXYb7_2;
	wire w_dff_B_vlnoy0995_2;
	wire w_dff_B_D3JC63K48_2;
	wire w_dff_B_PaiYz4uk8_2;
	wire w_dff_B_4dNax5Ww0_2;
	wire w_dff_B_QXnmCyxB3_2;
	wire w_dff_B_1OwSHxWC7_2;
	wire w_dff_B_K27QHcQL5_2;
	wire w_dff_B_dAPh4Opn0_2;
	wire w_dff_B_dAL4aXgJ4_2;
	wire w_dff_B_N9dgmGfc2_2;
	wire w_dff_B_ZWAQwnOr9_2;
	wire w_dff_B_PMFJBWlE4_2;
	wire w_dff_B_Z0oss8sb3_1;
	wire w_dff_B_Mwi8CdeB6_2;
	wire w_dff_B_z5EpUGAC6_2;
	wire w_dff_B_XH4IWRzp9_2;
	wire w_dff_B_K2wgqb1J8_2;
	wire w_dff_B_hbks4zt12_2;
	wire w_dff_B_qyTI3Nyt3_2;
	wire w_dff_B_Dyoe2unM8_2;
	wire w_dff_B_pBRBWnLh8_2;
	wire w_dff_B_QcXGHQf89_2;
	wire w_dff_B_Fw28KfIW4_2;
	wire w_dff_B_PIOMStCF6_2;
	wire w_dff_B_gShgcL5Z6_2;
	wire w_dff_B_rie49QFk7_2;
	wire w_dff_B_SuTYyFwc0_2;
	wire w_dff_B_3z9HK80M4_2;
	wire w_dff_B_riCzz8px7_2;
	wire w_dff_B_rWRAWtER1_2;
	wire w_dff_B_wxI1J3450_2;
	wire w_dff_B_3LSC9JC04_2;
	wire w_dff_B_H4NMfe866_2;
	wire w_dff_B_Be4zUztE7_2;
	wire w_dff_B_fnUFx6UZ3_2;
	wire w_dff_B_durrI5fz2_2;
	wire w_dff_B_AGj8QWtJ3_2;
	wire w_dff_B_70vRGkCI2_2;
	wire w_dff_B_RgH76awt7_2;
	wire w_dff_B_xFU6vod69_2;
	wire w_dff_B_SadRMwjg6_2;
	wire w_dff_B_vTxBxvLn4_2;
	wire w_dff_B_rM9QpD1R3_1;
	wire w_dff_B_5dAVkk415_2;
	wire w_dff_B_aEObCI7S3_2;
	wire w_dff_B_q4kr5DnY3_2;
	wire w_dff_B_TsoL5NO09_2;
	wire w_dff_B_w0g1rqsj8_2;
	wire w_dff_B_uz6FBTgE1_2;
	wire w_dff_B_ifSb8xnW1_2;
	wire w_dff_B_twNRafDj6_2;
	wire w_dff_B_RWbUv56y6_2;
	wire w_dff_B_wJEGs35L2_2;
	wire w_dff_B_wrFkDeYM7_2;
	wire w_dff_B_IDmoxZk77_2;
	wire w_dff_B_K1cx9ejt3_2;
	wire w_dff_B_Xz83PU8N3_2;
	wire w_dff_B_9MEZUAb25_2;
	wire w_dff_B_VJnHLuVn6_2;
	wire w_dff_B_u5l4rsjr6_2;
	wire w_dff_B_QLfIW2Nn0_2;
	wire w_dff_B_Tn4eHpk71_2;
	wire w_dff_B_pLlPYgku6_2;
	wire w_dff_B_1D5k8vXx1_2;
	wire w_dff_B_EkusFtkZ6_2;
	wire w_dff_B_7mTBadUp4_2;
	wire w_dff_B_gPHTXJU91_2;
	wire w_dff_B_eWwKaM8K4_2;
	wire w_dff_B_Bg6ghQej4_2;
	wire w_dff_B_QYADrKf36_1;
	wire w_dff_B_iqYUAous7_2;
	wire w_dff_B_IEgBySH99_2;
	wire w_dff_B_nmKsp4GW7_2;
	wire w_dff_B_sSrGumgj2_2;
	wire w_dff_B_2xqrFsFT3_2;
	wire w_dff_B_PeuKAcu55_2;
	wire w_dff_B_O6TyCTLV1_2;
	wire w_dff_B_V4O8t3vE8_2;
	wire w_dff_B_nh2rqO655_2;
	wire w_dff_B_tkHSC4hs7_2;
	wire w_dff_B_WVMS96HE7_2;
	wire w_dff_B_SklZIgxa3_2;
	wire w_dff_B_DqNHx9xf9_2;
	wire w_dff_B_Lc8xv4eH8_2;
	wire w_dff_B_0C8Y6kl37_2;
	wire w_dff_B_MusmQAan0_2;
	wire w_dff_B_2jQ2rd5G9_2;
	wire w_dff_B_bbKFYL1K1_2;
	wire w_dff_B_dGWY89kj9_2;
	wire w_dff_B_aUznYYAe2_2;
	wire w_dff_B_rGFNe1vY4_2;
	wire w_dff_B_mIlvcbW99_2;
	wire w_dff_B_GrOGSWfp7_2;
	wire w_dff_B_j9Ffr4DS0_1;
	wire w_dff_B_S7TvtqRR6_2;
	wire w_dff_B_wU3lPNwg6_2;
	wire w_dff_B_KvYMa5gq0_2;
	wire w_dff_B_JcfDtML31_2;
	wire w_dff_B_F6mLJgiV3_2;
	wire w_dff_B_HiaFSaBM4_2;
	wire w_dff_B_S2wL8ocN7_2;
	wire w_dff_B_6L2vsn9P1_2;
	wire w_dff_B_EXuGGKSs2_2;
	wire w_dff_B_j8iIcsy09_2;
	wire w_dff_B_8OE73jPJ3_2;
	wire w_dff_B_LPNmaUta7_2;
	wire w_dff_B_0gKLIgS97_2;
	wire w_dff_B_zJhJNn6o8_2;
	wire w_dff_B_f8npws4O8_2;
	wire w_dff_B_NJOTFBwo4_2;
	wire w_dff_B_PQd7iCdk7_2;
	wire w_dff_B_dgvqKwQl5_2;
	wire w_dff_B_9uQXoqq93_2;
	wire w_dff_B_BUOFNaTh0_2;
	wire w_dff_B_mW1TSD8L4_1;
	wire w_dff_B_WKBOTvv13_2;
	wire w_dff_B_sqn5zKLR6_2;
	wire w_dff_B_JV4GuYjx5_2;
	wire w_dff_B_69kkkViF9_2;
	wire w_dff_B_M0pxyStW1_2;
	wire w_dff_B_Es4cV7i55_2;
	wire w_dff_B_zMfhwVej3_2;
	wire w_dff_B_CtmUTiVC0_2;
	wire w_dff_B_zCyAhcLj0_2;
	wire w_dff_B_iKz7KXCa2_2;
	wire w_dff_B_a8n0zfU29_2;
	wire w_dff_B_PhDtRwzW1_2;
	wire w_dff_B_Dz0DTGEy6_2;
	wire w_dff_B_QU4yYePb4_2;
	wire w_dff_B_CS5SZ2Kk7_2;
	wire w_dff_B_ACczwGNs0_2;
	wire w_dff_B_8w35Olta4_2;
	wire w_dff_B_1jkOuCTe1_1;
	wire w_dff_B_UU0niQwW9_2;
	wire w_dff_B_KeVEyKMb1_2;
	wire w_dff_B_IfGQKgo49_2;
	wire w_dff_B_v8NkCyuF8_2;
	wire w_dff_B_DmBSNOsi5_2;
	wire w_dff_B_Bx2gnNGo9_2;
	wire w_dff_B_B5o8vsOp5_2;
	wire w_dff_B_8WFP1M3O3_2;
	wire w_dff_B_EtJZypqQ0_2;
	wire w_dff_B_2hTid2xz7_2;
	wire w_dff_B_wIPEjqCa4_2;
	wire w_dff_B_t2VXvQob3_2;
	wire w_dff_B_ugtxxaRF8_2;
	wire w_dff_B_4A2pXL0w9_2;
	wire w_dff_B_o1AElAy04_1;
	wire w_dff_B_yaTJdMX62_2;
	wire w_dff_B_0xzqZkN16_2;
	wire w_dff_B_x4Y8O32m2_2;
	wire w_dff_B_bjdxf3zh8_2;
	wire w_dff_B_QQPzpzg94_2;
	wire w_dff_B_Ygl76m6v6_2;
	wire w_dff_B_F1A8SqEE5_2;
	wire w_dff_B_9Ppv3XtM6_2;
	wire w_dff_B_csYC4KPe7_2;
	wire w_dff_B_REcqCrEE4_2;
	wire w_dff_B_t22o2eFd8_2;
	wire w_dff_B_1TPbLWoN5_2;
	wire w_dff_B_OO1D15tP2_1;
	wire w_dff_B_9zEPRubG3_2;
	wire w_dff_B_sqaADirs6_2;
	wire w_dff_B_fWKoUnXJ9_2;
	wire w_dff_B_QunNc8Us6_2;
	wire w_dff_B_feEC5aAb8_2;
	wire w_dff_B_ShoRSDqQ1_2;
	wire w_dff_B_xUKku5GK7_2;
	wire w_dff_B_03fXdbCs7_1;
	wire w_dff_B_wUHlHhtp4_2;
	wire w_dff_B_YPvNkcuG0_2;
	wire w_dff_B_gIDleT7U8_2;
	wire w_dff_B_InSP26yk6_2;
	wire w_dff_B_pBKm8eeb1_1;
	wire w_dff_A_ND5nyXI76_0;
	wire w_dff_A_Sleh7iQV6_1;
	wire w_dff_A_oB75lPv25_1;
	wire w_dff_B_dscEN8CP3_1;
	wire w_dff_B_gZs9LaEz2_2;
	wire w_dff_B_PGEfNWI99_2;
	wire w_dff_B_W1Ek9dO77_2;
	wire w_dff_B_DDxqsWXw0_2;
	wire w_dff_B_OIYPBMRb4_2;
	wire w_dff_B_3syitiH25_2;
	wire w_dff_B_X0r7ewxt6_2;
	wire w_dff_B_YVKeeVHG7_2;
	wire w_dff_B_0KiXGFQ22_2;
	wire w_dff_B_OrxITFSE4_2;
	wire w_dff_B_p5XSaOeV3_2;
	wire w_dff_B_gX0PHthV9_2;
	wire w_dff_B_tSmN1HZK4_2;
	wire w_dff_B_bCg1fvIv9_2;
	wire w_dff_B_4rhMCbdM3_2;
	wire w_dff_B_zKAIuavT5_2;
	wire w_dff_B_WcE5HeEP9_2;
	wire w_dff_B_3v0Yo8XO9_2;
	wire w_dff_B_qz1XyZz10_2;
	wire w_dff_B_up5Fvazq8_2;
	wire w_dff_B_v26EmyiN3_2;
	wire w_dff_B_ybA0UQjG3_2;
	wire w_dff_B_gF3nxzH06_2;
	wire w_dff_B_iAAMCwx31_2;
	wire w_dff_B_3MjKph8N1_2;
	wire w_dff_B_5RdFssbW6_2;
	wire w_dff_B_uJfkE8X17_2;
	wire w_dff_B_w5zmZzTC5_2;
	wire w_dff_B_1goNVmJf8_2;
	wire w_dff_B_RwHDKR2h5_2;
	wire w_dff_B_SsVQtzwa4_2;
	wire w_dff_B_TzmBMLPI6_2;
	wire w_dff_B_H094nLHV7_2;
	wire w_dff_B_YWili5MT2_2;
	wire w_dff_B_NXZJJkEl4_2;
	wire w_dff_B_eODnW7n96_2;
	wire w_dff_B_VVeJMVTu0_2;
	wire w_dff_B_AFw9awkp9_2;
	wire w_dff_B_F4SSRS5d3_2;
	wire w_dff_B_unPgbOLe3_2;
	wire w_dff_B_xC7olaV15_2;
	wire w_dff_B_oWqxCd2C4_2;
	wire w_dff_B_XnMTc3tc5_2;
	wire w_dff_B_0UDdrsng6_2;
	wire w_dff_B_OdFVZsp64_2;
	wire w_dff_B_CeQ2fuut0_2;
	wire w_dff_B_ePm4FQ1L1_2;
	wire w_dff_B_xVbS7BIv1_0;
	wire w_dff_A_NoaSoI4S5_1;
	wire w_dff_B_lQf6csxZ2_1;
	wire w_dff_B_K8kUTWgq2_2;
	wire w_dff_B_CedpvwHs7_2;
	wire w_dff_B_7r2aTGij9_2;
	wire w_dff_B_dLvlGtDV0_2;
	wire w_dff_B_CMj8XDe25_2;
	wire w_dff_B_Y5UX4S5g2_2;
	wire w_dff_B_fGnOEmCY6_2;
	wire w_dff_B_dFvKUDWG2_2;
	wire w_dff_B_LZLEP57y7_2;
	wire w_dff_B_mL2VAuwq7_2;
	wire w_dff_B_QiyUvBsP5_2;
	wire w_dff_B_8zxexqDf3_2;
	wire w_dff_B_6oIlwFf77_2;
	wire w_dff_B_QIeW735N2_2;
	wire w_dff_B_t8xIgAYJ0_2;
	wire w_dff_B_WjDxrsoN8_2;
	wire w_dff_B_RJ1DzOCD2_2;
	wire w_dff_B_dPpnypC14_2;
	wire w_dff_B_YtEO3TLT3_2;
	wire w_dff_B_UarUl7fZ6_2;
	wire w_dff_B_Sj5WLCgo6_2;
	wire w_dff_B_s5q85r9E2_2;
	wire w_dff_B_ALefSdLr9_2;
	wire w_dff_B_24P93rEn5_2;
	wire w_dff_B_DouM5BnR5_2;
	wire w_dff_B_XicY1ay78_2;
	wire w_dff_B_MpMpxdGa3_2;
	wire w_dff_B_8XS9pli16_2;
	wire w_dff_B_dfwLvLV80_2;
	wire w_dff_B_eMQrLM579_2;
	wire w_dff_B_0g7HKPQi8_2;
	wire w_dff_B_gmFrnxSi7_2;
	wire w_dff_B_LHpRKbC69_2;
	wire w_dff_B_W5N0RPnN5_2;
	wire w_dff_B_RUCj2EVl5_2;
	wire w_dff_B_lfATVw4Z2_2;
	wire w_dff_B_9OaOwsta5_2;
	wire w_dff_B_5TU4Zch19_2;
	wire w_dff_B_mNTGIM3g0_2;
	wire w_dff_B_BNmq484u1_2;
	wire w_dff_B_ld4nXSo43_2;
	wire w_dff_B_hnjWvXPB6_2;
	wire w_dff_B_yDwue3896_2;
	wire w_dff_B_GNK67qew6_1;
	wire w_dff_B_mjwuSWFV6_2;
	wire w_dff_B_U9B1suxo8_2;
	wire w_dff_B_gb66n7Gz7_2;
	wire w_dff_B_M8ox9jiE1_2;
	wire w_dff_B_N6QIAid07_2;
	wire w_dff_B_Lx054sw25_2;
	wire w_dff_B_FCemGsSY4_2;
	wire w_dff_B_KJFQD4d71_2;
	wire w_dff_B_2u4iloU37_2;
	wire w_dff_B_nOkojfNl0_2;
	wire w_dff_B_23B6pC2S5_2;
	wire w_dff_B_MLegzzsA6_2;
	wire w_dff_B_qfg5kSDx2_2;
	wire w_dff_B_1abGkJLL3_2;
	wire w_dff_B_kRKuTYsx8_2;
	wire w_dff_B_Ku8lmRN92_2;
	wire w_dff_B_063y1oDD3_2;
	wire w_dff_B_4dR0k1Pe3_2;
	wire w_dff_B_uI4duSeb9_2;
	wire w_dff_B_ekNn9Kd60_2;
	wire w_dff_B_eNOnXkzs7_2;
	wire w_dff_B_pQ9JVMvA4_2;
	wire w_dff_B_91m689Lr0_2;
	wire w_dff_B_FXH8UVvw0_2;
	wire w_dff_B_7C8x3nza3_2;
	wire w_dff_B_sW6OVQP58_2;
	wire w_dff_B_k6h6274F0_2;
	wire w_dff_B_eQ2z22vz5_2;
	wire w_dff_B_qwQc6bcR9_2;
	wire w_dff_B_Pl7K4qeE4_2;
	wire w_dff_B_kjwtRpYF9_2;
	wire w_dff_B_3rpmHdA50_2;
	wire w_dff_B_lmYWVv327_2;
	wire w_dff_B_ymBku5oQ0_2;
	wire w_dff_B_JAcND1yG6_2;
	wire w_dff_B_dGRTS4v79_2;
	wire w_dff_B_c8zPlz7S7_2;
	wire w_dff_B_WBr45EPs8_2;
	wire w_dff_B_6NUDczgV1_2;
	wire w_dff_B_9ek3H3DE0_2;
	wire w_dff_B_faBXe0Lc1_1;
	wire w_dff_B_Zy0EmF5c8_2;
	wire w_dff_B_wxkXcXhe5_2;
	wire w_dff_B_6UXazMBB8_2;
	wire w_dff_B_0OQ4zjqZ5_2;
	wire w_dff_B_M37svjXN3_2;
	wire w_dff_B_48SDdk871_2;
	wire w_dff_B_tDVM4FSx0_2;
	wire w_dff_B_RnRX0C9p1_2;
	wire w_dff_B_jKbWh6lA2_2;
	wire w_dff_B_z1aBQxpj9_2;
	wire w_dff_B_zyFaztIQ2_2;
	wire w_dff_B_cX9Q2pET6_2;
	wire w_dff_B_kHfSLF8B6_2;
	wire w_dff_B_D5kFYsyw9_2;
	wire w_dff_B_rDwStpPN5_2;
	wire w_dff_B_vF3hEizx7_2;
	wire w_dff_B_AI8jw5il9_2;
	wire w_dff_B_lIeYby8V8_2;
	wire w_dff_B_nw4ESBAx9_2;
	wire w_dff_B_6qvCuHvB9_2;
	wire w_dff_B_bTUEaydP0_2;
	wire w_dff_B_9TVk05s40_2;
	wire w_dff_B_IMPzkTTk6_2;
	wire w_dff_B_IciobQ9S3_2;
	wire w_dff_B_olRmnmKX5_2;
	wire w_dff_B_D0Fo8iyw5_2;
	wire w_dff_B_XZfn5ScZ8_2;
	wire w_dff_B_xGr38sAj9_2;
	wire w_dff_B_iRazComT1_2;
	wire w_dff_B_6LfYAUrp2_2;
	wire w_dff_B_tMTFfhlg1_2;
	wire w_dff_B_KIPhj9SK0_2;
	wire w_dff_B_B4Ub5xnK4_2;
	wire w_dff_B_hVnXmHOG6_2;
	wire w_dff_B_Szd2QzRz4_2;
	wire w_dff_B_wK63IE4k2_2;
	wire w_dff_B_cN1DcKVD7_2;
	wire w_dff_B_ImpNrGtm4_1;
	wire w_dff_B_tupij4Nv5_2;
	wire w_dff_B_sHKsTPx80_2;
	wire w_dff_B_6vke0d8c0_2;
	wire w_dff_B_VLIgPtqg2_2;
	wire w_dff_B_yISFIlMI7_2;
	wire w_dff_B_vCX7vl4r7_2;
	wire w_dff_B_ROeHYyK89_2;
	wire w_dff_B_j8JRjkZw1_2;
	wire w_dff_B_OWIr4lcW8_2;
	wire w_dff_B_ihePhkrq9_2;
	wire w_dff_B_GVr11g0U7_2;
	wire w_dff_B_TvSbY1429_2;
	wire w_dff_B_KPrejBD39_2;
	wire w_dff_B_wBdZKpMH2_2;
	wire w_dff_B_AvTnVext5_2;
	wire w_dff_B_P9gTtpwK6_2;
	wire w_dff_B_ov0xG9pm8_2;
	wire w_dff_B_VGXCQCUd0_2;
	wire w_dff_B_kXYsHOV08_2;
	wire w_dff_B_1MMKTMfP2_2;
	wire w_dff_B_Of4YOxQd3_2;
	wire w_dff_B_4A2sPORL6_2;
	wire w_dff_B_fIhypljW9_2;
	wire w_dff_B_jWP9SUZ06_2;
	wire w_dff_B_D5aerA2U8_2;
	wire w_dff_B_CLOCFoYJ4_2;
	wire w_dff_B_9hCzTUK42_2;
	wire w_dff_B_fFiVH1kG4_2;
	wire w_dff_B_FKVraEVe9_2;
	wire w_dff_B_r3FGNd2r9_2;
	wire w_dff_B_2Xm7Rslv6_2;
	wire w_dff_B_HT9VLYAA6_2;
	wire w_dff_B_iArFbLF42_2;
	wire w_dff_B_X8PXlsSu2_2;
	wire w_dff_B_0sSPHn4O8_1;
	wire w_dff_B_c3Vd6GrN3_2;
	wire w_dff_B_lf3zomKh8_2;
	wire w_dff_B_FqoalI5p1_2;
	wire w_dff_B_BUS2HOza9_2;
	wire w_dff_B_NqlTAb3O0_2;
	wire w_dff_B_aJA2haG50_2;
	wire w_dff_B_MXv2KJ0H9_2;
	wire w_dff_B_5dIt3qRJ9_2;
	wire w_dff_B_tzWFpcnl3_2;
	wire w_dff_B_UE1XYbw51_2;
	wire w_dff_B_M4LX79iD3_2;
	wire w_dff_B_pMOogKxM1_2;
	wire w_dff_B_jQLXLeSi6_2;
	wire w_dff_B_m0zmUcfS8_2;
	wire w_dff_B_Umklu2qo4_2;
	wire w_dff_B_iIqrvonK1_2;
	wire w_dff_B_pRCVsK5J0_2;
	wire w_dff_B_FNJztTfC8_2;
	wire w_dff_B_prQxtbgJ4_2;
	wire w_dff_B_EyfdXWdF9_2;
	wire w_dff_B_MLxzRiDT8_2;
	wire w_dff_B_Scpb4JCl2_2;
	wire w_dff_B_al9HdKIK0_2;
	wire w_dff_B_JbQX7Hbj0_2;
	wire w_dff_B_BhDPqHiN3_2;
	wire w_dff_B_KCug5COe5_2;
	wire w_dff_B_vf3dco6h5_2;
	wire w_dff_B_MlpgTR5Q3_2;
	wire w_dff_B_MjcPfnJp5_2;
	wire w_dff_B_tE3GPyAT6_2;
	wire w_dff_B_Ey1mCoSe0_2;
	wire w_dff_B_EU9fSBA64_1;
	wire w_dff_B_msWHd3oh5_2;
	wire w_dff_B_Neyv2mKd0_2;
	wire w_dff_B_R6CN6o1L5_2;
	wire w_dff_B_qzQiVGiQ8_2;
	wire w_dff_B_EKLGHIcV9_2;
	wire w_dff_B_plfNoSIO3_2;
	wire w_dff_B_1twOcQB14_2;
	wire w_dff_B_DOMXe3GP5_2;
	wire w_dff_B_BPq00AG38_2;
	wire w_dff_B_OwlEvNCk5_2;
	wire w_dff_B_9691XIaT6_2;
	wire w_dff_B_Evd8MDCF3_2;
	wire w_dff_B_EWB6sXBG3_2;
	wire w_dff_B_7kx7y9Xv3_2;
	wire w_dff_B_7YH5rV9f4_2;
	wire w_dff_B_ol5XeFAm4_2;
	wire w_dff_B_nxNUkvJm1_2;
	wire w_dff_B_HHso2Rpj0_2;
	wire w_dff_B_W0w5z7bF8_2;
	wire w_dff_B_jTzzGAYl7_2;
	wire w_dff_B_Xuak1bne9_2;
	wire w_dff_B_Y4K0I4uD3_2;
	wire w_dff_B_vYRFEYbL2_2;
	wire w_dff_B_IpURNv8y7_2;
	wire w_dff_B_P3FSdtuF0_2;
	wire w_dff_B_6GbxEZyg9_2;
	wire w_dff_B_9B0pqAp15_2;
	wire w_dff_B_odIEMLG73_2;
	wire w_dff_B_P00V99xF6_1;
	wire w_dff_B_WJAPKH9r4_2;
	wire w_dff_B_Be2y1eLw1_2;
	wire w_dff_B_PP4BbTAx4_2;
	wire w_dff_B_knzvl6E08_2;
	wire w_dff_B_4SrQ0URV1_2;
	wire w_dff_B_yAIpMIn73_2;
	wire w_dff_B_UfsHC1C33_2;
	wire w_dff_B_5deEPxUu2_2;
	wire w_dff_B_ZQlbNdte0_2;
	wire w_dff_B_8ganj8Pt3_2;
	wire w_dff_B_wLDMP53B3_2;
	wire w_dff_B_QC9oHw9t2_2;
	wire w_dff_B_tkkr1hc26_2;
	wire w_dff_B_PBbUxTOK4_2;
	wire w_dff_B_GheVLLBZ8_2;
	wire w_dff_B_ygMLiikt8_2;
	wire w_dff_B_q5NYwUsE9_2;
	wire w_dff_B_3uzTq3Az3_2;
	wire w_dff_B_Rjet8Wn75_2;
	wire w_dff_B_J1iPLDCX0_2;
	wire w_dff_B_eF9Tk66p4_2;
	wire w_dff_B_47ZRFloy8_2;
	wire w_dff_B_H2RfDcbU6_2;
	wire w_dff_B_W4fjIvWG8_2;
	wire w_dff_B_SqSzmfJI2_2;
	wire w_dff_B_FwUjwLpg3_1;
	wire w_dff_B_sbiRgiuq9_2;
	wire w_dff_B_2qFNidnc3_2;
	wire w_dff_B_s8IYWgUJ6_2;
	wire w_dff_B_bfVDU8DR9_2;
	wire w_dff_B_Zsg35E7T0_2;
	wire w_dff_B_NIuS8Gao2_2;
	wire w_dff_B_2R3SzqrG6_2;
	wire w_dff_B_RnlveGLs4_2;
	wire w_dff_B_yKvtNNbC3_2;
	wire w_dff_B_nJLfIOD81_2;
	wire w_dff_B_XJEfy2eA2_2;
	wire w_dff_B_MjUiPWYF1_2;
	wire w_dff_B_2xI6hlF41_2;
	wire w_dff_B_rSF8CSo16_2;
	wire w_dff_B_W0mRZfbF5_2;
	wire w_dff_B_B6eRyLYW2_2;
	wire w_dff_B_kEoxd8r45_2;
	wire w_dff_B_DNoRZaMs0_2;
	wire w_dff_B_amQhJ1rp8_2;
	wire w_dff_B_hfBLVgxm8_2;
	wire w_dff_B_NJq9Mwmv8_2;
	wire w_dff_B_9rJcZFO74_2;
	wire w_dff_B_aLCONApw9_1;
	wire w_dff_B_eTKLcG3n9_2;
	wire w_dff_B_R6UHHqcU8_2;
	wire w_dff_B_hXhFr7N95_2;
	wire w_dff_B_NRLcLJR19_2;
	wire w_dff_B_dUEnkPYr7_2;
	wire w_dff_B_XLvcjCws7_2;
	wire w_dff_B_icyC7InA1_2;
	wire w_dff_B_Uqk8bYov4_2;
	wire w_dff_B_MpLiHoPy2_2;
	wire w_dff_B_F2gVclQR0_2;
	wire w_dff_B_DQ9DLNxE3_2;
	wire w_dff_B_F6QBbcuy4_2;
	wire w_dff_B_QjgN8iEH3_2;
	wire w_dff_B_7TsXYrYs6_2;
	wire w_dff_B_azhVPQdI9_2;
	wire w_dff_B_hbH2dvgo3_2;
	wire w_dff_B_9lYNUB6v6_2;
	wire w_dff_B_sWjd90256_2;
	wire w_dff_B_RHR0rDDN0_2;
	wire w_dff_B_myZc1rch3_1;
	wire w_dff_B_Wk0729rd9_2;
	wire w_dff_B_9j2TjyNq2_2;
	wire w_dff_B_0zH9w3kZ5_2;
	wire w_dff_B_hzUDXxsE8_2;
	wire w_dff_B_fDnBT49Y9_2;
	wire w_dff_B_AVfeqjyG7_2;
	wire w_dff_B_4BuUGYnX4_2;
	wire w_dff_B_mtqPUI0T1_2;
	wire w_dff_B_Mpp5fT8p6_2;
	wire w_dff_B_TViT5sPd4_2;
	wire w_dff_B_eQU8pXQN6_2;
	wire w_dff_B_hB9y8UTf7_2;
	wire w_dff_B_8lRcB4fm6_2;
	wire w_dff_B_aXuJiYt90_2;
	wire w_dff_B_N4qhkeI07_2;
	wire w_dff_B_rldC3BJ47_2;
	wire w_dff_B_JXDGhtOe4_1;
	wire w_dff_B_2RydlANO8_2;
	wire w_dff_B_CIScbIBQ6_2;
	wire w_dff_B_zH8a4xVO4_2;
	wire w_dff_B_sDahNV6J7_2;
	wire w_dff_B_94Su4Wyr7_2;
	wire w_dff_B_RRUJDn0M0_2;
	wire w_dff_B_PC0IDieh3_2;
	wire w_dff_B_Hd6Dvm0S6_2;
	wire w_dff_B_vnDs6X5n0_2;
	wire w_dff_B_SpKWs8qL6_2;
	wire w_dff_B_deIYh7Pd5_2;
	wire w_dff_B_StDSFw8h8_2;
	wire w_dff_B_CVnLg0kR4_2;
	wire w_dff_B_fr234X5Q7_1;
	wire w_dff_B_6tT9T7Su6_2;
	wire w_dff_B_Wqu20p4v5_2;
	wire w_dff_B_A8a4HFKX5_2;
	wire w_dff_B_nnvA88J42_2;
	wire w_dff_B_48uXmbWc9_2;
	wire w_dff_B_8H9EKZis3_2;
	wire w_dff_B_hIDVNv4n8_2;
	wire w_dff_B_wmccnfO15_2;
	wire w_dff_B_j23U0sOR6_2;
	wire w_dff_B_DENUeDNg6_2;
	wire w_dff_B_ugK7QYqi7_2;
	wire w_dff_B_MYapCTdd2_1;
	wire w_dff_B_xgmph9Mx5_1;
	wire w_dff_B_9kdLMMw17_1;
	wire w_dff_B_ou4UUd8m9_1;
	wire w_dff_B_Eg0G2rQK4_1;
	wire w_dff_B_zin7EFie7_1;
	wire w_dff_B_ayM6OZZT9_0;
	wire w_dff_B_L41QrBO30_0;
	wire w_dff_A_TmYr42cC0_0;
	wire w_dff_A_v2T2r6Bw5_0;
	wire w_dff_A_CFnGIAnQ4_0;
	wire w_dff_B_AuDEaiwK0_1;
	wire w_dff_A_CWv4PehF4_0;
	wire w_dff_A_PldyxTtr0_1;
	wire w_dff_A_IQZnHAAl3_1;
	wire w_dff_A_jlCOkuN10_1;
	wire w_dff_A_Vzuu0Vkz3_1;
	wire w_dff_A_5iOY39rK3_1;
	wire w_dff_A_fYxLTpdA0_1;
	wire w_dff_A_vkF2PkVD2_1;
	wire w_dff_A_AlngDwTI8_1;
	wire w_dff_B_tmATA0839_2;
	wire w_dff_B_qO9LQxKl1_2;
	wire w_dff_B_mP2VrqKQ6_1;
	wire w_dff_B_plqLQFNf4_2;
	wire w_dff_B_FSU4Fl4o1_2;
	wire w_dff_B_YCffW1NN1_2;
	wire w_dff_B_tnMY8Ikd0_2;
	wire w_dff_B_aRbZ0vuq7_2;
	wire w_dff_B_XjtbQkA16_2;
	wire w_dff_B_SZmuMXNF5_2;
	wire w_dff_B_8NpBifyg5_2;
	wire w_dff_B_EmYtTHYT5_2;
	wire w_dff_B_QWZjE07A5_2;
	wire w_dff_B_48xUDhoj6_2;
	wire w_dff_B_Yh5tGfSY6_2;
	wire w_dff_B_z2ELHyry4_2;
	wire w_dff_B_qW6Bg2YV3_2;
	wire w_dff_B_t36SaB8O2_2;
	wire w_dff_B_RKhaZqiF6_2;
	wire w_dff_B_knm0k8Xg4_2;
	wire w_dff_B_yEHtgwAw9_2;
	wire w_dff_B_CBPGj1Xr9_2;
	wire w_dff_B_wfNlrhA39_2;
	wire w_dff_B_XZWc1MA07_2;
	wire w_dff_B_tjYOlqZm1_2;
	wire w_dff_B_hELfrm557_2;
	wire w_dff_B_EeHt7nf20_2;
	wire w_dff_B_PUVktDH65_2;
	wire w_dff_B_e8tfmy4u5_2;
	wire w_dff_B_DE1T8EcF2_2;
	wire w_dff_B_DbnIVGSV5_2;
	wire w_dff_B_Semw6xyf3_2;
	wire w_dff_B_6HL6TPZi0_2;
	wire w_dff_B_dKWFuJb32_2;
	wire w_dff_B_tQwvjZBp2_2;
	wire w_dff_B_O3rmj7Hd0_2;
	wire w_dff_B_bSnaak8k2_2;
	wire w_dff_B_C3SRLnC69_2;
	wire w_dff_B_70Xy8b0j3_2;
	wire w_dff_B_zmavL6419_2;
	wire w_dff_B_0wlAA0ud1_2;
	wire w_dff_B_ow3Kdl3O0_2;
	wire w_dff_B_IXcVz9od3_2;
	wire w_dff_B_UIupoNSA5_2;
	wire w_dff_B_IxFvomfa6_2;
	wire w_dff_B_uivDMDmA9_2;
	wire w_dff_B_vJbzwzhe9_2;
	wire w_dff_B_y9QMcpst5_2;
	wire w_dff_B_KEC61UbN7_2;
	wire w_dff_B_4gjy0nN20_2;
	wire w_dff_B_ewia6aDz7_1;
	wire w_dff_B_SPXqW2dm1_2;
	wire w_dff_B_kTykYwNQ1_2;
	wire w_dff_B_OC4OnPtO3_2;
	wire w_dff_B_H1ekknui1_2;
	wire w_dff_B_ey9eU7cV7_2;
	wire w_dff_B_n7EoCFBQ3_2;
	wire w_dff_B_msYtl1oB4_2;
	wire w_dff_B_DhnOhXgm6_2;
	wire w_dff_B_hPp4pb6m3_2;
	wire w_dff_B_NcOOZW1C0_2;
	wire w_dff_B_H9TtCYDc6_2;
	wire w_dff_B_04DJ5N5p2_2;
	wire w_dff_B_1VzuVgi55_2;
	wire w_dff_B_jI0d8bc10_2;
	wire w_dff_B_W0I0efQf8_2;
	wire w_dff_B_w8oH05OQ2_2;
	wire w_dff_B_DCvcBuH23_2;
	wire w_dff_B_PQ9kNBfv0_2;
	wire w_dff_B_02MewigC3_2;
	wire w_dff_B_567YfJb48_2;
	wire w_dff_B_mv94IPBP5_2;
	wire w_dff_B_Rvyk1bc65_2;
	wire w_dff_B_u2ZuBt3E8_2;
	wire w_dff_B_4WU0sOu84_2;
	wire w_dff_B_nltW59Ju1_2;
	wire w_dff_B_1ZNXYIwD0_2;
	wire w_dff_B_o7z3vP909_2;
	wire w_dff_B_pZPftn4o4_2;
	wire w_dff_B_nROt5SIt4_2;
	wire w_dff_B_ivCzFx8c8_2;
	wire w_dff_B_D8shVlpO4_2;
	wire w_dff_B_HAGUHgsz6_2;
	wire w_dff_B_ASSS5cmR7_2;
	wire w_dff_B_B8QSHjaK1_2;
	wire w_dff_B_pBJ2Dndp1_2;
	wire w_dff_B_TnpgL7Sz4_2;
	wire w_dff_B_ZFryTQeT9_2;
	wire w_dff_B_vpmIoObM3_2;
	wire w_dff_B_7lS39wSh8_2;
	wire w_dff_B_t4TYKUIV5_2;
	wire w_dff_B_rG0GDWV04_2;
	wire w_dff_B_2Dc2Cqqv3_2;
	wire w_dff_B_DhnMH88a8_2;
	wire w_dff_B_t36JFZHW4_1;
	wire w_dff_B_W2D9LgdN6_2;
	wire w_dff_B_0WMAt5ZJ9_2;
	wire w_dff_B_27gtSKIT6_2;
	wire w_dff_B_2yeudNdz7_2;
	wire w_dff_B_mH2dwj8j0_2;
	wire w_dff_B_4ykKdkSo1_2;
	wire w_dff_B_YQPuyVSy9_2;
	wire w_dff_B_vRmFT9vW7_2;
	wire w_dff_B_AQ32ZqUO8_2;
	wire w_dff_B_NAzTCZhW0_2;
	wire w_dff_B_Xw5Zjdo61_2;
	wire w_dff_B_aHC6WF8t9_2;
	wire w_dff_B_hsBo7oyx7_2;
	wire w_dff_B_vl4HxP8H4_2;
	wire w_dff_B_AZ8Uq0Je9_2;
	wire w_dff_B_c77SKypD8_2;
	wire w_dff_B_4J9yUMTh4_2;
	wire w_dff_B_Kc4qZdze1_2;
	wire w_dff_B_FUUV2IFK0_2;
	wire w_dff_B_4IaHg2y39_2;
	wire w_dff_B_tSxKbDZx9_2;
	wire w_dff_B_XsHjt4T17_2;
	wire w_dff_B_zgWTXqDe3_2;
	wire w_dff_B_aQLIWByr2_2;
	wire w_dff_B_vjhBhKZL7_2;
	wire w_dff_B_15SdAugp4_2;
	wire w_dff_B_eZaSc35B2_2;
	wire w_dff_B_s0s7SrLJ2_2;
	wire w_dff_B_Pf8NYs0X7_2;
	wire w_dff_B_JS6VDofc4_2;
	wire w_dff_B_MxlpbtEz8_2;
	wire w_dff_B_ryAZhdJc6_2;
	wire w_dff_B_T8fmoYTS6_2;
	wire w_dff_B_XVlVHmCQ4_2;
	wire w_dff_B_RNOVQFcl9_2;
	wire w_dff_B_dgOO3eT99_2;
	wire w_dff_B_cHGSWxIC0_2;
	wire w_dff_B_p9L3JcAh3_2;
	wire w_dff_B_Gzmv50DE8_2;
	wire w_dff_B_A3R2VAa63_2;
	wire w_dff_B_NTWXxtiL6_1;
	wire w_dff_B_RNJJNCz87_2;
	wire w_dff_B_Ao0pvMLT7_2;
	wire w_dff_B_m5IhTBR80_2;
	wire w_dff_B_Fv0nOfa90_2;
	wire w_dff_B_rkybG2kM7_2;
	wire w_dff_B_l6mnBk3Z3_2;
	wire w_dff_B_WTfkTDFu1_2;
	wire w_dff_B_8PNFX68G2_2;
	wire w_dff_B_237ECkMK0_2;
	wire w_dff_B_iMGYnLzT3_2;
	wire w_dff_B_WUTQDFVG2_2;
	wire w_dff_B_ZjXT7OBx5_2;
	wire w_dff_B_kAhla4n08_2;
	wire w_dff_B_tomTPd9y1_2;
	wire w_dff_B_CfCdbbvS2_2;
	wire w_dff_B_3OUYU2I74_2;
	wire w_dff_B_pbxAkWNd0_2;
	wire w_dff_B_R5nBeBZ59_2;
	wire w_dff_B_QNOqrJ0A8_2;
	wire w_dff_B_MoKvDhTo5_2;
	wire w_dff_B_J7i9nfDu3_2;
	wire w_dff_B_TobCk7kL6_2;
	wire w_dff_B_xcs9joq36_2;
	wire w_dff_B_ZVqcZxM41_2;
	wire w_dff_B_P4niPtod4_2;
	wire w_dff_B_v92yHpEa5_2;
	wire w_dff_B_kfOIsyGW9_2;
	wire w_dff_B_1LofYttv4_2;
	wire w_dff_B_qrJBSzC89_2;
	wire w_dff_B_PB6FJwQ53_2;
	wire w_dff_B_MwzE1mE58_2;
	wire w_dff_B_7BAifTpZ3_2;
	wire w_dff_B_eRUPqLDn5_2;
	wire w_dff_B_gEpaOo1z1_2;
	wire w_dff_B_vJylCD1i2_2;
	wire w_dff_B_aVwQOu5d0_2;
	wire w_dff_B_1ibA4IKY8_2;
	wire w_dff_B_sP4Ejq843_1;
	wire w_dff_B_UPfBcQpT9_2;
	wire w_dff_B_Z5Iv1g5Q9_2;
	wire w_dff_B_jdLlyNxj6_2;
	wire w_dff_B_G4MVYnug1_2;
	wire w_dff_B_J4zpvQO48_2;
	wire w_dff_B_iXrriSKA5_2;
	wire w_dff_B_IML1f4pw4_2;
	wire w_dff_B_RCo6VYIV9_2;
	wire w_dff_B_Y0hH1vEO4_2;
	wire w_dff_B_nzvBuzoc2_2;
	wire w_dff_B_YeruEgU76_2;
	wire w_dff_B_LeEsOAyE2_2;
	wire w_dff_B_64IjW4vJ1_2;
	wire w_dff_B_sAwzFx3z9_2;
	wire w_dff_B_eP4KJ1Ce8_2;
	wire w_dff_B_cycacQty7_2;
	wire w_dff_B_C3SbwQnh2_2;
	wire w_dff_B_Eyqr2xo32_2;
	wire w_dff_B_HLctiEbA8_2;
	wire w_dff_B_EEFVhxNg0_2;
	wire w_dff_B_LOoSonQp4_2;
	wire w_dff_B_djsuKSzd7_2;
	wire w_dff_B_ZOROOSvj7_2;
	wire w_dff_B_95KqB4Id8_2;
	wire w_dff_B_KVdZoxK02_2;
	wire w_dff_B_LcUsYLLa3_2;
	wire w_dff_B_dFmMhxME2_2;
	wire w_dff_B_G4v4cB765_2;
	wire w_dff_B_txscnVFt6_2;
	wire w_dff_B_b0KI3EAq2_2;
	wire w_dff_B_5ndnb7647_2;
	wire w_dff_B_xTxfJX3d8_2;
	wire w_dff_B_7R0lN1O60_2;
	wire w_dff_B_gBIJsM8w9_2;
	wire w_dff_B_OV7ggkl04_1;
	wire w_dff_B_q7OUFDbZ9_2;
	wire w_dff_B_EdsKtupo0_2;
	wire w_dff_B_bbHw0lxs0_2;
	wire w_dff_B_Nj5M3Epq0_2;
	wire w_dff_B_oaFW9q362_2;
	wire w_dff_B_Gp1rMAbZ4_2;
	wire w_dff_B_tOq3sVn01_2;
	wire w_dff_B_o67CCh235_2;
	wire w_dff_B_MzV4yTXU7_2;
	wire w_dff_B_74rA2ppH0_2;
	wire w_dff_B_Aovb1Zli7_2;
	wire w_dff_B_T6WNXiWJ1_2;
	wire w_dff_B_RscgG0iQ7_2;
	wire w_dff_B_JnOtgfc76_2;
	wire w_dff_B_IxwqDl0d7_2;
	wire w_dff_B_8hqdvpSS9_2;
	wire w_dff_B_PeXW10J35_2;
	wire w_dff_B_9dZ3Len40_2;
	wire w_dff_B_5xM2FZkd0_2;
	wire w_dff_B_E1Fw6C7v8_2;
	wire w_dff_B_7Q8qCMYt1_2;
	wire w_dff_B_p90lf7R15_2;
	wire w_dff_B_zHe1xKuS3_2;
	wire w_dff_B_8ojM9xyx8_2;
	wire w_dff_B_rjS4bj6V0_2;
	wire w_dff_B_aruJWUHh6_2;
	wire w_dff_B_Y0cRz4VG2_2;
	wire w_dff_B_MhuYKNBv9_2;
	wire w_dff_B_EhXr46m92_2;
	wire w_dff_B_WTHNYiGv2_2;
	wire w_dff_B_lnYCOwVq2_2;
	wire w_dff_B_uzd3W8qA3_1;
	wire w_dff_B_xjj871zb0_2;
	wire w_dff_B_BZQu8nka9_2;
	wire w_dff_B_c8yZwTfn0_2;
	wire w_dff_B_yv4d6TTA5_2;
	wire w_dff_B_WDPk0vP99_2;
	wire w_dff_B_BtEugkbS4_2;
	wire w_dff_B_8CIlX0JD2_2;
	wire w_dff_B_vDtilpDP2_2;
	wire w_dff_B_b2SqLpvp0_2;
	wire w_dff_B_icSYXwrt0_2;
	wire w_dff_B_GTN6xiao0_2;
	wire w_dff_B_IkiyTq7T5_2;
	wire w_dff_B_sBy8yfAK0_2;
	wire w_dff_B_ayjmuoYy3_2;
	wire w_dff_B_c4HkXHup8_2;
	wire w_dff_B_ewLgdc4O5_2;
	wire w_dff_B_0rz40acQ1_2;
	wire w_dff_B_pDr0YIfu4_2;
	wire w_dff_B_ArYQ0XeZ8_2;
	wire w_dff_B_M7tjpi6J9_2;
	wire w_dff_B_K1ETa2s77_2;
	wire w_dff_B_dUA6h99e5_2;
	wire w_dff_B_YoWvCeLF3_2;
	wire w_dff_B_I2RdSUql2_2;
	wire w_dff_B_mGmdX3Wl9_2;
	wire w_dff_B_Aq25DpYO1_2;
	wire w_dff_B_0zxA06rf9_2;
	wire w_dff_B_xeE0Cf714_2;
	wire w_dff_B_Xewy7ynQ2_1;
	wire w_dff_B_ILqYK7GA6_2;
	wire w_dff_B_KefUfuQX2_2;
	wire w_dff_B_vbYQ3d9e6_2;
	wire w_dff_B_FxTI3rpf0_2;
	wire w_dff_B_eaz4wfXi4_2;
	wire w_dff_B_jHkGQAW51_2;
	wire w_dff_B_OsQFIn089_2;
	wire w_dff_B_yMkFgDtb4_2;
	wire w_dff_B_oxnhuztm1_2;
	wire w_dff_B_soxTaaV85_2;
	wire w_dff_B_PLudMCF56_2;
	wire w_dff_B_G3qFdKgE6_2;
	wire w_dff_B_ShZ6kQEh3_2;
	wire w_dff_B_ynNPUrKu4_2;
	wire w_dff_B_PPTnP7aQ2_2;
	wire w_dff_B_HmDCQnBm7_2;
	wire w_dff_B_snohWNGp8_2;
	wire w_dff_B_9o4564HU1_2;
	wire w_dff_B_fV8OAf4n9_2;
	wire w_dff_B_xzvpndms1_2;
	wire w_dff_B_cAiJ0cTE5_2;
	wire w_dff_B_LglNHTVx1_2;
	wire w_dff_B_AguJD1uK1_2;
	wire w_dff_B_jwFo8Crr7_2;
	wire w_dff_B_srM51NvW5_2;
	wire w_dff_B_KizjIKLD4_1;
	wire w_dff_B_kJbx6HmA4_2;
	wire w_dff_B_B2LcDPZV8_2;
	wire w_dff_B_VVtjfoL76_2;
	wire w_dff_B_D6V39gPe4_2;
	wire w_dff_B_I7fehIHE4_2;
	wire w_dff_B_Xv1jmA005_2;
	wire w_dff_B_AzezYvDp3_2;
	wire w_dff_B_Lfu3r4Qc2_2;
	wire w_dff_B_Vxrn0VrF8_2;
	wire w_dff_B_joRcfVxS5_2;
	wire w_dff_B_GIy6Ni797_2;
	wire w_dff_B_tEBNFMUf8_2;
	wire w_dff_B_aQAknhHc8_2;
	wire w_dff_B_C3FlaVdQ2_2;
	wire w_dff_B_4rN7hxPq4_2;
	wire w_dff_B_oStUWTwr1_2;
	wire w_dff_B_1FcR4dni7_2;
	wire w_dff_B_whimdm246_2;
	wire w_dff_B_kwEysLM92_2;
	wire w_dff_B_5f3kWY4S0_2;
	wire w_dff_B_kYkqdPMr6_2;
	wire w_dff_B_JcBbMAdb9_2;
	wire w_dff_B_c8K0u9p28_1;
	wire w_dff_B_HqPS48kr8_2;
	wire w_dff_B_JBOVN3QN0_2;
	wire w_dff_B_7TY5rIS07_2;
	wire w_dff_B_nP7lwz5r2_2;
	wire w_dff_B_e4hR2Ggt0_2;
	wire w_dff_B_wfs4P79U9_2;
	wire w_dff_B_AnLpgX643_2;
	wire w_dff_B_EPu3zuoE4_2;
	wire w_dff_B_jk0muqlY7_2;
	wire w_dff_B_Dbv7Pg6n5_2;
	wire w_dff_B_EM1pjMts4_2;
	wire w_dff_B_32uSxC0p3_2;
	wire w_dff_B_CRrFrIAr8_2;
	wire w_dff_B_T16sNmeR3_2;
	wire w_dff_B_j2u7iEnl2_2;
	wire w_dff_B_qVFpwbDJ5_2;
	wire w_dff_B_vIE5lVX17_2;
	wire w_dff_B_BcXpF4rI7_2;
	wire w_dff_B_FgF8KqwX0_2;
	wire w_dff_B_gkIHDYrP0_1;
	wire w_dff_B_KPE4BNW90_2;
	wire w_dff_B_IxD6OlcQ7_2;
	wire w_dff_B_Q6TigjFH5_2;
	wire w_dff_B_ORohxeBL6_2;
	wire w_dff_B_xfRwrgGu7_2;
	wire w_dff_B_JRz79APs0_2;
	wire w_dff_B_vI6OPqDp0_2;
	wire w_dff_B_VQPOLqxI8_2;
	wire w_dff_B_n3VJb7os0_2;
	wire w_dff_B_PXpKiGS69_2;
	wire w_dff_B_0NrkS6646_2;
	wire w_dff_B_JAffA4Ep7_2;
	wire w_dff_B_qZizcAE34_2;
	wire w_dff_B_Pec7xNWs6_2;
	wire w_dff_B_TGg6KFiC7_2;
	wire w_dff_B_4fGVicy57_2;
	wire w_dff_B_6qB0P92B1_1;
	wire w_dff_B_7blUpne13_2;
	wire w_dff_B_C4QfKUdZ7_2;
	wire w_dff_B_ekc50hko6_2;
	wire w_dff_B_LJBvSjCD6_2;
	wire w_dff_B_aK4zCiUF0_2;
	wire w_dff_B_4L345AdN8_2;
	wire w_dff_B_ieqWtctJ7_2;
	wire w_dff_B_jBAJX7Gd4_2;
	wire w_dff_B_27o1vert5_2;
	wire w_dff_B_emLOxp1V6_2;
	wire w_dff_B_FXgapH284_2;
	wire w_dff_B_DbqvFnC43_2;
	wire w_dff_B_oy8umolf6_2;
	wire w_dff_B_rAYAdfFl2_1;
	wire w_dff_B_ja1CMELV8_2;
	wire w_dff_B_5qSuCpD44_2;
	wire w_dff_B_f8f72HM14_2;
	wire w_dff_B_L2PET60S9_2;
	wire w_dff_B_4bgFc24M3_2;
	wire w_dff_B_dSKmSjOY5_2;
	wire w_dff_B_yx21GZjs0_2;
	wire w_dff_B_NnjONBx14_2;
	wire w_dff_B_aWyavlEF5_2;
	wire w_dff_B_CmShW5m65_2;
	wire w_dff_B_QiWXyrP18_2;
	wire w_dff_B_okGvTIfp4_1;
	wire w_dff_B_Ovga210J9_1;
	wire w_dff_B_cfkcpT9w5_1;
	wire w_dff_B_DNOyaLVM2_1;
	wire w_dff_B_N1MTUlbu6_1;
	wire w_dff_B_Oo0S0JvP8_1;
	wire w_dff_B_2LjfKZ2q1_0;
	wire w_dff_B_fzZDPGCA0_0;
	wire w_dff_A_uHGO6zZS9_0;
	wire w_dff_A_qXO6zwHi7_0;
	wire w_dff_A_PzvLBQM62_0;
	wire w_dff_B_kfrBW14e5_1;
	wire w_dff_A_OqaIikFK2_0;
	wire w_dff_A_OSxUYutW3_1;
	wire w_dff_A_RVoeUevc7_1;
	wire w_dff_A_teBB2hqj4_1;
	wire w_dff_A_tV7cHCuR6_1;
	wire w_dff_A_MwvqcJvR8_1;
	wire w_dff_A_i0ZkdQHk1_1;
	wire w_dff_A_WrFDIzY00_1;
	wire w_dff_A_mAPv3Wu33_1;
	wire w_dff_B_3RnJicDM9_2;
	wire w_dff_B_VVOCdBKQ9_1;
	wire w_dff_B_rQGk3lVe3_2;
	wire w_dff_B_H1sxGiWm9_2;
	wire w_dff_B_SJ3sHZQ76_2;
	wire w_dff_B_vdXYDhFr4_2;
	wire w_dff_B_gwD71AgJ4_2;
	wire w_dff_B_FLBhM1gE1_2;
	wire w_dff_B_k97zJxyz8_2;
	wire w_dff_B_TIjQOkkX5_2;
	wire w_dff_B_C9K4kJzr3_2;
	wire w_dff_B_N4ORJPVi3_2;
	wire w_dff_B_Z0giA0840_2;
	wire w_dff_B_MFFiOSBY4_2;
	wire w_dff_B_MANj7Cr24_2;
	wire w_dff_B_K50yHLw83_2;
	wire w_dff_B_04MGH8kK4_2;
	wire w_dff_B_yKcc2K6C6_2;
	wire w_dff_B_oUwf0fKg8_2;
	wire w_dff_B_BboUODOo8_2;
	wire w_dff_B_SHciex9f9_2;
	wire w_dff_B_OoS0rA8j2_2;
	wire w_dff_B_4lqdVSLO9_2;
	wire w_dff_B_46iNrCSM2_2;
	wire w_dff_B_SyTGHSIE7_2;
	wire w_dff_B_JsB3ySxS8_2;
	wire w_dff_B_t0h8V9m91_2;
	wire w_dff_B_jZQQWcrI5_2;
	wire w_dff_B_HGM76Mk49_2;
	wire w_dff_B_DjSDpkoM1_2;
	wire w_dff_B_dc9NxKfl2_2;
	wire w_dff_B_WnYEq7mm6_2;
	wire w_dff_B_6E6uATDr7_2;
	wire w_dff_B_nB2Qk6472_2;
	wire w_dff_B_eBpkP9O22_2;
	wire w_dff_B_RtIma7D91_2;
	wire w_dff_B_GGChZvOx8_2;
	wire w_dff_B_yeOGpDpF3_2;
	wire w_dff_B_zGTN5gvK3_2;
	wire w_dff_B_MxzjAqhn0_2;
	wire w_dff_B_bigACyS58_2;
	wire w_dff_B_cOGu1qVi3_2;
	wire w_dff_B_dLX3NpNs7_2;
	wire w_dff_B_z1i7qGpa8_2;
	wire w_dff_B_vFbDe1Cc7_2;
	wire w_dff_B_L0r0AVv03_2;
	wire w_dff_B_iJxvJt2Q7_2;
	wire w_dff_B_Hxpq3uqt4_2;
	wire w_dff_B_DRCkAmS47_2;
	wire w_dff_B_oshq8HRc1_2;
	wire w_dff_B_8udX8bne1_2;
	wire w_dff_B_rqcdsL8S1_1;
	wire w_dff_A_4JJX4vbh2_1;
	wire w_dff_B_caV1Uciq4_1;
	wire w_dff_B_00vZXMjC9_2;
	wire w_dff_B_OMYvfEqK5_2;
	wire w_dff_B_DsR74SI38_2;
	wire w_dff_B_2Knia5NI5_2;
	wire w_dff_B_T6O79sgf8_2;
	wire w_dff_B_z9TPqOtJ6_2;
	wire w_dff_B_6Fef7Z8Z2_2;
	wire w_dff_B_TRGcbW495_2;
	wire w_dff_B_Ue3RsntW9_2;
	wire w_dff_B_474AUWGh0_2;
	wire w_dff_B_ajBr2uW02_2;
	wire w_dff_B_fRCweLPu0_2;
	wire w_dff_B_I7lrImhF5_2;
	wire w_dff_B_2XBlZWlG4_2;
	wire w_dff_B_tKsrIPLH9_2;
	wire w_dff_B_ICsQXzqu8_2;
	wire w_dff_B_6QXffW1I2_2;
	wire w_dff_B_5Av5Qla75_2;
	wire w_dff_B_SGU9ONIy9_2;
	wire w_dff_B_AScHc9bz7_2;
	wire w_dff_B_rIh4aMwv5_2;
	wire w_dff_B_78i17mhF0_2;
	wire w_dff_B_ptYBTz6k8_2;
	wire w_dff_B_lIpR6Luf5_2;
	wire w_dff_B_sa5nhSK93_2;
	wire w_dff_B_9vYERfv13_2;
	wire w_dff_B_AmwdL0Gj9_2;
	wire w_dff_B_XJk98zk63_2;
	wire w_dff_B_mc0IQvLR4_2;
	wire w_dff_B_t9UkyfRx6_2;
	wire w_dff_B_rxn0rczN1_2;
	wire w_dff_B_HQz4GrLV4_2;
	wire w_dff_B_P6z2MrgN2_2;
	wire w_dff_B_Q3l6Dwu72_2;
	wire w_dff_B_TQORNAjw3_2;
	wire w_dff_B_Ni5NJVNp1_2;
	wire w_dff_B_oLOv9SCj5_2;
	wire w_dff_B_ue0jFElA2_2;
	wire w_dff_B_4Jvsh2GY7_2;
	wire w_dff_B_lo3ZEi1K0_2;
	wire w_dff_B_lc7UO8933_2;
	wire w_dff_B_svI6uF3k7_2;
	wire w_dff_B_zYjooRPh7_2;
	wire w_dff_B_rKUlpOpo5_2;
	wire w_dff_B_OVFaeoJQ4_1;
	wire w_dff_B_dxyA2MqL0_2;
	wire w_dff_B_F0NMUvbu7_2;
	wire w_dff_B_jMvfmP3p5_2;
	wire w_dff_B_q5vBtwrN5_2;
	wire w_dff_B_AwtR4eou3_2;
	wire w_dff_B_q1W5I5cG8_2;
	wire w_dff_B_8DqNIZRW2_2;
	wire w_dff_B_dtoVpleY8_2;
	wire w_dff_B_KpsN6g3A3_2;
	wire w_dff_B_UUpkqryu9_2;
	wire w_dff_B_Z0mBabTw8_2;
	wire w_dff_B_70Vadccr9_2;
	wire w_dff_B_BkAydNWi0_2;
	wire w_dff_B_Kc7AVJjm8_2;
	wire w_dff_B_QoXqCVU15_2;
	wire w_dff_B_RkQ1Wc8J6_2;
	wire w_dff_B_KsuwzJpz1_2;
	wire w_dff_B_aEWQcq2K0_2;
	wire w_dff_B_TdSHs97D6_2;
	wire w_dff_B_ojYdJ6xP7_2;
	wire w_dff_B_2aqGnBmB3_2;
	wire w_dff_B_BY9jdHMx3_2;
	wire w_dff_B_G75FPiZ94_2;
	wire w_dff_B_KH1bkfDM3_2;
	wire w_dff_B_ZCw7RZE63_2;
	wire w_dff_B_O5R55zZc6_2;
	wire w_dff_B_CltihA214_2;
	wire w_dff_B_NFs8nu665_2;
	wire w_dff_B_dA59S4zW5_2;
	wire w_dff_B_wZS7RfwH9_2;
	wire w_dff_B_ekZVA6Pp4_2;
	wire w_dff_B_qDnt8Nwe4_2;
	wire w_dff_B_5gyJeHCz5_2;
	wire w_dff_B_7IOPICYw1_2;
	wire w_dff_B_3b8WpZfL0_2;
	wire w_dff_B_YnabyG0G3_2;
	wire w_dff_B_n77vf1nt9_2;
	wire w_dff_B_Vm42VOx80_2;
	wire w_dff_B_m0eMMI8i3_2;
	wire w_dff_B_ep9J85lm5_1;
	wire w_dff_B_NITjvwZO1_2;
	wire w_dff_B_pp1IcoEZ3_2;
	wire w_dff_B_yCg6xIBm2_2;
	wire w_dff_B_AXH3ceeX4_2;
	wire w_dff_B_hBxhxHyA9_2;
	wire w_dff_B_2VNxjfxP7_2;
	wire w_dff_B_jUKy0EVc6_2;
	wire w_dff_B_pVmGhPvx3_2;
	wire w_dff_B_uKayVfot0_2;
	wire w_dff_B_vvfc7eE66_2;
	wire w_dff_B_5hX1zHPV4_2;
	wire w_dff_B_dcXSkwkr4_2;
	wire w_dff_B_wirYtMQL7_2;
	wire w_dff_B_o6umcOOP8_2;
	wire w_dff_B_d9CUyejE7_2;
	wire w_dff_B_L8ISDlfd1_2;
	wire w_dff_B_j1J6srgp4_2;
	wire w_dff_B_VQnKRV0Y2_2;
	wire w_dff_B_rhduM2fl6_2;
	wire w_dff_B_lG6L7IyP0_2;
	wire w_dff_B_I4ezPKmf1_2;
	wire w_dff_B_I5Mn5VT17_2;
	wire w_dff_B_63fQgczl7_2;
	wire w_dff_B_stByCNqY7_2;
	wire w_dff_B_PQDJDI380_2;
	wire w_dff_B_zFRQ0nHT0_2;
	wire w_dff_B_ErKhzT9D7_2;
	wire w_dff_B_yXmbOzmP5_2;
	wire w_dff_B_T5upasdN9_2;
	wire w_dff_B_JtUGBNnw2_2;
	wire w_dff_B_hI6yFXJz7_2;
	wire w_dff_B_PNQIdWr74_2;
	wire w_dff_B_wjpq9D6j9_2;
	wire w_dff_B_vRvr2wr26_2;
	wire w_dff_B_Nk3AB6I91_2;
	wire w_dff_B_2ywxSxKj8_2;
	wire w_dff_B_HISQ8N1N8_2;
	wire w_dff_B_bc8EOeQJ5_1;
	wire w_dff_B_9dobeQkJ7_2;
	wire w_dff_B_jyVHoDC70_2;
	wire w_dff_B_m7F28Hkb4_2;
	wire w_dff_B_eMQ3XJKt9_2;
	wire w_dff_B_fTpM45iT8_2;
	wire w_dff_B_hhwn8Kaf2_2;
	wire w_dff_B_1gBks4D78_2;
	wire w_dff_B_EUu8PYPN4_2;
	wire w_dff_B_dRIsLWDc5_2;
	wire w_dff_B_okH6juCc3_2;
	wire w_dff_B_HZpdYgyn7_2;
	wire w_dff_B_Pj4hLcsP1_2;
	wire w_dff_B_NYENvobe8_2;
	wire w_dff_B_wzcWJJa17_2;
	wire w_dff_B_Y17Tzvel4_2;
	wire w_dff_B_OAL4d9VV7_2;
	wire w_dff_B_uFMc3xi21_2;
	wire w_dff_B_1CWtZyUO2_2;
	wire w_dff_B_6sOJFOLV6_2;
	wire w_dff_B_PLWr5jKS6_2;
	wire w_dff_B_74DTXMSh3_2;
	wire w_dff_B_ajl8NgPG4_2;
	wire w_dff_B_fMU1GJRk7_2;
	wire w_dff_B_hoNMd5JW0_2;
	wire w_dff_B_Yn3XMZPW3_2;
	wire w_dff_B_muVvpKeL8_2;
	wire w_dff_B_ownsU5WY6_2;
	wire w_dff_B_KaOcZpno8_2;
	wire w_dff_B_X3GzVAcQ1_2;
	wire w_dff_B_0u3Qh3XZ2_2;
	wire w_dff_B_5S0Pu4gx2_2;
	wire w_dff_B_gtqgsyJ29_2;
	wire w_dff_B_ytPP6zC89_2;
	wire w_dff_B_1JzL5Mq57_2;
	wire w_dff_B_WVn4gxIs4_1;
	wire w_dff_B_ip10Dipr1_2;
	wire w_dff_B_F6lJWV9g8_2;
	wire w_dff_B_ZeC5lp6w7_2;
	wire w_dff_B_Fe3noJUt0_2;
	wire w_dff_B_6rMTpEze6_2;
	wire w_dff_B_iHGDDPCs5_2;
	wire w_dff_B_qAzHfZTW8_2;
	wire w_dff_B_toU4PPUN8_2;
	wire w_dff_B_ncnBoFdE2_2;
	wire w_dff_B_skqtymb74_2;
	wire w_dff_B_0VPZXGuf9_2;
	wire w_dff_B_YBZzA1aF4_2;
	wire w_dff_B_apHUwt5q6_2;
	wire w_dff_B_9iGDo3O46_2;
	wire w_dff_B_iAabzOLN2_2;
	wire w_dff_B_64YivDpv3_2;
	wire w_dff_B_GIcp11qT1_2;
	wire w_dff_B_Rr24kxsg3_2;
	wire w_dff_B_oxBHb8iV9_2;
	wire w_dff_B_BEKKcG2v0_2;
	wire w_dff_B_uM1nMhGN2_2;
	wire w_dff_B_Z3txKOzB0_2;
	wire w_dff_B_NsuF8KsE1_2;
	wire w_dff_B_SAvm11bq7_2;
	wire w_dff_B_L8G6ABRI2_2;
	wire w_dff_B_oFuVGFgH8_2;
	wire w_dff_B_eFMZsobE9_2;
	wire w_dff_B_2YLg9TQ78_2;
	wire w_dff_B_T1HO2Rd15_2;
	wire w_dff_B_7zpv10YT7_2;
	wire w_dff_B_mADqmqP18_2;
	wire w_dff_B_nwJXkFV64_1;
	wire w_dff_B_LiWGV6py7_2;
	wire w_dff_B_We4PU8jH9_2;
	wire w_dff_B_lcrIB0qU5_2;
	wire w_dff_B_cjjx011v3_2;
	wire w_dff_B_rrpxWGx76_2;
	wire w_dff_B_zWgXi6xT9_2;
	wire w_dff_B_eAkQYT9l8_2;
	wire w_dff_B_K8jmrcin0_2;
	wire w_dff_B_Uqjnyzse5_2;
	wire w_dff_B_2fxMLfWK8_2;
	wire w_dff_B_jAXTuAWY0_2;
	wire w_dff_B_WrljdxqX4_2;
	wire w_dff_B_G8Sh7LQa3_2;
	wire w_dff_B_VyJhSFsX7_2;
	wire w_dff_B_n4fjb4Hx4_2;
	wire w_dff_B_ctJpDmhB3_2;
	wire w_dff_B_dKvI9GS99_2;
	wire w_dff_B_kzUkZZI13_2;
	wire w_dff_B_7ZeqhotU4_2;
	wire w_dff_B_FgEaB1x25_2;
	wire w_dff_B_M6ZF9rCk4_2;
	wire w_dff_B_mRnJoWnI9_2;
	wire w_dff_B_uCuvAqPS5_2;
	wire w_dff_B_aZ27IuzA5_2;
	wire w_dff_B_x8ueRvEL4_2;
	wire w_dff_B_V7vgzhww6_2;
	wire w_dff_B_44hlovNk6_2;
	wire w_dff_B_MsvinaVe8_2;
	wire w_dff_B_k0AmojMX2_1;
	wire w_dff_B_dBxrUPST0_2;
	wire w_dff_B_6FQvDauU0_2;
	wire w_dff_B_On3kuz2s7_2;
	wire w_dff_B_i4PD0MDB5_2;
	wire w_dff_B_ZAyC6yzB2_2;
	wire w_dff_B_ACqCUdJK3_2;
	wire w_dff_B_7wAoJzCG3_2;
	wire w_dff_B_5imdgR868_2;
	wire w_dff_B_ezW95HMd0_2;
	wire w_dff_B_2hjVwVmF8_2;
	wire w_dff_B_QBlXEqT10_2;
	wire w_dff_B_uAyDHpfw6_2;
	wire w_dff_B_zMbHL9B32_2;
	wire w_dff_B_598SblUx5_2;
	wire w_dff_B_FFHcRYqL3_2;
	wire w_dff_B_xkdNef0i0_2;
	wire w_dff_B_mKinpzrY2_2;
	wire w_dff_B_sVlZZoUM2_2;
	wire w_dff_B_wizdV6E65_2;
	wire w_dff_B_WmzQRrq68_2;
	wire w_dff_B_RfEcLeU20_2;
	wire w_dff_B_hpnRPkPl8_2;
	wire w_dff_B_BOHMR4jD0_2;
	wire w_dff_B_zmFlblHR9_2;
	wire w_dff_B_ArKrp9Jo9_2;
	wire w_dff_B_IHPr1Lw29_1;
	wire w_dff_B_tXrxXVHm9_2;
	wire w_dff_B_MrHLKQ150_2;
	wire w_dff_B_ibuG9Ba73_2;
	wire w_dff_B_naOkVaFF0_2;
	wire w_dff_B_UTSv0xFq2_2;
	wire w_dff_B_H2a9u2ng7_2;
	wire w_dff_B_ERHndalF5_2;
	wire w_dff_B_q2HbTIzh3_2;
	wire w_dff_B_wrcCZKqo9_2;
	wire w_dff_B_ZDwDkWAI9_2;
	wire w_dff_B_HWroxUo33_2;
	wire w_dff_B_g1Lf0It04_2;
	wire w_dff_B_e6WgFQ6R8_2;
	wire w_dff_B_kpoUAvar0_2;
	wire w_dff_B_5xcht1sV5_2;
	wire w_dff_B_LIuaEXWL2_2;
	wire w_dff_B_JpvsrTgi6_2;
	wire w_dff_B_j5B9MQpc4_2;
	wire w_dff_B_0d3qYfrT5_2;
	wire w_dff_B_NlFy0QL04_2;
	wire w_dff_B_AU6jyrFE3_2;
	wire w_dff_B_hOikBsCD4_2;
	wire w_dff_B_xA5TsFm41_1;
	wire w_dff_B_5Xu7gypW2_2;
	wire w_dff_B_VbfjyOeY5_2;
	wire w_dff_B_rPfXnYEv0_2;
	wire w_dff_B_Whxa2VIo9_2;
	wire w_dff_B_JbtUBMFH5_2;
	wire w_dff_B_eCibOGKe4_2;
	wire w_dff_B_SofNfQdv7_2;
	wire w_dff_B_DxpG3HVZ7_2;
	wire w_dff_B_UMPJEe397_2;
	wire w_dff_B_DEN1JuF13_2;
	wire w_dff_B_SvVeqdPa7_2;
	wire w_dff_B_jwUptlux1_2;
	wire w_dff_B_WFlrYD1e1_2;
	wire w_dff_B_jiy5FE7l9_2;
	wire w_dff_B_BeVZ6VZy0_2;
	wire w_dff_B_hipvSVQU7_2;
	wire w_dff_B_LkHXZCBK7_2;
	wire w_dff_B_pfabGU1z4_2;
	wire w_dff_B_n9EISm401_2;
	wire w_dff_B_HJQyML745_1;
	wire w_dff_B_wQfdFuV10_2;
	wire w_dff_B_o73wuKI98_2;
	wire w_dff_B_wmM4FHRy8_2;
	wire w_dff_B_3FrgMzfP3_2;
	wire w_dff_B_zzCFyGPl5_2;
	wire w_dff_B_CTrWC2XS6_2;
	wire w_dff_B_7bFV2QGw0_2;
	wire w_dff_B_NeFY834T1_2;
	wire w_dff_B_7VkI8jLT7_2;
	wire w_dff_B_i1IxUYqg2_2;
	wire w_dff_B_knIISLSD0_2;
	wire w_dff_B_lARREP0g7_2;
	wire w_dff_B_g7j7Yk6r6_2;
	wire w_dff_B_XkKe7h4n6_2;
	wire w_dff_B_dOQjWle73_2;
	wire w_dff_B_yEpiPgRN8_2;
	wire w_dff_B_bSQO3Iix9_1;
	wire w_dff_B_KbwQes492_2;
	wire w_dff_B_IXmf1d398_2;
	wire w_dff_B_ix1OoRRr9_2;
	wire w_dff_B_uCJoVFSw0_2;
	wire w_dff_B_5xjfZ3Wp0_2;
	wire w_dff_B_X1viEgLQ7_2;
	wire w_dff_B_YuiNqHBZ8_2;
	wire w_dff_B_YOyAP99l4_2;
	wire w_dff_B_Uk4p2vjt6_2;
	wire w_dff_B_oQsncDie8_2;
	wire w_dff_B_PqihfLAO8_2;
	wire w_dff_B_7W6IBFpX8_2;
	wire w_dff_B_Q5STwsBo3_2;
	wire w_dff_B_vavzs6245_1;
	wire w_dff_B_uFybdbnK0_2;
	wire w_dff_B_0LVi9f7f4_2;
	wire w_dff_B_ZR15t9k95_2;
	wire w_dff_B_uoKljbTd4_2;
	wire w_dff_B_GalnD0kl1_2;
	wire w_dff_B_ykNEyVAn8_2;
	wire w_dff_B_WjD1AETW3_2;
	wire w_dff_B_bsuqZ2859_2;
	wire w_dff_B_jZe4YHWU3_2;
	wire w_dff_B_OhS1WdKY6_2;
	wire w_dff_B_Y11zjUIr9_2;
	wire w_dff_B_2NBhPVEo0_1;
	wire w_dff_B_yhRwLhSl0_1;
	wire w_dff_B_h5csbh3Q4_1;
	wire w_dff_B_A6id4RZi6_1;
	wire w_dff_B_tz6VrQ7D8_1;
	wire w_dff_B_CbMh0etk8_1;
	wire w_dff_B_clarPqnr6_0;
	wire w_dff_B_5EYqdB1x0_0;
	wire w_dff_A_yizNcz2A1_0;
	wire w_dff_A_sFCCDAuD8_0;
	wire w_dff_A_BnbUiBaX3_0;
	wire w_dff_B_pIrr73m08_1;
	wire w_dff_A_VEjDMFPq4_0;
	wire w_dff_A_SAfrAM5U4_1;
	wire w_dff_A_DzAcwloZ4_1;
	wire w_dff_A_ajZXznoi4_1;
	wire w_dff_A_2oHCCgGu6_1;
	wire w_dff_A_BK8X57VK0_1;
	wire w_dff_A_PbKr4Kqu4_1;
	wire w_dff_A_0GWR2Htb6_1;
	wire w_dff_A_6STtgGwI6_1;
	wire w_dff_B_TCewL5c97_1;
	wire w_dff_A_gs11IcZb5_1;
	wire w_dff_B_ZNA61zx23_1;
	wire w_dff_B_TkY1yLGK6_2;
	wire w_dff_B_diW2C7mX8_2;
	wire w_dff_B_rE5T2yVe7_2;
	wire w_dff_B_CS8zggMj5_2;
	wire w_dff_B_b2mo3lKz6_2;
	wire w_dff_B_KLT5Lpxt9_2;
	wire w_dff_B_b3FesVu59_2;
	wire w_dff_B_Ph3YzaFY7_2;
	wire w_dff_B_ANayHqti9_2;
	wire w_dff_B_4JXILDJZ6_2;
	wire w_dff_B_CfMFsKap0_2;
	wire w_dff_B_RWGSRGPx5_2;
	wire w_dff_B_9K3JBp0j7_2;
	wire w_dff_B_zJqTLJr99_2;
	wire w_dff_B_99CbURTR4_2;
	wire w_dff_B_GI3UMVU34_2;
	wire w_dff_B_5KSbgHdb9_2;
	wire w_dff_B_eGCNUpTC8_2;
	wire w_dff_B_bu3eTSlq2_2;
	wire w_dff_B_9otfr0AT1_2;
	wire w_dff_B_eh42FrmY0_2;
	wire w_dff_B_rawarsQ76_2;
	wire w_dff_B_FgThDuMj4_2;
	wire w_dff_B_vGmS6IKl5_2;
	wire w_dff_B_0C2ytVHC6_2;
	wire w_dff_B_Jq9SG4xc0_2;
	wire w_dff_B_fmhu7x7C5_2;
	wire w_dff_B_rWFzzuz68_2;
	wire w_dff_B_F5bXzkmW5_2;
	wire w_dff_B_n9uHyAWm4_2;
	wire w_dff_B_UWOLfndn8_2;
	wire w_dff_B_oXm7oNef5_2;
	wire w_dff_B_CBNzjB7B2_2;
	wire w_dff_B_Syiaelsg1_2;
	wire w_dff_B_3zQJlg3H0_2;
	wire w_dff_B_JI51UZ669_2;
	wire w_dff_B_vzn2Bcph8_2;
	wire w_dff_B_ppiBzVLm1_2;
	wire w_dff_B_Mftj1Eta7_2;
	wire w_dff_B_O4UpiI2e8_2;
	wire w_dff_B_eRtSiULM4_2;
	wire w_dff_B_aspaOuBq0_2;
	wire w_dff_B_9a1SXeoi0_2;
	wire w_dff_B_lWuhQ7km8_2;
	wire w_dff_B_yP0Jf2nB5_2;
	wire w_dff_B_JNbSNTFf9_2;
	wire w_dff_B_mAJPjSWK4_2;
	wire w_dff_B_tcULOzcr5_2;
	wire w_dff_B_1pDKIZ093_2;
	wire w_dff_B_N2jdzGk90_2;
	wire w_dff_B_OD8zsOFz3_1;
	wire w_dff_B_Le2aNLXW1_2;
	wire w_dff_B_X940kKQk4_2;
	wire w_dff_B_WQWOCGvC2_2;
	wire w_dff_B_KKy3QRSz1_2;
	wire w_dff_B_Dbr6G2PZ9_2;
	wire w_dff_B_G0ADHMuC9_2;
	wire w_dff_B_oEcDhbXk8_2;
	wire w_dff_B_l0jqOEwI9_2;
	wire w_dff_B_NZYnER997_2;
	wire w_dff_B_9eFXj9rZ8_2;
	wire w_dff_B_lATkhR9x2_2;
	wire w_dff_B_fjW11Uiw8_2;
	wire w_dff_B_AWWjL4iO7_2;
	wire w_dff_B_9zkz70Iy8_2;
	wire w_dff_B_4JdnowO17_2;
	wire w_dff_B_PFUZM9UN2_2;
	wire w_dff_B_eNZAHqET7_2;
	wire w_dff_B_23GPd94w8_2;
	wire w_dff_B_U06PEwPw6_2;
	wire w_dff_B_svnKd5Hb2_2;
	wire w_dff_B_WolfQb4C1_2;
	wire w_dff_B_8sef5ni97_2;
	wire w_dff_B_COQEwRTS3_2;
	wire w_dff_B_eNKHHtb45_2;
	wire w_dff_B_vZM6LUyC7_2;
	wire w_dff_B_O9ovA19C0_2;
	wire w_dff_B_0ayl8ijC5_2;
	wire w_dff_B_B3NPte5y2_2;
	wire w_dff_B_pkTmhiov8_2;
	wire w_dff_B_bU4njUtF6_2;
	wire w_dff_B_h9EIukWF0_2;
	wire w_dff_B_Qh8KRF7c1_2;
	wire w_dff_B_MdxlzSYs3_2;
	wire w_dff_B_5ocVLUiB6_2;
	wire w_dff_B_qwmLDYlS5_2;
	wire w_dff_B_K8LkMMUf4_2;
	wire w_dff_B_3QpEcBYS5_2;
	wire w_dff_B_B68IbSmN4_2;
	wire w_dff_B_q2UG8rry9_2;
	wire w_dff_B_GWmTiUBi7_2;
	wire w_dff_B_6czhGHEI7_2;
	wire w_dff_B_0dWJxbfB1_2;
	wire w_dff_B_Wiglwtz19_2;
	wire w_dff_B_e4hHRO710_2;
	wire w_dff_B_t7NTSo022_2;
	wire w_dff_B_gEWZXbi90_2;
	wire w_dff_B_4DM503qx1_1;
	wire w_dff_B_XSj0W33P0_2;
	wire w_dff_B_mF69VJTT3_2;
	wire w_dff_B_ucASIHuc0_2;
	wire w_dff_B_Qftq9QV42_2;
	wire w_dff_B_et16hyLE3_2;
	wire w_dff_B_9Nd1Zc0o6_2;
	wire w_dff_B_QzZVqoBh7_2;
	wire w_dff_B_IkSMX9aT1_2;
	wire w_dff_B_vQHBgyYe9_2;
	wire w_dff_B_vvAv7Okf5_2;
	wire w_dff_B_5e5HsEMC4_2;
	wire w_dff_B_pEBgNAwd1_2;
	wire w_dff_B_Vuefmv1m0_2;
	wire w_dff_B_COoAiAtz7_2;
	wire w_dff_B_DnnAyAKx2_2;
	wire w_dff_B_muPSitCL1_2;
	wire w_dff_B_muLNuAq94_2;
	wire w_dff_B_CAX2kDuR4_2;
	wire w_dff_B_TWbd1d8b4_2;
	wire w_dff_B_JI8RnBij7_2;
	wire w_dff_B_p95ohL3o8_2;
	wire w_dff_B_TxH64Jd20_2;
	wire w_dff_B_vlsk8rsp8_2;
	wire w_dff_B_HWi3T1sR2_2;
	wire w_dff_B_syxz5Bew5_2;
	wire w_dff_B_ViomdNKI7_2;
	wire w_dff_B_B2IHkcjU0_2;
	wire w_dff_B_JFXiRL2v5_2;
	wire w_dff_B_qnOSOI3J0_2;
	wire w_dff_B_o0aGfLs23_2;
	wire w_dff_B_2ZGwtNOI0_2;
	wire w_dff_B_oYfWgQwj4_2;
	wire w_dff_B_vrHRwwY64_2;
	wire w_dff_B_w6MhnlCF4_2;
	wire w_dff_B_dLFBpsyn4_2;
	wire w_dff_B_lOrcylcN4_2;
	wire w_dff_B_NTf9Cb4h1_2;
	wire w_dff_B_1xK1Vb336_2;
	wire w_dff_B_k00PbxRh3_2;
	wire w_dff_B_shqddaeU0_2;
	wire w_dff_B_PlW01fJO6_2;
	wire w_dff_B_k6Z3dM301_2;
	wire w_dff_B_KWsj1w4I1_1;
	wire w_dff_B_fnADqmUn2_2;
	wire w_dff_B_HtyjzvXR0_2;
	wire w_dff_B_niEEAyfw3_2;
	wire w_dff_B_nkqB8I3H3_2;
	wire w_dff_B_MBEf3onO7_2;
	wire w_dff_B_xExIR2Qf8_2;
	wire w_dff_B_ZZj8lqqf6_2;
	wire w_dff_B_wDnhVLNH7_2;
	wire w_dff_B_N5r9Gnzo9_2;
	wire w_dff_B_dFgESHhn5_2;
	wire w_dff_B_I5XpsT1x0_2;
	wire w_dff_B_qxrLQuA97_2;
	wire w_dff_B_TwS7Su2d1_2;
	wire w_dff_B_TI4D2na19_2;
	wire w_dff_B_wdtrvRXi8_2;
	wire w_dff_B_GE6M4kkh9_2;
	wire w_dff_B_1v9xkd8r2_2;
	wire w_dff_B_c8p1SSMr9_2;
	wire w_dff_B_rG8uYtic6_2;
	wire w_dff_B_G2qFkAGH0_2;
	wire w_dff_B_BmlNWpeI1_2;
	wire w_dff_B_8s4SRJPV3_2;
	wire w_dff_B_hxYpHBWI4_2;
	wire w_dff_B_iqOqpiti7_2;
	wire w_dff_B_1ap5ySk98_2;
	wire w_dff_B_ThBV1DCF0_2;
	wire w_dff_B_7iAodSeq2_2;
	wire w_dff_B_wopjOCEN2_2;
	wire w_dff_B_1WI3EKo63_2;
	wire w_dff_B_NR4hBKQh4_2;
	wire w_dff_B_G5gHnXfc5_2;
	wire w_dff_B_QN5lWEbu1_2;
	wire w_dff_B_hL6rvXJP4_2;
	wire w_dff_B_Xcz8bQt79_2;
	wire w_dff_B_lrITYiHD2_2;
	wire w_dff_B_BHbMM9XM6_2;
	wire w_dff_B_2q0oM0jv1_2;
	wire w_dff_B_f4y5ryhm3_2;
	wire w_dff_B_QlXDA0Gs6_1;
	wire w_dff_B_HFuURorS5_2;
	wire w_dff_B_HYtwev9K1_2;
	wire w_dff_B_jsr3QjnB4_2;
	wire w_dff_B_KLGBzTgE6_2;
	wire w_dff_B_6ChZadHj3_2;
	wire w_dff_B_UbqCyEjC9_2;
	wire w_dff_B_Hhwahzwe4_2;
	wire w_dff_B_2iJvjgP80_2;
	wire w_dff_B_0rAaLXo55_2;
	wire w_dff_B_WKRz6zFz4_2;
	wire w_dff_B_mYj8hEJG2_2;
	wire w_dff_B_2tDofd421_2;
	wire w_dff_B_BrDCQca44_2;
	wire w_dff_B_ovWFeDIW3_2;
	wire w_dff_B_UFvFRXVG7_2;
	wire w_dff_B_dWjQTx6d2_2;
	wire w_dff_B_Z1pQawyx2_2;
	wire w_dff_B_2Mws1gYY1_2;
	wire w_dff_B_tviATJVO9_2;
	wire w_dff_B_GTeB3NYr8_2;
	wire w_dff_B_Y6j6lNRV8_2;
	wire w_dff_B_unFGG66d8_2;
	wire w_dff_B_7aIpXPD49_2;
	wire w_dff_B_V2ISwFEN5_2;
	wire w_dff_B_LJw5olb82_2;
	wire w_dff_B_Fx76HhxW5_2;
	wire w_dff_B_0u5xo9Bq9_2;
	wire w_dff_B_GmD0ky7j3_2;
	wire w_dff_B_n9K19JA90_2;
	wire w_dff_B_fMOdFGYu5_2;
	wire w_dff_B_y2k1Dz5Y5_2;
	wire w_dff_B_ogX3M0e88_2;
	wire w_dff_B_NIiP5MnK3_2;
	wire w_dff_B_0Ke26RMA9_1;
	wire w_dff_B_zdur0rHx6_2;
	wire w_dff_B_NHoRZHjM0_2;
	wire w_dff_B_8SYQqcns8_2;
	wire w_dff_B_YBcxg5414_2;
	wire w_dff_B_erQ4fIHP6_2;
	wire w_dff_B_4PuvGxbi5_2;
	wire w_dff_B_HMFb1ltr6_2;
	wire w_dff_B_Ife0iku81_2;
	wire w_dff_B_f8cjXL9Z2_2;
	wire w_dff_B_UiOIbgrz5_2;
	wire w_dff_B_7jUvcbn46_2;
	wire w_dff_B_EVeQGmWW3_2;
	wire w_dff_B_H9Ffuray3_2;
	wire w_dff_B_3akg4uhZ2_2;
	wire w_dff_B_qlAL7DbF5_2;
	wire w_dff_B_rcyTbpPx5_2;
	wire w_dff_B_Egp1LORW2_2;
	wire w_dff_B_W59M4nOI8_2;
	wire w_dff_B_bxryLyCT7_2;
	wire w_dff_B_7WUGfm5W9_2;
	wire w_dff_B_4Lb1V7ce6_2;
	wire w_dff_B_VoDIUlxA7_2;
	wire w_dff_B_XTgZh5318_2;
	wire w_dff_B_CL2iF2yL3_2;
	wire w_dff_B_k9owATDD3_2;
	wire w_dff_B_iyU4cppo5_2;
	wire w_dff_B_MsQzurds4_2;
	wire w_dff_B_TTTi2UUd8_2;
	wire w_dff_B_WJEV09jc6_2;
	wire w_dff_B_iqpIQTzU2_2;
	wire w_dff_B_2gb9Bxer1_2;
	wire w_dff_B_jkB5FMPY5_1;
	wire w_dff_B_EHNiVPGa5_2;
	wire w_dff_B_R53KKUYP0_2;
	wire w_dff_B_cZjVBzQE5_2;
	wire w_dff_B_4j4JNBkS9_2;
	wire w_dff_B_qudDM4mX8_2;
	wire w_dff_B_I2hQy2mV6_2;
	wire w_dff_B_GUVxetKd4_2;
	wire w_dff_B_WlH3N3xI3_2;
	wire w_dff_B_qaD0liny8_2;
	wire w_dff_B_pskPLXQP5_2;
	wire w_dff_B_RY5mHMTT7_2;
	wire w_dff_B_w31ARI7p5_2;
	wire w_dff_B_q0iaNeqA5_2;
	wire w_dff_B_Ktf7kmeC2_2;
	wire w_dff_B_DQnPTe6U1_2;
	wire w_dff_B_s3baH0L16_2;
	wire w_dff_B_smTXGo765_2;
	wire w_dff_B_wqyk9ScC3_2;
	wire w_dff_B_MOC4qZHb7_2;
	wire w_dff_B_ypz8S9Q79_2;
	wire w_dff_B_NMepsmpw3_2;
	wire w_dff_B_mbJAJiPN0_2;
	wire w_dff_B_yLgDWa1g2_2;
	wire w_dff_B_DO6sKrzx2_2;
	wire w_dff_B_SnAK9J960_2;
	wire w_dff_B_EeLLnJ7g4_2;
	wire w_dff_B_1Klk0tMV1_2;
	wire w_dff_B_OyczPD237_2;
	wire w_dff_B_IZsyeWf28_1;
	wire w_dff_B_L1gaHzF19_2;
	wire w_dff_B_cihPYqz81_2;
	wire w_dff_B_GbGbOR9e9_2;
	wire w_dff_B_zOOFACYH8_2;
	wire w_dff_B_NrA7s80c8_2;
	wire w_dff_B_HsfuJafL4_2;
	wire w_dff_B_z8Spxi6f9_2;
	wire w_dff_B_TMGb5HZq1_2;
	wire w_dff_B_icSf5HTl1_2;
	wire w_dff_B_EAbTJmvu8_2;
	wire w_dff_B_MqnxQ0SH0_2;
	wire w_dff_B_TTRDu9L52_2;
	wire w_dff_B_UTsSfrOG5_2;
	wire w_dff_B_YY5hh0fQ9_2;
	wire w_dff_B_DhV318ib4_2;
	wire w_dff_B_Lf99Nr2G0_2;
	wire w_dff_B_GMR7TjrY2_2;
	wire w_dff_B_JLZtvhgW5_2;
	wire w_dff_B_ih9TGE8T8_2;
	wire w_dff_B_2WOqcq8D2_2;
	wire w_dff_B_NxtaKpLL8_2;
	wire w_dff_B_2FGWKC1H9_2;
	wire w_dff_B_uomZ3BfG8_2;
	wire w_dff_B_vuesWQg10_2;
	wire w_dff_B_0ln7i3yv3_2;
	wire w_dff_B_teh9vl1E7_1;
	wire w_dff_B_52OESfC01_2;
	wire w_dff_B_nySWuDaB3_2;
	wire w_dff_B_0j5IJlxb1_2;
	wire w_dff_B_xUnWSZUa1_2;
	wire w_dff_B_q6Jh4Fqk1_2;
	wire w_dff_B_VqFUs14A8_2;
	wire w_dff_B_PEclydIw9_2;
	wire w_dff_B_dwJuQe8d3_2;
	wire w_dff_B_bEUvZqBd9_2;
	wire w_dff_B_kn7fbtFZ0_2;
	wire w_dff_B_LARXZbmT2_2;
	wire w_dff_B_6HOxNdgJ9_2;
	wire w_dff_B_aX6E68Rs5_2;
	wire w_dff_B_IfY7yqZW1_2;
	wire w_dff_B_qxKB7DB39_2;
	wire w_dff_B_KBa7162e0_2;
	wire w_dff_B_KHTrgNUI6_2;
	wire w_dff_B_iNU01zlk3_2;
	wire w_dff_B_Y66iCzaW2_2;
	wire w_dff_B_FIAq9V0Q4_2;
	wire w_dff_B_F7lIEWSj0_2;
	wire w_dff_B_HKVoNoEe3_2;
	wire w_dff_B_g9P1r5ym0_1;
	wire w_dff_B_xiWu0dwT2_2;
	wire w_dff_B_YHrjbzBw9_2;
	wire w_dff_B_LEWog6le3_2;
	wire w_dff_B_gx8vGpJf7_2;
	wire w_dff_B_iXjk25ko9_2;
	wire w_dff_B_QmnEWcnm7_2;
	wire w_dff_B_Tk30aquB3_2;
	wire w_dff_B_XUzeh79p2_2;
	wire w_dff_B_9RsS1pdi9_2;
	wire w_dff_B_PvucHwYW2_2;
	wire w_dff_B_aHsH2MyB5_2;
	wire w_dff_B_dlJ8ddlK4_2;
	wire w_dff_B_xtYAbrtG5_2;
	wire w_dff_B_ic7GWx239_2;
	wire w_dff_B_ezXa3Q176_2;
	wire w_dff_B_M7KNXDcu3_2;
	wire w_dff_B_E60SA92c5_2;
	wire w_dff_B_A61RqbDr9_2;
	wire w_dff_B_RcsfpYi26_2;
	wire w_dff_B_nYni0s4q4_1;
	wire w_dff_B_16wA4Tok1_2;
	wire w_dff_B_HcoFhwj94_2;
	wire w_dff_B_ssb5h6nL8_2;
	wire w_dff_B_WhAQoRf68_2;
	wire w_dff_B_1W6cgkrg1_2;
	wire w_dff_B_qcw6OwS11_2;
	wire w_dff_B_eBYhpD1m0_2;
	wire w_dff_B_5Y0gQePj7_2;
	wire w_dff_B_gqcx2evk1_2;
	wire w_dff_B_rmOU3GDN6_2;
	wire w_dff_B_z7giTpya6_2;
	wire w_dff_B_Z3acxj7O5_2;
	wire w_dff_B_SG9yeJir4_2;
	wire w_dff_B_f9xz1iH55_2;
	wire w_dff_B_JmAnH8nQ3_2;
	wire w_dff_B_Lcdxw4Xr7_2;
	wire w_dff_B_6TftSVYF7_1;
	wire w_dff_B_fOZFgnN18_2;
	wire w_dff_B_J6dWZeOp2_2;
	wire w_dff_B_NEtTj2Mq9_2;
	wire w_dff_B_S3EBGOoQ6_2;
	wire w_dff_B_y1VeWTxt8_2;
	wire w_dff_B_jOoHe2UU8_2;
	wire w_dff_B_gsI5fYDQ3_2;
	wire w_dff_B_NBf5rh7b4_2;
	wire w_dff_B_OydbojVv2_2;
	wire w_dff_B_XepdfhXy6_2;
	wire w_dff_B_r2F1US2v5_2;
	wire w_dff_B_Fx7TQE1T8_2;
	wire w_dff_B_tWtJj8lm3_2;
	wire w_dff_B_R12el6iH1_1;
	wire w_dff_B_tdkRVyET1_2;
	wire w_dff_B_Dw7Hi8SV3_2;
	wire w_dff_B_frbER5xA9_2;
	wire w_dff_B_rmnmQTaV7_2;
	wire w_dff_B_qIGRpHMu2_2;
	wire w_dff_B_3QBsWR8H1_2;
	wire w_dff_B_zqHIAowd4_2;
	wire w_dff_B_y05Obsgc0_2;
	wire w_dff_B_PumEGzma6_2;
	wire w_dff_B_yd2VpjQb7_2;
	wire w_dff_B_GTmP2KeA8_2;
	wire w_dff_B_Y7u0ICTY3_1;
	wire w_dff_B_vMOoao6P2_1;
	wire w_dff_B_6wM3bMd49_1;
	wire w_dff_B_GKLQP4Ta8_1;
	wire w_dff_B_pEl37SFF6_1;
	wire w_dff_B_w4rI4dlB8_1;
	wire w_dff_B_uvHwSihO4_0;
	wire w_dff_B_yeWItqQb4_0;
	wire w_dff_A_sMSki8O07_0;
	wire w_dff_A_mV1ETtr76_0;
	wire w_dff_A_DwgwG6gr1_0;
	wire w_dff_B_wtlWOni45_1;
	wire w_dff_A_8UhmKZc75_0;
	wire w_dff_A_TaYnXwFq7_1;
	wire w_dff_A_NfLo46A38_1;
	wire w_dff_A_lD78zEp75_1;
	wire w_dff_A_iRN75Ff71_1;
	wire w_dff_A_U1GsVckW9_1;
	wire w_dff_A_kf5tlb256_1;
	wire w_dff_A_9RwiuLbM9_1;
	wire w_dff_A_7lPIcV558_1;
	wire w_dff_B_swAYl7xU4_1;
	wire w_dff_A_WItlfLpC4_1;
	wire w_dff_B_LzPbpWEu3_1;
	wire w_dff_B_H6mtBv1K6_2;
	wire w_dff_B_9XvtSTpv6_2;
	wire w_dff_B_yb1kLai44_2;
	wire w_dff_B_9JzcRiYJ3_2;
	wire w_dff_B_kdxV89qc4_2;
	wire w_dff_B_1nr48IKx1_2;
	wire w_dff_B_anXGj3Lk6_2;
	wire w_dff_B_gP6AfZ4R5_2;
	wire w_dff_B_l7rqyiSV9_2;
	wire w_dff_B_ShfQ0cvR2_2;
	wire w_dff_B_svNpG9i57_2;
	wire w_dff_B_xp2N5JwY0_2;
	wire w_dff_B_jlivo5LI9_2;
	wire w_dff_B_ej2HIOCH3_2;
	wire w_dff_B_6jU6beEu7_2;
	wire w_dff_B_aEVKyXID7_2;
	wire w_dff_B_ZU662TJJ7_2;
	wire w_dff_B_4qnuRD3s8_2;
	wire w_dff_B_9Gx5wGeG1_2;
	wire w_dff_B_Yo0Vf7SH7_2;
	wire w_dff_B_LbMODvhb2_2;
	wire w_dff_B_wrDSOEST9_2;
	wire w_dff_B_EIvnxcR78_2;
	wire w_dff_B_5v8GyuaA4_2;
	wire w_dff_B_Yhoexs5x1_2;
	wire w_dff_B_OrtWqyKA3_2;
	wire w_dff_B_tgn7m4K28_2;
	wire w_dff_B_yJcC1C7Q1_2;
	wire w_dff_B_UPcYNmSS2_2;
	wire w_dff_B_RIwApUQW6_2;
	wire w_dff_B_bQfhKYo91_2;
	wire w_dff_B_fMkyXAsr2_2;
	wire w_dff_B_zsGQLSGN9_2;
	wire w_dff_B_9FlxtoOI5_2;
	wire w_dff_B_IQdKcivU4_2;
	wire w_dff_B_CUKrA4Cw9_2;
	wire w_dff_B_Y9PhFo438_2;
	wire w_dff_B_LzbBETMS3_2;
	wire w_dff_B_957WxHNJ7_2;
	wire w_dff_B_rqZ2L9jc4_2;
	wire w_dff_B_tdgePMaP4_2;
	wire w_dff_B_gUyDHGLI0_2;
	wire w_dff_B_9MgmbgsI1_2;
	wire w_dff_B_syFGDCgS1_2;
	wire w_dff_B_utdgoEAV1_2;
	wire w_dff_B_YSxTucuZ5_2;
	wire w_dff_B_j7cEDYbT1_2;
	wire w_dff_B_wcq1zbGT0_2;
	wire w_dff_B_umlEhmbA0_2;
	wire w_dff_B_8T0UyFxb2_2;
	wire w_dff_B_xe0e7oJ50_2;
	wire w_dff_B_bUQI7BuH1_2;
	wire w_dff_B_cbqqkSOt3_1;
	wire w_dff_B_4WuJtOWd5_2;
	wire w_dff_B_YOyTYtVv5_2;
	wire w_dff_B_d9tLDOwU8_2;
	wire w_dff_B_BqLPgxoY5_2;
	wire w_dff_B_a0WegON35_2;
	wire w_dff_B_0Z9Q4Un26_2;
	wire w_dff_B_N1F4fEdb1_2;
	wire w_dff_B_eTMkIJLa1_2;
	wire w_dff_B_djqRUxpN1_2;
	wire w_dff_B_o3iJ7W9p2_2;
	wire w_dff_B_QkBUDKmJ9_2;
	wire w_dff_B_HMeZxEat8_2;
	wire w_dff_B_VgB0xkrC5_2;
	wire w_dff_B_edFqKEm53_2;
	wire w_dff_B_fH4Oxttf8_2;
	wire w_dff_B_NOTK3CBt7_2;
	wire w_dff_B_dPVSB4Nc7_2;
	wire w_dff_B_aFdUhKba3_2;
	wire w_dff_B_qMp8mdia4_2;
	wire w_dff_B_RoXPRaTS4_2;
	wire w_dff_B_bJhY5KSt2_2;
	wire w_dff_B_EZ6E0mIH9_2;
	wire w_dff_B_LiOHpp0s8_2;
	wire w_dff_B_UvNqbsXi3_2;
	wire w_dff_B_ZYkrU6122_2;
	wire w_dff_B_kyw1KR4g9_2;
	wire w_dff_B_P62hqi5Z4_2;
	wire w_dff_B_txPKKbPr8_2;
	wire w_dff_B_41AylPxe4_2;
	wire w_dff_B_mOKvSalK5_2;
	wire w_dff_B_z47xiuzn1_2;
	wire w_dff_B_K2Habuhe4_2;
	wire w_dff_B_KRwvONfS6_2;
	wire w_dff_B_3NSyxBTa3_2;
	wire w_dff_B_ExW8D8dv7_2;
	wire w_dff_B_GnmsHfMT3_2;
	wire w_dff_B_GJ6aRfhb6_2;
	wire w_dff_B_yQM7XMqw2_2;
	wire w_dff_B_vBvVXIyN1_2;
	wire w_dff_B_EN9LNgMC8_2;
	wire w_dff_B_sg1tNUUs7_2;
	wire w_dff_B_FcxZ8jjA7_2;
	wire w_dff_B_Z0iUD3KS2_2;
	wire w_dff_B_GnLQSwgO7_2;
	wire w_dff_B_mYHW4hAb0_2;
	wire w_dff_B_5F8Eq4700_2;
	wire w_dff_B_nj4zgaFg1_2;
	wire w_dff_B_jVVl5q6J8_2;
	wire w_dff_B_YNu2zp3w3_1;
	wire w_dff_B_TUQ9DmFl3_2;
	wire w_dff_B_2OdILCNc6_2;
	wire w_dff_B_OjvU5On85_2;
	wire w_dff_B_mLQhD9fW2_2;
	wire w_dff_B_oWwDZk5Y7_2;
	wire w_dff_B_GoOhqLBZ2_2;
	wire w_dff_B_eizSrCK38_2;
	wire w_dff_B_bcoynlxS0_2;
	wire w_dff_B_3A4MX6ls7_2;
	wire w_dff_B_tWhHESrw8_2;
	wire w_dff_B_VIfc0kX26_2;
	wire w_dff_B_zEMQBD2f6_2;
	wire w_dff_B_BKvZJwyW9_2;
	wire w_dff_B_yNQHINSw0_2;
	wire w_dff_B_qfR2ewqZ8_2;
	wire w_dff_B_K5ZmDyLb1_2;
	wire w_dff_B_0YAJk6Uj1_2;
	wire w_dff_B_z8BhNc4j2_2;
	wire w_dff_B_Y3ZIg1M75_2;
	wire w_dff_B_YSqnfV811_2;
	wire w_dff_B_ai8j6rzt5_2;
	wire w_dff_B_a98vFQd63_2;
	wire w_dff_B_CsJ1R2Tr4_2;
	wire w_dff_B_aDMptzkZ5_2;
	wire w_dff_B_ZLN7o7mO9_2;
	wire w_dff_B_W97JhkRO2_2;
	wire w_dff_B_GUzZIFy88_2;
	wire w_dff_B_5vcJ02eG7_2;
	wire w_dff_B_LgymVEUt2_2;
	wire w_dff_B_SrU3J8Tn8_2;
	wire w_dff_B_90hJe6is0_2;
	wire w_dff_B_An0iTvcV8_2;
	wire w_dff_B_CV5w5Dn94_2;
	wire w_dff_B_TMIYBPzl7_2;
	wire w_dff_B_GfeaITEK3_2;
	wire w_dff_B_o6gHOwCh1_2;
	wire w_dff_B_N1nDXXcd8_2;
	wire w_dff_B_X9SB6rxh9_2;
	wire w_dff_B_AvYioCkM2_2;
	wire w_dff_B_9ONkPx6P2_2;
	wire w_dff_B_sS0vzrBr8_2;
	wire w_dff_B_hSEr7CFm3_2;
	wire w_dff_B_gg96ixUT7_2;
	wire w_dff_B_RlKTCuxy7_2;
	wire w_dff_B_jPDNsV4f5_1;
	wire w_dff_B_FWhxwsyp1_2;
	wire w_dff_B_hN6NoHL09_2;
	wire w_dff_B_LmcKsD8k2_2;
	wire w_dff_B_HEZbZo4H0_2;
	wire w_dff_B_a5JieUma1_2;
	wire w_dff_B_SZllBtwh5_2;
	wire w_dff_B_CWE7WaOw3_2;
	wire w_dff_B_T5ucWDJP3_2;
	wire w_dff_B_vUhUwuC36_2;
	wire w_dff_B_qWV9Z5bT0_2;
	wire w_dff_B_S8Pv2Su02_2;
	wire w_dff_B_vTyWXmq13_2;
	wire w_dff_B_bPFVtFv45_2;
	wire w_dff_B_N6U4zmN03_2;
	wire w_dff_B_SSUob3hE8_2;
	wire w_dff_B_NT6MnoK61_2;
	wire w_dff_B_5oPMN6Tr6_2;
	wire w_dff_B_fIFqLAVR8_2;
	wire w_dff_B_A35TbZZY1_2;
	wire w_dff_B_TuHtGioY2_2;
	wire w_dff_B_EenB9Ik38_2;
	wire w_dff_B_zcY1HmAm6_2;
	wire w_dff_B_9DLkRjS03_2;
	wire w_dff_B_vGgx5UOl8_2;
	wire w_dff_B_0ss9W9jf0_2;
	wire w_dff_B_sQzvEDJH0_2;
	wire w_dff_B_Hj9Y9dzq5_2;
	wire w_dff_B_RE2q9mKr2_2;
	wire w_dff_B_cgkKqhsh2_2;
	wire w_dff_B_IllvyTv35_2;
	wire w_dff_B_OzYlfES70_2;
	wire w_dff_B_CupDJq5Y7_2;
	wire w_dff_B_V3vfjcVw0_2;
	wire w_dff_B_Cfb4vqSe7_2;
	wire w_dff_B_4C0WKNQH4_2;
	wire w_dff_B_i96nFEU98_2;
	wire w_dff_B_ypZ51DHP7_2;
	wire w_dff_B_zk0hrgOT6_2;
	wire w_dff_B_fmCt4rpQ0_2;
	wire w_dff_B_Us3zuZTo6_2;
	wire w_dff_B_8o2FsipG4_1;
	wire w_dff_B_yvHiPnQw7_2;
	wire w_dff_B_jUVPFEwC2_2;
	wire w_dff_B_GJuLF0m44_2;
	wire w_dff_B_b12wuBNb6_2;
	wire w_dff_B_qay5OBGx1_2;
	wire w_dff_B_lP0gwImO0_2;
	wire w_dff_B_k7XucLjP3_2;
	wire w_dff_B_NqDDxPS28_2;
	wire w_dff_B_0JQlx2xx9_2;
	wire w_dff_B_dDyXOI5Y6_2;
	wire w_dff_B_3T4EUipr5_2;
	wire w_dff_B_EmAbx1th6_2;
	wire w_dff_B_zDFDPh4S8_2;
	wire w_dff_B_MmorXoxh8_2;
	wire w_dff_B_7aMezkkc7_2;
	wire w_dff_B_PZUNlUiX7_2;
	wire w_dff_B_C1bhB9y15_2;
	wire w_dff_B_wL0SRZO77_2;
	wire w_dff_B_PQmflSPZ8_2;
	wire w_dff_B_2bVdqd6s8_2;
	wire w_dff_B_DQ6r8t1B7_2;
	wire w_dff_B_cIbBd5qZ7_2;
	wire w_dff_B_RacqNaBe5_2;
	wire w_dff_B_nD6vQqlA2_2;
	wire w_dff_B_uNVs8MvF4_2;
	wire w_dff_B_JQlG46sZ5_2;
	wire w_dff_B_VGko9RUY8_2;
	wire w_dff_B_HTldysDF6_2;
	wire w_dff_B_JzVxaj0z2_2;
	wire w_dff_B_NyAFTD8h7_2;
	wire w_dff_B_H3rhAmjQ4_2;
	wire w_dff_B_SUOXQVS70_2;
	wire w_dff_B_9UqHuJWk3_2;
	wire w_dff_B_5af9HRqt5_2;
	wire w_dff_B_68ngA5Vo5_2;
	wire w_dff_B_OMES7jqo9_2;
	wire w_dff_B_u5IVoq2a4_1;
	wire w_dff_B_YcFCBFPO3_2;
	wire w_dff_B_w4zDWyvm6_2;
	wire w_dff_B_2JWSzrzO0_2;
	wire w_dff_B_oTIs4USt9_2;
	wire w_dff_B_3zipsOJY5_2;
	wire w_dff_B_YIFSJtrs0_2;
	wire w_dff_B_N4acTxeA6_2;
	wire w_dff_B_eXEd1Tmq8_2;
	wire w_dff_B_21cSfqmk9_2;
	wire w_dff_B_OydAEvk49_2;
	wire w_dff_B_zLqu2rxX3_2;
	wire w_dff_B_zXzp0jIM8_2;
	wire w_dff_B_anhUD9a27_2;
	wire w_dff_B_eE1Wg2bl5_2;
	wire w_dff_B_MDKR1x8E2_2;
	wire w_dff_B_2O9MIAMb3_2;
	wire w_dff_B_iNFgzxZ08_2;
	wire w_dff_B_U8aDgk9d7_2;
	wire w_dff_B_ufLv9hl44_2;
	wire w_dff_B_8vwtoFUA6_2;
	wire w_dff_B_n7xiUSD47_2;
	wire w_dff_B_kciiJgb55_2;
	wire w_dff_B_zEkxCo4z3_2;
	wire w_dff_B_pgNjoc4F8_2;
	wire w_dff_B_u9kmetFt3_2;
	wire w_dff_B_ltVj1MsD6_2;
	wire w_dff_B_W2YPltbM3_2;
	wire w_dff_B_2oCdhB3n3_2;
	wire w_dff_B_ajPvAAUC4_2;
	wire w_dff_B_jYZV3R8I4_2;
	wire w_dff_B_jjedWkFG1_2;
	wire w_dff_B_njPQvG9e8_2;
	wire w_dff_B_DeIbx7lP9_1;
	wire w_dff_B_8e4NqzHw4_2;
	wire w_dff_B_9Vh8Bn5K4_2;
	wire w_dff_B_yRa6JZ6l7_2;
	wire w_dff_B_zdwx9JsP5_2;
	wire w_dff_B_3RknptOY1_2;
	wire w_dff_B_AOVLuSwa7_2;
	wire w_dff_B_wrNpn0Rv4_2;
	wire w_dff_B_SuxR5NWe6_2;
	wire w_dff_B_9Vxltf1N5_2;
	wire w_dff_B_oSCyB8iY8_2;
	wire w_dff_B_yrycadkq0_2;
	wire w_dff_B_vIIsJsSq8_2;
	wire w_dff_B_TgSk8gGZ1_2;
	wire w_dff_B_TFTtsks27_2;
	wire w_dff_B_RvZnRIGG5_2;
	wire w_dff_B_QD4U42DU1_2;
	wire w_dff_B_0sF7O7788_2;
	wire w_dff_B_VaE4exiy4_2;
	wire w_dff_B_xy9r5xCJ6_2;
	wire w_dff_B_rrP0XZrv6_2;
	wire w_dff_B_EjHAvBwx7_2;
	wire w_dff_B_dbN2Nquh8_2;
	wire w_dff_B_e34QdL9G8_2;
	wire w_dff_B_8cxraynF3_2;
	wire w_dff_B_QbmdQVPc6_2;
	wire w_dff_B_ouMsuwRl7_2;
	wire w_dff_B_kHJAgOSm2_2;
	wire w_dff_B_g4zIW2PC4_1;
	wire w_dff_B_AYwQZKXF4_2;
	wire w_dff_B_xaBHkDI30_2;
	wire w_dff_B_jeOGttWN8_2;
	wire w_dff_B_dHIOjesb1_2;
	wire w_dff_B_ygGQLR5W8_2;
	wire w_dff_B_WynmUHo74_2;
	wire w_dff_B_7KpYrw5Z4_2;
	wire w_dff_B_UVypv7lh7_2;
	wire w_dff_B_Ol5CSGFC4_2;
	wire w_dff_B_LUr1MXYX4_2;
	wire w_dff_B_URSG0eUG4_2;
	wire w_dff_B_7Jq3Nyio3_2;
	wire w_dff_B_k5Q1N5zD2_2;
	wire w_dff_B_OYPcVGBD1_2;
	wire w_dff_B_qXnGpUXg3_2;
	wire w_dff_B_IPPbY5Lz0_2;
	wire w_dff_B_1rwHte9Y5_2;
	wire w_dff_B_Np6mHN2u7_2;
	wire w_dff_B_jslJltsU6_2;
	wire w_dff_B_prf6axQ95_2;
	wire w_dff_B_AoafReTF8_2;
	wire w_dff_B_ikuXHfzF8_2;
	wire w_dff_B_5rfyVuhh2_2;
	wire w_dff_B_bpkdk6rt2_2;
	wire w_dff_B_JJRZtfhZ9_2;
	wire w_dff_B_uZ7dF0Vi0_1;
	wire w_dff_B_NOQlrnEz4_2;
	wire w_dff_B_ivEGhaFx0_2;
	wire w_dff_B_GRbcs1Zq0_2;
	wire w_dff_B_COEcUgMw3_2;
	wire w_dff_B_gJR63a2E9_2;
	wire w_dff_B_GG8SLyLe1_2;
	wire w_dff_B_q7RnC2cO8_2;
	wire w_dff_B_qG4cZdZk7_2;
	wire w_dff_B_9R7Dz9iL9_2;
	wire w_dff_B_vYsibJJa3_2;
	wire w_dff_B_eu0eYM0b0_2;
	wire w_dff_B_8myywXnU8_2;
	wire w_dff_B_mOsJWtyd9_2;
	wire w_dff_B_bH83fHp69_2;
	wire w_dff_B_Fzu3Vkti7_2;
	wire w_dff_B_zByCkGqu9_2;
	wire w_dff_B_Tcx4Y4gi5_2;
	wire w_dff_B_JkexPaGh0_2;
	wire w_dff_B_o4Lc9StX7_2;
	wire w_dff_B_n4cbJXyH0_2;
	wire w_dff_B_eXoYxCfj8_2;
	wire w_dff_B_cMtgVFzy1_2;
	wire w_dff_B_kK2ESgpI4_1;
	wire w_dff_B_mHn6A1TG5_2;
	wire w_dff_B_1vwQrPGr6_2;
	wire w_dff_B_qlumm9ey3_2;
	wire w_dff_B_buLk5kNv1_2;
	wire w_dff_B_brqUSC524_2;
	wire w_dff_B_hmKDX2123_2;
	wire w_dff_B_7a6b6YKa7_2;
	wire w_dff_B_KfiuQHT62_2;
	wire w_dff_B_UX5K9AA02_2;
	wire w_dff_B_5xw0O59C9_2;
	wire w_dff_B_XaBd5fvY9_2;
	wire w_dff_B_4Ajmh4Hz1_2;
	wire w_dff_B_GeeD8kzF0_2;
	wire w_dff_B_nEMqyReq9_2;
	wire w_dff_B_jiPdFc5v4_2;
	wire w_dff_B_7nqQFFA68_2;
	wire w_dff_B_KYByy9QX1_2;
	wire w_dff_B_9eFiQyfl7_2;
	wire w_dff_B_hZ2lehh50_2;
	wire w_dff_B_yk5YtVJ65_1;
	wire w_dff_B_iFI0Jw5b8_2;
	wire w_dff_B_Kv4pRacZ1_2;
	wire w_dff_B_bLaoZtQK9_2;
	wire w_dff_B_Tk3tCumm3_2;
	wire w_dff_B_RIbb9lo81_2;
	wire w_dff_B_fNkKkKfD6_2;
	wire w_dff_B_zRxHkNoV3_2;
	wire w_dff_B_FNNAJWGs8_2;
	wire w_dff_B_uVu1qw1Q7_2;
	wire w_dff_B_4lKUbKg04_2;
	wire w_dff_B_Tmmw64Qi2_2;
	wire w_dff_B_paeWwoNP1_2;
	wire w_dff_B_vV0WF0t53_2;
	wire w_dff_B_blbVkEUT9_2;
	wire w_dff_B_bflIGW7s7_2;
	wire w_dff_B_i5sM6kEZ8_2;
	wire w_dff_B_SB7dlvBc6_1;
	wire w_dff_B_Sklpz0k90_2;
	wire w_dff_B_W4v6kaYt6_2;
	wire w_dff_B_E09KK3E12_2;
	wire w_dff_B_lPn8Wxfn7_2;
	wire w_dff_B_jxOpEzbY9_2;
	wire w_dff_B_aE7bPIxk7_2;
	wire w_dff_B_kEUTOeIR7_2;
	wire w_dff_B_v4S3pv8l4_2;
	wire w_dff_B_EhWVhiBI6_2;
	wire w_dff_B_LIaiFfNQ6_2;
	wire w_dff_B_uKetQiRC1_2;
	wire w_dff_B_yAr04H9W1_2;
	wire w_dff_B_QPpQGM361_2;
	wire w_dff_B_UNbWXrTi5_1;
	wire w_dff_B_C5q94eMr1_2;
	wire w_dff_B_irBegRFQ8_2;
	wire w_dff_B_qwRekFJZ8_2;
	wire w_dff_B_eb8W9Ta22_2;
	wire w_dff_B_l2EDcrU55_2;
	wire w_dff_B_85hhOQCy4_2;
	wire w_dff_B_qsBeduna3_2;
	wire w_dff_B_XGOvkdA66_2;
	wire w_dff_B_4LFn6EgN7_2;
	wire w_dff_B_6JFRe99A8_2;
	wire w_dff_B_nzwKRckY6_2;
	wire w_dff_B_F6KKqp0I8_1;
	wire w_dff_B_208H61nz4_1;
	wire w_dff_B_nfh0Anse2_1;
	wire w_dff_B_aGehSRJq9_1;
	wire w_dff_B_pK6cNqnY1_1;
	wire w_dff_B_ycQziHRj5_1;
	wire w_dff_B_ghKvLSbr0_0;
	wire w_dff_B_PYhFfXDa8_0;
	wire w_dff_A_Iuo8bC7C8_0;
	wire w_dff_A_UmkstwiT2_0;
	wire w_dff_A_LRlOYx2p2_0;
	wire w_dff_B_j6eUikvB2_1;
	wire w_dff_A_Ai6ny8Yz9_0;
	wire w_dff_A_sWnJlBNP2_1;
	wire w_dff_A_MUWNUiji3_1;
	wire w_dff_A_DKGW4iE87_1;
	wire w_dff_A_ZtDRweVm1_1;
	wire w_dff_A_3Pzw6UTd0_1;
	wire w_dff_A_1d6TTFCT0_1;
	wire w_dff_A_Ophfcl6M1_1;
	wire w_dff_A_bBP3iweD3_1;
	wire w_dff_B_NiRQ0XUX0_1;
	wire w_dff_A_yvPCCEoS2_1;
	wire w_dff_B_CTe4bPiS3_1;
	wire w_dff_B_4nIVDGd25_2;
	wire w_dff_B_QUfPRJAv6_2;
	wire w_dff_B_quiluQjn1_2;
	wire w_dff_B_Lwpwq0Rs1_2;
	wire w_dff_B_go08VVGf3_2;
	wire w_dff_B_r02VsDN50_2;
	wire w_dff_B_AD3YtUdT3_2;
	wire w_dff_B_YidBgOfN1_2;
	wire w_dff_B_Eh6HP9FU7_2;
	wire w_dff_B_aCqiNgN90_2;
	wire w_dff_B_O7uZei4a2_2;
	wire w_dff_B_KlPistLC0_2;
	wire w_dff_B_5Uci0xnl4_2;
	wire w_dff_B_tsTNUwdT8_2;
	wire w_dff_B_IhEt0xlD8_2;
	wire w_dff_B_R5eYr6q44_2;
	wire w_dff_B_HF8XaDwQ5_2;
	wire w_dff_B_eCZCoMfL5_2;
	wire w_dff_B_65c9tFPw6_2;
	wire w_dff_B_c7nY5kDD2_2;
	wire w_dff_B_aUv76SM82_2;
	wire w_dff_B_NjvE3s542_2;
	wire w_dff_B_BeEC1Zg71_2;
	wire w_dff_B_8o94F5ir9_2;
	wire w_dff_B_6jffrsIL3_2;
	wire w_dff_B_obcOtCP87_2;
	wire w_dff_B_hwvu0FLI9_2;
	wire w_dff_B_pbZRBvRS6_2;
	wire w_dff_B_SPRwxoXi1_2;
	wire w_dff_B_W5tD9vhU1_2;
	wire w_dff_B_gKsJZiiL0_2;
	wire w_dff_B_kiKmBUMo3_2;
	wire w_dff_B_tROCr7Qy1_2;
	wire w_dff_B_9DKHQsVB6_2;
	wire w_dff_B_lvIOlS5B8_2;
	wire w_dff_B_aULnmtzK4_2;
	wire w_dff_B_gICv0iZF9_2;
	wire w_dff_B_qNV9so0P2_2;
	wire w_dff_B_ymtchohA0_2;
	wire w_dff_B_hzjYATWG7_2;
	wire w_dff_B_mX3K5PLX2_2;
	wire w_dff_B_CxOv5dCV8_2;
	wire w_dff_B_N9peuzqX8_2;
	wire w_dff_B_ia8C6Jxo2_2;
	wire w_dff_B_4h1mvUyI5_2;
	wire w_dff_B_dFVoXNyH6_2;
	wire w_dff_B_R2Uyxj707_2;
	wire w_dff_B_t6OTknWa2_2;
	wire w_dff_B_KJSXHFsq9_2;
	wire w_dff_B_ZaTVUDFY8_2;
	wire w_dff_B_NrKguckG2_2;
	wire w_dff_B_slftNcig9_2;
	wire w_dff_B_Yzc9RcZh4_2;
	wire w_dff_B_2XG2nvNA2_2;
	wire w_dff_B_b90Z7vXn8_1;
	wire w_dff_B_KXCtdLDY9_2;
	wire w_dff_B_ZPMbSx675_2;
	wire w_dff_B_oabqylBl9_2;
	wire w_dff_B_A0AcWmW61_2;
	wire w_dff_B_3pAKkzOx4_2;
	wire w_dff_B_qUoeQIKv6_2;
	wire w_dff_B_s4PK1PJk0_2;
	wire w_dff_B_5qVeG1Dk9_2;
	wire w_dff_B_ZdHKM6qD3_2;
	wire w_dff_B_i9an8hkh6_2;
	wire w_dff_B_5sjCzV3N6_2;
	wire w_dff_B_gPof9vDJ0_2;
	wire w_dff_B_Aq0lgHlt0_2;
	wire w_dff_B_Tres6fIH3_2;
	wire w_dff_B_b7EvgEKd2_2;
	wire w_dff_B_9vI8bOzX1_2;
	wire w_dff_B_2RDqrGKY7_2;
	wire w_dff_B_5TwqCLW80_2;
	wire w_dff_B_woQAuOM94_2;
	wire w_dff_B_f2G8Qthw2_2;
	wire w_dff_B_PG6hOt2x3_2;
	wire w_dff_B_m0ipGKvO8_2;
	wire w_dff_B_lUtFYRnr3_2;
	wire w_dff_B_KebbMlSm5_2;
	wire w_dff_B_oNxnqqyu5_2;
	wire w_dff_B_1l8dkLAa2_2;
	wire w_dff_B_nCz172J18_2;
	wire w_dff_B_AxL68lvD9_2;
	wire w_dff_B_f5mxh1ET3_2;
	wire w_dff_B_o20zr0du2_2;
	wire w_dff_B_ZeIq7Lxt3_2;
	wire w_dff_B_3OKcia3V4_2;
	wire w_dff_B_x1Y6veYi8_2;
	wire w_dff_B_mrBya4Ue2_2;
	wire w_dff_B_1rR9e1Ob7_2;
	wire w_dff_B_VgSSCo7L6_2;
	wire w_dff_B_4Inb6VYI6_2;
	wire w_dff_B_iFlcSjGb2_2;
	wire w_dff_B_Uc3LKQd95_2;
	wire w_dff_B_7uSCX6Ej2_2;
	wire w_dff_B_VTXlkmTV2_2;
	wire w_dff_B_ta4tm3Ee2_2;
	wire w_dff_B_ETpWHW4o5_2;
	wire w_dff_B_2PiFW1EC3_2;
	wire w_dff_B_hXelHWkr4_2;
	wire w_dff_B_1YHFoZHD0_2;
	wire w_dff_B_xCbISSsD1_2;
	wire w_dff_B_MIp6UnZx6_2;
	wire w_dff_B_09FlSBNU8_2;
	wire w_dff_B_Hto6pA017_2;
	wire w_dff_B_GBFhlqJt1_1;
	wire w_dff_B_4UDLIoq55_2;
	wire w_dff_B_6W6ZzYxM6_2;
	wire w_dff_B_XH1xguaG7_2;
	wire w_dff_B_wEzATMU09_2;
	wire w_dff_B_nndZOcyO3_2;
	wire w_dff_B_DFfnGP5J9_2;
	wire w_dff_B_BLdlEHzf0_2;
	wire w_dff_B_mh1EG16L9_2;
	wire w_dff_B_k5sQI2H94_2;
	wire w_dff_B_gIS3kEDz2_2;
	wire w_dff_B_WuTXHVMW8_2;
	wire w_dff_B_tVhIJKlQ7_2;
	wire w_dff_B_cWNrJTbM5_2;
	wire w_dff_B_kbAsr9uR3_2;
	wire w_dff_B_NipPy7uN2_2;
	wire w_dff_B_eiXdaOvx5_2;
	wire w_dff_B_vLi2tK112_2;
	wire w_dff_B_ksl1FEt55_2;
	wire w_dff_B_9juIz4GK3_2;
	wire w_dff_B_87lSFLpn4_2;
	wire w_dff_B_uX0s9TIR7_2;
	wire w_dff_B_K6W7jNUc1_2;
	wire w_dff_B_xBMYqHLV8_2;
	wire w_dff_B_D1VcgLeh7_2;
	wire w_dff_B_Kc3U1Dgf5_2;
	wire w_dff_B_fS7xFAsa4_2;
	wire w_dff_B_hJgONq219_2;
	wire w_dff_B_7HZ5Uspp5_2;
	wire w_dff_B_lRMMQxUd3_2;
	wire w_dff_B_NUYPluOB9_2;
	wire w_dff_B_M4hO2AI63_2;
	wire w_dff_B_E38pZlid0_2;
	wire w_dff_B_v3RGeEgj5_2;
	wire w_dff_B_0IskqFG09_2;
	wire w_dff_B_s5JImO5R6_2;
	wire w_dff_B_IFDitTZ19_2;
	wire w_dff_B_zqvwS3iM5_2;
	wire w_dff_B_i1aIOw928_2;
	wire w_dff_B_Gdc5TsG35_2;
	wire w_dff_B_CqHiyiZY7_2;
	wire w_dff_B_LfEiPaCA7_2;
	wire w_dff_B_Gpze2ohh9_2;
	wire w_dff_B_4OrxLSvx8_2;
	wire w_dff_B_lb9kz3zq0_2;
	wire w_dff_B_icbpygs14_2;
	wire w_dff_B_CWjW9Ljq8_2;
	wire w_dff_B_IVGV1hWr7_1;
	wire w_dff_B_273ZWcL18_2;
	wire w_dff_B_gLWEgUOH6_2;
	wire w_dff_B_oco2Xphf9_2;
	wire w_dff_B_xZiyinH49_2;
	wire w_dff_B_QtSkH6op7_2;
	wire w_dff_B_n6Yh4seq7_2;
	wire w_dff_B_7MxdhzbH0_2;
	wire w_dff_B_g5a79xU07_2;
	wire w_dff_B_W0GnBM7v9_2;
	wire w_dff_B_ApJ9mZ5m1_2;
	wire w_dff_B_BeobT1ZP5_2;
	wire w_dff_B_vW33an8Q9_2;
	wire w_dff_B_QOIXrkTW8_2;
	wire w_dff_B_NtK0a0m25_2;
	wire w_dff_B_VCgPFZcq9_2;
	wire w_dff_B_g26D1fnS9_2;
	wire w_dff_B_cUQTFXfz3_2;
	wire w_dff_B_fc7bjt8A9_2;
	wire w_dff_B_QTttfCQz4_2;
	wire w_dff_B_dN2AR35P0_2;
	wire w_dff_B_TOHUYWdZ1_2;
	wire w_dff_B_q6qrVm9B0_2;
	wire w_dff_B_OihMuvS32_2;
	wire w_dff_B_ndJRK4Ir6_2;
	wire w_dff_B_if7qqmyu3_2;
	wire w_dff_B_pksl8QHj3_2;
	wire w_dff_B_i6IMqcDR0_2;
	wire w_dff_B_k2vqLwNI5_2;
	wire w_dff_B_JnDYOcxb6_2;
	wire w_dff_B_u2SVdbn26_2;
	wire w_dff_B_uyYZNR952_2;
	wire w_dff_B_CaS43xin0_2;
	wire w_dff_B_iTqTfpYg1_2;
	wire w_dff_B_JzbMjfsx6_2;
	wire w_dff_B_Qe7aWXeH0_2;
	wire w_dff_B_045T1oLg8_2;
	wire w_dff_B_URcjHMWH7_2;
	wire w_dff_B_hyrv6va34_2;
	wire w_dff_B_dnZ792338_2;
	wire w_dff_B_mFUXl2Vr0_2;
	wire w_dff_B_49g8mCix4_2;
	wire w_dff_B_D0oz23es3_2;
	wire w_dff_B_BceJ9HAg2_1;
	wire w_dff_B_XU1ib5pi4_2;
	wire w_dff_B_4Hf9CiEg8_2;
	wire w_dff_B_PQbTCk5t0_2;
	wire w_dff_B_JwZJKHav3_2;
	wire w_dff_B_IU07JJ6l8_2;
	wire w_dff_B_iQyohNPb5_2;
	wire w_dff_B_2syLQrTk8_2;
	wire w_dff_B_c6BjeoqK3_2;
	wire w_dff_B_5CWHnyk14_2;
	wire w_dff_B_1ev366XH7_2;
	wire w_dff_B_kAPCeusT6_2;
	wire w_dff_B_Ui9tzaJe3_2;
	wire w_dff_B_8hseRavn4_2;
	wire w_dff_B_1hIBzhWY4_2;
	wire w_dff_B_yPUbsZcR6_2;
	wire w_dff_B_0Yx81Hka1_2;
	wire w_dff_B_0iY5WYrK6_2;
	wire w_dff_B_vIluE7Hi3_2;
	wire w_dff_B_jO7epaEW3_2;
	wire w_dff_B_Qwxy4cgT8_2;
	wire w_dff_B_6P7mbnmE0_2;
	wire w_dff_B_T9lmb8lD4_2;
	wire w_dff_B_uBmoyWnJ8_2;
	wire w_dff_B_aXfjF8iJ7_2;
	wire w_dff_B_L5RnNB3u8_2;
	wire w_dff_B_F3I74PE33_2;
	wire w_dff_B_OSC9w5fH6_2;
	wire w_dff_B_7aV4A1kK0_2;
	wire w_dff_B_Vqb8uKpm7_2;
	wire w_dff_B_VZEGaTD22_2;
	wire w_dff_B_e2dWQ5mI9_2;
	wire w_dff_B_eWJ0iAyU8_2;
	wire w_dff_B_yTiDZGKA7_2;
	wire w_dff_B_BB7c8lP05_2;
	wire w_dff_B_9VhKkMOn9_2;
	wire w_dff_B_gBhgOVnT1_2;
	wire w_dff_B_89y1K2Xs8_2;
	wire w_dff_B_mk4QHZQS7_2;
	wire w_dff_B_SAOoRhsC9_1;
	wire w_dff_B_XjefX4721_2;
	wire w_dff_B_NolhAyI60_2;
	wire w_dff_B_5Ux9wGwm5_2;
	wire w_dff_B_LD6nPV3L0_2;
	wire w_dff_B_qi2cPUYf2_2;
	wire w_dff_B_EnY0yLLv9_2;
	wire w_dff_B_aKQqJcDg9_2;
	wire w_dff_B_ZClTf7qy1_2;
	wire w_dff_B_IpAfcqwl0_2;
	wire w_dff_B_mrKCDw2q9_2;
	wire w_dff_B_U08s84Q54_2;
	wire w_dff_B_YVAuNIrv0_2;
	wire w_dff_B_0LxnTeCw2_2;
	wire w_dff_B_9xHkYdKc0_2;
	wire w_dff_B_l4Mnnc7U8_2;
	wire w_dff_B_W0QLLP3E9_2;
	wire w_dff_B_kJ4UVvww1_2;
	wire w_dff_B_iYxINs7f7_2;
	wire w_dff_B_IS2dR1B27_2;
	wire w_dff_B_7k2RvW6g1_2;
	wire w_dff_B_v75OYDqx0_2;
	wire w_dff_B_f3JmymHX2_2;
	wire w_dff_B_xnqkOxxm0_2;
	wire w_dff_B_s6uW2cIn2_2;
	wire w_dff_B_XRBAfsxD8_2;
	wire w_dff_B_YwwbrA3T6_2;
	wire w_dff_B_ndj0dHNJ8_2;
	wire w_dff_B_6bjCgydK2_2;
	wire w_dff_B_vpcUPsY24_2;
	wire w_dff_B_3eIUFEBL4_2;
	wire w_dff_B_yz6ItiD02_2;
	wire w_dff_B_OYI5TTQ27_2;
	wire w_dff_B_sEVUrz8g0_2;
	wire w_dff_B_4P5mUltv6_2;
	wire w_dff_B_TCdl79rD8_1;
	wire w_dff_B_edWN1NhW4_2;
	wire w_dff_B_HHx47qXL1_2;
	wire w_dff_B_rc7qgt0a3_2;
	wire w_dff_B_dIWe51b91_2;
	wire w_dff_B_HHe1uSsr2_2;
	wire w_dff_B_UUMlViDm1_2;
	wire w_dff_B_FACeCpGh4_2;
	wire w_dff_B_FRwGckXt5_2;
	wire w_dff_B_1DapE0cs9_2;
	wire w_dff_B_JVZC70tZ0_2;
	wire w_dff_B_ljxaKdkG0_2;
	wire w_dff_B_VOthYxX98_2;
	wire w_dff_B_fdfOxRjd5_2;
	wire w_dff_B_XKiqIZ5r4_2;
	wire w_dff_B_NeSmKgSE2_2;
	wire w_dff_B_F3SclU8R3_2;
	wire w_dff_B_XSyHIbcY0_2;
	wire w_dff_B_4LHxSwYK3_2;
	wire w_dff_B_P187kyDT4_2;
	wire w_dff_B_v0lmHB5I7_2;
	wire w_dff_B_wVKtpP5L9_2;
	wire w_dff_B_vYdEo0Fz2_2;
	wire w_dff_B_hz8Uspyn5_2;
	wire w_dff_B_zRU4CEaB0_2;
	wire w_dff_B_5zbn9sFc5_2;
	wire w_dff_B_7ubZMhHE7_2;
	wire w_dff_B_7EEoPkXK2_2;
	wire w_dff_B_VsStI1L86_2;
	wire w_dff_B_hT9Ev7Vt9_2;
	wire w_dff_B_qdYNCKvA2_2;
	wire w_dff_B_QsPz98oR1_1;
	wire w_dff_B_GrRxEaNu6_2;
	wire w_dff_B_rEGRSoG71_2;
	wire w_dff_B_tGa8r5Lc4_2;
	wire w_dff_B_ejkEqu0H3_2;
	wire w_dff_B_2NN5B2kf0_2;
	wire w_dff_B_RHDjHqwB8_2;
	wire w_dff_B_QEiEL3mN7_2;
	wire w_dff_B_JJKIdqw52_2;
	wire w_dff_B_OUNeJMVY8_2;
	wire w_dff_B_xkoXLOF85_2;
	wire w_dff_B_Jed5Tjm11_2;
	wire w_dff_B_mp4F1oZH8_2;
	wire w_dff_B_eEJfo6TG8_2;
	wire w_dff_B_RO0EvG131_2;
	wire w_dff_B_0hbscURz9_2;
	wire w_dff_B_uErcEyIz3_2;
	wire w_dff_B_8wOoISR05_2;
	wire w_dff_B_fKU9188e7_2;
	wire w_dff_B_ZbKGSvYT9_2;
	wire w_dff_B_MqbE7NgF3_2;
	wire w_dff_B_OoAHvFgV5_2;
	wire w_dff_B_qf2DMypr4_2;
	wire w_dff_B_pMKCDJvG9_2;
	wire w_dff_B_VrZdiStE9_2;
	wire w_dff_B_7bdxXkSP7_2;
	wire w_dff_B_c1BRs3pm3_2;
	wire w_dff_B_f3NceXEh7_1;
	wire w_dff_B_lCx35bWy3_2;
	wire w_dff_B_AztIEZv59_2;
	wire w_dff_B_d7TUXjew0_2;
	wire w_dff_B_k9Jg1eEh3_2;
	wire w_dff_B_124TKauY1_2;
	wire w_dff_B_mOF0fu9Y5_2;
	wire w_dff_B_Kl3R1ejy5_2;
	wire w_dff_B_qfbSuO2U5_2;
	wire w_dff_B_iPLNtMfH4_2;
	wire w_dff_B_LFvrOSLM2_2;
	wire w_dff_B_y5xnIrsl7_2;
	wire w_dff_B_KiJengFT6_2;
	wire w_dff_B_Ha11kADe9_2;
	wire w_dff_B_UrtMm4fC2_2;
	wire w_dff_B_n98Zh5Uc4_2;
	wire w_dff_B_6BtnarNa7_2;
	wire w_dff_B_WIL0cb5J4_2;
	wire w_dff_B_NqJgbb3l5_2;
	wire w_dff_B_bPKMX1LZ2_2;
	wire w_dff_B_gOxNeTZb8_2;
	wire w_dff_B_3XfacPBE0_2;
	wire w_dff_B_Za8DoiXy7_1;
	wire w_dff_B_r5fzfAxf9_2;
	wire w_dff_B_ePE49Jzy5_2;
	wire w_dff_B_Ve2RcBtt0_2;
	wire w_dff_B_Mz06rtE93_2;
	wire w_dff_B_9CMdKNfD5_2;
	wire w_dff_B_b8GLL0Nk3_2;
	wire w_dff_B_h7pYsV878_2;
	wire w_dff_B_lE00m7Z73_2;
	wire w_dff_B_eRPL2gmp0_2;
	wire w_dff_B_a6kvGCiD9_2;
	wire w_dff_B_L9TnrSUB8_2;
	wire w_dff_B_baOIVWVp9_2;
	wire w_dff_B_R8slybch4_2;
	wire w_dff_B_6hbSk1TN9_2;
	wire w_dff_B_ddo9L6QE0_2;
	wire w_dff_B_MczcRKuC2_2;
	wire w_dff_B_nvfTUSFu6_2;
	wire w_dff_B_Xiu0xkK29_2;
	wire w_dff_B_msSltTL19_2;
	wire w_dff_B_af6URBAC0_1;
	wire w_dff_B_oYP1l3rM5_2;
	wire w_dff_B_gRf78oQM8_2;
	wire w_dff_B_tgN7iGGJ7_2;
	wire w_dff_B_l7CesZvX9_2;
	wire w_dff_B_ezaZEJrp5_2;
	wire w_dff_B_RfHQRe791_2;
	wire w_dff_B_dsUBNTIy8_2;
	wire w_dff_B_nWAzqlwX2_2;
	wire w_dff_B_RaF2pSzQ5_2;
	wire w_dff_B_VZxdJc120_2;
	wire w_dff_B_L5Z5gPi44_2;
	wire w_dff_B_Px5rwGni0_2;
	wire w_dff_B_sbDZY1tI2_2;
	wire w_dff_B_WtGIh4183_2;
	wire w_dff_B_9P0YEedD2_2;
	wire w_dff_B_RSnN9Bqc6_2;
	wire w_dff_B_GbnFbinF7_2;
	wire w_dff_B_JdMX0b1g2_1;
	wire w_dff_B_eeCbMqGg7_2;
	wire w_dff_B_z1LRiTOE0_2;
	wire w_dff_B_gv3NYn6P6_2;
	wire w_dff_B_1ENQgEHy7_2;
	wire w_dff_B_vijbYQq07_2;
	wire w_dff_B_BhQpaSSH3_2;
	wire w_dff_B_CBo7bbq76_2;
	wire w_dff_B_JYBkCv3n7_2;
	wire w_dff_B_edUcnAT04_2;
	wire w_dff_B_yHYHauRk5_2;
	wire w_dff_B_eCVnUcVL2_2;
	wire w_dff_B_RN7mN8hd4_2;
	wire w_dff_B_DOAQMQjL2_2;
	wire w_dff_B_QkUk3v3e1_2;
	wire w_dff_B_PJf0cWwu9_1;
	wire w_dff_B_h9kLTsBE7_2;
	wire w_dff_B_3IuYWM1f7_2;
	wire w_dff_B_ZSeLQX9n7_2;
	wire w_dff_B_nGXJ12E88_2;
	wire w_dff_B_HdZ7ZILy2_2;
	wire w_dff_B_xWtGqVjE0_2;
	wire w_dff_B_aTqj50vP2_2;
	wire w_dff_B_FKjZDHFt8_2;
	wire w_dff_B_PJROlhI89_2;
	wire w_dff_B_WNF3HEs58_2;
	wire w_dff_B_6IN4EJlK2_2;
	wire w_dff_B_sYNSHnuN6_2;
	wire w_dff_B_yTJ3of4o1_1;
	wire w_dff_B_7Qv96jdo5_1;
	wire w_dff_B_qojY8BTd6_1;
	wire w_dff_B_3WH9b8qn6_1;
	wire w_dff_B_l0OJj6WW6_1;
	wire w_dff_B_Q36U5tAt1_1;
	wire w_dff_B_UmxfwUrb4_0;
	wire w_dff_B_l1FIUshX7_0;
	wire w_dff_A_IZ0xkOZa6_0;
	wire w_dff_A_Vp1im4IS8_0;
	wire w_dff_A_xxdJDKKt3_0;
	wire w_dff_B_fexZ1vyZ4_1;
	wire w_dff_A_PWnxLbLl4_0;
	wire w_dff_A_sW6BxUtj5_1;
	wire w_dff_A_j2EXnS4j2_1;
	wire w_dff_A_Bng07JI51_1;
	wire w_dff_A_DMRk3z007_1;
	wire w_dff_A_FPrhdtpG5_1;
	wire w_dff_A_kH63j8y58_1;
	wire w_dff_A_N3X0YXy17_1;
	wire w_dff_A_YFE1FYKA7_1;
	wire w_dff_B_G1Be0w1L8_1;
	wire w_dff_B_BJk9Dbvo7_1;
	wire w_dff_B_AxN3HC4J1_1;
	wire w_dff_B_9vMD6hbD0_2;
	wire w_dff_B_iR3Wwocn7_2;
	wire w_dff_B_y2CLNKJg3_2;
	wire w_dff_B_thMdE1km3_2;
	wire w_dff_B_gqRyL4kK8_2;
	wire w_dff_B_2A6sBGJO0_2;
	wire w_dff_B_1FX43Tc53_2;
	wire w_dff_B_6x2Ex84T7_2;
	wire w_dff_B_LYPyE8tY2_2;
	wire w_dff_B_zVhitRX36_2;
	wire w_dff_B_mtiAUmNd6_2;
	wire w_dff_B_7SoSryC90_2;
	wire w_dff_B_fP3eqyak0_2;
	wire w_dff_B_njOaAzGI0_2;
	wire w_dff_B_7tPl8Cjy8_2;
	wire w_dff_B_v8BIbjAg8_2;
	wire w_dff_B_StLRGRLP9_2;
	wire w_dff_B_QfVDqDwH8_2;
	wire w_dff_B_B3KWInmO7_2;
	wire w_dff_B_M7DCY9k03_2;
	wire w_dff_B_rAUwfWYI2_2;
	wire w_dff_B_52iviQen5_2;
	wire w_dff_B_nYhK47Pe4_2;
	wire w_dff_B_ETSoEChk3_2;
	wire w_dff_B_wJZ6jOMz5_2;
	wire w_dff_B_MnNlc0Ou7_2;
	wire w_dff_B_tEmivrTT0_2;
	wire w_dff_B_cE7dGaTG7_2;
	wire w_dff_B_eBmY3vh63_2;
	wire w_dff_B_UqrvQW5a4_2;
	wire w_dff_B_9S1WPhc23_2;
	wire w_dff_B_sgCui1Oh6_2;
	wire w_dff_B_dFFw3xfX4_2;
	wire w_dff_B_KykwPUDp1_2;
	wire w_dff_B_6nFXMZBp9_2;
	wire w_dff_B_Q4CBMmkC9_2;
	wire w_dff_B_UC5kuJaV0_2;
	wire w_dff_B_1fdUktiK4_2;
	wire w_dff_B_Pmflzgv54_2;
	wire w_dff_B_zhUTe2rp2_2;
	wire w_dff_B_D2PBaTFe8_2;
	wire w_dff_B_sH9z1PyZ3_2;
	wire w_dff_B_MvYL5r789_2;
	wire w_dff_B_5BFebvs10_2;
	wire w_dff_B_PULcOqeB0_2;
	wire w_dff_B_gXqmDAeT8_2;
	wire w_dff_B_xgFFtDeH6_2;
	wire w_dff_B_3H1iyCRn6_2;
	wire w_dff_B_06s29llU5_2;
	wire w_dff_B_NCg4KGXy8_2;
	wire w_dff_B_aDtcJ0ba2_2;
	wire w_dff_B_DBu9MS8x8_2;
	wire w_dff_B_WqK2XOQa0_2;
	wire w_dff_B_K12XMtUH4_2;
	wire w_dff_B_NX47Qo9X3_2;
	wire w_dff_B_1EHsxoj72_2;
	wire w_dff_B_XFzugYOA1_2;
	wire w_dff_B_T28lCIe81_2;
	wire w_dff_B_wkflulbq7_2;
	wire w_dff_B_U5frjtpA6_2;
	wire w_dff_B_O6i7BYTM1_2;
	wire w_dff_B_rwByXSln1_2;
	wire w_dff_B_rtwrQ7Tv5_2;
	wire w_dff_B_HDbnImm39_2;
	wire w_dff_B_AaMS8tfn6_2;
	wire w_dff_B_pVk1HtIl5_2;
	wire w_dff_B_FAc6RLLw4_2;
	wire w_dff_B_1TFpC6D21_2;
	wire w_dff_B_PfAeb9oB3_2;
	wire w_dff_B_MVQii1Gd8_2;
	wire w_dff_B_Djsn6kpn7_2;
	wire w_dff_B_xexikIMK3_2;
	wire w_dff_B_ggMbpQ1Y0_2;
	wire w_dff_B_vCgWseQY3_2;
	wire w_dff_B_JdEPa84d2_2;
	wire w_dff_B_4BkPHsBH0_2;
	wire w_dff_B_vHAFnp5x2_2;
	wire w_dff_B_nBcdnM9J5_2;
	wire w_dff_B_mqHpdWmB4_2;
	wire w_dff_B_XxhIOBW03_2;
	wire w_dff_B_YerTaQ5M3_2;
	wire w_dff_B_5qeh0qTg4_2;
	wire w_dff_B_N5mK56Ne9_2;
	wire w_dff_B_YvHSALV81_2;
	wire w_dff_B_SVjep5Kl0_2;
	wire w_dff_B_i2mWbpK86_2;
	wire w_dff_B_FxwMyqUs3_2;
	wire w_dff_B_cxmOkPJ61_2;
	wire w_dff_B_dyIoaoXw8_2;
	wire w_dff_B_SflPcyWR9_2;
	wire w_dff_B_jrItXETU6_2;
	wire w_dff_B_WK2EgIWG3_2;
	wire w_dff_B_xFAOHMdw9_2;
	wire w_dff_B_dhnAj0hT9_2;
	wire w_dff_B_QTDhhjWn0_2;
	wire w_dff_B_lN3EfoVL0_2;
	wire w_dff_B_8s5o3v5U4_2;
	wire w_dff_B_qde6tAky2_2;
	wire w_dff_B_In3gVkjm5_2;
	wire w_dff_B_STu83squ6_2;
	wire w_dff_B_gfdF8Odu5_2;
	wire w_dff_B_oyiBnt7S7_2;
	wire w_dff_B_ix5DV3Pj9_2;
	wire w_dff_B_DQziWUWh7_2;
	wire w_dff_B_tKKdVf3h6_2;
	wire w_dff_B_ZnvyxNqF0_2;
	wire w_dff_B_bVUR7K3M1_2;
	wire w_dff_B_NfQ7qjpF1_2;
	wire w_dff_B_KvjGBq3E4_2;
	wire w_dff_B_PFWPYXhD6_2;
	wire w_dff_B_JwSfpbBe7_2;
	wire w_dff_B_JRF5aHui3_2;
	wire w_dff_B_n6ngT6Yo2_2;
	wire w_dff_B_eP2sF8fc1_2;
	wire w_dff_A_Gl0YM9RQ1_1;
	wire w_dff_B_mgjKK9GJ3_1;
	wire w_dff_B_SCL5FPKf3_2;
	wire w_dff_B_rzXmh0BJ1_2;
	wire w_dff_B_qeZt0Tgx5_2;
	wire w_dff_B_f3WvnnPU4_2;
	wire w_dff_B_NyTNzeqe7_2;
	wire w_dff_B_bu82JbmM1_2;
	wire w_dff_B_PtMZMIJq2_2;
	wire w_dff_B_iAqmL0DB6_2;
	wire w_dff_B_ljIttL9l9_2;
	wire w_dff_B_nxCSWGlt7_2;
	wire w_dff_B_qwNFtUbC2_2;
	wire w_dff_B_eX9ZyAfw3_2;
	wire w_dff_B_d40C5jOH5_2;
	wire w_dff_B_QYCke47w0_2;
	wire w_dff_B_O7ZtqB7H8_2;
	wire w_dff_B_buJwVWIL1_2;
	wire w_dff_B_4wdRDvXP7_2;
	wire w_dff_B_M027ArTJ2_2;
	wire w_dff_B_IgbOy04R6_2;
	wire w_dff_B_JKKOcUY14_2;
	wire w_dff_B_uOyyPRu64_2;
	wire w_dff_B_Qq5pQ5Py1_2;
	wire w_dff_B_RNL4Jt5w8_2;
	wire w_dff_B_mDVG1MSg6_2;
	wire w_dff_B_qPSvWAOh0_2;
	wire w_dff_B_0OTCxfDP5_2;
	wire w_dff_B_e3nTQoLs9_2;
	wire w_dff_B_tpHaKlcI8_2;
	wire w_dff_B_2ux7tTVC2_2;
	wire w_dff_B_pVz0MthM3_2;
	wire w_dff_B_xpITjV6J8_2;
	wire w_dff_B_zCFukkEW2_2;
	wire w_dff_B_6GVByEGo9_2;
	wire w_dff_B_PzF4wiI91_2;
	wire w_dff_B_PZRbMNPF1_2;
	wire w_dff_B_wE8M9pSE6_2;
	wire w_dff_B_sxF7Nnto4_2;
	wire w_dff_B_0s4hG60m4_2;
	wire w_dff_B_5h7NepSj5_2;
	wire w_dff_B_pop4QW1h9_2;
	wire w_dff_B_upAQuHGD9_2;
	wire w_dff_B_vnGnmv5D6_2;
	wire w_dff_B_WsEJNZR41_2;
	wire w_dff_B_t8NUpRFL8_2;
	wire w_dff_B_n4UBlc7K0_2;
	wire w_dff_B_9QpmV5qC5_2;
	wire w_dff_B_LTNHYBTm5_2;
	wire w_dff_B_yZxKMZrc0_2;
	wire w_dff_B_t5UhvOzR9_2;
	wire w_dff_B_u4xfTwzc5_2;
	wire w_dff_B_f5WMARNu2_2;
	wire w_dff_B_kqOINCaK6_2;
	wire w_dff_B_pZhfJMe73_2;
	wire w_dff_B_DDLXVTVi5_2;
	wire w_dff_B_iy3NUKPE5_2;
	wire w_dff_B_C5PFZR9b4_1;
	wire w_dff_B_HF7UIH5v7_1;
	wire w_dff_B_wHsykZ4H0_2;
	wire w_dff_B_zhuPOkfj8_2;
	wire w_dff_B_0XaTQvYi4_2;
	wire w_dff_B_yDLhR7300_2;
	wire w_dff_B_Eex5LyVM5_2;
	wire w_dff_B_6ZvvSzvv7_2;
	wire w_dff_B_U9JaiPV90_2;
	wire w_dff_B_3HEWHJvJ7_2;
	wire w_dff_B_5tC6oTRG6_2;
	wire w_dff_B_kaXIRbLv3_2;
	wire w_dff_B_CP6JXgNu9_2;
	wire w_dff_B_gzs4q0lq2_2;
	wire w_dff_B_3esntLel3_2;
	wire w_dff_B_V4mb45DA0_2;
	wire w_dff_B_BelUqyhy5_2;
	wire w_dff_B_6H5KFKj60_2;
	wire w_dff_B_s8QpbDgg2_2;
	wire w_dff_B_U7g7E0915_2;
	wire w_dff_B_HQwyle1y5_2;
	wire w_dff_B_0TwLzO5A5_2;
	wire w_dff_B_jmKALU6T0_2;
	wire w_dff_B_eBUFuLKM9_2;
	wire w_dff_B_33O9jhYA3_2;
	wire w_dff_B_YJDYGVz93_2;
	wire w_dff_B_pG3Im42M8_2;
	wire w_dff_B_IST5TWf49_2;
	wire w_dff_B_Tl1UPHVz1_2;
	wire w_dff_B_oNE4NWWT9_2;
	wire w_dff_B_lyFbzixm0_2;
	wire w_dff_B_TocHg3WY7_2;
	wire w_dff_B_3cBaZWW75_2;
	wire w_dff_B_SDyoQ5iT4_2;
	wire w_dff_B_64TKNjo47_2;
	wire w_dff_B_uyHq7NzC1_2;
	wire w_dff_B_ZoiUq8a02_2;
	wire w_dff_B_Ba850tM69_2;
	wire w_dff_B_mnXNmXzB8_2;
	wire w_dff_B_4gS6xnRA7_2;
	wire w_dff_B_EbhUxANj2_2;
	wire w_dff_B_vuE5VV8D4_2;
	wire w_dff_B_eT333xhz5_2;
	wire w_dff_B_467KL0ma9_2;
	wire w_dff_B_0qy5Wpy23_2;
	wire w_dff_B_eFqEJzwg6_2;
	wire w_dff_B_a8QS7p6D1_2;
	wire w_dff_B_QPsg3qiV0_2;
	wire w_dff_B_VjQUnkm02_2;
	wire w_dff_B_Xv7fqjh14_2;
	wire w_dff_B_KY5ozMdg9_2;
	wire w_dff_B_fD031rCq7_2;
	wire w_dff_B_E57eyS4L2_2;
	wire w_dff_B_qDLH0N856_2;
	wire w_dff_B_2fPJuVhx8_2;
	wire w_dff_B_7dzdvXTd5_2;
	wire w_dff_B_0VyNcSpR3_2;
	wire w_dff_B_1P0ZU3AO1_2;
	wire w_dff_B_9eR9o1238_2;
	wire w_dff_B_Lt9yd9Dk1_2;
	wire w_dff_B_UuhZQnPW4_2;
	wire w_dff_B_bYhuYC8K5_2;
	wire w_dff_B_tCOv0GtU3_2;
	wire w_dff_B_LkK62bDd0_2;
	wire w_dff_B_FdqfFCXn2_2;
	wire w_dff_B_hxVovnc37_2;
	wire w_dff_B_tFMXEZ056_2;
	wire w_dff_B_YG1uLtQO4_2;
	wire w_dff_B_NIhudi1f7_2;
	wire w_dff_B_FBxUjoSz5_2;
	wire w_dff_B_c7fpcYcG8_2;
	wire w_dff_B_5NAKAHfi0_2;
	wire w_dff_B_P6j1z3zi3_2;
	wire w_dff_B_eaU1Od7X3_2;
	wire w_dff_B_luTLKIV70_2;
	wire w_dff_B_czYanEhE8_2;
	wire w_dff_B_X6ighRgX3_2;
	wire w_dff_B_asnk09Ta4_2;
	wire w_dff_B_ijlB5QAU4_2;
	wire w_dff_B_hmkodBnU9_2;
	wire w_dff_B_9m5MlGyv0_2;
	wire w_dff_B_oEHLFViE1_2;
	wire w_dff_B_7IopQFbk8_2;
	wire w_dff_B_FJXngTPx4_2;
	wire w_dff_B_CcvmYj4K1_2;
	wire w_dff_B_IcljosVj9_2;
	wire w_dff_B_D3OS0tOl8_2;
	wire w_dff_B_vLq7xXXe6_2;
	wire w_dff_B_Cxlbn2YH1_2;
	wire w_dff_B_bYDkw8ey7_2;
	wire w_dff_B_YsVtuTww3_2;
	wire w_dff_B_zeQHvMfS1_2;
	wire w_dff_B_xh3h0ZTH5_2;
	wire w_dff_B_Bxbj5GNR9_2;
	wire w_dff_B_DDQoObtD0_2;
	wire w_dff_B_WPWPEX9p4_2;
	wire w_dff_B_qe5l42G07_2;
	wire w_dff_B_5NwC0zyT1_2;
	wire w_dff_B_XMJKtRfu1_2;
	wire w_dff_B_gPYNN6We1_2;
	wire w_dff_B_4X61qpGa9_2;
	wire w_dff_B_g88UkIkL3_2;
	wire w_dff_B_xm3ajwH93_2;
	wire w_dff_B_LgYseWrf1_2;
	wire w_dff_B_fwwxPM7b0_2;
	wire w_dff_B_oawvuwEe3_2;
	wire w_dff_B_smj7f7QK1_2;
	wire w_dff_B_eAyBbxsi5_2;
	wire w_dff_B_qwcLaNmX5_2;
	wire w_dff_B_DCVTibQ27_1;
	wire w_dff_B_mBr9zinK6_2;
	wire w_dff_B_LULJaJzn4_2;
	wire w_dff_B_sUAEr5C76_2;
	wire w_dff_B_7O0dQzBl7_2;
	wire w_dff_B_2bRqSR7K4_2;
	wire w_dff_B_9oiuXmBM5_2;
	wire w_dff_B_CWyPJmsp1_2;
	wire w_dff_B_JQClPjCb6_2;
	wire w_dff_B_vmLGuPmO0_2;
	wire w_dff_B_M3aP8gb95_2;
	wire w_dff_B_wV5zPB190_2;
	wire w_dff_B_sjcZzzYF5_2;
	wire w_dff_B_430T1Hu07_2;
	wire w_dff_B_W97Gox2J2_2;
	wire w_dff_B_y0f3K5dY3_2;
	wire w_dff_B_6msuEzT60_2;
	wire w_dff_B_b4ApuG0W5_2;
	wire w_dff_B_f0i7id6f0_2;
	wire w_dff_B_fy0ZoZUL7_2;
	wire w_dff_B_DjY4juBD1_2;
	wire w_dff_B_NP1GV6ld1_2;
	wire w_dff_B_paD3DpxO7_2;
	wire w_dff_B_sDHHtcpz7_2;
	wire w_dff_B_wjppf0Bc1_2;
	wire w_dff_B_lbLrs8LF4_2;
	wire w_dff_B_L0DmwOYo7_2;
	wire w_dff_B_Ft5TVyL50_2;
	wire w_dff_B_9aue72Ua0_2;
	wire w_dff_B_cIwxU3zM3_2;
	wire w_dff_B_RHqIKApR7_2;
	wire w_dff_B_ujN89r0g6_2;
	wire w_dff_B_wvxQYmri1_2;
	wire w_dff_B_ePiEQjG64_2;
	wire w_dff_B_GrU9M4Jm8_2;
	wire w_dff_B_6f4JRWgK8_2;
	wire w_dff_B_D5mwCWO32_2;
	wire w_dff_B_xl4p3TSt5_2;
	wire w_dff_B_9GkEsjpZ8_2;
	wire w_dff_B_lAUcFlBh4_2;
	wire w_dff_B_DOaNXmBB7_2;
	wire w_dff_B_2MlMu2sh8_2;
	wire w_dff_B_74oQAdo70_2;
	wire w_dff_B_3wHcWuwi0_2;
	wire w_dff_B_R67BSxLW1_2;
	wire w_dff_B_Vw8N4D9R7_2;
	wire w_dff_B_00ZDp0qO0_2;
	wire w_dff_B_52nWTJBW9_2;
	wire w_dff_B_gh6p9pkQ1_2;
	wire w_dff_B_ov1qn2jK9_2;
	wire w_dff_B_gKuxhXwY3_2;
	wire w_dff_B_KRSHZt2L9_2;
	wire w_dff_B_1pa574RV7_1;
	wire w_dff_B_ab685Q2h6_1;
	wire w_dff_B_ZTQGXS6I4_2;
	wire w_dff_B_Lx3mjdSi3_2;
	wire w_dff_B_2yMd3pmf8_2;
	wire w_dff_B_GvLXw1Dy4_2;
	wire w_dff_B_Y34VWZRz1_2;
	wire w_dff_B_ASvUhJ8E6_2;
	wire w_dff_B_0DR97vdd7_2;
	wire w_dff_B_mhEG4gnA9_2;
	wire w_dff_B_NiVKBVR14_2;
	wire w_dff_B_zg14c5Ki7_2;
	wire w_dff_B_KW35wHnr4_2;
	wire w_dff_B_Lr2extkt9_2;
	wire w_dff_B_dTuSMScV1_2;
	wire w_dff_B_HUyS1SZJ5_2;
	wire w_dff_B_wi4EoFSo0_2;
	wire w_dff_B_JBWjeKvm9_2;
	wire w_dff_B_nPHj5vVo7_2;
	wire w_dff_B_zboqbU9m7_2;
	wire w_dff_B_Dpr5pW0F1_2;
	wire w_dff_B_4Rt9FTG91_2;
	wire w_dff_B_poSUiAYG0_2;
	wire w_dff_B_kIyNPvVA4_2;
	wire w_dff_B_jTSwfXPJ8_2;
	wire w_dff_B_nOxYfUo26_2;
	wire w_dff_B_h8cPlX6y5_2;
	wire w_dff_B_WPqMUme29_2;
	wire w_dff_B_MI5UAQtl8_2;
	wire w_dff_B_WRtTMCzU1_2;
	wire w_dff_B_5n4V0OA64_2;
	wire w_dff_B_O4WLllGz5_2;
	wire w_dff_B_qP2Freca0_2;
	wire w_dff_B_aYAGfY9R4_2;
	wire w_dff_B_HQbZyGRz8_2;
	wire w_dff_B_6XQUihbW8_2;
	wire w_dff_B_Hn32oo9u0_2;
	wire w_dff_B_aYmWKJlS1_2;
	wire w_dff_B_RddqjjSj7_2;
	wire w_dff_B_KzTHHdTZ9_2;
	wire w_dff_B_LQMIU07m6_2;
	wire w_dff_B_ANxyz6Kb5_2;
	wire w_dff_B_NCvwvwDQ1_2;
	wire w_dff_B_8ZyEKesh8_2;
	wire w_dff_B_12TJV3oR1_2;
	wire w_dff_B_6pviUdXw0_2;
	wire w_dff_B_Lgp6UKpm6_2;
	wire w_dff_B_vPpUmE0L7_2;
	wire w_dff_B_JTOL4DZN6_2;
	wire w_dff_B_T0DnmlcE6_2;
	wire w_dff_B_UTRszQtn2_2;
	wire w_dff_B_Cr8357xq0_2;
	wire w_dff_B_QZf6fSZk6_2;
	wire w_dff_B_KPhStNhc8_2;
	wire w_dff_B_vWPu9wjV8_2;
	wire w_dff_B_YYYBmQsF7_2;
	wire w_dff_B_ePWIeJ7V6_2;
	wire w_dff_B_bzgpolVd7_2;
	wire w_dff_B_JbbDq3Bd9_2;
	wire w_dff_B_05NofmFR7_2;
	wire w_dff_B_grb6c2iX6_2;
	wire w_dff_B_3T42BwSA4_2;
	wire w_dff_B_6MX5TUvy2_2;
	wire w_dff_B_vhJlguC05_2;
	wire w_dff_B_e7b6DkQD1_2;
	wire w_dff_B_Jlhw6XOj4_2;
	wire w_dff_B_BztSFJGT6_2;
	wire w_dff_B_WCvndrbo4_2;
	wire w_dff_B_O0eLY8gG7_2;
	wire w_dff_B_XRz4o72X2_2;
	wire w_dff_B_gdE9GhUH5_2;
	wire w_dff_B_owaIawDw8_2;
	wire w_dff_B_4DSfg6gF5_2;
	wire w_dff_B_2NbcAh0T1_2;
	wire w_dff_B_gdSaeRLj7_2;
	wire w_dff_B_9HrCLUZ11_2;
	wire w_dff_B_pm2HzBRZ3_2;
	wire w_dff_B_bGsG0aH45_2;
	wire w_dff_B_4EO0Me7n0_2;
	wire w_dff_B_xAwSMO3D1_2;
	wire w_dff_B_z2EjJ4dY6_2;
	wire w_dff_B_WsrsDtnA7_2;
	wire w_dff_B_Njbn7fqq4_2;
	wire w_dff_B_5El2Biyu2_2;
	wire w_dff_B_bYCIXVhK1_2;
	wire w_dff_B_Yq0xn5UJ7_2;
	wire w_dff_B_Sxnc3k794_2;
	wire w_dff_B_WM4jHbNO0_2;
	wire w_dff_B_8k2UQPcp3_2;
	wire w_dff_B_CQGVIHtp5_2;
	wire w_dff_B_WqHq0ZFJ8_2;
	wire w_dff_B_awSFrf515_2;
	wire w_dff_B_rlXqutju2_2;
	wire w_dff_B_inKx7PGA4_2;
	wire w_dff_B_RWuu1e251_2;
	wire w_dff_B_5rGmhKVO8_2;
	wire w_dff_B_dzzTHMoz6_2;
	wire w_dff_B_eIn0hFC26_2;
	wire w_dff_B_DigdRgnJ2_2;
	wire w_dff_B_qFmd4odf4_2;
	wire w_dff_B_agF8t62T8_2;
	wire w_dff_B_3hVnrSk46_1;
	wire w_dff_B_5T2MMC6t4_2;
	wire w_dff_B_jHJYw1tZ2_2;
	wire w_dff_B_ipwt0XsT6_2;
	wire w_dff_B_1eZUEalB9_2;
	wire w_dff_B_ZLREOlSh2_2;
	wire w_dff_B_3WHtvTS26_2;
	wire w_dff_B_r3UPrdIk0_2;
	wire w_dff_B_30ZujImX2_2;
	wire w_dff_B_LuAgpGXj1_2;
	wire w_dff_B_CueCAGRS1_2;
	wire w_dff_B_rR8nMODP8_2;
	wire w_dff_B_vlA4WHrT9_2;
	wire w_dff_B_hNPXYkr54_2;
	wire w_dff_B_CbJP7g9z3_2;
	wire w_dff_B_l7GiGpvr5_2;
	wire w_dff_B_TlmxsKRL8_2;
	wire w_dff_B_9TkOdnhg8_2;
	wire w_dff_B_o0H4G08Y3_2;
	wire w_dff_B_XlcvIfD08_2;
	wire w_dff_B_Rmq9Dlrt6_2;
	wire w_dff_B_fu5VFzlx7_2;
	wire w_dff_B_wIA6K3Ev7_2;
	wire w_dff_B_ub2kmoWX3_2;
	wire w_dff_B_U2zk2YV07_2;
	wire w_dff_B_aYTXs1Rt6_2;
	wire w_dff_B_4RGwT7B56_2;
	wire w_dff_B_opA2uA8u9_2;
	wire w_dff_B_znimIONV6_2;
	wire w_dff_B_0Is8eCHY6_2;
	wire w_dff_B_tqvDZqSD6_2;
	wire w_dff_B_fO3nrgpd7_2;
	wire w_dff_B_bVnvuLRV5_2;
	wire w_dff_B_peI1zMN58_2;
	wire w_dff_B_uVS5ZH7X4_2;
	wire w_dff_B_m8kkNvOa9_2;
	wire w_dff_B_zMTkOWJj4_2;
	wire w_dff_B_4VO5xxc52_2;
	wire w_dff_B_rsDZjJQp9_2;
	wire w_dff_B_Xx1zgopg7_2;
	wire w_dff_B_UJiMHZ1T7_2;
	wire w_dff_B_CqfMuxuq4_2;
	wire w_dff_B_fQriyvUs6_2;
	wire w_dff_B_rbfuiNGA4_2;
	wire w_dff_B_0L2gbH7y8_2;
	wire w_dff_B_IQenXnjK5_2;
	wire w_dff_B_gVBE3rh19_2;
	wire w_dff_B_DyB1IKPC5_2;
	wire w_dff_B_qT5sAETC5_1;
	wire w_dff_B_ITq5ODvv5_1;
	wire w_dff_B_sqPDmQhi6_2;
	wire w_dff_B_XHC47qVA8_2;
	wire w_dff_B_Lcsrw7ZW2_2;
	wire w_dff_B_AghjpGzh2_2;
	wire w_dff_B_AsT0YJje5_2;
	wire w_dff_B_jMrePLeH8_2;
	wire w_dff_B_Ra7XznvX7_2;
	wire w_dff_B_sPrRGCIl5_2;
	wire w_dff_B_9m5DIBku3_2;
	wire w_dff_B_wd47nu722_2;
	wire w_dff_B_kOheLc7A8_2;
	wire w_dff_B_UBxZJgp13_2;
	wire w_dff_B_W3z5arOG0_2;
	wire w_dff_B_nEPJvcAE5_2;
	wire w_dff_B_e9AZpvSL1_2;
	wire w_dff_B_34hCClRC5_2;
	wire w_dff_B_QtxlQDeo3_2;
	wire w_dff_B_A5G1GQsU1_2;
	wire w_dff_B_Z6WgYcih9_2;
	wire w_dff_B_Un0gvM0A3_2;
	wire w_dff_B_cEG43IBd2_2;
	wire w_dff_B_UmiKB51T9_2;
	wire w_dff_B_vmejwXTn7_2;
	wire w_dff_B_fBUGWA7r4_2;
	wire w_dff_B_RybLmypm7_2;
	wire w_dff_B_TrRCfxIc6_2;
	wire w_dff_B_NudGuLI28_2;
	wire w_dff_B_Udft1zug1_2;
	wire w_dff_B_bndFKDjV2_2;
	wire w_dff_B_tRLHHMq32_2;
	wire w_dff_B_6oO5qoZ88_2;
	wire w_dff_B_PPkq81yt1_2;
	wire w_dff_B_Up27UF968_2;
	wire w_dff_B_h8i0gn0l5_2;
	wire w_dff_B_pa97XfOY7_2;
	wire w_dff_B_9G0AjUt00_2;
	wire w_dff_B_hDkgm3b39_2;
	wire w_dff_B_gRhSfi7Y4_2;
	wire w_dff_B_kFbdzq0O6_2;
	wire w_dff_B_Vk0OT2gT7_2;
	wire w_dff_B_0NfvmgbE2_2;
	wire w_dff_B_IQFjwthz5_2;
	wire w_dff_B_MgjlpJUQ4_2;
	wire w_dff_B_XccXmWny7_2;
	wire w_dff_B_bIda4Wl94_2;
	wire w_dff_B_D2cKQdCD6_2;
	wire w_dff_B_WOviowce3_2;
	wire w_dff_B_RtvW9lIH1_2;
	wire w_dff_B_ngoc9Dr45_2;
	wire w_dff_B_yM6Mq15k2_2;
	wire w_dff_B_YYC0TVfN6_2;
	wire w_dff_B_LcvQ6Vel9_2;
	wire w_dff_B_Gj7zbwEj5_2;
	wire w_dff_B_NIhRWEWa3_2;
	wire w_dff_B_6RhbpRHq5_2;
	wire w_dff_B_xrjWXvYI5_2;
	wire w_dff_B_nOwczB7i9_2;
	wire w_dff_B_sw9dZln41_2;
	wire w_dff_B_zBpaf05x4_2;
	wire w_dff_B_HPBngvMO2_2;
	wire w_dff_B_V2xOTHGb5_2;
	wire w_dff_B_M9SZ4K9n7_2;
	wire w_dff_B_BVMznqHk9_2;
	wire w_dff_B_c1B8b2oY8_2;
	wire w_dff_B_idg30Hq10_2;
	wire w_dff_B_2RjKTG4C6_2;
	wire w_dff_B_ro5LUE5u7_2;
	wire w_dff_B_COgsj6Jh5_2;
	wire w_dff_B_IyAuwlPp5_2;
	wire w_dff_B_Iz5CJ1uM3_2;
	wire w_dff_B_HlG3ISFt2_2;
	wire w_dff_B_Rd4TqUI25_2;
	wire w_dff_B_cDI7qBXs5_2;
	wire w_dff_B_EqfTcMKK7_2;
	wire w_dff_B_dCEUnK2t6_2;
	wire w_dff_B_8Lpohban6_2;
	wire w_dff_B_3mIoPgG90_2;
	wire w_dff_B_0gNR8ukV1_2;
	wire w_dff_B_ZOUbpQuz2_2;
	wire w_dff_B_zi9iEQlJ1_2;
	wire w_dff_B_P4LaNWa51_2;
	wire w_dff_B_KWCFnulf0_2;
	wire w_dff_B_FqOHMpem9_2;
	wire w_dff_B_2Xg4DstL1_2;
	wire w_dff_B_1B3fioXq4_2;
	wire w_dff_B_SlOPBWUG4_2;
	wire w_dff_B_ZlrO80Xt4_2;
	wire w_dff_B_o2rqvsZX4_2;
	wire w_dff_B_DAygf4x11_2;
	wire w_dff_B_B7RNIbNT7_2;
	wire w_dff_B_0wdXCfdC9_2;
	wire w_dff_B_UFVwRiwo2_1;
	wire w_dff_B_4CbQx41F9_2;
	wire w_dff_B_tOzd0Gtu8_2;
	wire w_dff_B_3RK9jRb23_2;
	wire w_dff_B_aHLVSmPo4_2;
	wire w_dff_B_njx5V7RV3_2;
	wire w_dff_B_AWLuKZf47_2;
	wire w_dff_B_8yo0YQbD7_2;
	wire w_dff_B_R1JKiXfl3_2;
	wire w_dff_B_hPiNVPYx9_2;
	wire w_dff_B_xRtlWB7b4_2;
	wire w_dff_B_7g4ARltO2_2;
	wire w_dff_B_cl3vqZW91_2;
	wire w_dff_B_aifoDLxY3_2;
	wire w_dff_B_WZ7VcjL10_2;
	wire w_dff_B_6HbPTyBX3_2;
	wire w_dff_B_UlcXload6_2;
	wire w_dff_B_DWbaprGE6_2;
	wire w_dff_B_0v5qJSuu3_2;
	wire w_dff_B_rt0SGGiy8_2;
	wire w_dff_B_uYwP1HhH2_2;
	wire w_dff_B_8Gn5FTjb7_2;
	wire w_dff_B_thXTg66f1_2;
	wire w_dff_B_1C367qgX9_2;
	wire w_dff_B_d8ORhABr8_2;
	wire w_dff_B_5ixPI9vT5_2;
	wire w_dff_B_s2XpSyNf3_2;
	wire w_dff_B_FPkc7MQy5_2;
	wire w_dff_B_Lfo6DpxF6_2;
	wire w_dff_B_dgD72bWa6_2;
	wire w_dff_B_BY1kU5Ct4_2;
	wire w_dff_B_eFP3B0QO9_2;
	wire w_dff_B_HJR4GMn03_2;
	wire w_dff_B_pV2aBFeC8_2;
	wire w_dff_B_UM4RUzm44_2;
	wire w_dff_B_zr5HyVi01_2;
	wire w_dff_B_z2ACCUCN5_2;
	wire w_dff_B_szGS4o266_2;
	wire w_dff_B_gLEu3eWy3_2;
	wire w_dff_B_BMMSSA753_2;
	wire w_dff_B_BBLcp6S29_2;
	wire w_dff_B_9MIUmrvb4_2;
	wire w_dff_B_WvOsFQZ35_2;
	wire w_dff_B_YpBZ67h04_2;
	wire w_dff_B_YXZvJO2k0_1;
	wire w_dff_B_sl9LlNAT0_1;
	wire w_dff_B_a60FCBK10_2;
	wire w_dff_B_s1t0Ne6l1_2;
	wire w_dff_B_8txMS7B40_2;
	wire w_dff_B_DX4hwEel0_2;
	wire w_dff_B_UALV2Nvv2_2;
	wire w_dff_B_rbZtHZzC4_2;
	wire w_dff_B_Mckbp9AA5_2;
	wire w_dff_B_LqIoFn6Q8_2;
	wire w_dff_B_f3VAqxAh7_2;
	wire w_dff_B_CnYgRNZE5_2;
	wire w_dff_B_pVWbBQ752_2;
	wire w_dff_B_lQkJtgS43_2;
	wire w_dff_B_OoVrgO5r5_2;
	wire w_dff_B_01azvw9k8_2;
	wire w_dff_B_vvHpNv2c6_2;
	wire w_dff_B_0Nxn7GMb3_2;
	wire w_dff_B_oJBPUXTm8_2;
	wire w_dff_B_jtkDR4jN2_2;
	wire w_dff_B_0QZrmuTs4_2;
	wire w_dff_B_4ONyxXPC6_2;
	wire w_dff_B_9DXOjNco4_2;
	wire w_dff_B_plsApLue3_2;
	wire w_dff_B_iZ8OwxC19_2;
	wire w_dff_B_P7ODU0VS2_2;
	wire w_dff_B_7XkJH0Kl6_2;
	wire w_dff_B_J2CyJSVW3_2;
	wire w_dff_B_awG32zrH7_2;
	wire w_dff_B_G4phLsEV1_2;
	wire w_dff_B_1sSPCddY0_2;
	wire w_dff_B_1KItqeoN9_2;
	wire w_dff_B_bjkQGqVN7_2;
	wire w_dff_B_GnKywHke3_2;
	wire w_dff_B_hcg06UVb7_2;
	wire w_dff_B_KMgVGQSX8_2;
	wire w_dff_B_m8TLvjHr8_2;
	wire w_dff_B_lBGh094G6_2;
	wire w_dff_B_A9W44fyG5_2;
	wire w_dff_B_ITUO9W679_2;
	wire w_dff_B_jubSsqcg2_2;
	wire w_dff_B_ftAC1Tv30_2;
	wire w_dff_B_lQcMoh2d5_2;
	wire w_dff_B_RzhjSOY79_2;
	wire w_dff_B_IVtF71gj1_2;
	wire w_dff_B_ne5l9KOw5_2;
	wire w_dff_B_LZv7m9H48_2;
	wire w_dff_B_xLPZGdPs7_2;
	wire w_dff_B_WpcYmYiE8_2;
	wire w_dff_B_Xe29gkP29_2;
	wire w_dff_B_X8q39fkN9_2;
	wire w_dff_B_qEs4RS6u6_2;
	wire w_dff_B_wu1PItlE7_2;
	wire w_dff_B_b7iuyeou2_2;
	wire w_dff_B_VMXC3PbE2_2;
	wire w_dff_B_mHuU6GOr7_2;
	wire w_dff_B_7fl2GvwK8_2;
	wire w_dff_B_4YiJLsiw6_2;
	wire w_dff_B_eP5FJVGW1_2;
	wire w_dff_B_d4gPjic42_2;
	wire w_dff_B_JOLA9J4w9_2;
	wire w_dff_B_c2lYvNJ78_2;
	wire w_dff_B_hODBv9zx5_2;
	wire w_dff_B_zNY6mDat2_2;
	wire w_dff_B_x8AeANCb1_2;
	wire w_dff_B_gqMnlbSj4_2;
	wire w_dff_B_QR4AWM4t6_2;
	wire w_dff_B_eoTPu0120_2;
	wire w_dff_B_KRrr06ro0_2;
	wire w_dff_B_yPDbsUSp2_2;
	wire w_dff_B_4D4VzV5M7_2;
	wire w_dff_B_iAMWRmag3_2;
	wire w_dff_B_i7GRGFgO4_2;
	wire w_dff_B_QEukstIO4_2;
	wire w_dff_B_Q5QgZt8i7_2;
	wire w_dff_B_89Bz2bgh5_2;
	wire w_dff_B_X7fyyJgm1_2;
	wire w_dff_B_pvEecekj9_2;
	wire w_dff_B_epgzQZn99_2;
	wire w_dff_B_WbEVTkPs8_2;
	wire w_dff_B_QDa8gHla1_2;
	wire w_dff_B_mEwxybiH7_2;
	wire w_dff_B_7lJ4oeRx8_2;
	wire w_dff_B_kv4gH2Zd2_2;
	wire w_dff_B_hrir7I2z8_2;
	wire w_dff_B_LD9XSOiS3_1;
	wire w_dff_B_IO8osC6D0_2;
	wire w_dff_B_5YZ5C6Kq6_2;
	wire w_dff_B_mt6k1Qos2_2;
	wire w_dff_B_jtmtyrZ36_2;
	wire w_dff_B_M5YPqomP5_2;
	wire w_dff_B_HgGLTEMa7_2;
	wire w_dff_B_2QcuSjtX7_2;
	wire w_dff_B_wmwHp6Js4_2;
	wire w_dff_B_zzYyRr8p3_2;
	wire w_dff_B_VO1JxMWh7_2;
	wire w_dff_B_AqsmNwUX4_2;
	wire w_dff_B_B9KIpRH98_2;
	wire w_dff_B_V2zO15AL1_2;
	wire w_dff_B_WGas6kLb8_2;
	wire w_dff_B_dxtI1b3L5_2;
	wire w_dff_B_BNkXoz4z2_2;
	wire w_dff_B_p6AAIeBf7_2;
	wire w_dff_B_loF9KRgF4_2;
	wire w_dff_B_55OKPuuj6_2;
	wire w_dff_B_D5tdWEfJ1_2;
	wire w_dff_B_uT3CuPGq1_2;
	wire w_dff_B_2YkQPLcm9_2;
	wire w_dff_B_7Ie72Y0Y4_2;
	wire w_dff_B_LQYwPaLL0_2;
	wire w_dff_B_LuE6FoXo9_2;
	wire w_dff_B_VeGAicis8_2;
	wire w_dff_B_OAZR1hcB0_2;
	wire w_dff_B_z6tL5lTR1_2;
	wire w_dff_B_3SOP35U57_2;
	wire w_dff_B_4ldaTvvg9_2;
	wire w_dff_B_E4V7pNm14_2;
	wire w_dff_B_GjkRbhM33_2;
	wire w_dff_B_8RUqxONn7_2;
	wire w_dff_B_rjemjsH95_2;
	wire w_dff_B_pXfP7u089_2;
	wire w_dff_B_6fugebGy4_2;
	wire w_dff_B_SuRv9RT48_2;
	wire w_dff_B_grxZZwjR0_2;
	wire w_dff_B_FH7jW32D5_2;
	wire w_dff_B_11h2mnBb6_1;
	wire w_dff_B_QnrhvDJ39_1;
	wire w_dff_B_OjtRWkz85_2;
	wire w_dff_B_H4sLWXAM1_2;
	wire w_dff_B_rhKgKYmg2_2;
	wire w_dff_B_PrcewLJg3_2;
	wire w_dff_B_ciMQANda1_2;
	wire w_dff_B_BsoIaXf27_2;
	wire w_dff_B_oQWgyVv40_2;
	wire w_dff_B_yB01E5nB4_2;
	wire w_dff_B_7FeFVmGh3_2;
	wire w_dff_B_Tmxh3YeH3_2;
	wire w_dff_B_yCsTGjWz8_2;
	wire w_dff_B_y9zwp4Az5_2;
	wire w_dff_B_YFiH6sbf2_2;
	wire w_dff_B_FnzaljUV9_2;
	wire w_dff_B_ix1L4zjC8_2;
	wire w_dff_B_VVQpPhB32_2;
	wire w_dff_B_sSgwnOrU2_2;
	wire w_dff_B_UJZ3Wht43_2;
	wire w_dff_B_S6OOM1Kq2_2;
	wire w_dff_B_dBV8XEuL1_2;
	wire w_dff_B_sxWOfH029_2;
	wire w_dff_B_uwtfZuaL3_2;
	wire w_dff_B_PRHyGlfj1_2;
	wire w_dff_B_NwBrKywE1_2;
	wire w_dff_B_mI0wTFno9_2;
	wire w_dff_B_hX6AAV445_2;
	wire w_dff_B_5CvxOZxv5_2;
	wire w_dff_B_7c00OjEb2_2;
	wire w_dff_B_MbRKR5KN5_2;
	wire w_dff_B_BkYHmE6V4_2;
	wire w_dff_B_YE2rx8cE6_2;
	wire w_dff_B_Q2Bm8MuR8_2;
	wire w_dff_B_5MqNYOMH4_2;
	wire w_dff_B_lnxo9GcD3_2;
	wire w_dff_B_dOovRSgX9_2;
	wire w_dff_B_gllUR0MF3_2;
	wire w_dff_B_XnR8pnxw7_2;
	wire w_dff_B_GR15E4pp6_2;
	wire w_dff_B_PCIhFuYQ6_2;
	wire w_dff_B_IKYZ6lqQ6_2;
	wire w_dff_B_E65ue60G1_2;
	wire w_dff_B_CuRHdUgE3_2;
	wire w_dff_B_vf1kuXxr8_2;
	wire w_dff_B_jnb87pNR1_2;
	wire w_dff_B_8X9VvcrN1_2;
	wire w_dff_B_nrCLN1p26_2;
	wire w_dff_B_yog6ln8E5_2;
	wire w_dff_B_pEmW8hLs0_2;
	wire w_dff_B_TkCdXKA67_2;
	wire w_dff_B_FW6cNoW11_2;
	wire w_dff_B_ehuOBwyZ0_2;
	wire w_dff_B_0ZrObZ2m1_2;
	wire w_dff_B_Eq7tGFbb8_2;
	wire w_dff_B_10mGnbdy4_2;
	wire w_dff_B_cJiyqwCu8_2;
	wire w_dff_B_CVoOe6WP7_2;
	wire w_dff_B_868FyOFP4_2;
	wire w_dff_B_Q08SRK5p4_2;
	wire w_dff_B_alGe5RtK7_2;
	wire w_dff_B_Zp6xdwHW2_2;
	wire w_dff_B_I8DUJgua2_2;
	wire w_dff_B_31Sj8Rt25_2;
	wire w_dff_B_JV0yl0MZ1_2;
	wire w_dff_B_j9x3Q7nm3_2;
	wire w_dff_B_GnXLaZHG8_2;
	wire w_dff_B_Z3pLEOEH0_2;
	wire w_dff_B_HbzwnA556_2;
	wire w_dff_B_dv1s7Ykx1_2;
	wire w_dff_B_ObRThRGk1_2;
	wire w_dff_B_XwJ5JWuj3_2;
	wire w_dff_B_2q4SW0fe1_2;
	wire w_dff_B_ocKxbxSA6_2;
	wire w_dff_B_9PAd5v7J8_2;
	wire w_dff_B_NufzxXYp2_2;
	wire w_dff_B_IGBSwx534_2;
	wire w_dff_B_PRIZboWh1_1;
	wire w_dff_B_NracL9LR4_2;
	wire w_dff_B_0NUeyTxa8_2;
	wire w_dff_B_zRK2UE0c0_2;
	wire w_dff_B_FN3IRPQl4_2;
	wire w_dff_B_jAv1NIka7_2;
	wire w_dff_B_teeeHzWr1_2;
	wire w_dff_B_6fvY58Yc2_2;
	wire w_dff_B_Qwudmptu0_2;
	wire w_dff_B_MCD9BKO21_2;
	wire w_dff_B_dgyQrOCl3_2;
	wire w_dff_B_caS2ihKx8_2;
	wire w_dff_B_sERGt8je2_2;
	wire w_dff_B_wse96MkP4_2;
	wire w_dff_B_YVoBk29T8_2;
	wire w_dff_B_rNnEPmTd7_2;
	wire w_dff_B_91DkQBZA9_2;
	wire w_dff_B_WzkmCQyW8_2;
	wire w_dff_B_2Mjyl81S8_2;
	wire w_dff_B_RQRhDMSc3_2;
	wire w_dff_B_xLWUme7f7_2;
	wire w_dff_B_M4pE5sV05_2;
	wire w_dff_B_FiRVVw5h1_2;
	wire w_dff_B_4mzbmJPp6_2;
	wire w_dff_B_AOlAwuXk7_2;
	wire w_dff_B_BTHarfsS1_2;
	wire w_dff_B_4UvEFnxN4_2;
	wire w_dff_B_TbSFipsC5_2;
	wire w_dff_B_qCxYuplw6_2;
	wire w_dff_B_02PCvWrG3_2;
	wire w_dff_B_TwB6wEks6_2;
	wire w_dff_B_FDz5upXD3_2;
	wire w_dff_B_SiabVybH4_2;
	wire w_dff_B_VraM9NXu3_2;
	wire w_dff_B_qJzGZ17T5_2;
	wire w_dff_B_poyiy4tx3_2;
	wire w_dff_B_o269yUIt0_1;
	wire w_dff_B_F8seNExg6_1;
	wire w_dff_B_CKhLp4CL1_2;
	wire w_dff_B_xRDHZbVN6_2;
	wire w_dff_B_oqi26wSG4_2;
	wire w_dff_B_9tYi3ZoF6_2;
	wire w_dff_B_wZVMEj6s0_2;
	wire w_dff_B_tJibNlXw0_2;
	wire w_dff_B_JbuW4FVZ4_2;
	wire w_dff_B_JMyUr2pa2_2;
	wire w_dff_B_spw74YZt9_2;
	wire w_dff_B_68BhCiDL5_2;
	wire w_dff_B_9pAHtDJY3_2;
	wire w_dff_B_tD8IOVpw4_2;
	wire w_dff_B_lFHHKp1E1_2;
	wire w_dff_B_sYNlZP2V8_2;
	wire w_dff_B_6fJPR5jL1_2;
	wire w_dff_B_Z1351Jwl1_2;
	wire w_dff_B_NAhqd4hB7_2;
	wire w_dff_B_uftwVYDF0_2;
	wire w_dff_B_YTM6FdhP4_2;
	wire w_dff_B_XT5l0IX35_2;
	wire w_dff_B_gfi2GPms9_2;
	wire w_dff_B_7LGXwjJU3_2;
	wire w_dff_B_9Bl4KFyY8_2;
	wire w_dff_B_P7fVqXY20_2;
	wire w_dff_B_bcNGexlG7_2;
	wire w_dff_B_qkyEtRzg8_2;
	wire w_dff_B_5zXY9Bby4_2;
	wire w_dff_B_I9nvUdiI9_2;
	wire w_dff_B_Wzt3jgkN5_2;
	wire w_dff_B_qa9CpgJ81_2;
	wire w_dff_B_4MP7TjJv7_2;
	wire w_dff_B_k33KKcJH0_2;
	wire w_dff_B_z5sIHDtl4_2;
	wire w_dff_B_ceOKQeDm3_2;
	wire w_dff_B_OIwOBmQ74_2;
	wire w_dff_B_3VDPHyRE7_2;
	wire w_dff_B_45xF50ic2_2;
	wire w_dff_B_OkN2jMdi2_2;
	wire w_dff_B_oH16Peh98_2;
	wire w_dff_B_LR98fBSb3_2;
	wire w_dff_B_m2VBFUQB9_2;
	wire w_dff_B_ofV171bt6_2;
	wire w_dff_B_y2q5XDX69_2;
	wire w_dff_B_XP0fBp7V2_2;
	wire w_dff_B_W8vqF5TY8_2;
	wire w_dff_B_ieeJvNcR6_2;
	wire w_dff_B_qfeuUqiQ7_2;
	wire w_dff_B_rCIUZCPg8_2;
	wire w_dff_B_RJ14PlcM2_2;
	wire w_dff_B_3ZsxmYPr5_2;
	wire w_dff_B_M8SpTF1E4_2;
	wire w_dff_B_cXHeC0i30_2;
	wire w_dff_B_3pZV89Ul7_2;
	wire w_dff_B_vKJCAfLp4_2;
	wire w_dff_B_YlPJwVTa2_2;
	wire w_dff_B_Ag52ToH48_2;
	wire w_dff_B_In1xradN7_2;
	wire w_dff_B_Ssv5yBim0_2;
	wire w_dff_B_eW05ITvY5_2;
	wire w_dff_B_VOxdsDCI2_2;
	wire w_dff_B_u4nTYRW40_2;
	wire w_dff_B_3WN5ZGwT8_2;
	wire w_dff_B_qENnCH9B0_2;
	wire w_dff_B_KU1oYdmK9_2;
	wire w_dff_B_PCSE2ZYu5_2;
	wire w_dff_B_Dk0tMq5b9_2;
	wire w_dff_B_896xBcra0_2;
	wire w_dff_B_McwKnVtr5_1;
	wire w_dff_B_bZ6WEBNu7_2;
	wire w_dff_B_xzEVptqB3_2;
	wire w_dff_B_ea4bv41s1_2;
	wire w_dff_B_EEK7yyOR7_2;
	wire w_dff_B_G5rB0ymr7_2;
	wire w_dff_B_GLf2xhsH2_2;
	wire w_dff_B_dXmZjGWX2_2;
	wire w_dff_B_3muGzQyA3_2;
	wire w_dff_B_2FDjoapF1_2;
	wire w_dff_B_KEI8AuKV3_2;
	wire w_dff_B_VDBAvZfu0_2;
	wire w_dff_B_NgLvRoqM9_2;
	wire w_dff_B_2ab4lZzW5_2;
	wire w_dff_B_BrQETskv6_2;
	wire w_dff_B_7Y5AYlhf9_2;
	wire w_dff_B_ewG0hSRH3_2;
	wire w_dff_B_WPS5zvIH6_2;
	wire w_dff_B_CBfMUNlC8_2;
	wire w_dff_B_Q7SK2WP14_2;
	wire w_dff_B_9RdwN7NJ2_2;
	wire w_dff_B_utU1DPPF8_2;
	wire w_dff_B_dCgsYsmP2_2;
	wire w_dff_B_MD0JMfIu9_2;
	wire w_dff_B_gBZwyyzt0_2;
	wire w_dff_B_AhXiICfe0_2;
	wire w_dff_B_v8yKt9CW2_2;
	wire w_dff_B_lMxW56rO1_2;
	wire w_dff_B_M4PoGaBP3_2;
	wire w_dff_B_XT0Pvyyn6_2;
	wire w_dff_B_ZOu315Ty6_2;
	wire w_dff_B_ugBGSNfa3_2;
	wire w_dff_B_qoDRJVxL7_1;
	wire w_dff_B_2ezTw40N3_1;
	wire w_dff_B_58UfveQP3_2;
	wire w_dff_B_ADp3j63K0_2;
	wire w_dff_B_i7itV8O29_2;
	wire w_dff_B_UAApKXy27_2;
	wire w_dff_B_ualVowA88_2;
	wire w_dff_B_QcDY9brj0_2;
	wire w_dff_B_GdyBCVIk3_2;
	wire w_dff_B_TiogwJfi9_2;
	wire w_dff_B_gPw2qPn51_2;
	wire w_dff_B_3lSYcOmN9_2;
	wire w_dff_B_RqrDtsIH9_2;
	wire w_dff_B_nqltyu9W7_2;
	wire w_dff_B_Llt5KdTM8_2;
	wire w_dff_B_Cbi5UaaD9_2;
	wire w_dff_B_Y1QeJM9E6_2;
	wire w_dff_B_dPpWhZ6g2_2;
	wire w_dff_B_qwjEigGV2_2;
	wire w_dff_B_8rUETevF1_2;
	wire w_dff_B_igXJoIem2_2;
	wire w_dff_B_uZnQPvYp7_2;
	wire w_dff_B_y8rwqxq31_2;
	wire w_dff_B_FKTrVXhZ8_2;
	wire w_dff_B_3nv21eCL6_2;
	wire w_dff_B_F19CCd8T2_2;
	wire w_dff_B_kFLHSc7L3_2;
	wire w_dff_B_VeEQDDQO3_2;
	wire w_dff_B_vzwqLw0d9_2;
	wire w_dff_B_7nodYucn0_2;
	wire w_dff_B_60a6Xq1l9_2;
	wire w_dff_B_hodZAB5S2_2;
	wire w_dff_B_KXkbuGap5_2;
	wire w_dff_B_q24DgdNX2_2;
	wire w_dff_B_lI9Asubr5_2;
	wire w_dff_B_C9nG3yxR4_2;
	wire w_dff_B_YcRguUlg1_2;
	wire w_dff_B_3vZBWnPc9_2;
	wire w_dff_B_pbwmV0Pd3_2;
	wire w_dff_B_N8ZhIHqc4_2;
	wire w_dff_B_f70K9my72_2;
	wire w_dff_B_irg1wuLv2_2;
	wire w_dff_B_z4IAjJXj2_2;
	wire w_dff_B_cbLsPkEf9_2;
	wire w_dff_B_BRob48bd0_2;
	wire w_dff_B_9uiwO0Nl7_2;
	wire w_dff_B_SLiuM5ML4_2;
	wire w_dff_B_KYcwbfYM0_2;
	wire w_dff_B_zRRdla247_2;
	wire w_dff_B_VYh0AFar9_2;
	wire w_dff_B_BvHwI7er9_2;
	wire w_dff_B_SSqH70Pr3_2;
	wire w_dff_B_s0avIIv43_2;
	wire w_dff_B_e6Yqgxd20_2;
	wire w_dff_B_C41PjQDs7_2;
	wire w_dff_B_voCVrfKC1_2;
	wire w_dff_B_Kf2JBVjW1_2;
	wire w_dff_B_oFa4G7VG1_2;
	wire w_dff_B_3CPhrYIH7_2;
	wire w_dff_B_8YzArT0w9_2;
	wire w_dff_B_jyCedYn23_2;
	wire w_dff_B_4ZGyLYI34_1;
	wire w_dff_B_qFNYwrEz8_2;
	wire w_dff_B_aPMWol1E1_2;
	wire w_dff_B_YHzQ0G6b9_2;
	wire w_dff_B_7x82HizO4_2;
	wire w_dff_B_trzPZ1DV9_2;
	wire w_dff_B_iTpLJomj2_2;
	wire w_dff_B_Noac6bpN9_2;
	wire w_dff_B_ziRsvjyZ2_2;
	wire w_dff_B_tY7iefEe6_2;
	wire w_dff_B_sTQAvUcs4_2;
	wire w_dff_B_mXctcUt55_2;
	wire w_dff_B_29Y4etSI2_2;
	wire w_dff_B_WuFtF8pK6_2;
	wire w_dff_B_zO4t1JEV1_2;
	wire w_dff_B_Hb4tDzjv1_2;
	wire w_dff_B_mnmD1hQL7_2;
	wire w_dff_B_mMfPWLG28_2;
	wire w_dff_B_F3GEOyI63_2;
	wire w_dff_B_QeSoVTIQ9_2;
	wire w_dff_B_PXKRWx8c6_2;
	wire w_dff_B_ofihC0d07_2;
	wire w_dff_B_c656eRfT1_2;
	wire w_dff_B_lOISoo5H7_2;
	wire w_dff_B_rPZS3WR15_2;
	wire w_dff_B_t3HreJNU1_2;
	wire w_dff_B_gN63ag3Z0_2;
	wire w_dff_B_FDLZUWT77_2;
	wire w_dff_B_VA2S6U9k3_1;
	wire w_dff_B_RSFFa2ch4_1;
	wire w_dff_B_qYTGGBHQ4_2;
	wire w_dff_B_DnQe1eps2_2;
	wire w_dff_B_wOc0NqTM3_2;
	wire w_dff_B_l2LCdCB09_2;
	wire w_dff_B_fMjO1sZz7_2;
	wire w_dff_B_D2krJ9sU8_2;
	wire w_dff_B_V3Tvob7D8_2;
	wire w_dff_B_aoBNOexl5_2;
	wire w_dff_B_Igy2xp7q7_2;
	wire w_dff_B_fPLs186h5_2;
	wire w_dff_B_ooSGm1Wu3_2;
	wire w_dff_B_EPIkemYa6_2;
	wire w_dff_B_0srqfk369_2;
	wire w_dff_B_mDjfZofs0_2;
	wire w_dff_B_ONRmRIjR0_2;
	wire w_dff_B_Fn0cynub1_2;
	wire w_dff_B_Cy1ke8qC5_2;
	wire w_dff_B_l3P9r0Z05_2;
	wire w_dff_B_tn8Bj7vT3_2;
	wire w_dff_B_ZZfgxB8n9_2;
	wire w_dff_B_inr8OxK96_2;
	wire w_dff_B_zqSBWBxZ4_2;
	wire w_dff_B_XdgUDHoV7_2;
	wire w_dff_B_qLO6wcXk4_2;
	wire w_dff_B_2GUUuvJi6_2;
	wire w_dff_B_BcUnDo3x0_2;
	wire w_dff_B_ZTUmweih7_2;
	wire w_dff_B_mnxWbeaS7_2;
	wire w_dff_B_mly1ZQ6m9_2;
	wire w_dff_B_DsxJIYWN8_2;
	wire w_dff_B_cSN5Cmro0_2;
	wire w_dff_B_CBPklAv78_2;
	wire w_dff_B_eYqCWvtK9_2;
	wire w_dff_B_JzIh3nX11_2;
	wire w_dff_B_R1tHNeA23_2;
	wire w_dff_B_y3sOlxXo1_2;
	wire w_dff_B_FQuTkHes5_2;
	wire w_dff_B_hF9g4pqb5_2;
	wire w_dff_B_hYx4OPiE9_2;
	wire w_dff_B_wqBGXGS29_2;
	wire w_dff_B_EVUWCY8u1_2;
	wire w_dff_B_AVD8uGbv5_2;
	wire w_dff_B_LZAS6Ncv7_2;
	wire w_dff_B_9Ezn80wH8_2;
	wire w_dff_B_drNNHBSY3_2;
	wire w_dff_B_40GxfDLh2_2;
	wire w_dff_B_hkNq5KuS4_2;
	wire w_dff_B_0jv3VXap9_2;
	wire w_dff_B_cx3cJiul8_2;
	wire w_dff_B_9HjdEJhl7_2;
	wire w_dff_B_jUVca4ae9_2;
	wire w_dff_B_QnmaqLHI3_1;
	wire w_dff_B_RTYpZfbk8_2;
	wire w_dff_B_1h5JXzJ86_2;
	wire w_dff_B_AcHC6nNx6_2;
	wire w_dff_B_ocXo9ELj4_2;
	wire w_dff_B_jKH6hJgT0_2;
	wire w_dff_B_ilvAowbK1_2;
	wire w_dff_B_VLPeSxyM5_2;
	wire w_dff_B_XU5Xcd4s4_2;
	wire w_dff_B_B89o1cIh6_2;
	wire w_dff_B_msrWJA2I1_2;
	wire w_dff_B_EzqXSzlB0_2;
	wire w_dff_B_GSA0RLq28_2;
	wire w_dff_B_yF99YuQj5_2;
	wire w_dff_B_myVQmF2v8_2;
	wire w_dff_B_H9CCqDaM9_2;
	wire w_dff_B_CITYv9zH7_2;
	wire w_dff_B_IqlDVPEu7_2;
	wire w_dff_B_k5spDBxP4_2;
	wire w_dff_B_hGmShCwr1_2;
	wire w_dff_B_9OR9JLkl7_2;
	wire w_dff_B_kehTNLxI5_2;
	wire w_dff_B_XzFRErpm5_2;
	wire w_dff_B_XOoBHcnR4_2;
	wire w_dff_B_5yASU09a7_1;
	wire w_dff_B_OLZWrOjp4_1;
	wire w_dff_B_olLFN9c87_2;
	wire w_dff_B_Oy1yACP37_2;
	wire w_dff_B_hILtbE4e4_2;
	wire w_dff_B_jAZ0UAPM5_2;
	wire w_dff_B_tD6kzMRP0_2;
	wire w_dff_B_9EfIgV226_2;
	wire w_dff_B_2sTwPaFB7_2;
	wire w_dff_B_LGlJ9LGR6_2;
	wire w_dff_B_Gy1z6sy28_2;
	wire w_dff_B_qil5CCJE2_2;
	wire w_dff_B_ugPp0WhU1_2;
	wire w_dff_B_fqUOMK534_2;
	wire w_dff_B_mhWh2Hty5_2;
	wire w_dff_B_v5OiShYa0_2;
	wire w_dff_B_wVN5XThm4_2;
	wire w_dff_B_XR9ue4V19_2;
	wire w_dff_B_bKVQjgk65_2;
	wire w_dff_B_P6lI9vI11_2;
	wire w_dff_B_zQGYo7ns2_2;
	wire w_dff_B_2TsNxkrJ7_2;
	wire w_dff_B_u4OSFqmP6_2;
	wire w_dff_B_nlfaaTG72_2;
	wire w_dff_B_VJVzxNCg7_2;
	wire w_dff_B_30SkPjq55_2;
	wire w_dff_B_uSQi8yFR7_2;
	wire w_dff_B_3Ahs3CHu0_2;
	wire w_dff_B_1jT8OPdh5_2;
	wire w_dff_B_5JuWZToz2_2;
	wire w_dff_B_VtPQUMxf3_2;
	wire w_dff_B_YH45DRSu7_2;
	wire w_dff_B_4APZnBpN8_2;
	wire w_dff_B_c0tyCitH7_2;
	wire w_dff_B_b4kjQ4vj9_2;
	wire w_dff_B_GtTC14yz3_2;
	wire w_dff_B_J9YPhhVi8_2;
	wire w_dff_B_ce6ZBtkp1_2;
	wire w_dff_B_EagJwI7z3_2;
	wire w_dff_B_x5wcMjqP2_2;
	wire w_dff_B_dz69GAil1_2;
	wire w_dff_B_USR9CEH27_2;
	wire w_dff_B_IVvOEBOt9_2;
	wire w_dff_B_IEOErc0A7_2;
	wire w_dff_B_fYYk5f3O9_2;
	wire w_dff_B_8PWg07E36_1;
	wire w_dff_B_OzHhAVOr8_2;
	wire w_dff_B_VKHez9Q05_2;
	wire w_dff_B_wSxZEkEG6_2;
	wire w_dff_B_bgpXZGrs1_2;
	wire w_dff_B_TQyk5DZu4_2;
	wire w_dff_B_iiZ26NXU0_2;
	wire w_dff_B_u3ZcPFKs5_2;
	wire w_dff_B_NH2bHgDY3_2;
	wire w_dff_B_KOPAkTZ98_2;
	wire w_dff_B_GJyHhEcH6_2;
	wire w_dff_B_H7y5d9bZ3_2;
	wire w_dff_B_tslGbXB79_2;
	wire w_dff_B_N1htLnBN3_2;
	wire w_dff_B_w00JVhEH6_2;
	wire w_dff_B_oZbSLAm03_2;
	wire w_dff_B_GFeb4tGH0_2;
	wire w_dff_B_2V2Ugc569_2;
	wire w_dff_B_VOrXH5oj5_2;
	wire w_dff_B_EGF4byLT4_2;
	wire w_dff_B_Qv0e2HCL2_1;
	wire w_dff_B_e2ET3Y1E7_1;
	wire w_dff_B_Y3Dj646E0_2;
	wire w_dff_B_7CvXI7ia0_2;
	wire w_dff_B_9xXQQOur9_2;
	wire w_dff_B_7HO27aZ45_2;
	wire w_dff_B_jJNuFAOp9_2;
	wire w_dff_B_cYqN30bH0_2;
	wire w_dff_B_DlhQfQlF8_2;
	wire w_dff_B_exE0wN6I5_2;
	wire w_dff_B_vuCazIXF0_2;
	wire w_dff_B_BKjuYlam2_2;
	wire w_dff_B_wD24toJc9_2;
	wire w_dff_B_MQpUhRpQ3_2;
	wire w_dff_B_ziTNQ1Cx2_2;
	wire w_dff_B_RkkV6wiZ3_2;
	wire w_dff_B_AxdOm1kF0_2;
	wire w_dff_B_7a6jpQSa0_2;
	wire w_dff_B_LFO4qeg28_2;
	wire w_dff_B_Mw2zSURz3_2;
	wire w_dff_B_BlHRHpQm6_2;
	wire w_dff_B_g23d2ye54_2;
	wire w_dff_B_HslQ4LMC2_2;
	wire w_dff_B_qFEL7Ce34_2;
	wire w_dff_B_NfJh0SOk3_2;
	wire w_dff_B_0kdqCHKs6_2;
	wire w_dff_B_RCXf0GSK9_2;
	wire w_dff_B_SbeIj4EA9_2;
	wire w_dff_B_oWCisUL88_2;
	wire w_dff_B_73KwR9kl1_2;
	wire w_dff_B_Ws0GHVFN2_2;
	wire w_dff_B_MSt4HiVG0_2;
	wire w_dff_B_yZAGZScQ3_2;
	wire w_dff_B_pM6Mmx3n7_2;
	wire w_dff_B_IjKhdoj22_2;
	wire w_dff_B_HNwucoHX8_2;
	wire w_dff_B_MWaXlhv09_2;
	wire w_dff_B_DZrKGAMs6_1;
	wire w_dff_B_szCQqSSU2_2;
	wire w_dff_B_lOEFlTU39_2;
	wire w_dff_B_Jqv4AdE23_2;
	wire w_dff_B_XiAMtTEU2_2;
	wire w_dff_B_cbUdpB1v5_2;
	wire w_dff_B_EZjbtMY64_2;
	wire w_dff_B_kCVwGTK17_2;
	wire w_dff_B_IM5IdGkX5_2;
	wire w_dff_B_EWB7lJfj3_2;
	wire w_dff_B_y4KSNL9q6_2;
	wire w_dff_B_BruesTkW2_2;
	wire w_dff_B_pgFTnIOK6_2;
	wire w_dff_B_xVlEOmrX7_2;
	wire w_dff_B_6J2NyFim8_2;
	wire w_dff_B_B9IrkPD37_2;
	wire w_dff_B_RntvHVY90_2;
	wire w_dff_B_fG3DPFL78_2;
	wire w_dff_B_utpFtmHA2_2;
	wire w_dff_B_NT2Q9DQR8_2;
	wire w_dff_B_0q3OCYoI2_2;
	wire w_dff_B_v2k9uez14_2;
	wire w_dff_B_5AdnHcnK5_2;
	wire w_dff_B_QqvYuJ5h8_2;
	wire w_dff_B_T2Q7Wbqm2_2;
	wire w_dff_B_mES2Qmt23_2;
	wire w_dff_B_fxYnfF0S9_2;
	wire w_dff_B_RqiMIXOz0_2;
	wire w_dff_B_wTSyRGBe8_2;
	wire w_dff_B_R7U1seq15_2;
	wire w_dff_B_Cnh3ALpc1_2;
	wire w_dff_B_wAlqMFZK2_2;
	wire w_dff_B_YmJ0rA5v8_2;
	wire w_dff_B_EqXigxnl2_2;
	wire w_dff_B_qEd7GUfv1_2;
	wire w_dff_B_USPE4sBL7_2;
	wire w_dff_B_9s7J8j272_2;
	wire w_dff_B_MW0mOvnW2_2;
	wire w_dff_B_uHG8XFyv3_2;
	wire w_dff_B_VSTZy9ar0_2;
	wire w_dff_B_5pvmsgAx2_2;
	wire w_dff_B_y5rNK1No5_2;
	wire w_dff_B_ZnJx9fZ55_2;
	wire w_dff_B_ekLgpStc5_1;
	wire w_dff_B_bStYKeD78_2;
	wire w_dff_B_tcQEwGcI6_2;
	wire w_dff_B_HzGCXw0e3_2;
	wire w_dff_B_o0zYhiyG4_2;
	wire w_dff_B_TI8ZuKjZ5_2;
	wire w_dff_B_TpDxDOgf3_2;
	wire w_dff_B_gXurmGlr9_2;
	wire w_dff_B_7IOOwjVc4_2;
	wire w_dff_B_R5OmwPa20_2;
	wire w_dff_B_lIu6VCdA5_2;
	wire w_dff_B_9lWhhvuT2_2;
	wire w_dff_A_Ajg6pi0s7_0;
	wire w_dff_A_AKZFsUKo0_0;
	wire w_dff_A_f2e2Ey2h5_0;
	wire w_dff_B_GDoq4Fl55_2;
	wire w_dff_B_35JBD6cT9_1;
	wire w_dff_B_mznpII4E5_1;
	wire w_dff_B_vwTQ4LEh0_1;
	wire w_dff_B_tLoMFTzR5_1;
	wire w_dff_B_pfb2HwpJ1_1;
	wire w_dff_B_B5JNyJST3_1;
	wire w_dff_B_PQHk8nW76_1;
	wire w_dff_B_IWVdypPc3_1;
	wire w_dff_A_TZ6tGNyO8_1;
	wire w_dff_A_4xiO9KTf8_1;
	wire w_dff_A_m2JdDYnS7_1;
	wire w_dff_A_XdPmzeat0_1;
	wire w_dff_A_vhJuOkKT5_1;
	wire w_dff_A_xXmrnfsi0_1;
	wire w_dff_A_TGokZRHD9_1;
	wire w_dff_B_RmMAyjat2_2;
	wire w_dff_B_39TboRSy1_2;
	wire w_dff_B_Ch6Yixrm2_2;
	wire w_dff_B_gZ8hmKrM8_2;
	wire w_dff_B_YNY4Uvzw2_2;
	wire w_dff_B_1yeDeOyg8_2;
	wire w_dff_B_dq8Y05WN7_2;
	wire w_dff_B_UC6AoPgJ6_2;
	wire w_dff_B_pKyIMzVa8_2;
	wire w_dff_B_cqFfBWP55_2;
	wire w_dff_B_cmfpmCl56_1;
	wire w_dff_B_X1hBfCeL4_2;
	wire w_dff_B_UfPsd2bc2_2;
	wire w_dff_B_yV00sn1Q7_2;
	wire w_dff_B_y9DjVUcg0_2;
	wire w_dff_B_jWFSNWq73_2;
	wire w_dff_B_JD0A8qP97_2;
	wire w_dff_B_snnwlZP56_2;
	wire w_dff_B_rvbvWtr08_2;
	wire w_dff_B_aMxbGL8a2_2;
	wire w_dff_B_WbleH03o3_2;
	wire w_dff_B_m1RCkkPH9_2;
	wire w_dff_B_Wp4tjeBe1_2;
	wire w_dff_B_rbubUt2i7_2;
	wire w_dff_A_U1HcrelJ0_0;
	wire w_dff_A_2ggyHQ8U6_0;
	wire w_dff_A_vaNofmMD7_0;
	wire w_dff_A_uVjBeraU8_0;
	wire w_dff_A_B5pqTIi46_1;
	wire w_dff_A_DIA0lUDf8_1;
	wire w_dff_B_5oDqQnFC4_1;
	wire w_dff_B_KZLhzZXj0_1;
	wire w_dff_B_YmpiVlK80_1;
	wire w_dff_B_bvM5pOaO1_1;
	wire w_dff_B_7ocKJlph9_1;
	wire w_dff_A_3tzYqdid4_0;
	wire w_dff_A_iPbA4AM20_0;
	wire w_dff_A_uLByc2El7_0;
	wire w_dff_A_f2OUeufa5_0;
	wire w_dff_A_0kBr7MwZ8_0;
	wire w_dff_A_VCHMQp1s7_0;
	wire w_dff_B_lLac3uo07_2;
	wire w_dff_A_HlqjyqD42_1;
	wire w_dff_A_z9GPjSto8_1;
	wire w_dff_A_PqR25d2d6_1;
	wire w_dff_A_LFZNbteQ8_1;
	wire w_dff_A_AhwbHvEf1_1;
	wire w_dff_A_rE4qmGgL3_1;
	wire w_dff_A_ZHjSjUI17_0;
	wire w_dff_A_a5FiIX6v2_0;
	wire w_dff_A_GjJySaNj3_0;
	wire w_dff_A_qNBEAGXc1_0;
	wire w_dff_A_BU4rTDgm3_0;
	wire w_dff_A_fGX7JfCv5_0;
	wire w_dff_A_pr6bOVe40_0;
	wire w_dff_A_fE7kvKyq3_0;
	wire w_dff_A_44kvQYtZ7_0;
	wire w_dff_A_Qu8OTBtf4_0;
	wire w_dff_A_A30gUBkh9_0;
	wire w_dff_A_sGgHrYJb0_0;
	wire w_dff_A_AlYXZySL1_0;
	wire w_dff_A_7eGlORmV1_0;
	wire w_dff_A_4IMo6afp9_0;
	wire w_dff_A_9l1niQwx9_0;
	wire w_dff_A_77ogvPP86_0;
	wire w_dff_A_BHSr3EmJ0_0;
	wire w_dff_A_bjAgsrpW0_0;
	wire w_dff_A_NrivGG2h2_0;
	wire w_dff_A_XYj3p9UF8_0;
	wire w_dff_A_J9yBLkpz7_0;
	wire w_dff_A_itn12WyD8_0;
	wire w_dff_A_xu7skIGf8_0;
	wire w_dff_A_JcuAN9sZ9_0;
	wire w_dff_A_UqtOzkKK3_0;
	wire w_dff_A_KdfBZQGv4_0;
	wire w_dff_A_6YgT5HmA5_0;
	wire w_dff_A_1TftoEOW8_0;
	wire w_dff_A_USQYQHf75_0;
	wire w_dff_A_1D1Y6BUd5_0;
	wire w_dff_A_AGJH553l7_0;
	wire w_dff_A_hwq5kgka2_0;
	wire w_dff_A_YN4nNPtx9_0;
	wire w_dff_A_mtZguglp8_0;
	wire w_dff_A_yJGhVhhl3_0;
	wire w_dff_A_548WKCsg9_0;
	wire w_dff_A_mLPPM5sn6_0;
	wire w_dff_A_nrufeGX17_0;
	wire w_dff_A_4MqFCvoH0_0;
	wire w_dff_A_2zk8f1AU5_0;
	wire w_dff_A_AguR2ECu4_0;
	wire w_dff_A_ny7PYMA96_0;
	wire w_dff_A_98ErYpfl4_0;
	wire w_dff_A_qce9Ezw64_0;
	wire w_dff_A_LvmED0907_0;
	wire w_dff_A_ZrwPCZx36_0;
	wire w_dff_A_6Fb6qF1p2_0;
	wire w_dff_A_TTH40hc38_0;
	wire w_dff_A_8qhQPsyN2_0;
	wire w_dff_A_slabGQfO5_0;
	wire w_dff_A_lEDkFNI38_0;
	wire w_dff_A_iYmAUuzm0_0;
	wire w_dff_A_OlYLz6wX1_0;
	wire w_dff_A_dALT4q3n8_0;
	wire w_dff_A_CgyGOVCN8_0;
	wire w_dff_A_5gfEFDge0_0;
	wire w_dff_A_s78YTkNL7_0;
	wire w_dff_A_kPG8ZVs28_0;
	wire w_dff_A_WAUmUw6U6_0;
	wire w_dff_A_NPgZlsW65_0;
	wire w_dff_A_jOaAEEDT2_0;
	wire w_dff_A_PWbMRYmD2_0;
	wire w_dff_A_LM1FenCm6_0;
	wire w_dff_A_qHIUtCQv8_0;
	wire w_dff_A_NTuBIZC16_0;
	wire w_dff_A_irNDFiMt4_0;
	wire w_dff_A_P4linBrj6_0;
	wire w_dff_A_Giinq9195_0;
	wire w_dff_A_cYf0crjQ1_0;
	wire w_dff_A_VBKTxnU93_0;
	wire w_dff_A_aumP3CjT5_0;
	wire w_dff_A_98G6dCIX3_0;
	wire w_dff_A_P7Rt7lic5_0;
	wire w_dff_A_YXiv6Yx23_2;
	wire w_dff_A_p64RLqHA6_0;
	wire w_dff_A_Kc8P7odh1_0;
	wire w_dff_A_SjmfjdMv9_0;
	wire w_dff_A_5RDbOpvM5_0;
	wire w_dff_A_peI4Grcg6_0;
	wire w_dff_A_or75KAGO6_0;
	wire w_dff_A_wGvRFbvr5_0;
	wire w_dff_A_8B23OrgM6_0;
	wire w_dff_A_H3ssAJR90_0;
	wire w_dff_A_fzAJolga8_0;
	wire w_dff_A_jDtwgd2i4_0;
	wire w_dff_A_W2yE3rvl0_0;
	wire w_dff_A_PFsb8Yf51_0;
	wire w_dff_A_p7puu2no7_0;
	wire w_dff_A_vfDdvrFO3_0;
	wire w_dff_A_TTeC5tV14_0;
	wire w_dff_A_jzfbyS4I7_0;
	wire w_dff_A_i9vzbcfc5_0;
	wire w_dff_A_ktjbljTE0_0;
	wire w_dff_A_LVV36kZL1_0;
	wire w_dff_A_6CjaYoLO1_0;
	wire w_dff_A_HxOUhU9n0_0;
	wire w_dff_A_By7SmI832_0;
	wire w_dff_A_zxKvatpL2_0;
	wire w_dff_A_5ameRFIA4_0;
	wire w_dff_A_YcFPflsI3_0;
	wire w_dff_A_FKECd3dk6_0;
	wire w_dff_A_FOjuWzTf0_0;
	wire w_dff_A_OMTNsVM81_0;
	wire w_dff_A_JkSPIyLB4_0;
	wire w_dff_A_merzZsE68_0;
	wire w_dff_A_cdYbLOH19_0;
	wire w_dff_A_JGeJVqJn3_0;
	wire w_dff_A_S0FYVG1S0_0;
	wire w_dff_A_xgRwYFbb3_0;
	wire w_dff_A_8yiAk4tD8_0;
	wire w_dff_A_kpXii2qt5_0;
	wire w_dff_A_kpY6t2RW1_0;
	wire w_dff_A_LFJqh0xF9_0;
	wire w_dff_A_Ct3URjSe1_0;
	wire w_dff_A_LpTzvMRc1_0;
	wire w_dff_A_agohsC0X8_0;
	wire w_dff_A_05f6D0SG2_0;
	wire w_dff_A_MHH2uqGI2_0;
	wire w_dff_A_M8fUQQ3i5_0;
	wire w_dff_A_SF7FExQW6_0;
	wire w_dff_A_khpJA9Vz3_0;
	wire w_dff_A_N8OZYB3v1_0;
	wire w_dff_A_7G07MALF0_0;
	wire w_dff_A_MXdsDW6I3_0;
	wire w_dff_A_1CBWRDSR3_0;
	wire w_dff_A_YerZPohO3_0;
	wire w_dff_A_BhZ3RtV71_0;
	wire w_dff_A_rY2wFcGx5_0;
	wire w_dff_A_NxZsVi9t8_0;
	wire w_dff_A_7ZVKcPhK8_0;
	wire w_dff_A_U4GUl6kQ8_0;
	wire w_dff_A_D1V1DfQ07_0;
	wire w_dff_A_35XEmrYb4_0;
	wire w_dff_A_RhiqKDrt0_0;
	wire w_dff_A_Ulr0o6TO5_0;
	wire w_dff_A_aligU5lK9_0;
	wire w_dff_A_FAYZJtDj5_0;
	wire w_dff_A_JWJAKf7Q0_0;
	wire w_dff_A_KseXWj2U4_0;
	wire w_dff_A_TQU6YDac1_0;
	wire w_dff_A_BvEGz6x93_0;
	wire w_dff_A_UpFK9dU44_0;
	wire w_dff_A_2Yd292y00_0;
	wire w_dff_A_NoShJDYn0_0;
	wire w_dff_A_7LlMToQR5_0;
	wire w_dff_A_bk66JIRc7_2;
	wire w_dff_A_IKCfQeGD9_0;
	wire w_dff_A_lC3t4jek6_0;
	wire w_dff_A_n57bBGQP3_0;
	wire w_dff_A_Dpyr2gKH1_0;
	wire w_dff_A_o8HRGzKQ7_0;
	wire w_dff_A_V99KVqkz2_0;
	wire w_dff_A_teGtxT7P7_0;
	wire w_dff_A_ee17YuJ77_0;
	wire w_dff_A_16J9Ltb47_0;
	wire w_dff_A_itTsayCO6_0;
	wire w_dff_A_1ScT891b9_0;
	wire w_dff_A_fiuBGqNA6_0;
	wire w_dff_A_J5JYw0Cg9_0;
	wire w_dff_A_n6lkNNPd0_0;
	wire w_dff_A_GjzVWqgl2_0;
	wire w_dff_A_OsT9bsmP2_0;
	wire w_dff_A_IsUssCpU0_0;
	wire w_dff_A_LZmai8il1_0;
	wire w_dff_A_X0r76xsS0_0;
	wire w_dff_A_R6ur1G3R4_0;
	wire w_dff_A_WSus9DQn2_0;
	wire w_dff_A_ue27BoMK0_0;
	wire w_dff_A_B5EsmqgE8_0;
	wire w_dff_A_tPS7lwTn4_0;
	wire w_dff_A_sxyqDQwb0_0;
	wire w_dff_A_fJDhVgOz5_0;
	wire w_dff_A_Gox6RqJK1_0;
	wire w_dff_A_yWfJCSsM6_0;
	wire w_dff_A_npB4fh242_0;
	wire w_dff_A_ZJOgWIsk0_0;
	wire w_dff_A_cdoOIn1i1_0;
	wire w_dff_A_cpQj61Q11_0;
	wire w_dff_A_8u57dXdM6_0;
	wire w_dff_A_m6TfIlGV0_0;
	wire w_dff_A_YfxDWxVz7_0;
	wire w_dff_A_0iddeGKK0_0;
	wire w_dff_A_rfogrGqH8_0;
	wire w_dff_A_DWnq424u4_0;
	wire w_dff_A_qLjqvj5B3_0;
	wire w_dff_A_RYFMtx8M8_0;
	wire w_dff_A_9rqH1VZm4_0;
	wire w_dff_A_wNigYBvw4_0;
	wire w_dff_A_tR05fWiy5_0;
	wire w_dff_A_Ia2f72Ci3_0;
	wire w_dff_A_Yqpxj6UB9_0;
	wire w_dff_A_K11Uetar0_0;
	wire w_dff_A_pIIYnlCH7_0;
	wire w_dff_A_P5yrAl677_0;
	wire w_dff_A_ATBUR3tj3_0;
	wire w_dff_A_nD9hgrCF5_0;
	wire w_dff_A_NTln6Xsz8_0;
	wire w_dff_A_G2CKQlSS9_0;
	wire w_dff_A_qqjCttYu8_0;
	wire w_dff_A_8eNjoxBn4_0;
	wire w_dff_A_JFGtlC5t4_0;
	wire w_dff_A_KgoDcpQ35_0;
	wire w_dff_A_zVR9oK5w1_0;
	wire w_dff_A_mBg5cCz30_0;
	wire w_dff_A_wCUZ1sVW6_0;
	wire w_dff_A_rYcqg5M32_0;
	wire w_dff_A_KGNYuGTP1_0;
	wire w_dff_A_1AMb7ab21_0;
	wire w_dff_A_1yl3Tr0K0_0;
	wire w_dff_A_MYeHyNuP9_0;
	wire w_dff_A_dA0i9buk1_0;
	wire w_dff_A_UwY88ub12_0;
	wire w_dff_A_QOUpQTe75_0;
	wire w_dff_A_ZO8vVKK11_0;
	wire w_dff_A_ihkYZoXx2_2;
	wire w_dff_A_SC53etb39_0;
	wire w_dff_A_GTMw07LJ7_0;
	wire w_dff_A_abpLbixo1_0;
	wire w_dff_A_g6MFUHP52_0;
	wire w_dff_A_dIuFx3vT5_0;
	wire w_dff_A_mwkUC4UP9_0;
	wire w_dff_A_dVLD3Ro47_0;
	wire w_dff_A_kWQRDeEs6_0;
	wire w_dff_A_C5iXU3DY6_0;
	wire w_dff_A_P9xwoMHP3_0;
	wire w_dff_A_188WxzeC5_0;
	wire w_dff_A_c37TLJfK1_0;
	wire w_dff_A_l58SNuKq3_0;
	wire w_dff_A_guS0juLC7_0;
	wire w_dff_A_kAcV4oxf0_0;
	wire w_dff_A_ZIiaFsVb2_0;
	wire w_dff_A_wHt4zteD1_0;
	wire w_dff_A_DHMaLv0r3_0;
	wire w_dff_A_xzotiHdE6_0;
	wire w_dff_A_OJlLLM5O7_0;
	wire w_dff_A_Yg4WvvCX9_0;
	wire w_dff_A_gYj8Sm3I7_0;
	wire w_dff_A_Gi9v8lA62_0;
	wire w_dff_A_DSpPYdNM5_0;
	wire w_dff_A_xly4i3pr4_0;
	wire w_dff_A_lBDkvRUu2_0;
	wire w_dff_A_zQgRC7OG7_0;
	wire w_dff_A_2QpKr6gk8_0;
	wire w_dff_A_yZmlUCb06_0;
	wire w_dff_A_ozZXWHbn6_0;
	wire w_dff_A_TglgS7hl8_0;
	wire w_dff_A_E6nEfCKl2_0;
	wire w_dff_A_WvDEKKvF0_0;
	wire w_dff_A_NhVoXUf70_0;
	wire w_dff_A_Tjw3eYba6_0;
	wire w_dff_A_Df4bkLAL2_0;
	wire w_dff_A_GwQLWlZ29_0;
	wire w_dff_A_kJPi2ieZ8_0;
	wire w_dff_A_6kIevxMP0_0;
	wire w_dff_A_yJZO6A449_0;
	wire w_dff_A_IXbyTuFa5_0;
	wire w_dff_A_q8X3NXYg4_0;
	wire w_dff_A_CuZuBnGt2_0;
	wire w_dff_A_aUujZGe54_0;
	wire w_dff_A_Q9mGDfoZ7_0;
	wire w_dff_A_EOe5qfW22_0;
	wire w_dff_A_FslfGcvR1_0;
	wire w_dff_A_fUn8xO5C3_0;
	wire w_dff_A_lJ3FDdwu0_0;
	wire w_dff_A_KHvpRFUN1_0;
	wire w_dff_A_hVdqspZl2_0;
	wire w_dff_A_u1mu6W740_0;
	wire w_dff_A_KCMgCse62_0;
	wire w_dff_A_TvsniWpr4_0;
	wire w_dff_A_K1YnwdvK1_0;
	wire w_dff_A_72m3X7Vd2_0;
	wire w_dff_A_CrKFiCqf1_0;
	wire w_dff_A_dahJqzWt9_0;
	wire w_dff_A_HkFVYLsx4_0;
	wire w_dff_A_U61jtEFG5_0;
	wire w_dff_A_G2CYWKhS2_0;
	wire w_dff_A_deKqIOxp6_0;
	wire w_dff_A_jTlifDtK4_0;
	wire w_dff_A_7E3bbe5x1_0;
	wire w_dff_A_49Gda4N82_0;
	wire w_dff_A_u59OK6MR6_2;
	wire w_dff_A_AUDRS8GG1_0;
	wire w_dff_A_EdpmgK5y6_0;
	wire w_dff_A_ZiAS5RSm0_0;
	wire w_dff_A_nBUqx7vL4_0;
	wire w_dff_A_Tcg6oiJu6_0;
	wire w_dff_A_z0wpr7zP6_0;
	wire w_dff_A_6gqQAzuL4_0;
	wire w_dff_A_APpQpcHi8_0;
	wire w_dff_A_nyLnwlWy9_0;
	wire w_dff_A_tbpEb7BY9_0;
	wire w_dff_A_rOIcZZDu9_0;
	wire w_dff_A_Ja78ZvCe2_0;
	wire w_dff_A_CXGxDzkH2_0;
	wire w_dff_A_pnrcnN4J1_0;
	wire w_dff_A_UGT5LskC9_0;
	wire w_dff_A_AeEhZNnb2_0;
	wire w_dff_A_hJBYENos7_0;
	wire w_dff_A_AjK0qOSk1_0;
	wire w_dff_A_GBYgOpBd7_0;
	wire w_dff_A_QnVD2dQL5_0;
	wire w_dff_A_Fl6TlHCf6_0;
	wire w_dff_A_FbLdgRgn8_0;
	wire w_dff_A_wZULdw2L9_0;
	wire w_dff_A_QFUs9Ila8_0;
	wire w_dff_A_wJOokmHS5_0;
	wire w_dff_A_dEmfk64u5_0;
	wire w_dff_A_FVKsp7M03_0;
	wire w_dff_A_MvLXYLxv5_0;
	wire w_dff_A_CFZpnAs40_0;
	wire w_dff_A_LD930DMu4_0;
	wire w_dff_A_40sP0Bmi0_0;
	wire w_dff_A_PY1Wxqvw7_0;
	wire w_dff_A_Nk71cV790_0;
	wire w_dff_A_EvxITJEX9_0;
	wire w_dff_A_Kqrr3aOs4_0;
	wire w_dff_A_uYbfkqNb0_0;
	wire w_dff_A_ysW22CG84_0;
	wire w_dff_A_io4ikEzF2_0;
	wire w_dff_A_R0kt95vW2_0;
	wire w_dff_A_3pPmDxCy2_0;
	wire w_dff_A_cS8XrOzc9_0;
	wire w_dff_A_G4B3b3nI4_0;
	wire w_dff_A_v8EUxYoE6_0;
	wire w_dff_A_W1ZfZD3z6_0;
	wire w_dff_A_MYsLJGFR8_0;
	wire w_dff_A_wR71dWOy1_0;
	wire w_dff_A_xFfKk3BB7_0;
	wire w_dff_A_EPvQzi5F2_0;
	wire w_dff_A_S1jL8bHB9_0;
	wire w_dff_A_HnpzXgXD2_0;
	wire w_dff_A_8AIsEPAw5_0;
	wire w_dff_A_qpXikVWH1_0;
	wire w_dff_A_09EW2rDW4_0;
	wire w_dff_A_fR8LNZsj5_0;
	wire w_dff_A_gArMwLcF2_0;
	wire w_dff_A_csHlvfVS8_0;
	wire w_dff_A_qaoRYh0E1_0;
	wire w_dff_A_Ocxo46xu6_0;
	wire w_dff_A_KGlUjaKO8_0;
	wire w_dff_A_gkNXnR409_0;
	wire w_dff_A_nbpHtQDg8_0;
	wire w_dff_A_xu0HXtiL9_0;
	wire w_dff_A_RUYPQsDY7_2;
	wire w_dff_A_FERBmCp34_0;
	wire w_dff_A_lSRreIfz1_0;
	wire w_dff_A_D8PKPrPK0_0;
	wire w_dff_A_Wgwibnsv3_0;
	wire w_dff_A_3c7oaCSD7_0;
	wire w_dff_A_i9vTsd9D9_0;
	wire w_dff_A_aYXvXpA00_0;
	wire w_dff_A_gqknKMfQ0_0;
	wire w_dff_A_fKVkzAPb6_0;
	wire w_dff_A_J1woOXAB6_0;
	wire w_dff_A_RDyDpIKL3_0;
	wire w_dff_A_tGrCqxOn3_0;
	wire w_dff_A_TNghpsKr9_0;
	wire w_dff_A_B9jwKtEi0_0;
	wire w_dff_A_Mh1ZkqB01_0;
	wire w_dff_A_zDZVouRh0_0;
	wire w_dff_A_yUimV0Bh9_0;
	wire w_dff_A_RAueuALN5_0;
	wire w_dff_A_AxMvzLU83_0;
	wire w_dff_A_3gSVC3rH2_0;
	wire w_dff_A_awNIhsVs6_0;
	wire w_dff_A_G3QlGVPr3_0;
	wire w_dff_A_RhKMlQyO5_0;
	wire w_dff_A_QQyIJLSQ3_0;
	wire w_dff_A_O1DAztnV3_0;
	wire w_dff_A_QxPjcjDw3_0;
	wire w_dff_A_8Uat7pf94_0;
	wire w_dff_A_r8XYs8Hd3_0;
	wire w_dff_A_BdxTEUHS9_0;
	wire w_dff_A_qpsctrvC1_0;
	wire w_dff_A_lpZGXu0y2_0;
	wire w_dff_A_19fCI6Zc0_0;
	wire w_dff_A_XybjtclJ7_0;
	wire w_dff_A_Czx8K6yD4_0;
	wire w_dff_A_R9sSCIk98_0;
	wire w_dff_A_dn38EZaj9_0;
	wire w_dff_A_uQOZSzyv7_0;
	wire w_dff_A_YKdDcgJM5_0;
	wire w_dff_A_Rj33y8Qg2_0;
	wire w_dff_A_H0xHfJn59_0;
	wire w_dff_A_joOw27Ci1_0;
	wire w_dff_A_SH4AX4Fe8_0;
	wire w_dff_A_YIkkrbas4_0;
	wire w_dff_A_bnRvhZUK2_0;
	wire w_dff_A_Np5uqXUX6_0;
	wire w_dff_A_xgSBFmNI2_0;
	wire w_dff_A_MD9CjD6p0_0;
	wire w_dff_A_IMUfPG2y2_0;
	wire w_dff_A_jz5MI4T16_0;
	wire w_dff_A_8MbgAvdt1_0;
	wire w_dff_A_hvHqZMJY9_0;
	wire w_dff_A_0kYKmnQE1_0;
	wire w_dff_A_3K3I5SLN9_0;
	wire w_dff_A_hsBftZC11_0;
	wire w_dff_A_fj6EaFpb0_0;
	wire w_dff_A_f4420IxB5_0;
	wire w_dff_A_wn5HowOg8_0;
	wire w_dff_A_I9IweMtn6_0;
	wire w_dff_A_XQpzOOFe4_0;
	wire w_dff_A_3cNNDt623_2;
	wire w_dff_A_OeD4kmTb0_0;
	wire w_dff_A_gbjDoEu50_0;
	wire w_dff_A_sti6URCX3_0;
	wire w_dff_A_Ixj4wH3s3_0;
	wire w_dff_A_zqHGa9GZ9_0;
	wire w_dff_A_A4V818kf7_0;
	wire w_dff_A_d8LqlvIK9_0;
	wire w_dff_A_incpz5RR2_0;
	wire w_dff_A_SDcD5pXx9_0;
	wire w_dff_A_UIl9BgcD5_0;
	wire w_dff_A_oZzv7tR73_0;
	wire w_dff_A_RwzAJwkD4_0;
	wire w_dff_A_z4swIlhP5_0;
	wire w_dff_A_ET5BbgDx8_0;
	wire w_dff_A_dLTlhKMU5_0;
	wire w_dff_A_EIOYCWZT6_0;
	wire w_dff_A_i55dgTbi1_0;
	wire w_dff_A_lv79t8RY6_0;
	wire w_dff_A_m3MsK69G3_0;
	wire w_dff_A_wWCHn3aI2_0;
	wire w_dff_A_QYU6znvH3_0;
	wire w_dff_A_Yf2eC9iE3_0;
	wire w_dff_A_x75KIasX8_0;
	wire w_dff_A_cGlLDSgH2_0;
	wire w_dff_A_4BGdnQu19_0;
	wire w_dff_A_aWzaHUEc1_0;
	wire w_dff_A_IMY3fq3d2_0;
	wire w_dff_A_TfhU36SW1_0;
	wire w_dff_A_8aFoTaVN9_0;
	wire w_dff_A_tZSNMhT42_0;
	wire w_dff_A_P5Laq6MP6_0;
	wire w_dff_A_XhvDV9rF2_0;
	wire w_dff_A_lcAp889A4_0;
	wire w_dff_A_urBqOGvO9_0;
	wire w_dff_A_h5UpJryP1_0;
	wire w_dff_A_V3mBh8Xe1_0;
	wire w_dff_A_VVRS5WCw3_0;
	wire w_dff_A_KQEBDqy60_0;
	wire w_dff_A_mGKEe4Tn7_0;
	wire w_dff_A_MdjoMgUH1_0;
	wire w_dff_A_GD3P4vfF6_0;
	wire w_dff_A_SPWjq15W3_0;
	wire w_dff_A_SuSjSHB70_0;
	wire w_dff_A_KOXpkjoS4_0;
	wire w_dff_A_rPFu5ZpZ8_0;
	wire w_dff_A_Y70DArRS4_0;
	wire w_dff_A_nagS59Gw5_0;
	wire w_dff_A_DBTLQpSv1_0;
	wire w_dff_A_BWCZocTP7_0;
	wire w_dff_A_qZ22fWx69_0;
	wire w_dff_A_XXBn1gv58_0;
	wire w_dff_A_z29R41yA9_0;
	wire w_dff_A_2oBeUSdY0_0;
	wire w_dff_A_XdntmXwb6_0;
	wire w_dff_A_1KEcECGy0_0;
	wire w_dff_A_yJ4EGLoz5_0;
	wire w_dff_A_AWpHub178_2;
	wire w_dff_A_k1paZK0Y2_0;
	wire w_dff_A_ijtJorKs5_0;
	wire w_dff_A_DQ4C7Sfr2_0;
	wire w_dff_A_Xxke3TNk9_0;
	wire w_dff_A_LOY1HQbs4_0;
	wire w_dff_A_n8Qrp2Vw8_0;
	wire w_dff_A_8teEXTp34_0;
	wire w_dff_A_iWRwJXu99_0;
	wire w_dff_A_npqPB1Q28_0;
	wire w_dff_A_oijkPitJ0_0;
	wire w_dff_A_vZkmqeXs2_0;
	wire w_dff_A_OU5mnSOI7_0;
	wire w_dff_A_0Ej9uaVS9_0;
	wire w_dff_A_hmWynH6E1_0;
	wire w_dff_A_IAEEHCxV1_0;
	wire w_dff_A_R06KiJGO1_0;
	wire w_dff_A_xgL3MgNv9_0;
	wire w_dff_A_BPh9lray7_0;
	wire w_dff_A_AxcYoavu9_0;
	wire w_dff_A_VHTLPc0a7_0;
	wire w_dff_A_AcMpOlLu9_0;
	wire w_dff_A_3mqbvP4W1_0;
	wire w_dff_A_lecah2h29_0;
	wire w_dff_A_0yWtDODy3_0;
	wire w_dff_A_roPLPGKs4_0;
	wire w_dff_A_rfVEkmun7_0;
	wire w_dff_A_9nAAV3iw0_0;
	wire w_dff_A_MbeVzEdF9_0;
	wire w_dff_A_oqXMtO5e1_0;
	wire w_dff_A_9iXITTRO2_0;
	wire w_dff_A_bW12ClKR0_0;
	wire w_dff_A_BglbO1Nb1_0;
	wire w_dff_A_ZKRWuKQ48_0;
	wire w_dff_A_gUA9l13G5_0;
	wire w_dff_A_rYLWwpsi5_0;
	wire w_dff_A_nNAihJVP2_0;
	wire w_dff_A_KpCWsgbB6_0;
	wire w_dff_A_5TP7WeBX6_0;
	wire w_dff_A_pwjGtfFN2_0;
	wire w_dff_A_Clh6yr2s4_0;
	wire w_dff_A_0bmlHtoQ2_0;
	wire w_dff_A_NEVy6wJg0_0;
	wire w_dff_A_AABDCGJa1_0;
	wire w_dff_A_DyDEiMTR9_0;
	wire w_dff_A_0CHITjur6_0;
	wire w_dff_A_NWFLROeL9_0;
	wire w_dff_A_PrqbpDdw6_0;
	wire w_dff_A_vBxmA6LB5_0;
	wire w_dff_A_YDg62S291_0;
	wire w_dff_A_tGZYoIwU7_0;
	wire w_dff_A_e41qEz0N0_0;
	wire w_dff_A_XFF46Scq2_0;
	wire w_dff_A_E6Tczljx8_0;
	wire w_dff_A_8gCK9mkA1_2;
	wire w_dff_A_gZhCNXNw1_0;
	wire w_dff_A_JAUFx1H55_0;
	wire w_dff_A_3vcoTw601_0;
	wire w_dff_A_5YmVidb34_0;
	wire w_dff_A_5J3Q3rFA6_0;
	wire w_dff_A_qAgfKp1R4_0;
	wire w_dff_A_d3KWg11b4_0;
	wire w_dff_A_vlL9DLbv4_0;
	wire w_dff_A_mRhjIvPZ4_0;
	wire w_dff_A_Bblxg0SQ5_0;
	wire w_dff_A_7wu4IHuK6_0;
	wire w_dff_A_rnXu5VpJ8_0;
	wire w_dff_A_KWfWl4Vb3_0;
	wire w_dff_A_WIJih7lt7_0;
	wire w_dff_A_MNG0GSFM8_0;
	wire w_dff_A_Hx307nNz5_0;
	wire w_dff_A_QSNsEGjp8_0;
	wire w_dff_A_IIaFWszV3_0;
	wire w_dff_A_6ljpBP196_0;
	wire w_dff_A_yzWhyFCM4_0;
	wire w_dff_A_79dKQcCA6_0;
	wire w_dff_A_OxNPGvac0_0;
	wire w_dff_A_jcMpPvlb7_0;
	wire w_dff_A_FiLwcXha9_0;
	wire w_dff_A_T1zyELv61_0;
	wire w_dff_A_uwXDEM0t8_0;
	wire w_dff_A_WO0q5qOl7_0;
	wire w_dff_A_fVChj8QF5_0;
	wire w_dff_A_u5lQ2RIG2_0;
	wire w_dff_A_bMyFap6R8_0;
	wire w_dff_A_9LJ5SVdU0_0;
	wire w_dff_A_7SpiseeD3_0;
	wire w_dff_A_cHyQKoF31_0;
	wire w_dff_A_PCqNBvVU8_0;
	wire w_dff_A_UyEANOgG7_0;
	wire w_dff_A_97w0fdhi5_0;
	wire w_dff_A_GCTuFQdP2_0;
	wire w_dff_A_8xKbKkRf2_0;
	wire w_dff_A_GJiTmOg07_0;
	wire w_dff_A_iWyeoXsu8_0;
	wire w_dff_A_vGZPtRr95_0;
	wire w_dff_A_v1wARnUV7_0;
	wire w_dff_A_d8ZKm9L55_0;
	wire w_dff_A_uUTRxxwB7_0;
	wire w_dff_A_1I2yB0dQ3_0;
	wire w_dff_A_5tWePsnQ5_0;
	wire w_dff_A_QGDy6GMk4_0;
	wire w_dff_A_WPod74vA5_0;
	wire w_dff_A_hZpcWkUB7_0;
	wire w_dff_A_G853ioWQ5_0;
	wire w_dff_A_mdcJ4ar90_2;
	wire w_dff_A_ucXRuTTy6_0;
	wire w_dff_A_8wzFp3Rz4_0;
	wire w_dff_A_2Q16xPir4_0;
	wire w_dff_A_RD4HbXrN3_0;
	wire w_dff_A_j0fwaono3_0;
	wire w_dff_A_ErXFPDHr2_0;
	wire w_dff_A_lNjD4OkO5_0;
	wire w_dff_A_Ytk9gg1e7_0;
	wire w_dff_A_EEAvtlMp8_0;
	wire w_dff_A_apc6Yn0R8_0;
	wire w_dff_A_SDwRpmoh6_0;
	wire w_dff_A_5rDcnqKM0_0;
	wire w_dff_A_ewKztJgs5_0;
	wire w_dff_A_TFdvfNZE4_0;
	wire w_dff_A_JMBMXPot0_0;
	wire w_dff_A_FjyxqxJR5_0;
	wire w_dff_A_v1cz1S526_0;
	wire w_dff_A_3U3ruLjg7_0;
	wire w_dff_A_kdfXz4xG5_0;
	wire w_dff_A_J6LhkjTI5_0;
	wire w_dff_A_kkd0xx6G5_0;
	wire w_dff_A_E2RjHl9D8_0;
	wire w_dff_A_mPavfK0m8_0;
	wire w_dff_A_C4PI9ZpR7_0;
	wire w_dff_A_VdZlvEUK6_0;
	wire w_dff_A_ZWZPEdqW4_0;
	wire w_dff_A_gS7FByvC2_0;
	wire w_dff_A_EKThDx0b3_0;
	wire w_dff_A_zsBQAZrm8_0;
	wire w_dff_A_w6tNTT3C9_0;
	wire w_dff_A_yfka91WD1_0;
	wire w_dff_A_YJElB5c46_0;
	wire w_dff_A_p3iF3YJn8_0;
	wire w_dff_A_UFeWtC3S0_0;
	wire w_dff_A_EsM5A4XG5_0;
	wire w_dff_A_C06t6JTJ2_0;
	wire w_dff_A_PAynWK271_0;
	wire w_dff_A_rIywPZc71_0;
	wire w_dff_A_O50fT2260_0;
	wire w_dff_A_SjRZRti05_0;
	wire w_dff_A_6c2Zg5Hw8_0;
	wire w_dff_A_qc3faVvK6_0;
	wire w_dff_A_d0TPnhfP7_0;
	wire w_dff_A_BCvXb6co5_0;
	wire w_dff_A_kGMURzPc5_0;
	wire w_dff_A_TD0rCCw76_0;
	wire w_dff_A_UElGlsnx8_0;
	wire w_dff_A_Phb6U75D9_2;
	wire w_dff_A_mR2Eva228_0;
	wire w_dff_A_iiBkQspR7_0;
	wire w_dff_A_q4LRSY5y5_0;
	wire w_dff_A_Y84AA9ZC1_0;
	wire w_dff_A_Llfmmfo59_0;
	wire w_dff_A_DUTLKYQL6_0;
	wire w_dff_A_9aQLkix55_0;
	wire w_dff_A_YpfIfAzr6_0;
	wire w_dff_A_KNsYc6qM1_0;
	wire w_dff_A_ngcDbCQN1_0;
	wire w_dff_A_LUg8UohJ2_0;
	wire w_dff_A_FB2kpki42_0;
	wire w_dff_A_MVtKYeAe9_0;
	wire w_dff_A_xEF2irEO8_0;
	wire w_dff_A_nGGdf9zh1_0;
	wire w_dff_A_cTZlejHs1_0;
	wire w_dff_A_0JAzP6X92_0;
	wire w_dff_A_TShY5e1Z7_0;
	wire w_dff_A_Vy2WT7NC9_0;
	wire w_dff_A_0de3tUVL0_0;
	wire w_dff_A_GpRypKlf2_0;
	wire w_dff_A_iuQwrsgM3_0;
	wire w_dff_A_PZD3Cajo7_0;
	wire w_dff_A_EPf5hEiT1_0;
	wire w_dff_A_GoxV6nt89_0;
	wire w_dff_A_hE0m3T3e9_0;
	wire w_dff_A_3tX2e9C44_0;
	wire w_dff_A_jNyxx1wT6_0;
	wire w_dff_A_QJEE8DWm4_0;
	wire w_dff_A_PuXQpVOz3_0;
	wire w_dff_A_7XI49bBE6_0;
	wire w_dff_A_6XOZBCHi0_0;
	wire w_dff_A_85U7jzTf1_0;
	wire w_dff_A_MnTObEKb6_0;
	wire w_dff_A_o8iwBowI6_0;
	wire w_dff_A_nhjQHZwh3_0;
	wire w_dff_A_Oa3dy7Jx0_0;
	wire w_dff_A_moRygh1K1_0;
	wire w_dff_A_J86AyhRy1_0;
	wire w_dff_A_zsMZny7A9_0;
	wire w_dff_A_9jyakfJn9_0;
	wire w_dff_A_YmCBS2ot5_0;
	wire w_dff_A_vsJcTJdJ4_0;
	wire w_dff_A_H8sTOo013_0;
	wire w_dff_A_x2APV6JE4_2;
	wire w_dff_A_4ZUMfstK2_0;
	wire w_dff_A_8isAp7KB2_0;
	wire w_dff_A_4Z7Lme3u0_0;
	wire w_dff_A_bXFsMF1j7_0;
	wire w_dff_A_4IEEwk6D1_0;
	wire w_dff_A_m8vhnz8X6_0;
	wire w_dff_A_HYP6mTaq8_0;
	wire w_dff_A_u2lVkaxh5_0;
	wire w_dff_A_AdqfIWAB0_0;
	wire w_dff_A_EWuIz2Yi1_0;
	wire w_dff_A_2kzbZG6l7_0;
	wire w_dff_A_DeGW5AQc1_0;
	wire w_dff_A_NiH8YMgt1_0;
	wire w_dff_A_CnZPTTrA1_0;
	wire w_dff_A_BNP7UCab2_0;
	wire w_dff_A_KvAm47Gq4_0;
	wire w_dff_A_bMRb5fEI9_0;
	wire w_dff_A_HBs1nnTQ8_0;
	wire w_dff_A_AxWT3cyQ6_0;
	wire w_dff_A_0yEshw0C5_0;
	wire w_dff_A_hgW0cZ6R3_0;
	wire w_dff_A_1FU2AFeo8_0;
	wire w_dff_A_38nBbQo59_0;
	wire w_dff_A_TxihdmPS3_0;
	wire w_dff_A_PhBFujKQ8_0;
	wire w_dff_A_5R1Urcqo2_0;
	wire w_dff_A_PlGwnbl21_0;
	wire w_dff_A_9dQXlluI7_0;
	wire w_dff_A_2Bc3iSTU2_0;
	wire w_dff_A_2GQKVBUa4_0;
	wire w_dff_A_9BaNkW873_0;
	wire w_dff_A_YKM56Nk35_0;
	wire w_dff_A_iMAxdH4P7_0;
	wire w_dff_A_BMI7anqQ5_0;
	wire w_dff_A_kVagMUbd2_0;
	wire w_dff_A_bc52apDh2_0;
	wire w_dff_A_dRqHU3vM2_0;
	wire w_dff_A_jBG6z9Zz6_0;
	wire w_dff_A_HbMaSnJb1_0;
	wire w_dff_A_sGerDx5E0_0;
	wire w_dff_A_xgDN7rc03_0;
	wire w_dff_A_7vyaZLbT9_2;
	wire w_dff_A_rBGM1luv2_0;
	wire w_dff_A_lSs1vlGz9_0;
	wire w_dff_A_96qz8p685_0;
	wire w_dff_A_gxl8MQ4C1_0;
	wire w_dff_A_6Zc0b0fZ8_0;
	wire w_dff_A_UKQhSSBv1_0;
	wire w_dff_A_0Uc7yspJ2_0;
	wire w_dff_A_p2BWwzJt9_0;
	wire w_dff_A_jgqmBM7u3_0;
	wire w_dff_A_TC6LzhCv1_0;
	wire w_dff_A_lWMirraW9_0;
	wire w_dff_A_2fBCdJA41_0;
	wire w_dff_A_AgMpUUJg0_0;
	wire w_dff_A_qFMdeTVf4_0;
	wire w_dff_A_LMHMNP2S0_0;
	wire w_dff_A_My7pE2MQ1_0;
	wire w_dff_A_18ITMQEf6_0;
	wire w_dff_A_AUUizrVk3_0;
	wire w_dff_A_cEGfUJgl3_0;
	wire w_dff_A_oJXbKlhp9_0;
	wire w_dff_A_R70apvjg6_0;
	wire w_dff_A_hxDU4T4v5_0;
	wire w_dff_A_y09MRX6l3_0;
	wire w_dff_A_TUn1Bpxd1_0;
	wire w_dff_A_xDZBgepc1_0;
	wire w_dff_A_Avkw0D2G0_0;
	wire w_dff_A_3yAZ8lbo1_0;
	wire w_dff_A_Vb4wSG9j9_0;
	wire w_dff_A_Yh73tfam1_0;
	wire w_dff_A_vROip8wM3_0;
	wire w_dff_A_u3M4koVj4_0;
	wire w_dff_A_1OqLBf1z9_0;
	wire w_dff_A_wjoisF5K4_0;
	wire w_dff_A_6Sybiw3c3_0;
	wire w_dff_A_2AMhb9GJ6_0;
	wire w_dff_A_xvKm44JZ0_0;
	wire w_dff_A_LQ7uLL3z4_0;
	wire w_dff_A_SCqH8zVk4_0;
	wire w_dff_A_TEKx8qT56_2;
	wire w_dff_A_5mbaOIAJ7_0;
	wire w_dff_A_EeD76MjA9_0;
	wire w_dff_A_LEiV6ZbY0_0;
	wire w_dff_A_k3IAA0DQ1_0;
	wire w_dff_A_hUJ43Mx16_0;
	wire w_dff_A_9IUh5jR18_0;
	wire w_dff_A_AhKosuqg5_0;
	wire w_dff_A_LPRA2KEJ1_0;
	wire w_dff_A_2RppvQGd1_0;
	wire w_dff_A_hhlbElyG8_0;
	wire w_dff_A_uzU0o8xR2_0;
	wire w_dff_A_UINZN4gY4_0;
	wire w_dff_A_8cLKzRYr0_0;
	wire w_dff_A_vKxdlqmx2_0;
	wire w_dff_A_gqh9o9Uh4_0;
	wire w_dff_A_24sZSyuT2_0;
	wire w_dff_A_NqdZPWQn1_0;
	wire w_dff_A_AiBYpJBN9_0;
	wire w_dff_A_D50d9q789_0;
	wire w_dff_A_ac4B31Zm5_0;
	wire w_dff_A_s2yProDA8_0;
	wire w_dff_A_brPQUTpK2_0;
	wire w_dff_A_0XnJtovy0_0;
	wire w_dff_A_lsm4iIuD7_0;
	wire w_dff_A_F6jGdstK4_0;
	wire w_dff_A_SVNBHzQj6_0;
	wire w_dff_A_kBXQzIa09_0;
	wire w_dff_A_r43YaIL49_0;
	wire w_dff_A_Ltom9Con4_0;
	wire w_dff_A_raTQam683_0;
	wire w_dff_A_TiehvIPe1_0;
	wire w_dff_A_Vx8PwlVK2_0;
	wire w_dff_A_lBGpUiJc3_0;
	wire w_dff_A_ezVCfewI6_0;
	wire w_dff_A_miMC25NO6_0;
	wire w_dff_A_ND5rrPHV5_2;
	wire w_dff_A_rnAfQz647_0;
	wire w_dff_A_ZoFID5zg1_0;
	wire w_dff_A_noM0juy98_0;
	wire w_dff_A_UD61nGIn5_0;
	wire w_dff_A_dCcWln6m4_0;
	wire w_dff_A_iSE9KQJO4_0;
	wire w_dff_A_6luKBhuP9_0;
	wire w_dff_A_uNvo4nFD0_0;
	wire w_dff_A_64uUHRJo8_0;
	wire w_dff_A_DlEzE1mQ8_0;
	wire w_dff_A_4oxaVBo92_0;
	wire w_dff_A_a6yGjMhT8_0;
	wire w_dff_A_3vS5ofQE4_0;
	wire w_dff_A_uO5GxKNN4_0;
	wire w_dff_A_QGzY2HHp8_0;
	wire w_dff_A_ctOe0XbO7_0;
	wire w_dff_A_seMU5cwB7_0;
	wire w_dff_A_fJ2ksThq7_0;
	wire w_dff_A_kNbLuFPy1_0;
	wire w_dff_A_tDwSXBuX8_0;
	wire w_dff_A_TkTttgAE7_0;
	wire w_dff_A_1MceHRts7_0;
	wire w_dff_A_6ri971VA8_0;
	wire w_dff_A_KIrgp2FT9_0;
	wire w_dff_A_FxLDEICg3_0;
	wire w_dff_A_Q7ZELAT24_0;
	wire w_dff_A_49v8goCE1_0;
	wire w_dff_A_hBHHZSBk0_0;
	wire w_dff_A_yhb5xtMo9_0;
	wire w_dff_A_fD7qzMXK6_0;
	wire w_dff_A_BwrTxgv56_0;
	wire w_dff_A_7zApRyyX4_0;
	wire w_dff_A_NtHJwKOW4_2;
	wire w_dff_A_tTAugpDu8_0;
	wire w_dff_A_YArGBafw5_0;
	wire w_dff_A_WFPPUgIw0_0;
	wire w_dff_A_13jcXOoq3_0;
	wire w_dff_A_CkGOUhHZ3_0;
	wire w_dff_A_xiSZTgnd1_0;
	wire w_dff_A_XaxNQUaZ9_0;
	wire w_dff_A_sxEwDzW34_0;
	wire w_dff_A_aWMd9Avm2_0;
	wire w_dff_A_IjeC78Q92_0;
	wire w_dff_A_ExpXmqPP2_0;
	wire w_dff_A_ChGizsMB3_0;
	wire w_dff_A_jMGqfSc36_0;
	wire w_dff_A_4c4B0fIt5_0;
	wire w_dff_A_O2DG3k1q4_0;
	wire w_dff_A_eUEtAQCo4_0;
	wire w_dff_A_4bLZjiLN2_0;
	wire w_dff_A_wBb23zsF9_0;
	wire w_dff_A_Mo48ahrG7_0;
	wire w_dff_A_4uVDk40k9_0;
	wire w_dff_A_QPJq0wl87_0;
	wire w_dff_A_RIzwbEFv3_0;
	wire w_dff_A_wW8DdkE31_0;
	wire w_dff_A_G9Hukp1N3_0;
	wire w_dff_A_RqIx8HCk4_0;
	wire w_dff_A_ALOEaoHQ2_0;
	wire w_dff_A_UG3LSBeI9_0;
	wire w_dff_A_slTLL1i85_0;
	wire w_dff_A_fvjl21Pj0_0;
	wire w_dff_A_GkoBMSiy7_2;
	wire w_dff_A_dFa2grTs5_0;
	wire w_dff_A_gJhzoAqT4_0;
	wire w_dff_A_wzQDPlfJ8_0;
	wire w_dff_A_79cZBL3i4_0;
	wire w_dff_A_2pjyHanq4_0;
	wire w_dff_A_OSRhVY1y6_0;
	wire w_dff_A_zwZK5P7g3_0;
	wire w_dff_A_ELBK5l5c3_0;
	wire w_dff_A_v22zptni0_0;
	wire w_dff_A_p3wQVyqS2_0;
	wire w_dff_A_YVwbXvNp5_0;
	wire w_dff_A_vSa1ery42_0;
	wire w_dff_A_gp0tKW2z2_0;
	wire w_dff_A_w2Cxhf6o2_0;
	wire w_dff_A_q04g2wjQ5_0;
	wire w_dff_A_8ywlq8QD5_0;
	wire w_dff_A_Po2kMWjL0_0;
	wire w_dff_A_BZaa3w2n4_0;
	wire w_dff_A_6tTqPnQr9_0;
	wire w_dff_A_1gZyF6l89_0;
	wire w_dff_A_mjBcYgBA6_0;
	wire w_dff_A_c2YqTHKU9_0;
	wire w_dff_A_Mig4cTnu4_0;
	wire w_dff_A_2l8yetws1_0;
	wire w_dff_A_Y7CuQ6JA8_0;
	wire w_dff_A_kQnOLAU39_0;
	wire w_dff_A_5SPcpRbO5_0;
	wire w_dff_A_fgq1tWlH0_2;
	wire w_dff_A_FMBJe05O9_0;
	wire w_dff_A_4CLg10dh8_0;
	wire w_dff_A_LVL9bFe91_0;
	wire w_dff_A_oppvS8j14_0;
	wire w_dff_A_OSQHFrAg1_0;
	wire w_dff_A_ryMO8kaz0_0;
	wire w_dff_A_rYofgzWO9_0;
	wire w_dff_A_mBkmDaAr7_0;
	wire w_dff_A_oYaKYWwJ3_0;
	wire w_dff_A_NEEFFIV93_0;
	wire w_dff_A_NKLITBXP5_0;
	wire w_dff_A_KiciQbBH1_0;
	wire w_dff_A_tCRfYsDX5_0;
	wire w_dff_A_XyVUbH8F1_0;
	wire w_dff_A_diXooZ1c8_0;
	wire w_dff_A_JYl2zW550_0;
	wire w_dff_A_ChMB0Ynx5_0;
	wire w_dff_A_tLXdZOYV8_0;
	wire w_dff_A_aPx83fBB0_0;
	wire w_dff_A_kiSBccT21_0;
	wire w_dff_A_9aIz1G115_0;
	wire w_dff_A_VrkgbPSv9_0;
	wire w_dff_A_VvnvkjsB7_0;
	wire w_dff_A_bPuLvC5u3_0;
	wire w_dff_A_K0VMRFxq2_0;
	wire w_dff_A_obuUdNIl2_2;
	wire w_dff_A_3LVBNeEx3_0;
	wire w_dff_A_Xouw1Ph47_0;
	wire w_dff_A_wX4PHBXr0_0;
	wire w_dff_A_uzrl6ITp3_0;
	wire w_dff_A_RbZnFsIQ5_0;
	wire w_dff_A_DggnEZFj7_0;
	wire w_dff_A_PFmNnG3k8_0;
	wire w_dff_A_K9dQJapv8_0;
	wire w_dff_A_jYnAtpYq3_0;
	wire w_dff_A_ISuhW5kz7_0;
	wire w_dff_A_j8rDyhVM4_0;
	wire w_dff_A_ofAzioCB2_0;
	wire w_dff_A_tbZj41kF9_0;
	wire w_dff_A_vlDewE9B9_0;
	wire w_dff_A_ZPeyBSXX7_0;
	wire w_dff_A_wK1dcayQ8_0;
	wire w_dff_A_WEVIotbk2_0;
	wire w_dff_A_oIOw8cGC7_0;
	wire w_dff_A_HvckR75J2_0;
	wire w_dff_A_LwNB3OKs1_0;
	wire w_dff_A_kFu9MVUT3_0;
	wire w_dff_A_gM8cknpP4_0;
	wire w_dff_A_ytUpiMlJ5_0;
	wire w_dff_A_wJ6PBTgs4_0;
	wire w_dff_A_XYc3sDAs5_2;
	wire w_dff_A_s8Lz3PP21_0;
	wire w_dff_A_Vl6XXqKR4_0;
	wire w_dff_A_mIRvBGgs2_0;
	wire w_dff_A_j61eup6U3_0;
	wire w_dff_A_XzSjgAJD4_0;
	wire w_dff_A_qN60RfzG1_0;
	wire w_dff_A_gc57QrSY6_0;
	wire w_dff_A_l0SLvcbN7_0;
	wire w_dff_A_DrbsFgqW9_0;
	wire w_dff_A_N4255XaA4_0;
	wire w_dff_A_9t9c2ZSL7_0;
	wire w_dff_A_TwcTavwt2_0;
	wire w_dff_A_gGj8T90x1_0;
	wire w_dff_A_gSEeBq5e7_0;
	wire w_dff_A_LYPqDeu10_0;
	wire w_dff_A_Eo0iLPBH0_0;
	wire w_dff_A_IulUPpmL5_0;
	wire w_dff_A_qHkWz9bX2_0;
	wire w_dff_A_FdyIXHAm7_0;
	wire w_dff_A_WwhykUhZ0_0;
	wire w_dff_A_2s2nWD7l1_0;
	wire w_dff_A_jIx7cOiV7_0;
	wire w_dff_A_0iZHqm6h1_2;
	wire w_dff_A_prtqAZc98_0;
	wire w_dff_A_YziWlVof8_0;
	wire w_dff_A_UiZcUW5a0_0;
	wire w_dff_A_W2hvF0zz0_0;
	wire w_dff_A_xjdaaH8o2_0;
	wire w_dff_A_UfmbiT5a1_0;
	wire w_dff_A_dWzIwmUM7_0;
	wire w_dff_A_138kPFry8_0;
	wire w_dff_A_gTtrjauN9_0;
	wire w_dff_A_bLdR2FXj9_0;
	wire w_dff_A_W7qz9fsH8_0;
	wire w_dff_A_CaEvomZQ3_0;
	wire w_dff_A_mHVkNbvH7_0;
	wire w_dff_A_kJMyCwVs3_0;
	wire w_dff_A_8jUGBtcG2_0;
	wire w_dff_A_bOQ97r6R4_0;
	wire w_dff_A_T6qWt4nx7_0;
	wire w_dff_A_ixdpxXyl9_0;
	wire w_dff_A_QDexrUex8_0;
	wire w_dff_A_4Tot9Ke45_0;
	wire w_dff_A_DbIDePej4_2;
	wire w_dff_A_mGau4jRS5_0;
	wire w_dff_A_aQIhDYMB0_0;
	wire w_dff_A_QVEmwyc12_0;
	wire w_dff_A_1vdIsrcS5_0;
	wire w_dff_A_nUyTD8ts3_0;
	wire w_dff_A_u2jthr0Z6_0;
	wire w_dff_A_qQ7jFv5L9_0;
	wire w_dff_A_4KyxBQfF9_0;
	wire w_dff_A_pzlp7gQm8_0;
	wire w_dff_A_gQCbsAhm6_0;
	wire w_dff_A_oTcZHgAl7_0;
	wire w_dff_A_Tfh6mXU79_0;
	wire w_dff_A_RiKmipjv3_0;
	wire w_dff_A_JSEHANbP2_0;
	wire w_dff_A_OS4F2H9T4_0;
	wire w_dff_A_nNDroKgT3_0;
	wire w_dff_A_ryZ5pVjc1_0;
	wire w_dff_A_CwF0X3Qt5_0;
	wire w_dff_A_IUYnNff39_2;
	wire w_dff_A_xQeTjuds5_0;
	wire w_dff_A_U1EP0ICI1_0;
	wire w_dff_A_XPescyqL8_0;
	wire w_dff_A_6lpCmimB2_0;
	wire w_dff_A_vYYr7qNX5_0;
	wire w_dff_A_taIrpx5f3_0;
	wire w_dff_A_xU2xglG99_0;
	wire w_dff_A_fr2ZZxGV7_0;
	wire w_dff_A_Yq6pLs3I3_0;
	wire w_dff_A_KxfVw64E6_0;
	wire w_dff_A_uTlf0yaM5_0;
	wire w_dff_A_b9Imky7T9_0;
	wire w_dff_A_ngYzzIIk4_0;
	wire w_dff_A_LHDF6mO28_0;
	wire w_dff_A_Wqx6ig220_0;
	wire w_dff_A_q0ovqedw9_0;
	wire w_dff_A_bLrqy25k9_2;
	wire w_dff_A_Zvp8zY511_0;
	wire w_dff_A_3phXYowu3_0;
	wire w_dff_A_93feg0hY2_0;
	wire w_dff_A_h9JzAGb39_0;
	wire w_dff_A_EvwOX0nf7_0;
	wire w_dff_A_csAyt3t46_0;
	wire w_dff_A_XiOyo2uX4_0;
	wire w_dff_A_p3fTEORF6_0;
	wire w_dff_A_TNemDBlJ5_0;
	wire w_dff_A_AidrJimb7_0;
	wire w_dff_A_zvqnxQ0t7_0;
	wire w_dff_A_ReOMoYRg9_0;
	wire w_dff_A_FhgJ3KMa0_0;
	wire w_dff_A_zFU6cqn04_0;
	wire w_dff_A_LmfDc3mX7_2;
	wire w_dff_A_hboK2Rm15_0;
	wire w_dff_A_At2BKpWp7_0;
	wire w_dff_A_QV3e7I3m6_0;
	wire w_dff_A_CltQHqxN1_0;
	wire w_dff_A_EP4Nrif76_0;
	wire w_dff_A_EDFDqcWu2_0;
	wire w_dff_A_C9lOJ36M2_0;
	wire w_dff_A_KMCrbG5i2_0;
	wire w_dff_A_B1mpiYQK7_0;
	wire w_dff_A_VxSjdbXL3_0;
	wire w_dff_A_jemr7PEt7_0;
	wire w_dff_A_tVYZQ0xk2_0;
	wire w_dff_A_hXEXHGJP4_2;
	wire w_dff_A_Jd6PsPPu4_0;
	wire w_dff_A_JL78wWS26_0;
	wire w_dff_A_BovAFiDd6_0;
	wire w_dff_A_S33jOICy7_0;
	wire w_dff_A_LK6wRUxT8_0;
	wire w_dff_A_dMe4vE8R8_0;
	wire w_dff_A_PFx33hNw4_0;
	wire w_dff_A_fwuPYOIa2_0;
	wire w_dff_A_O5HVrv8X7_0;
	wire w_dff_A_v64lkwQT4_0;
	wire w_dff_A_3iLVSEwm9_2;
	wire w_dff_A_4W1dVK516_0;
	wire w_dff_A_NaxIzPxG7_0;
	wire w_dff_A_EGkVELoi0_0;
	wire w_dff_A_dpmFDk4l4_0;
	wire w_dff_A_zWPEkxoE8_0;
	wire w_dff_A_S2fxXnOh9_0;
	wire w_dff_A_pUDoKapv1_0;
	wire w_dff_A_he6AWlgo8_0;
	wire w_dff_A_ItMjlGlT1_2;
	wire w_dff_A_C1CdSTLN7_0;
	wire w_dff_A_W6uKVywC5_0;
	wire w_dff_A_GG2KKa2p5_0;
	wire w_dff_A_QFPb4j7j6_0;
	wire w_dff_A_C1glzCQw2_0;
	wire w_dff_A_VtpZWgPZ6_0;
	wire w_dff_A_WJUS03tP8_2;
	wire w_dff_A_4TathcMT6_0;
	wire w_dff_A_ifSQI7J07_0;
	wire w_dff_A_6OgvdeOL1_0;
	wire w_dff_A_MHHB6UYJ2_0;
	wire w_dff_A_8IBM46XT7_2;
	wire w_dff_A_PeO9O6Ih5_0;
	wire w_dff_A_Axb5Z3Rn6_0;
	wire w_dff_A_Sal8trTP1_2;
	jand g0000(.dina(w_G273gat_7[2]),.dinb(w_G1gat_7[1]),.dout(G545gat_fa_),.clk(gclk));
	jand g0001(.dina(w_G273gat_7[1]),.dinb(w_G18gat_7[2]),.dout(n65),.clk(gclk));
	jand g0002(.dina(w_G290gat_7[2]),.dinb(w_G1gat_7[0]),.dout(n66),.clk(gclk));
	jor g0003(.dina(n66),.dinb(w_n65_0[1]),.dout(n67),.clk(gclk));
	jand g0004(.dina(w_G290gat_7[1]),.dinb(w_G18gat_7[1]),.dout(n68),.clk(gclk));
	jand g0005(.dina(n68),.dinb(w_G545gat_0),.dout(n69),.clk(gclk));
	jnot g0006(.din(w_n69_0[1]),.dout(n70),.clk(gclk));
	jand g0007(.dina(w_n70_0[1]),.dinb(w_dff_B_ORLY9DPs0_1),.dout(w_dff_A_YXiv6Yx23_2),.clk(gclk));
	jand g0008(.dina(w_G307gat_7[2]),.dinb(w_G1gat_6[2]),.dout(n72),.clk(gclk));
	jnot g0009(.din(w_n72_0[1]),.dout(n73),.clk(gclk));
	jnot g0010(.din(w_G18gat_7[0]),.dout(n74),.clk(gclk));
	jnot g0011(.din(w_G290gat_7[0]),.dout(n75),.clk(gclk));
	jor g0012(.dina(w_n75_0[1]),.dinb(n74),.dout(n76),.clk(gclk));
	jnot g0013(.din(w_G35gat_7[2]),.dout(n77),.clk(gclk));
	jnot g0014(.din(w_G273gat_7[0]),.dout(n78),.clk(gclk));
	jor g0015(.dina(w_n78_0[1]),.dinb(w_n77_0[1]),.dout(n79),.clk(gclk));
	jand g0016(.dina(n79),.dinb(n76),.dout(n80),.clk(gclk));
	jand g0017(.dina(w_G290gat_6[2]),.dinb(w_G35gat_7[1]),.dout(n81),.clk(gclk));
	jand g0018(.dina(w_n81_0[1]),.dinb(w_n65_0[0]),.dout(n82),.clk(gclk));
	jor g0019(.dina(w_n82_1[1]),.dinb(n80),.dout(n83),.clk(gclk));
	jand g0020(.dina(n83),.dinb(w_n70_0[0]),.dout(n84),.clk(gclk));
	jnot g0021(.din(w_n82_1[0]),.dout(n85),.clk(gclk));
	jand g0022(.dina(w_n85_0[1]),.dinb(w_n69_0[0]),.dout(n86),.clk(gclk));
	jor g0023(.dina(w_dff_B_CNllXBTv4_0),.dinb(w_n84_0[1]),.dout(n87),.clk(gclk));
	jxor g0024(.dina(w_n87_0[1]),.dinb(w_dff_B_G2992b235_1),.dout(w_dff_A_bk66JIRc7_2),.clk(gclk));
	jand g0025(.dina(w_G324gat_7[1]),.dinb(w_G1gat_6[1]),.dout(n89),.clk(gclk));
	jnot g0026(.din(w_n89_0[1]),.dout(n90),.clk(gclk));
	jnot g0027(.din(w_n84_0[0]),.dout(n91),.clk(gclk));
	jor g0028(.dina(w_n87_0[0]),.dinb(w_n72_0[0]),.dout(n92),.clk(gclk));
	jand g0029(.dina(n92),.dinb(w_dff_B_GUp30YFz8_1),.dout(n93),.clk(gclk));
	jand g0030(.dina(w_G307gat_7[1]),.dinb(w_G18gat_6[2]),.dout(n94),.clk(gclk));
	jnot g0031(.din(w_n94_0[1]),.dout(n95),.clk(gclk));
	jand g0032(.dina(w_G273gat_6[2]),.dinb(w_G52gat_7[2]),.dout(n96),.clk(gclk));
	jor g0033(.dina(w_n96_0[1]),.dinb(w_n81_0[0]),.dout(n97),.clk(gclk));
	jand g0034(.dina(w_G273gat_6[1]),.dinb(w_G35gat_7[0]),.dout(n98),.clk(gclk));
	jand g0035(.dina(w_G290gat_6[1]),.dinb(w_G52gat_7[1]),.dout(n99),.clk(gclk));
	jand g0036(.dina(w_n99_0[1]),.dinb(n98),.dout(n100),.clk(gclk));
	jnot g0037(.din(w_n100_1[1]),.dout(n101),.clk(gclk));
	jand g0038(.dina(w_n101_0[2]),.dinb(w_dff_B_GTzGY71r8_1),.dout(n102),.clk(gclk));
	jor g0039(.dina(n102),.dinb(w_n82_0[2]),.dout(n103),.clk(gclk));
	jand g0040(.dina(w_n101_0[1]),.dinb(w_n82_0[1]),.dout(n104),.clk(gclk));
	jnot g0041(.din(w_n104_0[1]),.dout(n105),.clk(gclk));
	jand g0042(.dina(n105),.dinb(w_n103_0[1]),.dout(n106),.clk(gclk));
	jxor g0043(.dina(n106),.dinb(w_dff_B_jffWmVSl8_1),.dout(n107),.clk(gclk));
	jxor g0044(.dina(w_n107_0[1]),.dinb(w_n93_0[1]),.dout(n108),.clk(gclk));
	jxor g0045(.dina(w_n108_0[1]),.dinb(w_dff_B_YgdLPBYN7_1),.dout(w_dff_A_ihkYZoXx2_2),.clk(gclk));
	jand g0046(.dina(w_G341gat_7[1]),.dinb(w_G1gat_6[0]),.dout(n110),.clk(gclk));
	jnot g0047(.din(w_n110_0[1]),.dout(n111),.clk(gclk));
	jnot g0048(.din(w_n107_0[0]),.dout(n112),.clk(gclk));
	jor g0049(.dina(n112),.dinb(w_n93_0[0]),.dout(n113),.clk(gclk));
	jor g0050(.dina(w_n108_0[0]),.dinb(w_n89_0[0]),.dout(n114),.clk(gclk));
	jand g0051(.dina(n114),.dinb(w_dff_B_1qvD8ff13_1),.dout(n115),.clk(gclk));
	jand g0052(.dina(w_G324gat_7[0]),.dinb(w_G18gat_6[1]),.dout(n116),.clk(gclk));
	jnot g0053(.din(w_n116_0[1]),.dout(n117),.clk(gclk));
	jor g0054(.dina(w_n75_0[0]),.dinb(w_n77_0[0]),.dout(n118),.clk(gclk));
	jnot g0055(.din(w_G52gat_7[0]),.dout(n119),.clk(gclk));
	jor g0056(.dina(w_n78_0[0]),.dinb(n119),.dout(n120),.clk(gclk));
	jand g0057(.dina(n120),.dinb(n118),.dout(n121),.clk(gclk));
	jor g0058(.dina(w_n100_1[0]),.dinb(n121),.dout(n122),.clk(gclk));
	jand g0059(.dina(n122),.dinb(w_n85_0[0]),.dout(n123),.clk(gclk));
	jor g0060(.dina(w_n104_0[0]),.dinb(n123),.dout(n124),.clk(gclk));
	jor g0061(.dina(n124),.dinb(w_n94_0[0]),.dout(n125),.clk(gclk));
	jand g0062(.dina(n125),.dinb(w_n103_0[0]),.dout(n126),.clk(gclk));
	jand g0063(.dina(w_G307gat_7[0]),.dinb(w_G35gat_6[2]),.dout(n127),.clk(gclk));
	jnot g0064(.din(n127),.dout(n128),.clk(gclk));
	jand g0065(.dina(w_G273gat_6[0]),.dinb(w_G69gat_7[1]),.dout(n129),.clk(gclk));
	jor g0066(.dina(w_n129_0[1]),.dinb(w_n99_0[0]),.dout(n130),.clk(gclk));
	jand g0067(.dina(w_G290gat_6[0]),.dinb(w_G69gat_7[0]),.dout(n131),.clk(gclk));
	jand g0068(.dina(w_n131_0[1]),.dinb(w_n96_0[0]),.dout(n132),.clk(gclk));
	jnot g0069(.din(w_n132_0[2]),.dout(n133),.clk(gclk));
	jand g0070(.dina(w_n133_0[2]),.dinb(w_n130_0[1]),.dout(n134),.clk(gclk));
	jor g0071(.dina(n134),.dinb(w_n100_0[2]),.dout(n135),.clk(gclk));
	jand g0072(.dina(w_n133_0[1]),.dinb(w_n100_0[1]),.dout(n136),.clk(gclk));
	jnot g0073(.din(n136),.dout(n137),.clk(gclk));
	jand g0074(.dina(n137),.dinb(n135),.dout(n138),.clk(gclk));
	jxor g0075(.dina(w_n138_0[1]),.dinb(w_n128_0[1]),.dout(n139),.clk(gclk));
	jnot g0076(.din(w_n139_0[1]),.dout(n140),.clk(gclk));
	jxor g0077(.dina(w_n140_0[1]),.dinb(w_n126_0[2]),.dout(n141),.clk(gclk));
	jxor g0078(.dina(n141),.dinb(w_dff_B_tBHNWRrm0_1),.dout(n142),.clk(gclk));
	jxor g0079(.dina(w_n142_0[1]),.dinb(w_n115_0[1]),.dout(n143),.clk(gclk));
	jxor g0080(.dina(w_n143_0[1]),.dinb(w_dff_B_M40SSfNW0_1),.dout(w_dff_A_u59OK6MR6_2),.clk(gclk));
	jand g0081(.dina(w_G358gat_7[1]),.dinb(w_G1gat_5[2]),.dout(n145),.clk(gclk));
	jnot g0082(.din(w_n145_0[1]),.dout(n146),.clk(gclk));
	jnot g0083(.din(w_n142_0[0]),.dout(n147),.clk(gclk));
	jor g0084(.dina(n147),.dinb(w_n115_0[0]),.dout(n148),.clk(gclk));
	jor g0085(.dina(w_n143_0[0]),.dinb(w_n110_0[0]),.dout(n149),.clk(gclk));
	jand g0086(.dina(n149),.dinb(w_dff_B_TKqaCuwG8_1),.dout(n150),.clk(gclk));
	jand g0087(.dina(w_G341gat_7[0]),.dinb(w_G18gat_6[0]),.dout(n151),.clk(gclk));
	jnot g0088(.din(w_n151_0[1]),.dout(n152),.clk(gclk));
	jor g0089(.dina(w_n140_0[0]),.dinb(w_n126_0[1]),.dout(n153),.clk(gclk));
	jxor g0090(.dina(w_n139_0[0]),.dinb(w_n126_0[0]),.dout(n154),.clk(gclk));
	jor g0091(.dina(n154),.dinb(w_n116_0[0]),.dout(n155),.clk(gclk));
	jand g0092(.dina(n155),.dinb(w_dff_B_Mhfr6fth5_1),.dout(n156),.clk(gclk));
	jand g0093(.dina(w_G324gat_6[2]),.dinb(w_G35gat_6[1]),.dout(n157),.clk(gclk));
	jnot g0094(.din(n157),.dout(n158),.clk(gclk));
	jnot g0095(.din(w_n130_0[0]),.dout(n159),.clk(gclk));
	jor g0096(.dina(w_n132_0[1]),.dinb(n159),.dout(n160),.clk(gclk));
	jand g0097(.dina(n160),.dinb(w_n101_0[0]),.dout(n161),.clk(gclk));
	jand g0098(.dina(w_n138_0[0]),.dinb(w_n128_0[0]),.dout(n162),.clk(gclk));
	jor g0099(.dina(n162),.dinb(w_dff_B_jyMdLAoA5_1),.dout(n163),.clk(gclk));
	jand g0100(.dina(w_G307gat_6[2]),.dinb(w_G52gat_6[2]),.dout(n164),.clk(gclk));
	jnot g0101(.din(n164),.dout(n165),.clk(gclk));
	jand g0102(.dina(w_G273gat_5[2]),.dinb(w_G86gat_7[1]),.dout(n166),.clk(gclk));
	jor g0103(.dina(w_n166_0[1]),.dinb(w_n131_0[0]),.dout(n167),.clk(gclk));
	jand g0104(.dina(w_G290gat_5[2]),.dinb(w_G86gat_7[0]),.dout(n168),.clk(gclk));
	jand g0105(.dina(w_n168_0[1]),.dinb(w_n129_0[0]),.dout(n169),.clk(gclk));
	jnot g0106(.din(w_n169_0[2]),.dout(n170),.clk(gclk));
	jand g0107(.dina(w_n170_0[1]),.dinb(w_dff_B_owZoKCNi7_1),.dout(n171),.clk(gclk));
	jor g0108(.dina(n171),.dinb(w_n132_0[0]),.dout(n172),.clk(gclk));
	jor g0109(.dina(w_n169_0[1]),.dinb(w_n133_0[0]),.dout(n173),.clk(gclk));
	jand g0110(.dina(w_dff_B_CraBrRg64_0),.dinb(w_n172_0[1]),.dout(n174),.clk(gclk));
	jxor g0111(.dina(w_n174_0[1]),.dinb(w_n165_0[1]),.dout(n175),.clk(gclk));
	jxor g0112(.dina(w_n175_0[1]),.dinb(w_n163_0[1]),.dout(n176),.clk(gclk));
	jxor g0113(.dina(w_n176_0[1]),.dinb(w_n158_0[1]),.dout(n177),.clk(gclk));
	jnot g0114(.din(w_n177_0[1]),.dout(n178),.clk(gclk));
	jxor g0115(.dina(w_n178_0[1]),.dinb(w_n156_0[2]),.dout(n179),.clk(gclk));
	jxor g0116(.dina(n179),.dinb(w_dff_B_Y7QU2Ebk7_1),.dout(n180),.clk(gclk));
	jxor g0117(.dina(w_n180_0[1]),.dinb(w_n150_0[1]),.dout(n181),.clk(gclk));
	jxor g0118(.dina(w_n181_0[1]),.dinb(w_dff_B_Blu890lS8_1),.dout(w_dff_A_RUYPQsDY7_2),.clk(gclk));
	jand g0119(.dina(w_G375gat_7[1]),.dinb(w_G1gat_5[1]),.dout(n183),.clk(gclk));
	jnot g0120(.din(w_n183_0[1]),.dout(n184),.clk(gclk));
	jnot g0121(.din(w_n180_0[0]),.dout(n185),.clk(gclk));
	jor g0122(.dina(n185),.dinb(w_n150_0[0]),.dout(n186),.clk(gclk));
	jor g0123(.dina(w_n181_0[0]),.dinb(w_n145_0[0]),.dout(n187),.clk(gclk));
	jand g0124(.dina(n187),.dinb(w_dff_B_AwKqnTL31_1),.dout(n188),.clk(gclk));
	jand g0125(.dina(w_G358gat_7[0]),.dinb(w_G18gat_5[2]),.dout(n189),.clk(gclk));
	jnot g0126(.din(w_n189_0[1]),.dout(n190),.clk(gclk));
	jor g0127(.dina(w_n178_0[0]),.dinb(w_n156_0[1]),.dout(n191),.clk(gclk));
	jxor g0128(.dina(w_n177_0[0]),.dinb(w_n156_0[0]),.dout(n192),.clk(gclk));
	jor g0129(.dina(n192),.dinb(w_n151_0[0]),.dout(n193),.clk(gclk));
	jand g0130(.dina(n193),.dinb(w_dff_B_5lD7qqqs3_1),.dout(n194),.clk(gclk));
	jand g0131(.dina(w_G341gat_6[2]),.dinb(w_G35gat_6[0]),.dout(n195),.clk(gclk));
	jnot g0132(.din(n195),.dout(n196),.clk(gclk));
	jand g0133(.dina(w_n175_0[0]),.dinb(w_n163_0[0]),.dout(n197),.clk(gclk));
	jand g0134(.dina(w_n176_0[0]),.dinb(w_n158_0[0]),.dout(n198),.clk(gclk));
	jor g0135(.dina(n198),.dinb(w_dff_B_Rn758qRw2_1),.dout(n199),.clk(gclk));
	jand g0136(.dina(w_G324gat_6[1]),.dinb(w_G52gat_6[1]),.dout(n200),.clk(gclk));
	jnot g0137(.din(n200),.dout(n201),.clk(gclk));
	jnot g0138(.din(w_n172_0[0]),.dout(n202),.clk(gclk));
	jand g0139(.dina(w_n174_0[0]),.dinb(w_n165_0[0]),.dout(n203),.clk(gclk));
	jor g0140(.dina(n203),.dinb(w_dff_B_7gwb7JRl2_1),.dout(n204),.clk(gclk));
	jand g0141(.dina(w_G307gat_6[1]),.dinb(w_G69gat_6[2]),.dout(n205),.clk(gclk));
	jnot g0142(.din(n205),.dout(n206),.clk(gclk));
	jand g0143(.dina(w_G273gat_5[1]),.dinb(w_G103gat_7[1]),.dout(n207),.clk(gclk));
	jor g0144(.dina(w_n207_0[1]),.dinb(w_n168_0[0]),.dout(n208),.clk(gclk));
	jand g0145(.dina(w_G290gat_5[1]),.dinb(w_G103gat_7[0]),.dout(n209),.clk(gclk));
	jand g0146(.dina(w_n209_0[1]),.dinb(w_n166_0[0]),.dout(n210),.clk(gclk));
	jnot g0147(.din(w_n210_1[1]),.dout(n211),.clk(gclk));
	jand g0148(.dina(n211),.dinb(w_dff_B_74u3CizV5_1),.dout(n212),.clk(gclk));
	jor g0149(.dina(n212),.dinb(w_n169_0[0]),.dout(n213),.clk(gclk));
	jor g0150(.dina(w_n210_1[0]),.dinb(w_n170_0[0]),.dout(n214),.clk(gclk));
	jand g0151(.dina(w_dff_B_fEsB0Ljq9_0),.dinb(w_n213_0[1]),.dout(n215),.clk(gclk));
	jxor g0152(.dina(w_n215_0[1]),.dinb(w_n206_0[1]),.dout(n216),.clk(gclk));
	jxor g0153(.dina(w_n216_0[1]),.dinb(w_n204_0[1]),.dout(n217),.clk(gclk));
	jxor g0154(.dina(w_n217_0[1]),.dinb(w_n201_0[1]),.dout(n218),.clk(gclk));
	jxor g0155(.dina(w_n218_0[1]),.dinb(w_n199_0[1]),.dout(n219),.clk(gclk));
	jxor g0156(.dina(w_n219_0[1]),.dinb(w_n196_0[1]),.dout(n220),.clk(gclk));
	jnot g0157(.din(w_n220_0[1]),.dout(n221),.clk(gclk));
	jxor g0158(.dina(w_n221_0[1]),.dinb(w_n194_0[2]),.dout(n222),.clk(gclk));
	jxor g0159(.dina(n222),.dinb(w_dff_B_AmcbYULr1_1),.dout(n223),.clk(gclk));
	jxor g0160(.dina(w_n223_0[1]),.dinb(w_n188_0[1]),.dout(n224),.clk(gclk));
	jxor g0161(.dina(w_n224_0[1]),.dinb(w_dff_B_tADF5loM5_1),.dout(w_dff_A_3cNNDt623_2),.clk(gclk));
	jand g0162(.dina(w_G392gat_7[1]),.dinb(w_G1gat_5[0]),.dout(n226),.clk(gclk));
	jnot g0163(.din(w_n226_0[1]),.dout(n227),.clk(gclk));
	jnot g0164(.din(w_n223_0[0]),.dout(n228),.clk(gclk));
	jor g0165(.dina(n228),.dinb(w_n188_0[0]),.dout(n229),.clk(gclk));
	jor g0166(.dina(w_n224_0[0]),.dinb(w_n183_0[0]),.dout(n230),.clk(gclk));
	jand g0167(.dina(n230),.dinb(w_dff_B_rd8mdpko9_1),.dout(n231),.clk(gclk));
	jand g0168(.dina(w_G375gat_7[0]),.dinb(w_G18gat_5[1]),.dout(n232),.clk(gclk));
	jnot g0169(.din(w_n232_0[1]),.dout(n233),.clk(gclk));
	jor g0170(.dina(w_n221_0[0]),.dinb(w_n194_0[1]),.dout(n234),.clk(gclk));
	jxor g0171(.dina(w_n220_0[0]),.dinb(w_n194_0[0]),.dout(n235),.clk(gclk));
	jor g0172(.dina(n235),.dinb(w_n189_0[0]),.dout(n236),.clk(gclk));
	jand g0173(.dina(n236),.dinb(w_dff_B_0Uuq0fZ45_1),.dout(n237),.clk(gclk));
	jand g0174(.dina(w_G358gat_6[2]),.dinb(w_G35gat_5[2]),.dout(n238),.clk(gclk));
	jnot g0175(.din(n238),.dout(n239),.clk(gclk));
	jand g0176(.dina(w_n218_0[0]),.dinb(w_n199_0[0]),.dout(n240),.clk(gclk));
	jand g0177(.dina(w_n219_0[0]),.dinb(w_n196_0[0]),.dout(n241),.clk(gclk));
	jor g0178(.dina(n241),.dinb(w_dff_B_ncfFgBcp6_1),.dout(n242),.clk(gclk));
	jand g0179(.dina(w_G341gat_6[1]),.dinb(w_G52gat_6[0]),.dout(n243),.clk(gclk));
	jnot g0180(.din(n243),.dout(n244),.clk(gclk));
	jand g0181(.dina(w_n216_0[0]),.dinb(w_n204_0[0]),.dout(n245),.clk(gclk));
	jand g0182(.dina(w_n217_0[0]),.dinb(w_n201_0[0]),.dout(n246),.clk(gclk));
	jor g0183(.dina(n246),.dinb(w_dff_B_CzRkLVTi9_1),.dout(n247),.clk(gclk));
	jand g0184(.dina(w_G324gat_6[0]),.dinb(w_G69gat_6[1]),.dout(n248),.clk(gclk));
	jnot g0185(.din(n248),.dout(n249),.clk(gclk));
	jnot g0186(.din(w_n213_0[0]),.dout(n250),.clk(gclk));
	jand g0187(.dina(w_n215_0[0]),.dinb(w_n206_0[0]),.dout(n251),.clk(gclk));
	jor g0188(.dina(n251),.dinb(w_dff_B_BmR3h8NF0_1),.dout(n252),.clk(gclk));
	jand g0189(.dina(w_G307gat_6[0]),.dinb(w_G86gat_6[2]),.dout(n253),.clk(gclk));
	jnot g0190(.din(n253),.dout(n254),.clk(gclk));
	jand g0191(.dina(w_G273gat_5[0]),.dinb(w_G120gat_7[1]),.dout(n255),.clk(gclk));
	jor g0192(.dina(w_n255_0[1]),.dinb(w_n209_0[0]),.dout(n256),.clk(gclk));
	jand g0193(.dina(w_G290gat_5[0]),.dinb(w_G120gat_7[0]),.dout(n257),.clk(gclk));
	jand g0194(.dina(w_n257_0[1]),.dinb(w_n207_0[0]),.dout(n258),.clk(gclk));
	jnot g0195(.din(w_n258_0[2]),.dout(n259),.clk(gclk));
	jand g0196(.dina(w_n259_0[1]),.dinb(w_dff_B_9IuVKnvE7_1),.dout(n260),.clk(gclk));
	jor g0197(.dina(n260),.dinb(w_n210_0[2]),.dout(n261),.clk(gclk));
	jand g0198(.dina(w_n259_0[0]),.dinb(w_n210_0[1]),.dout(n262),.clk(gclk));
	jnot g0199(.din(n262),.dout(n263),.clk(gclk));
	jand g0200(.dina(n263),.dinb(w_n261_0[1]),.dout(n264),.clk(gclk));
	jxor g0201(.dina(w_n264_0[1]),.dinb(w_n254_0[1]),.dout(n265),.clk(gclk));
	jxor g0202(.dina(w_n265_0[1]),.dinb(w_n252_0[1]),.dout(n266),.clk(gclk));
	jxor g0203(.dina(w_n266_0[1]),.dinb(w_n249_0[1]),.dout(n267),.clk(gclk));
	jxor g0204(.dina(w_n267_0[1]),.dinb(w_n247_0[1]),.dout(n268),.clk(gclk));
	jxor g0205(.dina(w_n268_0[1]),.dinb(w_n244_0[1]),.dout(n269),.clk(gclk));
	jxor g0206(.dina(w_n269_0[1]),.dinb(w_n242_0[1]),.dout(n270),.clk(gclk));
	jxor g0207(.dina(w_n270_0[1]),.dinb(w_n239_0[1]),.dout(n271),.clk(gclk));
	jnot g0208(.din(w_n271_0[1]),.dout(n272),.clk(gclk));
	jxor g0209(.dina(w_n272_0[1]),.dinb(w_n237_0[2]),.dout(n273),.clk(gclk));
	jxor g0210(.dina(n273),.dinb(w_dff_B_txgUulhx8_1),.dout(n274),.clk(gclk));
	jxor g0211(.dina(w_n274_0[1]),.dinb(w_n231_0[1]),.dout(n275),.clk(gclk));
	jxor g0212(.dina(w_n275_0[1]),.dinb(w_dff_B_Rstyn61Z1_1),.dout(w_dff_A_AWpHub178_2),.clk(gclk));
	jand g0213(.dina(w_G409gat_7[1]),.dinb(w_G1gat_4[2]),.dout(n277),.clk(gclk));
	jnot g0214(.din(w_n277_0[1]),.dout(n278),.clk(gclk));
	jnot g0215(.din(w_n274_0[0]),.dout(n279),.clk(gclk));
	jor g0216(.dina(n279),.dinb(w_n231_0[0]),.dout(n280),.clk(gclk));
	jor g0217(.dina(w_n275_0[0]),.dinb(w_n226_0[0]),.dout(n281),.clk(gclk));
	jand g0218(.dina(n281),.dinb(w_dff_B_pRSP3AEO9_1),.dout(n282),.clk(gclk));
	jand g0219(.dina(w_G392gat_7[0]),.dinb(w_G18gat_5[0]),.dout(n283),.clk(gclk));
	jnot g0220(.din(w_n283_0[1]),.dout(n284),.clk(gclk));
	jor g0221(.dina(w_n272_0[0]),.dinb(w_n237_0[1]),.dout(n285),.clk(gclk));
	jxor g0222(.dina(w_n271_0[0]),.dinb(w_n237_0[0]),.dout(n286),.clk(gclk));
	jor g0223(.dina(n286),.dinb(w_n232_0[0]),.dout(n287),.clk(gclk));
	jand g0224(.dina(n287),.dinb(w_dff_B_t7zGmDAA3_1),.dout(n288),.clk(gclk));
	jand g0225(.dina(w_G375gat_6[2]),.dinb(w_G35gat_5[1]),.dout(n289),.clk(gclk));
	jnot g0226(.din(n289),.dout(n290),.clk(gclk));
	jand g0227(.dina(w_n269_0[0]),.dinb(w_n242_0[0]),.dout(n291),.clk(gclk));
	jand g0228(.dina(w_n270_0[0]),.dinb(w_n239_0[0]),.dout(n292),.clk(gclk));
	jor g0229(.dina(n292),.dinb(w_dff_B_6Fhf9Eju8_1),.dout(n293),.clk(gclk));
	jand g0230(.dina(w_G358gat_6[1]),.dinb(w_G52gat_5[2]),.dout(n294),.clk(gclk));
	jnot g0231(.din(n294),.dout(n295),.clk(gclk));
	jand g0232(.dina(w_n267_0[0]),.dinb(w_n247_0[0]),.dout(n296),.clk(gclk));
	jand g0233(.dina(w_n268_0[0]),.dinb(w_n244_0[0]),.dout(n297),.clk(gclk));
	jor g0234(.dina(n297),.dinb(w_dff_B_emUlAaqO8_1),.dout(n298),.clk(gclk));
	jand g0235(.dina(w_G341gat_6[0]),.dinb(w_G69gat_6[0]),.dout(n299),.clk(gclk));
	jnot g0236(.din(n299),.dout(n300),.clk(gclk));
	jand g0237(.dina(w_n265_0[0]),.dinb(w_n252_0[0]),.dout(n301),.clk(gclk));
	jand g0238(.dina(w_n266_0[0]),.dinb(w_n249_0[0]),.dout(n302),.clk(gclk));
	jor g0239(.dina(n302),.dinb(w_dff_B_lIUTpAE80_1),.dout(n303),.clk(gclk));
	jand g0240(.dina(w_G324gat_5[2]),.dinb(w_G86gat_6[1]),.dout(n304),.clk(gclk));
	jnot g0241(.din(n304),.dout(n305),.clk(gclk));
	jnot g0242(.din(w_n261_0[0]),.dout(n306),.clk(gclk));
	jand g0243(.dina(w_n264_0[0]),.dinb(w_n254_0[0]),.dout(n307),.clk(gclk));
	jor g0244(.dina(n307),.dinb(w_dff_B_p983pDwu3_1),.dout(n308),.clk(gclk));
	jand g0245(.dina(w_G307gat_5[2]),.dinb(w_G103gat_6[2]),.dout(n309),.clk(gclk));
	jnot g0246(.din(n309),.dout(n310),.clk(gclk));
	jand g0247(.dina(w_G273gat_4[2]),.dinb(w_G137gat_7[1]),.dout(n311),.clk(gclk));
	jor g0248(.dina(w_n311_0[1]),.dinb(w_n257_0[0]),.dout(n312),.clk(gclk));
	jand g0249(.dina(w_G290gat_4[2]),.dinb(w_G137gat_7[0]),.dout(n313),.clk(gclk));
	jand g0250(.dina(w_n313_0[1]),.dinb(w_n255_0[0]),.dout(n314),.clk(gclk));
	jnot g0251(.din(w_n314_0[2]),.dout(n315),.clk(gclk));
	jand g0252(.dina(w_n315_0[1]),.dinb(w_dff_B_pBKm8eeb1_1),.dout(n316),.clk(gclk));
	jor g0253(.dina(n316),.dinb(w_n258_0[1]),.dout(n317),.clk(gclk));
	jand g0254(.dina(w_n315_0[0]),.dinb(w_n258_0[0]),.dout(n318),.clk(gclk));
	jnot g0255(.din(n318),.dout(n319),.clk(gclk));
	jand g0256(.dina(n319),.dinb(w_n317_0[1]),.dout(n320),.clk(gclk));
	jxor g0257(.dina(w_n320_0[1]),.dinb(w_n310_0[1]),.dout(n321),.clk(gclk));
	jxor g0258(.dina(w_n321_0[1]),.dinb(w_n308_0[1]),.dout(n322),.clk(gclk));
	jxor g0259(.dina(w_n322_0[1]),.dinb(w_n305_0[1]),.dout(n323),.clk(gclk));
	jxor g0260(.dina(w_n323_0[1]),.dinb(w_n303_0[1]),.dout(n324),.clk(gclk));
	jxor g0261(.dina(w_n324_0[1]),.dinb(w_n300_0[1]),.dout(n325),.clk(gclk));
	jxor g0262(.dina(w_n325_0[1]),.dinb(w_n298_0[1]),.dout(n326),.clk(gclk));
	jxor g0263(.dina(w_n326_0[1]),.dinb(w_n295_0[1]),.dout(n327),.clk(gclk));
	jxor g0264(.dina(w_n327_0[1]),.dinb(w_n293_0[1]),.dout(n328),.clk(gclk));
	jxor g0265(.dina(w_n328_0[1]),.dinb(w_n290_0[1]),.dout(n329),.clk(gclk));
	jnot g0266(.din(w_n329_0[1]),.dout(n330),.clk(gclk));
	jxor g0267(.dina(w_n330_0[1]),.dinb(w_n288_0[2]),.dout(n331),.clk(gclk));
	jxor g0268(.dina(n331),.dinb(w_dff_B_U0LQCSR08_1),.dout(n332),.clk(gclk));
	jxor g0269(.dina(w_n332_0[1]),.dinb(w_n282_0[1]),.dout(n333),.clk(gclk));
	jxor g0270(.dina(w_n333_0[1]),.dinb(w_dff_B_sWvwVGJZ8_1),.dout(w_dff_A_8gCK9mkA1_2),.clk(gclk));
	jand g0271(.dina(w_G426gat_7[1]),.dinb(w_G1gat_4[1]),.dout(n335),.clk(gclk));
	jnot g0272(.din(w_n335_0[1]),.dout(n336),.clk(gclk));
	jnot g0273(.din(w_n332_0[0]),.dout(n337),.clk(gclk));
	jor g0274(.dina(n337),.dinb(w_n282_0[0]),.dout(n338),.clk(gclk));
	jor g0275(.dina(w_n333_0[0]),.dinb(w_n277_0[0]),.dout(n339),.clk(gclk));
	jand g0276(.dina(n339),.dinb(w_dff_B_AjWbN0rr3_1),.dout(n340),.clk(gclk));
	jand g0277(.dina(w_G409gat_7[0]),.dinb(w_G18gat_4[2]),.dout(n341),.clk(gclk));
	jnot g0278(.din(w_n341_0[1]),.dout(n342),.clk(gclk));
	jor g0279(.dina(w_n330_0[0]),.dinb(w_n288_0[1]),.dout(n343),.clk(gclk));
	jxor g0280(.dina(w_n329_0[0]),.dinb(w_n288_0[0]),.dout(n344),.clk(gclk));
	jor g0281(.dina(n344),.dinb(w_n283_0[0]),.dout(n345),.clk(gclk));
	jand g0282(.dina(n345),.dinb(w_dff_B_YN9xniCe7_1),.dout(n346),.clk(gclk));
	jand g0283(.dina(w_G392gat_6[2]),.dinb(w_G35gat_5[0]),.dout(n347),.clk(gclk));
	jnot g0284(.din(n347),.dout(n348),.clk(gclk));
	jand g0285(.dina(w_n327_0[0]),.dinb(w_n293_0[0]),.dout(n349),.clk(gclk));
	jand g0286(.dina(w_n328_0[0]),.dinb(w_n290_0[0]),.dout(n350),.clk(gclk));
	jor g0287(.dina(n350),.dinb(w_dff_B_QhBkAYhP6_1),.dout(n351),.clk(gclk));
	jand g0288(.dina(w_G375gat_6[1]),.dinb(w_G52gat_5[1]),.dout(n352),.clk(gclk));
	jnot g0289(.din(n352),.dout(n353),.clk(gclk));
	jand g0290(.dina(w_n325_0[0]),.dinb(w_n298_0[0]),.dout(n354),.clk(gclk));
	jand g0291(.dina(w_n326_0[0]),.dinb(w_n295_0[0]),.dout(n355),.clk(gclk));
	jor g0292(.dina(n355),.dinb(w_dff_B_YZOkLI4o6_1),.dout(n356),.clk(gclk));
	jand g0293(.dina(w_G358gat_6[0]),.dinb(w_G69gat_5[2]),.dout(n357),.clk(gclk));
	jnot g0294(.din(n357),.dout(n358),.clk(gclk));
	jand g0295(.dina(w_n323_0[0]),.dinb(w_n303_0[0]),.dout(n359),.clk(gclk));
	jand g0296(.dina(w_n324_0[0]),.dinb(w_n300_0[0]),.dout(n360),.clk(gclk));
	jor g0297(.dina(n360),.dinb(w_dff_B_ztAH3VDi4_1),.dout(n361),.clk(gclk));
	jand g0298(.dina(w_G341gat_5[2]),.dinb(w_G86gat_6[0]),.dout(n362),.clk(gclk));
	jnot g0299(.din(n362),.dout(n363),.clk(gclk));
	jand g0300(.dina(w_n321_0[0]),.dinb(w_n308_0[0]),.dout(n364),.clk(gclk));
	jand g0301(.dina(w_n322_0[0]),.dinb(w_n305_0[0]),.dout(n365),.clk(gclk));
	jor g0302(.dina(n365),.dinb(w_dff_B_TK43nvRb3_1),.dout(n366),.clk(gclk));
	jand g0303(.dina(w_G324gat_5[1]),.dinb(w_G103gat_6[1]),.dout(n367),.clk(gclk));
	jnot g0304(.din(n367),.dout(n368),.clk(gclk));
	jnot g0305(.din(w_n317_0[0]),.dout(n369),.clk(gclk));
	jand g0306(.dina(w_n320_0[0]),.dinb(w_n310_0[0]),.dout(n370),.clk(gclk));
	jor g0307(.dina(n370),.dinb(w_dff_B_03fXdbCs7_1),.dout(n371),.clk(gclk));
	jand g0308(.dina(w_G307gat_5[1]),.dinb(w_G120gat_6[2]),.dout(n372),.clk(gclk));
	jand g0309(.dina(w_G273gat_4[1]),.dinb(w_G154gat_7[1]),.dout(n373),.clk(gclk));
	jor g0310(.dina(w_n373_0[1]),.dinb(w_n313_0[0]),.dout(n374),.clk(gclk));
	jand g0311(.dina(w_G290gat_4[1]),.dinb(w_G154gat_7[0]),.dout(n375),.clk(gclk));
	jand g0312(.dina(w_n375_0[1]),.dinb(w_n311_0[0]),.dout(n376),.clk(gclk));
	jnot g0313(.din(w_n376_0[2]),.dout(n377),.clk(gclk));
	jand g0314(.dina(w_n377_0[1]),.dinb(w_dff_B_AuDEaiwK0_1),.dout(n378),.clk(gclk));
	jor g0315(.dina(n378),.dinb(w_n314_0[1]),.dout(n379),.clk(gclk));
	jnot g0316(.din(n379),.dout(n380),.clk(gclk));
	jand g0317(.dina(w_n377_0[0]),.dinb(w_n314_0[0]),.dout(n381),.clk(gclk));
	jor g0318(.dina(w_dff_B_L41QrBO30_0),.dinb(w_n380_0[1]),.dout(n382),.clk(gclk));
	jxor g0319(.dina(w_n382_0[1]),.dinb(w_n372_0[1]),.dout(n383),.clk(gclk));
	jxor g0320(.dina(w_n383_0[1]),.dinb(w_n371_0[1]),.dout(n384),.clk(gclk));
	jxor g0321(.dina(w_n384_0[1]),.dinb(w_n368_0[1]),.dout(n385),.clk(gclk));
	jxor g0322(.dina(w_n385_0[1]),.dinb(w_n366_0[1]),.dout(n386),.clk(gclk));
	jxor g0323(.dina(w_n386_0[1]),.dinb(w_n363_0[1]),.dout(n387),.clk(gclk));
	jxor g0324(.dina(w_n387_0[1]),.dinb(w_n361_0[1]),.dout(n388),.clk(gclk));
	jxor g0325(.dina(w_n388_0[1]),.dinb(w_n358_0[1]),.dout(n389),.clk(gclk));
	jxor g0326(.dina(w_n389_0[1]),.dinb(w_n356_0[1]),.dout(n390),.clk(gclk));
	jxor g0327(.dina(w_n390_0[1]),.dinb(w_n353_0[1]),.dout(n391),.clk(gclk));
	jxor g0328(.dina(w_n391_0[1]),.dinb(w_n351_0[1]),.dout(n392),.clk(gclk));
	jxor g0329(.dina(w_n392_0[1]),.dinb(w_n348_0[1]),.dout(n393),.clk(gclk));
	jnot g0330(.din(w_n393_0[1]),.dout(n394),.clk(gclk));
	jxor g0331(.dina(w_n394_0[1]),.dinb(w_n346_0[2]),.dout(n395),.clk(gclk));
	jxor g0332(.dina(n395),.dinb(w_dff_B_v1w7e7PW8_1),.dout(n396),.clk(gclk));
	jxor g0333(.dina(w_n396_0[1]),.dinb(w_n340_0[1]),.dout(n397),.clk(gclk));
	jxor g0334(.dina(w_n397_0[1]),.dinb(w_dff_B_EdoSg5X52_1),.dout(w_dff_A_mdcJ4ar90_2),.clk(gclk));
	jand g0335(.dina(w_G443gat_7[1]),.dinb(w_G1gat_4[0]),.dout(n399),.clk(gclk));
	jnot g0336(.din(w_n399_0[1]),.dout(n400),.clk(gclk));
	jnot g0337(.din(w_n396_0[0]),.dout(n401),.clk(gclk));
	jor g0338(.dina(n401),.dinb(w_n340_0[0]),.dout(n402),.clk(gclk));
	jor g0339(.dina(w_n397_0[0]),.dinb(w_n335_0[0]),.dout(n403),.clk(gclk));
	jand g0340(.dina(n403),.dinb(w_dff_B_ZBjdgUM75_1),.dout(n404),.clk(gclk));
	jand g0341(.dina(w_G426gat_7[0]),.dinb(w_G18gat_4[1]),.dout(n405),.clk(gclk));
	jnot g0342(.din(w_n405_0[1]),.dout(n406),.clk(gclk));
	jor g0343(.dina(w_n394_0[0]),.dinb(w_n346_0[1]),.dout(n407),.clk(gclk));
	jxor g0344(.dina(w_n393_0[0]),.dinb(w_n346_0[0]),.dout(n408),.clk(gclk));
	jor g0345(.dina(n408),.dinb(w_n341_0[0]),.dout(n409),.clk(gclk));
	jand g0346(.dina(n409),.dinb(w_dff_B_cNZdpEw14_1),.dout(n410),.clk(gclk));
	jand g0347(.dina(w_G409gat_6[2]),.dinb(w_G35gat_4[2]),.dout(n411),.clk(gclk));
	jnot g0348(.din(n411),.dout(n412),.clk(gclk));
	jand g0349(.dina(w_n391_0[0]),.dinb(w_n351_0[0]),.dout(n413),.clk(gclk));
	jand g0350(.dina(w_n392_0[0]),.dinb(w_n348_0[0]),.dout(n414),.clk(gclk));
	jor g0351(.dina(n414),.dinb(w_dff_B_Ha01Stdo7_1),.dout(n415),.clk(gclk));
	jand g0352(.dina(w_G392gat_6[1]),.dinb(w_G52gat_5[0]),.dout(n416),.clk(gclk));
	jnot g0353(.din(n416),.dout(n417),.clk(gclk));
	jand g0354(.dina(w_n389_0[0]),.dinb(w_n356_0[0]),.dout(n418),.clk(gclk));
	jand g0355(.dina(w_n390_0[0]),.dinb(w_n353_0[0]),.dout(n419),.clk(gclk));
	jor g0356(.dina(n419),.dinb(w_dff_B_dq2zZtCe8_1),.dout(n420),.clk(gclk));
	jand g0357(.dina(w_G375gat_6[0]),.dinb(w_G69gat_5[1]),.dout(n421),.clk(gclk));
	jnot g0358(.din(n421),.dout(n422),.clk(gclk));
	jand g0359(.dina(w_n387_0[0]),.dinb(w_n361_0[0]),.dout(n423),.clk(gclk));
	jand g0360(.dina(w_n388_0[0]),.dinb(w_n358_0[0]),.dout(n424),.clk(gclk));
	jor g0361(.dina(n424),.dinb(w_dff_B_UaNQnCtd9_1),.dout(n425),.clk(gclk));
	jand g0362(.dina(w_G358gat_5[2]),.dinb(w_G86gat_5[2]),.dout(n426),.clk(gclk));
	jnot g0363(.din(n426),.dout(n427),.clk(gclk));
	jand g0364(.dina(w_n385_0[0]),.dinb(w_n366_0[0]),.dout(n428),.clk(gclk));
	jand g0365(.dina(w_n386_0[0]),.dinb(w_n363_0[0]),.dout(n429),.clk(gclk));
	jor g0366(.dina(n429),.dinb(w_dff_B_BnZj7UBm8_1),.dout(n430),.clk(gclk));
	jand g0367(.dina(w_G341gat_5[1]),.dinb(w_G103gat_6[0]),.dout(n431),.clk(gclk));
	jnot g0368(.din(n431),.dout(n432),.clk(gclk));
	jand g0369(.dina(w_n383_0[0]),.dinb(w_n371_0[0]),.dout(n433),.clk(gclk));
	jand g0370(.dina(w_n384_0[0]),.dinb(w_n368_0[0]),.dout(n434),.clk(gclk));
	jor g0371(.dina(n434),.dinb(w_dff_B_OO1D15tP2_1),.dout(n435),.clk(gclk));
	jand g0372(.dina(w_G324gat_5[0]),.dinb(w_G120gat_6[1]),.dout(n436),.clk(gclk));
	jnot g0373(.din(n436),.dout(n437),.clk(gclk));
	jnot g0374(.din(w_n372_0[0]),.dout(n438),.clk(gclk));
	jnot g0375(.din(w_n382_0[0]),.dout(n439),.clk(gclk));
	jand g0376(.dina(n439),.dinb(w_dff_B_zin7EFie7_1),.dout(n440),.clk(gclk));
	jor g0377(.dina(n440),.dinb(w_n380_0[0]),.dout(n441),.clk(gclk));
	jand g0378(.dina(w_G307gat_5[0]),.dinb(w_G137gat_6[2]),.dout(n442),.clk(gclk));
	jand g0379(.dina(w_G273gat_4[0]),.dinb(w_G171gat_7[1]),.dout(n443),.clk(gclk));
	jor g0380(.dina(w_n443_0[1]),.dinb(w_n375_0[0]),.dout(n444),.clk(gclk));
	jand g0381(.dina(w_G290gat_4[0]),.dinb(w_G171gat_7[0]),.dout(n445),.clk(gclk));
	jand g0382(.dina(w_n445_0[1]),.dinb(w_n373_0[0]),.dout(n446),.clk(gclk));
	jnot g0383(.din(w_n446_0[2]),.dout(n447),.clk(gclk));
	jand g0384(.dina(w_n447_0[1]),.dinb(w_dff_B_kfrBW14e5_1),.dout(n448),.clk(gclk));
	jor g0385(.dina(n448),.dinb(w_n376_0[1]),.dout(n449),.clk(gclk));
	jnot g0386(.din(n449),.dout(n450),.clk(gclk));
	jand g0387(.dina(w_n447_0[0]),.dinb(w_n376_0[0]),.dout(n451),.clk(gclk));
	jor g0388(.dina(w_dff_B_fzZDPGCA0_0),.dinb(w_n450_0[1]),.dout(n452),.clk(gclk));
	jxor g0389(.dina(w_n452_0[1]),.dinb(w_n442_0[1]),.dout(n453),.clk(gclk));
	jxor g0390(.dina(w_n453_0[1]),.dinb(w_n441_0[1]),.dout(n454),.clk(gclk));
	jxor g0391(.dina(w_n454_0[1]),.dinb(w_n437_0[1]),.dout(n455),.clk(gclk));
	jxor g0392(.dina(w_n455_0[1]),.dinb(w_n435_0[1]),.dout(n456),.clk(gclk));
	jxor g0393(.dina(w_n456_0[1]),.dinb(w_n432_0[1]),.dout(n457),.clk(gclk));
	jxor g0394(.dina(w_n457_0[1]),.dinb(w_n430_0[1]),.dout(n458),.clk(gclk));
	jxor g0395(.dina(w_n458_0[1]),.dinb(w_n427_0[1]),.dout(n459),.clk(gclk));
	jxor g0396(.dina(w_n459_0[1]),.dinb(w_n425_0[1]),.dout(n460),.clk(gclk));
	jxor g0397(.dina(w_n460_0[1]),.dinb(w_n422_0[1]),.dout(n461),.clk(gclk));
	jxor g0398(.dina(w_n461_0[1]),.dinb(w_n420_0[1]),.dout(n462),.clk(gclk));
	jxor g0399(.dina(w_n462_0[1]),.dinb(w_n417_0[1]),.dout(n463),.clk(gclk));
	jxor g0400(.dina(w_n463_0[1]),.dinb(w_n415_0[1]),.dout(n464),.clk(gclk));
	jxor g0401(.dina(w_n464_0[1]),.dinb(w_n412_0[1]),.dout(n465),.clk(gclk));
	jnot g0402(.din(w_n465_0[1]),.dout(n466),.clk(gclk));
	jxor g0403(.dina(w_n466_0[1]),.dinb(w_n410_0[2]),.dout(n467),.clk(gclk));
	jxor g0404(.dina(n467),.dinb(w_dff_B_wop3Ppbk9_1),.dout(n468),.clk(gclk));
	jxor g0405(.dina(w_n468_0[1]),.dinb(w_n404_0[1]),.dout(n469),.clk(gclk));
	jxor g0406(.dina(w_n469_0[1]),.dinb(w_dff_B_wgsWXVkt3_1),.dout(w_dff_A_Phb6U75D9_2),.clk(gclk));
	jand g0407(.dina(w_G460gat_7[1]),.dinb(w_G1gat_3[2]),.dout(n471),.clk(gclk));
	jnot g0408(.din(w_n471_0[1]),.dout(n472),.clk(gclk));
	jnot g0409(.din(w_n468_0[0]),.dout(n473),.clk(gclk));
	jor g0410(.dina(n473),.dinb(w_n404_0[0]),.dout(n474),.clk(gclk));
	jor g0411(.dina(w_n469_0[0]),.dinb(w_n399_0[0]),.dout(n475),.clk(gclk));
	jand g0412(.dina(n475),.dinb(w_dff_B_DQfbDQM90_1),.dout(n476),.clk(gclk));
	jand g0413(.dina(w_G443gat_7[0]),.dinb(w_G18gat_4[0]),.dout(n477),.clk(gclk));
	jnot g0414(.din(w_n477_0[1]),.dout(n478),.clk(gclk));
	jor g0415(.dina(w_n466_0[0]),.dinb(w_n410_0[1]),.dout(n479),.clk(gclk));
	jxor g0416(.dina(w_n465_0[0]),.dinb(w_n410_0[0]),.dout(n480),.clk(gclk));
	jor g0417(.dina(n480),.dinb(w_n405_0[0]),.dout(n481),.clk(gclk));
	jand g0418(.dina(n481),.dinb(w_dff_B_wkFc1ith2_1),.dout(n482),.clk(gclk));
	jand g0419(.dina(w_G426gat_6[2]),.dinb(w_G35gat_4[1]),.dout(n483),.clk(gclk));
	jnot g0420(.din(n483),.dout(n484),.clk(gclk));
	jand g0421(.dina(w_n463_0[0]),.dinb(w_n415_0[0]),.dout(n485),.clk(gclk));
	jand g0422(.dina(w_n464_0[0]),.dinb(w_n412_0[0]),.dout(n486),.clk(gclk));
	jor g0423(.dina(n486),.dinb(w_dff_B_VdB4vGKp5_1),.dout(n487),.clk(gclk));
	jand g0424(.dina(w_G409gat_6[1]),.dinb(w_G52gat_4[2]),.dout(n488),.clk(gclk));
	jnot g0425(.din(n488),.dout(n489),.clk(gclk));
	jand g0426(.dina(w_n461_0[0]),.dinb(w_n420_0[0]),.dout(n490),.clk(gclk));
	jand g0427(.dina(w_n462_0[0]),.dinb(w_n417_0[0]),.dout(n491),.clk(gclk));
	jor g0428(.dina(n491),.dinb(w_dff_B_P8KsRJix4_1),.dout(n492),.clk(gclk));
	jand g0429(.dina(w_G392gat_6[0]),.dinb(w_G69gat_5[0]),.dout(n493),.clk(gclk));
	jnot g0430(.din(n493),.dout(n494),.clk(gclk));
	jand g0431(.dina(w_n459_0[0]),.dinb(w_n425_0[0]),.dout(n495),.clk(gclk));
	jand g0432(.dina(w_n460_0[0]),.dinb(w_n422_0[0]),.dout(n496),.clk(gclk));
	jor g0433(.dina(n496),.dinb(w_dff_B_VvhQZ0NB6_1),.dout(n497),.clk(gclk));
	jand g0434(.dina(w_G375gat_5[2]),.dinb(w_G86gat_5[1]),.dout(n498),.clk(gclk));
	jnot g0435(.din(n498),.dout(n499),.clk(gclk));
	jand g0436(.dina(w_n457_0[0]),.dinb(w_n430_0[0]),.dout(n500),.clk(gclk));
	jand g0437(.dina(w_n458_0[0]),.dinb(w_n427_0[0]),.dout(n501),.clk(gclk));
	jor g0438(.dina(n501),.dinb(w_dff_B_qAkQqxEW1_1),.dout(n502),.clk(gclk));
	jand g0439(.dina(w_G358gat_5[1]),.dinb(w_G103gat_5[2]),.dout(n503),.clk(gclk));
	jnot g0440(.din(n503),.dout(n504),.clk(gclk));
	jand g0441(.dina(w_n455_0[0]),.dinb(w_n435_0[0]),.dout(n505),.clk(gclk));
	jand g0442(.dina(w_n456_0[0]),.dinb(w_n432_0[0]),.dout(n506),.clk(gclk));
	jor g0443(.dina(n506),.dinb(w_dff_B_o1AElAy04_1),.dout(n507),.clk(gclk));
	jand g0444(.dina(w_G341gat_5[0]),.dinb(w_G120gat_6[0]),.dout(n508),.clk(gclk));
	jnot g0445(.din(n508),.dout(n509),.clk(gclk));
	jand g0446(.dina(w_n453_0[0]),.dinb(w_n441_0[0]),.dout(n510),.clk(gclk));
	jand g0447(.dina(w_n454_0[0]),.dinb(w_n437_0[0]),.dout(n511),.clk(gclk));
	jor g0448(.dina(n511),.dinb(w_dff_B_fr234X5Q7_1),.dout(n512),.clk(gclk));
	jand g0449(.dina(w_G324gat_4[2]),.dinb(w_G137gat_6[1]),.dout(n513),.clk(gclk));
	jnot g0450(.din(n513),.dout(n514),.clk(gclk));
	jnot g0451(.din(w_n442_0[0]),.dout(n515),.clk(gclk));
	jnot g0452(.din(w_n452_0[0]),.dout(n516),.clk(gclk));
	jand g0453(.dina(n516),.dinb(w_dff_B_Oo0S0JvP8_1),.dout(n517),.clk(gclk));
	jor g0454(.dina(n517),.dinb(w_n450_0[0]),.dout(n518),.clk(gclk));
	jand g0455(.dina(w_G307gat_4[2]),.dinb(w_G154gat_6[2]),.dout(n519),.clk(gclk));
	jand g0456(.dina(w_G273gat_3[2]),.dinb(w_G188gat_7[1]),.dout(n520),.clk(gclk));
	jor g0457(.dina(w_n520_0[1]),.dinb(w_n445_0[0]),.dout(n521),.clk(gclk));
	jand g0458(.dina(w_G290gat_3[2]),.dinb(w_G188gat_7[0]),.dout(n522),.clk(gclk));
	jand g0459(.dina(w_n522_0[1]),.dinb(w_n443_0[0]),.dout(n523),.clk(gclk));
	jnot g0460(.din(w_n523_0[2]),.dout(n524),.clk(gclk));
	jand g0461(.dina(w_n524_0[1]),.dinb(w_dff_B_pIrr73m08_1),.dout(n525),.clk(gclk));
	jor g0462(.dina(n525),.dinb(w_n446_0[1]),.dout(n526),.clk(gclk));
	jnot g0463(.din(n526),.dout(n527),.clk(gclk));
	jand g0464(.dina(w_n524_0[0]),.dinb(w_n446_0[0]),.dout(n528),.clk(gclk));
	jor g0465(.dina(w_dff_B_5EYqdB1x0_0),.dinb(w_n527_0[1]),.dout(n529),.clk(gclk));
	jxor g0466(.dina(w_n529_0[1]),.dinb(w_n519_0[1]),.dout(n530),.clk(gclk));
	jxor g0467(.dina(w_n530_0[1]),.dinb(w_n518_0[1]),.dout(n531),.clk(gclk));
	jxor g0468(.dina(w_n531_0[1]),.dinb(w_n514_0[1]),.dout(n532),.clk(gclk));
	jxor g0469(.dina(w_n532_0[1]),.dinb(w_n512_0[1]),.dout(n533),.clk(gclk));
	jxor g0470(.dina(w_n533_0[1]),.dinb(w_n509_0[1]),.dout(n534),.clk(gclk));
	jxor g0471(.dina(w_n534_0[1]),.dinb(w_n507_0[1]),.dout(n535),.clk(gclk));
	jxor g0472(.dina(w_n535_0[1]),.dinb(w_n504_0[1]),.dout(n536),.clk(gclk));
	jxor g0473(.dina(w_n536_0[1]),.dinb(w_n502_0[1]),.dout(n537),.clk(gclk));
	jxor g0474(.dina(w_n537_0[1]),.dinb(w_n499_0[1]),.dout(n538),.clk(gclk));
	jxor g0475(.dina(w_n538_0[1]),.dinb(w_n497_0[1]),.dout(n539),.clk(gclk));
	jxor g0476(.dina(w_n539_0[1]),.dinb(w_n494_0[1]),.dout(n540),.clk(gclk));
	jxor g0477(.dina(w_n540_0[1]),.dinb(w_n492_0[1]),.dout(n541),.clk(gclk));
	jxor g0478(.dina(w_n541_0[1]),.dinb(w_n489_0[1]),.dout(n542),.clk(gclk));
	jxor g0479(.dina(w_n542_0[1]),.dinb(w_n487_0[1]),.dout(n543),.clk(gclk));
	jxor g0480(.dina(w_n543_0[1]),.dinb(w_n484_0[1]),.dout(n544),.clk(gclk));
	jnot g0481(.din(w_n544_0[1]),.dout(n545),.clk(gclk));
	jxor g0482(.dina(w_n545_0[1]),.dinb(w_n482_0[2]),.dout(n546),.clk(gclk));
	jxor g0483(.dina(n546),.dinb(w_dff_B_9nDqJSLu7_1),.dout(n547),.clk(gclk));
	jxor g0484(.dina(w_n547_0[1]),.dinb(w_n476_0[1]),.dout(n548),.clk(gclk));
	jxor g0485(.dina(w_n548_0[1]),.dinb(w_dff_B_g6Pg8PGz3_1),.dout(w_dff_A_x2APV6JE4_2),.clk(gclk));
	jand g0486(.dina(w_G477gat_7[1]),.dinb(w_G1gat_3[1]),.dout(n550),.clk(gclk));
	jnot g0487(.din(w_n550_0[1]),.dout(n551),.clk(gclk));
	jnot g0488(.din(w_n547_0[0]),.dout(n552),.clk(gclk));
	jor g0489(.dina(n552),.dinb(w_n476_0[0]),.dout(n553),.clk(gclk));
	jor g0490(.dina(w_n548_0[0]),.dinb(w_n471_0[0]),.dout(n554),.clk(gclk));
	jand g0491(.dina(n554),.dinb(w_dff_B_qOHS1r4z9_1),.dout(n555),.clk(gclk));
	jand g0492(.dina(w_G460gat_7[0]),.dinb(w_G18gat_3[2]),.dout(n556),.clk(gclk));
	jnot g0493(.din(w_n556_0[1]),.dout(n557),.clk(gclk));
	jor g0494(.dina(w_n545_0[0]),.dinb(w_n482_0[1]),.dout(n558),.clk(gclk));
	jxor g0495(.dina(w_n544_0[0]),.dinb(w_n482_0[0]),.dout(n559),.clk(gclk));
	jor g0496(.dina(n559),.dinb(w_n477_0[0]),.dout(n560),.clk(gclk));
	jand g0497(.dina(n560),.dinb(w_dff_B_SpoUZEwd0_1),.dout(n561),.clk(gclk));
	jand g0498(.dina(w_G443gat_6[2]),.dinb(w_G35gat_4[0]),.dout(n562),.clk(gclk));
	jnot g0499(.din(n562),.dout(n563),.clk(gclk));
	jand g0500(.dina(w_n542_0[0]),.dinb(w_n487_0[0]),.dout(n564),.clk(gclk));
	jand g0501(.dina(w_n543_0[0]),.dinb(w_n484_0[0]),.dout(n565),.clk(gclk));
	jor g0502(.dina(n565),.dinb(w_dff_B_LdbHXJz70_1),.dout(n566),.clk(gclk));
	jand g0503(.dina(w_G426gat_6[1]),.dinb(w_G52gat_4[1]),.dout(n567),.clk(gclk));
	jnot g0504(.din(n567),.dout(n568),.clk(gclk));
	jand g0505(.dina(w_n540_0[0]),.dinb(w_n492_0[0]),.dout(n569),.clk(gclk));
	jand g0506(.dina(w_n541_0[0]),.dinb(w_n489_0[0]),.dout(n570),.clk(gclk));
	jor g0507(.dina(n570),.dinb(w_dff_B_sfAyzdid9_1),.dout(n571),.clk(gclk));
	jand g0508(.dina(w_G409gat_6[0]),.dinb(w_G69gat_4[2]),.dout(n572),.clk(gclk));
	jnot g0509(.din(n572),.dout(n573),.clk(gclk));
	jand g0510(.dina(w_n538_0[0]),.dinb(w_n497_0[0]),.dout(n574),.clk(gclk));
	jand g0511(.dina(w_n539_0[0]),.dinb(w_n494_0[0]),.dout(n575),.clk(gclk));
	jor g0512(.dina(n575),.dinb(w_dff_B_WMEeveX70_1),.dout(n576),.clk(gclk));
	jand g0513(.dina(w_G392gat_5[2]),.dinb(w_G86gat_5[0]),.dout(n577),.clk(gclk));
	jnot g0514(.din(n577),.dout(n578),.clk(gclk));
	jand g0515(.dina(w_n536_0[0]),.dinb(w_n502_0[0]),.dout(n579),.clk(gclk));
	jand g0516(.dina(w_n537_0[0]),.dinb(w_n499_0[0]),.dout(n580),.clk(gclk));
	jor g0517(.dina(n580),.dinb(w_dff_B_s9Cd84hT8_1),.dout(n581),.clk(gclk));
	jand g0518(.dina(w_G375gat_5[1]),.dinb(w_G103gat_5[1]),.dout(n582),.clk(gclk));
	jnot g0519(.din(n582),.dout(n583),.clk(gclk));
	jand g0520(.dina(w_n534_0[0]),.dinb(w_n507_0[0]),.dout(n584),.clk(gclk));
	jand g0521(.dina(w_n535_0[0]),.dinb(w_n504_0[0]),.dout(n585),.clk(gclk));
	jor g0522(.dina(n585),.dinb(w_dff_B_1jkOuCTe1_1),.dout(n586),.clk(gclk));
	jand g0523(.dina(w_G358gat_5[0]),.dinb(w_G120gat_5[2]),.dout(n587),.clk(gclk));
	jnot g0524(.din(n587),.dout(n588),.clk(gclk));
	jand g0525(.dina(w_n532_0[0]),.dinb(w_n512_0[0]),.dout(n589),.clk(gclk));
	jand g0526(.dina(w_n533_0[0]),.dinb(w_n509_0[0]),.dout(n590),.clk(gclk));
	jor g0527(.dina(n590),.dinb(w_dff_B_JXDGhtOe4_1),.dout(n591),.clk(gclk));
	jand g0528(.dina(w_G341gat_4[2]),.dinb(w_G137gat_6[0]),.dout(n592),.clk(gclk));
	jnot g0529(.din(n592),.dout(n593),.clk(gclk));
	jand g0530(.dina(w_n530_0[0]),.dinb(w_n518_0[0]),.dout(n594),.clk(gclk));
	jand g0531(.dina(w_n531_0[0]),.dinb(w_n514_0[0]),.dout(n595),.clk(gclk));
	jor g0532(.dina(n595),.dinb(w_dff_B_rAYAdfFl2_1),.dout(n596),.clk(gclk));
	jand g0533(.dina(w_G324gat_4[1]),.dinb(w_G154gat_6[1]),.dout(n597),.clk(gclk));
	jnot g0534(.din(n597),.dout(n598),.clk(gclk));
	jnot g0535(.din(w_n519_0[0]),.dout(n599),.clk(gclk));
	jnot g0536(.din(w_n529_0[0]),.dout(n600),.clk(gclk));
	jand g0537(.dina(n600),.dinb(w_dff_B_CbMh0etk8_1),.dout(n601),.clk(gclk));
	jor g0538(.dina(n601),.dinb(w_n527_0[0]),.dout(n602),.clk(gclk));
	jand g0539(.dina(w_G307gat_4[1]),.dinb(w_G171gat_6[2]),.dout(n603),.clk(gclk));
	jand g0540(.dina(w_G273gat_3[1]),.dinb(w_G205gat_7[1]),.dout(n604),.clk(gclk));
	jor g0541(.dina(w_n604_0[1]),.dinb(w_n522_0[0]),.dout(n605),.clk(gclk));
	jand g0542(.dina(w_G290gat_3[1]),.dinb(w_G205gat_7[0]),.dout(n606),.clk(gclk));
	jand g0543(.dina(w_n606_0[1]),.dinb(w_n520_0[0]),.dout(n607),.clk(gclk));
	jnot g0544(.din(w_n607_0[2]),.dout(n608),.clk(gclk));
	jand g0545(.dina(w_n608_0[1]),.dinb(w_dff_B_wtlWOni45_1),.dout(n609),.clk(gclk));
	jor g0546(.dina(n609),.dinb(w_n523_0[1]),.dout(n610),.clk(gclk));
	jnot g0547(.din(n610),.dout(n611),.clk(gclk));
	jand g0548(.dina(w_n608_0[0]),.dinb(w_n523_0[0]),.dout(n612),.clk(gclk));
	jor g0549(.dina(w_dff_B_yeWItqQb4_0),.dinb(w_n611_0[1]),.dout(n613),.clk(gclk));
	jxor g0550(.dina(w_n613_0[1]),.dinb(w_n603_0[1]),.dout(n614),.clk(gclk));
	jxor g0551(.dina(w_n614_0[1]),.dinb(w_n602_0[1]),.dout(n615),.clk(gclk));
	jxor g0552(.dina(w_n615_0[1]),.dinb(w_n598_0[1]),.dout(n616),.clk(gclk));
	jxor g0553(.dina(w_n616_0[1]),.dinb(w_n596_0[1]),.dout(n617),.clk(gclk));
	jxor g0554(.dina(w_n617_0[1]),.dinb(w_n593_0[1]),.dout(n618),.clk(gclk));
	jxor g0555(.dina(w_n618_0[1]),.dinb(w_n591_0[1]),.dout(n619),.clk(gclk));
	jxor g0556(.dina(w_n619_0[1]),.dinb(w_n588_0[1]),.dout(n620),.clk(gclk));
	jxor g0557(.dina(w_n620_0[1]),.dinb(w_n586_0[1]),.dout(n621),.clk(gclk));
	jxor g0558(.dina(w_n621_0[1]),.dinb(w_n583_0[1]),.dout(n622),.clk(gclk));
	jxor g0559(.dina(w_n622_0[1]),.dinb(w_n581_0[1]),.dout(n623),.clk(gclk));
	jxor g0560(.dina(w_n623_0[1]),.dinb(w_n578_0[1]),.dout(n624),.clk(gclk));
	jxor g0561(.dina(w_n624_0[1]),.dinb(w_n576_0[1]),.dout(n625),.clk(gclk));
	jxor g0562(.dina(w_n625_0[1]),.dinb(w_n573_0[1]),.dout(n626),.clk(gclk));
	jxor g0563(.dina(w_n626_0[1]),.dinb(w_n571_0[1]),.dout(n627),.clk(gclk));
	jxor g0564(.dina(w_n627_0[1]),.dinb(w_n568_0[1]),.dout(n628),.clk(gclk));
	jxor g0565(.dina(w_n628_0[1]),.dinb(w_n566_0[1]),.dout(n629),.clk(gclk));
	jxor g0566(.dina(w_n629_0[1]),.dinb(w_n563_0[1]),.dout(n630),.clk(gclk));
	jnot g0567(.din(w_n630_0[1]),.dout(n631),.clk(gclk));
	jxor g0568(.dina(w_n631_0[1]),.dinb(w_n561_0[2]),.dout(n632),.clk(gclk));
	jxor g0569(.dina(n632),.dinb(w_dff_B_fSmRDmHs5_1),.dout(n633),.clk(gclk));
	jxor g0570(.dina(w_n633_0[1]),.dinb(w_n555_0[1]),.dout(n634),.clk(gclk));
	jxor g0571(.dina(w_n634_0[1]),.dinb(w_dff_B_I9nJ9Bc26_1),.dout(w_dff_A_7vyaZLbT9_2),.clk(gclk));
	jand g0572(.dina(w_G494gat_7[1]),.dinb(w_G1gat_3[0]),.dout(n636),.clk(gclk));
	jnot g0573(.din(w_n636_0[1]),.dout(n637),.clk(gclk));
	jnot g0574(.din(w_n633_0[0]),.dout(n638),.clk(gclk));
	jor g0575(.dina(n638),.dinb(w_n555_0[0]),.dout(n639),.clk(gclk));
	jor g0576(.dina(w_n634_0[0]),.dinb(w_n550_0[0]),.dout(n640),.clk(gclk));
	jand g0577(.dina(n640),.dinb(w_dff_B_ycRlJSps1_1),.dout(n641),.clk(gclk));
	jand g0578(.dina(w_G477gat_7[0]),.dinb(w_G18gat_3[1]),.dout(n642),.clk(gclk));
	jnot g0579(.din(w_n642_0[1]),.dout(n643),.clk(gclk));
	jor g0580(.dina(w_n631_0[0]),.dinb(w_n561_0[1]),.dout(n644),.clk(gclk));
	jxor g0581(.dina(w_n630_0[0]),.dinb(w_n561_0[0]),.dout(n645),.clk(gclk));
	jor g0582(.dina(n645),.dinb(w_n556_0[0]),.dout(n646),.clk(gclk));
	jand g0583(.dina(n646),.dinb(w_dff_B_T0JlXUcf3_1),.dout(n647),.clk(gclk));
	jand g0584(.dina(w_G460gat_6[2]),.dinb(w_G35gat_3[2]),.dout(n648),.clk(gclk));
	jnot g0585(.din(n648),.dout(n649),.clk(gclk));
	jand g0586(.dina(w_n628_0[0]),.dinb(w_n566_0[0]),.dout(n650),.clk(gclk));
	jand g0587(.dina(w_n629_0[0]),.dinb(w_n563_0[0]),.dout(n651),.clk(gclk));
	jor g0588(.dina(n651),.dinb(w_dff_B_p7A5tY8K4_1),.dout(n652),.clk(gclk));
	jand g0589(.dina(w_G443gat_6[1]),.dinb(w_G52gat_4[0]),.dout(n653),.clk(gclk));
	jnot g0590(.din(n653),.dout(n654),.clk(gclk));
	jand g0591(.dina(w_n626_0[0]),.dinb(w_n571_0[0]),.dout(n655),.clk(gclk));
	jand g0592(.dina(w_n627_0[0]),.dinb(w_n568_0[0]),.dout(n656),.clk(gclk));
	jor g0593(.dina(n656),.dinb(w_dff_B_yk77LfyS1_1),.dout(n657),.clk(gclk));
	jand g0594(.dina(w_G426gat_6[0]),.dinb(w_G69gat_4[1]),.dout(n658),.clk(gclk));
	jnot g0595(.din(n658),.dout(n659),.clk(gclk));
	jand g0596(.dina(w_n624_0[0]),.dinb(w_n576_0[0]),.dout(n660),.clk(gclk));
	jand g0597(.dina(w_n625_0[0]),.dinb(w_n573_0[0]),.dout(n661),.clk(gclk));
	jor g0598(.dina(n661),.dinb(w_dff_B_ygjs60Th7_1),.dout(n662),.clk(gclk));
	jand g0599(.dina(w_G409gat_5[2]),.dinb(w_G86gat_4[2]),.dout(n663),.clk(gclk));
	jnot g0600(.din(n663),.dout(n664),.clk(gclk));
	jand g0601(.dina(w_n622_0[0]),.dinb(w_n581_0[0]),.dout(n665),.clk(gclk));
	jand g0602(.dina(w_n623_0[0]),.dinb(w_n578_0[0]),.dout(n666),.clk(gclk));
	jor g0603(.dina(n666),.dinb(w_dff_B_9M5pmyQ40_1),.dout(n667),.clk(gclk));
	jand g0604(.dina(w_G392gat_5[1]),.dinb(w_G103gat_5[0]),.dout(n668),.clk(gclk));
	jnot g0605(.din(n668),.dout(n669),.clk(gclk));
	jand g0606(.dina(w_n620_0[0]),.dinb(w_n586_0[0]),.dout(n670),.clk(gclk));
	jand g0607(.dina(w_n621_0[0]),.dinb(w_n583_0[0]),.dout(n671),.clk(gclk));
	jor g0608(.dina(n671),.dinb(w_dff_B_mW1TSD8L4_1),.dout(n672),.clk(gclk));
	jand g0609(.dina(w_G375gat_5[0]),.dinb(w_G120gat_5[1]),.dout(n673),.clk(gclk));
	jnot g0610(.din(n673),.dout(n674),.clk(gclk));
	jand g0611(.dina(w_n618_0[0]),.dinb(w_n591_0[0]),.dout(n675),.clk(gclk));
	jand g0612(.dina(w_n619_0[0]),.dinb(w_n588_0[0]),.dout(n676),.clk(gclk));
	jor g0613(.dina(n676),.dinb(w_dff_B_myZc1rch3_1),.dout(n677),.clk(gclk));
	jand g0614(.dina(w_G358gat_4[2]),.dinb(w_G137gat_5[2]),.dout(n678),.clk(gclk));
	jnot g0615(.din(n678),.dout(n679),.clk(gclk));
	jand g0616(.dina(w_n616_0[0]),.dinb(w_n596_0[0]),.dout(n680),.clk(gclk));
	jand g0617(.dina(w_n617_0[0]),.dinb(w_n593_0[0]),.dout(n681),.clk(gclk));
	jor g0618(.dina(n681),.dinb(w_dff_B_6qB0P92B1_1),.dout(n682),.clk(gclk));
	jand g0619(.dina(w_G341gat_4[1]),.dinb(w_G154gat_6[0]),.dout(n683),.clk(gclk));
	jnot g0620(.din(n683),.dout(n684),.clk(gclk));
	jand g0621(.dina(w_n614_0[0]),.dinb(w_n602_0[0]),.dout(n685),.clk(gclk));
	jand g0622(.dina(w_n615_0[0]),.dinb(w_n598_0[0]),.dout(n686),.clk(gclk));
	jor g0623(.dina(n686),.dinb(w_dff_B_vavzs6245_1),.dout(n687),.clk(gclk));
	jand g0624(.dina(w_G324gat_4[0]),.dinb(w_G171gat_6[1]),.dout(n688),.clk(gclk));
	jnot g0625(.din(n688),.dout(n689),.clk(gclk));
	jnot g0626(.din(w_n603_0[0]),.dout(n690),.clk(gclk));
	jnot g0627(.din(w_n613_0[0]),.dout(n691),.clk(gclk));
	jand g0628(.dina(n691),.dinb(w_dff_B_w4rI4dlB8_1),.dout(n692),.clk(gclk));
	jor g0629(.dina(n692),.dinb(w_n611_0[0]),.dout(n693),.clk(gclk));
	jand g0630(.dina(w_G307gat_4[0]),.dinb(w_G188gat_6[2]),.dout(n694),.clk(gclk));
	jand g0631(.dina(w_G273gat_3[0]),.dinb(w_G222gat_7[1]),.dout(n695),.clk(gclk));
	jor g0632(.dina(w_n695_0[2]),.dinb(w_n606_0[0]),.dout(n696),.clk(gclk));
	jand g0633(.dina(w_G290gat_3[0]),.dinb(w_G222gat_7[0]),.dout(n697),.clk(gclk));
	jand g0634(.dina(w_n697_0[1]),.dinb(w_n604_0[0]),.dout(n698),.clk(gclk));
	jnot g0635(.din(w_n698_0[2]),.dout(n699),.clk(gclk));
	jand g0636(.dina(w_n699_0[1]),.dinb(w_dff_B_j6eUikvB2_1),.dout(n700),.clk(gclk));
	jor g0637(.dina(n700),.dinb(w_n607_0[1]),.dout(n701),.clk(gclk));
	jnot g0638(.din(n701),.dout(n702),.clk(gclk));
	jand g0639(.dina(w_n699_0[0]),.dinb(w_n607_0[0]),.dout(n703),.clk(gclk));
	jor g0640(.dina(w_dff_B_PYhFfXDa8_0),.dinb(w_n702_0[1]),.dout(n704),.clk(gclk));
	jxor g0641(.dina(w_n704_0[1]),.dinb(w_n694_0[1]),.dout(n705),.clk(gclk));
	jxor g0642(.dina(w_n705_0[1]),.dinb(w_n693_0[1]),.dout(n706),.clk(gclk));
	jxor g0643(.dina(w_n706_0[1]),.dinb(w_n689_0[1]),.dout(n707),.clk(gclk));
	jxor g0644(.dina(w_n707_0[1]),.dinb(w_n687_0[1]),.dout(n708),.clk(gclk));
	jxor g0645(.dina(w_n708_0[1]),.dinb(w_n684_0[1]),.dout(n709),.clk(gclk));
	jxor g0646(.dina(w_n709_0[1]),.dinb(w_n682_0[1]),.dout(n710),.clk(gclk));
	jxor g0647(.dina(w_n710_0[1]),.dinb(w_n679_0[1]),.dout(n711),.clk(gclk));
	jxor g0648(.dina(w_n711_0[1]),.dinb(w_n677_0[1]),.dout(n712),.clk(gclk));
	jxor g0649(.dina(w_n712_0[1]),.dinb(w_n674_0[1]),.dout(n713),.clk(gclk));
	jxor g0650(.dina(w_n713_0[1]),.dinb(w_n672_0[1]),.dout(n714),.clk(gclk));
	jxor g0651(.dina(w_n714_0[1]),.dinb(w_n669_0[1]),.dout(n715),.clk(gclk));
	jxor g0652(.dina(w_n715_0[1]),.dinb(w_n667_0[1]),.dout(n716),.clk(gclk));
	jxor g0653(.dina(w_n716_0[1]),.dinb(w_n664_0[1]),.dout(n717),.clk(gclk));
	jxor g0654(.dina(w_n717_0[1]),.dinb(w_n662_0[1]),.dout(n718),.clk(gclk));
	jxor g0655(.dina(w_n718_0[1]),.dinb(w_n659_0[1]),.dout(n719),.clk(gclk));
	jxor g0656(.dina(w_n719_0[1]),.dinb(w_n657_0[1]),.dout(n720),.clk(gclk));
	jxor g0657(.dina(w_n720_0[1]),.dinb(w_n654_0[1]),.dout(n721),.clk(gclk));
	jxor g0658(.dina(w_n721_0[1]),.dinb(w_n652_0[1]),.dout(n722),.clk(gclk));
	jxor g0659(.dina(w_n722_0[1]),.dinb(w_n649_0[1]),.dout(n723),.clk(gclk));
	jnot g0660(.din(w_n723_0[1]),.dout(n724),.clk(gclk));
	jxor g0661(.dina(w_n724_0[1]),.dinb(w_n647_0[2]),.dout(n725),.clk(gclk));
	jxor g0662(.dina(n725),.dinb(w_dff_B_gR0O5Ao48_1),.dout(n726),.clk(gclk));
	jxor g0663(.dina(w_n726_0[1]),.dinb(w_n641_0[1]),.dout(n727),.clk(gclk));
	jxor g0664(.dina(w_n727_0[1]),.dinb(w_dff_B_fX6XFwfv2_1),.dout(w_dff_A_TEKx8qT56_2),.clk(gclk));
	jand g0665(.dina(w_G511gat_7[1]),.dinb(w_G1gat_2[2]),.dout(n729),.clk(gclk));
	jnot g0666(.din(w_n729_0[1]),.dout(n730),.clk(gclk));
	jnot g0667(.din(w_n726_0[0]),.dout(n731),.clk(gclk));
	jor g0668(.dina(n731),.dinb(w_n641_0[0]),.dout(n732),.clk(gclk));
	jor g0669(.dina(w_n727_0[0]),.dinb(w_n636_0[0]),.dout(n733),.clk(gclk));
	jand g0670(.dina(n733),.dinb(w_dff_B_XehIwMva3_1),.dout(n734),.clk(gclk));
	jand g0671(.dina(w_G494gat_7[0]),.dinb(w_G18gat_3[0]),.dout(n735),.clk(gclk));
	jnot g0672(.din(w_n735_0[1]),.dout(n736),.clk(gclk));
	jor g0673(.dina(w_n724_0[0]),.dinb(w_n647_0[1]),.dout(n737),.clk(gclk));
	jxor g0674(.dina(w_n723_0[0]),.dinb(w_n647_0[0]),.dout(n738),.clk(gclk));
	jor g0675(.dina(n738),.dinb(w_n642_0[0]),.dout(n739),.clk(gclk));
	jand g0676(.dina(n739),.dinb(w_dff_B_n1qofQ7N6_1),.dout(n740),.clk(gclk));
	jand g0677(.dina(w_G477gat_6[2]),.dinb(w_G35gat_3[1]),.dout(n741),.clk(gclk));
	jnot g0678(.din(n741),.dout(n742),.clk(gclk));
	jand g0679(.dina(w_n721_0[0]),.dinb(w_n652_0[0]),.dout(n743),.clk(gclk));
	jand g0680(.dina(w_n722_0[0]),.dinb(w_n649_0[0]),.dout(n744),.clk(gclk));
	jor g0681(.dina(n744),.dinb(w_dff_B_YFGLmNff5_1),.dout(n745),.clk(gclk));
	jand g0682(.dina(w_G460gat_6[1]),.dinb(w_G52gat_3[2]),.dout(n746),.clk(gclk));
	jnot g0683(.din(n746),.dout(n747),.clk(gclk));
	jand g0684(.dina(w_n719_0[0]),.dinb(w_n657_0[0]),.dout(n748),.clk(gclk));
	jand g0685(.dina(w_n720_0[0]),.dinb(w_n654_0[0]),.dout(n749),.clk(gclk));
	jor g0686(.dina(n749),.dinb(w_dff_B_BJRhwV3R5_1),.dout(n750),.clk(gclk));
	jand g0687(.dina(w_G443gat_6[0]),.dinb(w_G69gat_4[0]),.dout(n751),.clk(gclk));
	jnot g0688(.din(n751),.dout(n752),.clk(gclk));
	jand g0689(.dina(w_n717_0[0]),.dinb(w_n662_0[0]),.dout(n753),.clk(gclk));
	jand g0690(.dina(w_n718_0[0]),.dinb(w_n659_0[0]),.dout(n754),.clk(gclk));
	jor g0691(.dina(n754),.dinb(w_dff_B_mxcrFEy75_1),.dout(n755),.clk(gclk));
	jand g0692(.dina(w_G426gat_5[2]),.dinb(w_G86gat_4[1]),.dout(n756),.clk(gclk));
	jnot g0693(.din(n756),.dout(n757),.clk(gclk));
	jand g0694(.dina(w_n715_0[0]),.dinb(w_n667_0[0]),.dout(n758),.clk(gclk));
	jand g0695(.dina(w_n716_0[0]),.dinb(w_n664_0[0]),.dout(n759),.clk(gclk));
	jor g0696(.dina(n759),.dinb(w_dff_B_F4vP9F4i6_1),.dout(n760),.clk(gclk));
	jand g0697(.dina(w_G409gat_5[1]),.dinb(w_G103gat_4[2]),.dout(n761),.clk(gclk));
	jnot g0698(.din(n761),.dout(n762),.clk(gclk));
	jand g0699(.dina(w_n713_0[0]),.dinb(w_n672_0[0]),.dout(n763),.clk(gclk));
	jand g0700(.dina(w_n714_0[0]),.dinb(w_n669_0[0]),.dout(n764),.clk(gclk));
	jor g0701(.dina(n764),.dinb(w_dff_B_j9Ffr4DS0_1),.dout(n765),.clk(gclk));
	jand g0702(.dina(w_G392gat_5[0]),.dinb(w_G120gat_5[0]),.dout(n766),.clk(gclk));
	jnot g0703(.din(n766),.dout(n767),.clk(gclk));
	jand g0704(.dina(w_n711_0[0]),.dinb(w_n677_0[0]),.dout(n768),.clk(gclk));
	jand g0705(.dina(w_n712_0[0]),.dinb(w_n674_0[0]),.dout(n769),.clk(gclk));
	jor g0706(.dina(n769),.dinb(w_dff_B_aLCONApw9_1),.dout(n770),.clk(gclk));
	jand g0707(.dina(w_G375gat_4[2]),.dinb(w_G137gat_5[1]),.dout(n771),.clk(gclk));
	jnot g0708(.din(n771),.dout(n772),.clk(gclk));
	jand g0709(.dina(w_n709_0[0]),.dinb(w_n682_0[0]),.dout(n773),.clk(gclk));
	jand g0710(.dina(w_n710_0[0]),.dinb(w_n679_0[0]),.dout(n774),.clk(gclk));
	jor g0711(.dina(n774),.dinb(w_dff_B_gkIHDYrP0_1),.dout(n775),.clk(gclk));
	jand g0712(.dina(w_G358gat_4[1]),.dinb(w_G154gat_5[2]),.dout(n776),.clk(gclk));
	jnot g0713(.din(n776),.dout(n777),.clk(gclk));
	jand g0714(.dina(w_n707_0[0]),.dinb(w_n687_0[0]),.dout(n778),.clk(gclk));
	jand g0715(.dina(w_n708_0[0]),.dinb(w_n684_0[0]),.dout(n779),.clk(gclk));
	jor g0716(.dina(n779),.dinb(w_dff_B_bSQO3Iix9_1),.dout(n780),.clk(gclk));
	jand g0717(.dina(w_G341gat_4[0]),.dinb(w_G171gat_6[0]),.dout(n781),.clk(gclk));
	jnot g0718(.din(n781),.dout(n782),.clk(gclk));
	jand g0719(.dina(w_n705_0[0]),.dinb(w_n693_0[0]),.dout(n783),.clk(gclk));
	jand g0720(.dina(w_n706_0[0]),.dinb(w_n689_0[0]),.dout(n784),.clk(gclk));
	jor g0721(.dina(n784),.dinb(w_dff_B_R12el6iH1_1),.dout(n785),.clk(gclk));
	jand g0722(.dina(w_G324gat_3[2]),.dinb(w_G188gat_6[1]),.dout(n786),.clk(gclk));
	jnot g0723(.din(n786),.dout(n787),.clk(gclk));
	jnot g0724(.din(w_n694_0[0]),.dout(n788),.clk(gclk));
	jnot g0725(.din(w_n704_0[0]),.dout(n789),.clk(gclk));
	jand g0726(.dina(n789),.dinb(w_dff_B_ycQziHRj5_1),.dout(n790),.clk(gclk));
	jor g0727(.dina(n790),.dinb(w_n702_0[0]),.dout(n791),.clk(gclk));
	jand g0728(.dina(w_G307gat_3[2]),.dinb(w_G205gat_6[2]),.dout(n792),.clk(gclk));
	jand g0729(.dina(w_G273gat_2[2]),.dinb(w_G239gat_7[1]),.dout(n793),.clk(gclk));
	jor g0730(.dina(w_n793_0[1]),.dinb(w_n697_0[0]),.dout(n794),.clk(gclk));
	jand g0731(.dina(w_G290gat_2[2]),.dinb(w_G239gat_7[0]),.dout(n795),.clk(gclk));
	jand g0732(.dina(w_n795_0[1]),.dinb(w_n695_0[1]),.dout(n796),.clk(gclk));
	jnot g0733(.din(n796),.dout(n797),.clk(gclk));
	jand g0734(.dina(w_n797_0[2]),.dinb(w_dff_B_fexZ1vyZ4_1),.dout(n798),.clk(gclk));
	jor g0735(.dina(n798),.dinb(w_n698_0[1]),.dout(n799),.clk(gclk));
	jnot g0736(.din(n799),.dout(n800),.clk(gclk));
	jand g0737(.dina(w_n797_0[1]),.dinb(w_n698_0[0]),.dout(n801),.clk(gclk));
	jor g0738(.dina(w_dff_B_l1FIUshX7_0),.dinb(w_n800_0[1]),.dout(n802),.clk(gclk));
	jxor g0739(.dina(w_n802_0[1]),.dinb(w_n792_0[1]),.dout(n803),.clk(gclk));
	jxor g0740(.dina(w_n803_0[1]),.dinb(w_n791_0[1]),.dout(n804),.clk(gclk));
	jxor g0741(.dina(w_n804_0[1]),.dinb(w_n787_0[1]),.dout(n805),.clk(gclk));
	jxor g0742(.dina(w_n805_0[1]),.dinb(w_n785_0[1]),.dout(n806),.clk(gclk));
	jxor g0743(.dina(w_n806_0[1]),.dinb(w_n782_0[1]),.dout(n807),.clk(gclk));
	jxor g0744(.dina(w_n807_0[1]),.dinb(w_n780_0[1]),.dout(n808),.clk(gclk));
	jxor g0745(.dina(w_n808_0[1]),.dinb(w_n777_0[1]),.dout(n809),.clk(gclk));
	jxor g0746(.dina(w_n809_0[1]),.dinb(w_n775_0[1]),.dout(n810),.clk(gclk));
	jxor g0747(.dina(w_n810_0[1]),.dinb(w_n772_0[1]),.dout(n811),.clk(gclk));
	jxor g0748(.dina(w_n811_0[1]),.dinb(w_n770_0[1]),.dout(n812),.clk(gclk));
	jxor g0749(.dina(w_n812_0[1]),.dinb(w_n767_0[1]),.dout(n813),.clk(gclk));
	jxor g0750(.dina(w_n813_0[1]),.dinb(w_n765_0[1]),.dout(n814),.clk(gclk));
	jxor g0751(.dina(w_n814_0[1]),.dinb(w_n762_0[1]),.dout(n815),.clk(gclk));
	jxor g0752(.dina(w_n815_0[1]),.dinb(w_n760_0[1]),.dout(n816),.clk(gclk));
	jxor g0753(.dina(w_n816_0[1]),.dinb(w_n757_0[1]),.dout(n817),.clk(gclk));
	jxor g0754(.dina(w_n817_0[1]),.dinb(w_n755_0[1]),.dout(n818),.clk(gclk));
	jxor g0755(.dina(w_n818_0[1]),.dinb(w_n752_0[1]),.dout(n819),.clk(gclk));
	jxor g0756(.dina(w_n819_0[1]),.dinb(w_n750_0[1]),.dout(n820),.clk(gclk));
	jxor g0757(.dina(w_n820_0[1]),.dinb(w_n747_0[1]),.dout(n821),.clk(gclk));
	jxor g0758(.dina(w_n821_0[1]),.dinb(w_n745_0[1]),.dout(n822),.clk(gclk));
	jxor g0759(.dina(w_n822_0[1]),.dinb(w_n742_0[1]),.dout(n823),.clk(gclk));
	jnot g0760(.din(w_n823_0[1]),.dout(n824),.clk(gclk));
	jxor g0761(.dina(w_n824_0[1]),.dinb(w_n740_0[2]),.dout(n825),.clk(gclk));
	jxor g0762(.dina(n825),.dinb(w_dff_B_6piPLQWx6_1),.dout(n826),.clk(gclk));
	jxor g0763(.dina(w_n826_0[1]),.dinb(w_n734_0[1]),.dout(n827),.clk(gclk));
	jxor g0764(.dina(w_n827_0[1]),.dinb(w_dff_B_P2cfAhMG6_1),.dout(w_dff_A_ND5rrPHV5_2),.clk(gclk));
	jand g0765(.dina(w_G528gat_7[1]),.dinb(w_G1gat_2[1]),.dout(n829),.clk(gclk));
	jnot g0766(.din(w_n829_0[1]),.dout(n830),.clk(gclk));
	jnot g0767(.din(w_n826_0[0]),.dout(n831),.clk(gclk));
	jor g0768(.dina(n831),.dinb(w_n734_0[0]),.dout(n832),.clk(gclk));
	jor g0769(.dina(w_n827_0[0]),.dinb(w_n729_0[0]),.dout(n833),.clk(gclk));
	jand g0770(.dina(n833),.dinb(w_dff_B_cm5qEtPD6_1),.dout(n834),.clk(gclk));
	jand g0771(.dina(w_G511gat_7[0]),.dinb(w_G18gat_2[2]),.dout(n835),.clk(gclk));
	jor g0772(.dina(w_n824_0[0]),.dinb(w_n740_0[1]),.dout(n836),.clk(gclk));
	jxor g0773(.dina(w_n823_0[0]),.dinb(w_n740_0[0]),.dout(n837),.clk(gclk));
	jor g0774(.dina(n837),.dinb(w_n735_0[0]),.dout(n838),.clk(gclk));
	jand g0775(.dina(n838),.dinb(w_dff_B_KpqY4Roc0_1),.dout(n839),.clk(gclk));
	jand g0776(.dina(w_G494gat_6[2]),.dinb(w_G35gat_3[0]),.dout(n840),.clk(gclk));
	jnot g0777(.din(w_n840_0[1]),.dout(n841),.clk(gclk));
	jand g0778(.dina(w_n821_0[0]),.dinb(w_n745_0[0]),.dout(n842),.clk(gclk));
	jand g0779(.dina(w_n822_0[0]),.dinb(w_n742_0[0]),.dout(n843),.clk(gclk));
	jor g0780(.dina(n843),.dinb(w_dff_B_pFzgrlqQ6_1),.dout(n844),.clk(gclk));
	jand g0781(.dina(w_G477gat_6[1]),.dinb(w_G52gat_3[1]),.dout(n845),.clk(gclk));
	jnot g0782(.din(n845),.dout(n846),.clk(gclk));
	jand g0783(.dina(w_n819_0[0]),.dinb(w_n750_0[0]),.dout(n847),.clk(gclk));
	jand g0784(.dina(w_n820_0[0]),.dinb(w_n747_0[0]),.dout(n848),.clk(gclk));
	jor g0785(.dina(n848),.dinb(w_dff_B_pkXP9ILj6_1),.dout(n849),.clk(gclk));
	jand g0786(.dina(w_G460gat_6[0]),.dinb(w_G69gat_3[2]),.dout(n850),.clk(gclk));
	jnot g0787(.din(n850),.dout(n851),.clk(gclk));
	jand g0788(.dina(w_n817_0[0]),.dinb(w_n755_0[0]),.dout(n852),.clk(gclk));
	jand g0789(.dina(w_n818_0[0]),.dinb(w_n752_0[0]),.dout(n853),.clk(gclk));
	jor g0790(.dina(n853),.dinb(w_dff_B_fWUgkO5b0_1),.dout(n854),.clk(gclk));
	jand g0791(.dina(w_G443gat_5[2]),.dinb(w_G86gat_4[0]),.dout(n855),.clk(gclk));
	jnot g0792(.din(n855),.dout(n856),.clk(gclk));
	jand g0793(.dina(w_n815_0[0]),.dinb(w_n760_0[0]),.dout(n857),.clk(gclk));
	jand g0794(.dina(w_n816_0[0]),.dinb(w_n757_0[0]),.dout(n858),.clk(gclk));
	jor g0795(.dina(n858),.dinb(w_dff_B_aOKnKsbI5_1),.dout(n859),.clk(gclk));
	jand g0796(.dina(w_G426gat_5[1]),.dinb(w_G103gat_4[1]),.dout(n860),.clk(gclk));
	jnot g0797(.din(n860),.dout(n861),.clk(gclk));
	jand g0798(.dina(w_n813_0[0]),.dinb(w_n765_0[0]),.dout(n862),.clk(gclk));
	jand g0799(.dina(w_n814_0[0]),.dinb(w_n762_0[0]),.dout(n863),.clk(gclk));
	jor g0800(.dina(n863),.dinb(w_dff_B_QYADrKf36_1),.dout(n864),.clk(gclk));
	jand g0801(.dina(w_G409gat_5[0]),.dinb(w_G120gat_4[2]),.dout(n865),.clk(gclk));
	jnot g0802(.din(n865),.dout(n866),.clk(gclk));
	jand g0803(.dina(w_n811_0[0]),.dinb(w_n770_0[0]),.dout(n867),.clk(gclk));
	jand g0804(.dina(w_n812_0[0]),.dinb(w_n767_0[0]),.dout(n868),.clk(gclk));
	jor g0805(.dina(n868),.dinb(w_dff_B_FwUjwLpg3_1),.dout(n869),.clk(gclk));
	jand g0806(.dina(w_G392gat_4[2]),.dinb(w_G137gat_5[0]),.dout(n870),.clk(gclk));
	jnot g0807(.din(n870),.dout(n871),.clk(gclk));
	jand g0808(.dina(w_n809_0[0]),.dinb(w_n775_0[0]),.dout(n872),.clk(gclk));
	jand g0809(.dina(w_n810_0[0]),.dinb(w_n772_0[0]),.dout(n873),.clk(gclk));
	jor g0810(.dina(n873),.dinb(w_dff_B_c8K0u9p28_1),.dout(n874),.clk(gclk));
	jand g0811(.dina(w_G375gat_4[1]),.dinb(w_G154gat_5[1]),.dout(n875),.clk(gclk));
	jnot g0812(.din(n875),.dout(n876),.clk(gclk));
	jand g0813(.dina(w_n807_0[0]),.dinb(w_n780_0[0]),.dout(n877),.clk(gclk));
	jand g0814(.dina(w_n808_0[0]),.dinb(w_n777_0[0]),.dout(n878),.clk(gclk));
	jor g0815(.dina(n878),.dinb(w_dff_B_HJQyML745_1),.dout(n879),.clk(gclk));
	jand g0816(.dina(w_G358gat_4[0]),.dinb(w_G171gat_5[2]),.dout(n880),.clk(gclk));
	jnot g0817(.din(n880),.dout(n881),.clk(gclk));
	jand g0818(.dina(w_n805_0[0]),.dinb(w_n785_0[0]),.dout(n882),.clk(gclk));
	jand g0819(.dina(w_n806_0[0]),.dinb(w_n782_0[0]),.dout(n883),.clk(gclk));
	jor g0820(.dina(n883),.dinb(w_dff_B_6TftSVYF7_1),.dout(n884),.clk(gclk));
	jand g0821(.dina(w_G341gat_3[2]),.dinb(w_G188gat_6[0]),.dout(n885),.clk(gclk));
	jnot g0822(.din(n885),.dout(n886),.clk(gclk));
	jand g0823(.dina(w_n803_0[0]),.dinb(w_n791_0[0]),.dout(n887),.clk(gclk));
	jand g0824(.dina(w_n804_0[0]),.dinb(w_n787_0[0]),.dout(n888),.clk(gclk));
	jor g0825(.dina(n888),.dinb(w_dff_B_UNbWXrTi5_1),.dout(n889),.clk(gclk));
	jand g0826(.dina(w_G324gat_3[1]),.dinb(w_G205gat_6[1]),.dout(n890),.clk(gclk));
	jnot g0827(.din(n890),.dout(n891),.clk(gclk));
	jnot g0828(.din(w_n792_0[0]),.dout(n892),.clk(gclk));
	jnot g0829(.din(w_n802_0[0]),.dout(n893),.clk(gclk));
	jand g0830(.dina(n893),.dinb(w_dff_B_Q36U5tAt1_1),.dout(n894),.clk(gclk));
	jor g0831(.dina(n894),.dinb(w_n800_0[0]),.dout(n895),.clk(gclk));
	jand g0832(.dina(w_G307gat_3[1]),.dinb(w_G222gat_6[2]),.dout(n896),.clk(gclk));
	jnot g0833(.din(w_n795_0[0]),.dout(n897),.clk(gclk));
	jand g0834(.dina(w_G273gat_2[1]),.dinb(w_G256gat_7[1]),.dout(n898),.clk(gclk));
	jand g0835(.dina(w_n898_0[1]),.dinb(w_n897_0[1]),.dout(n899),.clk(gclk));
	jnot g0836(.din(n899),.dout(n900),.clk(gclk));
	jor g0837(.dina(w_n898_0[0]),.dinb(w_n897_0[0]),.dout(n901),.clk(gclk));
	jand g0838(.dina(w_n901_0[1]),.dinb(w_n797_0[0]),.dout(n902),.clk(gclk));
	jand g0839(.dina(n902),.dinb(n900),.dout(n903),.clk(gclk));
	jnot g0840(.din(w_n901_0[0]),.dout(n904),.clk(gclk));
	jand g0841(.dina(n904),.dinb(w_n695_0[0]),.dout(n905),.clk(gclk));
	jor g0842(.dina(n905),.dinb(w_n903_0[1]),.dout(n906),.clk(gclk));
	jxor g0843(.dina(w_n906_0[1]),.dinb(w_n896_0[1]),.dout(n907),.clk(gclk));
	jxor g0844(.dina(w_n907_0[1]),.dinb(w_n895_0[1]),.dout(n908),.clk(gclk));
	jxor g0845(.dina(w_n908_0[1]),.dinb(w_n891_0[1]),.dout(n909),.clk(gclk));
	jxor g0846(.dina(w_n909_0[1]),.dinb(w_n889_0[1]),.dout(n910),.clk(gclk));
	jxor g0847(.dina(w_n910_0[1]),.dinb(w_n886_0[1]),.dout(n911),.clk(gclk));
	jxor g0848(.dina(w_n911_0[1]),.dinb(w_n884_0[1]),.dout(n912),.clk(gclk));
	jxor g0849(.dina(w_n912_0[1]),.dinb(w_n881_0[1]),.dout(n913),.clk(gclk));
	jxor g0850(.dina(w_n913_0[1]),.dinb(w_n879_0[1]),.dout(n914),.clk(gclk));
	jxor g0851(.dina(w_n914_0[1]),.dinb(w_n876_0[1]),.dout(n915),.clk(gclk));
	jxor g0852(.dina(w_n915_0[1]),.dinb(w_n874_0[1]),.dout(n916),.clk(gclk));
	jxor g0853(.dina(w_n916_0[1]),.dinb(w_n871_0[1]),.dout(n917),.clk(gclk));
	jxor g0854(.dina(w_n917_0[1]),.dinb(w_n869_0[1]),.dout(n918),.clk(gclk));
	jxor g0855(.dina(w_n918_0[1]),.dinb(w_n866_0[1]),.dout(n919),.clk(gclk));
	jxor g0856(.dina(w_n919_0[1]),.dinb(w_n864_0[1]),.dout(n920),.clk(gclk));
	jxor g0857(.dina(w_n920_0[1]),.dinb(w_n861_0[1]),.dout(n921),.clk(gclk));
	jxor g0858(.dina(w_n921_0[1]),.dinb(w_n859_0[1]),.dout(n922),.clk(gclk));
	jxor g0859(.dina(w_n922_0[1]),.dinb(w_n856_0[1]),.dout(n923),.clk(gclk));
	jxor g0860(.dina(w_n923_0[1]),.dinb(w_n854_0[1]),.dout(n924),.clk(gclk));
	jxor g0861(.dina(w_n924_0[1]),.dinb(w_n851_0[1]),.dout(n925),.clk(gclk));
	jxor g0862(.dina(w_n925_0[1]),.dinb(w_n849_0[1]),.dout(n926),.clk(gclk));
	jxor g0863(.dina(w_n926_0[1]),.dinb(w_n846_0[1]),.dout(n927),.clk(gclk));
	jxor g0864(.dina(w_n927_0[2]),.dinb(w_n844_0[2]),.dout(n928),.clk(gclk));
	jxor g0865(.dina(n928),.dinb(w_dff_B_VV2MIwFT6_1),.dout(n929),.clk(gclk));
	jxor g0866(.dina(w_n929_0[1]),.dinb(w_n839_0[1]),.dout(n930),.clk(gclk));
	jxor g0867(.dina(w_n930_0[1]),.dinb(w_n835_0[1]),.dout(n931),.clk(gclk));
	jxor g0868(.dina(w_n931_0[1]),.dinb(w_n834_0[1]),.dout(n932),.clk(gclk));
	jxor g0869(.dina(w_n932_0[1]),.dinb(w_dff_B_vYOXfILh7_1),.dout(w_dff_A_NtHJwKOW4_2),.clk(gclk));
	jnot g0870(.din(w_n931_0[0]),.dout(n934),.clk(gclk));
	jor g0871(.dina(n934),.dinb(w_n834_0[0]),.dout(n935),.clk(gclk));
	jor g0872(.dina(w_n932_0[0]),.dinb(w_n829_0[0]),.dout(n936),.clk(gclk));
	jand g0873(.dina(n936),.dinb(w_dff_B_uKVEnDbQ2_1),.dout(n937),.clk(gclk));
	jand g0874(.dina(w_G528gat_7[0]),.dinb(w_G18gat_2[1]),.dout(n938),.clk(gclk));
	jnot g0875(.din(w_n929_0[0]),.dout(n939),.clk(gclk));
	jor g0876(.dina(n939),.dinb(w_n839_0[0]),.dout(n940),.clk(gclk));
	jor g0877(.dina(w_n930_0[0]),.dinb(w_n835_0[0]),.dout(n941),.clk(gclk));
	jand g0878(.dina(n941),.dinb(w_dff_B_YU9Fs9yY9_1),.dout(n942),.clk(gclk));
	jand g0879(.dina(w_G511gat_6[2]),.dinb(w_G35gat_2[2]),.dout(n943),.clk(gclk));
	jand g0880(.dina(w_n927_0[1]),.dinb(w_n844_0[1]),.dout(n944),.clk(gclk));
	jnot g0881(.din(n944),.dout(n945),.clk(gclk));
	jnot g0882(.din(w_n927_0[0]),.dout(n946),.clk(gclk));
	jxor g0883(.dina(n946),.dinb(w_n844_0[0]),.dout(n947),.clk(gclk));
	jor g0884(.dina(n947),.dinb(w_n840_0[0]),.dout(n948),.clk(gclk));
	jand g0885(.dina(n948),.dinb(n945),.dout(n949),.clk(gclk));
	jand g0886(.dina(w_G494gat_6[1]),.dinb(w_G52gat_3[0]),.dout(n950),.clk(gclk));
	jnot g0887(.din(n950),.dout(n951),.clk(gclk));
	jand g0888(.dina(w_n925_0[0]),.dinb(w_n849_0[0]),.dout(n952),.clk(gclk));
	jand g0889(.dina(w_n926_0[0]),.dinb(w_n846_0[0]),.dout(n953),.clk(gclk));
	jor g0890(.dina(n953),.dinb(w_dff_B_vxmO1t5E1_1),.dout(n954),.clk(gclk));
	jand g0891(.dina(w_G477gat_6[0]),.dinb(w_G69gat_3[1]),.dout(n955),.clk(gclk));
	jnot g0892(.din(n955),.dout(n956),.clk(gclk));
	jand g0893(.dina(w_n923_0[0]),.dinb(w_n854_0[0]),.dout(n957),.clk(gclk));
	jand g0894(.dina(w_n924_0[0]),.dinb(w_n851_0[0]),.dout(n958),.clk(gclk));
	jor g0895(.dina(n958),.dinb(w_dff_B_Rb5srVo57_1),.dout(n959),.clk(gclk));
	jand g0896(.dina(w_G460gat_5[2]),.dinb(w_G86gat_3[2]),.dout(n960),.clk(gclk));
	jnot g0897(.din(n960),.dout(n961),.clk(gclk));
	jand g0898(.dina(w_n921_0[0]),.dinb(w_n859_0[0]),.dout(n962),.clk(gclk));
	jand g0899(.dina(w_n922_0[0]),.dinb(w_n856_0[0]),.dout(n963),.clk(gclk));
	jor g0900(.dina(n963),.dinb(w_dff_B_Ty6trjOr3_1),.dout(n964),.clk(gclk));
	jand g0901(.dina(w_G443gat_5[1]),.dinb(w_G103gat_4[0]),.dout(n965),.clk(gclk));
	jnot g0902(.din(n965),.dout(n966),.clk(gclk));
	jand g0903(.dina(w_n919_0[0]),.dinb(w_n864_0[0]),.dout(n967),.clk(gclk));
	jand g0904(.dina(w_n920_0[0]),.dinb(w_n861_0[0]),.dout(n968),.clk(gclk));
	jor g0905(.dina(n968),.dinb(w_dff_B_rM9QpD1R3_1),.dout(n969),.clk(gclk));
	jand g0906(.dina(w_G426gat_5[0]),.dinb(w_G120gat_4[1]),.dout(n970),.clk(gclk));
	jnot g0907(.din(n970),.dout(n971),.clk(gclk));
	jand g0908(.dina(w_n917_0[0]),.dinb(w_n869_0[0]),.dout(n972),.clk(gclk));
	jand g0909(.dina(w_n918_0[0]),.dinb(w_n866_0[0]),.dout(n973),.clk(gclk));
	jor g0910(.dina(n973),.dinb(w_dff_B_P00V99xF6_1),.dout(n974),.clk(gclk));
	jand g0911(.dina(w_G409gat_4[2]),.dinb(w_G137gat_4[2]),.dout(n975),.clk(gclk));
	jnot g0912(.din(n975),.dout(n976),.clk(gclk));
	jand g0913(.dina(w_n915_0[0]),.dinb(w_n874_0[0]),.dout(n977),.clk(gclk));
	jand g0914(.dina(w_n916_0[0]),.dinb(w_n871_0[0]),.dout(n978),.clk(gclk));
	jor g0915(.dina(n978),.dinb(w_dff_B_KizjIKLD4_1),.dout(n979),.clk(gclk));
	jand g0916(.dina(w_G392gat_4[1]),.dinb(w_G154gat_5[0]),.dout(n980),.clk(gclk));
	jnot g0917(.din(n980),.dout(n981),.clk(gclk));
	jand g0918(.dina(w_n913_0[0]),.dinb(w_n879_0[0]),.dout(n982),.clk(gclk));
	jand g0919(.dina(w_n914_0[0]),.dinb(w_n876_0[0]),.dout(n983),.clk(gclk));
	jor g0920(.dina(n983),.dinb(w_dff_B_xA5TsFm41_1),.dout(n984),.clk(gclk));
	jand g0921(.dina(w_G375gat_4[0]),.dinb(w_G171gat_5[1]),.dout(n985),.clk(gclk));
	jnot g0922(.din(n985),.dout(n986),.clk(gclk));
	jand g0923(.dina(w_n911_0[0]),.dinb(w_n884_0[0]),.dout(n987),.clk(gclk));
	jand g0924(.dina(w_n912_0[0]),.dinb(w_n881_0[0]),.dout(n988),.clk(gclk));
	jor g0925(.dina(n988),.dinb(w_dff_B_nYni0s4q4_1),.dout(n989),.clk(gclk));
	jand g0926(.dina(w_G358gat_3[2]),.dinb(w_G188gat_5[2]),.dout(n990),.clk(gclk));
	jnot g0927(.din(n990),.dout(n991),.clk(gclk));
	jand g0928(.dina(w_n909_0[0]),.dinb(w_n889_0[0]),.dout(n992),.clk(gclk));
	jand g0929(.dina(w_n910_0[0]),.dinb(w_n886_0[0]),.dout(n993),.clk(gclk));
	jor g0930(.dina(n993),.dinb(w_dff_B_SB7dlvBc6_1),.dout(n994),.clk(gclk));
	jand g0931(.dina(w_G341gat_3[1]),.dinb(w_G205gat_6[0]),.dout(n995),.clk(gclk));
	jnot g0932(.din(n995),.dout(n996),.clk(gclk));
	jand g0933(.dina(w_n907_0[0]),.dinb(w_n895_0[0]),.dout(n997),.clk(gclk));
	jand g0934(.dina(w_n908_0[0]),.dinb(w_n891_0[0]),.dout(n998),.clk(gclk));
	jor g0935(.dina(n998),.dinb(w_dff_B_PJf0cWwu9_1),.dout(n999),.clk(gclk));
	jand g0936(.dina(w_G324gat_3[0]),.dinb(w_G222gat_6[1]),.dout(n1000),.clk(gclk));
	jnot g0937(.din(n1000),.dout(n1001),.clk(gclk));
	jnot g0938(.din(w_n896_0[0]),.dout(n1002),.clk(gclk));
	jnot g0939(.din(w_n906_0[0]),.dout(n1003),.clk(gclk));
	jand g0940(.dina(n1003),.dinb(w_dff_B_7ocKJlph9_1),.dout(n1004),.clk(gclk));
	jor g0941(.dina(n1004),.dinb(w_n903_0[0]),.dout(n1005),.clk(gclk));
	jand g0942(.dina(w_G307gat_3[0]),.dinb(w_G239gat_6[2]),.dout(n1006),.clk(gclk));
	jand g0943(.dina(w_G290gat_2[1]),.dinb(w_G256gat_7[0]),.dout(n1007),.clk(gclk));
	jnot g0944(.din(n1007),.dout(n1008),.clk(gclk));
	jor g0945(.dina(w_n1008_0[1]),.dinb(w_n793_0[0]),.dout(n1009),.clk(gclk));
	jxor g0946(.dina(w_n1009_0[1]),.dinb(w_n1006_0[1]),.dout(n1010),.clk(gclk));
	jxor g0947(.dina(w_n1010_0[1]),.dinb(w_n1005_0[1]),.dout(n1011),.clk(gclk));
	jxor g0948(.dina(w_n1011_0[1]),.dinb(w_n1001_0[1]),.dout(n1012),.clk(gclk));
	jxor g0949(.dina(w_n1012_0[1]),.dinb(w_n999_0[1]),.dout(n1013),.clk(gclk));
	jxor g0950(.dina(w_n1013_0[1]),.dinb(w_n996_0[1]),.dout(n1014),.clk(gclk));
	jxor g0951(.dina(w_n1014_0[1]),.dinb(w_n994_0[1]),.dout(n1015),.clk(gclk));
	jxor g0952(.dina(w_n1015_0[1]),.dinb(w_n991_0[1]),.dout(n1016),.clk(gclk));
	jxor g0953(.dina(w_n1016_0[1]),.dinb(w_n989_0[1]),.dout(n1017),.clk(gclk));
	jxor g0954(.dina(w_n1017_0[1]),.dinb(w_n986_0[1]),.dout(n1018),.clk(gclk));
	jxor g0955(.dina(w_n1018_0[1]),.dinb(w_n984_0[1]),.dout(n1019),.clk(gclk));
	jxor g0956(.dina(w_n1019_0[1]),.dinb(w_n981_0[1]),.dout(n1020),.clk(gclk));
	jxor g0957(.dina(w_n1020_0[1]),.dinb(w_n979_0[1]),.dout(n1021),.clk(gclk));
	jxor g0958(.dina(w_n1021_0[1]),.dinb(w_n976_0[1]),.dout(n1022),.clk(gclk));
	jxor g0959(.dina(w_n1022_0[1]),.dinb(w_n974_0[1]),.dout(n1023),.clk(gclk));
	jxor g0960(.dina(w_n1023_0[1]),.dinb(w_n971_0[1]),.dout(n1024),.clk(gclk));
	jxor g0961(.dina(w_n1024_0[1]),.dinb(w_n969_0[1]),.dout(n1025),.clk(gclk));
	jxor g0962(.dina(w_n1025_0[1]),.dinb(w_n966_0[1]),.dout(n1026),.clk(gclk));
	jxor g0963(.dina(w_n1026_0[1]),.dinb(w_n964_0[1]),.dout(n1027),.clk(gclk));
	jxor g0964(.dina(w_n1027_0[1]),.dinb(w_n961_0[1]),.dout(n1028),.clk(gclk));
	jxor g0965(.dina(w_n1028_0[1]),.dinb(w_n959_0[1]),.dout(n1029),.clk(gclk));
	jxor g0966(.dina(w_n1029_0[1]),.dinb(w_n956_0[1]),.dout(n1030),.clk(gclk));
	jxor g0967(.dina(w_n1030_0[1]),.dinb(w_n954_0[1]),.dout(n1031),.clk(gclk));
	jxor g0968(.dina(w_n1031_0[1]),.dinb(w_n951_0[1]),.dout(n1032),.clk(gclk));
	jxor g0969(.dina(w_n1032_0[1]),.dinb(w_n949_0[1]),.dout(n1033),.clk(gclk));
	jxor g0970(.dina(w_n1033_0[1]),.dinb(w_n943_0[1]),.dout(n1034),.clk(gclk));
	jnot g0971(.din(w_n1034_0[1]),.dout(n1035),.clk(gclk));
	jxor g0972(.dina(w_n1035_0[1]),.dinb(w_n942_0[2]),.dout(n1036),.clk(gclk));
	jxor g0973(.dina(n1036),.dinb(w_n938_0[1]),.dout(n1037),.clk(gclk));
	jxor g0974(.dina(w_n1037_0[1]),.dinb(w_n937_0[1]),.dout(w_dff_A_GkoBMSiy7_2),.clk(gclk));
	jand g0975(.dina(w_n1037_0[0]),.dinb(w_n937_0[0]),.dout(n1039),.clk(gclk));
	jor g0976(.dina(w_n1035_0[0]),.dinb(w_n942_0[1]),.dout(n1040),.clk(gclk));
	jxor g0977(.dina(w_n1034_0[0]),.dinb(w_n942_0[0]),.dout(n1041),.clk(gclk));
	jor g0978(.dina(n1041),.dinb(w_n938_0[0]),.dout(n1042),.clk(gclk));
	jand g0979(.dina(n1042),.dinb(w_dff_B_oFoXuBJi1_1),.dout(n1043),.clk(gclk));
	jand g0980(.dina(w_G528gat_6[2]),.dinb(w_G35gat_2[1]),.dout(n1044),.clk(gclk));
	jnot g0981(.din(w_n1032_0[0]),.dout(n1045),.clk(gclk));
	jor g0982(.dina(n1045),.dinb(w_n949_0[0]),.dout(n1046),.clk(gclk));
	jor g0983(.dina(w_n1033_0[0]),.dinb(w_n943_0[0]),.dout(n1047),.clk(gclk));
	jand g0984(.dina(n1047),.dinb(w_dff_B_ixj7yUiC0_1),.dout(n1048),.clk(gclk));
	jand g0985(.dina(w_G511gat_6[1]),.dinb(w_G52gat_2[2]),.dout(n1049),.clk(gclk));
	jand g0986(.dina(w_n1030_0[0]),.dinb(w_n954_0[0]),.dout(n1050),.clk(gclk));
	jand g0987(.dina(w_n1031_0[0]),.dinb(w_n951_0[0]),.dout(n1051),.clk(gclk));
	jor g0988(.dina(n1051),.dinb(w_dff_B_877gKBVH1_1),.dout(n1052),.clk(gclk));
	jand g0989(.dina(w_G494gat_6[0]),.dinb(w_G69gat_3[0]),.dout(n1053),.clk(gclk));
	jnot g0990(.din(n1053),.dout(n1054),.clk(gclk));
	jand g0991(.dina(w_n1028_0[0]),.dinb(w_n959_0[0]),.dout(n1055),.clk(gclk));
	jand g0992(.dina(w_n1029_0[0]),.dinb(w_n956_0[0]),.dout(n1056),.clk(gclk));
	jor g0993(.dina(n1056),.dinb(w_dff_B_eCtGb53e0_1),.dout(n1057),.clk(gclk));
	jand g0994(.dina(w_G477gat_5[2]),.dinb(w_G86gat_3[1]),.dout(n1058),.clk(gclk));
	jnot g0995(.din(n1058),.dout(n1059),.clk(gclk));
	jand g0996(.dina(w_n1026_0[0]),.dinb(w_n964_0[0]),.dout(n1060),.clk(gclk));
	jand g0997(.dina(w_n1027_0[0]),.dinb(w_n961_0[0]),.dout(n1061),.clk(gclk));
	jor g0998(.dina(n1061),.dinb(w_dff_B_UhIogdie1_1),.dout(n1062),.clk(gclk));
	jand g0999(.dina(w_G460gat_5[1]),.dinb(w_G103gat_3[2]),.dout(n1063),.clk(gclk));
	jnot g1000(.din(n1063),.dout(n1064),.clk(gclk));
	jand g1001(.dina(w_n1024_0[0]),.dinb(w_n969_0[0]),.dout(n1065),.clk(gclk));
	jand g1002(.dina(w_n1025_0[0]),.dinb(w_n966_0[0]),.dout(n1066),.clk(gclk));
	jor g1003(.dina(n1066),.dinb(w_dff_B_Z0oss8sb3_1),.dout(n1067),.clk(gclk));
	jand g1004(.dina(w_G443gat_5[0]),.dinb(w_G120gat_4[0]),.dout(n1068),.clk(gclk));
	jnot g1005(.din(n1068),.dout(n1069),.clk(gclk));
	jand g1006(.dina(w_n1022_0[0]),.dinb(w_n974_0[0]),.dout(n1070),.clk(gclk));
	jand g1007(.dina(w_n1023_0[0]),.dinb(w_n971_0[0]),.dout(n1071),.clk(gclk));
	jor g1008(.dina(n1071),.dinb(w_dff_B_EU9fSBA64_1),.dout(n1072),.clk(gclk));
	jand g1009(.dina(w_G426gat_4[2]),.dinb(w_G137gat_4[1]),.dout(n1073),.clk(gclk));
	jnot g1010(.din(n1073),.dout(n1074),.clk(gclk));
	jand g1011(.dina(w_n1020_0[0]),.dinb(w_n979_0[0]),.dout(n1075),.clk(gclk));
	jand g1012(.dina(w_n1021_0[0]),.dinb(w_n976_0[0]),.dout(n1076),.clk(gclk));
	jor g1013(.dina(n1076),.dinb(w_dff_B_Xewy7ynQ2_1),.dout(n1077),.clk(gclk));
	jand g1014(.dina(w_G409gat_4[1]),.dinb(w_G154gat_4[2]),.dout(n1078),.clk(gclk));
	jnot g1015(.din(n1078),.dout(n1079),.clk(gclk));
	jand g1016(.dina(w_n1018_0[0]),.dinb(w_n984_0[0]),.dout(n1080),.clk(gclk));
	jand g1017(.dina(w_n1019_0[0]),.dinb(w_n981_0[0]),.dout(n1081),.clk(gclk));
	jor g1018(.dina(n1081),.dinb(w_dff_B_IHPr1Lw29_1),.dout(n1082),.clk(gclk));
	jand g1019(.dina(w_G392gat_4[0]),.dinb(w_G171gat_5[0]),.dout(n1083),.clk(gclk));
	jnot g1020(.din(n1083),.dout(n1084),.clk(gclk));
	jand g1021(.dina(w_n1016_0[0]),.dinb(w_n989_0[0]),.dout(n1085),.clk(gclk));
	jand g1022(.dina(w_n1017_0[0]),.dinb(w_n986_0[0]),.dout(n1086),.clk(gclk));
	jor g1023(.dina(n1086),.dinb(w_dff_B_g9P1r5ym0_1),.dout(n1087),.clk(gclk));
	jand g1024(.dina(w_G375gat_3[2]),.dinb(w_G188gat_5[1]),.dout(n1088),.clk(gclk));
	jnot g1025(.din(n1088),.dout(n1089),.clk(gclk));
	jand g1026(.dina(w_n1014_0[0]),.dinb(w_n994_0[0]),.dout(n1090),.clk(gclk));
	jand g1027(.dina(w_n1015_0[0]),.dinb(w_n991_0[0]),.dout(n1091),.clk(gclk));
	jor g1028(.dina(n1091),.dinb(w_dff_B_yk5YtVJ65_1),.dout(n1092),.clk(gclk));
	jand g1029(.dina(w_G358gat_3[1]),.dinb(w_G205gat_5[2]),.dout(n1093),.clk(gclk));
	jnot g1030(.din(n1093),.dout(n1094),.clk(gclk));
	jand g1031(.dina(w_n1012_0[0]),.dinb(w_n999_0[0]),.dout(n1095),.clk(gclk));
	jand g1032(.dina(w_n1013_0[0]),.dinb(w_n996_0[0]),.dout(n1096),.clk(gclk));
	jor g1033(.dina(n1096),.dinb(w_dff_B_JdMX0b1g2_1),.dout(n1097),.clk(gclk));
	jand g1034(.dina(w_G341gat_3[0]),.dinb(w_G222gat_6[0]),.dout(n1098),.clk(gclk));
	jnot g1035(.din(n1098),.dout(n1099),.clk(gclk));
	jand g1036(.dina(w_n1010_0[0]),.dinb(w_n1005_0[0]),.dout(n1100),.clk(gclk));
	jand g1037(.dina(w_n1011_0[0]),.dinb(w_n1001_0[0]),.dout(n1101),.clk(gclk));
	jor g1038(.dina(n1101),.dinb(w_dff_B_cmfpmCl56_1),.dout(n1102),.clk(gclk));
	jand g1039(.dina(w_G324gat_2[2]),.dinb(w_G239gat_6[1]),.dout(n1103),.clk(gclk));
	jand g1040(.dina(w_G307gat_2[2]),.dinb(w_G256gat_6[2]),.dout(n1104),.clk(gclk));
	jnot g1041(.din(w_n1006_0[0]),.dout(n1105),.clk(gclk));
	jnot g1042(.din(w_n1009_0[0]),.dout(n1106),.clk(gclk));
	jand g1043(.dina(n1106),.dinb(w_dff_B_IWVdypPc3_1),.dout(n1107),.clk(gclk));
	jor g1044(.dina(n1107),.dinb(w_n1008_0[0]),.dout(n1108),.clk(gclk));
	jnot g1045(.din(n1108),.dout(n1109),.clk(gclk));
	jor g1046(.dina(w_n1109_0[1]),.dinb(w_dff_B_B5JNyJST3_1),.dout(n1110),.clk(gclk));
	jand g1047(.dina(w_n1109_0[0]),.dinb(w_G307gat_2[1]),.dout(n1111),.clk(gclk));
	jnot g1048(.din(n1111),.dout(n1112),.clk(gclk));
	jand g1049(.dina(n1112),.dinb(w_n1110_0[1]),.dout(n1113),.clk(gclk));
	jnot g1050(.din(n1113),.dout(n1114),.clk(gclk));
	jxor g1051(.dina(w_n1114_0[1]),.dinb(w_n1103_0[1]),.dout(n1115),.clk(gclk));
	jxor g1052(.dina(w_n1115_0[1]),.dinb(w_n1102_0[1]),.dout(n1116),.clk(gclk));
	jxor g1053(.dina(w_n1116_0[1]),.dinb(w_n1099_0[1]),.dout(n1117),.clk(gclk));
	jxor g1054(.dina(w_n1117_0[1]),.dinb(w_n1097_0[1]),.dout(n1118),.clk(gclk));
	jxor g1055(.dina(w_n1118_0[1]),.dinb(w_n1094_0[1]),.dout(n1119),.clk(gclk));
	jxor g1056(.dina(w_n1119_0[1]),.dinb(w_n1092_0[1]),.dout(n1120),.clk(gclk));
	jxor g1057(.dina(w_n1120_0[1]),.dinb(w_n1089_0[1]),.dout(n1121),.clk(gclk));
	jxor g1058(.dina(w_n1121_0[1]),.dinb(w_n1087_0[1]),.dout(n1122),.clk(gclk));
	jxor g1059(.dina(w_n1122_0[1]),.dinb(w_n1084_0[1]),.dout(n1123),.clk(gclk));
	jxor g1060(.dina(w_n1123_0[1]),.dinb(w_n1082_0[1]),.dout(n1124),.clk(gclk));
	jxor g1061(.dina(w_n1124_0[1]),.dinb(w_n1079_0[1]),.dout(n1125),.clk(gclk));
	jxor g1062(.dina(w_n1125_0[1]),.dinb(w_n1077_0[1]),.dout(n1126),.clk(gclk));
	jxor g1063(.dina(w_n1126_0[1]),.dinb(w_n1074_0[1]),.dout(n1127),.clk(gclk));
	jxor g1064(.dina(w_n1127_0[1]),.dinb(w_n1072_0[1]),.dout(n1128),.clk(gclk));
	jxor g1065(.dina(w_n1128_0[1]),.dinb(w_n1069_0[1]),.dout(n1129),.clk(gclk));
	jxor g1066(.dina(w_n1129_0[1]),.dinb(w_n1067_0[1]),.dout(n1130),.clk(gclk));
	jxor g1067(.dina(w_n1130_0[1]),.dinb(w_n1064_0[1]),.dout(n1131),.clk(gclk));
	jxor g1068(.dina(w_n1131_0[1]),.dinb(w_n1062_0[1]),.dout(n1132),.clk(gclk));
	jxor g1069(.dina(w_n1132_0[1]),.dinb(w_n1059_0[1]),.dout(n1133),.clk(gclk));
	jxor g1070(.dina(w_n1133_0[1]),.dinb(w_n1057_0[1]),.dout(n1134),.clk(gclk));
	jxor g1071(.dina(w_n1134_0[1]),.dinb(w_n1054_0[1]),.dout(n1135),.clk(gclk));
	jxor g1072(.dina(w_n1135_0[1]),.dinb(w_n1052_0[1]),.dout(n1136),.clk(gclk));
	jnot g1073(.din(n1136),.dout(n1137),.clk(gclk));
	jxor g1074(.dina(w_n1137_0[1]),.dinb(w_n1049_0[1]),.dout(n1138),.clk(gclk));
	jxor g1075(.dina(w_n1138_0[1]),.dinb(w_n1048_0[1]),.dout(n1139),.clk(gclk));
	jxor g1076(.dina(w_n1139_0[1]),.dinb(w_n1044_0[1]),.dout(n1140),.clk(gclk));
	jxor g1077(.dina(w_n1140_0[1]),.dinb(w_n1043_0[1]),.dout(n1141),.clk(gclk));
	jnot g1078(.din(w_n1141_0[1]),.dout(n1142),.clk(gclk));
	jxor g1079(.dina(n1142),.dinb(w_n1039_0[1]),.dout(w_dff_A_fgq1tWlH0_2),.clk(gclk));
	jnot g1080(.din(w_n1140_0[0]),.dout(n1144),.clk(gclk));
	jor g1081(.dina(n1144),.dinb(w_n1043_0[0]),.dout(n1145),.clk(gclk));
	jor g1082(.dina(w_n1141_0[0]),.dinb(w_n1039_0[0]),.dout(n1146),.clk(gclk));
	jand g1083(.dina(n1146),.dinb(w_dff_B_YxY9L11J6_1),.dout(n1147),.clk(gclk));
	jnot g1084(.din(w_n1138_0[0]),.dout(n1148),.clk(gclk));
	jor g1085(.dina(n1148),.dinb(w_n1048_0[0]),.dout(n1149),.clk(gclk));
	jor g1086(.dina(w_n1139_0[0]),.dinb(w_n1044_0[0]),.dout(n1150),.clk(gclk));
	jand g1087(.dina(n1150),.dinb(n1149),.dout(n1151),.clk(gclk));
	jand g1088(.dina(w_G528gat_6[1]),.dinb(w_G52gat_2[1]),.dout(n1152),.clk(gclk));
	jand g1089(.dina(w_n1135_0[0]),.dinb(w_n1052_0[0]),.dout(n1153),.clk(gclk));
	jnot g1090(.din(n1153),.dout(n1154),.clk(gclk));
	jor g1091(.dina(w_n1137_0[0]),.dinb(w_n1049_0[0]),.dout(n1155),.clk(gclk));
	jand g1092(.dina(n1155),.dinb(w_dff_B_KiUGehzL6_1),.dout(n1156),.clk(gclk));
	jand g1093(.dina(w_G511gat_6[0]),.dinb(w_G69gat_2[2]),.dout(n1157),.clk(gclk));
	jnot g1094(.din(n1157),.dout(n1158),.clk(gclk));
	jand g1095(.dina(w_n1133_0[0]),.dinb(w_n1057_0[0]),.dout(n1159),.clk(gclk));
	jand g1096(.dina(w_n1134_0[0]),.dinb(w_n1054_0[0]),.dout(n1160),.clk(gclk));
	jor g1097(.dina(n1160),.dinb(w_dff_B_lOSBJ7tE3_1),.dout(n1161),.clk(gclk));
	jand g1098(.dina(w_G494gat_5[2]),.dinb(w_G86gat_3[0]),.dout(n1162),.clk(gclk));
	jnot g1099(.din(n1162),.dout(n1163),.clk(gclk));
	jand g1100(.dina(w_n1131_0[0]),.dinb(w_n1062_0[0]),.dout(n1164),.clk(gclk));
	jand g1101(.dina(w_n1132_0[0]),.dinb(w_n1059_0[0]),.dout(n1165),.clk(gclk));
	jor g1102(.dina(n1165),.dinb(w_dff_B_uOEOZObL3_1),.dout(n1166),.clk(gclk));
	jand g1103(.dina(w_G477gat_5[1]),.dinb(w_G103gat_3[1]),.dout(n1167),.clk(gclk));
	jnot g1104(.din(n1167),.dout(n1168),.clk(gclk));
	jand g1105(.dina(w_n1129_0[0]),.dinb(w_n1067_0[0]),.dout(n1169),.clk(gclk));
	jand g1106(.dina(w_n1130_0[0]),.dinb(w_n1064_0[0]),.dout(n1170),.clk(gclk));
	jor g1107(.dina(n1170),.dinb(w_dff_B_Ow6XnM5z2_1),.dout(n1171),.clk(gclk));
	jand g1108(.dina(w_G460gat_5[0]),.dinb(w_G120gat_3[2]),.dout(n1172),.clk(gclk));
	jnot g1109(.din(n1172),.dout(n1173),.clk(gclk));
	jand g1110(.dina(w_n1127_0[0]),.dinb(w_n1072_0[0]),.dout(n1174),.clk(gclk));
	jand g1111(.dina(w_n1128_0[0]),.dinb(w_n1069_0[0]),.dout(n1175),.clk(gclk));
	jor g1112(.dina(n1175),.dinb(w_dff_B_0sSPHn4O8_1),.dout(n1176),.clk(gclk));
	jand g1113(.dina(w_G443gat_4[2]),.dinb(w_G137gat_4[0]),.dout(n1177),.clk(gclk));
	jnot g1114(.din(n1177),.dout(n1178),.clk(gclk));
	jand g1115(.dina(w_n1125_0[0]),.dinb(w_n1077_0[0]),.dout(n1179),.clk(gclk));
	jand g1116(.dina(w_n1126_0[0]),.dinb(w_n1074_0[0]),.dout(n1180),.clk(gclk));
	jor g1117(.dina(n1180),.dinb(w_dff_B_uzd3W8qA3_1),.dout(n1181),.clk(gclk));
	jand g1118(.dina(w_G426gat_4[1]),.dinb(w_G154gat_4[1]),.dout(n1182),.clk(gclk));
	jnot g1119(.din(n1182),.dout(n1183),.clk(gclk));
	jand g1120(.dina(w_n1123_0[0]),.dinb(w_n1082_0[0]),.dout(n1184),.clk(gclk));
	jand g1121(.dina(w_n1124_0[0]),.dinb(w_n1079_0[0]),.dout(n1185),.clk(gclk));
	jor g1122(.dina(n1185),.dinb(w_dff_B_k0AmojMX2_1),.dout(n1186),.clk(gclk));
	jand g1123(.dina(w_G409gat_4[0]),.dinb(w_G171gat_4[2]),.dout(n1187),.clk(gclk));
	jnot g1124(.din(n1187),.dout(n1188),.clk(gclk));
	jand g1125(.dina(w_n1121_0[0]),.dinb(w_n1087_0[0]),.dout(n1189),.clk(gclk));
	jand g1126(.dina(w_n1122_0[0]),.dinb(w_n1084_0[0]),.dout(n1190),.clk(gclk));
	jor g1127(.dina(n1190),.dinb(w_dff_B_teh9vl1E7_1),.dout(n1191),.clk(gclk));
	jand g1128(.dina(w_G392gat_3[2]),.dinb(w_G188gat_5[0]),.dout(n1192),.clk(gclk));
	jnot g1129(.din(n1192),.dout(n1193),.clk(gclk));
	jand g1130(.dina(w_n1119_0[0]),.dinb(w_n1092_0[0]),.dout(n1194),.clk(gclk));
	jand g1131(.dina(w_n1120_0[0]),.dinb(w_n1089_0[0]),.dout(n1195),.clk(gclk));
	jor g1132(.dina(n1195),.dinb(w_dff_B_kK2ESgpI4_1),.dout(n1196),.clk(gclk));
	jand g1133(.dina(w_G375gat_3[1]),.dinb(w_G205gat_5[1]),.dout(n1197),.clk(gclk));
	jnot g1134(.din(n1197),.dout(n1198),.clk(gclk));
	jand g1135(.dina(w_n1117_0[0]),.dinb(w_n1097_0[0]),.dout(n1199),.clk(gclk));
	jand g1136(.dina(w_n1118_0[0]),.dinb(w_n1094_0[0]),.dout(n1200),.clk(gclk));
	jor g1137(.dina(n1200),.dinb(w_dff_B_af6URBAC0_1),.dout(n1201),.clk(gclk));
	jand g1138(.dina(w_G358gat_3[0]),.dinb(w_G222gat_5[2]),.dout(n1202),.clk(gclk));
	jnot g1139(.din(n1202),.dout(n1203),.clk(gclk));
	jand g1140(.dina(w_n1115_0[0]),.dinb(w_n1102_0[0]),.dout(n1204),.clk(gclk));
	jand g1141(.dina(w_n1116_0[0]),.dinb(w_n1099_0[0]),.dout(n1205),.clk(gclk));
	jor g1142(.dina(n1205),.dinb(w_dff_B_ekLgpStc5_1),.dout(n1206),.clk(gclk));
	jand g1143(.dina(w_G341gat_2[2]),.dinb(w_G239gat_6[0]),.dout(n1207),.clk(gclk));
	jand g1144(.dina(w_G324gat_2[1]),.dinb(w_G256gat_6[1]),.dout(n1208),.clk(gclk));
	jor g1145(.dina(w_n1114_0[0]),.dinb(w_n1103_0[0]),.dout(n1209),.clk(gclk));
	jand g1146(.dina(n1209),.dinb(w_n1110_0[0]),.dout(n1210),.clk(gclk));
	jxor g1147(.dina(w_n1210_0[1]),.dinb(w_n1208_0[1]),.dout(n1211),.clk(gclk));
	jnot g1148(.din(n1211),.dout(n1212),.clk(gclk));
	jxor g1149(.dina(w_n1212_0[1]),.dinb(w_n1207_0[1]),.dout(n1213),.clk(gclk));
	jxor g1150(.dina(w_n1213_0[1]),.dinb(w_n1206_0[1]),.dout(n1214),.clk(gclk));
	jxor g1151(.dina(w_n1214_0[1]),.dinb(w_n1203_0[1]),.dout(n1215),.clk(gclk));
	jxor g1152(.dina(w_n1215_0[1]),.dinb(w_n1201_0[1]),.dout(n1216),.clk(gclk));
	jxor g1153(.dina(w_n1216_0[1]),.dinb(w_n1198_0[1]),.dout(n1217),.clk(gclk));
	jxor g1154(.dina(w_n1217_0[1]),.dinb(w_n1196_0[1]),.dout(n1218),.clk(gclk));
	jxor g1155(.dina(w_n1218_0[1]),.dinb(w_n1193_0[1]),.dout(n1219),.clk(gclk));
	jxor g1156(.dina(w_n1219_0[1]),.dinb(w_n1191_0[1]),.dout(n1220),.clk(gclk));
	jxor g1157(.dina(w_n1220_0[1]),.dinb(w_n1188_0[1]),.dout(n1221),.clk(gclk));
	jxor g1158(.dina(w_n1221_0[1]),.dinb(w_n1186_0[1]),.dout(n1222),.clk(gclk));
	jxor g1159(.dina(w_n1222_0[1]),.dinb(w_n1183_0[1]),.dout(n1223),.clk(gclk));
	jxor g1160(.dina(w_n1223_0[1]),.dinb(w_n1181_0[1]),.dout(n1224),.clk(gclk));
	jxor g1161(.dina(w_n1224_0[1]),.dinb(w_n1178_0[1]),.dout(n1225),.clk(gclk));
	jxor g1162(.dina(w_n1225_0[1]),.dinb(w_n1176_0[1]),.dout(n1226),.clk(gclk));
	jxor g1163(.dina(w_n1226_0[1]),.dinb(w_n1173_0[1]),.dout(n1227),.clk(gclk));
	jxor g1164(.dina(w_n1227_0[1]),.dinb(w_n1171_0[1]),.dout(n1228),.clk(gclk));
	jxor g1165(.dina(w_n1228_0[1]),.dinb(w_n1168_0[1]),.dout(n1229),.clk(gclk));
	jxor g1166(.dina(w_n1229_0[1]),.dinb(w_n1166_0[1]),.dout(n1230),.clk(gclk));
	jxor g1167(.dina(w_n1230_0[1]),.dinb(w_n1163_0[1]),.dout(n1231),.clk(gclk));
	jxor g1168(.dina(w_n1231_0[1]),.dinb(w_n1161_0[1]),.dout(n1232),.clk(gclk));
	jxor g1169(.dina(w_n1232_0[1]),.dinb(w_n1158_0[1]),.dout(n1233),.clk(gclk));
	jnot g1170(.din(n1233),.dout(n1234),.clk(gclk));
	jxor g1171(.dina(w_n1234_0[1]),.dinb(w_n1156_0[1]),.dout(n1235),.clk(gclk));
	jnot g1172(.din(n1235),.dout(n1236),.clk(gclk));
	jxor g1173(.dina(w_n1236_0[1]),.dinb(w_n1152_0[1]),.dout(n1237),.clk(gclk));
	jxor g1174(.dina(w_n1237_0[1]),.dinb(w_n1151_0[1]),.dout(n1238),.clk(gclk));
	jnot g1175(.din(w_n1238_0[1]),.dout(n1239),.clk(gclk));
	jxor g1176(.dina(n1239),.dinb(w_n1147_0[1]),.dout(w_dff_A_obuUdNIl2_2),.clk(gclk));
	jnot g1177(.din(w_n1237_0[0]),.dout(n1241),.clk(gclk));
	jor g1178(.dina(n1241),.dinb(w_n1151_0[0]),.dout(n1242),.clk(gclk));
	jor g1179(.dina(w_n1238_0[0]),.dinb(w_n1147_0[0]),.dout(n1243),.clk(gclk));
	jand g1180(.dina(n1243),.dinb(w_dff_B_BFNl21zT8_1),.dout(n1244),.clk(gclk));
	jor g1181(.dina(w_n1234_0[0]),.dinb(w_n1156_0[0]),.dout(n1245),.clk(gclk));
	jor g1182(.dina(w_n1236_0[0]),.dinb(w_n1152_0[0]),.dout(n1246),.clk(gclk));
	jand g1183(.dina(n1246),.dinb(w_dff_B_Xe2jUCZn7_1),.dout(n1247),.clk(gclk));
	jand g1184(.dina(w_G528gat_6[0]),.dinb(w_G69gat_2[1]),.dout(n1248),.clk(gclk));
	jand g1185(.dina(w_n1231_0[0]),.dinb(w_n1161_0[0]),.dout(n1249),.clk(gclk));
	jand g1186(.dina(w_n1232_0[0]),.dinb(w_n1158_0[0]),.dout(n1250),.clk(gclk));
	jor g1187(.dina(n1250),.dinb(w_dff_B_JQvbpp403_1),.dout(n1251),.clk(gclk));
	jand g1188(.dina(w_G511gat_5[2]),.dinb(w_G86gat_2[2]),.dout(n1252),.clk(gclk));
	jnot g1189(.din(n1252),.dout(n1253),.clk(gclk));
	jand g1190(.dina(w_n1229_0[0]),.dinb(w_n1166_0[0]),.dout(n1254),.clk(gclk));
	jand g1191(.dina(w_n1230_0[0]),.dinb(w_n1163_0[0]),.dout(n1255),.clk(gclk));
	jor g1192(.dina(n1255),.dinb(w_dff_B_veZHBUJv1_1),.dout(n1256),.clk(gclk));
	jand g1193(.dina(w_G494gat_5[1]),.dinb(w_G103gat_3[0]),.dout(n1257),.clk(gclk));
	jnot g1194(.din(n1257),.dout(n1258),.clk(gclk));
	jand g1195(.dina(w_n1227_0[0]),.dinb(w_n1171_0[0]),.dout(n1259),.clk(gclk));
	jand g1196(.dina(w_n1228_0[0]),.dinb(w_n1168_0[0]),.dout(n1260),.clk(gclk));
	jor g1197(.dina(n1260),.dinb(w_dff_B_9SfuAkYY9_1),.dout(n1261),.clk(gclk));
	jand g1198(.dina(w_G477gat_5[0]),.dinb(w_G120gat_3[1]),.dout(n1262),.clk(gclk));
	jnot g1199(.din(n1262),.dout(n1263),.clk(gclk));
	jand g1200(.dina(w_n1225_0[0]),.dinb(w_n1176_0[0]),.dout(n1264),.clk(gclk));
	jand g1201(.dina(w_n1226_0[0]),.dinb(w_n1173_0[0]),.dout(n1265),.clk(gclk));
	jor g1202(.dina(n1265),.dinb(w_dff_B_ImpNrGtm4_1),.dout(n1266),.clk(gclk));
	jand g1203(.dina(w_G460gat_4[2]),.dinb(w_G137gat_3[2]),.dout(n1267),.clk(gclk));
	jnot g1204(.din(n1267),.dout(n1268),.clk(gclk));
	jand g1205(.dina(w_n1223_0[0]),.dinb(w_n1181_0[0]),.dout(n1269),.clk(gclk));
	jand g1206(.dina(w_n1224_0[0]),.dinb(w_n1178_0[0]),.dout(n1270),.clk(gclk));
	jor g1207(.dina(n1270),.dinb(w_dff_B_OV7ggkl04_1),.dout(n1271),.clk(gclk));
	jand g1208(.dina(w_G443gat_4[1]),.dinb(w_G154gat_4[0]),.dout(n1272),.clk(gclk));
	jnot g1209(.din(n1272),.dout(n1273),.clk(gclk));
	jand g1210(.dina(w_n1221_0[0]),.dinb(w_n1186_0[0]),.dout(n1274),.clk(gclk));
	jand g1211(.dina(w_n1222_0[0]),.dinb(w_n1183_0[0]),.dout(n1275),.clk(gclk));
	jor g1212(.dina(n1275),.dinb(w_dff_B_nwJXkFV64_1),.dout(n1276),.clk(gclk));
	jand g1213(.dina(w_G426gat_4[0]),.dinb(w_G171gat_4[1]),.dout(n1277),.clk(gclk));
	jnot g1214(.din(n1277),.dout(n1278),.clk(gclk));
	jand g1215(.dina(w_n1219_0[0]),.dinb(w_n1191_0[0]),.dout(n1279),.clk(gclk));
	jand g1216(.dina(w_n1220_0[0]),.dinb(w_n1188_0[0]),.dout(n1280),.clk(gclk));
	jor g1217(.dina(n1280),.dinb(w_dff_B_IZsyeWf28_1),.dout(n1281),.clk(gclk));
	jand g1218(.dina(w_G409gat_3[2]),.dinb(w_G188gat_4[2]),.dout(n1282),.clk(gclk));
	jnot g1219(.din(n1282),.dout(n1283),.clk(gclk));
	jand g1220(.dina(w_n1217_0[0]),.dinb(w_n1196_0[0]),.dout(n1284),.clk(gclk));
	jand g1221(.dina(w_n1218_0[0]),.dinb(w_n1193_0[0]),.dout(n1285),.clk(gclk));
	jor g1222(.dina(n1285),.dinb(w_dff_B_uZ7dF0Vi0_1),.dout(n1286),.clk(gclk));
	jand g1223(.dina(w_G392gat_3[1]),.dinb(w_G205gat_5[0]),.dout(n1287),.clk(gclk));
	jnot g1224(.din(n1287),.dout(n1288),.clk(gclk));
	jand g1225(.dina(w_n1215_0[0]),.dinb(w_n1201_0[0]),.dout(n1289),.clk(gclk));
	jand g1226(.dina(w_n1216_0[0]),.dinb(w_n1198_0[0]),.dout(n1290),.clk(gclk));
	jor g1227(.dina(n1290),.dinb(w_dff_B_Za8DoiXy7_1),.dout(n1291),.clk(gclk));
	jand g1228(.dina(w_G375gat_3[0]),.dinb(w_G222gat_5[1]),.dout(n1292),.clk(gclk));
	jnot g1229(.din(n1292),.dout(n1293),.clk(gclk));
	jand g1230(.dina(w_n1213_0[0]),.dinb(w_n1206_0[0]),.dout(n1294),.clk(gclk));
	jand g1231(.dina(w_n1214_0[0]),.dinb(w_n1203_0[0]),.dout(n1295),.clk(gclk));
	jor g1232(.dina(n1295),.dinb(w_dff_B_DZrKGAMs6_1),.dout(n1296),.clk(gclk));
	jand g1233(.dina(w_G358gat_2[2]),.dinb(w_G239gat_5[2]),.dout(n1297),.clk(gclk));
	jand g1234(.dina(w_G341gat_2[1]),.dinb(w_G256gat_6[0]),.dout(n1298),.clk(gclk));
	jor g1235(.dina(w_n1210_0[0]),.dinb(w_n1208_0[0]),.dout(n1299),.clk(gclk));
	jor g1236(.dina(w_n1212_0[0]),.dinb(w_n1207_0[0]),.dout(n1300),.clk(gclk));
	jand g1237(.dina(n1300),.dinb(w_dff_B_e2ET3Y1E7_1),.dout(n1301),.clk(gclk));
	jxor g1238(.dina(w_n1301_0[1]),.dinb(w_n1298_0[1]),.dout(n1302),.clk(gclk));
	jnot g1239(.din(n1302),.dout(n1303),.clk(gclk));
	jxor g1240(.dina(w_n1303_0[1]),.dinb(w_n1297_0[1]),.dout(n1304),.clk(gclk));
	jxor g1241(.dina(w_n1304_0[1]),.dinb(w_n1296_0[1]),.dout(n1305),.clk(gclk));
	jxor g1242(.dina(w_n1305_0[1]),.dinb(w_n1293_0[1]),.dout(n1306),.clk(gclk));
	jxor g1243(.dina(w_n1306_0[1]),.dinb(w_n1291_0[1]),.dout(n1307),.clk(gclk));
	jxor g1244(.dina(w_n1307_0[1]),.dinb(w_n1288_0[1]),.dout(n1308),.clk(gclk));
	jxor g1245(.dina(w_n1308_0[1]),.dinb(w_n1286_0[1]),.dout(n1309),.clk(gclk));
	jxor g1246(.dina(w_n1309_0[1]),.dinb(w_n1283_0[1]),.dout(n1310),.clk(gclk));
	jxor g1247(.dina(w_n1310_0[1]),.dinb(w_n1281_0[1]),.dout(n1311),.clk(gclk));
	jxor g1248(.dina(w_n1311_0[1]),.dinb(w_n1278_0[1]),.dout(n1312),.clk(gclk));
	jxor g1249(.dina(w_n1312_0[1]),.dinb(w_n1276_0[1]),.dout(n1313),.clk(gclk));
	jxor g1250(.dina(w_n1313_0[1]),.dinb(w_n1273_0[1]),.dout(n1314),.clk(gclk));
	jxor g1251(.dina(w_n1314_0[1]),.dinb(w_n1271_0[1]),.dout(n1315),.clk(gclk));
	jxor g1252(.dina(w_n1315_0[1]),.dinb(w_n1268_0[1]),.dout(n1316),.clk(gclk));
	jxor g1253(.dina(w_n1316_0[1]),.dinb(w_n1266_0[1]),.dout(n1317),.clk(gclk));
	jxor g1254(.dina(w_n1317_0[1]),.dinb(w_n1263_0[1]),.dout(n1318),.clk(gclk));
	jxor g1255(.dina(w_n1318_0[1]),.dinb(w_n1261_0[1]),.dout(n1319),.clk(gclk));
	jxor g1256(.dina(w_n1319_0[1]),.dinb(w_n1258_0[1]),.dout(n1320),.clk(gclk));
	jxor g1257(.dina(w_n1320_0[1]),.dinb(w_n1256_0[1]),.dout(n1321),.clk(gclk));
	jxor g1258(.dina(w_n1321_0[1]),.dinb(w_n1253_0[1]),.dout(n1322),.clk(gclk));
	jxor g1259(.dina(w_n1322_0[1]),.dinb(w_n1251_0[1]),.dout(n1323),.clk(gclk));
	jnot g1260(.din(n1323),.dout(n1324),.clk(gclk));
	jxor g1261(.dina(w_n1324_0[1]),.dinb(w_n1248_0[1]),.dout(n1325),.clk(gclk));
	jxor g1262(.dina(w_n1325_0[1]),.dinb(w_n1247_0[1]),.dout(n1326),.clk(gclk));
	jnot g1263(.din(w_n1326_0[1]),.dout(n1327),.clk(gclk));
	jxor g1264(.dina(w_dff_B_fMoeLlFX7_0),.dinb(w_n1244_0[1]),.dout(w_dff_A_XYc3sDAs5_2),.clk(gclk));
	jnot g1265(.din(w_n1325_0[0]),.dout(n1329),.clk(gclk));
	jor g1266(.dina(w_dff_B_iWR1jGX20_0),.dinb(w_n1247_0[0]),.dout(n1330),.clk(gclk));
	jor g1267(.dina(w_n1326_0[0]),.dinb(w_n1244_0[0]),.dout(n1331),.clk(gclk));
	jand g1268(.dina(n1331),.dinb(w_dff_B_3s0PRdKJ2_1),.dout(n1332),.clk(gclk));
	jnot g1269(.din(w_n1251_0[0]),.dout(n1333),.clk(gclk));
	jnot g1270(.din(w_n1322_0[0]),.dout(n1334),.clk(gclk));
	jor g1271(.dina(w_dff_B_RhxBNb8P7_0),.dinb(n1333),.dout(n1335),.clk(gclk));
	jor g1272(.dina(w_n1324_0[0]),.dinb(w_n1248_0[0]),.dout(n1336),.clk(gclk));
	jand g1273(.dina(n1336),.dinb(w_dff_B_xI4KtHss7_1),.dout(n1337),.clk(gclk));
	jand g1274(.dina(w_G528gat_5[2]),.dinb(w_G86gat_2[1]),.dout(n1338),.clk(gclk));
	jand g1275(.dina(w_n1320_0[0]),.dinb(w_n1256_0[0]),.dout(n1339),.clk(gclk));
	jand g1276(.dina(w_n1321_0[0]),.dinb(w_n1253_0[0]),.dout(n1340),.clk(gclk));
	jor g1277(.dina(n1340),.dinb(w_dff_B_Y7cEae5U1_1),.dout(n1341),.clk(gclk));
	jand g1278(.dina(w_G511gat_5[1]),.dinb(w_G103gat_2[2]),.dout(n1342),.clk(gclk));
	jnot g1279(.din(n1342),.dout(n1343),.clk(gclk));
	jand g1280(.dina(w_n1318_0[0]),.dinb(w_n1261_0[0]),.dout(n1344),.clk(gclk));
	jand g1281(.dina(w_n1319_0[0]),.dinb(w_n1258_0[0]),.dout(n1345),.clk(gclk));
	jor g1282(.dina(n1345),.dinb(w_dff_B_1csLnxFv0_1),.dout(n1346),.clk(gclk));
	jand g1283(.dina(w_G494gat_5[0]),.dinb(w_G120gat_3[0]),.dout(n1347),.clk(gclk));
	jnot g1284(.din(n1347),.dout(n1348),.clk(gclk));
	jand g1285(.dina(w_n1316_0[0]),.dinb(w_n1266_0[0]),.dout(n1349),.clk(gclk));
	jand g1286(.dina(w_n1317_0[0]),.dinb(w_n1263_0[0]),.dout(n1350),.clk(gclk));
	jor g1287(.dina(n1350),.dinb(w_dff_B_faBXe0Lc1_1),.dout(n1351),.clk(gclk));
	jand g1288(.dina(w_G477gat_4[2]),.dinb(w_G137gat_3[1]),.dout(n1352),.clk(gclk));
	jnot g1289(.din(n1352),.dout(n1353),.clk(gclk));
	jand g1290(.dina(w_n1314_0[0]),.dinb(w_n1271_0[0]),.dout(n1354),.clk(gclk));
	jand g1291(.dina(w_n1315_0[0]),.dinb(w_n1268_0[0]),.dout(n1355),.clk(gclk));
	jor g1292(.dina(n1355),.dinb(w_dff_B_sP4Ejq843_1),.dout(n1356),.clk(gclk));
	jand g1293(.dina(w_G460gat_4[1]),.dinb(w_G154gat_3[2]),.dout(n1357),.clk(gclk));
	jnot g1294(.din(n1357),.dout(n1358),.clk(gclk));
	jand g1295(.dina(w_n1312_0[0]),.dinb(w_n1276_0[0]),.dout(n1359),.clk(gclk));
	jand g1296(.dina(w_n1313_0[0]),.dinb(w_n1273_0[0]),.dout(n1360),.clk(gclk));
	jor g1297(.dina(n1360),.dinb(w_dff_B_WVn4gxIs4_1),.dout(n1361),.clk(gclk));
	jand g1298(.dina(w_G443gat_4[0]),.dinb(w_G171gat_4[0]),.dout(n1362),.clk(gclk));
	jnot g1299(.din(n1362),.dout(n1363),.clk(gclk));
	jand g1300(.dina(w_n1310_0[0]),.dinb(w_n1281_0[0]),.dout(n1364),.clk(gclk));
	jand g1301(.dina(w_n1311_0[0]),.dinb(w_n1278_0[0]),.dout(n1365),.clk(gclk));
	jor g1302(.dina(n1365),.dinb(w_dff_B_jkB5FMPY5_1),.dout(n1366),.clk(gclk));
	jand g1303(.dina(w_G426gat_3[2]),.dinb(w_G188gat_4[1]),.dout(n1367),.clk(gclk));
	jnot g1304(.din(n1367),.dout(n1368),.clk(gclk));
	jand g1305(.dina(w_n1308_0[0]),.dinb(w_n1286_0[0]),.dout(n1369),.clk(gclk));
	jand g1306(.dina(w_n1309_0[0]),.dinb(w_n1283_0[0]),.dout(n1370),.clk(gclk));
	jor g1307(.dina(n1370),.dinb(w_dff_B_g4zIW2PC4_1),.dout(n1371),.clk(gclk));
	jand g1308(.dina(w_G409gat_3[1]),.dinb(w_G205gat_4[2]),.dout(n1372),.clk(gclk));
	jnot g1309(.din(n1372),.dout(n1373),.clk(gclk));
	jand g1310(.dina(w_n1306_0[0]),.dinb(w_n1291_0[0]),.dout(n1374),.clk(gclk));
	jand g1311(.dina(w_n1307_0[0]),.dinb(w_n1288_0[0]),.dout(n1375),.clk(gclk));
	jor g1312(.dina(n1375),.dinb(w_dff_B_f3NceXEh7_1),.dout(n1376),.clk(gclk));
	jand g1313(.dina(w_G392gat_3[0]),.dinb(w_G222gat_5[0]),.dout(n1377),.clk(gclk));
	jnot g1314(.din(n1377),.dout(n1378),.clk(gclk));
	jand g1315(.dina(w_n1304_0[0]),.dinb(w_n1296_0[0]),.dout(n1379),.clk(gclk));
	jand g1316(.dina(w_n1305_0[0]),.dinb(w_n1293_0[0]),.dout(n1380),.clk(gclk));
	jor g1317(.dina(n1380),.dinb(w_dff_B_8PWg07E36_1),.dout(n1381),.clk(gclk));
	jand g1318(.dina(w_G375gat_2[2]),.dinb(w_G239gat_5[1]),.dout(n1382),.clk(gclk));
	jand g1319(.dina(w_G358gat_2[1]),.dinb(w_G256gat_5[2]),.dout(n1383),.clk(gclk));
	jor g1320(.dina(w_n1301_0[0]),.dinb(w_n1298_0[0]),.dout(n1384),.clk(gclk));
	jor g1321(.dina(w_n1303_0[0]),.dinb(w_n1297_0[0]),.dout(n1385),.clk(gclk));
	jand g1322(.dina(n1385),.dinb(w_dff_B_OLZWrOjp4_1),.dout(n1386),.clk(gclk));
	jxor g1323(.dina(w_n1386_0[1]),.dinb(w_n1383_0[1]),.dout(n1387),.clk(gclk));
	jnot g1324(.din(n1387),.dout(n1388),.clk(gclk));
	jxor g1325(.dina(w_n1388_0[1]),.dinb(w_n1382_0[1]),.dout(n1389),.clk(gclk));
	jxor g1326(.dina(w_n1389_0[1]),.dinb(w_n1381_0[1]),.dout(n1390),.clk(gclk));
	jxor g1327(.dina(w_n1390_0[1]),.dinb(w_n1378_0[1]),.dout(n1391),.clk(gclk));
	jxor g1328(.dina(w_n1391_0[1]),.dinb(w_n1376_0[1]),.dout(n1392),.clk(gclk));
	jxor g1329(.dina(w_n1392_0[1]),.dinb(w_n1373_0[1]),.dout(n1393),.clk(gclk));
	jxor g1330(.dina(w_n1393_0[1]),.dinb(w_n1371_0[1]),.dout(n1394),.clk(gclk));
	jxor g1331(.dina(w_n1394_0[1]),.dinb(w_n1368_0[1]),.dout(n1395),.clk(gclk));
	jxor g1332(.dina(w_n1395_0[1]),.dinb(w_n1366_0[1]),.dout(n1396),.clk(gclk));
	jxor g1333(.dina(w_n1396_0[1]),.dinb(w_n1363_0[1]),.dout(n1397),.clk(gclk));
	jxor g1334(.dina(w_n1397_0[1]),.dinb(w_n1361_0[1]),.dout(n1398),.clk(gclk));
	jxor g1335(.dina(w_n1398_0[1]),.dinb(w_n1358_0[1]),.dout(n1399),.clk(gclk));
	jxor g1336(.dina(w_n1399_0[1]),.dinb(w_n1356_0[1]),.dout(n1400),.clk(gclk));
	jxor g1337(.dina(w_n1400_0[1]),.dinb(w_n1353_0[1]),.dout(n1401),.clk(gclk));
	jxor g1338(.dina(w_n1401_0[1]),.dinb(w_n1351_0[1]),.dout(n1402),.clk(gclk));
	jxor g1339(.dina(w_n1402_0[1]),.dinb(w_n1348_0[1]),.dout(n1403),.clk(gclk));
	jxor g1340(.dina(w_n1403_0[1]),.dinb(w_n1346_0[1]),.dout(n1404),.clk(gclk));
	jxor g1341(.dina(w_n1404_0[1]),.dinb(w_n1343_0[1]),.dout(n1405),.clk(gclk));
	jxor g1342(.dina(w_n1405_0[1]),.dinb(w_n1341_0[1]),.dout(n1406),.clk(gclk));
	jnot g1343(.din(n1406),.dout(n1407),.clk(gclk));
	jxor g1344(.dina(w_n1407_0[1]),.dinb(w_n1338_0[1]),.dout(n1408),.clk(gclk));
	jnot g1345(.din(n1408),.dout(n1409),.clk(gclk));
	jxor g1346(.dina(w_n1409_0[1]),.dinb(w_n1337_0[1]),.dout(n1410),.clk(gclk));
	jxor g1347(.dina(w_n1410_0[1]),.dinb(w_n1332_0[1]),.dout(w_dff_A_0iZHqm6h1_2),.clk(gclk));
	jor g1348(.dina(w_n1409_0[0]),.dinb(w_n1337_0[0]),.dout(n1412),.clk(gclk));
	jnot g1349(.din(w_n1410_0[0]),.dout(n1413),.clk(gclk));
	jor g1350(.dina(w_dff_B_RMHEEMGh8_0),.dinb(w_n1332_0[0]),.dout(n1414),.clk(gclk));
	jand g1351(.dina(n1414),.dinb(w_dff_B_WWr6rpmz9_1),.dout(n1415),.clk(gclk));
	jnot g1352(.din(w_n1341_0[0]),.dout(n1416),.clk(gclk));
	jnot g1353(.din(w_n1405_0[0]),.dout(n1417),.clk(gclk));
	jor g1354(.dina(n1417),.dinb(n1416),.dout(n1418),.clk(gclk));
	jor g1355(.dina(w_n1407_0[0]),.dinb(w_n1338_0[0]),.dout(n1419),.clk(gclk));
	jand g1356(.dina(n1419),.dinb(w_dff_B_2YkkQ9rd3_1),.dout(n1420),.clk(gclk));
	jand g1357(.dina(w_G528gat_5[1]),.dinb(w_G103gat_2[1]),.dout(n1421),.clk(gclk));
	jand g1358(.dina(w_n1403_0[0]),.dinb(w_n1346_0[0]),.dout(n1422),.clk(gclk));
	jand g1359(.dina(w_n1404_0[0]),.dinb(w_n1343_0[0]),.dout(n1423),.clk(gclk));
	jor g1360(.dina(n1423),.dinb(w_dff_B_sIuJ0ldn2_1),.dout(n1424),.clk(gclk));
	jand g1361(.dina(w_G511gat_5[0]),.dinb(w_G120gat_2[2]),.dout(n1425),.clk(gclk));
	jnot g1362(.din(n1425),.dout(n1426),.clk(gclk));
	jand g1363(.dina(w_n1401_0[0]),.dinb(w_n1351_0[0]),.dout(n1427),.clk(gclk));
	jand g1364(.dina(w_n1402_0[0]),.dinb(w_n1348_0[0]),.dout(n1428),.clk(gclk));
	jor g1365(.dina(n1428),.dinb(w_dff_B_GNK67qew6_1),.dout(n1429),.clk(gclk));
	jand g1366(.dina(w_G494gat_4[2]),.dinb(w_G137gat_3[0]),.dout(n1430),.clk(gclk));
	jnot g1367(.din(n1430),.dout(n1431),.clk(gclk));
	jand g1368(.dina(w_n1399_0[0]),.dinb(w_n1356_0[0]),.dout(n1432),.clk(gclk));
	jand g1369(.dina(w_n1400_0[0]),.dinb(w_n1353_0[0]),.dout(n1433),.clk(gclk));
	jor g1370(.dina(n1433),.dinb(w_dff_B_NTWXxtiL6_1),.dout(n1434),.clk(gclk));
	jand g1371(.dina(w_G477gat_4[1]),.dinb(w_G154gat_3[1]),.dout(n1435),.clk(gclk));
	jnot g1372(.din(n1435),.dout(n1436),.clk(gclk));
	jand g1373(.dina(w_n1397_0[0]),.dinb(w_n1361_0[0]),.dout(n1437),.clk(gclk));
	jand g1374(.dina(w_n1398_0[0]),.dinb(w_n1358_0[0]),.dout(n1438),.clk(gclk));
	jor g1375(.dina(n1438),.dinb(w_dff_B_bc8EOeQJ5_1),.dout(n1439),.clk(gclk));
	jand g1376(.dina(w_G460gat_4[0]),.dinb(w_G171gat_3[2]),.dout(n1440),.clk(gclk));
	jnot g1377(.din(n1440),.dout(n1441),.clk(gclk));
	jand g1378(.dina(w_n1395_0[0]),.dinb(w_n1366_0[0]),.dout(n1442),.clk(gclk));
	jand g1379(.dina(w_n1396_0[0]),.dinb(w_n1363_0[0]),.dout(n1443),.clk(gclk));
	jor g1380(.dina(n1443),.dinb(w_dff_B_0Ke26RMA9_1),.dout(n1444),.clk(gclk));
	jand g1381(.dina(w_G443gat_3[2]),.dinb(w_G188gat_4[0]),.dout(n1445),.clk(gclk));
	jnot g1382(.din(n1445),.dout(n1446),.clk(gclk));
	jand g1383(.dina(w_n1393_0[0]),.dinb(w_n1371_0[0]),.dout(n1447),.clk(gclk));
	jand g1384(.dina(w_n1394_0[0]),.dinb(w_n1368_0[0]),.dout(n1448),.clk(gclk));
	jor g1385(.dina(n1448),.dinb(w_dff_B_DeIbx7lP9_1),.dout(n1449),.clk(gclk));
	jand g1386(.dina(w_G426gat_3[1]),.dinb(w_G205gat_4[1]),.dout(n1450),.clk(gclk));
	jnot g1387(.din(n1450),.dout(n1451),.clk(gclk));
	jand g1388(.dina(w_n1391_0[0]),.dinb(w_n1376_0[0]),.dout(n1452),.clk(gclk));
	jand g1389(.dina(w_n1392_0[0]),.dinb(w_n1373_0[0]),.dout(n1453),.clk(gclk));
	jor g1390(.dina(n1453),.dinb(w_dff_B_QsPz98oR1_1),.dout(n1454),.clk(gclk));
	jand g1391(.dina(w_G409gat_3[0]),.dinb(w_G222gat_4[2]),.dout(n1455),.clk(gclk));
	jnot g1392(.din(n1455),.dout(n1456),.clk(gclk));
	jand g1393(.dina(w_n1389_0[0]),.dinb(w_n1381_0[0]),.dout(n1457),.clk(gclk));
	jand g1394(.dina(w_n1390_0[0]),.dinb(w_n1378_0[0]),.dout(n1458),.clk(gclk));
	jor g1395(.dina(n1458),.dinb(w_dff_B_QnmaqLHI3_1),.dout(n1459),.clk(gclk));
	jand g1396(.dina(w_G392gat_2[2]),.dinb(w_G239gat_5[0]),.dout(n1460),.clk(gclk));
	jand g1397(.dina(w_G375gat_2[1]),.dinb(w_G256gat_5[1]),.dout(n1461),.clk(gclk));
	jor g1398(.dina(w_n1386_0[0]),.dinb(w_n1383_0[0]),.dout(n1462),.clk(gclk));
	jor g1399(.dina(w_n1388_0[0]),.dinb(w_n1382_0[0]),.dout(n1463),.clk(gclk));
	jand g1400(.dina(n1463),.dinb(w_dff_B_RSFFa2ch4_1),.dout(n1464),.clk(gclk));
	jxor g1401(.dina(w_n1464_0[1]),.dinb(w_n1461_0[1]),.dout(n1465),.clk(gclk));
	jnot g1402(.din(n1465),.dout(n1466),.clk(gclk));
	jxor g1403(.dina(w_n1466_0[1]),.dinb(w_n1460_0[1]),.dout(n1467),.clk(gclk));
	jxor g1404(.dina(w_n1467_0[1]),.dinb(w_n1459_0[1]),.dout(n1468),.clk(gclk));
	jxor g1405(.dina(w_n1468_0[1]),.dinb(w_n1456_0[1]),.dout(n1469),.clk(gclk));
	jxor g1406(.dina(w_n1469_0[1]),.dinb(w_n1454_0[1]),.dout(n1470),.clk(gclk));
	jxor g1407(.dina(w_n1470_0[1]),.dinb(w_n1451_0[1]),.dout(n1471),.clk(gclk));
	jxor g1408(.dina(w_n1471_0[1]),.dinb(w_n1449_0[1]),.dout(n1472),.clk(gclk));
	jxor g1409(.dina(w_n1472_0[1]),.dinb(w_n1446_0[1]),.dout(n1473),.clk(gclk));
	jxor g1410(.dina(w_n1473_0[1]),.dinb(w_n1444_0[1]),.dout(n1474),.clk(gclk));
	jxor g1411(.dina(w_n1474_0[1]),.dinb(w_n1441_0[1]),.dout(n1475),.clk(gclk));
	jxor g1412(.dina(w_n1475_0[1]),.dinb(w_n1439_0[1]),.dout(n1476),.clk(gclk));
	jxor g1413(.dina(w_n1476_0[1]),.dinb(w_n1436_0[1]),.dout(n1477),.clk(gclk));
	jxor g1414(.dina(w_n1477_0[1]),.dinb(w_n1434_0[1]),.dout(n1478),.clk(gclk));
	jxor g1415(.dina(w_n1478_0[1]),.dinb(w_n1431_0[1]),.dout(n1479),.clk(gclk));
	jxor g1416(.dina(w_n1479_0[1]),.dinb(w_n1429_0[1]),.dout(n1480),.clk(gclk));
	jxor g1417(.dina(w_n1480_0[1]),.dinb(w_n1426_0[1]),.dout(n1481),.clk(gclk));
	jxor g1418(.dina(w_n1481_0[1]),.dinb(w_n1424_0[1]),.dout(n1482),.clk(gclk));
	jnot g1419(.din(n1482),.dout(n1483),.clk(gclk));
	jxor g1420(.dina(w_n1483_0[1]),.dinb(w_n1421_0[1]),.dout(n1484),.clk(gclk));
	jnot g1421(.din(n1484),.dout(n1485),.clk(gclk));
	jxor g1422(.dina(w_n1485_0[1]),.dinb(w_n1420_0[1]),.dout(n1486),.clk(gclk));
	jxor g1423(.dina(w_n1486_0[1]),.dinb(w_n1415_0[1]),.dout(w_dff_A_DbIDePej4_2),.clk(gclk));
	jor g1424(.dina(w_n1485_0[0]),.dinb(w_n1420_0[0]),.dout(n1488),.clk(gclk));
	jnot g1425(.din(w_n1486_0[0]),.dout(n1489),.clk(gclk));
	jor g1426(.dina(w_dff_B_fW2lPW9w3_0),.dinb(w_n1415_0[0]),.dout(n1490),.clk(gclk));
	jand g1427(.dina(n1490),.dinb(w_dff_B_uM7kyvMl1_1),.dout(n1491),.clk(gclk));
	jnot g1428(.din(w_n1424_0[0]),.dout(n1492),.clk(gclk));
	jnot g1429(.din(w_n1481_0[0]),.dout(n1493),.clk(gclk));
	jor g1430(.dina(n1493),.dinb(n1492),.dout(n1494),.clk(gclk));
	jor g1431(.dina(w_n1483_0[0]),.dinb(w_n1421_0[0]),.dout(n1495),.clk(gclk));
	jand g1432(.dina(n1495),.dinb(w_dff_B_RRuD0sth9_1),.dout(n1496),.clk(gclk));
	jand g1433(.dina(w_G528gat_5[0]),.dinb(w_G120gat_2[1]),.dout(n1497),.clk(gclk));
	jand g1434(.dina(w_n1479_0[0]),.dinb(w_n1429_0[0]),.dout(n1498),.clk(gclk));
	jand g1435(.dina(w_n1480_0[0]),.dinb(w_n1426_0[0]),.dout(n1499),.clk(gclk));
	jor g1436(.dina(n1499),.dinb(w_dff_B_lQf6csxZ2_1),.dout(n1500),.clk(gclk));
	jand g1437(.dina(w_G511gat_4[2]),.dinb(w_G137gat_2[2]),.dout(n1501),.clk(gclk));
	jnot g1438(.din(n1501),.dout(n1502),.clk(gclk));
	jand g1439(.dina(w_n1477_0[0]),.dinb(w_n1434_0[0]),.dout(n1503),.clk(gclk));
	jand g1440(.dina(w_n1478_0[0]),.dinb(w_n1431_0[0]),.dout(n1504),.clk(gclk));
	jor g1441(.dina(n1504),.dinb(w_dff_B_t36JFZHW4_1),.dout(n1505),.clk(gclk));
	jand g1442(.dina(w_G494gat_4[1]),.dinb(w_G154gat_3[0]),.dout(n1506),.clk(gclk));
	jnot g1443(.din(n1506),.dout(n1507),.clk(gclk));
	jand g1444(.dina(w_n1475_0[0]),.dinb(w_n1439_0[0]),.dout(n1508),.clk(gclk));
	jand g1445(.dina(w_n1476_0[0]),.dinb(w_n1436_0[0]),.dout(n1509),.clk(gclk));
	jor g1446(.dina(n1509),.dinb(w_dff_B_ep9J85lm5_1),.dout(n1510),.clk(gclk));
	jand g1447(.dina(w_G477gat_4[0]),.dinb(w_G171gat_3[1]),.dout(n1511),.clk(gclk));
	jnot g1448(.din(n1511),.dout(n1512),.clk(gclk));
	jand g1449(.dina(w_n1473_0[0]),.dinb(w_n1444_0[0]),.dout(n1513),.clk(gclk));
	jand g1450(.dina(w_n1474_0[0]),.dinb(w_n1441_0[0]),.dout(n1514),.clk(gclk));
	jor g1451(.dina(n1514),.dinb(w_dff_B_QlXDA0Gs6_1),.dout(n1515),.clk(gclk));
	jand g1452(.dina(w_G460gat_3[2]),.dinb(w_G188gat_3[2]),.dout(n1516),.clk(gclk));
	jnot g1453(.din(n1516),.dout(n1517),.clk(gclk));
	jand g1454(.dina(w_n1471_0[0]),.dinb(w_n1449_0[0]),.dout(n1518),.clk(gclk));
	jand g1455(.dina(w_n1472_0[0]),.dinb(w_n1446_0[0]),.dout(n1519),.clk(gclk));
	jor g1456(.dina(n1519),.dinb(w_dff_B_u5IVoq2a4_1),.dout(n1520),.clk(gclk));
	jand g1457(.dina(w_G443gat_3[1]),.dinb(w_G205gat_4[0]),.dout(n1521),.clk(gclk));
	jnot g1458(.din(n1521),.dout(n1522),.clk(gclk));
	jand g1459(.dina(w_n1469_0[0]),.dinb(w_n1454_0[0]),.dout(n1523),.clk(gclk));
	jand g1460(.dina(w_n1470_0[0]),.dinb(w_n1451_0[0]),.dout(n1524),.clk(gclk));
	jor g1461(.dina(n1524),.dinb(w_dff_B_TCdl79rD8_1),.dout(n1525),.clk(gclk));
	jand g1462(.dina(w_G426gat_3[0]),.dinb(w_G222gat_4[1]),.dout(n1526),.clk(gclk));
	jnot g1463(.din(n1526),.dout(n1527),.clk(gclk));
	jand g1464(.dina(w_n1467_0[0]),.dinb(w_n1459_0[0]),.dout(n1528),.clk(gclk));
	jand g1465(.dina(w_n1468_0[0]),.dinb(w_n1456_0[0]),.dout(n1529),.clk(gclk));
	jor g1466(.dina(n1529),.dinb(w_dff_B_4ZGyLYI34_1),.dout(n1530),.clk(gclk));
	jand g1467(.dina(w_G409gat_2[2]),.dinb(w_G239gat_4[2]),.dout(n1531),.clk(gclk));
	jand g1468(.dina(w_G392gat_2[1]),.dinb(w_G256gat_5[0]),.dout(n1532),.clk(gclk));
	jor g1469(.dina(w_n1464_0[0]),.dinb(w_n1461_0[0]),.dout(n1533),.clk(gclk));
	jor g1470(.dina(w_n1466_0[0]),.dinb(w_n1460_0[0]),.dout(n1534),.clk(gclk));
	jand g1471(.dina(n1534),.dinb(w_dff_B_2ezTw40N3_1),.dout(n1535),.clk(gclk));
	jxor g1472(.dina(w_n1535_0[1]),.dinb(w_n1532_0[1]),.dout(n1536),.clk(gclk));
	jnot g1473(.din(n1536),.dout(n1537),.clk(gclk));
	jxor g1474(.dina(w_n1537_0[1]),.dinb(w_n1531_0[1]),.dout(n1538),.clk(gclk));
	jxor g1475(.dina(w_n1538_0[1]),.dinb(w_n1530_0[1]),.dout(n1539),.clk(gclk));
	jxor g1476(.dina(w_n1539_0[1]),.dinb(w_n1527_0[1]),.dout(n1540),.clk(gclk));
	jxor g1477(.dina(w_n1540_0[1]),.dinb(w_n1525_0[1]),.dout(n1541),.clk(gclk));
	jxor g1478(.dina(w_n1541_0[1]),.dinb(w_n1522_0[1]),.dout(n1542),.clk(gclk));
	jxor g1479(.dina(w_n1542_0[1]),.dinb(w_n1520_0[1]),.dout(n1543),.clk(gclk));
	jxor g1480(.dina(w_n1543_0[1]),.dinb(w_n1517_0[1]),.dout(n1544),.clk(gclk));
	jxor g1481(.dina(w_n1544_0[1]),.dinb(w_n1515_0[1]),.dout(n1545),.clk(gclk));
	jxor g1482(.dina(w_n1545_0[1]),.dinb(w_n1512_0[1]),.dout(n1546),.clk(gclk));
	jxor g1483(.dina(w_n1546_0[1]),.dinb(w_n1510_0[1]),.dout(n1547),.clk(gclk));
	jxor g1484(.dina(w_n1547_0[1]),.dinb(w_n1507_0[1]),.dout(n1548),.clk(gclk));
	jxor g1485(.dina(w_n1548_0[1]),.dinb(w_n1505_0[1]),.dout(n1549),.clk(gclk));
	jxor g1486(.dina(w_n1549_0[1]),.dinb(w_n1502_0[1]),.dout(n1550),.clk(gclk));
	jxor g1487(.dina(w_n1550_0[1]),.dinb(w_n1500_0[1]),.dout(n1551),.clk(gclk));
	jnot g1488(.din(n1551),.dout(n1552),.clk(gclk));
	jxor g1489(.dina(w_n1552_0[1]),.dinb(w_n1497_0[1]),.dout(n1553),.clk(gclk));
	jnot g1490(.din(n1553),.dout(n1554),.clk(gclk));
	jxor g1491(.dina(w_n1554_0[1]),.dinb(w_n1496_0[1]),.dout(n1555),.clk(gclk));
	jxor g1492(.dina(w_n1555_0[1]),.dinb(w_n1491_0[1]),.dout(w_dff_A_IUYnNff39_2),.clk(gclk));
	jor g1493(.dina(w_n1554_0[0]),.dinb(w_n1496_0[0]),.dout(n1557),.clk(gclk));
	jnot g1494(.din(w_n1555_0[0]),.dout(n1558),.clk(gclk));
	jor g1495(.dina(w_dff_B_qqrw33Vf4_0),.dinb(w_n1491_0[0]),.dout(n1559),.clk(gclk));
	jand g1496(.dina(n1559),.dinb(w_dff_B_PaiXs0mt7_1),.dout(n1560),.clk(gclk));
	jnot g1497(.din(w_n1500_0[0]),.dout(n1561),.clk(gclk));
	jnot g1498(.din(w_n1550_0[0]),.dout(n1562),.clk(gclk));
	jor g1499(.dina(w_dff_B_xVbS7BIv1_0),.dinb(n1561),.dout(n1563),.clk(gclk));
	jor g1500(.dina(w_n1552_0[0]),.dinb(w_n1497_0[0]),.dout(n1564),.clk(gclk));
	jand g1501(.dina(n1564),.dinb(w_dff_B_dscEN8CP3_1),.dout(n1565),.clk(gclk));
	jand g1502(.dina(w_G528gat_4[2]),.dinb(w_G137gat_2[1]),.dout(n1566),.clk(gclk));
	jand g1503(.dina(w_n1548_0[0]),.dinb(w_n1505_0[0]),.dout(n1567),.clk(gclk));
	jand g1504(.dina(w_n1549_0[0]),.dinb(w_n1502_0[0]),.dout(n1568),.clk(gclk));
	jor g1505(.dina(n1568),.dinb(w_dff_B_ewia6aDz7_1),.dout(n1569),.clk(gclk));
	jand g1506(.dina(w_G511gat_4[1]),.dinb(w_G154gat_2[2]),.dout(n1570),.clk(gclk));
	jnot g1507(.din(n1570),.dout(n1571),.clk(gclk));
	jand g1508(.dina(w_n1546_0[0]),.dinb(w_n1510_0[0]),.dout(n1572),.clk(gclk));
	jand g1509(.dina(w_n1547_0[0]),.dinb(w_n1507_0[0]),.dout(n1573),.clk(gclk));
	jor g1510(.dina(n1573),.dinb(w_dff_B_OVFaeoJQ4_1),.dout(n1574),.clk(gclk));
	jand g1511(.dina(w_G494gat_4[0]),.dinb(w_G171gat_3[0]),.dout(n1575),.clk(gclk));
	jnot g1512(.din(n1575),.dout(n1576),.clk(gclk));
	jand g1513(.dina(w_n1544_0[0]),.dinb(w_n1515_0[0]),.dout(n1577),.clk(gclk));
	jand g1514(.dina(w_n1545_0[0]),.dinb(w_n1512_0[0]),.dout(n1578),.clk(gclk));
	jor g1515(.dina(n1578),.dinb(w_dff_B_KWsj1w4I1_1),.dout(n1579),.clk(gclk));
	jand g1516(.dina(w_G477gat_3[2]),.dinb(w_G188gat_3[1]),.dout(n1580),.clk(gclk));
	jnot g1517(.din(n1580),.dout(n1581),.clk(gclk));
	jand g1518(.dina(w_n1542_0[0]),.dinb(w_n1520_0[0]),.dout(n1582),.clk(gclk));
	jand g1519(.dina(w_n1543_0[0]),.dinb(w_n1517_0[0]),.dout(n1583),.clk(gclk));
	jor g1520(.dina(n1583),.dinb(w_dff_B_8o2FsipG4_1),.dout(n1584),.clk(gclk));
	jand g1521(.dina(w_G460gat_3[1]),.dinb(w_G205gat_3[2]),.dout(n1585),.clk(gclk));
	jnot g1522(.din(n1585),.dout(n1586),.clk(gclk));
	jand g1523(.dina(w_n1540_0[0]),.dinb(w_n1525_0[0]),.dout(n1587),.clk(gclk));
	jand g1524(.dina(w_n1541_0[0]),.dinb(w_n1522_0[0]),.dout(n1588),.clk(gclk));
	jor g1525(.dina(n1588),.dinb(w_dff_B_SAOoRhsC9_1),.dout(n1589),.clk(gclk));
	jand g1526(.dina(w_G443gat_3[0]),.dinb(w_G222gat_4[0]),.dout(n1590),.clk(gclk));
	jnot g1527(.din(n1590),.dout(n1591),.clk(gclk));
	jand g1528(.dina(w_n1538_0[0]),.dinb(w_n1530_0[0]),.dout(n1592),.clk(gclk));
	jand g1529(.dina(w_n1539_0[0]),.dinb(w_n1527_0[0]),.dout(n1593),.clk(gclk));
	jor g1530(.dina(n1593),.dinb(w_dff_B_McwKnVtr5_1),.dout(n1594),.clk(gclk));
	jand g1531(.dina(w_G426gat_2[2]),.dinb(w_G239gat_4[1]),.dout(n1595),.clk(gclk));
	jand g1532(.dina(w_G409gat_2[1]),.dinb(w_G256gat_4[2]),.dout(n1596),.clk(gclk));
	jor g1533(.dina(w_n1535_0[0]),.dinb(w_n1532_0[0]),.dout(n1597),.clk(gclk));
	jor g1534(.dina(w_n1537_0[0]),.dinb(w_n1531_0[0]),.dout(n1598),.clk(gclk));
	jand g1535(.dina(n1598),.dinb(w_dff_B_F8seNExg6_1),.dout(n1599),.clk(gclk));
	jxor g1536(.dina(w_n1599_0[1]),.dinb(w_n1596_0[1]),.dout(n1600),.clk(gclk));
	jnot g1537(.din(n1600),.dout(n1601),.clk(gclk));
	jxor g1538(.dina(w_n1601_0[1]),.dinb(w_n1595_0[1]),.dout(n1602),.clk(gclk));
	jxor g1539(.dina(w_n1602_0[1]),.dinb(w_n1594_0[1]),.dout(n1603),.clk(gclk));
	jxor g1540(.dina(w_n1603_0[1]),.dinb(w_n1591_0[1]),.dout(n1604),.clk(gclk));
	jxor g1541(.dina(w_n1604_0[1]),.dinb(w_n1589_0[1]),.dout(n1605),.clk(gclk));
	jxor g1542(.dina(w_n1605_0[1]),.dinb(w_n1586_0[1]),.dout(n1606),.clk(gclk));
	jxor g1543(.dina(w_n1606_0[1]),.dinb(w_n1584_0[1]),.dout(n1607),.clk(gclk));
	jxor g1544(.dina(w_n1607_0[1]),.dinb(w_n1581_0[1]),.dout(n1608),.clk(gclk));
	jxor g1545(.dina(w_n1608_0[1]),.dinb(w_n1579_0[1]),.dout(n1609),.clk(gclk));
	jxor g1546(.dina(w_n1609_0[1]),.dinb(w_n1576_0[1]),.dout(n1610),.clk(gclk));
	jxor g1547(.dina(w_n1610_0[1]),.dinb(w_n1574_0[1]),.dout(n1611),.clk(gclk));
	jxor g1548(.dina(w_n1611_0[1]),.dinb(w_n1571_0[1]),.dout(n1612),.clk(gclk));
	jxor g1549(.dina(w_n1612_0[1]),.dinb(w_n1569_0[1]),.dout(n1613),.clk(gclk));
	jnot g1550(.din(n1613),.dout(n1614),.clk(gclk));
	jxor g1551(.dina(w_n1614_0[1]),.dinb(w_n1566_0[1]),.dout(n1615),.clk(gclk));
	jnot g1552(.din(n1615),.dout(n1616),.clk(gclk));
	jxor g1553(.dina(w_n1616_0[1]),.dinb(w_n1565_0[1]),.dout(n1617),.clk(gclk));
	jxor g1554(.dina(w_n1617_0[1]),.dinb(w_n1560_0[1]),.dout(w_dff_A_bLrqy25k9_2),.clk(gclk));
	jor g1555(.dina(w_n1616_0[0]),.dinb(w_n1565_0[0]),.dout(n1619),.clk(gclk));
	jnot g1556(.din(w_n1617_0[0]),.dout(n1620),.clk(gclk));
	jor g1557(.dina(w_dff_B_UtgNrEWs9_0),.dinb(w_n1560_0[0]),.dout(n1621),.clk(gclk));
	jand g1558(.dina(n1621),.dinb(w_dff_B_LL8oMdvo3_1),.dout(n1622),.clk(gclk));
	jnot g1559(.din(w_n1569_0[0]),.dout(n1623),.clk(gclk));
	jnot g1560(.din(w_n1612_0[0]),.dout(n1624),.clk(gclk));
	jor g1561(.dina(n1624),.dinb(n1623),.dout(n1625),.clk(gclk));
	jor g1562(.dina(w_n1614_0[0]),.dinb(w_n1566_0[0]),.dout(n1626),.clk(gclk));
	jand g1563(.dina(n1626),.dinb(w_dff_B_mP2VrqKQ6_1),.dout(n1627),.clk(gclk));
	jand g1564(.dina(w_G528gat_4[1]),.dinb(w_G154gat_2[1]),.dout(n1628),.clk(gclk));
	jand g1565(.dina(w_n1610_0[0]),.dinb(w_n1574_0[0]),.dout(n1629),.clk(gclk));
	jand g1566(.dina(w_n1611_0[0]),.dinb(w_n1571_0[0]),.dout(n1630),.clk(gclk));
	jor g1567(.dina(n1630),.dinb(w_dff_B_caV1Uciq4_1),.dout(n1631),.clk(gclk));
	jand g1568(.dina(w_G511gat_4[0]),.dinb(w_G171gat_2[2]),.dout(n1632),.clk(gclk));
	jnot g1569(.din(n1632),.dout(n1633),.clk(gclk));
	jand g1570(.dina(w_n1608_0[0]),.dinb(w_n1579_0[0]),.dout(n1634),.clk(gclk));
	jand g1571(.dina(w_n1609_0[0]),.dinb(w_n1576_0[0]),.dout(n1635),.clk(gclk));
	jor g1572(.dina(n1635),.dinb(w_dff_B_4DM503qx1_1),.dout(n1636),.clk(gclk));
	jand g1573(.dina(w_G494gat_3[2]),.dinb(w_G188gat_3[0]),.dout(n1637),.clk(gclk));
	jnot g1574(.din(n1637),.dout(n1638),.clk(gclk));
	jand g1575(.dina(w_n1606_0[0]),.dinb(w_n1584_0[0]),.dout(n1639),.clk(gclk));
	jand g1576(.dina(w_n1607_0[0]),.dinb(w_n1581_0[0]),.dout(n1640),.clk(gclk));
	jor g1577(.dina(n1640),.dinb(w_dff_B_jPDNsV4f5_1),.dout(n1641),.clk(gclk));
	jand g1578(.dina(w_G477gat_3[1]),.dinb(w_G205gat_3[1]),.dout(n1642),.clk(gclk));
	jnot g1579(.din(n1642),.dout(n1643),.clk(gclk));
	jand g1580(.dina(w_n1604_0[0]),.dinb(w_n1589_0[0]),.dout(n1644),.clk(gclk));
	jand g1581(.dina(w_n1605_0[0]),.dinb(w_n1586_0[0]),.dout(n1645),.clk(gclk));
	jor g1582(.dina(n1645),.dinb(w_dff_B_BceJ9HAg2_1),.dout(n1646),.clk(gclk));
	jand g1583(.dina(w_G460gat_3[0]),.dinb(w_G222gat_3[2]),.dout(n1647),.clk(gclk));
	jnot g1584(.din(n1647),.dout(n1648),.clk(gclk));
	jand g1585(.dina(w_n1602_0[0]),.dinb(w_n1594_0[0]),.dout(n1649),.clk(gclk));
	jand g1586(.dina(w_n1603_0[0]),.dinb(w_n1591_0[0]),.dout(n1650),.clk(gclk));
	jor g1587(.dina(n1650),.dinb(w_dff_B_PRIZboWh1_1),.dout(n1651),.clk(gclk));
	jand g1588(.dina(w_G443gat_2[2]),.dinb(w_G239gat_4[0]),.dout(n1652),.clk(gclk));
	jand g1589(.dina(w_G426gat_2[1]),.dinb(w_G256gat_4[1]),.dout(n1653),.clk(gclk));
	jor g1590(.dina(w_n1599_0[0]),.dinb(w_n1596_0[0]),.dout(n1654),.clk(gclk));
	jor g1591(.dina(w_n1601_0[0]),.dinb(w_n1595_0[0]),.dout(n1655),.clk(gclk));
	jand g1592(.dina(n1655),.dinb(w_dff_B_QnrhvDJ39_1),.dout(n1656),.clk(gclk));
	jxor g1593(.dina(w_n1656_0[1]),.dinb(w_n1653_0[1]),.dout(n1657),.clk(gclk));
	jnot g1594(.din(n1657),.dout(n1658),.clk(gclk));
	jxor g1595(.dina(w_n1658_0[1]),.dinb(w_n1652_0[1]),.dout(n1659),.clk(gclk));
	jxor g1596(.dina(w_n1659_0[1]),.dinb(w_n1651_0[1]),.dout(n1660),.clk(gclk));
	jxor g1597(.dina(w_n1660_0[1]),.dinb(w_n1648_0[1]),.dout(n1661),.clk(gclk));
	jxor g1598(.dina(w_n1661_0[1]),.dinb(w_n1646_0[1]),.dout(n1662),.clk(gclk));
	jxor g1599(.dina(w_n1662_0[1]),.dinb(w_n1643_0[1]),.dout(n1663),.clk(gclk));
	jxor g1600(.dina(w_n1663_0[1]),.dinb(w_n1641_0[1]),.dout(n1664),.clk(gclk));
	jxor g1601(.dina(w_n1664_0[1]),.dinb(w_n1638_0[1]),.dout(n1665),.clk(gclk));
	jxor g1602(.dina(w_n1665_0[1]),.dinb(w_n1636_0[1]),.dout(n1666),.clk(gclk));
	jxor g1603(.dina(w_n1666_0[1]),.dinb(w_n1633_0[1]),.dout(n1667),.clk(gclk));
	jxor g1604(.dina(w_n1667_0[1]),.dinb(w_n1631_0[1]),.dout(n1668),.clk(gclk));
	jnot g1605(.din(n1668),.dout(n1669),.clk(gclk));
	jxor g1606(.dina(w_n1669_0[1]),.dinb(w_n1628_0[1]),.dout(n1670),.clk(gclk));
	jnot g1607(.din(n1670),.dout(n1671),.clk(gclk));
	jxor g1608(.dina(w_n1671_0[1]),.dinb(w_n1627_0[1]),.dout(n1672),.clk(gclk));
	jxor g1609(.dina(w_n1672_0[1]),.dinb(w_n1622_0[1]),.dout(w_dff_A_LmfDc3mX7_2),.clk(gclk));
	jor g1610(.dina(w_n1671_0[0]),.dinb(w_n1627_0[0]),.dout(n1674),.clk(gclk));
	jnot g1611(.din(w_n1672_0[0]),.dout(n1675),.clk(gclk));
	jor g1612(.dina(w_dff_B_hwj8yCsY3_0),.dinb(w_n1622_0[0]),.dout(n1676),.clk(gclk));
	jand g1613(.dina(n1676),.dinb(w_dff_B_J3ei1HvP0_1),.dout(n1677),.clk(gclk));
	jnot g1614(.din(w_n1631_0[0]),.dout(n1678),.clk(gclk));
	jnot g1615(.din(w_n1667_0[0]),.dout(n1679),.clk(gclk));
	jor g1616(.dina(n1679),.dinb(w_dff_B_rqcdsL8S1_1),.dout(n1680),.clk(gclk));
	jor g1617(.dina(w_n1669_0[0]),.dinb(w_n1628_0[0]),.dout(n1681),.clk(gclk));
	jand g1618(.dina(n1681),.dinb(w_dff_B_VVOCdBKQ9_1),.dout(n1682),.clk(gclk));
	jand g1619(.dina(w_G528gat_4[0]),.dinb(w_G171gat_2[1]),.dout(n1683),.clk(gclk));
	jnot g1620(.din(n1683),.dout(n1684),.clk(gclk));
	jand g1621(.dina(w_n1665_0[0]),.dinb(w_n1636_0[0]),.dout(n1685),.clk(gclk));
	jand g1622(.dina(w_n1666_0[0]),.dinb(w_n1633_0[0]),.dout(n1686),.clk(gclk));
	jor g1623(.dina(n1686),.dinb(w_dff_B_OD8zsOFz3_1),.dout(n1687),.clk(gclk));
	jand g1624(.dina(w_G511gat_3[2]),.dinb(w_G188gat_2[2]),.dout(n1688),.clk(gclk));
	jnot g1625(.din(n1688),.dout(n1689),.clk(gclk));
	jand g1626(.dina(w_n1663_0[0]),.dinb(w_n1641_0[0]),.dout(n1690),.clk(gclk));
	jand g1627(.dina(w_n1664_0[0]),.dinb(w_n1638_0[0]),.dout(n1691),.clk(gclk));
	jor g1628(.dina(n1691),.dinb(w_dff_B_YNu2zp3w3_1),.dout(n1692),.clk(gclk));
	jand g1629(.dina(w_G494gat_3[1]),.dinb(w_G205gat_3[0]),.dout(n1693),.clk(gclk));
	jnot g1630(.din(n1693),.dout(n1694),.clk(gclk));
	jand g1631(.dina(w_n1661_0[0]),.dinb(w_n1646_0[0]),.dout(n1695),.clk(gclk));
	jand g1632(.dina(w_n1662_0[0]),.dinb(w_n1643_0[0]),.dout(n1696),.clk(gclk));
	jor g1633(.dina(n1696),.dinb(w_dff_B_IVGV1hWr7_1),.dout(n1697),.clk(gclk));
	jand g1634(.dina(w_G477gat_3[0]),.dinb(w_G222gat_3[1]),.dout(n1698),.clk(gclk));
	jnot g1635(.din(n1698),.dout(n1699),.clk(gclk));
	jand g1636(.dina(w_n1659_0[0]),.dinb(w_n1651_0[0]),.dout(n1700),.clk(gclk));
	jand g1637(.dina(w_n1660_0[0]),.dinb(w_n1648_0[0]),.dout(n1701),.clk(gclk));
	jor g1638(.dina(n1701),.dinb(w_dff_B_LD9XSOiS3_1),.dout(n1702),.clk(gclk));
	jand g1639(.dina(w_G460gat_2[2]),.dinb(w_G239gat_3[2]),.dout(n1703),.clk(gclk));
	jand g1640(.dina(w_G443gat_2[1]),.dinb(w_G256gat_4[0]),.dout(n1704),.clk(gclk));
	jor g1641(.dina(w_n1656_0[0]),.dinb(w_n1653_0[0]),.dout(n1705),.clk(gclk));
	jor g1642(.dina(w_n1658_0[0]),.dinb(w_n1652_0[0]),.dout(n1706),.clk(gclk));
	jand g1643(.dina(n1706),.dinb(w_dff_B_sl9LlNAT0_1),.dout(n1707),.clk(gclk));
	jxor g1644(.dina(w_n1707_0[1]),.dinb(w_n1704_0[1]),.dout(n1708),.clk(gclk));
	jnot g1645(.din(n1708),.dout(n1709),.clk(gclk));
	jxor g1646(.dina(w_n1709_0[1]),.dinb(w_n1703_0[1]),.dout(n1710),.clk(gclk));
	jxor g1647(.dina(w_n1710_0[1]),.dinb(w_n1702_0[1]),.dout(n1711),.clk(gclk));
	jxor g1648(.dina(w_n1711_0[1]),.dinb(w_n1699_0[1]),.dout(n1712),.clk(gclk));
	jxor g1649(.dina(w_n1712_0[1]),.dinb(w_n1697_0[1]),.dout(n1713),.clk(gclk));
	jxor g1650(.dina(w_n1713_0[1]),.dinb(w_n1694_0[1]),.dout(n1714),.clk(gclk));
	jxor g1651(.dina(w_n1714_0[1]),.dinb(w_n1692_0[1]),.dout(n1715),.clk(gclk));
	jxor g1652(.dina(w_n1715_0[1]),.dinb(w_n1689_0[1]),.dout(n1716),.clk(gclk));
	jxor g1653(.dina(w_n1716_0[1]),.dinb(w_n1687_0[1]),.dout(n1717),.clk(gclk));
	jxor g1654(.dina(w_n1717_0[1]),.dinb(w_n1684_0[1]),.dout(n1718),.clk(gclk));
	jnot g1655(.din(n1718),.dout(n1719),.clk(gclk));
	jxor g1656(.dina(w_n1719_0[1]),.dinb(w_n1682_0[1]),.dout(n1720),.clk(gclk));
	jxor g1657(.dina(w_n1720_0[1]),.dinb(w_n1677_0[1]),.dout(w_dff_A_hXEXHGJP4_2),.clk(gclk));
	jor g1658(.dina(w_n1719_0[0]),.dinb(w_n1682_0[0]),.dout(n1722),.clk(gclk));
	jnot g1659(.din(w_n1720_0[0]),.dout(n1723),.clk(gclk));
	jor g1660(.dina(w_dff_B_plAUKf9m5_0),.dinb(w_n1677_0[0]),.dout(n1724),.clk(gclk));
	jand g1661(.dina(n1724),.dinb(w_dff_B_j8qeHvjW3_1),.dout(n1725),.clk(gclk));
	jand g1662(.dina(w_n1716_0[0]),.dinb(w_n1687_0[0]),.dout(n1726),.clk(gclk));
	jand g1663(.dina(w_n1717_0[0]),.dinb(w_n1684_0[0]),.dout(n1727),.clk(gclk));
	jor g1664(.dina(n1727),.dinb(w_dff_B_ZNA61zx23_1),.dout(n1728),.clk(gclk));
	jand g1665(.dina(w_G528gat_3[2]),.dinb(w_G188gat_2[1]),.dout(n1729),.clk(gclk));
	jnot g1666(.din(n1729),.dout(n1730),.clk(gclk));
	jand g1667(.dina(w_n1714_0[0]),.dinb(w_n1692_0[0]),.dout(n1731),.clk(gclk));
	jand g1668(.dina(w_n1715_0[0]),.dinb(w_n1689_0[0]),.dout(n1732),.clk(gclk));
	jor g1669(.dina(n1732),.dinb(w_dff_B_cbqqkSOt3_1),.dout(n1733),.clk(gclk));
	jand g1670(.dina(w_G511gat_3[1]),.dinb(w_G205gat_2[2]),.dout(n1734),.clk(gclk));
	jnot g1671(.din(n1734),.dout(n1735),.clk(gclk));
	jand g1672(.dina(w_n1712_0[0]),.dinb(w_n1697_0[0]),.dout(n1736),.clk(gclk));
	jand g1673(.dina(w_n1713_0[0]),.dinb(w_n1694_0[0]),.dout(n1737),.clk(gclk));
	jor g1674(.dina(n1737),.dinb(w_dff_B_GBFhlqJt1_1),.dout(n1738),.clk(gclk));
	jand g1675(.dina(w_G494gat_3[0]),.dinb(w_G222gat_3[0]),.dout(n1739),.clk(gclk));
	jnot g1676(.din(n1739),.dout(n1740),.clk(gclk));
	jand g1677(.dina(w_n1710_0[0]),.dinb(w_n1702_0[0]),.dout(n1741),.clk(gclk));
	jand g1678(.dina(w_n1711_0[0]),.dinb(w_n1699_0[0]),.dout(n1742),.clk(gclk));
	jor g1679(.dina(n1742),.dinb(w_dff_B_UFVwRiwo2_1),.dout(n1743),.clk(gclk));
	jand g1680(.dina(w_G477gat_2[2]),.dinb(w_G239gat_3[1]),.dout(n1744),.clk(gclk));
	jand g1681(.dina(w_G460gat_2[1]),.dinb(w_G256gat_3[2]),.dout(n1745),.clk(gclk));
	jor g1682(.dina(w_n1707_0[0]),.dinb(w_n1704_0[0]),.dout(n1746),.clk(gclk));
	jor g1683(.dina(w_n1709_0[0]),.dinb(w_n1703_0[0]),.dout(n1747),.clk(gclk));
	jand g1684(.dina(n1747),.dinb(w_dff_B_ITq5ODvv5_1),.dout(n1748),.clk(gclk));
	jxor g1685(.dina(w_n1748_0[1]),.dinb(w_n1745_0[1]),.dout(n1749),.clk(gclk));
	jnot g1686(.din(n1749),.dout(n1750),.clk(gclk));
	jxor g1687(.dina(w_n1750_0[1]),.dinb(w_n1744_0[1]),.dout(n1751),.clk(gclk));
	jxor g1688(.dina(w_n1751_0[1]),.dinb(w_n1743_0[1]),.dout(n1752),.clk(gclk));
	jxor g1689(.dina(w_n1752_0[1]),.dinb(w_n1740_0[1]),.dout(n1753),.clk(gclk));
	jxor g1690(.dina(w_n1753_0[1]),.dinb(w_n1738_0[1]),.dout(n1754),.clk(gclk));
	jxor g1691(.dina(w_n1754_0[1]),.dinb(w_n1735_0[1]),.dout(n1755),.clk(gclk));
	jxor g1692(.dina(w_n1755_0[1]),.dinb(w_n1733_0[1]),.dout(n1756),.clk(gclk));
	jxor g1693(.dina(w_n1756_0[1]),.dinb(w_n1730_0[1]),.dout(n1757),.clk(gclk));
	jxor g1694(.dina(w_n1757_0[1]),.dinb(w_n1728_0[1]),.dout(n1758),.clk(gclk));
	jxor g1695(.dina(w_n1758_0[1]),.dinb(w_n1725_0[1]),.dout(w_dff_A_3iLVSEwm9_2),.clk(gclk));
	jnot g1696(.din(w_n1728_0[0]),.dout(n1760),.clk(gclk));
	jnot g1697(.din(w_n1757_0[0]),.dout(n1761),.clk(gclk));
	jor g1698(.dina(n1761),.dinb(w_dff_B_TCewL5c97_1),.dout(n1762),.clk(gclk));
	jnot g1699(.din(w_n1758_0[0]),.dout(n1763),.clk(gclk));
	jor g1700(.dina(w_dff_B_pS6Cq4dI7_0),.dinb(w_n1725_0[0]),.dout(n1764),.clk(gclk));
	jand g1701(.dina(n1764),.dinb(w_dff_B_wn5H5gc59_1),.dout(n1765),.clk(gclk));
	jand g1702(.dina(w_n1755_0[0]),.dinb(w_n1733_0[0]),.dout(n1766),.clk(gclk));
	jand g1703(.dina(w_n1756_0[0]),.dinb(w_n1730_0[0]),.dout(n1767),.clk(gclk));
	jor g1704(.dina(n1767),.dinb(w_dff_B_LzPbpWEu3_1),.dout(n1768),.clk(gclk));
	jand g1705(.dina(w_G528gat_3[1]),.dinb(w_G205gat_2[1]),.dout(n1769),.clk(gclk));
	jnot g1706(.din(n1769),.dout(n1770),.clk(gclk));
	jand g1707(.dina(w_n1753_0[0]),.dinb(w_n1738_0[0]),.dout(n1771),.clk(gclk));
	jand g1708(.dina(w_n1754_0[0]),.dinb(w_n1735_0[0]),.dout(n1772),.clk(gclk));
	jor g1709(.dina(n1772),.dinb(w_dff_B_b90Z7vXn8_1),.dout(n1773),.clk(gclk));
	jand g1710(.dina(w_G511gat_3[0]),.dinb(w_G222gat_2[2]),.dout(n1774),.clk(gclk));
	jnot g1711(.din(n1774),.dout(n1775),.clk(gclk));
	jand g1712(.dina(w_n1751_0[0]),.dinb(w_n1743_0[0]),.dout(n1776),.clk(gclk));
	jand g1713(.dina(w_n1752_0[0]),.dinb(w_n1740_0[0]),.dout(n1777),.clk(gclk));
	jor g1714(.dina(n1777),.dinb(w_dff_B_3hVnrSk46_1),.dout(n1778),.clk(gclk));
	jand g1715(.dina(w_G494gat_2[2]),.dinb(w_G239gat_3[0]),.dout(n1779),.clk(gclk));
	jand g1716(.dina(w_G477gat_2[1]),.dinb(w_G256gat_3[1]),.dout(n1780),.clk(gclk));
	jor g1717(.dina(w_n1748_0[0]),.dinb(w_n1745_0[0]),.dout(n1781),.clk(gclk));
	jor g1718(.dina(w_n1750_0[0]),.dinb(w_n1744_0[0]),.dout(n1782),.clk(gclk));
	jand g1719(.dina(n1782),.dinb(w_dff_B_ab685Q2h6_1),.dout(n1783),.clk(gclk));
	jxor g1720(.dina(w_n1783_0[1]),.dinb(w_n1780_0[1]),.dout(n1784),.clk(gclk));
	jnot g1721(.din(n1784),.dout(n1785),.clk(gclk));
	jxor g1722(.dina(w_n1785_0[1]),.dinb(w_n1779_0[1]),.dout(n1786),.clk(gclk));
	jxor g1723(.dina(w_n1786_0[1]),.dinb(w_n1778_0[1]),.dout(n1787),.clk(gclk));
	jxor g1724(.dina(w_n1787_0[1]),.dinb(w_n1775_0[1]),.dout(n1788),.clk(gclk));
	jxor g1725(.dina(w_n1788_0[1]),.dinb(w_n1773_0[1]),.dout(n1789),.clk(gclk));
	jxor g1726(.dina(w_n1789_0[1]),.dinb(w_n1770_0[1]),.dout(n1790),.clk(gclk));
	jxor g1727(.dina(w_n1790_0[1]),.dinb(w_n1768_0[1]),.dout(n1791),.clk(gclk));
	jxor g1728(.dina(w_n1791_0[1]),.dinb(w_n1765_0[1]),.dout(w_dff_A_ItMjlGlT1_2),.clk(gclk));
	jnot g1729(.din(w_n1768_0[0]),.dout(n1793),.clk(gclk));
	jnot g1730(.din(w_n1790_0[0]),.dout(n1794),.clk(gclk));
	jor g1731(.dina(n1794),.dinb(w_dff_B_swAYl7xU4_1),.dout(n1795),.clk(gclk));
	jnot g1732(.din(w_n1791_0[0]),.dout(n1796),.clk(gclk));
	jor g1733(.dina(w_dff_B_uo9daJrs0_0),.dinb(w_n1765_0[0]),.dout(n1797),.clk(gclk));
	jand g1734(.dina(n1797),.dinb(w_dff_B_2lTowDer4_1),.dout(n1798),.clk(gclk));
	jand g1735(.dina(w_n1788_0[0]),.dinb(w_n1773_0[0]),.dout(n1799),.clk(gclk));
	jand g1736(.dina(w_n1789_0[0]),.dinb(w_n1770_0[0]),.dout(n1800),.clk(gclk));
	jor g1737(.dina(n1800),.dinb(w_dff_B_CTe4bPiS3_1),.dout(n1801),.clk(gclk));
	jand g1738(.dina(w_G528gat_3[0]),.dinb(w_G222gat_2[1]),.dout(n1802),.clk(gclk));
	jnot g1739(.din(n1802),.dout(n1803),.clk(gclk));
	jand g1740(.dina(w_n1786_0[0]),.dinb(w_n1778_0[0]),.dout(n1804),.clk(gclk));
	jand g1741(.dina(w_n1787_0[0]),.dinb(w_n1775_0[0]),.dout(n1805),.clk(gclk));
	jor g1742(.dina(n1805),.dinb(w_dff_B_DCVTibQ27_1),.dout(n1806),.clk(gclk));
	jand g1743(.dina(w_G511gat_2[2]),.dinb(w_G239gat_2[2]),.dout(n1807),.clk(gclk));
	jand g1744(.dina(w_G494gat_2[1]),.dinb(w_G256gat_3[0]),.dout(n1808),.clk(gclk));
	jor g1745(.dina(w_n1783_0[0]),.dinb(w_n1780_0[0]),.dout(n1809),.clk(gclk));
	jor g1746(.dina(w_n1785_0[0]),.dinb(w_n1779_0[0]),.dout(n1810),.clk(gclk));
	jand g1747(.dina(n1810),.dinb(w_dff_B_HF7UIH5v7_1),.dout(n1811),.clk(gclk));
	jxor g1748(.dina(w_n1811_0[1]),.dinb(w_n1808_0[1]),.dout(n1812),.clk(gclk));
	jnot g1749(.din(n1812),.dout(n1813),.clk(gclk));
	jxor g1750(.dina(w_n1813_0[1]),.dinb(w_n1807_0[1]),.dout(n1814),.clk(gclk));
	jxor g1751(.dina(w_n1814_0[1]),.dinb(w_n1806_0[1]),.dout(n1815),.clk(gclk));
	jxor g1752(.dina(w_n1815_0[1]),.dinb(w_n1803_0[1]),.dout(n1816),.clk(gclk));
	jxor g1753(.dina(w_n1816_0[1]),.dinb(w_n1801_0[1]),.dout(n1817),.clk(gclk));
	jxor g1754(.dina(w_n1817_0[1]),.dinb(w_n1798_0[1]),.dout(w_dff_A_WJUS03tP8_2),.clk(gclk));
	jnot g1755(.din(w_n1801_0[0]),.dout(n1819),.clk(gclk));
	jnot g1756(.din(w_n1816_0[0]),.dout(n1820),.clk(gclk));
	jor g1757(.dina(n1820),.dinb(w_dff_B_NiRQ0XUX0_1),.dout(n1821),.clk(gclk));
	jnot g1758(.din(w_n1817_0[0]),.dout(n1822),.clk(gclk));
	jor g1759(.dina(w_dff_B_k03xV37X7_0),.dinb(w_n1798_0[0]),.dout(n1823),.clk(gclk));
	jand g1760(.dina(n1823),.dinb(w_dff_B_V4tVImYF3_1),.dout(n1824),.clk(gclk));
	jand g1761(.dina(w_n1814_0[0]),.dinb(w_n1806_0[0]),.dout(n1825),.clk(gclk));
	jand g1762(.dina(w_n1815_0[0]),.dinb(w_n1803_0[0]),.dout(n1826),.clk(gclk));
	jor g1763(.dina(n1826),.dinb(w_dff_B_mgjKK9GJ3_1),.dout(n1827),.clk(gclk));
	jand g1764(.dina(w_G528gat_2[2]),.dinb(w_G239gat_2[1]),.dout(n1828),.clk(gclk));
	jand g1765(.dina(w_G511gat_2[1]),.dinb(w_G256gat_2[2]),.dout(n1829),.clk(gclk));
	jor g1766(.dina(w_n1811_0[0]),.dinb(w_n1808_0[0]),.dout(n1830),.clk(gclk));
	jor g1767(.dina(w_n1813_0[0]),.dinb(w_n1807_0[0]),.dout(n1831),.clk(gclk));
	jand g1768(.dina(n1831),.dinb(w_dff_B_AxN3HC4J1_1),.dout(n1832),.clk(gclk));
	jxor g1769(.dina(w_n1832_0[1]),.dinb(w_n1829_0[1]),.dout(n1833),.clk(gclk));
	jnot g1770(.din(n1833),.dout(n1834),.clk(gclk));
	jxor g1771(.dina(w_n1834_0[1]),.dinb(w_n1828_0[1]),.dout(n1835),.clk(gclk));
	jxor g1772(.dina(w_n1835_0[1]),.dinb(w_n1827_0[1]),.dout(n1836),.clk(gclk));
	jxor g1773(.dina(w_n1836_0[1]),.dinb(w_n1824_0[1]),.dout(w_dff_A_8IBM46XT7_2),.clk(gclk));
	jand g1774(.dina(w_G528gat_2[1]),.dinb(w_G256gat_2[1]),.dout(n1838),.clk(gclk));
	jor g1775(.dina(w_n1832_0[0]),.dinb(w_n1829_0[0]),.dout(n1839),.clk(gclk));
	jor g1776(.dina(w_n1834_0[0]),.dinb(w_n1828_0[0]),.dout(n1840),.clk(gclk));
	jand g1777(.dina(n1840),.dinb(w_dff_B_l8E1hQ3o8_1),.dout(n1841),.clk(gclk));
	jor g1778(.dina(w_n1841_0[1]),.dinb(w_n1838_0[1]),.dout(n1842),.clk(gclk));
	jnot g1779(.din(w_n1827_0[0]),.dout(n1843),.clk(gclk));
	jnot g1780(.din(w_n1835_0[0]),.dout(n1844),.clk(gclk));
	jor g1781(.dina(n1844),.dinb(w_dff_B_G1Be0w1L8_1),.dout(n1845),.clk(gclk));
	jnot g1782(.din(w_n1836_0[0]),.dout(n1846),.clk(gclk));
	jor g1783(.dina(w_dff_B_4MdSaJGN5_0),.dinb(w_n1824_0[0]),.dout(n1847),.clk(gclk));
	jand g1784(.dina(n1847),.dinb(w_dff_B_wJhP7oj49_1),.dout(n1848),.clk(gclk));
	jxor g1785(.dina(w_n1841_0[0]),.dinb(w_n1838_0[0]),.dout(n1849),.clk(gclk));
	jnot g1786(.din(w_n1849_0[1]),.dout(n1850),.clk(gclk));
	jor g1787(.dina(w_dff_B_lO57ET7m6_0),.dinb(w_n1848_0[1]),.dout(n1851),.clk(gclk));
	jand g1788(.dina(n1851),.dinb(w_dff_B_tEIzL6Si8_1),.dout(G6287gat),.clk(gclk));
	jxor g1789(.dina(w_n1849_0[0]),.dinb(w_n1848_0[0]),.dout(w_dff_A_Sal8trTP1_2),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_G1gat_0[0]),.doutb(w_G1gat_0[1]),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G1gat_1(.douta(w_G1gat_1[0]),.doutb(w_G1gat_1[1]),.doutc(w_G1gat_1[2]),.din(w_G1gat_0[0]));
	jspl3 jspl3_w_G1gat_2(.douta(w_G1gat_2[0]),.doutb(w_G1gat_2[1]),.doutc(w_G1gat_2[2]),.din(w_G1gat_0[1]));
	jspl3 jspl3_w_G1gat_3(.douta(w_G1gat_3[0]),.doutb(w_G1gat_3[1]),.doutc(w_G1gat_3[2]),.din(w_G1gat_0[2]));
	jspl3 jspl3_w_G1gat_4(.douta(w_G1gat_4[0]),.doutb(w_G1gat_4[1]),.doutc(w_G1gat_4[2]),.din(w_G1gat_1[0]));
	jspl3 jspl3_w_G1gat_5(.douta(w_G1gat_5[0]),.doutb(w_G1gat_5[1]),.doutc(w_G1gat_5[2]),.din(w_G1gat_1[1]));
	jspl3 jspl3_w_G1gat_6(.douta(w_G1gat_6[0]),.doutb(w_G1gat_6[1]),.doutc(w_G1gat_6[2]),.din(w_G1gat_1[2]));
	jspl jspl_w_G1gat_7(.douta(w_G1gat_7[0]),.doutb(w_G1gat_7[1]),.din(w_G1gat_2[0]));
	jspl3 jspl3_w_G18gat_0(.douta(w_G18gat_0[0]),.doutb(w_G18gat_0[1]),.doutc(w_G18gat_0[2]),.din(G18gat));
	jspl3 jspl3_w_G18gat_1(.douta(w_G18gat_1[0]),.doutb(w_G18gat_1[1]),.doutc(w_G18gat_1[2]),.din(w_G18gat_0[0]));
	jspl3 jspl3_w_G18gat_2(.douta(w_G18gat_2[0]),.doutb(w_G18gat_2[1]),.doutc(w_G18gat_2[2]),.din(w_G18gat_0[1]));
	jspl3 jspl3_w_G18gat_3(.douta(w_G18gat_3[0]),.doutb(w_G18gat_3[1]),.doutc(w_G18gat_3[2]),.din(w_G18gat_0[2]));
	jspl3 jspl3_w_G18gat_4(.douta(w_G18gat_4[0]),.doutb(w_G18gat_4[1]),.doutc(w_G18gat_4[2]),.din(w_G18gat_1[0]));
	jspl3 jspl3_w_G18gat_5(.douta(w_G18gat_5[0]),.doutb(w_G18gat_5[1]),.doutc(w_G18gat_5[2]),.din(w_G18gat_1[1]));
	jspl3 jspl3_w_G18gat_6(.douta(w_G18gat_6[0]),.doutb(w_G18gat_6[1]),.doutc(w_G18gat_6[2]),.din(w_G18gat_1[2]));
	jspl3 jspl3_w_G18gat_7(.douta(w_G18gat_7[0]),.doutb(w_G18gat_7[1]),.doutc(w_G18gat_7[2]),.din(w_G18gat_2[0]));
	jspl3 jspl3_w_G35gat_0(.douta(w_G35gat_0[0]),.doutb(w_G35gat_0[1]),.doutc(w_G35gat_0[2]),.din(G35gat));
	jspl3 jspl3_w_G35gat_1(.douta(w_G35gat_1[0]),.doutb(w_G35gat_1[1]),.doutc(w_G35gat_1[2]),.din(w_G35gat_0[0]));
	jspl3 jspl3_w_G35gat_2(.douta(w_G35gat_2[0]),.doutb(w_G35gat_2[1]),.doutc(w_G35gat_2[2]),.din(w_G35gat_0[1]));
	jspl3 jspl3_w_G35gat_3(.douta(w_G35gat_3[0]),.doutb(w_G35gat_3[1]),.doutc(w_G35gat_3[2]),.din(w_G35gat_0[2]));
	jspl3 jspl3_w_G35gat_4(.douta(w_G35gat_4[0]),.doutb(w_G35gat_4[1]),.doutc(w_G35gat_4[2]),.din(w_G35gat_1[0]));
	jspl3 jspl3_w_G35gat_5(.douta(w_G35gat_5[0]),.doutb(w_G35gat_5[1]),.doutc(w_G35gat_5[2]),.din(w_G35gat_1[1]));
	jspl3 jspl3_w_G35gat_6(.douta(w_G35gat_6[0]),.doutb(w_G35gat_6[1]),.doutc(w_G35gat_6[2]),.din(w_G35gat_1[2]));
	jspl3 jspl3_w_G35gat_7(.douta(w_G35gat_7[0]),.doutb(w_G35gat_7[1]),.doutc(w_G35gat_7[2]),.din(w_G35gat_2[0]));
	jspl3 jspl3_w_G52gat_0(.douta(w_G52gat_0[0]),.doutb(w_G52gat_0[1]),.doutc(w_G52gat_0[2]),.din(G52gat));
	jspl3 jspl3_w_G52gat_1(.douta(w_G52gat_1[0]),.doutb(w_G52gat_1[1]),.doutc(w_G52gat_1[2]),.din(w_G52gat_0[0]));
	jspl3 jspl3_w_G52gat_2(.douta(w_G52gat_2[0]),.doutb(w_G52gat_2[1]),.doutc(w_G52gat_2[2]),.din(w_G52gat_0[1]));
	jspl3 jspl3_w_G52gat_3(.douta(w_G52gat_3[0]),.doutb(w_G52gat_3[1]),.doutc(w_G52gat_3[2]),.din(w_G52gat_0[2]));
	jspl3 jspl3_w_G52gat_4(.douta(w_G52gat_4[0]),.doutb(w_G52gat_4[1]),.doutc(w_G52gat_4[2]),.din(w_G52gat_1[0]));
	jspl3 jspl3_w_G52gat_5(.douta(w_G52gat_5[0]),.doutb(w_G52gat_5[1]),.doutc(w_G52gat_5[2]),.din(w_G52gat_1[1]));
	jspl3 jspl3_w_G52gat_6(.douta(w_G52gat_6[0]),.doutb(w_G52gat_6[1]),.doutc(w_G52gat_6[2]),.din(w_G52gat_1[2]));
	jspl3 jspl3_w_G52gat_7(.douta(w_G52gat_7[0]),.doutb(w_G52gat_7[1]),.doutc(w_G52gat_7[2]),.din(w_G52gat_2[0]));
	jspl3 jspl3_w_G69gat_0(.douta(w_G69gat_0[0]),.doutb(w_G69gat_0[1]),.doutc(w_G69gat_0[2]),.din(G69gat));
	jspl3 jspl3_w_G69gat_1(.douta(w_G69gat_1[0]),.doutb(w_G69gat_1[1]),.doutc(w_G69gat_1[2]),.din(w_G69gat_0[0]));
	jspl3 jspl3_w_G69gat_2(.douta(w_G69gat_2[0]),.doutb(w_G69gat_2[1]),.doutc(w_G69gat_2[2]),.din(w_G69gat_0[1]));
	jspl3 jspl3_w_G69gat_3(.douta(w_G69gat_3[0]),.doutb(w_G69gat_3[1]),.doutc(w_G69gat_3[2]),.din(w_G69gat_0[2]));
	jspl3 jspl3_w_G69gat_4(.douta(w_G69gat_4[0]),.doutb(w_G69gat_4[1]),.doutc(w_G69gat_4[2]),.din(w_G69gat_1[0]));
	jspl3 jspl3_w_G69gat_5(.douta(w_G69gat_5[0]),.doutb(w_G69gat_5[1]),.doutc(w_G69gat_5[2]),.din(w_G69gat_1[1]));
	jspl3 jspl3_w_G69gat_6(.douta(w_G69gat_6[0]),.doutb(w_G69gat_6[1]),.doutc(w_G69gat_6[2]),.din(w_G69gat_1[2]));
	jspl jspl_w_G69gat_7(.douta(w_G69gat_7[0]),.doutb(w_G69gat_7[1]),.din(w_G69gat_2[0]));
	jspl3 jspl3_w_G86gat_0(.douta(w_G86gat_0[0]),.doutb(w_G86gat_0[1]),.doutc(w_G86gat_0[2]),.din(G86gat));
	jspl3 jspl3_w_G86gat_1(.douta(w_G86gat_1[0]),.doutb(w_G86gat_1[1]),.doutc(w_G86gat_1[2]),.din(w_G86gat_0[0]));
	jspl3 jspl3_w_G86gat_2(.douta(w_G86gat_2[0]),.doutb(w_G86gat_2[1]),.doutc(w_G86gat_2[2]),.din(w_G86gat_0[1]));
	jspl3 jspl3_w_G86gat_3(.douta(w_G86gat_3[0]),.doutb(w_G86gat_3[1]),.doutc(w_G86gat_3[2]),.din(w_G86gat_0[2]));
	jspl3 jspl3_w_G86gat_4(.douta(w_G86gat_4[0]),.doutb(w_G86gat_4[1]),.doutc(w_G86gat_4[2]),.din(w_G86gat_1[0]));
	jspl3 jspl3_w_G86gat_5(.douta(w_G86gat_5[0]),.doutb(w_G86gat_5[1]),.doutc(w_G86gat_5[2]),.din(w_G86gat_1[1]));
	jspl3 jspl3_w_G86gat_6(.douta(w_G86gat_6[0]),.doutb(w_G86gat_6[1]),.doutc(w_G86gat_6[2]),.din(w_G86gat_1[2]));
	jspl jspl_w_G86gat_7(.douta(w_G86gat_7[0]),.doutb(w_G86gat_7[1]),.din(w_G86gat_2[0]));
	jspl3 jspl3_w_G103gat_0(.douta(w_G103gat_0[0]),.doutb(w_G103gat_0[1]),.doutc(w_G103gat_0[2]),.din(G103gat));
	jspl3 jspl3_w_G103gat_1(.douta(w_G103gat_1[0]),.doutb(w_G103gat_1[1]),.doutc(w_G103gat_1[2]),.din(w_G103gat_0[0]));
	jspl3 jspl3_w_G103gat_2(.douta(w_G103gat_2[0]),.doutb(w_G103gat_2[1]),.doutc(w_G103gat_2[2]),.din(w_G103gat_0[1]));
	jspl3 jspl3_w_G103gat_3(.douta(w_G103gat_3[0]),.doutb(w_G103gat_3[1]),.doutc(w_G103gat_3[2]),.din(w_G103gat_0[2]));
	jspl3 jspl3_w_G103gat_4(.douta(w_G103gat_4[0]),.doutb(w_G103gat_4[1]),.doutc(w_G103gat_4[2]),.din(w_G103gat_1[0]));
	jspl3 jspl3_w_G103gat_5(.douta(w_G103gat_5[0]),.doutb(w_G103gat_5[1]),.doutc(w_G103gat_5[2]),.din(w_G103gat_1[1]));
	jspl3 jspl3_w_G103gat_6(.douta(w_G103gat_6[0]),.doutb(w_G103gat_6[1]),.doutc(w_G103gat_6[2]),.din(w_G103gat_1[2]));
	jspl jspl_w_G103gat_7(.douta(w_G103gat_7[0]),.doutb(w_G103gat_7[1]),.din(w_G103gat_2[0]));
	jspl3 jspl3_w_G120gat_0(.douta(w_G120gat_0[0]),.doutb(w_G120gat_0[1]),.doutc(w_G120gat_0[2]),.din(G120gat));
	jspl3 jspl3_w_G120gat_1(.douta(w_G120gat_1[0]),.doutb(w_G120gat_1[1]),.doutc(w_G120gat_1[2]),.din(w_G120gat_0[0]));
	jspl3 jspl3_w_G120gat_2(.douta(w_G120gat_2[0]),.doutb(w_G120gat_2[1]),.doutc(w_G120gat_2[2]),.din(w_G120gat_0[1]));
	jspl3 jspl3_w_G120gat_3(.douta(w_G120gat_3[0]),.doutb(w_G120gat_3[1]),.doutc(w_G120gat_3[2]),.din(w_G120gat_0[2]));
	jspl3 jspl3_w_G120gat_4(.douta(w_G120gat_4[0]),.doutb(w_G120gat_4[1]),.doutc(w_G120gat_4[2]),.din(w_G120gat_1[0]));
	jspl3 jspl3_w_G120gat_5(.douta(w_G120gat_5[0]),.doutb(w_G120gat_5[1]),.doutc(w_G120gat_5[2]),.din(w_G120gat_1[1]));
	jspl3 jspl3_w_G120gat_6(.douta(w_G120gat_6[0]),.doutb(w_G120gat_6[1]),.doutc(w_G120gat_6[2]),.din(w_G120gat_1[2]));
	jspl jspl_w_G120gat_7(.douta(w_G120gat_7[0]),.doutb(w_G120gat_7[1]),.din(w_G120gat_2[0]));
	jspl3 jspl3_w_G137gat_0(.douta(w_G137gat_0[0]),.doutb(w_G137gat_0[1]),.doutc(w_G137gat_0[2]),.din(G137gat));
	jspl3 jspl3_w_G137gat_1(.douta(w_G137gat_1[0]),.doutb(w_G137gat_1[1]),.doutc(w_G137gat_1[2]),.din(w_G137gat_0[0]));
	jspl3 jspl3_w_G137gat_2(.douta(w_G137gat_2[0]),.doutb(w_G137gat_2[1]),.doutc(w_G137gat_2[2]),.din(w_G137gat_0[1]));
	jspl3 jspl3_w_G137gat_3(.douta(w_G137gat_3[0]),.doutb(w_G137gat_3[1]),.doutc(w_G137gat_3[2]),.din(w_G137gat_0[2]));
	jspl3 jspl3_w_G137gat_4(.douta(w_G137gat_4[0]),.doutb(w_G137gat_4[1]),.doutc(w_G137gat_4[2]),.din(w_G137gat_1[0]));
	jspl3 jspl3_w_G137gat_5(.douta(w_G137gat_5[0]),.doutb(w_G137gat_5[1]),.doutc(w_G137gat_5[2]),.din(w_G137gat_1[1]));
	jspl3 jspl3_w_G137gat_6(.douta(w_G137gat_6[0]),.doutb(w_G137gat_6[1]),.doutc(w_G137gat_6[2]),.din(w_G137gat_1[2]));
	jspl jspl_w_G137gat_7(.douta(w_G137gat_7[0]),.doutb(w_G137gat_7[1]),.din(w_G137gat_2[0]));
	jspl3 jspl3_w_G154gat_0(.douta(w_G154gat_0[0]),.doutb(w_G154gat_0[1]),.doutc(w_G154gat_0[2]),.din(G154gat));
	jspl3 jspl3_w_G154gat_1(.douta(w_G154gat_1[0]),.doutb(w_G154gat_1[1]),.doutc(w_G154gat_1[2]),.din(w_G154gat_0[0]));
	jspl3 jspl3_w_G154gat_2(.douta(w_G154gat_2[0]),.doutb(w_G154gat_2[1]),.doutc(w_G154gat_2[2]),.din(w_G154gat_0[1]));
	jspl3 jspl3_w_G154gat_3(.douta(w_G154gat_3[0]),.doutb(w_G154gat_3[1]),.doutc(w_G154gat_3[2]),.din(w_G154gat_0[2]));
	jspl3 jspl3_w_G154gat_4(.douta(w_G154gat_4[0]),.doutb(w_G154gat_4[1]),.doutc(w_G154gat_4[2]),.din(w_G154gat_1[0]));
	jspl3 jspl3_w_G154gat_5(.douta(w_G154gat_5[0]),.doutb(w_G154gat_5[1]),.doutc(w_G154gat_5[2]),.din(w_G154gat_1[1]));
	jspl3 jspl3_w_G154gat_6(.douta(w_G154gat_6[0]),.doutb(w_G154gat_6[1]),.doutc(w_G154gat_6[2]),.din(w_G154gat_1[2]));
	jspl jspl_w_G154gat_7(.douta(w_G154gat_7[0]),.doutb(w_G154gat_7[1]),.din(w_G154gat_2[0]));
	jspl3 jspl3_w_G171gat_0(.douta(w_G171gat_0[0]),.doutb(w_G171gat_0[1]),.doutc(w_G171gat_0[2]),.din(G171gat));
	jspl3 jspl3_w_G171gat_1(.douta(w_G171gat_1[0]),.doutb(w_G171gat_1[1]),.doutc(w_G171gat_1[2]),.din(w_G171gat_0[0]));
	jspl3 jspl3_w_G171gat_2(.douta(w_G171gat_2[0]),.doutb(w_G171gat_2[1]),.doutc(w_G171gat_2[2]),.din(w_G171gat_0[1]));
	jspl3 jspl3_w_G171gat_3(.douta(w_G171gat_3[0]),.doutb(w_G171gat_3[1]),.doutc(w_G171gat_3[2]),.din(w_G171gat_0[2]));
	jspl3 jspl3_w_G171gat_4(.douta(w_G171gat_4[0]),.doutb(w_G171gat_4[1]),.doutc(w_G171gat_4[2]),.din(w_G171gat_1[0]));
	jspl3 jspl3_w_G171gat_5(.douta(w_G171gat_5[0]),.doutb(w_G171gat_5[1]),.doutc(w_G171gat_5[2]),.din(w_G171gat_1[1]));
	jspl3 jspl3_w_G171gat_6(.douta(w_G171gat_6[0]),.doutb(w_G171gat_6[1]),.doutc(w_G171gat_6[2]),.din(w_G171gat_1[2]));
	jspl jspl_w_G171gat_7(.douta(w_G171gat_7[0]),.doutb(w_G171gat_7[1]),.din(w_G171gat_2[0]));
	jspl3 jspl3_w_G188gat_0(.douta(w_G188gat_0[0]),.doutb(w_G188gat_0[1]),.doutc(w_G188gat_0[2]),.din(G188gat));
	jspl3 jspl3_w_G188gat_1(.douta(w_G188gat_1[0]),.doutb(w_G188gat_1[1]),.doutc(w_G188gat_1[2]),.din(w_G188gat_0[0]));
	jspl3 jspl3_w_G188gat_2(.douta(w_G188gat_2[0]),.doutb(w_G188gat_2[1]),.doutc(w_G188gat_2[2]),.din(w_G188gat_0[1]));
	jspl3 jspl3_w_G188gat_3(.douta(w_G188gat_3[0]),.doutb(w_G188gat_3[1]),.doutc(w_G188gat_3[2]),.din(w_G188gat_0[2]));
	jspl3 jspl3_w_G188gat_4(.douta(w_G188gat_4[0]),.doutb(w_G188gat_4[1]),.doutc(w_G188gat_4[2]),.din(w_G188gat_1[0]));
	jspl3 jspl3_w_G188gat_5(.douta(w_G188gat_5[0]),.doutb(w_G188gat_5[1]),.doutc(w_G188gat_5[2]),.din(w_G188gat_1[1]));
	jspl3 jspl3_w_G188gat_6(.douta(w_G188gat_6[0]),.doutb(w_G188gat_6[1]),.doutc(w_G188gat_6[2]),.din(w_G188gat_1[2]));
	jspl jspl_w_G188gat_7(.douta(w_G188gat_7[0]),.doutb(w_G188gat_7[1]),.din(w_G188gat_2[0]));
	jspl3 jspl3_w_G205gat_0(.douta(w_G205gat_0[0]),.doutb(w_G205gat_0[1]),.doutc(w_G205gat_0[2]),.din(G205gat));
	jspl3 jspl3_w_G205gat_1(.douta(w_G205gat_1[0]),.doutb(w_G205gat_1[1]),.doutc(w_G205gat_1[2]),.din(w_G205gat_0[0]));
	jspl3 jspl3_w_G205gat_2(.douta(w_G205gat_2[0]),.doutb(w_G205gat_2[1]),.doutc(w_G205gat_2[2]),.din(w_G205gat_0[1]));
	jspl3 jspl3_w_G205gat_3(.douta(w_G205gat_3[0]),.doutb(w_G205gat_3[1]),.doutc(w_G205gat_3[2]),.din(w_G205gat_0[2]));
	jspl3 jspl3_w_G205gat_4(.douta(w_G205gat_4[0]),.doutb(w_G205gat_4[1]),.doutc(w_G205gat_4[2]),.din(w_G205gat_1[0]));
	jspl3 jspl3_w_G205gat_5(.douta(w_G205gat_5[0]),.doutb(w_G205gat_5[1]),.doutc(w_G205gat_5[2]),.din(w_G205gat_1[1]));
	jspl3 jspl3_w_G205gat_6(.douta(w_G205gat_6[0]),.doutb(w_G205gat_6[1]),.doutc(w_G205gat_6[2]),.din(w_G205gat_1[2]));
	jspl jspl_w_G205gat_7(.douta(w_G205gat_7[0]),.doutb(w_G205gat_7[1]),.din(w_G205gat_2[0]));
	jspl3 jspl3_w_G222gat_0(.douta(w_G222gat_0[0]),.doutb(w_G222gat_0[1]),.doutc(w_G222gat_0[2]),.din(G222gat));
	jspl3 jspl3_w_G222gat_1(.douta(w_G222gat_1[0]),.doutb(w_G222gat_1[1]),.doutc(w_G222gat_1[2]),.din(w_G222gat_0[0]));
	jspl3 jspl3_w_G222gat_2(.douta(w_G222gat_2[0]),.doutb(w_G222gat_2[1]),.doutc(w_G222gat_2[2]),.din(w_G222gat_0[1]));
	jspl3 jspl3_w_G222gat_3(.douta(w_G222gat_3[0]),.doutb(w_G222gat_3[1]),.doutc(w_G222gat_3[2]),.din(w_G222gat_0[2]));
	jspl3 jspl3_w_G222gat_4(.douta(w_G222gat_4[0]),.doutb(w_G222gat_4[1]),.doutc(w_G222gat_4[2]),.din(w_G222gat_1[0]));
	jspl3 jspl3_w_G222gat_5(.douta(w_G222gat_5[0]),.doutb(w_G222gat_5[1]),.doutc(w_G222gat_5[2]),.din(w_G222gat_1[1]));
	jspl3 jspl3_w_G222gat_6(.douta(w_G222gat_6[0]),.doutb(w_G222gat_6[1]),.doutc(w_G222gat_6[2]),.din(w_G222gat_1[2]));
	jspl jspl_w_G222gat_7(.douta(w_G222gat_7[0]),.doutb(w_G222gat_7[1]),.din(w_G222gat_2[0]));
	jspl3 jspl3_w_G239gat_0(.douta(w_G239gat_0[0]),.doutb(w_G239gat_0[1]),.doutc(w_G239gat_0[2]),.din(G239gat));
	jspl3 jspl3_w_G239gat_1(.douta(w_G239gat_1[0]),.doutb(w_G239gat_1[1]),.doutc(w_G239gat_1[2]),.din(w_G239gat_0[0]));
	jspl3 jspl3_w_G239gat_2(.douta(w_G239gat_2[0]),.doutb(w_G239gat_2[1]),.doutc(w_G239gat_2[2]),.din(w_G239gat_0[1]));
	jspl3 jspl3_w_G239gat_3(.douta(w_G239gat_3[0]),.doutb(w_G239gat_3[1]),.doutc(w_G239gat_3[2]),.din(w_G239gat_0[2]));
	jspl3 jspl3_w_G239gat_4(.douta(w_G239gat_4[0]),.doutb(w_G239gat_4[1]),.doutc(w_G239gat_4[2]),.din(w_G239gat_1[0]));
	jspl3 jspl3_w_G239gat_5(.douta(w_G239gat_5[0]),.doutb(w_G239gat_5[1]),.doutc(w_G239gat_5[2]),.din(w_G239gat_1[1]));
	jspl3 jspl3_w_G239gat_6(.douta(w_G239gat_6[0]),.doutb(w_G239gat_6[1]),.doutc(w_G239gat_6[2]),.din(w_G239gat_1[2]));
	jspl jspl_w_G239gat_7(.douta(w_G239gat_7[0]),.doutb(w_G239gat_7[1]),.din(w_G239gat_2[0]));
	jspl3 jspl3_w_G256gat_0(.douta(w_G256gat_0[0]),.doutb(w_G256gat_0[1]),.doutc(w_G256gat_0[2]),.din(G256gat));
	jspl3 jspl3_w_G256gat_1(.douta(w_G256gat_1[0]),.doutb(w_G256gat_1[1]),.doutc(w_G256gat_1[2]),.din(w_G256gat_0[0]));
	jspl3 jspl3_w_G256gat_2(.douta(w_G256gat_2[0]),.doutb(w_G256gat_2[1]),.doutc(w_G256gat_2[2]),.din(w_G256gat_0[1]));
	jspl3 jspl3_w_G256gat_3(.douta(w_G256gat_3[0]),.doutb(w_G256gat_3[1]),.doutc(w_G256gat_3[2]),.din(w_G256gat_0[2]));
	jspl3 jspl3_w_G256gat_4(.douta(w_G256gat_4[0]),.doutb(w_G256gat_4[1]),.doutc(w_G256gat_4[2]),.din(w_G256gat_1[0]));
	jspl3 jspl3_w_G256gat_5(.douta(w_G256gat_5[0]),.doutb(w_G256gat_5[1]),.doutc(w_G256gat_5[2]),.din(w_G256gat_1[1]));
	jspl3 jspl3_w_G256gat_6(.douta(w_G256gat_6[0]),.doutb(w_G256gat_6[1]),.doutc(w_G256gat_6[2]),.din(w_G256gat_1[2]));
	jspl jspl_w_G256gat_7(.douta(w_G256gat_7[0]),.doutb(w_G256gat_7[1]),.din(w_G256gat_2[0]));
	jspl3 jspl3_w_G273gat_0(.douta(w_G273gat_0[0]),.doutb(w_G273gat_0[1]),.doutc(w_G273gat_0[2]),.din(G273gat));
	jspl3 jspl3_w_G273gat_1(.douta(w_G273gat_1[0]),.doutb(w_G273gat_1[1]),.doutc(w_G273gat_1[2]),.din(w_G273gat_0[0]));
	jspl3 jspl3_w_G273gat_2(.douta(w_G273gat_2[0]),.doutb(w_G273gat_2[1]),.doutc(w_G273gat_2[2]),.din(w_G273gat_0[1]));
	jspl3 jspl3_w_G273gat_3(.douta(w_G273gat_3[0]),.doutb(w_G273gat_3[1]),.doutc(w_G273gat_3[2]),.din(w_G273gat_0[2]));
	jspl3 jspl3_w_G273gat_4(.douta(w_G273gat_4[0]),.doutb(w_G273gat_4[1]),.doutc(w_G273gat_4[2]),.din(w_G273gat_1[0]));
	jspl3 jspl3_w_G273gat_5(.douta(w_G273gat_5[0]),.doutb(w_G273gat_5[1]),.doutc(w_G273gat_5[2]),.din(w_G273gat_1[1]));
	jspl3 jspl3_w_G273gat_6(.douta(w_G273gat_6[0]),.doutb(w_G273gat_6[1]),.doutc(w_G273gat_6[2]),.din(w_G273gat_1[2]));
	jspl3 jspl3_w_G273gat_7(.douta(w_G273gat_7[0]),.doutb(w_G273gat_7[1]),.doutc(w_G273gat_7[2]),.din(w_G273gat_2[0]));
	jspl3 jspl3_w_G290gat_0(.douta(w_G290gat_0[0]),.doutb(w_G290gat_0[1]),.doutc(w_G290gat_0[2]),.din(G290gat));
	jspl3 jspl3_w_G290gat_1(.douta(w_G290gat_1[0]),.doutb(w_G290gat_1[1]),.doutc(w_G290gat_1[2]),.din(w_G290gat_0[0]));
	jspl3 jspl3_w_G290gat_2(.douta(w_G290gat_2[0]),.doutb(w_G290gat_2[1]),.doutc(w_G290gat_2[2]),.din(w_G290gat_0[1]));
	jspl3 jspl3_w_G290gat_3(.douta(w_G290gat_3[0]),.doutb(w_G290gat_3[1]),.doutc(w_G290gat_3[2]),.din(w_G290gat_0[2]));
	jspl3 jspl3_w_G290gat_4(.douta(w_G290gat_4[0]),.doutb(w_G290gat_4[1]),.doutc(w_G290gat_4[2]),.din(w_G290gat_1[0]));
	jspl3 jspl3_w_G290gat_5(.douta(w_G290gat_5[0]),.doutb(w_G290gat_5[1]),.doutc(w_G290gat_5[2]),.din(w_G290gat_1[1]));
	jspl3 jspl3_w_G290gat_6(.douta(w_G290gat_6[0]),.doutb(w_G290gat_6[1]),.doutc(w_G290gat_6[2]),.din(w_G290gat_1[2]));
	jspl3 jspl3_w_G290gat_7(.douta(w_G290gat_7[0]),.doutb(w_G290gat_7[1]),.doutc(w_G290gat_7[2]),.din(w_G290gat_2[0]));
	jspl3 jspl3_w_G307gat_0(.douta(w_G307gat_0[0]),.doutb(w_G307gat_0[1]),.doutc(w_G307gat_0[2]),.din(G307gat));
	jspl3 jspl3_w_G307gat_1(.douta(w_G307gat_1[0]),.doutb(w_G307gat_1[1]),.doutc(w_G307gat_1[2]),.din(w_G307gat_0[0]));
	jspl3 jspl3_w_G307gat_2(.douta(w_G307gat_2[0]),.doutb(w_dff_A_TGokZRHD9_1),.doutc(w_G307gat_2[2]),.din(w_G307gat_0[1]));
	jspl3 jspl3_w_G307gat_3(.douta(w_G307gat_3[0]),.doutb(w_G307gat_3[1]),.doutc(w_G307gat_3[2]),.din(w_G307gat_0[2]));
	jspl3 jspl3_w_G307gat_4(.douta(w_G307gat_4[0]),.doutb(w_G307gat_4[1]),.doutc(w_G307gat_4[2]),.din(w_G307gat_1[0]));
	jspl3 jspl3_w_G307gat_5(.douta(w_G307gat_5[0]),.doutb(w_G307gat_5[1]),.doutc(w_G307gat_5[2]),.din(w_G307gat_1[1]));
	jspl3 jspl3_w_G307gat_6(.douta(w_G307gat_6[0]),.doutb(w_G307gat_6[1]),.doutc(w_G307gat_6[2]),.din(w_G307gat_1[2]));
	jspl3 jspl3_w_G307gat_7(.douta(w_G307gat_7[0]),.doutb(w_G307gat_7[1]),.doutc(w_G307gat_7[2]),.din(w_G307gat_2[0]));
	jspl3 jspl3_w_G324gat_0(.douta(w_G324gat_0[0]),.doutb(w_G324gat_0[1]),.doutc(w_G324gat_0[2]),.din(G324gat));
	jspl3 jspl3_w_G324gat_1(.douta(w_G324gat_1[0]),.doutb(w_G324gat_1[1]),.doutc(w_G324gat_1[2]),.din(w_G324gat_0[0]));
	jspl3 jspl3_w_G324gat_2(.douta(w_G324gat_2[0]),.doutb(w_G324gat_2[1]),.doutc(w_G324gat_2[2]),.din(w_G324gat_0[1]));
	jspl3 jspl3_w_G324gat_3(.douta(w_G324gat_3[0]),.doutb(w_G324gat_3[1]),.doutc(w_G324gat_3[2]),.din(w_G324gat_0[2]));
	jspl3 jspl3_w_G324gat_4(.douta(w_G324gat_4[0]),.doutb(w_G324gat_4[1]),.doutc(w_G324gat_4[2]),.din(w_G324gat_1[0]));
	jspl3 jspl3_w_G324gat_5(.douta(w_G324gat_5[0]),.doutb(w_G324gat_5[1]),.doutc(w_G324gat_5[2]),.din(w_G324gat_1[1]));
	jspl3 jspl3_w_G324gat_6(.douta(w_G324gat_6[0]),.doutb(w_G324gat_6[1]),.doutc(w_G324gat_6[2]),.din(w_G324gat_1[2]));
	jspl jspl_w_G324gat_7(.douta(w_G324gat_7[0]),.doutb(w_G324gat_7[1]),.din(w_G324gat_2[0]));
	jspl3 jspl3_w_G341gat_0(.douta(w_G341gat_0[0]),.doutb(w_G341gat_0[1]),.doutc(w_G341gat_0[2]),.din(G341gat));
	jspl3 jspl3_w_G341gat_1(.douta(w_G341gat_1[0]),.doutb(w_G341gat_1[1]),.doutc(w_G341gat_1[2]),.din(w_G341gat_0[0]));
	jspl3 jspl3_w_G341gat_2(.douta(w_G341gat_2[0]),.doutb(w_G341gat_2[1]),.doutc(w_G341gat_2[2]),.din(w_G341gat_0[1]));
	jspl3 jspl3_w_G341gat_3(.douta(w_G341gat_3[0]),.doutb(w_G341gat_3[1]),.doutc(w_G341gat_3[2]),.din(w_G341gat_0[2]));
	jspl3 jspl3_w_G341gat_4(.douta(w_G341gat_4[0]),.doutb(w_G341gat_4[1]),.doutc(w_G341gat_4[2]),.din(w_G341gat_1[0]));
	jspl3 jspl3_w_G341gat_5(.douta(w_G341gat_5[0]),.doutb(w_G341gat_5[1]),.doutc(w_G341gat_5[2]),.din(w_G341gat_1[1]));
	jspl3 jspl3_w_G341gat_6(.douta(w_G341gat_6[0]),.doutb(w_G341gat_6[1]),.doutc(w_G341gat_6[2]),.din(w_G341gat_1[2]));
	jspl jspl_w_G341gat_7(.douta(w_G341gat_7[0]),.doutb(w_G341gat_7[1]),.din(w_G341gat_2[0]));
	jspl3 jspl3_w_G358gat_0(.douta(w_G358gat_0[0]),.doutb(w_G358gat_0[1]),.doutc(w_G358gat_0[2]),.din(G358gat));
	jspl3 jspl3_w_G358gat_1(.douta(w_G358gat_1[0]),.doutb(w_G358gat_1[1]),.doutc(w_G358gat_1[2]),.din(w_G358gat_0[0]));
	jspl3 jspl3_w_G358gat_2(.douta(w_G358gat_2[0]),.doutb(w_G358gat_2[1]),.doutc(w_G358gat_2[2]),.din(w_G358gat_0[1]));
	jspl3 jspl3_w_G358gat_3(.douta(w_G358gat_3[0]),.doutb(w_G358gat_3[1]),.doutc(w_G358gat_3[2]),.din(w_G358gat_0[2]));
	jspl3 jspl3_w_G358gat_4(.douta(w_G358gat_4[0]),.doutb(w_G358gat_4[1]),.doutc(w_G358gat_4[2]),.din(w_G358gat_1[0]));
	jspl3 jspl3_w_G358gat_5(.douta(w_G358gat_5[0]),.doutb(w_G358gat_5[1]),.doutc(w_G358gat_5[2]),.din(w_G358gat_1[1]));
	jspl3 jspl3_w_G358gat_6(.douta(w_G358gat_6[0]),.doutb(w_G358gat_6[1]),.doutc(w_G358gat_6[2]),.din(w_G358gat_1[2]));
	jspl jspl_w_G358gat_7(.douta(w_G358gat_7[0]),.doutb(w_G358gat_7[1]),.din(w_G358gat_2[0]));
	jspl3 jspl3_w_G375gat_0(.douta(w_G375gat_0[0]),.doutb(w_G375gat_0[1]),.doutc(w_G375gat_0[2]),.din(G375gat));
	jspl3 jspl3_w_G375gat_1(.douta(w_G375gat_1[0]),.doutb(w_G375gat_1[1]),.doutc(w_G375gat_1[2]),.din(w_G375gat_0[0]));
	jspl3 jspl3_w_G375gat_2(.douta(w_G375gat_2[0]),.doutb(w_G375gat_2[1]),.doutc(w_G375gat_2[2]),.din(w_G375gat_0[1]));
	jspl3 jspl3_w_G375gat_3(.douta(w_G375gat_3[0]),.doutb(w_G375gat_3[1]),.doutc(w_G375gat_3[2]),.din(w_G375gat_0[2]));
	jspl3 jspl3_w_G375gat_4(.douta(w_G375gat_4[0]),.doutb(w_G375gat_4[1]),.doutc(w_G375gat_4[2]),.din(w_G375gat_1[0]));
	jspl3 jspl3_w_G375gat_5(.douta(w_G375gat_5[0]),.doutb(w_G375gat_5[1]),.doutc(w_G375gat_5[2]),.din(w_G375gat_1[1]));
	jspl3 jspl3_w_G375gat_6(.douta(w_G375gat_6[0]),.doutb(w_G375gat_6[1]),.doutc(w_G375gat_6[2]),.din(w_G375gat_1[2]));
	jspl jspl_w_G375gat_7(.douta(w_G375gat_7[0]),.doutb(w_G375gat_7[1]),.din(w_G375gat_2[0]));
	jspl3 jspl3_w_G392gat_0(.douta(w_G392gat_0[0]),.doutb(w_G392gat_0[1]),.doutc(w_G392gat_0[2]),.din(G392gat));
	jspl3 jspl3_w_G392gat_1(.douta(w_G392gat_1[0]),.doutb(w_G392gat_1[1]),.doutc(w_G392gat_1[2]),.din(w_G392gat_0[0]));
	jspl3 jspl3_w_G392gat_2(.douta(w_G392gat_2[0]),.doutb(w_G392gat_2[1]),.doutc(w_G392gat_2[2]),.din(w_G392gat_0[1]));
	jspl3 jspl3_w_G392gat_3(.douta(w_G392gat_3[0]),.doutb(w_G392gat_3[1]),.doutc(w_G392gat_3[2]),.din(w_G392gat_0[2]));
	jspl3 jspl3_w_G392gat_4(.douta(w_G392gat_4[0]),.doutb(w_G392gat_4[1]),.doutc(w_G392gat_4[2]),.din(w_G392gat_1[0]));
	jspl3 jspl3_w_G392gat_5(.douta(w_G392gat_5[0]),.doutb(w_G392gat_5[1]),.doutc(w_G392gat_5[2]),.din(w_G392gat_1[1]));
	jspl3 jspl3_w_G392gat_6(.douta(w_G392gat_6[0]),.doutb(w_G392gat_6[1]),.doutc(w_G392gat_6[2]),.din(w_G392gat_1[2]));
	jspl jspl_w_G392gat_7(.douta(w_G392gat_7[0]),.doutb(w_G392gat_7[1]),.din(w_G392gat_2[0]));
	jspl3 jspl3_w_G409gat_0(.douta(w_G409gat_0[0]),.doutb(w_G409gat_0[1]),.doutc(w_G409gat_0[2]),.din(G409gat));
	jspl3 jspl3_w_G409gat_1(.douta(w_G409gat_1[0]),.doutb(w_G409gat_1[1]),.doutc(w_G409gat_1[2]),.din(w_G409gat_0[0]));
	jspl3 jspl3_w_G409gat_2(.douta(w_G409gat_2[0]),.doutb(w_G409gat_2[1]),.doutc(w_G409gat_2[2]),.din(w_G409gat_0[1]));
	jspl3 jspl3_w_G409gat_3(.douta(w_G409gat_3[0]),.doutb(w_G409gat_3[1]),.doutc(w_G409gat_3[2]),.din(w_G409gat_0[2]));
	jspl3 jspl3_w_G409gat_4(.douta(w_G409gat_4[0]),.doutb(w_G409gat_4[1]),.doutc(w_G409gat_4[2]),.din(w_G409gat_1[0]));
	jspl3 jspl3_w_G409gat_5(.douta(w_G409gat_5[0]),.doutb(w_G409gat_5[1]),.doutc(w_G409gat_5[2]),.din(w_G409gat_1[1]));
	jspl3 jspl3_w_G409gat_6(.douta(w_G409gat_6[0]),.doutb(w_G409gat_6[1]),.doutc(w_G409gat_6[2]),.din(w_G409gat_1[2]));
	jspl jspl_w_G409gat_7(.douta(w_G409gat_7[0]),.doutb(w_G409gat_7[1]),.din(w_G409gat_2[0]));
	jspl3 jspl3_w_G426gat_0(.douta(w_G426gat_0[0]),.doutb(w_G426gat_0[1]),.doutc(w_G426gat_0[2]),.din(G426gat));
	jspl3 jspl3_w_G426gat_1(.douta(w_G426gat_1[0]),.doutb(w_G426gat_1[1]),.doutc(w_G426gat_1[2]),.din(w_G426gat_0[0]));
	jspl3 jspl3_w_G426gat_2(.douta(w_G426gat_2[0]),.doutb(w_G426gat_2[1]),.doutc(w_G426gat_2[2]),.din(w_G426gat_0[1]));
	jspl3 jspl3_w_G426gat_3(.douta(w_G426gat_3[0]),.doutb(w_G426gat_3[1]),.doutc(w_G426gat_3[2]),.din(w_G426gat_0[2]));
	jspl3 jspl3_w_G426gat_4(.douta(w_G426gat_4[0]),.doutb(w_G426gat_4[1]),.doutc(w_G426gat_4[2]),.din(w_G426gat_1[0]));
	jspl3 jspl3_w_G426gat_5(.douta(w_G426gat_5[0]),.doutb(w_G426gat_5[1]),.doutc(w_G426gat_5[2]),.din(w_G426gat_1[1]));
	jspl3 jspl3_w_G426gat_6(.douta(w_G426gat_6[0]),.doutb(w_G426gat_6[1]),.doutc(w_G426gat_6[2]),.din(w_G426gat_1[2]));
	jspl jspl_w_G426gat_7(.douta(w_G426gat_7[0]),.doutb(w_G426gat_7[1]),.din(w_G426gat_2[0]));
	jspl3 jspl3_w_G443gat_0(.douta(w_G443gat_0[0]),.doutb(w_G443gat_0[1]),.doutc(w_G443gat_0[2]),.din(G443gat));
	jspl3 jspl3_w_G443gat_1(.douta(w_G443gat_1[0]),.doutb(w_G443gat_1[1]),.doutc(w_G443gat_1[2]),.din(w_G443gat_0[0]));
	jspl3 jspl3_w_G443gat_2(.douta(w_G443gat_2[0]),.doutb(w_G443gat_2[1]),.doutc(w_G443gat_2[2]),.din(w_G443gat_0[1]));
	jspl3 jspl3_w_G443gat_3(.douta(w_G443gat_3[0]),.doutb(w_G443gat_3[1]),.doutc(w_G443gat_3[2]),.din(w_G443gat_0[2]));
	jspl3 jspl3_w_G443gat_4(.douta(w_G443gat_4[0]),.doutb(w_G443gat_4[1]),.doutc(w_G443gat_4[2]),.din(w_G443gat_1[0]));
	jspl3 jspl3_w_G443gat_5(.douta(w_G443gat_5[0]),.doutb(w_G443gat_5[1]),.doutc(w_G443gat_5[2]),.din(w_G443gat_1[1]));
	jspl3 jspl3_w_G443gat_6(.douta(w_G443gat_6[0]),.doutb(w_G443gat_6[1]),.doutc(w_G443gat_6[2]),.din(w_G443gat_1[2]));
	jspl jspl_w_G443gat_7(.douta(w_G443gat_7[0]),.doutb(w_G443gat_7[1]),.din(w_G443gat_2[0]));
	jspl3 jspl3_w_G460gat_0(.douta(w_G460gat_0[0]),.doutb(w_G460gat_0[1]),.doutc(w_G460gat_0[2]),.din(G460gat));
	jspl3 jspl3_w_G460gat_1(.douta(w_G460gat_1[0]),.doutb(w_G460gat_1[1]),.doutc(w_G460gat_1[2]),.din(w_G460gat_0[0]));
	jspl3 jspl3_w_G460gat_2(.douta(w_G460gat_2[0]),.doutb(w_G460gat_2[1]),.doutc(w_G460gat_2[2]),.din(w_G460gat_0[1]));
	jspl3 jspl3_w_G460gat_3(.douta(w_G460gat_3[0]),.doutb(w_G460gat_3[1]),.doutc(w_G460gat_3[2]),.din(w_G460gat_0[2]));
	jspl3 jspl3_w_G460gat_4(.douta(w_G460gat_4[0]),.doutb(w_G460gat_4[1]),.doutc(w_G460gat_4[2]),.din(w_G460gat_1[0]));
	jspl3 jspl3_w_G460gat_5(.douta(w_G460gat_5[0]),.doutb(w_G460gat_5[1]),.doutc(w_G460gat_5[2]),.din(w_G460gat_1[1]));
	jspl3 jspl3_w_G460gat_6(.douta(w_G460gat_6[0]),.doutb(w_G460gat_6[1]),.doutc(w_G460gat_6[2]),.din(w_G460gat_1[2]));
	jspl jspl_w_G460gat_7(.douta(w_G460gat_7[0]),.doutb(w_G460gat_7[1]),.din(w_G460gat_2[0]));
	jspl3 jspl3_w_G477gat_0(.douta(w_G477gat_0[0]),.doutb(w_G477gat_0[1]),.doutc(w_G477gat_0[2]),.din(G477gat));
	jspl3 jspl3_w_G477gat_1(.douta(w_G477gat_1[0]),.doutb(w_G477gat_1[1]),.doutc(w_G477gat_1[2]),.din(w_G477gat_0[0]));
	jspl3 jspl3_w_G477gat_2(.douta(w_G477gat_2[0]),.doutb(w_G477gat_2[1]),.doutc(w_G477gat_2[2]),.din(w_G477gat_0[1]));
	jspl3 jspl3_w_G477gat_3(.douta(w_G477gat_3[0]),.doutb(w_G477gat_3[1]),.doutc(w_G477gat_3[2]),.din(w_G477gat_0[2]));
	jspl3 jspl3_w_G477gat_4(.douta(w_G477gat_4[0]),.doutb(w_G477gat_4[1]),.doutc(w_G477gat_4[2]),.din(w_G477gat_1[0]));
	jspl3 jspl3_w_G477gat_5(.douta(w_G477gat_5[0]),.doutb(w_G477gat_5[1]),.doutc(w_G477gat_5[2]),.din(w_G477gat_1[1]));
	jspl3 jspl3_w_G477gat_6(.douta(w_G477gat_6[0]),.doutb(w_G477gat_6[1]),.doutc(w_G477gat_6[2]),.din(w_G477gat_1[2]));
	jspl jspl_w_G477gat_7(.douta(w_G477gat_7[0]),.doutb(w_G477gat_7[1]),.din(w_G477gat_2[0]));
	jspl3 jspl3_w_G494gat_0(.douta(w_G494gat_0[0]),.doutb(w_G494gat_0[1]),.doutc(w_G494gat_0[2]),.din(G494gat));
	jspl3 jspl3_w_G494gat_1(.douta(w_G494gat_1[0]),.doutb(w_G494gat_1[1]),.doutc(w_G494gat_1[2]),.din(w_G494gat_0[0]));
	jspl3 jspl3_w_G494gat_2(.douta(w_G494gat_2[0]),.doutb(w_G494gat_2[1]),.doutc(w_G494gat_2[2]),.din(w_G494gat_0[1]));
	jspl3 jspl3_w_G494gat_3(.douta(w_G494gat_3[0]),.doutb(w_G494gat_3[1]),.doutc(w_G494gat_3[2]),.din(w_G494gat_0[2]));
	jspl3 jspl3_w_G494gat_4(.douta(w_G494gat_4[0]),.doutb(w_G494gat_4[1]),.doutc(w_G494gat_4[2]),.din(w_G494gat_1[0]));
	jspl3 jspl3_w_G494gat_5(.douta(w_G494gat_5[0]),.doutb(w_G494gat_5[1]),.doutc(w_G494gat_5[2]),.din(w_G494gat_1[1]));
	jspl3 jspl3_w_G494gat_6(.douta(w_G494gat_6[0]),.doutb(w_G494gat_6[1]),.doutc(w_G494gat_6[2]),.din(w_G494gat_1[2]));
	jspl jspl_w_G494gat_7(.douta(w_G494gat_7[0]),.doutb(w_G494gat_7[1]),.din(w_G494gat_2[0]));
	jspl3 jspl3_w_G511gat_0(.douta(w_G511gat_0[0]),.doutb(w_G511gat_0[1]),.doutc(w_G511gat_0[2]),.din(G511gat));
	jspl3 jspl3_w_G511gat_1(.douta(w_G511gat_1[0]),.doutb(w_G511gat_1[1]),.doutc(w_G511gat_1[2]),.din(w_G511gat_0[0]));
	jspl3 jspl3_w_G511gat_2(.douta(w_G511gat_2[0]),.doutb(w_G511gat_2[1]),.doutc(w_G511gat_2[2]),.din(w_G511gat_0[1]));
	jspl3 jspl3_w_G511gat_3(.douta(w_G511gat_3[0]),.doutb(w_G511gat_3[1]),.doutc(w_G511gat_3[2]),.din(w_G511gat_0[2]));
	jspl3 jspl3_w_G511gat_4(.douta(w_G511gat_4[0]),.doutb(w_G511gat_4[1]),.doutc(w_G511gat_4[2]),.din(w_G511gat_1[0]));
	jspl3 jspl3_w_G511gat_5(.douta(w_G511gat_5[0]),.doutb(w_G511gat_5[1]),.doutc(w_G511gat_5[2]),.din(w_G511gat_1[1]));
	jspl3 jspl3_w_G511gat_6(.douta(w_G511gat_6[0]),.doutb(w_G511gat_6[1]),.doutc(w_G511gat_6[2]),.din(w_G511gat_1[2]));
	jspl jspl_w_G511gat_7(.douta(w_G511gat_7[0]),.doutb(w_G511gat_7[1]),.din(w_G511gat_2[0]));
	jspl3 jspl3_w_G528gat_0(.douta(w_G528gat_0[0]),.doutb(w_G528gat_0[1]),.doutc(w_G528gat_0[2]),.din(G528gat));
	jspl3 jspl3_w_G528gat_1(.douta(w_G528gat_1[0]),.doutb(w_G528gat_1[1]),.doutc(w_G528gat_1[2]),.din(w_G528gat_0[0]));
	jspl3 jspl3_w_G528gat_2(.douta(w_G528gat_2[0]),.doutb(w_G528gat_2[1]),.doutc(w_G528gat_2[2]),.din(w_G528gat_0[1]));
	jspl3 jspl3_w_G528gat_3(.douta(w_G528gat_3[0]),.doutb(w_G528gat_3[1]),.doutc(w_G528gat_3[2]),.din(w_G528gat_0[2]));
	jspl3 jspl3_w_G528gat_4(.douta(w_G528gat_4[0]),.doutb(w_G528gat_4[1]),.doutc(w_G528gat_4[2]),.din(w_G528gat_1[0]));
	jspl3 jspl3_w_G528gat_5(.douta(w_G528gat_5[0]),.doutb(w_G528gat_5[1]),.doutc(w_G528gat_5[2]),.din(w_G528gat_1[1]));
	jspl3 jspl3_w_G528gat_6(.douta(w_G528gat_6[0]),.doutb(w_G528gat_6[1]),.doutc(w_G528gat_6[2]),.din(w_G528gat_1[2]));
	jspl jspl_w_G528gat_7(.douta(w_G528gat_7[0]),.doutb(w_G528gat_7[1]),.din(w_G528gat_2[0]));
	jspl jspl_w_G545gat_0(.douta(w_G545gat_0),.doutb(w_dff_A_rE4qmGgL3_1),.din(G545gat_fa_));
	jspl jspl_w_n65_0(.douta(w_n65_0[0]),.doutb(w_n65_0[1]),.din(n65));
	jspl jspl_w_n69_0(.douta(w_dff_A_uhOhIG0A7_0),.doutb(w_n69_0[1]),.din(n69));
	jspl jspl_w_n70_0(.douta(w_dff_A_nYOTDYLC5_0),.doutb(w_n70_0[1]),.din(n70));
	jspl jspl_w_n72_0(.douta(w_dff_A_MuhjVLNl5_0),.doutb(w_n72_0[1]),.din(n72));
	jspl jspl_w_n75_0(.douta(w_n75_0[0]),.doutb(w_n75_0[1]),.din(n75));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl jspl_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.din(n78));
	jspl jspl_w_n81_0(.douta(w_n81_0[0]),.doutb(w_n81_0[1]),.din(n81));
	jspl3 jspl3_w_n82_0(.douta(w_n82_0[0]),.doutb(w_dff_A_JJnjh7cr5_1),.doutc(w_dff_A_129vUXF14_2),.din(n82));
	jspl jspl_w_n82_1(.douta(w_n82_1[0]),.doutb(w_dff_A_3cslWXqh6_1),.din(w_n82_0[0]));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n85_0(.douta(w_dff_A_bcA037ij8_0),.doutb(w_n85_0[1]),.din(n85));
	jspl jspl_w_n87_0(.douta(w_n87_0[0]),.doutb(w_n87_0[1]),.din(n87));
	jspl jspl_w_n89_0(.douta(w_dff_A_JUvwpQwb8_0),.doutb(w_n89_0[1]),.din(n89));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl jspl_w_n94_0(.douta(w_dff_A_K0SsOrCV3_0),.doutb(w_n94_0[1]),.din(n94));
	jspl jspl_w_n96_0(.douta(w_n96_0[0]),.doutb(w_n96_0[1]),.din(n96));
	jspl jspl_w_n99_0(.douta(w_n99_0[0]),.doutb(w_n99_0[1]),.din(n99));
	jspl3 jspl3_w_n100_0(.douta(w_n100_0[0]),.doutb(w_dff_A_ixNCcfTv9_1),.doutc(w_dff_A_srC73IwU0_2),.din(n100));
	jspl jspl_w_n100_1(.douta(w_dff_A_avonoj9j1_0),.doutb(w_n100_1[1]),.din(w_n100_0[0]));
	jspl3 jspl3_w_n101_0(.douta(w_dff_A_1G0AuNFk3_0),.doutb(w_n101_0[1]),.doutc(w_n101_0[2]),.din(n101));
	jspl jspl_w_n103_0(.douta(w_dff_A_QvvnFDEe2_0),.doutb(w_n103_0[1]),.din(n103));
	jspl jspl_w_n104_0(.douta(w_dff_A_ykQi1sID8_0),.doutb(w_n104_0[1]),.din(n104));
	jspl jspl_w_n107_0(.douta(w_n107_0[0]),.doutb(w_dff_A_YXMU8p9c8_1),.din(n107));
	jspl jspl_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n110_0(.douta(w_dff_A_Tooep5n49_0),.doutb(w_n110_0[1]),.din(n110));
	jspl jspl_w_n115_0(.douta(w_n115_0[0]),.doutb(w_n115_0[1]),.din(n115));
	jspl jspl_w_n116_0(.douta(w_dff_A_lF7GCaFH7_0),.doutb(w_n116_0[1]),.din(n116));
	jspl3 jspl3_w_n126_0(.douta(w_n126_0[0]),.doutb(w_n126_0[1]),.doutc(w_n126_0[2]),.din(n126));
	jspl jspl_w_n128_0(.douta(w_n128_0[0]),.doutb(w_n128_0[1]),.din(w_dff_B_uXlhIgzZ4_2));
	jspl jspl_w_n129_0(.douta(w_n129_0[0]),.doutb(w_n129_0[1]),.din(n129));
	jspl jspl_w_n130_0(.douta(w_n130_0[0]),.doutb(w_dff_A_bcg8oVQH4_1),.din(n130));
	jspl jspl_w_n131_0(.douta(w_n131_0[0]),.doutb(w_n131_0[1]),.din(n131));
	jspl3 jspl3_w_n132_0(.douta(w_dff_A_g6UKxOzF8_0),.doutb(w_dff_A_5rzIXust7_1),.doutc(w_n132_0[2]),.din(n132));
	jspl3 jspl3_w_n133_0(.douta(w_n133_0[0]),.doutb(w_n133_0[1]),.doutc(w_n133_0[2]),.din(n133));
	jspl jspl_w_n138_0(.douta(w_n138_0[0]),.doutb(w_n138_0[1]),.din(n138));
	jspl jspl_w_n139_0(.douta(w_dff_A_SZD2cvwN7_0),.doutb(w_n139_0[1]),.din(n139));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl jspl_w_n142_0(.douta(w_n142_0[0]),.doutb(w_dff_A_VpV1Wt6x7_1),.din(n142));
	jspl jspl_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.din(n143));
	jspl jspl_w_n145_0(.douta(w_dff_A_0h3CobnG1_0),.doutb(w_n145_0[1]),.din(n145));
	jspl jspl_w_n150_0(.douta(w_n150_0[0]),.doutb(w_n150_0[1]),.din(n150));
	jspl jspl_w_n151_0(.douta(w_dff_A_VWcmwtMh6_0),.doutb(w_n151_0[1]),.din(n151));
	jspl3 jspl3_w_n156_0(.douta(w_n156_0[0]),.doutb(w_n156_0[1]),.doutc(w_n156_0[2]),.din(n156));
	jspl jspl_w_n158_0(.douta(w_n158_0[0]),.doutb(w_n158_0[1]),.din(w_dff_B_E9bULjDw7_2));
	jspl jspl_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.din(n163));
	jspl jspl_w_n165_0(.douta(w_n165_0[0]),.doutb(w_n165_0[1]),.din(w_dff_B_LYuZZ2cD3_2));
	jspl jspl_w_n166_0(.douta(w_n166_0[0]),.doutb(w_n166_0[1]),.din(n166));
	jspl jspl_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.din(n168));
	jspl3 jspl3_w_n169_0(.douta(w_dff_A_g6U8xrxE7_0),.doutb(w_dff_A_IX8YLItY8_1),.doutc(w_n169_0[2]),.din(n169));
	jspl jspl_w_n170_0(.douta(w_n170_0[0]),.doutb(w_n170_0[1]),.din(n170));
	jspl jspl_w_n172_0(.douta(w_n172_0[0]),.doutb(w_n172_0[1]),.din(n172));
	jspl jspl_w_n174_0(.douta(w_n174_0[0]),.doutb(w_n174_0[1]),.din(n174));
	jspl jspl_w_n175_0(.douta(w_n175_0[0]),.doutb(w_n175_0[1]),.din(w_dff_B_U2AtfufT8_2));
	jspl jspl_w_n176_0(.douta(w_n176_0[0]),.doutb(w_n176_0[1]),.din(n176));
	jspl jspl_w_n177_0(.douta(w_dff_A_m59HVWWN7_0),.doutb(w_n177_0[1]),.din(n177));
	jspl jspl_w_n178_0(.douta(w_n178_0[0]),.doutb(w_n178_0[1]),.din(n178));
	jspl jspl_w_n180_0(.douta(w_n180_0[0]),.doutb(w_dff_A_kqbN4kqC7_1),.din(n180));
	jspl jspl_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.din(n181));
	jspl jspl_w_n183_0(.douta(w_dff_A_Ond58uNP5_0),.doutb(w_n183_0[1]),.din(n183));
	jspl jspl_w_n188_0(.douta(w_n188_0[0]),.doutb(w_n188_0[1]),.din(n188));
	jspl jspl_w_n189_0(.douta(w_dff_A_E3uuICfZ1_0),.doutb(w_n189_0[1]),.din(n189));
	jspl3 jspl3_w_n194_0(.douta(w_n194_0[0]),.doutb(w_n194_0[1]),.doutc(w_n194_0[2]),.din(n194));
	jspl jspl_w_n196_0(.douta(w_n196_0[0]),.doutb(w_n196_0[1]),.din(w_dff_B_2BHgDr6f3_2));
	jspl jspl_w_n199_0(.douta(w_n199_0[0]),.doutb(w_n199_0[1]),.din(n199));
	jspl jspl_w_n201_0(.douta(w_n201_0[0]),.doutb(w_n201_0[1]),.din(w_dff_B_1YazrMbv9_2));
	jspl jspl_w_n204_0(.douta(w_n204_0[0]),.doutb(w_n204_0[1]),.din(n204));
	jspl jspl_w_n206_0(.douta(w_n206_0[0]),.doutb(w_n206_0[1]),.din(w_dff_B_psp5KmyI1_2));
	jspl jspl_w_n207_0(.douta(w_n207_0[0]),.doutb(w_n207_0[1]),.din(n207));
	jspl jspl_w_n209_0(.douta(w_n209_0[0]),.doutb(w_n209_0[1]),.din(n209));
	jspl3 jspl3_w_n210_0(.douta(w_n210_0[0]),.doutb(w_dff_A_pnxRAwe47_1),.doutc(w_dff_A_MHJ6KRGP1_2),.din(n210));
	jspl jspl_w_n210_1(.douta(w_dff_A_lY35Gf6q5_0),.doutb(w_n210_1[1]),.din(w_n210_0[0]));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_n213_0[1]),.din(n213));
	jspl jspl_w_n215_0(.douta(w_n215_0[0]),.doutb(w_n215_0[1]),.din(n215));
	jspl jspl_w_n216_0(.douta(w_n216_0[0]),.doutb(w_n216_0[1]),.din(w_dff_B_eHQGTVDo8_2));
	jspl jspl_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.din(n217));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.din(w_dff_B_Hwp7sJGy6_2));
	jspl jspl_w_n219_0(.douta(w_n219_0[0]),.doutb(w_n219_0[1]),.din(n219));
	jspl jspl_w_n220_0(.douta(w_dff_A_AGyhUYPC7_0),.doutb(w_n220_0[1]),.din(n220));
	jspl jspl_w_n221_0(.douta(w_n221_0[0]),.doutb(w_n221_0[1]),.din(n221));
	jspl jspl_w_n223_0(.douta(w_n223_0[0]),.doutb(w_dff_A_iWmMC9ts3_1),.din(n223));
	jspl jspl_w_n224_0(.douta(w_n224_0[0]),.doutb(w_n224_0[1]),.din(n224));
	jspl jspl_w_n226_0(.douta(w_dff_A_edGf9AFJ6_0),.doutb(w_n226_0[1]),.din(n226));
	jspl jspl_w_n231_0(.douta(w_n231_0[0]),.doutb(w_n231_0[1]),.din(n231));
	jspl jspl_w_n232_0(.douta(w_dff_A_Q4WRj3c35_0),.doutb(w_n232_0[1]),.din(n232));
	jspl3 jspl3_w_n237_0(.douta(w_n237_0[0]),.doutb(w_n237_0[1]),.doutc(w_n237_0[2]),.din(n237));
	jspl jspl_w_n239_0(.douta(w_n239_0[0]),.doutb(w_n239_0[1]),.din(w_dff_B_7t7VuDNg2_2));
	jspl jspl_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.din(n242));
	jspl jspl_w_n244_0(.douta(w_n244_0[0]),.doutb(w_n244_0[1]),.din(w_dff_B_Eevn5yIO0_2));
	jspl jspl_w_n247_0(.douta(w_n247_0[0]),.doutb(w_n247_0[1]),.din(n247));
	jspl jspl_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.din(w_dff_B_9cmf9K3G9_2));
	jspl jspl_w_n252_0(.douta(w_n252_0[0]),.doutb(w_n252_0[1]),.din(n252));
	jspl jspl_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.din(w_dff_B_Cjc6iVEW9_2));
	jspl jspl_w_n255_0(.douta(w_n255_0[0]),.doutb(w_n255_0[1]),.din(n255));
	jspl jspl_w_n257_0(.douta(w_n257_0[0]),.doutb(w_n257_0[1]),.din(n257));
	jspl3 jspl3_w_n258_0(.douta(w_dff_A_ND5nyXI76_0),.doutb(w_dff_A_oB75lPv25_1),.doutc(w_n258_0[2]),.din(n258));
	jspl jspl_w_n259_0(.douta(w_n259_0[0]),.doutb(w_n259_0[1]),.din(n259));
	jspl jspl_w_n261_0(.douta(w_n261_0[0]),.doutb(w_n261_0[1]),.din(n261));
	jspl jspl_w_n264_0(.douta(w_n264_0[0]),.doutb(w_n264_0[1]),.din(n264));
	jspl jspl_w_n265_0(.douta(w_n265_0[0]),.doutb(w_n265_0[1]),.din(w_dff_B_nalj3afZ5_2));
	jspl jspl_w_n266_0(.douta(w_n266_0[0]),.doutb(w_n266_0[1]),.din(n266));
	jspl jspl_w_n267_0(.douta(w_n267_0[0]),.doutb(w_n267_0[1]),.din(w_dff_B_HK1uxouA2_2));
	jspl jspl_w_n268_0(.douta(w_n268_0[0]),.doutb(w_n268_0[1]),.din(n268));
	jspl jspl_w_n269_0(.douta(w_n269_0[0]),.doutb(w_n269_0[1]),.din(w_dff_B_5WzUuFtq7_2));
	jspl jspl_w_n270_0(.douta(w_n270_0[0]),.doutb(w_n270_0[1]),.din(n270));
	jspl jspl_w_n271_0(.douta(w_dff_A_AoFzQpzy8_0),.doutb(w_n271_0[1]),.din(n271));
	jspl jspl_w_n272_0(.douta(w_n272_0[0]),.doutb(w_n272_0[1]),.din(n272));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_dff_A_tZxpkrLk3_1),.din(n274));
	jspl jspl_w_n275_0(.douta(w_n275_0[0]),.doutb(w_n275_0[1]),.din(n275));
	jspl jspl_w_n277_0(.douta(w_dff_A_eUbJdN5F3_0),.doutb(w_n277_0[1]),.din(n277));
	jspl jspl_w_n282_0(.douta(w_n282_0[0]),.doutb(w_n282_0[1]),.din(n282));
	jspl jspl_w_n283_0(.douta(w_dff_A_bWWMFQmV5_0),.doutb(w_n283_0[1]),.din(n283));
	jspl3 jspl3_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.doutc(w_n288_0[2]),.din(n288));
	jspl jspl_w_n290_0(.douta(w_n290_0[0]),.doutb(w_n290_0[1]),.din(w_dff_B_OnVhSGaU0_2));
	jspl jspl_w_n293_0(.douta(w_n293_0[0]),.doutb(w_n293_0[1]),.din(n293));
	jspl jspl_w_n295_0(.douta(w_n295_0[0]),.doutb(w_n295_0[1]),.din(w_dff_B_ZT1o73KG3_2));
	jspl jspl_w_n298_0(.douta(w_n298_0[0]),.doutb(w_n298_0[1]),.din(n298));
	jspl jspl_w_n300_0(.douta(w_n300_0[0]),.doutb(w_n300_0[1]),.din(w_dff_B_BMfrFhAf7_2));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.din(n303));
	jspl jspl_w_n305_0(.douta(w_n305_0[0]),.doutb(w_n305_0[1]),.din(w_dff_B_JqLKAmu29_2));
	jspl jspl_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.din(n308));
	jspl jspl_w_n310_0(.douta(w_n310_0[0]),.doutb(w_n310_0[1]),.din(w_dff_B_InSP26yk6_2));
	jspl jspl_w_n311_0(.douta(w_n311_0[0]),.doutb(w_n311_0[1]),.din(n311));
	jspl jspl_w_n313_0(.douta(w_n313_0[0]),.doutb(w_n313_0[1]),.din(n313));
	jspl3 jspl3_w_n314_0(.douta(w_dff_A_CWv4PehF4_0),.doutb(w_dff_A_IQZnHAAl3_1),.doutc(w_n314_0[2]),.din(n314));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl jspl_w_n317_0(.douta(w_n317_0[0]),.doutb(w_n317_0[1]),.din(n317));
	jspl jspl_w_n320_0(.douta(w_n320_0[0]),.doutb(w_n320_0[1]),.din(n320));
	jspl jspl_w_n321_0(.douta(w_n321_0[0]),.doutb(w_n321_0[1]),.din(w_dff_B_NxEO5AfJ9_2));
	jspl jspl_w_n322_0(.douta(w_n322_0[0]),.doutb(w_n322_0[1]),.din(n322));
	jspl jspl_w_n323_0(.douta(w_n323_0[0]),.doutb(w_n323_0[1]),.din(w_dff_B_cFedhM6m6_2));
	jspl jspl_w_n324_0(.douta(w_n324_0[0]),.doutb(w_n324_0[1]),.din(n324));
	jspl jspl_w_n325_0(.douta(w_n325_0[0]),.doutb(w_n325_0[1]),.din(w_dff_B_Pwl0RWjL6_2));
	jspl jspl_w_n326_0(.douta(w_n326_0[0]),.doutb(w_n326_0[1]),.din(n326));
	jspl jspl_w_n327_0(.douta(w_n327_0[0]),.doutb(w_n327_0[1]),.din(w_dff_B_Flxa6Eko8_2));
	jspl jspl_w_n328_0(.douta(w_n328_0[0]),.doutb(w_n328_0[1]),.din(n328));
	jspl jspl_w_n329_0(.douta(w_dff_A_vOuZa3lL8_0),.doutb(w_n329_0[1]),.din(n329));
	jspl jspl_w_n330_0(.douta(w_n330_0[0]),.doutb(w_n330_0[1]),.din(n330));
	jspl jspl_w_n332_0(.douta(w_n332_0[0]),.doutb(w_dff_A_peHk2qng5_1),.din(n332));
	jspl jspl_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.din(n333));
	jspl jspl_w_n335_0(.douta(w_dff_A_t8tAzgMp1_0),.doutb(w_n335_0[1]),.din(n335));
	jspl jspl_w_n340_0(.douta(w_n340_0[0]),.doutb(w_n340_0[1]),.din(n340));
	jspl jspl_w_n341_0(.douta(w_dff_A_F7GGot049_0),.doutb(w_n341_0[1]),.din(n341));
	jspl3 jspl3_w_n346_0(.douta(w_n346_0[0]),.doutb(w_n346_0[1]),.doutc(w_n346_0[2]),.din(n346));
	jspl jspl_w_n348_0(.douta(w_n348_0[0]),.doutb(w_n348_0[1]),.din(w_dff_B_Jv3A2qaZ9_2));
	jspl jspl_w_n351_0(.douta(w_n351_0[0]),.doutb(w_n351_0[1]),.din(n351));
	jspl jspl_w_n353_0(.douta(w_n353_0[0]),.doutb(w_n353_0[1]),.din(w_dff_B_VzlPzLz94_2));
	jspl jspl_w_n356_0(.douta(w_n356_0[0]),.doutb(w_n356_0[1]),.din(n356));
	jspl jspl_w_n358_0(.douta(w_n358_0[0]),.doutb(w_n358_0[1]),.din(w_dff_B_TCa8Nxe60_2));
	jspl jspl_w_n361_0(.douta(w_n361_0[0]),.doutb(w_n361_0[1]),.din(n361));
	jspl jspl_w_n363_0(.douta(w_n363_0[0]),.doutb(w_n363_0[1]),.din(w_dff_B_wVO3rB1a0_2));
	jspl jspl_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.din(n366));
	jspl jspl_w_n368_0(.douta(w_n368_0[0]),.doutb(w_n368_0[1]),.din(w_dff_B_xUKku5GK7_2));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.din(n371));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_dff_A_AlngDwTI8_1),.din(n372));
	jspl jspl_w_n373_0(.douta(w_n373_0[0]),.doutb(w_n373_0[1]),.din(n373));
	jspl jspl_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.din(n375));
	jspl3 jspl3_w_n376_0(.douta(w_dff_A_OqaIikFK2_0),.doutb(w_dff_A_RVoeUevc7_1),.doutc(w_n376_0[2]),.din(n376));
	jspl jspl_w_n377_0(.douta(w_n377_0[0]),.doutb(w_n377_0[1]),.din(n377));
	jspl jspl_w_n380_0(.douta(w_dff_A_CFnGIAnQ4_0),.doutb(w_n380_0[1]),.din(n380));
	jspl jspl_w_n382_0(.douta(w_n382_0[0]),.doutb(w_n382_0[1]),.din(n382));
	jspl jspl_w_n383_0(.douta(w_n383_0[0]),.doutb(w_n383_0[1]),.din(n383));
	jspl jspl_w_n384_0(.douta(w_n384_0[0]),.doutb(w_n384_0[1]),.din(n384));
	jspl jspl_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.din(w_dff_B_OOIwGHPY4_2));
	jspl jspl_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.din(n386));
	jspl jspl_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.din(w_dff_B_nnVOysn11_2));
	jspl jspl_w_n388_0(.douta(w_n388_0[0]),.doutb(w_n388_0[1]),.din(n388));
	jspl jspl_w_n389_0(.douta(w_n389_0[0]),.doutb(w_n389_0[1]),.din(w_dff_B_eVcoFSmM5_2));
	jspl jspl_w_n390_0(.douta(w_n390_0[0]),.doutb(w_n390_0[1]),.din(n390));
	jspl jspl_w_n391_0(.douta(w_n391_0[0]),.doutb(w_n391_0[1]),.din(w_dff_B_rbZL3TVO2_2));
	jspl jspl_w_n392_0(.douta(w_n392_0[0]),.doutb(w_n392_0[1]),.din(n392));
	jspl jspl_w_n393_0(.douta(w_dff_A_H5a6kMnc7_0),.doutb(w_n393_0[1]),.din(n393));
	jspl jspl_w_n394_0(.douta(w_n394_0[0]),.doutb(w_n394_0[1]),.din(n394));
	jspl jspl_w_n396_0(.douta(w_n396_0[0]),.doutb(w_dff_A_CHZGfPAc5_1),.din(n396));
	jspl jspl_w_n397_0(.douta(w_n397_0[0]),.doutb(w_n397_0[1]),.din(n397));
	jspl jspl_w_n399_0(.douta(w_dff_A_Bh1ZRL9E6_0),.doutb(w_n399_0[1]),.din(n399));
	jspl jspl_w_n404_0(.douta(w_n404_0[0]),.doutb(w_n404_0[1]),.din(n404));
	jspl jspl_w_n405_0(.douta(w_dff_A_pPk0ZHij9_0),.doutb(w_n405_0[1]),.din(n405));
	jspl3 jspl3_w_n410_0(.douta(w_n410_0[0]),.doutb(w_n410_0[1]),.doutc(w_n410_0[2]),.din(n410));
	jspl jspl_w_n412_0(.douta(w_n412_0[0]),.doutb(w_n412_0[1]),.din(w_dff_B_B1MHIwkE4_2));
	jspl jspl_w_n415_0(.douta(w_n415_0[0]),.doutb(w_n415_0[1]),.din(n415));
	jspl jspl_w_n417_0(.douta(w_n417_0[0]),.doutb(w_n417_0[1]),.din(w_dff_B_OMGyWvRk1_2));
	jspl jspl_w_n420_0(.douta(w_n420_0[0]),.doutb(w_n420_0[1]),.din(n420));
	jspl jspl_w_n422_0(.douta(w_n422_0[0]),.doutb(w_n422_0[1]),.din(w_dff_B_RNkWNosq9_2));
	jspl jspl_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.din(n425));
	jspl jspl_w_n427_0(.douta(w_n427_0[0]),.doutb(w_n427_0[1]),.din(w_dff_B_WVEh5NPZ2_2));
	jspl jspl_w_n430_0(.douta(w_n430_0[0]),.doutb(w_n430_0[1]),.din(n430));
	jspl jspl_w_n432_0(.douta(w_n432_0[0]),.doutb(w_n432_0[1]),.din(w_dff_B_t22o2eFd8_2));
	jspl jspl_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.din(w_dff_B_1TPbLWoN5_2));
	jspl jspl_w_n437_0(.douta(w_n437_0[0]),.doutb(w_n437_0[1]),.din(w_dff_B_j23U0sOR6_2));
	jspl jspl_w_n441_0(.douta(w_n441_0[0]),.doutb(w_n441_0[1]),.din(n441));
	jspl jspl_w_n442_0(.douta(w_n442_0[0]),.doutb(w_dff_A_mAPv3Wu33_1),.din(n442));
	jspl jspl_w_n443_0(.douta(w_n443_0[0]),.doutb(w_n443_0[1]),.din(n443));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl3 jspl3_w_n446_0(.douta(w_dff_A_VEjDMFPq4_0),.doutb(w_dff_A_DzAcwloZ4_1),.doutc(w_n446_0[2]),.din(n446));
	jspl jspl_w_n447_0(.douta(w_n447_0[0]),.doutb(w_n447_0[1]),.din(n447));
	jspl jspl_w_n450_0(.douta(w_dff_A_PzvLBQM62_0),.doutb(w_n450_0[1]),.din(n450));
	jspl jspl_w_n452_0(.douta(w_n452_0[0]),.doutb(w_n452_0[1]),.din(n452));
	jspl jspl_w_n453_0(.douta(w_n453_0[0]),.doutb(w_n453_0[1]),.din(w_dff_B_ugK7QYqi7_2));
	jspl jspl_w_n454_0(.douta(w_n454_0[0]),.doutb(w_n454_0[1]),.din(n454));
	jspl jspl_w_n455_0(.douta(w_n455_0[0]),.doutb(w_n455_0[1]),.din(n455));
	jspl jspl_w_n456_0(.douta(w_n456_0[0]),.doutb(w_n456_0[1]),.din(n456));
	jspl jspl_w_n457_0(.douta(w_n457_0[0]),.doutb(w_n457_0[1]),.din(n457));
	jspl jspl_w_n458_0(.douta(w_n458_0[0]),.doutb(w_n458_0[1]),.din(n458));
	jspl jspl_w_n459_0(.douta(w_n459_0[0]),.doutb(w_n459_0[1]),.din(w_dff_B_J6QBkd1c4_2));
	jspl jspl_w_n460_0(.douta(w_n460_0[0]),.doutb(w_n460_0[1]),.din(n460));
	jspl jspl_w_n461_0(.douta(w_n461_0[0]),.doutb(w_n461_0[1]),.din(w_dff_B_oiv1Ej0a7_2));
	jspl jspl_w_n462_0(.douta(w_n462_0[0]),.doutb(w_n462_0[1]),.din(n462));
	jspl jspl_w_n463_0(.douta(w_n463_0[0]),.doutb(w_n463_0[1]),.din(w_dff_B_oai99Er00_2));
	jspl jspl_w_n464_0(.douta(w_n464_0[0]),.doutb(w_n464_0[1]),.din(n464));
	jspl jspl_w_n465_0(.douta(w_dff_A_w7T9nth90_0),.doutb(w_n465_0[1]),.din(n465));
	jspl jspl_w_n466_0(.douta(w_n466_0[0]),.doutb(w_n466_0[1]),.din(n466));
	jspl jspl_w_n468_0(.douta(w_n468_0[0]),.doutb(w_dff_A_CjzJvrro2_1),.din(n468));
	jspl jspl_w_n469_0(.douta(w_n469_0[0]),.doutb(w_n469_0[1]),.din(n469));
	jspl jspl_w_n471_0(.douta(w_dff_A_QyYqNGcL2_0),.doutb(w_n471_0[1]),.din(n471));
	jspl jspl_w_n476_0(.douta(w_n476_0[0]),.doutb(w_n476_0[1]),.din(n476));
	jspl jspl_w_n477_0(.douta(w_dff_A_UZ7DrGWN9_0),.doutb(w_n477_0[1]),.din(n477));
	jspl3 jspl3_w_n482_0(.douta(w_n482_0[0]),.doutb(w_n482_0[1]),.doutc(w_n482_0[2]),.din(n482));
	jspl jspl_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.din(w_dff_B_YZsqRtp03_2));
	jspl jspl_w_n487_0(.douta(w_n487_0[0]),.doutb(w_n487_0[1]),.din(n487));
	jspl jspl_w_n489_0(.douta(w_n489_0[0]),.doutb(w_n489_0[1]),.din(w_dff_B_fS3wTcsS6_2));
	jspl jspl_w_n492_0(.douta(w_n492_0[0]),.doutb(w_n492_0[1]),.din(n492));
	jspl jspl_w_n494_0(.douta(w_n494_0[0]),.doutb(w_n494_0[1]),.din(w_dff_B_A3MxRWOn7_2));
	jspl jspl_w_n497_0(.douta(w_n497_0[0]),.doutb(w_n497_0[1]),.din(n497));
	jspl jspl_w_n499_0(.douta(w_n499_0[0]),.doutb(w_n499_0[1]),.din(w_dff_B_1WJwsVqu8_2));
	jspl jspl_w_n502_0(.douta(w_n502_0[0]),.doutb(w_n502_0[1]),.din(n502));
	jspl jspl_w_n504_0(.douta(w_n504_0[0]),.doutb(w_n504_0[1]),.din(w_dff_B_4A2pXL0w9_2));
	jspl jspl_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.din(n507));
	jspl jspl_w_n509_0(.douta(w_n509_0[0]),.doutb(w_n509_0[1]),.din(w_dff_B_StDSFw8h8_2));
	jspl jspl_w_n512_0(.douta(w_n512_0[0]),.doutb(w_n512_0[1]),.din(n512));
	jspl jspl_w_n514_0(.douta(w_n514_0[0]),.doutb(w_n514_0[1]),.din(w_dff_B_aWyavlEF5_2));
	jspl jspl_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.din(n518));
	jspl jspl_w_n519_0(.douta(w_n519_0[0]),.doutb(w_dff_A_6STtgGwI6_1),.din(n519));
	jspl jspl_w_n520_0(.douta(w_n520_0[0]),.doutb(w_n520_0[1]),.din(n520));
	jspl jspl_w_n522_0(.douta(w_n522_0[0]),.doutb(w_n522_0[1]),.din(n522));
	jspl3 jspl3_w_n523_0(.douta(w_dff_A_8UhmKZc75_0),.doutb(w_dff_A_NfLo46A38_1),.doutc(w_n523_0[2]),.din(n523));
	jspl jspl_w_n524_0(.douta(w_n524_0[0]),.doutb(w_n524_0[1]),.din(n524));
	jspl jspl_w_n527_0(.douta(w_dff_A_BnbUiBaX3_0),.doutb(w_n527_0[1]),.din(n527));
	jspl jspl_w_n529_0(.douta(w_n529_0[0]),.doutb(w_n529_0[1]),.din(n529));
	jspl jspl_w_n530_0(.douta(w_n530_0[0]),.doutb(w_n530_0[1]),.din(w_dff_B_QiWXyrP18_2));
	jspl jspl_w_n531_0(.douta(w_n531_0[0]),.doutb(w_n531_0[1]),.din(n531));
	jspl jspl_w_n532_0(.douta(w_n532_0[0]),.doutb(w_n532_0[1]),.din(w_dff_B_CVnLg0kR4_2));
	jspl jspl_w_n533_0(.douta(w_n533_0[0]),.doutb(w_n533_0[1]),.din(n533));
	jspl jspl_w_n534_0(.douta(w_n534_0[0]),.doutb(w_n534_0[1]),.din(n534));
	jspl jspl_w_n535_0(.douta(w_n535_0[0]),.doutb(w_n535_0[1]),.din(n535));
	jspl jspl_w_n536_0(.douta(w_n536_0[0]),.doutb(w_n536_0[1]),.din(n536));
	jspl jspl_w_n537_0(.douta(w_n537_0[0]),.doutb(w_n537_0[1]),.din(n537));
	jspl jspl_w_n538_0(.douta(w_n538_0[0]),.doutb(w_n538_0[1]),.din(w_dff_B_DFyyoA0N0_2));
	jspl jspl_w_n539_0(.douta(w_n539_0[0]),.doutb(w_n539_0[1]),.din(n539));
	jspl jspl_w_n540_0(.douta(w_n540_0[0]),.doutb(w_n540_0[1]),.din(w_dff_B_SXqyNsLN2_2));
	jspl jspl_w_n541_0(.douta(w_n541_0[0]),.doutb(w_n541_0[1]),.din(n541));
	jspl jspl_w_n542_0(.douta(w_n542_0[0]),.doutb(w_n542_0[1]),.din(w_dff_B_ahnDQaUE2_2));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_n543_0[1]),.din(n543));
	jspl jspl_w_n544_0(.douta(w_dff_A_8tiOknIL2_0),.doutb(w_n544_0[1]),.din(n544));
	jspl jspl_w_n545_0(.douta(w_n545_0[0]),.doutb(w_n545_0[1]),.din(n545));
	jspl jspl_w_n547_0(.douta(w_n547_0[0]),.doutb(w_dff_A_y52OnWIm4_1),.din(n547));
	jspl jspl_w_n548_0(.douta(w_n548_0[0]),.doutb(w_n548_0[1]),.din(n548));
	jspl jspl_w_n550_0(.douta(w_dff_A_U6tTMT4n6_0),.doutb(w_n550_0[1]),.din(n550));
	jspl jspl_w_n555_0(.douta(w_n555_0[0]),.doutb(w_n555_0[1]),.din(n555));
	jspl jspl_w_n556_0(.douta(w_dff_A_4Sqb3nNa1_0),.doutb(w_n556_0[1]),.din(n556));
	jspl3 jspl3_w_n561_0(.douta(w_n561_0[0]),.doutb(w_n561_0[1]),.doutc(w_n561_0[2]),.din(n561));
	jspl jspl_w_n563_0(.douta(w_n563_0[0]),.doutb(w_n563_0[1]),.din(w_dff_B_IqjvnNs23_2));
	jspl jspl_w_n566_0(.douta(w_n566_0[0]),.doutb(w_n566_0[1]),.din(n566));
	jspl jspl_w_n568_0(.douta(w_n568_0[0]),.doutb(w_n568_0[1]),.din(w_dff_B_tVGUx8Nc5_2));
	jspl jspl_w_n571_0(.douta(w_n571_0[0]),.doutb(w_n571_0[1]),.din(n571));
	jspl jspl_w_n573_0(.douta(w_n573_0[0]),.doutb(w_n573_0[1]),.din(w_dff_B_DGBVxjsn9_2));
	jspl jspl_w_n576_0(.douta(w_n576_0[0]),.doutb(w_n576_0[1]),.din(n576));
	jspl jspl_w_n578_0(.douta(w_n578_0[0]),.doutb(w_n578_0[1]),.din(w_dff_B_qqduDE2g4_2));
	jspl jspl_w_n581_0(.douta(w_n581_0[0]),.doutb(w_n581_0[1]),.din(n581));
	jspl jspl_w_n583_0(.douta(w_n583_0[0]),.doutb(w_n583_0[1]),.din(w_dff_B_8w35Olta4_2));
	jspl jspl_w_n586_0(.douta(w_n586_0[0]),.doutb(w_n586_0[1]),.din(n586));
	jspl jspl_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.din(w_dff_B_N4qhkeI07_2));
	jspl jspl_w_n591_0(.douta(w_n591_0[0]),.doutb(w_n591_0[1]),.din(n591));
	jspl jspl_w_n593_0(.douta(w_n593_0[0]),.doutb(w_n593_0[1]),.din(w_dff_B_DbqvFnC43_2));
	jspl jspl_w_n596_0(.douta(w_n596_0[0]),.doutb(w_n596_0[1]),.din(n596));
	jspl jspl_w_n598_0(.douta(w_n598_0[0]),.doutb(w_n598_0[1]),.din(w_dff_B_jZe4YHWU3_2));
	jspl jspl_w_n602_0(.douta(w_n602_0[0]),.doutb(w_n602_0[1]),.din(n602));
	jspl jspl_w_n603_0(.douta(w_n603_0[0]),.doutb(w_dff_A_7lPIcV558_1),.din(n603));
	jspl jspl_w_n604_0(.douta(w_n604_0[0]),.doutb(w_n604_0[1]),.din(n604));
	jspl jspl_w_n606_0(.douta(w_n606_0[0]),.doutb(w_n606_0[1]),.din(n606));
	jspl3 jspl3_w_n607_0(.douta(w_dff_A_Ai6ny8Yz9_0),.doutb(w_dff_A_MUWNUiji3_1),.doutc(w_n607_0[2]),.din(n607));
	jspl jspl_w_n608_0(.douta(w_n608_0[0]),.doutb(w_n608_0[1]),.din(n608));
	jspl jspl_w_n611_0(.douta(w_dff_A_DwgwG6gr1_0),.doutb(w_n611_0[1]),.din(n611));
	jspl jspl_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.din(n613));
	jspl jspl_w_n614_0(.douta(w_n614_0[0]),.doutb(w_n614_0[1]),.din(w_dff_B_Y11zjUIr9_2));
	jspl jspl_w_n615_0(.douta(w_n615_0[0]),.doutb(w_n615_0[1]),.din(n615));
	jspl jspl_w_n616_0(.douta(w_n616_0[0]),.doutb(w_n616_0[1]),.din(w_dff_B_oy8umolf6_2));
	jspl jspl_w_n617_0(.douta(w_n617_0[0]),.doutb(w_n617_0[1]),.din(n617));
	jspl jspl_w_n618_0(.douta(w_n618_0[0]),.doutb(w_n618_0[1]),.din(w_dff_B_rldC3BJ47_2));
	jspl jspl_w_n619_0(.douta(w_n619_0[0]),.doutb(w_n619_0[1]),.din(n619));
	jspl jspl_w_n620_0(.douta(w_n620_0[0]),.doutb(w_n620_0[1]),.din(n620));
	jspl jspl_w_n621_0(.douta(w_n621_0[0]),.doutb(w_n621_0[1]),.din(n621));
	jspl jspl_w_n622_0(.douta(w_n622_0[0]),.doutb(w_n622_0[1]),.din(n622));
	jspl jspl_w_n623_0(.douta(w_n623_0[0]),.doutb(w_n623_0[1]),.din(n623));
	jspl jspl_w_n624_0(.douta(w_n624_0[0]),.doutb(w_n624_0[1]),.din(w_dff_B_vZ6KDoV16_2));
	jspl jspl_w_n625_0(.douta(w_n625_0[0]),.doutb(w_n625_0[1]),.din(n625));
	jspl jspl_w_n626_0(.douta(w_n626_0[0]),.doutb(w_n626_0[1]),.din(w_dff_B_KPzLWWr84_2));
	jspl jspl_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.din(n627));
	jspl jspl_w_n628_0(.douta(w_n628_0[0]),.doutb(w_n628_0[1]),.din(w_dff_B_A0EP2u038_2));
	jspl jspl_w_n629_0(.douta(w_n629_0[0]),.doutb(w_n629_0[1]),.din(n629));
	jspl jspl_w_n630_0(.douta(w_dff_A_5WYeOW9D8_0),.doutb(w_n630_0[1]),.din(n630));
	jspl jspl_w_n631_0(.douta(w_n631_0[0]),.doutb(w_n631_0[1]),.din(n631));
	jspl jspl_w_n633_0(.douta(w_n633_0[0]),.doutb(w_dff_A_aPxlJXc64_1),.din(n633));
	jspl jspl_w_n634_0(.douta(w_n634_0[0]),.doutb(w_n634_0[1]),.din(n634));
	jspl jspl_w_n636_0(.douta(w_dff_A_MyPZGV0G3_0),.doutb(w_n636_0[1]),.din(n636));
	jspl jspl_w_n641_0(.douta(w_n641_0[0]),.doutb(w_n641_0[1]),.din(n641));
	jspl jspl_w_n642_0(.douta(w_dff_A_1KDVfjr33_0),.doutb(w_n642_0[1]),.din(n642));
	jspl3 jspl3_w_n647_0(.douta(w_n647_0[0]),.doutb(w_n647_0[1]),.doutc(w_n647_0[2]),.din(n647));
	jspl jspl_w_n649_0(.douta(w_n649_0[0]),.doutb(w_n649_0[1]),.din(w_dff_B_ZYWG448Y6_2));
	jspl jspl_w_n652_0(.douta(w_n652_0[0]),.doutb(w_n652_0[1]),.din(n652));
	jspl jspl_w_n654_0(.douta(w_n654_0[0]),.doutb(w_n654_0[1]),.din(w_dff_B_ovFfKiA53_2));
	jspl jspl_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.din(n657));
	jspl jspl_w_n659_0(.douta(w_n659_0[0]),.doutb(w_n659_0[1]),.din(w_dff_B_UDGVpLg17_2));
	jspl jspl_w_n662_0(.douta(w_n662_0[0]),.doutb(w_n662_0[1]),.din(n662));
	jspl jspl_w_n664_0(.douta(w_n664_0[0]),.doutb(w_n664_0[1]),.din(w_dff_B_QpjVlIc90_2));
	jspl jspl_w_n667_0(.douta(w_n667_0[0]),.doutb(w_n667_0[1]),.din(n667));
	jspl jspl_w_n669_0(.douta(w_n669_0[0]),.doutb(w_n669_0[1]),.din(w_dff_B_BUOFNaTh0_2));
	jspl jspl_w_n672_0(.douta(w_n672_0[0]),.doutb(w_n672_0[1]),.din(n672));
	jspl jspl_w_n674_0(.douta(w_n674_0[0]),.doutb(w_n674_0[1]),.din(w_dff_B_sWjd90256_2));
	jspl jspl_w_n677_0(.douta(w_n677_0[0]),.doutb(w_n677_0[1]),.din(n677));
	jspl jspl_w_n679_0(.douta(w_n679_0[0]),.doutb(w_n679_0[1]),.din(w_dff_B_TGg6KFiC7_2));
	jspl jspl_w_n682_0(.douta(w_n682_0[0]),.doutb(w_n682_0[1]),.din(n682));
	jspl jspl_w_n684_0(.douta(w_n684_0[0]),.doutb(w_n684_0[1]),.din(w_dff_B_7W6IBFpX8_2));
	jspl jspl_w_n687_0(.douta(w_n687_0[0]),.doutb(w_n687_0[1]),.din(n687));
	jspl jspl_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.din(w_dff_B_PumEGzma6_2));
	jspl jspl_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.din(n693));
	jspl jspl_w_n694_0(.douta(w_n694_0[0]),.doutb(w_dff_A_bBP3iweD3_1),.din(n694));
	jspl3 jspl3_w_n695_0(.douta(w_dff_A_VCHMQp1s7_0),.doutb(w_n695_0[1]),.doutc(w_n695_0[2]),.din(n695));
	jspl jspl_w_n697_0(.douta(w_n697_0[0]),.doutb(w_n697_0[1]),.din(n697));
	jspl3 jspl3_w_n698_0(.douta(w_dff_A_PWnxLbLl4_0),.doutb(w_dff_A_j2EXnS4j2_1),.doutc(w_n698_0[2]),.din(n698));
	jspl jspl_w_n699_0(.douta(w_n699_0[0]),.doutb(w_n699_0[1]),.din(n699));
	jspl jspl_w_n702_0(.douta(w_dff_A_LRlOYx2p2_0),.doutb(w_n702_0[1]),.din(n702));
	jspl jspl_w_n704_0(.douta(w_n704_0[0]),.doutb(w_n704_0[1]),.din(n704));
	jspl jspl_w_n705_0(.douta(w_n705_0[0]),.doutb(w_n705_0[1]),.din(w_dff_B_GTmP2KeA8_2));
	jspl jspl_w_n706_0(.douta(w_n706_0[0]),.doutb(w_n706_0[1]),.din(n706));
	jspl jspl_w_n707_0(.douta(w_n707_0[0]),.doutb(w_n707_0[1]),.din(w_dff_B_Q5STwsBo3_2));
	jspl jspl_w_n708_0(.douta(w_n708_0[0]),.doutb(w_n708_0[1]),.din(n708));
	jspl jspl_w_n709_0(.douta(w_n709_0[0]),.doutb(w_n709_0[1]),.din(w_dff_B_4fGVicy57_2));
	jspl jspl_w_n710_0(.douta(w_n710_0[0]),.doutb(w_n710_0[1]),.din(n710));
	jspl jspl_w_n711_0(.douta(w_n711_0[0]),.doutb(w_n711_0[1]),.din(w_dff_B_RHR0rDDN0_2));
	jspl jspl_w_n712_0(.douta(w_n712_0[0]),.doutb(w_n712_0[1]),.din(n712));
	jspl jspl_w_n713_0(.douta(w_n713_0[0]),.doutb(w_n713_0[1]),.din(n713));
	jspl jspl_w_n714_0(.douta(w_n714_0[0]),.doutb(w_n714_0[1]),.din(n714));
	jspl jspl_w_n715_0(.douta(w_n715_0[0]),.doutb(w_n715_0[1]),.din(n715));
	jspl jspl_w_n716_0(.douta(w_n716_0[0]),.doutb(w_n716_0[1]),.din(n716));
	jspl jspl_w_n717_0(.douta(w_n717_0[0]),.doutb(w_n717_0[1]),.din(w_dff_B_ycB40T2b3_2));
	jspl jspl_w_n718_0(.douta(w_n718_0[0]),.doutb(w_n718_0[1]),.din(n718));
	jspl jspl_w_n719_0(.douta(w_n719_0[0]),.doutb(w_n719_0[1]),.din(w_dff_B_LjFoFNip1_2));
	jspl jspl_w_n720_0(.douta(w_n720_0[0]),.doutb(w_n720_0[1]),.din(n720));
	jspl jspl_w_n721_0(.douta(w_n721_0[0]),.doutb(w_n721_0[1]),.din(w_dff_B_XMyO4VcL9_2));
	jspl jspl_w_n722_0(.douta(w_n722_0[0]),.doutb(w_n722_0[1]),.din(n722));
	jspl jspl_w_n723_0(.douta(w_dff_A_OgeeSzwv6_0),.doutb(w_n723_0[1]),.din(n723));
	jspl jspl_w_n724_0(.douta(w_n724_0[0]),.doutb(w_n724_0[1]),.din(n724));
	jspl jspl_w_n726_0(.douta(w_n726_0[0]),.doutb(w_dff_A_hATT4C2w2_1),.din(n726));
	jspl jspl_w_n727_0(.douta(w_n727_0[0]),.doutb(w_n727_0[1]),.din(n727));
	jspl jspl_w_n729_0(.douta(w_dff_A_O44AF8rm8_0),.doutb(w_n729_0[1]),.din(n729));
	jspl jspl_w_n734_0(.douta(w_n734_0[0]),.doutb(w_n734_0[1]),.din(n734));
	jspl jspl_w_n735_0(.douta(w_dff_A_7YxzHdl95_0),.doutb(w_n735_0[1]),.din(n735));
	jspl3 jspl3_w_n740_0(.douta(w_n740_0[0]),.doutb(w_n740_0[1]),.doutc(w_n740_0[2]),.din(n740));
	jspl jspl_w_n742_0(.douta(w_n742_0[0]),.doutb(w_n742_0[1]),.din(w_dff_B_CGzaqclw9_2));
	jspl jspl_w_n745_0(.douta(w_n745_0[0]),.doutb(w_n745_0[1]),.din(n745));
	jspl jspl_w_n747_0(.douta(w_n747_0[0]),.doutb(w_n747_0[1]),.din(w_dff_B_HMm1T04d9_2));
	jspl jspl_w_n750_0(.douta(w_n750_0[0]),.doutb(w_n750_0[1]),.din(n750));
	jspl jspl_w_n752_0(.douta(w_n752_0[0]),.doutb(w_n752_0[1]),.din(w_dff_B_fj8Vgs8k0_2));
	jspl jspl_w_n755_0(.douta(w_n755_0[0]),.doutb(w_n755_0[1]),.din(n755));
	jspl jspl_w_n757_0(.douta(w_n757_0[0]),.doutb(w_n757_0[1]),.din(w_dff_B_zR9qlZKD4_2));
	jspl jspl_w_n760_0(.douta(w_n760_0[0]),.doutb(w_n760_0[1]),.din(n760));
	jspl jspl_w_n762_0(.douta(w_n762_0[0]),.doutb(w_n762_0[1]),.din(w_dff_B_GrOGSWfp7_2));
	jspl jspl_w_n765_0(.douta(w_n765_0[0]),.doutb(w_n765_0[1]),.din(n765));
	jspl jspl_w_n767_0(.douta(w_n767_0[0]),.doutb(w_n767_0[1]),.din(w_dff_B_NJq9Mwmv8_2));
	jspl jspl_w_n770_0(.douta(w_n770_0[0]),.doutb(w_n770_0[1]),.din(n770));
	jspl jspl_w_n772_0(.douta(w_n772_0[0]),.doutb(w_n772_0[1]),.din(w_dff_B_BcXpF4rI7_2));
	jspl jspl_w_n775_0(.douta(w_n775_0[0]),.doutb(w_n775_0[1]),.din(n775));
	jspl jspl_w_n777_0(.douta(w_n777_0[0]),.doutb(w_n777_0[1]),.din(w_dff_B_dOQjWle73_2));
	jspl jspl_w_n780_0(.douta(w_n780_0[0]),.doutb(w_n780_0[1]),.din(n780));
	jspl jspl_w_n782_0(.douta(w_n782_0[0]),.doutb(w_n782_0[1]),.din(w_dff_B_Fx7TQE1T8_2));
	jspl jspl_w_n785_0(.douta(w_n785_0[0]),.doutb(w_n785_0[1]),.din(n785));
	jspl jspl_w_n787_0(.douta(w_n787_0[0]),.doutb(w_n787_0[1]),.din(w_dff_B_4LFn6EgN7_2));
	jspl jspl_w_n791_0(.douta(w_n791_0[0]),.doutb(w_n791_0[1]),.din(n791));
	jspl jspl_w_n792_0(.douta(w_n792_0[0]),.doutb(w_dff_A_YFE1FYKA7_1),.din(n792));
	jspl jspl_w_n793_0(.douta(w_dff_A_uVjBeraU8_0),.doutb(w_n793_0[1]),.din(n793));
	jspl jspl_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.din(n795));
	jspl3 jspl3_w_n797_0(.douta(w_n797_0[0]),.doutb(w_n797_0[1]),.doutc(w_n797_0[2]),.din(n797));
	jspl jspl_w_n800_0(.douta(w_dff_A_xxdJDKKt3_0),.doutb(w_n800_0[1]),.din(n800));
	jspl jspl_w_n802_0(.douta(w_n802_0[0]),.doutb(w_n802_0[1]),.din(n802));
	jspl jspl_w_n803_0(.douta(w_n803_0[0]),.doutb(w_n803_0[1]),.din(w_dff_B_nzwKRckY6_2));
	jspl jspl_w_n804_0(.douta(w_n804_0[0]),.doutb(w_n804_0[1]),.din(n804));
	jspl jspl_w_n805_0(.douta(w_n805_0[0]),.doutb(w_n805_0[1]),.din(w_dff_B_tWtJj8lm3_2));
	jspl jspl_w_n806_0(.douta(w_n806_0[0]),.doutb(w_n806_0[1]),.din(n806));
	jspl jspl_w_n807_0(.douta(w_n807_0[0]),.doutb(w_n807_0[1]),.din(w_dff_B_yEpiPgRN8_2));
	jspl jspl_w_n808_0(.douta(w_n808_0[0]),.doutb(w_n808_0[1]),.din(n808));
	jspl jspl_w_n809_0(.douta(w_n809_0[0]),.doutb(w_n809_0[1]),.din(w_dff_B_FgF8KqwX0_2));
	jspl jspl_w_n810_0(.douta(w_n810_0[0]),.doutb(w_n810_0[1]),.din(n810));
	jspl jspl_w_n811_0(.douta(w_n811_0[0]),.doutb(w_n811_0[1]),.din(w_dff_B_9rJcZFO74_2));
	jspl jspl_w_n812_0(.douta(w_n812_0[0]),.doutb(w_n812_0[1]),.din(n812));
	jspl jspl_w_n813_0(.douta(w_n813_0[0]),.doutb(w_n813_0[1]),.din(n813));
	jspl jspl_w_n814_0(.douta(w_n814_0[0]),.doutb(w_n814_0[1]),.din(n814));
	jspl jspl_w_n815_0(.douta(w_n815_0[0]),.doutb(w_n815_0[1]),.din(n815));
	jspl jspl_w_n816_0(.douta(w_n816_0[0]),.doutb(w_n816_0[1]),.din(n816));
	jspl jspl_w_n817_0(.douta(w_n817_0[0]),.doutb(w_n817_0[1]),.din(w_dff_B_c0w64E9o7_2));
	jspl jspl_w_n818_0(.douta(w_n818_0[0]),.doutb(w_n818_0[1]),.din(n818));
	jspl jspl_w_n819_0(.douta(w_n819_0[0]),.doutb(w_n819_0[1]),.din(w_dff_B_pf4x7cqt6_2));
	jspl jspl_w_n820_0(.douta(w_n820_0[0]),.doutb(w_n820_0[1]),.din(n820));
	jspl jspl_w_n821_0(.douta(w_n821_0[0]),.doutb(w_n821_0[1]),.din(w_dff_B_lsaBQh7J8_2));
	jspl jspl_w_n822_0(.douta(w_n822_0[0]),.doutb(w_n822_0[1]),.din(n822));
	jspl jspl_w_n823_0(.douta(w_dff_A_CZ2jEFdf6_0),.doutb(w_n823_0[1]),.din(n823));
	jspl jspl_w_n824_0(.douta(w_n824_0[0]),.doutb(w_n824_0[1]),.din(n824));
	jspl jspl_w_n826_0(.douta(w_n826_0[0]),.doutb(w_dff_A_ve3QpJuC3_1),.din(n826));
	jspl jspl_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.din(n827));
	jspl jspl_w_n829_0(.douta(w_dff_A_4Cy19Jzl6_0),.doutb(w_n829_0[1]),.din(n829));
	jspl jspl_w_n834_0(.douta(w_n834_0[0]),.doutb(w_n834_0[1]),.din(n834));
	jspl jspl_w_n835_0(.douta(w_n835_0[0]),.doutb(w_n835_0[1]),.din(w_dff_B_N6d7RHoj3_2));
	jspl jspl_w_n839_0(.douta(w_n839_0[0]),.doutb(w_n839_0[1]),.din(n839));
	jspl jspl_w_n840_0(.douta(w_dff_A_PXYu4tFF2_0),.doutb(w_n840_0[1]),.din(n840));
	jspl3 jspl3_w_n844_0(.douta(w_n844_0[0]),.doutb(w_n844_0[1]),.doutc(w_n844_0[2]),.din(n844));
	jspl jspl_w_n846_0(.douta(w_n846_0[0]),.doutb(w_n846_0[1]),.din(w_dff_B_X2kT5Udq3_2));
	jspl jspl_w_n849_0(.douta(w_n849_0[0]),.doutb(w_n849_0[1]),.din(n849));
	jspl jspl_w_n851_0(.douta(w_n851_0[0]),.doutb(w_n851_0[1]),.din(w_dff_B_E2Lm7Htj4_2));
	jspl jspl_w_n854_0(.douta(w_n854_0[0]),.doutb(w_n854_0[1]),.din(n854));
	jspl jspl_w_n856_0(.douta(w_n856_0[0]),.doutb(w_n856_0[1]),.din(w_dff_B_j1yGSPFY8_2));
	jspl jspl_w_n859_0(.douta(w_n859_0[0]),.doutb(w_n859_0[1]),.din(n859));
	jspl jspl_w_n861_0(.douta(w_n861_0[0]),.doutb(w_n861_0[1]),.din(w_dff_B_Bg6ghQej4_2));
	jspl jspl_w_n864_0(.douta(w_n864_0[0]),.doutb(w_n864_0[1]),.din(n864));
	jspl jspl_w_n866_0(.douta(w_n866_0[0]),.doutb(w_n866_0[1]),.din(w_dff_B_W4fjIvWG8_2));
	jspl jspl_w_n869_0(.douta(w_n869_0[0]),.doutb(w_n869_0[1]),.din(n869));
	jspl jspl_w_n871_0(.douta(w_n871_0[0]),.doutb(w_n871_0[1]),.din(w_dff_B_kYkqdPMr6_2));
	jspl jspl_w_n874_0(.douta(w_n874_0[0]),.doutb(w_n874_0[1]),.din(n874));
	jspl jspl_w_n876_0(.douta(w_n876_0[0]),.doutb(w_n876_0[1]),.din(w_dff_B_pfabGU1z4_2));
	jspl jspl_w_n879_0(.douta(w_n879_0[0]),.doutb(w_n879_0[1]),.din(n879));
	jspl jspl_w_n881_0(.douta(w_n881_0[0]),.doutb(w_n881_0[1]),.din(w_dff_B_JmAnH8nQ3_2));
	jspl jspl_w_n884_0(.douta(w_n884_0[0]),.doutb(w_n884_0[1]),.din(n884));
	jspl jspl_w_n886_0(.douta(w_n886_0[0]),.doutb(w_n886_0[1]),.din(w_dff_B_yAr04H9W1_2));
	jspl jspl_w_n889_0(.douta(w_n889_0[0]),.doutb(w_n889_0[1]),.din(n889));
	jspl jspl_w_n891_0(.douta(w_n891_0[0]),.doutb(w_n891_0[1]),.din(w_dff_B_PJROlhI89_2));
	jspl jspl_w_n895_0(.douta(w_n895_0[0]),.doutb(w_n895_0[1]),.din(n895));
	jspl jspl_w_n896_0(.douta(w_n896_0[0]),.doutb(w_dff_A_AhwbHvEf1_1),.din(n896));
	jspl jspl_w_n897_0(.douta(w_n897_0[0]),.doutb(w_n897_0[1]),.din(n897));
	jspl jspl_w_n898_0(.douta(w_n898_0[0]),.doutb(w_n898_0[1]),.din(w_dff_B_lLac3uo07_2));
	jspl jspl_w_n901_0(.douta(w_n901_0[0]),.doutb(w_n901_0[1]),.din(n901));
	jspl jspl_w_n903_0(.douta(w_dff_A_uLByc2El7_0),.doutb(w_n903_0[1]),.din(n903));
	jspl jspl_w_n906_0(.douta(w_n906_0[0]),.doutb(w_n906_0[1]),.din(n906));
	jspl jspl_w_n907_0(.douta(w_n907_0[0]),.doutb(w_n907_0[1]),.din(w_dff_B_sYNSHnuN6_2));
	jspl jspl_w_n908_0(.douta(w_n908_0[0]),.doutb(w_n908_0[1]),.din(n908));
	jspl jspl_w_n909_0(.douta(w_n909_0[0]),.doutb(w_n909_0[1]),.din(w_dff_B_QPpQGM361_2));
	jspl jspl_w_n910_0(.douta(w_n910_0[0]),.doutb(w_n910_0[1]),.din(n910));
	jspl jspl_w_n911_0(.douta(w_n911_0[0]),.doutb(w_n911_0[1]),.din(w_dff_B_Lcdxw4Xr7_2));
	jspl jspl_w_n912_0(.douta(w_n912_0[0]),.doutb(w_n912_0[1]),.din(n912));
	jspl jspl_w_n913_0(.douta(w_n913_0[0]),.doutb(w_n913_0[1]),.din(w_dff_B_n9EISm401_2));
	jspl jspl_w_n914_0(.douta(w_n914_0[0]),.doutb(w_n914_0[1]),.din(n914));
	jspl jspl_w_n915_0(.douta(w_n915_0[0]),.doutb(w_n915_0[1]),.din(w_dff_B_JcBbMAdb9_2));
	jspl jspl_w_n916_0(.douta(w_n916_0[0]),.doutb(w_n916_0[1]),.din(n916));
	jspl jspl_w_n917_0(.douta(w_n917_0[0]),.doutb(w_n917_0[1]),.din(w_dff_B_SqSzmfJI2_2));
	jspl jspl_w_n918_0(.douta(w_n918_0[0]),.doutb(w_n918_0[1]),.din(n918));
	jspl jspl_w_n919_0(.douta(w_n919_0[0]),.doutb(w_n919_0[1]),.din(n919));
	jspl jspl_w_n920_0(.douta(w_n920_0[0]),.doutb(w_n920_0[1]),.din(n920));
	jspl jspl_w_n921_0(.douta(w_n921_0[0]),.doutb(w_n921_0[1]),.din(n921));
	jspl jspl_w_n922_0(.douta(w_n922_0[0]),.doutb(w_n922_0[1]),.din(n922));
	jspl jspl_w_n923_0(.douta(w_n923_0[0]),.doutb(w_n923_0[1]),.din(w_dff_B_eZBfBava6_2));
	jspl jspl_w_n924_0(.douta(w_n924_0[0]),.doutb(w_n924_0[1]),.din(n924));
	jspl jspl_w_n925_0(.douta(w_n925_0[0]),.doutb(w_n925_0[1]),.din(w_dff_B_6Gtr6lbk5_2));
	jspl jspl_w_n926_0(.douta(w_n926_0[0]),.doutb(w_n926_0[1]),.din(n926));
	jspl3 jspl3_w_n927_0(.douta(w_n927_0[0]),.doutb(w_dff_A_rNhfqppf1_1),.doutc(w_dff_A_ERUtKZw50_2),.din(n927));
	jspl jspl_w_n929_0(.douta(w_n929_0[0]),.doutb(w_dff_A_hHU6UceV1_1),.din(n929));
	jspl jspl_w_n930_0(.douta(w_n930_0[0]),.doutb(w_n930_0[1]),.din(n930));
	jspl jspl_w_n931_0(.douta(w_n931_0[0]),.doutb(w_dff_A_nNe7f8Xx0_1),.din(n931));
	jspl jspl_w_n932_0(.douta(w_n932_0[0]),.doutb(w_n932_0[1]),.din(n932));
	jspl jspl_w_n937_0(.douta(w_n937_0[0]),.doutb(w_n937_0[1]),.din(n937));
	jspl jspl_w_n938_0(.douta(w_n938_0[0]),.doutb(w_n938_0[1]),.din(w_dff_B_OUTFygTT9_2));
	jspl3 jspl3_w_n942_0(.douta(w_n942_0[0]),.doutb(w_n942_0[1]),.doutc(w_n942_0[2]),.din(n942));
	jspl jspl_w_n943_0(.douta(w_n943_0[0]),.doutb(w_n943_0[1]),.din(w_dff_B_0RTT3rWU7_2));
	jspl jspl_w_n949_0(.douta(w_n949_0[0]),.doutb(w_n949_0[1]),.din(n949));
	jspl jspl_w_n951_0(.douta(w_n951_0[0]),.doutb(w_n951_0[1]),.din(w_dff_B_zFBisT5P4_2));
	jspl jspl_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.din(n954));
	jspl jspl_w_n956_0(.douta(w_n956_0[0]),.doutb(w_n956_0[1]),.din(w_dff_B_vZdHmVoe7_2));
	jspl jspl_w_n959_0(.douta(w_n959_0[0]),.doutb(w_n959_0[1]),.din(n959));
	jspl jspl_w_n961_0(.douta(w_n961_0[0]),.doutb(w_n961_0[1]),.din(w_dff_B_eSqY2FEm1_2));
	jspl jspl_w_n964_0(.douta(w_n964_0[0]),.doutb(w_n964_0[1]),.din(n964));
	jspl jspl_w_n966_0(.douta(w_n966_0[0]),.doutb(w_n966_0[1]),.din(w_dff_B_vTxBxvLn4_2));
	jspl jspl_w_n969_0(.douta(w_n969_0[0]),.doutb(w_n969_0[1]),.din(n969));
	jspl jspl_w_n971_0(.douta(w_n971_0[0]),.doutb(w_n971_0[1]),.din(w_dff_B_9B0pqAp15_2));
	jspl jspl_w_n974_0(.douta(w_n974_0[0]),.doutb(w_n974_0[1]),.din(n974));
	jspl jspl_w_n976_0(.douta(w_n976_0[0]),.doutb(w_n976_0[1]),.din(w_dff_B_jwFo8Crr7_2));
	jspl jspl_w_n979_0(.douta(w_n979_0[0]),.doutb(w_n979_0[1]),.din(n979));
	jspl jspl_w_n981_0(.douta(w_n981_0[0]),.doutb(w_n981_0[1]),.din(w_dff_B_AU6jyrFE3_2));
	jspl jspl_w_n984_0(.douta(w_n984_0[0]),.doutb(w_n984_0[1]),.din(n984));
	jspl jspl_w_n986_0(.douta(w_n986_0[0]),.doutb(w_n986_0[1]),.din(w_dff_B_A61RqbDr9_2));
	jspl jspl_w_n989_0(.douta(w_n989_0[0]),.doutb(w_n989_0[1]),.din(n989));
	jspl jspl_w_n991_0(.douta(w_n991_0[0]),.doutb(w_n991_0[1]),.din(w_dff_B_bflIGW7s7_2));
	jspl jspl_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.din(n994));
	jspl jspl_w_n996_0(.douta(w_n996_0[0]),.doutb(w_n996_0[1]),.din(w_dff_B_RN7mN8hd4_2));
	jspl jspl_w_n999_0(.douta(w_n999_0[0]),.doutb(w_n999_0[1]),.din(n999));
	jspl jspl_w_n1001_0(.douta(w_n1001_0[0]),.doutb(w_n1001_0[1]),.din(w_dff_B_rvbvWtr08_2));
	jspl jspl_w_n1005_0(.douta(w_n1005_0[0]),.doutb(w_n1005_0[1]),.din(n1005));
	jspl jspl_w_n1006_0(.douta(w_n1006_0[0]),.doutb(w_dff_A_DIA0lUDf8_1),.din(n1006));
	jspl jspl_w_n1008_0(.douta(w_dff_A_vaNofmMD7_0),.doutb(w_n1008_0[1]),.din(n1008));
	jspl jspl_w_n1009_0(.douta(w_n1009_0[0]),.doutb(w_n1009_0[1]),.din(n1009));
	jspl jspl_w_n1010_0(.douta(w_n1010_0[0]),.doutb(w_n1010_0[1]),.din(w_dff_B_rbubUt2i7_2));
	jspl jspl_w_n1011_0(.douta(w_n1011_0[0]),.doutb(w_n1011_0[1]),.din(n1011));
	jspl jspl_w_n1012_0(.douta(w_n1012_0[0]),.doutb(w_n1012_0[1]),.din(w_dff_B_QkUk3v3e1_2));
	jspl jspl_w_n1013_0(.douta(w_n1013_0[0]),.doutb(w_n1013_0[1]),.din(n1013));
	jspl jspl_w_n1014_0(.douta(w_n1014_0[0]),.doutb(w_n1014_0[1]),.din(w_dff_B_i5sM6kEZ8_2));
	jspl jspl_w_n1015_0(.douta(w_n1015_0[0]),.doutb(w_n1015_0[1]),.din(n1015));
	jspl jspl_w_n1016_0(.douta(w_n1016_0[0]),.doutb(w_n1016_0[1]),.din(w_dff_B_RcsfpYi26_2));
	jspl jspl_w_n1017_0(.douta(w_n1017_0[0]),.doutb(w_n1017_0[1]),.din(n1017));
	jspl jspl_w_n1018_0(.douta(w_n1018_0[0]),.doutb(w_n1018_0[1]),.din(w_dff_B_hOikBsCD4_2));
	jspl jspl_w_n1019_0(.douta(w_n1019_0[0]),.doutb(w_n1019_0[1]),.din(n1019));
	jspl jspl_w_n1020_0(.douta(w_n1020_0[0]),.doutb(w_n1020_0[1]),.din(w_dff_B_srM51NvW5_2));
	jspl jspl_w_n1021_0(.douta(w_n1021_0[0]),.doutb(w_n1021_0[1]),.din(n1021));
	jspl jspl_w_n1022_0(.douta(w_n1022_0[0]),.doutb(w_n1022_0[1]),.din(w_dff_B_odIEMLG73_2));
	jspl jspl_w_n1023_0(.douta(w_n1023_0[0]),.doutb(w_n1023_0[1]),.din(n1023));
	jspl jspl_w_n1024_0(.douta(w_n1024_0[0]),.doutb(w_n1024_0[1]),.din(n1024));
	jspl jspl_w_n1025_0(.douta(w_n1025_0[0]),.doutb(w_n1025_0[1]),.din(n1025));
	jspl jspl_w_n1026_0(.douta(w_n1026_0[0]),.doutb(w_n1026_0[1]),.din(n1026));
	jspl jspl_w_n1027_0(.douta(w_n1027_0[0]),.doutb(w_n1027_0[1]),.din(n1027));
	jspl jspl_w_n1028_0(.douta(w_n1028_0[0]),.doutb(w_n1028_0[1]),.din(w_dff_B_pV0mhRZL3_2));
	jspl jspl_w_n1029_0(.douta(w_n1029_0[0]),.doutb(w_n1029_0[1]),.din(n1029));
	jspl jspl_w_n1030_0(.douta(w_n1030_0[0]),.doutb(w_n1030_0[1]),.din(w_dff_B_lwCdysTz7_2));
	jspl jspl_w_n1031_0(.douta(w_n1031_0[0]),.doutb(w_n1031_0[1]),.din(n1031));
	jspl jspl_w_n1032_0(.douta(w_n1032_0[0]),.doutb(w_dff_A_LiLLaKQ70_1),.din(n1032));
	jspl jspl_w_n1033_0(.douta(w_n1033_0[0]),.doutb(w_n1033_0[1]),.din(n1033));
	jspl jspl_w_n1034_0(.douta(w_dff_A_8FZFsssn1_0),.doutb(w_n1034_0[1]),.din(n1034));
	jspl jspl_w_n1035_0(.douta(w_n1035_0[0]),.doutb(w_n1035_0[1]),.din(n1035));
	jspl jspl_w_n1037_0(.douta(w_n1037_0[0]),.doutb(w_n1037_0[1]),.din(w_dff_B_6NEy3HGz2_2));
	jspl jspl_w_n1039_0(.douta(w_n1039_0[0]),.doutb(w_dff_A_BLchi0CF4_1),.din(n1039));
	jspl jspl_w_n1043_0(.douta(w_n1043_0[0]),.doutb(w_n1043_0[1]),.din(n1043));
	jspl jspl_w_n1044_0(.douta(w_n1044_0[0]),.doutb(w_n1044_0[1]),.din(w_dff_B_A3hoYYku9_2));
	jspl jspl_w_n1048_0(.douta(w_dff_A_0WP8bNhx8_0),.doutb(w_n1048_0[1]),.din(n1048));
	jspl jspl_w_n1049_0(.douta(w_n1049_0[0]),.doutb(w_n1049_0[1]),.din(w_dff_B_LLAZKhDn3_2));
	jspl jspl_w_n1052_0(.douta(w_n1052_0[0]),.doutb(w_n1052_0[1]),.din(n1052));
	jspl jspl_w_n1054_0(.douta(w_n1054_0[0]),.doutb(w_n1054_0[1]),.din(w_dff_B_SzYlsXIl7_2));
	jspl jspl_w_n1057_0(.douta(w_n1057_0[0]),.doutb(w_n1057_0[1]),.din(n1057));
	jspl jspl_w_n1059_0(.douta(w_n1059_0[0]),.doutb(w_n1059_0[1]),.din(w_dff_B_4P83CbSp6_2));
	jspl jspl_w_n1062_0(.douta(w_n1062_0[0]),.doutb(w_n1062_0[1]),.din(n1062));
	jspl jspl_w_n1064_0(.douta(w_n1064_0[0]),.doutb(w_n1064_0[1]),.din(w_dff_B_PMFJBWlE4_2));
	jspl jspl_w_n1067_0(.douta(w_n1067_0[0]),.doutb(w_n1067_0[1]),.din(n1067));
	jspl jspl_w_n1069_0(.douta(w_n1069_0[0]),.doutb(w_n1069_0[1]),.din(w_dff_B_tE3GPyAT6_2));
	jspl jspl_w_n1072_0(.douta(w_n1072_0[0]),.doutb(w_n1072_0[1]),.din(n1072));
	jspl jspl_w_n1074_0(.douta(w_n1074_0[0]),.doutb(w_n1074_0[1]),.din(w_dff_B_0zxA06rf9_2));
	jspl jspl_w_n1077_0(.douta(w_n1077_0[0]),.doutb(w_n1077_0[1]),.din(n1077));
	jspl jspl_w_n1079_0(.douta(w_n1079_0[0]),.doutb(w_n1079_0[1]),.din(w_dff_B_zmFlblHR9_2));
	jspl jspl_w_n1082_0(.douta(w_n1082_0[0]),.doutb(w_n1082_0[1]),.din(n1082));
	jspl jspl_w_n1084_0(.douta(w_n1084_0[0]),.doutb(w_n1084_0[1]),.din(w_dff_B_F7lIEWSj0_2));
	jspl jspl_w_n1087_0(.douta(w_n1087_0[0]),.doutb(w_n1087_0[1]),.din(n1087));
	jspl jspl_w_n1089_0(.douta(w_n1089_0[0]),.doutb(w_n1089_0[1]),.din(w_dff_B_9eFiQyfl7_2));
	jspl jspl_w_n1092_0(.douta(w_n1092_0[0]),.doutb(w_n1092_0[1]),.din(n1092));
	jspl jspl_w_n1094_0(.douta(w_n1094_0[0]),.doutb(w_n1094_0[1]),.din(w_dff_B_9P0YEedD2_2));
	jspl jspl_w_n1097_0(.douta(w_n1097_0[0]),.doutb(w_n1097_0[1]),.din(n1097));
	jspl jspl_w_n1099_0(.douta(w_n1099_0[0]),.doutb(w_n1099_0[1]),.din(w_dff_B_9lWhhvuT2_2));
	jspl jspl_w_n1102_0(.douta(w_n1102_0[0]),.doutb(w_n1102_0[1]),.din(n1102));
	jspl jspl_w_n1103_0(.douta(w_n1103_0[0]),.doutb(w_n1103_0[1]),.din(w_dff_B_cqFfBWP55_2));
	jspl jspl_w_n1109_0(.douta(w_n1109_0[0]),.doutb(w_n1109_0[1]),.din(n1109));
	jspl jspl_w_n1110_0(.douta(w_dff_A_f2e2Ey2h5_0),.doutb(w_n1110_0[1]),.din(w_dff_B_GDoq4Fl55_2));
	jspl jspl_w_n1114_0(.douta(w_n1114_0[0]),.doutb(w_n1114_0[1]),.din(n1114));
	jspl jspl_w_n1115_0(.douta(w_n1115_0[0]),.doutb(w_n1115_0[1]),.din(n1115));
	jspl jspl_w_n1116_0(.douta(w_n1116_0[0]),.doutb(w_n1116_0[1]),.din(n1116));
	jspl jspl_w_n1117_0(.douta(w_n1117_0[0]),.doutb(w_n1117_0[1]),.din(w_dff_B_GbnFbinF7_2));
	jspl jspl_w_n1118_0(.douta(w_n1118_0[0]),.doutb(w_n1118_0[1]),.din(n1118));
	jspl jspl_w_n1119_0(.douta(w_n1119_0[0]),.doutb(w_n1119_0[1]),.din(w_dff_B_hZ2lehh50_2));
	jspl jspl_w_n1120_0(.douta(w_n1120_0[0]),.doutb(w_n1120_0[1]),.din(n1120));
	jspl jspl_w_n1121_0(.douta(w_n1121_0[0]),.doutb(w_n1121_0[1]),.din(w_dff_B_HKVoNoEe3_2));
	jspl jspl_w_n1122_0(.douta(w_n1122_0[0]),.doutb(w_n1122_0[1]),.din(n1122));
	jspl jspl_w_n1123_0(.douta(w_n1123_0[0]),.doutb(w_n1123_0[1]),.din(w_dff_B_ArKrp9Jo9_2));
	jspl jspl_w_n1124_0(.douta(w_n1124_0[0]),.doutb(w_n1124_0[1]),.din(n1124));
	jspl jspl_w_n1125_0(.douta(w_n1125_0[0]),.doutb(w_n1125_0[1]),.din(w_dff_B_xeE0Cf714_2));
	jspl jspl_w_n1126_0(.douta(w_n1126_0[0]),.doutb(w_n1126_0[1]),.din(n1126));
	jspl jspl_w_n1127_0(.douta(w_n1127_0[0]),.doutb(w_n1127_0[1]),.din(w_dff_B_Ey1mCoSe0_2));
	jspl jspl_w_n1128_0(.douta(w_n1128_0[0]),.doutb(w_n1128_0[1]),.din(n1128));
	jspl jspl_w_n1129_0(.douta(w_n1129_0[0]),.doutb(w_n1129_0[1]),.din(n1129));
	jspl jspl_w_n1130_0(.douta(w_n1130_0[0]),.doutb(w_n1130_0[1]),.din(n1130));
	jspl jspl_w_n1131_0(.douta(w_n1131_0[0]),.doutb(w_n1131_0[1]),.din(n1131));
	jspl jspl_w_n1132_0(.douta(w_n1132_0[0]),.doutb(w_n1132_0[1]),.din(n1132));
	jspl jspl_w_n1133_0(.douta(w_n1133_0[0]),.doutb(w_n1133_0[1]),.din(w_dff_B_dQDJWevx9_2));
	jspl jspl_w_n1134_0(.douta(w_n1134_0[0]),.doutb(w_n1134_0[1]),.din(n1134));
	jspl jspl_w_n1135_0(.douta(w_n1135_0[0]),.doutb(w_n1135_0[1]),.din(w_dff_B_4OqqlQj08_2));
	jspl jspl_w_n1137_0(.douta(w_n1137_0[0]),.doutb(w_n1137_0[1]),.din(n1137));
	jspl jspl_w_n1138_0(.douta(w_n1138_0[0]),.doutb(w_n1138_0[1]),.din(n1138));
	jspl jspl_w_n1139_0(.douta(w_n1139_0[0]),.doutb(w_n1139_0[1]),.din(n1139));
	jspl jspl_w_n1140_0(.douta(w_n1140_0[0]),.doutb(w_dff_A_HyISg1en7_1),.din(n1140));
	jspl jspl_w_n1141_0(.douta(w_n1141_0[0]),.doutb(w_n1141_0[1]),.din(n1141));
	jspl jspl_w_n1147_0(.douta(w_n1147_0[0]),.doutb(w_n1147_0[1]),.din(n1147));
	jspl jspl_w_n1151_0(.douta(w_dff_A_58oNjSm74_0),.doutb(w_n1151_0[1]),.din(w_dff_B_Xfkd7YaU7_2));
	jspl jspl_w_n1152_0(.douta(w_n1152_0[0]),.doutb(w_n1152_0[1]),.din(w_dff_B_la2T5edW5_2));
	jspl jspl_w_n1156_0(.douta(w_n1156_0[0]),.doutb(w_n1156_0[1]),.din(n1156));
	jspl jspl_w_n1158_0(.douta(w_n1158_0[0]),.doutb(w_n1158_0[1]),.din(w_dff_B_Iuv5wbIc7_2));
	jspl jspl_w_n1161_0(.douta(w_n1161_0[0]),.doutb(w_n1161_0[1]),.din(n1161));
	jspl jspl_w_n1163_0(.douta(w_n1163_0[0]),.doutb(w_n1163_0[1]),.din(w_dff_B_WFUfie7T9_2));
	jspl jspl_w_n1166_0(.douta(w_n1166_0[0]),.doutb(w_n1166_0[1]),.din(n1166));
	jspl jspl_w_n1168_0(.douta(w_n1168_0[0]),.doutb(w_n1168_0[1]),.din(w_dff_B_22AifnwD9_2));
	jspl jspl_w_n1171_0(.douta(w_n1171_0[0]),.doutb(w_n1171_0[1]),.din(n1171));
	jspl jspl_w_n1173_0(.douta(w_n1173_0[0]),.doutb(w_n1173_0[1]),.din(w_dff_B_iArFbLF42_2));
	jspl jspl_w_n1176_0(.douta(w_n1176_0[0]),.doutb(w_n1176_0[1]),.din(n1176));
	jspl jspl_w_n1178_0(.douta(w_n1178_0[0]),.doutb(w_n1178_0[1]),.din(w_dff_B_WTHNYiGv2_2));
	jspl jspl_w_n1181_0(.douta(w_n1181_0[0]),.doutb(w_n1181_0[1]),.din(n1181));
	jspl jspl_w_n1183_0(.douta(w_n1183_0[0]),.doutb(w_n1183_0[1]),.din(w_dff_B_44hlovNk6_2));
	jspl jspl_w_n1186_0(.douta(w_n1186_0[0]),.doutb(w_n1186_0[1]),.din(n1186));
	jspl jspl_w_n1188_0(.douta(w_n1188_0[0]),.doutb(w_n1188_0[1]),.din(w_dff_B_vuesWQg10_2));
	jspl jspl_w_n1191_0(.douta(w_n1191_0[0]),.doutb(w_n1191_0[1]),.din(n1191));
	jspl jspl_w_n1193_0(.douta(w_n1193_0[0]),.doutb(w_n1193_0[1]),.din(w_dff_B_eXoYxCfj8_2));
	jspl jspl_w_n1196_0(.douta(w_n1196_0[0]),.doutb(w_n1196_0[1]),.din(n1196));
	jspl jspl_w_n1198_0(.douta(w_n1198_0[0]),.doutb(w_n1198_0[1]),.din(w_dff_B_Xiu0xkK29_2));
	jspl jspl_w_n1201_0(.douta(w_n1201_0[0]),.doutb(w_n1201_0[1]),.din(n1201));
	jspl jspl_w_n1203_0(.douta(w_n1203_0[0]),.doutb(w_n1203_0[1]),.din(w_dff_B_B9IrkPD37_2));
	jspl jspl_w_n1206_0(.douta(w_n1206_0[0]),.doutb(w_n1206_0[1]),.din(w_dff_B_ZnJx9fZ55_2));
	jspl jspl_w_n1207_0(.douta(w_n1207_0[0]),.doutb(w_n1207_0[1]),.din(w_dff_B_y5rNK1No5_2));
	jspl jspl_w_n1208_0(.douta(w_n1208_0[0]),.doutb(w_n1208_0[1]),.din(w_dff_B_RqiMIXOz0_2));
	jspl jspl_w_n1210_0(.douta(w_n1210_0[0]),.doutb(w_n1210_0[1]),.din(n1210));
	jspl jspl_w_n1212_0(.douta(w_n1212_0[0]),.doutb(w_n1212_0[1]),.din(n1212));
	jspl jspl_w_n1213_0(.douta(w_n1213_0[0]),.doutb(w_n1213_0[1]),.din(n1213));
	jspl jspl_w_n1214_0(.douta(w_n1214_0[0]),.doutb(w_n1214_0[1]),.din(n1214));
	jspl jspl_w_n1215_0(.douta(w_n1215_0[0]),.doutb(w_n1215_0[1]),.din(w_dff_B_msSltTL19_2));
	jspl jspl_w_n1216_0(.douta(w_n1216_0[0]),.doutb(w_n1216_0[1]),.din(n1216));
	jspl jspl_w_n1217_0(.douta(w_n1217_0[0]),.doutb(w_n1217_0[1]),.din(w_dff_B_cMtgVFzy1_2));
	jspl jspl_w_n1218_0(.douta(w_n1218_0[0]),.doutb(w_n1218_0[1]),.din(n1218));
	jspl jspl_w_n1219_0(.douta(w_n1219_0[0]),.doutb(w_n1219_0[1]),.din(w_dff_B_0ln7i3yv3_2));
	jspl jspl_w_n1220_0(.douta(w_n1220_0[0]),.doutb(w_n1220_0[1]),.din(n1220));
	jspl jspl_w_n1221_0(.douta(w_n1221_0[0]),.doutb(w_n1221_0[1]),.din(w_dff_B_MsvinaVe8_2));
	jspl jspl_w_n1222_0(.douta(w_n1222_0[0]),.doutb(w_n1222_0[1]),.din(n1222));
	jspl jspl_w_n1223_0(.douta(w_n1223_0[0]),.doutb(w_n1223_0[1]),.din(w_dff_B_lnYCOwVq2_2));
	jspl jspl_w_n1224_0(.douta(w_n1224_0[0]),.doutb(w_n1224_0[1]),.din(n1224));
	jspl jspl_w_n1225_0(.douta(w_n1225_0[0]),.doutb(w_n1225_0[1]),.din(w_dff_B_X8PXlsSu2_2));
	jspl jspl_w_n1226_0(.douta(w_n1226_0[0]),.doutb(w_n1226_0[1]),.din(n1226));
	jspl jspl_w_n1227_0(.douta(w_n1227_0[0]),.doutb(w_n1227_0[1]),.din(n1227));
	jspl jspl_w_n1228_0(.douta(w_n1228_0[0]),.doutb(w_n1228_0[1]),.din(n1228));
	jspl jspl_w_n1229_0(.douta(w_n1229_0[0]),.doutb(w_n1229_0[1]),.din(n1229));
	jspl jspl_w_n1230_0(.douta(w_n1230_0[0]),.doutb(w_n1230_0[1]),.din(n1230));
	jspl jspl_w_n1231_0(.douta(w_n1231_0[0]),.doutb(w_n1231_0[1]),.din(w_dff_B_O1NHPjoB7_2));
	jspl jspl_w_n1232_0(.douta(w_n1232_0[0]),.doutb(w_n1232_0[1]),.din(n1232));
	jspl jspl_w_n1234_0(.douta(w_n1234_0[0]),.doutb(w_n1234_0[1]),.din(w_dff_B_GIJup5jm6_2));
	jspl jspl_w_n1236_0(.douta(w_n1236_0[0]),.doutb(w_n1236_0[1]),.din(n1236));
	jspl jspl_w_n1237_0(.douta(w_n1237_0[0]),.doutb(w_n1237_0[1]),.din(n1237));
	jspl jspl_w_n1238_0(.douta(w_dff_A_8LRjp0fZ3_0),.doutb(w_n1238_0[1]),.din(n1238));
	jspl jspl_w_n1244_0(.douta(w_n1244_0[0]),.doutb(w_n1244_0[1]),.din(n1244));
	jspl jspl_w_n1247_0(.douta(w_n1247_0[0]),.doutb(w_n1247_0[1]),.din(n1247));
	jspl jspl_w_n1248_0(.douta(w_n1248_0[0]),.doutb(w_n1248_0[1]),.din(w_dff_B_aULq1Jt46_2));
	jspl jspl_w_n1251_0(.douta(w_n1251_0[0]),.doutb(w_n1251_0[1]),.din(n1251));
	jspl jspl_w_n1253_0(.douta(w_n1253_0[0]),.doutb(w_n1253_0[1]),.din(w_dff_B_zS3qZF2g9_2));
	jspl jspl_w_n1256_0(.douta(w_n1256_0[0]),.doutb(w_n1256_0[1]),.din(n1256));
	jspl jspl_w_n1258_0(.douta(w_n1258_0[0]),.doutb(w_n1258_0[1]),.din(w_dff_B_qyzV3BIc3_2));
	jspl jspl_w_n1261_0(.douta(w_n1261_0[0]),.doutb(w_n1261_0[1]),.din(n1261));
	jspl jspl_w_n1263_0(.douta(w_n1263_0[0]),.doutb(w_n1263_0[1]),.din(w_dff_B_wK63IE4k2_2));
	jspl jspl_w_n1266_0(.douta(w_n1266_0[0]),.doutb(w_n1266_0[1]),.din(n1266));
	jspl jspl_w_n1268_0(.douta(w_n1268_0[0]),.doutb(w_n1268_0[1]),.din(w_dff_B_7R0lN1O60_2));
	jspl jspl_w_n1271_0(.douta(w_n1271_0[0]),.doutb(w_n1271_0[1]),.din(n1271));
	jspl jspl_w_n1273_0(.douta(w_n1273_0[0]),.doutb(w_n1273_0[1]),.din(w_dff_B_7zpv10YT7_2));
	jspl jspl_w_n1276_0(.douta(w_n1276_0[0]),.doutb(w_n1276_0[1]),.din(n1276));
	jspl jspl_w_n1278_0(.douta(w_n1278_0[0]),.doutb(w_n1278_0[1]),.din(w_dff_B_1Klk0tMV1_2));
	jspl jspl_w_n1281_0(.douta(w_n1281_0[0]),.doutb(w_n1281_0[1]),.din(n1281));
	jspl jspl_w_n1283_0(.douta(w_n1283_0[0]),.doutb(w_n1283_0[1]),.din(w_dff_B_bpkdk6rt2_2));
	jspl jspl_w_n1286_0(.douta(w_n1286_0[0]),.doutb(w_n1286_0[1]),.din(n1286));
	jspl jspl_w_n1288_0(.douta(w_n1288_0[0]),.doutb(w_n1288_0[1]),.din(w_dff_B_3XfacPBE0_2));
	jspl jspl_w_n1291_0(.douta(w_n1291_0[0]),.doutb(w_n1291_0[1]),.din(n1291));
	jspl jspl_w_n1293_0(.douta(w_n1293_0[0]),.doutb(w_n1293_0[1]),.din(w_dff_B_EGF4byLT4_2));
	jspl jspl_w_n1296_0(.douta(w_n1296_0[0]),.doutb(w_n1296_0[1]),.din(w_dff_B_MWaXlhv09_2));
	jspl jspl_w_n1297_0(.douta(w_n1297_0[0]),.doutb(w_n1297_0[1]),.din(w_dff_B_HNwucoHX8_2));
	jspl jspl_w_n1298_0(.douta(w_n1298_0[0]),.doutb(w_n1298_0[1]),.din(w_dff_B_7a6jpQSa0_2));
	jspl jspl_w_n1301_0(.douta(w_n1301_0[0]),.doutb(w_n1301_0[1]),.din(n1301));
	jspl jspl_w_n1303_0(.douta(w_n1303_0[0]),.doutb(w_n1303_0[1]),.din(n1303));
	jspl jspl_w_n1304_0(.douta(w_n1304_0[0]),.doutb(w_n1304_0[1]),.din(n1304));
	jspl jspl_w_n1305_0(.douta(w_n1305_0[0]),.doutb(w_n1305_0[1]),.din(n1305));
	jspl jspl_w_n1306_0(.douta(w_n1306_0[0]),.doutb(w_n1306_0[1]),.din(n1306));
	jspl jspl_w_n1307_0(.douta(w_n1307_0[0]),.doutb(w_n1307_0[1]),.din(n1307));
	jspl jspl_w_n1308_0(.douta(w_n1308_0[0]),.doutb(w_n1308_0[1]),.din(w_dff_B_JJRZtfhZ9_2));
	jspl jspl_w_n1309_0(.douta(w_n1309_0[0]),.doutb(w_n1309_0[1]),.din(n1309));
	jspl jspl_w_n1310_0(.douta(w_n1310_0[0]),.doutb(w_n1310_0[1]),.din(w_dff_B_OyczPD237_2));
	jspl jspl_w_n1311_0(.douta(w_n1311_0[0]),.doutb(w_n1311_0[1]),.din(n1311));
	jspl jspl_w_n1312_0(.douta(w_n1312_0[0]),.doutb(w_n1312_0[1]),.din(w_dff_B_mADqmqP18_2));
	jspl jspl_w_n1313_0(.douta(w_n1313_0[0]),.doutb(w_n1313_0[1]),.din(n1313));
	jspl jspl_w_n1314_0(.douta(w_n1314_0[0]),.doutb(w_n1314_0[1]),.din(w_dff_B_gBIJsM8w9_2));
	jspl jspl_w_n1315_0(.douta(w_n1315_0[0]),.doutb(w_n1315_0[1]),.din(n1315));
	jspl jspl_w_n1316_0(.douta(w_n1316_0[0]),.doutb(w_n1316_0[1]),.din(w_dff_B_cN1DcKVD7_2));
	jspl jspl_w_n1317_0(.douta(w_n1317_0[0]),.doutb(w_n1317_0[1]),.din(n1317));
	jspl jspl_w_n1318_0(.douta(w_n1318_0[0]),.doutb(w_n1318_0[1]),.din(n1318));
	jspl jspl_w_n1319_0(.douta(w_n1319_0[0]),.doutb(w_n1319_0[1]),.din(n1319));
	jspl jspl_w_n1320_0(.douta(w_n1320_0[0]),.doutb(w_n1320_0[1]),.din(n1320));
	jspl jspl_w_n1321_0(.douta(w_n1321_0[0]),.doutb(w_n1321_0[1]),.din(n1321));
	jspl jspl_w_n1322_0(.douta(w_n1322_0[0]),.doutb(w_dff_A_LfO3RIHK7_1),.din(n1322));
	jspl jspl_w_n1324_0(.douta(w_n1324_0[0]),.doutb(w_n1324_0[1]),.din(n1324));
	jspl jspl_w_n1325_0(.douta(w_n1325_0[0]),.doutb(w_dff_A_nsNq7sN28_1),.din(n1325));
	jspl jspl_w_n1326_0(.douta(w_dff_A_K4ToNhLz9_0),.doutb(w_n1326_0[1]),.din(n1326));
	jspl jspl_w_n1332_0(.douta(w_n1332_0[0]),.doutb(w_n1332_0[1]),.din(n1332));
	jspl jspl_w_n1337_0(.douta(w_n1337_0[0]),.doutb(w_n1337_0[1]),.din(n1337));
	jspl jspl_w_n1338_0(.douta(w_n1338_0[0]),.doutb(w_n1338_0[1]),.din(w_dff_B_mJ9wVZH48_2));
	jspl jspl_w_n1341_0(.douta(w_n1341_0[0]),.doutb(w_n1341_0[1]),.din(n1341));
	jspl jspl_w_n1343_0(.douta(w_n1343_0[0]),.doutb(w_n1343_0[1]),.din(w_dff_B_Cg2CwX5J4_2));
	jspl jspl_w_n1346_0(.douta(w_n1346_0[0]),.doutb(w_n1346_0[1]),.din(n1346));
	jspl jspl_w_n1348_0(.douta(w_n1348_0[0]),.doutb(w_n1348_0[1]),.din(w_dff_B_6NUDczgV1_2));
	jspl jspl_w_n1351_0(.douta(w_n1351_0[0]),.doutb(w_n1351_0[1]),.din(n1351));
	jspl jspl_w_n1353_0(.douta(w_n1353_0[0]),.doutb(w_n1353_0[1]),.din(w_dff_B_aVwQOu5d0_2));
	jspl jspl_w_n1356_0(.douta(w_n1356_0[0]),.doutb(w_n1356_0[1]),.din(n1356));
	jspl jspl_w_n1358_0(.douta(w_n1358_0[0]),.doutb(w_n1358_0[1]),.din(w_dff_B_ytPP6zC89_2));
	jspl jspl_w_n1361_0(.douta(w_n1361_0[0]),.doutb(w_n1361_0[1]),.din(n1361));
	jspl jspl_w_n1363_0(.douta(w_n1363_0[0]),.doutb(w_n1363_0[1]),.din(w_dff_B_iqpIQTzU2_2));
	jspl jspl_w_n1366_0(.douta(w_n1366_0[0]),.doutb(w_n1366_0[1]),.din(n1366));
	jspl jspl_w_n1368_0(.douta(w_n1368_0[0]),.doutb(w_n1368_0[1]),.din(w_dff_B_kHJAgOSm2_2));
	jspl jspl_w_n1371_0(.douta(w_n1371_0[0]),.doutb(w_n1371_0[1]),.din(n1371));
	jspl jspl_w_n1373_0(.douta(w_n1373_0[0]),.doutb(w_n1373_0[1]),.din(w_dff_B_7bdxXkSP7_2));
	jspl jspl_w_n1376_0(.douta(w_n1376_0[0]),.doutb(w_n1376_0[1]),.din(w_dff_B_c1BRs3pm3_2));
	jspl jspl_w_n1378_0(.douta(w_n1378_0[0]),.doutb(w_n1378_0[1]),.din(w_dff_B_XOoBHcnR4_2));
	jspl jspl_w_n1381_0(.douta(w_n1381_0[0]),.doutb(w_n1381_0[1]),.din(w_dff_B_fYYk5f3O9_2));
	jspl jspl_w_n1382_0(.douta(w_n1382_0[0]),.doutb(w_n1382_0[1]),.din(w_dff_B_IEOErc0A7_2));
	jspl jspl_w_n1383_0(.douta(w_n1383_0[0]),.doutb(w_n1383_0[1]),.din(w_dff_B_2TsNxkrJ7_2));
	jspl jspl_w_n1386_0(.douta(w_n1386_0[0]),.doutb(w_n1386_0[1]),.din(n1386));
	jspl jspl_w_n1388_0(.douta(w_n1388_0[0]),.doutb(w_n1388_0[1]),.din(n1388));
	jspl jspl_w_n1389_0(.douta(w_n1389_0[0]),.doutb(w_n1389_0[1]),.din(n1389));
	jspl jspl_w_n1390_0(.douta(w_n1390_0[0]),.doutb(w_n1390_0[1]),.din(n1390));
	jspl jspl_w_n1391_0(.douta(w_n1391_0[0]),.doutb(w_n1391_0[1]),.din(n1391));
	jspl jspl_w_n1392_0(.douta(w_n1392_0[0]),.doutb(w_n1392_0[1]),.din(n1392));
	jspl jspl_w_n1393_0(.douta(w_n1393_0[0]),.doutb(w_n1393_0[1]),.din(n1393));
	jspl jspl_w_n1394_0(.douta(w_n1394_0[0]),.doutb(w_n1394_0[1]),.din(n1394));
	jspl jspl_w_n1395_0(.douta(w_n1395_0[0]),.doutb(w_n1395_0[1]),.din(w_dff_B_2gb9Bxer1_2));
	jspl jspl_w_n1396_0(.douta(w_n1396_0[0]),.doutb(w_n1396_0[1]),.din(n1396));
	jspl jspl_w_n1397_0(.douta(w_n1397_0[0]),.doutb(w_n1397_0[1]),.din(w_dff_B_1JzL5Mq57_2));
	jspl jspl_w_n1398_0(.douta(w_n1398_0[0]),.doutb(w_n1398_0[1]),.din(n1398));
	jspl jspl_w_n1399_0(.douta(w_n1399_0[0]),.doutb(w_n1399_0[1]),.din(w_dff_B_1ibA4IKY8_2));
	jspl jspl_w_n1400_0(.douta(w_n1400_0[0]),.doutb(w_n1400_0[1]),.din(n1400));
	jspl jspl_w_n1401_0(.douta(w_n1401_0[0]),.doutb(w_n1401_0[1]),.din(w_dff_B_9ek3H3DE0_2));
	jspl jspl_w_n1402_0(.douta(w_n1402_0[0]),.doutb(w_n1402_0[1]),.din(n1402));
	jspl jspl_w_n1403_0(.douta(w_n1403_0[0]),.doutb(w_n1403_0[1]),.din(n1403));
	jspl jspl_w_n1404_0(.douta(w_n1404_0[0]),.doutb(w_n1404_0[1]),.din(n1404));
	jspl jspl_w_n1405_0(.douta(w_n1405_0[0]),.doutb(w_n1405_0[1]),.din(n1405));
	jspl jspl_w_n1407_0(.douta(w_n1407_0[0]),.doutb(w_n1407_0[1]),.din(n1407));
	jspl jspl_w_n1409_0(.douta(w_n1409_0[0]),.doutb(w_n1409_0[1]),.din(n1409));
	jspl jspl_w_n1410_0(.douta(w_n1410_0[0]),.doutb(w_dff_A_VznJHwpx9_1),.din(n1410));
	jspl jspl_w_n1415_0(.douta(w_n1415_0[0]),.doutb(w_n1415_0[1]),.din(n1415));
	jspl jspl_w_n1420_0(.douta(w_n1420_0[0]),.doutb(w_n1420_0[1]),.din(w_dff_B_5P4pp9zh5_2));
	jspl jspl_w_n1421_0(.douta(w_n1421_0[0]),.doutb(w_n1421_0[1]),.din(w_dff_B_wthlQ4w61_2));
	jspl jspl_w_n1424_0(.douta(w_n1424_0[0]),.doutb(w_n1424_0[1]),.din(n1424));
	jspl jspl_w_n1426_0(.douta(w_n1426_0[0]),.doutb(w_n1426_0[1]),.din(w_dff_B_hnjWvXPB6_2));
	jspl jspl_w_n1429_0(.douta(w_n1429_0[0]),.doutb(w_n1429_0[1]),.din(n1429));
	jspl jspl_w_n1431_0(.douta(w_n1431_0[0]),.doutb(w_n1431_0[1]),.din(w_dff_B_Gzmv50DE8_2));
	jspl jspl_w_n1434_0(.douta(w_n1434_0[0]),.doutb(w_n1434_0[1]),.din(n1434));
	jspl jspl_w_n1436_0(.douta(w_n1436_0[0]),.doutb(w_n1436_0[1]),.din(w_dff_B_2ywxSxKj8_2));
	jspl jspl_w_n1439_0(.douta(w_n1439_0[0]),.doutb(w_n1439_0[1]),.din(n1439));
	jspl jspl_w_n1441_0(.douta(w_n1441_0[0]),.doutb(w_n1441_0[1]),.din(w_dff_B_NIiP5MnK3_2));
	jspl jspl_w_n1444_0(.douta(w_n1444_0[0]),.doutb(w_n1444_0[1]),.din(n1444));
	jspl jspl_w_n1446_0(.douta(w_n1446_0[0]),.doutb(w_n1446_0[1]),.din(w_dff_B_jjedWkFG1_2));
	jspl jspl_w_n1449_0(.douta(w_n1449_0[0]),.doutb(w_n1449_0[1]),.din(w_dff_B_njPQvG9e8_2));
	jspl jspl_w_n1451_0(.douta(w_n1451_0[0]),.doutb(w_n1451_0[1]),.din(w_dff_B_hT9Ev7Vt9_2));
	jspl jspl_w_n1454_0(.douta(w_n1454_0[0]),.doutb(w_n1454_0[1]),.din(w_dff_B_qdYNCKvA2_2));
	jspl jspl_w_n1456_0(.douta(w_n1456_0[0]),.doutb(w_n1456_0[1]),.din(w_dff_B_FDLZUWT77_2));
	jspl jspl_w_n1459_0(.douta(w_n1459_0[0]),.doutb(w_n1459_0[1]),.din(w_dff_B_jUVca4ae9_2));
	jspl jspl_w_n1460_0(.douta(w_n1460_0[0]),.doutb(w_n1460_0[1]),.din(w_dff_B_9HjdEJhl7_2));
	jspl jspl_w_n1461_0(.douta(w_n1461_0[0]),.doutb(w_n1461_0[1]),.din(w_dff_B_qLO6wcXk4_2));
	jspl jspl_w_n1464_0(.douta(w_n1464_0[0]),.doutb(w_n1464_0[1]),.din(n1464));
	jspl jspl_w_n1466_0(.douta(w_n1466_0[0]),.doutb(w_n1466_0[1]),.din(n1466));
	jspl jspl_w_n1467_0(.douta(w_n1467_0[0]),.doutb(w_n1467_0[1]),.din(n1467));
	jspl jspl_w_n1468_0(.douta(w_n1468_0[0]),.doutb(w_n1468_0[1]),.din(n1468));
	jspl jspl_w_n1469_0(.douta(w_n1469_0[0]),.doutb(w_n1469_0[1]),.din(n1469));
	jspl jspl_w_n1470_0(.douta(w_n1470_0[0]),.doutb(w_n1470_0[1]),.din(n1470));
	jspl jspl_w_n1471_0(.douta(w_n1471_0[0]),.doutb(w_n1471_0[1]),.din(n1471));
	jspl jspl_w_n1472_0(.douta(w_n1472_0[0]),.doutb(w_n1472_0[1]),.din(n1472));
	jspl jspl_w_n1473_0(.douta(w_n1473_0[0]),.doutb(w_n1473_0[1]),.din(n1473));
	jspl jspl_w_n1474_0(.douta(w_n1474_0[0]),.doutb(w_n1474_0[1]),.din(n1474));
	jspl jspl_w_n1475_0(.douta(w_n1475_0[0]),.doutb(w_n1475_0[1]),.din(w_dff_B_HISQ8N1N8_2));
	jspl jspl_w_n1476_0(.douta(w_n1476_0[0]),.doutb(w_n1476_0[1]),.din(n1476));
	jspl jspl_w_n1477_0(.douta(w_n1477_0[0]),.doutb(w_n1477_0[1]),.din(w_dff_B_A3R2VAa63_2));
	jspl jspl_w_n1478_0(.douta(w_n1478_0[0]),.doutb(w_n1478_0[1]),.din(n1478));
	jspl jspl_w_n1479_0(.douta(w_n1479_0[0]),.doutb(w_n1479_0[1]),.din(w_dff_B_yDwue3896_2));
	jspl jspl_w_n1480_0(.douta(w_n1480_0[0]),.doutb(w_n1480_0[1]),.din(n1480));
	jspl jspl_w_n1481_0(.douta(w_n1481_0[0]),.doutb(w_n1481_0[1]),.din(n1481));
	jspl jspl_w_n1483_0(.douta(w_n1483_0[0]),.doutb(w_n1483_0[1]),.din(n1483));
	jspl jspl_w_n1485_0(.douta(w_n1485_0[0]),.doutb(w_n1485_0[1]),.din(n1485));
	jspl jspl_w_n1486_0(.douta(w_n1486_0[0]),.doutb(w_dff_A_aEBeq1PX8_1),.din(n1486));
	jspl jspl_w_n1491_0(.douta(w_n1491_0[0]),.doutb(w_n1491_0[1]),.din(n1491));
	jspl jspl_w_n1496_0(.douta(w_n1496_0[0]),.doutb(w_n1496_0[1]),.din(w_dff_B_1PbYWcAW4_2));
	jspl jspl_w_n1497_0(.douta(w_n1497_0[0]),.doutb(w_n1497_0[1]),.din(w_dff_B_ePm4FQ1L1_2));
	jspl jspl_w_n1500_0(.douta(w_n1500_0[0]),.doutb(w_n1500_0[1]),.din(n1500));
	jspl jspl_w_n1502_0(.douta(w_n1502_0[0]),.doutb(w_n1502_0[1]),.din(w_dff_B_2Dc2Cqqv3_2));
	jspl jspl_w_n1505_0(.douta(w_n1505_0[0]),.doutb(w_n1505_0[1]),.din(n1505));
	jspl jspl_w_n1507_0(.douta(w_n1507_0[0]),.doutb(w_n1507_0[1]),.din(w_dff_B_m0eMMI8i3_2));
	jspl jspl_w_n1510_0(.douta(w_n1510_0[0]),.doutb(w_n1510_0[1]),.din(n1510));
	jspl jspl_w_n1512_0(.douta(w_n1512_0[0]),.doutb(w_n1512_0[1]),.din(w_dff_B_2q0oM0jv1_2));
	jspl jspl_w_n1515_0(.douta(w_n1515_0[0]),.doutb(w_n1515_0[1]),.din(w_dff_B_f4y5ryhm3_2));
	jspl jspl_w_n1517_0(.douta(w_n1517_0[0]),.doutb(w_n1517_0[1]),.din(w_dff_B_68ngA5Vo5_2));
	jspl jspl_w_n1520_0(.douta(w_n1520_0[0]),.doutb(w_n1520_0[1]),.din(w_dff_B_OMES7jqo9_2));
	jspl jspl_w_n1522_0(.douta(w_n1522_0[0]),.doutb(w_n1522_0[1]),.din(w_dff_B_sEVUrz8g0_2));
	jspl jspl_w_n1525_0(.douta(w_n1525_0[0]),.doutb(w_n1525_0[1]),.din(w_dff_B_4P5mUltv6_2));
	jspl jspl_w_n1527_0(.douta(w_n1527_0[0]),.doutb(w_n1527_0[1]),.din(w_dff_B_ugBGSNfa3_2));
	jspl jspl_w_n1530_0(.douta(w_n1530_0[0]),.doutb(w_n1530_0[1]),.din(w_dff_B_jyCedYn23_2));
	jspl jspl_w_n1531_0(.douta(w_n1531_0[0]),.doutb(w_n1531_0[1]),.din(w_dff_B_8YzArT0w9_2));
	jspl jspl_w_n1532_0(.douta(w_n1532_0[0]),.doutb(w_n1532_0[1]),.din(w_dff_B_7nodYucn0_2));
	jspl jspl_w_n1535_0(.douta(w_n1535_0[0]),.doutb(w_n1535_0[1]),.din(n1535));
	jspl jspl_w_n1537_0(.douta(w_n1537_0[0]),.doutb(w_n1537_0[1]),.din(n1537));
	jspl jspl_w_n1538_0(.douta(w_n1538_0[0]),.doutb(w_n1538_0[1]),.din(n1538));
	jspl jspl_w_n1539_0(.douta(w_n1539_0[0]),.doutb(w_n1539_0[1]),.din(n1539));
	jspl jspl_w_n1540_0(.douta(w_n1540_0[0]),.doutb(w_n1540_0[1]),.din(n1540));
	jspl jspl_w_n1541_0(.douta(w_n1541_0[0]),.doutb(w_n1541_0[1]),.din(n1541));
	jspl jspl_w_n1542_0(.douta(w_n1542_0[0]),.doutb(w_n1542_0[1]),.din(n1542));
	jspl jspl_w_n1543_0(.douta(w_n1543_0[0]),.doutb(w_n1543_0[1]),.din(n1543));
	jspl jspl_w_n1544_0(.douta(w_n1544_0[0]),.doutb(w_n1544_0[1]),.din(n1544));
	jspl jspl_w_n1545_0(.douta(w_n1545_0[0]),.doutb(w_n1545_0[1]),.din(n1545));
	jspl jspl_w_n1546_0(.douta(w_n1546_0[0]),.doutb(w_n1546_0[1]),.din(n1546));
	jspl jspl_w_n1547_0(.douta(w_n1547_0[0]),.doutb(w_n1547_0[1]),.din(n1547));
	jspl jspl_w_n1548_0(.douta(w_n1548_0[0]),.doutb(w_n1548_0[1]),.din(w_dff_B_DhnMH88a8_2));
	jspl jspl_w_n1549_0(.douta(w_n1549_0[0]),.doutb(w_n1549_0[1]),.din(n1549));
	jspl jspl_w_n1550_0(.douta(w_n1550_0[0]),.doutb(w_dff_A_NoaSoI4S5_1),.din(n1550));
	jspl jspl_w_n1552_0(.douta(w_n1552_0[0]),.doutb(w_n1552_0[1]),.din(n1552));
	jspl jspl_w_n1554_0(.douta(w_n1554_0[0]),.doutb(w_n1554_0[1]),.din(n1554));
	jspl jspl_w_n1555_0(.douta(w_n1555_0[0]),.doutb(w_dff_A_0GFTuX1r9_1),.din(n1555));
	jspl jspl_w_n1560_0(.douta(w_n1560_0[0]),.doutb(w_n1560_0[1]),.din(n1560));
	jspl jspl_w_n1565_0(.douta(w_n1565_0[0]),.doutb(w_n1565_0[1]),.din(n1565));
	jspl jspl_w_n1566_0(.douta(w_n1566_0[0]),.doutb(w_n1566_0[1]),.din(w_dff_B_4gjy0nN20_2));
	jspl jspl_w_n1569_0(.douta(w_n1569_0[0]),.doutb(w_n1569_0[1]),.din(n1569));
	jspl jspl_w_n1571_0(.douta(w_n1571_0[0]),.doutb(w_n1571_0[1]),.din(w_dff_B_zYjooRPh7_2));
	jspl jspl_w_n1574_0(.douta(w_n1574_0[0]),.doutb(w_n1574_0[1]),.din(w_dff_B_rKUlpOpo5_2));
	jspl jspl_w_n1576_0(.douta(w_n1576_0[0]),.doutb(w_n1576_0[1]),.din(w_dff_B_PlW01fJO6_2));
	jspl jspl_w_n1579_0(.douta(w_n1579_0[0]),.doutb(w_n1579_0[1]),.din(w_dff_B_k6Z3dM301_2));
	jspl jspl_w_n1581_0(.douta(w_n1581_0[0]),.doutb(w_n1581_0[1]),.din(w_dff_B_fmCt4rpQ0_2));
	jspl jspl_w_n1584_0(.douta(w_n1584_0[0]),.doutb(w_n1584_0[1]),.din(w_dff_B_Us3zuZTo6_2));
	jspl jspl_w_n1586_0(.douta(w_n1586_0[0]),.doutb(w_n1586_0[1]),.din(w_dff_B_89y1K2Xs8_2));
	jspl jspl_w_n1589_0(.douta(w_n1589_0[0]),.doutb(w_n1589_0[1]),.din(w_dff_B_mk4QHZQS7_2));
	jspl jspl_w_n1591_0(.douta(w_n1591_0[0]),.doutb(w_n1591_0[1]),.din(w_dff_B_poyiy4tx3_2));
	jspl jspl_w_n1594_0(.douta(w_n1594_0[0]),.doutb(w_n1594_0[1]),.din(w_dff_B_896xBcra0_2));
	jspl jspl_w_n1595_0(.douta(w_n1595_0[0]),.doutb(w_n1595_0[1]),.din(w_dff_B_Dk0tMq5b9_2));
	jspl jspl_w_n1596_0(.douta(w_n1596_0[0]),.doutb(w_n1596_0[1]),.din(w_dff_B_k33KKcJH0_2));
	jspl jspl_w_n1599_0(.douta(w_n1599_0[0]),.doutb(w_n1599_0[1]),.din(n1599));
	jspl jspl_w_n1601_0(.douta(w_n1601_0[0]),.doutb(w_n1601_0[1]),.din(n1601));
	jspl jspl_w_n1602_0(.douta(w_n1602_0[0]),.doutb(w_n1602_0[1]),.din(n1602));
	jspl jspl_w_n1603_0(.douta(w_n1603_0[0]),.doutb(w_n1603_0[1]),.din(n1603));
	jspl jspl_w_n1604_0(.douta(w_n1604_0[0]),.doutb(w_n1604_0[1]),.din(n1604));
	jspl jspl_w_n1605_0(.douta(w_n1605_0[0]),.doutb(w_n1605_0[1]),.din(n1605));
	jspl jspl_w_n1606_0(.douta(w_n1606_0[0]),.doutb(w_n1606_0[1]),.din(n1606));
	jspl jspl_w_n1607_0(.douta(w_n1607_0[0]),.doutb(w_n1607_0[1]),.din(n1607));
	jspl jspl_w_n1608_0(.douta(w_n1608_0[0]),.doutb(w_n1608_0[1]),.din(n1608));
	jspl jspl_w_n1609_0(.douta(w_n1609_0[0]),.doutb(w_n1609_0[1]),.din(n1609));
	jspl jspl_w_n1610_0(.douta(w_n1610_0[0]),.doutb(w_n1610_0[1]),.din(n1610));
	jspl jspl_w_n1611_0(.douta(w_n1611_0[0]),.doutb(w_n1611_0[1]),.din(n1611));
	jspl jspl_w_n1612_0(.douta(w_n1612_0[0]),.doutb(w_n1612_0[1]),.din(n1612));
	jspl jspl_w_n1614_0(.douta(w_n1614_0[0]),.doutb(w_n1614_0[1]),.din(n1614));
	jspl jspl_w_n1616_0(.douta(w_n1616_0[0]),.doutb(w_n1616_0[1]),.din(n1616));
	jspl jspl_w_n1617_0(.douta(w_n1617_0[0]),.doutb(w_dff_A_1K1g5fbW6_1),.din(n1617));
	jspl jspl_w_n1622_0(.douta(w_n1622_0[0]),.doutb(w_n1622_0[1]),.din(n1622));
	jspl jspl_w_n1627_0(.douta(w_n1627_0[0]),.doutb(w_n1627_0[1]),.din(w_dff_B_qO9LQxKl1_2));
	jspl jspl_w_n1628_0(.douta(w_n1628_0[0]),.doutb(w_n1628_0[1]),.din(w_dff_B_8udX8bne1_2));
	jspl jspl_w_n1631_0(.douta(w_n1631_0[0]),.doutb(w_dff_A_4JJX4vbh2_1),.din(n1631));
	jspl jspl_w_n1633_0(.douta(w_n1633_0[0]),.doutb(w_n1633_0[1]),.din(w_dff_B_t7NTSo022_2));
	jspl jspl_w_n1636_0(.douta(w_n1636_0[0]),.doutb(w_n1636_0[1]),.din(w_dff_B_gEWZXbi90_2));
	jspl jspl_w_n1638_0(.douta(w_n1638_0[0]),.doutb(w_n1638_0[1]),.din(w_dff_B_gg96ixUT7_2));
	jspl jspl_w_n1641_0(.douta(w_n1641_0[0]),.doutb(w_n1641_0[1]),.din(w_dff_B_RlKTCuxy7_2));
	jspl jspl_w_n1643_0(.douta(w_n1643_0[0]),.doutb(w_n1643_0[1]),.din(w_dff_B_49g8mCix4_2));
	jspl jspl_w_n1646_0(.douta(w_n1646_0[0]),.doutb(w_n1646_0[1]),.din(w_dff_B_D0oz23es3_2));
	jspl jspl_w_n1648_0(.douta(w_n1648_0[0]),.doutb(w_n1648_0[1]),.din(w_dff_B_FH7jW32D5_2));
	jspl jspl_w_n1651_0(.douta(w_n1651_0[0]),.doutb(w_n1651_0[1]),.din(w_dff_B_IGBSwx534_2));
	jspl jspl_w_n1652_0(.douta(w_n1652_0[0]),.doutb(w_n1652_0[1]),.din(w_dff_B_NufzxXYp2_2));
	jspl jspl_w_n1653_0(.douta(w_n1653_0[0]),.doutb(w_n1653_0[1]),.din(w_dff_B_gllUR0MF3_2));
	jspl jspl_w_n1656_0(.douta(w_n1656_0[0]),.doutb(w_n1656_0[1]),.din(n1656));
	jspl jspl_w_n1658_0(.douta(w_n1658_0[0]),.doutb(w_n1658_0[1]),.din(n1658));
	jspl jspl_w_n1659_0(.douta(w_n1659_0[0]),.doutb(w_n1659_0[1]),.din(n1659));
	jspl jspl_w_n1660_0(.douta(w_n1660_0[0]),.doutb(w_n1660_0[1]),.din(n1660));
	jspl jspl_w_n1661_0(.douta(w_n1661_0[0]),.doutb(w_n1661_0[1]),.din(n1661));
	jspl jspl_w_n1662_0(.douta(w_n1662_0[0]),.doutb(w_n1662_0[1]),.din(n1662));
	jspl jspl_w_n1663_0(.douta(w_n1663_0[0]),.doutb(w_n1663_0[1]),.din(n1663));
	jspl jspl_w_n1664_0(.douta(w_n1664_0[0]),.doutb(w_n1664_0[1]),.din(n1664));
	jspl jspl_w_n1665_0(.douta(w_n1665_0[0]),.doutb(w_n1665_0[1]),.din(n1665));
	jspl jspl_w_n1666_0(.douta(w_n1666_0[0]),.doutb(w_n1666_0[1]),.din(n1666));
	jspl jspl_w_n1667_0(.douta(w_n1667_0[0]),.doutb(w_n1667_0[1]),.din(n1667));
	jspl jspl_w_n1669_0(.douta(w_n1669_0[0]),.doutb(w_n1669_0[1]),.din(n1669));
	jspl jspl_w_n1671_0(.douta(w_n1671_0[0]),.doutb(w_n1671_0[1]),.din(n1671));
	jspl jspl_w_n1672_0(.douta(w_n1672_0[0]),.doutb(w_dff_A_alqW54nR6_1),.din(n1672));
	jspl jspl_w_n1677_0(.douta(w_n1677_0[0]),.doutb(w_n1677_0[1]),.din(n1677));
	jspl jspl_w_n1682_0(.douta(w_n1682_0[0]),.doutb(w_n1682_0[1]),.din(w_dff_B_3RnJicDM9_2));
	jspl jspl_w_n1684_0(.douta(w_n1684_0[0]),.doutb(w_n1684_0[1]),.din(w_dff_B_1pDKIZ093_2));
	jspl jspl_w_n1687_0(.douta(w_n1687_0[0]),.doutb(w_n1687_0[1]),.din(w_dff_B_N2jdzGk90_2));
	jspl jspl_w_n1689_0(.douta(w_n1689_0[0]),.doutb(w_n1689_0[1]),.din(w_dff_B_nj4zgaFg1_2));
	jspl jspl_w_n1692_0(.douta(w_n1692_0[0]),.doutb(w_n1692_0[1]),.din(w_dff_B_jVVl5q6J8_2));
	jspl jspl_w_n1694_0(.douta(w_n1694_0[0]),.doutb(w_n1694_0[1]),.din(w_dff_B_icbpygs14_2));
	jspl jspl_w_n1697_0(.douta(w_n1697_0[0]),.doutb(w_n1697_0[1]),.din(w_dff_B_CWjW9Ljq8_2));
	jspl jspl_w_n1699_0(.douta(w_n1699_0[0]),.doutb(w_n1699_0[1]),.din(w_dff_B_YpBZ67h04_2));
	jspl jspl_w_n1702_0(.douta(w_n1702_0[0]),.doutb(w_n1702_0[1]),.din(w_dff_B_hrir7I2z8_2));
	jspl jspl_w_n1703_0(.douta(w_n1703_0[0]),.doutb(w_n1703_0[1]),.din(w_dff_B_kv4gH2Zd2_2));
	jspl jspl_w_n1704_0(.douta(w_n1704_0[0]),.doutb(w_n1704_0[1]),.din(w_dff_B_ftAC1Tv30_2));
	jspl jspl_w_n1707_0(.douta(w_n1707_0[0]),.doutb(w_n1707_0[1]),.din(n1707));
	jspl jspl_w_n1709_0(.douta(w_n1709_0[0]),.doutb(w_n1709_0[1]),.din(n1709));
	jspl jspl_w_n1710_0(.douta(w_n1710_0[0]),.doutb(w_n1710_0[1]),.din(n1710));
	jspl jspl_w_n1711_0(.douta(w_n1711_0[0]),.doutb(w_n1711_0[1]),.din(n1711));
	jspl jspl_w_n1712_0(.douta(w_n1712_0[0]),.doutb(w_n1712_0[1]),.din(n1712));
	jspl jspl_w_n1713_0(.douta(w_n1713_0[0]),.doutb(w_n1713_0[1]),.din(n1713));
	jspl jspl_w_n1714_0(.douta(w_n1714_0[0]),.doutb(w_n1714_0[1]),.din(n1714));
	jspl jspl_w_n1715_0(.douta(w_n1715_0[0]),.doutb(w_n1715_0[1]),.din(n1715));
	jspl jspl_w_n1716_0(.douta(w_n1716_0[0]),.doutb(w_n1716_0[1]),.din(n1716));
	jspl jspl_w_n1717_0(.douta(w_n1717_0[0]),.doutb(w_n1717_0[1]),.din(n1717));
	jspl jspl_w_n1719_0(.douta(w_n1719_0[0]),.doutb(w_n1719_0[1]),.din(n1719));
	jspl jspl_w_n1720_0(.douta(w_n1720_0[0]),.doutb(w_dff_A_mHhCd8B79_1),.din(n1720));
	jspl jspl_w_n1725_0(.douta(w_n1725_0[0]),.doutb(w_n1725_0[1]),.din(n1725));
	jspl jspl_w_n1728_0(.douta(w_n1728_0[0]),.doutb(w_dff_A_gs11IcZb5_1),.din(n1728));
	jspl jspl_w_n1730_0(.douta(w_n1730_0[0]),.doutb(w_n1730_0[1]),.din(w_dff_B_xe0e7oJ50_2));
	jspl jspl_w_n1733_0(.douta(w_n1733_0[0]),.doutb(w_n1733_0[1]),.din(w_dff_B_bUQI7BuH1_2));
	jspl jspl_w_n1735_0(.douta(w_n1735_0[0]),.doutb(w_n1735_0[1]),.din(w_dff_B_09FlSBNU8_2));
	jspl jspl_w_n1738_0(.douta(w_n1738_0[0]),.doutb(w_n1738_0[1]),.din(w_dff_B_Hto6pA017_2));
	jspl jspl_w_n1740_0(.douta(w_n1740_0[0]),.doutb(w_n1740_0[1]),.din(w_dff_B_DyB1IKPC5_2));
	jspl jspl_w_n1743_0(.douta(w_n1743_0[0]),.doutb(w_n1743_0[1]),.din(w_dff_B_0wdXCfdC9_2));
	jspl jspl_w_n1744_0(.douta(w_n1744_0[0]),.doutb(w_n1744_0[1]),.din(w_dff_B_B7RNIbNT7_2));
	jspl jspl_w_n1745_0(.douta(w_n1745_0[0]),.doutb(w_n1745_0[1]),.din(w_dff_B_XccXmWny7_2));
	jspl jspl_w_n1748_0(.douta(w_n1748_0[0]),.doutb(w_n1748_0[1]),.din(n1748));
	jspl jspl_w_n1750_0(.douta(w_n1750_0[0]),.doutb(w_n1750_0[1]),.din(n1750));
	jspl jspl_w_n1751_0(.douta(w_n1751_0[0]),.doutb(w_n1751_0[1]),.din(n1751));
	jspl jspl_w_n1752_0(.douta(w_n1752_0[0]),.doutb(w_n1752_0[1]),.din(n1752));
	jspl jspl_w_n1753_0(.douta(w_n1753_0[0]),.doutb(w_n1753_0[1]),.din(n1753));
	jspl jspl_w_n1754_0(.douta(w_n1754_0[0]),.doutb(w_n1754_0[1]),.din(n1754));
	jspl jspl_w_n1755_0(.douta(w_n1755_0[0]),.doutb(w_n1755_0[1]),.din(n1755));
	jspl jspl_w_n1756_0(.douta(w_n1756_0[0]),.doutb(w_n1756_0[1]),.din(n1756));
	jspl jspl_w_n1757_0(.douta(w_n1757_0[0]),.doutb(w_n1757_0[1]),.din(n1757));
	jspl jspl_w_n1758_0(.douta(w_n1758_0[0]),.doutb(w_dff_A_RlkqRC6Q9_1),.din(n1758));
	jspl jspl_w_n1765_0(.douta(w_n1765_0[0]),.doutb(w_n1765_0[1]),.din(n1765));
	jspl jspl_w_n1768_0(.douta(w_n1768_0[0]),.doutb(w_dff_A_WItlfLpC4_1),.din(n1768));
	jspl jspl_w_n1770_0(.douta(w_n1770_0[0]),.doutb(w_n1770_0[1]),.din(w_dff_B_Yzc9RcZh4_2));
	jspl jspl_w_n1773_0(.douta(w_n1773_0[0]),.doutb(w_n1773_0[1]),.din(w_dff_B_2XG2nvNA2_2));
	jspl jspl_w_n1775_0(.douta(w_n1775_0[0]),.doutb(w_n1775_0[1]),.din(w_dff_B_KRSHZt2L9_2));
	jspl jspl_w_n1778_0(.douta(w_n1778_0[0]),.doutb(w_n1778_0[1]),.din(w_dff_B_agF8t62T8_2));
	jspl jspl_w_n1779_0(.douta(w_n1779_0[0]),.doutb(w_n1779_0[1]),.din(w_dff_B_qFmd4odf4_2));
	jspl jspl_w_n1780_0(.douta(w_n1780_0[0]),.doutb(w_n1780_0[1]),.din(w_dff_B_T0DnmlcE6_2));
	jspl jspl_w_n1783_0(.douta(w_n1783_0[0]),.doutb(w_n1783_0[1]),.din(n1783));
	jspl jspl_w_n1785_0(.douta(w_n1785_0[0]),.doutb(w_n1785_0[1]),.din(n1785));
	jspl jspl_w_n1786_0(.douta(w_n1786_0[0]),.doutb(w_n1786_0[1]),.din(n1786));
	jspl jspl_w_n1787_0(.douta(w_n1787_0[0]),.doutb(w_n1787_0[1]),.din(n1787));
	jspl jspl_w_n1788_0(.douta(w_n1788_0[0]),.doutb(w_n1788_0[1]),.din(n1788));
	jspl jspl_w_n1789_0(.douta(w_n1789_0[0]),.doutb(w_n1789_0[1]),.din(n1789));
	jspl jspl_w_n1790_0(.douta(w_n1790_0[0]),.doutb(w_n1790_0[1]),.din(n1790));
	jspl jspl_w_n1791_0(.douta(w_n1791_0[0]),.doutb(w_dff_A_DbyttkQU3_1),.din(n1791));
	jspl jspl_w_n1798_0(.douta(w_n1798_0[0]),.doutb(w_n1798_0[1]),.din(n1798));
	jspl jspl_w_n1801_0(.douta(w_n1801_0[0]),.doutb(w_dff_A_yvPCCEoS2_1),.din(n1801));
	jspl jspl_w_n1803_0(.douta(w_n1803_0[0]),.doutb(w_n1803_0[1]),.din(w_dff_B_iy3NUKPE5_2));
	jspl jspl_w_n1806_0(.douta(w_n1806_0[0]),.doutb(w_n1806_0[1]),.din(w_dff_B_qwcLaNmX5_2));
	jspl jspl_w_n1807_0(.douta(w_n1807_0[0]),.doutb(w_n1807_0[1]),.din(w_dff_B_eAyBbxsi5_2));
	jspl jspl_w_n1808_0(.douta(w_n1808_0[0]),.doutb(w_n1808_0[1]),.din(w_dff_B_qDLH0N856_2));
	jspl jspl_w_n1811_0(.douta(w_n1811_0[0]),.doutb(w_n1811_0[1]),.din(n1811));
	jspl jspl_w_n1813_0(.douta(w_n1813_0[0]),.doutb(w_n1813_0[1]),.din(n1813));
	jspl jspl_w_n1814_0(.douta(w_n1814_0[0]),.doutb(w_n1814_0[1]),.din(n1814));
	jspl jspl_w_n1815_0(.douta(w_n1815_0[0]),.doutb(w_n1815_0[1]),.din(n1815));
	jspl jspl_w_n1816_0(.douta(w_n1816_0[0]),.doutb(w_n1816_0[1]),.din(n1816));
	jspl jspl_w_n1817_0(.douta(w_n1817_0[0]),.doutb(w_dff_A_axlC0KEc6_1),.din(n1817));
	jspl jspl_w_n1824_0(.douta(w_n1824_0[0]),.doutb(w_n1824_0[1]),.din(n1824));
	jspl jspl_w_n1827_0(.douta(w_n1827_0[0]),.doutb(w_dff_A_Gl0YM9RQ1_1),.din(n1827));
	jspl jspl_w_n1828_0(.douta(w_n1828_0[0]),.doutb(w_n1828_0[1]),.din(w_dff_B_eP2sF8fc1_2));
	jspl jspl_w_n1829_0(.douta(w_n1829_0[0]),.doutb(w_n1829_0[1]),.din(w_dff_B_1EHsxoj72_2));
	jspl jspl_w_n1832_0(.douta(w_n1832_0[0]),.doutb(w_n1832_0[1]),.din(n1832));
	jspl jspl_w_n1834_0(.douta(w_n1834_0[0]),.doutb(w_n1834_0[1]),.din(n1834));
	jspl jspl_w_n1835_0(.douta(w_n1835_0[0]),.doutb(w_n1835_0[1]),.din(n1835));
	jspl jspl_w_n1836_0(.douta(w_n1836_0[0]),.doutb(w_dff_A_TxFnIYqv4_1),.din(n1836));
	jspl jspl_w_n1838_0(.douta(w_n1838_0[0]),.doutb(w_n1838_0[1]),.din(w_dff_B_g4xoyXVp5_2));
	jspl jspl_w_n1841_0(.douta(w_n1841_0[0]),.doutb(w_n1841_0[1]),.din(n1841));
	jspl jspl_w_n1848_0(.douta(w_n1848_0[0]),.doutb(w_n1848_0[1]),.din(n1848));
	jspl jspl_w_n1849_0(.douta(w_dff_A_AfYw5laX3_0),.doutb(w_n1849_0[1]),.din(n1849));
	jdff dff_B_ORLY9DPs0_1(.din(n67),.dout(w_dff_B_ORLY9DPs0_1),.clk(gclk));
	jdff dff_B_oZHNDDvI5_1(.din(n73),.dout(w_dff_B_oZHNDDvI5_1),.clk(gclk));
	jdff dff_B_Ij8bIAet5_1(.din(w_dff_B_oZHNDDvI5_1),.dout(w_dff_B_Ij8bIAet5_1),.clk(gclk));
	jdff dff_B_LNzalzae9_1(.din(w_dff_B_Ij8bIAet5_1),.dout(w_dff_B_LNzalzae9_1),.clk(gclk));
	jdff dff_B_G2992b235_1(.din(w_dff_B_LNzalzae9_1),.dout(w_dff_B_G2992b235_1),.clk(gclk));
	jdff dff_B_Y9xjsZpf4_1(.din(n90),.dout(w_dff_B_Y9xjsZpf4_1),.clk(gclk));
	jdff dff_B_cB49q0lG3_1(.din(w_dff_B_Y9xjsZpf4_1),.dout(w_dff_B_cB49q0lG3_1),.clk(gclk));
	jdff dff_B_w7BFs5Bb5_1(.din(w_dff_B_cB49q0lG3_1),.dout(w_dff_B_w7BFs5Bb5_1),.clk(gclk));
	jdff dff_B_gK2wT7JT1_1(.din(w_dff_B_w7BFs5Bb5_1),.dout(w_dff_B_gK2wT7JT1_1),.clk(gclk));
	jdff dff_B_eri50NwL8_1(.din(w_dff_B_gK2wT7JT1_1),.dout(w_dff_B_eri50NwL8_1),.clk(gclk));
	jdff dff_B_sHtfu03p8_1(.din(w_dff_B_eri50NwL8_1),.dout(w_dff_B_sHtfu03p8_1),.clk(gclk));
	jdff dff_B_YgdLPBYN7_1(.din(w_dff_B_sHtfu03p8_1),.dout(w_dff_B_YgdLPBYN7_1),.clk(gclk));
	jdff dff_B_7odUktbF4_1(.din(n111),.dout(w_dff_B_7odUktbF4_1),.clk(gclk));
	jdff dff_B_AIe7hqhN6_1(.din(w_dff_B_7odUktbF4_1),.dout(w_dff_B_AIe7hqhN6_1),.clk(gclk));
	jdff dff_B_LtMhjqtt0_1(.din(w_dff_B_AIe7hqhN6_1),.dout(w_dff_B_LtMhjqtt0_1),.clk(gclk));
	jdff dff_B_E8jnQa4e2_1(.din(w_dff_B_LtMhjqtt0_1),.dout(w_dff_B_E8jnQa4e2_1),.clk(gclk));
	jdff dff_B_k0vSFOZe6_1(.din(w_dff_B_E8jnQa4e2_1),.dout(w_dff_B_k0vSFOZe6_1),.clk(gclk));
	jdff dff_B_KTFb8unQ6_1(.din(w_dff_B_k0vSFOZe6_1),.dout(w_dff_B_KTFb8unQ6_1),.clk(gclk));
	jdff dff_B_JaqLzDzK5_1(.din(w_dff_B_KTFb8unQ6_1),.dout(w_dff_B_JaqLzDzK5_1),.clk(gclk));
	jdff dff_B_UaZUS7uq1_1(.din(w_dff_B_JaqLzDzK5_1),.dout(w_dff_B_UaZUS7uq1_1),.clk(gclk));
	jdff dff_B_Gw3gHxAU9_1(.din(w_dff_B_UaZUS7uq1_1),.dout(w_dff_B_Gw3gHxAU9_1),.clk(gclk));
	jdff dff_B_M40SSfNW0_1(.din(w_dff_B_Gw3gHxAU9_1),.dout(w_dff_B_M40SSfNW0_1),.clk(gclk));
	jdff dff_B_k9xHOgEo2_1(.din(n146),.dout(w_dff_B_k9xHOgEo2_1),.clk(gclk));
	jdff dff_B_EBqLY7Wb5_1(.din(w_dff_B_k9xHOgEo2_1),.dout(w_dff_B_EBqLY7Wb5_1),.clk(gclk));
	jdff dff_B_r2MimJxL5_1(.din(w_dff_B_EBqLY7Wb5_1),.dout(w_dff_B_r2MimJxL5_1),.clk(gclk));
	jdff dff_B_IuaNMIbD0_1(.din(w_dff_B_r2MimJxL5_1),.dout(w_dff_B_IuaNMIbD0_1),.clk(gclk));
	jdff dff_B_IX9gG3S53_1(.din(w_dff_B_IuaNMIbD0_1),.dout(w_dff_B_IX9gG3S53_1),.clk(gclk));
	jdff dff_B_LRtb1ykq6_1(.din(w_dff_B_IX9gG3S53_1),.dout(w_dff_B_LRtb1ykq6_1),.clk(gclk));
	jdff dff_B_JDdX9bxa1_1(.din(w_dff_B_LRtb1ykq6_1),.dout(w_dff_B_JDdX9bxa1_1),.clk(gclk));
	jdff dff_B_g2lSI0ru0_1(.din(w_dff_B_JDdX9bxa1_1),.dout(w_dff_B_g2lSI0ru0_1),.clk(gclk));
	jdff dff_B_QBhLXg9E7_1(.din(w_dff_B_g2lSI0ru0_1),.dout(w_dff_B_QBhLXg9E7_1),.clk(gclk));
	jdff dff_B_6ndOoDWP9_1(.din(w_dff_B_QBhLXg9E7_1),.dout(w_dff_B_6ndOoDWP9_1),.clk(gclk));
	jdff dff_B_xCeUiCs86_1(.din(w_dff_B_6ndOoDWP9_1),.dout(w_dff_B_xCeUiCs86_1),.clk(gclk));
	jdff dff_B_oAZrojAF4_1(.din(w_dff_B_xCeUiCs86_1),.dout(w_dff_B_oAZrojAF4_1),.clk(gclk));
	jdff dff_B_Blu890lS8_1(.din(w_dff_B_oAZrojAF4_1),.dout(w_dff_B_Blu890lS8_1),.clk(gclk));
	jdff dff_B_XmDg2Ir85_1(.din(n184),.dout(w_dff_B_XmDg2Ir85_1),.clk(gclk));
	jdff dff_B_sWBqXna13_1(.din(w_dff_B_XmDg2Ir85_1),.dout(w_dff_B_sWBqXna13_1),.clk(gclk));
	jdff dff_B_eH6mOT2k8_1(.din(w_dff_B_sWBqXna13_1),.dout(w_dff_B_eH6mOT2k8_1),.clk(gclk));
	jdff dff_B_h6aemqzt4_1(.din(w_dff_B_eH6mOT2k8_1),.dout(w_dff_B_h6aemqzt4_1),.clk(gclk));
	jdff dff_B_zCAitGh83_1(.din(w_dff_B_h6aemqzt4_1),.dout(w_dff_B_zCAitGh83_1),.clk(gclk));
	jdff dff_B_yFASLsDr1_1(.din(w_dff_B_zCAitGh83_1),.dout(w_dff_B_yFASLsDr1_1),.clk(gclk));
	jdff dff_B_IJSxLSEe1_1(.din(w_dff_B_yFASLsDr1_1),.dout(w_dff_B_IJSxLSEe1_1),.clk(gclk));
	jdff dff_B_PFVS4DSZ5_1(.din(w_dff_B_IJSxLSEe1_1),.dout(w_dff_B_PFVS4DSZ5_1),.clk(gclk));
	jdff dff_B_n6Xnw4qU0_1(.din(w_dff_B_PFVS4DSZ5_1),.dout(w_dff_B_n6Xnw4qU0_1),.clk(gclk));
	jdff dff_B_0AmiNKMU8_1(.din(w_dff_B_n6Xnw4qU0_1),.dout(w_dff_B_0AmiNKMU8_1),.clk(gclk));
	jdff dff_B_dopvKpGm6_1(.din(w_dff_B_0AmiNKMU8_1),.dout(w_dff_B_dopvKpGm6_1),.clk(gclk));
	jdff dff_B_rkGExKL76_1(.din(w_dff_B_dopvKpGm6_1),.dout(w_dff_B_rkGExKL76_1),.clk(gclk));
	jdff dff_B_vaHARmQP2_1(.din(w_dff_B_rkGExKL76_1),.dout(w_dff_B_vaHARmQP2_1),.clk(gclk));
	jdff dff_B_EOhZpgfC5_1(.din(w_dff_B_vaHARmQP2_1),.dout(w_dff_B_EOhZpgfC5_1),.clk(gclk));
	jdff dff_B_1N97qTn32_1(.din(w_dff_B_EOhZpgfC5_1),.dout(w_dff_B_1N97qTn32_1),.clk(gclk));
	jdff dff_B_tADF5loM5_1(.din(w_dff_B_1N97qTn32_1),.dout(w_dff_B_tADF5loM5_1),.clk(gclk));
	jdff dff_B_oz165xF91_1(.din(n227),.dout(w_dff_B_oz165xF91_1),.clk(gclk));
	jdff dff_B_7xNgGFpp8_1(.din(w_dff_B_oz165xF91_1),.dout(w_dff_B_7xNgGFpp8_1),.clk(gclk));
	jdff dff_B_tRx9jQr35_1(.din(w_dff_B_7xNgGFpp8_1),.dout(w_dff_B_tRx9jQr35_1),.clk(gclk));
	jdff dff_B_Ryqjbisa9_1(.din(w_dff_B_tRx9jQr35_1),.dout(w_dff_B_Ryqjbisa9_1),.clk(gclk));
	jdff dff_B_Y3zQrAZz4_1(.din(w_dff_B_Ryqjbisa9_1),.dout(w_dff_B_Y3zQrAZz4_1),.clk(gclk));
	jdff dff_B_FqB3WI4q8_1(.din(w_dff_B_Y3zQrAZz4_1),.dout(w_dff_B_FqB3WI4q8_1),.clk(gclk));
	jdff dff_B_to8w4a7x0_1(.din(w_dff_B_FqB3WI4q8_1),.dout(w_dff_B_to8w4a7x0_1),.clk(gclk));
	jdff dff_B_OU0FYghf6_1(.din(w_dff_B_to8w4a7x0_1),.dout(w_dff_B_OU0FYghf6_1),.clk(gclk));
	jdff dff_B_H5DkQQS58_1(.din(w_dff_B_OU0FYghf6_1),.dout(w_dff_B_H5DkQQS58_1),.clk(gclk));
	jdff dff_B_0lzxZQvI1_1(.din(w_dff_B_H5DkQQS58_1),.dout(w_dff_B_0lzxZQvI1_1),.clk(gclk));
	jdff dff_B_sGY503si0_1(.din(w_dff_B_0lzxZQvI1_1),.dout(w_dff_B_sGY503si0_1),.clk(gclk));
	jdff dff_B_N40UKXNQ2_1(.din(w_dff_B_sGY503si0_1),.dout(w_dff_B_N40UKXNQ2_1),.clk(gclk));
	jdff dff_B_hNRrtrSy6_1(.din(w_dff_B_N40UKXNQ2_1),.dout(w_dff_B_hNRrtrSy6_1),.clk(gclk));
	jdff dff_B_kCq1Pjjp4_1(.din(w_dff_B_hNRrtrSy6_1),.dout(w_dff_B_kCq1Pjjp4_1),.clk(gclk));
	jdff dff_B_5hSiQmj88_1(.din(w_dff_B_kCq1Pjjp4_1),.dout(w_dff_B_5hSiQmj88_1),.clk(gclk));
	jdff dff_B_53B8NZmX8_1(.din(w_dff_B_5hSiQmj88_1),.dout(w_dff_B_53B8NZmX8_1),.clk(gclk));
	jdff dff_B_sVGJtqzn0_1(.din(w_dff_B_53B8NZmX8_1),.dout(w_dff_B_sVGJtqzn0_1),.clk(gclk));
	jdff dff_B_R1c7Z2Ac4_1(.din(w_dff_B_sVGJtqzn0_1),.dout(w_dff_B_R1c7Z2Ac4_1),.clk(gclk));
	jdff dff_B_Rstyn61Z1_1(.din(w_dff_B_R1c7Z2Ac4_1),.dout(w_dff_B_Rstyn61Z1_1),.clk(gclk));
	jdff dff_B_VB1NPt8j4_1(.din(n278),.dout(w_dff_B_VB1NPt8j4_1),.clk(gclk));
	jdff dff_B_ZXGd2pai9_1(.din(w_dff_B_VB1NPt8j4_1),.dout(w_dff_B_ZXGd2pai9_1),.clk(gclk));
	jdff dff_B_HpRRLtSh1_1(.din(w_dff_B_ZXGd2pai9_1),.dout(w_dff_B_HpRRLtSh1_1),.clk(gclk));
	jdff dff_B_BP6dCCub8_1(.din(w_dff_B_HpRRLtSh1_1),.dout(w_dff_B_BP6dCCub8_1),.clk(gclk));
	jdff dff_B_7EYqV7Xu1_1(.din(w_dff_B_BP6dCCub8_1),.dout(w_dff_B_7EYqV7Xu1_1),.clk(gclk));
	jdff dff_B_W4LGGPQG0_1(.din(w_dff_B_7EYqV7Xu1_1),.dout(w_dff_B_W4LGGPQG0_1),.clk(gclk));
	jdff dff_B_9mt1mbrt9_1(.din(w_dff_B_W4LGGPQG0_1),.dout(w_dff_B_9mt1mbrt9_1),.clk(gclk));
	jdff dff_B_MeN2bBFT2_1(.din(w_dff_B_9mt1mbrt9_1),.dout(w_dff_B_MeN2bBFT2_1),.clk(gclk));
	jdff dff_B_MNcptmay2_1(.din(w_dff_B_MeN2bBFT2_1),.dout(w_dff_B_MNcptmay2_1),.clk(gclk));
	jdff dff_B_80TRIpfk9_1(.din(w_dff_B_MNcptmay2_1),.dout(w_dff_B_80TRIpfk9_1),.clk(gclk));
	jdff dff_B_YMAcT9ym8_1(.din(w_dff_B_80TRIpfk9_1),.dout(w_dff_B_YMAcT9ym8_1),.clk(gclk));
	jdff dff_B_dnK0GQsU2_1(.din(w_dff_B_YMAcT9ym8_1),.dout(w_dff_B_dnK0GQsU2_1),.clk(gclk));
	jdff dff_B_Tpuf8Jvi6_1(.din(w_dff_B_dnK0GQsU2_1),.dout(w_dff_B_Tpuf8Jvi6_1),.clk(gclk));
	jdff dff_B_piRrKy2c2_1(.din(w_dff_B_Tpuf8Jvi6_1),.dout(w_dff_B_piRrKy2c2_1),.clk(gclk));
	jdff dff_B_r4gZneIh8_1(.din(w_dff_B_piRrKy2c2_1),.dout(w_dff_B_r4gZneIh8_1),.clk(gclk));
	jdff dff_B_ZDLBo6Uh5_1(.din(w_dff_B_r4gZneIh8_1),.dout(w_dff_B_ZDLBo6Uh5_1),.clk(gclk));
	jdff dff_B_WzugrBuw6_1(.din(w_dff_B_ZDLBo6Uh5_1),.dout(w_dff_B_WzugrBuw6_1),.clk(gclk));
	jdff dff_B_vQoBen6M1_1(.din(w_dff_B_WzugrBuw6_1),.dout(w_dff_B_vQoBen6M1_1),.clk(gclk));
	jdff dff_B_ZqgtYdFw3_1(.din(w_dff_B_vQoBen6M1_1),.dout(w_dff_B_ZqgtYdFw3_1),.clk(gclk));
	jdff dff_B_Cq3OTBLI9_1(.din(w_dff_B_ZqgtYdFw3_1),.dout(w_dff_B_Cq3OTBLI9_1),.clk(gclk));
	jdff dff_B_By0i8jzb1_1(.din(w_dff_B_Cq3OTBLI9_1),.dout(w_dff_B_By0i8jzb1_1),.clk(gclk));
	jdff dff_B_sWvwVGJZ8_1(.din(w_dff_B_By0i8jzb1_1),.dout(w_dff_B_sWvwVGJZ8_1),.clk(gclk));
	jdff dff_B_VoQ6TS7b0_1(.din(n336),.dout(w_dff_B_VoQ6TS7b0_1),.clk(gclk));
	jdff dff_B_Wle8A4Yf0_1(.din(w_dff_B_VoQ6TS7b0_1),.dout(w_dff_B_Wle8A4Yf0_1),.clk(gclk));
	jdff dff_B_UQQW8iTz5_1(.din(w_dff_B_Wle8A4Yf0_1),.dout(w_dff_B_UQQW8iTz5_1),.clk(gclk));
	jdff dff_B_itdCWixZ0_1(.din(w_dff_B_UQQW8iTz5_1),.dout(w_dff_B_itdCWixZ0_1),.clk(gclk));
	jdff dff_B_V5JRKZ0E7_1(.din(w_dff_B_itdCWixZ0_1),.dout(w_dff_B_V5JRKZ0E7_1),.clk(gclk));
	jdff dff_B_nuTxSf3V6_1(.din(w_dff_B_V5JRKZ0E7_1),.dout(w_dff_B_nuTxSf3V6_1),.clk(gclk));
	jdff dff_B_NsCMPFEu6_1(.din(w_dff_B_nuTxSf3V6_1),.dout(w_dff_B_NsCMPFEu6_1),.clk(gclk));
	jdff dff_B_VTRLNAiW9_1(.din(w_dff_B_NsCMPFEu6_1),.dout(w_dff_B_VTRLNAiW9_1),.clk(gclk));
	jdff dff_B_MKOKdvzz0_1(.din(w_dff_B_VTRLNAiW9_1),.dout(w_dff_B_MKOKdvzz0_1),.clk(gclk));
	jdff dff_B_rLdClAAR1_1(.din(w_dff_B_MKOKdvzz0_1),.dout(w_dff_B_rLdClAAR1_1),.clk(gclk));
	jdff dff_B_tjssuTd70_1(.din(w_dff_B_rLdClAAR1_1),.dout(w_dff_B_tjssuTd70_1),.clk(gclk));
	jdff dff_B_OLX31m4k8_1(.din(w_dff_B_tjssuTd70_1),.dout(w_dff_B_OLX31m4k8_1),.clk(gclk));
	jdff dff_B_aIeLOVwR2_1(.din(w_dff_B_OLX31m4k8_1),.dout(w_dff_B_aIeLOVwR2_1),.clk(gclk));
	jdff dff_B_uC8AU9eC6_1(.din(w_dff_B_aIeLOVwR2_1),.dout(w_dff_B_uC8AU9eC6_1),.clk(gclk));
	jdff dff_B_IQ226zB29_1(.din(w_dff_B_uC8AU9eC6_1),.dout(w_dff_B_IQ226zB29_1),.clk(gclk));
	jdff dff_B_G9jovtSI4_1(.din(w_dff_B_IQ226zB29_1),.dout(w_dff_B_G9jovtSI4_1),.clk(gclk));
	jdff dff_B_mmDSTvj04_1(.din(w_dff_B_G9jovtSI4_1),.dout(w_dff_B_mmDSTvj04_1),.clk(gclk));
	jdff dff_B_mDnqxGGm3_1(.din(w_dff_B_mmDSTvj04_1),.dout(w_dff_B_mDnqxGGm3_1),.clk(gclk));
	jdff dff_B_BPQLcRlU0_1(.din(w_dff_B_mDnqxGGm3_1),.dout(w_dff_B_BPQLcRlU0_1),.clk(gclk));
	jdff dff_B_aiGt8Dic1_1(.din(w_dff_B_BPQLcRlU0_1),.dout(w_dff_B_aiGt8Dic1_1),.clk(gclk));
	jdff dff_B_s52Nu9LV3_1(.din(w_dff_B_aiGt8Dic1_1),.dout(w_dff_B_s52Nu9LV3_1),.clk(gclk));
	jdff dff_B_bSVOMIX40_1(.din(w_dff_B_s52Nu9LV3_1),.dout(w_dff_B_bSVOMIX40_1),.clk(gclk));
	jdff dff_B_BJLX2naj7_1(.din(w_dff_B_bSVOMIX40_1),.dout(w_dff_B_BJLX2naj7_1),.clk(gclk));
	jdff dff_B_vcPR8CNy8_1(.din(w_dff_B_BJLX2naj7_1),.dout(w_dff_B_vcPR8CNy8_1),.clk(gclk));
	jdff dff_B_EdoSg5X52_1(.din(w_dff_B_vcPR8CNy8_1),.dout(w_dff_B_EdoSg5X52_1),.clk(gclk));
	jdff dff_B_4gsK11Xq9_1(.din(n400),.dout(w_dff_B_4gsK11Xq9_1),.clk(gclk));
	jdff dff_B_RiXaZqSO7_1(.din(w_dff_B_4gsK11Xq9_1),.dout(w_dff_B_RiXaZqSO7_1),.clk(gclk));
	jdff dff_B_YEdKv2G26_1(.din(w_dff_B_RiXaZqSO7_1),.dout(w_dff_B_YEdKv2G26_1),.clk(gclk));
	jdff dff_B_MqDQFoRb5_1(.din(w_dff_B_YEdKv2G26_1),.dout(w_dff_B_MqDQFoRb5_1),.clk(gclk));
	jdff dff_B_XAk9Ie3e6_1(.din(w_dff_B_MqDQFoRb5_1),.dout(w_dff_B_XAk9Ie3e6_1),.clk(gclk));
	jdff dff_B_ZcCR1UC79_1(.din(w_dff_B_XAk9Ie3e6_1),.dout(w_dff_B_ZcCR1UC79_1),.clk(gclk));
	jdff dff_B_RYAcUgtn8_1(.din(w_dff_B_ZcCR1UC79_1),.dout(w_dff_B_RYAcUgtn8_1),.clk(gclk));
	jdff dff_B_6U4SpEKA3_1(.din(w_dff_B_RYAcUgtn8_1),.dout(w_dff_B_6U4SpEKA3_1),.clk(gclk));
	jdff dff_B_1W6La1mW7_1(.din(w_dff_B_6U4SpEKA3_1),.dout(w_dff_B_1W6La1mW7_1),.clk(gclk));
	jdff dff_B_U3NVz7Gm3_1(.din(w_dff_B_1W6La1mW7_1),.dout(w_dff_B_U3NVz7Gm3_1),.clk(gclk));
	jdff dff_B_uqQY5foB5_1(.din(w_dff_B_U3NVz7Gm3_1),.dout(w_dff_B_uqQY5foB5_1),.clk(gclk));
	jdff dff_B_f8Wxk0BQ4_1(.din(w_dff_B_uqQY5foB5_1),.dout(w_dff_B_f8Wxk0BQ4_1),.clk(gclk));
	jdff dff_B_FdNtK8LV3_1(.din(w_dff_B_f8Wxk0BQ4_1),.dout(w_dff_B_FdNtK8LV3_1),.clk(gclk));
	jdff dff_B_nk4NLpLZ7_1(.din(w_dff_B_FdNtK8LV3_1),.dout(w_dff_B_nk4NLpLZ7_1),.clk(gclk));
	jdff dff_B_uwf0iG056_1(.din(w_dff_B_nk4NLpLZ7_1),.dout(w_dff_B_uwf0iG056_1),.clk(gclk));
	jdff dff_B_NfkAaFSp9_1(.din(w_dff_B_uwf0iG056_1),.dout(w_dff_B_NfkAaFSp9_1),.clk(gclk));
	jdff dff_B_FzXvi16b5_1(.din(w_dff_B_NfkAaFSp9_1),.dout(w_dff_B_FzXvi16b5_1),.clk(gclk));
	jdff dff_B_ssy4zHjc9_1(.din(w_dff_B_FzXvi16b5_1),.dout(w_dff_B_ssy4zHjc9_1),.clk(gclk));
	jdff dff_B_M4pUayoG1_1(.din(w_dff_B_ssy4zHjc9_1),.dout(w_dff_B_M4pUayoG1_1),.clk(gclk));
	jdff dff_B_Cr8Iu6sw6_1(.din(w_dff_B_M4pUayoG1_1),.dout(w_dff_B_Cr8Iu6sw6_1),.clk(gclk));
	jdff dff_B_y9oGrr659_1(.din(w_dff_B_Cr8Iu6sw6_1),.dout(w_dff_B_y9oGrr659_1),.clk(gclk));
	jdff dff_B_leFj1xjK8_1(.din(w_dff_B_y9oGrr659_1),.dout(w_dff_B_leFj1xjK8_1),.clk(gclk));
	jdff dff_B_1SPpOoKH7_1(.din(w_dff_B_leFj1xjK8_1),.dout(w_dff_B_1SPpOoKH7_1),.clk(gclk));
	jdff dff_B_yxOTRkff3_1(.din(w_dff_B_1SPpOoKH7_1),.dout(w_dff_B_yxOTRkff3_1),.clk(gclk));
	jdff dff_B_NXBs2v549_1(.din(w_dff_B_yxOTRkff3_1),.dout(w_dff_B_NXBs2v549_1),.clk(gclk));
	jdff dff_B_QxvYgTXT7_1(.din(w_dff_B_NXBs2v549_1),.dout(w_dff_B_QxvYgTXT7_1),.clk(gclk));
	jdff dff_B_7nDGrMEn4_1(.din(w_dff_B_QxvYgTXT7_1),.dout(w_dff_B_7nDGrMEn4_1),.clk(gclk));
	jdff dff_B_wgsWXVkt3_1(.din(w_dff_B_7nDGrMEn4_1),.dout(w_dff_B_wgsWXVkt3_1),.clk(gclk));
	jdff dff_B_Ng7TGNCt8_1(.din(n472),.dout(w_dff_B_Ng7TGNCt8_1),.clk(gclk));
	jdff dff_B_eBBkXGyg4_1(.din(w_dff_B_Ng7TGNCt8_1),.dout(w_dff_B_eBBkXGyg4_1),.clk(gclk));
	jdff dff_B_5oeXDePC1_1(.din(w_dff_B_eBBkXGyg4_1),.dout(w_dff_B_5oeXDePC1_1),.clk(gclk));
	jdff dff_B_WNVXoER12_1(.din(w_dff_B_5oeXDePC1_1),.dout(w_dff_B_WNVXoER12_1),.clk(gclk));
	jdff dff_B_Uh2Azmw13_1(.din(w_dff_B_WNVXoER12_1),.dout(w_dff_B_Uh2Azmw13_1),.clk(gclk));
	jdff dff_B_LB5rLVW66_1(.din(w_dff_B_Uh2Azmw13_1),.dout(w_dff_B_LB5rLVW66_1),.clk(gclk));
	jdff dff_B_Q251MPaq6_1(.din(w_dff_B_LB5rLVW66_1),.dout(w_dff_B_Q251MPaq6_1),.clk(gclk));
	jdff dff_B_FxOmnJYt7_1(.din(w_dff_B_Q251MPaq6_1),.dout(w_dff_B_FxOmnJYt7_1),.clk(gclk));
	jdff dff_B_b4tasGne0_1(.din(w_dff_B_FxOmnJYt7_1),.dout(w_dff_B_b4tasGne0_1),.clk(gclk));
	jdff dff_B_RQpEWAFG6_1(.din(w_dff_B_b4tasGne0_1),.dout(w_dff_B_RQpEWAFG6_1),.clk(gclk));
	jdff dff_B_udbH2LjQ4_1(.din(w_dff_B_RQpEWAFG6_1),.dout(w_dff_B_udbH2LjQ4_1),.clk(gclk));
	jdff dff_B_e6tXLClc7_1(.din(w_dff_B_udbH2LjQ4_1),.dout(w_dff_B_e6tXLClc7_1),.clk(gclk));
	jdff dff_B_k5wDjoX28_1(.din(w_dff_B_e6tXLClc7_1),.dout(w_dff_B_k5wDjoX28_1),.clk(gclk));
	jdff dff_B_7n3OBNNV4_1(.din(w_dff_B_k5wDjoX28_1),.dout(w_dff_B_7n3OBNNV4_1),.clk(gclk));
	jdff dff_B_AlWaHE5r6_1(.din(w_dff_B_7n3OBNNV4_1),.dout(w_dff_B_AlWaHE5r6_1),.clk(gclk));
	jdff dff_B_MuIFzA4v1_1(.din(w_dff_B_AlWaHE5r6_1),.dout(w_dff_B_MuIFzA4v1_1),.clk(gclk));
	jdff dff_B_xpKQQ4mf8_1(.din(w_dff_B_MuIFzA4v1_1),.dout(w_dff_B_xpKQQ4mf8_1),.clk(gclk));
	jdff dff_B_TSMfxi0V4_1(.din(w_dff_B_xpKQQ4mf8_1),.dout(w_dff_B_TSMfxi0V4_1),.clk(gclk));
	jdff dff_B_3Tyoumh72_1(.din(w_dff_B_TSMfxi0V4_1),.dout(w_dff_B_3Tyoumh72_1),.clk(gclk));
	jdff dff_B_l8S7gwAd0_1(.din(w_dff_B_3Tyoumh72_1),.dout(w_dff_B_l8S7gwAd0_1),.clk(gclk));
	jdff dff_B_teFzx1jm2_1(.din(w_dff_B_l8S7gwAd0_1),.dout(w_dff_B_teFzx1jm2_1),.clk(gclk));
	jdff dff_B_Mb96YJlx9_1(.din(w_dff_B_teFzx1jm2_1),.dout(w_dff_B_Mb96YJlx9_1),.clk(gclk));
	jdff dff_B_8r7Z6t1f5_1(.din(w_dff_B_Mb96YJlx9_1),.dout(w_dff_B_8r7Z6t1f5_1),.clk(gclk));
	jdff dff_B_7Cm8J7323_1(.din(w_dff_B_8r7Z6t1f5_1),.dout(w_dff_B_7Cm8J7323_1),.clk(gclk));
	jdff dff_B_YO0GtC4U2_1(.din(w_dff_B_7Cm8J7323_1),.dout(w_dff_B_YO0GtC4U2_1),.clk(gclk));
	jdff dff_B_L1iFFo4V1_1(.din(w_dff_B_YO0GtC4U2_1),.dout(w_dff_B_L1iFFo4V1_1),.clk(gclk));
	jdff dff_B_DPvSa2gd6_1(.din(w_dff_B_L1iFFo4V1_1),.dout(w_dff_B_DPvSa2gd6_1),.clk(gclk));
	jdff dff_B_NsC6prcU0_1(.din(w_dff_B_DPvSa2gd6_1),.dout(w_dff_B_NsC6prcU0_1),.clk(gclk));
	jdff dff_B_7ROqNocH2_1(.din(w_dff_B_NsC6prcU0_1),.dout(w_dff_B_7ROqNocH2_1),.clk(gclk));
	jdff dff_B_QHokTbzR1_1(.din(w_dff_B_7ROqNocH2_1),.dout(w_dff_B_QHokTbzR1_1),.clk(gclk));
	jdff dff_B_g6Pg8PGz3_1(.din(w_dff_B_QHokTbzR1_1),.dout(w_dff_B_g6Pg8PGz3_1),.clk(gclk));
	jdff dff_B_o02MqCH97_1(.din(n551),.dout(w_dff_B_o02MqCH97_1),.clk(gclk));
	jdff dff_B_rzPZ16kv6_1(.din(w_dff_B_o02MqCH97_1),.dout(w_dff_B_rzPZ16kv6_1),.clk(gclk));
	jdff dff_B_MKEs9oF78_1(.din(w_dff_B_rzPZ16kv6_1),.dout(w_dff_B_MKEs9oF78_1),.clk(gclk));
	jdff dff_B_NeRT2TyM7_1(.din(w_dff_B_MKEs9oF78_1),.dout(w_dff_B_NeRT2TyM7_1),.clk(gclk));
	jdff dff_B_vjBECOxd6_1(.din(w_dff_B_NeRT2TyM7_1),.dout(w_dff_B_vjBECOxd6_1),.clk(gclk));
	jdff dff_B_1i8tbPKA3_1(.din(w_dff_B_vjBECOxd6_1),.dout(w_dff_B_1i8tbPKA3_1),.clk(gclk));
	jdff dff_B_843t3xRY4_1(.din(w_dff_B_1i8tbPKA3_1),.dout(w_dff_B_843t3xRY4_1),.clk(gclk));
	jdff dff_B_bdqLC7vo9_1(.din(w_dff_B_843t3xRY4_1),.dout(w_dff_B_bdqLC7vo9_1),.clk(gclk));
	jdff dff_B_TNcI5eRw5_1(.din(w_dff_B_bdqLC7vo9_1),.dout(w_dff_B_TNcI5eRw5_1),.clk(gclk));
	jdff dff_B_LwTHwz5h1_1(.din(w_dff_B_TNcI5eRw5_1),.dout(w_dff_B_LwTHwz5h1_1),.clk(gclk));
	jdff dff_B_ogKjg4TT7_1(.din(w_dff_B_LwTHwz5h1_1),.dout(w_dff_B_ogKjg4TT7_1),.clk(gclk));
	jdff dff_B_1tnGRLsd5_1(.din(w_dff_B_ogKjg4TT7_1),.dout(w_dff_B_1tnGRLsd5_1),.clk(gclk));
	jdff dff_B_VX77IbmL3_1(.din(w_dff_B_1tnGRLsd5_1),.dout(w_dff_B_VX77IbmL3_1),.clk(gclk));
	jdff dff_B_OYPlSZWi4_1(.din(w_dff_B_VX77IbmL3_1),.dout(w_dff_B_OYPlSZWi4_1),.clk(gclk));
	jdff dff_B_ZyFnTC5A9_1(.din(w_dff_B_OYPlSZWi4_1),.dout(w_dff_B_ZyFnTC5A9_1),.clk(gclk));
	jdff dff_B_Bq9AfCGp8_1(.din(w_dff_B_ZyFnTC5A9_1),.dout(w_dff_B_Bq9AfCGp8_1),.clk(gclk));
	jdff dff_B_FBymBW7n1_1(.din(w_dff_B_Bq9AfCGp8_1),.dout(w_dff_B_FBymBW7n1_1),.clk(gclk));
	jdff dff_B_MBqbtgjv8_1(.din(w_dff_B_FBymBW7n1_1),.dout(w_dff_B_MBqbtgjv8_1),.clk(gclk));
	jdff dff_B_atvdlYe82_1(.din(w_dff_B_MBqbtgjv8_1),.dout(w_dff_B_atvdlYe82_1),.clk(gclk));
	jdff dff_B_wuJiLk3f0_1(.din(w_dff_B_atvdlYe82_1),.dout(w_dff_B_wuJiLk3f0_1),.clk(gclk));
	jdff dff_B_f8wiba432_1(.din(w_dff_B_wuJiLk3f0_1),.dout(w_dff_B_f8wiba432_1),.clk(gclk));
	jdff dff_B_iarYdNOs8_1(.din(w_dff_B_f8wiba432_1),.dout(w_dff_B_iarYdNOs8_1),.clk(gclk));
	jdff dff_B_SUNnvvs75_1(.din(w_dff_B_iarYdNOs8_1),.dout(w_dff_B_SUNnvvs75_1),.clk(gclk));
	jdff dff_B_p8pivOpx2_1(.din(w_dff_B_SUNnvvs75_1),.dout(w_dff_B_p8pivOpx2_1),.clk(gclk));
	jdff dff_B_WrnvBMAh0_1(.din(w_dff_B_p8pivOpx2_1),.dout(w_dff_B_WrnvBMAh0_1),.clk(gclk));
	jdff dff_B_OMVFAJ2a6_1(.din(w_dff_B_WrnvBMAh0_1),.dout(w_dff_B_OMVFAJ2a6_1),.clk(gclk));
	jdff dff_B_YElUZzDf9_1(.din(w_dff_B_OMVFAJ2a6_1),.dout(w_dff_B_YElUZzDf9_1),.clk(gclk));
	jdff dff_B_U1mmLwCZ0_1(.din(w_dff_B_YElUZzDf9_1),.dout(w_dff_B_U1mmLwCZ0_1),.clk(gclk));
	jdff dff_B_4oTRfwQr8_1(.din(w_dff_B_U1mmLwCZ0_1),.dout(w_dff_B_4oTRfwQr8_1),.clk(gclk));
	jdff dff_B_dKRgVAHZ8_1(.din(w_dff_B_4oTRfwQr8_1),.dout(w_dff_B_dKRgVAHZ8_1),.clk(gclk));
	jdff dff_B_UrxQXydp3_1(.din(w_dff_B_dKRgVAHZ8_1),.dout(w_dff_B_UrxQXydp3_1),.clk(gclk));
	jdff dff_B_5wtEYjLL2_1(.din(w_dff_B_UrxQXydp3_1),.dout(w_dff_B_5wtEYjLL2_1),.clk(gclk));
	jdff dff_B_4lb9XoRh5_1(.din(w_dff_B_5wtEYjLL2_1),.dout(w_dff_B_4lb9XoRh5_1),.clk(gclk));
	jdff dff_B_I9nJ9Bc26_1(.din(w_dff_B_4lb9XoRh5_1),.dout(w_dff_B_I9nJ9Bc26_1),.clk(gclk));
	jdff dff_B_ba7yHDor7_1(.din(n637),.dout(w_dff_B_ba7yHDor7_1),.clk(gclk));
	jdff dff_B_1v9PejCt4_1(.din(w_dff_B_ba7yHDor7_1),.dout(w_dff_B_1v9PejCt4_1),.clk(gclk));
	jdff dff_B_E6K7aPBy9_1(.din(w_dff_B_1v9PejCt4_1),.dout(w_dff_B_E6K7aPBy9_1),.clk(gclk));
	jdff dff_B_kjU0WIxU8_1(.din(w_dff_B_E6K7aPBy9_1),.dout(w_dff_B_kjU0WIxU8_1),.clk(gclk));
	jdff dff_B_m5VZ61L67_1(.din(w_dff_B_kjU0WIxU8_1),.dout(w_dff_B_m5VZ61L67_1),.clk(gclk));
	jdff dff_B_hoJsCj2k7_1(.din(w_dff_B_m5VZ61L67_1),.dout(w_dff_B_hoJsCj2k7_1),.clk(gclk));
	jdff dff_B_YNt5KqTj9_1(.din(w_dff_B_hoJsCj2k7_1),.dout(w_dff_B_YNt5KqTj9_1),.clk(gclk));
	jdff dff_B_KrtjcLqM4_1(.din(w_dff_B_YNt5KqTj9_1),.dout(w_dff_B_KrtjcLqM4_1),.clk(gclk));
	jdff dff_B_cjyca7w44_1(.din(w_dff_B_KrtjcLqM4_1),.dout(w_dff_B_cjyca7w44_1),.clk(gclk));
	jdff dff_B_LMGnYrWV7_1(.din(w_dff_B_cjyca7w44_1),.dout(w_dff_B_LMGnYrWV7_1),.clk(gclk));
	jdff dff_B_D0n8gG373_1(.din(w_dff_B_LMGnYrWV7_1),.dout(w_dff_B_D0n8gG373_1),.clk(gclk));
	jdff dff_B_xustH9JN0_1(.din(w_dff_B_D0n8gG373_1),.dout(w_dff_B_xustH9JN0_1),.clk(gclk));
	jdff dff_B_AdciMGAg0_1(.din(w_dff_B_xustH9JN0_1),.dout(w_dff_B_AdciMGAg0_1),.clk(gclk));
	jdff dff_B_YgVZMix71_1(.din(w_dff_B_AdciMGAg0_1),.dout(w_dff_B_YgVZMix71_1),.clk(gclk));
	jdff dff_B_2x8z9CsQ3_1(.din(w_dff_B_YgVZMix71_1),.dout(w_dff_B_2x8z9CsQ3_1),.clk(gclk));
	jdff dff_B_3R5MpDEX5_1(.din(w_dff_B_2x8z9CsQ3_1),.dout(w_dff_B_3R5MpDEX5_1),.clk(gclk));
	jdff dff_B_MAphkkXz6_1(.din(w_dff_B_3R5MpDEX5_1),.dout(w_dff_B_MAphkkXz6_1),.clk(gclk));
	jdff dff_B_tBGD9mXy0_1(.din(w_dff_B_MAphkkXz6_1),.dout(w_dff_B_tBGD9mXy0_1),.clk(gclk));
	jdff dff_B_nxywcEQT7_1(.din(w_dff_B_tBGD9mXy0_1),.dout(w_dff_B_nxywcEQT7_1),.clk(gclk));
	jdff dff_B_43c16sot3_1(.din(w_dff_B_nxywcEQT7_1),.dout(w_dff_B_43c16sot3_1),.clk(gclk));
	jdff dff_B_YOI6Kdlw6_1(.din(w_dff_B_43c16sot3_1),.dout(w_dff_B_YOI6Kdlw6_1),.clk(gclk));
	jdff dff_B_4vog6DFp5_1(.din(w_dff_B_YOI6Kdlw6_1),.dout(w_dff_B_4vog6DFp5_1),.clk(gclk));
	jdff dff_B_HLRyeS8Z6_1(.din(w_dff_B_4vog6DFp5_1),.dout(w_dff_B_HLRyeS8Z6_1),.clk(gclk));
	jdff dff_B_YPLgVBAv6_1(.din(w_dff_B_HLRyeS8Z6_1),.dout(w_dff_B_YPLgVBAv6_1),.clk(gclk));
	jdff dff_B_EnAH4Js65_1(.din(w_dff_B_YPLgVBAv6_1),.dout(w_dff_B_EnAH4Js65_1),.clk(gclk));
	jdff dff_B_xvFx4mJ55_1(.din(w_dff_B_EnAH4Js65_1),.dout(w_dff_B_xvFx4mJ55_1),.clk(gclk));
	jdff dff_B_TTSwfGcV1_1(.din(w_dff_B_xvFx4mJ55_1),.dout(w_dff_B_TTSwfGcV1_1),.clk(gclk));
	jdff dff_B_5a35RJUv5_1(.din(w_dff_B_TTSwfGcV1_1),.dout(w_dff_B_5a35RJUv5_1),.clk(gclk));
	jdff dff_B_IkHbgszW1_1(.din(w_dff_B_5a35RJUv5_1),.dout(w_dff_B_IkHbgszW1_1),.clk(gclk));
	jdff dff_B_OHLiR9ce0_1(.din(w_dff_B_IkHbgszW1_1),.dout(w_dff_B_OHLiR9ce0_1),.clk(gclk));
	jdff dff_B_aQJSDXwv1_1(.din(w_dff_B_OHLiR9ce0_1),.dout(w_dff_B_aQJSDXwv1_1),.clk(gclk));
	jdff dff_B_KEclRy8v4_1(.din(w_dff_B_aQJSDXwv1_1),.dout(w_dff_B_KEclRy8v4_1),.clk(gclk));
	jdff dff_B_J6hTIKWU6_1(.din(w_dff_B_KEclRy8v4_1),.dout(w_dff_B_J6hTIKWU6_1),.clk(gclk));
	jdff dff_B_1xGOBdgR8_1(.din(w_dff_B_J6hTIKWU6_1),.dout(w_dff_B_1xGOBdgR8_1),.clk(gclk));
	jdff dff_B_4I22MR9j5_1(.din(w_dff_B_1xGOBdgR8_1),.dout(w_dff_B_4I22MR9j5_1),.clk(gclk));
	jdff dff_B_l9Znp2i90_1(.din(w_dff_B_4I22MR9j5_1),.dout(w_dff_B_l9Znp2i90_1),.clk(gclk));
	jdff dff_B_fX6XFwfv2_1(.din(w_dff_B_l9Znp2i90_1),.dout(w_dff_B_fX6XFwfv2_1),.clk(gclk));
	jdff dff_B_bhERwpZM9_1(.din(n730),.dout(w_dff_B_bhERwpZM9_1),.clk(gclk));
	jdff dff_B_vounQEKF0_1(.din(w_dff_B_bhERwpZM9_1),.dout(w_dff_B_vounQEKF0_1),.clk(gclk));
	jdff dff_B_iEe7ZKqG0_1(.din(w_dff_B_vounQEKF0_1),.dout(w_dff_B_iEe7ZKqG0_1),.clk(gclk));
	jdff dff_B_E0LBWgmp0_1(.din(w_dff_B_iEe7ZKqG0_1),.dout(w_dff_B_E0LBWgmp0_1),.clk(gclk));
	jdff dff_B_fckmYLXb9_1(.din(w_dff_B_E0LBWgmp0_1),.dout(w_dff_B_fckmYLXb9_1),.clk(gclk));
	jdff dff_B_ojD4jv0Q0_1(.din(w_dff_B_fckmYLXb9_1),.dout(w_dff_B_ojD4jv0Q0_1),.clk(gclk));
	jdff dff_B_0lII4XEZ5_1(.din(w_dff_B_ojD4jv0Q0_1),.dout(w_dff_B_0lII4XEZ5_1),.clk(gclk));
	jdff dff_B_1yEjaGtF8_1(.din(w_dff_B_0lII4XEZ5_1),.dout(w_dff_B_1yEjaGtF8_1),.clk(gclk));
	jdff dff_B_16CiTP473_1(.din(w_dff_B_1yEjaGtF8_1),.dout(w_dff_B_16CiTP473_1),.clk(gclk));
	jdff dff_B_GPpO06U95_1(.din(w_dff_B_16CiTP473_1),.dout(w_dff_B_GPpO06U95_1),.clk(gclk));
	jdff dff_B_ywCLCs4H4_1(.din(w_dff_B_GPpO06U95_1),.dout(w_dff_B_ywCLCs4H4_1),.clk(gclk));
	jdff dff_B_cd6ipKFb5_1(.din(w_dff_B_ywCLCs4H4_1),.dout(w_dff_B_cd6ipKFb5_1),.clk(gclk));
	jdff dff_B_zxKrJ2Hg1_1(.din(w_dff_B_cd6ipKFb5_1),.dout(w_dff_B_zxKrJ2Hg1_1),.clk(gclk));
	jdff dff_B_4yU7EuX57_1(.din(w_dff_B_zxKrJ2Hg1_1),.dout(w_dff_B_4yU7EuX57_1),.clk(gclk));
	jdff dff_B_TP0usAbO3_1(.din(w_dff_B_4yU7EuX57_1),.dout(w_dff_B_TP0usAbO3_1),.clk(gclk));
	jdff dff_B_sAXTRqGj2_1(.din(w_dff_B_TP0usAbO3_1),.dout(w_dff_B_sAXTRqGj2_1),.clk(gclk));
	jdff dff_B_5ZVIeCy01_1(.din(w_dff_B_sAXTRqGj2_1),.dout(w_dff_B_5ZVIeCy01_1),.clk(gclk));
	jdff dff_B_gKeN94ss9_1(.din(w_dff_B_5ZVIeCy01_1),.dout(w_dff_B_gKeN94ss9_1),.clk(gclk));
	jdff dff_B_mYQ91xFU0_1(.din(w_dff_B_gKeN94ss9_1),.dout(w_dff_B_mYQ91xFU0_1),.clk(gclk));
	jdff dff_B_dqyaHDPz6_1(.din(w_dff_B_mYQ91xFU0_1),.dout(w_dff_B_dqyaHDPz6_1),.clk(gclk));
	jdff dff_B_83rQTowt2_1(.din(w_dff_B_dqyaHDPz6_1),.dout(w_dff_B_83rQTowt2_1),.clk(gclk));
	jdff dff_B_gGVYeCIU3_1(.din(w_dff_B_83rQTowt2_1),.dout(w_dff_B_gGVYeCIU3_1),.clk(gclk));
	jdff dff_B_qegBv0gk7_1(.din(w_dff_B_gGVYeCIU3_1),.dout(w_dff_B_qegBv0gk7_1),.clk(gclk));
	jdff dff_B_ljCYe4Mi5_1(.din(w_dff_B_qegBv0gk7_1),.dout(w_dff_B_ljCYe4Mi5_1),.clk(gclk));
	jdff dff_B_eERNXww16_1(.din(w_dff_B_ljCYe4Mi5_1),.dout(w_dff_B_eERNXww16_1),.clk(gclk));
	jdff dff_B_1j0PqywI6_1(.din(w_dff_B_eERNXww16_1),.dout(w_dff_B_1j0PqywI6_1),.clk(gclk));
	jdff dff_B_Fp4hZQj24_1(.din(w_dff_B_1j0PqywI6_1),.dout(w_dff_B_Fp4hZQj24_1),.clk(gclk));
	jdff dff_B_Bzd4Gd4G7_1(.din(w_dff_B_Fp4hZQj24_1),.dout(w_dff_B_Bzd4Gd4G7_1),.clk(gclk));
	jdff dff_B_IOkKtf9i2_1(.din(w_dff_B_Bzd4Gd4G7_1),.dout(w_dff_B_IOkKtf9i2_1),.clk(gclk));
	jdff dff_B_I0WggfyD7_1(.din(w_dff_B_IOkKtf9i2_1),.dout(w_dff_B_I0WggfyD7_1),.clk(gclk));
	jdff dff_B_fonbVM4p5_1(.din(w_dff_B_I0WggfyD7_1),.dout(w_dff_B_fonbVM4p5_1),.clk(gclk));
	jdff dff_B_vaq0t36y3_1(.din(w_dff_B_fonbVM4p5_1),.dout(w_dff_B_vaq0t36y3_1),.clk(gclk));
	jdff dff_B_gorOyYwL1_1(.din(w_dff_B_vaq0t36y3_1),.dout(w_dff_B_gorOyYwL1_1),.clk(gclk));
	jdff dff_B_9aONanXf9_1(.din(w_dff_B_gorOyYwL1_1),.dout(w_dff_B_9aONanXf9_1),.clk(gclk));
	jdff dff_B_VfrXnsV62_1(.din(w_dff_B_9aONanXf9_1),.dout(w_dff_B_VfrXnsV62_1),.clk(gclk));
	jdff dff_B_Qvl9bDzk3_1(.din(w_dff_B_VfrXnsV62_1),.dout(w_dff_B_Qvl9bDzk3_1),.clk(gclk));
	jdff dff_B_A2DRuLiV4_1(.din(w_dff_B_Qvl9bDzk3_1),.dout(w_dff_B_A2DRuLiV4_1),.clk(gclk));
	jdff dff_B_pjxF3ZmG0_1(.din(w_dff_B_A2DRuLiV4_1),.dout(w_dff_B_pjxF3ZmG0_1),.clk(gclk));
	jdff dff_B_pCPX82E15_1(.din(w_dff_B_pjxF3ZmG0_1),.dout(w_dff_B_pCPX82E15_1),.clk(gclk));
	jdff dff_B_P2cfAhMG6_1(.din(w_dff_B_pCPX82E15_1),.dout(w_dff_B_P2cfAhMG6_1),.clk(gclk));
	jdff dff_B_EcYzZ6w71_1(.din(n830),.dout(w_dff_B_EcYzZ6w71_1),.clk(gclk));
	jdff dff_B_wIr2XIFU7_1(.din(w_dff_B_EcYzZ6w71_1),.dout(w_dff_B_wIr2XIFU7_1),.clk(gclk));
	jdff dff_B_furpVV9k1_1(.din(w_dff_B_wIr2XIFU7_1),.dout(w_dff_B_furpVV9k1_1),.clk(gclk));
	jdff dff_B_QvHf1xwY0_1(.din(w_dff_B_furpVV9k1_1),.dout(w_dff_B_QvHf1xwY0_1),.clk(gclk));
	jdff dff_B_o4u3vI5k6_1(.din(w_dff_B_QvHf1xwY0_1),.dout(w_dff_B_o4u3vI5k6_1),.clk(gclk));
	jdff dff_B_kHPkxqTA9_1(.din(w_dff_B_o4u3vI5k6_1),.dout(w_dff_B_kHPkxqTA9_1),.clk(gclk));
	jdff dff_B_obd657vg8_1(.din(w_dff_B_kHPkxqTA9_1),.dout(w_dff_B_obd657vg8_1),.clk(gclk));
	jdff dff_B_33mIoTbk8_1(.din(w_dff_B_obd657vg8_1),.dout(w_dff_B_33mIoTbk8_1),.clk(gclk));
	jdff dff_B_yxBmnghK9_1(.din(w_dff_B_33mIoTbk8_1),.dout(w_dff_B_yxBmnghK9_1),.clk(gclk));
	jdff dff_B_eXX13Pqf2_1(.din(w_dff_B_yxBmnghK9_1),.dout(w_dff_B_eXX13Pqf2_1),.clk(gclk));
	jdff dff_B_0ueVHSbU3_1(.din(w_dff_B_eXX13Pqf2_1),.dout(w_dff_B_0ueVHSbU3_1),.clk(gclk));
	jdff dff_B_k8P4wljZ5_1(.din(w_dff_B_0ueVHSbU3_1),.dout(w_dff_B_k8P4wljZ5_1),.clk(gclk));
	jdff dff_B_xLEamzwr9_1(.din(w_dff_B_k8P4wljZ5_1),.dout(w_dff_B_xLEamzwr9_1),.clk(gclk));
	jdff dff_B_zURI3Hdu6_1(.din(w_dff_B_xLEamzwr9_1),.dout(w_dff_B_zURI3Hdu6_1),.clk(gclk));
	jdff dff_B_kYeKGal02_1(.din(w_dff_B_zURI3Hdu6_1),.dout(w_dff_B_kYeKGal02_1),.clk(gclk));
	jdff dff_B_wnEDff3J9_1(.din(w_dff_B_kYeKGal02_1),.dout(w_dff_B_wnEDff3J9_1),.clk(gclk));
	jdff dff_B_vU0e0Ijl7_1(.din(w_dff_B_wnEDff3J9_1),.dout(w_dff_B_vU0e0Ijl7_1),.clk(gclk));
	jdff dff_B_TjK5C9pn3_1(.din(w_dff_B_vU0e0Ijl7_1),.dout(w_dff_B_TjK5C9pn3_1),.clk(gclk));
	jdff dff_B_leCVotMu8_1(.din(w_dff_B_TjK5C9pn3_1),.dout(w_dff_B_leCVotMu8_1),.clk(gclk));
	jdff dff_B_Ocyxqbgr9_1(.din(w_dff_B_leCVotMu8_1),.dout(w_dff_B_Ocyxqbgr9_1),.clk(gclk));
	jdff dff_B_3u7UaqNw8_1(.din(w_dff_B_Ocyxqbgr9_1),.dout(w_dff_B_3u7UaqNw8_1),.clk(gclk));
	jdff dff_B_2SKH4sBb5_1(.din(w_dff_B_3u7UaqNw8_1),.dout(w_dff_B_2SKH4sBb5_1),.clk(gclk));
	jdff dff_B_xPcaFZLU2_1(.din(w_dff_B_2SKH4sBb5_1),.dout(w_dff_B_xPcaFZLU2_1),.clk(gclk));
	jdff dff_B_8S3jPgSq7_1(.din(w_dff_B_xPcaFZLU2_1),.dout(w_dff_B_8S3jPgSq7_1),.clk(gclk));
	jdff dff_B_vGd5woqt0_1(.din(w_dff_B_8S3jPgSq7_1),.dout(w_dff_B_vGd5woqt0_1),.clk(gclk));
	jdff dff_B_ZTvQ8cOR8_1(.din(w_dff_B_vGd5woqt0_1),.dout(w_dff_B_ZTvQ8cOR8_1),.clk(gclk));
	jdff dff_B_PirkwQWd4_1(.din(w_dff_B_ZTvQ8cOR8_1),.dout(w_dff_B_PirkwQWd4_1),.clk(gclk));
	jdff dff_B_jpzYNZOM2_1(.din(w_dff_B_PirkwQWd4_1),.dout(w_dff_B_jpzYNZOM2_1),.clk(gclk));
	jdff dff_B_Lg15YytX8_1(.din(w_dff_B_jpzYNZOM2_1),.dout(w_dff_B_Lg15YytX8_1),.clk(gclk));
	jdff dff_B_C37td1dx7_1(.din(w_dff_B_Lg15YytX8_1),.dout(w_dff_B_C37td1dx7_1),.clk(gclk));
	jdff dff_B_L6WtZiIo4_1(.din(w_dff_B_C37td1dx7_1),.dout(w_dff_B_L6WtZiIo4_1),.clk(gclk));
	jdff dff_B_n3S53RUV4_1(.din(w_dff_B_L6WtZiIo4_1),.dout(w_dff_B_n3S53RUV4_1),.clk(gclk));
	jdff dff_B_hupLYL7c3_1(.din(w_dff_B_n3S53RUV4_1),.dout(w_dff_B_hupLYL7c3_1),.clk(gclk));
	jdff dff_B_gmBAj38L4_1(.din(w_dff_B_hupLYL7c3_1),.dout(w_dff_B_gmBAj38L4_1),.clk(gclk));
	jdff dff_B_qLJbvFUF3_1(.din(w_dff_B_gmBAj38L4_1),.dout(w_dff_B_qLJbvFUF3_1),.clk(gclk));
	jdff dff_B_lMpFMA492_1(.din(w_dff_B_qLJbvFUF3_1),.dout(w_dff_B_lMpFMA492_1),.clk(gclk));
	jdff dff_B_DMuZ9GNp9_1(.din(w_dff_B_lMpFMA492_1),.dout(w_dff_B_DMuZ9GNp9_1),.clk(gclk));
	jdff dff_B_eN08a2vV8_1(.din(w_dff_B_DMuZ9GNp9_1),.dout(w_dff_B_eN08a2vV8_1),.clk(gclk));
	jdff dff_B_TZVngQF69_1(.din(w_dff_B_eN08a2vV8_1),.dout(w_dff_B_TZVngQF69_1),.clk(gclk));
	jdff dff_B_5aFT5H7H8_1(.din(w_dff_B_TZVngQF69_1),.dout(w_dff_B_5aFT5H7H8_1),.clk(gclk));
	jdff dff_B_AH6MrSp94_1(.din(w_dff_B_5aFT5H7H8_1),.dout(w_dff_B_AH6MrSp94_1),.clk(gclk));
	jdff dff_B_fxHsrPUf6_1(.din(w_dff_B_AH6MrSp94_1),.dout(w_dff_B_fxHsrPUf6_1),.clk(gclk));
	jdff dff_B_vYOXfILh7_1(.din(w_dff_B_fxHsrPUf6_1),.dout(w_dff_B_vYOXfILh7_1),.clk(gclk));
	jdff dff_B_fMoeLlFX7_0(.din(n1327),.dout(w_dff_B_fMoeLlFX7_0),.clk(gclk));
	jdff dff_B_sbFeo1EI5_1(.din(n1842),.dout(w_dff_B_sbFeo1EI5_1),.clk(gclk));
	jdff dff_B_2INyUXAH4_1(.din(w_dff_B_sbFeo1EI5_1),.dout(w_dff_B_2INyUXAH4_1),.clk(gclk));
	jdff dff_B_zTW8EAQk9_1(.din(w_dff_B_2INyUXAH4_1),.dout(w_dff_B_zTW8EAQk9_1),.clk(gclk));
	jdff dff_B_kcolGlWG7_1(.din(w_dff_B_zTW8EAQk9_1),.dout(w_dff_B_kcolGlWG7_1),.clk(gclk));
	jdff dff_B_bmKLUEvh2_1(.din(w_dff_B_kcolGlWG7_1),.dout(w_dff_B_bmKLUEvh2_1),.clk(gclk));
	jdff dff_B_RwqUbpFi6_1(.din(w_dff_B_bmKLUEvh2_1),.dout(w_dff_B_RwqUbpFi6_1),.clk(gclk));
	jdff dff_B_ReuhXnQ20_1(.din(w_dff_B_RwqUbpFi6_1),.dout(w_dff_B_ReuhXnQ20_1),.clk(gclk));
	jdff dff_B_pAVLRkq43_1(.din(w_dff_B_ReuhXnQ20_1),.dout(w_dff_B_pAVLRkq43_1),.clk(gclk));
	jdff dff_B_pihkHoxr6_1(.din(w_dff_B_pAVLRkq43_1),.dout(w_dff_B_pihkHoxr6_1),.clk(gclk));
	jdff dff_B_6xtnLTau1_1(.din(w_dff_B_pihkHoxr6_1),.dout(w_dff_B_6xtnLTau1_1),.clk(gclk));
	jdff dff_B_bna7xfMG2_1(.din(w_dff_B_6xtnLTau1_1),.dout(w_dff_B_bna7xfMG2_1),.clk(gclk));
	jdff dff_B_qeId6v1Q8_1(.din(w_dff_B_bna7xfMG2_1),.dout(w_dff_B_qeId6v1Q8_1),.clk(gclk));
	jdff dff_B_tEIzL6Si8_1(.din(w_dff_B_qeId6v1Q8_1),.dout(w_dff_B_tEIzL6Si8_1),.clk(gclk));
	jdff dff_B_hQicRh9g9_0(.din(n1850),.dout(w_dff_B_hQicRh9g9_0),.clk(gclk));
	jdff dff_B_Zsh8d9J27_0(.din(w_dff_B_hQicRh9g9_0),.dout(w_dff_B_Zsh8d9J27_0),.clk(gclk));
	jdff dff_B_EJ1uPLOd7_0(.din(w_dff_B_Zsh8d9J27_0),.dout(w_dff_B_EJ1uPLOd7_0),.clk(gclk));
	jdff dff_B_49lDF8be5_0(.din(w_dff_B_EJ1uPLOd7_0),.dout(w_dff_B_49lDF8be5_0),.clk(gclk));
	jdff dff_B_oubJSXAn0_0(.din(w_dff_B_49lDF8be5_0),.dout(w_dff_B_oubJSXAn0_0),.clk(gclk));
	jdff dff_B_AgpVtZNU5_0(.din(w_dff_B_oubJSXAn0_0),.dout(w_dff_B_AgpVtZNU5_0),.clk(gclk));
	jdff dff_B_aqxE7IaL6_0(.din(w_dff_B_AgpVtZNU5_0),.dout(w_dff_B_aqxE7IaL6_0),.clk(gclk));
	jdff dff_B_z2OGlrf04_0(.din(w_dff_B_aqxE7IaL6_0),.dout(w_dff_B_z2OGlrf04_0),.clk(gclk));
	jdff dff_B_gMnJwXhg9_0(.din(w_dff_B_z2OGlrf04_0),.dout(w_dff_B_gMnJwXhg9_0),.clk(gclk));
	jdff dff_B_MHn6vCaL1_0(.din(w_dff_B_gMnJwXhg9_0),.dout(w_dff_B_MHn6vCaL1_0),.clk(gclk));
	jdff dff_B_lO57ET7m6_0(.din(w_dff_B_MHn6vCaL1_0),.dout(w_dff_B_lO57ET7m6_0),.clk(gclk));
	jdff dff_A_m0JjNuvI8_0(.dout(w_n1849_0[0]),.din(w_dff_A_m0JjNuvI8_0),.clk(gclk));
	jdff dff_A_XyLHhIko8_0(.dout(w_dff_A_m0JjNuvI8_0),.din(w_dff_A_XyLHhIko8_0),.clk(gclk));
	jdff dff_A_YZyxKGH84_0(.dout(w_dff_A_XyLHhIko8_0),.din(w_dff_A_YZyxKGH84_0),.clk(gclk));
	jdff dff_A_zNE32iKI2_0(.dout(w_dff_A_YZyxKGH84_0),.din(w_dff_A_zNE32iKI2_0),.clk(gclk));
	jdff dff_A_J6oD1eTw0_0(.dout(w_dff_A_zNE32iKI2_0),.din(w_dff_A_J6oD1eTw0_0),.clk(gclk));
	jdff dff_A_RzBZ9N197_0(.dout(w_dff_A_J6oD1eTw0_0),.din(w_dff_A_RzBZ9N197_0),.clk(gclk));
	jdff dff_A_PbKFL8IP9_0(.dout(w_dff_A_RzBZ9N197_0),.din(w_dff_A_PbKFL8IP9_0),.clk(gclk));
	jdff dff_A_w5ljE4UP8_0(.dout(w_dff_A_PbKFL8IP9_0),.din(w_dff_A_w5ljE4UP8_0),.clk(gclk));
	jdff dff_A_ldpsVJv72_0(.dout(w_dff_A_w5ljE4UP8_0),.din(w_dff_A_ldpsVJv72_0),.clk(gclk));
	jdff dff_A_BIR0T2Er1_0(.dout(w_dff_A_ldpsVJv72_0),.din(w_dff_A_BIR0T2Er1_0),.clk(gclk));
	jdff dff_A_UOZBiI5q7_0(.dout(w_dff_A_BIR0T2Er1_0),.din(w_dff_A_UOZBiI5q7_0),.clk(gclk));
	jdff dff_A_AfYw5laX3_0(.dout(w_dff_A_UOZBiI5q7_0),.din(w_dff_A_AfYw5laX3_0),.clk(gclk));
	jdff dff_B_tWoZIzdD1_1(.din(n1839),.dout(w_dff_B_tWoZIzdD1_1),.clk(gclk));
	jdff dff_B_l8E1hQ3o8_1(.din(w_dff_B_tWoZIzdD1_1),.dout(w_dff_B_l8E1hQ3o8_1),.clk(gclk));
	jdff dff_B_iz9aTgB08_2(.din(n1838),.dout(w_dff_B_iz9aTgB08_2),.clk(gclk));
	jdff dff_B_bV3ZWcCp4_2(.din(w_dff_B_iz9aTgB08_2),.dout(w_dff_B_bV3ZWcCp4_2),.clk(gclk));
	jdff dff_B_qTkMv25N4_2(.din(w_dff_B_bV3ZWcCp4_2),.dout(w_dff_B_qTkMv25N4_2),.clk(gclk));
	jdff dff_B_qYKJNjHM8_2(.din(w_dff_B_qTkMv25N4_2),.dout(w_dff_B_qYKJNjHM8_2),.clk(gclk));
	jdff dff_B_ZE0PLiXw4_2(.din(w_dff_B_qYKJNjHM8_2),.dout(w_dff_B_ZE0PLiXw4_2),.clk(gclk));
	jdff dff_B_e7JmlJml1_2(.din(w_dff_B_ZE0PLiXw4_2),.dout(w_dff_B_e7JmlJml1_2),.clk(gclk));
	jdff dff_B_pSibLW3N1_2(.din(w_dff_B_e7JmlJml1_2),.dout(w_dff_B_pSibLW3N1_2),.clk(gclk));
	jdff dff_B_Xb5OxJb10_2(.din(w_dff_B_pSibLW3N1_2),.dout(w_dff_B_Xb5OxJb10_2),.clk(gclk));
	jdff dff_B_2fv4WZuu7_2(.din(w_dff_B_Xb5OxJb10_2),.dout(w_dff_B_2fv4WZuu7_2),.clk(gclk));
	jdff dff_B_aU7SC2Mt6_2(.din(w_dff_B_2fv4WZuu7_2),.dout(w_dff_B_aU7SC2Mt6_2),.clk(gclk));
	jdff dff_B_AMl8UHIt8_2(.din(w_dff_B_aU7SC2Mt6_2),.dout(w_dff_B_AMl8UHIt8_2),.clk(gclk));
	jdff dff_B_zqxapdLY1_2(.din(w_dff_B_AMl8UHIt8_2),.dout(w_dff_B_zqxapdLY1_2),.clk(gclk));
	jdff dff_B_r1kE9BxB6_2(.din(w_dff_B_zqxapdLY1_2),.dout(w_dff_B_r1kE9BxB6_2),.clk(gclk));
	jdff dff_B_QatLuJBO0_2(.din(w_dff_B_r1kE9BxB6_2),.dout(w_dff_B_QatLuJBO0_2),.clk(gclk));
	jdff dff_B_xgMpC9re1_2(.din(w_dff_B_QatLuJBO0_2),.dout(w_dff_B_xgMpC9re1_2),.clk(gclk));
	jdff dff_B_4XrfGHGV8_2(.din(w_dff_B_xgMpC9re1_2),.dout(w_dff_B_4XrfGHGV8_2),.clk(gclk));
	jdff dff_B_tBJTXV7x1_2(.din(w_dff_B_4XrfGHGV8_2),.dout(w_dff_B_tBJTXV7x1_2),.clk(gclk));
	jdff dff_B_MR6tEHgC4_2(.din(w_dff_B_tBJTXV7x1_2),.dout(w_dff_B_MR6tEHgC4_2),.clk(gclk));
	jdff dff_B_e34WTH2O3_2(.din(w_dff_B_MR6tEHgC4_2),.dout(w_dff_B_e34WTH2O3_2),.clk(gclk));
	jdff dff_B_hUnFkNs61_2(.din(w_dff_B_e34WTH2O3_2),.dout(w_dff_B_hUnFkNs61_2),.clk(gclk));
	jdff dff_B_RnZXvcQH5_2(.din(w_dff_B_hUnFkNs61_2),.dout(w_dff_B_RnZXvcQH5_2),.clk(gclk));
	jdff dff_B_7ADFwLpP0_2(.din(w_dff_B_RnZXvcQH5_2),.dout(w_dff_B_7ADFwLpP0_2),.clk(gclk));
	jdff dff_B_wXScGgMg6_2(.din(w_dff_B_7ADFwLpP0_2),.dout(w_dff_B_wXScGgMg6_2),.clk(gclk));
	jdff dff_B_A3sTDcJI9_2(.din(w_dff_B_wXScGgMg6_2),.dout(w_dff_B_A3sTDcJI9_2),.clk(gclk));
	jdff dff_B_AUuzRjLB8_2(.din(w_dff_B_A3sTDcJI9_2),.dout(w_dff_B_AUuzRjLB8_2),.clk(gclk));
	jdff dff_B_3LPsbA4d6_2(.din(w_dff_B_AUuzRjLB8_2),.dout(w_dff_B_3LPsbA4d6_2),.clk(gclk));
	jdff dff_B_m28lmXxm5_2(.din(w_dff_B_3LPsbA4d6_2),.dout(w_dff_B_m28lmXxm5_2),.clk(gclk));
	jdff dff_B_vGvo1yPu8_2(.din(w_dff_B_m28lmXxm5_2),.dout(w_dff_B_vGvo1yPu8_2),.clk(gclk));
	jdff dff_B_orcXzQlX1_2(.din(w_dff_B_vGvo1yPu8_2),.dout(w_dff_B_orcXzQlX1_2),.clk(gclk));
	jdff dff_B_TW4Lygyl1_2(.din(w_dff_B_orcXzQlX1_2),.dout(w_dff_B_TW4Lygyl1_2),.clk(gclk));
	jdff dff_B_NehRVWgf9_2(.din(w_dff_B_TW4Lygyl1_2),.dout(w_dff_B_NehRVWgf9_2),.clk(gclk));
	jdff dff_B_k6lnXCH26_2(.din(w_dff_B_NehRVWgf9_2),.dout(w_dff_B_k6lnXCH26_2),.clk(gclk));
	jdff dff_B_mtTvTe6Y9_2(.din(w_dff_B_k6lnXCH26_2),.dout(w_dff_B_mtTvTe6Y9_2),.clk(gclk));
	jdff dff_B_1Qyk3WNZ6_2(.din(w_dff_B_mtTvTe6Y9_2),.dout(w_dff_B_1Qyk3WNZ6_2),.clk(gclk));
	jdff dff_B_CtmDnbP80_2(.din(w_dff_B_1Qyk3WNZ6_2),.dout(w_dff_B_CtmDnbP80_2),.clk(gclk));
	jdff dff_B_3t6dei1P1_2(.din(w_dff_B_CtmDnbP80_2),.dout(w_dff_B_3t6dei1P1_2),.clk(gclk));
	jdff dff_B_7uNCo4D26_2(.din(w_dff_B_3t6dei1P1_2),.dout(w_dff_B_7uNCo4D26_2),.clk(gclk));
	jdff dff_B_T8ejGtNS7_2(.din(w_dff_B_7uNCo4D26_2),.dout(w_dff_B_T8ejGtNS7_2),.clk(gclk));
	jdff dff_B_Yak9Udtk2_2(.din(w_dff_B_T8ejGtNS7_2),.dout(w_dff_B_Yak9Udtk2_2),.clk(gclk));
	jdff dff_B_R0LIlpBN7_2(.din(w_dff_B_Yak9Udtk2_2),.dout(w_dff_B_R0LIlpBN7_2),.clk(gclk));
	jdff dff_B_5SzAzHYS9_2(.din(w_dff_B_R0LIlpBN7_2),.dout(w_dff_B_5SzAzHYS9_2),.clk(gclk));
	jdff dff_B_ICHowvGj6_2(.din(w_dff_B_5SzAzHYS9_2),.dout(w_dff_B_ICHowvGj6_2),.clk(gclk));
	jdff dff_B_J7UtQFDH1_2(.din(w_dff_B_ICHowvGj6_2),.dout(w_dff_B_J7UtQFDH1_2),.clk(gclk));
	jdff dff_B_D6Ik5QjN1_2(.din(w_dff_B_J7UtQFDH1_2),.dout(w_dff_B_D6Ik5QjN1_2),.clk(gclk));
	jdff dff_B_PMAbDxLz8_2(.din(w_dff_B_D6Ik5QjN1_2),.dout(w_dff_B_PMAbDxLz8_2),.clk(gclk));
	jdff dff_B_ImRoXffv4_2(.din(w_dff_B_PMAbDxLz8_2),.dout(w_dff_B_ImRoXffv4_2),.clk(gclk));
	jdff dff_B_Pftahw966_2(.din(w_dff_B_ImRoXffv4_2),.dout(w_dff_B_Pftahw966_2),.clk(gclk));
	jdff dff_B_lG50ej0b4_2(.din(w_dff_B_Pftahw966_2),.dout(w_dff_B_lG50ej0b4_2),.clk(gclk));
	jdff dff_B_r4AF2vQW2_2(.din(w_dff_B_lG50ej0b4_2),.dout(w_dff_B_r4AF2vQW2_2),.clk(gclk));
	jdff dff_B_uBLBvLJo3_2(.din(w_dff_B_r4AF2vQW2_2),.dout(w_dff_B_uBLBvLJo3_2),.clk(gclk));
	jdff dff_B_fOJhEY0Y2_2(.din(w_dff_B_uBLBvLJo3_2),.dout(w_dff_B_fOJhEY0Y2_2),.clk(gclk));
	jdff dff_B_ktcPXAgr7_2(.din(w_dff_B_fOJhEY0Y2_2),.dout(w_dff_B_ktcPXAgr7_2),.clk(gclk));
	jdff dff_B_4OKefqFS1_2(.din(w_dff_B_ktcPXAgr7_2),.dout(w_dff_B_4OKefqFS1_2),.clk(gclk));
	jdff dff_B_mF1Ktk8h2_2(.din(w_dff_B_4OKefqFS1_2),.dout(w_dff_B_mF1Ktk8h2_2),.clk(gclk));
	jdff dff_B_FhwPWVkg5_2(.din(w_dff_B_mF1Ktk8h2_2),.dout(w_dff_B_FhwPWVkg5_2),.clk(gclk));
	jdff dff_B_ZRuRRZd25_2(.din(w_dff_B_FhwPWVkg5_2),.dout(w_dff_B_ZRuRRZd25_2),.clk(gclk));
	jdff dff_B_IgwhY4ht2_2(.din(w_dff_B_ZRuRRZd25_2),.dout(w_dff_B_IgwhY4ht2_2),.clk(gclk));
	jdff dff_B_rgzkUHGt0_2(.din(w_dff_B_IgwhY4ht2_2),.dout(w_dff_B_rgzkUHGt0_2),.clk(gclk));
	jdff dff_B_jAPfrKB49_2(.din(w_dff_B_rgzkUHGt0_2),.dout(w_dff_B_jAPfrKB49_2),.clk(gclk));
	jdff dff_B_g4xoyXVp5_2(.din(w_dff_B_jAPfrKB49_2),.dout(w_dff_B_g4xoyXVp5_2),.clk(gclk));
	jdff dff_B_YAyryhwi7_1(.din(n1845),.dout(w_dff_B_YAyryhwi7_1),.clk(gclk));
	jdff dff_B_n8wgVtZu5_1(.din(w_dff_B_YAyryhwi7_1),.dout(w_dff_B_n8wgVtZu5_1),.clk(gclk));
	jdff dff_B_CEZXvmhg5_1(.din(w_dff_B_n8wgVtZu5_1),.dout(w_dff_B_CEZXvmhg5_1),.clk(gclk));
	jdff dff_B_iE86Ry8q4_1(.din(w_dff_B_CEZXvmhg5_1),.dout(w_dff_B_iE86Ry8q4_1),.clk(gclk));
	jdff dff_B_5Gr5F1uv0_1(.din(w_dff_B_iE86Ry8q4_1),.dout(w_dff_B_5Gr5F1uv0_1),.clk(gclk));
	jdff dff_B_AjkQlkJc1_1(.din(w_dff_B_5Gr5F1uv0_1),.dout(w_dff_B_AjkQlkJc1_1),.clk(gclk));
	jdff dff_B_lVVVOTHN7_1(.din(w_dff_B_AjkQlkJc1_1),.dout(w_dff_B_lVVVOTHN7_1),.clk(gclk));
	jdff dff_B_YjTJqmDs0_1(.din(w_dff_B_lVVVOTHN7_1),.dout(w_dff_B_YjTJqmDs0_1),.clk(gclk));
	jdff dff_B_OztWx61B7_1(.din(w_dff_B_YjTJqmDs0_1),.dout(w_dff_B_OztWx61B7_1),.clk(gclk));
	jdff dff_B_GCPIvll60_1(.din(w_dff_B_OztWx61B7_1),.dout(w_dff_B_GCPIvll60_1),.clk(gclk));
	jdff dff_B_wJhP7oj49_1(.din(w_dff_B_GCPIvll60_1),.dout(w_dff_B_wJhP7oj49_1),.clk(gclk));
	jdff dff_B_EMOiCLTU2_0(.din(n1846),.dout(w_dff_B_EMOiCLTU2_0),.clk(gclk));
	jdff dff_B_VZTT7cji8_0(.din(w_dff_B_EMOiCLTU2_0),.dout(w_dff_B_VZTT7cji8_0),.clk(gclk));
	jdff dff_B_DC8U9q976_0(.din(w_dff_B_VZTT7cji8_0),.dout(w_dff_B_DC8U9q976_0),.clk(gclk));
	jdff dff_B_3YqqsRiB0_0(.din(w_dff_B_DC8U9q976_0),.dout(w_dff_B_3YqqsRiB0_0),.clk(gclk));
	jdff dff_B_t7nv8bQi1_0(.din(w_dff_B_3YqqsRiB0_0),.dout(w_dff_B_t7nv8bQi1_0),.clk(gclk));
	jdff dff_B_I0yUCq319_0(.din(w_dff_B_t7nv8bQi1_0),.dout(w_dff_B_I0yUCq319_0),.clk(gclk));
	jdff dff_B_7Uv01WtP1_0(.din(w_dff_B_I0yUCq319_0),.dout(w_dff_B_7Uv01WtP1_0),.clk(gclk));
	jdff dff_B_LzStQ3BC8_0(.din(w_dff_B_7Uv01WtP1_0),.dout(w_dff_B_LzStQ3BC8_0),.clk(gclk));
	jdff dff_B_WmBNDTAf5_0(.din(w_dff_B_LzStQ3BC8_0),.dout(w_dff_B_WmBNDTAf5_0),.clk(gclk));
	jdff dff_B_4MdSaJGN5_0(.din(w_dff_B_WmBNDTAf5_0),.dout(w_dff_B_4MdSaJGN5_0),.clk(gclk));
	jdff dff_A_fmIwcrek3_1(.dout(w_n1836_0[1]),.din(w_dff_A_fmIwcrek3_1),.clk(gclk));
	jdff dff_A_IdGKqR6F6_1(.dout(w_dff_A_fmIwcrek3_1),.din(w_dff_A_IdGKqR6F6_1),.clk(gclk));
	jdff dff_A_xkn4FbBm7_1(.dout(w_dff_A_IdGKqR6F6_1),.din(w_dff_A_xkn4FbBm7_1),.clk(gclk));
	jdff dff_A_sJ43ChCR0_1(.dout(w_dff_A_xkn4FbBm7_1),.din(w_dff_A_sJ43ChCR0_1),.clk(gclk));
	jdff dff_A_Jnu1htZZ2_1(.dout(w_dff_A_sJ43ChCR0_1),.din(w_dff_A_Jnu1htZZ2_1),.clk(gclk));
	jdff dff_A_2yfFXLks2_1(.dout(w_dff_A_Jnu1htZZ2_1),.din(w_dff_A_2yfFXLks2_1),.clk(gclk));
	jdff dff_A_ewtxhN3X2_1(.dout(w_dff_A_2yfFXLks2_1),.din(w_dff_A_ewtxhN3X2_1),.clk(gclk));
	jdff dff_A_FQo0tz0n9_1(.dout(w_dff_A_ewtxhN3X2_1),.din(w_dff_A_FQo0tz0n9_1),.clk(gclk));
	jdff dff_A_TaYisTDI2_1(.dout(w_dff_A_FQo0tz0n9_1),.din(w_dff_A_TaYisTDI2_1),.clk(gclk));
	jdff dff_A_JC7YBa092_1(.dout(w_dff_A_TaYisTDI2_1),.din(w_dff_A_JC7YBa092_1),.clk(gclk));
	jdff dff_A_TxFnIYqv4_1(.dout(w_dff_A_JC7YBa092_1),.din(w_dff_A_TxFnIYqv4_1),.clk(gclk));
	jdff dff_B_q6Qq8Sg23_1(.din(n1821),.dout(w_dff_B_q6Qq8Sg23_1),.clk(gclk));
	jdff dff_B_Ay8glTj51_1(.din(w_dff_B_q6Qq8Sg23_1),.dout(w_dff_B_Ay8glTj51_1),.clk(gclk));
	jdff dff_B_b8Ma6md70_1(.din(w_dff_B_Ay8glTj51_1),.dout(w_dff_B_b8Ma6md70_1),.clk(gclk));
	jdff dff_B_aQi1gvLr0_1(.din(w_dff_B_b8Ma6md70_1),.dout(w_dff_B_aQi1gvLr0_1),.clk(gclk));
	jdff dff_B_Ldv37RNC9_1(.din(w_dff_B_aQi1gvLr0_1),.dout(w_dff_B_Ldv37RNC9_1),.clk(gclk));
	jdff dff_B_4Nq2UBo37_1(.din(w_dff_B_Ldv37RNC9_1),.dout(w_dff_B_4Nq2UBo37_1),.clk(gclk));
	jdff dff_B_7vTiqso71_1(.din(w_dff_B_4Nq2UBo37_1),.dout(w_dff_B_7vTiqso71_1),.clk(gclk));
	jdff dff_B_gnm77Bmi3_1(.din(w_dff_B_7vTiqso71_1),.dout(w_dff_B_gnm77Bmi3_1),.clk(gclk));
	jdff dff_B_fO3h4D8N1_1(.din(w_dff_B_gnm77Bmi3_1),.dout(w_dff_B_fO3h4D8N1_1),.clk(gclk));
	jdff dff_B_OClDH2tm0_1(.din(w_dff_B_fO3h4D8N1_1),.dout(w_dff_B_OClDH2tm0_1),.clk(gclk));
	jdff dff_B_V4tVImYF3_1(.din(w_dff_B_OClDH2tm0_1),.dout(w_dff_B_V4tVImYF3_1),.clk(gclk));
	jdff dff_B_m15yRGzY6_0(.din(n1822),.dout(w_dff_B_m15yRGzY6_0),.clk(gclk));
	jdff dff_B_UBlVmbjq0_0(.din(w_dff_B_m15yRGzY6_0),.dout(w_dff_B_UBlVmbjq0_0),.clk(gclk));
	jdff dff_B_uNkVxzEa5_0(.din(w_dff_B_UBlVmbjq0_0),.dout(w_dff_B_uNkVxzEa5_0),.clk(gclk));
	jdff dff_B_KJL4lO9v3_0(.din(w_dff_B_uNkVxzEa5_0),.dout(w_dff_B_KJL4lO9v3_0),.clk(gclk));
	jdff dff_B_aPw0MuTd1_0(.din(w_dff_B_KJL4lO9v3_0),.dout(w_dff_B_aPw0MuTd1_0),.clk(gclk));
	jdff dff_B_rcNnLJ2S1_0(.din(w_dff_B_aPw0MuTd1_0),.dout(w_dff_B_rcNnLJ2S1_0),.clk(gclk));
	jdff dff_B_j4djZjDh0_0(.din(w_dff_B_rcNnLJ2S1_0),.dout(w_dff_B_j4djZjDh0_0),.clk(gclk));
	jdff dff_B_82Yeytqs9_0(.din(w_dff_B_j4djZjDh0_0),.dout(w_dff_B_82Yeytqs9_0),.clk(gclk));
	jdff dff_B_qkz65yQF3_0(.din(w_dff_B_82Yeytqs9_0),.dout(w_dff_B_qkz65yQF3_0),.clk(gclk));
	jdff dff_B_k03xV37X7_0(.din(w_dff_B_qkz65yQF3_0),.dout(w_dff_B_k03xV37X7_0),.clk(gclk));
	jdff dff_A_Yy2ZexX11_1(.dout(w_n1817_0[1]),.din(w_dff_A_Yy2ZexX11_1),.clk(gclk));
	jdff dff_A_6sBrAL3t7_1(.dout(w_dff_A_Yy2ZexX11_1),.din(w_dff_A_6sBrAL3t7_1),.clk(gclk));
	jdff dff_A_9BRfZH5s0_1(.dout(w_dff_A_6sBrAL3t7_1),.din(w_dff_A_9BRfZH5s0_1),.clk(gclk));
	jdff dff_A_L9cWyI3p3_1(.dout(w_dff_A_9BRfZH5s0_1),.din(w_dff_A_L9cWyI3p3_1),.clk(gclk));
	jdff dff_A_nIyoYqLH8_1(.dout(w_dff_A_L9cWyI3p3_1),.din(w_dff_A_nIyoYqLH8_1),.clk(gclk));
	jdff dff_A_dQdlcR7G4_1(.dout(w_dff_A_nIyoYqLH8_1),.din(w_dff_A_dQdlcR7G4_1),.clk(gclk));
	jdff dff_A_etzBS0ph8_1(.dout(w_dff_A_dQdlcR7G4_1),.din(w_dff_A_etzBS0ph8_1),.clk(gclk));
	jdff dff_A_b1nMr4uH3_1(.dout(w_dff_A_etzBS0ph8_1),.din(w_dff_A_b1nMr4uH3_1),.clk(gclk));
	jdff dff_A_LTxjtvaL4_1(.dout(w_dff_A_b1nMr4uH3_1),.din(w_dff_A_LTxjtvaL4_1),.clk(gclk));
	jdff dff_A_PfRSPYNF2_1(.dout(w_dff_A_LTxjtvaL4_1),.din(w_dff_A_PfRSPYNF2_1),.clk(gclk));
	jdff dff_A_axlC0KEc6_1(.dout(w_dff_A_PfRSPYNF2_1),.din(w_dff_A_axlC0KEc6_1),.clk(gclk));
	jdff dff_B_kVPEUSYw5_1(.din(n1795),.dout(w_dff_B_kVPEUSYw5_1),.clk(gclk));
	jdff dff_B_5l0iSaGZ3_1(.din(w_dff_B_kVPEUSYw5_1),.dout(w_dff_B_5l0iSaGZ3_1),.clk(gclk));
	jdff dff_B_IIk8IVHM1_1(.din(w_dff_B_5l0iSaGZ3_1),.dout(w_dff_B_IIk8IVHM1_1),.clk(gclk));
	jdff dff_B_OrVwB2EW5_1(.din(w_dff_B_IIk8IVHM1_1),.dout(w_dff_B_OrVwB2EW5_1),.clk(gclk));
	jdff dff_B_jC1WHUIe7_1(.din(w_dff_B_OrVwB2EW5_1),.dout(w_dff_B_jC1WHUIe7_1),.clk(gclk));
	jdff dff_B_JynPFKln8_1(.din(w_dff_B_jC1WHUIe7_1),.dout(w_dff_B_JynPFKln8_1),.clk(gclk));
	jdff dff_B_KvA4F5B44_1(.din(w_dff_B_JynPFKln8_1),.dout(w_dff_B_KvA4F5B44_1),.clk(gclk));
	jdff dff_B_aYfYaXIp1_1(.din(w_dff_B_KvA4F5B44_1),.dout(w_dff_B_aYfYaXIp1_1),.clk(gclk));
	jdff dff_B_1bzdDDi43_1(.din(w_dff_B_aYfYaXIp1_1),.dout(w_dff_B_1bzdDDi43_1),.clk(gclk));
	jdff dff_B_IuZmrOTp9_1(.din(w_dff_B_1bzdDDi43_1),.dout(w_dff_B_IuZmrOTp9_1),.clk(gclk));
	jdff dff_B_2lTowDer4_1(.din(w_dff_B_IuZmrOTp9_1),.dout(w_dff_B_2lTowDer4_1),.clk(gclk));
	jdff dff_B_C8qvizap8_0(.din(n1796),.dout(w_dff_B_C8qvizap8_0),.clk(gclk));
	jdff dff_B_lBnjesKo5_0(.din(w_dff_B_C8qvizap8_0),.dout(w_dff_B_lBnjesKo5_0),.clk(gclk));
	jdff dff_B_jz1RhArz6_0(.din(w_dff_B_lBnjesKo5_0),.dout(w_dff_B_jz1RhArz6_0),.clk(gclk));
	jdff dff_B_CuB6WOtN4_0(.din(w_dff_B_jz1RhArz6_0),.dout(w_dff_B_CuB6WOtN4_0),.clk(gclk));
	jdff dff_B_zjvUSenK3_0(.din(w_dff_B_CuB6WOtN4_0),.dout(w_dff_B_zjvUSenK3_0),.clk(gclk));
	jdff dff_B_23I54xxa7_0(.din(w_dff_B_zjvUSenK3_0),.dout(w_dff_B_23I54xxa7_0),.clk(gclk));
	jdff dff_B_LPvYyFpm3_0(.din(w_dff_B_23I54xxa7_0),.dout(w_dff_B_LPvYyFpm3_0),.clk(gclk));
	jdff dff_B_C3nCA6dU3_0(.din(w_dff_B_LPvYyFpm3_0),.dout(w_dff_B_C3nCA6dU3_0),.clk(gclk));
	jdff dff_B_Y22ZQXVl8_0(.din(w_dff_B_C3nCA6dU3_0),.dout(w_dff_B_Y22ZQXVl8_0),.clk(gclk));
	jdff dff_B_uo9daJrs0_0(.din(w_dff_B_Y22ZQXVl8_0),.dout(w_dff_B_uo9daJrs0_0),.clk(gclk));
	jdff dff_A_1wWc61pi3_1(.dout(w_n1791_0[1]),.din(w_dff_A_1wWc61pi3_1),.clk(gclk));
	jdff dff_A_yQ3s8HxE3_1(.dout(w_dff_A_1wWc61pi3_1),.din(w_dff_A_yQ3s8HxE3_1),.clk(gclk));
	jdff dff_A_bZZlQ63Z6_1(.dout(w_dff_A_yQ3s8HxE3_1),.din(w_dff_A_bZZlQ63Z6_1),.clk(gclk));
	jdff dff_A_sJz3lPCI2_1(.dout(w_dff_A_bZZlQ63Z6_1),.din(w_dff_A_sJz3lPCI2_1),.clk(gclk));
	jdff dff_A_AeVnl6g52_1(.dout(w_dff_A_sJz3lPCI2_1),.din(w_dff_A_AeVnl6g52_1),.clk(gclk));
	jdff dff_A_ujEWTp711_1(.dout(w_dff_A_AeVnl6g52_1),.din(w_dff_A_ujEWTp711_1),.clk(gclk));
	jdff dff_A_CjsMYCwH0_1(.dout(w_dff_A_ujEWTp711_1),.din(w_dff_A_CjsMYCwH0_1),.clk(gclk));
	jdff dff_A_3I90hbjW0_1(.dout(w_dff_A_CjsMYCwH0_1),.din(w_dff_A_3I90hbjW0_1),.clk(gclk));
	jdff dff_A_P6IelWAb2_1(.dout(w_dff_A_3I90hbjW0_1),.din(w_dff_A_P6IelWAb2_1),.clk(gclk));
	jdff dff_A_6NepZbbQ7_1(.dout(w_dff_A_P6IelWAb2_1),.din(w_dff_A_6NepZbbQ7_1),.clk(gclk));
	jdff dff_A_DbyttkQU3_1(.dout(w_dff_A_6NepZbbQ7_1),.din(w_dff_A_DbyttkQU3_1),.clk(gclk));
	jdff dff_B_5IpxAz8Z3_1(.din(n1762),.dout(w_dff_B_5IpxAz8Z3_1),.clk(gclk));
	jdff dff_B_vmnqg6ss9_1(.din(w_dff_B_5IpxAz8Z3_1),.dout(w_dff_B_vmnqg6ss9_1),.clk(gclk));
	jdff dff_B_a0HmcnQt4_1(.din(w_dff_B_vmnqg6ss9_1),.dout(w_dff_B_a0HmcnQt4_1),.clk(gclk));
	jdff dff_B_GDNd8PaH0_1(.din(w_dff_B_a0HmcnQt4_1),.dout(w_dff_B_GDNd8PaH0_1),.clk(gclk));
	jdff dff_B_Dx47z0606_1(.din(w_dff_B_GDNd8PaH0_1),.dout(w_dff_B_Dx47z0606_1),.clk(gclk));
	jdff dff_B_7y7VD2tk1_1(.din(w_dff_B_Dx47z0606_1),.dout(w_dff_B_7y7VD2tk1_1),.clk(gclk));
	jdff dff_B_RhgaHpNV8_1(.din(w_dff_B_7y7VD2tk1_1),.dout(w_dff_B_RhgaHpNV8_1),.clk(gclk));
	jdff dff_B_2eVIsDYU4_1(.din(w_dff_B_RhgaHpNV8_1),.dout(w_dff_B_2eVIsDYU4_1),.clk(gclk));
	jdff dff_B_LpGSaLql7_1(.din(w_dff_B_2eVIsDYU4_1),.dout(w_dff_B_LpGSaLql7_1),.clk(gclk));
	jdff dff_B_B6zPzUqH3_1(.din(w_dff_B_LpGSaLql7_1),.dout(w_dff_B_B6zPzUqH3_1),.clk(gclk));
	jdff dff_B_wn5H5gc59_1(.din(w_dff_B_B6zPzUqH3_1),.dout(w_dff_B_wn5H5gc59_1),.clk(gclk));
	jdff dff_B_SNWo6Qzh0_0(.din(n1763),.dout(w_dff_B_SNWo6Qzh0_0),.clk(gclk));
	jdff dff_B_JCohFOdw7_0(.din(w_dff_B_SNWo6Qzh0_0),.dout(w_dff_B_JCohFOdw7_0),.clk(gclk));
	jdff dff_B_dBnURjkZ9_0(.din(w_dff_B_JCohFOdw7_0),.dout(w_dff_B_dBnURjkZ9_0),.clk(gclk));
	jdff dff_B_KKfS702Q7_0(.din(w_dff_B_dBnURjkZ9_0),.dout(w_dff_B_KKfS702Q7_0),.clk(gclk));
	jdff dff_B_SLl5u2BT3_0(.din(w_dff_B_KKfS702Q7_0),.dout(w_dff_B_SLl5u2BT3_0),.clk(gclk));
	jdff dff_B_HcmqYFwf9_0(.din(w_dff_B_SLl5u2BT3_0),.dout(w_dff_B_HcmqYFwf9_0),.clk(gclk));
	jdff dff_B_6ZEM32JD3_0(.din(w_dff_B_HcmqYFwf9_0),.dout(w_dff_B_6ZEM32JD3_0),.clk(gclk));
	jdff dff_B_2mWIb39J0_0(.din(w_dff_B_6ZEM32JD3_0),.dout(w_dff_B_2mWIb39J0_0),.clk(gclk));
	jdff dff_B_nnnlgVky2_0(.din(w_dff_B_2mWIb39J0_0),.dout(w_dff_B_nnnlgVky2_0),.clk(gclk));
	jdff dff_B_pS6Cq4dI7_0(.din(w_dff_B_nnnlgVky2_0),.dout(w_dff_B_pS6Cq4dI7_0),.clk(gclk));
	jdff dff_A_BL7JtSMX2_1(.dout(w_n1758_0[1]),.din(w_dff_A_BL7JtSMX2_1),.clk(gclk));
	jdff dff_A_gVAvQkw08_1(.dout(w_dff_A_BL7JtSMX2_1),.din(w_dff_A_gVAvQkw08_1),.clk(gclk));
	jdff dff_A_OA5pJVT69_1(.dout(w_dff_A_gVAvQkw08_1),.din(w_dff_A_OA5pJVT69_1),.clk(gclk));
	jdff dff_A_19h8PTCo1_1(.dout(w_dff_A_OA5pJVT69_1),.din(w_dff_A_19h8PTCo1_1),.clk(gclk));
	jdff dff_A_L7S2zJkL2_1(.dout(w_dff_A_19h8PTCo1_1),.din(w_dff_A_L7S2zJkL2_1),.clk(gclk));
	jdff dff_A_0knXNdyO8_1(.dout(w_dff_A_L7S2zJkL2_1),.din(w_dff_A_0knXNdyO8_1),.clk(gclk));
	jdff dff_A_XLhx0YIo9_1(.dout(w_dff_A_0knXNdyO8_1),.din(w_dff_A_XLhx0YIo9_1),.clk(gclk));
	jdff dff_A_DjUE5ZZc0_1(.dout(w_dff_A_XLhx0YIo9_1),.din(w_dff_A_DjUE5ZZc0_1),.clk(gclk));
	jdff dff_A_8xz9VRPK9_1(.dout(w_dff_A_DjUE5ZZc0_1),.din(w_dff_A_8xz9VRPK9_1),.clk(gclk));
	jdff dff_A_mHSJJKXo5_1(.dout(w_dff_A_8xz9VRPK9_1),.din(w_dff_A_mHSJJKXo5_1),.clk(gclk));
	jdff dff_A_RlkqRC6Q9_1(.dout(w_dff_A_mHSJJKXo5_1),.din(w_dff_A_RlkqRC6Q9_1),.clk(gclk));
	jdff dff_B_v6IhuskW6_1(.din(n1722),.dout(w_dff_B_v6IhuskW6_1),.clk(gclk));
	jdff dff_B_63Mcjvni8_1(.din(w_dff_B_v6IhuskW6_1),.dout(w_dff_B_63Mcjvni8_1),.clk(gclk));
	jdff dff_B_wWKuo2wb4_1(.din(w_dff_B_63Mcjvni8_1),.dout(w_dff_B_wWKuo2wb4_1),.clk(gclk));
	jdff dff_B_Bdhejcms1_1(.din(w_dff_B_wWKuo2wb4_1),.dout(w_dff_B_Bdhejcms1_1),.clk(gclk));
	jdff dff_B_E5cBadYg7_1(.din(w_dff_B_Bdhejcms1_1),.dout(w_dff_B_E5cBadYg7_1),.clk(gclk));
	jdff dff_B_kvA1IVVx7_1(.din(w_dff_B_E5cBadYg7_1),.dout(w_dff_B_kvA1IVVx7_1),.clk(gclk));
	jdff dff_B_KTiaSrYS3_1(.din(w_dff_B_kvA1IVVx7_1),.dout(w_dff_B_KTiaSrYS3_1),.clk(gclk));
	jdff dff_B_gdbnzCQD1_1(.din(w_dff_B_KTiaSrYS3_1),.dout(w_dff_B_gdbnzCQD1_1),.clk(gclk));
	jdff dff_B_YncGPHfT1_1(.din(w_dff_B_gdbnzCQD1_1),.dout(w_dff_B_YncGPHfT1_1),.clk(gclk));
	jdff dff_B_g1SETCA08_1(.din(w_dff_B_YncGPHfT1_1),.dout(w_dff_B_g1SETCA08_1),.clk(gclk));
	jdff dff_B_j8qeHvjW3_1(.din(w_dff_B_g1SETCA08_1),.dout(w_dff_B_j8qeHvjW3_1),.clk(gclk));
	jdff dff_B_NMCqCl6C4_0(.din(n1723),.dout(w_dff_B_NMCqCl6C4_0),.clk(gclk));
	jdff dff_B_6NwIBqkQ4_0(.din(w_dff_B_NMCqCl6C4_0),.dout(w_dff_B_6NwIBqkQ4_0),.clk(gclk));
	jdff dff_B_C65pYUIX2_0(.din(w_dff_B_6NwIBqkQ4_0),.dout(w_dff_B_C65pYUIX2_0),.clk(gclk));
	jdff dff_B_VrInQc6Q7_0(.din(w_dff_B_C65pYUIX2_0),.dout(w_dff_B_VrInQc6Q7_0),.clk(gclk));
	jdff dff_B_qAXq7WAD6_0(.din(w_dff_B_VrInQc6Q7_0),.dout(w_dff_B_qAXq7WAD6_0),.clk(gclk));
	jdff dff_B_T8MwLudp5_0(.din(w_dff_B_qAXq7WAD6_0),.dout(w_dff_B_T8MwLudp5_0),.clk(gclk));
	jdff dff_B_dDKNL7hr7_0(.din(w_dff_B_T8MwLudp5_0),.dout(w_dff_B_dDKNL7hr7_0),.clk(gclk));
	jdff dff_B_NYILoQxo0_0(.din(w_dff_B_dDKNL7hr7_0),.dout(w_dff_B_NYILoQxo0_0),.clk(gclk));
	jdff dff_B_plAUKf9m5_0(.din(w_dff_B_NYILoQxo0_0),.dout(w_dff_B_plAUKf9m5_0),.clk(gclk));
	jdff dff_A_JDqsIVPy3_1(.dout(w_n1720_0[1]),.din(w_dff_A_JDqsIVPy3_1),.clk(gclk));
	jdff dff_A_9Rl5Nb2Z0_1(.dout(w_dff_A_JDqsIVPy3_1),.din(w_dff_A_9Rl5Nb2Z0_1),.clk(gclk));
	jdff dff_A_3yhR6Yn71_1(.dout(w_dff_A_9Rl5Nb2Z0_1),.din(w_dff_A_3yhR6Yn71_1),.clk(gclk));
	jdff dff_A_FZKJHNdz8_1(.dout(w_dff_A_3yhR6Yn71_1),.din(w_dff_A_FZKJHNdz8_1),.clk(gclk));
	jdff dff_A_pe6LVOie1_1(.dout(w_dff_A_FZKJHNdz8_1),.din(w_dff_A_pe6LVOie1_1),.clk(gclk));
	jdff dff_A_PRTjnTu04_1(.dout(w_dff_A_pe6LVOie1_1),.din(w_dff_A_PRTjnTu04_1),.clk(gclk));
	jdff dff_A_mwh0BfB78_1(.dout(w_dff_A_PRTjnTu04_1),.din(w_dff_A_mwh0BfB78_1),.clk(gclk));
	jdff dff_A_ho26mdp31_1(.dout(w_dff_A_mwh0BfB78_1),.din(w_dff_A_ho26mdp31_1),.clk(gclk));
	jdff dff_A_G9YDQs7A9_1(.dout(w_dff_A_ho26mdp31_1),.din(w_dff_A_G9YDQs7A9_1),.clk(gclk));
	jdff dff_A_mHhCd8B79_1(.dout(w_dff_A_G9YDQs7A9_1),.din(w_dff_A_mHhCd8B79_1),.clk(gclk));
	jdff dff_B_wn7ZCnbN9_1(.din(n1674),.dout(w_dff_B_wn7ZCnbN9_1),.clk(gclk));
	jdff dff_B_dn4JiUK64_1(.din(w_dff_B_wn7ZCnbN9_1),.dout(w_dff_B_dn4JiUK64_1),.clk(gclk));
	jdff dff_B_VUJCs6ZS0_1(.din(w_dff_B_dn4JiUK64_1),.dout(w_dff_B_VUJCs6ZS0_1),.clk(gclk));
	jdff dff_B_OrD85vZy6_1(.din(w_dff_B_VUJCs6ZS0_1),.dout(w_dff_B_OrD85vZy6_1),.clk(gclk));
	jdff dff_B_zEJMwPul2_1(.din(w_dff_B_OrD85vZy6_1),.dout(w_dff_B_zEJMwPul2_1),.clk(gclk));
	jdff dff_B_OWdu6gAX7_1(.din(w_dff_B_zEJMwPul2_1),.dout(w_dff_B_OWdu6gAX7_1),.clk(gclk));
	jdff dff_B_w5AIDrQX9_1(.din(w_dff_B_OWdu6gAX7_1),.dout(w_dff_B_w5AIDrQX9_1),.clk(gclk));
	jdff dff_B_4mhNrqrI1_1(.din(w_dff_B_w5AIDrQX9_1),.dout(w_dff_B_4mhNrqrI1_1),.clk(gclk));
	jdff dff_B_OK4ySXev2_1(.din(w_dff_B_4mhNrqrI1_1),.dout(w_dff_B_OK4ySXev2_1),.clk(gclk));
	jdff dff_B_J3ei1HvP0_1(.din(w_dff_B_OK4ySXev2_1),.dout(w_dff_B_J3ei1HvP0_1),.clk(gclk));
	jdff dff_B_zqYyVafT0_0(.din(n1675),.dout(w_dff_B_zqYyVafT0_0),.clk(gclk));
	jdff dff_B_yFBrxJni0_0(.din(w_dff_B_zqYyVafT0_0),.dout(w_dff_B_yFBrxJni0_0),.clk(gclk));
	jdff dff_B_UQIfRW0B4_0(.din(w_dff_B_yFBrxJni0_0),.dout(w_dff_B_UQIfRW0B4_0),.clk(gclk));
	jdff dff_B_73QqV5xQ9_0(.din(w_dff_B_UQIfRW0B4_0),.dout(w_dff_B_73QqV5xQ9_0),.clk(gclk));
	jdff dff_B_U7IAGtya2_0(.din(w_dff_B_73QqV5xQ9_0),.dout(w_dff_B_U7IAGtya2_0),.clk(gclk));
	jdff dff_B_T6fUOHGE2_0(.din(w_dff_B_U7IAGtya2_0),.dout(w_dff_B_T6fUOHGE2_0),.clk(gclk));
	jdff dff_B_Qh64Slzd2_0(.din(w_dff_B_T6fUOHGE2_0),.dout(w_dff_B_Qh64Slzd2_0),.clk(gclk));
	jdff dff_B_hwj8yCsY3_0(.din(w_dff_B_Qh64Slzd2_0),.dout(w_dff_B_hwj8yCsY3_0),.clk(gclk));
	jdff dff_A_PEMtf3vg5_1(.dout(w_n1672_0[1]),.din(w_dff_A_PEMtf3vg5_1),.clk(gclk));
	jdff dff_A_Cdu3USMO5_1(.dout(w_dff_A_PEMtf3vg5_1),.din(w_dff_A_Cdu3USMO5_1),.clk(gclk));
	jdff dff_A_zhX2MfbU8_1(.dout(w_dff_A_Cdu3USMO5_1),.din(w_dff_A_zhX2MfbU8_1),.clk(gclk));
	jdff dff_A_LFvGuECz9_1(.dout(w_dff_A_zhX2MfbU8_1),.din(w_dff_A_LFvGuECz9_1),.clk(gclk));
	jdff dff_A_niCj6BqO6_1(.dout(w_dff_A_LFvGuECz9_1),.din(w_dff_A_niCj6BqO6_1),.clk(gclk));
	jdff dff_A_jxK1qrBp5_1(.dout(w_dff_A_niCj6BqO6_1),.din(w_dff_A_jxK1qrBp5_1),.clk(gclk));
	jdff dff_A_eQCJCu5d0_1(.dout(w_dff_A_jxK1qrBp5_1),.din(w_dff_A_eQCJCu5d0_1),.clk(gclk));
	jdff dff_A_uuOsS5Nl6_1(.dout(w_dff_A_eQCJCu5d0_1),.din(w_dff_A_uuOsS5Nl6_1),.clk(gclk));
	jdff dff_A_alqW54nR6_1(.dout(w_dff_A_uuOsS5Nl6_1),.din(w_dff_A_alqW54nR6_1),.clk(gclk));
	jdff dff_B_hDIJRorC0_1(.din(n1619),.dout(w_dff_B_hDIJRorC0_1),.clk(gclk));
	jdff dff_B_XYhI3q5R6_1(.din(w_dff_B_hDIJRorC0_1),.dout(w_dff_B_XYhI3q5R6_1),.clk(gclk));
	jdff dff_B_IT6zoV182_1(.din(w_dff_B_XYhI3q5R6_1),.dout(w_dff_B_IT6zoV182_1),.clk(gclk));
	jdff dff_B_91PgArA15_1(.din(w_dff_B_IT6zoV182_1),.dout(w_dff_B_91PgArA15_1),.clk(gclk));
	jdff dff_B_hREdb58u6_1(.din(w_dff_B_91PgArA15_1),.dout(w_dff_B_hREdb58u6_1),.clk(gclk));
	jdff dff_B_MWc4OmHJ5_1(.din(w_dff_B_hREdb58u6_1),.dout(w_dff_B_MWc4OmHJ5_1),.clk(gclk));
	jdff dff_B_rK8WkAaj8_1(.din(w_dff_B_MWc4OmHJ5_1),.dout(w_dff_B_rK8WkAaj8_1),.clk(gclk));
	jdff dff_B_BN5B8V2h3_1(.din(w_dff_B_rK8WkAaj8_1),.dout(w_dff_B_BN5B8V2h3_1),.clk(gclk));
	jdff dff_B_QPdpzU6K2_1(.din(w_dff_B_BN5B8V2h3_1),.dout(w_dff_B_QPdpzU6K2_1),.clk(gclk));
	jdff dff_B_LL8oMdvo3_1(.din(w_dff_B_QPdpzU6K2_1),.dout(w_dff_B_LL8oMdvo3_1),.clk(gclk));
	jdff dff_B_IYlB5aSd1_0(.din(n1620),.dout(w_dff_B_IYlB5aSd1_0),.clk(gclk));
	jdff dff_B_ZTaSJ6TW1_0(.din(w_dff_B_IYlB5aSd1_0),.dout(w_dff_B_ZTaSJ6TW1_0),.clk(gclk));
	jdff dff_B_jdmB6ANR4_0(.din(w_dff_B_ZTaSJ6TW1_0),.dout(w_dff_B_jdmB6ANR4_0),.clk(gclk));
	jdff dff_B_3PQFhNu23_0(.din(w_dff_B_jdmB6ANR4_0),.dout(w_dff_B_3PQFhNu23_0),.clk(gclk));
	jdff dff_B_Y0oZyQIu9_0(.din(w_dff_B_3PQFhNu23_0),.dout(w_dff_B_Y0oZyQIu9_0),.clk(gclk));
	jdff dff_B_N3LBxeXa8_0(.din(w_dff_B_Y0oZyQIu9_0),.dout(w_dff_B_N3LBxeXa8_0),.clk(gclk));
	jdff dff_B_YGbr3H580_0(.din(w_dff_B_N3LBxeXa8_0),.dout(w_dff_B_YGbr3H580_0),.clk(gclk));
	jdff dff_B_UtgNrEWs9_0(.din(w_dff_B_YGbr3H580_0),.dout(w_dff_B_UtgNrEWs9_0),.clk(gclk));
	jdff dff_A_vqWjPbkR0_1(.dout(w_n1617_0[1]),.din(w_dff_A_vqWjPbkR0_1),.clk(gclk));
	jdff dff_A_fQ4eruGN5_1(.dout(w_dff_A_vqWjPbkR0_1),.din(w_dff_A_fQ4eruGN5_1),.clk(gclk));
	jdff dff_A_5M2X4v0J2_1(.dout(w_dff_A_fQ4eruGN5_1),.din(w_dff_A_5M2X4v0J2_1),.clk(gclk));
	jdff dff_A_2OamhUUX4_1(.dout(w_dff_A_5M2X4v0J2_1),.din(w_dff_A_2OamhUUX4_1),.clk(gclk));
	jdff dff_A_iwFPN9Lb6_1(.dout(w_dff_A_2OamhUUX4_1),.din(w_dff_A_iwFPN9Lb6_1),.clk(gclk));
	jdff dff_A_OHdBHNXF9_1(.dout(w_dff_A_iwFPN9Lb6_1),.din(w_dff_A_OHdBHNXF9_1),.clk(gclk));
	jdff dff_A_l60AQmtu6_1(.dout(w_dff_A_OHdBHNXF9_1),.din(w_dff_A_l60AQmtu6_1),.clk(gclk));
	jdff dff_A_kro1kpmS6_1(.dout(w_dff_A_l60AQmtu6_1),.din(w_dff_A_kro1kpmS6_1),.clk(gclk));
	jdff dff_A_1K1g5fbW6_1(.dout(w_dff_A_kro1kpmS6_1),.din(w_dff_A_1K1g5fbW6_1),.clk(gclk));
	jdff dff_B_qThZXVAS5_1(.din(n1557),.dout(w_dff_B_qThZXVAS5_1),.clk(gclk));
	jdff dff_B_4KsNT68r4_1(.din(w_dff_B_qThZXVAS5_1),.dout(w_dff_B_4KsNT68r4_1),.clk(gclk));
	jdff dff_B_m0321h2C0_1(.din(w_dff_B_4KsNT68r4_1),.dout(w_dff_B_m0321h2C0_1),.clk(gclk));
	jdff dff_B_AtHV9SqQ6_1(.din(w_dff_B_m0321h2C0_1),.dout(w_dff_B_AtHV9SqQ6_1),.clk(gclk));
	jdff dff_B_1taZFBdh8_1(.din(w_dff_B_AtHV9SqQ6_1),.dout(w_dff_B_1taZFBdh8_1),.clk(gclk));
	jdff dff_B_ZuRuUN8X6_1(.din(w_dff_B_1taZFBdh8_1),.dout(w_dff_B_ZuRuUN8X6_1),.clk(gclk));
	jdff dff_B_RNNhOt3S1_1(.din(w_dff_B_ZuRuUN8X6_1),.dout(w_dff_B_RNNhOt3S1_1),.clk(gclk));
	jdff dff_B_PaiXs0mt7_1(.din(w_dff_B_RNNhOt3S1_1),.dout(w_dff_B_PaiXs0mt7_1),.clk(gclk));
	jdff dff_B_tH6DKS5D0_0(.din(n1558),.dout(w_dff_B_tH6DKS5D0_0),.clk(gclk));
	jdff dff_B_wAzPyPXZ1_0(.din(w_dff_B_tH6DKS5D0_0),.dout(w_dff_B_wAzPyPXZ1_0),.clk(gclk));
	jdff dff_B_453u6ucA1_0(.din(w_dff_B_wAzPyPXZ1_0),.dout(w_dff_B_453u6ucA1_0),.clk(gclk));
	jdff dff_B_KBA9Z8uR9_0(.din(w_dff_B_453u6ucA1_0),.dout(w_dff_B_KBA9Z8uR9_0),.clk(gclk));
	jdff dff_B_eK1Ui84y8_0(.din(w_dff_B_KBA9Z8uR9_0),.dout(w_dff_B_eK1Ui84y8_0),.clk(gclk));
	jdff dff_B_qqrw33Vf4_0(.din(w_dff_B_eK1Ui84y8_0),.dout(w_dff_B_qqrw33Vf4_0),.clk(gclk));
	jdff dff_A_sBMcs55T8_1(.dout(w_n1555_0[1]),.din(w_dff_A_sBMcs55T8_1),.clk(gclk));
	jdff dff_A_fyj4QY1o3_1(.dout(w_dff_A_sBMcs55T8_1),.din(w_dff_A_fyj4QY1o3_1),.clk(gclk));
	jdff dff_A_oxyUvhSv3_1(.dout(w_dff_A_fyj4QY1o3_1),.din(w_dff_A_oxyUvhSv3_1),.clk(gclk));
	jdff dff_A_aaetnem01_1(.dout(w_dff_A_oxyUvhSv3_1),.din(w_dff_A_aaetnem01_1),.clk(gclk));
	jdff dff_A_Bw5tnDwG9_1(.dout(w_dff_A_aaetnem01_1),.din(w_dff_A_Bw5tnDwG9_1),.clk(gclk));
	jdff dff_A_vFKT07tG1_1(.dout(w_dff_A_Bw5tnDwG9_1),.din(w_dff_A_vFKT07tG1_1),.clk(gclk));
	jdff dff_A_0GFTuX1r9_1(.dout(w_dff_A_vFKT07tG1_1),.din(w_dff_A_0GFTuX1r9_1),.clk(gclk));
	jdff dff_B_89zGTgIV5_1(.din(n1488),.dout(w_dff_B_89zGTgIV5_1),.clk(gclk));
	jdff dff_B_tbNkuEda9_1(.din(w_dff_B_89zGTgIV5_1),.dout(w_dff_B_tbNkuEda9_1),.clk(gclk));
	jdff dff_B_Lf1hSQTd4_1(.din(w_dff_B_tbNkuEda9_1),.dout(w_dff_B_Lf1hSQTd4_1),.clk(gclk));
	jdff dff_B_B7Y8Xqzg5_1(.din(w_dff_B_Lf1hSQTd4_1),.dout(w_dff_B_B7Y8Xqzg5_1),.clk(gclk));
	jdff dff_B_sipoZOv55_1(.din(w_dff_B_B7Y8Xqzg5_1),.dout(w_dff_B_sipoZOv55_1),.clk(gclk));
	jdff dff_B_I6yWBDMP5_1(.din(w_dff_B_sipoZOv55_1),.dout(w_dff_B_I6yWBDMP5_1),.clk(gclk));
	jdff dff_B_uM7kyvMl1_1(.din(w_dff_B_I6yWBDMP5_1),.dout(w_dff_B_uM7kyvMl1_1),.clk(gclk));
	jdff dff_B_BOAjz2Gm4_0(.din(n1489),.dout(w_dff_B_BOAjz2Gm4_0),.clk(gclk));
	jdff dff_B_NlqWlu6X0_0(.din(w_dff_B_BOAjz2Gm4_0),.dout(w_dff_B_NlqWlu6X0_0),.clk(gclk));
	jdff dff_B_NBYt3pqa5_0(.din(w_dff_B_NlqWlu6X0_0),.dout(w_dff_B_NBYt3pqa5_0),.clk(gclk));
	jdff dff_B_WfTwraRJ8_0(.din(w_dff_B_NBYt3pqa5_0),.dout(w_dff_B_WfTwraRJ8_0),.clk(gclk));
	jdff dff_B_fW2lPW9w3_0(.din(w_dff_B_WfTwraRJ8_0),.dout(w_dff_B_fW2lPW9w3_0),.clk(gclk));
	jdff dff_A_YyE8LCpd2_1(.dout(w_n1486_0[1]),.din(w_dff_A_YyE8LCpd2_1),.clk(gclk));
	jdff dff_A_kyqDLJ360_1(.dout(w_dff_A_YyE8LCpd2_1),.din(w_dff_A_kyqDLJ360_1),.clk(gclk));
	jdff dff_A_yVVeluAA9_1(.dout(w_dff_A_kyqDLJ360_1),.din(w_dff_A_yVVeluAA9_1),.clk(gclk));
	jdff dff_A_BK3FG69W3_1(.dout(w_dff_A_yVVeluAA9_1),.din(w_dff_A_BK3FG69W3_1),.clk(gclk));
	jdff dff_A_bd6lX0Qc8_1(.dout(w_dff_A_BK3FG69W3_1),.din(w_dff_A_bd6lX0Qc8_1),.clk(gclk));
	jdff dff_A_aEBeq1PX8_1(.dout(w_dff_A_bd6lX0Qc8_1),.din(w_dff_A_aEBeq1PX8_1),.clk(gclk));
	jdff dff_B_7YPz0EEJ5_1(.din(n1412),.dout(w_dff_B_7YPz0EEJ5_1),.clk(gclk));
	jdff dff_B_vSqMAagr0_1(.din(w_dff_B_7YPz0EEJ5_1),.dout(w_dff_B_vSqMAagr0_1),.clk(gclk));
	jdff dff_B_g1EjlE8T9_1(.din(w_dff_B_vSqMAagr0_1),.dout(w_dff_B_g1EjlE8T9_1),.clk(gclk));
	jdff dff_B_UukhTS6B9_1(.din(w_dff_B_g1EjlE8T9_1),.dout(w_dff_B_UukhTS6B9_1),.clk(gclk));
	jdff dff_B_TnCH5q7Z6_1(.din(w_dff_B_UukhTS6B9_1),.dout(w_dff_B_TnCH5q7Z6_1),.clk(gclk));
	jdff dff_B_WWr6rpmz9_1(.din(w_dff_B_TnCH5q7Z6_1),.dout(w_dff_B_WWr6rpmz9_1),.clk(gclk));
	jdff dff_B_fwtVPQSN3_0(.din(n1413),.dout(w_dff_B_fwtVPQSN3_0),.clk(gclk));
	jdff dff_B_od5UusqG5_0(.din(w_dff_B_fwtVPQSN3_0),.dout(w_dff_B_od5UusqG5_0),.clk(gclk));
	jdff dff_B_L58Alc1U3_0(.din(w_dff_B_od5UusqG5_0),.dout(w_dff_B_L58Alc1U3_0),.clk(gclk));
	jdff dff_B_RMHEEMGh8_0(.din(w_dff_B_L58Alc1U3_0),.dout(w_dff_B_RMHEEMGh8_0),.clk(gclk));
	jdff dff_A_icapOvkN0_1(.dout(w_n1410_0[1]),.din(w_dff_A_icapOvkN0_1),.clk(gclk));
	jdff dff_A_Dh0iTn9n1_1(.dout(w_dff_A_icapOvkN0_1),.din(w_dff_A_Dh0iTn9n1_1),.clk(gclk));
	jdff dff_A_00RSsezR6_1(.dout(w_dff_A_Dh0iTn9n1_1),.din(w_dff_A_00RSsezR6_1),.clk(gclk));
	jdff dff_A_adH5Mp8P7_1(.dout(w_dff_A_00RSsezR6_1),.din(w_dff_A_adH5Mp8P7_1),.clk(gclk));
	jdff dff_A_VznJHwpx9_1(.dout(w_dff_A_adH5Mp8P7_1),.din(w_dff_A_VznJHwpx9_1),.clk(gclk));
	jdff dff_B_EaACql833_1(.din(n1330),.dout(w_dff_B_EaACql833_1),.clk(gclk));
	jdff dff_B_CNq2ygGW5_1(.din(w_dff_B_EaACql833_1),.dout(w_dff_B_CNq2ygGW5_1),.clk(gclk));
	jdff dff_B_3s0PRdKJ2_1(.din(w_dff_B_CNq2ygGW5_1),.dout(w_dff_B_3s0PRdKJ2_1),.clk(gclk));
	jdff dff_A_MOiX7ir23_0(.dout(w_n1326_0[0]),.din(w_dff_A_MOiX7ir23_0),.clk(gclk));
	jdff dff_A_K4ToNhLz9_0(.dout(w_dff_A_MOiX7ir23_0),.din(w_dff_A_K4ToNhLz9_0),.clk(gclk));
	jdff dff_B_BFNl21zT8_1(.din(n1242),.dout(w_dff_B_BFNl21zT8_1),.clk(gclk));
	jdff dff_A_8LRjp0fZ3_0(.dout(w_n1238_0[0]),.din(w_dff_A_8LRjp0fZ3_0),.clk(gclk));
	jdff dff_B_YxY9L11J6_1(.din(n1145),.dout(w_dff_B_YxY9L11J6_1),.clk(gclk));
	jdff dff_A_BLchi0CF4_1(.dout(w_n1039_0[1]),.din(w_dff_A_BLchi0CF4_1),.clk(gclk));
	jdff dff_B_6NEy3HGz2_2(.din(n1037),.dout(w_dff_B_6NEy3HGz2_2),.clk(gclk));
	jdff dff_B_uKVEnDbQ2_1(.din(n935),.dout(w_dff_B_uKVEnDbQ2_1),.clk(gclk));
	jdff dff_A_6V7hrwzn6_0(.dout(w_n829_0[0]),.din(w_dff_A_6V7hrwzn6_0),.clk(gclk));
	jdff dff_A_fNxtcm6l6_0(.dout(w_dff_A_6V7hrwzn6_0),.din(w_dff_A_fNxtcm6l6_0),.clk(gclk));
	jdff dff_A_6F0XgFpA4_0(.dout(w_dff_A_fNxtcm6l6_0),.din(w_dff_A_6F0XgFpA4_0),.clk(gclk));
	jdff dff_A_J44bVdcI7_0(.dout(w_dff_A_6F0XgFpA4_0),.din(w_dff_A_J44bVdcI7_0),.clk(gclk));
	jdff dff_A_psvP85Nc8_0(.dout(w_dff_A_J44bVdcI7_0),.din(w_dff_A_psvP85Nc8_0),.clk(gclk));
	jdff dff_A_svKF7qMX4_0(.dout(w_dff_A_psvP85Nc8_0),.din(w_dff_A_svKF7qMX4_0),.clk(gclk));
	jdff dff_A_ceoaJjlg4_0(.dout(w_dff_A_svKF7qMX4_0),.din(w_dff_A_ceoaJjlg4_0),.clk(gclk));
	jdff dff_A_uMh3wmh43_0(.dout(w_dff_A_ceoaJjlg4_0),.din(w_dff_A_uMh3wmh43_0),.clk(gclk));
	jdff dff_A_W9TbWtlx1_0(.dout(w_dff_A_uMh3wmh43_0),.din(w_dff_A_W9TbWtlx1_0),.clk(gclk));
	jdff dff_A_56uq5eD56_0(.dout(w_dff_A_W9TbWtlx1_0),.din(w_dff_A_56uq5eD56_0),.clk(gclk));
	jdff dff_A_pk7oJCgU3_0(.dout(w_dff_A_56uq5eD56_0),.din(w_dff_A_pk7oJCgU3_0),.clk(gclk));
	jdff dff_A_OWeYt4PU1_0(.dout(w_dff_A_pk7oJCgU3_0),.din(w_dff_A_OWeYt4PU1_0),.clk(gclk));
	jdff dff_A_BRlYgQwf5_0(.dout(w_dff_A_OWeYt4PU1_0),.din(w_dff_A_BRlYgQwf5_0),.clk(gclk));
	jdff dff_A_lXeA3x2S5_0(.dout(w_dff_A_BRlYgQwf5_0),.din(w_dff_A_lXeA3x2S5_0),.clk(gclk));
	jdff dff_A_izlyF6sL0_0(.dout(w_dff_A_lXeA3x2S5_0),.din(w_dff_A_izlyF6sL0_0),.clk(gclk));
	jdff dff_A_8v87OChG1_0(.dout(w_dff_A_izlyF6sL0_0),.din(w_dff_A_8v87OChG1_0),.clk(gclk));
	jdff dff_A_Q37cT2OV6_0(.dout(w_dff_A_8v87OChG1_0),.din(w_dff_A_Q37cT2OV6_0),.clk(gclk));
	jdff dff_A_8lR8qIBP6_0(.dout(w_dff_A_Q37cT2OV6_0),.din(w_dff_A_8lR8qIBP6_0),.clk(gclk));
	jdff dff_A_f2ymBBmN9_0(.dout(w_dff_A_8lR8qIBP6_0),.din(w_dff_A_f2ymBBmN9_0),.clk(gclk));
	jdff dff_A_uwxDyZH07_0(.dout(w_dff_A_f2ymBBmN9_0),.din(w_dff_A_uwxDyZH07_0),.clk(gclk));
	jdff dff_A_TaJiwgA97_0(.dout(w_dff_A_uwxDyZH07_0),.din(w_dff_A_TaJiwgA97_0),.clk(gclk));
	jdff dff_A_JsTOEFvp2_0(.dout(w_dff_A_TaJiwgA97_0),.din(w_dff_A_JsTOEFvp2_0),.clk(gclk));
	jdff dff_A_5XoUr31V9_0(.dout(w_dff_A_JsTOEFvp2_0),.din(w_dff_A_5XoUr31V9_0),.clk(gclk));
	jdff dff_A_s2FCC40a3_0(.dout(w_dff_A_5XoUr31V9_0),.din(w_dff_A_s2FCC40a3_0),.clk(gclk));
	jdff dff_A_rCDjsYt57_0(.dout(w_dff_A_s2FCC40a3_0),.din(w_dff_A_rCDjsYt57_0),.clk(gclk));
	jdff dff_A_6XcoHjrL7_0(.dout(w_dff_A_rCDjsYt57_0),.din(w_dff_A_6XcoHjrL7_0),.clk(gclk));
	jdff dff_A_plIe5c5R0_0(.dout(w_dff_A_6XcoHjrL7_0),.din(w_dff_A_plIe5c5R0_0),.clk(gclk));
	jdff dff_A_lXIm4D0B8_0(.dout(w_dff_A_plIe5c5R0_0),.din(w_dff_A_lXIm4D0B8_0),.clk(gclk));
	jdff dff_A_cjOmuz7j2_0(.dout(w_dff_A_lXIm4D0B8_0),.din(w_dff_A_cjOmuz7j2_0),.clk(gclk));
	jdff dff_A_MQJ1NTqI4_0(.dout(w_dff_A_cjOmuz7j2_0),.din(w_dff_A_MQJ1NTqI4_0),.clk(gclk));
	jdff dff_A_6pA4xgLf6_0(.dout(w_dff_A_MQJ1NTqI4_0),.din(w_dff_A_6pA4xgLf6_0),.clk(gclk));
	jdff dff_A_AVj3Kxvt1_0(.dout(w_dff_A_6pA4xgLf6_0),.din(w_dff_A_AVj3Kxvt1_0),.clk(gclk));
	jdff dff_A_riwt5X847_0(.dout(w_dff_A_AVj3Kxvt1_0),.din(w_dff_A_riwt5X847_0),.clk(gclk));
	jdff dff_A_hQVe51HY8_0(.dout(w_dff_A_riwt5X847_0),.din(w_dff_A_hQVe51HY8_0),.clk(gclk));
	jdff dff_A_CT7W2dHd3_0(.dout(w_dff_A_hQVe51HY8_0),.din(w_dff_A_CT7W2dHd3_0),.clk(gclk));
	jdff dff_A_lHUiqZYq7_0(.dout(w_dff_A_CT7W2dHd3_0),.din(w_dff_A_lHUiqZYq7_0),.clk(gclk));
	jdff dff_A_0DwLaxM29_0(.dout(w_dff_A_lHUiqZYq7_0),.din(w_dff_A_0DwLaxM29_0),.clk(gclk));
	jdff dff_A_cvpYQpNF5_0(.dout(w_dff_A_0DwLaxM29_0),.din(w_dff_A_cvpYQpNF5_0),.clk(gclk));
	jdff dff_A_K5Az5ea85_0(.dout(w_dff_A_cvpYQpNF5_0),.din(w_dff_A_K5Az5ea85_0),.clk(gclk));
	jdff dff_A_9jw0b8U63_0(.dout(w_dff_A_K5Az5ea85_0),.din(w_dff_A_9jw0b8U63_0),.clk(gclk));
	jdff dff_A_UJ9I5hKy2_0(.dout(w_dff_A_9jw0b8U63_0),.din(w_dff_A_UJ9I5hKy2_0),.clk(gclk));
	jdff dff_A_0ZD60s2I6_0(.dout(w_dff_A_UJ9I5hKy2_0),.din(w_dff_A_0ZD60s2I6_0),.clk(gclk));
	jdff dff_A_6Qm3LNbZ2_0(.dout(w_dff_A_0ZD60s2I6_0),.din(w_dff_A_6Qm3LNbZ2_0),.clk(gclk));
	jdff dff_A_4Cy19Jzl6_0(.dout(w_dff_A_6Qm3LNbZ2_0),.din(w_dff_A_4Cy19Jzl6_0),.clk(gclk));
	jdff dff_A_nNe7f8Xx0_1(.dout(w_n931_0[1]),.din(w_dff_A_nNe7f8Xx0_1),.clk(gclk));
	jdff dff_B_cm5qEtPD6_1(.din(n832),.dout(w_dff_B_cm5qEtPD6_1),.clk(gclk));
	jdff dff_A_hpkQO7MK5_0(.dout(w_n729_0[0]),.din(w_dff_A_hpkQO7MK5_0),.clk(gclk));
	jdff dff_A_S0gkK6by2_0(.dout(w_dff_A_hpkQO7MK5_0),.din(w_dff_A_S0gkK6by2_0),.clk(gclk));
	jdff dff_A_wv30d5M87_0(.dout(w_dff_A_S0gkK6by2_0),.din(w_dff_A_wv30d5M87_0),.clk(gclk));
	jdff dff_A_l5LiC6On9_0(.dout(w_dff_A_wv30d5M87_0),.din(w_dff_A_l5LiC6On9_0),.clk(gclk));
	jdff dff_A_x8gfXW7k9_0(.dout(w_dff_A_l5LiC6On9_0),.din(w_dff_A_x8gfXW7k9_0),.clk(gclk));
	jdff dff_A_sZ1guD3X8_0(.dout(w_dff_A_x8gfXW7k9_0),.din(w_dff_A_sZ1guD3X8_0),.clk(gclk));
	jdff dff_A_AMEnIHwt7_0(.dout(w_dff_A_sZ1guD3X8_0),.din(w_dff_A_AMEnIHwt7_0),.clk(gclk));
	jdff dff_A_XOlSkgMJ2_0(.dout(w_dff_A_AMEnIHwt7_0),.din(w_dff_A_XOlSkgMJ2_0),.clk(gclk));
	jdff dff_A_BYrGcG2S3_0(.dout(w_dff_A_XOlSkgMJ2_0),.din(w_dff_A_BYrGcG2S3_0),.clk(gclk));
	jdff dff_A_QEu5ft5c4_0(.dout(w_dff_A_BYrGcG2S3_0),.din(w_dff_A_QEu5ft5c4_0),.clk(gclk));
	jdff dff_A_4dHJ5FnO9_0(.dout(w_dff_A_QEu5ft5c4_0),.din(w_dff_A_4dHJ5FnO9_0),.clk(gclk));
	jdff dff_A_0qZAWYTK7_0(.dout(w_dff_A_4dHJ5FnO9_0),.din(w_dff_A_0qZAWYTK7_0),.clk(gclk));
	jdff dff_A_uF596t8g2_0(.dout(w_dff_A_0qZAWYTK7_0),.din(w_dff_A_uF596t8g2_0),.clk(gclk));
	jdff dff_A_ijqfPpKd9_0(.dout(w_dff_A_uF596t8g2_0),.din(w_dff_A_ijqfPpKd9_0),.clk(gclk));
	jdff dff_A_Ug3QQrpa5_0(.dout(w_dff_A_ijqfPpKd9_0),.din(w_dff_A_Ug3QQrpa5_0),.clk(gclk));
	jdff dff_A_ZR61NCGG8_0(.dout(w_dff_A_Ug3QQrpa5_0),.din(w_dff_A_ZR61NCGG8_0),.clk(gclk));
	jdff dff_A_v4Ozbc4b5_0(.dout(w_dff_A_ZR61NCGG8_0),.din(w_dff_A_v4Ozbc4b5_0),.clk(gclk));
	jdff dff_A_WwPIPAVl7_0(.dout(w_dff_A_v4Ozbc4b5_0),.din(w_dff_A_WwPIPAVl7_0),.clk(gclk));
	jdff dff_A_gb66Bs6G0_0(.dout(w_dff_A_WwPIPAVl7_0),.din(w_dff_A_gb66Bs6G0_0),.clk(gclk));
	jdff dff_A_uFyblmZr5_0(.dout(w_dff_A_gb66Bs6G0_0),.din(w_dff_A_uFyblmZr5_0),.clk(gclk));
	jdff dff_A_jzHJH7ng6_0(.dout(w_dff_A_uFyblmZr5_0),.din(w_dff_A_jzHJH7ng6_0),.clk(gclk));
	jdff dff_A_kvrYy2i36_0(.dout(w_dff_A_jzHJH7ng6_0),.din(w_dff_A_kvrYy2i36_0),.clk(gclk));
	jdff dff_A_5bfFOKNy9_0(.dout(w_dff_A_kvrYy2i36_0),.din(w_dff_A_5bfFOKNy9_0),.clk(gclk));
	jdff dff_A_YTXbspCj6_0(.dout(w_dff_A_5bfFOKNy9_0),.din(w_dff_A_YTXbspCj6_0),.clk(gclk));
	jdff dff_A_QbgmQ9GR0_0(.dout(w_dff_A_YTXbspCj6_0),.din(w_dff_A_QbgmQ9GR0_0),.clk(gclk));
	jdff dff_A_DWtzE9Lg9_0(.dout(w_dff_A_QbgmQ9GR0_0),.din(w_dff_A_DWtzE9Lg9_0),.clk(gclk));
	jdff dff_A_rD2ES1qK5_0(.dout(w_dff_A_DWtzE9Lg9_0),.din(w_dff_A_rD2ES1qK5_0),.clk(gclk));
	jdff dff_A_M8jWDMan9_0(.dout(w_dff_A_rD2ES1qK5_0),.din(w_dff_A_M8jWDMan9_0),.clk(gclk));
	jdff dff_A_D9l9qJ8J3_0(.dout(w_dff_A_M8jWDMan9_0),.din(w_dff_A_D9l9qJ8J3_0),.clk(gclk));
	jdff dff_A_hd2BDvex8_0(.dout(w_dff_A_D9l9qJ8J3_0),.din(w_dff_A_hd2BDvex8_0),.clk(gclk));
	jdff dff_A_pQIeJ1yR6_0(.dout(w_dff_A_hd2BDvex8_0),.din(w_dff_A_pQIeJ1yR6_0),.clk(gclk));
	jdff dff_A_3nxdof6H0_0(.dout(w_dff_A_pQIeJ1yR6_0),.din(w_dff_A_3nxdof6H0_0),.clk(gclk));
	jdff dff_A_j3UuPga36_0(.dout(w_dff_A_3nxdof6H0_0),.din(w_dff_A_j3UuPga36_0),.clk(gclk));
	jdff dff_A_jnYUxKz76_0(.dout(w_dff_A_j3UuPga36_0),.din(w_dff_A_jnYUxKz76_0),.clk(gclk));
	jdff dff_A_s9qkdFRi6_0(.dout(w_dff_A_jnYUxKz76_0),.din(w_dff_A_s9qkdFRi6_0),.clk(gclk));
	jdff dff_A_0Qx3SRCO8_0(.dout(w_dff_A_s9qkdFRi6_0),.din(w_dff_A_0Qx3SRCO8_0),.clk(gclk));
	jdff dff_A_uknZAKxN2_0(.dout(w_dff_A_0Qx3SRCO8_0),.din(w_dff_A_uknZAKxN2_0),.clk(gclk));
	jdff dff_A_jIWh811E7_0(.dout(w_dff_A_uknZAKxN2_0),.din(w_dff_A_jIWh811E7_0),.clk(gclk));
	jdff dff_A_CDbqx1dQ0_0(.dout(w_dff_A_jIWh811E7_0),.din(w_dff_A_CDbqx1dQ0_0),.clk(gclk));
	jdff dff_A_zTPZjg254_0(.dout(w_dff_A_CDbqx1dQ0_0),.din(w_dff_A_zTPZjg254_0),.clk(gclk));
	jdff dff_A_O44AF8rm8_0(.dout(w_dff_A_zTPZjg254_0),.din(w_dff_A_O44AF8rm8_0),.clk(gclk));
	jdff dff_A_ve3QpJuC3_1(.dout(w_n826_0[1]),.din(w_dff_A_ve3QpJuC3_1),.clk(gclk));
	jdff dff_B_L99dMJIv6_1(.din(n736),.dout(w_dff_B_L99dMJIv6_1),.clk(gclk));
	jdff dff_B_KKp1gkxY3_1(.din(w_dff_B_L99dMJIv6_1),.dout(w_dff_B_KKp1gkxY3_1),.clk(gclk));
	jdff dff_B_OprdLYLo0_1(.din(w_dff_B_KKp1gkxY3_1),.dout(w_dff_B_OprdLYLo0_1),.clk(gclk));
	jdff dff_B_76Lwyahd0_1(.din(w_dff_B_OprdLYLo0_1),.dout(w_dff_B_76Lwyahd0_1),.clk(gclk));
	jdff dff_B_bwVhD8xL5_1(.din(w_dff_B_76Lwyahd0_1),.dout(w_dff_B_bwVhD8xL5_1),.clk(gclk));
	jdff dff_B_c9FhlcRE6_1(.din(w_dff_B_bwVhD8xL5_1),.dout(w_dff_B_c9FhlcRE6_1),.clk(gclk));
	jdff dff_B_db3vdHwX2_1(.din(w_dff_B_c9FhlcRE6_1),.dout(w_dff_B_db3vdHwX2_1),.clk(gclk));
	jdff dff_B_TzrojeaV2_1(.din(w_dff_B_db3vdHwX2_1),.dout(w_dff_B_TzrojeaV2_1),.clk(gclk));
	jdff dff_B_OdyuZ8aR4_1(.din(w_dff_B_TzrojeaV2_1),.dout(w_dff_B_OdyuZ8aR4_1),.clk(gclk));
	jdff dff_B_OtluU48w3_1(.din(w_dff_B_OdyuZ8aR4_1),.dout(w_dff_B_OtluU48w3_1),.clk(gclk));
	jdff dff_B_1rwJXIys4_1(.din(w_dff_B_OtluU48w3_1),.dout(w_dff_B_1rwJXIys4_1),.clk(gclk));
	jdff dff_B_yNTuvNMC9_1(.din(w_dff_B_1rwJXIys4_1),.dout(w_dff_B_yNTuvNMC9_1),.clk(gclk));
	jdff dff_B_O7B3LFZ33_1(.din(w_dff_B_yNTuvNMC9_1),.dout(w_dff_B_O7B3LFZ33_1),.clk(gclk));
	jdff dff_B_Dt2BYe0z8_1(.din(w_dff_B_O7B3LFZ33_1),.dout(w_dff_B_Dt2BYe0z8_1),.clk(gclk));
	jdff dff_B_bph5RScJ6_1(.din(w_dff_B_Dt2BYe0z8_1),.dout(w_dff_B_bph5RScJ6_1),.clk(gclk));
	jdff dff_B_srYuAKkj3_1(.din(w_dff_B_bph5RScJ6_1),.dout(w_dff_B_srYuAKkj3_1),.clk(gclk));
	jdff dff_B_22bIZSn63_1(.din(w_dff_B_srYuAKkj3_1),.dout(w_dff_B_22bIZSn63_1),.clk(gclk));
	jdff dff_B_lYRTQzSs5_1(.din(w_dff_B_22bIZSn63_1),.dout(w_dff_B_lYRTQzSs5_1),.clk(gclk));
	jdff dff_B_hcq8z5Yw5_1(.din(w_dff_B_lYRTQzSs5_1),.dout(w_dff_B_hcq8z5Yw5_1),.clk(gclk));
	jdff dff_B_5PdSpXBM8_1(.din(w_dff_B_hcq8z5Yw5_1),.dout(w_dff_B_5PdSpXBM8_1),.clk(gclk));
	jdff dff_B_o3oBp1mo1_1(.din(w_dff_B_5PdSpXBM8_1),.dout(w_dff_B_o3oBp1mo1_1),.clk(gclk));
	jdff dff_B_eEfCfQXT7_1(.din(w_dff_B_o3oBp1mo1_1),.dout(w_dff_B_eEfCfQXT7_1),.clk(gclk));
	jdff dff_B_HTVDmjNe4_1(.din(w_dff_B_eEfCfQXT7_1),.dout(w_dff_B_HTVDmjNe4_1),.clk(gclk));
	jdff dff_B_bA9Iry2k2_1(.din(w_dff_B_HTVDmjNe4_1),.dout(w_dff_B_bA9Iry2k2_1),.clk(gclk));
	jdff dff_B_xcpF8nml9_1(.din(w_dff_B_bA9Iry2k2_1),.dout(w_dff_B_xcpF8nml9_1),.clk(gclk));
	jdff dff_B_OyxFWTsp4_1(.din(w_dff_B_xcpF8nml9_1),.dout(w_dff_B_OyxFWTsp4_1),.clk(gclk));
	jdff dff_B_qoWgq2Zp2_1(.din(w_dff_B_OyxFWTsp4_1),.dout(w_dff_B_qoWgq2Zp2_1),.clk(gclk));
	jdff dff_B_u6EardZn0_1(.din(w_dff_B_qoWgq2Zp2_1),.dout(w_dff_B_u6EardZn0_1),.clk(gclk));
	jdff dff_B_of8g8xc52_1(.din(w_dff_B_u6EardZn0_1),.dout(w_dff_B_of8g8xc52_1),.clk(gclk));
	jdff dff_B_Qasj3y822_1(.din(w_dff_B_of8g8xc52_1),.dout(w_dff_B_Qasj3y822_1),.clk(gclk));
	jdff dff_B_g0HV2ilx8_1(.din(w_dff_B_Qasj3y822_1),.dout(w_dff_B_g0HV2ilx8_1),.clk(gclk));
	jdff dff_B_A5sm3Avt5_1(.din(w_dff_B_g0HV2ilx8_1),.dout(w_dff_B_A5sm3Avt5_1),.clk(gclk));
	jdff dff_B_xuTN1zfU2_1(.din(w_dff_B_A5sm3Avt5_1),.dout(w_dff_B_xuTN1zfU2_1),.clk(gclk));
	jdff dff_B_0NtVP1NK5_1(.din(w_dff_B_xuTN1zfU2_1),.dout(w_dff_B_0NtVP1NK5_1),.clk(gclk));
	jdff dff_B_gZlEn6vm6_1(.din(w_dff_B_0NtVP1NK5_1),.dout(w_dff_B_gZlEn6vm6_1),.clk(gclk));
	jdff dff_B_VyAkWJzf9_1(.din(w_dff_B_gZlEn6vm6_1),.dout(w_dff_B_VyAkWJzf9_1),.clk(gclk));
	jdff dff_B_6piPLQWx6_1(.din(w_dff_B_VyAkWJzf9_1),.dout(w_dff_B_6piPLQWx6_1),.clk(gclk));
	jdff dff_B_XehIwMva3_1(.din(n732),.dout(w_dff_B_XehIwMva3_1),.clk(gclk));
	jdff dff_A_dkFBMNyd3_0(.dout(w_n636_0[0]),.din(w_dff_A_dkFBMNyd3_0),.clk(gclk));
	jdff dff_A_IYbI70kl3_0(.dout(w_dff_A_dkFBMNyd3_0),.din(w_dff_A_IYbI70kl3_0),.clk(gclk));
	jdff dff_A_RV4KjewY1_0(.dout(w_dff_A_IYbI70kl3_0),.din(w_dff_A_RV4KjewY1_0),.clk(gclk));
	jdff dff_A_AD3xpUNw8_0(.dout(w_dff_A_RV4KjewY1_0),.din(w_dff_A_AD3xpUNw8_0),.clk(gclk));
	jdff dff_A_pZk4GdOh0_0(.dout(w_dff_A_AD3xpUNw8_0),.din(w_dff_A_pZk4GdOh0_0),.clk(gclk));
	jdff dff_A_T0CF8oMq8_0(.dout(w_dff_A_pZk4GdOh0_0),.din(w_dff_A_T0CF8oMq8_0),.clk(gclk));
	jdff dff_A_eUxaKqhA6_0(.dout(w_dff_A_T0CF8oMq8_0),.din(w_dff_A_eUxaKqhA6_0),.clk(gclk));
	jdff dff_A_FHxmToAu5_0(.dout(w_dff_A_eUxaKqhA6_0),.din(w_dff_A_FHxmToAu5_0),.clk(gclk));
	jdff dff_A_QsmErd6W4_0(.dout(w_dff_A_FHxmToAu5_0),.din(w_dff_A_QsmErd6W4_0),.clk(gclk));
	jdff dff_A_MnpNT35V7_0(.dout(w_dff_A_QsmErd6W4_0),.din(w_dff_A_MnpNT35V7_0),.clk(gclk));
	jdff dff_A_aQIKJJWY2_0(.dout(w_dff_A_MnpNT35V7_0),.din(w_dff_A_aQIKJJWY2_0),.clk(gclk));
	jdff dff_A_51EP7Rqb8_0(.dout(w_dff_A_aQIKJJWY2_0),.din(w_dff_A_51EP7Rqb8_0),.clk(gclk));
	jdff dff_A_DPrAYKxd9_0(.dout(w_dff_A_51EP7Rqb8_0),.din(w_dff_A_DPrAYKxd9_0),.clk(gclk));
	jdff dff_A_BJjSs7Ka8_0(.dout(w_dff_A_DPrAYKxd9_0),.din(w_dff_A_BJjSs7Ka8_0),.clk(gclk));
	jdff dff_A_6lMKKesw8_0(.dout(w_dff_A_BJjSs7Ka8_0),.din(w_dff_A_6lMKKesw8_0),.clk(gclk));
	jdff dff_A_oII8ASb93_0(.dout(w_dff_A_6lMKKesw8_0),.din(w_dff_A_oII8ASb93_0),.clk(gclk));
	jdff dff_A_5vYfnKTv1_0(.dout(w_dff_A_oII8ASb93_0),.din(w_dff_A_5vYfnKTv1_0),.clk(gclk));
	jdff dff_A_TObYhCgW7_0(.dout(w_dff_A_5vYfnKTv1_0),.din(w_dff_A_TObYhCgW7_0),.clk(gclk));
	jdff dff_A_0DYMsleC5_0(.dout(w_dff_A_TObYhCgW7_0),.din(w_dff_A_0DYMsleC5_0),.clk(gclk));
	jdff dff_A_fhKsflu15_0(.dout(w_dff_A_0DYMsleC5_0),.din(w_dff_A_fhKsflu15_0),.clk(gclk));
	jdff dff_A_6DrtfXqu5_0(.dout(w_dff_A_fhKsflu15_0),.din(w_dff_A_6DrtfXqu5_0),.clk(gclk));
	jdff dff_A_yL4F9Vsb6_0(.dout(w_dff_A_6DrtfXqu5_0),.din(w_dff_A_yL4F9Vsb6_0),.clk(gclk));
	jdff dff_A_waY3hmgA8_0(.dout(w_dff_A_yL4F9Vsb6_0),.din(w_dff_A_waY3hmgA8_0),.clk(gclk));
	jdff dff_A_KBExpihi0_0(.dout(w_dff_A_waY3hmgA8_0),.din(w_dff_A_KBExpihi0_0),.clk(gclk));
	jdff dff_A_YskG4wLk4_0(.dout(w_dff_A_KBExpihi0_0),.din(w_dff_A_YskG4wLk4_0),.clk(gclk));
	jdff dff_A_qpxTXPI91_0(.dout(w_dff_A_YskG4wLk4_0),.din(w_dff_A_qpxTXPI91_0),.clk(gclk));
	jdff dff_A_QwLV5MNt0_0(.dout(w_dff_A_qpxTXPI91_0),.din(w_dff_A_QwLV5MNt0_0),.clk(gclk));
	jdff dff_A_xzuvi9cr1_0(.dout(w_dff_A_QwLV5MNt0_0),.din(w_dff_A_xzuvi9cr1_0),.clk(gclk));
	jdff dff_A_deE9DqQJ7_0(.dout(w_dff_A_xzuvi9cr1_0),.din(w_dff_A_deE9DqQJ7_0),.clk(gclk));
	jdff dff_A_KaBZbPk31_0(.dout(w_dff_A_deE9DqQJ7_0),.din(w_dff_A_KaBZbPk31_0),.clk(gclk));
	jdff dff_A_OkqWzp1N0_0(.dout(w_dff_A_KaBZbPk31_0),.din(w_dff_A_OkqWzp1N0_0),.clk(gclk));
	jdff dff_A_Ofu4lpNa4_0(.dout(w_dff_A_OkqWzp1N0_0),.din(w_dff_A_Ofu4lpNa4_0),.clk(gclk));
	jdff dff_A_MQKVLyyw0_0(.dout(w_dff_A_Ofu4lpNa4_0),.din(w_dff_A_MQKVLyyw0_0),.clk(gclk));
	jdff dff_A_I2smT1Jo3_0(.dout(w_dff_A_MQKVLyyw0_0),.din(w_dff_A_I2smT1Jo3_0),.clk(gclk));
	jdff dff_A_W7hnBpyI7_0(.dout(w_dff_A_I2smT1Jo3_0),.din(w_dff_A_W7hnBpyI7_0),.clk(gclk));
	jdff dff_A_bLF0rPgD2_0(.dout(w_dff_A_W7hnBpyI7_0),.din(w_dff_A_bLF0rPgD2_0),.clk(gclk));
	jdff dff_A_4iRi0tfL7_0(.dout(w_dff_A_bLF0rPgD2_0),.din(w_dff_A_4iRi0tfL7_0),.clk(gclk));
	jdff dff_A_MyPZGV0G3_0(.dout(w_dff_A_4iRi0tfL7_0),.din(w_dff_A_MyPZGV0G3_0),.clk(gclk));
	jdff dff_A_hATT4C2w2_1(.dout(w_n726_0[1]),.din(w_dff_A_hATT4C2w2_1),.clk(gclk));
	jdff dff_B_YKDZx7fy4_1(.din(n643),.dout(w_dff_B_YKDZx7fy4_1),.clk(gclk));
	jdff dff_B_30CAmLrj8_1(.din(w_dff_B_YKDZx7fy4_1),.dout(w_dff_B_30CAmLrj8_1),.clk(gclk));
	jdff dff_B_0YaJDvfN2_1(.din(w_dff_B_30CAmLrj8_1),.dout(w_dff_B_0YaJDvfN2_1),.clk(gclk));
	jdff dff_B_xYO3EXLV4_1(.din(w_dff_B_0YaJDvfN2_1),.dout(w_dff_B_xYO3EXLV4_1),.clk(gclk));
	jdff dff_B_YRhavu0M3_1(.din(w_dff_B_xYO3EXLV4_1),.dout(w_dff_B_YRhavu0M3_1),.clk(gclk));
	jdff dff_B_gWiVubG23_1(.din(w_dff_B_YRhavu0M3_1),.dout(w_dff_B_gWiVubG23_1),.clk(gclk));
	jdff dff_B_h6IxwEcD2_1(.din(w_dff_B_gWiVubG23_1),.dout(w_dff_B_h6IxwEcD2_1),.clk(gclk));
	jdff dff_B_o8F9vjcx2_1(.din(w_dff_B_h6IxwEcD2_1),.dout(w_dff_B_o8F9vjcx2_1),.clk(gclk));
	jdff dff_B_rd95D0NW5_1(.din(w_dff_B_o8F9vjcx2_1),.dout(w_dff_B_rd95D0NW5_1),.clk(gclk));
	jdff dff_B_f2dDuNHD4_1(.din(w_dff_B_rd95D0NW5_1),.dout(w_dff_B_f2dDuNHD4_1),.clk(gclk));
	jdff dff_B_6UVGXx0J7_1(.din(w_dff_B_f2dDuNHD4_1),.dout(w_dff_B_6UVGXx0J7_1),.clk(gclk));
	jdff dff_B_zzhPxBZM3_1(.din(w_dff_B_6UVGXx0J7_1),.dout(w_dff_B_zzhPxBZM3_1),.clk(gclk));
	jdff dff_B_Le6VQwOB4_1(.din(w_dff_B_zzhPxBZM3_1),.dout(w_dff_B_Le6VQwOB4_1),.clk(gclk));
	jdff dff_B_ViuBbaOd0_1(.din(w_dff_B_Le6VQwOB4_1),.dout(w_dff_B_ViuBbaOd0_1),.clk(gclk));
	jdff dff_B_8AZluf0v6_1(.din(w_dff_B_ViuBbaOd0_1),.dout(w_dff_B_8AZluf0v6_1),.clk(gclk));
	jdff dff_B_JUi4qjU18_1(.din(w_dff_B_8AZluf0v6_1),.dout(w_dff_B_JUi4qjU18_1),.clk(gclk));
	jdff dff_B_JtZdrjT47_1(.din(w_dff_B_JUi4qjU18_1),.dout(w_dff_B_JtZdrjT47_1),.clk(gclk));
	jdff dff_B_B4lfhRrp4_1(.din(w_dff_B_JtZdrjT47_1),.dout(w_dff_B_B4lfhRrp4_1),.clk(gclk));
	jdff dff_B_ebo5fi4h9_1(.din(w_dff_B_B4lfhRrp4_1),.dout(w_dff_B_ebo5fi4h9_1),.clk(gclk));
	jdff dff_B_Zr7omRJh7_1(.din(w_dff_B_ebo5fi4h9_1),.dout(w_dff_B_Zr7omRJh7_1),.clk(gclk));
	jdff dff_B_2K1G3JGf0_1(.din(w_dff_B_Zr7omRJh7_1),.dout(w_dff_B_2K1G3JGf0_1),.clk(gclk));
	jdff dff_B_UuRafueM8_1(.din(w_dff_B_2K1G3JGf0_1),.dout(w_dff_B_UuRafueM8_1),.clk(gclk));
	jdff dff_B_jkTLqjWb8_1(.din(w_dff_B_UuRafueM8_1),.dout(w_dff_B_jkTLqjWb8_1),.clk(gclk));
	jdff dff_B_hMUURlBV9_1(.din(w_dff_B_jkTLqjWb8_1),.dout(w_dff_B_hMUURlBV9_1),.clk(gclk));
	jdff dff_B_WbWycBrW8_1(.din(w_dff_B_hMUURlBV9_1),.dout(w_dff_B_WbWycBrW8_1),.clk(gclk));
	jdff dff_B_ItSywzld8_1(.din(w_dff_B_WbWycBrW8_1),.dout(w_dff_B_ItSywzld8_1),.clk(gclk));
	jdff dff_B_ItYAKeDP6_1(.din(w_dff_B_ItSywzld8_1),.dout(w_dff_B_ItYAKeDP6_1),.clk(gclk));
	jdff dff_B_ogltcAiF7_1(.din(w_dff_B_ItYAKeDP6_1),.dout(w_dff_B_ogltcAiF7_1),.clk(gclk));
	jdff dff_B_sz1Trnej1_1(.din(w_dff_B_ogltcAiF7_1),.dout(w_dff_B_sz1Trnej1_1),.clk(gclk));
	jdff dff_B_Tqtrvtr68_1(.din(w_dff_B_sz1Trnej1_1),.dout(w_dff_B_Tqtrvtr68_1),.clk(gclk));
	jdff dff_B_5KlUi48L2_1(.din(w_dff_B_Tqtrvtr68_1),.dout(w_dff_B_5KlUi48L2_1),.clk(gclk));
	jdff dff_B_mFQJulWB4_1(.din(w_dff_B_5KlUi48L2_1),.dout(w_dff_B_mFQJulWB4_1),.clk(gclk));
	jdff dff_B_MA7cwNGm2_1(.din(w_dff_B_mFQJulWB4_1),.dout(w_dff_B_MA7cwNGm2_1),.clk(gclk));
	jdff dff_B_gR0O5Ao48_1(.din(w_dff_B_MA7cwNGm2_1),.dout(w_dff_B_gR0O5Ao48_1),.clk(gclk));
	jdff dff_B_ycRlJSps1_1(.din(n639),.dout(w_dff_B_ycRlJSps1_1),.clk(gclk));
	jdff dff_A_p7GUuktE2_0(.dout(w_n550_0[0]),.din(w_dff_A_p7GUuktE2_0),.clk(gclk));
	jdff dff_A_WHpTdWff5_0(.dout(w_dff_A_p7GUuktE2_0),.din(w_dff_A_WHpTdWff5_0),.clk(gclk));
	jdff dff_A_XCfgdy1a4_0(.dout(w_dff_A_WHpTdWff5_0),.din(w_dff_A_XCfgdy1a4_0),.clk(gclk));
	jdff dff_A_DRj5AaGN2_0(.dout(w_dff_A_XCfgdy1a4_0),.din(w_dff_A_DRj5AaGN2_0),.clk(gclk));
	jdff dff_A_94I3XL4l4_0(.dout(w_dff_A_DRj5AaGN2_0),.din(w_dff_A_94I3XL4l4_0),.clk(gclk));
	jdff dff_A_yy9zWcg31_0(.dout(w_dff_A_94I3XL4l4_0),.din(w_dff_A_yy9zWcg31_0),.clk(gclk));
	jdff dff_A_JeXyUzJI4_0(.dout(w_dff_A_yy9zWcg31_0),.din(w_dff_A_JeXyUzJI4_0),.clk(gclk));
	jdff dff_A_p4iV8HMX0_0(.dout(w_dff_A_JeXyUzJI4_0),.din(w_dff_A_p4iV8HMX0_0),.clk(gclk));
	jdff dff_A_fPsliYym6_0(.dout(w_dff_A_p4iV8HMX0_0),.din(w_dff_A_fPsliYym6_0),.clk(gclk));
	jdff dff_A_ZKMmuNkq9_0(.dout(w_dff_A_fPsliYym6_0),.din(w_dff_A_ZKMmuNkq9_0),.clk(gclk));
	jdff dff_A_gwudE4ZE6_0(.dout(w_dff_A_ZKMmuNkq9_0),.din(w_dff_A_gwudE4ZE6_0),.clk(gclk));
	jdff dff_A_9io5mtJi6_0(.dout(w_dff_A_gwudE4ZE6_0),.din(w_dff_A_9io5mtJi6_0),.clk(gclk));
	jdff dff_A_yYey6hKF0_0(.dout(w_dff_A_9io5mtJi6_0),.din(w_dff_A_yYey6hKF0_0),.clk(gclk));
	jdff dff_A_ZC2toaYY2_0(.dout(w_dff_A_yYey6hKF0_0),.din(w_dff_A_ZC2toaYY2_0),.clk(gclk));
	jdff dff_A_I5CCOEl28_0(.dout(w_dff_A_ZC2toaYY2_0),.din(w_dff_A_I5CCOEl28_0),.clk(gclk));
	jdff dff_A_Q1PIakiP2_0(.dout(w_dff_A_I5CCOEl28_0),.din(w_dff_A_Q1PIakiP2_0),.clk(gclk));
	jdff dff_A_HoZCIjjc0_0(.dout(w_dff_A_Q1PIakiP2_0),.din(w_dff_A_HoZCIjjc0_0),.clk(gclk));
	jdff dff_A_gBioCk720_0(.dout(w_dff_A_HoZCIjjc0_0),.din(w_dff_A_gBioCk720_0),.clk(gclk));
	jdff dff_A_fiU2mHFd9_0(.dout(w_dff_A_gBioCk720_0),.din(w_dff_A_fiU2mHFd9_0),.clk(gclk));
	jdff dff_A_Gb6RctpV2_0(.dout(w_dff_A_fiU2mHFd9_0),.din(w_dff_A_Gb6RctpV2_0),.clk(gclk));
	jdff dff_A_A3rKjPti5_0(.dout(w_dff_A_Gb6RctpV2_0),.din(w_dff_A_A3rKjPti5_0),.clk(gclk));
	jdff dff_A_8ueIGBPZ8_0(.dout(w_dff_A_A3rKjPti5_0),.din(w_dff_A_8ueIGBPZ8_0),.clk(gclk));
	jdff dff_A_MhypBxVz4_0(.dout(w_dff_A_8ueIGBPZ8_0),.din(w_dff_A_MhypBxVz4_0),.clk(gclk));
	jdff dff_A_PXkaP1gN3_0(.dout(w_dff_A_MhypBxVz4_0),.din(w_dff_A_PXkaP1gN3_0),.clk(gclk));
	jdff dff_A_lTvnh4hg6_0(.dout(w_dff_A_PXkaP1gN3_0),.din(w_dff_A_lTvnh4hg6_0),.clk(gclk));
	jdff dff_A_401zNE1z2_0(.dout(w_dff_A_lTvnh4hg6_0),.din(w_dff_A_401zNE1z2_0),.clk(gclk));
	jdff dff_A_HiI0Rbrh6_0(.dout(w_dff_A_401zNE1z2_0),.din(w_dff_A_HiI0Rbrh6_0),.clk(gclk));
	jdff dff_A_yB0SWjtR4_0(.dout(w_dff_A_HiI0Rbrh6_0),.din(w_dff_A_yB0SWjtR4_0),.clk(gclk));
	jdff dff_A_BtnbUn9A9_0(.dout(w_dff_A_yB0SWjtR4_0),.din(w_dff_A_BtnbUn9A9_0),.clk(gclk));
	jdff dff_A_wYQVAkQO0_0(.dout(w_dff_A_BtnbUn9A9_0),.din(w_dff_A_wYQVAkQO0_0),.clk(gclk));
	jdff dff_A_CyWGjM0H9_0(.dout(w_dff_A_wYQVAkQO0_0),.din(w_dff_A_CyWGjM0H9_0),.clk(gclk));
	jdff dff_A_KQhmwlZn2_0(.dout(w_dff_A_CyWGjM0H9_0),.din(w_dff_A_KQhmwlZn2_0),.clk(gclk));
	jdff dff_A_3WzrqVap0_0(.dout(w_dff_A_KQhmwlZn2_0),.din(w_dff_A_3WzrqVap0_0),.clk(gclk));
	jdff dff_A_AS5QDOLL6_0(.dout(w_dff_A_3WzrqVap0_0),.din(w_dff_A_AS5QDOLL6_0),.clk(gclk));
	jdff dff_A_U6tTMT4n6_0(.dout(w_dff_A_AS5QDOLL6_0),.din(w_dff_A_U6tTMT4n6_0),.clk(gclk));
	jdff dff_A_aPxlJXc64_1(.dout(w_n633_0[1]),.din(w_dff_A_aPxlJXc64_1),.clk(gclk));
	jdff dff_B_iy31NKBE3_1(.din(n557),.dout(w_dff_B_iy31NKBE3_1),.clk(gclk));
	jdff dff_B_RTB9HEF04_1(.din(w_dff_B_iy31NKBE3_1),.dout(w_dff_B_RTB9HEF04_1),.clk(gclk));
	jdff dff_B_I7c2d6g67_1(.din(w_dff_B_RTB9HEF04_1),.dout(w_dff_B_I7c2d6g67_1),.clk(gclk));
	jdff dff_B_gBizV6y55_1(.din(w_dff_B_I7c2d6g67_1),.dout(w_dff_B_gBizV6y55_1),.clk(gclk));
	jdff dff_B_a2aYoDrQ9_1(.din(w_dff_B_gBizV6y55_1),.dout(w_dff_B_a2aYoDrQ9_1),.clk(gclk));
	jdff dff_B_TBDvLm7N3_1(.din(w_dff_B_a2aYoDrQ9_1),.dout(w_dff_B_TBDvLm7N3_1),.clk(gclk));
	jdff dff_B_IqOAo8VR3_1(.din(w_dff_B_TBDvLm7N3_1),.dout(w_dff_B_IqOAo8VR3_1),.clk(gclk));
	jdff dff_B_OSVZOmad4_1(.din(w_dff_B_IqOAo8VR3_1),.dout(w_dff_B_OSVZOmad4_1),.clk(gclk));
	jdff dff_B_zCNee9JC4_1(.din(w_dff_B_OSVZOmad4_1),.dout(w_dff_B_zCNee9JC4_1),.clk(gclk));
	jdff dff_B_4ver7lNm3_1(.din(w_dff_B_zCNee9JC4_1),.dout(w_dff_B_4ver7lNm3_1),.clk(gclk));
	jdff dff_B_uiigXH6p4_1(.din(w_dff_B_4ver7lNm3_1),.dout(w_dff_B_uiigXH6p4_1),.clk(gclk));
	jdff dff_B_8VcGRPQe1_1(.din(w_dff_B_uiigXH6p4_1),.dout(w_dff_B_8VcGRPQe1_1),.clk(gclk));
	jdff dff_B_Vxa46z4X8_1(.din(w_dff_B_8VcGRPQe1_1),.dout(w_dff_B_Vxa46z4X8_1),.clk(gclk));
	jdff dff_B_nnl1cWl62_1(.din(w_dff_B_Vxa46z4X8_1),.dout(w_dff_B_nnl1cWl62_1),.clk(gclk));
	jdff dff_B_SEmewUDT4_1(.din(w_dff_B_nnl1cWl62_1),.dout(w_dff_B_SEmewUDT4_1),.clk(gclk));
	jdff dff_B_T4XHIcec4_1(.din(w_dff_B_SEmewUDT4_1),.dout(w_dff_B_T4XHIcec4_1),.clk(gclk));
	jdff dff_B_sKOzv35U8_1(.din(w_dff_B_T4XHIcec4_1),.dout(w_dff_B_sKOzv35U8_1),.clk(gclk));
	jdff dff_B_yEvHS9qk0_1(.din(w_dff_B_sKOzv35U8_1),.dout(w_dff_B_yEvHS9qk0_1),.clk(gclk));
	jdff dff_B_Ips5b0QF2_1(.din(w_dff_B_yEvHS9qk0_1),.dout(w_dff_B_Ips5b0QF2_1),.clk(gclk));
	jdff dff_B_UWKtcUi81_1(.din(w_dff_B_Ips5b0QF2_1),.dout(w_dff_B_UWKtcUi81_1),.clk(gclk));
	jdff dff_B_L4HA2sbK5_1(.din(w_dff_B_UWKtcUi81_1),.dout(w_dff_B_L4HA2sbK5_1),.clk(gclk));
	jdff dff_B_YydlJqw35_1(.din(w_dff_B_L4HA2sbK5_1),.dout(w_dff_B_YydlJqw35_1),.clk(gclk));
	jdff dff_B_bZESkjES9_1(.din(w_dff_B_YydlJqw35_1),.dout(w_dff_B_bZESkjES9_1),.clk(gclk));
	jdff dff_B_5Uifv4636_1(.din(w_dff_B_bZESkjES9_1),.dout(w_dff_B_5Uifv4636_1),.clk(gclk));
	jdff dff_B_nyAcTbUx9_1(.din(w_dff_B_5Uifv4636_1),.dout(w_dff_B_nyAcTbUx9_1),.clk(gclk));
	jdff dff_B_quG33DA47_1(.din(w_dff_B_nyAcTbUx9_1),.dout(w_dff_B_quG33DA47_1),.clk(gclk));
	jdff dff_B_DagU8vkE8_1(.din(w_dff_B_quG33DA47_1),.dout(w_dff_B_DagU8vkE8_1),.clk(gclk));
	jdff dff_B_NdnLBpy36_1(.din(w_dff_B_DagU8vkE8_1),.dout(w_dff_B_NdnLBpy36_1),.clk(gclk));
	jdff dff_B_qzLi7wxI0_1(.din(w_dff_B_NdnLBpy36_1),.dout(w_dff_B_qzLi7wxI0_1),.clk(gclk));
	jdff dff_B_vFSrm8xK7_1(.din(w_dff_B_qzLi7wxI0_1),.dout(w_dff_B_vFSrm8xK7_1),.clk(gclk));
	jdff dff_B_fSmRDmHs5_1(.din(w_dff_B_vFSrm8xK7_1),.dout(w_dff_B_fSmRDmHs5_1),.clk(gclk));
	jdff dff_B_qOHS1r4z9_1(.din(n553),.dout(w_dff_B_qOHS1r4z9_1),.clk(gclk));
	jdff dff_A_25J1ABlK1_0(.dout(w_n471_0[0]),.din(w_dff_A_25J1ABlK1_0),.clk(gclk));
	jdff dff_A_dN3XHPRR1_0(.dout(w_dff_A_25J1ABlK1_0),.din(w_dff_A_dN3XHPRR1_0),.clk(gclk));
	jdff dff_A_xhb7EiLO9_0(.dout(w_dff_A_dN3XHPRR1_0),.din(w_dff_A_xhb7EiLO9_0),.clk(gclk));
	jdff dff_A_fiM37NNF6_0(.dout(w_dff_A_xhb7EiLO9_0),.din(w_dff_A_fiM37NNF6_0),.clk(gclk));
	jdff dff_A_Vt79zmtK1_0(.dout(w_dff_A_fiM37NNF6_0),.din(w_dff_A_Vt79zmtK1_0),.clk(gclk));
	jdff dff_A_X86iegjD5_0(.dout(w_dff_A_Vt79zmtK1_0),.din(w_dff_A_X86iegjD5_0),.clk(gclk));
	jdff dff_A_1GqdSVGj9_0(.dout(w_dff_A_X86iegjD5_0),.din(w_dff_A_1GqdSVGj9_0),.clk(gclk));
	jdff dff_A_vNkKSNx74_0(.dout(w_dff_A_1GqdSVGj9_0),.din(w_dff_A_vNkKSNx74_0),.clk(gclk));
	jdff dff_A_At5yY3qr4_0(.dout(w_dff_A_vNkKSNx74_0),.din(w_dff_A_At5yY3qr4_0),.clk(gclk));
	jdff dff_A_GGZLjlkr5_0(.dout(w_dff_A_At5yY3qr4_0),.din(w_dff_A_GGZLjlkr5_0),.clk(gclk));
	jdff dff_A_JQnaDncF0_0(.dout(w_dff_A_GGZLjlkr5_0),.din(w_dff_A_JQnaDncF0_0),.clk(gclk));
	jdff dff_A_gHGlTTdY7_0(.dout(w_dff_A_JQnaDncF0_0),.din(w_dff_A_gHGlTTdY7_0),.clk(gclk));
	jdff dff_A_jEfy5eT24_0(.dout(w_dff_A_gHGlTTdY7_0),.din(w_dff_A_jEfy5eT24_0),.clk(gclk));
	jdff dff_A_6IQDB7TZ7_0(.dout(w_dff_A_jEfy5eT24_0),.din(w_dff_A_6IQDB7TZ7_0),.clk(gclk));
	jdff dff_A_E7tr3AmN3_0(.dout(w_dff_A_6IQDB7TZ7_0),.din(w_dff_A_E7tr3AmN3_0),.clk(gclk));
	jdff dff_A_hleiiF2t2_0(.dout(w_dff_A_E7tr3AmN3_0),.din(w_dff_A_hleiiF2t2_0),.clk(gclk));
	jdff dff_A_eqLjgLOn4_0(.dout(w_dff_A_hleiiF2t2_0),.din(w_dff_A_eqLjgLOn4_0),.clk(gclk));
	jdff dff_A_91W6l9NE5_0(.dout(w_dff_A_eqLjgLOn4_0),.din(w_dff_A_91W6l9NE5_0),.clk(gclk));
	jdff dff_A_9e2Mw5bp3_0(.dout(w_dff_A_91W6l9NE5_0),.din(w_dff_A_9e2Mw5bp3_0),.clk(gclk));
	jdff dff_A_Bulf4hA77_0(.dout(w_dff_A_9e2Mw5bp3_0),.din(w_dff_A_Bulf4hA77_0),.clk(gclk));
	jdff dff_A_7HAxMaP98_0(.dout(w_dff_A_Bulf4hA77_0),.din(w_dff_A_7HAxMaP98_0),.clk(gclk));
	jdff dff_A_53WWlr557_0(.dout(w_dff_A_7HAxMaP98_0),.din(w_dff_A_53WWlr557_0),.clk(gclk));
	jdff dff_A_VJ9VPnRZ1_0(.dout(w_dff_A_53WWlr557_0),.din(w_dff_A_VJ9VPnRZ1_0),.clk(gclk));
	jdff dff_A_1mR2f2WZ5_0(.dout(w_dff_A_VJ9VPnRZ1_0),.din(w_dff_A_1mR2f2WZ5_0),.clk(gclk));
	jdff dff_A_pAYbq8Wm4_0(.dout(w_dff_A_1mR2f2WZ5_0),.din(w_dff_A_pAYbq8Wm4_0),.clk(gclk));
	jdff dff_A_vpfnu7Zo2_0(.dout(w_dff_A_pAYbq8Wm4_0),.din(w_dff_A_vpfnu7Zo2_0),.clk(gclk));
	jdff dff_A_8QmlS4kl5_0(.dout(w_dff_A_vpfnu7Zo2_0),.din(w_dff_A_8QmlS4kl5_0),.clk(gclk));
	jdff dff_A_YVshM2O80_0(.dout(w_dff_A_8QmlS4kl5_0),.din(w_dff_A_YVshM2O80_0),.clk(gclk));
	jdff dff_A_BbvnutCV7_0(.dout(w_dff_A_YVshM2O80_0),.din(w_dff_A_BbvnutCV7_0),.clk(gclk));
	jdff dff_A_9bNkaOUZ7_0(.dout(w_dff_A_BbvnutCV7_0),.din(w_dff_A_9bNkaOUZ7_0),.clk(gclk));
	jdff dff_A_3Z9gBS8J2_0(.dout(w_dff_A_9bNkaOUZ7_0),.din(w_dff_A_3Z9gBS8J2_0),.clk(gclk));
	jdff dff_A_QyYqNGcL2_0(.dout(w_dff_A_3Z9gBS8J2_0),.din(w_dff_A_QyYqNGcL2_0),.clk(gclk));
	jdff dff_A_y52OnWIm4_1(.dout(w_n547_0[1]),.din(w_dff_A_y52OnWIm4_1),.clk(gclk));
	jdff dff_B_03OhajKk6_1(.din(n478),.dout(w_dff_B_03OhajKk6_1),.clk(gclk));
	jdff dff_B_78yyYrFy9_1(.din(w_dff_B_03OhajKk6_1),.dout(w_dff_B_78yyYrFy9_1),.clk(gclk));
	jdff dff_B_gP9qIGun5_1(.din(w_dff_B_78yyYrFy9_1),.dout(w_dff_B_gP9qIGun5_1),.clk(gclk));
	jdff dff_B_a0D0ATka5_1(.din(w_dff_B_gP9qIGun5_1),.dout(w_dff_B_a0D0ATka5_1),.clk(gclk));
	jdff dff_B_r5GjRDuH9_1(.din(w_dff_B_a0D0ATka5_1),.dout(w_dff_B_r5GjRDuH9_1),.clk(gclk));
	jdff dff_B_uyfJ7Mt46_1(.din(w_dff_B_r5GjRDuH9_1),.dout(w_dff_B_uyfJ7Mt46_1),.clk(gclk));
	jdff dff_B_vEwSBPt70_1(.din(w_dff_B_uyfJ7Mt46_1),.dout(w_dff_B_vEwSBPt70_1),.clk(gclk));
	jdff dff_B_shnxaGXY8_1(.din(w_dff_B_vEwSBPt70_1),.dout(w_dff_B_shnxaGXY8_1),.clk(gclk));
	jdff dff_B_sjrSdDmm3_1(.din(w_dff_B_shnxaGXY8_1),.dout(w_dff_B_sjrSdDmm3_1),.clk(gclk));
	jdff dff_B_WpSDGyFr8_1(.din(w_dff_B_sjrSdDmm3_1),.dout(w_dff_B_WpSDGyFr8_1),.clk(gclk));
	jdff dff_B_YSayJaUO7_1(.din(w_dff_B_WpSDGyFr8_1),.dout(w_dff_B_YSayJaUO7_1),.clk(gclk));
	jdff dff_B_L1y1wUmA7_1(.din(w_dff_B_YSayJaUO7_1),.dout(w_dff_B_L1y1wUmA7_1),.clk(gclk));
	jdff dff_B_DhnnIlKP4_1(.din(w_dff_B_L1y1wUmA7_1),.dout(w_dff_B_DhnnIlKP4_1),.clk(gclk));
	jdff dff_B_aPPAH2Ah1_1(.din(w_dff_B_DhnnIlKP4_1),.dout(w_dff_B_aPPAH2Ah1_1),.clk(gclk));
	jdff dff_B_CbCL1So65_1(.din(w_dff_B_aPPAH2Ah1_1),.dout(w_dff_B_CbCL1So65_1),.clk(gclk));
	jdff dff_B_tF0PQgSd6_1(.din(w_dff_B_CbCL1So65_1),.dout(w_dff_B_tF0PQgSd6_1),.clk(gclk));
	jdff dff_B_W1EZMm6m4_1(.din(w_dff_B_tF0PQgSd6_1),.dout(w_dff_B_W1EZMm6m4_1),.clk(gclk));
	jdff dff_B_HBH1vVDM0_1(.din(w_dff_B_W1EZMm6m4_1),.dout(w_dff_B_HBH1vVDM0_1),.clk(gclk));
	jdff dff_B_GobGod4P7_1(.din(w_dff_B_HBH1vVDM0_1),.dout(w_dff_B_GobGod4P7_1),.clk(gclk));
	jdff dff_B_lg1clGu56_1(.din(w_dff_B_GobGod4P7_1),.dout(w_dff_B_lg1clGu56_1),.clk(gclk));
	jdff dff_B_VGX2ImSY9_1(.din(w_dff_B_lg1clGu56_1),.dout(w_dff_B_VGX2ImSY9_1),.clk(gclk));
	jdff dff_B_old76uYA3_1(.din(w_dff_B_VGX2ImSY9_1),.dout(w_dff_B_old76uYA3_1),.clk(gclk));
	jdff dff_B_WLCDqwmH1_1(.din(w_dff_B_old76uYA3_1),.dout(w_dff_B_WLCDqwmH1_1),.clk(gclk));
	jdff dff_B_OiiVPp338_1(.din(w_dff_B_WLCDqwmH1_1),.dout(w_dff_B_OiiVPp338_1),.clk(gclk));
	jdff dff_B_TzjhTPpi6_1(.din(w_dff_B_OiiVPp338_1),.dout(w_dff_B_TzjhTPpi6_1),.clk(gclk));
	jdff dff_B_SMsTbFdw7_1(.din(w_dff_B_TzjhTPpi6_1),.dout(w_dff_B_SMsTbFdw7_1),.clk(gclk));
	jdff dff_B_rrKbl2Oz7_1(.din(w_dff_B_SMsTbFdw7_1),.dout(w_dff_B_rrKbl2Oz7_1),.clk(gclk));
	jdff dff_B_9nDqJSLu7_1(.din(w_dff_B_rrKbl2Oz7_1),.dout(w_dff_B_9nDqJSLu7_1),.clk(gclk));
	jdff dff_B_DQfbDQM90_1(.din(n474),.dout(w_dff_B_DQfbDQM90_1),.clk(gclk));
	jdff dff_A_koecHf197_0(.dout(w_n399_0[0]),.din(w_dff_A_koecHf197_0),.clk(gclk));
	jdff dff_A_88of4Y3H2_0(.dout(w_dff_A_koecHf197_0),.din(w_dff_A_88of4Y3H2_0),.clk(gclk));
	jdff dff_A_zUKI2ipk6_0(.dout(w_dff_A_88of4Y3H2_0),.din(w_dff_A_zUKI2ipk6_0),.clk(gclk));
	jdff dff_A_Mg1QMq1y0_0(.dout(w_dff_A_zUKI2ipk6_0),.din(w_dff_A_Mg1QMq1y0_0),.clk(gclk));
	jdff dff_A_KO8gUpMt8_0(.dout(w_dff_A_Mg1QMq1y0_0),.din(w_dff_A_KO8gUpMt8_0),.clk(gclk));
	jdff dff_A_bZyjf5QM0_0(.dout(w_dff_A_KO8gUpMt8_0),.din(w_dff_A_bZyjf5QM0_0),.clk(gclk));
	jdff dff_A_Jp87AN728_0(.dout(w_dff_A_bZyjf5QM0_0),.din(w_dff_A_Jp87AN728_0),.clk(gclk));
	jdff dff_A_Vw0XLAzK7_0(.dout(w_dff_A_Jp87AN728_0),.din(w_dff_A_Vw0XLAzK7_0),.clk(gclk));
	jdff dff_A_j1sNWFGB9_0(.dout(w_dff_A_Vw0XLAzK7_0),.din(w_dff_A_j1sNWFGB9_0),.clk(gclk));
	jdff dff_A_nX2OLA8t1_0(.dout(w_dff_A_j1sNWFGB9_0),.din(w_dff_A_nX2OLA8t1_0),.clk(gclk));
	jdff dff_A_3bBkmYjL4_0(.dout(w_dff_A_nX2OLA8t1_0),.din(w_dff_A_3bBkmYjL4_0),.clk(gclk));
	jdff dff_A_GeiHwEMD0_0(.dout(w_dff_A_3bBkmYjL4_0),.din(w_dff_A_GeiHwEMD0_0),.clk(gclk));
	jdff dff_A_WZnIHl6l9_0(.dout(w_dff_A_GeiHwEMD0_0),.din(w_dff_A_WZnIHl6l9_0),.clk(gclk));
	jdff dff_A_p5kFz4gF7_0(.dout(w_dff_A_WZnIHl6l9_0),.din(w_dff_A_p5kFz4gF7_0),.clk(gclk));
	jdff dff_A_sx8ig0DO6_0(.dout(w_dff_A_p5kFz4gF7_0),.din(w_dff_A_sx8ig0DO6_0),.clk(gclk));
	jdff dff_A_mYZKCLuz6_0(.dout(w_dff_A_sx8ig0DO6_0),.din(w_dff_A_mYZKCLuz6_0),.clk(gclk));
	jdff dff_A_1oFOzSW69_0(.dout(w_dff_A_mYZKCLuz6_0),.din(w_dff_A_1oFOzSW69_0),.clk(gclk));
	jdff dff_A_uGPvtTVX7_0(.dout(w_dff_A_1oFOzSW69_0),.din(w_dff_A_uGPvtTVX7_0),.clk(gclk));
	jdff dff_A_zZu1xyvL2_0(.dout(w_dff_A_uGPvtTVX7_0),.din(w_dff_A_zZu1xyvL2_0),.clk(gclk));
	jdff dff_A_VybmS4eT2_0(.dout(w_dff_A_zZu1xyvL2_0),.din(w_dff_A_VybmS4eT2_0),.clk(gclk));
	jdff dff_A_j5yhgpTH9_0(.dout(w_dff_A_VybmS4eT2_0),.din(w_dff_A_j5yhgpTH9_0),.clk(gclk));
	jdff dff_A_VW0iDvQY7_0(.dout(w_dff_A_j5yhgpTH9_0),.din(w_dff_A_VW0iDvQY7_0),.clk(gclk));
	jdff dff_A_lVUI89H38_0(.dout(w_dff_A_VW0iDvQY7_0),.din(w_dff_A_lVUI89H38_0),.clk(gclk));
	jdff dff_A_vcBEXZuq6_0(.dout(w_dff_A_lVUI89H38_0),.din(w_dff_A_vcBEXZuq6_0),.clk(gclk));
	jdff dff_A_QF69uTUZ8_0(.dout(w_dff_A_vcBEXZuq6_0),.din(w_dff_A_QF69uTUZ8_0),.clk(gclk));
	jdff dff_A_iaD0Ui6t2_0(.dout(w_dff_A_QF69uTUZ8_0),.din(w_dff_A_iaD0Ui6t2_0),.clk(gclk));
	jdff dff_A_E4NDaTF07_0(.dout(w_dff_A_iaD0Ui6t2_0),.din(w_dff_A_E4NDaTF07_0),.clk(gclk));
	jdff dff_A_3CQsH5Ge1_0(.dout(w_dff_A_E4NDaTF07_0),.din(w_dff_A_3CQsH5Ge1_0),.clk(gclk));
	jdff dff_A_Bh1ZRL9E6_0(.dout(w_dff_A_3CQsH5Ge1_0),.din(w_dff_A_Bh1ZRL9E6_0),.clk(gclk));
	jdff dff_A_CjzJvrro2_1(.dout(w_n468_0[1]),.din(w_dff_A_CjzJvrro2_1),.clk(gclk));
	jdff dff_B_jPf9d1437_1(.din(n406),.dout(w_dff_B_jPf9d1437_1),.clk(gclk));
	jdff dff_B_PMZhOHfG5_1(.din(w_dff_B_jPf9d1437_1),.dout(w_dff_B_PMZhOHfG5_1),.clk(gclk));
	jdff dff_B_7m5Ljs6L5_1(.din(w_dff_B_PMZhOHfG5_1),.dout(w_dff_B_7m5Ljs6L5_1),.clk(gclk));
	jdff dff_B_91Eq0bsZ1_1(.din(w_dff_B_7m5Ljs6L5_1),.dout(w_dff_B_91Eq0bsZ1_1),.clk(gclk));
	jdff dff_B_caNJuHBv3_1(.din(w_dff_B_91Eq0bsZ1_1),.dout(w_dff_B_caNJuHBv3_1),.clk(gclk));
	jdff dff_B_uq5XLDR71_1(.din(w_dff_B_caNJuHBv3_1),.dout(w_dff_B_uq5XLDR71_1),.clk(gclk));
	jdff dff_B_7sdbKtDC6_1(.din(w_dff_B_uq5XLDR71_1),.dout(w_dff_B_7sdbKtDC6_1),.clk(gclk));
	jdff dff_B_Hhdpf7DE2_1(.din(w_dff_B_7sdbKtDC6_1),.dout(w_dff_B_Hhdpf7DE2_1),.clk(gclk));
	jdff dff_B_6UqegZxt9_1(.din(w_dff_B_Hhdpf7DE2_1),.dout(w_dff_B_6UqegZxt9_1),.clk(gclk));
	jdff dff_B_sU8svXl31_1(.din(w_dff_B_6UqegZxt9_1),.dout(w_dff_B_sU8svXl31_1),.clk(gclk));
	jdff dff_B_Stgp5cb35_1(.din(w_dff_B_sU8svXl31_1),.dout(w_dff_B_Stgp5cb35_1),.clk(gclk));
	jdff dff_B_qngqHhWW7_1(.din(w_dff_B_Stgp5cb35_1),.dout(w_dff_B_qngqHhWW7_1),.clk(gclk));
	jdff dff_B_tZVYjBeh0_1(.din(w_dff_B_qngqHhWW7_1),.dout(w_dff_B_tZVYjBeh0_1),.clk(gclk));
	jdff dff_B_Ar81sFvH3_1(.din(w_dff_B_tZVYjBeh0_1),.dout(w_dff_B_Ar81sFvH3_1),.clk(gclk));
	jdff dff_B_3P3blIMd6_1(.din(w_dff_B_Ar81sFvH3_1),.dout(w_dff_B_3P3blIMd6_1),.clk(gclk));
	jdff dff_B_tGnemvza7_1(.din(w_dff_B_3P3blIMd6_1),.dout(w_dff_B_tGnemvza7_1),.clk(gclk));
	jdff dff_B_TSPrvUGD6_1(.din(w_dff_B_tGnemvza7_1),.dout(w_dff_B_TSPrvUGD6_1),.clk(gclk));
	jdff dff_B_FdpkVCvy7_1(.din(w_dff_B_TSPrvUGD6_1),.dout(w_dff_B_FdpkVCvy7_1),.clk(gclk));
	jdff dff_B_cLibVtUJ7_1(.din(w_dff_B_FdpkVCvy7_1),.dout(w_dff_B_cLibVtUJ7_1),.clk(gclk));
	jdff dff_B_hra5wWkj4_1(.din(w_dff_B_cLibVtUJ7_1),.dout(w_dff_B_hra5wWkj4_1),.clk(gclk));
	jdff dff_B_L4Z2YD5P5_1(.din(w_dff_B_hra5wWkj4_1),.dout(w_dff_B_L4Z2YD5P5_1),.clk(gclk));
	jdff dff_B_zBbDLL0r2_1(.din(w_dff_B_L4Z2YD5P5_1),.dout(w_dff_B_zBbDLL0r2_1),.clk(gclk));
	jdff dff_B_V8cBGbxW4_1(.din(w_dff_B_zBbDLL0r2_1),.dout(w_dff_B_V8cBGbxW4_1),.clk(gclk));
	jdff dff_B_cUpVF8kC7_1(.din(w_dff_B_V8cBGbxW4_1),.dout(w_dff_B_cUpVF8kC7_1),.clk(gclk));
	jdff dff_B_wop3Ppbk9_1(.din(w_dff_B_cUpVF8kC7_1),.dout(w_dff_B_wop3Ppbk9_1),.clk(gclk));
	jdff dff_B_ZBjdgUM75_1(.din(n402),.dout(w_dff_B_ZBjdgUM75_1),.clk(gclk));
	jdff dff_A_4yTvoOGG4_0(.dout(w_n335_0[0]),.din(w_dff_A_4yTvoOGG4_0),.clk(gclk));
	jdff dff_A_f4aJ6Dam8_0(.dout(w_dff_A_4yTvoOGG4_0),.din(w_dff_A_f4aJ6Dam8_0),.clk(gclk));
	jdff dff_A_lH0gg2iX6_0(.dout(w_dff_A_f4aJ6Dam8_0),.din(w_dff_A_lH0gg2iX6_0),.clk(gclk));
	jdff dff_A_zUAKggiq6_0(.dout(w_dff_A_lH0gg2iX6_0),.din(w_dff_A_zUAKggiq6_0),.clk(gclk));
	jdff dff_A_vNUFrGXP7_0(.dout(w_dff_A_zUAKggiq6_0),.din(w_dff_A_vNUFrGXP7_0),.clk(gclk));
	jdff dff_A_UfxBdeRD1_0(.dout(w_dff_A_vNUFrGXP7_0),.din(w_dff_A_UfxBdeRD1_0),.clk(gclk));
	jdff dff_A_VdQzMsFY8_0(.dout(w_dff_A_UfxBdeRD1_0),.din(w_dff_A_VdQzMsFY8_0),.clk(gclk));
	jdff dff_A_GhDlmh643_0(.dout(w_dff_A_VdQzMsFY8_0),.din(w_dff_A_GhDlmh643_0),.clk(gclk));
	jdff dff_A_6B1Ba9kp1_0(.dout(w_dff_A_GhDlmh643_0),.din(w_dff_A_6B1Ba9kp1_0),.clk(gclk));
	jdff dff_A_Orz0hikz5_0(.dout(w_dff_A_6B1Ba9kp1_0),.din(w_dff_A_Orz0hikz5_0),.clk(gclk));
	jdff dff_A_t472kEWT1_0(.dout(w_dff_A_Orz0hikz5_0),.din(w_dff_A_t472kEWT1_0),.clk(gclk));
	jdff dff_A_r2bAcMBp7_0(.dout(w_dff_A_t472kEWT1_0),.din(w_dff_A_r2bAcMBp7_0),.clk(gclk));
	jdff dff_A_kuDJKgVV6_0(.dout(w_dff_A_r2bAcMBp7_0),.din(w_dff_A_kuDJKgVV6_0),.clk(gclk));
	jdff dff_A_4EAKvhJF0_0(.dout(w_dff_A_kuDJKgVV6_0),.din(w_dff_A_4EAKvhJF0_0),.clk(gclk));
	jdff dff_A_ScwgxVOV1_0(.dout(w_dff_A_4EAKvhJF0_0),.din(w_dff_A_ScwgxVOV1_0),.clk(gclk));
	jdff dff_A_xDNSVloW3_0(.dout(w_dff_A_ScwgxVOV1_0),.din(w_dff_A_xDNSVloW3_0),.clk(gclk));
	jdff dff_A_mJ4UpHWR6_0(.dout(w_dff_A_xDNSVloW3_0),.din(w_dff_A_mJ4UpHWR6_0),.clk(gclk));
	jdff dff_A_FQBlAXKf7_0(.dout(w_dff_A_mJ4UpHWR6_0),.din(w_dff_A_FQBlAXKf7_0),.clk(gclk));
	jdff dff_A_2rVn07hh8_0(.dout(w_dff_A_FQBlAXKf7_0),.din(w_dff_A_2rVn07hh8_0),.clk(gclk));
	jdff dff_A_xaaj5BxM3_0(.dout(w_dff_A_2rVn07hh8_0),.din(w_dff_A_xaaj5BxM3_0),.clk(gclk));
	jdff dff_A_ApncF34F8_0(.dout(w_dff_A_xaaj5BxM3_0),.din(w_dff_A_ApncF34F8_0),.clk(gclk));
	jdff dff_A_HfF4ygvD2_0(.dout(w_dff_A_ApncF34F8_0),.din(w_dff_A_HfF4ygvD2_0),.clk(gclk));
	jdff dff_A_TwrHOL4N2_0(.dout(w_dff_A_HfF4ygvD2_0),.din(w_dff_A_TwrHOL4N2_0),.clk(gclk));
	jdff dff_A_WBeW4mnR4_0(.dout(w_dff_A_TwrHOL4N2_0),.din(w_dff_A_WBeW4mnR4_0),.clk(gclk));
	jdff dff_A_f5dVDaYY7_0(.dout(w_dff_A_WBeW4mnR4_0),.din(w_dff_A_f5dVDaYY7_0),.clk(gclk));
	jdff dff_A_t8tAzgMp1_0(.dout(w_dff_A_f5dVDaYY7_0),.din(w_dff_A_t8tAzgMp1_0),.clk(gclk));
	jdff dff_A_CHZGfPAc5_1(.dout(w_n396_0[1]),.din(w_dff_A_CHZGfPAc5_1),.clk(gclk));
	jdff dff_B_uPooh4ko2_1(.din(n342),.dout(w_dff_B_uPooh4ko2_1),.clk(gclk));
	jdff dff_B_jB9bx6RJ4_1(.din(w_dff_B_uPooh4ko2_1),.dout(w_dff_B_jB9bx6RJ4_1),.clk(gclk));
	jdff dff_B_rEj5h7iN0_1(.din(w_dff_B_jB9bx6RJ4_1),.dout(w_dff_B_rEj5h7iN0_1),.clk(gclk));
	jdff dff_B_y2Bpli1n5_1(.din(w_dff_B_rEj5h7iN0_1),.dout(w_dff_B_y2Bpli1n5_1),.clk(gclk));
	jdff dff_B_z1Cb8xDh4_1(.din(w_dff_B_y2Bpli1n5_1),.dout(w_dff_B_z1Cb8xDh4_1),.clk(gclk));
	jdff dff_B_fg0i13d87_1(.din(w_dff_B_z1Cb8xDh4_1),.dout(w_dff_B_fg0i13d87_1),.clk(gclk));
	jdff dff_B_KXGIOptQ6_1(.din(w_dff_B_fg0i13d87_1),.dout(w_dff_B_KXGIOptQ6_1),.clk(gclk));
	jdff dff_B_jcuzs3am8_1(.din(w_dff_B_KXGIOptQ6_1),.dout(w_dff_B_jcuzs3am8_1),.clk(gclk));
	jdff dff_B_mSXkN6kp4_1(.din(w_dff_B_jcuzs3am8_1),.dout(w_dff_B_mSXkN6kp4_1),.clk(gclk));
	jdff dff_B_noNM6B8J1_1(.din(w_dff_B_mSXkN6kp4_1),.dout(w_dff_B_noNM6B8J1_1),.clk(gclk));
	jdff dff_B_O0RoGiIr8_1(.din(w_dff_B_noNM6B8J1_1),.dout(w_dff_B_O0RoGiIr8_1),.clk(gclk));
	jdff dff_B_VDCUgvIi3_1(.din(w_dff_B_O0RoGiIr8_1),.dout(w_dff_B_VDCUgvIi3_1),.clk(gclk));
	jdff dff_B_GnCt8pN18_1(.din(w_dff_B_VDCUgvIi3_1),.dout(w_dff_B_GnCt8pN18_1),.clk(gclk));
	jdff dff_B_V9ew3Jy92_1(.din(w_dff_B_GnCt8pN18_1),.dout(w_dff_B_V9ew3Jy92_1),.clk(gclk));
	jdff dff_B_i0ViKzR78_1(.din(w_dff_B_V9ew3Jy92_1),.dout(w_dff_B_i0ViKzR78_1),.clk(gclk));
	jdff dff_B_6ylNFGro7_1(.din(w_dff_B_i0ViKzR78_1),.dout(w_dff_B_6ylNFGro7_1),.clk(gclk));
	jdff dff_B_ACRkX0KM3_1(.din(w_dff_B_6ylNFGro7_1),.dout(w_dff_B_ACRkX0KM3_1),.clk(gclk));
	jdff dff_B_LZbVOwwh8_1(.din(w_dff_B_ACRkX0KM3_1),.dout(w_dff_B_LZbVOwwh8_1),.clk(gclk));
	jdff dff_B_IH4X7iGM9_1(.din(w_dff_B_LZbVOwwh8_1),.dout(w_dff_B_IH4X7iGM9_1),.clk(gclk));
	jdff dff_B_yu6bXgS87_1(.din(w_dff_B_IH4X7iGM9_1),.dout(w_dff_B_yu6bXgS87_1),.clk(gclk));
	jdff dff_B_k6SXAJtP2_1(.din(w_dff_B_yu6bXgS87_1),.dout(w_dff_B_k6SXAJtP2_1),.clk(gclk));
	jdff dff_B_v1w7e7PW8_1(.din(w_dff_B_k6SXAJtP2_1),.dout(w_dff_B_v1w7e7PW8_1),.clk(gclk));
	jdff dff_B_AjWbN0rr3_1(.din(n338),.dout(w_dff_B_AjWbN0rr3_1),.clk(gclk));
	jdff dff_A_6PiLb6KC4_0(.dout(w_n277_0[0]),.din(w_dff_A_6PiLb6KC4_0),.clk(gclk));
	jdff dff_A_Bb9UfAdB0_0(.dout(w_dff_A_6PiLb6KC4_0),.din(w_dff_A_Bb9UfAdB0_0),.clk(gclk));
	jdff dff_A_HPwUAGCC3_0(.dout(w_dff_A_Bb9UfAdB0_0),.din(w_dff_A_HPwUAGCC3_0),.clk(gclk));
	jdff dff_A_dFCAAs831_0(.dout(w_dff_A_HPwUAGCC3_0),.din(w_dff_A_dFCAAs831_0),.clk(gclk));
	jdff dff_A_Iy9sInHu9_0(.dout(w_dff_A_dFCAAs831_0),.din(w_dff_A_Iy9sInHu9_0),.clk(gclk));
	jdff dff_A_VclKgW8m9_0(.dout(w_dff_A_Iy9sInHu9_0),.din(w_dff_A_VclKgW8m9_0),.clk(gclk));
	jdff dff_A_qI9EW8fy2_0(.dout(w_dff_A_VclKgW8m9_0),.din(w_dff_A_qI9EW8fy2_0),.clk(gclk));
	jdff dff_A_xyJySTWb1_0(.dout(w_dff_A_qI9EW8fy2_0),.din(w_dff_A_xyJySTWb1_0),.clk(gclk));
	jdff dff_A_JSmQBqyU7_0(.dout(w_dff_A_xyJySTWb1_0),.din(w_dff_A_JSmQBqyU7_0),.clk(gclk));
	jdff dff_A_TtAhHQGa5_0(.dout(w_dff_A_JSmQBqyU7_0),.din(w_dff_A_TtAhHQGa5_0),.clk(gclk));
	jdff dff_A_RSrEA1wc2_0(.dout(w_dff_A_TtAhHQGa5_0),.din(w_dff_A_RSrEA1wc2_0),.clk(gclk));
	jdff dff_A_2eu7Rc9D6_0(.dout(w_dff_A_RSrEA1wc2_0),.din(w_dff_A_2eu7Rc9D6_0),.clk(gclk));
	jdff dff_A_ke2CuF9w4_0(.dout(w_dff_A_2eu7Rc9D6_0),.din(w_dff_A_ke2CuF9w4_0),.clk(gclk));
	jdff dff_A_DmWln3eR4_0(.dout(w_dff_A_ke2CuF9w4_0),.din(w_dff_A_DmWln3eR4_0),.clk(gclk));
	jdff dff_A_JLIO5ySW8_0(.dout(w_dff_A_DmWln3eR4_0),.din(w_dff_A_JLIO5ySW8_0),.clk(gclk));
	jdff dff_A_QR3vwlDf0_0(.dout(w_dff_A_JLIO5ySW8_0),.din(w_dff_A_QR3vwlDf0_0),.clk(gclk));
	jdff dff_A_lYlufg023_0(.dout(w_dff_A_QR3vwlDf0_0),.din(w_dff_A_lYlufg023_0),.clk(gclk));
	jdff dff_A_k4nutc9v4_0(.dout(w_dff_A_lYlufg023_0),.din(w_dff_A_k4nutc9v4_0),.clk(gclk));
	jdff dff_A_vpDUgNWM4_0(.dout(w_dff_A_k4nutc9v4_0),.din(w_dff_A_vpDUgNWM4_0),.clk(gclk));
	jdff dff_A_xMXRsrhP8_0(.dout(w_dff_A_vpDUgNWM4_0),.din(w_dff_A_xMXRsrhP8_0),.clk(gclk));
	jdff dff_A_naWIhevA7_0(.dout(w_dff_A_xMXRsrhP8_0),.din(w_dff_A_naWIhevA7_0),.clk(gclk));
	jdff dff_A_V1cu7Egm0_0(.dout(w_dff_A_naWIhevA7_0),.din(w_dff_A_V1cu7Egm0_0),.clk(gclk));
	jdff dff_A_eUbJdN5F3_0(.dout(w_dff_A_V1cu7Egm0_0),.din(w_dff_A_eUbJdN5F3_0),.clk(gclk));
	jdff dff_A_peHk2qng5_1(.dout(w_n332_0[1]),.din(w_dff_A_peHk2qng5_1),.clk(gclk));
	jdff dff_B_3jm1LoUs7_1(.din(n284),.dout(w_dff_B_3jm1LoUs7_1),.clk(gclk));
	jdff dff_B_5OHO6uYD6_1(.din(w_dff_B_3jm1LoUs7_1),.dout(w_dff_B_5OHO6uYD6_1),.clk(gclk));
	jdff dff_B_YdpCmWmt5_1(.din(w_dff_B_5OHO6uYD6_1),.dout(w_dff_B_YdpCmWmt5_1),.clk(gclk));
	jdff dff_B_d2BgRoeI9_1(.din(w_dff_B_YdpCmWmt5_1),.dout(w_dff_B_d2BgRoeI9_1),.clk(gclk));
	jdff dff_B_XfRatf0y3_1(.din(w_dff_B_d2BgRoeI9_1),.dout(w_dff_B_XfRatf0y3_1),.clk(gclk));
	jdff dff_B_zgYCR2wc2_1(.din(w_dff_B_XfRatf0y3_1),.dout(w_dff_B_zgYCR2wc2_1),.clk(gclk));
	jdff dff_B_3nhwhcBJ4_1(.din(w_dff_B_zgYCR2wc2_1),.dout(w_dff_B_3nhwhcBJ4_1),.clk(gclk));
	jdff dff_B_6ETBEvVU5_1(.din(w_dff_B_3nhwhcBJ4_1),.dout(w_dff_B_6ETBEvVU5_1),.clk(gclk));
	jdff dff_B_JKJeDhBx4_1(.din(w_dff_B_6ETBEvVU5_1),.dout(w_dff_B_JKJeDhBx4_1),.clk(gclk));
	jdff dff_B_z2UOf6LZ5_1(.din(w_dff_B_JKJeDhBx4_1),.dout(w_dff_B_z2UOf6LZ5_1),.clk(gclk));
	jdff dff_B_3Tk7LKh01_1(.din(w_dff_B_z2UOf6LZ5_1),.dout(w_dff_B_3Tk7LKh01_1),.clk(gclk));
	jdff dff_B_5MH3Oeh13_1(.din(w_dff_B_3Tk7LKh01_1),.dout(w_dff_B_5MH3Oeh13_1),.clk(gclk));
	jdff dff_B_t99yLnjP3_1(.din(w_dff_B_5MH3Oeh13_1),.dout(w_dff_B_t99yLnjP3_1),.clk(gclk));
	jdff dff_B_ECHD0jid6_1(.din(w_dff_B_t99yLnjP3_1),.dout(w_dff_B_ECHD0jid6_1),.clk(gclk));
	jdff dff_B_lksvYya75_1(.din(w_dff_B_ECHD0jid6_1),.dout(w_dff_B_lksvYya75_1),.clk(gclk));
	jdff dff_B_jqsJEwL29_1(.din(w_dff_B_lksvYya75_1),.dout(w_dff_B_jqsJEwL29_1),.clk(gclk));
	jdff dff_B_g0eg8jXV5_1(.din(w_dff_B_jqsJEwL29_1),.dout(w_dff_B_g0eg8jXV5_1),.clk(gclk));
	jdff dff_B_umj1hFfn6_1(.din(w_dff_B_g0eg8jXV5_1),.dout(w_dff_B_umj1hFfn6_1),.clk(gclk));
	jdff dff_B_U0LQCSR08_1(.din(w_dff_B_umj1hFfn6_1),.dout(w_dff_B_U0LQCSR08_1),.clk(gclk));
	jdff dff_B_pRSP3AEO9_1(.din(n280),.dout(w_dff_B_pRSP3AEO9_1),.clk(gclk));
	jdff dff_A_9DNkYF7O1_0(.dout(w_n226_0[0]),.din(w_dff_A_9DNkYF7O1_0),.clk(gclk));
	jdff dff_A_MTW7eLSF3_0(.dout(w_dff_A_9DNkYF7O1_0),.din(w_dff_A_MTW7eLSF3_0),.clk(gclk));
	jdff dff_A_XOaFlA969_0(.dout(w_dff_A_MTW7eLSF3_0),.din(w_dff_A_XOaFlA969_0),.clk(gclk));
	jdff dff_A_vW6bK1cy4_0(.dout(w_dff_A_XOaFlA969_0),.din(w_dff_A_vW6bK1cy4_0),.clk(gclk));
	jdff dff_A_Db1PgHsM6_0(.dout(w_dff_A_vW6bK1cy4_0),.din(w_dff_A_Db1PgHsM6_0),.clk(gclk));
	jdff dff_A_wXTeGHmP5_0(.dout(w_dff_A_Db1PgHsM6_0),.din(w_dff_A_wXTeGHmP5_0),.clk(gclk));
	jdff dff_A_57S724kv0_0(.dout(w_dff_A_wXTeGHmP5_0),.din(w_dff_A_57S724kv0_0),.clk(gclk));
	jdff dff_A_cHuF6PXi2_0(.dout(w_dff_A_57S724kv0_0),.din(w_dff_A_cHuF6PXi2_0),.clk(gclk));
	jdff dff_A_lIFHSSwv1_0(.dout(w_dff_A_cHuF6PXi2_0),.din(w_dff_A_lIFHSSwv1_0),.clk(gclk));
	jdff dff_A_UW6i24ke9_0(.dout(w_dff_A_lIFHSSwv1_0),.din(w_dff_A_UW6i24ke9_0),.clk(gclk));
	jdff dff_A_hz9fPhRz7_0(.dout(w_dff_A_UW6i24ke9_0),.din(w_dff_A_hz9fPhRz7_0),.clk(gclk));
	jdff dff_A_7RfluJ9C7_0(.dout(w_dff_A_hz9fPhRz7_0),.din(w_dff_A_7RfluJ9C7_0),.clk(gclk));
	jdff dff_A_2CBO0o5u6_0(.dout(w_dff_A_7RfluJ9C7_0),.din(w_dff_A_2CBO0o5u6_0),.clk(gclk));
	jdff dff_A_wPxwHqT10_0(.dout(w_dff_A_2CBO0o5u6_0),.din(w_dff_A_wPxwHqT10_0),.clk(gclk));
	jdff dff_A_TQfBR9oN4_0(.dout(w_dff_A_wPxwHqT10_0),.din(w_dff_A_TQfBR9oN4_0),.clk(gclk));
	jdff dff_A_WyQ6RYTx7_0(.dout(w_dff_A_TQfBR9oN4_0),.din(w_dff_A_WyQ6RYTx7_0),.clk(gclk));
	jdff dff_A_eCWI2sTG8_0(.dout(w_dff_A_WyQ6RYTx7_0),.din(w_dff_A_eCWI2sTG8_0),.clk(gclk));
	jdff dff_A_S0RWZkCc7_0(.dout(w_dff_A_eCWI2sTG8_0),.din(w_dff_A_S0RWZkCc7_0),.clk(gclk));
	jdff dff_A_5eQzsYTy1_0(.dout(w_dff_A_S0RWZkCc7_0),.din(w_dff_A_5eQzsYTy1_0),.clk(gclk));
	jdff dff_A_edGf9AFJ6_0(.dout(w_dff_A_5eQzsYTy1_0),.din(w_dff_A_edGf9AFJ6_0),.clk(gclk));
	jdff dff_A_tZxpkrLk3_1(.dout(w_n274_0[1]),.din(w_dff_A_tZxpkrLk3_1),.clk(gclk));
	jdff dff_B_h6JbXv9q1_1(.din(n233),.dout(w_dff_B_h6JbXv9q1_1),.clk(gclk));
	jdff dff_B_5pF6I5F77_1(.din(w_dff_B_h6JbXv9q1_1),.dout(w_dff_B_5pF6I5F77_1),.clk(gclk));
	jdff dff_B_vVA7RSmo9_1(.din(w_dff_B_5pF6I5F77_1),.dout(w_dff_B_vVA7RSmo9_1),.clk(gclk));
	jdff dff_B_mARE0DzF5_1(.din(w_dff_B_vVA7RSmo9_1),.dout(w_dff_B_mARE0DzF5_1),.clk(gclk));
	jdff dff_B_jZnpDUjS2_1(.din(w_dff_B_mARE0DzF5_1),.dout(w_dff_B_jZnpDUjS2_1),.clk(gclk));
	jdff dff_B_MBIWsY8n5_1(.din(w_dff_B_jZnpDUjS2_1),.dout(w_dff_B_MBIWsY8n5_1),.clk(gclk));
	jdff dff_B_JebC4doU8_1(.din(w_dff_B_MBIWsY8n5_1),.dout(w_dff_B_JebC4doU8_1),.clk(gclk));
	jdff dff_B_0k6QPpgW6_1(.din(w_dff_B_JebC4doU8_1),.dout(w_dff_B_0k6QPpgW6_1),.clk(gclk));
	jdff dff_B_0K1i2wLI0_1(.din(w_dff_B_0k6QPpgW6_1),.dout(w_dff_B_0K1i2wLI0_1),.clk(gclk));
	jdff dff_B_8ETZk4Mc5_1(.din(w_dff_B_0K1i2wLI0_1),.dout(w_dff_B_8ETZk4Mc5_1),.clk(gclk));
	jdff dff_B_DqYHRLOG4_1(.din(w_dff_B_8ETZk4Mc5_1),.dout(w_dff_B_DqYHRLOG4_1),.clk(gclk));
	jdff dff_B_VOnfjZ3w1_1(.din(w_dff_B_DqYHRLOG4_1),.dout(w_dff_B_VOnfjZ3w1_1),.clk(gclk));
	jdff dff_B_k9OxSITD3_1(.din(w_dff_B_VOnfjZ3w1_1),.dout(w_dff_B_k9OxSITD3_1),.clk(gclk));
	jdff dff_B_CjOzhyUA6_1(.din(w_dff_B_k9OxSITD3_1),.dout(w_dff_B_CjOzhyUA6_1),.clk(gclk));
	jdff dff_B_wpjKZvYm1_1(.din(w_dff_B_CjOzhyUA6_1),.dout(w_dff_B_wpjKZvYm1_1),.clk(gclk));
	jdff dff_B_txgUulhx8_1(.din(w_dff_B_wpjKZvYm1_1),.dout(w_dff_B_txgUulhx8_1),.clk(gclk));
	jdff dff_B_rd8mdpko9_1(.din(n229),.dout(w_dff_B_rd8mdpko9_1),.clk(gclk));
	jdff dff_A_jFTrrHOP4_0(.dout(w_n183_0[0]),.din(w_dff_A_jFTrrHOP4_0),.clk(gclk));
	jdff dff_A_HnMp1a7O1_0(.dout(w_dff_A_jFTrrHOP4_0),.din(w_dff_A_HnMp1a7O1_0),.clk(gclk));
	jdff dff_A_QOFFq5fX4_0(.dout(w_dff_A_HnMp1a7O1_0),.din(w_dff_A_QOFFq5fX4_0),.clk(gclk));
	jdff dff_A_YsTdaKn61_0(.dout(w_dff_A_QOFFq5fX4_0),.din(w_dff_A_YsTdaKn61_0),.clk(gclk));
	jdff dff_A_55FDEM2a4_0(.dout(w_dff_A_YsTdaKn61_0),.din(w_dff_A_55FDEM2a4_0),.clk(gclk));
	jdff dff_A_0MrTwIOG1_0(.dout(w_dff_A_55FDEM2a4_0),.din(w_dff_A_0MrTwIOG1_0),.clk(gclk));
	jdff dff_A_wLDUqIBe9_0(.dout(w_dff_A_0MrTwIOG1_0),.din(w_dff_A_wLDUqIBe9_0),.clk(gclk));
	jdff dff_A_GCZtswWN6_0(.dout(w_dff_A_wLDUqIBe9_0),.din(w_dff_A_GCZtswWN6_0),.clk(gclk));
	jdff dff_A_0h0x7GFn7_0(.dout(w_dff_A_GCZtswWN6_0),.din(w_dff_A_0h0x7GFn7_0),.clk(gclk));
	jdff dff_A_kXcckj9G0_0(.dout(w_dff_A_0h0x7GFn7_0),.din(w_dff_A_kXcckj9G0_0),.clk(gclk));
	jdff dff_A_qLW1G1338_0(.dout(w_dff_A_kXcckj9G0_0),.din(w_dff_A_qLW1G1338_0),.clk(gclk));
	jdff dff_A_a3wbc89U7_0(.dout(w_dff_A_qLW1G1338_0),.din(w_dff_A_a3wbc89U7_0),.clk(gclk));
	jdff dff_A_UoZYWiHc9_0(.dout(w_dff_A_a3wbc89U7_0),.din(w_dff_A_UoZYWiHc9_0),.clk(gclk));
	jdff dff_A_HDQ0hPqB8_0(.dout(w_dff_A_UoZYWiHc9_0),.din(w_dff_A_HDQ0hPqB8_0),.clk(gclk));
	jdff dff_A_SJPEAaCf7_0(.dout(w_dff_A_HDQ0hPqB8_0),.din(w_dff_A_SJPEAaCf7_0),.clk(gclk));
	jdff dff_A_OV18yayR5_0(.dout(w_dff_A_SJPEAaCf7_0),.din(w_dff_A_OV18yayR5_0),.clk(gclk));
	jdff dff_A_Ond58uNP5_0(.dout(w_dff_A_OV18yayR5_0),.din(w_dff_A_Ond58uNP5_0),.clk(gclk));
	jdff dff_A_iWmMC9ts3_1(.dout(w_n223_0[1]),.din(w_dff_A_iWmMC9ts3_1),.clk(gclk));
	jdff dff_B_bbmCodpv9_1(.din(n190),.dout(w_dff_B_bbmCodpv9_1),.clk(gclk));
	jdff dff_B_T3DLMfQa1_1(.din(w_dff_B_bbmCodpv9_1),.dout(w_dff_B_T3DLMfQa1_1),.clk(gclk));
	jdff dff_B_ZGze8S695_1(.din(w_dff_B_T3DLMfQa1_1),.dout(w_dff_B_ZGze8S695_1),.clk(gclk));
	jdff dff_B_KelZoE8Z9_1(.din(w_dff_B_ZGze8S695_1),.dout(w_dff_B_KelZoE8Z9_1),.clk(gclk));
	jdff dff_B_WZqPo0yc3_1(.din(w_dff_B_KelZoE8Z9_1),.dout(w_dff_B_WZqPo0yc3_1),.clk(gclk));
	jdff dff_B_u1qfyp3f0_1(.din(w_dff_B_WZqPo0yc3_1),.dout(w_dff_B_u1qfyp3f0_1),.clk(gclk));
	jdff dff_B_VZCzrF6J2_1(.din(w_dff_B_u1qfyp3f0_1),.dout(w_dff_B_VZCzrF6J2_1),.clk(gclk));
	jdff dff_B_ld2M7Io84_1(.din(w_dff_B_VZCzrF6J2_1),.dout(w_dff_B_ld2M7Io84_1),.clk(gclk));
	jdff dff_B_ej3hterM9_1(.din(w_dff_B_ld2M7Io84_1),.dout(w_dff_B_ej3hterM9_1),.clk(gclk));
	jdff dff_B_BNA27gul1_1(.din(w_dff_B_ej3hterM9_1),.dout(w_dff_B_BNA27gul1_1),.clk(gclk));
	jdff dff_B_1dBIy7716_1(.din(w_dff_B_BNA27gul1_1),.dout(w_dff_B_1dBIy7716_1),.clk(gclk));
	jdff dff_B_9B6EDUzt7_1(.din(w_dff_B_1dBIy7716_1),.dout(w_dff_B_9B6EDUzt7_1),.clk(gclk));
	jdff dff_B_AmcbYULr1_1(.din(w_dff_B_9B6EDUzt7_1),.dout(w_dff_B_AmcbYULr1_1),.clk(gclk));
	jdff dff_B_AwKqnTL31_1(.din(n186),.dout(w_dff_B_AwKqnTL31_1),.clk(gclk));
	jdff dff_A_DJjqOhdm7_0(.dout(w_n145_0[0]),.din(w_dff_A_DJjqOhdm7_0),.clk(gclk));
	jdff dff_A_YvHKOKcx4_0(.dout(w_dff_A_DJjqOhdm7_0),.din(w_dff_A_YvHKOKcx4_0),.clk(gclk));
	jdff dff_A_eVvSIuyt5_0(.dout(w_dff_A_YvHKOKcx4_0),.din(w_dff_A_eVvSIuyt5_0),.clk(gclk));
	jdff dff_A_TroSCxah7_0(.dout(w_dff_A_eVvSIuyt5_0),.din(w_dff_A_TroSCxah7_0),.clk(gclk));
	jdff dff_A_9WzLxNoc4_0(.dout(w_dff_A_TroSCxah7_0),.din(w_dff_A_9WzLxNoc4_0),.clk(gclk));
	jdff dff_A_0DsPOaC91_0(.dout(w_dff_A_9WzLxNoc4_0),.din(w_dff_A_0DsPOaC91_0),.clk(gclk));
	jdff dff_A_SUaqs6Qk8_0(.dout(w_dff_A_0DsPOaC91_0),.din(w_dff_A_SUaqs6Qk8_0),.clk(gclk));
	jdff dff_A_vedmNpOY1_0(.dout(w_dff_A_SUaqs6Qk8_0),.din(w_dff_A_vedmNpOY1_0),.clk(gclk));
	jdff dff_A_hzU4Gapk7_0(.dout(w_dff_A_vedmNpOY1_0),.din(w_dff_A_hzU4Gapk7_0),.clk(gclk));
	jdff dff_A_DU3UOxV42_0(.dout(w_dff_A_hzU4Gapk7_0),.din(w_dff_A_DU3UOxV42_0),.clk(gclk));
	jdff dff_A_9hV77ayo2_0(.dout(w_dff_A_DU3UOxV42_0),.din(w_dff_A_9hV77ayo2_0),.clk(gclk));
	jdff dff_A_T6AGU7rH3_0(.dout(w_dff_A_9hV77ayo2_0),.din(w_dff_A_T6AGU7rH3_0),.clk(gclk));
	jdff dff_A_CCzX6Ho66_0(.dout(w_dff_A_T6AGU7rH3_0),.din(w_dff_A_CCzX6Ho66_0),.clk(gclk));
	jdff dff_A_0h3CobnG1_0(.dout(w_dff_A_CCzX6Ho66_0),.din(w_dff_A_0h3CobnG1_0),.clk(gclk));
	jdff dff_A_kqbN4kqC7_1(.dout(w_n180_0[1]),.din(w_dff_A_kqbN4kqC7_1),.clk(gclk));
	jdff dff_B_WDHxITla2_1(.din(n152),.dout(w_dff_B_WDHxITla2_1),.clk(gclk));
	jdff dff_B_YHInVKxR8_1(.din(w_dff_B_WDHxITla2_1),.dout(w_dff_B_YHInVKxR8_1),.clk(gclk));
	jdff dff_B_zeOKIsAd7_1(.din(w_dff_B_YHInVKxR8_1),.dout(w_dff_B_zeOKIsAd7_1),.clk(gclk));
	jdff dff_B_fdAkYsbd6_1(.din(w_dff_B_zeOKIsAd7_1),.dout(w_dff_B_fdAkYsbd6_1),.clk(gclk));
	jdff dff_B_rndcK6l50_1(.din(w_dff_B_fdAkYsbd6_1),.dout(w_dff_B_rndcK6l50_1),.clk(gclk));
	jdff dff_B_5Mq1T8Oi4_1(.din(w_dff_B_rndcK6l50_1),.dout(w_dff_B_5Mq1T8Oi4_1),.clk(gclk));
	jdff dff_B_nBl7lXVE3_1(.din(w_dff_B_5Mq1T8Oi4_1),.dout(w_dff_B_nBl7lXVE3_1),.clk(gclk));
	jdff dff_B_EdRrC5GC0_1(.din(w_dff_B_nBl7lXVE3_1),.dout(w_dff_B_EdRrC5GC0_1),.clk(gclk));
	jdff dff_B_0vCdFfoY2_1(.din(w_dff_B_EdRrC5GC0_1),.dout(w_dff_B_0vCdFfoY2_1),.clk(gclk));
	jdff dff_B_Y7QU2Ebk7_1(.din(w_dff_B_0vCdFfoY2_1),.dout(w_dff_B_Y7QU2Ebk7_1),.clk(gclk));
	jdff dff_B_TKqaCuwG8_1(.din(n148),.dout(w_dff_B_TKqaCuwG8_1),.clk(gclk));
	jdff dff_A_8kpIdcK42_0(.dout(w_n110_0[0]),.din(w_dff_A_8kpIdcK42_0),.clk(gclk));
	jdff dff_A_8D7AhApE5_0(.dout(w_dff_A_8kpIdcK42_0),.din(w_dff_A_8D7AhApE5_0),.clk(gclk));
	jdff dff_A_h55Xr0L76_0(.dout(w_dff_A_8D7AhApE5_0),.din(w_dff_A_h55Xr0L76_0),.clk(gclk));
	jdff dff_A_BcyEWGfB6_0(.dout(w_dff_A_h55Xr0L76_0),.din(w_dff_A_BcyEWGfB6_0),.clk(gclk));
	jdff dff_A_uo5N9op78_0(.dout(w_dff_A_BcyEWGfB6_0),.din(w_dff_A_uo5N9op78_0),.clk(gclk));
	jdff dff_A_22USeGXd2_0(.dout(w_dff_A_uo5N9op78_0),.din(w_dff_A_22USeGXd2_0),.clk(gclk));
	jdff dff_A_HducLP3S1_0(.dout(w_dff_A_22USeGXd2_0),.din(w_dff_A_HducLP3S1_0),.clk(gclk));
	jdff dff_A_NOebkhnB5_0(.dout(w_dff_A_HducLP3S1_0),.din(w_dff_A_NOebkhnB5_0),.clk(gclk));
	jdff dff_A_zww6rqlG3_0(.dout(w_dff_A_NOebkhnB5_0),.din(w_dff_A_zww6rqlG3_0),.clk(gclk));
	jdff dff_A_r6DPxvsI5_0(.dout(w_dff_A_zww6rqlG3_0),.din(w_dff_A_r6DPxvsI5_0),.clk(gclk));
	jdff dff_A_Tooep5n49_0(.dout(w_dff_A_r6DPxvsI5_0),.din(w_dff_A_Tooep5n49_0),.clk(gclk));
	jdff dff_A_VpV1Wt6x7_1(.dout(w_n142_0[1]),.din(w_dff_A_VpV1Wt6x7_1),.clk(gclk));
	jdff dff_B_FxJTXI7R9_1(.din(n117),.dout(w_dff_B_FxJTXI7R9_1),.clk(gclk));
	jdff dff_B_y8vDRHA60_1(.din(w_dff_B_FxJTXI7R9_1),.dout(w_dff_B_y8vDRHA60_1),.clk(gclk));
	jdff dff_B_63Slu4xQ8_1(.din(w_dff_B_y8vDRHA60_1),.dout(w_dff_B_63Slu4xQ8_1),.clk(gclk));
	jdff dff_B_Rf2K9rdr8_1(.din(w_dff_B_63Slu4xQ8_1),.dout(w_dff_B_Rf2K9rdr8_1),.clk(gclk));
	jdff dff_B_42yb08Af2_1(.din(w_dff_B_Rf2K9rdr8_1),.dout(w_dff_B_42yb08Af2_1),.clk(gclk));
	jdff dff_B_19nrQdrO5_1(.din(w_dff_B_42yb08Af2_1),.dout(w_dff_B_19nrQdrO5_1),.clk(gclk));
	jdff dff_B_tBHNWRrm0_1(.din(w_dff_B_19nrQdrO5_1),.dout(w_dff_B_tBHNWRrm0_1),.clk(gclk));
	jdff dff_B_1qvD8ff13_1(.din(n113),.dout(w_dff_B_1qvD8ff13_1),.clk(gclk));
	jdff dff_A_dTyP0f7L8_0(.dout(w_n89_0[0]),.din(w_dff_A_dTyP0f7L8_0),.clk(gclk));
	jdff dff_A_bV00JtyD4_0(.dout(w_dff_A_dTyP0f7L8_0),.din(w_dff_A_bV00JtyD4_0),.clk(gclk));
	jdff dff_A_U1trpJOS5_0(.dout(w_dff_A_bV00JtyD4_0),.din(w_dff_A_U1trpJOS5_0),.clk(gclk));
	jdff dff_A_ePo85IVu4_0(.dout(w_dff_A_U1trpJOS5_0),.din(w_dff_A_ePo85IVu4_0),.clk(gclk));
	jdff dff_A_ruNAtg1E0_0(.dout(w_dff_A_ePo85IVu4_0),.din(w_dff_A_ruNAtg1E0_0),.clk(gclk));
	jdff dff_A_aYd37mFd2_0(.dout(w_dff_A_ruNAtg1E0_0),.din(w_dff_A_aYd37mFd2_0),.clk(gclk));
	jdff dff_A_BE4QZEcY8_0(.dout(w_dff_A_aYd37mFd2_0),.din(w_dff_A_BE4QZEcY8_0),.clk(gclk));
	jdff dff_A_JUvwpQwb8_0(.dout(w_dff_A_BE4QZEcY8_0),.din(w_dff_A_JUvwpQwb8_0),.clk(gclk));
	jdff dff_A_YXMU8p9c8_1(.dout(w_n107_0[1]),.din(w_dff_A_YXMU8p9c8_1),.clk(gclk));
	jdff dff_B_6LZmB3Gn3_1(.din(n95),.dout(w_dff_B_6LZmB3Gn3_1),.clk(gclk));
	jdff dff_B_012J1un06_1(.din(w_dff_B_6LZmB3Gn3_1),.dout(w_dff_B_012J1un06_1),.clk(gclk));
	jdff dff_B_OxwRlb8w7_1(.din(w_dff_B_012J1un06_1),.dout(w_dff_B_OxwRlb8w7_1),.clk(gclk));
	jdff dff_B_jffWmVSl8_1(.din(w_dff_B_OxwRlb8w7_1),.dout(w_dff_B_jffWmVSl8_1),.clk(gclk));
	jdff dff_B_GUp30YFz8_1(.din(n91),.dout(w_dff_B_GUp30YFz8_1),.clk(gclk));
	jdff dff_B_CNllXBTv4_0(.din(n86),.dout(w_dff_B_CNllXBTv4_0),.clk(gclk));
	jdff dff_A_gix6zsfO9_0(.dout(w_n72_0[0]),.din(w_dff_A_gix6zsfO9_0),.clk(gclk));
	jdff dff_A_IN8XLFiq7_0(.dout(w_dff_A_gix6zsfO9_0),.din(w_dff_A_IN8XLFiq7_0),.clk(gclk));
	jdff dff_A_OgaaY1J50_0(.dout(w_dff_A_IN8XLFiq7_0),.din(w_dff_A_OgaaY1J50_0),.clk(gclk));
	jdff dff_A_FLj6H75i3_0(.dout(w_dff_A_OgaaY1J50_0),.din(w_dff_A_FLj6H75i3_0),.clk(gclk));
	jdff dff_A_MuhjVLNl5_0(.dout(w_dff_A_FLj6H75i3_0),.din(w_dff_A_MuhjVLNl5_0),.clk(gclk));
	jdff dff_A_nYOTDYLC5_0(.dout(w_n70_0[0]),.din(w_dff_A_nYOTDYLC5_0),.clk(gclk));
	jdff dff_A_uhOhIG0A7_0(.dout(w_n69_0[0]),.din(w_dff_A_uhOhIG0A7_0),.clk(gclk));
	jdff dff_A_HyISg1en7_1(.dout(w_n1140_0[1]),.din(w_dff_A_HyISg1en7_1),.clk(gclk));
	jdff dff_B_oFoXuBJi1_1(.din(n1040),.dout(w_dff_B_oFoXuBJi1_1),.clk(gclk));
	jdff dff_B_uu5s7mxV8_2(.din(n938),.dout(w_dff_B_uu5s7mxV8_2),.clk(gclk));
	jdff dff_B_RrcJzKsF4_2(.din(w_dff_B_uu5s7mxV8_2),.dout(w_dff_B_RrcJzKsF4_2),.clk(gclk));
	jdff dff_B_RM9G0PvZ0_2(.din(w_dff_B_RrcJzKsF4_2),.dout(w_dff_B_RM9G0PvZ0_2),.clk(gclk));
	jdff dff_B_s4PasYeV7_2(.din(w_dff_B_RM9G0PvZ0_2),.dout(w_dff_B_s4PasYeV7_2),.clk(gclk));
	jdff dff_B_vxw4WpAf9_2(.din(w_dff_B_s4PasYeV7_2),.dout(w_dff_B_vxw4WpAf9_2),.clk(gclk));
	jdff dff_B_CIWvcv9n0_2(.din(w_dff_B_vxw4WpAf9_2),.dout(w_dff_B_CIWvcv9n0_2),.clk(gclk));
	jdff dff_B_zrqvvdgs2_2(.din(w_dff_B_CIWvcv9n0_2),.dout(w_dff_B_zrqvvdgs2_2),.clk(gclk));
	jdff dff_B_ibP34pDL5_2(.din(w_dff_B_zrqvvdgs2_2),.dout(w_dff_B_ibP34pDL5_2),.clk(gclk));
	jdff dff_B_KvdxSQg76_2(.din(w_dff_B_ibP34pDL5_2),.dout(w_dff_B_KvdxSQg76_2),.clk(gclk));
	jdff dff_B_qS1V03CX0_2(.din(w_dff_B_KvdxSQg76_2),.dout(w_dff_B_qS1V03CX0_2),.clk(gclk));
	jdff dff_B_Z0CElkhq4_2(.din(w_dff_B_qS1V03CX0_2),.dout(w_dff_B_Z0CElkhq4_2),.clk(gclk));
	jdff dff_B_Z4oX2eZC2_2(.din(w_dff_B_Z0CElkhq4_2),.dout(w_dff_B_Z4oX2eZC2_2),.clk(gclk));
	jdff dff_B_mmnzgVYX2_2(.din(w_dff_B_Z4oX2eZC2_2),.dout(w_dff_B_mmnzgVYX2_2),.clk(gclk));
	jdff dff_B_nIFa6QTK4_2(.din(w_dff_B_mmnzgVYX2_2),.dout(w_dff_B_nIFa6QTK4_2),.clk(gclk));
	jdff dff_B_jmxhQi6B0_2(.din(w_dff_B_nIFa6QTK4_2),.dout(w_dff_B_jmxhQi6B0_2),.clk(gclk));
	jdff dff_B_TCn8qOCJ0_2(.din(w_dff_B_jmxhQi6B0_2),.dout(w_dff_B_TCn8qOCJ0_2),.clk(gclk));
	jdff dff_B_5LFSMMoA6_2(.din(w_dff_B_TCn8qOCJ0_2),.dout(w_dff_B_5LFSMMoA6_2),.clk(gclk));
	jdff dff_B_VltZJW6A5_2(.din(w_dff_B_5LFSMMoA6_2),.dout(w_dff_B_VltZJW6A5_2),.clk(gclk));
	jdff dff_B_N1Y9uENj0_2(.din(w_dff_B_VltZJW6A5_2),.dout(w_dff_B_N1Y9uENj0_2),.clk(gclk));
	jdff dff_B_sYSfSS3X1_2(.din(w_dff_B_N1Y9uENj0_2),.dout(w_dff_B_sYSfSS3X1_2),.clk(gclk));
	jdff dff_B_GgAsFdPT7_2(.din(w_dff_B_sYSfSS3X1_2),.dout(w_dff_B_GgAsFdPT7_2),.clk(gclk));
	jdff dff_B_wFhOb4C65_2(.din(w_dff_B_GgAsFdPT7_2),.dout(w_dff_B_wFhOb4C65_2),.clk(gclk));
	jdff dff_B_ESdU0vGh2_2(.din(w_dff_B_wFhOb4C65_2),.dout(w_dff_B_ESdU0vGh2_2),.clk(gclk));
	jdff dff_B_3V9cVasK4_2(.din(w_dff_B_ESdU0vGh2_2),.dout(w_dff_B_3V9cVasK4_2),.clk(gclk));
	jdff dff_B_0cHK6SdN2_2(.din(w_dff_B_3V9cVasK4_2),.dout(w_dff_B_0cHK6SdN2_2),.clk(gclk));
	jdff dff_B_5mXlmx2L3_2(.din(w_dff_B_0cHK6SdN2_2),.dout(w_dff_B_5mXlmx2L3_2),.clk(gclk));
	jdff dff_B_wGCg2bAy6_2(.din(w_dff_B_5mXlmx2L3_2),.dout(w_dff_B_wGCg2bAy6_2),.clk(gclk));
	jdff dff_B_RVQJ6Jm35_2(.din(w_dff_B_wGCg2bAy6_2),.dout(w_dff_B_RVQJ6Jm35_2),.clk(gclk));
	jdff dff_B_ja9cWSXL8_2(.din(w_dff_B_RVQJ6Jm35_2),.dout(w_dff_B_ja9cWSXL8_2),.clk(gclk));
	jdff dff_B_Se2B2VG83_2(.din(w_dff_B_ja9cWSXL8_2),.dout(w_dff_B_Se2B2VG83_2),.clk(gclk));
	jdff dff_B_IiGk1jLN6_2(.din(w_dff_B_Se2B2VG83_2),.dout(w_dff_B_IiGk1jLN6_2),.clk(gclk));
	jdff dff_B_4VFrOGka8_2(.din(w_dff_B_IiGk1jLN6_2),.dout(w_dff_B_4VFrOGka8_2),.clk(gclk));
	jdff dff_B_zSN1oP7s0_2(.din(w_dff_B_4VFrOGka8_2),.dout(w_dff_B_zSN1oP7s0_2),.clk(gclk));
	jdff dff_B_SzOasAmJ6_2(.din(w_dff_B_zSN1oP7s0_2),.dout(w_dff_B_SzOasAmJ6_2),.clk(gclk));
	jdff dff_B_Sn72WNp93_2(.din(w_dff_B_SzOasAmJ6_2),.dout(w_dff_B_Sn72WNp93_2),.clk(gclk));
	jdff dff_B_aUPtDaFI0_2(.din(w_dff_B_Sn72WNp93_2),.dout(w_dff_B_aUPtDaFI0_2),.clk(gclk));
	jdff dff_B_DJwCsm9G0_2(.din(w_dff_B_aUPtDaFI0_2),.dout(w_dff_B_DJwCsm9G0_2),.clk(gclk));
	jdff dff_B_iBTf6qWn7_2(.din(w_dff_B_DJwCsm9G0_2),.dout(w_dff_B_iBTf6qWn7_2),.clk(gclk));
	jdff dff_B_LSnm5eJl7_2(.din(w_dff_B_iBTf6qWn7_2),.dout(w_dff_B_LSnm5eJl7_2),.clk(gclk));
	jdff dff_B_pBlO0dTg7_2(.din(w_dff_B_LSnm5eJl7_2),.dout(w_dff_B_pBlO0dTg7_2),.clk(gclk));
	jdff dff_B_mtHqs9xD2_2(.din(w_dff_B_pBlO0dTg7_2),.dout(w_dff_B_mtHqs9xD2_2),.clk(gclk));
	jdff dff_B_bvKCUuvs3_2(.din(w_dff_B_mtHqs9xD2_2),.dout(w_dff_B_bvKCUuvs3_2),.clk(gclk));
	jdff dff_B_QGnr771I8_2(.din(w_dff_B_bvKCUuvs3_2),.dout(w_dff_B_QGnr771I8_2),.clk(gclk));
	jdff dff_B_OUTFygTT9_2(.din(w_dff_B_QGnr771I8_2),.dout(w_dff_B_OUTFygTT9_2),.clk(gclk));
	jdff dff_A_8FZFsssn1_0(.dout(w_n1034_0[0]),.din(w_dff_A_8FZFsssn1_0),.clk(gclk));
	jdff dff_B_YU9Fs9yY9_1(.din(n940),.dout(w_dff_B_YU9Fs9yY9_1),.clk(gclk));
	jdff dff_B_Cmju4XkZ6_2(.din(n835),.dout(w_dff_B_Cmju4XkZ6_2),.clk(gclk));
	jdff dff_B_XKJLECiX2_2(.din(w_dff_B_Cmju4XkZ6_2),.dout(w_dff_B_XKJLECiX2_2),.clk(gclk));
	jdff dff_B_9iJPZpOG0_2(.din(w_dff_B_XKJLECiX2_2),.dout(w_dff_B_9iJPZpOG0_2),.clk(gclk));
	jdff dff_B_riD7Hhbp0_2(.din(w_dff_B_9iJPZpOG0_2),.dout(w_dff_B_riD7Hhbp0_2),.clk(gclk));
	jdff dff_B_MUBFnhlV8_2(.din(w_dff_B_riD7Hhbp0_2),.dout(w_dff_B_MUBFnhlV8_2),.clk(gclk));
	jdff dff_B_oWvVhCi61_2(.din(w_dff_B_MUBFnhlV8_2),.dout(w_dff_B_oWvVhCi61_2),.clk(gclk));
	jdff dff_B_244JvJfI4_2(.din(w_dff_B_oWvVhCi61_2),.dout(w_dff_B_244JvJfI4_2),.clk(gclk));
	jdff dff_B_smPeRvbF6_2(.din(w_dff_B_244JvJfI4_2),.dout(w_dff_B_smPeRvbF6_2),.clk(gclk));
	jdff dff_B_144CYuEf9_2(.din(w_dff_B_smPeRvbF6_2),.dout(w_dff_B_144CYuEf9_2),.clk(gclk));
	jdff dff_B_VUKIUUqr1_2(.din(w_dff_B_144CYuEf9_2),.dout(w_dff_B_VUKIUUqr1_2),.clk(gclk));
	jdff dff_B_89P51siD4_2(.din(w_dff_B_VUKIUUqr1_2),.dout(w_dff_B_89P51siD4_2),.clk(gclk));
	jdff dff_B_53acqq0B2_2(.din(w_dff_B_89P51siD4_2),.dout(w_dff_B_53acqq0B2_2),.clk(gclk));
	jdff dff_B_QZyI493c2_2(.din(w_dff_B_53acqq0B2_2),.dout(w_dff_B_QZyI493c2_2),.clk(gclk));
	jdff dff_B_ieQuILvB7_2(.din(w_dff_B_QZyI493c2_2),.dout(w_dff_B_ieQuILvB7_2),.clk(gclk));
	jdff dff_B_9XVzMyIm3_2(.din(w_dff_B_ieQuILvB7_2),.dout(w_dff_B_9XVzMyIm3_2),.clk(gclk));
	jdff dff_B_CBSWQztz5_2(.din(w_dff_B_9XVzMyIm3_2),.dout(w_dff_B_CBSWQztz5_2),.clk(gclk));
	jdff dff_B_rLPlqZ4P8_2(.din(w_dff_B_CBSWQztz5_2),.dout(w_dff_B_rLPlqZ4P8_2),.clk(gclk));
	jdff dff_B_V0N7pwgU0_2(.din(w_dff_B_rLPlqZ4P8_2),.dout(w_dff_B_V0N7pwgU0_2),.clk(gclk));
	jdff dff_B_mJkgIjw38_2(.din(w_dff_B_V0N7pwgU0_2),.dout(w_dff_B_mJkgIjw38_2),.clk(gclk));
	jdff dff_B_7JTOvEP82_2(.din(w_dff_B_mJkgIjw38_2),.dout(w_dff_B_7JTOvEP82_2),.clk(gclk));
	jdff dff_B_PexFvD751_2(.din(w_dff_B_7JTOvEP82_2),.dout(w_dff_B_PexFvD751_2),.clk(gclk));
	jdff dff_B_cONiCm715_2(.din(w_dff_B_PexFvD751_2),.dout(w_dff_B_cONiCm715_2),.clk(gclk));
	jdff dff_B_1rjeMho76_2(.din(w_dff_B_cONiCm715_2),.dout(w_dff_B_1rjeMho76_2),.clk(gclk));
	jdff dff_B_53CgxPdn7_2(.din(w_dff_B_1rjeMho76_2),.dout(w_dff_B_53CgxPdn7_2),.clk(gclk));
	jdff dff_B_HFO9JKgM9_2(.din(w_dff_B_53CgxPdn7_2),.dout(w_dff_B_HFO9JKgM9_2),.clk(gclk));
	jdff dff_B_gNeO94Sq5_2(.din(w_dff_B_HFO9JKgM9_2),.dout(w_dff_B_gNeO94Sq5_2),.clk(gclk));
	jdff dff_B_8ZKoRUde3_2(.din(w_dff_B_gNeO94Sq5_2),.dout(w_dff_B_8ZKoRUde3_2),.clk(gclk));
	jdff dff_B_Kce3qLiA4_2(.din(w_dff_B_8ZKoRUde3_2),.dout(w_dff_B_Kce3qLiA4_2),.clk(gclk));
	jdff dff_B_N0iyvKSp3_2(.din(w_dff_B_Kce3qLiA4_2),.dout(w_dff_B_N0iyvKSp3_2),.clk(gclk));
	jdff dff_B_7hRlI4ES7_2(.din(w_dff_B_N0iyvKSp3_2),.dout(w_dff_B_7hRlI4ES7_2),.clk(gclk));
	jdff dff_B_KpSFj8zI0_2(.din(w_dff_B_7hRlI4ES7_2),.dout(w_dff_B_KpSFj8zI0_2),.clk(gclk));
	jdff dff_B_hFDt0Kgj7_2(.din(w_dff_B_KpSFj8zI0_2),.dout(w_dff_B_hFDt0Kgj7_2),.clk(gclk));
	jdff dff_B_uIG9bSch6_2(.din(w_dff_B_hFDt0Kgj7_2),.dout(w_dff_B_uIG9bSch6_2),.clk(gclk));
	jdff dff_B_MO1mBpfc0_2(.din(w_dff_B_uIG9bSch6_2),.dout(w_dff_B_MO1mBpfc0_2),.clk(gclk));
	jdff dff_B_PpjVTIOw8_2(.din(w_dff_B_MO1mBpfc0_2),.dout(w_dff_B_PpjVTIOw8_2),.clk(gclk));
	jdff dff_B_5MoCXwDb0_2(.din(w_dff_B_PpjVTIOw8_2),.dout(w_dff_B_5MoCXwDb0_2),.clk(gclk));
	jdff dff_B_wR1jJcqr2_2(.din(w_dff_B_5MoCXwDb0_2),.dout(w_dff_B_wR1jJcqr2_2),.clk(gclk));
	jdff dff_B_exRrguur1_2(.din(w_dff_B_wR1jJcqr2_2),.dout(w_dff_B_exRrguur1_2),.clk(gclk));
	jdff dff_B_wcFWD4uh4_2(.din(w_dff_B_exRrguur1_2),.dout(w_dff_B_wcFWD4uh4_2),.clk(gclk));
	jdff dff_B_RRR1lM4Q7_2(.din(w_dff_B_wcFWD4uh4_2),.dout(w_dff_B_RRR1lM4Q7_2),.clk(gclk));
	jdff dff_B_N6d7RHoj3_2(.din(w_dff_B_RRR1lM4Q7_2),.dout(w_dff_B_N6d7RHoj3_2),.clk(gclk));
	jdff dff_A_hHU6UceV1_1(.dout(w_n929_0[1]),.din(w_dff_A_hHU6UceV1_1),.clk(gclk));
	jdff dff_B_fzzOmr8J1_1(.din(n841),.dout(w_dff_B_fzzOmr8J1_1),.clk(gclk));
	jdff dff_B_yIf3oAeV5_1(.din(w_dff_B_fzzOmr8J1_1),.dout(w_dff_B_yIf3oAeV5_1),.clk(gclk));
	jdff dff_B_n1ODXD237_1(.din(w_dff_B_yIf3oAeV5_1),.dout(w_dff_B_n1ODXD237_1),.clk(gclk));
	jdff dff_B_wsJVEs0y7_1(.din(w_dff_B_n1ODXD237_1),.dout(w_dff_B_wsJVEs0y7_1),.clk(gclk));
	jdff dff_B_E0fa8WJR7_1(.din(w_dff_B_wsJVEs0y7_1),.dout(w_dff_B_E0fa8WJR7_1),.clk(gclk));
	jdff dff_B_4P9o2Dp96_1(.din(w_dff_B_E0fa8WJR7_1),.dout(w_dff_B_4P9o2Dp96_1),.clk(gclk));
	jdff dff_B_xnWLgX6V4_1(.din(w_dff_B_4P9o2Dp96_1),.dout(w_dff_B_xnWLgX6V4_1),.clk(gclk));
	jdff dff_B_UY0riLX37_1(.din(w_dff_B_xnWLgX6V4_1),.dout(w_dff_B_UY0riLX37_1),.clk(gclk));
	jdff dff_B_3BS2JmOQ3_1(.din(w_dff_B_UY0riLX37_1),.dout(w_dff_B_3BS2JmOQ3_1),.clk(gclk));
	jdff dff_B_GSLimxgR9_1(.din(w_dff_B_3BS2JmOQ3_1),.dout(w_dff_B_GSLimxgR9_1),.clk(gclk));
	jdff dff_B_xlxmilYB6_1(.din(w_dff_B_GSLimxgR9_1),.dout(w_dff_B_xlxmilYB6_1),.clk(gclk));
	jdff dff_B_g0smN5WD2_1(.din(w_dff_B_xlxmilYB6_1),.dout(w_dff_B_g0smN5WD2_1),.clk(gclk));
	jdff dff_B_pZCtFNNp6_1(.din(w_dff_B_g0smN5WD2_1),.dout(w_dff_B_pZCtFNNp6_1),.clk(gclk));
	jdff dff_B_YwwKu8VX9_1(.din(w_dff_B_pZCtFNNp6_1),.dout(w_dff_B_YwwKu8VX9_1),.clk(gclk));
	jdff dff_B_reuRlGSb4_1(.din(w_dff_B_YwwKu8VX9_1),.dout(w_dff_B_reuRlGSb4_1),.clk(gclk));
	jdff dff_B_LDMW8fnj0_1(.din(w_dff_B_reuRlGSb4_1),.dout(w_dff_B_LDMW8fnj0_1),.clk(gclk));
	jdff dff_B_ldAQpglH3_1(.din(w_dff_B_LDMW8fnj0_1),.dout(w_dff_B_ldAQpglH3_1),.clk(gclk));
	jdff dff_B_U8ofqQwm2_1(.din(w_dff_B_ldAQpglH3_1),.dout(w_dff_B_U8ofqQwm2_1),.clk(gclk));
	jdff dff_B_rsk4C2hf8_1(.din(w_dff_B_U8ofqQwm2_1),.dout(w_dff_B_rsk4C2hf8_1),.clk(gclk));
	jdff dff_B_0kIq5otZ5_1(.din(w_dff_B_rsk4C2hf8_1),.dout(w_dff_B_0kIq5otZ5_1),.clk(gclk));
	jdff dff_B_KghDC9zd6_1(.din(w_dff_B_0kIq5otZ5_1),.dout(w_dff_B_KghDC9zd6_1),.clk(gclk));
	jdff dff_B_mcbKVaae7_1(.din(w_dff_B_KghDC9zd6_1),.dout(w_dff_B_mcbKVaae7_1),.clk(gclk));
	jdff dff_B_3jhVv5In6_1(.din(w_dff_B_mcbKVaae7_1),.dout(w_dff_B_3jhVv5In6_1),.clk(gclk));
	jdff dff_B_b8eEDtjU1_1(.din(w_dff_B_3jhVv5In6_1),.dout(w_dff_B_b8eEDtjU1_1),.clk(gclk));
	jdff dff_B_iqDhQZyc2_1(.din(w_dff_B_b8eEDtjU1_1),.dout(w_dff_B_iqDhQZyc2_1),.clk(gclk));
	jdff dff_B_8xbn7ygX3_1(.din(w_dff_B_iqDhQZyc2_1),.dout(w_dff_B_8xbn7ygX3_1),.clk(gclk));
	jdff dff_B_SOSxbKXV8_1(.din(w_dff_B_8xbn7ygX3_1),.dout(w_dff_B_SOSxbKXV8_1),.clk(gclk));
	jdff dff_B_FGd2q3r20_1(.din(w_dff_B_SOSxbKXV8_1),.dout(w_dff_B_FGd2q3r20_1),.clk(gclk));
	jdff dff_B_MAUVOqBM6_1(.din(w_dff_B_FGd2q3r20_1),.dout(w_dff_B_MAUVOqBM6_1),.clk(gclk));
	jdff dff_B_hzdiH5tC3_1(.din(w_dff_B_MAUVOqBM6_1),.dout(w_dff_B_hzdiH5tC3_1),.clk(gclk));
	jdff dff_B_wQDkuLSQ2_1(.din(w_dff_B_hzdiH5tC3_1),.dout(w_dff_B_wQDkuLSQ2_1),.clk(gclk));
	jdff dff_B_gnZ80UEL4_1(.din(w_dff_B_wQDkuLSQ2_1),.dout(w_dff_B_gnZ80UEL4_1),.clk(gclk));
	jdff dff_B_6RSExyqG0_1(.din(w_dff_B_gnZ80UEL4_1),.dout(w_dff_B_6RSExyqG0_1),.clk(gclk));
	jdff dff_B_TEwbDJuc7_1(.din(w_dff_B_6RSExyqG0_1),.dout(w_dff_B_TEwbDJuc7_1),.clk(gclk));
	jdff dff_B_xxvzGOjw8_1(.din(w_dff_B_TEwbDJuc7_1),.dout(w_dff_B_xxvzGOjw8_1),.clk(gclk));
	jdff dff_B_k2Occ9hC0_1(.din(w_dff_B_xxvzGOjw8_1),.dout(w_dff_B_k2Occ9hC0_1),.clk(gclk));
	jdff dff_B_VV2MIwFT6_1(.din(w_dff_B_k2Occ9hC0_1),.dout(w_dff_B_VV2MIwFT6_1),.clk(gclk));
	jdff dff_B_KpqY4Roc0_1(.din(n836),.dout(w_dff_B_KpqY4Roc0_1),.clk(gclk));
	jdff dff_A_0x7sXd5j0_0(.dout(w_n735_0[0]),.din(w_dff_A_0x7sXd5j0_0),.clk(gclk));
	jdff dff_A_1t0KfLDD4_0(.dout(w_dff_A_0x7sXd5j0_0),.din(w_dff_A_1t0KfLDD4_0),.clk(gclk));
	jdff dff_A_c1C5p1y66_0(.dout(w_dff_A_1t0KfLDD4_0),.din(w_dff_A_c1C5p1y66_0),.clk(gclk));
	jdff dff_A_OEpCSvpc2_0(.dout(w_dff_A_c1C5p1y66_0),.din(w_dff_A_OEpCSvpc2_0),.clk(gclk));
	jdff dff_A_HboQAD2X9_0(.dout(w_dff_A_OEpCSvpc2_0),.din(w_dff_A_HboQAD2X9_0),.clk(gclk));
	jdff dff_A_VSaBkZhR9_0(.dout(w_dff_A_HboQAD2X9_0),.din(w_dff_A_VSaBkZhR9_0),.clk(gclk));
	jdff dff_A_tx41zBWz7_0(.dout(w_dff_A_VSaBkZhR9_0),.din(w_dff_A_tx41zBWz7_0),.clk(gclk));
	jdff dff_A_ar4OMavj3_0(.dout(w_dff_A_tx41zBWz7_0),.din(w_dff_A_ar4OMavj3_0),.clk(gclk));
	jdff dff_A_3kyOvU4F9_0(.dout(w_dff_A_ar4OMavj3_0),.din(w_dff_A_3kyOvU4F9_0),.clk(gclk));
	jdff dff_A_QqCw3m452_0(.dout(w_dff_A_3kyOvU4F9_0),.din(w_dff_A_QqCw3m452_0),.clk(gclk));
	jdff dff_A_2TVhhPhf6_0(.dout(w_dff_A_QqCw3m452_0),.din(w_dff_A_2TVhhPhf6_0),.clk(gclk));
	jdff dff_A_eQ9CyBdA7_0(.dout(w_dff_A_2TVhhPhf6_0),.din(w_dff_A_eQ9CyBdA7_0),.clk(gclk));
	jdff dff_A_Q6Bpm4h13_0(.dout(w_dff_A_eQ9CyBdA7_0),.din(w_dff_A_Q6Bpm4h13_0),.clk(gclk));
	jdff dff_A_zz8k9yHb4_0(.dout(w_dff_A_Q6Bpm4h13_0),.din(w_dff_A_zz8k9yHb4_0),.clk(gclk));
	jdff dff_A_itMEMbUa8_0(.dout(w_dff_A_zz8k9yHb4_0),.din(w_dff_A_itMEMbUa8_0),.clk(gclk));
	jdff dff_A_gP9gCfzn7_0(.dout(w_dff_A_itMEMbUa8_0),.din(w_dff_A_gP9gCfzn7_0),.clk(gclk));
	jdff dff_A_EPexjiHt3_0(.dout(w_dff_A_gP9gCfzn7_0),.din(w_dff_A_EPexjiHt3_0),.clk(gclk));
	jdff dff_A_gpcO4scG3_0(.dout(w_dff_A_EPexjiHt3_0),.din(w_dff_A_gpcO4scG3_0),.clk(gclk));
	jdff dff_A_hISEMg0b2_0(.dout(w_dff_A_gpcO4scG3_0),.din(w_dff_A_hISEMg0b2_0),.clk(gclk));
	jdff dff_A_AErJsgPT6_0(.dout(w_dff_A_hISEMg0b2_0),.din(w_dff_A_AErJsgPT6_0),.clk(gclk));
	jdff dff_A_XnsgTuen7_0(.dout(w_dff_A_AErJsgPT6_0),.din(w_dff_A_XnsgTuen7_0),.clk(gclk));
	jdff dff_A_gSUsSpUM9_0(.dout(w_dff_A_XnsgTuen7_0),.din(w_dff_A_gSUsSpUM9_0),.clk(gclk));
	jdff dff_A_xJh2KpoY8_0(.dout(w_dff_A_gSUsSpUM9_0),.din(w_dff_A_xJh2KpoY8_0),.clk(gclk));
	jdff dff_A_aqHw9f9o2_0(.dout(w_dff_A_xJh2KpoY8_0),.din(w_dff_A_aqHw9f9o2_0),.clk(gclk));
	jdff dff_A_Z1OQV4rR3_0(.dout(w_dff_A_aqHw9f9o2_0),.din(w_dff_A_Z1OQV4rR3_0),.clk(gclk));
	jdff dff_A_aW88qQaB0_0(.dout(w_dff_A_Z1OQV4rR3_0),.din(w_dff_A_aW88qQaB0_0),.clk(gclk));
	jdff dff_A_dBKO5jgt7_0(.dout(w_dff_A_aW88qQaB0_0),.din(w_dff_A_dBKO5jgt7_0),.clk(gclk));
	jdff dff_A_tvTL01T53_0(.dout(w_dff_A_dBKO5jgt7_0),.din(w_dff_A_tvTL01T53_0),.clk(gclk));
	jdff dff_A_0NIWXbRw4_0(.dout(w_dff_A_tvTL01T53_0),.din(w_dff_A_0NIWXbRw4_0),.clk(gclk));
	jdff dff_A_RF6jJ1qM4_0(.dout(w_dff_A_0NIWXbRw4_0),.din(w_dff_A_RF6jJ1qM4_0),.clk(gclk));
	jdff dff_A_wpKf0Pax1_0(.dout(w_dff_A_RF6jJ1qM4_0),.din(w_dff_A_wpKf0Pax1_0),.clk(gclk));
	jdff dff_A_cSGwaseN9_0(.dout(w_dff_A_wpKf0Pax1_0),.din(w_dff_A_cSGwaseN9_0),.clk(gclk));
	jdff dff_A_IqWGRieV0_0(.dout(w_dff_A_cSGwaseN9_0),.din(w_dff_A_IqWGRieV0_0),.clk(gclk));
	jdff dff_A_MquVKvAs7_0(.dout(w_dff_A_IqWGRieV0_0),.din(w_dff_A_MquVKvAs7_0),.clk(gclk));
	jdff dff_A_iK6EvYbl7_0(.dout(w_dff_A_MquVKvAs7_0),.din(w_dff_A_iK6EvYbl7_0),.clk(gclk));
	jdff dff_A_ojtGVxro0_0(.dout(w_dff_A_iK6EvYbl7_0),.din(w_dff_A_ojtGVxro0_0),.clk(gclk));
	jdff dff_A_VdfbowkM1_0(.dout(w_dff_A_ojtGVxro0_0),.din(w_dff_A_VdfbowkM1_0),.clk(gclk));
	jdff dff_A_7YxzHdl95_0(.dout(w_dff_A_VdfbowkM1_0),.din(w_dff_A_7YxzHdl95_0),.clk(gclk));
	jdff dff_A_CZ2jEFdf6_0(.dout(w_n823_0[0]),.din(w_dff_A_CZ2jEFdf6_0),.clk(gclk));
	jdff dff_B_n1qofQ7N6_1(.din(n737),.dout(w_dff_B_n1qofQ7N6_1),.clk(gclk));
	jdff dff_A_To4CQYwR5_0(.dout(w_n642_0[0]),.din(w_dff_A_To4CQYwR5_0),.clk(gclk));
	jdff dff_A_ggh7op5Z7_0(.dout(w_dff_A_To4CQYwR5_0),.din(w_dff_A_ggh7op5Z7_0),.clk(gclk));
	jdff dff_A_yxOIQ4lR2_0(.dout(w_dff_A_ggh7op5Z7_0),.din(w_dff_A_yxOIQ4lR2_0),.clk(gclk));
	jdff dff_A_FrkpCw5a8_0(.dout(w_dff_A_yxOIQ4lR2_0),.din(w_dff_A_FrkpCw5a8_0),.clk(gclk));
	jdff dff_A_JElZmtGa1_0(.dout(w_dff_A_FrkpCw5a8_0),.din(w_dff_A_JElZmtGa1_0),.clk(gclk));
	jdff dff_A_3mFIzyLZ1_0(.dout(w_dff_A_JElZmtGa1_0),.din(w_dff_A_3mFIzyLZ1_0),.clk(gclk));
	jdff dff_A_3HmzR6yy1_0(.dout(w_dff_A_3mFIzyLZ1_0),.din(w_dff_A_3HmzR6yy1_0),.clk(gclk));
	jdff dff_A_RlOVBzJF3_0(.dout(w_dff_A_3HmzR6yy1_0),.din(w_dff_A_RlOVBzJF3_0),.clk(gclk));
	jdff dff_A_eCWTqBit2_0(.dout(w_dff_A_RlOVBzJF3_0),.din(w_dff_A_eCWTqBit2_0),.clk(gclk));
	jdff dff_A_smlIJURR8_0(.dout(w_dff_A_eCWTqBit2_0),.din(w_dff_A_smlIJURR8_0),.clk(gclk));
	jdff dff_A_Aeraraba3_0(.dout(w_dff_A_smlIJURR8_0),.din(w_dff_A_Aeraraba3_0),.clk(gclk));
	jdff dff_A_WbXmNPCy1_0(.dout(w_dff_A_Aeraraba3_0),.din(w_dff_A_WbXmNPCy1_0),.clk(gclk));
	jdff dff_A_fzBGNR4C0_0(.dout(w_dff_A_WbXmNPCy1_0),.din(w_dff_A_fzBGNR4C0_0),.clk(gclk));
	jdff dff_A_pDscmNUD6_0(.dout(w_dff_A_fzBGNR4C0_0),.din(w_dff_A_pDscmNUD6_0),.clk(gclk));
	jdff dff_A_1rabCNHB7_0(.dout(w_dff_A_pDscmNUD6_0),.din(w_dff_A_1rabCNHB7_0),.clk(gclk));
	jdff dff_A_tEb8e0M24_0(.dout(w_dff_A_1rabCNHB7_0),.din(w_dff_A_tEb8e0M24_0),.clk(gclk));
	jdff dff_A_EWJSBKE89_0(.dout(w_dff_A_tEb8e0M24_0),.din(w_dff_A_EWJSBKE89_0),.clk(gclk));
	jdff dff_A_GMdCjHzv1_0(.dout(w_dff_A_EWJSBKE89_0),.din(w_dff_A_GMdCjHzv1_0),.clk(gclk));
	jdff dff_A_8DzFQCZx0_0(.dout(w_dff_A_GMdCjHzv1_0),.din(w_dff_A_8DzFQCZx0_0),.clk(gclk));
	jdff dff_A_5gg0W96i4_0(.dout(w_dff_A_8DzFQCZx0_0),.din(w_dff_A_5gg0W96i4_0),.clk(gclk));
	jdff dff_A_mF2BH9hX5_0(.dout(w_dff_A_5gg0W96i4_0),.din(w_dff_A_mF2BH9hX5_0),.clk(gclk));
	jdff dff_A_6qLITpxo1_0(.dout(w_dff_A_mF2BH9hX5_0),.din(w_dff_A_6qLITpxo1_0),.clk(gclk));
	jdff dff_A_gvQuIHqD6_0(.dout(w_dff_A_6qLITpxo1_0),.din(w_dff_A_gvQuIHqD6_0),.clk(gclk));
	jdff dff_A_np2AACK71_0(.dout(w_dff_A_gvQuIHqD6_0),.din(w_dff_A_np2AACK71_0),.clk(gclk));
	jdff dff_A_dSSqv5el9_0(.dout(w_dff_A_np2AACK71_0),.din(w_dff_A_dSSqv5el9_0),.clk(gclk));
	jdff dff_A_6ZcnzBpi8_0(.dout(w_dff_A_dSSqv5el9_0),.din(w_dff_A_6ZcnzBpi8_0),.clk(gclk));
	jdff dff_A_9TJo8J1h8_0(.dout(w_dff_A_6ZcnzBpi8_0),.din(w_dff_A_9TJo8J1h8_0),.clk(gclk));
	jdff dff_A_A3svwYQ96_0(.dout(w_dff_A_9TJo8J1h8_0),.din(w_dff_A_A3svwYQ96_0),.clk(gclk));
	jdff dff_A_wgUbjRhB2_0(.dout(w_dff_A_A3svwYQ96_0),.din(w_dff_A_wgUbjRhB2_0),.clk(gclk));
	jdff dff_A_7HSPdK1j0_0(.dout(w_dff_A_wgUbjRhB2_0),.din(w_dff_A_7HSPdK1j0_0),.clk(gclk));
	jdff dff_A_htXIfznG4_0(.dout(w_dff_A_7HSPdK1j0_0),.din(w_dff_A_htXIfznG4_0),.clk(gclk));
	jdff dff_A_WKGGiWb44_0(.dout(w_dff_A_htXIfznG4_0),.din(w_dff_A_WKGGiWb44_0),.clk(gclk));
	jdff dff_A_XareqLXt0_0(.dout(w_dff_A_WKGGiWb44_0),.din(w_dff_A_XareqLXt0_0),.clk(gclk));
	jdff dff_A_gM7V1X5D8_0(.dout(w_dff_A_XareqLXt0_0),.din(w_dff_A_gM7V1X5D8_0),.clk(gclk));
	jdff dff_A_1KDVfjr33_0(.dout(w_dff_A_gM7V1X5D8_0),.din(w_dff_A_1KDVfjr33_0),.clk(gclk));
	jdff dff_A_OgeeSzwv6_0(.dout(w_n723_0[0]),.din(w_dff_A_OgeeSzwv6_0),.clk(gclk));
	jdff dff_B_T0JlXUcf3_1(.din(n644),.dout(w_dff_B_T0JlXUcf3_1),.clk(gclk));
	jdff dff_A_1FBtlnJd4_0(.dout(w_n556_0[0]),.din(w_dff_A_1FBtlnJd4_0),.clk(gclk));
	jdff dff_A_YRhvihQA6_0(.dout(w_dff_A_1FBtlnJd4_0),.din(w_dff_A_YRhvihQA6_0),.clk(gclk));
	jdff dff_A_2u9NoB241_0(.dout(w_dff_A_YRhvihQA6_0),.din(w_dff_A_2u9NoB241_0),.clk(gclk));
	jdff dff_A_qw0GAhjs9_0(.dout(w_dff_A_2u9NoB241_0),.din(w_dff_A_qw0GAhjs9_0),.clk(gclk));
	jdff dff_A_QDn77CaY5_0(.dout(w_dff_A_qw0GAhjs9_0),.din(w_dff_A_QDn77CaY5_0),.clk(gclk));
	jdff dff_A_voPjoagP0_0(.dout(w_dff_A_QDn77CaY5_0),.din(w_dff_A_voPjoagP0_0),.clk(gclk));
	jdff dff_A_FJAaoLIb1_0(.dout(w_dff_A_voPjoagP0_0),.din(w_dff_A_FJAaoLIb1_0),.clk(gclk));
	jdff dff_A_GLoNUQPe4_0(.dout(w_dff_A_FJAaoLIb1_0),.din(w_dff_A_GLoNUQPe4_0),.clk(gclk));
	jdff dff_A_hvLyiykL5_0(.dout(w_dff_A_GLoNUQPe4_0),.din(w_dff_A_hvLyiykL5_0),.clk(gclk));
	jdff dff_A_6E27U3Vr7_0(.dout(w_dff_A_hvLyiykL5_0),.din(w_dff_A_6E27U3Vr7_0),.clk(gclk));
	jdff dff_A_kZyClB2W3_0(.dout(w_dff_A_6E27U3Vr7_0),.din(w_dff_A_kZyClB2W3_0),.clk(gclk));
	jdff dff_A_szql5YIY2_0(.dout(w_dff_A_kZyClB2W3_0),.din(w_dff_A_szql5YIY2_0),.clk(gclk));
	jdff dff_A_dhUrHtm81_0(.dout(w_dff_A_szql5YIY2_0),.din(w_dff_A_dhUrHtm81_0),.clk(gclk));
	jdff dff_A_uVzSUWcq3_0(.dout(w_dff_A_dhUrHtm81_0),.din(w_dff_A_uVzSUWcq3_0),.clk(gclk));
	jdff dff_A_6OhY4Zcq0_0(.dout(w_dff_A_uVzSUWcq3_0),.din(w_dff_A_6OhY4Zcq0_0),.clk(gclk));
	jdff dff_A_jlwv0Zhf6_0(.dout(w_dff_A_6OhY4Zcq0_0),.din(w_dff_A_jlwv0Zhf6_0),.clk(gclk));
	jdff dff_A_9AwAA0PN1_0(.dout(w_dff_A_jlwv0Zhf6_0),.din(w_dff_A_9AwAA0PN1_0),.clk(gclk));
	jdff dff_A_jMPHnMES8_0(.dout(w_dff_A_9AwAA0PN1_0),.din(w_dff_A_jMPHnMES8_0),.clk(gclk));
	jdff dff_A_STtMjR668_0(.dout(w_dff_A_jMPHnMES8_0),.din(w_dff_A_STtMjR668_0),.clk(gclk));
	jdff dff_A_i4fnA0FW5_0(.dout(w_dff_A_STtMjR668_0),.din(w_dff_A_i4fnA0FW5_0),.clk(gclk));
	jdff dff_A_9ca1J4kT0_0(.dout(w_dff_A_i4fnA0FW5_0),.din(w_dff_A_9ca1J4kT0_0),.clk(gclk));
	jdff dff_A_4KZVR7Fb3_0(.dout(w_dff_A_9ca1J4kT0_0),.din(w_dff_A_4KZVR7Fb3_0),.clk(gclk));
	jdff dff_A_OY8XUwl90_0(.dout(w_dff_A_4KZVR7Fb3_0),.din(w_dff_A_OY8XUwl90_0),.clk(gclk));
	jdff dff_A_qWRvH4Bx0_0(.dout(w_dff_A_OY8XUwl90_0),.din(w_dff_A_qWRvH4Bx0_0),.clk(gclk));
	jdff dff_A_Vp8wa24D0_0(.dout(w_dff_A_qWRvH4Bx0_0),.din(w_dff_A_Vp8wa24D0_0),.clk(gclk));
	jdff dff_A_wVfnTa6n8_0(.dout(w_dff_A_Vp8wa24D0_0),.din(w_dff_A_wVfnTa6n8_0),.clk(gclk));
	jdff dff_A_ZVuLWI3g9_0(.dout(w_dff_A_wVfnTa6n8_0),.din(w_dff_A_ZVuLWI3g9_0),.clk(gclk));
	jdff dff_A_ctXthAzv4_0(.dout(w_dff_A_ZVuLWI3g9_0),.din(w_dff_A_ctXthAzv4_0),.clk(gclk));
	jdff dff_A_iQzNwUYQ3_0(.dout(w_dff_A_ctXthAzv4_0),.din(w_dff_A_iQzNwUYQ3_0),.clk(gclk));
	jdff dff_A_pB3OO0pO7_0(.dout(w_dff_A_iQzNwUYQ3_0),.din(w_dff_A_pB3OO0pO7_0),.clk(gclk));
	jdff dff_A_w2rvrd2E6_0(.dout(w_dff_A_pB3OO0pO7_0),.din(w_dff_A_w2rvrd2E6_0),.clk(gclk));
	jdff dff_A_4Sqb3nNa1_0(.dout(w_dff_A_w2rvrd2E6_0),.din(w_dff_A_4Sqb3nNa1_0),.clk(gclk));
	jdff dff_A_5WYeOW9D8_0(.dout(w_n630_0[0]),.din(w_dff_A_5WYeOW9D8_0),.clk(gclk));
	jdff dff_B_SpoUZEwd0_1(.din(n558),.dout(w_dff_B_SpoUZEwd0_1),.clk(gclk));
	jdff dff_A_BonLGtCS7_0(.dout(w_n477_0[0]),.din(w_dff_A_BonLGtCS7_0),.clk(gclk));
	jdff dff_A_qXCCAQEi7_0(.dout(w_dff_A_BonLGtCS7_0),.din(w_dff_A_qXCCAQEi7_0),.clk(gclk));
	jdff dff_A_hvhrF0bn2_0(.dout(w_dff_A_qXCCAQEi7_0),.din(w_dff_A_hvhrF0bn2_0),.clk(gclk));
	jdff dff_A_hZ6uZVYi5_0(.dout(w_dff_A_hvhrF0bn2_0),.din(w_dff_A_hZ6uZVYi5_0),.clk(gclk));
	jdff dff_A_FpERn6Cd7_0(.dout(w_dff_A_hZ6uZVYi5_0),.din(w_dff_A_FpERn6Cd7_0),.clk(gclk));
	jdff dff_A_KEBm57gp9_0(.dout(w_dff_A_FpERn6Cd7_0),.din(w_dff_A_KEBm57gp9_0),.clk(gclk));
	jdff dff_A_Ff4uTXqb2_0(.dout(w_dff_A_KEBm57gp9_0),.din(w_dff_A_Ff4uTXqb2_0),.clk(gclk));
	jdff dff_A_4KQt9KZB9_0(.dout(w_dff_A_Ff4uTXqb2_0),.din(w_dff_A_4KQt9KZB9_0),.clk(gclk));
	jdff dff_A_aSzd3V5y7_0(.dout(w_dff_A_4KQt9KZB9_0),.din(w_dff_A_aSzd3V5y7_0),.clk(gclk));
	jdff dff_A_eQBooRoZ2_0(.dout(w_dff_A_aSzd3V5y7_0),.din(w_dff_A_eQBooRoZ2_0),.clk(gclk));
	jdff dff_A_9EjCucF43_0(.dout(w_dff_A_eQBooRoZ2_0),.din(w_dff_A_9EjCucF43_0),.clk(gclk));
	jdff dff_A_rnB0gZ014_0(.dout(w_dff_A_9EjCucF43_0),.din(w_dff_A_rnB0gZ014_0),.clk(gclk));
	jdff dff_A_D8avDmqJ8_0(.dout(w_dff_A_rnB0gZ014_0),.din(w_dff_A_D8avDmqJ8_0),.clk(gclk));
	jdff dff_A_zjAVnxuZ6_0(.dout(w_dff_A_D8avDmqJ8_0),.din(w_dff_A_zjAVnxuZ6_0),.clk(gclk));
	jdff dff_A_QgM4FMme2_0(.dout(w_dff_A_zjAVnxuZ6_0),.din(w_dff_A_QgM4FMme2_0),.clk(gclk));
	jdff dff_A_6jVIJBg65_0(.dout(w_dff_A_QgM4FMme2_0),.din(w_dff_A_6jVIJBg65_0),.clk(gclk));
	jdff dff_A_iSLGsF3h3_0(.dout(w_dff_A_6jVIJBg65_0),.din(w_dff_A_iSLGsF3h3_0),.clk(gclk));
	jdff dff_A_FHou2Rh10_0(.dout(w_dff_A_iSLGsF3h3_0),.din(w_dff_A_FHou2Rh10_0),.clk(gclk));
	jdff dff_A_GQCklcge3_0(.dout(w_dff_A_FHou2Rh10_0),.din(w_dff_A_GQCklcge3_0),.clk(gclk));
	jdff dff_A_oSYctBLT9_0(.dout(w_dff_A_GQCklcge3_0),.din(w_dff_A_oSYctBLT9_0),.clk(gclk));
	jdff dff_A_jFsyfJ843_0(.dout(w_dff_A_oSYctBLT9_0),.din(w_dff_A_jFsyfJ843_0),.clk(gclk));
	jdff dff_A_eAmjjxs99_0(.dout(w_dff_A_jFsyfJ843_0),.din(w_dff_A_eAmjjxs99_0),.clk(gclk));
	jdff dff_A_Oa5q03m06_0(.dout(w_dff_A_eAmjjxs99_0),.din(w_dff_A_Oa5q03m06_0),.clk(gclk));
	jdff dff_A_slspMlqY1_0(.dout(w_dff_A_Oa5q03m06_0),.din(w_dff_A_slspMlqY1_0),.clk(gclk));
	jdff dff_A_cSBYrpul6_0(.dout(w_dff_A_slspMlqY1_0),.din(w_dff_A_cSBYrpul6_0),.clk(gclk));
	jdff dff_A_lzmXifd79_0(.dout(w_dff_A_cSBYrpul6_0),.din(w_dff_A_lzmXifd79_0),.clk(gclk));
	jdff dff_A_InnUBaSo2_0(.dout(w_dff_A_lzmXifd79_0),.din(w_dff_A_InnUBaSo2_0),.clk(gclk));
	jdff dff_A_E2J9lZA42_0(.dout(w_dff_A_InnUBaSo2_0),.din(w_dff_A_E2J9lZA42_0),.clk(gclk));
	jdff dff_A_UZ7DrGWN9_0(.dout(w_dff_A_E2J9lZA42_0),.din(w_dff_A_UZ7DrGWN9_0),.clk(gclk));
	jdff dff_A_8tiOknIL2_0(.dout(w_n544_0[0]),.din(w_dff_A_8tiOknIL2_0),.clk(gclk));
	jdff dff_B_wkFc1ith2_1(.din(n479),.dout(w_dff_B_wkFc1ith2_1),.clk(gclk));
	jdff dff_A_Z0qkaj588_0(.dout(w_n405_0[0]),.din(w_dff_A_Z0qkaj588_0),.clk(gclk));
	jdff dff_A_Mgna3mO74_0(.dout(w_dff_A_Z0qkaj588_0),.din(w_dff_A_Mgna3mO74_0),.clk(gclk));
	jdff dff_A_0K0H1mcN6_0(.dout(w_dff_A_Mgna3mO74_0),.din(w_dff_A_0K0H1mcN6_0),.clk(gclk));
	jdff dff_A_U8uKCunH7_0(.dout(w_dff_A_0K0H1mcN6_0),.din(w_dff_A_U8uKCunH7_0),.clk(gclk));
	jdff dff_A_ZCcxNhSW5_0(.dout(w_dff_A_U8uKCunH7_0),.din(w_dff_A_ZCcxNhSW5_0),.clk(gclk));
	jdff dff_A_Vq4Igk4k9_0(.dout(w_dff_A_ZCcxNhSW5_0),.din(w_dff_A_Vq4Igk4k9_0),.clk(gclk));
	jdff dff_A_leSBSrue9_0(.dout(w_dff_A_Vq4Igk4k9_0),.din(w_dff_A_leSBSrue9_0),.clk(gclk));
	jdff dff_A_a1D3WmsL1_0(.dout(w_dff_A_leSBSrue9_0),.din(w_dff_A_a1D3WmsL1_0),.clk(gclk));
	jdff dff_A_97FYEoeL1_0(.dout(w_dff_A_a1D3WmsL1_0),.din(w_dff_A_97FYEoeL1_0),.clk(gclk));
	jdff dff_A_NeaUB9Zu6_0(.dout(w_dff_A_97FYEoeL1_0),.din(w_dff_A_NeaUB9Zu6_0),.clk(gclk));
	jdff dff_A_wLEdSDoS0_0(.dout(w_dff_A_NeaUB9Zu6_0),.din(w_dff_A_wLEdSDoS0_0),.clk(gclk));
	jdff dff_A_AZ733hQx0_0(.dout(w_dff_A_wLEdSDoS0_0),.din(w_dff_A_AZ733hQx0_0),.clk(gclk));
	jdff dff_A_owYA2bLA9_0(.dout(w_dff_A_AZ733hQx0_0),.din(w_dff_A_owYA2bLA9_0),.clk(gclk));
	jdff dff_A_h1BVIcgu9_0(.dout(w_dff_A_owYA2bLA9_0),.din(w_dff_A_h1BVIcgu9_0),.clk(gclk));
	jdff dff_A_OKGD1lo05_0(.dout(w_dff_A_h1BVIcgu9_0),.din(w_dff_A_OKGD1lo05_0),.clk(gclk));
	jdff dff_A_L2wyClKZ6_0(.dout(w_dff_A_OKGD1lo05_0),.din(w_dff_A_L2wyClKZ6_0),.clk(gclk));
	jdff dff_A_1pTA4NV72_0(.dout(w_dff_A_L2wyClKZ6_0),.din(w_dff_A_1pTA4NV72_0),.clk(gclk));
	jdff dff_A_sulAL0da8_0(.dout(w_dff_A_1pTA4NV72_0),.din(w_dff_A_sulAL0da8_0),.clk(gclk));
	jdff dff_A_jKqVXPEE7_0(.dout(w_dff_A_sulAL0da8_0),.din(w_dff_A_jKqVXPEE7_0),.clk(gclk));
	jdff dff_A_5ZzBjgKr7_0(.dout(w_dff_A_jKqVXPEE7_0),.din(w_dff_A_5ZzBjgKr7_0),.clk(gclk));
	jdff dff_A_fh5MXxQN3_0(.dout(w_dff_A_5ZzBjgKr7_0),.din(w_dff_A_fh5MXxQN3_0),.clk(gclk));
	jdff dff_A_kCwfeBfB8_0(.dout(w_dff_A_fh5MXxQN3_0),.din(w_dff_A_kCwfeBfB8_0),.clk(gclk));
	jdff dff_A_Se7yCc9P7_0(.dout(w_dff_A_kCwfeBfB8_0),.din(w_dff_A_Se7yCc9P7_0),.clk(gclk));
	jdff dff_A_alDo3FBj1_0(.dout(w_dff_A_Se7yCc9P7_0),.din(w_dff_A_alDo3FBj1_0),.clk(gclk));
	jdff dff_A_jw9LVS7v8_0(.dout(w_dff_A_alDo3FBj1_0),.din(w_dff_A_jw9LVS7v8_0),.clk(gclk));
	jdff dff_A_pPk0ZHij9_0(.dout(w_dff_A_jw9LVS7v8_0),.din(w_dff_A_pPk0ZHij9_0),.clk(gclk));
	jdff dff_A_w7T9nth90_0(.dout(w_n465_0[0]),.din(w_dff_A_w7T9nth90_0),.clk(gclk));
	jdff dff_B_cNZdpEw14_1(.din(n407),.dout(w_dff_B_cNZdpEw14_1),.clk(gclk));
	jdff dff_A_dDbcnEjY4_0(.dout(w_n341_0[0]),.din(w_dff_A_dDbcnEjY4_0),.clk(gclk));
	jdff dff_A_JIpFM2TJ9_0(.dout(w_dff_A_dDbcnEjY4_0),.din(w_dff_A_JIpFM2TJ9_0),.clk(gclk));
	jdff dff_A_UivY7Xvx2_0(.dout(w_dff_A_JIpFM2TJ9_0),.din(w_dff_A_UivY7Xvx2_0),.clk(gclk));
	jdff dff_A_66jSKIFW0_0(.dout(w_dff_A_UivY7Xvx2_0),.din(w_dff_A_66jSKIFW0_0),.clk(gclk));
	jdff dff_A_c7SNGAbI1_0(.dout(w_dff_A_66jSKIFW0_0),.din(w_dff_A_c7SNGAbI1_0),.clk(gclk));
	jdff dff_A_Qn1WG3OA6_0(.dout(w_dff_A_c7SNGAbI1_0),.din(w_dff_A_Qn1WG3OA6_0),.clk(gclk));
	jdff dff_A_UX79hV7d6_0(.dout(w_dff_A_Qn1WG3OA6_0),.din(w_dff_A_UX79hV7d6_0),.clk(gclk));
	jdff dff_A_3QMeQRYx4_0(.dout(w_dff_A_UX79hV7d6_0),.din(w_dff_A_3QMeQRYx4_0),.clk(gclk));
	jdff dff_A_AkiNZV2m3_0(.dout(w_dff_A_3QMeQRYx4_0),.din(w_dff_A_AkiNZV2m3_0),.clk(gclk));
	jdff dff_A_4GLBo9I30_0(.dout(w_dff_A_AkiNZV2m3_0),.din(w_dff_A_4GLBo9I30_0),.clk(gclk));
	jdff dff_A_C6znERXG9_0(.dout(w_dff_A_4GLBo9I30_0),.din(w_dff_A_C6znERXG9_0),.clk(gclk));
	jdff dff_A_OTrDjAso9_0(.dout(w_dff_A_C6znERXG9_0),.din(w_dff_A_OTrDjAso9_0),.clk(gclk));
	jdff dff_A_M9TN7u1o8_0(.dout(w_dff_A_OTrDjAso9_0),.din(w_dff_A_M9TN7u1o8_0),.clk(gclk));
	jdff dff_A_SpNUAerN7_0(.dout(w_dff_A_M9TN7u1o8_0),.din(w_dff_A_SpNUAerN7_0),.clk(gclk));
	jdff dff_A_Li1BxMt35_0(.dout(w_dff_A_SpNUAerN7_0),.din(w_dff_A_Li1BxMt35_0),.clk(gclk));
	jdff dff_A_hVARLdF90_0(.dout(w_dff_A_Li1BxMt35_0),.din(w_dff_A_hVARLdF90_0),.clk(gclk));
	jdff dff_A_KOyFnJ6P3_0(.dout(w_dff_A_hVARLdF90_0),.din(w_dff_A_KOyFnJ6P3_0),.clk(gclk));
	jdff dff_A_heyaKFTt6_0(.dout(w_dff_A_KOyFnJ6P3_0),.din(w_dff_A_heyaKFTt6_0),.clk(gclk));
	jdff dff_A_IfoL8a475_0(.dout(w_dff_A_heyaKFTt6_0),.din(w_dff_A_IfoL8a475_0),.clk(gclk));
	jdff dff_A_qzKxelDI9_0(.dout(w_dff_A_IfoL8a475_0),.din(w_dff_A_qzKxelDI9_0),.clk(gclk));
	jdff dff_A_wrjPjiGi8_0(.dout(w_dff_A_qzKxelDI9_0),.din(w_dff_A_wrjPjiGi8_0),.clk(gclk));
	jdff dff_A_U06rrlK61_0(.dout(w_dff_A_wrjPjiGi8_0),.din(w_dff_A_U06rrlK61_0),.clk(gclk));
	jdff dff_A_F7GGot049_0(.dout(w_dff_A_U06rrlK61_0),.din(w_dff_A_F7GGot049_0),.clk(gclk));
	jdff dff_A_H5a6kMnc7_0(.dout(w_n393_0[0]),.din(w_dff_A_H5a6kMnc7_0),.clk(gclk));
	jdff dff_B_YN9xniCe7_1(.din(n343),.dout(w_dff_B_YN9xniCe7_1),.clk(gclk));
	jdff dff_A_B3WQpwTl4_0(.dout(w_n283_0[0]),.din(w_dff_A_B3WQpwTl4_0),.clk(gclk));
	jdff dff_A_0YemFUP72_0(.dout(w_dff_A_B3WQpwTl4_0),.din(w_dff_A_0YemFUP72_0),.clk(gclk));
	jdff dff_A_KRiL7IEK0_0(.dout(w_dff_A_0YemFUP72_0),.din(w_dff_A_KRiL7IEK0_0),.clk(gclk));
	jdff dff_A_GBy94EUE8_0(.dout(w_dff_A_KRiL7IEK0_0),.din(w_dff_A_GBy94EUE8_0),.clk(gclk));
	jdff dff_A_zaQIbnIG7_0(.dout(w_dff_A_GBy94EUE8_0),.din(w_dff_A_zaQIbnIG7_0),.clk(gclk));
	jdff dff_A_TRKK8lrZ0_0(.dout(w_dff_A_zaQIbnIG7_0),.din(w_dff_A_TRKK8lrZ0_0),.clk(gclk));
	jdff dff_A_fHLYcBzl5_0(.dout(w_dff_A_TRKK8lrZ0_0),.din(w_dff_A_fHLYcBzl5_0),.clk(gclk));
	jdff dff_A_jeGCbEct3_0(.dout(w_dff_A_fHLYcBzl5_0),.din(w_dff_A_jeGCbEct3_0),.clk(gclk));
	jdff dff_A_xwjJ8Hl73_0(.dout(w_dff_A_jeGCbEct3_0),.din(w_dff_A_xwjJ8Hl73_0),.clk(gclk));
	jdff dff_A_l0S9gEMM7_0(.dout(w_dff_A_xwjJ8Hl73_0),.din(w_dff_A_l0S9gEMM7_0),.clk(gclk));
	jdff dff_A_4eGXOV3D3_0(.dout(w_dff_A_l0S9gEMM7_0),.din(w_dff_A_4eGXOV3D3_0),.clk(gclk));
	jdff dff_A_A5zXeENM3_0(.dout(w_dff_A_4eGXOV3D3_0),.din(w_dff_A_A5zXeENM3_0),.clk(gclk));
	jdff dff_A_pH1V3gBq1_0(.dout(w_dff_A_A5zXeENM3_0),.din(w_dff_A_pH1V3gBq1_0),.clk(gclk));
	jdff dff_A_O5YybVCM4_0(.dout(w_dff_A_pH1V3gBq1_0),.din(w_dff_A_O5YybVCM4_0),.clk(gclk));
	jdff dff_A_AYkCkQii3_0(.dout(w_dff_A_O5YybVCM4_0),.din(w_dff_A_AYkCkQii3_0),.clk(gclk));
	jdff dff_A_E8GAXqDH7_0(.dout(w_dff_A_AYkCkQii3_0),.din(w_dff_A_E8GAXqDH7_0),.clk(gclk));
	jdff dff_A_6XWz6aFm8_0(.dout(w_dff_A_E8GAXqDH7_0),.din(w_dff_A_6XWz6aFm8_0),.clk(gclk));
	jdff dff_A_cC0z3G040_0(.dout(w_dff_A_6XWz6aFm8_0),.din(w_dff_A_cC0z3G040_0),.clk(gclk));
	jdff dff_A_5pWPVmoE9_0(.dout(w_dff_A_cC0z3G040_0),.din(w_dff_A_5pWPVmoE9_0),.clk(gclk));
	jdff dff_A_bWWMFQmV5_0(.dout(w_dff_A_5pWPVmoE9_0),.din(w_dff_A_bWWMFQmV5_0),.clk(gclk));
	jdff dff_A_vOuZa3lL8_0(.dout(w_n329_0[0]),.din(w_dff_A_vOuZa3lL8_0),.clk(gclk));
	jdff dff_B_t7zGmDAA3_1(.din(n285),.dout(w_dff_B_t7zGmDAA3_1),.clk(gclk));
	jdff dff_A_2UkcZ4Vf5_0(.dout(w_n232_0[0]),.din(w_dff_A_2UkcZ4Vf5_0),.clk(gclk));
	jdff dff_A_3tkynaLc6_0(.dout(w_dff_A_2UkcZ4Vf5_0),.din(w_dff_A_3tkynaLc6_0),.clk(gclk));
	jdff dff_A_Bn60p0gt6_0(.dout(w_dff_A_3tkynaLc6_0),.din(w_dff_A_Bn60p0gt6_0),.clk(gclk));
	jdff dff_A_LBSeKYrW7_0(.dout(w_dff_A_Bn60p0gt6_0),.din(w_dff_A_LBSeKYrW7_0),.clk(gclk));
	jdff dff_A_ktP54q1O9_0(.dout(w_dff_A_LBSeKYrW7_0),.din(w_dff_A_ktP54q1O9_0),.clk(gclk));
	jdff dff_A_oKlHnjZ98_0(.dout(w_dff_A_ktP54q1O9_0),.din(w_dff_A_oKlHnjZ98_0),.clk(gclk));
	jdff dff_A_5fnwKwEV0_0(.dout(w_dff_A_oKlHnjZ98_0),.din(w_dff_A_5fnwKwEV0_0),.clk(gclk));
	jdff dff_A_28cwp9BN3_0(.dout(w_dff_A_5fnwKwEV0_0),.din(w_dff_A_28cwp9BN3_0),.clk(gclk));
	jdff dff_A_TZyYsELy1_0(.dout(w_dff_A_28cwp9BN3_0),.din(w_dff_A_TZyYsELy1_0),.clk(gclk));
	jdff dff_A_PdIZnOZs0_0(.dout(w_dff_A_TZyYsELy1_0),.din(w_dff_A_PdIZnOZs0_0),.clk(gclk));
	jdff dff_A_qu5JsAQ68_0(.dout(w_dff_A_PdIZnOZs0_0),.din(w_dff_A_qu5JsAQ68_0),.clk(gclk));
	jdff dff_A_iIdUagJN7_0(.dout(w_dff_A_qu5JsAQ68_0),.din(w_dff_A_iIdUagJN7_0),.clk(gclk));
	jdff dff_A_7DmEP9vG1_0(.dout(w_dff_A_iIdUagJN7_0),.din(w_dff_A_7DmEP9vG1_0),.clk(gclk));
	jdff dff_A_QHMsashP2_0(.dout(w_dff_A_7DmEP9vG1_0),.din(w_dff_A_QHMsashP2_0),.clk(gclk));
	jdff dff_A_Z335YrJW3_0(.dout(w_dff_A_QHMsashP2_0),.din(w_dff_A_Z335YrJW3_0),.clk(gclk));
	jdff dff_A_YzF7m0cY7_0(.dout(w_dff_A_Z335YrJW3_0),.din(w_dff_A_YzF7m0cY7_0),.clk(gclk));
	jdff dff_A_Q4WRj3c35_0(.dout(w_dff_A_YzF7m0cY7_0),.din(w_dff_A_Q4WRj3c35_0),.clk(gclk));
	jdff dff_A_AoFzQpzy8_0(.dout(w_n271_0[0]),.din(w_dff_A_AoFzQpzy8_0),.clk(gclk));
	jdff dff_B_0Uuq0fZ45_1(.din(n234),.dout(w_dff_B_0Uuq0fZ45_1),.clk(gclk));
	jdff dff_A_2QI3qJVS2_0(.dout(w_n189_0[0]),.din(w_dff_A_2QI3qJVS2_0),.clk(gclk));
	jdff dff_A_4TwJTyUU2_0(.dout(w_dff_A_2QI3qJVS2_0),.din(w_dff_A_4TwJTyUU2_0),.clk(gclk));
	jdff dff_A_zxDsxLGi9_0(.dout(w_dff_A_4TwJTyUU2_0),.din(w_dff_A_zxDsxLGi9_0),.clk(gclk));
	jdff dff_A_lCKEQrTs5_0(.dout(w_dff_A_zxDsxLGi9_0),.din(w_dff_A_lCKEQrTs5_0),.clk(gclk));
	jdff dff_A_D7FM4cfR4_0(.dout(w_dff_A_lCKEQrTs5_0),.din(w_dff_A_D7FM4cfR4_0),.clk(gclk));
	jdff dff_A_bh17kYxA5_0(.dout(w_dff_A_D7FM4cfR4_0),.din(w_dff_A_bh17kYxA5_0),.clk(gclk));
	jdff dff_A_Y0CCq4A94_0(.dout(w_dff_A_bh17kYxA5_0),.din(w_dff_A_Y0CCq4A94_0),.clk(gclk));
	jdff dff_A_NK5EfVlx2_0(.dout(w_dff_A_Y0CCq4A94_0),.din(w_dff_A_NK5EfVlx2_0),.clk(gclk));
	jdff dff_A_dLqodMmE1_0(.dout(w_dff_A_NK5EfVlx2_0),.din(w_dff_A_dLqodMmE1_0),.clk(gclk));
	jdff dff_A_sagg0vuS4_0(.dout(w_dff_A_dLqodMmE1_0),.din(w_dff_A_sagg0vuS4_0),.clk(gclk));
	jdff dff_A_0LFcPuXD3_0(.dout(w_dff_A_sagg0vuS4_0),.din(w_dff_A_0LFcPuXD3_0),.clk(gclk));
	jdff dff_A_cKBBEiH61_0(.dout(w_dff_A_0LFcPuXD3_0),.din(w_dff_A_cKBBEiH61_0),.clk(gclk));
	jdff dff_A_NB7t1PsP8_0(.dout(w_dff_A_cKBBEiH61_0),.din(w_dff_A_NB7t1PsP8_0),.clk(gclk));
	jdff dff_A_E3uuICfZ1_0(.dout(w_dff_A_NB7t1PsP8_0),.din(w_dff_A_E3uuICfZ1_0),.clk(gclk));
	jdff dff_A_AGyhUYPC7_0(.dout(w_n220_0[0]),.din(w_dff_A_AGyhUYPC7_0),.clk(gclk));
	jdff dff_B_5lD7qqqs3_1(.din(n191),.dout(w_dff_B_5lD7qqqs3_1),.clk(gclk));
	jdff dff_A_AeuZPtDG8_0(.dout(w_n151_0[0]),.din(w_dff_A_AeuZPtDG8_0),.clk(gclk));
	jdff dff_A_vrALIgrq6_0(.dout(w_dff_A_AeuZPtDG8_0),.din(w_dff_A_vrALIgrq6_0),.clk(gclk));
	jdff dff_A_qH8KSHAO7_0(.dout(w_dff_A_vrALIgrq6_0),.din(w_dff_A_qH8KSHAO7_0),.clk(gclk));
	jdff dff_A_ilmxlb7E5_0(.dout(w_dff_A_qH8KSHAO7_0),.din(w_dff_A_ilmxlb7E5_0),.clk(gclk));
	jdff dff_A_ke8BPedF2_0(.dout(w_dff_A_ilmxlb7E5_0),.din(w_dff_A_ke8BPedF2_0),.clk(gclk));
	jdff dff_A_inHWBLTv5_0(.dout(w_dff_A_ke8BPedF2_0),.din(w_dff_A_inHWBLTv5_0),.clk(gclk));
	jdff dff_A_pccu4gh62_0(.dout(w_dff_A_inHWBLTv5_0),.din(w_dff_A_pccu4gh62_0),.clk(gclk));
	jdff dff_A_IbKovbYn7_0(.dout(w_dff_A_pccu4gh62_0),.din(w_dff_A_IbKovbYn7_0),.clk(gclk));
	jdff dff_A_fu6aqHvG5_0(.dout(w_dff_A_IbKovbYn7_0),.din(w_dff_A_fu6aqHvG5_0),.clk(gclk));
	jdff dff_A_0EY2T5k61_0(.dout(w_dff_A_fu6aqHvG5_0),.din(w_dff_A_0EY2T5k61_0),.clk(gclk));
	jdff dff_A_VWcmwtMh6_0(.dout(w_dff_A_0EY2T5k61_0),.din(w_dff_A_VWcmwtMh6_0),.clk(gclk));
	jdff dff_A_m59HVWWN7_0(.dout(w_n177_0[0]),.din(w_dff_A_m59HVWWN7_0),.clk(gclk));
	jdff dff_B_Mhfr6fth5_1(.din(n153),.dout(w_dff_B_Mhfr6fth5_1),.clk(gclk));
	jdff dff_A_hyLvjgaq0_0(.dout(w_n116_0[0]),.din(w_dff_A_hyLvjgaq0_0),.clk(gclk));
	jdff dff_A_fBk1XXtD8_0(.dout(w_dff_A_hyLvjgaq0_0),.din(w_dff_A_fBk1XXtD8_0),.clk(gclk));
	jdff dff_A_zOV19tar9_0(.dout(w_dff_A_fBk1XXtD8_0),.din(w_dff_A_zOV19tar9_0),.clk(gclk));
	jdff dff_A_cxfpP6D50_0(.dout(w_dff_A_zOV19tar9_0),.din(w_dff_A_cxfpP6D50_0),.clk(gclk));
	jdff dff_A_e9mREQgc5_0(.dout(w_dff_A_cxfpP6D50_0),.din(w_dff_A_e9mREQgc5_0),.clk(gclk));
	jdff dff_A_dDUC5QbX1_0(.dout(w_dff_A_e9mREQgc5_0),.din(w_dff_A_dDUC5QbX1_0),.clk(gclk));
	jdff dff_A_HeV4VCqy0_0(.dout(w_dff_A_dDUC5QbX1_0),.din(w_dff_A_HeV4VCqy0_0),.clk(gclk));
	jdff dff_A_lF7GCaFH7_0(.dout(w_dff_A_HeV4VCqy0_0),.din(w_dff_A_lF7GCaFH7_0),.clk(gclk));
	jdff dff_A_SZD2cvwN7_0(.dout(w_n139_0[0]),.din(w_dff_A_SZD2cvwN7_0),.clk(gclk));
	jdff dff_A_ykQi1sID8_0(.dout(w_n104_0[0]),.din(w_dff_A_ykQi1sID8_0),.clk(gclk));
	jdff dff_A_bcA037ij8_0(.dout(w_n85_0[0]),.din(w_dff_A_bcA037ij8_0),.clk(gclk));
	jdff dff_A_3cslWXqh6_1(.dout(w_n82_1[1]),.din(w_dff_A_3cslWXqh6_1),.clk(gclk));
	jdff dff_A_FWT5Eskw0_0(.dout(w_n94_0[0]),.din(w_dff_A_FWT5Eskw0_0),.clk(gclk));
	jdff dff_A_100ztZiO3_0(.dout(w_dff_A_FWT5Eskw0_0),.din(w_dff_A_100ztZiO3_0),.clk(gclk));
	jdff dff_A_rKcGLXn78_0(.dout(w_dff_A_100ztZiO3_0),.din(w_dff_A_rKcGLXn78_0),.clk(gclk));
	jdff dff_A_zmkCMecj4_0(.dout(w_dff_A_rKcGLXn78_0),.din(w_dff_A_zmkCMecj4_0),.clk(gclk));
	jdff dff_A_K0SsOrCV3_0(.dout(w_dff_A_zmkCMecj4_0),.din(w_dff_A_K0SsOrCV3_0),.clk(gclk));
	jdff dff_A_dpwNAxEi6_0(.dout(w_n103_0[0]),.din(w_dff_A_dpwNAxEi6_0),.clk(gclk));
	jdff dff_A_QvvnFDEe2_0(.dout(w_dff_A_dpwNAxEi6_0),.din(w_dff_A_QvvnFDEe2_0),.clk(gclk));
	jdff dff_B_GTzGY71r8_1(.din(n97),.dout(w_dff_B_GTzGY71r8_1),.clk(gclk));
	jdff dff_A_JJnjh7cr5_1(.dout(w_n82_0[1]),.din(w_dff_A_JJnjh7cr5_1),.clk(gclk));
	jdff dff_A_O3sEcoDA0_2(.dout(w_n82_0[2]),.din(w_dff_A_O3sEcoDA0_2),.clk(gclk));
	jdff dff_A_129vUXF14_2(.dout(w_dff_A_O3sEcoDA0_2),.din(w_dff_A_129vUXF14_2),.clk(gclk));
	jdff dff_A_58oNjSm74_0(.dout(w_n1151_0[0]),.din(w_dff_A_58oNjSm74_0),.clk(gclk));
	jdff dff_B_Xfkd7YaU7_2(.din(n1151),.dout(w_dff_B_Xfkd7YaU7_2),.clk(gclk));
	jdff dff_B_XYCnbEGk1_2(.din(n1044),.dout(w_dff_B_XYCnbEGk1_2),.clk(gclk));
	jdff dff_B_ALEJVILM3_2(.din(w_dff_B_XYCnbEGk1_2),.dout(w_dff_B_ALEJVILM3_2),.clk(gclk));
	jdff dff_B_hfXJN78t0_2(.din(w_dff_B_ALEJVILM3_2),.dout(w_dff_B_hfXJN78t0_2),.clk(gclk));
	jdff dff_B_IzVQw3Tg1_2(.din(w_dff_B_hfXJN78t0_2),.dout(w_dff_B_IzVQw3Tg1_2),.clk(gclk));
	jdff dff_B_86eJopzj1_2(.din(w_dff_B_IzVQw3Tg1_2),.dout(w_dff_B_86eJopzj1_2),.clk(gclk));
	jdff dff_B_z0CKpGcV5_2(.din(w_dff_B_86eJopzj1_2),.dout(w_dff_B_z0CKpGcV5_2),.clk(gclk));
	jdff dff_B_VQGFMzn25_2(.din(w_dff_B_z0CKpGcV5_2),.dout(w_dff_B_VQGFMzn25_2),.clk(gclk));
	jdff dff_B_pMLI55rQ1_2(.din(w_dff_B_VQGFMzn25_2),.dout(w_dff_B_pMLI55rQ1_2),.clk(gclk));
	jdff dff_B_W07sIFpL5_2(.din(w_dff_B_pMLI55rQ1_2),.dout(w_dff_B_W07sIFpL5_2),.clk(gclk));
	jdff dff_B_b4GITiFx9_2(.din(w_dff_B_W07sIFpL5_2),.dout(w_dff_B_b4GITiFx9_2),.clk(gclk));
	jdff dff_B_7vqDzFke6_2(.din(w_dff_B_b4GITiFx9_2),.dout(w_dff_B_7vqDzFke6_2),.clk(gclk));
	jdff dff_B_AFOV77Yp9_2(.din(w_dff_B_7vqDzFke6_2),.dout(w_dff_B_AFOV77Yp9_2),.clk(gclk));
	jdff dff_B_LLMZEDco8_2(.din(w_dff_B_AFOV77Yp9_2),.dout(w_dff_B_LLMZEDco8_2),.clk(gclk));
	jdff dff_B_IHcIAwtU1_2(.din(w_dff_B_LLMZEDco8_2),.dout(w_dff_B_IHcIAwtU1_2),.clk(gclk));
	jdff dff_B_SX5AH0VY9_2(.din(w_dff_B_IHcIAwtU1_2),.dout(w_dff_B_SX5AH0VY9_2),.clk(gclk));
	jdff dff_B_skJe9Cz49_2(.din(w_dff_B_SX5AH0VY9_2),.dout(w_dff_B_skJe9Cz49_2),.clk(gclk));
	jdff dff_B_GJkn4qjp1_2(.din(w_dff_B_skJe9Cz49_2),.dout(w_dff_B_GJkn4qjp1_2),.clk(gclk));
	jdff dff_B_klc7ieDe0_2(.din(w_dff_B_GJkn4qjp1_2),.dout(w_dff_B_klc7ieDe0_2),.clk(gclk));
	jdff dff_B_wwrrlaah7_2(.din(w_dff_B_klc7ieDe0_2),.dout(w_dff_B_wwrrlaah7_2),.clk(gclk));
	jdff dff_B_8JFqXxNQ4_2(.din(w_dff_B_wwrrlaah7_2),.dout(w_dff_B_8JFqXxNQ4_2),.clk(gclk));
	jdff dff_B_GXl8i9xh2_2(.din(w_dff_B_8JFqXxNQ4_2),.dout(w_dff_B_GXl8i9xh2_2),.clk(gclk));
	jdff dff_B_1XnU7mGy5_2(.din(w_dff_B_GXl8i9xh2_2),.dout(w_dff_B_1XnU7mGy5_2),.clk(gclk));
	jdff dff_B_7yYzIjPa6_2(.din(w_dff_B_1XnU7mGy5_2),.dout(w_dff_B_7yYzIjPa6_2),.clk(gclk));
	jdff dff_B_E2v58dEj9_2(.din(w_dff_B_7yYzIjPa6_2),.dout(w_dff_B_E2v58dEj9_2),.clk(gclk));
	jdff dff_B_GGvRfait7_2(.din(w_dff_B_E2v58dEj9_2),.dout(w_dff_B_GGvRfait7_2),.clk(gclk));
	jdff dff_B_8421x3Dt3_2(.din(w_dff_B_GGvRfait7_2),.dout(w_dff_B_8421x3Dt3_2),.clk(gclk));
	jdff dff_B_rIQAlWVs4_2(.din(w_dff_B_8421x3Dt3_2),.dout(w_dff_B_rIQAlWVs4_2),.clk(gclk));
	jdff dff_B_FV3ApBIe9_2(.din(w_dff_B_rIQAlWVs4_2),.dout(w_dff_B_FV3ApBIe9_2),.clk(gclk));
	jdff dff_B_9QeiNDJJ8_2(.din(w_dff_B_FV3ApBIe9_2),.dout(w_dff_B_9QeiNDJJ8_2),.clk(gclk));
	jdff dff_B_3Jm3eYIe2_2(.din(w_dff_B_9QeiNDJJ8_2),.dout(w_dff_B_3Jm3eYIe2_2),.clk(gclk));
	jdff dff_B_JaCMRJUa7_2(.din(w_dff_B_3Jm3eYIe2_2),.dout(w_dff_B_JaCMRJUa7_2),.clk(gclk));
	jdff dff_B_7gh0oi4N6_2(.din(w_dff_B_JaCMRJUa7_2),.dout(w_dff_B_7gh0oi4N6_2),.clk(gclk));
	jdff dff_B_YrVzFK9A7_2(.din(w_dff_B_7gh0oi4N6_2),.dout(w_dff_B_YrVzFK9A7_2),.clk(gclk));
	jdff dff_B_LseRDJ8k7_2(.din(w_dff_B_YrVzFK9A7_2),.dout(w_dff_B_LseRDJ8k7_2),.clk(gclk));
	jdff dff_B_aYL9nx0e2_2(.din(w_dff_B_LseRDJ8k7_2),.dout(w_dff_B_aYL9nx0e2_2),.clk(gclk));
	jdff dff_B_77BJru3w1_2(.din(w_dff_B_aYL9nx0e2_2),.dout(w_dff_B_77BJru3w1_2),.clk(gclk));
	jdff dff_B_210xLPz89_2(.din(w_dff_B_77BJru3w1_2),.dout(w_dff_B_210xLPz89_2),.clk(gclk));
	jdff dff_B_ai8Za3sR0_2(.din(w_dff_B_210xLPz89_2),.dout(w_dff_B_ai8Za3sR0_2),.clk(gclk));
	jdff dff_B_7stG2Ylw7_2(.din(w_dff_B_ai8Za3sR0_2),.dout(w_dff_B_7stG2Ylw7_2),.clk(gclk));
	jdff dff_B_rD4XypI92_2(.din(w_dff_B_7stG2Ylw7_2),.dout(w_dff_B_rD4XypI92_2),.clk(gclk));
	jdff dff_B_9k8wHymZ8_2(.din(w_dff_B_rD4XypI92_2),.dout(w_dff_B_9k8wHymZ8_2),.clk(gclk));
	jdff dff_B_si7ZQzf03_2(.din(w_dff_B_9k8wHymZ8_2),.dout(w_dff_B_si7ZQzf03_2),.clk(gclk));
	jdff dff_B_4MuhyZz56_2(.din(w_dff_B_si7ZQzf03_2),.dout(w_dff_B_4MuhyZz56_2),.clk(gclk));
	jdff dff_B_A3hoYYku9_2(.din(w_dff_B_4MuhyZz56_2),.dout(w_dff_B_A3hoYYku9_2),.clk(gclk));
	jdff dff_A_0WP8bNhx8_0(.dout(w_n1048_0[0]),.din(w_dff_A_0WP8bNhx8_0),.clk(gclk));
	jdff dff_B_ixj7yUiC0_1(.din(n1046),.dout(w_dff_B_ixj7yUiC0_1),.clk(gclk));
	jdff dff_B_RdEFjcEE0_2(.din(n943),.dout(w_dff_B_RdEFjcEE0_2),.clk(gclk));
	jdff dff_B_MV4bqQJz9_2(.din(w_dff_B_RdEFjcEE0_2),.dout(w_dff_B_MV4bqQJz9_2),.clk(gclk));
	jdff dff_B_ClRaOHsw9_2(.din(w_dff_B_MV4bqQJz9_2),.dout(w_dff_B_ClRaOHsw9_2),.clk(gclk));
	jdff dff_B_UHV0fyxY3_2(.din(w_dff_B_ClRaOHsw9_2),.dout(w_dff_B_UHV0fyxY3_2),.clk(gclk));
	jdff dff_B_dygcDZ8r6_2(.din(w_dff_B_UHV0fyxY3_2),.dout(w_dff_B_dygcDZ8r6_2),.clk(gclk));
	jdff dff_B_6TgLpY779_2(.din(w_dff_B_dygcDZ8r6_2),.dout(w_dff_B_6TgLpY779_2),.clk(gclk));
	jdff dff_B_ir36mJq39_2(.din(w_dff_B_6TgLpY779_2),.dout(w_dff_B_ir36mJq39_2),.clk(gclk));
	jdff dff_B_8JZxrxqd7_2(.din(w_dff_B_ir36mJq39_2),.dout(w_dff_B_8JZxrxqd7_2),.clk(gclk));
	jdff dff_B_qmho1tvv5_2(.din(w_dff_B_8JZxrxqd7_2),.dout(w_dff_B_qmho1tvv5_2),.clk(gclk));
	jdff dff_B_eA36qhs15_2(.din(w_dff_B_qmho1tvv5_2),.dout(w_dff_B_eA36qhs15_2),.clk(gclk));
	jdff dff_B_vKHAUT8B3_2(.din(w_dff_B_eA36qhs15_2),.dout(w_dff_B_vKHAUT8B3_2),.clk(gclk));
	jdff dff_B_NHDgziGL8_2(.din(w_dff_B_vKHAUT8B3_2),.dout(w_dff_B_NHDgziGL8_2),.clk(gclk));
	jdff dff_B_U12dkmG22_2(.din(w_dff_B_NHDgziGL8_2),.dout(w_dff_B_U12dkmG22_2),.clk(gclk));
	jdff dff_B_qYCAoU1x6_2(.din(w_dff_B_U12dkmG22_2),.dout(w_dff_B_qYCAoU1x6_2),.clk(gclk));
	jdff dff_B_P1FziXA14_2(.din(w_dff_B_qYCAoU1x6_2),.dout(w_dff_B_P1FziXA14_2),.clk(gclk));
	jdff dff_B_KtVatRyz5_2(.din(w_dff_B_P1FziXA14_2),.dout(w_dff_B_KtVatRyz5_2),.clk(gclk));
	jdff dff_B_manjh1NZ5_2(.din(w_dff_B_KtVatRyz5_2),.dout(w_dff_B_manjh1NZ5_2),.clk(gclk));
	jdff dff_B_QTwQ1JIM6_2(.din(w_dff_B_manjh1NZ5_2),.dout(w_dff_B_QTwQ1JIM6_2),.clk(gclk));
	jdff dff_B_9F3Cheqa6_2(.din(w_dff_B_QTwQ1JIM6_2),.dout(w_dff_B_9F3Cheqa6_2),.clk(gclk));
	jdff dff_B_wYumgaWL6_2(.din(w_dff_B_9F3Cheqa6_2),.dout(w_dff_B_wYumgaWL6_2),.clk(gclk));
	jdff dff_B_pCSDMmHc2_2(.din(w_dff_B_wYumgaWL6_2),.dout(w_dff_B_pCSDMmHc2_2),.clk(gclk));
	jdff dff_B_WLlRa5yB2_2(.din(w_dff_B_pCSDMmHc2_2),.dout(w_dff_B_WLlRa5yB2_2),.clk(gclk));
	jdff dff_B_RlF98wIe1_2(.din(w_dff_B_WLlRa5yB2_2),.dout(w_dff_B_RlF98wIe1_2),.clk(gclk));
	jdff dff_B_gSOEA2j56_2(.din(w_dff_B_RlF98wIe1_2),.dout(w_dff_B_gSOEA2j56_2),.clk(gclk));
	jdff dff_B_VXDqMmki5_2(.din(w_dff_B_gSOEA2j56_2),.dout(w_dff_B_VXDqMmki5_2),.clk(gclk));
	jdff dff_B_n8gUi5QA1_2(.din(w_dff_B_VXDqMmki5_2),.dout(w_dff_B_n8gUi5QA1_2),.clk(gclk));
	jdff dff_B_PX2sR0uv3_2(.din(w_dff_B_n8gUi5QA1_2),.dout(w_dff_B_PX2sR0uv3_2),.clk(gclk));
	jdff dff_B_ZQyEPytw4_2(.din(w_dff_B_PX2sR0uv3_2),.dout(w_dff_B_ZQyEPytw4_2),.clk(gclk));
	jdff dff_B_9bhBoudj2_2(.din(w_dff_B_ZQyEPytw4_2),.dout(w_dff_B_9bhBoudj2_2),.clk(gclk));
	jdff dff_B_CEJjXlkA2_2(.din(w_dff_B_9bhBoudj2_2),.dout(w_dff_B_CEJjXlkA2_2),.clk(gclk));
	jdff dff_B_irtCtgqt4_2(.din(w_dff_B_CEJjXlkA2_2),.dout(w_dff_B_irtCtgqt4_2),.clk(gclk));
	jdff dff_B_NtCTb9NO3_2(.din(w_dff_B_irtCtgqt4_2),.dout(w_dff_B_NtCTb9NO3_2),.clk(gclk));
	jdff dff_B_QAMRhUhQ1_2(.din(w_dff_B_NtCTb9NO3_2),.dout(w_dff_B_QAMRhUhQ1_2),.clk(gclk));
	jdff dff_B_L3KJJBar3_2(.din(w_dff_B_QAMRhUhQ1_2),.dout(w_dff_B_L3KJJBar3_2),.clk(gclk));
	jdff dff_B_X3hmDc9U0_2(.din(w_dff_B_L3KJJBar3_2),.dout(w_dff_B_X3hmDc9U0_2),.clk(gclk));
	jdff dff_B_t8a7mpJc1_2(.din(w_dff_B_X3hmDc9U0_2),.dout(w_dff_B_t8a7mpJc1_2),.clk(gclk));
	jdff dff_B_eakJ78K88_2(.din(w_dff_B_t8a7mpJc1_2),.dout(w_dff_B_eakJ78K88_2),.clk(gclk));
	jdff dff_B_7Stnel8r1_2(.din(w_dff_B_eakJ78K88_2),.dout(w_dff_B_7Stnel8r1_2),.clk(gclk));
	jdff dff_B_qFncmWYE3_2(.din(w_dff_B_7Stnel8r1_2),.dout(w_dff_B_qFncmWYE3_2),.clk(gclk));
	jdff dff_B_NK1cGy002_2(.din(w_dff_B_qFncmWYE3_2),.dout(w_dff_B_NK1cGy002_2),.clk(gclk));
	jdff dff_B_0RTT3rWU7_2(.din(w_dff_B_NK1cGy002_2),.dout(w_dff_B_0RTT3rWU7_2),.clk(gclk));
	jdff dff_A_LiLLaKQ70_1(.dout(w_n1032_0[1]),.din(w_dff_A_LiLLaKQ70_1),.clk(gclk));
	jdff dff_A_JVFZYS5k2_0(.dout(w_n840_0[0]),.din(w_dff_A_JVFZYS5k2_0),.clk(gclk));
	jdff dff_A_ThE4032i7_0(.dout(w_dff_A_JVFZYS5k2_0),.din(w_dff_A_ThE4032i7_0),.clk(gclk));
	jdff dff_A_b8dyL3Gc7_0(.dout(w_dff_A_ThE4032i7_0),.din(w_dff_A_b8dyL3Gc7_0),.clk(gclk));
	jdff dff_A_MFmMa0Sk5_0(.dout(w_dff_A_b8dyL3Gc7_0),.din(w_dff_A_MFmMa0Sk5_0),.clk(gclk));
	jdff dff_A_hNVLQOt59_0(.dout(w_dff_A_MFmMa0Sk5_0),.din(w_dff_A_hNVLQOt59_0),.clk(gclk));
	jdff dff_A_aNJzPPnh5_0(.dout(w_dff_A_hNVLQOt59_0),.din(w_dff_A_aNJzPPnh5_0),.clk(gclk));
	jdff dff_A_sTza9uYR8_0(.dout(w_dff_A_aNJzPPnh5_0),.din(w_dff_A_sTza9uYR8_0),.clk(gclk));
	jdff dff_A_ucZrvFil5_0(.dout(w_dff_A_sTza9uYR8_0),.din(w_dff_A_ucZrvFil5_0),.clk(gclk));
	jdff dff_A_rujyZHXO7_0(.dout(w_dff_A_ucZrvFil5_0),.din(w_dff_A_rujyZHXO7_0),.clk(gclk));
	jdff dff_A_BTuUOtKP4_0(.dout(w_dff_A_rujyZHXO7_0),.din(w_dff_A_BTuUOtKP4_0),.clk(gclk));
	jdff dff_A_oicvysoX1_0(.dout(w_dff_A_BTuUOtKP4_0),.din(w_dff_A_oicvysoX1_0),.clk(gclk));
	jdff dff_A_tmZXjUZJ1_0(.dout(w_dff_A_oicvysoX1_0),.din(w_dff_A_tmZXjUZJ1_0),.clk(gclk));
	jdff dff_A_OP2JCiGM7_0(.dout(w_dff_A_tmZXjUZJ1_0),.din(w_dff_A_OP2JCiGM7_0),.clk(gclk));
	jdff dff_A_X51ycMFW3_0(.dout(w_dff_A_OP2JCiGM7_0),.din(w_dff_A_X51ycMFW3_0),.clk(gclk));
	jdff dff_A_ulWJkAd52_0(.dout(w_dff_A_X51ycMFW3_0),.din(w_dff_A_ulWJkAd52_0),.clk(gclk));
	jdff dff_A_wBkthbbs3_0(.dout(w_dff_A_ulWJkAd52_0),.din(w_dff_A_wBkthbbs3_0),.clk(gclk));
	jdff dff_A_efQbvt229_0(.dout(w_dff_A_wBkthbbs3_0),.din(w_dff_A_efQbvt229_0),.clk(gclk));
	jdff dff_A_QeXAeT9f6_0(.dout(w_dff_A_efQbvt229_0),.din(w_dff_A_QeXAeT9f6_0),.clk(gclk));
	jdff dff_A_s7D7sebC2_0(.dout(w_dff_A_QeXAeT9f6_0),.din(w_dff_A_s7D7sebC2_0),.clk(gclk));
	jdff dff_A_x885c7Ue6_0(.dout(w_dff_A_s7D7sebC2_0),.din(w_dff_A_x885c7Ue6_0),.clk(gclk));
	jdff dff_A_wiavjYbC8_0(.dout(w_dff_A_x885c7Ue6_0),.din(w_dff_A_wiavjYbC8_0),.clk(gclk));
	jdff dff_A_qLhJBFLE0_0(.dout(w_dff_A_wiavjYbC8_0),.din(w_dff_A_qLhJBFLE0_0),.clk(gclk));
	jdff dff_A_1kIhnF6k7_0(.dout(w_dff_A_qLhJBFLE0_0),.din(w_dff_A_1kIhnF6k7_0),.clk(gclk));
	jdff dff_A_Z84DsC3x1_0(.dout(w_dff_A_1kIhnF6k7_0),.din(w_dff_A_Z84DsC3x1_0),.clk(gclk));
	jdff dff_A_O8e5PD9S4_0(.dout(w_dff_A_Z84DsC3x1_0),.din(w_dff_A_O8e5PD9S4_0),.clk(gclk));
	jdff dff_A_mxB2yEn90_0(.dout(w_dff_A_O8e5PD9S4_0),.din(w_dff_A_mxB2yEn90_0),.clk(gclk));
	jdff dff_A_VLDufczS1_0(.dout(w_dff_A_mxB2yEn90_0),.din(w_dff_A_VLDufczS1_0),.clk(gclk));
	jdff dff_A_tyScGpDV5_0(.dout(w_dff_A_VLDufczS1_0),.din(w_dff_A_tyScGpDV5_0),.clk(gclk));
	jdff dff_A_CrJ0yvYZ5_0(.dout(w_dff_A_tyScGpDV5_0),.din(w_dff_A_CrJ0yvYZ5_0),.clk(gclk));
	jdff dff_A_RrkunfDu4_0(.dout(w_dff_A_CrJ0yvYZ5_0),.din(w_dff_A_RrkunfDu4_0),.clk(gclk));
	jdff dff_A_BZnmWBMG8_0(.dout(w_dff_A_RrkunfDu4_0),.din(w_dff_A_BZnmWBMG8_0),.clk(gclk));
	jdff dff_A_JpAY9JLX4_0(.dout(w_dff_A_BZnmWBMG8_0),.din(w_dff_A_JpAY9JLX4_0),.clk(gclk));
	jdff dff_A_NN1WPiiH7_0(.dout(w_dff_A_JpAY9JLX4_0),.din(w_dff_A_NN1WPiiH7_0),.clk(gclk));
	jdff dff_A_ElRliAgJ8_0(.dout(w_dff_A_NN1WPiiH7_0),.din(w_dff_A_ElRliAgJ8_0),.clk(gclk));
	jdff dff_A_DqnCeYFm4_0(.dout(w_dff_A_ElRliAgJ8_0),.din(w_dff_A_DqnCeYFm4_0),.clk(gclk));
	jdff dff_A_Zrw86vAk2_0(.dout(w_dff_A_DqnCeYFm4_0),.din(w_dff_A_Zrw86vAk2_0),.clk(gclk));
	jdff dff_A_dfoK9Vu36_0(.dout(w_dff_A_Zrw86vAk2_0),.din(w_dff_A_dfoK9Vu36_0),.clk(gclk));
	jdff dff_A_PXYu4tFF2_0(.dout(w_dff_A_dfoK9Vu36_0),.din(w_dff_A_PXYu4tFF2_0),.clk(gclk));
	jdff dff_A_rNhfqppf1_1(.dout(w_n927_0[1]),.din(w_dff_A_rNhfqppf1_1),.clk(gclk));
	jdff dff_A_ERUtKZw50_2(.dout(w_n927_0[2]),.din(w_dff_A_ERUtKZw50_2),.clk(gclk));
	jdff dff_B_pFzgrlqQ6_1(.din(n842),.dout(w_dff_B_pFzgrlqQ6_1),.clk(gclk));
	jdff dff_B_aqLqSVbb5_2(.din(n742),.dout(w_dff_B_aqLqSVbb5_2),.clk(gclk));
	jdff dff_B_8TtlUCFZ6_2(.din(w_dff_B_aqLqSVbb5_2),.dout(w_dff_B_8TtlUCFZ6_2),.clk(gclk));
	jdff dff_B_fGoWAijM3_2(.din(w_dff_B_8TtlUCFZ6_2),.dout(w_dff_B_fGoWAijM3_2),.clk(gclk));
	jdff dff_B_LX6g5d3q0_2(.din(w_dff_B_fGoWAijM3_2),.dout(w_dff_B_LX6g5d3q0_2),.clk(gclk));
	jdff dff_B_OxgyoqTX1_2(.din(w_dff_B_LX6g5d3q0_2),.dout(w_dff_B_OxgyoqTX1_2),.clk(gclk));
	jdff dff_B_ePUgQZSz9_2(.din(w_dff_B_OxgyoqTX1_2),.dout(w_dff_B_ePUgQZSz9_2),.clk(gclk));
	jdff dff_B_855WPIpP8_2(.din(w_dff_B_ePUgQZSz9_2),.dout(w_dff_B_855WPIpP8_2),.clk(gclk));
	jdff dff_B_1SLzG1sJ8_2(.din(w_dff_B_855WPIpP8_2),.dout(w_dff_B_1SLzG1sJ8_2),.clk(gclk));
	jdff dff_B_ZONFmFUc2_2(.din(w_dff_B_1SLzG1sJ8_2),.dout(w_dff_B_ZONFmFUc2_2),.clk(gclk));
	jdff dff_B_zgrMX4vu2_2(.din(w_dff_B_ZONFmFUc2_2),.dout(w_dff_B_zgrMX4vu2_2),.clk(gclk));
	jdff dff_B_CWoryAm58_2(.din(w_dff_B_zgrMX4vu2_2),.dout(w_dff_B_CWoryAm58_2),.clk(gclk));
	jdff dff_B_8PI4HxTW1_2(.din(w_dff_B_CWoryAm58_2),.dout(w_dff_B_8PI4HxTW1_2),.clk(gclk));
	jdff dff_B_W565hlja3_2(.din(w_dff_B_8PI4HxTW1_2),.dout(w_dff_B_W565hlja3_2),.clk(gclk));
	jdff dff_B_goC2GtdM8_2(.din(w_dff_B_W565hlja3_2),.dout(w_dff_B_goC2GtdM8_2),.clk(gclk));
	jdff dff_B_zglewjTh2_2(.din(w_dff_B_goC2GtdM8_2),.dout(w_dff_B_zglewjTh2_2),.clk(gclk));
	jdff dff_B_NCfsaHxY3_2(.din(w_dff_B_zglewjTh2_2),.dout(w_dff_B_NCfsaHxY3_2),.clk(gclk));
	jdff dff_B_izzFwD9P7_2(.din(w_dff_B_NCfsaHxY3_2),.dout(w_dff_B_izzFwD9P7_2),.clk(gclk));
	jdff dff_B_jcVvnAzP3_2(.din(w_dff_B_izzFwD9P7_2),.dout(w_dff_B_jcVvnAzP3_2),.clk(gclk));
	jdff dff_B_V8ljW9QM2_2(.din(w_dff_B_jcVvnAzP3_2),.dout(w_dff_B_V8ljW9QM2_2),.clk(gclk));
	jdff dff_B_RiDZEjDY7_2(.din(w_dff_B_V8ljW9QM2_2),.dout(w_dff_B_RiDZEjDY7_2),.clk(gclk));
	jdff dff_B_PiUefMaQ9_2(.din(w_dff_B_RiDZEjDY7_2),.dout(w_dff_B_PiUefMaQ9_2),.clk(gclk));
	jdff dff_B_l17r3wle0_2(.din(w_dff_B_PiUefMaQ9_2),.dout(w_dff_B_l17r3wle0_2),.clk(gclk));
	jdff dff_B_pjpfPEhq9_2(.din(w_dff_B_l17r3wle0_2),.dout(w_dff_B_pjpfPEhq9_2),.clk(gclk));
	jdff dff_B_DVx2s3wq5_2(.din(w_dff_B_pjpfPEhq9_2),.dout(w_dff_B_DVx2s3wq5_2),.clk(gclk));
	jdff dff_B_73GQfmpV4_2(.din(w_dff_B_DVx2s3wq5_2),.dout(w_dff_B_73GQfmpV4_2),.clk(gclk));
	jdff dff_B_iiZJ8oQK7_2(.din(w_dff_B_73GQfmpV4_2),.dout(w_dff_B_iiZJ8oQK7_2),.clk(gclk));
	jdff dff_B_ETLGqHFC0_2(.din(w_dff_B_iiZJ8oQK7_2),.dout(w_dff_B_ETLGqHFC0_2),.clk(gclk));
	jdff dff_B_wuc06J5x0_2(.din(w_dff_B_ETLGqHFC0_2),.dout(w_dff_B_wuc06J5x0_2),.clk(gclk));
	jdff dff_B_2mWbSJ3u6_2(.din(w_dff_B_wuc06J5x0_2),.dout(w_dff_B_2mWbSJ3u6_2),.clk(gclk));
	jdff dff_B_UVLb67d54_2(.din(w_dff_B_2mWbSJ3u6_2),.dout(w_dff_B_UVLb67d54_2),.clk(gclk));
	jdff dff_B_dXYrXhlm3_2(.din(w_dff_B_UVLb67d54_2),.dout(w_dff_B_dXYrXhlm3_2),.clk(gclk));
	jdff dff_B_sNZ6qBcz6_2(.din(w_dff_B_dXYrXhlm3_2),.dout(w_dff_B_sNZ6qBcz6_2),.clk(gclk));
	jdff dff_B_GSt3l0oj2_2(.din(w_dff_B_sNZ6qBcz6_2),.dout(w_dff_B_GSt3l0oj2_2),.clk(gclk));
	jdff dff_B_CGzaqclw9_2(.din(w_dff_B_GSt3l0oj2_2),.dout(w_dff_B_CGzaqclw9_2),.clk(gclk));
	jdff dff_B_lsaBQh7J8_2(.din(n821),.dout(w_dff_B_lsaBQh7J8_2),.clk(gclk));
	jdff dff_B_YFGLmNff5_1(.din(n743),.dout(w_dff_B_YFGLmNff5_1),.clk(gclk));
	jdff dff_B_qjeV4zON2_2(.din(n649),.dout(w_dff_B_qjeV4zON2_2),.clk(gclk));
	jdff dff_B_8R7Ti3qY2_2(.din(w_dff_B_qjeV4zON2_2),.dout(w_dff_B_8R7Ti3qY2_2),.clk(gclk));
	jdff dff_B_84YqnIUj2_2(.din(w_dff_B_8R7Ti3qY2_2),.dout(w_dff_B_84YqnIUj2_2),.clk(gclk));
	jdff dff_B_IJnCaoWh3_2(.din(w_dff_B_84YqnIUj2_2),.dout(w_dff_B_IJnCaoWh3_2),.clk(gclk));
	jdff dff_B_0OEM80xx5_2(.din(w_dff_B_IJnCaoWh3_2),.dout(w_dff_B_0OEM80xx5_2),.clk(gclk));
	jdff dff_B_uV6ZS0iu8_2(.din(w_dff_B_0OEM80xx5_2),.dout(w_dff_B_uV6ZS0iu8_2),.clk(gclk));
	jdff dff_B_6Y0S37xe5_2(.din(w_dff_B_uV6ZS0iu8_2),.dout(w_dff_B_6Y0S37xe5_2),.clk(gclk));
	jdff dff_B_lHV9p9xl7_2(.din(w_dff_B_6Y0S37xe5_2),.dout(w_dff_B_lHV9p9xl7_2),.clk(gclk));
	jdff dff_B_8REZEnvQ1_2(.din(w_dff_B_lHV9p9xl7_2),.dout(w_dff_B_8REZEnvQ1_2),.clk(gclk));
	jdff dff_B_VqROLeH34_2(.din(w_dff_B_8REZEnvQ1_2),.dout(w_dff_B_VqROLeH34_2),.clk(gclk));
	jdff dff_B_ogbzXqZ74_2(.din(w_dff_B_VqROLeH34_2),.dout(w_dff_B_ogbzXqZ74_2),.clk(gclk));
	jdff dff_B_t8uPvq429_2(.din(w_dff_B_ogbzXqZ74_2),.dout(w_dff_B_t8uPvq429_2),.clk(gclk));
	jdff dff_B_JaALiz3y5_2(.din(w_dff_B_t8uPvq429_2),.dout(w_dff_B_JaALiz3y5_2),.clk(gclk));
	jdff dff_B_nRCTL3CB6_2(.din(w_dff_B_JaALiz3y5_2),.dout(w_dff_B_nRCTL3CB6_2),.clk(gclk));
	jdff dff_B_rZWLath03_2(.din(w_dff_B_nRCTL3CB6_2),.dout(w_dff_B_rZWLath03_2),.clk(gclk));
	jdff dff_B_8235HZRe8_2(.din(w_dff_B_rZWLath03_2),.dout(w_dff_B_8235HZRe8_2),.clk(gclk));
	jdff dff_B_vj6GeHQl1_2(.din(w_dff_B_8235HZRe8_2),.dout(w_dff_B_vj6GeHQl1_2),.clk(gclk));
	jdff dff_B_wWrx1rJ38_2(.din(w_dff_B_vj6GeHQl1_2),.dout(w_dff_B_wWrx1rJ38_2),.clk(gclk));
	jdff dff_B_fYft93dk1_2(.din(w_dff_B_wWrx1rJ38_2),.dout(w_dff_B_fYft93dk1_2),.clk(gclk));
	jdff dff_B_3JYrxhaL4_2(.din(w_dff_B_fYft93dk1_2),.dout(w_dff_B_3JYrxhaL4_2),.clk(gclk));
	jdff dff_B_wNm6FKIX1_2(.din(w_dff_B_3JYrxhaL4_2),.dout(w_dff_B_wNm6FKIX1_2),.clk(gclk));
	jdff dff_B_2itOObFF4_2(.din(w_dff_B_wNm6FKIX1_2),.dout(w_dff_B_2itOObFF4_2),.clk(gclk));
	jdff dff_B_Rzkg6iNm6_2(.din(w_dff_B_2itOObFF4_2),.dout(w_dff_B_Rzkg6iNm6_2),.clk(gclk));
	jdff dff_B_MkZbSH8v5_2(.din(w_dff_B_Rzkg6iNm6_2),.dout(w_dff_B_MkZbSH8v5_2),.clk(gclk));
	jdff dff_B_LwCJR8VV8_2(.din(w_dff_B_MkZbSH8v5_2),.dout(w_dff_B_LwCJR8VV8_2),.clk(gclk));
	jdff dff_B_oPY21CCQ4_2(.din(w_dff_B_LwCJR8VV8_2),.dout(w_dff_B_oPY21CCQ4_2),.clk(gclk));
	jdff dff_B_vMqCSAr18_2(.din(w_dff_B_oPY21CCQ4_2),.dout(w_dff_B_vMqCSAr18_2),.clk(gclk));
	jdff dff_B_vkit0yNc5_2(.din(w_dff_B_vMqCSAr18_2),.dout(w_dff_B_vkit0yNc5_2),.clk(gclk));
	jdff dff_B_LoFVokDw9_2(.din(w_dff_B_vkit0yNc5_2),.dout(w_dff_B_LoFVokDw9_2),.clk(gclk));
	jdff dff_B_JaDhI1AO8_2(.din(w_dff_B_LoFVokDw9_2),.dout(w_dff_B_JaDhI1AO8_2),.clk(gclk));
	jdff dff_B_ZYWG448Y6_2(.din(w_dff_B_JaDhI1AO8_2),.dout(w_dff_B_ZYWG448Y6_2),.clk(gclk));
	jdff dff_B_XMyO4VcL9_2(.din(n721),.dout(w_dff_B_XMyO4VcL9_2),.clk(gclk));
	jdff dff_B_p7A5tY8K4_1(.din(n650),.dout(w_dff_B_p7A5tY8K4_1),.clk(gclk));
	jdff dff_B_SWE7pXwo9_2(.din(n563),.dout(w_dff_B_SWE7pXwo9_2),.clk(gclk));
	jdff dff_B_lOav3PfN0_2(.din(w_dff_B_SWE7pXwo9_2),.dout(w_dff_B_lOav3PfN0_2),.clk(gclk));
	jdff dff_B_wFYf2lav8_2(.din(w_dff_B_lOav3PfN0_2),.dout(w_dff_B_wFYf2lav8_2),.clk(gclk));
	jdff dff_B_HZIKFsvb9_2(.din(w_dff_B_wFYf2lav8_2),.dout(w_dff_B_HZIKFsvb9_2),.clk(gclk));
	jdff dff_B_R488Rsjb9_2(.din(w_dff_B_HZIKFsvb9_2),.dout(w_dff_B_R488Rsjb9_2),.clk(gclk));
	jdff dff_B_098UAozT5_2(.din(w_dff_B_R488Rsjb9_2),.dout(w_dff_B_098UAozT5_2),.clk(gclk));
	jdff dff_B_iFUaAVA13_2(.din(w_dff_B_098UAozT5_2),.dout(w_dff_B_iFUaAVA13_2),.clk(gclk));
	jdff dff_B_IWrhjz9Z0_2(.din(w_dff_B_iFUaAVA13_2),.dout(w_dff_B_IWrhjz9Z0_2),.clk(gclk));
	jdff dff_B_4J5QOlcx4_2(.din(w_dff_B_IWrhjz9Z0_2),.dout(w_dff_B_4J5QOlcx4_2),.clk(gclk));
	jdff dff_B_xfOBvoTR5_2(.din(w_dff_B_4J5QOlcx4_2),.dout(w_dff_B_xfOBvoTR5_2),.clk(gclk));
	jdff dff_B_03J3pO6K2_2(.din(w_dff_B_xfOBvoTR5_2),.dout(w_dff_B_03J3pO6K2_2),.clk(gclk));
	jdff dff_B_aZn31KFm0_2(.din(w_dff_B_03J3pO6K2_2),.dout(w_dff_B_aZn31KFm0_2),.clk(gclk));
	jdff dff_B_226Xofee5_2(.din(w_dff_B_aZn31KFm0_2),.dout(w_dff_B_226Xofee5_2),.clk(gclk));
	jdff dff_B_lhKvZDVA2_2(.din(w_dff_B_226Xofee5_2),.dout(w_dff_B_lhKvZDVA2_2),.clk(gclk));
	jdff dff_B_itQyYcEO2_2(.din(w_dff_B_lhKvZDVA2_2),.dout(w_dff_B_itQyYcEO2_2),.clk(gclk));
	jdff dff_B_v2OoYA8f8_2(.din(w_dff_B_itQyYcEO2_2),.dout(w_dff_B_v2OoYA8f8_2),.clk(gclk));
	jdff dff_B_w06hzSZz7_2(.din(w_dff_B_v2OoYA8f8_2),.dout(w_dff_B_w06hzSZz7_2),.clk(gclk));
	jdff dff_B_TVmd71Bt5_2(.din(w_dff_B_w06hzSZz7_2),.dout(w_dff_B_TVmd71Bt5_2),.clk(gclk));
	jdff dff_B_gAUP2gyM6_2(.din(w_dff_B_TVmd71Bt5_2),.dout(w_dff_B_gAUP2gyM6_2),.clk(gclk));
	jdff dff_B_pGZDE7MI4_2(.din(w_dff_B_gAUP2gyM6_2),.dout(w_dff_B_pGZDE7MI4_2),.clk(gclk));
	jdff dff_B_FF3Y9FHH8_2(.din(w_dff_B_pGZDE7MI4_2),.dout(w_dff_B_FF3Y9FHH8_2),.clk(gclk));
	jdff dff_B_TlxNAIKP7_2(.din(w_dff_B_FF3Y9FHH8_2),.dout(w_dff_B_TlxNAIKP7_2),.clk(gclk));
	jdff dff_B_uSV59Dl34_2(.din(w_dff_B_TlxNAIKP7_2),.dout(w_dff_B_uSV59Dl34_2),.clk(gclk));
	jdff dff_B_r445SAU90_2(.din(w_dff_B_uSV59Dl34_2),.dout(w_dff_B_r445SAU90_2),.clk(gclk));
	jdff dff_B_pWXeHk9R5_2(.din(w_dff_B_r445SAU90_2),.dout(w_dff_B_pWXeHk9R5_2),.clk(gclk));
	jdff dff_B_sVujVXx70_2(.din(w_dff_B_pWXeHk9R5_2),.dout(w_dff_B_sVujVXx70_2),.clk(gclk));
	jdff dff_B_IvwcZuZ52_2(.din(w_dff_B_sVujVXx70_2),.dout(w_dff_B_IvwcZuZ52_2),.clk(gclk));
	jdff dff_B_IqjvnNs23_2(.din(w_dff_B_IvwcZuZ52_2),.dout(w_dff_B_IqjvnNs23_2),.clk(gclk));
	jdff dff_B_A0EP2u038_2(.din(n628),.dout(w_dff_B_A0EP2u038_2),.clk(gclk));
	jdff dff_B_LdbHXJz70_1(.din(n564),.dout(w_dff_B_LdbHXJz70_1),.clk(gclk));
	jdff dff_B_remLdU3W7_2(.din(n484),.dout(w_dff_B_remLdU3W7_2),.clk(gclk));
	jdff dff_B_nSCTjnSp5_2(.din(w_dff_B_remLdU3W7_2),.dout(w_dff_B_nSCTjnSp5_2),.clk(gclk));
	jdff dff_B_EmZUjoei5_2(.din(w_dff_B_nSCTjnSp5_2),.dout(w_dff_B_EmZUjoei5_2),.clk(gclk));
	jdff dff_B_kzvdLuxQ4_2(.din(w_dff_B_EmZUjoei5_2),.dout(w_dff_B_kzvdLuxQ4_2),.clk(gclk));
	jdff dff_B_j0nqz0qI3_2(.din(w_dff_B_kzvdLuxQ4_2),.dout(w_dff_B_j0nqz0qI3_2),.clk(gclk));
	jdff dff_B_UF4stipx1_2(.din(w_dff_B_j0nqz0qI3_2),.dout(w_dff_B_UF4stipx1_2),.clk(gclk));
	jdff dff_B_Ong0mR9n3_2(.din(w_dff_B_UF4stipx1_2),.dout(w_dff_B_Ong0mR9n3_2),.clk(gclk));
	jdff dff_B_BoG9dJsj3_2(.din(w_dff_B_Ong0mR9n3_2),.dout(w_dff_B_BoG9dJsj3_2),.clk(gclk));
	jdff dff_B_4l8CMNvt4_2(.din(w_dff_B_BoG9dJsj3_2),.dout(w_dff_B_4l8CMNvt4_2),.clk(gclk));
	jdff dff_B_0AtmG2Cn7_2(.din(w_dff_B_4l8CMNvt4_2),.dout(w_dff_B_0AtmG2Cn7_2),.clk(gclk));
	jdff dff_B_vaaTdudL8_2(.din(w_dff_B_0AtmG2Cn7_2),.dout(w_dff_B_vaaTdudL8_2),.clk(gclk));
	jdff dff_B_fJqk2wzJ0_2(.din(w_dff_B_vaaTdudL8_2),.dout(w_dff_B_fJqk2wzJ0_2),.clk(gclk));
	jdff dff_B_FPlSDfho2_2(.din(w_dff_B_fJqk2wzJ0_2),.dout(w_dff_B_FPlSDfho2_2),.clk(gclk));
	jdff dff_B_FukND1Vq8_2(.din(w_dff_B_FPlSDfho2_2),.dout(w_dff_B_FukND1Vq8_2),.clk(gclk));
	jdff dff_B_g0Om3uaU4_2(.din(w_dff_B_FukND1Vq8_2),.dout(w_dff_B_g0Om3uaU4_2),.clk(gclk));
	jdff dff_B_Pj0dZwwN3_2(.din(w_dff_B_g0Om3uaU4_2),.dout(w_dff_B_Pj0dZwwN3_2),.clk(gclk));
	jdff dff_B_Bh7jb3Mx6_2(.din(w_dff_B_Pj0dZwwN3_2),.dout(w_dff_B_Bh7jb3Mx6_2),.clk(gclk));
	jdff dff_B_ffTQWIFS5_2(.din(w_dff_B_Bh7jb3Mx6_2),.dout(w_dff_B_ffTQWIFS5_2),.clk(gclk));
	jdff dff_B_wLMNGDU23_2(.din(w_dff_B_ffTQWIFS5_2),.dout(w_dff_B_wLMNGDU23_2),.clk(gclk));
	jdff dff_B_A3BrkMmV3_2(.din(w_dff_B_wLMNGDU23_2),.dout(w_dff_B_A3BrkMmV3_2),.clk(gclk));
	jdff dff_B_gSujsVYH1_2(.din(w_dff_B_A3BrkMmV3_2),.dout(w_dff_B_gSujsVYH1_2),.clk(gclk));
	jdff dff_B_qErqbt8q0_2(.din(w_dff_B_gSujsVYH1_2),.dout(w_dff_B_qErqbt8q0_2),.clk(gclk));
	jdff dff_B_fOtmj0Vl2_2(.din(w_dff_B_qErqbt8q0_2),.dout(w_dff_B_fOtmj0Vl2_2),.clk(gclk));
	jdff dff_B_G3PK9Dmz9_2(.din(w_dff_B_fOtmj0Vl2_2),.dout(w_dff_B_G3PK9Dmz9_2),.clk(gclk));
	jdff dff_B_YZsqRtp03_2(.din(w_dff_B_G3PK9Dmz9_2),.dout(w_dff_B_YZsqRtp03_2),.clk(gclk));
	jdff dff_B_ahnDQaUE2_2(.din(n542),.dout(w_dff_B_ahnDQaUE2_2),.clk(gclk));
	jdff dff_B_VdB4vGKp5_1(.din(n485),.dout(w_dff_B_VdB4vGKp5_1),.clk(gclk));
	jdff dff_B_2VwStOel9_2(.din(n412),.dout(w_dff_B_2VwStOel9_2),.clk(gclk));
	jdff dff_B_kLxdcguU7_2(.din(w_dff_B_2VwStOel9_2),.dout(w_dff_B_kLxdcguU7_2),.clk(gclk));
	jdff dff_B_7jOyGxjd9_2(.din(w_dff_B_kLxdcguU7_2),.dout(w_dff_B_7jOyGxjd9_2),.clk(gclk));
	jdff dff_B_iAYneITv0_2(.din(w_dff_B_7jOyGxjd9_2),.dout(w_dff_B_iAYneITv0_2),.clk(gclk));
	jdff dff_B_7W1gMF8E6_2(.din(w_dff_B_iAYneITv0_2),.dout(w_dff_B_7W1gMF8E6_2),.clk(gclk));
	jdff dff_B_4heQCxFT6_2(.din(w_dff_B_7W1gMF8E6_2),.dout(w_dff_B_4heQCxFT6_2),.clk(gclk));
	jdff dff_B_BmKSXrJd4_2(.din(w_dff_B_4heQCxFT6_2),.dout(w_dff_B_BmKSXrJd4_2),.clk(gclk));
	jdff dff_B_YIhP0J3W2_2(.din(w_dff_B_BmKSXrJd4_2),.dout(w_dff_B_YIhP0J3W2_2),.clk(gclk));
	jdff dff_B_DxH8y57k0_2(.din(w_dff_B_YIhP0J3W2_2),.dout(w_dff_B_DxH8y57k0_2),.clk(gclk));
	jdff dff_B_DxkGXL4K2_2(.din(w_dff_B_DxH8y57k0_2),.dout(w_dff_B_DxkGXL4K2_2),.clk(gclk));
	jdff dff_B_LG1DRUM75_2(.din(w_dff_B_DxkGXL4K2_2),.dout(w_dff_B_LG1DRUM75_2),.clk(gclk));
	jdff dff_B_gwkAKuOX3_2(.din(w_dff_B_LG1DRUM75_2),.dout(w_dff_B_gwkAKuOX3_2),.clk(gclk));
	jdff dff_B_HZIXzl9R1_2(.din(w_dff_B_gwkAKuOX3_2),.dout(w_dff_B_HZIXzl9R1_2),.clk(gclk));
	jdff dff_B_t0YiUaOj3_2(.din(w_dff_B_HZIXzl9R1_2),.dout(w_dff_B_t0YiUaOj3_2),.clk(gclk));
	jdff dff_B_XaEkSQOJ5_2(.din(w_dff_B_t0YiUaOj3_2),.dout(w_dff_B_XaEkSQOJ5_2),.clk(gclk));
	jdff dff_B_Ieuytx2k1_2(.din(w_dff_B_XaEkSQOJ5_2),.dout(w_dff_B_Ieuytx2k1_2),.clk(gclk));
	jdff dff_B_rVH2xRnM3_2(.din(w_dff_B_Ieuytx2k1_2),.dout(w_dff_B_rVH2xRnM3_2),.clk(gclk));
	jdff dff_B_MNSiRIMK9_2(.din(w_dff_B_rVH2xRnM3_2),.dout(w_dff_B_MNSiRIMK9_2),.clk(gclk));
	jdff dff_B_gIFGXc919_2(.din(w_dff_B_MNSiRIMK9_2),.dout(w_dff_B_gIFGXc919_2),.clk(gclk));
	jdff dff_B_CrCxR1cm2_2(.din(w_dff_B_gIFGXc919_2),.dout(w_dff_B_CrCxR1cm2_2),.clk(gclk));
	jdff dff_B_gQ6syMS02_2(.din(w_dff_B_CrCxR1cm2_2),.dout(w_dff_B_gQ6syMS02_2),.clk(gclk));
	jdff dff_B_B1MHIwkE4_2(.din(w_dff_B_gQ6syMS02_2),.dout(w_dff_B_B1MHIwkE4_2),.clk(gclk));
	jdff dff_B_oai99Er00_2(.din(n463),.dout(w_dff_B_oai99Er00_2),.clk(gclk));
	jdff dff_B_Ha01Stdo7_1(.din(n413),.dout(w_dff_B_Ha01Stdo7_1),.clk(gclk));
	jdff dff_B_kPzXdT731_2(.din(n348),.dout(w_dff_B_kPzXdT731_2),.clk(gclk));
	jdff dff_B_rtyGdkVm1_2(.din(w_dff_B_kPzXdT731_2),.dout(w_dff_B_rtyGdkVm1_2),.clk(gclk));
	jdff dff_B_vhAZV4Tc4_2(.din(w_dff_B_rtyGdkVm1_2),.dout(w_dff_B_vhAZV4Tc4_2),.clk(gclk));
	jdff dff_B_gWd43pn36_2(.din(w_dff_B_vhAZV4Tc4_2),.dout(w_dff_B_gWd43pn36_2),.clk(gclk));
	jdff dff_B_ZdFhonGr4_2(.din(w_dff_B_gWd43pn36_2),.dout(w_dff_B_ZdFhonGr4_2),.clk(gclk));
	jdff dff_B_Rtwqnh0h5_2(.din(w_dff_B_ZdFhonGr4_2),.dout(w_dff_B_Rtwqnh0h5_2),.clk(gclk));
	jdff dff_B_HNe5PlZm0_2(.din(w_dff_B_Rtwqnh0h5_2),.dout(w_dff_B_HNe5PlZm0_2),.clk(gclk));
	jdff dff_B_3SxQLx4g3_2(.din(w_dff_B_HNe5PlZm0_2),.dout(w_dff_B_3SxQLx4g3_2),.clk(gclk));
	jdff dff_B_okHSrSDq9_2(.din(w_dff_B_3SxQLx4g3_2),.dout(w_dff_B_okHSrSDq9_2),.clk(gclk));
	jdff dff_B_3B9sHaTO1_2(.din(w_dff_B_okHSrSDq9_2),.dout(w_dff_B_3B9sHaTO1_2),.clk(gclk));
	jdff dff_B_jpsQrg4H5_2(.din(w_dff_B_3B9sHaTO1_2),.dout(w_dff_B_jpsQrg4H5_2),.clk(gclk));
	jdff dff_B_DsHnBPqt4_2(.din(w_dff_B_jpsQrg4H5_2),.dout(w_dff_B_DsHnBPqt4_2),.clk(gclk));
	jdff dff_B_jZdjHIib2_2(.din(w_dff_B_DsHnBPqt4_2),.dout(w_dff_B_jZdjHIib2_2),.clk(gclk));
	jdff dff_B_DBAuNXme7_2(.din(w_dff_B_jZdjHIib2_2),.dout(w_dff_B_DBAuNXme7_2),.clk(gclk));
	jdff dff_B_Z1xPljwx3_2(.din(w_dff_B_DBAuNXme7_2),.dout(w_dff_B_Z1xPljwx3_2),.clk(gclk));
	jdff dff_B_a779KKf65_2(.din(w_dff_B_Z1xPljwx3_2),.dout(w_dff_B_a779KKf65_2),.clk(gclk));
	jdff dff_B_t1I5GBDE3_2(.din(w_dff_B_a779KKf65_2),.dout(w_dff_B_t1I5GBDE3_2),.clk(gclk));
	jdff dff_B_pLjYX2P31_2(.din(w_dff_B_t1I5GBDE3_2),.dout(w_dff_B_pLjYX2P31_2),.clk(gclk));
	jdff dff_B_Jv3A2qaZ9_2(.din(w_dff_B_pLjYX2P31_2),.dout(w_dff_B_Jv3A2qaZ9_2),.clk(gclk));
	jdff dff_B_rbZL3TVO2_2(.din(n391),.dout(w_dff_B_rbZL3TVO2_2),.clk(gclk));
	jdff dff_B_QhBkAYhP6_1(.din(n349),.dout(w_dff_B_QhBkAYhP6_1),.clk(gclk));
	jdff dff_B_3yKfvuf39_2(.din(n290),.dout(w_dff_B_3yKfvuf39_2),.clk(gclk));
	jdff dff_B_QAyCvtyq7_2(.din(w_dff_B_3yKfvuf39_2),.dout(w_dff_B_QAyCvtyq7_2),.clk(gclk));
	jdff dff_B_Ob3yL81s1_2(.din(w_dff_B_QAyCvtyq7_2),.dout(w_dff_B_Ob3yL81s1_2),.clk(gclk));
	jdff dff_B_SW0GfjWC1_2(.din(w_dff_B_Ob3yL81s1_2),.dout(w_dff_B_SW0GfjWC1_2),.clk(gclk));
	jdff dff_B_pdfeUBWc5_2(.din(w_dff_B_SW0GfjWC1_2),.dout(w_dff_B_pdfeUBWc5_2),.clk(gclk));
	jdff dff_B_bzFlRNgb6_2(.din(w_dff_B_pdfeUBWc5_2),.dout(w_dff_B_bzFlRNgb6_2),.clk(gclk));
	jdff dff_B_reD8dfdd1_2(.din(w_dff_B_bzFlRNgb6_2),.dout(w_dff_B_reD8dfdd1_2),.clk(gclk));
	jdff dff_B_HlnvGXCL2_2(.din(w_dff_B_reD8dfdd1_2),.dout(w_dff_B_HlnvGXCL2_2),.clk(gclk));
	jdff dff_B_9R9D6Qrj3_2(.din(w_dff_B_HlnvGXCL2_2),.dout(w_dff_B_9R9D6Qrj3_2),.clk(gclk));
	jdff dff_B_685BWqiP9_2(.din(w_dff_B_9R9D6Qrj3_2),.dout(w_dff_B_685BWqiP9_2),.clk(gclk));
	jdff dff_B_OjdGeNKJ3_2(.din(w_dff_B_685BWqiP9_2),.dout(w_dff_B_OjdGeNKJ3_2),.clk(gclk));
	jdff dff_B_ryEQoQyp0_2(.din(w_dff_B_OjdGeNKJ3_2),.dout(w_dff_B_ryEQoQyp0_2),.clk(gclk));
	jdff dff_B_snitgZz50_2(.din(w_dff_B_ryEQoQyp0_2),.dout(w_dff_B_snitgZz50_2),.clk(gclk));
	jdff dff_B_2EI7hVaw4_2(.din(w_dff_B_snitgZz50_2),.dout(w_dff_B_2EI7hVaw4_2),.clk(gclk));
	jdff dff_B_1Huhmroh3_2(.din(w_dff_B_2EI7hVaw4_2),.dout(w_dff_B_1Huhmroh3_2),.clk(gclk));
	jdff dff_B_OnVhSGaU0_2(.din(w_dff_B_1Huhmroh3_2),.dout(w_dff_B_OnVhSGaU0_2),.clk(gclk));
	jdff dff_B_Flxa6Eko8_2(.din(n327),.dout(w_dff_B_Flxa6Eko8_2),.clk(gclk));
	jdff dff_B_6Fhf9Eju8_1(.din(n291),.dout(w_dff_B_6Fhf9Eju8_1),.clk(gclk));
	jdff dff_B_7OpAxnXt7_2(.din(n239),.dout(w_dff_B_7OpAxnXt7_2),.clk(gclk));
	jdff dff_B_j0cy7ffD7_2(.din(w_dff_B_7OpAxnXt7_2),.dout(w_dff_B_j0cy7ffD7_2),.clk(gclk));
	jdff dff_B_Peeqc6VE0_2(.din(w_dff_B_j0cy7ffD7_2),.dout(w_dff_B_Peeqc6VE0_2),.clk(gclk));
	jdff dff_B_3ekBNrqu2_2(.din(w_dff_B_Peeqc6VE0_2),.dout(w_dff_B_3ekBNrqu2_2),.clk(gclk));
	jdff dff_B_Tvh1sZvk8_2(.din(w_dff_B_3ekBNrqu2_2),.dout(w_dff_B_Tvh1sZvk8_2),.clk(gclk));
	jdff dff_B_iKrspdTh0_2(.din(w_dff_B_Tvh1sZvk8_2),.dout(w_dff_B_iKrspdTh0_2),.clk(gclk));
	jdff dff_B_NT2WauMy1_2(.din(w_dff_B_iKrspdTh0_2),.dout(w_dff_B_NT2WauMy1_2),.clk(gclk));
	jdff dff_B_OW93GX1A8_2(.din(w_dff_B_NT2WauMy1_2),.dout(w_dff_B_OW93GX1A8_2),.clk(gclk));
	jdff dff_B_wPlQyK8K5_2(.din(w_dff_B_OW93GX1A8_2),.dout(w_dff_B_wPlQyK8K5_2),.clk(gclk));
	jdff dff_B_3gwdVvUv7_2(.din(w_dff_B_wPlQyK8K5_2),.dout(w_dff_B_3gwdVvUv7_2),.clk(gclk));
	jdff dff_B_QcrKqKi74_2(.din(w_dff_B_3gwdVvUv7_2),.dout(w_dff_B_QcrKqKi74_2),.clk(gclk));
	jdff dff_B_7XhZKsfy9_2(.din(w_dff_B_QcrKqKi74_2),.dout(w_dff_B_7XhZKsfy9_2),.clk(gclk));
	jdff dff_B_7t7VuDNg2_2(.din(w_dff_B_7XhZKsfy9_2),.dout(w_dff_B_7t7VuDNg2_2),.clk(gclk));
	jdff dff_B_5WzUuFtq7_2(.din(n269),.dout(w_dff_B_5WzUuFtq7_2),.clk(gclk));
	jdff dff_B_ncfFgBcp6_1(.din(n240),.dout(w_dff_B_ncfFgBcp6_1),.clk(gclk));
	jdff dff_B_1SQv2chZ3_2(.din(n196),.dout(w_dff_B_1SQv2chZ3_2),.clk(gclk));
	jdff dff_B_kaNBOWuF6_2(.din(w_dff_B_1SQv2chZ3_2),.dout(w_dff_B_kaNBOWuF6_2),.clk(gclk));
	jdff dff_B_pMy8k2Y10_2(.din(w_dff_B_kaNBOWuF6_2),.dout(w_dff_B_pMy8k2Y10_2),.clk(gclk));
	jdff dff_B_CPnvODoO8_2(.din(w_dff_B_pMy8k2Y10_2),.dout(w_dff_B_CPnvODoO8_2),.clk(gclk));
	jdff dff_B_BsS1fQvf8_2(.din(w_dff_B_CPnvODoO8_2),.dout(w_dff_B_BsS1fQvf8_2),.clk(gclk));
	jdff dff_B_4KO8A3aG2_2(.din(w_dff_B_BsS1fQvf8_2),.dout(w_dff_B_4KO8A3aG2_2),.clk(gclk));
	jdff dff_B_WoJonN7K9_2(.din(w_dff_B_4KO8A3aG2_2),.dout(w_dff_B_WoJonN7K9_2),.clk(gclk));
	jdff dff_B_cFRAFIlK7_2(.din(w_dff_B_WoJonN7K9_2),.dout(w_dff_B_cFRAFIlK7_2),.clk(gclk));
	jdff dff_B_sE7s3cCi0_2(.din(w_dff_B_cFRAFIlK7_2),.dout(w_dff_B_sE7s3cCi0_2),.clk(gclk));
	jdff dff_B_2BHgDr6f3_2(.din(w_dff_B_sE7s3cCi0_2),.dout(w_dff_B_2BHgDr6f3_2),.clk(gclk));
	jdff dff_B_Hwp7sJGy6_2(.din(n218),.dout(w_dff_B_Hwp7sJGy6_2),.clk(gclk));
	jdff dff_B_Rn758qRw2_1(.din(n197),.dout(w_dff_B_Rn758qRw2_1),.clk(gclk));
	jdff dff_B_245dB2Vj1_2(.din(n158),.dout(w_dff_B_245dB2Vj1_2),.clk(gclk));
	jdff dff_B_GxmnUU2i9_2(.din(w_dff_B_245dB2Vj1_2),.dout(w_dff_B_GxmnUU2i9_2),.clk(gclk));
	jdff dff_B_qMjk9fbg4_2(.din(w_dff_B_GxmnUU2i9_2),.dout(w_dff_B_qMjk9fbg4_2),.clk(gclk));
	jdff dff_B_HfWphmhP3_2(.din(w_dff_B_qMjk9fbg4_2),.dout(w_dff_B_HfWphmhP3_2),.clk(gclk));
	jdff dff_B_QZE1CIaw1_2(.din(w_dff_B_HfWphmhP3_2),.dout(w_dff_B_QZE1CIaw1_2),.clk(gclk));
	jdff dff_B_ht3rygSr0_2(.din(w_dff_B_QZE1CIaw1_2),.dout(w_dff_B_ht3rygSr0_2),.clk(gclk));
	jdff dff_B_E9bULjDw7_2(.din(w_dff_B_ht3rygSr0_2),.dout(w_dff_B_E9bULjDw7_2),.clk(gclk));
	jdff dff_B_U2AtfufT8_2(.din(n175),.dout(w_dff_B_U2AtfufT8_2),.clk(gclk));
	jdff dff_B_6BySlTG00_1(.din(n161),.dout(w_dff_B_6BySlTG00_1),.clk(gclk));
	jdff dff_B_jyMdLAoA5_1(.din(w_dff_B_6BySlTG00_1),.dout(w_dff_B_jyMdLAoA5_1),.clk(gclk));
	jdff dff_B_55AhhSfT5_2(.din(n128),.dout(w_dff_B_55AhhSfT5_2),.clk(gclk));
	jdff dff_B_AR0OBn1x1_2(.din(w_dff_B_55AhhSfT5_2),.dout(w_dff_B_AR0OBn1x1_2),.clk(gclk));
	jdff dff_B_SKN6sspX6_2(.din(w_dff_B_AR0OBn1x1_2),.dout(w_dff_B_SKN6sspX6_2),.clk(gclk));
	jdff dff_B_uXlhIgzZ4_2(.din(w_dff_B_SKN6sspX6_2),.dout(w_dff_B_uXlhIgzZ4_2),.clk(gclk));
	jdff dff_A_bcg8oVQH4_1(.dout(w_n130_0[1]),.din(w_dff_A_bcg8oVQH4_1),.clk(gclk));
	jdff dff_A_1G0AuNFk3_0(.dout(w_n101_0[0]),.din(w_dff_A_1G0AuNFk3_0),.clk(gclk));
	jdff dff_A_avonoj9j1_0(.dout(w_n100_1[0]),.din(w_dff_A_avonoj9j1_0),.clk(gclk));
	jdff dff_A_ixNCcfTv9_1(.dout(w_n100_0[1]),.din(w_dff_A_ixNCcfTv9_1),.clk(gclk));
	jdff dff_A_ir0jkoTy5_2(.dout(w_n100_0[2]),.din(w_dff_A_ir0jkoTy5_2),.clk(gclk));
	jdff dff_A_srC73IwU0_2(.dout(w_dff_A_ir0jkoTy5_2),.din(w_dff_A_srC73IwU0_2),.clk(gclk));
	jdff dff_B_iWR1jGX20_0(.din(n1329),.dout(w_dff_B_iWR1jGX20_0),.clk(gclk));
	jdff dff_A_vNJLJ28L9_1(.dout(w_n1325_0[1]),.din(w_dff_A_vNJLJ28L9_1),.clk(gclk));
	jdff dff_A_nsNq7sN28_1(.dout(w_dff_A_vNJLJ28L9_1),.din(w_dff_A_nsNq7sN28_1),.clk(gclk));
	jdff dff_B_YGmA32BL2_1(.din(n1245),.dout(w_dff_B_YGmA32BL2_1),.clk(gclk));
	jdff dff_B_Xe2jUCZn7_1(.din(w_dff_B_YGmA32BL2_1),.dout(w_dff_B_Xe2jUCZn7_1),.clk(gclk));
	jdff dff_B_VrfINGLF2_2(.din(n1152),.dout(w_dff_B_VrfINGLF2_2),.clk(gclk));
	jdff dff_B_XRfA1XNS1_2(.din(w_dff_B_VrfINGLF2_2),.dout(w_dff_B_XRfA1XNS1_2),.clk(gclk));
	jdff dff_B_OcDoaZCJ1_2(.din(w_dff_B_XRfA1XNS1_2),.dout(w_dff_B_OcDoaZCJ1_2),.clk(gclk));
	jdff dff_B_TgjGHPTz1_2(.din(w_dff_B_OcDoaZCJ1_2),.dout(w_dff_B_TgjGHPTz1_2),.clk(gclk));
	jdff dff_B_uirphLHQ6_2(.din(w_dff_B_TgjGHPTz1_2),.dout(w_dff_B_uirphLHQ6_2),.clk(gclk));
	jdff dff_B_pXrGjQ6a9_2(.din(w_dff_B_uirphLHQ6_2),.dout(w_dff_B_pXrGjQ6a9_2),.clk(gclk));
	jdff dff_B_z75aXurF5_2(.din(w_dff_B_pXrGjQ6a9_2),.dout(w_dff_B_z75aXurF5_2),.clk(gclk));
	jdff dff_B_gMdAcu1U7_2(.din(w_dff_B_z75aXurF5_2),.dout(w_dff_B_gMdAcu1U7_2),.clk(gclk));
	jdff dff_B_SAinsTPC1_2(.din(w_dff_B_gMdAcu1U7_2),.dout(w_dff_B_SAinsTPC1_2),.clk(gclk));
	jdff dff_B_Vz6fifrE0_2(.din(w_dff_B_SAinsTPC1_2),.dout(w_dff_B_Vz6fifrE0_2),.clk(gclk));
	jdff dff_B_G7rr8G725_2(.din(w_dff_B_Vz6fifrE0_2),.dout(w_dff_B_G7rr8G725_2),.clk(gclk));
	jdff dff_B_I2mQM6LX9_2(.din(w_dff_B_G7rr8G725_2),.dout(w_dff_B_I2mQM6LX9_2),.clk(gclk));
	jdff dff_B_QUJcTRdT2_2(.din(w_dff_B_I2mQM6LX9_2),.dout(w_dff_B_QUJcTRdT2_2),.clk(gclk));
	jdff dff_B_2BGDN8B65_2(.din(w_dff_B_QUJcTRdT2_2),.dout(w_dff_B_2BGDN8B65_2),.clk(gclk));
	jdff dff_B_hBQWltrx1_2(.din(w_dff_B_2BGDN8B65_2),.dout(w_dff_B_hBQWltrx1_2),.clk(gclk));
	jdff dff_B_TdXrTcUA7_2(.din(w_dff_B_hBQWltrx1_2),.dout(w_dff_B_TdXrTcUA7_2),.clk(gclk));
	jdff dff_B_IpKsEiml0_2(.din(w_dff_B_TdXrTcUA7_2),.dout(w_dff_B_IpKsEiml0_2),.clk(gclk));
	jdff dff_B_VgYxqRs84_2(.din(w_dff_B_IpKsEiml0_2),.dout(w_dff_B_VgYxqRs84_2),.clk(gclk));
	jdff dff_B_Jr4pzSBm6_2(.din(w_dff_B_VgYxqRs84_2),.dout(w_dff_B_Jr4pzSBm6_2),.clk(gclk));
	jdff dff_B_9v4AewAA1_2(.din(w_dff_B_Jr4pzSBm6_2),.dout(w_dff_B_9v4AewAA1_2),.clk(gclk));
	jdff dff_B_sUyJAQLP2_2(.din(w_dff_B_9v4AewAA1_2),.dout(w_dff_B_sUyJAQLP2_2),.clk(gclk));
	jdff dff_B_iIaN59k97_2(.din(w_dff_B_sUyJAQLP2_2),.dout(w_dff_B_iIaN59k97_2),.clk(gclk));
	jdff dff_B_7STjTvPY6_2(.din(w_dff_B_iIaN59k97_2),.dout(w_dff_B_7STjTvPY6_2),.clk(gclk));
	jdff dff_B_SrNRAmR12_2(.din(w_dff_B_7STjTvPY6_2),.dout(w_dff_B_SrNRAmR12_2),.clk(gclk));
	jdff dff_B_O8jpz1An2_2(.din(w_dff_B_SrNRAmR12_2),.dout(w_dff_B_O8jpz1An2_2),.clk(gclk));
	jdff dff_B_7T1mB0cm9_2(.din(w_dff_B_O8jpz1An2_2),.dout(w_dff_B_7T1mB0cm9_2),.clk(gclk));
	jdff dff_B_DmaFqNAH0_2(.din(w_dff_B_7T1mB0cm9_2),.dout(w_dff_B_DmaFqNAH0_2),.clk(gclk));
	jdff dff_B_WobrmUQu2_2(.din(w_dff_B_DmaFqNAH0_2),.dout(w_dff_B_WobrmUQu2_2),.clk(gclk));
	jdff dff_B_D2JmnkdL1_2(.din(w_dff_B_WobrmUQu2_2),.dout(w_dff_B_D2JmnkdL1_2),.clk(gclk));
	jdff dff_B_tpgvJ9CA8_2(.din(w_dff_B_D2JmnkdL1_2),.dout(w_dff_B_tpgvJ9CA8_2),.clk(gclk));
	jdff dff_B_BSOTueR98_2(.din(w_dff_B_tpgvJ9CA8_2),.dout(w_dff_B_BSOTueR98_2),.clk(gclk));
	jdff dff_B_VQH5x6mD1_2(.din(w_dff_B_BSOTueR98_2),.dout(w_dff_B_VQH5x6mD1_2),.clk(gclk));
	jdff dff_B_EbjNuSer1_2(.din(w_dff_B_VQH5x6mD1_2),.dout(w_dff_B_EbjNuSer1_2),.clk(gclk));
	jdff dff_B_ka8jStj19_2(.din(w_dff_B_EbjNuSer1_2),.dout(w_dff_B_ka8jStj19_2),.clk(gclk));
	jdff dff_B_kNTlWiqX7_2(.din(w_dff_B_ka8jStj19_2),.dout(w_dff_B_kNTlWiqX7_2),.clk(gclk));
	jdff dff_B_afMCcITk5_2(.din(w_dff_B_kNTlWiqX7_2),.dout(w_dff_B_afMCcITk5_2),.clk(gclk));
	jdff dff_B_bpOdG4iR4_2(.din(w_dff_B_afMCcITk5_2),.dout(w_dff_B_bpOdG4iR4_2),.clk(gclk));
	jdff dff_B_EH4SD5so8_2(.din(w_dff_B_bpOdG4iR4_2),.dout(w_dff_B_EH4SD5so8_2),.clk(gclk));
	jdff dff_B_ebJun9CI7_2(.din(w_dff_B_EH4SD5so8_2),.dout(w_dff_B_ebJun9CI7_2),.clk(gclk));
	jdff dff_B_Rk1dtwek0_2(.din(w_dff_B_ebJun9CI7_2),.dout(w_dff_B_Rk1dtwek0_2),.clk(gclk));
	jdff dff_B_71HUwSnK0_2(.din(w_dff_B_Rk1dtwek0_2),.dout(w_dff_B_71HUwSnK0_2),.clk(gclk));
	jdff dff_B_dZZyLqHf4_2(.din(w_dff_B_71HUwSnK0_2),.dout(w_dff_B_dZZyLqHf4_2),.clk(gclk));
	jdff dff_B_QSRCM4is5_2(.din(w_dff_B_dZZyLqHf4_2),.dout(w_dff_B_QSRCM4is5_2),.clk(gclk));
	jdff dff_B_yiuIGVGX8_2(.din(w_dff_B_QSRCM4is5_2),.dout(w_dff_B_yiuIGVGX8_2),.clk(gclk));
	jdff dff_B_fZaMNZMF5_2(.din(w_dff_B_yiuIGVGX8_2),.dout(w_dff_B_fZaMNZMF5_2),.clk(gclk));
	jdff dff_B_la2T5edW5_2(.din(w_dff_B_fZaMNZMF5_2),.dout(w_dff_B_la2T5edW5_2),.clk(gclk));
	jdff dff_B_GIJup5jm6_2(.din(n1234),.dout(w_dff_B_GIJup5jm6_2),.clk(gclk));
	jdff dff_B_KiUGehzL6_1(.din(n1154),.dout(w_dff_B_KiUGehzL6_1),.clk(gclk));
	jdff dff_B_rewq4jsN8_2(.din(n1049),.dout(w_dff_B_rewq4jsN8_2),.clk(gclk));
	jdff dff_B_FsJAHL7T8_2(.din(w_dff_B_rewq4jsN8_2),.dout(w_dff_B_FsJAHL7T8_2),.clk(gclk));
	jdff dff_B_DxbEk9Do7_2(.din(w_dff_B_FsJAHL7T8_2),.dout(w_dff_B_DxbEk9Do7_2),.clk(gclk));
	jdff dff_B_qk9p5GUp6_2(.din(w_dff_B_DxbEk9Do7_2),.dout(w_dff_B_qk9p5GUp6_2),.clk(gclk));
	jdff dff_B_HZN6197g9_2(.din(w_dff_B_qk9p5GUp6_2),.dout(w_dff_B_HZN6197g9_2),.clk(gclk));
	jdff dff_B_ItHsGKyE2_2(.din(w_dff_B_HZN6197g9_2),.dout(w_dff_B_ItHsGKyE2_2),.clk(gclk));
	jdff dff_B_hRMkurKu0_2(.din(w_dff_B_ItHsGKyE2_2),.dout(w_dff_B_hRMkurKu0_2),.clk(gclk));
	jdff dff_B_10g616Fd4_2(.din(w_dff_B_hRMkurKu0_2),.dout(w_dff_B_10g616Fd4_2),.clk(gclk));
	jdff dff_B_AjD8ZvoK2_2(.din(w_dff_B_10g616Fd4_2),.dout(w_dff_B_AjD8ZvoK2_2),.clk(gclk));
	jdff dff_B_EsPpHUED9_2(.din(w_dff_B_AjD8ZvoK2_2),.dout(w_dff_B_EsPpHUED9_2),.clk(gclk));
	jdff dff_B_z4QvrVIP4_2(.din(w_dff_B_EsPpHUED9_2),.dout(w_dff_B_z4QvrVIP4_2),.clk(gclk));
	jdff dff_B_EdUwjeuf8_2(.din(w_dff_B_z4QvrVIP4_2),.dout(w_dff_B_EdUwjeuf8_2),.clk(gclk));
	jdff dff_B_nYnp5rFQ8_2(.din(w_dff_B_EdUwjeuf8_2),.dout(w_dff_B_nYnp5rFQ8_2),.clk(gclk));
	jdff dff_B_aRSQi7JQ7_2(.din(w_dff_B_nYnp5rFQ8_2),.dout(w_dff_B_aRSQi7JQ7_2),.clk(gclk));
	jdff dff_B_5C1Bkj3z8_2(.din(w_dff_B_aRSQi7JQ7_2),.dout(w_dff_B_5C1Bkj3z8_2),.clk(gclk));
	jdff dff_B_FNBeGY117_2(.din(w_dff_B_5C1Bkj3z8_2),.dout(w_dff_B_FNBeGY117_2),.clk(gclk));
	jdff dff_B_TQGFwaNc2_2(.din(w_dff_B_FNBeGY117_2),.dout(w_dff_B_TQGFwaNc2_2),.clk(gclk));
	jdff dff_B_nMaRYxcD2_2(.din(w_dff_B_TQGFwaNc2_2),.dout(w_dff_B_nMaRYxcD2_2),.clk(gclk));
	jdff dff_B_EqTgjE9Q8_2(.din(w_dff_B_nMaRYxcD2_2),.dout(w_dff_B_EqTgjE9Q8_2),.clk(gclk));
	jdff dff_B_wSvHJhfE2_2(.din(w_dff_B_EqTgjE9Q8_2),.dout(w_dff_B_wSvHJhfE2_2),.clk(gclk));
	jdff dff_B_Cm294iTF6_2(.din(w_dff_B_wSvHJhfE2_2),.dout(w_dff_B_Cm294iTF6_2),.clk(gclk));
	jdff dff_B_xmhdO6RH9_2(.din(w_dff_B_Cm294iTF6_2),.dout(w_dff_B_xmhdO6RH9_2),.clk(gclk));
	jdff dff_B_xtH2xk4b5_2(.din(w_dff_B_xmhdO6RH9_2),.dout(w_dff_B_xtH2xk4b5_2),.clk(gclk));
	jdff dff_B_9c9MD8zi2_2(.din(w_dff_B_xtH2xk4b5_2),.dout(w_dff_B_9c9MD8zi2_2),.clk(gclk));
	jdff dff_B_yRBYk8Oe2_2(.din(w_dff_B_9c9MD8zi2_2),.dout(w_dff_B_yRBYk8Oe2_2),.clk(gclk));
	jdff dff_B_MGHYPV087_2(.din(w_dff_B_yRBYk8Oe2_2),.dout(w_dff_B_MGHYPV087_2),.clk(gclk));
	jdff dff_B_yE4eQ1Uh3_2(.din(w_dff_B_MGHYPV087_2),.dout(w_dff_B_yE4eQ1Uh3_2),.clk(gclk));
	jdff dff_B_TqRH4DC72_2(.din(w_dff_B_yE4eQ1Uh3_2),.dout(w_dff_B_TqRH4DC72_2),.clk(gclk));
	jdff dff_B_QTy9EYpY8_2(.din(w_dff_B_TqRH4DC72_2),.dout(w_dff_B_QTy9EYpY8_2),.clk(gclk));
	jdff dff_B_LR2IAJHR2_2(.din(w_dff_B_QTy9EYpY8_2),.dout(w_dff_B_LR2IAJHR2_2),.clk(gclk));
	jdff dff_B_u2lXHmpz3_2(.din(w_dff_B_LR2IAJHR2_2),.dout(w_dff_B_u2lXHmpz3_2),.clk(gclk));
	jdff dff_B_9sNQnnWr0_2(.din(w_dff_B_u2lXHmpz3_2),.dout(w_dff_B_9sNQnnWr0_2),.clk(gclk));
	jdff dff_B_JvxBIJkd5_2(.din(w_dff_B_9sNQnnWr0_2),.dout(w_dff_B_JvxBIJkd5_2),.clk(gclk));
	jdff dff_B_bdNK3aFA1_2(.din(w_dff_B_JvxBIJkd5_2),.dout(w_dff_B_bdNK3aFA1_2),.clk(gclk));
	jdff dff_B_OXb66QLL0_2(.din(w_dff_B_bdNK3aFA1_2),.dout(w_dff_B_OXb66QLL0_2),.clk(gclk));
	jdff dff_B_ui7AadZK3_2(.din(w_dff_B_OXb66QLL0_2),.dout(w_dff_B_ui7AadZK3_2),.clk(gclk));
	jdff dff_B_acAocIjr2_2(.din(w_dff_B_ui7AadZK3_2),.dout(w_dff_B_acAocIjr2_2),.clk(gclk));
	jdff dff_B_uObjiOEf1_2(.din(w_dff_B_acAocIjr2_2),.dout(w_dff_B_uObjiOEf1_2),.clk(gclk));
	jdff dff_B_RP3MClyb5_2(.din(w_dff_B_uObjiOEf1_2),.dout(w_dff_B_RP3MClyb5_2),.clk(gclk));
	jdff dff_B_6ZcaJYfa8_2(.din(w_dff_B_RP3MClyb5_2),.dout(w_dff_B_6ZcaJYfa8_2),.clk(gclk));
	jdff dff_B_hSsYxRe46_2(.din(w_dff_B_6ZcaJYfa8_2),.dout(w_dff_B_hSsYxRe46_2),.clk(gclk));
	jdff dff_B_LLAZKhDn3_2(.din(w_dff_B_hSsYxRe46_2),.dout(w_dff_B_LLAZKhDn3_2),.clk(gclk));
	jdff dff_B_4OqqlQj08_2(.din(n1135),.dout(w_dff_B_4OqqlQj08_2),.clk(gclk));
	jdff dff_B_877gKBVH1_1(.din(n1050),.dout(w_dff_B_877gKBVH1_1),.clk(gclk));
	jdff dff_B_5jft2Vwy6_2(.din(n951),.dout(w_dff_B_5jft2Vwy6_2),.clk(gclk));
	jdff dff_B_ZN8TJwuQ8_2(.din(w_dff_B_5jft2Vwy6_2),.dout(w_dff_B_ZN8TJwuQ8_2),.clk(gclk));
	jdff dff_B_zTZjp51P1_2(.din(w_dff_B_ZN8TJwuQ8_2),.dout(w_dff_B_zTZjp51P1_2),.clk(gclk));
	jdff dff_B_hUvwZgQR1_2(.din(w_dff_B_zTZjp51P1_2),.dout(w_dff_B_hUvwZgQR1_2),.clk(gclk));
	jdff dff_B_FVNmkt943_2(.din(w_dff_B_hUvwZgQR1_2),.dout(w_dff_B_FVNmkt943_2),.clk(gclk));
	jdff dff_B_sXLylmgx7_2(.din(w_dff_B_FVNmkt943_2),.dout(w_dff_B_sXLylmgx7_2),.clk(gclk));
	jdff dff_B_WANgA7vs3_2(.din(w_dff_B_sXLylmgx7_2),.dout(w_dff_B_WANgA7vs3_2),.clk(gclk));
	jdff dff_B_fCC3zs2y6_2(.din(w_dff_B_WANgA7vs3_2),.dout(w_dff_B_fCC3zs2y6_2),.clk(gclk));
	jdff dff_B_x2qKhbFB6_2(.din(w_dff_B_fCC3zs2y6_2),.dout(w_dff_B_x2qKhbFB6_2),.clk(gclk));
	jdff dff_B_GUNSKsCY0_2(.din(w_dff_B_x2qKhbFB6_2),.dout(w_dff_B_GUNSKsCY0_2),.clk(gclk));
	jdff dff_B_iQmc28Lc0_2(.din(w_dff_B_GUNSKsCY0_2),.dout(w_dff_B_iQmc28Lc0_2),.clk(gclk));
	jdff dff_B_uY4a52hs4_2(.din(w_dff_B_iQmc28Lc0_2),.dout(w_dff_B_uY4a52hs4_2),.clk(gclk));
	jdff dff_B_3iCrlnnm9_2(.din(w_dff_B_uY4a52hs4_2),.dout(w_dff_B_3iCrlnnm9_2),.clk(gclk));
	jdff dff_B_LJLGwmyK7_2(.din(w_dff_B_3iCrlnnm9_2),.dout(w_dff_B_LJLGwmyK7_2),.clk(gclk));
	jdff dff_B_NV4ochvg1_2(.din(w_dff_B_LJLGwmyK7_2),.dout(w_dff_B_NV4ochvg1_2),.clk(gclk));
	jdff dff_B_cTAZdZuN9_2(.din(w_dff_B_NV4ochvg1_2),.dout(w_dff_B_cTAZdZuN9_2),.clk(gclk));
	jdff dff_B_PrHX0WOD4_2(.din(w_dff_B_cTAZdZuN9_2),.dout(w_dff_B_PrHX0WOD4_2),.clk(gclk));
	jdff dff_B_rxkKwHsc1_2(.din(w_dff_B_PrHX0WOD4_2),.dout(w_dff_B_rxkKwHsc1_2),.clk(gclk));
	jdff dff_B_8rmTXVCC1_2(.din(w_dff_B_rxkKwHsc1_2),.dout(w_dff_B_8rmTXVCC1_2),.clk(gclk));
	jdff dff_B_6nCHpHQ83_2(.din(w_dff_B_8rmTXVCC1_2),.dout(w_dff_B_6nCHpHQ83_2),.clk(gclk));
	jdff dff_B_v9bxAY7j3_2(.din(w_dff_B_6nCHpHQ83_2),.dout(w_dff_B_v9bxAY7j3_2),.clk(gclk));
	jdff dff_B_dkFlagy72_2(.din(w_dff_B_v9bxAY7j3_2),.dout(w_dff_B_dkFlagy72_2),.clk(gclk));
	jdff dff_B_aXPHQdB68_2(.din(w_dff_B_dkFlagy72_2),.dout(w_dff_B_aXPHQdB68_2),.clk(gclk));
	jdff dff_B_dnoxVV8M8_2(.din(w_dff_B_aXPHQdB68_2),.dout(w_dff_B_dnoxVV8M8_2),.clk(gclk));
	jdff dff_B_siVuMN1S1_2(.din(w_dff_B_dnoxVV8M8_2),.dout(w_dff_B_siVuMN1S1_2),.clk(gclk));
	jdff dff_B_OvKBIR2v5_2(.din(w_dff_B_siVuMN1S1_2),.dout(w_dff_B_OvKBIR2v5_2),.clk(gclk));
	jdff dff_B_VGwR5a5V8_2(.din(w_dff_B_OvKBIR2v5_2),.dout(w_dff_B_VGwR5a5V8_2),.clk(gclk));
	jdff dff_B_PfZATf5Z7_2(.din(w_dff_B_VGwR5a5V8_2),.dout(w_dff_B_PfZATf5Z7_2),.clk(gclk));
	jdff dff_B_JO5e3owO8_2(.din(w_dff_B_PfZATf5Z7_2),.dout(w_dff_B_JO5e3owO8_2),.clk(gclk));
	jdff dff_B_QOIGMBCv0_2(.din(w_dff_B_JO5e3owO8_2),.dout(w_dff_B_QOIGMBCv0_2),.clk(gclk));
	jdff dff_B_cOEeJdOO5_2(.din(w_dff_B_QOIGMBCv0_2),.dout(w_dff_B_cOEeJdOO5_2),.clk(gclk));
	jdff dff_B_bLVjfL3e5_2(.din(w_dff_B_cOEeJdOO5_2),.dout(w_dff_B_bLVjfL3e5_2),.clk(gclk));
	jdff dff_B_RaWgKTIy8_2(.din(w_dff_B_bLVjfL3e5_2),.dout(w_dff_B_RaWgKTIy8_2),.clk(gclk));
	jdff dff_B_l22DOOKi2_2(.din(w_dff_B_RaWgKTIy8_2),.dout(w_dff_B_l22DOOKi2_2),.clk(gclk));
	jdff dff_B_0GbXCiTa4_2(.din(w_dff_B_l22DOOKi2_2),.dout(w_dff_B_0GbXCiTa4_2),.clk(gclk));
	jdff dff_B_ET3KHaJ89_2(.din(w_dff_B_0GbXCiTa4_2),.dout(w_dff_B_ET3KHaJ89_2),.clk(gclk));
	jdff dff_B_zFBisT5P4_2(.din(w_dff_B_ET3KHaJ89_2),.dout(w_dff_B_zFBisT5P4_2),.clk(gclk));
	jdff dff_B_lwCdysTz7_2(.din(n1030),.dout(w_dff_B_lwCdysTz7_2),.clk(gclk));
	jdff dff_B_vxmO1t5E1_1(.din(n952),.dout(w_dff_B_vxmO1t5E1_1),.clk(gclk));
	jdff dff_B_KgNEIDdg7_2(.din(n846),.dout(w_dff_B_KgNEIDdg7_2),.clk(gclk));
	jdff dff_B_DyOciAqY6_2(.din(w_dff_B_KgNEIDdg7_2),.dout(w_dff_B_DyOciAqY6_2),.clk(gclk));
	jdff dff_B_AO610JJm0_2(.din(w_dff_B_DyOciAqY6_2),.dout(w_dff_B_AO610JJm0_2),.clk(gclk));
	jdff dff_B_4Bx7eUcR0_2(.din(w_dff_B_AO610JJm0_2),.dout(w_dff_B_4Bx7eUcR0_2),.clk(gclk));
	jdff dff_B_Dce8WUZR6_2(.din(w_dff_B_4Bx7eUcR0_2),.dout(w_dff_B_Dce8WUZR6_2),.clk(gclk));
	jdff dff_B_NTm7gPf28_2(.din(w_dff_B_Dce8WUZR6_2),.dout(w_dff_B_NTm7gPf28_2),.clk(gclk));
	jdff dff_B_fU6SomYh0_2(.din(w_dff_B_NTm7gPf28_2),.dout(w_dff_B_fU6SomYh0_2),.clk(gclk));
	jdff dff_B_OdaSii8Z4_2(.din(w_dff_B_fU6SomYh0_2),.dout(w_dff_B_OdaSii8Z4_2),.clk(gclk));
	jdff dff_B_1niVhtcy2_2(.din(w_dff_B_OdaSii8Z4_2),.dout(w_dff_B_1niVhtcy2_2),.clk(gclk));
	jdff dff_B_GstPYLjk1_2(.din(w_dff_B_1niVhtcy2_2),.dout(w_dff_B_GstPYLjk1_2),.clk(gclk));
	jdff dff_B_T8Spe6jd9_2(.din(w_dff_B_GstPYLjk1_2),.dout(w_dff_B_T8Spe6jd9_2),.clk(gclk));
	jdff dff_B_lPRBVp1C3_2(.din(w_dff_B_T8Spe6jd9_2),.dout(w_dff_B_lPRBVp1C3_2),.clk(gclk));
	jdff dff_B_pwA5AzaO2_2(.din(w_dff_B_lPRBVp1C3_2),.dout(w_dff_B_pwA5AzaO2_2),.clk(gclk));
	jdff dff_B_BI5zecxF9_2(.din(w_dff_B_pwA5AzaO2_2),.dout(w_dff_B_BI5zecxF9_2),.clk(gclk));
	jdff dff_B_Rf3UPpIJ2_2(.din(w_dff_B_BI5zecxF9_2),.dout(w_dff_B_Rf3UPpIJ2_2),.clk(gclk));
	jdff dff_B_NJz4azqW1_2(.din(w_dff_B_Rf3UPpIJ2_2),.dout(w_dff_B_NJz4azqW1_2),.clk(gclk));
	jdff dff_B_NfQ241217_2(.din(w_dff_B_NJz4azqW1_2),.dout(w_dff_B_NfQ241217_2),.clk(gclk));
	jdff dff_B_awfMdEK42_2(.din(w_dff_B_NfQ241217_2),.dout(w_dff_B_awfMdEK42_2),.clk(gclk));
	jdff dff_B_0PeRm2hj5_2(.din(w_dff_B_awfMdEK42_2),.dout(w_dff_B_0PeRm2hj5_2),.clk(gclk));
	jdff dff_B_Qmg3mdtc5_2(.din(w_dff_B_0PeRm2hj5_2),.dout(w_dff_B_Qmg3mdtc5_2),.clk(gclk));
	jdff dff_B_wG7tUDtG6_2(.din(w_dff_B_Qmg3mdtc5_2),.dout(w_dff_B_wG7tUDtG6_2),.clk(gclk));
	jdff dff_B_oB2hDlLM6_2(.din(w_dff_B_wG7tUDtG6_2),.dout(w_dff_B_oB2hDlLM6_2),.clk(gclk));
	jdff dff_B_P7fByLw52_2(.din(w_dff_B_oB2hDlLM6_2),.dout(w_dff_B_P7fByLw52_2),.clk(gclk));
	jdff dff_B_4lr70A8b7_2(.din(w_dff_B_P7fByLw52_2),.dout(w_dff_B_4lr70A8b7_2),.clk(gclk));
	jdff dff_B_dhwmhWxF1_2(.din(w_dff_B_4lr70A8b7_2),.dout(w_dff_B_dhwmhWxF1_2),.clk(gclk));
	jdff dff_B_jl7oPzYT6_2(.din(w_dff_B_dhwmhWxF1_2),.dout(w_dff_B_jl7oPzYT6_2),.clk(gclk));
	jdff dff_B_2extvQgJ6_2(.din(w_dff_B_jl7oPzYT6_2),.dout(w_dff_B_2extvQgJ6_2),.clk(gclk));
	jdff dff_B_AuJWx6rf1_2(.din(w_dff_B_2extvQgJ6_2),.dout(w_dff_B_AuJWx6rf1_2),.clk(gclk));
	jdff dff_B_tLaxWX5T1_2(.din(w_dff_B_AuJWx6rf1_2),.dout(w_dff_B_tLaxWX5T1_2),.clk(gclk));
	jdff dff_B_bBV8Rk6E4_2(.din(w_dff_B_tLaxWX5T1_2),.dout(w_dff_B_bBV8Rk6E4_2),.clk(gclk));
	jdff dff_B_HpW7zvZH0_2(.din(w_dff_B_bBV8Rk6E4_2),.dout(w_dff_B_HpW7zvZH0_2),.clk(gclk));
	jdff dff_B_EipvCePu1_2(.din(w_dff_B_HpW7zvZH0_2),.dout(w_dff_B_EipvCePu1_2),.clk(gclk));
	jdff dff_B_l7FlFbyc1_2(.din(w_dff_B_EipvCePu1_2),.dout(w_dff_B_l7FlFbyc1_2),.clk(gclk));
	jdff dff_B_X2kT5Udq3_2(.din(w_dff_B_l7FlFbyc1_2),.dout(w_dff_B_X2kT5Udq3_2),.clk(gclk));
	jdff dff_B_6Gtr6lbk5_2(.din(n925),.dout(w_dff_B_6Gtr6lbk5_2),.clk(gclk));
	jdff dff_B_pkXP9ILj6_1(.din(n847),.dout(w_dff_B_pkXP9ILj6_1),.clk(gclk));
	jdff dff_B_7T2LisQI8_2(.din(n747),.dout(w_dff_B_7T2LisQI8_2),.clk(gclk));
	jdff dff_B_83iD7Qxu4_2(.din(w_dff_B_7T2LisQI8_2),.dout(w_dff_B_83iD7Qxu4_2),.clk(gclk));
	jdff dff_B_4jDij4Gy4_2(.din(w_dff_B_83iD7Qxu4_2),.dout(w_dff_B_4jDij4Gy4_2),.clk(gclk));
	jdff dff_B_7JujXeVW3_2(.din(w_dff_B_4jDij4Gy4_2),.dout(w_dff_B_7JujXeVW3_2),.clk(gclk));
	jdff dff_B_Y591g1cA7_2(.din(w_dff_B_7JujXeVW3_2),.dout(w_dff_B_Y591g1cA7_2),.clk(gclk));
	jdff dff_B_OPsknhG53_2(.din(w_dff_B_Y591g1cA7_2),.dout(w_dff_B_OPsknhG53_2),.clk(gclk));
	jdff dff_B_Oet3mOMN6_2(.din(w_dff_B_OPsknhG53_2),.dout(w_dff_B_Oet3mOMN6_2),.clk(gclk));
	jdff dff_B_dzqTfCik5_2(.din(w_dff_B_Oet3mOMN6_2),.dout(w_dff_B_dzqTfCik5_2),.clk(gclk));
	jdff dff_B_5eDO5SmG6_2(.din(w_dff_B_dzqTfCik5_2),.dout(w_dff_B_5eDO5SmG6_2),.clk(gclk));
	jdff dff_B_jPoroVdG8_2(.din(w_dff_B_5eDO5SmG6_2),.dout(w_dff_B_jPoroVdG8_2),.clk(gclk));
	jdff dff_B_iIynPmaY5_2(.din(w_dff_B_jPoroVdG8_2),.dout(w_dff_B_iIynPmaY5_2),.clk(gclk));
	jdff dff_B_4aihdRmi2_2(.din(w_dff_B_iIynPmaY5_2),.dout(w_dff_B_4aihdRmi2_2),.clk(gclk));
	jdff dff_B_O3vtcIue1_2(.din(w_dff_B_4aihdRmi2_2),.dout(w_dff_B_O3vtcIue1_2),.clk(gclk));
	jdff dff_B_GinTlZ4E5_2(.din(w_dff_B_O3vtcIue1_2),.dout(w_dff_B_GinTlZ4E5_2),.clk(gclk));
	jdff dff_B_8hOLKX822_2(.din(w_dff_B_GinTlZ4E5_2),.dout(w_dff_B_8hOLKX822_2),.clk(gclk));
	jdff dff_B_D4wy2Okt0_2(.din(w_dff_B_8hOLKX822_2),.dout(w_dff_B_D4wy2Okt0_2),.clk(gclk));
	jdff dff_B_zogtRBeB2_2(.din(w_dff_B_D4wy2Okt0_2),.dout(w_dff_B_zogtRBeB2_2),.clk(gclk));
	jdff dff_B_kcYT7JJE9_2(.din(w_dff_B_zogtRBeB2_2),.dout(w_dff_B_kcYT7JJE9_2),.clk(gclk));
	jdff dff_B_h74PmwWU9_2(.din(w_dff_B_kcYT7JJE9_2),.dout(w_dff_B_h74PmwWU9_2),.clk(gclk));
	jdff dff_B_fxamom8A5_2(.din(w_dff_B_h74PmwWU9_2),.dout(w_dff_B_fxamom8A5_2),.clk(gclk));
	jdff dff_B_7plIDstX4_2(.din(w_dff_B_fxamom8A5_2),.dout(w_dff_B_7plIDstX4_2),.clk(gclk));
	jdff dff_B_zwt3KlqH6_2(.din(w_dff_B_7plIDstX4_2),.dout(w_dff_B_zwt3KlqH6_2),.clk(gclk));
	jdff dff_B_F0e8ypID5_2(.din(w_dff_B_zwt3KlqH6_2),.dout(w_dff_B_F0e8ypID5_2),.clk(gclk));
	jdff dff_B_INyCAKn87_2(.din(w_dff_B_F0e8ypID5_2),.dout(w_dff_B_INyCAKn87_2),.clk(gclk));
	jdff dff_B_bG8EAJce6_2(.din(w_dff_B_INyCAKn87_2),.dout(w_dff_B_bG8EAJce6_2),.clk(gclk));
	jdff dff_B_zqeQsN1F0_2(.din(w_dff_B_bG8EAJce6_2),.dout(w_dff_B_zqeQsN1F0_2),.clk(gclk));
	jdff dff_B_vGlcpdYO4_2(.din(w_dff_B_zqeQsN1F0_2),.dout(w_dff_B_vGlcpdYO4_2),.clk(gclk));
	jdff dff_B_EGrDx8bY8_2(.din(w_dff_B_vGlcpdYO4_2),.dout(w_dff_B_EGrDx8bY8_2),.clk(gclk));
	jdff dff_B_M3k35jO77_2(.din(w_dff_B_EGrDx8bY8_2),.dout(w_dff_B_M3k35jO77_2),.clk(gclk));
	jdff dff_B_V8sBfmYO8_2(.din(w_dff_B_M3k35jO77_2),.dout(w_dff_B_V8sBfmYO8_2),.clk(gclk));
	jdff dff_B_HMm1T04d9_2(.din(w_dff_B_V8sBfmYO8_2),.dout(w_dff_B_HMm1T04d9_2),.clk(gclk));
	jdff dff_B_pf4x7cqt6_2(.din(n819),.dout(w_dff_B_pf4x7cqt6_2),.clk(gclk));
	jdff dff_B_BJRhwV3R5_1(.din(n748),.dout(w_dff_B_BJRhwV3R5_1),.clk(gclk));
	jdff dff_B_BQnm9l3F7_2(.din(n654),.dout(w_dff_B_BQnm9l3F7_2),.clk(gclk));
	jdff dff_B_0fs6jalb2_2(.din(w_dff_B_BQnm9l3F7_2),.dout(w_dff_B_0fs6jalb2_2),.clk(gclk));
	jdff dff_B_tWegmQyn5_2(.din(w_dff_B_0fs6jalb2_2),.dout(w_dff_B_tWegmQyn5_2),.clk(gclk));
	jdff dff_B_c8BeTa936_2(.din(w_dff_B_tWegmQyn5_2),.dout(w_dff_B_c8BeTa936_2),.clk(gclk));
	jdff dff_B_UT333E6g5_2(.din(w_dff_B_c8BeTa936_2),.dout(w_dff_B_UT333E6g5_2),.clk(gclk));
	jdff dff_B_7aK2YLmc4_2(.din(w_dff_B_UT333E6g5_2),.dout(w_dff_B_7aK2YLmc4_2),.clk(gclk));
	jdff dff_B_YSRAgxvZ2_2(.din(w_dff_B_7aK2YLmc4_2),.dout(w_dff_B_YSRAgxvZ2_2),.clk(gclk));
	jdff dff_B_hZO859T94_2(.din(w_dff_B_YSRAgxvZ2_2),.dout(w_dff_B_hZO859T94_2),.clk(gclk));
	jdff dff_B_Rjud5mMf3_2(.din(w_dff_B_hZO859T94_2),.dout(w_dff_B_Rjud5mMf3_2),.clk(gclk));
	jdff dff_B_jKvJFixD2_2(.din(w_dff_B_Rjud5mMf3_2),.dout(w_dff_B_jKvJFixD2_2),.clk(gclk));
	jdff dff_B_o2SywZtH9_2(.din(w_dff_B_jKvJFixD2_2),.dout(w_dff_B_o2SywZtH9_2),.clk(gclk));
	jdff dff_B_3K0e5WII4_2(.din(w_dff_B_o2SywZtH9_2),.dout(w_dff_B_3K0e5WII4_2),.clk(gclk));
	jdff dff_B_FM3HVfhi8_2(.din(w_dff_B_3K0e5WII4_2),.dout(w_dff_B_FM3HVfhi8_2),.clk(gclk));
	jdff dff_B_zWDUI0Me3_2(.din(w_dff_B_FM3HVfhi8_2),.dout(w_dff_B_zWDUI0Me3_2),.clk(gclk));
	jdff dff_B_avZ27p1p6_2(.din(w_dff_B_zWDUI0Me3_2),.dout(w_dff_B_avZ27p1p6_2),.clk(gclk));
	jdff dff_B_NEm5x4Wc3_2(.din(w_dff_B_avZ27p1p6_2),.dout(w_dff_B_NEm5x4Wc3_2),.clk(gclk));
	jdff dff_B_C5PNdhBg2_2(.din(w_dff_B_NEm5x4Wc3_2),.dout(w_dff_B_C5PNdhBg2_2),.clk(gclk));
	jdff dff_B_VKCtOqN43_2(.din(w_dff_B_C5PNdhBg2_2),.dout(w_dff_B_VKCtOqN43_2),.clk(gclk));
	jdff dff_B_lUwmlAeX7_2(.din(w_dff_B_VKCtOqN43_2),.dout(w_dff_B_lUwmlAeX7_2),.clk(gclk));
	jdff dff_B_Fbiezlze8_2(.din(w_dff_B_lUwmlAeX7_2),.dout(w_dff_B_Fbiezlze8_2),.clk(gclk));
	jdff dff_B_nufP5pcR3_2(.din(w_dff_B_Fbiezlze8_2),.dout(w_dff_B_nufP5pcR3_2),.clk(gclk));
	jdff dff_B_uakW9DrU9_2(.din(w_dff_B_nufP5pcR3_2),.dout(w_dff_B_uakW9DrU9_2),.clk(gclk));
	jdff dff_B_p9UZvedm1_2(.din(w_dff_B_uakW9DrU9_2),.dout(w_dff_B_p9UZvedm1_2),.clk(gclk));
	jdff dff_B_eucCY8Co8_2(.din(w_dff_B_p9UZvedm1_2),.dout(w_dff_B_eucCY8Co8_2),.clk(gclk));
	jdff dff_B_HTzDBLQN1_2(.din(w_dff_B_eucCY8Co8_2),.dout(w_dff_B_HTzDBLQN1_2),.clk(gclk));
	jdff dff_B_LJb31AHq0_2(.din(w_dff_B_HTzDBLQN1_2),.dout(w_dff_B_LJb31AHq0_2),.clk(gclk));
	jdff dff_B_DzISyPcN3_2(.din(w_dff_B_LJb31AHq0_2),.dout(w_dff_B_DzISyPcN3_2),.clk(gclk));
	jdff dff_B_ovFfKiA53_2(.din(w_dff_B_DzISyPcN3_2),.dout(w_dff_B_ovFfKiA53_2),.clk(gclk));
	jdff dff_B_LjFoFNip1_2(.din(n719),.dout(w_dff_B_LjFoFNip1_2),.clk(gclk));
	jdff dff_B_yk77LfyS1_1(.din(n655),.dout(w_dff_B_yk77LfyS1_1),.clk(gclk));
	jdff dff_B_vX247xk67_2(.din(n568),.dout(w_dff_B_vX247xk67_2),.clk(gclk));
	jdff dff_B_sokSTcOG0_2(.din(w_dff_B_vX247xk67_2),.dout(w_dff_B_sokSTcOG0_2),.clk(gclk));
	jdff dff_B_Au02DbKr4_2(.din(w_dff_B_sokSTcOG0_2),.dout(w_dff_B_Au02DbKr4_2),.clk(gclk));
	jdff dff_B_xAKdDGgk1_2(.din(w_dff_B_Au02DbKr4_2),.dout(w_dff_B_xAKdDGgk1_2),.clk(gclk));
	jdff dff_B_CKOuBb2H3_2(.din(w_dff_B_xAKdDGgk1_2),.dout(w_dff_B_CKOuBb2H3_2),.clk(gclk));
	jdff dff_B_J4gbxKKz7_2(.din(w_dff_B_CKOuBb2H3_2),.dout(w_dff_B_J4gbxKKz7_2),.clk(gclk));
	jdff dff_B_HmJft7fe1_2(.din(w_dff_B_J4gbxKKz7_2),.dout(w_dff_B_HmJft7fe1_2),.clk(gclk));
	jdff dff_B_0o4AMnh69_2(.din(w_dff_B_HmJft7fe1_2),.dout(w_dff_B_0o4AMnh69_2),.clk(gclk));
	jdff dff_B_uotRdzng1_2(.din(w_dff_B_0o4AMnh69_2),.dout(w_dff_B_uotRdzng1_2),.clk(gclk));
	jdff dff_B_7k9pINyR9_2(.din(w_dff_B_uotRdzng1_2),.dout(w_dff_B_7k9pINyR9_2),.clk(gclk));
	jdff dff_B_yzGc4yFe4_2(.din(w_dff_B_7k9pINyR9_2),.dout(w_dff_B_yzGc4yFe4_2),.clk(gclk));
	jdff dff_B_nNtGhztX6_2(.din(w_dff_B_yzGc4yFe4_2),.dout(w_dff_B_nNtGhztX6_2),.clk(gclk));
	jdff dff_B_C3pVjf5o5_2(.din(w_dff_B_nNtGhztX6_2),.dout(w_dff_B_C3pVjf5o5_2),.clk(gclk));
	jdff dff_B_SiadrbWM7_2(.din(w_dff_B_C3pVjf5o5_2),.dout(w_dff_B_SiadrbWM7_2),.clk(gclk));
	jdff dff_B_VByJf3059_2(.din(w_dff_B_SiadrbWM7_2),.dout(w_dff_B_VByJf3059_2),.clk(gclk));
	jdff dff_B_yH2hGQCi7_2(.din(w_dff_B_VByJf3059_2),.dout(w_dff_B_yH2hGQCi7_2),.clk(gclk));
	jdff dff_B_PHYtLVdL3_2(.din(w_dff_B_yH2hGQCi7_2),.dout(w_dff_B_PHYtLVdL3_2),.clk(gclk));
	jdff dff_B_aWFLV4zV8_2(.din(w_dff_B_PHYtLVdL3_2),.dout(w_dff_B_aWFLV4zV8_2),.clk(gclk));
	jdff dff_B_VreCK2Zn9_2(.din(w_dff_B_aWFLV4zV8_2),.dout(w_dff_B_VreCK2Zn9_2),.clk(gclk));
	jdff dff_B_vhbocJP33_2(.din(w_dff_B_VreCK2Zn9_2),.dout(w_dff_B_vhbocJP33_2),.clk(gclk));
	jdff dff_B_b36eqfI50_2(.din(w_dff_B_vhbocJP33_2),.dout(w_dff_B_b36eqfI50_2),.clk(gclk));
	jdff dff_B_tsznxY1O7_2(.din(w_dff_B_b36eqfI50_2),.dout(w_dff_B_tsznxY1O7_2),.clk(gclk));
	jdff dff_B_cqMgiee46_2(.din(w_dff_B_tsznxY1O7_2),.dout(w_dff_B_cqMgiee46_2),.clk(gclk));
	jdff dff_B_euIm4nAl6_2(.din(w_dff_B_cqMgiee46_2),.dout(w_dff_B_euIm4nAl6_2),.clk(gclk));
	jdff dff_B_tVGUx8Nc5_2(.din(w_dff_B_euIm4nAl6_2),.dout(w_dff_B_tVGUx8Nc5_2),.clk(gclk));
	jdff dff_B_KPzLWWr84_2(.din(n626),.dout(w_dff_B_KPzLWWr84_2),.clk(gclk));
	jdff dff_B_sfAyzdid9_1(.din(n569),.dout(w_dff_B_sfAyzdid9_1),.clk(gclk));
	jdff dff_B_tBziSE9s9_2(.din(n489),.dout(w_dff_B_tBziSE9s9_2),.clk(gclk));
	jdff dff_B_E3WiGHgg3_2(.din(w_dff_B_tBziSE9s9_2),.dout(w_dff_B_E3WiGHgg3_2),.clk(gclk));
	jdff dff_B_3odx0bRh1_2(.din(w_dff_B_E3WiGHgg3_2),.dout(w_dff_B_3odx0bRh1_2),.clk(gclk));
	jdff dff_B_5xvwF1AJ0_2(.din(w_dff_B_3odx0bRh1_2),.dout(w_dff_B_5xvwF1AJ0_2),.clk(gclk));
	jdff dff_B_PXwsmNAp1_2(.din(w_dff_B_5xvwF1AJ0_2),.dout(w_dff_B_PXwsmNAp1_2),.clk(gclk));
	jdff dff_B_EPR7Gnig5_2(.din(w_dff_B_PXwsmNAp1_2),.dout(w_dff_B_EPR7Gnig5_2),.clk(gclk));
	jdff dff_B_BdDlnazm5_2(.din(w_dff_B_EPR7Gnig5_2),.dout(w_dff_B_BdDlnazm5_2),.clk(gclk));
	jdff dff_B_MNrxvM1N4_2(.din(w_dff_B_BdDlnazm5_2),.dout(w_dff_B_MNrxvM1N4_2),.clk(gclk));
	jdff dff_B_FktG2pVH6_2(.din(w_dff_B_MNrxvM1N4_2),.dout(w_dff_B_FktG2pVH6_2),.clk(gclk));
	jdff dff_B_QO1tV3ur3_2(.din(w_dff_B_FktG2pVH6_2),.dout(w_dff_B_QO1tV3ur3_2),.clk(gclk));
	jdff dff_B_cHrW7Fv70_2(.din(w_dff_B_QO1tV3ur3_2),.dout(w_dff_B_cHrW7Fv70_2),.clk(gclk));
	jdff dff_B_WpCoG4pw2_2(.din(w_dff_B_cHrW7Fv70_2),.dout(w_dff_B_WpCoG4pw2_2),.clk(gclk));
	jdff dff_B_hRKP4OTP6_2(.din(w_dff_B_WpCoG4pw2_2),.dout(w_dff_B_hRKP4OTP6_2),.clk(gclk));
	jdff dff_B_aMKpDt5s2_2(.din(w_dff_B_hRKP4OTP6_2),.dout(w_dff_B_aMKpDt5s2_2),.clk(gclk));
	jdff dff_B_SBAQuFqy8_2(.din(w_dff_B_aMKpDt5s2_2),.dout(w_dff_B_SBAQuFqy8_2),.clk(gclk));
	jdff dff_B_KfWZey4c7_2(.din(w_dff_B_SBAQuFqy8_2),.dout(w_dff_B_KfWZey4c7_2),.clk(gclk));
	jdff dff_B_1sSUDwjL5_2(.din(w_dff_B_KfWZey4c7_2),.dout(w_dff_B_1sSUDwjL5_2),.clk(gclk));
	jdff dff_B_kRM71OWs1_2(.din(w_dff_B_1sSUDwjL5_2),.dout(w_dff_B_kRM71OWs1_2),.clk(gclk));
	jdff dff_B_L7Re6p556_2(.din(w_dff_B_kRM71OWs1_2),.dout(w_dff_B_L7Re6p556_2),.clk(gclk));
	jdff dff_B_RLZ1sl8P5_2(.din(w_dff_B_L7Re6p556_2),.dout(w_dff_B_RLZ1sl8P5_2),.clk(gclk));
	jdff dff_B_j7Hhtgq99_2(.din(w_dff_B_RLZ1sl8P5_2),.dout(w_dff_B_j7Hhtgq99_2),.clk(gclk));
	jdff dff_B_fS3wTcsS6_2(.din(w_dff_B_j7Hhtgq99_2),.dout(w_dff_B_fS3wTcsS6_2),.clk(gclk));
	jdff dff_B_SXqyNsLN2_2(.din(n540),.dout(w_dff_B_SXqyNsLN2_2),.clk(gclk));
	jdff dff_B_P8KsRJix4_1(.din(n490),.dout(w_dff_B_P8KsRJix4_1),.clk(gclk));
	jdff dff_B_ivtSATeg6_2(.din(n417),.dout(w_dff_B_ivtSATeg6_2),.clk(gclk));
	jdff dff_B_bSck8pg16_2(.din(w_dff_B_ivtSATeg6_2),.dout(w_dff_B_bSck8pg16_2),.clk(gclk));
	jdff dff_B_PPlnoxLt1_2(.din(w_dff_B_bSck8pg16_2),.dout(w_dff_B_PPlnoxLt1_2),.clk(gclk));
	jdff dff_B_gVRRjAkj5_2(.din(w_dff_B_PPlnoxLt1_2),.dout(w_dff_B_gVRRjAkj5_2),.clk(gclk));
	jdff dff_B_yXvRq2zm9_2(.din(w_dff_B_gVRRjAkj5_2),.dout(w_dff_B_yXvRq2zm9_2),.clk(gclk));
	jdff dff_B_udWu3Xpw1_2(.din(w_dff_B_yXvRq2zm9_2),.dout(w_dff_B_udWu3Xpw1_2),.clk(gclk));
	jdff dff_B_HPD2iSFG7_2(.din(w_dff_B_udWu3Xpw1_2),.dout(w_dff_B_HPD2iSFG7_2),.clk(gclk));
	jdff dff_B_3wR3YO3U4_2(.din(w_dff_B_HPD2iSFG7_2),.dout(w_dff_B_3wR3YO3U4_2),.clk(gclk));
	jdff dff_B_tjZYPU2Z4_2(.din(w_dff_B_3wR3YO3U4_2),.dout(w_dff_B_tjZYPU2Z4_2),.clk(gclk));
	jdff dff_B_WQXKZcJ65_2(.din(w_dff_B_tjZYPU2Z4_2),.dout(w_dff_B_WQXKZcJ65_2),.clk(gclk));
	jdff dff_B_cbevVVP57_2(.din(w_dff_B_WQXKZcJ65_2),.dout(w_dff_B_cbevVVP57_2),.clk(gclk));
	jdff dff_B_q1NKHPOc8_2(.din(w_dff_B_cbevVVP57_2),.dout(w_dff_B_q1NKHPOc8_2),.clk(gclk));
	jdff dff_B_DAKdFrKw1_2(.din(w_dff_B_q1NKHPOc8_2),.dout(w_dff_B_DAKdFrKw1_2),.clk(gclk));
	jdff dff_B_kSqrz5ax3_2(.din(w_dff_B_DAKdFrKw1_2),.dout(w_dff_B_kSqrz5ax3_2),.clk(gclk));
	jdff dff_B_jT95uDpE4_2(.din(w_dff_B_kSqrz5ax3_2),.dout(w_dff_B_jT95uDpE4_2),.clk(gclk));
	jdff dff_B_tWTx0CE57_2(.din(w_dff_B_jT95uDpE4_2),.dout(w_dff_B_tWTx0CE57_2),.clk(gclk));
	jdff dff_B_OTXhif4F3_2(.din(w_dff_B_tWTx0CE57_2),.dout(w_dff_B_OTXhif4F3_2),.clk(gclk));
	jdff dff_B_2CSl2zK59_2(.din(w_dff_B_OTXhif4F3_2),.dout(w_dff_B_2CSl2zK59_2),.clk(gclk));
	jdff dff_B_OMGyWvRk1_2(.din(w_dff_B_2CSl2zK59_2),.dout(w_dff_B_OMGyWvRk1_2),.clk(gclk));
	jdff dff_B_oiv1Ej0a7_2(.din(n461),.dout(w_dff_B_oiv1Ej0a7_2),.clk(gclk));
	jdff dff_B_dq2zZtCe8_1(.din(n418),.dout(w_dff_B_dq2zZtCe8_1),.clk(gclk));
	jdff dff_B_xM74ADJ29_2(.din(n353),.dout(w_dff_B_xM74ADJ29_2),.clk(gclk));
	jdff dff_B_3eiP6WyV9_2(.din(w_dff_B_xM74ADJ29_2),.dout(w_dff_B_3eiP6WyV9_2),.clk(gclk));
	jdff dff_B_wwcWKxWg0_2(.din(w_dff_B_3eiP6WyV9_2),.dout(w_dff_B_wwcWKxWg0_2),.clk(gclk));
	jdff dff_B_6JXvXZL78_2(.din(w_dff_B_wwcWKxWg0_2),.dout(w_dff_B_6JXvXZL78_2),.clk(gclk));
	jdff dff_B_nhQwA36v6_2(.din(w_dff_B_6JXvXZL78_2),.dout(w_dff_B_nhQwA36v6_2),.clk(gclk));
	jdff dff_B_tKbfhqnV1_2(.din(w_dff_B_nhQwA36v6_2),.dout(w_dff_B_tKbfhqnV1_2),.clk(gclk));
	jdff dff_B_u3mx4Fm42_2(.din(w_dff_B_tKbfhqnV1_2),.dout(w_dff_B_u3mx4Fm42_2),.clk(gclk));
	jdff dff_B_AHTXeoLm0_2(.din(w_dff_B_u3mx4Fm42_2),.dout(w_dff_B_AHTXeoLm0_2),.clk(gclk));
	jdff dff_B_AC2GPz4U2_2(.din(w_dff_B_AHTXeoLm0_2),.dout(w_dff_B_AC2GPz4U2_2),.clk(gclk));
	jdff dff_B_1m42DFdN0_2(.din(w_dff_B_AC2GPz4U2_2),.dout(w_dff_B_1m42DFdN0_2),.clk(gclk));
	jdff dff_B_M8rU20jP3_2(.din(w_dff_B_1m42DFdN0_2),.dout(w_dff_B_M8rU20jP3_2),.clk(gclk));
	jdff dff_B_D2qZE4Ho3_2(.din(w_dff_B_M8rU20jP3_2),.dout(w_dff_B_D2qZE4Ho3_2),.clk(gclk));
	jdff dff_B_0hHmznac2_2(.din(w_dff_B_D2qZE4Ho3_2),.dout(w_dff_B_0hHmznac2_2),.clk(gclk));
	jdff dff_B_qIOTDY6n4_2(.din(w_dff_B_0hHmznac2_2),.dout(w_dff_B_qIOTDY6n4_2),.clk(gclk));
	jdff dff_B_EBfLEmbc8_2(.din(w_dff_B_qIOTDY6n4_2),.dout(w_dff_B_EBfLEmbc8_2),.clk(gclk));
	jdff dff_B_VzlPzLz94_2(.din(w_dff_B_EBfLEmbc8_2),.dout(w_dff_B_VzlPzLz94_2),.clk(gclk));
	jdff dff_B_eVcoFSmM5_2(.din(n389),.dout(w_dff_B_eVcoFSmM5_2),.clk(gclk));
	jdff dff_B_YZOkLI4o6_1(.din(n354),.dout(w_dff_B_YZOkLI4o6_1),.clk(gclk));
	jdff dff_B_xuWjU0ax0_2(.din(n295),.dout(w_dff_B_xuWjU0ax0_2),.clk(gclk));
	jdff dff_B_udVe7QZu4_2(.din(w_dff_B_xuWjU0ax0_2),.dout(w_dff_B_udVe7QZu4_2),.clk(gclk));
	jdff dff_B_Klc1olYN9_2(.din(w_dff_B_udVe7QZu4_2),.dout(w_dff_B_Klc1olYN9_2),.clk(gclk));
	jdff dff_B_7yt3SJo93_2(.din(w_dff_B_Klc1olYN9_2),.dout(w_dff_B_7yt3SJo93_2),.clk(gclk));
	jdff dff_B_X0RUb1Vg3_2(.din(w_dff_B_7yt3SJo93_2),.dout(w_dff_B_X0RUb1Vg3_2),.clk(gclk));
	jdff dff_B_khSBdDmA2_2(.din(w_dff_B_X0RUb1Vg3_2),.dout(w_dff_B_khSBdDmA2_2),.clk(gclk));
	jdff dff_B_gmVkOzqQ9_2(.din(w_dff_B_khSBdDmA2_2),.dout(w_dff_B_gmVkOzqQ9_2),.clk(gclk));
	jdff dff_B_PJFu1ViR8_2(.din(w_dff_B_gmVkOzqQ9_2),.dout(w_dff_B_PJFu1ViR8_2),.clk(gclk));
	jdff dff_B_HwKhKumH7_2(.din(w_dff_B_PJFu1ViR8_2),.dout(w_dff_B_HwKhKumH7_2),.clk(gclk));
	jdff dff_B_OVKJk7MB5_2(.din(w_dff_B_HwKhKumH7_2),.dout(w_dff_B_OVKJk7MB5_2),.clk(gclk));
	jdff dff_B_kFgG7cQJ0_2(.din(w_dff_B_OVKJk7MB5_2),.dout(w_dff_B_kFgG7cQJ0_2),.clk(gclk));
	jdff dff_B_CgvGs1og2_2(.din(w_dff_B_kFgG7cQJ0_2),.dout(w_dff_B_CgvGs1og2_2),.clk(gclk));
	jdff dff_B_ZT1o73KG3_2(.din(w_dff_B_CgvGs1og2_2),.dout(w_dff_B_ZT1o73KG3_2),.clk(gclk));
	jdff dff_B_Pwl0RWjL6_2(.din(n325),.dout(w_dff_B_Pwl0RWjL6_2),.clk(gclk));
	jdff dff_B_emUlAaqO8_1(.din(n296),.dout(w_dff_B_emUlAaqO8_1),.clk(gclk));
	jdff dff_B_VhQFQa4L7_2(.din(n244),.dout(w_dff_B_VhQFQa4L7_2),.clk(gclk));
	jdff dff_B_mI8afoDC6_2(.din(w_dff_B_VhQFQa4L7_2),.dout(w_dff_B_mI8afoDC6_2),.clk(gclk));
	jdff dff_B_lD2EsLUg4_2(.din(w_dff_B_mI8afoDC6_2),.dout(w_dff_B_lD2EsLUg4_2),.clk(gclk));
	jdff dff_B_hAofEnzJ7_2(.din(w_dff_B_lD2EsLUg4_2),.dout(w_dff_B_hAofEnzJ7_2),.clk(gclk));
	jdff dff_B_2jUyhUpQ3_2(.din(w_dff_B_hAofEnzJ7_2),.dout(w_dff_B_2jUyhUpQ3_2),.clk(gclk));
	jdff dff_B_mEOz2IDu0_2(.din(w_dff_B_2jUyhUpQ3_2),.dout(w_dff_B_mEOz2IDu0_2),.clk(gclk));
	jdff dff_B_21cavMbj0_2(.din(w_dff_B_mEOz2IDu0_2),.dout(w_dff_B_21cavMbj0_2),.clk(gclk));
	jdff dff_B_tOik5Oue3_2(.din(w_dff_B_21cavMbj0_2),.dout(w_dff_B_tOik5Oue3_2),.clk(gclk));
	jdff dff_B_lfRjL2Zh3_2(.din(w_dff_B_tOik5Oue3_2),.dout(w_dff_B_lfRjL2Zh3_2),.clk(gclk));
	jdff dff_B_Eevn5yIO0_2(.din(w_dff_B_lfRjL2Zh3_2),.dout(w_dff_B_Eevn5yIO0_2),.clk(gclk));
	jdff dff_B_HK1uxouA2_2(.din(n267),.dout(w_dff_B_HK1uxouA2_2),.clk(gclk));
	jdff dff_B_CzRkLVTi9_1(.din(n245),.dout(w_dff_B_CzRkLVTi9_1),.clk(gclk));
	jdff dff_B_7w8WipcE5_2(.din(n201),.dout(w_dff_B_7w8WipcE5_2),.clk(gclk));
	jdff dff_B_dyrzvjCK6_2(.din(w_dff_B_7w8WipcE5_2),.dout(w_dff_B_dyrzvjCK6_2),.clk(gclk));
	jdff dff_B_c4k9w88Y8_2(.din(w_dff_B_dyrzvjCK6_2),.dout(w_dff_B_c4k9w88Y8_2),.clk(gclk));
	jdff dff_B_KUDyAe7b5_2(.din(w_dff_B_c4k9w88Y8_2),.dout(w_dff_B_KUDyAe7b5_2),.clk(gclk));
	jdff dff_B_edYnSJi39_2(.din(w_dff_B_KUDyAe7b5_2),.dout(w_dff_B_edYnSJi39_2),.clk(gclk));
	jdff dff_B_Z1h68yYY9_2(.din(w_dff_B_edYnSJi39_2),.dout(w_dff_B_Z1h68yYY9_2),.clk(gclk));
	jdff dff_B_1YazrMbv9_2(.din(w_dff_B_Z1h68yYY9_2),.dout(w_dff_B_1YazrMbv9_2),.clk(gclk));
	jdff dff_B_eHQGTVDo8_2(.din(n216),.dout(w_dff_B_eHQGTVDo8_2),.clk(gclk));
	jdff dff_B_7gwb7JRl2_1(.din(n202),.dout(w_dff_B_7gwb7JRl2_1),.clk(gclk));
	jdff dff_B_CraBrRg64_0(.din(n173),.dout(w_dff_B_CraBrRg64_0),.clk(gclk));
	jdff dff_B_BzYavjYu2_2(.din(n165),.dout(w_dff_B_BzYavjYu2_2),.clk(gclk));
	jdff dff_B_uynEtcs31_2(.din(w_dff_B_BzYavjYu2_2),.dout(w_dff_B_uynEtcs31_2),.clk(gclk));
	jdff dff_B_VjiOsel71_2(.din(w_dff_B_uynEtcs31_2),.dout(w_dff_B_VjiOsel71_2),.clk(gclk));
	jdff dff_B_LYuZZ2cD3_2(.din(w_dff_B_VjiOsel71_2),.dout(w_dff_B_LYuZZ2cD3_2),.clk(gclk));
	jdff dff_B_owZoKCNi7_1(.din(n167),.dout(w_dff_B_owZoKCNi7_1),.clk(gclk));
	jdff dff_A_HULXV26v8_0(.dout(w_n132_0[0]),.din(w_dff_A_HULXV26v8_0),.clk(gclk));
	jdff dff_A_g6UKxOzF8_0(.dout(w_dff_A_HULXV26v8_0),.din(w_dff_A_g6UKxOzF8_0),.clk(gclk));
	jdff dff_A_5rzIXust7_1(.dout(w_n132_0[1]),.din(w_dff_A_5rzIXust7_1),.clk(gclk));
	jdff dff_B_xI4KtHss7_1(.din(n1335),.dout(w_dff_B_xI4KtHss7_1),.clk(gclk));
	jdff dff_B_UZHohOxC7_2(.din(n1248),.dout(w_dff_B_UZHohOxC7_2),.clk(gclk));
	jdff dff_B_TPMAldQH1_2(.din(w_dff_B_UZHohOxC7_2),.dout(w_dff_B_TPMAldQH1_2),.clk(gclk));
	jdff dff_B_5umnd9nw4_2(.din(w_dff_B_TPMAldQH1_2),.dout(w_dff_B_5umnd9nw4_2),.clk(gclk));
	jdff dff_B_0BLSgGkg2_2(.din(w_dff_B_5umnd9nw4_2),.dout(w_dff_B_0BLSgGkg2_2),.clk(gclk));
	jdff dff_B_OXUIaxMq9_2(.din(w_dff_B_0BLSgGkg2_2),.dout(w_dff_B_OXUIaxMq9_2),.clk(gclk));
	jdff dff_B_S9W9NEpu2_2(.din(w_dff_B_OXUIaxMq9_2),.dout(w_dff_B_S9W9NEpu2_2),.clk(gclk));
	jdff dff_B_5LMjWyT50_2(.din(w_dff_B_S9W9NEpu2_2),.dout(w_dff_B_5LMjWyT50_2),.clk(gclk));
	jdff dff_B_UEMTtNBy1_2(.din(w_dff_B_5LMjWyT50_2),.dout(w_dff_B_UEMTtNBy1_2),.clk(gclk));
	jdff dff_B_eD72nMjZ9_2(.din(w_dff_B_UEMTtNBy1_2),.dout(w_dff_B_eD72nMjZ9_2),.clk(gclk));
	jdff dff_B_oNjwemyX7_2(.din(w_dff_B_eD72nMjZ9_2),.dout(w_dff_B_oNjwemyX7_2),.clk(gclk));
	jdff dff_B_Bd2jz3141_2(.din(w_dff_B_oNjwemyX7_2),.dout(w_dff_B_Bd2jz3141_2),.clk(gclk));
	jdff dff_B_h9VDgHHg6_2(.din(w_dff_B_Bd2jz3141_2),.dout(w_dff_B_h9VDgHHg6_2),.clk(gclk));
	jdff dff_B_hunrCV1g8_2(.din(w_dff_B_h9VDgHHg6_2),.dout(w_dff_B_hunrCV1g8_2),.clk(gclk));
	jdff dff_B_Oip8vEve4_2(.din(w_dff_B_hunrCV1g8_2),.dout(w_dff_B_Oip8vEve4_2),.clk(gclk));
	jdff dff_B_CGb7fR6C3_2(.din(w_dff_B_Oip8vEve4_2),.dout(w_dff_B_CGb7fR6C3_2),.clk(gclk));
	jdff dff_B_lhU3fi1G5_2(.din(w_dff_B_CGb7fR6C3_2),.dout(w_dff_B_lhU3fi1G5_2),.clk(gclk));
	jdff dff_B_LMRqX8TV9_2(.din(w_dff_B_lhU3fi1G5_2),.dout(w_dff_B_LMRqX8TV9_2),.clk(gclk));
	jdff dff_B_gbUfhRb91_2(.din(w_dff_B_LMRqX8TV9_2),.dout(w_dff_B_gbUfhRb91_2),.clk(gclk));
	jdff dff_B_gTW28RTb5_2(.din(w_dff_B_gbUfhRb91_2),.dout(w_dff_B_gTW28RTb5_2),.clk(gclk));
	jdff dff_B_JzFV2ONK0_2(.din(w_dff_B_gTW28RTb5_2),.dout(w_dff_B_JzFV2ONK0_2),.clk(gclk));
	jdff dff_B_wZ2WsLoG4_2(.din(w_dff_B_JzFV2ONK0_2),.dout(w_dff_B_wZ2WsLoG4_2),.clk(gclk));
	jdff dff_B_32evhavQ6_2(.din(w_dff_B_wZ2WsLoG4_2),.dout(w_dff_B_32evhavQ6_2),.clk(gclk));
	jdff dff_B_zRNwHgyq7_2(.din(w_dff_B_32evhavQ6_2),.dout(w_dff_B_zRNwHgyq7_2),.clk(gclk));
	jdff dff_B_CSIE9nZD5_2(.din(w_dff_B_zRNwHgyq7_2),.dout(w_dff_B_CSIE9nZD5_2),.clk(gclk));
	jdff dff_B_Hw8v52VP5_2(.din(w_dff_B_CSIE9nZD5_2),.dout(w_dff_B_Hw8v52VP5_2),.clk(gclk));
	jdff dff_B_Z0XSY5sY1_2(.din(w_dff_B_Hw8v52VP5_2),.dout(w_dff_B_Z0XSY5sY1_2),.clk(gclk));
	jdff dff_B_hr8K6DLV8_2(.din(w_dff_B_Z0XSY5sY1_2),.dout(w_dff_B_hr8K6DLV8_2),.clk(gclk));
	jdff dff_B_CpslQAyj1_2(.din(w_dff_B_hr8K6DLV8_2),.dout(w_dff_B_CpslQAyj1_2),.clk(gclk));
	jdff dff_B_RY8Tk1dv4_2(.din(w_dff_B_CpslQAyj1_2),.dout(w_dff_B_RY8Tk1dv4_2),.clk(gclk));
	jdff dff_B_GBUU6KTQ5_2(.din(w_dff_B_RY8Tk1dv4_2),.dout(w_dff_B_GBUU6KTQ5_2),.clk(gclk));
	jdff dff_B_DjKzZ8ih2_2(.din(w_dff_B_GBUU6KTQ5_2),.dout(w_dff_B_DjKzZ8ih2_2),.clk(gclk));
	jdff dff_B_Novj0s5f8_2(.din(w_dff_B_DjKzZ8ih2_2),.dout(w_dff_B_Novj0s5f8_2),.clk(gclk));
	jdff dff_B_xk6Kvhft1_2(.din(w_dff_B_Novj0s5f8_2),.dout(w_dff_B_xk6Kvhft1_2),.clk(gclk));
	jdff dff_B_OAoSmCH78_2(.din(w_dff_B_xk6Kvhft1_2),.dout(w_dff_B_OAoSmCH78_2),.clk(gclk));
	jdff dff_B_apBZy1Lr3_2(.din(w_dff_B_OAoSmCH78_2),.dout(w_dff_B_apBZy1Lr3_2),.clk(gclk));
	jdff dff_B_6vvQA9U62_2(.din(w_dff_B_apBZy1Lr3_2),.dout(w_dff_B_6vvQA9U62_2),.clk(gclk));
	jdff dff_B_MZft0Rpa3_2(.din(w_dff_B_6vvQA9U62_2),.dout(w_dff_B_MZft0Rpa3_2),.clk(gclk));
	jdff dff_B_Mlm0szhn8_2(.din(w_dff_B_MZft0Rpa3_2),.dout(w_dff_B_Mlm0szhn8_2),.clk(gclk));
	jdff dff_B_WmvtQHks0_2(.din(w_dff_B_Mlm0szhn8_2),.dout(w_dff_B_WmvtQHks0_2),.clk(gclk));
	jdff dff_B_Hyy1Rhgv9_2(.din(w_dff_B_WmvtQHks0_2),.dout(w_dff_B_Hyy1Rhgv9_2),.clk(gclk));
	jdff dff_B_vRqrLQ890_2(.din(w_dff_B_Hyy1Rhgv9_2),.dout(w_dff_B_vRqrLQ890_2),.clk(gclk));
	jdff dff_B_4nmjdSV93_2(.din(w_dff_B_vRqrLQ890_2),.dout(w_dff_B_4nmjdSV93_2),.clk(gclk));
	jdff dff_B_GfL5xMsK7_2(.din(w_dff_B_4nmjdSV93_2),.dout(w_dff_B_GfL5xMsK7_2),.clk(gclk));
	jdff dff_B_ZCZqkJND0_2(.din(w_dff_B_GfL5xMsK7_2),.dout(w_dff_B_ZCZqkJND0_2),.clk(gclk));
	jdff dff_B_aULq1Jt46_2(.din(w_dff_B_ZCZqkJND0_2),.dout(w_dff_B_aULq1Jt46_2),.clk(gclk));
	jdff dff_B_RhxBNb8P7_0(.din(n1334),.dout(w_dff_B_RhxBNb8P7_0),.clk(gclk));
	jdff dff_A_LfO3RIHK7_1(.dout(w_n1322_0[1]),.din(w_dff_A_LfO3RIHK7_1),.clk(gclk));
	jdff dff_B_JQvbpp403_1(.din(n1249),.dout(w_dff_B_JQvbpp403_1),.clk(gclk));
	jdff dff_B_U90uMvAa1_2(.din(n1158),.dout(w_dff_B_U90uMvAa1_2),.clk(gclk));
	jdff dff_B_NoiBQRiJ2_2(.din(w_dff_B_U90uMvAa1_2),.dout(w_dff_B_NoiBQRiJ2_2),.clk(gclk));
	jdff dff_B_tL1mZXxV9_2(.din(w_dff_B_NoiBQRiJ2_2),.dout(w_dff_B_tL1mZXxV9_2),.clk(gclk));
	jdff dff_B_enHzjiiw8_2(.din(w_dff_B_tL1mZXxV9_2),.dout(w_dff_B_enHzjiiw8_2),.clk(gclk));
	jdff dff_B_rZPNWW4h8_2(.din(w_dff_B_enHzjiiw8_2),.dout(w_dff_B_rZPNWW4h8_2),.clk(gclk));
	jdff dff_B_5d4oZ88T3_2(.din(w_dff_B_rZPNWW4h8_2),.dout(w_dff_B_5d4oZ88T3_2),.clk(gclk));
	jdff dff_B_LF8NBnL16_2(.din(w_dff_B_5d4oZ88T3_2),.dout(w_dff_B_LF8NBnL16_2),.clk(gclk));
	jdff dff_B_aZ6ugA3w1_2(.din(w_dff_B_LF8NBnL16_2),.dout(w_dff_B_aZ6ugA3w1_2),.clk(gclk));
	jdff dff_B_6tSuWOSC7_2(.din(w_dff_B_aZ6ugA3w1_2),.dout(w_dff_B_6tSuWOSC7_2),.clk(gclk));
	jdff dff_B_7VPh3tWa7_2(.din(w_dff_B_6tSuWOSC7_2),.dout(w_dff_B_7VPh3tWa7_2),.clk(gclk));
	jdff dff_B_IYxYnHIB6_2(.din(w_dff_B_7VPh3tWa7_2),.dout(w_dff_B_IYxYnHIB6_2),.clk(gclk));
	jdff dff_B_ZfUC2LkC6_2(.din(w_dff_B_IYxYnHIB6_2),.dout(w_dff_B_ZfUC2LkC6_2),.clk(gclk));
	jdff dff_B_bJUgQ1XH8_2(.din(w_dff_B_ZfUC2LkC6_2),.dout(w_dff_B_bJUgQ1XH8_2),.clk(gclk));
	jdff dff_B_1nfqEaHb5_2(.din(w_dff_B_bJUgQ1XH8_2),.dout(w_dff_B_1nfqEaHb5_2),.clk(gclk));
	jdff dff_B_HHn9aFlQ1_2(.din(w_dff_B_1nfqEaHb5_2),.dout(w_dff_B_HHn9aFlQ1_2),.clk(gclk));
	jdff dff_B_GGXcCVo58_2(.din(w_dff_B_HHn9aFlQ1_2),.dout(w_dff_B_GGXcCVo58_2),.clk(gclk));
	jdff dff_B_Uuexpj197_2(.din(w_dff_B_GGXcCVo58_2),.dout(w_dff_B_Uuexpj197_2),.clk(gclk));
	jdff dff_B_qmZSuspL3_2(.din(w_dff_B_Uuexpj197_2),.dout(w_dff_B_qmZSuspL3_2),.clk(gclk));
	jdff dff_B_ujEsUb5c8_2(.din(w_dff_B_qmZSuspL3_2),.dout(w_dff_B_ujEsUb5c8_2),.clk(gclk));
	jdff dff_B_WaY0OldU3_2(.din(w_dff_B_ujEsUb5c8_2),.dout(w_dff_B_WaY0OldU3_2),.clk(gclk));
	jdff dff_B_8gIcdXQJ8_2(.din(w_dff_B_WaY0OldU3_2),.dout(w_dff_B_8gIcdXQJ8_2),.clk(gclk));
	jdff dff_B_XAq5HCEW5_2(.din(w_dff_B_8gIcdXQJ8_2),.dout(w_dff_B_XAq5HCEW5_2),.clk(gclk));
	jdff dff_B_b152A6lN0_2(.din(w_dff_B_XAq5HCEW5_2),.dout(w_dff_B_b152A6lN0_2),.clk(gclk));
	jdff dff_B_k5sYsebK4_2(.din(w_dff_B_b152A6lN0_2),.dout(w_dff_B_k5sYsebK4_2),.clk(gclk));
	jdff dff_B_p5e0Aezl2_2(.din(w_dff_B_k5sYsebK4_2),.dout(w_dff_B_p5e0Aezl2_2),.clk(gclk));
	jdff dff_B_mIXScm0Q0_2(.din(w_dff_B_p5e0Aezl2_2),.dout(w_dff_B_mIXScm0Q0_2),.clk(gclk));
	jdff dff_B_pkiogah55_2(.din(w_dff_B_mIXScm0Q0_2),.dout(w_dff_B_pkiogah55_2),.clk(gclk));
	jdff dff_B_y6dWHmgG4_2(.din(w_dff_B_pkiogah55_2),.dout(w_dff_B_y6dWHmgG4_2),.clk(gclk));
	jdff dff_B_m9hCgzYF4_2(.din(w_dff_B_y6dWHmgG4_2),.dout(w_dff_B_m9hCgzYF4_2),.clk(gclk));
	jdff dff_B_QPQHOcDJ8_2(.din(w_dff_B_m9hCgzYF4_2),.dout(w_dff_B_QPQHOcDJ8_2),.clk(gclk));
	jdff dff_B_Dm8NMg9V0_2(.din(w_dff_B_QPQHOcDJ8_2),.dout(w_dff_B_Dm8NMg9V0_2),.clk(gclk));
	jdff dff_B_5NYVmpA13_2(.din(w_dff_B_Dm8NMg9V0_2),.dout(w_dff_B_5NYVmpA13_2),.clk(gclk));
	jdff dff_B_QteqSDU96_2(.din(w_dff_B_5NYVmpA13_2),.dout(w_dff_B_QteqSDU96_2),.clk(gclk));
	jdff dff_B_t2oKy07e8_2(.din(w_dff_B_QteqSDU96_2),.dout(w_dff_B_t2oKy07e8_2),.clk(gclk));
	jdff dff_B_2a6sqRoH9_2(.din(w_dff_B_t2oKy07e8_2),.dout(w_dff_B_2a6sqRoH9_2),.clk(gclk));
	jdff dff_B_AFtX9sIe1_2(.din(w_dff_B_2a6sqRoH9_2),.dout(w_dff_B_AFtX9sIe1_2),.clk(gclk));
	jdff dff_B_mv30Dwhi6_2(.din(w_dff_B_AFtX9sIe1_2),.dout(w_dff_B_mv30Dwhi6_2),.clk(gclk));
	jdff dff_B_YQa0O84W7_2(.din(w_dff_B_mv30Dwhi6_2),.dout(w_dff_B_YQa0O84W7_2),.clk(gclk));
	jdff dff_B_Ot77QrI62_2(.din(w_dff_B_YQa0O84W7_2),.dout(w_dff_B_Ot77QrI62_2),.clk(gclk));
	jdff dff_B_Iuv5wbIc7_2(.din(w_dff_B_Ot77QrI62_2),.dout(w_dff_B_Iuv5wbIc7_2),.clk(gclk));
	jdff dff_B_O1NHPjoB7_2(.din(n1231),.dout(w_dff_B_O1NHPjoB7_2),.clk(gclk));
	jdff dff_B_lOSBJ7tE3_1(.din(n1159),.dout(w_dff_B_lOSBJ7tE3_1),.clk(gclk));
	jdff dff_B_9RJNcfrF2_2(.din(n1054),.dout(w_dff_B_9RJNcfrF2_2),.clk(gclk));
	jdff dff_B_aEoizBxe3_2(.din(w_dff_B_9RJNcfrF2_2),.dout(w_dff_B_aEoizBxe3_2),.clk(gclk));
	jdff dff_B_HUhjX3n13_2(.din(w_dff_B_aEoizBxe3_2),.dout(w_dff_B_HUhjX3n13_2),.clk(gclk));
	jdff dff_B_FAnE5Wis5_2(.din(w_dff_B_HUhjX3n13_2),.dout(w_dff_B_FAnE5Wis5_2),.clk(gclk));
	jdff dff_B_inS0zxTF9_2(.din(w_dff_B_FAnE5Wis5_2),.dout(w_dff_B_inS0zxTF9_2),.clk(gclk));
	jdff dff_B_ocxw3Y8Y4_2(.din(w_dff_B_inS0zxTF9_2),.dout(w_dff_B_ocxw3Y8Y4_2),.clk(gclk));
	jdff dff_B_jKQ9Slxc5_2(.din(w_dff_B_ocxw3Y8Y4_2),.dout(w_dff_B_jKQ9Slxc5_2),.clk(gclk));
	jdff dff_B_K6n4O5zN0_2(.din(w_dff_B_jKQ9Slxc5_2),.dout(w_dff_B_K6n4O5zN0_2),.clk(gclk));
	jdff dff_B_qOSioDeL5_2(.din(w_dff_B_K6n4O5zN0_2),.dout(w_dff_B_qOSioDeL5_2),.clk(gclk));
	jdff dff_B_sqONaICq0_2(.din(w_dff_B_qOSioDeL5_2),.dout(w_dff_B_sqONaICq0_2),.clk(gclk));
	jdff dff_B_Sn6e1hcZ3_2(.din(w_dff_B_sqONaICq0_2),.dout(w_dff_B_Sn6e1hcZ3_2),.clk(gclk));
	jdff dff_B_SeW8fSQC5_2(.din(w_dff_B_Sn6e1hcZ3_2),.dout(w_dff_B_SeW8fSQC5_2),.clk(gclk));
	jdff dff_B_HBLe2pbK5_2(.din(w_dff_B_SeW8fSQC5_2),.dout(w_dff_B_HBLe2pbK5_2),.clk(gclk));
	jdff dff_B_LW4q84Ob7_2(.din(w_dff_B_HBLe2pbK5_2),.dout(w_dff_B_LW4q84Ob7_2),.clk(gclk));
	jdff dff_B_SZByWkeP9_2(.din(w_dff_B_LW4q84Ob7_2),.dout(w_dff_B_SZByWkeP9_2),.clk(gclk));
	jdff dff_B_efFwplAt5_2(.din(w_dff_B_SZByWkeP9_2),.dout(w_dff_B_efFwplAt5_2),.clk(gclk));
	jdff dff_B_b34dtNXc7_2(.din(w_dff_B_efFwplAt5_2),.dout(w_dff_B_b34dtNXc7_2),.clk(gclk));
	jdff dff_B_hUPtkb717_2(.din(w_dff_B_b34dtNXc7_2),.dout(w_dff_B_hUPtkb717_2),.clk(gclk));
	jdff dff_B_iagk97iy3_2(.din(w_dff_B_hUPtkb717_2),.dout(w_dff_B_iagk97iy3_2),.clk(gclk));
	jdff dff_B_eEyigFEQ2_2(.din(w_dff_B_iagk97iy3_2),.dout(w_dff_B_eEyigFEQ2_2),.clk(gclk));
	jdff dff_B_Y2XLB0bw4_2(.din(w_dff_B_eEyigFEQ2_2),.dout(w_dff_B_Y2XLB0bw4_2),.clk(gclk));
	jdff dff_B_upcuLzjl5_2(.din(w_dff_B_Y2XLB0bw4_2),.dout(w_dff_B_upcuLzjl5_2),.clk(gclk));
	jdff dff_B_Es71zjQl3_2(.din(w_dff_B_upcuLzjl5_2),.dout(w_dff_B_Es71zjQl3_2),.clk(gclk));
	jdff dff_B_CDVgHeAy7_2(.din(w_dff_B_Es71zjQl3_2),.dout(w_dff_B_CDVgHeAy7_2),.clk(gclk));
	jdff dff_B_duaNfMR90_2(.din(w_dff_B_CDVgHeAy7_2),.dout(w_dff_B_duaNfMR90_2),.clk(gclk));
	jdff dff_B_PK063A7o8_2(.din(w_dff_B_duaNfMR90_2),.dout(w_dff_B_PK063A7o8_2),.clk(gclk));
	jdff dff_B_cavtLJ0J7_2(.din(w_dff_B_PK063A7o8_2),.dout(w_dff_B_cavtLJ0J7_2),.clk(gclk));
	jdff dff_B_Ta4lBXkR2_2(.din(w_dff_B_cavtLJ0J7_2),.dout(w_dff_B_Ta4lBXkR2_2),.clk(gclk));
	jdff dff_B_nys8lKOj7_2(.din(w_dff_B_Ta4lBXkR2_2),.dout(w_dff_B_nys8lKOj7_2),.clk(gclk));
	jdff dff_B_K8vOuI1A7_2(.din(w_dff_B_nys8lKOj7_2),.dout(w_dff_B_K8vOuI1A7_2),.clk(gclk));
	jdff dff_B_kcgKCWXT9_2(.din(w_dff_B_K8vOuI1A7_2),.dout(w_dff_B_kcgKCWXT9_2),.clk(gclk));
	jdff dff_B_w3iLftcQ4_2(.din(w_dff_B_kcgKCWXT9_2),.dout(w_dff_B_w3iLftcQ4_2),.clk(gclk));
	jdff dff_B_wyRUFoPh9_2(.din(w_dff_B_w3iLftcQ4_2),.dout(w_dff_B_wyRUFoPh9_2),.clk(gclk));
	jdff dff_B_XNdGnwWX0_2(.din(w_dff_B_wyRUFoPh9_2),.dout(w_dff_B_XNdGnwWX0_2),.clk(gclk));
	jdff dff_B_skBhd1sh3_2(.din(w_dff_B_XNdGnwWX0_2),.dout(w_dff_B_skBhd1sh3_2),.clk(gclk));
	jdff dff_B_3azMdPCw2_2(.din(w_dff_B_skBhd1sh3_2),.dout(w_dff_B_3azMdPCw2_2),.clk(gclk));
	jdff dff_B_SzYlsXIl7_2(.din(w_dff_B_3azMdPCw2_2),.dout(w_dff_B_SzYlsXIl7_2),.clk(gclk));
	jdff dff_B_dQDJWevx9_2(.din(n1133),.dout(w_dff_B_dQDJWevx9_2),.clk(gclk));
	jdff dff_B_eCtGb53e0_1(.din(n1055),.dout(w_dff_B_eCtGb53e0_1),.clk(gclk));
	jdff dff_B_TJ0XPJ058_2(.din(n956),.dout(w_dff_B_TJ0XPJ058_2),.clk(gclk));
	jdff dff_B_LFISirk68_2(.din(w_dff_B_TJ0XPJ058_2),.dout(w_dff_B_LFISirk68_2),.clk(gclk));
	jdff dff_B_jKk0oP377_2(.din(w_dff_B_LFISirk68_2),.dout(w_dff_B_jKk0oP377_2),.clk(gclk));
	jdff dff_B_42TnxQTR1_2(.din(w_dff_B_jKk0oP377_2),.dout(w_dff_B_42TnxQTR1_2),.clk(gclk));
	jdff dff_B_eBVbqtvU6_2(.din(w_dff_B_42TnxQTR1_2),.dout(w_dff_B_eBVbqtvU6_2),.clk(gclk));
	jdff dff_B_fmejP46P8_2(.din(w_dff_B_eBVbqtvU6_2),.dout(w_dff_B_fmejP46P8_2),.clk(gclk));
	jdff dff_B_P5Q0hKUW1_2(.din(w_dff_B_fmejP46P8_2),.dout(w_dff_B_P5Q0hKUW1_2),.clk(gclk));
	jdff dff_B_tFj8JxWy3_2(.din(w_dff_B_P5Q0hKUW1_2),.dout(w_dff_B_tFj8JxWy3_2),.clk(gclk));
	jdff dff_B_8kmoOYdH1_2(.din(w_dff_B_tFj8JxWy3_2),.dout(w_dff_B_8kmoOYdH1_2),.clk(gclk));
	jdff dff_B_xpmmf9ZZ5_2(.din(w_dff_B_8kmoOYdH1_2),.dout(w_dff_B_xpmmf9ZZ5_2),.clk(gclk));
	jdff dff_B_vVzBuWer4_2(.din(w_dff_B_xpmmf9ZZ5_2),.dout(w_dff_B_vVzBuWer4_2),.clk(gclk));
	jdff dff_B_ia0jNExX5_2(.din(w_dff_B_vVzBuWer4_2),.dout(w_dff_B_ia0jNExX5_2),.clk(gclk));
	jdff dff_B_OxSmDrYf1_2(.din(w_dff_B_ia0jNExX5_2),.dout(w_dff_B_OxSmDrYf1_2),.clk(gclk));
	jdff dff_B_yjNFD4bk2_2(.din(w_dff_B_OxSmDrYf1_2),.dout(w_dff_B_yjNFD4bk2_2),.clk(gclk));
	jdff dff_B_iN8QNmSG1_2(.din(w_dff_B_yjNFD4bk2_2),.dout(w_dff_B_iN8QNmSG1_2),.clk(gclk));
	jdff dff_B_DuOCbTw32_2(.din(w_dff_B_iN8QNmSG1_2),.dout(w_dff_B_DuOCbTw32_2),.clk(gclk));
	jdff dff_B_v2omJpgm9_2(.din(w_dff_B_DuOCbTw32_2),.dout(w_dff_B_v2omJpgm9_2),.clk(gclk));
	jdff dff_B_9sJXtV8b3_2(.din(w_dff_B_v2omJpgm9_2),.dout(w_dff_B_9sJXtV8b3_2),.clk(gclk));
	jdff dff_B_HyIdw98L7_2(.din(w_dff_B_9sJXtV8b3_2),.dout(w_dff_B_HyIdw98L7_2),.clk(gclk));
	jdff dff_B_EmupylG62_2(.din(w_dff_B_HyIdw98L7_2),.dout(w_dff_B_EmupylG62_2),.clk(gclk));
	jdff dff_B_QFbOzZc40_2(.din(w_dff_B_EmupylG62_2),.dout(w_dff_B_QFbOzZc40_2),.clk(gclk));
	jdff dff_B_ECWOHVdg0_2(.din(w_dff_B_QFbOzZc40_2),.dout(w_dff_B_ECWOHVdg0_2),.clk(gclk));
	jdff dff_B_Rw1BSHKQ9_2(.din(w_dff_B_ECWOHVdg0_2),.dout(w_dff_B_Rw1BSHKQ9_2),.clk(gclk));
	jdff dff_B_O5WmV9b73_2(.din(w_dff_B_Rw1BSHKQ9_2),.dout(w_dff_B_O5WmV9b73_2),.clk(gclk));
	jdff dff_B_GxUPNd4x8_2(.din(w_dff_B_O5WmV9b73_2),.dout(w_dff_B_GxUPNd4x8_2),.clk(gclk));
	jdff dff_B_vtbgzxZ13_2(.din(w_dff_B_GxUPNd4x8_2),.dout(w_dff_B_vtbgzxZ13_2),.clk(gclk));
	jdff dff_B_zpW5bKD34_2(.din(w_dff_B_vtbgzxZ13_2),.dout(w_dff_B_zpW5bKD34_2),.clk(gclk));
	jdff dff_B_IJr7b9Kn5_2(.din(w_dff_B_zpW5bKD34_2),.dout(w_dff_B_IJr7b9Kn5_2),.clk(gclk));
	jdff dff_B_jpvW04FO2_2(.din(w_dff_B_IJr7b9Kn5_2),.dout(w_dff_B_jpvW04FO2_2),.clk(gclk));
	jdff dff_B_zcdynVVv1_2(.din(w_dff_B_jpvW04FO2_2),.dout(w_dff_B_zcdynVVv1_2),.clk(gclk));
	jdff dff_B_SOxiC8ch5_2(.din(w_dff_B_zcdynVVv1_2),.dout(w_dff_B_SOxiC8ch5_2),.clk(gclk));
	jdff dff_B_yfTvDbjC5_2(.din(w_dff_B_SOxiC8ch5_2),.dout(w_dff_B_yfTvDbjC5_2),.clk(gclk));
	jdff dff_B_r9psN4dq6_2(.din(w_dff_B_yfTvDbjC5_2),.dout(w_dff_B_r9psN4dq6_2),.clk(gclk));
	jdff dff_B_vZdHmVoe7_2(.din(w_dff_B_r9psN4dq6_2),.dout(w_dff_B_vZdHmVoe7_2),.clk(gclk));
	jdff dff_B_pV0mhRZL3_2(.din(n1028),.dout(w_dff_B_pV0mhRZL3_2),.clk(gclk));
	jdff dff_B_Rb5srVo57_1(.din(n957),.dout(w_dff_B_Rb5srVo57_1),.clk(gclk));
	jdff dff_B_lZn9UF0Q4_2(.din(n851),.dout(w_dff_B_lZn9UF0Q4_2),.clk(gclk));
	jdff dff_B_15z3pBvV7_2(.din(w_dff_B_lZn9UF0Q4_2),.dout(w_dff_B_15z3pBvV7_2),.clk(gclk));
	jdff dff_B_v8TT3key1_2(.din(w_dff_B_15z3pBvV7_2),.dout(w_dff_B_v8TT3key1_2),.clk(gclk));
	jdff dff_B_3WxeF3as2_2(.din(w_dff_B_v8TT3key1_2),.dout(w_dff_B_3WxeF3as2_2),.clk(gclk));
	jdff dff_B_cW4lRg5Y5_2(.din(w_dff_B_3WxeF3as2_2),.dout(w_dff_B_cW4lRg5Y5_2),.clk(gclk));
	jdff dff_B_on5C6lik6_2(.din(w_dff_B_cW4lRg5Y5_2),.dout(w_dff_B_on5C6lik6_2),.clk(gclk));
	jdff dff_B_poWIt2H63_2(.din(w_dff_B_on5C6lik6_2),.dout(w_dff_B_poWIt2H63_2),.clk(gclk));
	jdff dff_B_keKaoNRj2_2(.din(w_dff_B_poWIt2H63_2),.dout(w_dff_B_keKaoNRj2_2),.clk(gclk));
	jdff dff_B_YPAGzvB34_2(.din(w_dff_B_keKaoNRj2_2),.dout(w_dff_B_YPAGzvB34_2),.clk(gclk));
	jdff dff_B_sKfDDsa15_2(.din(w_dff_B_YPAGzvB34_2),.dout(w_dff_B_sKfDDsa15_2),.clk(gclk));
	jdff dff_B_145WmUMG5_2(.din(w_dff_B_sKfDDsa15_2),.dout(w_dff_B_145WmUMG5_2),.clk(gclk));
	jdff dff_B_IDhYC0Mq0_2(.din(w_dff_B_145WmUMG5_2),.dout(w_dff_B_IDhYC0Mq0_2),.clk(gclk));
	jdff dff_B_ltG2fnaH3_2(.din(w_dff_B_IDhYC0Mq0_2),.dout(w_dff_B_ltG2fnaH3_2),.clk(gclk));
	jdff dff_B_fcwqtJuG0_2(.din(w_dff_B_ltG2fnaH3_2),.dout(w_dff_B_fcwqtJuG0_2),.clk(gclk));
	jdff dff_B_3iixEj0N7_2(.din(w_dff_B_fcwqtJuG0_2),.dout(w_dff_B_3iixEj0N7_2),.clk(gclk));
	jdff dff_B_WrM8pzZb8_2(.din(w_dff_B_3iixEj0N7_2),.dout(w_dff_B_WrM8pzZb8_2),.clk(gclk));
	jdff dff_B_4tTfQJlb0_2(.din(w_dff_B_WrM8pzZb8_2),.dout(w_dff_B_4tTfQJlb0_2),.clk(gclk));
	jdff dff_B_olsGP0uP6_2(.din(w_dff_B_4tTfQJlb0_2),.dout(w_dff_B_olsGP0uP6_2),.clk(gclk));
	jdff dff_B_HoZJEgBU2_2(.din(w_dff_B_olsGP0uP6_2),.dout(w_dff_B_HoZJEgBU2_2),.clk(gclk));
	jdff dff_B_26PZ9btN9_2(.din(w_dff_B_HoZJEgBU2_2),.dout(w_dff_B_26PZ9btN9_2),.clk(gclk));
	jdff dff_B_wn9pbkMV8_2(.din(w_dff_B_26PZ9btN9_2),.dout(w_dff_B_wn9pbkMV8_2),.clk(gclk));
	jdff dff_B_IKMYJJjS8_2(.din(w_dff_B_wn9pbkMV8_2),.dout(w_dff_B_IKMYJJjS8_2),.clk(gclk));
	jdff dff_B_0d4yX2xg0_2(.din(w_dff_B_IKMYJJjS8_2),.dout(w_dff_B_0d4yX2xg0_2),.clk(gclk));
	jdff dff_B_3XdOFMFu8_2(.din(w_dff_B_0d4yX2xg0_2),.dout(w_dff_B_3XdOFMFu8_2),.clk(gclk));
	jdff dff_B_WPiWKbN28_2(.din(w_dff_B_3XdOFMFu8_2),.dout(w_dff_B_WPiWKbN28_2),.clk(gclk));
	jdff dff_B_3L6vqFYl4_2(.din(w_dff_B_WPiWKbN28_2),.dout(w_dff_B_3L6vqFYl4_2),.clk(gclk));
	jdff dff_B_OtpxpA1G4_2(.din(w_dff_B_3L6vqFYl4_2),.dout(w_dff_B_OtpxpA1G4_2),.clk(gclk));
	jdff dff_B_5o0b8ZpA8_2(.din(w_dff_B_OtpxpA1G4_2),.dout(w_dff_B_5o0b8ZpA8_2),.clk(gclk));
	jdff dff_B_pyChaReD3_2(.din(w_dff_B_5o0b8ZpA8_2),.dout(w_dff_B_pyChaReD3_2),.clk(gclk));
	jdff dff_B_djIcuisx9_2(.din(w_dff_B_pyChaReD3_2),.dout(w_dff_B_djIcuisx9_2),.clk(gclk));
	jdff dff_B_E2Lm7Htj4_2(.din(w_dff_B_djIcuisx9_2),.dout(w_dff_B_E2Lm7Htj4_2),.clk(gclk));
	jdff dff_B_eZBfBava6_2(.din(n923),.dout(w_dff_B_eZBfBava6_2),.clk(gclk));
	jdff dff_B_fWUgkO5b0_1(.din(n852),.dout(w_dff_B_fWUgkO5b0_1),.clk(gclk));
	jdff dff_B_6iUBDZHj4_2(.din(n752),.dout(w_dff_B_6iUBDZHj4_2),.clk(gclk));
	jdff dff_B_Fd0MyKka5_2(.din(w_dff_B_6iUBDZHj4_2),.dout(w_dff_B_Fd0MyKka5_2),.clk(gclk));
	jdff dff_B_ND8OBbwC0_2(.din(w_dff_B_Fd0MyKka5_2),.dout(w_dff_B_ND8OBbwC0_2),.clk(gclk));
	jdff dff_B_nErpmHl18_2(.din(w_dff_B_ND8OBbwC0_2),.dout(w_dff_B_nErpmHl18_2),.clk(gclk));
	jdff dff_B_2tEclMAK1_2(.din(w_dff_B_nErpmHl18_2),.dout(w_dff_B_2tEclMAK1_2),.clk(gclk));
	jdff dff_B_lA9v8wsM5_2(.din(w_dff_B_2tEclMAK1_2),.dout(w_dff_B_lA9v8wsM5_2),.clk(gclk));
	jdff dff_B_KnaG4l6K5_2(.din(w_dff_B_lA9v8wsM5_2),.dout(w_dff_B_KnaG4l6K5_2),.clk(gclk));
	jdff dff_B_m0I4GfXp4_2(.din(w_dff_B_KnaG4l6K5_2),.dout(w_dff_B_m0I4GfXp4_2),.clk(gclk));
	jdff dff_B_dwd3x7Ia6_2(.din(w_dff_B_m0I4GfXp4_2),.dout(w_dff_B_dwd3x7Ia6_2),.clk(gclk));
	jdff dff_B_klRcr3bk7_2(.din(w_dff_B_dwd3x7Ia6_2),.dout(w_dff_B_klRcr3bk7_2),.clk(gclk));
	jdff dff_B_rl1m2nHq1_2(.din(w_dff_B_klRcr3bk7_2),.dout(w_dff_B_rl1m2nHq1_2),.clk(gclk));
	jdff dff_B_gO1gN7Ik5_2(.din(w_dff_B_rl1m2nHq1_2),.dout(w_dff_B_gO1gN7Ik5_2),.clk(gclk));
	jdff dff_B_GHym1I754_2(.din(w_dff_B_gO1gN7Ik5_2),.dout(w_dff_B_GHym1I754_2),.clk(gclk));
	jdff dff_B_jl9Ge0LM5_2(.din(w_dff_B_GHym1I754_2),.dout(w_dff_B_jl9Ge0LM5_2),.clk(gclk));
	jdff dff_B_x0QUaPVo7_2(.din(w_dff_B_jl9Ge0LM5_2),.dout(w_dff_B_x0QUaPVo7_2),.clk(gclk));
	jdff dff_B_4qNuKCMZ4_2(.din(w_dff_B_x0QUaPVo7_2),.dout(w_dff_B_4qNuKCMZ4_2),.clk(gclk));
	jdff dff_B_wWjawONr7_2(.din(w_dff_B_4qNuKCMZ4_2),.dout(w_dff_B_wWjawONr7_2),.clk(gclk));
	jdff dff_B_YrfYcJyl0_2(.din(w_dff_B_wWjawONr7_2),.dout(w_dff_B_YrfYcJyl0_2),.clk(gclk));
	jdff dff_B_ALQWyxbg3_2(.din(w_dff_B_YrfYcJyl0_2),.dout(w_dff_B_ALQWyxbg3_2),.clk(gclk));
	jdff dff_B_VxcZ4zR37_2(.din(w_dff_B_ALQWyxbg3_2),.dout(w_dff_B_VxcZ4zR37_2),.clk(gclk));
	jdff dff_B_3SSxB3xy1_2(.din(w_dff_B_VxcZ4zR37_2),.dout(w_dff_B_3SSxB3xy1_2),.clk(gclk));
	jdff dff_B_r00RNczI8_2(.din(w_dff_B_3SSxB3xy1_2),.dout(w_dff_B_r00RNczI8_2),.clk(gclk));
	jdff dff_B_6TmPeOpD3_2(.din(w_dff_B_r00RNczI8_2),.dout(w_dff_B_6TmPeOpD3_2),.clk(gclk));
	jdff dff_B_QQGQvHcR2_2(.din(w_dff_B_6TmPeOpD3_2),.dout(w_dff_B_QQGQvHcR2_2),.clk(gclk));
	jdff dff_B_uwyEBFDM8_2(.din(w_dff_B_QQGQvHcR2_2),.dout(w_dff_B_uwyEBFDM8_2),.clk(gclk));
	jdff dff_B_PWGYKLKY5_2(.din(w_dff_B_uwyEBFDM8_2),.dout(w_dff_B_PWGYKLKY5_2),.clk(gclk));
	jdff dff_B_e6K5chWS2_2(.din(w_dff_B_PWGYKLKY5_2),.dout(w_dff_B_e6K5chWS2_2),.clk(gclk));
	jdff dff_B_fj8Vgs8k0_2(.din(w_dff_B_e6K5chWS2_2),.dout(w_dff_B_fj8Vgs8k0_2),.clk(gclk));
	jdff dff_B_c0w64E9o7_2(.din(n817),.dout(w_dff_B_c0w64E9o7_2),.clk(gclk));
	jdff dff_B_mxcrFEy75_1(.din(n753),.dout(w_dff_B_mxcrFEy75_1),.clk(gclk));
	jdff dff_B_4OMtVokv1_2(.din(n659),.dout(w_dff_B_4OMtVokv1_2),.clk(gclk));
	jdff dff_B_acoRmwt28_2(.din(w_dff_B_4OMtVokv1_2),.dout(w_dff_B_acoRmwt28_2),.clk(gclk));
	jdff dff_B_9KkUNVVI6_2(.din(w_dff_B_acoRmwt28_2),.dout(w_dff_B_9KkUNVVI6_2),.clk(gclk));
	jdff dff_B_G1Bo0LPI7_2(.din(w_dff_B_9KkUNVVI6_2),.dout(w_dff_B_G1Bo0LPI7_2),.clk(gclk));
	jdff dff_B_JICtEKpQ8_2(.din(w_dff_B_G1Bo0LPI7_2),.dout(w_dff_B_JICtEKpQ8_2),.clk(gclk));
	jdff dff_B_pEUGoxrz8_2(.din(w_dff_B_JICtEKpQ8_2),.dout(w_dff_B_pEUGoxrz8_2),.clk(gclk));
	jdff dff_B_N306hy2O3_2(.din(w_dff_B_pEUGoxrz8_2),.dout(w_dff_B_N306hy2O3_2),.clk(gclk));
	jdff dff_B_lceEbzHj3_2(.din(w_dff_B_N306hy2O3_2),.dout(w_dff_B_lceEbzHj3_2),.clk(gclk));
	jdff dff_B_gFD0s3mq0_2(.din(w_dff_B_lceEbzHj3_2),.dout(w_dff_B_gFD0s3mq0_2),.clk(gclk));
	jdff dff_B_2lffssTC4_2(.din(w_dff_B_gFD0s3mq0_2),.dout(w_dff_B_2lffssTC4_2),.clk(gclk));
	jdff dff_B_Yxr7O1Uj6_2(.din(w_dff_B_2lffssTC4_2),.dout(w_dff_B_Yxr7O1Uj6_2),.clk(gclk));
	jdff dff_B_5YMx5so30_2(.din(w_dff_B_Yxr7O1Uj6_2),.dout(w_dff_B_5YMx5so30_2),.clk(gclk));
	jdff dff_B_oexpnFcj0_2(.din(w_dff_B_5YMx5so30_2),.dout(w_dff_B_oexpnFcj0_2),.clk(gclk));
	jdff dff_B_AQJqsCTT4_2(.din(w_dff_B_oexpnFcj0_2),.dout(w_dff_B_AQJqsCTT4_2),.clk(gclk));
	jdff dff_B_4psAA1UQ1_2(.din(w_dff_B_AQJqsCTT4_2),.dout(w_dff_B_4psAA1UQ1_2),.clk(gclk));
	jdff dff_B_0eo6v2GS3_2(.din(w_dff_B_4psAA1UQ1_2),.dout(w_dff_B_0eo6v2GS3_2),.clk(gclk));
	jdff dff_B_297USJ0g9_2(.din(w_dff_B_0eo6v2GS3_2),.dout(w_dff_B_297USJ0g9_2),.clk(gclk));
	jdff dff_B_mAYcP06y0_2(.din(w_dff_B_297USJ0g9_2),.dout(w_dff_B_mAYcP06y0_2),.clk(gclk));
	jdff dff_B_NGHXSi535_2(.din(w_dff_B_mAYcP06y0_2),.dout(w_dff_B_NGHXSi535_2),.clk(gclk));
	jdff dff_B_lU1WgcM25_2(.din(w_dff_B_NGHXSi535_2),.dout(w_dff_B_lU1WgcM25_2),.clk(gclk));
	jdff dff_B_phJ4JOgn2_2(.din(w_dff_B_lU1WgcM25_2),.dout(w_dff_B_phJ4JOgn2_2),.clk(gclk));
	jdff dff_B_6Lz8YEo09_2(.din(w_dff_B_phJ4JOgn2_2),.dout(w_dff_B_6Lz8YEo09_2),.clk(gclk));
	jdff dff_B_q7GzRp9T7_2(.din(w_dff_B_6Lz8YEo09_2),.dout(w_dff_B_q7GzRp9T7_2),.clk(gclk));
	jdff dff_B_43Y1xxIr5_2(.din(w_dff_B_q7GzRp9T7_2),.dout(w_dff_B_43Y1xxIr5_2),.clk(gclk));
	jdff dff_B_UDGVpLg17_2(.din(w_dff_B_43Y1xxIr5_2),.dout(w_dff_B_UDGVpLg17_2),.clk(gclk));
	jdff dff_B_ycB40T2b3_2(.din(n717),.dout(w_dff_B_ycB40T2b3_2),.clk(gclk));
	jdff dff_B_ygjs60Th7_1(.din(n660),.dout(w_dff_B_ygjs60Th7_1),.clk(gclk));
	jdff dff_B_Z0Duo9dV0_2(.din(n573),.dout(w_dff_B_Z0Duo9dV0_2),.clk(gclk));
	jdff dff_B_VRnX6mHH9_2(.din(w_dff_B_Z0Duo9dV0_2),.dout(w_dff_B_VRnX6mHH9_2),.clk(gclk));
	jdff dff_B_hXfiWR3P6_2(.din(w_dff_B_VRnX6mHH9_2),.dout(w_dff_B_hXfiWR3P6_2),.clk(gclk));
	jdff dff_B_3jIfXF6T0_2(.din(w_dff_B_hXfiWR3P6_2),.dout(w_dff_B_3jIfXF6T0_2),.clk(gclk));
	jdff dff_B_vdyx2JQE5_2(.din(w_dff_B_3jIfXF6T0_2),.dout(w_dff_B_vdyx2JQE5_2),.clk(gclk));
	jdff dff_B_lOPKwDuT8_2(.din(w_dff_B_vdyx2JQE5_2),.dout(w_dff_B_lOPKwDuT8_2),.clk(gclk));
	jdff dff_B_l3MrveyU8_2(.din(w_dff_B_lOPKwDuT8_2),.dout(w_dff_B_l3MrveyU8_2),.clk(gclk));
	jdff dff_B_4NWA4bwp0_2(.din(w_dff_B_l3MrveyU8_2),.dout(w_dff_B_4NWA4bwp0_2),.clk(gclk));
	jdff dff_B_eOjGzMjl3_2(.din(w_dff_B_4NWA4bwp0_2),.dout(w_dff_B_eOjGzMjl3_2),.clk(gclk));
	jdff dff_B_x5te0b223_2(.din(w_dff_B_eOjGzMjl3_2),.dout(w_dff_B_x5te0b223_2),.clk(gclk));
	jdff dff_B_ynbAoZOU9_2(.din(w_dff_B_x5te0b223_2),.dout(w_dff_B_ynbAoZOU9_2),.clk(gclk));
	jdff dff_B_oaA6cAh42_2(.din(w_dff_B_ynbAoZOU9_2),.dout(w_dff_B_oaA6cAh42_2),.clk(gclk));
	jdff dff_B_yBxAq33v3_2(.din(w_dff_B_oaA6cAh42_2),.dout(w_dff_B_yBxAq33v3_2),.clk(gclk));
	jdff dff_B_5faZdRXQ3_2(.din(w_dff_B_yBxAq33v3_2),.dout(w_dff_B_5faZdRXQ3_2),.clk(gclk));
	jdff dff_B_DyBzSxvy7_2(.din(w_dff_B_5faZdRXQ3_2),.dout(w_dff_B_DyBzSxvy7_2),.clk(gclk));
	jdff dff_B_b2UQyiTc7_2(.din(w_dff_B_DyBzSxvy7_2),.dout(w_dff_B_b2UQyiTc7_2),.clk(gclk));
	jdff dff_B_EjFXhMjI9_2(.din(w_dff_B_b2UQyiTc7_2),.dout(w_dff_B_EjFXhMjI9_2),.clk(gclk));
	jdff dff_B_O4ZLzo7Q7_2(.din(w_dff_B_EjFXhMjI9_2),.dout(w_dff_B_O4ZLzo7Q7_2),.clk(gclk));
	jdff dff_B_OEPcdrkb7_2(.din(w_dff_B_O4ZLzo7Q7_2),.dout(w_dff_B_OEPcdrkb7_2),.clk(gclk));
	jdff dff_B_arWQVsp99_2(.din(w_dff_B_OEPcdrkb7_2),.dout(w_dff_B_arWQVsp99_2),.clk(gclk));
	jdff dff_B_xctT5K701_2(.din(w_dff_B_arWQVsp99_2),.dout(w_dff_B_xctT5K701_2),.clk(gclk));
	jdff dff_B_DGBVxjsn9_2(.din(w_dff_B_xctT5K701_2),.dout(w_dff_B_DGBVxjsn9_2),.clk(gclk));
	jdff dff_B_vZ6KDoV16_2(.din(n624),.dout(w_dff_B_vZ6KDoV16_2),.clk(gclk));
	jdff dff_B_WMEeveX70_1(.din(n574),.dout(w_dff_B_WMEeveX70_1),.clk(gclk));
	jdff dff_B_8xYkexNR0_2(.din(n494),.dout(w_dff_B_8xYkexNR0_2),.clk(gclk));
	jdff dff_B_XchKCJZz6_2(.din(w_dff_B_8xYkexNR0_2),.dout(w_dff_B_XchKCJZz6_2),.clk(gclk));
	jdff dff_B_BcqWLi289_2(.din(w_dff_B_XchKCJZz6_2),.dout(w_dff_B_BcqWLi289_2),.clk(gclk));
	jdff dff_B_7Ixca6yZ6_2(.din(w_dff_B_BcqWLi289_2),.dout(w_dff_B_7Ixca6yZ6_2),.clk(gclk));
	jdff dff_B_GfjppUmw8_2(.din(w_dff_B_7Ixca6yZ6_2),.dout(w_dff_B_GfjppUmw8_2),.clk(gclk));
	jdff dff_B_TL87T78e5_2(.din(w_dff_B_GfjppUmw8_2),.dout(w_dff_B_TL87T78e5_2),.clk(gclk));
	jdff dff_B_c6ACRB5u9_2(.din(w_dff_B_TL87T78e5_2),.dout(w_dff_B_c6ACRB5u9_2),.clk(gclk));
	jdff dff_B_7NIqPGV22_2(.din(w_dff_B_c6ACRB5u9_2),.dout(w_dff_B_7NIqPGV22_2),.clk(gclk));
	jdff dff_B_648NKTum2_2(.din(w_dff_B_7NIqPGV22_2),.dout(w_dff_B_648NKTum2_2),.clk(gclk));
	jdff dff_B_uf0MxER77_2(.din(w_dff_B_648NKTum2_2),.dout(w_dff_B_uf0MxER77_2),.clk(gclk));
	jdff dff_B_zrLxTw9F9_2(.din(w_dff_B_uf0MxER77_2),.dout(w_dff_B_zrLxTw9F9_2),.clk(gclk));
	jdff dff_B_8H5kqOg08_2(.din(w_dff_B_zrLxTw9F9_2),.dout(w_dff_B_8H5kqOg08_2),.clk(gclk));
	jdff dff_B_lCivCT015_2(.din(w_dff_B_8H5kqOg08_2),.dout(w_dff_B_lCivCT015_2),.clk(gclk));
	jdff dff_B_qMyG07dM2_2(.din(w_dff_B_lCivCT015_2),.dout(w_dff_B_qMyG07dM2_2),.clk(gclk));
	jdff dff_B_TGb8nIso0_2(.din(w_dff_B_qMyG07dM2_2),.dout(w_dff_B_TGb8nIso0_2),.clk(gclk));
	jdff dff_B_HDWsRIIj2_2(.din(w_dff_B_TGb8nIso0_2),.dout(w_dff_B_HDWsRIIj2_2),.clk(gclk));
	jdff dff_B_DsXCdJIH8_2(.din(w_dff_B_HDWsRIIj2_2),.dout(w_dff_B_DsXCdJIH8_2),.clk(gclk));
	jdff dff_B_sKSNMA531_2(.din(w_dff_B_DsXCdJIH8_2),.dout(w_dff_B_sKSNMA531_2),.clk(gclk));
	jdff dff_B_A3MxRWOn7_2(.din(w_dff_B_sKSNMA531_2),.dout(w_dff_B_A3MxRWOn7_2),.clk(gclk));
	jdff dff_B_DFyyoA0N0_2(.din(n538),.dout(w_dff_B_DFyyoA0N0_2),.clk(gclk));
	jdff dff_B_VvhQZ0NB6_1(.din(n495),.dout(w_dff_B_VvhQZ0NB6_1),.clk(gclk));
	jdff dff_B_pgbrNAnr1_2(.din(n422),.dout(w_dff_B_pgbrNAnr1_2),.clk(gclk));
	jdff dff_B_bEdYUBvI7_2(.din(w_dff_B_pgbrNAnr1_2),.dout(w_dff_B_bEdYUBvI7_2),.clk(gclk));
	jdff dff_B_zugL85Ye3_2(.din(w_dff_B_bEdYUBvI7_2),.dout(w_dff_B_zugL85Ye3_2),.clk(gclk));
	jdff dff_B_i48PGo582_2(.din(w_dff_B_zugL85Ye3_2),.dout(w_dff_B_i48PGo582_2),.clk(gclk));
	jdff dff_B_te4HLu1p9_2(.din(w_dff_B_i48PGo582_2),.dout(w_dff_B_te4HLu1p9_2),.clk(gclk));
	jdff dff_B_hwMFpPo93_2(.din(w_dff_B_te4HLu1p9_2),.dout(w_dff_B_hwMFpPo93_2),.clk(gclk));
	jdff dff_B_A60vuWWt2_2(.din(w_dff_B_hwMFpPo93_2),.dout(w_dff_B_A60vuWWt2_2),.clk(gclk));
	jdff dff_B_EQBRvvYW5_2(.din(w_dff_B_A60vuWWt2_2),.dout(w_dff_B_EQBRvvYW5_2),.clk(gclk));
	jdff dff_B_QIrZ9R2b6_2(.din(w_dff_B_EQBRvvYW5_2),.dout(w_dff_B_QIrZ9R2b6_2),.clk(gclk));
	jdff dff_B_aDMKBFu62_2(.din(w_dff_B_QIrZ9R2b6_2),.dout(w_dff_B_aDMKBFu62_2),.clk(gclk));
	jdff dff_B_HTRPVf4C5_2(.din(w_dff_B_aDMKBFu62_2),.dout(w_dff_B_HTRPVf4C5_2),.clk(gclk));
	jdff dff_B_ziCjGJz67_2(.din(w_dff_B_HTRPVf4C5_2),.dout(w_dff_B_ziCjGJz67_2),.clk(gclk));
	jdff dff_B_eIRFFKhB0_2(.din(w_dff_B_ziCjGJz67_2),.dout(w_dff_B_eIRFFKhB0_2),.clk(gclk));
	jdff dff_B_txtJm3rF6_2(.din(w_dff_B_eIRFFKhB0_2),.dout(w_dff_B_txtJm3rF6_2),.clk(gclk));
	jdff dff_B_k4XIAjuc1_2(.din(w_dff_B_txtJm3rF6_2),.dout(w_dff_B_k4XIAjuc1_2),.clk(gclk));
	jdff dff_B_RNkWNosq9_2(.din(w_dff_B_k4XIAjuc1_2),.dout(w_dff_B_RNkWNosq9_2),.clk(gclk));
	jdff dff_B_J6QBkd1c4_2(.din(n459),.dout(w_dff_B_J6QBkd1c4_2),.clk(gclk));
	jdff dff_B_UaNQnCtd9_1(.din(n423),.dout(w_dff_B_UaNQnCtd9_1),.clk(gclk));
	jdff dff_B_dighet794_2(.din(n358),.dout(w_dff_B_dighet794_2),.clk(gclk));
	jdff dff_B_XMXdOW4Z5_2(.din(w_dff_B_dighet794_2),.dout(w_dff_B_XMXdOW4Z5_2),.clk(gclk));
	jdff dff_B_vKmnixM04_2(.din(w_dff_B_XMXdOW4Z5_2),.dout(w_dff_B_vKmnixM04_2),.clk(gclk));
	jdff dff_B_MoWautym2_2(.din(w_dff_B_vKmnixM04_2),.dout(w_dff_B_MoWautym2_2),.clk(gclk));
	jdff dff_B_758aSQuj9_2(.din(w_dff_B_MoWautym2_2),.dout(w_dff_B_758aSQuj9_2),.clk(gclk));
	jdff dff_B_dFY0FqmX0_2(.din(w_dff_B_758aSQuj9_2),.dout(w_dff_B_dFY0FqmX0_2),.clk(gclk));
	jdff dff_B_ht9z6Nlz5_2(.din(w_dff_B_dFY0FqmX0_2),.dout(w_dff_B_ht9z6Nlz5_2),.clk(gclk));
	jdff dff_B_6LLvWaqw6_2(.din(w_dff_B_ht9z6Nlz5_2),.dout(w_dff_B_6LLvWaqw6_2),.clk(gclk));
	jdff dff_B_neqTqmG74_2(.din(w_dff_B_6LLvWaqw6_2),.dout(w_dff_B_neqTqmG74_2),.clk(gclk));
	jdff dff_B_NsYz8Tbc1_2(.din(w_dff_B_neqTqmG74_2),.dout(w_dff_B_NsYz8Tbc1_2),.clk(gclk));
	jdff dff_B_0bhSfjpg3_2(.din(w_dff_B_NsYz8Tbc1_2),.dout(w_dff_B_0bhSfjpg3_2),.clk(gclk));
	jdff dff_B_WSbE96bQ3_2(.din(w_dff_B_0bhSfjpg3_2),.dout(w_dff_B_WSbE96bQ3_2),.clk(gclk));
	jdff dff_B_TCa8Nxe60_2(.din(w_dff_B_WSbE96bQ3_2),.dout(w_dff_B_TCa8Nxe60_2),.clk(gclk));
	jdff dff_B_nnVOysn11_2(.din(n387),.dout(w_dff_B_nnVOysn11_2),.clk(gclk));
	jdff dff_B_ztAH3VDi4_1(.din(n359),.dout(w_dff_B_ztAH3VDi4_1),.clk(gclk));
	jdff dff_B_mwJc1BeS3_2(.din(n300),.dout(w_dff_B_mwJc1BeS3_2),.clk(gclk));
	jdff dff_B_3sxCiYtf9_2(.din(w_dff_B_mwJc1BeS3_2),.dout(w_dff_B_3sxCiYtf9_2),.clk(gclk));
	jdff dff_B_RLpQhle37_2(.din(w_dff_B_3sxCiYtf9_2),.dout(w_dff_B_RLpQhle37_2),.clk(gclk));
	jdff dff_B_b01OVPTv4_2(.din(w_dff_B_RLpQhle37_2),.dout(w_dff_B_b01OVPTv4_2),.clk(gclk));
	jdff dff_B_YVIsgybR5_2(.din(w_dff_B_b01OVPTv4_2),.dout(w_dff_B_YVIsgybR5_2),.clk(gclk));
	jdff dff_B_B7qquJtX8_2(.din(w_dff_B_YVIsgybR5_2),.dout(w_dff_B_B7qquJtX8_2),.clk(gclk));
	jdff dff_B_Ea8Tq7lI1_2(.din(w_dff_B_B7qquJtX8_2),.dout(w_dff_B_Ea8Tq7lI1_2),.clk(gclk));
	jdff dff_B_qcWevvG74_2(.din(w_dff_B_Ea8Tq7lI1_2),.dout(w_dff_B_qcWevvG74_2),.clk(gclk));
	jdff dff_B_5s5oyIZD3_2(.din(w_dff_B_qcWevvG74_2),.dout(w_dff_B_5s5oyIZD3_2),.clk(gclk));
	jdff dff_B_BMfrFhAf7_2(.din(w_dff_B_5s5oyIZD3_2),.dout(w_dff_B_BMfrFhAf7_2),.clk(gclk));
	jdff dff_B_cFedhM6m6_2(.din(n323),.dout(w_dff_B_cFedhM6m6_2),.clk(gclk));
	jdff dff_B_lIUTpAE80_1(.din(n301),.dout(w_dff_B_lIUTpAE80_1),.clk(gclk));
	jdff dff_B_uL5pjgHx5_2(.din(n249),.dout(w_dff_B_uL5pjgHx5_2),.clk(gclk));
	jdff dff_B_tHoIgdej0_2(.din(w_dff_B_uL5pjgHx5_2),.dout(w_dff_B_tHoIgdej0_2),.clk(gclk));
	jdff dff_B_VQfOBjtP3_2(.din(w_dff_B_tHoIgdej0_2),.dout(w_dff_B_VQfOBjtP3_2),.clk(gclk));
	jdff dff_B_xiJINwsA5_2(.din(w_dff_B_VQfOBjtP3_2),.dout(w_dff_B_xiJINwsA5_2),.clk(gclk));
	jdff dff_B_3ZyEqvnH6_2(.din(w_dff_B_xiJINwsA5_2),.dout(w_dff_B_3ZyEqvnH6_2),.clk(gclk));
	jdff dff_B_BG0lSzJ73_2(.din(w_dff_B_3ZyEqvnH6_2),.dout(w_dff_B_BG0lSzJ73_2),.clk(gclk));
	jdff dff_B_9cmf9K3G9_2(.din(w_dff_B_BG0lSzJ73_2),.dout(w_dff_B_9cmf9K3G9_2),.clk(gclk));
	jdff dff_B_nalj3afZ5_2(.din(n265),.dout(w_dff_B_nalj3afZ5_2),.clk(gclk));
	jdff dff_B_BmR3h8NF0_1(.din(n250),.dout(w_dff_B_BmR3h8NF0_1),.clk(gclk));
	jdff dff_B_fEsB0Ljq9_0(.din(n214),.dout(w_dff_B_fEsB0Ljq9_0),.clk(gclk));
	jdff dff_B_Su4WFigI8_2(.din(n206),.dout(w_dff_B_Su4WFigI8_2),.clk(gclk));
	jdff dff_B_jnLnM26k1_2(.din(w_dff_B_Su4WFigI8_2),.dout(w_dff_B_jnLnM26k1_2),.clk(gclk));
	jdff dff_B_nHW52yND5_2(.din(w_dff_B_jnLnM26k1_2),.dout(w_dff_B_nHW52yND5_2),.clk(gclk));
	jdff dff_B_psp5KmyI1_2(.din(w_dff_B_nHW52yND5_2),.dout(w_dff_B_psp5KmyI1_2),.clk(gclk));
	jdff dff_B_74u3CizV5_1(.din(n208),.dout(w_dff_B_74u3CizV5_1),.clk(gclk));
	jdff dff_A_lY35Gf6q5_0(.dout(w_n210_1[0]),.din(w_dff_A_lY35Gf6q5_0),.clk(gclk));
	jdff dff_A_4KBjmpb35_0(.dout(w_n169_0[0]),.din(w_dff_A_4KBjmpb35_0),.clk(gclk));
	jdff dff_A_g6U8xrxE7_0(.dout(w_dff_A_4KBjmpb35_0),.din(w_dff_A_g6U8xrxE7_0),.clk(gclk));
	jdff dff_A_IX8YLItY8_1(.dout(w_n169_0[1]),.din(w_dff_A_IX8YLItY8_1),.clk(gclk));
	jdff dff_B_5P4pp9zh5_2(.din(n1420),.dout(w_dff_B_5P4pp9zh5_2),.clk(gclk));
	jdff dff_B_2YkkQ9rd3_1(.din(n1418),.dout(w_dff_B_2YkkQ9rd3_1),.clk(gclk));
	jdff dff_B_JuqYWJY15_2(.din(n1338),.dout(w_dff_B_JuqYWJY15_2),.clk(gclk));
	jdff dff_B_MFOTu59Z4_2(.din(w_dff_B_JuqYWJY15_2),.dout(w_dff_B_MFOTu59Z4_2),.clk(gclk));
	jdff dff_B_pUrciEDZ6_2(.din(w_dff_B_MFOTu59Z4_2),.dout(w_dff_B_pUrciEDZ6_2),.clk(gclk));
	jdff dff_B_ae0rn1Vl9_2(.din(w_dff_B_pUrciEDZ6_2),.dout(w_dff_B_ae0rn1Vl9_2),.clk(gclk));
	jdff dff_B_QQMrrVrk5_2(.din(w_dff_B_ae0rn1Vl9_2),.dout(w_dff_B_QQMrrVrk5_2),.clk(gclk));
	jdff dff_B_4kSfgJ1w5_2(.din(w_dff_B_QQMrrVrk5_2),.dout(w_dff_B_4kSfgJ1w5_2),.clk(gclk));
	jdff dff_B_lm8Xe7PB3_2(.din(w_dff_B_4kSfgJ1w5_2),.dout(w_dff_B_lm8Xe7PB3_2),.clk(gclk));
	jdff dff_B_oohCaw863_2(.din(w_dff_B_lm8Xe7PB3_2),.dout(w_dff_B_oohCaw863_2),.clk(gclk));
	jdff dff_B_ZKqaoZ7F4_2(.din(w_dff_B_oohCaw863_2),.dout(w_dff_B_ZKqaoZ7F4_2),.clk(gclk));
	jdff dff_B_9n80JxzK0_2(.din(w_dff_B_ZKqaoZ7F4_2),.dout(w_dff_B_9n80JxzK0_2),.clk(gclk));
	jdff dff_B_9GOdYVMe1_2(.din(w_dff_B_9n80JxzK0_2),.dout(w_dff_B_9GOdYVMe1_2),.clk(gclk));
	jdff dff_B_W0HuBbm93_2(.din(w_dff_B_9GOdYVMe1_2),.dout(w_dff_B_W0HuBbm93_2),.clk(gclk));
	jdff dff_B_2WXWACs30_2(.din(w_dff_B_W0HuBbm93_2),.dout(w_dff_B_2WXWACs30_2),.clk(gclk));
	jdff dff_B_ItzjVcsw5_2(.din(w_dff_B_2WXWACs30_2),.dout(w_dff_B_ItzjVcsw5_2),.clk(gclk));
	jdff dff_B_jSscDheQ5_2(.din(w_dff_B_ItzjVcsw5_2),.dout(w_dff_B_jSscDheQ5_2),.clk(gclk));
	jdff dff_B_IFADsWC58_2(.din(w_dff_B_jSscDheQ5_2),.dout(w_dff_B_IFADsWC58_2),.clk(gclk));
	jdff dff_B_X2amMj6X1_2(.din(w_dff_B_IFADsWC58_2),.dout(w_dff_B_X2amMj6X1_2),.clk(gclk));
	jdff dff_B_hz0cZMFW7_2(.din(w_dff_B_X2amMj6X1_2),.dout(w_dff_B_hz0cZMFW7_2),.clk(gclk));
	jdff dff_B_R3E6d6yl4_2(.din(w_dff_B_hz0cZMFW7_2),.dout(w_dff_B_R3E6d6yl4_2),.clk(gclk));
	jdff dff_B_Jtl4fyGM1_2(.din(w_dff_B_R3E6d6yl4_2),.dout(w_dff_B_Jtl4fyGM1_2),.clk(gclk));
	jdff dff_B_0iPHElpd8_2(.din(w_dff_B_Jtl4fyGM1_2),.dout(w_dff_B_0iPHElpd8_2),.clk(gclk));
	jdff dff_B_sCXxBtso0_2(.din(w_dff_B_0iPHElpd8_2),.dout(w_dff_B_sCXxBtso0_2),.clk(gclk));
	jdff dff_B_hgajkR5L3_2(.din(w_dff_B_sCXxBtso0_2),.dout(w_dff_B_hgajkR5L3_2),.clk(gclk));
	jdff dff_B_MflVSr1N3_2(.din(w_dff_B_hgajkR5L3_2),.dout(w_dff_B_MflVSr1N3_2),.clk(gclk));
	jdff dff_B_uFbs19s49_2(.din(w_dff_B_MflVSr1N3_2),.dout(w_dff_B_uFbs19s49_2),.clk(gclk));
	jdff dff_B_JdRzqbq86_2(.din(w_dff_B_uFbs19s49_2),.dout(w_dff_B_JdRzqbq86_2),.clk(gclk));
	jdff dff_B_uEbBayz01_2(.din(w_dff_B_JdRzqbq86_2),.dout(w_dff_B_uEbBayz01_2),.clk(gclk));
	jdff dff_B_966hOrhk2_2(.din(w_dff_B_uEbBayz01_2),.dout(w_dff_B_966hOrhk2_2),.clk(gclk));
	jdff dff_B_TG4B0ySn7_2(.din(w_dff_B_966hOrhk2_2),.dout(w_dff_B_TG4B0ySn7_2),.clk(gclk));
	jdff dff_B_vUJgjzdo4_2(.din(w_dff_B_TG4B0ySn7_2),.dout(w_dff_B_vUJgjzdo4_2),.clk(gclk));
	jdff dff_B_1Zqukoio1_2(.din(w_dff_B_vUJgjzdo4_2),.dout(w_dff_B_1Zqukoio1_2),.clk(gclk));
	jdff dff_B_QgioRiTJ3_2(.din(w_dff_B_1Zqukoio1_2),.dout(w_dff_B_QgioRiTJ3_2),.clk(gclk));
	jdff dff_B_m8IPSO2E5_2(.din(w_dff_B_QgioRiTJ3_2),.dout(w_dff_B_m8IPSO2E5_2),.clk(gclk));
	jdff dff_B_z0uyovCq3_2(.din(w_dff_B_m8IPSO2E5_2),.dout(w_dff_B_z0uyovCq3_2),.clk(gclk));
	jdff dff_B_6P9Ru5e75_2(.din(w_dff_B_z0uyovCq3_2),.dout(w_dff_B_6P9Ru5e75_2),.clk(gclk));
	jdff dff_B_Mf8FdXk30_2(.din(w_dff_B_6P9Ru5e75_2),.dout(w_dff_B_Mf8FdXk30_2),.clk(gclk));
	jdff dff_B_2vxJTD2u6_2(.din(w_dff_B_Mf8FdXk30_2),.dout(w_dff_B_2vxJTD2u6_2),.clk(gclk));
	jdff dff_B_zKVWfg8V0_2(.din(w_dff_B_2vxJTD2u6_2),.dout(w_dff_B_zKVWfg8V0_2),.clk(gclk));
	jdff dff_B_tzpUw0ad2_2(.din(w_dff_B_zKVWfg8V0_2),.dout(w_dff_B_tzpUw0ad2_2),.clk(gclk));
	jdff dff_B_SicE7c7A6_2(.din(w_dff_B_tzpUw0ad2_2),.dout(w_dff_B_SicE7c7A6_2),.clk(gclk));
	jdff dff_B_uumtACLN2_2(.din(w_dff_B_SicE7c7A6_2),.dout(w_dff_B_uumtACLN2_2),.clk(gclk));
	jdff dff_B_FZ6IXBKU5_2(.din(w_dff_B_uumtACLN2_2),.dout(w_dff_B_FZ6IXBKU5_2),.clk(gclk));
	jdff dff_B_cSvpNLU87_2(.din(w_dff_B_FZ6IXBKU5_2),.dout(w_dff_B_cSvpNLU87_2),.clk(gclk));
	jdff dff_B_GjTXKUHD5_2(.din(w_dff_B_cSvpNLU87_2),.dout(w_dff_B_GjTXKUHD5_2),.clk(gclk));
	jdff dff_B_mJ9wVZH48_2(.din(w_dff_B_GjTXKUHD5_2),.dout(w_dff_B_mJ9wVZH48_2),.clk(gclk));
	jdff dff_B_Y7cEae5U1_1(.din(n1339),.dout(w_dff_B_Y7cEae5U1_1),.clk(gclk));
	jdff dff_B_R0URrd2P3_2(.din(n1253),.dout(w_dff_B_R0URrd2P3_2),.clk(gclk));
	jdff dff_B_hwqMBUsx1_2(.din(w_dff_B_R0URrd2P3_2),.dout(w_dff_B_hwqMBUsx1_2),.clk(gclk));
	jdff dff_B_YErTvJtL1_2(.din(w_dff_B_hwqMBUsx1_2),.dout(w_dff_B_YErTvJtL1_2),.clk(gclk));
	jdff dff_B_zut8PZZn6_2(.din(w_dff_B_YErTvJtL1_2),.dout(w_dff_B_zut8PZZn6_2),.clk(gclk));
	jdff dff_B_UbOtM6RN0_2(.din(w_dff_B_zut8PZZn6_2),.dout(w_dff_B_UbOtM6RN0_2),.clk(gclk));
	jdff dff_B_wieL0KOK9_2(.din(w_dff_B_UbOtM6RN0_2),.dout(w_dff_B_wieL0KOK9_2),.clk(gclk));
	jdff dff_B_pej1ijAG6_2(.din(w_dff_B_wieL0KOK9_2),.dout(w_dff_B_pej1ijAG6_2),.clk(gclk));
	jdff dff_B_8IfK4BbJ0_2(.din(w_dff_B_pej1ijAG6_2),.dout(w_dff_B_8IfK4BbJ0_2),.clk(gclk));
	jdff dff_B_wzqxTmUW5_2(.din(w_dff_B_8IfK4BbJ0_2),.dout(w_dff_B_wzqxTmUW5_2),.clk(gclk));
	jdff dff_B_3zUfbgfe6_2(.din(w_dff_B_wzqxTmUW5_2),.dout(w_dff_B_3zUfbgfe6_2),.clk(gclk));
	jdff dff_B_9u2PPMPm8_2(.din(w_dff_B_3zUfbgfe6_2),.dout(w_dff_B_9u2PPMPm8_2),.clk(gclk));
	jdff dff_B_somNHLV52_2(.din(w_dff_B_9u2PPMPm8_2),.dout(w_dff_B_somNHLV52_2),.clk(gclk));
	jdff dff_B_wL41hHxW5_2(.din(w_dff_B_somNHLV52_2),.dout(w_dff_B_wL41hHxW5_2),.clk(gclk));
	jdff dff_B_j9GT010h3_2(.din(w_dff_B_wL41hHxW5_2),.dout(w_dff_B_j9GT010h3_2),.clk(gclk));
	jdff dff_B_cX1W1JIx9_2(.din(w_dff_B_j9GT010h3_2),.dout(w_dff_B_cX1W1JIx9_2),.clk(gclk));
	jdff dff_B_8jhoHevL2_2(.din(w_dff_B_cX1W1JIx9_2),.dout(w_dff_B_8jhoHevL2_2),.clk(gclk));
	jdff dff_B_uC7tnTzC1_2(.din(w_dff_B_8jhoHevL2_2),.dout(w_dff_B_uC7tnTzC1_2),.clk(gclk));
	jdff dff_B_EbtojuWS9_2(.din(w_dff_B_uC7tnTzC1_2),.dout(w_dff_B_EbtojuWS9_2),.clk(gclk));
	jdff dff_B_ev9XnmBM8_2(.din(w_dff_B_EbtojuWS9_2),.dout(w_dff_B_ev9XnmBM8_2),.clk(gclk));
	jdff dff_B_wOC6kAbp3_2(.din(w_dff_B_ev9XnmBM8_2),.dout(w_dff_B_wOC6kAbp3_2),.clk(gclk));
	jdff dff_B_rgSopqSd3_2(.din(w_dff_B_wOC6kAbp3_2),.dout(w_dff_B_rgSopqSd3_2),.clk(gclk));
	jdff dff_B_4LkbpIWS1_2(.din(w_dff_B_rgSopqSd3_2),.dout(w_dff_B_4LkbpIWS1_2),.clk(gclk));
	jdff dff_B_Cd3jsIgJ2_2(.din(w_dff_B_4LkbpIWS1_2),.dout(w_dff_B_Cd3jsIgJ2_2),.clk(gclk));
	jdff dff_B_Jzi6yvEP6_2(.din(w_dff_B_Cd3jsIgJ2_2),.dout(w_dff_B_Jzi6yvEP6_2),.clk(gclk));
	jdff dff_B_fF6d4owR2_2(.din(w_dff_B_Jzi6yvEP6_2),.dout(w_dff_B_fF6d4owR2_2),.clk(gclk));
	jdff dff_B_CBEP8Hgy4_2(.din(w_dff_B_fF6d4owR2_2),.dout(w_dff_B_CBEP8Hgy4_2),.clk(gclk));
	jdff dff_B_eEsFpIIl4_2(.din(w_dff_B_CBEP8Hgy4_2),.dout(w_dff_B_eEsFpIIl4_2),.clk(gclk));
	jdff dff_B_b2m5Bg1A5_2(.din(w_dff_B_eEsFpIIl4_2),.dout(w_dff_B_b2m5Bg1A5_2),.clk(gclk));
	jdff dff_B_h6bXhJra1_2(.din(w_dff_B_b2m5Bg1A5_2),.dout(w_dff_B_h6bXhJra1_2),.clk(gclk));
	jdff dff_B_PAMu7WGB0_2(.din(w_dff_B_h6bXhJra1_2),.dout(w_dff_B_PAMu7WGB0_2),.clk(gclk));
	jdff dff_B_2Bnc9tCI2_2(.din(w_dff_B_PAMu7WGB0_2),.dout(w_dff_B_2Bnc9tCI2_2),.clk(gclk));
	jdff dff_B_NyIK2i0x2_2(.din(w_dff_B_2Bnc9tCI2_2),.dout(w_dff_B_NyIK2i0x2_2),.clk(gclk));
	jdff dff_B_KJkA6zte2_2(.din(w_dff_B_NyIK2i0x2_2),.dout(w_dff_B_KJkA6zte2_2),.clk(gclk));
	jdff dff_B_DCwdtyls8_2(.din(w_dff_B_KJkA6zte2_2),.dout(w_dff_B_DCwdtyls8_2),.clk(gclk));
	jdff dff_B_nYNWCZCP3_2(.din(w_dff_B_DCwdtyls8_2),.dout(w_dff_B_nYNWCZCP3_2),.clk(gclk));
	jdff dff_B_3jzPG3fB9_2(.din(w_dff_B_nYNWCZCP3_2),.dout(w_dff_B_3jzPG3fB9_2),.clk(gclk));
	jdff dff_B_fzmUEzNP9_2(.din(w_dff_B_3jzPG3fB9_2),.dout(w_dff_B_fzmUEzNP9_2),.clk(gclk));
	jdff dff_B_Krivrsg29_2(.din(w_dff_B_fzmUEzNP9_2),.dout(w_dff_B_Krivrsg29_2),.clk(gclk));
	jdff dff_B_MIEuH8hx6_2(.din(w_dff_B_Krivrsg29_2),.dout(w_dff_B_MIEuH8hx6_2),.clk(gclk));
	jdff dff_B_zS3qZF2g9_2(.din(w_dff_B_MIEuH8hx6_2),.dout(w_dff_B_zS3qZF2g9_2),.clk(gclk));
	jdff dff_B_veZHBUJv1_1(.din(n1254),.dout(w_dff_B_veZHBUJv1_1),.clk(gclk));
	jdff dff_B_lLeaJOqU6_2(.din(n1163),.dout(w_dff_B_lLeaJOqU6_2),.clk(gclk));
	jdff dff_B_Gpc8TddJ5_2(.din(w_dff_B_lLeaJOqU6_2),.dout(w_dff_B_Gpc8TddJ5_2),.clk(gclk));
	jdff dff_B_3dtFcCsZ5_2(.din(w_dff_B_Gpc8TddJ5_2),.dout(w_dff_B_3dtFcCsZ5_2),.clk(gclk));
	jdff dff_B_NgCwOr0u0_2(.din(w_dff_B_3dtFcCsZ5_2),.dout(w_dff_B_NgCwOr0u0_2),.clk(gclk));
	jdff dff_B_4oDTmw7D5_2(.din(w_dff_B_NgCwOr0u0_2),.dout(w_dff_B_4oDTmw7D5_2),.clk(gclk));
	jdff dff_B_HJtdDzz43_2(.din(w_dff_B_4oDTmw7D5_2),.dout(w_dff_B_HJtdDzz43_2),.clk(gclk));
	jdff dff_B_VEuFlud65_2(.din(w_dff_B_HJtdDzz43_2),.dout(w_dff_B_VEuFlud65_2),.clk(gclk));
	jdff dff_B_JW6v6wyL5_2(.din(w_dff_B_VEuFlud65_2),.dout(w_dff_B_JW6v6wyL5_2),.clk(gclk));
	jdff dff_B_r83ELxry2_2(.din(w_dff_B_JW6v6wyL5_2),.dout(w_dff_B_r83ELxry2_2),.clk(gclk));
	jdff dff_B_LOIXOIv78_2(.din(w_dff_B_r83ELxry2_2),.dout(w_dff_B_LOIXOIv78_2),.clk(gclk));
	jdff dff_B_F6yoJNjV6_2(.din(w_dff_B_LOIXOIv78_2),.dout(w_dff_B_F6yoJNjV6_2),.clk(gclk));
	jdff dff_B_zLLd9rv06_2(.din(w_dff_B_F6yoJNjV6_2),.dout(w_dff_B_zLLd9rv06_2),.clk(gclk));
	jdff dff_B_2BhHRQih1_2(.din(w_dff_B_zLLd9rv06_2),.dout(w_dff_B_2BhHRQih1_2),.clk(gclk));
	jdff dff_B_JB3k6geG3_2(.din(w_dff_B_2BhHRQih1_2),.dout(w_dff_B_JB3k6geG3_2),.clk(gclk));
	jdff dff_B_5q3NxEkH7_2(.din(w_dff_B_JB3k6geG3_2),.dout(w_dff_B_5q3NxEkH7_2),.clk(gclk));
	jdff dff_B_eSBQStM02_2(.din(w_dff_B_5q3NxEkH7_2),.dout(w_dff_B_eSBQStM02_2),.clk(gclk));
	jdff dff_B_Y8TEAzYS5_2(.din(w_dff_B_eSBQStM02_2),.dout(w_dff_B_Y8TEAzYS5_2),.clk(gclk));
	jdff dff_B_p9w5r6di2_2(.din(w_dff_B_Y8TEAzYS5_2),.dout(w_dff_B_p9w5r6di2_2),.clk(gclk));
	jdff dff_B_o7hHWP8Z2_2(.din(w_dff_B_p9w5r6di2_2),.dout(w_dff_B_o7hHWP8Z2_2),.clk(gclk));
	jdff dff_B_Nn3vFM4n8_2(.din(w_dff_B_o7hHWP8Z2_2),.dout(w_dff_B_Nn3vFM4n8_2),.clk(gclk));
	jdff dff_B_tSw5WrnD2_2(.din(w_dff_B_Nn3vFM4n8_2),.dout(w_dff_B_tSw5WrnD2_2),.clk(gclk));
	jdff dff_B_61w3WLDm2_2(.din(w_dff_B_tSw5WrnD2_2),.dout(w_dff_B_61w3WLDm2_2),.clk(gclk));
	jdff dff_B_P17ohZkU7_2(.din(w_dff_B_61w3WLDm2_2),.dout(w_dff_B_P17ohZkU7_2),.clk(gclk));
	jdff dff_B_RjHV7ITZ0_2(.din(w_dff_B_P17ohZkU7_2),.dout(w_dff_B_RjHV7ITZ0_2),.clk(gclk));
	jdff dff_B_9Tz4lley7_2(.din(w_dff_B_RjHV7ITZ0_2),.dout(w_dff_B_9Tz4lley7_2),.clk(gclk));
	jdff dff_B_QkGmoXMf7_2(.din(w_dff_B_9Tz4lley7_2),.dout(w_dff_B_QkGmoXMf7_2),.clk(gclk));
	jdff dff_B_6sVUDqCe5_2(.din(w_dff_B_QkGmoXMf7_2),.dout(w_dff_B_6sVUDqCe5_2),.clk(gclk));
	jdff dff_B_VwWx60VY1_2(.din(w_dff_B_6sVUDqCe5_2),.dout(w_dff_B_VwWx60VY1_2),.clk(gclk));
	jdff dff_B_czw2cOJi9_2(.din(w_dff_B_VwWx60VY1_2),.dout(w_dff_B_czw2cOJi9_2),.clk(gclk));
	jdff dff_B_NZD7xLZ20_2(.din(w_dff_B_czw2cOJi9_2),.dout(w_dff_B_NZD7xLZ20_2),.clk(gclk));
	jdff dff_B_bXjCGVl78_2(.din(w_dff_B_NZD7xLZ20_2),.dout(w_dff_B_bXjCGVl78_2),.clk(gclk));
	jdff dff_B_ViKNaZDL6_2(.din(w_dff_B_bXjCGVl78_2),.dout(w_dff_B_ViKNaZDL6_2),.clk(gclk));
	jdff dff_B_xm6oSMuN9_2(.din(w_dff_B_ViKNaZDL6_2),.dout(w_dff_B_xm6oSMuN9_2),.clk(gclk));
	jdff dff_B_w1Q7IhUT5_2(.din(w_dff_B_xm6oSMuN9_2),.dout(w_dff_B_w1Q7IhUT5_2),.clk(gclk));
	jdff dff_B_g0wfKieS7_2(.din(w_dff_B_w1Q7IhUT5_2),.dout(w_dff_B_g0wfKieS7_2),.clk(gclk));
	jdff dff_B_yb8ttNkF6_2(.din(w_dff_B_g0wfKieS7_2),.dout(w_dff_B_yb8ttNkF6_2),.clk(gclk));
	jdff dff_B_WFUfie7T9_2(.din(w_dff_B_yb8ttNkF6_2),.dout(w_dff_B_WFUfie7T9_2),.clk(gclk));
	jdff dff_B_uOEOZObL3_1(.din(n1164),.dout(w_dff_B_uOEOZObL3_1),.clk(gclk));
	jdff dff_B_1ojTqbuu5_2(.din(n1059),.dout(w_dff_B_1ojTqbuu5_2),.clk(gclk));
	jdff dff_B_Mu1h62B41_2(.din(w_dff_B_1ojTqbuu5_2),.dout(w_dff_B_Mu1h62B41_2),.clk(gclk));
	jdff dff_B_h48RORwK8_2(.din(w_dff_B_Mu1h62B41_2),.dout(w_dff_B_h48RORwK8_2),.clk(gclk));
	jdff dff_B_M8KCaOh65_2(.din(w_dff_B_h48RORwK8_2),.dout(w_dff_B_M8KCaOh65_2),.clk(gclk));
	jdff dff_B_id2XqKqF6_2(.din(w_dff_B_M8KCaOh65_2),.dout(w_dff_B_id2XqKqF6_2),.clk(gclk));
	jdff dff_B_477vbMIP6_2(.din(w_dff_B_id2XqKqF6_2),.dout(w_dff_B_477vbMIP6_2),.clk(gclk));
	jdff dff_B_YARh4HJy9_2(.din(w_dff_B_477vbMIP6_2),.dout(w_dff_B_YARh4HJy9_2),.clk(gclk));
	jdff dff_B_iaZlrNcx3_2(.din(w_dff_B_YARh4HJy9_2),.dout(w_dff_B_iaZlrNcx3_2),.clk(gclk));
	jdff dff_B_cXwSHk198_2(.din(w_dff_B_iaZlrNcx3_2),.dout(w_dff_B_cXwSHk198_2),.clk(gclk));
	jdff dff_B_RUWyyqcD6_2(.din(w_dff_B_cXwSHk198_2),.dout(w_dff_B_RUWyyqcD6_2),.clk(gclk));
	jdff dff_B_Z0uOcxay9_2(.din(w_dff_B_RUWyyqcD6_2),.dout(w_dff_B_Z0uOcxay9_2),.clk(gclk));
	jdff dff_B_iYnFwR0M6_2(.din(w_dff_B_Z0uOcxay9_2),.dout(w_dff_B_iYnFwR0M6_2),.clk(gclk));
	jdff dff_B_kyLjDg9w9_2(.din(w_dff_B_iYnFwR0M6_2),.dout(w_dff_B_kyLjDg9w9_2),.clk(gclk));
	jdff dff_B_pVeZ9JKP0_2(.din(w_dff_B_kyLjDg9w9_2),.dout(w_dff_B_pVeZ9JKP0_2),.clk(gclk));
	jdff dff_B_LMlpdPGc4_2(.din(w_dff_B_pVeZ9JKP0_2),.dout(w_dff_B_LMlpdPGc4_2),.clk(gclk));
	jdff dff_B_0pEm2brJ7_2(.din(w_dff_B_LMlpdPGc4_2),.dout(w_dff_B_0pEm2brJ7_2),.clk(gclk));
	jdff dff_B_caSTd6PM9_2(.din(w_dff_B_0pEm2brJ7_2),.dout(w_dff_B_caSTd6PM9_2),.clk(gclk));
	jdff dff_B_PePFdTAP5_2(.din(w_dff_B_caSTd6PM9_2),.dout(w_dff_B_PePFdTAP5_2),.clk(gclk));
	jdff dff_B_jsD4HgHt8_2(.din(w_dff_B_PePFdTAP5_2),.dout(w_dff_B_jsD4HgHt8_2),.clk(gclk));
	jdff dff_B_Sg1wUg0H2_2(.din(w_dff_B_jsD4HgHt8_2),.dout(w_dff_B_Sg1wUg0H2_2),.clk(gclk));
	jdff dff_B_yF28aubg9_2(.din(w_dff_B_Sg1wUg0H2_2),.dout(w_dff_B_yF28aubg9_2),.clk(gclk));
	jdff dff_B_tvAuubX99_2(.din(w_dff_B_yF28aubg9_2),.dout(w_dff_B_tvAuubX99_2),.clk(gclk));
	jdff dff_B_4BqsZZHS4_2(.din(w_dff_B_tvAuubX99_2),.dout(w_dff_B_4BqsZZHS4_2),.clk(gclk));
	jdff dff_B_A81Y95J23_2(.din(w_dff_B_4BqsZZHS4_2),.dout(w_dff_B_A81Y95J23_2),.clk(gclk));
	jdff dff_B_kPfcUBLB3_2(.din(w_dff_B_A81Y95J23_2),.dout(w_dff_B_kPfcUBLB3_2),.clk(gclk));
	jdff dff_B_g2enGmPe7_2(.din(w_dff_B_kPfcUBLB3_2),.dout(w_dff_B_g2enGmPe7_2),.clk(gclk));
	jdff dff_B_fZHCOcL76_2(.din(w_dff_B_g2enGmPe7_2),.dout(w_dff_B_fZHCOcL76_2),.clk(gclk));
	jdff dff_B_53SXnkVu4_2(.din(w_dff_B_fZHCOcL76_2),.dout(w_dff_B_53SXnkVu4_2),.clk(gclk));
	jdff dff_B_kCbt8Nyg5_2(.din(w_dff_B_53SXnkVu4_2),.dout(w_dff_B_kCbt8Nyg5_2),.clk(gclk));
	jdff dff_B_fJoq84PA2_2(.din(w_dff_B_kCbt8Nyg5_2),.dout(w_dff_B_fJoq84PA2_2),.clk(gclk));
	jdff dff_B_cRtX1KIi2_2(.din(w_dff_B_fJoq84PA2_2),.dout(w_dff_B_cRtX1KIi2_2),.clk(gclk));
	jdff dff_B_TMcWbaYf7_2(.din(w_dff_B_cRtX1KIi2_2),.dout(w_dff_B_TMcWbaYf7_2),.clk(gclk));
	jdff dff_B_GOyUKeLb9_2(.din(w_dff_B_TMcWbaYf7_2),.dout(w_dff_B_GOyUKeLb9_2),.clk(gclk));
	jdff dff_B_4P83CbSp6_2(.din(w_dff_B_GOyUKeLb9_2),.dout(w_dff_B_4P83CbSp6_2),.clk(gclk));
	jdff dff_B_UhIogdie1_1(.din(n1060),.dout(w_dff_B_UhIogdie1_1),.clk(gclk));
	jdff dff_B_ar28uOhU3_2(.din(n961),.dout(w_dff_B_ar28uOhU3_2),.clk(gclk));
	jdff dff_B_Mbxc45If8_2(.din(w_dff_B_ar28uOhU3_2),.dout(w_dff_B_Mbxc45If8_2),.clk(gclk));
	jdff dff_B_IRIz1hRJ5_2(.din(w_dff_B_Mbxc45If8_2),.dout(w_dff_B_IRIz1hRJ5_2),.clk(gclk));
	jdff dff_B_sAwZzgXI3_2(.din(w_dff_B_IRIz1hRJ5_2),.dout(w_dff_B_sAwZzgXI3_2),.clk(gclk));
	jdff dff_B_Su7aprlm6_2(.din(w_dff_B_sAwZzgXI3_2),.dout(w_dff_B_Su7aprlm6_2),.clk(gclk));
	jdff dff_B_0uBCu5Mm2_2(.din(w_dff_B_Su7aprlm6_2),.dout(w_dff_B_0uBCu5Mm2_2),.clk(gclk));
	jdff dff_B_zevdaLSW5_2(.din(w_dff_B_0uBCu5Mm2_2),.dout(w_dff_B_zevdaLSW5_2),.clk(gclk));
	jdff dff_B_Q7unzoo97_2(.din(w_dff_B_zevdaLSW5_2),.dout(w_dff_B_Q7unzoo97_2),.clk(gclk));
	jdff dff_B_mjsYeI5S9_2(.din(w_dff_B_Q7unzoo97_2),.dout(w_dff_B_mjsYeI5S9_2),.clk(gclk));
	jdff dff_B_3un0WgMB5_2(.din(w_dff_B_mjsYeI5S9_2),.dout(w_dff_B_3un0WgMB5_2),.clk(gclk));
	jdff dff_B_J0Da3LgN1_2(.din(w_dff_B_3un0WgMB5_2),.dout(w_dff_B_J0Da3LgN1_2),.clk(gclk));
	jdff dff_B_u054pjDB7_2(.din(w_dff_B_J0Da3LgN1_2),.dout(w_dff_B_u054pjDB7_2),.clk(gclk));
	jdff dff_B_k3aJothM2_2(.din(w_dff_B_u054pjDB7_2),.dout(w_dff_B_k3aJothM2_2),.clk(gclk));
	jdff dff_B_C2ncuhDq0_2(.din(w_dff_B_k3aJothM2_2),.dout(w_dff_B_C2ncuhDq0_2),.clk(gclk));
	jdff dff_B_U3SgzjHC2_2(.din(w_dff_B_C2ncuhDq0_2),.dout(w_dff_B_U3SgzjHC2_2),.clk(gclk));
	jdff dff_B_Fuqn5Uxb5_2(.din(w_dff_B_U3SgzjHC2_2),.dout(w_dff_B_Fuqn5Uxb5_2),.clk(gclk));
	jdff dff_B_4jyMa10R5_2(.din(w_dff_B_Fuqn5Uxb5_2),.dout(w_dff_B_4jyMa10R5_2),.clk(gclk));
	jdff dff_B_coKJHB6e8_2(.din(w_dff_B_4jyMa10R5_2),.dout(w_dff_B_coKJHB6e8_2),.clk(gclk));
	jdff dff_B_rmaE43Yd5_2(.din(w_dff_B_coKJHB6e8_2),.dout(w_dff_B_rmaE43Yd5_2),.clk(gclk));
	jdff dff_B_j4sQzHwf7_2(.din(w_dff_B_rmaE43Yd5_2),.dout(w_dff_B_j4sQzHwf7_2),.clk(gclk));
	jdff dff_B_dN0cZSOu0_2(.din(w_dff_B_j4sQzHwf7_2),.dout(w_dff_B_dN0cZSOu0_2),.clk(gclk));
	jdff dff_B_UaO0raDX3_2(.din(w_dff_B_dN0cZSOu0_2),.dout(w_dff_B_UaO0raDX3_2),.clk(gclk));
	jdff dff_B_zAux4gZk5_2(.din(w_dff_B_UaO0raDX3_2),.dout(w_dff_B_zAux4gZk5_2),.clk(gclk));
	jdff dff_B_lKn1YUqf5_2(.din(w_dff_B_zAux4gZk5_2),.dout(w_dff_B_lKn1YUqf5_2),.clk(gclk));
	jdff dff_B_386CQtn60_2(.din(w_dff_B_lKn1YUqf5_2),.dout(w_dff_B_386CQtn60_2),.clk(gclk));
	jdff dff_B_rpCfMSGh8_2(.din(w_dff_B_386CQtn60_2),.dout(w_dff_B_rpCfMSGh8_2),.clk(gclk));
	jdff dff_B_Sivw5WCI8_2(.din(w_dff_B_rpCfMSGh8_2),.dout(w_dff_B_Sivw5WCI8_2),.clk(gclk));
	jdff dff_B_h1mTn8qL8_2(.din(w_dff_B_Sivw5WCI8_2),.dout(w_dff_B_h1mTn8qL8_2),.clk(gclk));
	jdff dff_B_zQTzwlJ39_2(.din(w_dff_B_h1mTn8qL8_2),.dout(w_dff_B_zQTzwlJ39_2),.clk(gclk));
	jdff dff_B_wHbRWiRb4_2(.din(w_dff_B_zQTzwlJ39_2),.dout(w_dff_B_wHbRWiRb4_2),.clk(gclk));
	jdff dff_B_eSqY2FEm1_2(.din(w_dff_B_wHbRWiRb4_2),.dout(w_dff_B_eSqY2FEm1_2),.clk(gclk));
	jdff dff_B_Ty6trjOr3_1(.din(n962),.dout(w_dff_B_Ty6trjOr3_1),.clk(gclk));
	jdff dff_B_zyptDpkY2_2(.din(n856),.dout(w_dff_B_zyptDpkY2_2),.clk(gclk));
	jdff dff_B_y4Ube5an2_2(.din(w_dff_B_zyptDpkY2_2),.dout(w_dff_B_y4Ube5an2_2),.clk(gclk));
	jdff dff_B_I4zNbDoI3_2(.din(w_dff_B_y4Ube5an2_2),.dout(w_dff_B_I4zNbDoI3_2),.clk(gclk));
	jdff dff_B_iC6EmDSr4_2(.din(w_dff_B_I4zNbDoI3_2),.dout(w_dff_B_iC6EmDSr4_2),.clk(gclk));
	jdff dff_B_MrZ7h7iX8_2(.din(w_dff_B_iC6EmDSr4_2),.dout(w_dff_B_MrZ7h7iX8_2),.clk(gclk));
	jdff dff_B_9C48Tz4M7_2(.din(w_dff_B_MrZ7h7iX8_2),.dout(w_dff_B_9C48Tz4M7_2),.clk(gclk));
	jdff dff_B_eY43w6qp7_2(.din(w_dff_B_9C48Tz4M7_2),.dout(w_dff_B_eY43w6qp7_2),.clk(gclk));
	jdff dff_B_94bRS6Zc3_2(.din(w_dff_B_eY43w6qp7_2),.dout(w_dff_B_94bRS6Zc3_2),.clk(gclk));
	jdff dff_B_MnxwYbbG6_2(.din(w_dff_B_94bRS6Zc3_2),.dout(w_dff_B_MnxwYbbG6_2),.clk(gclk));
	jdff dff_B_FcPa4WaH5_2(.din(w_dff_B_MnxwYbbG6_2),.dout(w_dff_B_FcPa4WaH5_2),.clk(gclk));
	jdff dff_B_yTvnrMGf7_2(.din(w_dff_B_FcPa4WaH5_2),.dout(w_dff_B_yTvnrMGf7_2),.clk(gclk));
	jdff dff_B_tmnxWpXx3_2(.din(w_dff_B_yTvnrMGf7_2),.dout(w_dff_B_tmnxWpXx3_2),.clk(gclk));
	jdff dff_B_mP67yWkI7_2(.din(w_dff_B_tmnxWpXx3_2),.dout(w_dff_B_mP67yWkI7_2),.clk(gclk));
	jdff dff_B_ZVEW2Wgg7_2(.din(w_dff_B_mP67yWkI7_2),.dout(w_dff_B_ZVEW2Wgg7_2),.clk(gclk));
	jdff dff_B_jEqc3vX75_2(.din(w_dff_B_ZVEW2Wgg7_2),.dout(w_dff_B_jEqc3vX75_2),.clk(gclk));
	jdff dff_B_meSBabrK2_2(.din(w_dff_B_jEqc3vX75_2),.dout(w_dff_B_meSBabrK2_2),.clk(gclk));
	jdff dff_B_js3dBYcS8_2(.din(w_dff_B_meSBabrK2_2),.dout(w_dff_B_js3dBYcS8_2),.clk(gclk));
	jdff dff_B_BNKNvkt61_2(.din(w_dff_B_js3dBYcS8_2),.dout(w_dff_B_BNKNvkt61_2),.clk(gclk));
	jdff dff_B_0xtg43hz4_2(.din(w_dff_B_BNKNvkt61_2),.dout(w_dff_B_0xtg43hz4_2),.clk(gclk));
	jdff dff_B_lgd5mQvA2_2(.din(w_dff_B_0xtg43hz4_2),.dout(w_dff_B_lgd5mQvA2_2),.clk(gclk));
	jdff dff_B_sCW2FjgQ1_2(.din(w_dff_B_lgd5mQvA2_2),.dout(w_dff_B_sCW2FjgQ1_2),.clk(gclk));
	jdff dff_B_hMKtJyxY7_2(.din(w_dff_B_sCW2FjgQ1_2),.dout(w_dff_B_hMKtJyxY7_2),.clk(gclk));
	jdff dff_B_SgOIII2a1_2(.din(w_dff_B_hMKtJyxY7_2),.dout(w_dff_B_SgOIII2a1_2),.clk(gclk));
	jdff dff_B_LwYy6BIU8_2(.din(w_dff_B_SgOIII2a1_2),.dout(w_dff_B_LwYy6BIU8_2),.clk(gclk));
	jdff dff_B_NdHpaAPw4_2(.din(w_dff_B_LwYy6BIU8_2),.dout(w_dff_B_NdHpaAPw4_2),.clk(gclk));
	jdff dff_B_na7o3CWK8_2(.din(w_dff_B_NdHpaAPw4_2),.dout(w_dff_B_na7o3CWK8_2),.clk(gclk));
	jdff dff_B_o4fmtzml8_2(.din(w_dff_B_na7o3CWK8_2),.dout(w_dff_B_o4fmtzml8_2),.clk(gclk));
	jdff dff_B_j1yGSPFY8_2(.din(w_dff_B_o4fmtzml8_2),.dout(w_dff_B_j1yGSPFY8_2),.clk(gclk));
	jdff dff_B_aOKnKsbI5_1(.din(n857),.dout(w_dff_B_aOKnKsbI5_1),.clk(gclk));
	jdff dff_B_t8WFISp08_2(.din(n757),.dout(w_dff_B_t8WFISp08_2),.clk(gclk));
	jdff dff_B_44nP9i2V4_2(.din(w_dff_B_t8WFISp08_2),.dout(w_dff_B_44nP9i2V4_2),.clk(gclk));
	jdff dff_B_5bAK6Yg66_2(.din(w_dff_B_44nP9i2V4_2),.dout(w_dff_B_5bAK6Yg66_2),.clk(gclk));
	jdff dff_B_wihg9dZv6_2(.din(w_dff_B_5bAK6Yg66_2),.dout(w_dff_B_wihg9dZv6_2),.clk(gclk));
	jdff dff_B_y7sptAQY7_2(.din(w_dff_B_wihg9dZv6_2),.dout(w_dff_B_y7sptAQY7_2),.clk(gclk));
	jdff dff_B_r347IwI28_2(.din(w_dff_B_y7sptAQY7_2),.dout(w_dff_B_r347IwI28_2),.clk(gclk));
	jdff dff_B_OyhCjVUy9_2(.din(w_dff_B_r347IwI28_2),.dout(w_dff_B_OyhCjVUy9_2),.clk(gclk));
	jdff dff_B_Ab5EYeQs5_2(.din(w_dff_B_OyhCjVUy9_2),.dout(w_dff_B_Ab5EYeQs5_2),.clk(gclk));
	jdff dff_B_5E4cWV1U8_2(.din(w_dff_B_Ab5EYeQs5_2),.dout(w_dff_B_5E4cWV1U8_2),.clk(gclk));
	jdff dff_B_usSTADm85_2(.din(w_dff_B_5E4cWV1U8_2),.dout(w_dff_B_usSTADm85_2),.clk(gclk));
	jdff dff_B_C9OMeGqX5_2(.din(w_dff_B_usSTADm85_2),.dout(w_dff_B_C9OMeGqX5_2),.clk(gclk));
	jdff dff_B_EVQJ2NAe5_2(.din(w_dff_B_C9OMeGqX5_2),.dout(w_dff_B_EVQJ2NAe5_2),.clk(gclk));
	jdff dff_B_zaFgKXCb5_2(.din(w_dff_B_EVQJ2NAe5_2),.dout(w_dff_B_zaFgKXCb5_2),.clk(gclk));
	jdff dff_B_B9iZeQ1Q6_2(.din(w_dff_B_zaFgKXCb5_2),.dout(w_dff_B_B9iZeQ1Q6_2),.clk(gclk));
	jdff dff_B_76jpFiPs1_2(.din(w_dff_B_B9iZeQ1Q6_2),.dout(w_dff_B_76jpFiPs1_2),.clk(gclk));
	jdff dff_B_GMAX2RNd1_2(.din(w_dff_B_76jpFiPs1_2),.dout(w_dff_B_GMAX2RNd1_2),.clk(gclk));
	jdff dff_B_oYUp9omq1_2(.din(w_dff_B_GMAX2RNd1_2),.dout(w_dff_B_oYUp9omq1_2),.clk(gclk));
	jdff dff_B_qFhHMkon7_2(.din(w_dff_B_oYUp9omq1_2),.dout(w_dff_B_qFhHMkon7_2),.clk(gclk));
	jdff dff_B_o3ablrzL1_2(.din(w_dff_B_qFhHMkon7_2),.dout(w_dff_B_o3ablrzL1_2),.clk(gclk));
	jdff dff_B_UQv29VuB1_2(.din(w_dff_B_o3ablrzL1_2),.dout(w_dff_B_UQv29VuB1_2),.clk(gclk));
	jdff dff_B_M7jLzGgz1_2(.din(w_dff_B_UQv29VuB1_2),.dout(w_dff_B_M7jLzGgz1_2),.clk(gclk));
	jdff dff_B_PwLVjtrM8_2(.din(w_dff_B_M7jLzGgz1_2),.dout(w_dff_B_PwLVjtrM8_2),.clk(gclk));
	jdff dff_B_KYXnVwUT0_2(.din(w_dff_B_PwLVjtrM8_2),.dout(w_dff_B_KYXnVwUT0_2),.clk(gclk));
	jdff dff_B_kmKD18UZ3_2(.din(w_dff_B_KYXnVwUT0_2),.dout(w_dff_B_kmKD18UZ3_2),.clk(gclk));
	jdff dff_B_zR9qlZKD4_2(.din(w_dff_B_kmKD18UZ3_2),.dout(w_dff_B_zR9qlZKD4_2),.clk(gclk));
	jdff dff_B_F4vP9F4i6_1(.din(n758),.dout(w_dff_B_F4vP9F4i6_1),.clk(gclk));
	jdff dff_B_1p18hD567_2(.din(n664),.dout(w_dff_B_1p18hD567_2),.clk(gclk));
	jdff dff_B_MLapcce12_2(.din(w_dff_B_1p18hD567_2),.dout(w_dff_B_MLapcce12_2),.clk(gclk));
	jdff dff_B_EBSLFvWC5_2(.din(w_dff_B_MLapcce12_2),.dout(w_dff_B_EBSLFvWC5_2),.clk(gclk));
	jdff dff_B_APz24RGh2_2(.din(w_dff_B_EBSLFvWC5_2),.dout(w_dff_B_APz24RGh2_2),.clk(gclk));
	jdff dff_B_6mYl2Ci25_2(.din(w_dff_B_APz24RGh2_2),.dout(w_dff_B_6mYl2Ci25_2),.clk(gclk));
	jdff dff_B_AKhJBG480_2(.din(w_dff_B_6mYl2Ci25_2),.dout(w_dff_B_AKhJBG480_2),.clk(gclk));
	jdff dff_B_5i0imjQS0_2(.din(w_dff_B_AKhJBG480_2),.dout(w_dff_B_5i0imjQS0_2),.clk(gclk));
	jdff dff_B_NUXUo0vc7_2(.din(w_dff_B_5i0imjQS0_2),.dout(w_dff_B_NUXUo0vc7_2),.clk(gclk));
	jdff dff_B_spQShVNE1_2(.din(w_dff_B_NUXUo0vc7_2),.dout(w_dff_B_spQShVNE1_2),.clk(gclk));
	jdff dff_B_EQeg9lbJ2_2(.din(w_dff_B_spQShVNE1_2),.dout(w_dff_B_EQeg9lbJ2_2),.clk(gclk));
	jdff dff_B_tLQFADPr9_2(.din(w_dff_B_EQeg9lbJ2_2),.dout(w_dff_B_tLQFADPr9_2),.clk(gclk));
	jdff dff_B_EP7XPJMF7_2(.din(w_dff_B_tLQFADPr9_2),.dout(w_dff_B_EP7XPJMF7_2),.clk(gclk));
	jdff dff_B_l5VjWV6J7_2(.din(w_dff_B_EP7XPJMF7_2),.dout(w_dff_B_l5VjWV6J7_2),.clk(gclk));
	jdff dff_B_EhiQJxor2_2(.din(w_dff_B_l5VjWV6J7_2),.dout(w_dff_B_EhiQJxor2_2),.clk(gclk));
	jdff dff_B_HoUupqzo8_2(.din(w_dff_B_EhiQJxor2_2),.dout(w_dff_B_HoUupqzo8_2),.clk(gclk));
	jdff dff_B_8xTQIdKM1_2(.din(w_dff_B_HoUupqzo8_2),.dout(w_dff_B_8xTQIdKM1_2),.clk(gclk));
	jdff dff_B_eXlfqz2o1_2(.din(w_dff_B_8xTQIdKM1_2),.dout(w_dff_B_eXlfqz2o1_2),.clk(gclk));
	jdff dff_B_FRfXUKr84_2(.din(w_dff_B_eXlfqz2o1_2),.dout(w_dff_B_FRfXUKr84_2),.clk(gclk));
	jdff dff_B_9KiotzSZ4_2(.din(w_dff_B_FRfXUKr84_2),.dout(w_dff_B_9KiotzSZ4_2),.clk(gclk));
	jdff dff_B_W62zzIzD4_2(.din(w_dff_B_9KiotzSZ4_2),.dout(w_dff_B_W62zzIzD4_2),.clk(gclk));
	jdff dff_B_3KK4QQkq5_2(.din(w_dff_B_W62zzIzD4_2),.dout(w_dff_B_3KK4QQkq5_2),.clk(gclk));
	jdff dff_B_QpjVlIc90_2(.din(w_dff_B_3KK4QQkq5_2),.dout(w_dff_B_QpjVlIc90_2),.clk(gclk));
	jdff dff_B_9M5pmyQ40_1(.din(n665),.dout(w_dff_B_9M5pmyQ40_1),.clk(gclk));
	jdff dff_B_3Oy4zAc83_2(.din(n578),.dout(w_dff_B_3Oy4zAc83_2),.clk(gclk));
	jdff dff_B_RbVCnQe98_2(.din(w_dff_B_3Oy4zAc83_2),.dout(w_dff_B_RbVCnQe98_2),.clk(gclk));
	jdff dff_B_1pczOuZR7_2(.din(w_dff_B_RbVCnQe98_2),.dout(w_dff_B_1pczOuZR7_2),.clk(gclk));
	jdff dff_B_6yB0xafJ0_2(.din(w_dff_B_1pczOuZR7_2),.dout(w_dff_B_6yB0xafJ0_2),.clk(gclk));
	jdff dff_B_SuSjQcXD1_2(.din(w_dff_B_6yB0xafJ0_2),.dout(w_dff_B_SuSjQcXD1_2),.clk(gclk));
	jdff dff_B_DxiDnaAc5_2(.din(w_dff_B_SuSjQcXD1_2),.dout(w_dff_B_DxiDnaAc5_2),.clk(gclk));
	jdff dff_B_qiywJnVB2_2(.din(w_dff_B_DxiDnaAc5_2),.dout(w_dff_B_qiywJnVB2_2),.clk(gclk));
	jdff dff_B_WVtFyks58_2(.din(w_dff_B_qiywJnVB2_2),.dout(w_dff_B_WVtFyks58_2),.clk(gclk));
	jdff dff_B_16hPDcOk3_2(.din(w_dff_B_WVtFyks58_2),.dout(w_dff_B_16hPDcOk3_2),.clk(gclk));
	jdff dff_B_GIDQdYSE8_2(.din(w_dff_B_16hPDcOk3_2),.dout(w_dff_B_GIDQdYSE8_2),.clk(gclk));
	jdff dff_B_hjY8zbRe0_2(.din(w_dff_B_GIDQdYSE8_2),.dout(w_dff_B_hjY8zbRe0_2),.clk(gclk));
	jdff dff_B_flV9nWky7_2(.din(w_dff_B_hjY8zbRe0_2),.dout(w_dff_B_flV9nWky7_2),.clk(gclk));
	jdff dff_B_f6MA30B28_2(.din(w_dff_B_flV9nWky7_2),.dout(w_dff_B_f6MA30B28_2),.clk(gclk));
	jdff dff_B_rtRNaiLF9_2(.din(w_dff_B_f6MA30B28_2),.dout(w_dff_B_rtRNaiLF9_2),.clk(gclk));
	jdff dff_B_Weew9LTl7_2(.din(w_dff_B_rtRNaiLF9_2),.dout(w_dff_B_Weew9LTl7_2),.clk(gclk));
	jdff dff_B_sPbCZpbO2_2(.din(w_dff_B_Weew9LTl7_2),.dout(w_dff_B_sPbCZpbO2_2),.clk(gclk));
	jdff dff_B_UX0a4oAJ7_2(.din(w_dff_B_sPbCZpbO2_2),.dout(w_dff_B_UX0a4oAJ7_2),.clk(gclk));
	jdff dff_B_ifbYKzyJ1_2(.din(w_dff_B_UX0a4oAJ7_2),.dout(w_dff_B_ifbYKzyJ1_2),.clk(gclk));
	jdff dff_B_qqduDE2g4_2(.din(w_dff_B_ifbYKzyJ1_2),.dout(w_dff_B_qqduDE2g4_2),.clk(gclk));
	jdff dff_B_s9Cd84hT8_1(.din(n579),.dout(w_dff_B_s9Cd84hT8_1),.clk(gclk));
	jdff dff_B_ZSz19q7P4_2(.din(n499),.dout(w_dff_B_ZSz19q7P4_2),.clk(gclk));
	jdff dff_B_Lq2hAwIk1_2(.din(w_dff_B_ZSz19q7P4_2),.dout(w_dff_B_Lq2hAwIk1_2),.clk(gclk));
	jdff dff_B_R58AkyAS8_2(.din(w_dff_B_Lq2hAwIk1_2),.dout(w_dff_B_R58AkyAS8_2),.clk(gclk));
	jdff dff_B_2bS28fJ98_2(.din(w_dff_B_R58AkyAS8_2),.dout(w_dff_B_2bS28fJ98_2),.clk(gclk));
	jdff dff_B_X2Svo9sr2_2(.din(w_dff_B_2bS28fJ98_2),.dout(w_dff_B_X2Svo9sr2_2),.clk(gclk));
	jdff dff_B_JEo17NHy5_2(.din(w_dff_B_X2Svo9sr2_2),.dout(w_dff_B_JEo17NHy5_2),.clk(gclk));
	jdff dff_B_SgkybFcA6_2(.din(w_dff_B_JEo17NHy5_2),.dout(w_dff_B_SgkybFcA6_2),.clk(gclk));
	jdff dff_B_LY8odb8R5_2(.din(w_dff_B_SgkybFcA6_2),.dout(w_dff_B_LY8odb8R5_2),.clk(gclk));
	jdff dff_B_rVpjdAN79_2(.din(w_dff_B_LY8odb8R5_2),.dout(w_dff_B_rVpjdAN79_2),.clk(gclk));
	jdff dff_B_lyJmV2WD3_2(.din(w_dff_B_rVpjdAN79_2),.dout(w_dff_B_lyJmV2WD3_2),.clk(gclk));
	jdff dff_B_yUNS7d8j9_2(.din(w_dff_B_lyJmV2WD3_2),.dout(w_dff_B_yUNS7d8j9_2),.clk(gclk));
	jdff dff_B_So8gVGsf1_2(.din(w_dff_B_yUNS7d8j9_2),.dout(w_dff_B_So8gVGsf1_2),.clk(gclk));
	jdff dff_B_E31YnTJc1_2(.din(w_dff_B_So8gVGsf1_2),.dout(w_dff_B_E31YnTJc1_2),.clk(gclk));
	jdff dff_B_SeWOF00b6_2(.din(w_dff_B_E31YnTJc1_2),.dout(w_dff_B_SeWOF00b6_2),.clk(gclk));
	jdff dff_B_1g9pyNQd0_2(.din(w_dff_B_SeWOF00b6_2),.dout(w_dff_B_1g9pyNQd0_2),.clk(gclk));
	jdff dff_B_1WJwsVqu8_2(.din(w_dff_B_1g9pyNQd0_2),.dout(w_dff_B_1WJwsVqu8_2),.clk(gclk));
	jdff dff_B_qAkQqxEW1_1(.din(n500),.dout(w_dff_B_qAkQqxEW1_1),.clk(gclk));
	jdff dff_B_DRRdmiDW3_2(.din(n427),.dout(w_dff_B_DRRdmiDW3_2),.clk(gclk));
	jdff dff_B_urIvva7L5_2(.din(w_dff_B_DRRdmiDW3_2),.dout(w_dff_B_urIvva7L5_2),.clk(gclk));
	jdff dff_B_MuWDCOfI2_2(.din(w_dff_B_urIvva7L5_2),.dout(w_dff_B_MuWDCOfI2_2),.clk(gclk));
	jdff dff_B_IKxz5faF8_2(.din(w_dff_B_MuWDCOfI2_2),.dout(w_dff_B_IKxz5faF8_2),.clk(gclk));
	jdff dff_B_MUQ3CgdL6_2(.din(w_dff_B_IKxz5faF8_2),.dout(w_dff_B_MUQ3CgdL6_2),.clk(gclk));
	jdff dff_B_atjKpGNi7_2(.din(w_dff_B_MUQ3CgdL6_2),.dout(w_dff_B_atjKpGNi7_2),.clk(gclk));
	jdff dff_B_OXNf1yG70_2(.din(w_dff_B_atjKpGNi7_2),.dout(w_dff_B_OXNf1yG70_2),.clk(gclk));
	jdff dff_B_1UWUrrwO9_2(.din(w_dff_B_OXNf1yG70_2),.dout(w_dff_B_1UWUrrwO9_2),.clk(gclk));
	jdff dff_B_qce8hfQB1_2(.din(w_dff_B_1UWUrrwO9_2),.dout(w_dff_B_qce8hfQB1_2),.clk(gclk));
	jdff dff_B_mGHPOroW1_2(.din(w_dff_B_qce8hfQB1_2),.dout(w_dff_B_mGHPOroW1_2),.clk(gclk));
	jdff dff_B_mHDzVxhK5_2(.din(w_dff_B_mGHPOroW1_2),.dout(w_dff_B_mHDzVxhK5_2),.clk(gclk));
	jdff dff_B_Vu6i6Fll3_2(.din(w_dff_B_mHDzVxhK5_2),.dout(w_dff_B_Vu6i6Fll3_2),.clk(gclk));
	jdff dff_B_WVEh5NPZ2_2(.din(w_dff_B_Vu6i6Fll3_2),.dout(w_dff_B_WVEh5NPZ2_2),.clk(gclk));
	jdff dff_B_BnZj7UBm8_1(.din(n428),.dout(w_dff_B_BnZj7UBm8_1),.clk(gclk));
	jdff dff_B_4QyvSVSR8_2(.din(n363),.dout(w_dff_B_4QyvSVSR8_2),.clk(gclk));
	jdff dff_B_IIx56gXe0_2(.din(w_dff_B_4QyvSVSR8_2),.dout(w_dff_B_IIx56gXe0_2),.clk(gclk));
	jdff dff_B_6wZH7Ok81_2(.din(w_dff_B_IIx56gXe0_2),.dout(w_dff_B_6wZH7Ok81_2),.clk(gclk));
	jdff dff_B_gkNvJvQH7_2(.din(w_dff_B_6wZH7Ok81_2),.dout(w_dff_B_gkNvJvQH7_2),.clk(gclk));
	jdff dff_B_PUvLPEbX8_2(.din(w_dff_B_gkNvJvQH7_2),.dout(w_dff_B_PUvLPEbX8_2),.clk(gclk));
	jdff dff_B_613AM2O79_2(.din(w_dff_B_PUvLPEbX8_2),.dout(w_dff_B_613AM2O79_2),.clk(gclk));
	jdff dff_B_xrCZWvcG0_2(.din(w_dff_B_613AM2O79_2),.dout(w_dff_B_xrCZWvcG0_2),.clk(gclk));
	jdff dff_B_ly6g3P1U1_2(.din(w_dff_B_xrCZWvcG0_2),.dout(w_dff_B_ly6g3P1U1_2),.clk(gclk));
	jdff dff_B_QaJT2DOY0_2(.din(w_dff_B_ly6g3P1U1_2),.dout(w_dff_B_QaJT2DOY0_2),.clk(gclk));
	jdff dff_B_wVO3rB1a0_2(.din(w_dff_B_QaJT2DOY0_2),.dout(w_dff_B_wVO3rB1a0_2),.clk(gclk));
	jdff dff_B_OOIwGHPY4_2(.din(n385),.dout(w_dff_B_OOIwGHPY4_2),.clk(gclk));
	jdff dff_B_TK43nvRb3_1(.din(n364),.dout(w_dff_B_TK43nvRb3_1),.clk(gclk));
	jdff dff_B_L7G2pKg59_2(.din(n305),.dout(w_dff_B_L7G2pKg59_2),.clk(gclk));
	jdff dff_B_0KwACUyX9_2(.din(w_dff_B_L7G2pKg59_2),.dout(w_dff_B_0KwACUyX9_2),.clk(gclk));
	jdff dff_B_kIK5WVBH9_2(.din(w_dff_B_0KwACUyX9_2),.dout(w_dff_B_kIK5WVBH9_2),.clk(gclk));
	jdff dff_B_8YKbz1RU8_2(.din(w_dff_B_kIK5WVBH9_2),.dout(w_dff_B_8YKbz1RU8_2),.clk(gclk));
	jdff dff_B_F5ySW75Y5_2(.din(w_dff_B_8YKbz1RU8_2),.dout(w_dff_B_F5ySW75Y5_2),.clk(gclk));
	jdff dff_B_ffnSJ3H53_2(.din(w_dff_B_F5ySW75Y5_2),.dout(w_dff_B_ffnSJ3H53_2),.clk(gclk));
	jdff dff_B_JqLKAmu29_2(.din(w_dff_B_ffnSJ3H53_2),.dout(w_dff_B_JqLKAmu29_2),.clk(gclk));
	jdff dff_B_NxEO5AfJ9_2(.din(n321),.dout(w_dff_B_NxEO5AfJ9_2),.clk(gclk));
	jdff dff_B_p983pDwu3_1(.din(n306),.dout(w_dff_B_p983pDwu3_1),.clk(gclk));
	jdff dff_B_Lj5YMUYh5_2(.din(n254),.dout(w_dff_B_Lj5YMUYh5_2),.clk(gclk));
	jdff dff_B_xBmmamQh7_2(.din(w_dff_B_Lj5YMUYh5_2),.dout(w_dff_B_xBmmamQh7_2),.clk(gclk));
	jdff dff_B_JlmFxbUl8_2(.din(w_dff_B_xBmmamQh7_2),.dout(w_dff_B_JlmFxbUl8_2),.clk(gclk));
	jdff dff_B_Cjc6iVEW9_2(.din(w_dff_B_JlmFxbUl8_2),.dout(w_dff_B_Cjc6iVEW9_2),.clk(gclk));
	jdff dff_B_9IuVKnvE7_1(.din(n256),.dout(w_dff_B_9IuVKnvE7_1),.clk(gclk));
	jdff dff_A_pnxRAwe47_1(.dout(w_n210_0[1]),.din(w_dff_A_pnxRAwe47_1),.clk(gclk));
	jdff dff_A_bReyMFdL4_2(.dout(w_n210_0[2]),.din(w_dff_A_bReyMFdL4_2),.clk(gclk));
	jdff dff_A_MHJ6KRGP1_2(.dout(w_dff_A_bReyMFdL4_2),.din(w_dff_A_MHJ6KRGP1_2),.clk(gclk));
	jdff dff_B_1PbYWcAW4_2(.din(n1496),.dout(w_dff_B_1PbYWcAW4_2),.clk(gclk));
	jdff dff_B_RRuD0sth9_1(.din(n1494),.dout(w_dff_B_RRuD0sth9_1),.clk(gclk));
	jdff dff_B_phbo0j6D0_2(.din(n1421),.dout(w_dff_B_phbo0j6D0_2),.clk(gclk));
	jdff dff_B_8YVilGzq5_2(.din(w_dff_B_phbo0j6D0_2),.dout(w_dff_B_8YVilGzq5_2),.clk(gclk));
	jdff dff_B_BmzU59om7_2(.din(w_dff_B_8YVilGzq5_2),.dout(w_dff_B_BmzU59om7_2),.clk(gclk));
	jdff dff_B_YVIktdGg6_2(.din(w_dff_B_BmzU59om7_2),.dout(w_dff_B_YVIktdGg6_2),.clk(gclk));
	jdff dff_B_8ydDYcP81_2(.din(w_dff_B_YVIktdGg6_2),.dout(w_dff_B_8ydDYcP81_2),.clk(gclk));
	jdff dff_B_OQgfeYhR3_2(.din(w_dff_B_8ydDYcP81_2),.dout(w_dff_B_OQgfeYhR3_2),.clk(gclk));
	jdff dff_B_G11Lskv29_2(.din(w_dff_B_OQgfeYhR3_2),.dout(w_dff_B_G11Lskv29_2),.clk(gclk));
	jdff dff_B_CQCWSLBS8_2(.din(w_dff_B_G11Lskv29_2),.dout(w_dff_B_CQCWSLBS8_2),.clk(gclk));
	jdff dff_B_sUEr4TXq0_2(.din(w_dff_B_CQCWSLBS8_2),.dout(w_dff_B_sUEr4TXq0_2),.clk(gclk));
	jdff dff_B_7MbSH3721_2(.din(w_dff_B_sUEr4TXq0_2),.dout(w_dff_B_7MbSH3721_2),.clk(gclk));
	jdff dff_B_SePz8io24_2(.din(w_dff_B_7MbSH3721_2),.dout(w_dff_B_SePz8io24_2),.clk(gclk));
	jdff dff_B_NGQ8Tdl15_2(.din(w_dff_B_SePz8io24_2),.dout(w_dff_B_NGQ8Tdl15_2),.clk(gclk));
	jdff dff_B_lt75ed062_2(.din(w_dff_B_NGQ8Tdl15_2),.dout(w_dff_B_lt75ed062_2),.clk(gclk));
	jdff dff_B_VWqlhZly4_2(.din(w_dff_B_lt75ed062_2),.dout(w_dff_B_VWqlhZly4_2),.clk(gclk));
	jdff dff_B_ntIG5aVD8_2(.din(w_dff_B_VWqlhZly4_2),.dout(w_dff_B_ntIG5aVD8_2),.clk(gclk));
	jdff dff_B_W8LSHsh81_2(.din(w_dff_B_ntIG5aVD8_2),.dout(w_dff_B_W8LSHsh81_2),.clk(gclk));
	jdff dff_B_tSTUgfPQ8_2(.din(w_dff_B_W8LSHsh81_2),.dout(w_dff_B_tSTUgfPQ8_2),.clk(gclk));
	jdff dff_B_upkqrRwu6_2(.din(w_dff_B_tSTUgfPQ8_2),.dout(w_dff_B_upkqrRwu6_2),.clk(gclk));
	jdff dff_B_jy1WydnB1_2(.din(w_dff_B_upkqrRwu6_2),.dout(w_dff_B_jy1WydnB1_2),.clk(gclk));
	jdff dff_B_ohhgsH8T8_2(.din(w_dff_B_jy1WydnB1_2),.dout(w_dff_B_ohhgsH8T8_2),.clk(gclk));
	jdff dff_B_stsMYuIm9_2(.din(w_dff_B_ohhgsH8T8_2),.dout(w_dff_B_stsMYuIm9_2),.clk(gclk));
	jdff dff_B_U1tVEron5_2(.din(w_dff_B_stsMYuIm9_2),.dout(w_dff_B_U1tVEron5_2),.clk(gclk));
	jdff dff_B_ZiUT98Jd3_2(.din(w_dff_B_U1tVEron5_2),.dout(w_dff_B_ZiUT98Jd3_2),.clk(gclk));
	jdff dff_B_LaBPyo2r3_2(.din(w_dff_B_ZiUT98Jd3_2),.dout(w_dff_B_LaBPyo2r3_2),.clk(gclk));
	jdff dff_B_GkAN6Om21_2(.din(w_dff_B_LaBPyo2r3_2),.dout(w_dff_B_GkAN6Om21_2),.clk(gclk));
	jdff dff_B_tejtAvzC6_2(.din(w_dff_B_GkAN6Om21_2),.dout(w_dff_B_tejtAvzC6_2),.clk(gclk));
	jdff dff_B_cVencumn7_2(.din(w_dff_B_tejtAvzC6_2),.dout(w_dff_B_cVencumn7_2),.clk(gclk));
	jdff dff_B_IpnrKMFN1_2(.din(w_dff_B_cVencumn7_2),.dout(w_dff_B_IpnrKMFN1_2),.clk(gclk));
	jdff dff_B_LjnXAPnO4_2(.din(w_dff_B_IpnrKMFN1_2),.dout(w_dff_B_LjnXAPnO4_2),.clk(gclk));
	jdff dff_B_INSiJQO72_2(.din(w_dff_B_LjnXAPnO4_2),.dout(w_dff_B_INSiJQO72_2),.clk(gclk));
	jdff dff_B_hKsAMLUP0_2(.din(w_dff_B_INSiJQO72_2),.dout(w_dff_B_hKsAMLUP0_2),.clk(gclk));
	jdff dff_B_oEVqmzXk3_2(.din(w_dff_B_hKsAMLUP0_2),.dout(w_dff_B_oEVqmzXk3_2),.clk(gclk));
	jdff dff_B_684SEqpv1_2(.din(w_dff_B_oEVqmzXk3_2),.dout(w_dff_B_684SEqpv1_2),.clk(gclk));
	jdff dff_B_SZaKRMyP0_2(.din(w_dff_B_684SEqpv1_2),.dout(w_dff_B_SZaKRMyP0_2),.clk(gclk));
	jdff dff_B_b7TOsfdU2_2(.din(w_dff_B_SZaKRMyP0_2),.dout(w_dff_B_b7TOsfdU2_2),.clk(gclk));
	jdff dff_B_GRC7YGEg7_2(.din(w_dff_B_b7TOsfdU2_2),.dout(w_dff_B_GRC7YGEg7_2),.clk(gclk));
	jdff dff_B_wBGrFOu90_2(.din(w_dff_B_GRC7YGEg7_2),.dout(w_dff_B_wBGrFOu90_2),.clk(gclk));
	jdff dff_B_2ld1AzU40_2(.din(w_dff_B_wBGrFOu90_2),.dout(w_dff_B_2ld1AzU40_2),.clk(gclk));
	jdff dff_B_inHNCpSI0_2(.din(w_dff_B_2ld1AzU40_2),.dout(w_dff_B_inHNCpSI0_2),.clk(gclk));
	jdff dff_B_Q5QfrRvA9_2(.din(w_dff_B_inHNCpSI0_2),.dout(w_dff_B_Q5QfrRvA9_2),.clk(gclk));
	jdff dff_B_4HYX0Wkp9_2(.din(w_dff_B_Q5QfrRvA9_2),.dout(w_dff_B_4HYX0Wkp9_2),.clk(gclk));
	jdff dff_B_Z7CtsIPD6_2(.din(w_dff_B_4HYX0Wkp9_2),.dout(w_dff_B_Z7CtsIPD6_2),.clk(gclk));
	jdff dff_B_VF1cx7eZ3_2(.din(w_dff_B_Z7CtsIPD6_2),.dout(w_dff_B_VF1cx7eZ3_2),.clk(gclk));
	jdff dff_B_fExNCCvN4_2(.din(w_dff_B_VF1cx7eZ3_2),.dout(w_dff_B_fExNCCvN4_2),.clk(gclk));
	jdff dff_B_QRalWrY44_2(.din(w_dff_B_fExNCCvN4_2),.dout(w_dff_B_QRalWrY44_2),.clk(gclk));
	jdff dff_B_wthlQ4w61_2(.din(w_dff_B_QRalWrY44_2),.dout(w_dff_B_wthlQ4w61_2),.clk(gclk));
	jdff dff_B_sIuJ0ldn2_1(.din(n1422),.dout(w_dff_B_sIuJ0ldn2_1),.clk(gclk));
	jdff dff_B_6KJiEFqY2_2(.din(n1343),.dout(w_dff_B_6KJiEFqY2_2),.clk(gclk));
	jdff dff_B_mw3p6vg57_2(.din(w_dff_B_6KJiEFqY2_2),.dout(w_dff_B_mw3p6vg57_2),.clk(gclk));
	jdff dff_B_g5ipnwXZ8_2(.din(w_dff_B_mw3p6vg57_2),.dout(w_dff_B_g5ipnwXZ8_2),.clk(gclk));
	jdff dff_B_B7gmGxNR2_2(.din(w_dff_B_g5ipnwXZ8_2),.dout(w_dff_B_B7gmGxNR2_2),.clk(gclk));
	jdff dff_B_Ti3DIU192_2(.din(w_dff_B_B7gmGxNR2_2),.dout(w_dff_B_Ti3DIU192_2),.clk(gclk));
	jdff dff_B_lXKsN52i6_2(.din(w_dff_B_Ti3DIU192_2),.dout(w_dff_B_lXKsN52i6_2),.clk(gclk));
	jdff dff_B_1W4sHzwi9_2(.din(w_dff_B_lXKsN52i6_2),.dout(w_dff_B_1W4sHzwi9_2),.clk(gclk));
	jdff dff_B_RAn4t7HL8_2(.din(w_dff_B_1W4sHzwi9_2),.dout(w_dff_B_RAn4t7HL8_2),.clk(gclk));
	jdff dff_B_ELJ6mODA6_2(.din(w_dff_B_RAn4t7HL8_2),.dout(w_dff_B_ELJ6mODA6_2),.clk(gclk));
	jdff dff_B_dwQbV2VH6_2(.din(w_dff_B_ELJ6mODA6_2),.dout(w_dff_B_dwQbV2VH6_2),.clk(gclk));
	jdff dff_B_O7zE7Wi63_2(.din(w_dff_B_dwQbV2VH6_2),.dout(w_dff_B_O7zE7Wi63_2),.clk(gclk));
	jdff dff_B_FtPLZGxp7_2(.din(w_dff_B_O7zE7Wi63_2),.dout(w_dff_B_FtPLZGxp7_2),.clk(gclk));
	jdff dff_B_649zuP3T6_2(.din(w_dff_B_FtPLZGxp7_2),.dout(w_dff_B_649zuP3T6_2),.clk(gclk));
	jdff dff_B_cFneH57W6_2(.din(w_dff_B_649zuP3T6_2),.dout(w_dff_B_cFneH57W6_2),.clk(gclk));
	jdff dff_B_DqeffqpD8_2(.din(w_dff_B_cFneH57W6_2),.dout(w_dff_B_DqeffqpD8_2),.clk(gclk));
	jdff dff_B_bvBe0FNz4_2(.din(w_dff_B_DqeffqpD8_2),.dout(w_dff_B_bvBe0FNz4_2),.clk(gclk));
	jdff dff_B_tywvN8aH2_2(.din(w_dff_B_bvBe0FNz4_2),.dout(w_dff_B_tywvN8aH2_2),.clk(gclk));
	jdff dff_B_gLWEqJuP2_2(.din(w_dff_B_tywvN8aH2_2),.dout(w_dff_B_gLWEqJuP2_2),.clk(gclk));
	jdff dff_B_6gYaM4J94_2(.din(w_dff_B_gLWEqJuP2_2),.dout(w_dff_B_6gYaM4J94_2),.clk(gclk));
	jdff dff_B_RT9Hkvei7_2(.din(w_dff_B_6gYaM4J94_2),.dout(w_dff_B_RT9Hkvei7_2),.clk(gclk));
	jdff dff_B_Zxgv8LjW3_2(.din(w_dff_B_RT9Hkvei7_2),.dout(w_dff_B_Zxgv8LjW3_2),.clk(gclk));
	jdff dff_B_ZFv2T1Bh8_2(.din(w_dff_B_Zxgv8LjW3_2),.dout(w_dff_B_ZFv2T1Bh8_2),.clk(gclk));
	jdff dff_B_DeWHq8RW5_2(.din(w_dff_B_ZFv2T1Bh8_2),.dout(w_dff_B_DeWHq8RW5_2),.clk(gclk));
	jdff dff_B_Fn2Kytrg2_2(.din(w_dff_B_DeWHq8RW5_2),.dout(w_dff_B_Fn2Kytrg2_2),.clk(gclk));
	jdff dff_B_fOcOOTkF3_2(.din(w_dff_B_Fn2Kytrg2_2),.dout(w_dff_B_fOcOOTkF3_2),.clk(gclk));
	jdff dff_B_wqZknIfA0_2(.din(w_dff_B_fOcOOTkF3_2),.dout(w_dff_B_wqZknIfA0_2),.clk(gclk));
	jdff dff_B_XqwC3bhT1_2(.din(w_dff_B_wqZknIfA0_2),.dout(w_dff_B_XqwC3bhT1_2),.clk(gclk));
	jdff dff_B_jiJk4psO8_2(.din(w_dff_B_XqwC3bhT1_2),.dout(w_dff_B_jiJk4psO8_2),.clk(gclk));
	jdff dff_B_i43SwWRs6_2(.din(w_dff_B_jiJk4psO8_2),.dout(w_dff_B_i43SwWRs6_2),.clk(gclk));
	jdff dff_B_dXh13j5K4_2(.din(w_dff_B_i43SwWRs6_2),.dout(w_dff_B_dXh13j5K4_2),.clk(gclk));
	jdff dff_B_Kc0wYyDf7_2(.din(w_dff_B_dXh13j5K4_2),.dout(w_dff_B_Kc0wYyDf7_2),.clk(gclk));
	jdff dff_B_EvRJKgDR7_2(.din(w_dff_B_Kc0wYyDf7_2),.dout(w_dff_B_EvRJKgDR7_2),.clk(gclk));
	jdff dff_B_NjoHizA18_2(.din(w_dff_B_EvRJKgDR7_2),.dout(w_dff_B_NjoHizA18_2),.clk(gclk));
	jdff dff_B_lotqe8Oh9_2(.din(w_dff_B_NjoHizA18_2),.dout(w_dff_B_lotqe8Oh9_2),.clk(gclk));
	jdff dff_B_AXmoDAIb4_2(.din(w_dff_B_lotqe8Oh9_2),.dout(w_dff_B_AXmoDAIb4_2),.clk(gclk));
	jdff dff_B_eLZ0OLec7_2(.din(w_dff_B_AXmoDAIb4_2),.dout(w_dff_B_eLZ0OLec7_2),.clk(gclk));
	jdff dff_B_wAglXE6F0_2(.din(w_dff_B_eLZ0OLec7_2),.dout(w_dff_B_wAglXE6F0_2),.clk(gclk));
	jdff dff_B_UrBfy7n78_2(.din(w_dff_B_wAglXE6F0_2),.dout(w_dff_B_UrBfy7n78_2),.clk(gclk));
	jdff dff_B_odXcaD7i8_2(.din(w_dff_B_UrBfy7n78_2),.dout(w_dff_B_odXcaD7i8_2),.clk(gclk));
	jdff dff_B_M0LYrLI80_2(.din(w_dff_B_odXcaD7i8_2),.dout(w_dff_B_M0LYrLI80_2),.clk(gclk));
	jdff dff_B_Cg2CwX5J4_2(.din(w_dff_B_M0LYrLI80_2),.dout(w_dff_B_Cg2CwX5J4_2),.clk(gclk));
	jdff dff_B_1csLnxFv0_1(.din(n1344),.dout(w_dff_B_1csLnxFv0_1),.clk(gclk));
	jdff dff_B_b4kl91Zv3_2(.din(n1258),.dout(w_dff_B_b4kl91Zv3_2),.clk(gclk));
	jdff dff_B_QsZYzkpk1_2(.din(w_dff_B_b4kl91Zv3_2),.dout(w_dff_B_QsZYzkpk1_2),.clk(gclk));
	jdff dff_B_tNrblsGQ5_2(.din(w_dff_B_QsZYzkpk1_2),.dout(w_dff_B_tNrblsGQ5_2),.clk(gclk));
	jdff dff_B_XxOCstFK5_2(.din(w_dff_B_tNrblsGQ5_2),.dout(w_dff_B_XxOCstFK5_2),.clk(gclk));
	jdff dff_B_5ws6GyMH6_2(.din(w_dff_B_XxOCstFK5_2),.dout(w_dff_B_5ws6GyMH6_2),.clk(gclk));
	jdff dff_B_XiBkvPrz0_2(.din(w_dff_B_5ws6GyMH6_2),.dout(w_dff_B_XiBkvPrz0_2),.clk(gclk));
	jdff dff_B_ANZU9JIL9_2(.din(w_dff_B_XiBkvPrz0_2),.dout(w_dff_B_ANZU9JIL9_2),.clk(gclk));
	jdff dff_B_S7iFtZF05_2(.din(w_dff_B_ANZU9JIL9_2),.dout(w_dff_B_S7iFtZF05_2),.clk(gclk));
	jdff dff_B_G8OgqTJ99_2(.din(w_dff_B_S7iFtZF05_2),.dout(w_dff_B_G8OgqTJ99_2),.clk(gclk));
	jdff dff_B_nNTVIRhW9_2(.din(w_dff_B_G8OgqTJ99_2),.dout(w_dff_B_nNTVIRhW9_2),.clk(gclk));
	jdff dff_B_Fq3mlY0W3_2(.din(w_dff_B_nNTVIRhW9_2),.dout(w_dff_B_Fq3mlY0W3_2),.clk(gclk));
	jdff dff_B_42xAzjpx3_2(.din(w_dff_B_Fq3mlY0W3_2),.dout(w_dff_B_42xAzjpx3_2),.clk(gclk));
	jdff dff_B_PBaV0l5S1_2(.din(w_dff_B_42xAzjpx3_2),.dout(w_dff_B_PBaV0l5S1_2),.clk(gclk));
	jdff dff_B_uNJs50bg3_2(.din(w_dff_B_PBaV0l5S1_2),.dout(w_dff_B_uNJs50bg3_2),.clk(gclk));
	jdff dff_B_nJdHJFwc2_2(.din(w_dff_B_uNJs50bg3_2),.dout(w_dff_B_nJdHJFwc2_2),.clk(gclk));
	jdff dff_B_UTjvwtPY6_2(.din(w_dff_B_nJdHJFwc2_2),.dout(w_dff_B_UTjvwtPY6_2),.clk(gclk));
	jdff dff_B_IjWk86Bp9_2(.din(w_dff_B_UTjvwtPY6_2),.dout(w_dff_B_IjWk86Bp9_2),.clk(gclk));
	jdff dff_B_pnuPGRxD0_2(.din(w_dff_B_IjWk86Bp9_2),.dout(w_dff_B_pnuPGRxD0_2),.clk(gclk));
	jdff dff_B_x8cpswUn2_2(.din(w_dff_B_pnuPGRxD0_2),.dout(w_dff_B_x8cpswUn2_2),.clk(gclk));
	jdff dff_B_fGzF0AhU7_2(.din(w_dff_B_x8cpswUn2_2),.dout(w_dff_B_fGzF0AhU7_2),.clk(gclk));
	jdff dff_B_bFI6WgSD4_2(.din(w_dff_B_fGzF0AhU7_2),.dout(w_dff_B_bFI6WgSD4_2),.clk(gclk));
	jdff dff_B_095JIYNe4_2(.din(w_dff_B_bFI6WgSD4_2),.dout(w_dff_B_095JIYNe4_2),.clk(gclk));
	jdff dff_B_EiJlTDHF4_2(.din(w_dff_B_095JIYNe4_2),.dout(w_dff_B_EiJlTDHF4_2),.clk(gclk));
	jdff dff_B_bQNSlO170_2(.din(w_dff_B_EiJlTDHF4_2),.dout(w_dff_B_bQNSlO170_2),.clk(gclk));
	jdff dff_B_NB2NLA2v6_2(.din(w_dff_B_bQNSlO170_2),.dout(w_dff_B_NB2NLA2v6_2),.clk(gclk));
	jdff dff_B_MGxVDMPn2_2(.din(w_dff_B_NB2NLA2v6_2),.dout(w_dff_B_MGxVDMPn2_2),.clk(gclk));
	jdff dff_B_ZXh3Z5mH3_2(.din(w_dff_B_MGxVDMPn2_2),.dout(w_dff_B_ZXh3Z5mH3_2),.clk(gclk));
	jdff dff_B_lqvgRkIg5_2(.din(w_dff_B_ZXh3Z5mH3_2),.dout(w_dff_B_lqvgRkIg5_2),.clk(gclk));
	jdff dff_B_Ec17dfrk4_2(.din(w_dff_B_lqvgRkIg5_2),.dout(w_dff_B_Ec17dfrk4_2),.clk(gclk));
	jdff dff_B_ASikrecF2_2(.din(w_dff_B_Ec17dfrk4_2),.dout(w_dff_B_ASikrecF2_2),.clk(gclk));
	jdff dff_B_oUB0YSab3_2(.din(w_dff_B_ASikrecF2_2),.dout(w_dff_B_oUB0YSab3_2),.clk(gclk));
	jdff dff_B_rR8EqmPP1_2(.din(w_dff_B_oUB0YSab3_2),.dout(w_dff_B_rR8EqmPP1_2),.clk(gclk));
	jdff dff_B_zjR6gQcK8_2(.din(w_dff_B_rR8EqmPP1_2),.dout(w_dff_B_zjR6gQcK8_2),.clk(gclk));
	jdff dff_B_OwcYP0uH8_2(.din(w_dff_B_zjR6gQcK8_2),.dout(w_dff_B_OwcYP0uH8_2),.clk(gclk));
	jdff dff_B_3d7wCdrG2_2(.din(w_dff_B_OwcYP0uH8_2),.dout(w_dff_B_3d7wCdrG2_2),.clk(gclk));
	jdff dff_B_mahCikNx5_2(.din(w_dff_B_3d7wCdrG2_2),.dout(w_dff_B_mahCikNx5_2),.clk(gclk));
	jdff dff_B_si4xxSjr1_2(.din(w_dff_B_mahCikNx5_2),.dout(w_dff_B_si4xxSjr1_2),.clk(gclk));
	jdff dff_B_qyzV3BIc3_2(.din(w_dff_B_si4xxSjr1_2),.dout(w_dff_B_qyzV3BIc3_2),.clk(gclk));
	jdff dff_B_9SfuAkYY9_1(.din(n1259),.dout(w_dff_B_9SfuAkYY9_1),.clk(gclk));
	jdff dff_B_FsMcM0tO7_2(.din(n1168),.dout(w_dff_B_FsMcM0tO7_2),.clk(gclk));
	jdff dff_B_2ED1pqdD9_2(.din(w_dff_B_FsMcM0tO7_2),.dout(w_dff_B_2ED1pqdD9_2),.clk(gclk));
	jdff dff_B_jzNsQ8RR5_2(.din(w_dff_B_2ED1pqdD9_2),.dout(w_dff_B_jzNsQ8RR5_2),.clk(gclk));
	jdff dff_B_PRx9EmQN4_2(.din(w_dff_B_jzNsQ8RR5_2),.dout(w_dff_B_PRx9EmQN4_2),.clk(gclk));
	jdff dff_B_GtqUXrql6_2(.din(w_dff_B_PRx9EmQN4_2),.dout(w_dff_B_GtqUXrql6_2),.clk(gclk));
	jdff dff_B_JnZ8EYwP5_2(.din(w_dff_B_GtqUXrql6_2),.dout(w_dff_B_JnZ8EYwP5_2),.clk(gclk));
	jdff dff_B_5tNGFGjg9_2(.din(w_dff_B_JnZ8EYwP5_2),.dout(w_dff_B_5tNGFGjg9_2),.clk(gclk));
	jdff dff_B_ddYVAcUU7_2(.din(w_dff_B_5tNGFGjg9_2),.dout(w_dff_B_ddYVAcUU7_2),.clk(gclk));
	jdff dff_B_5YFqgaWt4_2(.din(w_dff_B_ddYVAcUU7_2),.dout(w_dff_B_5YFqgaWt4_2),.clk(gclk));
	jdff dff_B_oUbmb7iS9_2(.din(w_dff_B_5YFqgaWt4_2),.dout(w_dff_B_oUbmb7iS9_2),.clk(gclk));
	jdff dff_B_Kqs9sEQy3_2(.din(w_dff_B_oUbmb7iS9_2),.dout(w_dff_B_Kqs9sEQy3_2),.clk(gclk));
	jdff dff_B_o7EUY3su9_2(.din(w_dff_B_Kqs9sEQy3_2),.dout(w_dff_B_o7EUY3su9_2),.clk(gclk));
	jdff dff_B_mFHopx8k7_2(.din(w_dff_B_o7EUY3su9_2),.dout(w_dff_B_mFHopx8k7_2),.clk(gclk));
	jdff dff_B_vPeapwCx7_2(.din(w_dff_B_mFHopx8k7_2),.dout(w_dff_B_vPeapwCx7_2),.clk(gclk));
	jdff dff_B_LntdU5Z96_2(.din(w_dff_B_vPeapwCx7_2),.dout(w_dff_B_LntdU5Z96_2),.clk(gclk));
	jdff dff_B_LlkzF4AE4_2(.din(w_dff_B_LntdU5Z96_2),.dout(w_dff_B_LlkzF4AE4_2),.clk(gclk));
	jdff dff_B_UoDF4jVm3_2(.din(w_dff_B_LlkzF4AE4_2),.dout(w_dff_B_UoDF4jVm3_2),.clk(gclk));
	jdff dff_B_mlborhS82_2(.din(w_dff_B_UoDF4jVm3_2),.dout(w_dff_B_mlborhS82_2),.clk(gclk));
	jdff dff_B_kv6fnce34_2(.din(w_dff_B_mlborhS82_2),.dout(w_dff_B_kv6fnce34_2),.clk(gclk));
	jdff dff_B_F5EZnrfI6_2(.din(w_dff_B_kv6fnce34_2),.dout(w_dff_B_F5EZnrfI6_2),.clk(gclk));
	jdff dff_B_hg5VPneE7_2(.din(w_dff_B_F5EZnrfI6_2),.dout(w_dff_B_hg5VPneE7_2),.clk(gclk));
	jdff dff_B_Zc12SvIE2_2(.din(w_dff_B_hg5VPneE7_2),.dout(w_dff_B_Zc12SvIE2_2),.clk(gclk));
	jdff dff_B_9JW8665k2_2(.din(w_dff_B_Zc12SvIE2_2),.dout(w_dff_B_9JW8665k2_2),.clk(gclk));
	jdff dff_B_GC3jK5Dl2_2(.din(w_dff_B_9JW8665k2_2),.dout(w_dff_B_GC3jK5Dl2_2),.clk(gclk));
	jdff dff_B_g7K8x2lD0_2(.din(w_dff_B_GC3jK5Dl2_2),.dout(w_dff_B_g7K8x2lD0_2),.clk(gclk));
	jdff dff_B_9zfFNM3v5_2(.din(w_dff_B_g7K8x2lD0_2),.dout(w_dff_B_9zfFNM3v5_2),.clk(gclk));
	jdff dff_B_vfkppYBB0_2(.din(w_dff_B_9zfFNM3v5_2),.dout(w_dff_B_vfkppYBB0_2),.clk(gclk));
	jdff dff_B_JWG6VLI99_2(.din(w_dff_B_vfkppYBB0_2),.dout(w_dff_B_JWG6VLI99_2),.clk(gclk));
	jdff dff_B_xwEi4aM58_2(.din(w_dff_B_JWG6VLI99_2),.dout(w_dff_B_xwEi4aM58_2),.clk(gclk));
	jdff dff_B_m2V0cs3H6_2(.din(w_dff_B_xwEi4aM58_2),.dout(w_dff_B_m2V0cs3H6_2),.clk(gclk));
	jdff dff_B_uhzNH2U43_2(.din(w_dff_B_m2V0cs3H6_2),.dout(w_dff_B_uhzNH2U43_2),.clk(gclk));
	jdff dff_B_y8yadeKv2_2(.din(w_dff_B_uhzNH2U43_2),.dout(w_dff_B_y8yadeKv2_2),.clk(gclk));
	jdff dff_B_J8TzKbhy6_2(.din(w_dff_B_y8yadeKv2_2),.dout(w_dff_B_J8TzKbhy6_2),.clk(gclk));
	jdff dff_B_v8I2cg8R8_2(.din(w_dff_B_J8TzKbhy6_2),.dout(w_dff_B_v8I2cg8R8_2),.clk(gclk));
	jdff dff_B_22AifnwD9_2(.din(w_dff_B_v8I2cg8R8_2),.dout(w_dff_B_22AifnwD9_2),.clk(gclk));
	jdff dff_B_Ow6XnM5z2_1(.din(n1169),.dout(w_dff_B_Ow6XnM5z2_1),.clk(gclk));
	jdff dff_B_fXdVR7Yh4_2(.din(n1064),.dout(w_dff_B_fXdVR7Yh4_2),.clk(gclk));
	jdff dff_B_P4h4V8Nh2_2(.din(w_dff_B_fXdVR7Yh4_2),.dout(w_dff_B_P4h4V8Nh2_2),.clk(gclk));
	jdff dff_B_HxI3PnX11_2(.din(w_dff_B_P4h4V8Nh2_2),.dout(w_dff_B_HxI3PnX11_2),.clk(gclk));
	jdff dff_B_KWBjY2yn2_2(.din(w_dff_B_HxI3PnX11_2),.dout(w_dff_B_KWBjY2yn2_2),.clk(gclk));
	jdff dff_B_mKkk714A4_2(.din(w_dff_B_KWBjY2yn2_2),.dout(w_dff_B_mKkk714A4_2),.clk(gclk));
	jdff dff_B_qJJthC0G1_2(.din(w_dff_B_mKkk714A4_2),.dout(w_dff_B_qJJthC0G1_2),.clk(gclk));
	jdff dff_B_mxh4hOpr8_2(.din(w_dff_B_qJJthC0G1_2),.dout(w_dff_B_mxh4hOpr8_2),.clk(gclk));
	jdff dff_B_M77jESMV4_2(.din(w_dff_B_mxh4hOpr8_2),.dout(w_dff_B_M77jESMV4_2),.clk(gclk));
	jdff dff_B_mW368jgu3_2(.din(w_dff_B_M77jESMV4_2),.dout(w_dff_B_mW368jgu3_2),.clk(gclk));
	jdff dff_B_3CodNuHe9_2(.din(w_dff_B_mW368jgu3_2),.dout(w_dff_B_3CodNuHe9_2),.clk(gclk));
	jdff dff_B_qmSuJsmC7_2(.din(w_dff_B_3CodNuHe9_2),.dout(w_dff_B_qmSuJsmC7_2),.clk(gclk));
	jdff dff_B_cOYrjpoi4_2(.din(w_dff_B_qmSuJsmC7_2),.dout(w_dff_B_cOYrjpoi4_2),.clk(gclk));
	jdff dff_B_Z18h3vrZ8_2(.din(w_dff_B_cOYrjpoi4_2),.dout(w_dff_B_Z18h3vrZ8_2),.clk(gclk));
	jdff dff_B_lYFzWjRi4_2(.din(w_dff_B_Z18h3vrZ8_2),.dout(w_dff_B_lYFzWjRi4_2),.clk(gclk));
	jdff dff_B_qvJ3F9DW2_2(.din(w_dff_B_lYFzWjRi4_2),.dout(w_dff_B_qvJ3F9DW2_2),.clk(gclk));
	jdff dff_B_Hf6gstuf4_2(.din(w_dff_B_qvJ3F9DW2_2),.dout(w_dff_B_Hf6gstuf4_2),.clk(gclk));
	jdff dff_B_C5NwgdrA5_2(.din(w_dff_B_Hf6gstuf4_2),.dout(w_dff_B_C5NwgdrA5_2),.clk(gclk));
	jdff dff_B_YvHI9ZI63_2(.din(w_dff_B_C5NwgdrA5_2),.dout(w_dff_B_YvHI9ZI63_2),.clk(gclk));
	jdff dff_B_P5xYgdSi5_2(.din(w_dff_B_YvHI9ZI63_2),.dout(w_dff_B_P5xYgdSi5_2),.clk(gclk));
	jdff dff_B_W5nzsXYb7_2(.din(w_dff_B_P5xYgdSi5_2),.dout(w_dff_B_W5nzsXYb7_2),.clk(gclk));
	jdff dff_B_vlnoy0995_2(.din(w_dff_B_W5nzsXYb7_2),.dout(w_dff_B_vlnoy0995_2),.clk(gclk));
	jdff dff_B_D3JC63K48_2(.din(w_dff_B_vlnoy0995_2),.dout(w_dff_B_D3JC63K48_2),.clk(gclk));
	jdff dff_B_PaiYz4uk8_2(.din(w_dff_B_D3JC63K48_2),.dout(w_dff_B_PaiYz4uk8_2),.clk(gclk));
	jdff dff_B_4dNax5Ww0_2(.din(w_dff_B_PaiYz4uk8_2),.dout(w_dff_B_4dNax5Ww0_2),.clk(gclk));
	jdff dff_B_QXnmCyxB3_2(.din(w_dff_B_4dNax5Ww0_2),.dout(w_dff_B_QXnmCyxB3_2),.clk(gclk));
	jdff dff_B_1OwSHxWC7_2(.din(w_dff_B_QXnmCyxB3_2),.dout(w_dff_B_1OwSHxWC7_2),.clk(gclk));
	jdff dff_B_K27QHcQL5_2(.din(w_dff_B_1OwSHxWC7_2),.dout(w_dff_B_K27QHcQL5_2),.clk(gclk));
	jdff dff_B_dAPh4Opn0_2(.din(w_dff_B_K27QHcQL5_2),.dout(w_dff_B_dAPh4Opn0_2),.clk(gclk));
	jdff dff_B_dAL4aXgJ4_2(.din(w_dff_B_dAPh4Opn0_2),.dout(w_dff_B_dAL4aXgJ4_2),.clk(gclk));
	jdff dff_B_N9dgmGfc2_2(.din(w_dff_B_dAL4aXgJ4_2),.dout(w_dff_B_N9dgmGfc2_2),.clk(gclk));
	jdff dff_B_ZWAQwnOr9_2(.din(w_dff_B_N9dgmGfc2_2),.dout(w_dff_B_ZWAQwnOr9_2),.clk(gclk));
	jdff dff_B_PMFJBWlE4_2(.din(w_dff_B_ZWAQwnOr9_2),.dout(w_dff_B_PMFJBWlE4_2),.clk(gclk));
	jdff dff_B_Z0oss8sb3_1(.din(n1065),.dout(w_dff_B_Z0oss8sb3_1),.clk(gclk));
	jdff dff_B_Mwi8CdeB6_2(.din(n966),.dout(w_dff_B_Mwi8CdeB6_2),.clk(gclk));
	jdff dff_B_z5EpUGAC6_2(.din(w_dff_B_Mwi8CdeB6_2),.dout(w_dff_B_z5EpUGAC6_2),.clk(gclk));
	jdff dff_B_XH4IWRzp9_2(.din(w_dff_B_z5EpUGAC6_2),.dout(w_dff_B_XH4IWRzp9_2),.clk(gclk));
	jdff dff_B_K2wgqb1J8_2(.din(w_dff_B_XH4IWRzp9_2),.dout(w_dff_B_K2wgqb1J8_2),.clk(gclk));
	jdff dff_B_hbks4zt12_2(.din(w_dff_B_K2wgqb1J8_2),.dout(w_dff_B_hbks4zt12_2),.clk(gclk));
	jdff dff_B_qyTI3Nyt3_2(.din(w_dff_B_hbks4zt12_2),.dout(w_dff_B_qyTI3Nyt3_2),.clk(gclk));
	jdff dff_B_Dyoe2unM8_2(.din(w_dff_B_qyTI3Nyt3_2),.dout(w_dff_B_Dyoe2unM8_2),.clk(gclk));
	jdff dff_B_pBRBWnLh8_2(.din(w_dff_B_Dyoe2unM8_2),.dout(w_dff_B_pBRBWnLh8_2),.clk(gclk));
	jdff dff_B_QcXGHQf89_2(.din(w_dff_B_pBRBWnLh8_2),.dout(w_dff_B_QcXGHQf89_2),.clk(gclk));
	jdff dff_B_Fw28KfIW4_2(.din(w_dff_B_QcXGHQf89_2),.dout(w_dff_B_Fw28KfIW4_2),.clk(gclk));
	jdff dff_B_PIOMStCF6_2(.din(w_dff_B_Fw28KfIW4_2),.dout(w_dff_B_PIOMStCF6_2),.clk(gclk));
	jdff dff_B_gShgcL5Z6_2(.din(w_dff_B_PIOMStCF6_2),.dout(w_dff_B_gShgcL5Z6_2),.clk(gclk));
	jdff dff_B_rie49QFk7_2(.din(w_dff_B_gShgcL5Z6_2),.dout(w_dff_B_rie49QFk7_2),.clk(gclk));
	jdff dff_B_SuTYyFwc0_2(.din(w_dff_B_rie49QFk7_2),.dout(w_dff_B_SuTYyFwc0_2),.clk(gclk));
	jdff dff_B_3z9HK80M4_2(.din(w_dff_B_SuTYyFwc0_2),.dout(w_dff_B_3z9HK80M4_2),.clk(gclk));
	jdff dff_B_riCzz8px7_2(.din(w_dff_B_3z9HK80M4_2),.dout(w_dff_B_riCzz8px7_2),.clk(gclk));
	jdff dff_B_rWRAWtER1_2(.din(w_dff_B_riCzz8px7_2),.dout(w_dff_B_rWRAWtER1_2),.clk(gclk));
	jdff dff_B_wxI1J3450_2(.din(w_dff_B_rWRAWtER1_2),.dout(w_dff_B_wxI1J3450_2),.clk(gclk));
	jdff dff_B_3LSC9JC04_2(.din(w_dff_B_wxI1J3450_2),.dout(w_dff_B_3LSC9JC04_2),.clk(gclk));
	jdff dff_B_H4NMfe866_2(.din(w_dff_B_3LSC9JC04_2),.dout(w_dff_B_H4NMfe866_2),.clk(gclk));
	jdff dff_B_Be4zUztE7_2(.din(w_dff_B_H4NMfe866_2),.dout(w_dff_B_Be4zUztE7_2),.clk(gclk));
	jdff dff_B_fnUFx6UZ3_2(.din(w_dff_B_Be4zUztE7_2),.dout(w_dff_B_fnUFx6UZ3_2),.clk(gclk));
	jdff dff_B_durrI5fz2_2(.din(w_dff_B_fnUFx6UZ3_2),.dout(w_dff_B_durrI5fz2_2),.clk(gclk));
	jdff dff_B_AGj8QWtJ3_2(.din(w_dff_B_durrI5fz2_2),.dout(w_dff_B_AGj8QWtJ3_2),.clk(gclk));
	jdff dff_B_70vRGkCI2_2(.din(w_dff_B_AGj8QWtJ3_2),.dout(w_dff_B_70vRGkCI2_2),.clk(gclk));
	jdff dff_B_RgH76awt7_2(.din(w_dff_B_70vRGkCI2_2),.dout(w_dff_B_RgH76awt7_2),.clk(gclk));
	jdff dff_B_xFU6vod69_2(.din(w_dff_B_RgH76awt7_2),.dout(w_dff_B_xFU6vod69_2),.clk(gclk));
	jdff dff_B_SadRMwjg6_2(.din(w_dff_B_xFU6vod69_2),.dout(w_dff_B_SadRMwjg6_2),.clk(gclk));
	jdff dff_B_vTxBxvLn4_2(.din(w_dff_B_SadRMwjg6_2),.dout(w_dff_B_vTxBxvLn4_2),.clk(gclk));
	jdff dff_B_rM9QpD1R3_1(.din(n967),.dout(w_dff_B_rM9QpD1R3_1),.clk(gclk));
	jdff dff_B_5dAVkk415_2(.din(n861),.dout(w_dff_B_5dAVkk415_2),.clk(gclk));
	jdff dff_B_aEObCI7S3_2(.din(w_dff_B_5dAVkk415_2),.dout(w_dff_B_aEObCI7S3_2),.clk(gclk));
	jdff dff_B_q4kr5DnY3_2(.din(w_dff_B_aEObCI7S3_2),.dout(w_dff_B_q4kr5DnY3_2),.clk(gclk));
	jdff dff_B_TsoL5NO09_2(.din(w_dff_B_q4kr5DnY3_2),.dout(w_dff_B_TsoL5NO09_2),.clk(gclk));
	jdff dff_B_w0g1rqsj8_2(.din(w_dff_B_TsoL5NO09_2),.dout(w_dff_B_w0g1rqsj8_2),.clk(gclk));
	jdff dff_B_uz6FBTgE1_2(.din(w_dff_B_w0g1rqsj8_2),.dout(w_dff_B_uz6FBTgE1_2),.clk(gclk));
	jdff dff_B_ifSb8xnW1_2(.din(w_dff_B_uz6FBTgE1_2),.dout(w_dff_B_ifSb8xnW1_2),.clk(gclk));
	jdff dff_B_twNRafDj6_2(.din(w_dff_B_ifSb8xnW1_2),.dout(w_dff_B_twNRafDj6_2),.clk(gclk));
	jdff dff_B_RWbUv56y6_2(.din(w_dff_B_twNRafDj6_2),.dout(w_dff_B_RWbUv56y6_2),.clk(gclk));
	jdff dff_B_wJEGs35L2_2(.din(w_dff_B_RWbUv56y6_2),.dout(w_dff_B_wJEGs35L2_2),.clk(gclk));
	jdff dff_B_wrFkDeYM7_2(.din(w_dff_B_wJEGs35L2_2),.dout(w_dff_B_wrFkDeYM7_2),.clk(gclk));
	jdff dff_B_IDmoxZk77_2(.din(w_dff_B_wrFkDeYM7_2),.dout(w_dff_B_IDmoxZk77_2),.clk(gclk));
	jdff dff_B_K1cx9ejt3_2(.din(w_dff_B_IDmoxZk77_2),.dout(w_dff_B_K1cx9ejt3_2),.clk(gclk));
	jdff dff_B_Xz83PU8N3_2(.din(w_dff_B_K1cx9ejt3_2),.dout(w_dff_B_Xz83PU8N3_2),.clk(gclk));
	jdff dff_B_9MEZUAb25_2(.din(w_dff_B_Xz83PU8N3_2),.dout(w_dff_B_9MEZUAb25_2),.clk(gclk));
	jdff dff_B_VJnHLuVn6_2(.din(w_dff_B_9MEZUAb25_2),.dout(w_dff_B_VJnHLuVn6_2),.clk(gclk));
	jdff dff_B_u5l4rsjr6_2(.din(w_dff_B_VJnHLuVn6_2),.dout(w_dff_B_u5l4rsjr6_2),.clk(gclk));
	jdff dff_B_QLfIW2Nn0_2(.din(w_dff_B_u5l4rsjr6_2),.dout(w_dff_B_QLfIW2Nn0_2),.clk(gclk));
	jdff dff_B_Tn4eHpk71_2(.din(w_dff_B_QLfIW2Nn0_2),.dout(w_dff_B_Tn4eHpk71_2),.clk(gclk));
	jdff dff_B_pLlPYgku6_2(.din(w_dff_B_Tn4eHpk71_2),.dout(w_dff_B_pLlPYgku6_2),.clk(gclk));
	jdff dff_B_1D5k8vXx1_2(.din(w_dff_B_pLlPYgku6_2),.dout(w_dff_B_1D5k8vXx1_2),.clk(gclk));
	jdff dff_B_EkusFtkZ6_2(.din(w_dff_B_1D5k8vXx1_2),.dout(w_dff_B_EkusFtkZ6_2),.clk(gclk));
	jdff dff_B_7mTBadUp4_2(.din(w_dff_B_EkusFtkZ6_2),.dout(w_dff_B_7mTBadUp4_2),.clk(gclk));
	jdff dff_B_gPHTXJU91_2(.din(w_dff_B_7mTBadUp4_2),.dout(w_dff_B_gPHTXJU91_2),.clk(gclk));
	jdff dff_B_eWwKaM8K4_2(.din(w_dff_B_gPHTXJU91_2),.dout(w_dff_B_eWwKaM8K4_2),.clk(gclk));
	jdff dff_B_Bg6ghQej4_2(.din(w_dff_B_eWwKaM8K4_2),.dout(w_dff_B_Bg6ghQej4_2),.clk(gclk));
	jdff dff_B_QYADrKf36_1(.din(n862),.dout(w_dff_B_QYADrKf36_1),.clk(gclk));
	jdff dff_B_iqYUAous7_2(.din(n762),.dout(w_dff_B_iqYUAous7_2),.clk(gclk));
	jdff dff_B_IEgBySH99_2(.din(w_dff_B_iqYUAous7_2),.dout(w_dff_B_IEgBySH99_2),.clk(gclk));
	jdff dff_B_nmKsp4GW7_2(.din(w_dff_B_IEgBySH99_2),.dout(w_dff_B_nmKsp4GW7_2),.clk(gclk));
	jdff dff_B_sSrGumgj2_2(.din(w_dff_B_nmKsp4GW7_2),.dout(w_dff_B_sSrGumgj2_2),.clk(gclk));
	jdff dff_B_2xqrFsFT3_2(.din(w_dff_B_sSrGumgj2_2),.dout(w_dff_B_2xqrFsFT3_2),.clk(gclk));
	jdff dff_B_PeuKAcu55_2(.din(w_dff_B_2xqrFsFT3_2),.dout(w_dff_B_PeuKAcu55_2),.clk(gclk));
	jdff dff_B_O6TyCTLV1_2(.din(w_dff_B_PeuKAcu55_2),.dout(w_dff_B_O6TyCTLV1_2),.clk(gclk));
	jdff dff_B_V4O8t3vE8_2(.din(w_dff_B_O6TyCTLV1_2),.dout(w_dff_B_V4O8t3vE8_2),.clk(gclk));
	jdff dff_B_nh2rqO655_2(.din(w_dff_B_V4O8t3vE8_2),.dout(w_dff_B_nh2rqO655_2),.clk(gclk));
	jdff dff_B_tkHSC4hs7_2(.din(w_dff_B_nh2rqO655_2),.dout(w_dff_B_tkHSC4hs7_2),.clk(gclk));
	jdff dff_B_WVMS96HE7_2(.din(w_dff_B_tkHSC4hs7_2),.dout(w_dff_B_WVMS96HE7_2),.clk(gclk));
	jdff dff_B_SklZIgxa3_2(.din(w_dff_B_WVMS96HE7_2),.dout(w_dff_B_SklZIgxa3_2),.clk(gclk));
	jdff dff_B_DqNHx9xf9_2(.din(w_dff_B_SklZIgxa3_2),.dout(w_dff_B_DqNHx9xf9_2),.clk(gclk));
	jdff dff_B_Lc8xv4eH8_2(.din(w_dff_B_DqNHx9xf9_2),.dout(w_dff_B_Lc8xv4eH8_2),.clk(gclk));
	jdff dff_B_0C8Y6kl37_2(.din(w_dff_B_Lc8xv4eH8_2),.dout(w_dff_B_0C8Y6kl37_2),.clk(gclk));
	jdff dff_B_MusmQAan0_2(.din(w_dff_B_0C8Y6kl37_2),.dout(w_dff_B_MusmQAan0_2),.clk(gclk));
	jdff dff_B_2jQ2rd5G9_2(.din(w_dff_B_MusmQAan0_2),.dout(w_dff_B_2jQ2rd5G9_2),.clk(gclk));
	jdff dff_B_bbKFYL1K1_2(.din(w_dff_B_2jQ2rd5G9_2),.dout(w_dff_B_bbKFYL1K1_2),.clk(gclk));
	jdff dff_B_dGWY89kj9_2(.din(w_dff_B_bbKFYL1K1_2),.dout(w_dff_B_dGWY89kj9_2),.clk(gclk));
	jdff dff_B_aUznYYAe2_2(.din(w_dff_B_dGWY89kj9_2),.dout(w_dff_B_aUznYYAe2_2),.clk(gclk));
	jdff dff_B_rGFNe1vY4_2(.din(w_dff_B_aUznYYAe2_2),.dout(w_dff_B_rGFNe1vY4_2),.clk(gclk));
	jdff dff_B_mIlvcbW99_2(.din(w_dff_B_rGFNe1vY4_2),.dout(w_dff_B_mIlvcbW99_2),.clk(gclk));
	jdff dff_B_GrOGSWfp7_2(.din(w_dff_B_mIlvcbW99_2),.dout(w_dff_B_GrOGSWfp7_2),.clk(gclk));
	jdff dff_B_j9Ffr4DS0_1(.din(n763),.dout(w_dff_B_j9Ffr4DS0_1),.clk(gclk));
	jdff dff_B_S7TvtqRR6_2(.din(n669),.dout(w_dff_B_S7TvtqRR6_2),.clk(gclk));
	jdff dff_B_wU3lPNwg6_2(.din(w_dff_B_S7TvtqRR6_2),.dout(w_dff_B_wU3lPNwg6_2),.clk(gclk));
	jdff dff_B_KvYMa5gq0_2(.din(w_dff_B_wU3lPNwg6_2),.dout(w_dff_B_KvYMa5gq0_2),.clk(gclk));
	jdff dff_B_JcfDtML31_2(.din(w_dff_B_KvYMa5gq0_2),.dout(w_dff_B_JcfDtML31_2),.clk(gclk));
	jdff dff_B_F6mLJgiV3_2(.din(w_dff_B_JcfDtML31_2),.dout(w_dff_B_F6mLJgiV3_2),.clk(gclk));
	jdff dff_B_HiaFSaBM4_2(.din(w_dff_B_F6mLJgiV3_2),.dout(w_dff_B_HiaFSaBM4_2),.clk(gclk));
	jdff dff_B_S2wL8ocN7_2(.din(w_dff_B_HiaFSaBM4_2),.dout(w_dff_B_S2wL8ocN7_2),.clk(gclk));
	jdff dff_B_6L2vsn9P1_2(.din(w_dff_B_S2wL8ocN7_2),.dout(w_dff_B_6L2vsn9P1_2),.clk(gclk));
	jdff dff_B_EXuGGKSs2_2(.din(w_dff_B_6L2vsn9P1_2),.dout(w_dff_B_EXuGGKSs2_2),.clk(gclk));
	jdff dff_B_j8iIcsy09_2(.din(w_dff_B_EXuGGKSs2_2),.dout(w_dff_B_j8iIcsy09_2),.clk(gclk));
	jdff dff_B_8OE73jPJ3_2(.din(w_dff_B_j8iIcsy09_2),.dout(w_dff_B_8OE73jPJ3_2),.clk(gclk));
	jdff dff_B_LPNmaUta7_2(.din(w_dff_B_8OE73jPJ3_2),.dout(w_dff_B_LPNmaUta7_2),.clk(gclk));
	jdff dff_B_0gKLIgS97_2(.din(w_dff_B_LPNmaUta7_2),.dout(w_dff_B_0gKLIgS97_2),.clk(gclk));
	jdff dff_B_zJhJNn6o8_2(.din(w_dff_B_0gKLIgS97_2),.dout(w_dff_B_zJhJNn6o8_2),.clk(gclk));
	jdff dff_B_f8npws4O8_2(.din(w_dff_B_zJhJNn6o8_2),.dout(w_dff_B_f8npws4O8_2),.clk(gclk));
	jdff dff_B_NJOTFBwo4_2(.din(w_dff_B_f8npws4O8_2),.dout(w_dff_B_NJOTFBwo4_2),.clk(gclk));
	jdff dff_B_PQd7iCdk7_2(.din(w_dff_B_NJOTFBwo4_2),.dout(w_dff_B_PQd7iCdk7_2),.clk(gclk));
	jdff dff_B_dgvqKwQl5_2(.din(w_dff_B_PQd7iCdk7_2),.dout(w_dff_B_dgvqKwQl5_2),.clk(gclk));
	jdff dff_B_9uQXoqq93_2(.din(w_dff_B_dgvqKwQl5_2),.dout(w_dff_B_9uQXoqq93_2),.clk(gclk));
	jdff dff_B_BUOFNaTh0_2(.din(w_dff_B_9uQXoqq93_2),.dout(w_dff_B_BUOFNaTh0_2),.clk(gclk));
	jdff dff_B_mW1TSD8L4_1(.din(n670),.dout(w_dff_B_mW1TSD8L4_1),.clk(gclk));
	jdff dff_B_WKBOTvv13_2(.din(n583),.dout(w_dff_B_WKBOTvv13_2),.clk(gclk));
	jdff dff_B_sqn5zKLR6_2(.din(w_dff_B_WKBOTvv13_2),.dout(w_dff_B_sqn5zKLR6_2),.clk(gclk));
	jdff dff_B_JV4GuYjx5_2(.din(w_dff_B_sqn5zKLR6_2),.dout(w_dff_B_JV4GuYjx5_2),.clk(gclk));
	jdff dff_B_69kkkViF9_2(.din(w_dff_B_JV4GuYjx5_2),.dout(w_dff_B_69kkkViF9_2),.clk(gclk));
	jdff dff_B_M0pxyStW1_2(.din(w_dff_B_69kkkViF9_2),.dout(w_dff_B_M0pxyStW1_2),.clk(gclk));
	jdff dff_B_Es4cV7i55_2(.din(w_dff_B_M0pxyStW1_2),.dout(w_dff_B_Es4cV7i55_2),.clk(gclk));
	jdff dff_B_zMfhwVej3_2(.din(w_dff_B_Es4cV7i55_2),.dout(w_dff_B_zMfhwVej3_2),.clk(gclk));
	jdff dff_B_CtmUTiVC0_2(.din(w_dff_B_zMfhwVej3_2),.dout(w_dff_B_CtmUTiVC0_2),.clk(gclk));
	jdff dff_B_zCyAhcLj0_2(.din(w_dff_B_CtmUTiVC0_2),.dout(w_dff_B_zCyAhcLj0_2),.clk(gclk));
	jdff dff_B_iKz7KXCa2_2(.din(w_dff_B_zCyAhcLj0_2),.dout(w_dff_B_iKz7KXCa2_2),.clk(gclk));
	jdff dff_B_a8n0zfU29_2(.din(w_dff_B_iKz7KXCa2_2),.dout(w_dff_B_a8n0zfU29_2),.clk(gclk));
	jdff dff_B_PhDtRwzW1_2(.din(w_dff_B_a8n0zfU29_2),.dout(w_dff_B_PhDtRwzW1_2),.clk(gclk));
	jdff dff_B_Dz0DTGEy6_2(.din(w_dff_B_PhDtRwzW1_2),.dout(w_dff_B_Dz0DTGEy6_2),.clk(gclk));
	jdff dff_B_QU4yYePb4_2(.din(w_dff_B_Dz0DTGEy6_2),.dout(w_dff_B_QU4yYePb4_2),.clk(gclk));
	jdff dff_B_CS5SZ2Kk7_2(.din(w_dff_B_QU4yYePb4_2),.dout(w_dff_B_CS5SZ2Kk7_2),.clk(gclk));
	jdff dff_B_ACczwGNs0_2(.din(w_dff_B_CS5SZ2Kk7_2),.dout(w_dff_B_ACczwGNs0_2),.clk(gclk));
	jdff dff_B_8w35Olta4_2(.din(w_dff_B_ACczwGNs0_2),.dout(w_dff_B_8w35Olta4_2),.clk(gclk));
	jdff dff_B_1jkOuCTe1_1(.din(n584),.dout(w_dff_B_1jkOuCTe1_1),.clk(gclk));
	jdff dff_B_UU0niQwW9_2(.din(n504),.dout(w_dff_B_UU0niQwW9_2),.clk(gclk));
	jdff dff_B_KeVEyKMb1_2(.din(w_dff_B_UU0niQwW9_2),.dout(w_dff_B_KeVEyKMb1_2),.clk(gclk));
	jdff dff_B_IfGQKgo49_2(.din(w_dff_B_KeVEyKMb1_2),.dout(w_dff_B_IfGQKgo49_2),.clk(gclk));
	jdff dff_B_v8NkCyuF8_2(.din(w_dff_B_IfGQKgo49_2),.dout(w_dff_B_v8NkCyuF8_2),.clk(gclk));
	jdff dff_B_DmBSNOsi5_2(.din(w_dff_B_v8NkCyuF8_2),.dout(w_dff_B_DmBSNOsi5_2),.clk(gclk));
	jdff dff_B_Bx2gnNGo9_2(.din(w_dff_B_DmBSNOsi5_2),.dout(w_dff_B_Bx2gnNGo9_2),.clk(gclk));
	jdff dff_B_B5o8vsOp5_2(.din(w_dff_B_Bx2gnNGo9_2),.dout(w_dff_B_B5o8vsOp5_2),.clk(gclk));
	jdff dff_B_8WFP1M3O3_2(.din(w_dff_B_B5o8vsOp5_2),.dout(w_dff_B_8WFP1M3O3_2),.clk(gclk));
	jdff dff_B_EtJZypqQ0_2(.din(w_dff_B_8WFP1M3O3_2),.dout(w_dff_B_EtJZypqQ0_2),.clk(gclk));
	jdff dff_B_2hTid2xz7_2(.din(w_dff_B_EtJZypqQ0_2),.dout(w_dff_B_2hTid2xz7_2),.clk(gclk));
	jdff dff_B_wIPEjqCa4_2(.din(w_dff_B_2hTid2xz7_2),.dout(w_dff_B_wIPEjqCa4_2),.clk(gclk));
	jdff dff_B_t2VXvQob3_2(.din(w_dff_B_wIPEjqCa4_2),.dout(w_dff_B_t2VXvQob3_2),.clk(gclk));
	jdff dff_B_ugtxxaRF8_2(.din(w_dff_B_t2VXvQob3_2),.dout(w_dff_B_ugtxxaRF8_2),.clk(gclk));
	jdff dff_B_4A2pXL0w9_2(.din(w_dff_B_ugtxxaRF8_2),.dout(w_dff_B_4A2pXL0w9_2),.clk(gclk));
	jdff dff_B_o1AElAy04_1(.din(n505),.dout(w_dff_B_o1AElAy04_1),.clk(gclk));
	jdff dff_B_yaTJdMX62_2(.din(n432),.dout(w_dff_B_yaTJdMX62_2),.clk(gclk));
	jdff dff_B_0xzqZkN16_2(.din(w_dff_B_yaTJdMX62_2),.dout(w_dff_B_0xzqZkN16_2),.clk(gclk));
	jdff dff_B_x4Y8O32m2_2(.din(w_dff_B_0xzqZkN16_2),.dout(w_dff_B_x4Y8O32m2_2),.clk(gclk));
	jdff dff_B_bjdxf3zh8_2(.din(w_dff_B_x4Y8O32m2_2),.dout(w_dff_B_bjdxf3zh8_2),.clk(gclk));
	jdff dff_B_QQPzpzg94_2(.din(w_dff_B_bjdxf3zh8_2),.dout(w_dff_B_QQPzpzg94_2),.clk(gclk));
	jdff dff_B_Ygl76m6v6_2(.din(w_dff_B_QQPzpzg94_2),.dout(w_dff_B_Ygl76m6v6_2),.clk(gclk));
	jdff dff_B_F1A8SqEE5_2(.din(w_dff_B_Ygl76m6v6_2),.dout(w_dff_B_F1A8SqEE5_2),.clk(gclk));
	jdff dff_B_9Ppv3XtM6_2(.din(w_dff_B_F1A8SqEE5_2),.dout(w_dff_B_9Ppv3XtM6_2),.clk(gclk));
	jdff dff_B_csYC4KPe7_2(.din(w_dff_B_9Ppv3XtM6_2),.dout(w_dff_B_csYC4KPe7_2),.clk(gclk));
	jdff dff_B_REcqCrEE4_2(.din(w_dff_B_csYC4KPe7_2),.dout(w_dff_B_REcqCrEE4_2),.clk(gclk));
	jdff dff_B_t22o2eFd8_2(.din(w_dff_B_REcqCrEE4_2),.dout(w_dff_B_t22o2eFd8_2),.clk(gclk));
	jdff dff_B_1TPbLWoN5_2(.din(n435),.dout(w_dff_B_1TPbLWoN5_2),.clk(gclk));
	jdff dff_B_OO1D15tP2_1(.din(n433),.dout(w_dff_B_OO1D15tP2_1),.clk(gclk));
	jdff dff_B_9zEPRubG3_2(.din(n368),.dout(w_dff_B_9zEPRubG3_2),.clk(gclk));
	jdff dff_B_sqaADirs6_2(.din(w_dff_B_9zEPRubG3_2),.dout(w_dff_B_sqaADirs6_2),.clk(gclk));
	jdff dff_B_fWKoUnXJ9_2(.din(w_dff_B_sqaADirs6_2),.dout(w_dff_B_fWKoUnXJ9_2),.clk(gclk));
	jdff dff_B_QunNc8Us6_2(.din(w_dff_B_fWKoUnXJ9_2),.dout(w_dff_B_QunNc8Us6_2),.clk(gclk));
	jdff dff_B_feEC5aAb8_2(.din(w_dff_B_QunNc8Us6_2),.dout(w_dff_B_feEC5aAb8_2),.clk(gclk));
	jdff dff_B_ShoRSDqQ1_2(.din(w_dff_B_feEC5aAb8_2),.dout(w_dff_B_ShoRSDqQ1_2),.clk(gclk));
	jdff dff_B_xUKku5GK7_2(.din(w_dff_B_ShoRSDqQ1_2),.dout(w_dff_B_xUKku5GK7_2),.clk(gclk));
	jdff dff_B_03fXdbCs7_1(.din(n369),.dout(w_dff_B_03fXdbCs7_1),.clk(gclk));
	jdff dff_B_wUHlHhtp4_2(.din(n310),.dout(w_dff_B_wUHlHhtp4_2),.clk(gclk));
	jdff dff_B_YPvNkcuG0_2(.din(w_dff_B_wUHlHhtp4_2),.dout(w_dff_B_YPvNkcuG0_2),.clk(gclk));
	jdff dff_B_gIDleT7U8_2(.din(w_dff_B_YPvNkcuG0_2),.dout(w_dff_B_gIDleT7U8_2),.clk(gclk));
	jdff dff_B_InSP26yk6_2(.din(w_dff_B_gIDleT7U8_2),.dout(w_dff_B_InSP26yk6_2),.clk(gclk));
	jdff dff_B_pBKm8eeb1_1(.din(n312),.dout(w_dff_B_pBKm8eeb1_1),.clk(gclk));
	jdff dff_A_ND5nyXI76_0(.dout(w_n258_0[0]),.din(w_dff_A_ND5nyXI76_0),.clk(gclk));
	jdff dff_A_Sleh7iQV6_1(.dout(w_n258_0[1]),.din(w_dff_A_Sleh7iQV6_1),.clk(gclk));
	jdff dff_A_oB75lPv25_1(.dout(w_dff_A_Sleh7iQV6_1),.din(w_dff_A_oB75lPv25_1),.clk(gclk));
	jdff dff_B_dscEN8CP3_1(.din(n1563),.dout(w_dff_B_dscEN8CP3_1),.clk(gclk));
	jdff dff_B_gZs9LaEz2_2(.din(n1497),.dout(w_dff_B_gZs9LaEz2_2),.clk(gclk));
	jdff dff_B_PGEfNWI99_2(.din(w_dff_B_gZs9LaEz2_2),.dout(w_dff_B_PGEfNWI99_2),.clk(gclk));
	jdff dff_B_W1Ek9dO77_2(.din(w_dff_B_PGEfNWI99_2),.dout(w_dff_B_W1Ek9dO77_2),.clk(gclk));
	jdff dff_B_DDxqsWXw0_2(.din(w_dff_B_W1Ek9dO77_2),.dout(w_dff_B_DDxqsWXw0_2),.clk(gclk));
	jdff dff_B_OIYPBMRb4_2(.din(w_dff_B_DDxqsWXw0_2),.dout(w_dff_B_OIYPBMRb4_2),.clk(gclk));
	jdff dff_B_3syitiH25_2(.din(w_dff_B_OIYPBMRb4_2),.dout(w_dff_B_3syitiH25_2),.clk(gclk));
	jdff dff_B_X0r7ewxt6_2(.din(w_dff_B_3syitiH25_2),.dout(w_dff_B_X0r7ewxt6_2),.clk(gclk));
	jdff dff_B_YVKeeVHG7_2(.din(w_dff_B_X0r7ewxt6_2),.dout(w_dff_B_YVKeeVHG7_2),.clk(gclk));
	jdff dff_B_0KiXGFQ22_2(.din(w_dff_B_YVKeeVHG7_2),.dout(w_dff_B_0KiXGFQ22_2),.clk(gclk));
	jdff dff_B_OrxITFSE4_2(.din(w_dff_B_0KiXGFQ22_2),.dout(w_dff_B_OrxITFSE4_2),.clk(gclk));
	jdff dff_B_p5XSaOeV3_2(.din(w_dff_B_OrxITFSE4_2),.dout(w_dff_B_p5XSaOeV3_2),.clk(gclk));
	jdff dff_B_gX0PHthV9_2(.din(w_dff_B_p5XSaOeV3_2),.dout(w_dff_B_gX0PHthV9_2),.clk(gclk));
	jdff dff_B_tSmN1HZK4_2(.din(w_dff_B_gX0PHthV9_2),.dout(w_dff_B_tSmN1HZK4_2),.clk(gclk));
	jdff dff_B_bCg1fvIv9_2(.din(w_dff_B_tSmN1HZK4_2),.dout(w_dff_B_bCg1fvIv9_2),.clk(gclk));
	jdff dff_B_4rhMCbdM3_2(.din(w_dff_B_bCg1fvIv9_2),.dout(w_dff_B_4rhMCbdM3_2),.clk(gclk));
	jdff dff_B_zKAIuavT5_2(.din(w_dff_B_4rhMCbdM3_2),.dout(w_dff_B_zKAIuavT5_2),.clk(gclk));
	jdff dff_B_WcE5HeEP9_2(.din(w_dff_B_zKAIuavT5_2),.dout(w_dff_B_WcE5HeEP9_2),.clk(gclk));
	jdff dff_B_3v0Yo8XO9_2(.din(w_dff_B_WcE5HeEP9_2),.dout(w_dff_B_3v0Yo8XO9_2),.clk(gclk));
	jdff dff_B_qz1XyZz10_2(.din(w_dff_B_3v0Yo8XO9_2),.dout(w_dff_B_qz1XyZz10_2),.clk(gclk));
	jdff dff_B_up5Fvazq8_2(.din(w_dff_B_qz1XyZz10_2),.dout(w_dff_B_up5Fvazq8_2),.clk(gclk));
	jdff dff_B_v26EmyiN3_2(.din(w_dff_B_up5Fvazq8_2),.dout(w_dff_B_v26EmyiN3_2),.clk(gclk));
	jdff dff_B_ybA0UQjG3_2(.din(w_dff_B_v26EmyiN3_2),.dout(w_dff_B_ybA0UQjG3_2),.clk(gclk));
	jdff dff_B_gF3nxzH06_2(.din(w_dff_B_ybA0UQjG3_2),.dout(w_dff_B_gF3nxzH06_2),.clk(gclk));
	jdff dff_B_iAAMCwx31_2(.din(w_dff_B_gF3nxzH06_2),.dout(w_dff_B_iAAMCwx31_2),.clk(gclk));
	jdff dff_B_3MjKph8N1_2(.din(w_dff_B_iAAMCwx31_2),.dout(w_dff_B_3MjKph8N1_2),.clk(gclk));
	jdff dff_B_5RdFssbW6_2(.din(w_dff_B_3MjKph8N1_2),.dout(w_dff_B_5RdFssbW6_2),.clk(gclk));
	jdff dff_B_uJfkE8X17_2(.din(w_dff_B_5RdFssbW6_2),.dout(w_dff_B_uJfkE8X17_2),.clk(gclk));
	jdff dff_B_w5zmZzTC5_2(.din(w_dff_B_uJfkE8X17_2),.dout(w_dff_B_w5zmZzTC5_2),.clk(gclk));
	jdff dff_B_1goNVmJf8_2(.din(w_dff_B_w5zmZzTC5_2),.dout(w_dff_B_1goNVmJf8_2),.clk(gclk));
	jdff dff_B_RwHDKR2h5_2(.din(w_dff_B_1goNVmJf8_2),.dout(w_dff_B_RwHDKR2h5_2),.clk(gclk));
	jdff dff_B_SsVQtzwa4_2(.din(w_dff_B_RwHDKR2h5_2),.dout(w_dff_B_SsVQtzwa4_2),.clk(gclk));
	jdff dff_B_TzmBMLPI6_2(.din(w_dff_B_SsVQtzwa4_2),.dout(w_dff_B_TzmBMLPI6_2),.clk(gclk));
	jdff dff_B_H094nLHV7_2(.din(w_dff_B_TzmBMLPI6_2),.dout(w_dff_B_H094nLHV7_2),.clk(gclk));
	jdff dff_B_YWili5MT2_2(.din(w_dff_B_H094nLHV7_2),.dout(w_dff_B_YWili5MT2_2),.clk(gclk));
	jdff dff_B_NXZJJkEl4_2(.din(w_dff_B_YWili5MT2_2),.dout(w_dff_B_NXZJJkEl4_2),.clk(gclk));
	jdff dff_B_eODnW7n96_2(.din(w_dff_B_NXZJJkEl4_2),.dout(w_dff_B_eODnW7n96_2),.clk(gclk));
	jdff dff_B_VVeJMVTu0_2(.din(w_dff_B_eODnW7n96_2),.dout(w_dff_B_VVeJMVTu0_2),.clk(gclk));
	jdff dff_B_AFw9awkp9_2(.din(w_dff_B_VVeJMVTu0_2),.dout(w_dff_B_AFw9awkp9_2),.clk(gclk));
	jdff dff_B_F4SSRS5d3_2(.din(w_dff_B_AFw9awkp9_2),.dout(w_dff_B_F4SSRS5d3_2),.clk(gclk));
	jdff dff_B_unPgbOLe3_2(.din(w_dff_B_F4SSRS5d3_2),.dout(w_dff_B_unPgbOLe3_2),.clk(gclk));
	jdff dff_B_xC7olaV15_2(.din(w_dff_B_unPgbOLe3_2),.dout(w_dff_B_xC7olaV15_2),.clk(gclk));
	jdff dff_B_oWqxCd2C4_2(.din(w_dff_B_xC7olaV15_2),.dout(w_dff_B_oWqxCd2C4_2),.clk(gclk));
	jdff dff_B_XnMTc3tc5_2(.din(w_dff_B_oWqxCd2C4_2),.dout(w_dff_B_XnMTc3tc5_2),.clk(gclk));
	jdff dff_B_0UDdrsng6_2(.din(w_dff_B_XnMTc3tc5_2),.dout(w_dff_B_0UDdrsng6_2),.clk(gclk));
	jdff dff_B_OdFVZsp64_2(.din(w_dff_B_0UDdrsng6_2),.dout(w_dff_B_OdFVZsp64_2),.clk(gclk));
	jdff dff_B_CeQ2fuut0_2(.din(w_dff_B_OdFVZsp64_2),.dout(w_dff_B_CeQ2fuut0_2),.clk(gclk));
	jdff dff_B_ePm4FQ1L1_2(.din(w_dff_B_CeQ2fuut0_2),.dout(w_dff_B_ePm4FQ1L1_2),.clk(gclk));
	jdff dff_B_xVbS7BIv1_0(.din(n1562),.dout(w_dff_B_xVbS7BIv1_0),.clk(gclk));
	jdff dff_A_NoaSoI4S5_1(.dout(w_n1550_0[1]),.din(w_dff_A_NoaSoI4S5_1),.clk(gclk));
	jdff dff_B_lQf6csxZ2_1(.din(n1498),.dout(w_dff_B_lQf6csxZ2_1),.clk(gclk));
	jdff dff_B_K8kUTWgq2_2(.din(n1426),.dout(w_dff_B_K8kUTWgq2_2),.clk(gclk));
	jdff dff_B_CedpvwHs7_2(.din(w_dff_B_K8kUTWgq2_2),.dout(w_dff_B_CedpvwHs7_2),.clk(gclk));
	jdff dff_B_7r2aTGij9_2(.din(w_dff_B_CedpvwHs7_2),.dout(w_dff_B_7r2aTGij9_2),.clk(gclk));
	jdff dff_B_dLvlGtDV0_2(.din(w_dff_B_7r2aTGij9_2),.dout(w_dff_B_dLvlGtDV0_2),.clk(gclk));
	jdff dff_B_CMj8XDe25_2(.din(w_dff_B_dLvlGtDV0_2),.dout(w_dff_B_CMj8XDe25_2),.clk(gclk));
	jdff dff_B_Y5UX4S5g2_2(.din(w_dff_B_CMj8XDe25_2),.dout(w_dff_B_Y5UX4S5g2_2),.clk(gclk));
	jdff dff_B_fGnOEmCY6_2(.din(w_dff_B_Y5UX4S5g2_2),.dout(w_dff_B_fGnOEmCY6_2),.clk(gclk));
	jdff dff_B_dFvKUDWG2_2(.din(w_dff_B_fGnOEmCY6_2),.dout(w_dff_B_dFvKUDWG2_2),.clk(gclk));
	jdff dff_B_LZLEP57y7_2(.din(w_dff_B_dFvKUDWG2_2),.dout(w_dff_B_LZLEP57y7_2),.clk(gclk));
	jdff dff_B_mL2VAuwq7_2(.din(w_dff_B_LZLEP57y7_2),.dout(w_dff_B_mL2VAuwq7_2),.clk(gclk));
	jdff dff_B_QiyUvBsP5_2(.din(w_dff_B_mL2VAuwq7_2),.dout(w_dff_B_QiyUvBsP5_2),.clk(gclk));
	jdff dff_B_8zxexqDf3_2(.din(w_dff_B_QiyUvBsP5_2),.dout(w_dff_B_8zxexqDf3_2),.clk(gclk));
	jdff dff_B_6oIlwFf77_2(.din(w_dff_B_8zxexqDf3_2),.dout(w_dff_B_6oIlwFf77_2),.clk(gclk));
	jdff dff_B_QIeW735N2_2(.din(w_dff_B_6oIlwFf77_2),.dout(w_dff_B_QIeW735N2_2),.clk(gclk));
	jdff dff_B_t8xIgAYJ0_2(.din(w_dff_B_QIeW735N2_2),.dout(w_dff_B_t8xIgAYJ0_2),.clk(gclk));
	jdff dff_B_WjDxrsoN8_2(.din(w_dff_B_t8xIgAYJ0_2),.dout(w_dff_B_WjDxrsoN8_2),.clk(gclk));
	jdff dff_B_RJ1DzOCD2_2(.din(w_dff_B_WjDxrsoN8_2),.dout(w_dff_B_RJ1DzOCD2_2),.clk(gclk));
	jdff dff_B_dPpnypC14_2(.din(w_dff_B_RJ1DzOCD2_2),.dout(w_dff_B_dPpnypC14_2),.clk(gclk));
	jdff dff_B_YtEO3TLT3_2(.din(w_dff_B_dPpnypC14_2),.dout(w_dff_B_YtEO3TLT3_2),.clk(gclk));
	jdff dff_B_UarUl7fZ6_2(.din(w_dff_B_YtEO3TLT3_2),.dout(w_dff_B_UarUl7fZ6_2),.clk(gclk));
	jdff dff_B_Sj5WLCgo6_2(.din(w_dff_B_UarUl7fZ6_2),.dout(w_dff_B_Sj5WLCgo6_2),.clk(gclk));
	jdff dff_B_s5q85r9E2_2(.din(w_dff_B_Sj5WLCgo6_2),.dout(w_dff_B_s5q85r9E2_2),.clk(gclk));
	jdff dff_B_ALefSdLr9_2(.din(w_dff_B_s5q85r9E2_2),.dout(w_dff_B_ALefSdLr9_2),.clk(gclk));
	jdff dff_B_24P93rEn5_2(.din(w_dff_B_ALefSdLr9_2),.dout(w_dff_B_24P93rEn5_2),.clk(gclk));
	jdff dff_B_DouM5BnR5_2(.din(w_dff_B_24P93rEn5_2),.dout(w_dff_B_DouM5BnR5_2),.clk(gclk));
	jdff dff_B_XicY1ay78_2(.din(w_dff_B_DouM5BnR5_2),.dout(w_dff_B_XicY1ay78_2),.clk(gclk));
	jdff dff_B_MpMpxdGa3_2(.din(w_dff_B_XicY1ay78_2),.dout(w_dff_B_MpMpxdGa3_2),.clk(gclk));
	jdff dff_B_8XS9pli16_2(.din(w_dff_B_MpMpxdGa3_2),.dout(w_dff_B_8XS9pli16_2),.clk(gclk));
	jdff dff_B_dfwLvLV80_2(.din(w_dff_B_8XS9pli16_2),.dout(w_dff_B_dfwLvLV80_2),.clk(gclk));
	jdff dff_B_eMQrLM579_2(.din(w_dff_B_dfwLvLV80_2),.dout(w_dff_B_eMQrLM579_2),.clk(gclk));
	jdff dff_B_0g7HKPQi8_2(.din(w_dff_B_eMQrLM579_2),.dout(w_dff_B_0g7HKPQi8_2),.clk(gclk));
	jdff dff_B_gmFrnxSi7_2(.din(w_dff_B_0g7HKPQi8_2),.dout(w_dff_B_gmFrnxSi7_2),.clk(gclk));
	jdff dff_B_LHpRKbC69_2(.din(w_dff_B_gmFrnxSi7_2),.dout(w_dff_B_LHpRKbC69_2),.clk(gclk));
	jdff dff_B_W5N0RPnN5_2(.din(w_dff_B_LHpRKbC69_2),.dout(w_dff_B_W5N0RPnN5_2),.clk(gclk));
	jdff dff_B_RUCj2EVl5_2(.din(w_dff_B_W5N0RPnN5_2),.dout(w_dff_B_RUCj2EVl5_2),.clk(gclk));
	jdff dff_B_lfATVw4Z2_2(.din(w_dff_B_RUCj2EVl5_2),.dout(w_dff_B_lfATVw4Z2_2),.clk(gclk));
	jdff dff_B_9OaOwsta5_2(.din(w_dff_B_lfATVw4Z2_2),.dout(w_dff_B_9OaOwsta5_2),.clk(gclk));
	jdff dff_B_5TU4Zch19_2(.din(w_dff_B_9OaOwsta5_2),.dout(w_dff_B_5TU4Zch19_2),.clk(gclk));
	jdff dff_B_mNTGIM3g0_2(.din(w_dff_B_5TU4Zch19_2),.dout(w_dff_B_mNTGIM3g0_2),.clk(gclk));
	jdff dff_B_BNmq484u1_2(.din(w_dff_B_mNTGIM3g0_2),.dout(w_dff_B_BNmq484u1_2),.clk(gclk));
	jdff dff_B_ld4nXSo43_2(.din(w_dff_B_BNmq484u1_2),.dout(w_dff_B_ld4nXSo43_2),.clk(gclk));
	jdff dff_B_hnjWvXPB6_2(.din(w_dff_B_ld4nXSo43_2),.dout(w_dff_B_hnjWvXPB6_2),.clk(gclk));
	jdff dff_B_yDwue3896_2(.din(n1479),.dout(w_dff_B_yDwue3896_2),.clk(gclk));
	jdff dff_B_GNK67qew6_1(.din(n1427),.dout(w_dff_B_GNK67qew6_1),.clk(gclk));
	jdff dff_B_mjwuSWFV6_2(.din(n1348),.dout(w_dff_B_mjwuSWFV6_2),.clk(gclk));
	jdff dff_B_U9B1suxo8_2(.din(w_dff_B_mjwuSWFV6_2),.dout(w_dff_B_U9B1suxo8_2),.clk(gclk));
	jdff dff_B_gb66n7Gz7_2(.din(w_dff_B_U9B1suxo8_2),.dout(w_dff_B_gb66n7Gz7_2),.clk(gclk));
	jdff dff_B_M8ox9jiE1_2(.din(w_dff_B_gb66n7Gz7_2),.dout(w_dff_B_M8ox9jiE1_2),.clk(gclk));
	jdff dff_B_N6QIAid07_2(.din(w_dff_B_M8ox9jiE1_2),.dout(w_dff_B_N6QIAid07_2),.clk(gclk));
	jdff dff_B_Lx054sw25_2(.din(w_dff_B_N6QIAid07_2),.dout(w_dff_B_Lx054sw25_2),.clk(gclk));
	jdff dff_B_FCemGsSY4_2(.din(w_dff_B_Lx054sw25_2),.dout(w_dff_B_FCemGsSY4_2),.clk(gclk));
	jdff dff_B_KJFQD4d71_2(.din(w_dff_B_FCemGsSY4_2),.dout(w_dff_B_KJFQD4d71_2),.clk(gclk));
	jdff dff_B_2u4iloU37_2(.din(w_dff_B_KJFQD4d71_2),.dout(w_dff_B_2u4iloU37_2),.clk(gclk));
	jdff dff_B_nOkojfNl0_2(.din(w_dff_B_2u4iloU37_2),.dout(w_dff_B_nOkojfNl0_2),.clk(gclk));
	jdff dff_B_23B6pC2S5_2(.din(w_dff_B_nOkojfNl0_2),.dout(w_dff_B_23B6pC2S5_2),.clk(gclk));
	jdff dff_B_MLegzzsA6_2(.din(w_dff_B_23B6pC2S5_2),.dout(w_dff_B_MLegzzsA6_2),.clk(gclk));
	jdff dff_B_qfg5kSDx2_2(.din(w_dff_B_MLegzzsA6_2),.dout(w_dff_B_qfg5kSDx2_2),.clk(gclk));
	jdff dff_B_1abGkJLL3_2(.din(w_dff_B_qfg5kSDx2_2),.dout(w_dff_B_1abGkJLL3_2),.clk(gclk));
	jdff dff_B_kRKuTYsx8_2(.din(w_dff_B_1abGkJLL3_2),.dout(w_dff_B_kRKuTYsx8_2),.clk(gclk));
	jdff dff_B_Ku8lmRN92_2(.din(w_dff_B_kRKuTYsx8_2),.dout(w_dff_B_Ku8lmRN92_2),.clk(gclk));
	jdff dff_B_063y1oDD3_2(.din(w_dff_B_Ku8lmRN92_2),.dout(w_dff_B_063y1oDD3_2),.clk(gclk));
	jdff dff_B_4dR0k1Pe3_2(.din(w_dff_B_063y1oDD3_2),.dout(w_dff_B_4dR0k1Pe3_2),.clk(gclk));
	jdff dff_B_uI4duSeb9_2(.din(w_dff_B_4dR0k1Pe3_2),.dout(w_dff_B_uI4duSeb9_2),.clk(gclk));
	jdff dff_B_ekNn9Kd60_2(.din(w_dff_B_uI4duSeb9_2),.dout(w_dff_B_ekNn9Kd60_2),.clk(gclk));
	jdff dff_B_eNOnXkzs7_2(.din(w_dff_B_ekNn9Kd60_2),.dout(w_dff_B_eNOnXkzs7_2),.clk(gclk));
	jdff dff_B_pQ9JVMvA4_2(.din(w_dff_B_eNOnXkzs7_2),.dout(w_dff_B_pQ9JVMvA4_2),.clk(gclk));
	jdff dff_B_91m689Lr0_2(.din(w_dff_B_pQ9JVMvA4_2),.dout(w_dff_B_91m689Lr0_2),.clk(gclk));
	jdff dff_B_FXH8UVvw0_2(.din(w_dff_B_91m689Lr0_2),.dout(w_dff_B_FXH8UVvw0_2),.clk(gclk));
	jdff dff_B_7C8x3nza3_2(.din(w_dff_B_FXH8UVvw0_2),.dout(w_dff_B_7C8x3nza3_2),.clk(gclk));
	jdff dff_B_sW6OVQP58_2(.din(w_dff_B_7C8x3nza3_2),.dout(w_dff_B_sW6OVQP58_2),.clk(gclk));
	jdff dff_B_k6h6274F0_2(.din(w_dff_B_sW6OVQP58_2),.dout(w_dff_B_k6h6274F0_2),.clk(gclk));
	jdff dff_B_eQ2z22vz5_2(.din(w_dff_B_k6h6274F0_2),.dout(w_dff_B_eQ2z22vz5_2),.clk(gclk));
	jdff dff_B_qwQc6bcR9_2(.din(w_dff_B_eQ2z22vz5_2),.dout(w_dff_B_qwQc6bcR9_2),.clk(gclk));
	jdff dff_B_Pl7K4qeE4_2(.din(w_dff_B_qwQc6bcR9_2),.dout(w_dff_B_Pl7K4qeE4_2),.clk(gclk));
	jdff dff_B_kjwtRpYF9_2(.din(w_dff_B_Pl7K4qeE4_2),.dout(w_dff_B_kjwtRpYF9_2),.clk(gclk));
	jdff dff_B_3rpmHdA50_2(.din(w_dff_B_kjwtRpYF9_2),.dout(w_dff_B_3rpmHdA50_2),.clk(gclk));
	jdff dff_B_lmYWVv327_2(.din(w_dff_B_3rpmHdA50_2),.dout(w_dff_B_lmYWVv327_2),.clk(gclk));
	jdff dff_B_ymBku5oQ0_2(.din(w_dff_B_lmYWVv327_2),.dout(w_dff_B_ymBku5oQ0_2),.clk(gclk));
	jdff dff_B_JAcND1yG6_2(.din(w_dff_B_ymBku5oQ0_2),.dout(w_dff_B_JAcND1yG6_2),.clk(gclk));
	jdff dff_B_dGRTS4v79_2(.din(w_dff_B_JAcND1yG6_2),.dout(w_dff_B_dGRTS4v79_2),.clk(gclk));
	jdff dff_B_c8zPlz7S7_2(.din(w_dff_B_dGRTS4v79_2),.dout(w_dff_B_c8zPlz7S7_2),.clk(gclk));
	jdff dff_B_WBr45EPs8_2(.din(w_dff_B_c8zPlz7S7_2),.dout(w_dff_B_WBr45EPs8_2),.clk(gclk));
	jdff dff_B_6NUDczgV1_2(.din(w_dff_B_WBr45EPs8_2),.dout(w_dff_B_6NUDczgV1_2),.clk(gclk));
	jdff dff_B_9ek3H3DE0_2(.din(n1401),.dout(w_dff_B_9ek3H3DE0_2),.clk(gclk));
	jdff dff_B_faBXe0Lc1_1(.din(n1349),.dout(w_dff_B_faBXe0Lc1_1),.clk(gclk));
	jdff dff_B_Zy0EmF5c8_2(.din(n1263),.dout(w_dff_B_Zy0EmF5c8_2),.clk(gclk));
	jdff dff_B_wxkXcXhe5_2(.din(w_dff_B_Zy0EmF5c8_2),.dout(w_dff_B_wxkXcXhe5_2),.clk(gclk));
	jdff dff_B_6UXazMBB8_2(.din(w_dff_B_wxkXcXhe5_2),.dout(w_dff_B_6UXazMBB8_2),.clk(gclk));
	jdff dff_B_0OQ4zjqZ5_2(.din(w_dff_B_6UXazMBB8_2),.dout(w_dff_B_0OQ4zjqZ5_2),.clk(gclk));
	jdff dff_B_M37svjXN3_2(.din(w_dff_B_0OQ4zjqZ5_2),.dout(w_dff_B_M37svjXN3_2),.clk(gclk));
	jdff dff_B_48SDdk871_2(.din(w_dff_B_M37svjXN3_2),.dout(w_dff_B_48SDdk871_2),.clk(gclk));
	jdff dff_B_tDVM4FSx0_2(.din(w_dff_B_48SDdk871_2),.dout(w_dff_B_tDVM4FSx0_2),.clk(gclk));
	jdff dff_B_RnRX0C9p1_2(.din(w_dff_B_tDVM4FSx0_2),.dout(w_dff_B_RnRX0C9p1_2),.clk(gclk));
	jdff dff_B_jKbWh6lA2_2(.din(w_dff_B_RnRX0C9p1_2),.dout(w_dff_B_jKbWh6lA2_2),.clk(gclk));
	jdff dff_B_z1aBQxpj9_2(.din(w_dff_B_jKbWh6lA2_2),.dout(w_dff_B_z1aBQxpj9_2),.clk(gclk));
	jdff dff_B_zyFaztIQ2_2(.din(w_dff_B_z1aBQxpj9_2),.dout(w_dff_B_zyFaztIQ2_2),.clk(gclk));
	jdff dff_B_cX9Q2pET6_2(.din(w_dff_B_zyFaztIQ2_2),.dout(w_dff_B_cX9Q2pET6_2),.clk(gclk));
	jdff dff_B_kHfSLF8B6_2(.din(w_dff_B_cX9Q2pET6_2),.dout(w_dff_B_kHfSLF8B6_2),.clk(gclk));
	jdff dff_B_D5kFYsyw9_2(.din(w_dff_B_kHfSLF8B6_2),.dout(w_dff_B_D5kFYsyw9_2),.clk(gclk));
	jdff dff_B_rDwStpPN5_2(.din(w_dff_B_D5kFYsyw9_2),.dout(w_dff_B_rDwStpPN5_2),.clk(gclk));
	jdff dff_B_vF3hEizx7_2(.din(w_dff_B_rDwStpPN5_2),.dout(w_dff_B_vF3hEizx7_2),.clk(gclk));
	jdff dff_B_AI8jw5il9_2(.din(w_dff_B_vF3hEizx7_2),.dout(w_dff_B_AI8jw5il9_2),.clk(gclk));
	jdff dff_B_lIeYby8V8_2(.din(w_dff_B_AI8jw5il9_2),.dout(w_dff_B_lIeYby8V8_2),.clk(gclk));
	jdff dff_B_nw4ESBAx9_2(.din(w_dff_B_lIeYby8V8_2),.dout(w_dff_B_nw4ESBAx9_2),.clk(gclk));
	jdff dff_B_6qvCuHvB9_2(.din(w_dff_B_nw4ESBAx9_2),.dout(w_dff_B_6qvCuHvB9_2),.clk(gclk));
	jdff dff_B_bTUEaydP0_2(.din(w_dff_B_6qvCuHvB9_2),.dout(w_dff_B_bTUEaydP0_2),.clk(gclk));
	jdff dff_B_9TVk05s40_2(.din(w_dff_B_bTUEaydP0_2),.dout(w_dff_B_9TVk05s40_2),.clk(gclk));
	jdff dff_B_IMPzkTTk6_2(.din(w_dff_B_9TVk05s40_2),.dout(w_dff_B_IMPzkTTk6_2),.clk(gclk));
	jdff dff_B_IciobQ9S3_2(.din(w_dff_B_IMPzkTTk6_2),.dout(w_dff_B_IciobQ9S3_2),.clk(gclk));
	jdff dff_B_olRmnmKX5_2(.din(w_dff_B_IciobQ9S3_2),.dout(w_dff_B_olRmnmKX5_2),.clk(gclk));
	jdff dff_B_D0Fo8iyw5_2(.din(w_dff_B_olRmnmKX5_2),.dout(w_dff_B_D0Fo8iyw5_2),.clk(gclk));
	jdff dff_B_XZfn5ScZ8_2(.din(w_dff_B_D0Fo8iyw5_2),.dout(w_dff_B_XZfn5ScZ8_2),.clk(gclk));
	jdff dff_B_xGr38sAj9_2(.din(w_dff_B_XZfn5ScZ8_2),.dout(w_dff_B_xGr38sAj9_2),.clk(gclk));
	jdff dff_B_iRazComT1_2(.din(w_dff_B_xGr38sAj9_2),.dout(w_dff_B_iRazComT1_2),.clk(gclk));
	jdff dff_B_6LfYAUrp2_2(.din(w_dff_B_iRazComT1_2),.dout(w_dff_B_6LfYAUrp2_2),.clk(gclk));
	jdff dff_B_tMTFfhlg1_2(.din(w_dff_B_6LfYAUrp2_2),.dout(w_dff_B_tMTFfhlg1_2),.clk(gclk));
	jdff dff_B_KIPhj9SK0_2(.din(w_dff_B_tMTFfhlg1_2),.dout(w_dff_B_KIPhj9SK0_2),.clk(gclk));
	jdff dff_B_B4Ub5xnK4_2(.din(w_dff_B_KIPhj9SK0_2),.dout(w_dff_B_B4Ub5xnK4_2),.clk(gclk));
	jdff dff_B_hVnXmHOG6_2(.din(w_dff_B_B4Ub5xnK4_2),.dout(w_dff_B_hVnXmHOG6_2),.clk(gclk));
	jdff dff_B_Szd2QzRz4_2(.din(w_dff_B_hVnXmHOG6_2),.dout(w_dff_B_Szd2QzRz4_2),.clk(gclk));
	jdff dff_B_wK63IE4k2_2(.din(w_dff_B_Szd2QzRz4_2),.dout(w_dff_B_wK63IE4k2_2),.clk(gclk));
	jdff dff_B_cN1DcKVD7_2(.din(n1316),.dout(w_dff_B_cN1DcKVD7_2),.clk(gclk));
	jdff dff_B_ImpNrGtm4_1(.din(n1264),.dout(w_dff_B_ImpNrGtm4_1),.clk(gclk));
	jdff dff_B_tupij4Nv5_2(.din(n1173),.dout(w_dff_B_tupij4Nv5_2),.clk(gclk));
	jdff dff_B_sHKsTPx80_2(.din(w_dff_B_tupij4Nv5_2),.dout(w_dff_B_sHKsTPx80_2),.clk(gclk));
	jdff dff_B_6vke0d8c0_2(.din(w_dff_B_sHKsTPx80_2),.dout(w_dff_B_6vke0d8c0_2),.clk(gclk));
	jdff dff_B_VLIgPtqg2_2(.din(w_dff_B_6vke0d8c0_2),.dout(w_dff_B_VLIgPtqg2_2),.clk(gclk));
	jdff dff_B_yISFIlMI7_2(.din(w_dff_B_VLIgPtqg2_2),.dout(w_dff_B_yISFIlMI7_2),.clk(gclk));
	jdff dff_B_vCX7vl4r7_2(.din(w_dff_B_yISFIlMI7_2),.dout(w_dff_B_vCX7vl4r7_2),.clk(gclk));
	jdff dff_B_ROeHYyK89_2(.din(w_dff_B_vCX7vl4r7_2),.dout(w_dff_B_ROeHYyK89_2),.clk(gclk));
	jdff dff_B_j8JRjkZw1_2(.din(w_dff_B_ROeHYyK89_2),.dout(w_dff_B_j8JRjkZw1_2),.clk(gclk));
	jdff dff_B_OWIr4lcW8_2(.din(w_dff_B_j8JRjkZw1_2),.dout(w_dff_B_OWIr4lcW8_2),.clk(gclk));
	jdff dff_B_ihePhkrq9_2(.din(w_dff_B_OWIr4lcW8_2),.dout(w_dff_B_ihePhkrq9_2),.clk(gclk));
	jdff dff_B_GVr11g0U7_2(.din(w_dff_B_ihePhkrq9_2),.dout(w_dff_B_GVr11g0U7_2),.clk(gclk));
	jdff dff_B_TvSbY1429_2(.din(w_dff_B_GVr11g0U7_2),.dout(w_dff_B_TvSbY1429_2),.clk(gclk));
	jdff dff_B_KPrejBD39_2(.din(w_dff_B_TvSbY1429_2),.dout(w_dff_B_KPrejBD39_2),.clk(gclk));
	jdff dff_B_wBdZKpMH2_2(.din(w_dff_B_KPrejBD39_2),.dout(w_dff_B_wBdZKpMH2_2),.clk(gclk));
	jdff dff_B_AvTnVext5_2(.din(w_dff_B_wBdZKpMH2_2),.dout(w_dff_B_AvTnVext5_2),.clk(gclk));
	jdff dff_B_P9gTtpwK6_2(.din(w_dff_B_AvTnVext5_2),.dout(w_dff_B_P9gTtpwK6_2),.clk(gclk));
	jdff dff_B_ov0xG9pm8_2(.din(w_dff_B_P9gTtpwK6_2),.dout(w_dff_B_ov0xG9pm8_2),.clk(gclk));
	jdff dff_B_VGXCQCUd0_2(.din(w_dff_B_ov0xG9pm8_2),.dout(w_dff_B_VGXCQCUd0_2),.clk(gclk));
	jdff dff_B_kXYsHOV08_2(.din(w_dff_B_VGXCQCUd0_2),.dout(w_dff_B_kXYsHOV08_2),.clk(gclk));
	jdff dff_B_1MMKTMfP2_2(.din(w_dff_B_kXYsHOV08_2),.dout(w_dff_B_1MMKTMfP2_2),.clk(gclk));
	jdff dff_B_Of4YOxQd3_2(.din(w_dff_B_1MMKTMfP2_2),.dout(w_dff_B_Of4YOxQd3_2),.clk(gclk));
	jdff dff_B_4A2sPORL6_2(.din(w_dff_B_Of4YOxQd3_2),.dout(w_dff_B_4A2sPORL6_2),.clk(gclk));
	jdff dff_B_fIhypljW9_2(.din(w_dff_B_4A2sPORL6_2),.dout(w_dff_B_fIhypljW9_2),.clk(gclk));
	jdff dff_B_jWP9SUZ06_2(.din(w_dff_B_fIhypljW9_2),.dout(w_dff_B_jWP9SUZ06_2),.clk(gclk));
	jdff dff_B_D5aerA2U8_2(.din(w_dff_B_jWP9SUZ06_2),.dout(w_dff_B_D5aerA2U8_2),.clk(gclk));
	jdff dff_B_CLOCFoYJ4_2(.din(w_dff_B_D5aerA2U8_2),.dout(w_dff_B_CLOCFoYJ4_2),.clk(gclk));
	jdff dff_B_9hCzTUK42_2(.din(w_dff_B_CLOCFoYJ4_2),.dout(w_dff_B_9hCzTUK42_2),.clk(gclk));
	jdff dff_B_fFiVH1kG4_2(.din(w_dff_B_9hCzTUK42_2),.dout(w_dff_B_fFiVH1kG4_2),.clk(gclk));
	jdff dff_B_FKVraEVe9_2(.din(w_dff_B_fFiVH1kG4_2),.dout(w_dff_B_FKVraEVe9_2),.clk(gclk));
	jdff dff_B_r3FGNd2r9_2(.din(w_dff_B_FKVraEVe9_2),.dout(w_dff_B_r3FGNd2r9_2),.clk(gclk));
	jdff dff_B_2Xm7Rslv6_2(.din(w_dff_B_r3FGNd2r9_2),.dout(w_dff_B_2Xm7Rslv6_2),.clk(gclk));
	jdff dff_B_HT9VLYAA6_2(.din(w_dff_B_2Xm7Rslv6_2),.dout(w_dff_B_HT9VLYAA6_2),.clk(gclk));
	jdff dff_B_iArFbLF42_2(.din(w_dff_B_HT9VLYAA6_2),.dout(w_dff_B_iArFbLF42_2),.clk(gclk));
	jdff dff_B_X8PXlsSu2_2(.din(n1225),.dout(w_dff_B_X8PXlsSu2_2),.clk(gclk));
	jdff dff_B_0sSPHn4O8_1(.din(n1174),.dout(w_dff_B_0sSPHn4O8_1),.clk(gclk));
	jdff dff_B_c3Vd6GrN3_2(.din(n1069),.dout(w_dff_B_c3Vd6GrN3_2),.clk(gclk));
	jdff dff_B_lf3zomKh8_2(.din(w_dff_B_c3Vd6GrN3_2),.dout(w_dff_B_lf3zomKh8_2),.clk(gclk));
	jdff dff_B_FqoalI5p1_2(.din(w_dff_B_lf3zomKh8_2),.dout(w_dff_B_FqoalI5p1_2),.clk(gclk));
	jdff dff_B_BUS2HOza9_2(.din(w_dff_B_FqoalI5p1_2),.dout(w_dff_B_BUS2HOza9_2),.clk(gclk));
	jdff dff_B_NqlTAb3O0_2(.din(w_dff_B_BUS2HOza9_2),.dout(w_dff_B_NqlTAb3O0_2),.clk(gclk));
	jdff dff_B_aJA2haG50_2(.din(w_dff_B_NqlTAb3O0_2),.dout(w_dff_B_aJA2haG50_2),.clk(gclk));
	jdff dff_B_MXv2KJ0H9_2(.din(w_dff_B_aJA2haG50_2),.dout(w_dff_B_MXv2KJ0H9_2),.clk(gclk));
	jdff dff_B_5dIt3qRJ9_2(.din(w_dff_B_MXv2KJ0H9_2),.dout(w_dff_B_5dIt3qRJ9_2),.clk(gclk));
	jdff dff_B_tzWFpcnl3_2(.din(w_dff_B_5dIt3qRJ9_2),.dout(w_dff_B_tzWFpcnl3_2),.clk(gclk));
	jdff dff_B_UE1XYbw51_2(.din(w_dff_B_tzWFpcnl3_2),.dout(w_dff_B_UE1XYbw51_2),.clk(gclk));
	jdff dff_B_M4LX79iD3_2(.din(w_dff_B_UE1XYbw51_2),.dout(w_dff_B_M4LX79iD3_2),.clk(gclk));
	jdff dff_B_pMOogKxM1_2(.din(w_dff_B_M4LX79iD3_2),.dout(w_dff_B_pMOogKxM1_2),.clk(gclk));
	jdff dff_B_jQLXLeSi6_2(.din(w_dff_B_pMOogKxM1_2),.dout(w_dff_B_jQLXLeSi6_2),.clk(gclk));
	jdff dff_B_m0zmUcfS8_2(.din(w_dff_B_jQLXLeSi6_2),.dout(w_dff_B_m0zmUcfS8_2),.clk(gclk));
	jdff dff_B_Umklu2qo4_2(.din(w_dff_B_m0zmUcfS8_2),.dout(w_dff_B_Umklu2qo4_2),.clk(gclk));
	jdff dff_B_iIqrvonK1_2(.din(w_dff_B_Umklu2qo4_2),.dout(w_dff_B_iIqrvonK1_2),.clk(gclk));
	jdff dff_B_pRCVsK5J0_2(.din(w_dff_B_iIqrvonK1_2),.dout(w_dff_B_pRCVsK5J0_2),.clk(gclk));
	jdff dff_B_FNJztTfC8_2(.din(w_dff_B_pRCVsK5J0_2),.dout(w_dff_B_FNJztTfC8_2),.clk(gclk));
	jdff dff_B_prQxtbgJ4_2(.din(w_dff_B_FNJztTfC8_2),.dout(w_dff_B_prQxtbgJ4_2),.clk(gclk));
	jdff dff_B_EyfdXWdF9_2(.din(w_dff_B_prQxtbgJ4_2),.dout(w_dff_B_EyfdXWdF9_2),.clk(gclk));
	jdff dff_B_MLxzRiDT8_2(.din(w_dff_B_EyfdXWdF9_2),.dout(w_dff_B_MLxzRiDT8_2),.clk(gclk));
	jdff dff_B_Scpb4JCl2_2(.din(w_dff_B_MLxzRiDT8_2),.dout(w_dff_B_Scpb4JCl2_2),.clk(gclk));
	jdff dff_B_al9HdKIK0_2(.din(w_dff_B_Scpb4JCl2_2),.dout(w_dff_B_al9HdKIK0_2),.clk(gclk));
	jdff dff_B_JbQX7Hbj0_2(.din(w_dff_B_al9HdKIK0_2),.dout(w_dff_B_JbQX7Hbj0_2),.clk(gclk));
	jdff dff_B_BhDPqHiN3_2(.din(w_dff_B_JbQX7Hbj0_2),.dout(w_dff_B_BhDPqHiN3_2),.clk(gclk));
	jdff dff_B_KCug5COe5_2(.din(w_dff_B_BhDPqHiN3_2),.dout(w_dff_B_KCug5COe5_2),.clk(gclk));
	jdff dff_B_vf3dco6h5_2(.din(w_dff_B_KCug5COe5_2),.dout(w_dff_B_vf3dco6h5_2),.clk(gclk));
	jdff dff_B_MlpgTR5Q3_2(.din(w_dff_B_vf3dco6h5_2),.dout(w_dff_B_MlpgTR5Q3_2),.clk(gclk));
	jdff dff_B_MjcPfnJp5_2(.din(w_dff_B_MlpgTR5Q3_2),.dout(w_dff_B_MjcPfnJp5_2),.clk(gclk));
	jdff dff_B_tE3GPyAT6_2(.din(w_dff_B_MjcPfnJp5_2),.dout(w_dff_B_tE3GPyAT6_2),.clk(gclk));
	jdff dff_B_Ey1mCoSe0_2(.din(n1127),.dout(w_dff_B_Ey1mCoSe0_2),.clk(gclk));
	jdff dff_B_EU9fSBA64_1(.din(n1070),.dout(w_dff_B_EU9fSBA64_1),.clk(gclk));
	jdff dff_B_msWHd3oh5_2(.din(n971),.dout(w_dff_B_msWHd3oh5_2),.clk(gclk));
	jdff dff_B_Neyv2mKd0_2(.din(w_dff_B_msWHd3oh5_2),.dout(w_dff_B_Neyv2mKd0_2),.clk(gclk));
	jdff dff_B_R6CN6o1L5_2(.din(w_dff_B_Neyv2mKd0_2),.dout(w_dff_B_R6CN6o1L5_2),.clk(gclk));
	jdff dff_B_qzQiVGiQ8_2(.din(w_dff_B_R6CN6o1L5_2),.dout(w_dff_B_qzQiVGiQ8_2),.clk(gclk));
	jdff dff_B_EKLGHIcV9_2(.din(w_dff_B_qzQiVGiQ8_2),.dout(w_dff_B_EKLGHIcV9_2),.clk(gclk));
	jdff dff_B_plfNoSIO3_2(.din(w_dff_B_EKLGHIcV9_2),.dout(w_dff_B_plfNoSIO3_2),.clk(gclk));
	jdff dff_B_1twOcQB14_2(.din(w_dff_B_plfNoSIO3_2),.dout(w_dff_B_1twOcQB14_2),.clk(gclk));
	jdff dff_B_DOMXe3GP5_2(.din(w_dff_B_1twOcQB14_2),.dout(w_dff_B_DOMXe3GP5_2),.clk(gclk));
	jdff dff_B_BPq00AG38_2(.din(w_dff_B_DOMXe3GP5_2),.dout(w_dff_B_BPq00AG38_2),.clk(gclk));
	jdff dff_B_OwlEvNCk5_2(.din(w_dff_B_BPq00AG38_2),.dout(w_dff_B_OwlEvNCk5_2),.clk(gclk));
	jdff dff_B_9691XIaT6_2(.din(w_dff_B_OwlEvNCk5_2),.dout(w_dff_B_9691XIaT6_2),.clk(gclk));
	jdff dff_B_Evd8MDCF3_2(.din(w_dff_B_9691XIaT6_2),.dout(w_dff_B_Evd8MDCF3_2),.clk(gclk));
	jdff dff_B_EWB6sXBG3_2(.din(w_dff_B_Evd8MDCF3_2),.dout(w_dff_B_EWB6sXBG3_2),.clk(gclk));
	jdff dff_B_7kx7y9Xv3_2(.din(w_dff_B_EWB6sXBG3_2),.dout(w_dff_B_7kx7y9Xv3_2),.clk(gclk));
	jdff dff_B_7YH5rV9f4_2(.din(w_dff_B_7kx7y9Xv3_2),.dout(w_dff_B_7YH5rV9f4_2),.clk(gclk));
	jdff dff_B_ol5XeFAm4_2(.din(w_dff_B_7YH5rV9f4_2),.dout(w_dff_B_ol5XeFAm4_2),.clk(gclk));
	jdff dff_B_nxNUkvJm1_2(.din(w_dff_B_ol5XeFAm4_2),.dout(w_dff_B_nxNUkvJm1_2),.clk(gclk));
	jdff dff_B_HHso2Rpj0_2(.din(w_dff_B_nxNUkvJm1_2),.dout(w_dff_B_HHso2Rpj0_2),.clk(gclk));
	jdff dff_B_W0w5z7bF8_2(.din(w_dff_B_HHso2Rpj0_2),.dout(w_dff_B_W0w5z7bF8_2),.clk(gclk));
	jdff dff_B_jTzzGAYl7_2(.din(w_dff_B_W0w5z7bF8_2),.dout(w_dff_B_jTzzGAYl7_2),.clk(gclk));
	jdff dff_B_Xuak1bne9_2(.din(w_dff_B_jTzzGAYl7_2),.dout(w_dff_B_Xuak1bne9_2),.clk(gclk));
	jdff dff_B_Y4K0I4uD3_2(.din(w_dff_B_Xuak1bne9_2),.dout(w_dff_B_Y4K0I4uD3_2),.clk(gclk));
	jdff dff_B_vYRFEYbL2_2(.din(w_dff_B_Y4K0I4uD3_2),.dout(w_dff_B_vYRFEYbL2_2),.clk(gclk));
	jdff dff_B_IpURNv8y7_2(.din(w_dff_B_vYRFEYbL2_2),.dout(w_dff_B_IpURNv8y7_2),.clk(gclk));
	jdff dff_B_P3FSdtuF0_2(.din(w_dff_B_IpURNv8y7_2),.dout(w_dff_B_P3FSdtuF0_2),.clk(gclk));
	jdff dff_B_6GbxEZyg9_2(.din(w_dff_B_P3FSdtuF0_2),.dout(w_dff_B_6GbxEZyg9_2),.clk(gclk));
	jdff dff_B_9B0pqAp15_2(.din(w_dff_B_6GbxEZyg9_2),.dout(w_dff_B_9B0pqAp15_2),.clk(gclk));
	jdff dff_B_odIEMLG73_2(.din(n1022),.dout(w_dff_B_odIEMLG73_2),.clk(gclk));
	jdff dff_B_P00V99xF6_1(.din(n972),.dout(w_dff_B_P00V99xF6_1),.clk(gclk));
	jdff dff_B_WJAPKH9r4_2(.din(n866),.dout(w_dff_B_WJAPKH9r4_2),.clk(gclk));
	jdff dff_B_Be2y1eLw1_2(.din(w_dff_B_WJAPKH9r4_2),.dout(w_dff_B_Be2y1eLw1_2),.clk(gclk));
	jdff dff_B_PP4BbTAx4_2(.din(w_dff_B_Be2y1eLw1_2),.dout(w_dff_B_PP4BbTAx4_2),.clk(gclk));
	jdff dff_B_knzvl6E08_2(.din(w_dff_B_PP4BbTAx4_2),.dout(w_dff_B_knzvl6E08_2),.clk(gclk));
	jdff dff_B_4SrQ0URV1_2(.din(w_dff_B_knzvl6E08_2),.dout(w_dff_B_4SrQ0URV1_2),.clk(gclk));
	jdff dff_B_yAIpMIn73_2(.din(w_dff_B_4SrQ0URV1_2),.dout(w_dff_B_yAIpMIn73_2),.clk(gclk));
	jdff dff_B_UfsHC1C33_2(.din(w_dff_B_yAIpMIn73_2),.dout(w_dff_B_UfsHC1C33_2),.clk(gclk));
	jdff dff_B_5deEPxUu2_2(.din(w_dff_B_UfsHC1C33_2),.dout(w_dff_B_5deEPxUu2_2),.clk(gclk));
	jdff dff_B_ZQlbNdte0_2(.din(w_dff_B_5deEPxUu2_2),.dout(w_dff_B_ZQlbNdte0_2),.clk(gclk));
	jdff dff_B_8ganj8Pt3_2(.din(w_dff_B_ZQlbNdte0_2),.dout(w_dff_B_8ganj8Pt3_2),.clk(gclk));
	jdff dff_B_wLDMP53B3_2(.din(w_dff_B_8ganj8Pt3_2),.dout(w_dff_B_wLDMP53B3_2),.clk(gclk));
	jdff dff_B_QC9oHw9t2_2(.din(w_dff_B_wLDMP53B3_2),.dout(w_dff_B_QC9oHw9t2_2),.clk(gclk));
	jdff dff_B_tkkr1hc26_2(.din(w_dff_B_QC9oHw9t2_2),.dout(w_dff_B_tkkr1hc26_2),.clk(gclk));
	jdff dff_B_PBbUxTOK4_2(.din(w_dff_B_tkkr1hc26_2),.dout(w_dff_B_PBbUxTOK4_2),.clk(gclk));
	jdff dff_B_GheVLLBZ8_2(.din(w_dff_B_PBbUxTOK4_2),.dout(w_dff_B_GheVLLBZ8_2),.clk(gclk));
	jdff dff_B_ygMLiikt8_2(.din(w_dff_B_GheVLLBZ8_2),.dout(w_dff_B_ygMLiikt8_2),.clk(gclk));
	jdff dff_B_q5NYwUsE9_2(.din(w_dff_B_ygMLiikt8_2),.dout(w_dff_B_q5NYwUsE9_2),.clk(gclk));
	jdff dff_B_3uzTq3Az3_2(.din(w_dff_B_q5NYwUsE9_2),.dout(w_dff_B_3uzTq3Az3_2),.clk(gclk));
	jdff dff_B_Rjet8Wn75_2(.din(w_dff_B_3uzTq3Az3_2),.dout(w_dff_B_Rjet8Wn75_2),.clk(gclk));
	jdff dff_B_J1iPLDCX0_2(.din(w_dff_B_Rjet8Wn75_2),.dout(w_dff_B_J1iPLDCX0_2),.clk(gclk));
	jdff dff_B_eF9Tk66p4_2(.din(w_dff_B_J1iPLDCX0_2),.dout(w_dff_B_eF9Tk66p4_2),.clk(gclk));
	jdff dff_B_47ZRFloy8_2(.din(w_dff_B_eF9Tk66p4_2),.dout(w_dff_B_47ZRFloy8_2),.clk(gclk));
	jdff dff_B_H2RfDcbU6_2(.din(w_dff_B_47ZRFloy8_2),.dout(w_dff_B_H2RfDcbU6_2),.clk(gclk));
	jdff dff_B_W4fjIvWG8_2(.din(w_dff_B_H2RfDcbU6_2),.dout(w_dff_B_W4fjIvWG8_2),.clk(gclk));
	jdff dff_B_SqSzmfJI2_2(.din(n917),.dout(w_dff_B_SqSzmfJI2_2),.clk(gclk));
	jdff dff_B_FwUjwLpg3_1(.din(n867),.dout(w_dff_B_FwUjwLpg3_1),.clk(gclk));
	jdff dff_B_sbiRgiuq9_2(.din(n767),.dout(w_dff_B_sbiRgiuq9_2),.clk(gclk));
	jdff dff_B_2qFNidnc3_2(.din(w_dff_B_sbiRgiuq9_2),.dout(w_dff_B_2qFNidnc3_2),.clk(gclk));
	jdff dff_B_s8IYWgUJ6_2(.din(w_dff_B_2qFNidnc3_2),.dout(w_dff_B_s8IYWgUJ6_2),.clk(gclk));
	jdff dff_B_bfVDU8DR9_2(.din(w_dff_B_s8IYWgUJ6_2),.dout(w_dff_B_bfVDU8DR9_2),.clk(gclk));
	jdff dff_B_Zsg35E7T0_2(.din(w_dff_B_bfVDU8DR9_2),.dout(w_dff_B_Zsg35E7T0_2),.clk(gclk));
	jdff dff_B_NIuS8Gao2_2(.din(w_dff_B_Zsg35E7T0_2),.dout(w_dff_B_NIuS8Gao2_2),.clk(gclk));
	jdff dff_B_2R3SzqrG6_2(.din(w_dff_B_NIuS8Gao2_2),.dout(w_dff_B_2R3SzqrG6_2),.clk(gclk));
	jdff dff_B_RnlveGLs4_2(.din(w_dff_B_2R3SzqrG6_2),.dout(w_dff_B_RnlveGLs4_2),.clk(gclk));
	jdff dff_B_yKvtNNbC3_2(.din(w_dff_B_RnlveGLs4_2),.dout(w_dff_B_yKvtNNbC3_2),.clk(gclk));
	jdff dff_B_nJLfIOD81_2(.din(w_dff_B_yKvtNNbC3_2),.dout(w_dff_B_nJLfIOD81_2),.clk(gclk));
	jdff dff_B_XJEfy2eA2_2(.din(w_dff_B_nJLfIOD81_2),.dout(w_dff_B_XJEfy2eA2_2),.clk(gclk));
	jdff dff_B_MjUiPWYF1_2(.din(w_dff_B_XJEfy2eA2_2),.dout(w_dff_B_MjUiPWYF1_2),.clk(gclk));
	jdff dff_B_2xI6hlF41_2(.din(w_dff_B_MjUiPWYF1_2),.dout(w_dff_B_2xI6hlF41_2),.clk(gclk));
	jdff dff_B_rSF8CSo16_2(.din(w_dff_B_2xI6hlF41_2),.dout(w_dff_B_rSF8CSo16_2),.clk(gclk));
	jdff dff_B_W0mRZfbF5_2(.din(w_dff_B_rSF8CSo16_2),.dout(w_dff_B_W0mRZfbF5_2),.clk(gclk));
	jdff dff_B_B6eRyLYW2_2(.din(w_dff_B_W0mRZfbF5_2),.dout(w_dff_B_B6eRyLYW2_2),.clk(gclk));
	jdff dff_B_kEoxd8r45_2(.din(w_dff_B_B6eRyLYW2_2),.dout(w_dff_B_kEoxd8r45_2),.clk(gclk));
	jdff dff_B_DNoRZaMs0_2(.din(w_dff_B_kEoxd8r45_2),.dout(w_dff_B_DNoRZaMs0_2),.clk(gclk));
	jdff dff_B_amQhJ1rp8_2(.din(w_dff_B_DNoRZaMs0_2),.dout(w_dff_B_amQhJ1rp8_2),.clk(gclk));
	jdff dff_B_hfBLVgxm8_2(.din(w_dff_B_amQhJ1rp8_2),.dout(w_dff_B_hfBLVgxm8_2),.clk(gclk));
	jdff dff_B_NJq9Mwmv8_2(.din(w_dff_B_hfBLVgxm8_2),.dout(w_dff_B_NJq9Mwmv8_2),.clk(gclk));
	jdff dff_B_9rJcZFO74_2(.din(n811),.dout(w_dff_B_9rJcZFO74_2),.clk(gclk));
	jdff dff_B_aLCONApw9_1(.din(n768),.dout(w_dff_B_aLCONApw9_1),.clk(gclk));
	jdff dff_B_eTKLcG3n9_2(.din(n674),.dout(w_dff_B_eTKLcG3n9_2),.clk(gclk));
	jdff dff_B_R6UHHqcU8_2(.din(w_dff_B_eTKLcG3n9_2),.dout(w_dff_B_R6UHHqcU8_2),.clk(gclk));
	jdff dff_B_hXhFr7N95_2(.din(w_dff_B_R6UHHqcU8_2),.dout(w_dff_B_hXhFr7N95_2),.clk(gclk));
	jdff dff_B_NRLcLJR19_2(.din(w_dff_B_hXhFr7N95_2),.dout(w_dff_B_NRLcLJR19_2),.clk(gclk));
	jdff dff_B_dUEnkPYr7_2(.din(w_dff_B_NRLcLJR19_2),.dout(w_dff_B_dUEnkPYr7_2),.clk(gclk));
	jdff dff_B_XLvcjCws7_2(.din(w_dff_B_dUEnkPYr7_2),.dout(w_dff_B_XLvcjCws7_2),.clk(gclk));
	jdff dff_B_icyC7InA1_2(.din(w_dff_B_XLvcjCws7_2),.dout(w_dff_B_icyC7InA1_2),.clk(gclk));
	jdff dff_B_Uqk8bYov4_2(.din(w_dff_B_icyC7InA1_2),.dout(w_dff_B_Uqk8bYov4_2),.clk(gclk));
	jdff dff_B_MpLiHoPy2_2(.din(w_dff_B_Uqk8bYov4_2),.dout(w_dff_B_MpLiHoPy2_2),.clk(gclk));
	jdff dff_B_F2gVclQR0_2(.din(w_dff_B_MpLiHoPy2_2),.dout(w_dff_B_F2gVclQR0_2),.clk(gclk));
	jdff dff_B_DQ9DLNxE3_2(.din(w_dff_B_F2gVclQR0_2),.dout(w_dff_B_DQ9DLNxE3_2),.clk(gclk));
	jdff dff_B_F6QBbcuy4_2(.din(w_dff_B_DQ9DLNxE3_2),.dout(w_dff_B_F6QBbcuy4_2),.clk(gclk));
	jdff dff_B_QjgN8iEH3_2(.din(w_dff_B_F6QBbcuy4_2),.dout(w_dff_B_QjgN8iEH3_2),.clk(gclk));
	jdff dff_B_7TsXYrYs6_2(.din(w_dff_B_QjgN8iEH3_2),.dout(w_dff_B_7TsXYrYs6_2),.clk(gclk));
	jdff dff_B_azhVPQdI9_2(.din(w_dff_B_7TsXYrYs6_2),.dout(w_dff_B_azhVPQdI9_2),.clk(gclk));
	jdff dff_B_hbH2dvgo3_2(.din(w_dff_B_azhVPQdI9_2),.dout(w_dff_B_hbH2dvgo3_2),.clk(gclk));
	jdff dff_B_9lYNUB6v6_2(.din(w_dff_B_hbH2dvgo3_2),.dout(w_dff_B_9lYNUB6v6_2),.clk(gclk));
	jdff dff_B_sWjd90256_2(.din(w_dff_B_9lYNUB6v6_2),.dout(w_dff_B_sWjd90256_2),.clk(gclk));
	jdff dff_B_RHR0rDDN0_2(.din(n711),.dout(w_dff_B_RHR0rDDN0_2),.clk(gclk));
	jdff dff_B_myZc1rch3_1(.din(n675),.dout(w_dff_B_myZc1rch3_1),.clk(gclk));
	jdff dff_B_Wk0729rd9_2(.din(n588),.dout(w_dff_B_Wk0729rd9_2),.clk(gclk));
	jdff dff_B_9j2TjyNq2_2(.din(w_dff_B_Wk0729rd9_2),.dout(w_dff_B_9j2TjyNq2_2),.clk(gclk));
	jdff dff_B_0zH9w3kZ5_2(.din(w_dff_B_9j2TjyNq2_2),.dout(w_dff_B_0zH9w3kZ5_2),.clk(gclk));
	jdff dff_B_hzUDXxsE8_2(.din(w_dff_B_0zH9w3kZ5_2),.dout(w_dff_B_hzUDXxsE8_2),.clk(gclk));
	jdff dff_B_fDnBT49Y9_2(.din(w_dff_B_hzUDXxsE8_2),.dout(w_dff_B_fDnBT49Y9_2),.clk(gclk));
	jdff dff_B_AVfeqjyG7_2(.din(w_dff_B_fDnBT49Y9_2),.dout(w_dff_B_AVfeqjyG7_2),.clk(gclk));
	jdff dff_B_4BuUGYnX4_2(.din(w_dff_B_AVfeqjyG7_2),.dout(w_dff_B_4BuUGYnX4_2),.clk(gclk));
	jdff dff_B_mtqPUI0T1_2(.din(w_dff_B_4BuUGYnX4_2),.dout(w_dff_B_mtqPUI0T1_2),.clk(gclk));
	jdff dff_B_Mpp5fT8p6_2(.din(w_dff_B_mtqPUI0T1_2),.dout(w_dff_B_Mpp5fT8p6_2),.clk(gclk));
	jdff dff_B_TViT5sPd4_2(.din(w_dff_B_Mpp5fT8p6_2),.dout(w_dff_B_TViT5sPd4_2),.clk(gclk));
	jdff dff_B_eQU8pXQN6_2(.din(w_dff_B_TViT5sPd4_2),.dout(w_dff_B_eQU8pXQN6_2),.clk(gclk));
	jdff dff_B_hB9y8UTf7_2(.din(w_dff_B_eQU8pXQN6_2),.dout(w_dff_B_hB9y8UTf7_2),.clk(gclk));
	jdff dff_B_8lRcB4fm6_2(.din(w_dff_B_hB9y8UTf7_2),.dout(w_dff_B_8lRcB4fm6_2),.clk(gclk));
	jdff dff_B_aXuJiYt90_2(.din(w_dff_B_8lRcB4fm6_2),.dout(w_dff_B_aXuJiYt90_2),.clk(gclk));
	jdff dff_B_N4qhkeI07_2(.din(w_dff_B_aXuJiYt90_2),.dout(w_dff_B_N4qhkeI07_2),.clk(gclk));
	jdff dff_B_rldC3BJ47_2(.din(n618),.dout(w_dff_B_rldC3BJ47_2),.clk(gclk));
	jdff dff_B_JXDGhtOe4_1(.din(n589),.dout(w_dff_B_JXDGhtOe4_1),.clk(gclk));
	jdff dff_B_2RydlANO8_2(.din(n509),.dout(w_dff_B_2RydlANO8_2),.clk(gclk));
	jdff dff_B_CIScbIBQ6_2(.din(w_dff_B_2RydlANO8_2),.dout(w_dff_B_CIScbIBQ6_2),.clk(gclk));
	jdff dff_B_zH8a4xVO4_2(.din(w_dff_B_CIScbIBQ6_2),.dout(w_dff_B_zH8a4xVO4_2),.clk(gclk));
	jdff dff_B_sDahNV6J7_2(.din(w_dff_B_zH8a4xVO4_2),.dout(w_dff_B_sDahNV6J7_2),.clk(gclk));
	jdff dff_B_94Su4Wyr7_2(.din(w_dff_B_sDahNV6J7_2),.dout(w_dff_B_94Su4Wyr7_2),.clk(gclk));
	jdff dff_B_RRUJDn0M0_2(.din(w_dff_B_94Su4Wyr7_2),.dout(w_dff_B_RRUJDn0M0_2),.clk(gclk));
	jdff dff_B_PC0IDieh3_2(.din(w_dff_B_RRUJDn0M0_2),.dout(w_dff_B_PC0IDieh3_2),.clk(gclk));
	jdff dff_B_Hd6Dvm0S6_2(.din(w_dff_B_PC0IDieh3_2),.dout(w_dff_B_Hd6Dvm0S6_2),.clk(gclk));
	jdff dff_B_vnDs6X5n0_2(.din(w_dff_B_Hd6Dvm0S6_2),.dout(w_dff_B_vnDs6X5n0_2),.clk(gclk));
	jdff dff_B_SpKWs8qL6_2(.din(w_dff_B_vnDs6X5n0_2),.dout(w_dff_B_SpKWs8qL6_2),.clk(gclk));
	jdff dff_B_deIYh7Pd5_2(.din(w_dff_B_SpKWs8qL6_2),.dout(w_dff_B_deIYh7Pd5_2),.clk(gclk));
	jdff dff_B_StDSFw8h8_2(.din(w_dff_B_deIYh7Pd5_2),.dout(w_dff_B_StDSFw8h8_2),.clk(gclk));
	jdff dff_B_CVnLg0kR4_2(.din(n532),.dout(w_dff_B_CVnLg0kR4_2),.clk(gclk));
	jdff dff_B_fr234X5Q7_1(.din(n510),.dout(w_dff_B_fr234X5Q7_1),.clk(gclk));
	jdff dff_B_6tT9T7Su6_2(.din(n437),.dout(w_dff_B_6tT9T7Su6_2),.clk(gclk));
	jdff dff_B_Wqu20p4v5_2(.din(w_dff_B_6tT9T7Su6_2),.dout(w_dff_B_Wqu20p4v5_2),.clk(gclk));
	jdff dff_B_A8a4HFKX5_2(.din(w_dff_B_Wqu20p4v5_2),.dout(w_dff_B_A8a4HFKX5_2),.clk(gclk));
	jdff dff_B_nnvA88J42_2(.din(w_dff_B_A8a4HFKX5_2),.dout(w_dff_B_nnvA88J42_2),.clk(gclk));
	jdff dff_B_48uXmbWc9_2(.din(w_dff_B_nnvA88J42_2),.dout(w_dff_B_48uXmbWc9_2),.clk(gclk));
	jdff dff_B_8H9EKZis3_2(.din(w_dff_B_48uXmbWc9_2),.dout(w_dff_B_8H9EKZis3_2),.clk(gclk));
	jdff dff_B_hIDVNv4n8_2(.din(w_dff_B_8H9EKZis3_2),.dout(w_dff_B_hIDVNv4n8_2),.clk(gclk));
	jdff dff_B_wmccnfO15_2(.din(w_dff_B_hIDVNv4n8_2),.dout(w_dff_B_wmccnfO15_2),.clk(gclk));
	jdff dff_B_j23U0sOR6_2(.din(w_dff_B_wmccnfO15_2),.dout(w_dff_B_j23U0sOR6_2),.clk(gclk));
	jdff dff_B_DENUeDNg6_2(.din(n453),.dout(w_dff_B_DENUeDNg6_2),.clk(gclk));
	jdff dff_B_ugK7QYqi7_2(.din(w_dff_B_DENUeDNg6_2),.dout(w_dff_B_ugK7QYqi7_2),.clk(gclk));
	jdff dff_B_MYapCTdd2_1(.din(n438),.dout(w_dff_B_MYapCTdd2_1),.clk(gclk));
	jdff dff_B_xgmph9Mx5_1(.din(w_dff_B_MYapCTdd2_1),.dout(w_dff_B_xgmph9Mx5_1),.clk(gclk));
	jdff dff_B_9kdLMMw17_1(.din(w_dff_B_xgmph9Mx5_1),.dout(w_dff_B_9kdLMMw17_1),.clk(gclk));
	jdff dff_B_ou4UUd8m9_1(.din(w_dff_B_9kdLMMw17_1),.dout(w_dff_B_ou4UUd8m9_1),.clk(gclk));
	jdff dff_B_Eg0G2rQK4_1(.din(w_dff_B_ou4UUd8m9_1),.dout(w_dff_B_Eg0G2rQK4_1),.clk(gclk));
	jdff dff_B_zin7EFie7_1(.din(w_dff_B_Eg0G2rQK4_1),.dout(w_dff_B_zin7EFie7_1),.clk(gclk));
	jdff dff_B_ayM6OZZT9_0(.din(n381),.dout(w_dff_B_ayM6OZZT9_0),.clk(gclk));
	jdff dff_B_L41QrBO30_0(.din(w_dff_B_ayM6OZZT9_0),.dout(w_dff_B_L41QrBO30_0),.clk(gclk));
	jdff dff_A_TmYr42cC0_0(.dout(w_n380_0[0]),.din(w_dff_A_TmYr42cC0_0),.clk(gclk));
	jdff dff_A_v2T2r6Bw5_0(.dout(w_dff_A_TmYr42cC0_0),.din(w_dff_A_v2T2r6Bw5_0),.clk(gclk));
	jdff dff_A_CFnGIAnQ4_0(.dout(w_dff_A_v2T2r6Bw5_0),.din(w_dff_A_CFnGIAnQ4_0),.clk(gclk));
	jdff dff_B_AuDEaiwK0_1(.din(n374),.dout(w_dff_B_AuDEaiwK0_1),.clk(gclk));
	jdff dff_A_CWv4PehF4_0(.dout(w_n314_0[0]),.din(w_dff_A_CWv4PehF4_0),.clk(gclk));
	jdff dff_A_PldyxTtr0_1(.dout(w_n314_0[1]),.din(w_dff_A_PldyxTtr0_1),.clk(gclk));
	jdff dff_A_IQZnHAAl3_1(.dout(w_dff_A_PldyxTtr0_1),.din(w_dff_A_IQZnHAAl3_1),.clk(gclk));
	jdff dff_A_jlCOkuN10_1(.dout(w_n372_0[1]),.din(w_dff_A_jlCOkuN10_1),.clk(gclk));
	jdff dff_A_Vzuu0Vkz3_1(.dout(w_dff_A_jlCOkuN10_1),.din(w_dff_A_Vzuu0Vkz3_1),.clk(gclk));
	jdff dff_A_5iOY39rK3_1(.dout(w_dff_A_Vzuu0Vkz3_1),.din(w_dff_A_5iOY39rK3_1),.clk(gclk));
	jdff dff_A_fYxLTpdA0_1(.dout(w_dff_A_5iOY39rK3_1),.din(w_dff_A_fYxLTpdA0_1),.clk(gclk));
	jdff dff_A_vkF2PkVD2_1(.dout(w_dff_A_fYxLTpdA0_1),.din(w_dff_A_vkF2PkVD2_1),.clk(gclk));
	jdff dff_A_AlngDwTI8_1(.dout(w_dff_A_vkF2PkVD2_1),.din(w_dff_A_AlngDwTI8_1),.clk(gclk));
	jdff dff_B_tmATA0839_2(.din(n1627),.dout(w_dff_B_tmATA0839_2),.clk(gclk));
	jdff dff_B_qO9LQxKl1_2(.din(w_dff_B_tmATA0839_2),.dout(w_dff_B_qO9LQxKl1_2),.clk(gclk));
	jdff dff_B_mP2VrqKQ6_1(.din(n1625),.dout(w_dff_B_mP2VrqKQ6_1),.clk(gclk));
	jdff dff_B_plqLQFNf4_2(.din(n1566),.dout(w_dff_B_plqLQFNf4_2),.clk(gclk));
	jdff dff_B_FSU4Fl4o1_2(.din(w_dff_B_plqLQFNf4_2),.dout(w_dff_B_FSU4Fl4o1_2),.clk(gclk));
	jdff dff_B_YCffW1NN1_2(.din(w_dff_B_FSU4Fl4o1_2),.dout(w_dff_B_YCffW1NN1_2),.clk(gclk));
	jdff dff_B_tnMY8Ikd0_2(.din(w_dff_B_YCffW1NN1_2),.dout(w_dff_B_tnMY8Ikd0_2),.clk(gclk));
	jdff dff_B_aRbZ0vuq7_2(.din(w_dff_B_tnMY8Ikd0_2),.dout(w_dff_B_aRbZ0vuq7_2),.clk(gclk));
	jdff dff_B_XjtbQkA16_2(.din(w_dff_B_aRbZ0vuq7_2),.dout(w_dff_B_XjtbQkA16_2),.clk(gclk));
	jdff dff_B_SZmuMXNF5_2(.din(w_dff_B_XjtbQkA16_2),.dout(w_dff_B_SZmuMXNF5_2),.clk(gclk));
	jdff dff_B_8NpBifyg5_2(.din(w_dff_B_SZmuMXNF5_2),.dout(w_dff_B_8NpBifyg5_2),.clk(gclk));
	jdff dff_B_EmYtTHYT5_2(.din(w_dff_B_8NpBifyg5_2),.dout(w_dff_B_EmYtTHYT5_2),.clk(gclk));
	jdff dff_B_QWZjE07A5_2(.din(w_dff_B_EmYtTHYT5_2),.dout(w_dff_B_QWZjE07A5_2),.clk(gclk));
	jdff dff_B_48xUDhoj6_2(.din(w_dff_B_QWZjE07A5_2),.dout(w_dff_B_48xUDhoj6_2),.clk(gclk));
	jdff dff_B_Yh5tGfSY6_2(.din(w_dff_B_48xUDhoj6_2),.dout(w_dff_B_Yh5tGfSY6_2),.clk(gclk));
	jdff dff_B_z2ELHyry4_2(.din(w_dff_B_Yh5tGfSY6_2),.dout(w_dff_B_z2ELHyry4_2),.clk(gclk));
	jdff dff_B_qW6Bg2YV3_2(.din(w_dff_B_z2ELHyry4_2),.dout(w_dff_B_qW6Bg2YV3_2),.clk(gclk));
	jdff dff_B_t36SaB8O2_2(.din(w_dff_B_qW6Bg2YV3_2),.dout(w_dff_B_t36SaB8O2_2),.clk(gclk));
	jdff dff_B_RKhaZqiF6_2(.din(w_dff_B_t36SaB8O2_2),.dout(w_dff_B_RKhaZqiF6_2),.clk(gclk));
	jdff dff_B_knm0k8Xg4_2(.din(w_dff_B_RKhaZqiF6_2),.dout(w_dff_B_knm0k8Xg4_2),.clk(gclk));
	jdff dff_B_yEHtgwAw9_2(.din(w_dff_B_knm0k8Xg4_2),.dout(w_dff_B_yEHtgwAw9_2),.clk(gclk));
	jdff dff_B_CBPGj1Xr9_2(.din(w_dff_B_yEHtgwAw9_2),.dout(w_dff_B_CBPGj1Xr9_2),.clk(gclk));
	jdff dff_B_wfNlrhA39_2(.din(w_dff_B_CBPGj1Xr9_2),.dout(w_dff_B_wfNlrhA39_2),.clk(gclk));
	jdff dff_B_XZWc1MA07_2(.din(w_dff_B_wfNlrhA39_2),.dout(w_dff_B_XZWc1MA07_2),.clk(gclk));
	jdff dff_B_tjYOlqZm1_2(.din(w_dff_B_XZWc1MA07_2),.dout(w_dff_B_tjYOlqZm1_2),.clk(gclk));
	jdff dff_B_hELfrm557_2(.din(w_dff_B_tjYOlqZm1_2),.dout(w_dff_B_hELfrm557_2),.clk(gclk));
	jdff dff_B_EeHt7nf20_2(.din(w_dff_B_hELfrm557_2),.dout(w_dff_B_EeHt7nf20_2),.clk(gclk));
	jdff dff_B_PUVktDH65_2(.din(w_dff_B_EeHt7nf20_2),.dout(w_dff_B_PUVktDH65_2),.clk(gclk));
	jdff dff_B_e8tfmy4u5_2(.din(w_dff_B_PUVktDH65_2),.dout(w_dff_B_e8tfmy4u5_2),.clk(gclk));
	jdff dff_B_DE1T8EcF2_2(.din(w_dff_B_e8tfmy4u5_2),.dout(w_dff_B_DE1T8EcF2_2),.clk(gclk));
	jdff dff_B_DbnIVGSV5_2(.din(w_dff_B_DE1T8EcF2_2),.dout(w_dff_B_DbnIVGSV5_2),.clk(gclk));
	jdff dff_B_Semw6xyf3_2(.din(w_dff_B_DbnIVGSV5_2),.dout(w_dff_B_Semw6xyf3_2),.clk(gclk));
	jdff dff_B_6HL6TPZi0_2(.din(w_dff_B_Semw6xyf3_2),.dout(w_dff_B_6HL6TPZi0_2),.clk(gclk));
	jdff dff_B_dKWFuJb32_2(.din(w_dff_B_6HL6TPZi0_2),.dout(w_dff_B_dKWFuJb32_2),.clk(gclk));
	jdff dff_B_tQwvjZBp2_2(.din(w_dff_B_dKWFuJb32_2),.dout(w_dff_B_tQwvjZBp2_2),.clk(gclk));
	jdff dff_B_O3rmj7Hd0_2(.din(w_dff_B_tQwvjZBp2_2),.dout(w_dff_B_O3rmj7Hd0_2),.clk(gclk));
	jdff dff_B_bSnaak8k2_2(.din(w_dff_B_O3rmj7Hd0_2),.dout(w_dff_B_bSnaak8k2_2),.clk(gclk));
	jdff dff_B_C3SRLnC69_2(.din(w_dff_B_bSnaak8k2_2),.dout(w_dff_B_C3SRLnC69_2),.clk(gclk));
	jdff dff_B_70Xy8b0j3_2(.din(w_dff_B_C3SRLnC69_2),.dout(w_dff_B_70Xy8b0j3_2),.clk(gclk));
	jdff dff_B_zmavL6419_2(.din(w_dff_B_70Xy8b0j3_2),.dout(w_dff_B_zmavL6419_2),.clk(gclk));
	jdff dff_B_0wlAA0ud1_2(.din(w_dff_B_zmavL6419_2),.dout(w_dff_B_0wlAA0ud1_2),.clk(gclk));
	jdff dff_B_ow3Kdl3O0_2(.din(w_dff_B_0wlAA0ud1_2),.dout(w_dff_B_ow3Kdl3O0_2),.clk(gclk));
	jdff dff_B_IXcVz9od3_2(.din(w_dff_B_ow3Kdl3O0_2),.dout(w_dff_B_IXcVz9od3_2),.clk(gclk));
	jdff dff_B_UIupoNSA5_2(.din(w_dff_B_IXcVz9od3_2),.dout(w_dff_B_UIupoNSA5_2),.clk(gclk));
	jdff dff_B_IxFvomfa6_2(.din(w_dff_B_UIupoNSA5_2),.dout(w_dff_B_IxFvomfa6_2),.clk(gclk));
	jdff dff_B_uivDMDmA9_2(.din(w_dff_B_IxFvomfa6_2),.dout(w_dff_B_uivDMDmA9_2),.clk(gclk));
	jdff dff_B_vJbzwzhe9_2(.din(w_dff_B_uivDMDmA9_2),.dout(w_dff_B_vJbzwzhe9_2),.clk(gclk));
	jdff dff_B_y9QMcpst5_2(.din(w_dff_B_vJbzwzhe9_2),.dout(w_dff_B_y9QMcpst5_2),.clk(gclk));
	jdff dff_B_KEC61UbN7_2(.din(w_dff_B_y9QMcpst5_2),.dout(w_dff_B_KEC61UbN7_2),.clk(gclk));
	jdff dff_B_4gjy0nN20_2(.din(w_dff_B_KEC61UbN7_2),.dout(w_dff_B_4gjy0nN20_2),.clk(gclk));
	jdff dff_B_ewia6aDz7_1(.din(n1567),.dout(w_dff_B_ewia6aDz7_1),.clk(gclk));
	jdff dff_B_SPXqW2dm1_2(.din(n1502),.dout(w_dff_B_SPXqW2dm1_2),.clk(gclk));
	jdff dff_B_kTykYwNQ1_2(.din(w_dff_B_SPXqW2dm1_2),.dout(w_dff_B_kTykYwNQ1_2),.clk(gclk));
	jdff dff_B_OC4OnPtO3_2(.din(w_dff_B_kTykYwNQ1_2),.dout(w_dff_B_OC4OnPtO3_2),.clk(gclk));
	jdff dff_B_H1ekknui1_2(.din(w_dff_B_OC4OnPtO3_2),.dout(w_dff_B_H1ekknui1_2),.clk(gclk));
	jdff dff_B_ey9eU7cV7_2(.din(w_dff_B_H1ekknui1_2),.dout(w_dff_B_ey9eU7cV7_2),.clk(gclk));
	jdff dff_B_n7EoCFBQ3_2(.din(w_dff_B_ey9eU7cV7_2),.dout(w_dff_B_n7EoCFBQ3_2),.clk(gclk));
	jdff dff_B_msYtl1oB4_2(.din(w_dff_B_n7EoCFBQ3_2),.dout(w_dff_B_msYtl1oB4_2),.clk(gclk));
	jdff dff_B_DhnOhXgm6_2(.din(w_dff_B_msYtl1oB4_2),.dout(w_dff_B_DhnOhXgm6_2),.clk(gclk));
	jdff dff_B_hPp4pb6m3_2(.din(w_dff_B_DhnOhXgm6_2),.dout(w_dff_B_hPp4pb6m3_2),.clk(gclk));
	jdff dff_B_NcOOZW1C0_2(.din(w_dff_B_hPp4pb6m3_2),.dout(w_dff_B_NcOOZW1C0_2),.clk(gclk));
	jdff dff_B_H9TtCYDc6_2(.din(w_dff_B_NcOOZW1C0_2),.dout(w_dff_B_H9TtCYDc6_2),.clk(gclk));
	jdff dff_B_04DJ5N5p2_2(.din(w_dff_B_H9TtCYDc6_2),.dout(w_dff_B_04DJ5N5p2_2),.clk(gclk));
	jdff dff_B_1VzuVgi55_2(.din(w_dff_B_04DJ5N5p2_2),.dout(w_dff_B_1VzuVgi55_2),.clk(gclk));
	jdff dff_B_jI0d8bc10_2(.din(w_dff_B_1VzuVgi55_2),.dout(w_dff_B_jI0d8bc10_2),.clk(gclk));
	jdff dff_B_W0I0efQf8_2(.din(w_dff_B_jI0d8bc10_2),.dout(w_dff_B_W0I0efQf8_2),.clk(gclk));
	jdff dff_B_w8oH05OQ2_2(.din(w_dff_B_W0I0efQf8_2),.dout(w_dff_B_w8oH05OQ2_2),.clk(gclk));
	jdff dff_B_DCvcBuH23_2(.din(w_dff_B_w8oH05OQ2_2),.dout(w_dff_B_DCvcBuH23_2),.clk(gclk));
	jdff dff_B_PQ9kNBfv0_2(.din(w_dff_B_DCvcBuH23_2),.dout(w_dff_B_PQ9kNBfv0_2),.clk(gclk));
	jdff dff_B_02MewigC3_2(.din(w_dff_B_PQ9kNBfv0_2),.dout(w_dff_B_02MewigC3_2),.clk(gclk));
	jdff dff_B_567YfJb48_2(.din(w_dff_B_02MewigC3_2),.dout(w_dff_B_567YfJb48_2),.clk(gclk));
	jdff dff_B_mv94IPBP5_2(.din(w_dff_B_567YfJb48_2),.dout(w_dff_B_mv94IPBP5_2),.clk(gclk));
	jdff dff_B_Rvyk1bc65_2(.din(w_dff_B_mv94IPBP5_2),.dout(w_dff_B_Rvyk1bc65_2),.clk(gclk));
	jdff dff_B_u2ZuBt3E8_2(.din(w_dff_B_Rvyk1bc65_2),.dout(w_dff_B_u2ZuBt3E8_2),.clk(gclk));
	jdff dff_B_4WU0sOu84_2(.din(w_dff_B_u2ZuBt3E8_2),.dout(w_dff_B_4WU0sOu84_2),.clk(gclk));
	jdff dff_B_nltW59Ju1_2(.din(w_dff_B_4WU0sOu84_2),.dout(w_dff_B_nltW59Ju1_2),.clk(gclk));
	jdff dff_B_1ZNXYIwD0_2(.din(w_dff_B_nltW59Ju1_2),.dout(w_dff_B_1ZNXYIwD0_2),.clk(gclk));
	jdff dff_B_o7z3vP909_2(.din(w_dff_B_1ZNXYIwD0_2),.dout(w_dff_B_o7z3vP909_2),.clk(gclk));
	jdff dff_B_pZPftn4o4_2(.din(w_dff_B_o7z3vP909_2),.dout(w_dff_B_pZPftn4o4_2),.clk(gclk));
	jdff dff_B_nROt5SIt4_2(.din(w_dff_B_pZPftn4o4_2),.dout(w_dff_B_nROt5SIt4_2),.clk(gclk));
	jdff dff_B_ivCzFx8c8_2(.din(w_dff_B_nROt5SIt4_2),.dout(w_dff_B_ivCzFx8c8_2),.clk(gclk));
	jdff dff_B_D8shVlpO4_2(.din(w_dff_B_ivCzFx8c8_2),.dout(w_dff_B_D8shVlpO4_2),.clk(gclk));
	jdff dff_B_HAGUHgsz6_2(.din(w_dff_B_D8shVlpO4_2),.dout(w_dff_B_HAGUHgsz6_2),.clk(gclk));
	jdff dff_B_ASSS5cmR7_2(.din(w_dff_B_HAGUHgsz6_2),.dout(w_dff_B_ASSS5cmR7_2),.clk(gclk));
	jdff dff_B_B8QSHjaK1_2(.din(w_dff_B_ASSS5cmR7_2),.dout(w_dff_B_B8QSHjaK1_2),.clk(gclk));
	jdff dff_B_pBJ2Dndp1_2(.din(w_dff_B_B8QSHjaK1_2),.dout(w_dff_B_pBJ2Dndp1_2),.clk(gclk));
	jdff dff_B_TnpgL7Sz4_2(.din(w_dff_B_pBJ2Dndp1_2),.dout(w_dff_B_TnpgL7Sz4_2),.clk(gclk));
	jdff dff_B_ZFryTQeT9_2(.din(w_dff_B_TnpgL7Sz4_2),.dout(w_dff_B_ZFryTQeT9_2),.clk(gclk));
	jdff dff_B_vpmIoObM3_2(.din(w_dff_B_ZFryTQeT9_2),.dout(w_dff_B_vpmIoObM3_2),.clk(gclk));
	jdff dff_B_7lS39wSh8_2(.din(w_dff_B_vpmIoObM3_2),.dout(w_dff_B_7lS39wSh8_2),.clk(gclk));
	jdff dff_B_t4TYKUIV5_2(.din(w_dff_B_7lS39wSh8_2),.dout(w_dff_B_t4TYKUIV5_2),.clk(gclk));
	jdff dff_B_rG0GDWV04_2(.din(w_dff_B_t4TYKUIV5_2),.dout(w_dff_B_rG0GDWV04_2),.clk(gclk));
	jdff dff_B_2Dc2Cqqv3_2(.din(w_dff_B_rG0GDWV04_2),.dout(w_dff_B_2Dc2Cqqv3_2),.clk(gclk));
	jdff dff_B_DhnMH88a8_2(.din(n1548),.dout(w_dff_B_DhnMH88a8_2),.clk(gclk));
	jdff dff_B_t36JFZHW4_1(.din(n1503),.dout(w_dff_B_t36JFZHW4_1),.clk(gclk));
	jdff dff_B_W2D9LgdN6_2(.din(n1431),.dout(w_dff_B_W2D9LgdN6_2),.clk(gclk));
	jdff dff_B_0WMAt5ZJ9_2(.din(w_dff_B_W2D9LgdN6_2),.dout(w_dff_B_0WMAt5ZJ9_2),.clk(gclk));
	jdff dff_B_27gtSKIT6_2(.din(w_dff_B_0WMAt5ZJ9_2),.dout(w_dff_B_27gtSKIT6_2),.clk(gclk));
	jdff dff_B_2yeudNdz7_2(.din(w_dff_B_27gtSKIT6_2),.dout(w_dff_B_2yeudNdz7_2),.clk(gclk));
	jdff dff_B_mH2dwj8j0_2(.din(w_dff_B_2yeudNdz7_2),.dout(w_dff_B_mH2dwj8j0_2),.clk(gclk));
	jdff dff_B_4ykKdkSo1_2(.din(w_dff_B_mH2dwj8j0_2),.dout(w_dff_B_4ykKdkSo1_2),.clk(gclk));
	jdff dff_B_YQPuyVSy9_2(.din(w_dff_B_4ykKdkSo1_2),.dout(w_dff_B_YQPuyVSy9_2),.clk(gclk));
	jdff dff_B_vRmFT9vW7_2(.din(w_dff_B_YQPuyVSy9_2),.dout(w_dff_B_vRmFT9vW7_2),.clk(gclk));
	jdff dff_B_AQ32ZqUO8_2(.din(w_dff_B_vRmFT9vW7_2),.dout(w_dff_B_AQ32ZqUO8_2),.clk(gclk));
	jdff dff_B_NAzTCZhW0_2(.din(w_dff_B_AQ32ZqUO8_2),.dout(w_dff_B_NAzTCZhW0_2),.clk(gclk));
	jdff dff_B_Xw5Zjdo61_2(.din(w_dff_B_NAzTCZhW0_2),.dout(w_dff_B_Xw5Zjdo61_2),.clk(gclk));
	jdff dff_B_aHC6WF8t9_2(.din(w_dff_B_Xw5Zjdo61_2),.dout(w_dff_B_aHC6WF8t9_2),.clk(gclk));
	jdff dff_B_hsBo7oyx7_2(.din(w_dff_B_aHC6WF8t9_2),.dout(w_dff_B_hsBo7oyx7_2),.clk(gclk));
	jdff dff_B_vl4HxP8H4_2(.din(w_dff_B_hsBo7oyx7_2),.dout(w_dff_B_vl4HxP8H4_2),.clk(gclk));
	jdff dff_B_AZ8Uq0Je9_2(.din(w_dff_B_vl4HxP8H4_2),.dout(w_dff_B_AZ8Uq0Je9_2),.clk(gclk));
	jdff dff_B_c77SKypD8_2(.din(w_dff_B_AZ8Uq0Je9_2),.dout(w_dff_B_c77SKypD8_2),.clk(gclk));
	jdff dff_B_4J9yUMTh4_2(.din(w_dff_B_c77SKypD8_2),.dout(w_dff_B_4J9yUMTh4_2),.clk(gclk));
	jdff dff_B_Kc4qZdze1_2(.din(w_dff_B_4J9yUMTh4_2),.dout(w_dff_B_Kc4qZdze1_2),.clk(gclk));
	jdff dff_B_FUUV2IFK0_2(.din(w_dff_B_Kc4qZdze1_2),.dout(w_dff_B_FUUV2IFK0_2),.clk(gclk));
	jdff dff_B_4IaHg2y39_2(.din(w_dff_B_FUUV2IFK0_2),.dout(w_dff_B_4IaHg2y39_2),.clk(gclk));
	jdff dff_B_tSxKbDZx9_2(.din(w_dff_B_4IaHg2y39_2),.dout(w_dff_B_tSxKbDZx9_2),.clk(gclk));
	jdff dff_B_XsHjt4T17_2(.din(w_dff_B_tSxKbDZx9_2),.dout(w_dff_B_XsHjt4T17_2),.clk(gclk));
	jdff dff_B_zgWTXqDe3_2(.din(w_dff_B_XsHjt4T17_2),.dout(w_dff_B_zgWTXqDe3_2),.clk(gclk));
	jdff dff_B_aQLIWByr2_2(.din(w_dff_B_zgWTXqDe3_2),.dout(w_dff_B_aQLIWByr2_2),.clk(gclk));
	jdff dff_B_vjhBhKZL7_2(.din(w_dff_B_aQLIWByr2_2),.dout(w_dff_B_vjhBhKZL7_2),.clk(gclk));
	jdff dff_B_15SdAugp4_2(.din(w_dff_B_vjhBhKZL7_2),.dout(w_dff_B_15SdAugp4_2),.clk(gclk));
	jdff dff_B_eZaSc35B2_2(.din(w_dff_B_15SdAugp4_2),.dout(w_dff_B_eZaSc35B2_2),.clk(gclk));
	jdff dff_B_s0s7SrLJ2_2(.din(w_dff_B_eZaSc35B2_2),.dout(w_dff_B_s0s7SrLJ2_2),.clk(gclk));
	jdff dff_B_Pf8NYs0X7_2(.din(w_dff_B_s0s7SrLJ2_2),.dout(w_dff_B_Pf8NYs0X7_2),.clk(gclk));
	jdff dff_B_JS6VDofc4_2(.din(w_dff_B_Pf8NYs0X7_2),.dout(w_dff_B_JS6VDofc4_2),.clk(gclk));
	jdff dff_B_MxlpbtEz8_2(.din(w_dff_B_JS6VDofc4_2),.dout(w_dff_B_MxlpbtEz8_2),.clk(gclk));
	jdff dff_B_ryAZhdJc6_2(.din(w_dff_B_MxlpbtEz8_2),.dout(w_dff_B_ryAZhdJc6_2),.clk(gclk));
	jdff dff_B_T8fmoYTS6_2(.din(w_dff_B_ryAZhdJc6_2),.dout(w_dff_B_T8fmoYTS6_2),.clk(gclk));
	jdff dff_B_XVlVHmCQ4_2(.din(w_dff_B_T8fmoYTS6_2),.dout(w_dff_B_XVlVHmCQ4_2),.clk(gclk));
	jdff dff_B_RNOVQFcl9_2(.din(w_dff_B_XVlVHmCQ4_2),.dout(w_dff_B_RNOVQFcl9_2),.clk(gclk));
	jdff dff_B_dgOO3eT99_2(.din(w_dff_B_RNOVQFcl9_2),.dout(w_dff_B_dgOO3eT99_2),.clk(gclk));
	jdff dff_B_cHGSWxIC0_2(.din(w_dff_B_dgOO3eT99_2),.dout(w_dff_B_cHGSWxIC0_2),.clk(gclk));
	jdff dff_B_p9L3JcAh3_2(.din(w_dff_B_cHGSWxIC0_2),.dout(w_dff_B_p9L3JcAh3_2),.clk(gclk));
	jdff dff_B_Gzmv50DE8_2(.din(w_dff_B_p9L3JcAh3_2),.dout(w_dff_B_Gzmv50DE8_2),.clk(gclk));
	jdff dff_B_A3R2VAa63_2(.din(n1477),.dout(w_dff_B_A3R2VAa63_2),.clk(gclk));
	jdff dff_B_NTWXxtiL6_1(.din(n1432),.dout(w_dff_B_NTWXxtiL6_1),.clk(gclk));
	jdff dff_B_RNJJNCz87_2(.din(n1353),.dout(w_dff_B_RNJJNCz87_2),.clk(gclk));
	jdff dff_B_Ao0pvMLT7_2(.din(w_dff_B_RNJJNCz87_2),.dout(w_dff_B_Ao0pvMLT7_2),.clk(gclk));
	jdff dff_B_m5IhTBR80_2(.din(w_dff_B_Ao0pvMLT7_2),.dout(w_dff_B_m5IhTBR80_2),.clk(gclk));
	jdff dff_B_Fv0nOfa90_2(.din(w_dff_B_m5IhTBR80_2),.dout(w_dff_B_Fv0nOfa90_2),.clk(gclk));
	jdff dff_B_rkybG2kM7_2(.din(w_dff_B_Fv0nOfa90_2),.dout(w_dff_B_rkybG2kM7_2),.clk(gclk));
	jdff dff_B_l6mnBk3Z3_2(.din(w_dff_B_rkybG2kM7_2),.dout(w_dff_B_l6mnBk3Z3_2),.clk(gclk));
	jdff dff_B_WTfkTDFu1_2(.din(w_dff_B_l6mnBk3Z3_2),.dout(w_dff_B_WTfkTDFu1_2),.clk(gclk));
	jdff dff_B_8PNFX68G2_2(.din(w_dff_B_WTfkTDFu1_2),.dout(w_dff_B_8PNFX68G2_2),.clk(gclk));
	jdff dff_B_237ECkMK0_2(.din(w_dff_B_8PNFX68G2_2),.dout(w_dff_B_237ECkMK0_2),.clk(gclk));
	jdff dff_B_iMGYnLzT3_2(.din(w_dff_B_237ECkMK0_2),.dout(w_dff_B_iMGYnLzT3_2),.clk(gclk));
	jdff dff_B_WUTQDFVG2_2(.din(w_dff_B_iMGYnLzT3_2),.dout(w_dff_B_WUTQDFVG2_2),.clk(gclk));
	jdff dff_B_ZjXT7OBx5_2(.din(w_dff_B_WUTQDFVG2_2),.dout(w_dff_B_ZjXT7OBx5_2),.clk(gclk));
	jdff dff_B_kAhla4n08_2(.din(w_dff_B_ZjXT7OBx5_2),.dout(w_dff_B_kAhla4n08_2),.clk(gclk));
	jdff dff_B_tomTPd9y1_2(.din(w_dff_B_kAhla4n08_2),.dout(w_dff_B_tomTPd9y1_2),.clk(gclk));
	jdff dff_B_CfCdbbvS2_2(.din(w_dff_B_tomTPd9y1_2),.dout(w_dff_B_CfCdbbvS2_2),.clk(gclk));
	jdff dff_B_3OUYU2I74_2(.din(w_dff_B_CfCdbbvS2_2),.dout(w_dff_B_3OUYU2I74_2),.clk(gclk));
	jdff dff_B_pbxAkWNd0_2(.din(w_dff_B_3OUYU2I74_2),.dout(w_dff_B_pbxAkWNd0_2),.clk(gclk));
	jdff dff_B_R5nBeBZ59_2(.din(w_dff_B_pbxAkWNd0_2),.dout(w_dff_B_R5nBeBZ59_2),.clk(gclk));
	jdff dff_B_QNOqrJ0A8_2(.din(w_dff_B_R5nBeBZ59_2),.dout(w_dff_B_QNOqrJ0A8_2),.clk(gclk));
	jdff dff_B_MoKvDhTo5_2(.din(w_dff_B_QNOqrJ0A8_2),.dout(w_dff_B_MoKvDhTo5_2),.clk(gclk));
	jdff dff_B_J7i9nfDu3_2(.din(w_dff_B_MoKvDhTo5_2),.dout(w_dff_B_J7i9nfDu3_2),.clk(gclk));
	jdff dff_B_TobCk7kL6_2(.din(w_dff_B_J7i9nfDu3_2),.dout(w_dff_B_TobCk7kL6_2),.clk(gclk));
	jdff dff_B_xcs9joq36_2(.din(w_dff_B_TobCk7kL6_2),.dout(w_dff_B_xcs9joq36_2),.clk(gclk));
	jdff dff_B_ZVqcZxM41_2(.din(w_dff_B_xcs9joq36_2),.dout(w_dff_B_ZVqcZxM41_2),.clk(gclk));
	jdff dff_B_P4niPtod4_2(.din(w_dff_B_ZVqcZxM41_2),.dout(w_dff_B_P4niPtod4_2),.clk(gclk));
	jdff dff_B_v92yHpEa5_2(.din(w_dff_B_P4niPtod4_2),.dout(w_dff_B_v92yHpEa5_2),.clk(gclk));
	jdff dff_B_kfOIsyGW9_2(.din(w_dff_B_v92yHpEa5_2),.dout(w_dff_B_kfOIsyGW9_2),.clk(gclk));
	jdff dff_B_1LofYttv4_2(.din(w_dff_B_kfOIsyGW9_2),.dout(w_dff_B_1LofYttv4_2),.clk(gclk));
	jdff dff_B_qrJBSzC89_2(.din(w_dff_B_1LofYttv4_2),.dout(w_dff_B_qrJBSzC89_2),.clk(gclk));
	jdff dff_B_PB6FJwQ53_2(.din(w_dff_B_qrJBSzC89_2),.dout(w_dff_B_PB6FJwQ53_2),.clk(gclk));
	jdff dff_B_MwzE1mE58_2(.din(w_dff_B_PB6FJwQ53_2),.dout(w_dff_B_MwzE1mE58_2),.clk(gclk));
	jdff dff_B_7BAifTpZ3_2(.din(w_dff_B_MwzE1mE58_2),.dout(w_dff_B_7BAifTpZ3_2),.clk(gclk));
	jdff dff_B_eRUPqLDn5_2(.din(w_dff_B_7BAifTpZ3_2),.dout(w_dff_B_eRUPqLDn5_2),.clk(gclk));
	jdff dff_B_gEpaOo1z1_2(.din(w_dff_B_eRUPqLDn5_2),.dout(w_dff_B_gEpaOo1z1_2),.clk(gclk));
	jdff dff_B_vJylCD1i2_2(.din(w_dff_B_gEpaOo1z1_2),.dout(w_dff_B_vJylCD1i2_2),.clk(gclk));
	jdff dff_B_aVwQOu5d0_2(.din(w_dff_B_vJylCD1i2_2),.dout(w_dff_B_aVwQOu5d0_2),.clk(gclk));
	jdff dff_B_1ibA4IKY8_2(.din(n1399),.dout(w_dff_B_1ibA4IKY8_2),.clk(gclk));
	jdff dff_B_sP4Ejq843_1(.din(n1354),.dout(w_dff_B_sP4Ejq843_1),.clk(gclk));
	jdff dff_B_UPfBcQpT9_2(.din(n1268),.dout(w_dff_B_UPfBcQpT9_2),.clk(gclk));
	jdff dff_B_Z5Iv1g5Q9_2(.din(w_dff_B_UPfBcQpT9_2),.dout(w_dff_B_Z5Iv1g5Q9_2),.clk(gclk));
	jdff dff_B_jdLlyNxj6_2(.din(w_dff_B_Z5Iv1g5Q9_2),.dout(w_dff_B_jdLlyNxj6_2),.clk(gclk));
	jdff dff_B_G4MVYnug1_2(.din(w_dff_B_jdLlyNxj6_2),.dout(w_dff_B_G4MVYnug1_2),.clk(gclk));
	jdff dff_B_J4zpvQO48_2(.din(w_dff_B_G4MVYnug1_2),.dout(w_dff_B_J4zpvQO48_2),.clk(gclk));
	jdff dff_B_iXrriSKA5_2(.din(w_dff_B_J4zpvQO48_2),.dout(w_dff_B_iXrriSKA5_2),.clk(gclk));
	jdff dff_B_IML1f4pw4_2(.din(w_dff_B_iXrriSKA5_2),.dout(w_dff_B_IML1f4pw4_2),.clk(gclk));
	jdff dff_B_RCo6VYIV9_2(.din(w_dff_B_IML1f4pw4_2),.dout(w_dff_B_RCo6VYIV9_2),.clk(gclk));
	jdff dff_B_Y0hH1vEO4_2(.din(w_dff_B_RCo6VYIV9_2),.dout(w_dff_B_Y0hH1vEO4_2),.clk(gclk));
	jdff dff_B_nzvBuzoc2_2(.din(w_dff_B_Y0hH1vEO4_2),.dout(w_dff_B_nzvBuzoc2_2),.clk(gclk));
	jdff dff_B_YeruEgU76_2(.din(w_dff_B_nzvBuzoc2_2),.dout(w_dff_B_YeruEgU76_2),.clk(gclk));
	jdff dff_B_LeEsOAyE2_2(.din(w_dff_B_YeruEgU76_2),.dout(w_dff_B_LeEsOAyE2_2),.clk(gclk));
	jdff dff_B_64IjW4vJ1_2(.din(w_dff_B_LeEsOAyE2_2),.dout(w_dff_B_64IjW4vJ1_2),.clk(gclk));
	jdff dff_B_sAwzFx3z9_2(.din(w_dff_B_64IjW4vJ1_2),.dout(w_dff_B_sAwzFx3z9_2),.clk(gclk));
	jdff dff_B_eP4KJ1Ce8_2(.din(w_dff_B_sAwzFx3z9_2),.dout(w_dff_B_eP4KJ1Ce8_2),.clk(gclk));
	jdff dff_B_cycacQty7_2(.din(w_dff_B_eP4KJ1Ce8_2),.dout(w_dff_B_cycacQty7_2),.clk(gclk));
	jdff dff_B_C3SbwQnh2_2(.din(w_dff_B_cycacQty7_2),.dout(w_dff_B_C3SbwQnh2_2),.clk(gclk));
	jdff dff_B_Eyqr2xo32_2(.din(w_dff_B_C3SbwQnh2_2),.dout(w_dff_B_Eyqr2xo32_2),.clk(gclk));
	jdff dff_B_HLctiEbA8_2(.din(w_dff_B_Eyqr2xo32_2),.dout(w_dff_B_HLctiEbA8_2),.clk(gclk));
	jdff dff_B_EEFVhxNg0_2(.din(w_dff_B_HLctiEbA8_2),.dout(w_dff_B_EEFVhxNg0_2),.clk(gclk));
	jdff dff_B_LOoSonQp4_2(.din(w_dff_B_EEFVhxNg0_2),.dout(w_dff_B_LOoSonQp4_2),.clk(gclk));
	jdff dff_B_djsuKSzd7_2(.din(w_dff_B_LOoSonQp4_2),.dout(w_dff_B_djsuKSzd7_2),.clk(gclk));
	jdff dff_B_ZOROOSvj7_2(.din(w_dff_B_djsuKSzd7_2),.dout(w_dff_B_ZOROOSvj7_2),.clk(gclk));
	jdff dff_B_95KqB4Id8_2(.din(w_dff_B_ZOROOSvj7_2),.dout(w_dff_B_95KqB4Id8_2),.clk(gclk));
	jdff dff_B_KVdZoxK02_2(.din(w_dff_B_95KqB4Id8_2),.dout(w_dff_B_KVdZoxK02_2),.clk(gclk));
	jdff dff_B_LcUsYLLa3_2(.din(w_dff_B_KVdZoxK02_2),.dout(w_dff_B_LcUsYLLa3_2),.clk(gclk));
	jdff dff_B_dFmMhxME2_2(.din(w_dff_B_LcUsYLLa3_2),.dout(w_dff_B_dFmMhxME2_2),.clk(gclk));
	jdff dff_B_G4v4cB765_2(.din(w_dff_B_dFmMhxME2_2),.dout(w_dff_B_G4v4cB765_2),.clk(gclk));
	jdff dff_B_txscnVFt6_2(.din(w_dff_B_G4v4cB765_2),.dout(w_dff_B_txscnVFt6_2),.clk(gclk));
	jdff dff_B_b0KI3EAq2_2(.din(w_dff_B_txscnVFt6_2),.dout(w_dff_B_b0KI3EAq2_2),.clk(gclk));
	jdff dff_B_5ndnb7647_2(.din(w_dff_B_b0KI3EAq2_2),.dout(w_dff_B_5ndnb7647_2),.clk(gclk));
	jdff dff_B_xTxfJX3d8_2(.din(w_dff_B_5ndnb7647_2),.dout(w_dff_B_xTxfJX3d8_2),.clk(gclk));
	jdff dff_B_7R0lN1O60_2(.din(w_dff_B_xTxfJX3d8_2),.dout(w_dff_B_7R0lN1O60_2),.clk(gclk));
	jdff dff_B_gBIJsM8w9_2(.din(n1314),.dout(w_dff_B_gBIJsM8w9_2),.clk(gclk));
	jdff dff_B_OV7ggkl04_1(.din(n1269),.dout(w_dff_B_OV7ggkl04_1),.clk(gclk));
	jdff dff_B_q7OUFDbZ9_2(.din(n1178),.dout(w_dff_B_q7OUFDbZ9_2),.clk(gclk));
	jdff dff_B_EdsKtupo0_2(.din(w_dff_B_q7OUFDbZ9_2),.dout(w_dff_B_EdsKtupo0_2),.clk(gclk));
	jdff dff_B_bbHw0lxs0_2(.din(w_dff_B_EdsKtupo0_2),.dout(w_dff_B_bbHw0lxs0_2),.clk(gclk));
	jdff dff_B_Nj5M3Epq0_2(.din(w_dff_B_bbHw0lxs0_2),.dout(w_dff_B_Nj5M3Epq0_2),.clk(gclk));
	jdff dff_B_oaFW9q362_2(.din(w_dff_B_Nj5M3Epq0_2),.dout(w_dff_B_oaFW9q362_2),.clk(gclk));
	jdff dff_B_Gp1rMAbZ4_2(.din(w_dff_B_oaFW9q362_2),.dout(w_dff_B_Gp1rMAbZ4_2),.clk(gclk));
	jdff dff_B_tOq3sVn01_2(.din(w_dff_B_Gp1rMAbZ4_2),.dout(w_dff_B_tOq3sVn01_2),.clk(gclk));
	jdff dff_B_o67CCh235_2(.din(w_dff_B_tOq3sVn01_2),.dout(w_dff_B_o67CCh235_2),.clk(gclk));
	jdff dff_B_MzV4yTXU7_2(.din(w_dff_B_o67CCh235_2),.dout(w_dff_B_MzV4yTXU7_2),.clk(gclk));
	jdff dff_B_74rA2ppH0_2(.din(w_dff_B_MzV4yTXU7_2),.dout(w_dff_B_74rA2ppH0_2),.clk(gclk));
	jdff dff_B_Aovb1Zli7_2(.din(w_dff_B_74rA2ppH0_2),.dout(w_dff_B_Aovb1Zli7_2),.clk(gclk));
	jdff dff_B_T6WNXiWJ1_2(.din(w_dff_B_Aovb1Zli7_2),.dout(w_dff_B_T6WNXiWJ1_2),.clk(gclk));
	jdff dff_B_RscgG0iQ7_2(.din(w_dff_B_T6WNXiWJ1_2),.dout(w_dff_B_RscgG0iQ7_2),.clk(gclk));
	jdff dff_B_JnOtgfc76_2(.din(w_dff_B_RscgG0iQ7_2),.dout(w_dff_B_JnOtgfc76_2),.clk(gclk));
	jdff dff_B_IxwqDl0d7_2(.din(w_dff_B_JnOtgfc76_2),.dout(w_dff_B_IxwqDl0d7_2),.clk(gclk));
	jdff dff_B_8hqdvpSS9_2(.din(w_dff_B_IxwqDl0d7_2),.dout(w_dff_B_8hqdvpSS9_2),.clk(gclk));
	jdff dff_B_PeXW10J35_2(.din(w_dff_B_8hqdvpSS9_2),.dout(w_dff_B_PeXW10J35_2),.clk(gclk));
	jdff dff_B_9dZ3Len40_2(.din(w_dff_B_PeXW10J35_2),.dout(w_dff_B_9dZ3Len40_2),.clk(gclk));
	jdff dff_B_5xM2FZkd0_2(.din(w_dff_B_9dZ3Len40_2),.dout(w_dff_B_5xM2FZkd0_2),.clk(gclk));
	jdff dff_B_E1Fw6C7v8_2(.din(w_dff_B_5xM2FZkd0_2),.dout(w_dff_B_E1Fw6C7v8_2),.clk(gclk));
	jdff dff_B_7Q8qCMYt1_2(.din(w_dff_B_E1Fw6C7v8_2),.dout(w_dff_B_7Q8qCMYt1_2),.clk(gclk));
	jdff dff_B_p90lf7R15_2(.din(w_dff_B_7Q8qCMYt1_2),.dout(w_dff_B_p90lf7R15_2),.clk(gclk));
	jdff dff_B_zHe1xKuS3_2(.din(w_dff_B_p90lf7R15_2),.dout(w_dff_B_zHe1xKuS3_2),.clk(gclk));
	jdff dff_B_8ojM9xyx8_2(.din(w_dff_B_zHe1xKuS3_2),.dout(w_dff_B_8ojM9xyx8_2),.clk(gclk));
	jdff dff_B_rjS4bj6V0_2(.din(w_dff_B_8ojM9xyx8_2),.dout(w_dff_B_rjS4bj6V0_2),.clk(gclk));
	jdff dff_B_aruJWUHh6_2(.din(w_dff_B_rjS4bj6V0_2),.dout(w_dff_B_aruJWUHh6_2),.clk(gclk));
	jdff dff_B_Y0cRz4VG2_2(.din(w_dff_B_aruJWUHh6_2),.dout(w_dff_B_Y0cRz4VG2_2),.clk(gclk));
	jdff dff_B_MhuYKNBv9_2(.din(w_dff_B_Y0cRz4VG2_2),.dout(w_dff_B_MhuYKNBv9_2),.clk(gclk));
	jdff dff_B_EhXr46m92_2(.din(w_dff_B_MhuYKNBv9_2),.dout(w_dff_B_EhXr46m92_2),.clk(gclk));
	jdff dff_B_WTHNYiGv2_2(.din(w_dff_B_EhXr46m92_2),.dout(w_dff_B_WTHNYiGv2_2),.clk(gclk));
	jdff dff_B_lnYCOwVq2_2(.din(n1223),.dout(w_dff_B_lnYCOwVq2_2),.clk(gclk));
	jdff dff_B_uzd3W8qA3_1(.din(n1179),.dout(w_dff_B_uzd3W8qA3_1),.clk(gclk));
	jdff dff_B_xjj871zb0_2(.din(n1074),.dout(w_dff_B_xjj871zb0_2),.clk(gclk));
	jdff dff_B_BZQu8nka9_2(.din(w_dff_B_xjj871zb0_2),.dout(w_dff_B_BZQu8nka9_2),.clk(gclk));
	jdff dff_B_c8yZwTfn0_2(.din(w_dff_B_BZQu8nka9_2),.dout(w_dff_B_c8yZwTfn0_2),.clk(gclk));
	jdff dff_B_yv4d6TTA5_2(.din(w_dff_B_c8yZwTfn0_2),.dout(w_dff_B_yv4d6TTA5_2),.clk(gclk));
	jdff dff_B_WDPk0vP99_2(.din(w_dff_B_yv4d6TTA5_2),.dout(w_dff_B_WDPk0vP99_2),.clk(gclk));
	jdff dff_B_BtEugkbS4_2(.din(w_dff_B_WDPk0vP99_2),.dout(w_dff_B_BtEugkbS4_2),.clk(gclk));
	jdff dff_B_8CIlX0JD2_2(.din(w_dff_B_BtEugkbS4_2),.dout(w_dff_B_8CIlX0JD2_2),.clk(gclk));
	jdff dff_B_vDtilpDP2_2(.din(w_dff_B_8CIlX0JD2_2),.dout(w_dff_B_vDtilpDP2_2),.clk(gclk));
	jdff dff_B_b2SqLpvp0_2(.din(w_dff_B_vDtilpDP2_2),.dout(w_dff_B_b2SqLpvp0_2),.clk(gclk));
	jdff dff_B_icSYXwrt0_2(.din(w_dff_B_b2SqLpvp0_2),.dout(w_dff_B_icSYXwrt0_2),.clk(gclk));
	jdff dff_B_GTN6xiao0_2(.din(w_dff_B_icSYXwrt0_2),.dout(w_dff_B_GTN6xiao0_2),.clk(gclk));
	jdff dff_B_IkiyTq7T5_2(.din(w_dff_B_GTN6xiao0_2),.dout(w_dff_B_IkiyTq7T5_2),.clk(gclk));
	jdff dff_B_sBy8yfAK0_2(.din(w_dff_B_IkiyTq7T5_2),.dout(w_dff_B_sBy8yfAK0_2),.clk(gclk));
	jdff dff_B_ayjmuoYy3_2(.din(w_dff_B_sBy8yfAK0_2),.dout(w_dff_B_ayjmuoYy3_2),.clk(gclk));
	jdff dff_B_c4HkXHup8_2(.din(w_dff_B_ayjmuoYy3_2),.dout(w_dff_B_c4HkXHup8_2),.clk(gclk));
	jdff dff_B_ewLgdc4O5_2(.din(w_dff_B_c4HkXHup8_2),.dout(w_dff_B_ewLgdc4O5_2),.clk(gclk));
	jdff dff_B_0rz40acQ1_2(.din(w_dff_B_ewLgdc4O5_2),.dout(w_dff_B_0rz40acQ1_2),.clk(gclk));
	jdff dff_B_pDr0YIfu4_2(.din(w_dff_B_0rz40acQ1_2),.dout(w_dff_B_pDr0YIfu4_2),.clk(gclk));
	jdff dff_B_ArYQ0XeZ8_2(.din(w_dff_B_pDr0YIfu4_2),.dout(w_dff_B_ArYQ0XeZ8_2),.clk(gclk));
	jdff dff_B_M7tjpi6J9_2(.din(w_dff_B_ArYQ0XeZ8_2),.dout(w_dff_B_M7tjpi6J9_2),.clk(gclk));
	jdff dff_B_K1ETa2s77_2(.din(w_dff_B_M7tjpi6J9_2),.dout(w_dff_B_K1ETa2s77_2),.clk(gclk));
	jdff dff_B_dUA6h99e5_2(.din(w_dff_B_K1ETa2s77_2),.dout(w_dff_B_dUA6h99e5_2),.clk(gclk));
	jdff dff_B_YoWvCeLF3_2(.din(w_dff_B_dUA6h99e5_2),.dout(w_dff_B_YoWvCeLF3_2),.clk(gclk));
	jdff dff_B_I2RdSUql2_2(.din(w_dff_B_YoWvCeLF3_2),.dout(w_dff_B_I2RdSUql2_2),.clk(gclk));
	jdff dff_B_mGmdX3Wl9_2(.din(w_dff_B_I2RdSUql2_2),.dout(w_dff_B_mGmdX3Wl9_2),.clk(gclk));
	jdff dff_B_Aq25DpYO1_2(.din(w_dff_B_mGmdX3Wl9_2),.dout(w_dff_B_Aq25DpYO1_2),.clk(gclk));
	jdff dff_B_0zxA06rf9_2(.din(w_dff_B_Aq25DpYO1_2),.dout(w_dff_B_0zxA06rf9_2),.clk(gclk));
	jdff dff_B_xeE0Cf714_2(.din(n1125),.dout(w_dff_B_xeE0Cf714_2),.clk(gclk));
	jdff dff_B_Xewy7ynQ2_1(.din(n1075),.dout(w_dff_B_Xewy7ynQ2_1),.clk(gclk));
	jdff dff_B_ILqYK7GA6_2(.din(n976),.dout(w_dff_B_ILqYK7GA6_2),.clk(gclk));
	jdff dff_B_KefUfuQX2_2(.din(w_dff_B_ILqYK7GA6_2),.dout(w_dff_B_KefUfuQX2_2),.clk(gclk));
	jdff dff_B_vbYQ3d9e6_2(.din(w_dff_B_KefUfuQX2_2),.dout(w_dff_B_vbYQ3d9e6_2),.clk(gclk));
	jdff dff_B_FxTI3rpf0_2(.din(w_dff_B_vbYQ3d9e6_2),.dout(w_dff_B_FxTI3rpf0_2),.clk(gclk));
	jdff dff_B_eaz4wfXi4_2(.din(w_dff_B_FxTI3rpf0_2),.dout(w_dff_B_eaz4wfXi4_2),.clk(gclk));
	jdff dff_B_jHkGQAW51_2(.din(w_dff_B_eaz4wfXi4_2),.dout(w_dff_B_jHkGQAW51_2),.clk(gclk));
	jdff dff_B_OsQFIn089_2(.din(w_dff_B_jHkGQAW51_2),.dout(w_dff_B_OsQFIn089_2),.clk(gclk));
	jdff dff_B_yMkFgDtb4_2(.din(w_dff_B_OsQFIn089_2),.dout(w_dff_B_yMkFgDtb4_2),.clk(gclk));
	jdff dff_B_oxnhuztm1_2(.din(w_dff_B_yMkFgDtb4_2),.dout(w_dff_B_oxnhuztm1_2),.clk(gclk));
	jdff dff_B_soxTaaV85_2(.din(w_dff_B_oxnhuztm1_2),.dout(w_dff_B_soxTaaV85_2),.clk(gclk));
	jdff dff_B_PLudMCF56_2(.din(w_dff_B_soxTaaV85_2),.dout(w_dff_B_PLudMCF56_2),.clk(gclk));
	jdff dff_B_G3qFdKgE6_2(.din(w_dff_B_PLudMCF56_2),.dout(w_dff_B_G3qFdKgE6_2),.clk(gclk));
	jdff dff_B_ShZ6kQEh3_2(.din(w_dff_B_G3qFdKgE6_2),.dout(w_dff_B_ShZ6kQEh3_2),.clk(gclk));
	jdff dff_B_ynNPUrKu4_2(.din(w_dff_B_ShZ6kQEh3_2),.dout(w_dff_B_ynNPUrKu4_2),.clk(gclk));
	jdff dff_B_PPTnP7aQ2_2(.din(w_dff_B_ynNPUrKu4_2),.dout(w_dff_B_PPTnP7aQ2_2),.clk(gclk));
	jdff dff_B_HmDCQnBm7_2(.din(w_dff_B_PPTnP7aQ2_2),.dout(w_dff_B_HmDCQnBm7_2),.clk(gclk));
	jdff dff_B_snohWNGp8_2(.din(w_dff_B_HmDCQnBm7_2),.dout(w_dff_B_snohWNGp8_2),.clk(gclk));
	jdff dff_B_9o4564HU1_2(.din(w_dff_B_snohWNGp8_2),.dout(w_dff_B_9o4564HU1_2),.clk(gclk));
	jdff dff_B_fV8OAf4n9_2(.din(w_dff_B_9o4564HU1_2),.dout(w_dff_B_fV8OAf4n9_2),.clk(gclk));
	jdff dff_B_xzvpndms1_2(.din(w_dff_B_fV8OAf4n9_2),.dout(w_dff_B_xzvpndms1_2),.clk(gclk));
	jdff dff_B_cAiJ0cTE5_2(.din(w_dff_B_xzvpndms1_2),.dout(w_dff_B_cAiJ0cTE5_2),.clk(gclk));
	jdff dff_B_LglNHTVx1_2(.din(w_dff_B_cAiJ0cTE5_2),.dout(w_dff_B_LglNHTVx1_2),.clk(gclk));
	jdff dff_B_AguJD1uK1_2(.din(w_dff_B_LglNHTVx1_2),.dout(w_dff_B_AguJD1uK1_2),.clk(gclk));
	jdff dff_B_jwFo8Crr7_2(.din(w_dff_B_AguJD1uK1_2),.dout(w_dff_B_jwFo8Crr7_2),.clk(gclk));
	jdff dff_B_srM51NvW5_2(.din(n1020),.dout(w_dff_B_srM51NvW5_2),.clk(gclk));
	jdff dff_B_KizjIKLD4_1(.din(n977),.dout(w_dff_B_KizjIKLD4_1),.clk(gclk));
	jdff dff_B_kJbx6HmA4_2(.din(n871),.dout(w_dff_B_kJbx6HmA4_2),.clk(gclk));
	jdff dff_B_B2LcDPZV8_2(.din(w_dff_B_kJbx6HmA4_2),.dout(w_dff_B_B2LcDPZV8_2),.clk(gclk));
	jdff dff_B_VVtjfoL76_2(.din(w_dff_B_B2LcDPZV8_2),.dout(w_dff_B_VVtjfoL76_2),.clk(gclk));
	jdff dff_B_D6V39gPe4_2(.din(w_dff_B_VVtjfoL76_2),.dout(w_dff_B_D6V39gPe4_2),.clk(gclk));
	jdff dff_B_I7fehIHE4_2(.din(w_dff_B_D6V39gPe4_2),.dout(w_dff_B_I7fehIHE4_2),.clk(gclk));
	jdff dff_B_Xv1jmA005_2(.din(w_dff_B_I7fehIHE4_2),.dout(w_dff_B_Xv1jmA005_2),.clk(gclk));
	jdff dff_B_AzezYvDp3_2(.din(w_dff_B_Xv1jmA005_2),.dout(w_dff_B_AzezYvDp3_2),.clk(gclk));
	jdff dff_B_Lfu3r4Qc2_2(.din(w_dff_B_AzezYvDp3_2),.dout(w_dff_B_Lfu3r4Qc2_2),.clk(gclk));
	jdff dff_B_Vxrn0VrF8_2(.din(w_dff_B_Lfu3r4Qc2_2),.dout(w_dff_B_Vxrn0VrF8_2),.clk(gclk));
	jdff dff_B_joRcfVxS5_2(.din(w_dff_B_Vxrn0VrF8_2),.dout(w_dff_B_joRcfVxS5_2),.clk(gclk));
	jdff dff_B_GIy6Ni797_2(.din(w_dff_B_joRcfVxS5_2),.dout(w_dff_B_GIy6Ni797_2),.clk(gclk));
	jdff dff_B_tEBNFMUf8_2(.din(w_dff_B_GIy6Ni797_2),.dout(w_dff_B_tEBNFMUf8_2),.clk(gclk));
	jdff dff_B_aQAknhHc8_2(.din(w_dff_B_tEBNFMUf8_2),.dout(w_dff_B_aQAknhHc8_2),.clk(gclk));
	jdff dff_B_C3FlaVdQ2_2(.din(w_dff_B_aQAknhHc8_2),.dout(w_dff_B_C3FlaVdQ2_2),.clk(gclk));
	jdff dff_B_4rN7hxPq4_2(.din(w_dff_B_C3FlaVdQ2_2),.dout(w_dff_B_4rN7hxPq4_2),.clk(gclk));
	jdff dff_B_oStUWTwr1_2(.din(w_dff_B_4rN7hxPq4_2),.dout(w_dff_B_oStUWTwr1_2),.clk(gclk));
	jdff dff_B_1FcR4dni7_2(.din(w_dff_B_oStUWTwr1_2),.dout(w_dff_B_1FcR4dni7_2),.clk(gclk));
	jdff dff_B_whimdm246_2(.din(w_dff_B_1FcR4dni7_2),.dout(w_dff_B_whimdm246_2),.clk(gclk));
	jdff dff_B_kwEysLM92_2(.din(w_dff_B_whimdm246_2),.dout(w_dff_B_kwEysLM92_2),.clk(gclk));
	jdff dff_B_5f3kWY4S0_2(.din(w_dff_B_kwEysLM92_2),.dout(w_dff_B_5f3kWY4S0_2),.clk(gclk));
	jdff dff_B_kYkqdPMr6_2(.din(w_dff_B_5f3kWY4S0_2),.dout(w_dff_B_kYkqdPMr6_2),.clk(gclk));
	jdff dff_B_JcBbMAdb9_2(.din(n915),.dout(w_dff_B_JcBbMAdb9_2),.clk(gclk));
	jdff dff_B_c8K0u9p28_1(.din(n872),.dout(w_dff_B_c8K0u9p28_1),.clk(gclk));
	jdff dff_B_HqPS48kr8_2(.din(n772),.dout(w_dff_B_HqPS48kr8_2),.clk(gclk));
	jdff dff_B_JBOVN3QN0_2(.din(w_dff_B_HqPS48kr8_2),.dout(w_dff_B_JBOVN3QN0_2),.clk(gclk));
	jdff dff_B_7TY5rIS07_2(.din(w_dff_B_JBOVN3QN0_2),.dout(w_dff_B_7TY5rIS07_2),.clk(gclk));
	jdff dff_B_nP7lwz5r2_2(.din(w_dff_B_7TY5rIS07_2),.dout(w_dff_B_nP7lwz5r2_2),.clk(gclk));
	jdff dff_B_e4hR2Ggt0_2(.din(w_dff_B_nP7lwz5r2_2),.dout(w_dff_B_e4hR2Ggt0_2),.clk(gclk));
	jdff dff_B_wfs4P79U9_2(.din(w_dff_B_e4hR2Ggt0_2),.dout(w_dff_B_wfs4P79U9_2),.clk(gclk));
	jdff dff_B_AnLpgX643_2(.din(w_dff_B_wfs4P79U9_2),.dout(w_dff_B_AnLpgX643_2),.clk(gclk));
	jdff dff_B_EPu3zuoE4_2(.din(w_dff_B_AnLpgX643_2),.dout(w_dff_B_EPu3zuoE4_2),.clk(gclk));
	jdff dff_B_jk0muqlY7_2(.din(w_dff_B_EPu3zuoE4_2),.dout(w_dff_B_jk0muqlY7_2),.clk(gclk));
	jdff dff_B_Dbv7Pg6n5_2(.din(w_dff_B_jk0muqlY7_2),.dout(w_dff_B_Dbv7Pg6n5_2),.clk(gclk));
	jdff dff_B_EM1pjMts4_2(.din(w_dff_B_Dbv7Pg6n5_2),.dout(w_dff_B_EM1pjMts4_2),.clk(gclk));
	jdff dff_B_32uSxC0p3_2(.din(w_dff_B_EM1pjMts4_2),.dout(w_dff_B_32uSxC0p3_2),.clk(gclk));
	jdff dff_B_CRrFrIAr8_2(.din(w_dff_B_32uSxC0p3_2),.dout(w_dff_B_CRrFrIAr8_2),.clk(gclk));
	jdff dff_B_T16sNmeR3_2(.din(w_dff_B_CRrFrIAr8_2),.dout(w_dff_B_T16sNmeR3_2),.clk(gclk));
	jdff dff_B_j2u7iEnl2_2(.din(w_dff_B_T16sNmeR3_2),.dout(w_dff_B_j2u7iEnl2_2),.clk(gclk));
	jdff dff_B_qVFpwbDJ5_2(.din(w_dff_B_j2u7iEnl2_2),.dout(w_dff_B_qVFpwbDJ5_2),.clk(gclk));
	jdff dff_B_vIE5lVX17_2(.din(w_dff_B_qVFpwbDJ5_2),.dout(w_dff_B_vIE5lVX17_2),.clk(gclk));
	jdff dff_B_BcXpF4rI7_2(.din(w_dff_B_vIE5lVX17_2),.dout(w_dff_B_BcXpF4rI7_2),.clk(gclk));
	jdff dff_B_FgF8KqwX0_2(.din(n809),.dout(w_dff_B_FgF8KqwX0_2),.clk(gclk));
	jdff dff_B_gkIHDYrP0_1(.din(n773),.dout(w_dff_B_gkIHDYrP0_1),.clk(gclk));
	jdff dff_B_KPE4BNW90_2(.din(n679),.dout(w_dff_B_KPE4BNW90_2),.clk(gclk));
	jdff dff_B_IxD6OlcQ7_2(.din(w_dff_B_KPE4BNW90_2),.dout(w_dff_B_IxD6OlcQ7_2),.clk(gclk));
	jdff dff_B_Q6TigjFH5_2(.din(w_dff_B_IxD6OlcQ7_2),.dout(w_dff_B_Q6TigjFH5_2),.clk(gclk));
	jdff dff_B_ORohxeBL6_2(.din(w_dff_B_Q6TigjFH5_2),.dout(w_dff_B_ORohxeBL6_2),.clk(gclk));
	jdff dff_B_xfRwrgGu7_2(.din(w_dff_B_ORohxeBL6_2),.dout(w_dff_B_xfRwrgGu7_2),.clk(gclk));
	jdff dff_B_JRz79APs0_2(.din(w_dff_B_xfRwrgGu7_2),.dout(w_dff_B_JRz79APs0_2),.clk(gclk));
	jdff dff_B_vI6OPqDp0_2(.din(w_dff_B_JRz79APs0_2),.dout(w_dff_B_vI6OPqDp0_2),.clk(gclk));
	jdff dff_B_VQPOLqxI8_2(.din(w_dff_B_vI6OPqDp0_2),.dout(w_dff_B_VQPOLqxI8_2),.clk(gclk));
	jdff dff_B_n3VJb7os0_2(.din(w_dff_B_VQPOLqxI8_2),.dout(w_dff_B_n3VJb7os0_2),.clk(gclk));
	jdff dff_B_PXpKiGS69_2(.din(w_dff_B_n3VJb7os0_2),.dout(w_dff_B_PXpKiGS69_2),.clk(gclk));
	jdff dff_B_0NrkS6646_2(.din(w_dff_B_PXpKiGS69_2),.dout(w_dff_B_0NrkS6646_2),.clk(gclk));
	jdff dff_B_JAffA4Ep7_2(.din(w_dff_B_0NrkS6646_2),.dout(w_dff_B_JAffA4Ep7_2),.clk(gclk));
	jdff dff_B_qZizcAE34_2(.din(w_dff_B_JAffA4Ep7_2),.dout(w_dff_B_qZizcAE34_2),.clk(gclk));
	jdff dff_B_Pec7xNWs6_2(.din(w_dff_B_qZizcAE34_2),.dout(w_dff_B_Pec7xNWs6_2),.clk(gclk));
	jdff dff_B_TGg6KFiC7_2(.din(w_dff_B_Pec7xNWs6_2),.dout(w_dff_B_TGg6KFiC7_2),.clk(gclk));
	jdff dff_B_4fGVicy57_2(.din(n709),.dout(w_dff_B_4fGVicy57_2),.clk(gclk));
	jdff dff_B_6qB0P92B1_1(.din(n680),.dout(w_dff_B_6qB0P92B1_1),.clk(gclk));
	jdff dff_B_7blUpne13_2(.din(n593),.dout(w_dff_B_7blUpne13_2),.clk(gclk));
	jdff dff_B_C4QfKUdZ7_2(.din(w_dff_B_7blUpne13_2),.dout(w_dff_B_C4QfKUdZ7_2),.clk(gclk));
	jdff dff_B_ekc50hko6_2(.din(w_dff_B_C4QfKUdZ7_2),.dout(w_dff_B_ekc50hko6_2),.clk(gclk));
	jdff dff_B_LJBvSjCD6_2(.din(w_dff_B_ekc50hko6_2),.dout(w_dff_B_LJBvSjCD6_2),.clk(gclk));
	jdff dff_B_aK4zCiUF0_2(.din(w_dff_B_LJBvSjCD6_2),.dout(w_dff_B_aK4zCiUF0_2),.clk(gclk));
	jdff dff_B_4L345AdN8_2(.din(w_dff_B_aK4zCiUF0_2),.dout(w_dff_B_4L345AdN8_2),.clk(gclk));
	jdff dff_B_ieqWtctJ7_2(.din(w_dff_B_4L345AdN8_2),.dout(w_dff_B_ieqWtctJ7_2),.clk(gclk));
	jdff dff_B_jBAJX7Gd4_2(.din(w_dff_B_ieqWtctJ7_2),.dout(w_dff_B_jBAJX7Gd4_2),.clk(gclk));
	jdff dff_B_27o1vert5_2(.din(w_dff_B_jBAJX7Gd4_2),.dout(w_dff_B_27o1vert5_2),.clk(gclk));
	jdff dff_B_emLOxp1V6_2(.din(w_dff_B_27o1vert5_2),.dout(w_dff_B_emLOxp1V6_2),.clk(gclk));
	jdff dff_B_FXgapH284_2(.din(w_dff_B_emLOxp1V6_2),.dout(w_dff_B_FXgapH284_2),.clk(gclk));
	jdff dff_B_DbqvFnC43_2(.din(w_dff_B_FXgapH284_2),.dout(w_dff_B_DbqvFnC43_2),.clk(gclk));
	jdff dff_B_oy8umolf6_2(.din(n616),.dout(w_dff_B_oy8umolf6_2),.clk(gclk));
	jdff dff_B_rAYAdfFl2_1(.din(n594),.dout(w_dff_B_rAYAdfFl2_1),.clk(gclk));
	jdff dff_B_ja1CMELV8_2(.din(n514),.dout(w_dff_B_ja1CMELV8_2),.clk(gclk));
	jdff dff_B_5qSuCpD44_2(.din(w_dff_B_ja1CMELV8_2),.dout(w_dff_B_5qSuCpD44_2),.clk(gclk));
	jdff dff_B_f8f72HM14_2(.din(w_dff_B_5qSuCpD44_2),.dout(w_dff_B_f8f72HM14_2),.clk(gclk));
	jdff dff_B_L2PET60S9_2(.din(w_dff_B_f8f72HM14_2),.dout(w_dff_B_L2PET60S9_2),.clk(gclk));
	jdff dff_B_4bgFc24M3_2(.din(w_dff_B_L2PET60S9_2),.dout(w_dff_B_4bgFc24M3_2),.clk(gclk));
	jdff dff_B_dSKmSjOY5_2(.din(w_dff_B_4bgFc24M3_2),.dout(w_dff_B_dSKmSjOY5_2),.clk(gclk));
	jdff dff_B_yx21GZjs0_2(.din(w_dff_B_dSKmSjOY5_2),.dout(w_dff_B_yx21GZjs0_2),.clk(gclk));
	jdff dff_B_NnjONBx14_2(.din(w_dff_B_yx21GZjs0_2),.dout(w_dff_B_NnjONBx14_2),.clk(gclk));
	jdff dff_B_aWyavlEF5_2(.din(w_dff_B_NnjONBx14_2),.dout(w_dff_B_aWyavlEF5_2),.clk(gclk));
	jdff dff_B_CmShW5m65_2(.din(n530),.dout(w_dff_B_CmShW5m65_2),.clk(gclk));
	jdff dff_B_QiWXyrP18_2(.din(w_dff_B_CmShW5m65_2),.dout(w_dff_B_QiWXyrP18_2),.clk(gclk));
	jdff dff_B_okGvTIfp4_1(.din(n515),.dout(w_dff_B_okGvTIfp4_1),.clk(gclk));
	jdff dff_B_Ovga210J9_1(.din(w_dff_B_okGvTIfp4_1),.dout(w_dff_B_Ovga210J9_1),.clk(gclk));
	jdff dff_B_cfkcpT9w5_1(.din(w_dff_B_Ovga210J9_1),.dout(w_dff_B_cfkcpT9w5_1),.clk(gclk));
	jdff dff_B_DNOyaLVM2_1(.din(w_dff_B_cfkcpT9w5_1),.dout(w_dff_B_DNOyaLVM2_1),.clk(gclk));
	jdff dff_B_N1MTUlbu6_1(.din(w_dff_B_DNOyaLVM2_1),.dout(w_dff_B_N1MTUlbu6_1),.clk(gclk));
	jdff dff_B_Oo0S0JvP8_1(.din(w_dff_B_N1MTUlbu6_1),.dout(w_dff_B_Oo0S0JvP8_1),.clk(gclk));
	jdff dff_B_2LjfKZ2q1_0(.din(n451),.dout(w_dff_B_2LjfKZ2q1_0),.clk(gclk));
	jdff dff_B_fzZDPGCA0_0(.din(w_dff_B_2LjfKZ2q1_0),.dout(w_dff_B_fzZDPGCA0_0),.clk(gclk));
	jdff dff_A_uHGO6zZS9_0(.dout(w_n450_0[0]),.din(w_dff_A_uHGO6zZS9_0),.clk(gclk));
	jdff dff_A_qXO6zwHi7_0(.dout(w_dff_A_uHGO6zZS9_0),.din(w_dff_A_qXO6zwHi7_0),.clk(gclk));
	jdff dff_A_PzvLBQM62_0(.dout(w_dff_A_qXO6zwHi7_0),.din(w_dff_A_PzvLBQM62_0),.clk(gclk));
	jdff dff_B_kfrBW14e5_1(.din(n444),.dout(w_dff_B_kfrBW14e5_1),.clk(gclk));
	jdff dff_A_OqaIikFK2_0(.dout(w_n376_0[0]),.din(w_dff_A_OqaIikFK2_0),.clk(gclk));
	jdff dff_A_OSxUYutW3_1(.dout(w_n376_0[1]),.din(w_dff_A_OSxUYutW3_1),.clk(gclk));
	jdff dff_A_RVoeUevc7_1(.dout(w_dff_A_OSxUYutW3_1),.din(w_dff_A_RVoeUevc7_1),.clk(gclk));
	jdff dff_A_teBB2hqj4_1(.dout(w_n442_0[1]),.din(w_dff_A_teBB2hqj4_1),.clk(gclk));
	jdff dff_A_tV7cHCuR6_1(.dout(w_dff_A_teBB2hqj4_1),.din(w_dff_A_tV7cHCuR6_1),.clk(gclk));
	jdff dff_A_MwvqcJvR8_1(.dout(w_dff_A_tV7cHCuR6_1),.din(w_dff_A_MwvqcJvR8_1),.clk(gclk));
	jdff dff_A_i0ZkdQHk1_1(.dout(w_dff_A_MwvqcJvR8_1),.din(w_dff_A_i0ZkdQHk1_1),.clk(gclk));
	jdff dff_A_WrFDIzY00_1(.dout(w_dff_A_i0ZkdQHk1_1),.din(w_dff_A_WrFDIzY00_1),.clk(gclk));
	jdff dff_A_mAPv3Wu33_1(.dout(w_dff_A_WrFDIzY00_1),.din(w_dff_A_mAPv3Wu33_1),.clk(gclk));
	jdff dff_B_3RnJicDM9_2(.din(n1682),.dout(w_dff_B_3RnJicDM9_2),.clk(gclk));
	jdff dff_B_VVOCdBKQ9_1(.din(n1680),.dout(w_dff_B_VVOCdBKQ9_1),.clk(gclk));
	jdff dff_B_rQGk3lVe3_2(.din(n1628),.dout(w_dff_B_rQGk3lVe3_2),.clk(gclk));
	jdff dff_B_H1sxGiWm9_2(.din(w_dff_B_rQGk3lVe3_2),.dout(w_dff_B_H1sxGiWm9_2),.clk(gclk));
	jdff dff_B_SJ3sHZQ76_2(.din(w_dff_B_H1sxGiWm9_2),.dout(w_dff_B_SJ3sHZQ76_2),.clk(gclk));
	jdff dff_B_vdXYDhFr4_2(.din(w_dff_B_SJ3sHZQ76_2),.dout(w_dff_B_vdXYDhFr4_2),.clk(gclk));
	jdff dff_B_gwD71AgJ4_2(.din(w_dff_B_vdXYDhFr4_2),.dout(w_dff_B_gwD71AgJ4_2),.clk(gclk));
	jdff dff_B_FLBhM1gE1_2(.din(w_dff_B_gwD71AgJ4_2),.dout(w_dff_B_FLBhM1gE1_2),.clk(gclk));
	jdff dff_B_k97zJxyz8_2(.din(w_dff_B_FLBhM1gE1_2),.dout(w_dff_B_k97zJxyz8_2),.clk(gclk));
	jdff dff_B_TIjQOkkX5_2(.din(w_dff_B_k97zJxyz8_2),.dout(w_dff_B_TIjQOkkX5_2),.clk(gclk));
	jdff dff_B_C9K4kJzr3_2(.din(w_dff_B_TIjQOkkX5_2),.dout(w_dff_B_C9K4kJzr3_2),.clk(gclk));
	jdff dff_B_N4ORJPVi3_2(.din(w_dff_B_C9K4kJzr3_2),.dout(w_dff_B_N4ORJPVi3_2),.clk(gclk));
	jdff dff_B_Z0giA0840_2(.din(w_dff_B_N4ORJPVi3_2),.dout(w_dff_B_Z0giA0840_2),.clk(gclk));
	jdff dff_B_MFFiOSBY4_2(.din(w_dff_B_Z0giA0840_2),.dout(w_dff_B_MFFiOSBY4_2),.clk(gclk));
	jdff dff_B_MANj7Cr24_2(.din(w_dff_B_MFFiOSBY4_2),.dout(w_dff_B_MANj7Cr24_2),.clk(gclk));
	jdff dff_B_K50yHLw83_2(.din(w_dff_B_MANj7Cr24_2),.dout(w_dff_B_K50yHLw83_2),.clk(gclk));
	jdff dff_B_04MGH8kK4_2(.din(w_dff_B_K50yHLw83_2),.dout(w_dff_B_04MGH8kK4_2),.clk(gclk));
	jdff dff_B_yKcc2K6C6_2(.din(w_dff_B_04MGH8kK4_2),.dout(w_dff_B_yKcc2K6C6_2),.clk(gclk));
	jdff dff_B_oUwf0fKg8_2(.din(w_dff_B_yKcc2K6C6_2),.dout(w_dff_B_oUwf0fKg8_2),.clk(gclk));
	jdff dff_B_BboUODOo8_2(.din(w_dff_B_oUwf0fKg8_2),.dout(w_dff_B_BboUODOo8_2),.clk(gclk));
	jdff dff_B_SHciex9f9_2(.din(w_dff_B_BboUODOo8_2),.dout(w_dff_B_SHciex9f9_2),.clk(gclk));
	jdff dff_B_OoS0rA8j2_2(.din(w_dff_B_SHciex9f9_2),.dout(w_dff_B_OoS0rA8j2_2),.clk(gclk));
	jdff dff_B_4lqdVSLO9_2(.din(w_dff_B_OoS0rA8j2_2),.dout(w_dff_B_4lqdVSLO9_2),.clk(gclk));
	jdff dff_B_46iNrCSM2_2(.din(w_dff_B_4lqdVSLO9_2),.dout(w_dff_B_46iNrCSM2_2),.clk(gclk));
	jdff dff_B_SyTGHSIE7_2(.din(w_dff_B_46iNrCSM2_2),.dout(w_dff_B_SyTGHSIE7_2),.clk(gclk));
	jdff dff_B_JsB3ySxS8_2(.din(w_dff_B_SyTGHSIE7_2),.dout(w_dff_B_JsB3ySxS8_2),.clk(gclk));
	jdff dff_B_t0h8V9m91_2(.din(w_dff_B_JsB3ySxS8_2),.dout(w_dff_B_t0h8V9m91_2),.clk(gclk));
	jdff dff_B_jZQQWcrI5_2(.din(w_dff_B_t0h8V9m91_2),.dout(w_dff_B_jZQQWcrI5_2),.clk(gclk));
	jdff dff_B_HGM76Mk49_2(.din(w_dff_B_jZQQWcrI5_2),.dout(w_dff_B_HGM76Mk49_2),.clk(gclk));
	jdff dff_B_DjSDpkoM1_2(.din(w_dff_B_HGM76Mk49_2),.dout(w_dff_B_DjSDpkoM1_2),.clk(gclk));
	jdff dff_B_dc9NxKfl2_2(.din(w_dff_B_DjSDpkoM1_2),.dout(w_dff_B_dc9NxKfl2_2),.clk(gclk));
	jdff dff_B_WnYEq7mm6_2(.din(w_dff_B_dc9NxKfl2_2),.dout(w_dff_B_WnYEq7mm6_2),.clk(gclk));
	jdff dff_B_6E6uATDr7_2(.din(w_dff_B_WnYEq7mm6_2),.dout(w_dff_B_6E6uATDr7_2),.clk(gclk));
	jdff dff_B_nB2Qk6472_2(.din(w_dff_B_6E6uATDr7_2),.dout(w_dff_B_nB2Qk6472_2),.clk(gclk));
	jdff dff_B_eBpkP9O22_2(.din(w_dff_B_nB2Qk6472_2),.dout(w_dff_B_eBpkP9O22_2),.clk(gclk));
	jdff dff_B_RtIma7D91_2(.din(w_dff_B_eBpkP9O22_2),.dout(w_dff_B_RtIma7D91_2),.clk(gclk));
	jdff dff_B_GGChZvOx8_2(.din(w_dff_B_RtIma7D91_2),.dout(w_dff_B_GGChZvOx8_2),.clk(gclk));
	jdff dff_B_yeOGpDpF3_2(.din(w_dff_B_GGChZvOx8_2),.dout(w_dff_B_yeOGpDpF3_2),.clk(gclk));
	jdff dff_B_zGTN5gvK3_2(.din(w_dff_B_yeOGpDpF3_2),.dout(w_dff_B_zGTN5gvK3_2),.clk(gclk));
	jdff dff_B_MxzjAqhn0_2(.din(w_dff_B_zGTN5gvK3_2),.dout(w_dff_B_MxzjAqhn0_2),.clk(gclk));
	jdff dff_B_bigACyS58_2(.din(w_dff_B_MxzjAqhn0_2),.dout(w_dff_B_bigACyS58_2),.clk(gclk));
	jdff dff_B_cOGu1qVi3_2(.din(w_dff_B_bigACyS58_2),.dout(w_dff_B_cOGu1qVi3_2),.clk(gclk));
	jdff dff_B_dLX3NpNs7_2(.din(w_dff_B_cOGu1qVi3_2),.dout(w_dff_B_dLX3NpNs7_2),.clk(gclk));
	jdff dff_B_z1i7qGpa8_2(.din(w_dff_B_dLX3NpNs7_2),.dout(w_dff_B_z1i7qGpa8_2),.clk(gclk));
	jdff dff_B_vFbDe1Cc7_2(.din(w_dff_B_z1i7qGpa8_2),.dout(w_dff_B_vFbDe1Cc7_2),.clk(gclk));
	jdff dff_B_L0r0AVv03_2(.din(w_dff_B_vFbDe1Cc7_2),.dout(w_dff_B_L0r0AVv03_2),.clk(gclk));
	jdff dff_B_iJxvJt2Q7_2(.din(w_dff_B_L0r0AVv03_2),.dout(w_dff_B_iJxvJt2Q7_2),.clk(gclk));
	jdff dff_B_Hxpq3uqt4_2(.din(w_dff_B_iJxvJt2Q7_2),.dout(w_dff_B_Hxpq3uqt4_2),.clk(gclk));
	jdff dff_B_DRCkAmS47_2(.din(w_dff_B_Hxpq3uqt4_2),.dout(w_dff_B_DRCkAmS47_2),.clk(gclk));
	jdff dff_B_oshq8HRc1_2(.din(w_dff_B_DRCkAmS47_2),.dout(w_dff_B_oshq8HRc1_2),.clk(gclk));
	jdff dff_B_8udX8bne1_2(.din(w_dff_B_oshq8HRc1_2),.dout(w_dff_B_8udX8bne1_2),.clk(gclk));
	jdff dff_B_rqcdsL8S1_1(.din(n1678),.dout(w_dff_B_rqcdsL8S1_1),.clk(gclk));
	jdff dff_A_4JJX4vbh2_1(.dout(w_n1631_0[1]),.din(w_dff_A_4JJX4vbh2_1),.clk(gclk));
	jdff dff_B_caV1Uciq4_1(.din(n1629),.dout(w_dff_B_caV1Uciq4_1),.clk(gclk));
	jdff dff_B_00vZXMjC9_2(.din(n1571),.dout(w_dff_B_00vZXMjC9_2),.clk(gclk));
	jdff dff_B_OMYvfEqK5_2(.din(w_dff_B_00vZXMjC9_2),.dout(w_dff_B_OMYvfEqK5_2),.clk(gclk));
	jdff dff_B_DsR74SI38_2(.din(w_dff_B_OMYvfEqK5_2),.dout(w_dff_B_DsR74SI38_2),.clk(gclk));
	jdff dff_B_2Knia5NI5_2(.din(w_dff_B_DsR74SI38_2),.dout(w_dff_B_2Knia5NI5_2),.clk(gclk));
	jdff dff_B_T6O79sgf8_2(.din(w_dff_B_2Knia5NI5_2),.dout(w_dff_B_T6O79sgf8_2),.clk(gclk));
	jdff dff_B_z9TPqOtJ6_2(.din(w_dff_B_T6O79sgf8_2),.dout(w_dff_B_z9TPqOtJ6_2),.clk(gclk));
	jdff dff_B_6Fef7Z8Z2_2(.din(w_dff_B_z9TPqOtJ6_2),.dout(w_dff_B_6Fef7Z8Z2_2),.clk(gclk));
	jdff dff_B_TRGcbW495_2(.din(w_dff_B_6Fef7Z8Z2_2),.dout(w_dff_B_TRGcbW495_2),.clk(gclk));
	jdff dff_B_Ue3RsntW9_2(.din(w_dff_B_TRGcbW495_2),.dout(w_dff_B_Ue3RsntW9_2),.clk(gclk));
	jdff dff_B_474AUWGh0_2(.din(w_dff_B_Ue3RsntW9_2),.dout(w_dff_B_474AUWGh0_2),.clk(gclk));
	jdff dff_B_ajBr2uW02_2(.din(w_dff_B_474AUWGh0_2),.dout(w_dff_B_ajBr2uW02_2),.clk(gclk));
	jdff dff_B_fRCweLPu0_2(.din(w_dff_B_ajBr2uW02_2),.dout(w_dff_B_fRCweLPu0_2),.clk(gclk));
	jdff dff_B_I7lrImhF5_2(.din(w_dff_B_fRCweLPu0_2),.dout(w_dff_B_I7lrImhF5_2),.clk(gclk));
	jdff dff_B_2XBlZWlG4_2(.din(w_dff_B_I7lrImhF5_2),.dout(w_dff_B_2XBlZWlG4_2),.clk(gclk));
	jdff dff_B_tKsrIPLH9_2(.din(w_dff_B_2XBlZWlG4_2),.dout(w_dff_B_tKsrIPLH9_2),.clk(gclk));
	jdff dff_B_ICsQXzqu8_2(.din(w_dff_B_tKsrIPLH9_2),.dout(w_dff_B_ICsQXzqu8_2),.clk(gclk));
	jdff dff_B_6QXffW1I2_2(.din(w_dff_B_ICsQXzqu8_2),.dout(w_dff_B_6QXffW1I2_2),.clk(gclk));
	jdff dff_B_5Av5Qla75_2(.din(w_dff_B_6QXffW1I2_2),.dout(w_dff_B_5Av5Qla75_2),.clk(gclk));
	jdff dff_B_SGU9ONIy9_2(.din(w_dff_B_5Av5Qla75_2),.dout(w_dff_B_SGU9ONIy9_2),.clk(gclk));
	jdff dff_B_AScHc9bz7_2(.din(w_dff_B_SGU9ONIy9_2),.dout(w_dff_B_AScHc9bz7_2),.clk(gclk));
	jdff dff_B_rIh4aMwv5_2(.din(w_dff_B_AScHc9bz7_2),.dout(w_dff_B_rIh4aMwv5_2),.clk(gclk));
	jdff dff_B_78i17mhF0_2(.din(w_dff_B_rIh4aMwv5_2),.dout(w_dff_B_78i17mhF0_2),.clk(gclk));
	jdff dff_B_ptYBTz6k8_2(.din(w_dff_B_78i17mhF0_2),.dout(w_dff_B_ptYBTz6k8_2),.clk(gclk));
	jdff dff_B_lIpR6Luf5_2(.din(w_dff_B_ptYBTz6k8_2),.dout(w_dff_B_lIpR6Luf5_2),.clk(gclk));
	jdff dff_B_sa5nhSK93_2(.din(w_dff_B_lIpR6Luf5_2),.dout(w_dff_B_sa5nhSK93_2),.clk(gclk));
	jdff dff_B_9vYERfv13_2(.din(w_dff_B_sa5nhSK93_2),.dout(w_dff_B_9vYERfv13_2),.clk(gclk));
	jdff dff_B_AmwdL0Gj9_2(.din(w_dff_B_9vYERfv13_2),.dout(w_dff_B_AmwdL0Gj9_2),.clk(gclk));
	jdff dff_B_XJk98zk63_2(.din(w_dff_B_AmwdL0Gj9_2),.dout(w_dff_B_XJk98zk63_2),.clk(gclk));
	jdff dff_B_mc0IQvLR4_2(.din(w_dff_B_XJk98zk63_2),.dout(w_dff_B_mc0IQvLR4_2),.clk(gclk));
	jdff dff_B_t9UkyfRx6_2(.din(w_dff_B_mc0IQvLR4_2),.dout(w_dff_B_t9UkyfRx6_2),.clk(gclk));
	jdff dff_B_rxn0rczN1_2(.din(w_dff_B_t9UkyfRx6_2),.dout(w_dff_B_rxn0rczN1_2),.clk(gclk));
	jdff dff_B_HQz4GrLV4_2(.din(w_dff_B_rxn0rczN1_2),.dout(w_dff_B_HQz4GrLV4_2),.clk(gclk));
	jdff dff_B_P6z2MrgN2_2(.din(w_dff_B_HQz4GrLV4_2),.dout(w_dff_B_P6z2MrgN2_2),.clk(gclk));
	jdff dff_B_Q3l6Dwu72_2(.din(w_dff_B_P6z2MrgN2_2),.dout(w_dff_B_Q3l6Dwu72_2),.clk(gclk));
	jdff dff_B_TQORNAjw3_2(.din(w_dff_B_Q3l6Dwu72_2),.dout(w_dff_B_TQORNAjw3_2),.clk(gclk));
	jdff dff_B_Ni5NJVNp1_2(.din(w_dff_B_TQORNAjw3_2),.dout(w_dff_B_Ni5NJVNp1_2),.clk(gclk));
	jdff dff_B_oLOv9SCj5_2(.din(w_dff_B_Ni5NJVNp1_2),.dout(w_dff_B_oLOv9SCj5_2),.clk(gclk));
	jdff dff_B_ue0jFElA2_2(.din(w_dff_B_oLOv9SCj5_2),.dout(w_dff_B_ue0jFElA2_2),.clk(gclk));
	jdff dff_B_4Jvsh2GY7_2(.din(w_dff_B_ue0jFElA2_2),.dout(w_dff_B_4Jvsh2GY7_2),.clk(gclk));
	jdff dff_B_lo3ZEi1K0_2(.din(w_dff_B_4Jvsh2GY7_2),.dout(w_dff_B_lo3ZEi1K0_2),.clk(gclk));
	jdff dff_B_lc7UO8933_2(.din(w_dff_B_lo3ZEi1K0_2),.dout(w_dff_B_lc7UO8933_2),.clk(gclk));
	jdff dff_B_svI6uF3k7_2(.din(w_dff_B_lc7UO8933_2),.dout(w_dff_B_svI6uF3k7_2),.clk(gclk));
	jdff dff_B_zYjooRPh7_2(.din(w_dff_B_svI6uF3k7_2),.dout(w_dff_B_zYjooRPh7_2),.clk(gclk));
	jdff dff_B_rKUlpOpo5_2(.din(n1574),.dout(w_dff_B_rKUlpOpo5_2),.clk(gclk));
	jdff dff_B_OVFaeoJQ4_1(.din(n1572),.dout(w_dff_B_OVFaeoJQ4_1),.clk(gclk));
	jdff dff_B_dxyA2MqL0_2(.din(n1507),.dout(w_dff_B_dxyA2MqL0_2),.clk(gclk));
	jdff dff_B_F0NMUvbu7_2(.din(w_dff_B_dxyA2MqL0_2),.dout(w_dff_B_F0NMUvbu7_2),.clk(gclk));
	jdff dff_B_jMvfmP3p5_2(.din(w_dff_B_F0NMUvbu7_2),.dout(w_dff_B_jMvfmP3p5_2),.clk(gclk));
	jdff dff_B_q5vBtwrN5_2(.din(w_dff_B_jMvfmP3p5_2),.dout(w_dff_B_q5vBtwrN5_2),.clk(gclk));
	jdff dff_B_AwtR4eou3_2(.din(w_dff_B_q5vBtwrN5_2),.dout(w_dff_B_AwtR4eou3_2),.clk(gclk));
	jdff dff_B_q1W5I5cG8_2(.din(w_dff_B_AwtR4eou3_2),.dout(w_dff_B_q1W5I5cG8_2),.clk(gclk));
	jdff dff_B_8DqNIZRW2_2(.din(w_dff_B_q1W5I5cG8_2),.dout(w_dff_B_8DqNIZRW2_2),.clk(gclk));
	jdff dff_B_dtoVpleY8_2(.din(w_dff_B_8DqNIZRW2_2),.dout(w_dff_B_dtoVpleY8_2),.clk(gclk));
	jdff dff_B_KpsN6g3A3_2(.din(w_dff_B_dtoVpleY8_2),.dout(w_dff_B_KpsN6g3A3_2),.clk(gclk));
	jdff dff_B_UUpkqryu9_2(.din(w_dff_B_KpsN6g3A3_2),.dout(w_dff_B_UUpkqryu9_2),.clk(gclk));
	jdff dff_B_Z0mBabTw8_2(.din(w_dff_B_UUpkqryu9_2),.dout(w_dff_B_Z0mBabTw8_2),.clk(gclk));
	jdff dff_B_70Vadccr9_2(.din(w_dff_B_Z0mBabTw8_2),.dout(w_dff_B_70Vadccr9_2),.clk(gclk));
	jdff dff_B_BkAydNWi0_2(.din(w_dff_B_70Vadccr9_2),.dout(w_dff_B_BkAydNWi0_2),.clk(gclk));
	jdff dff_B_Kc7AVJjm8_2(.din(w_dff_B_BkAydNWi0_2),.dout(w_dff_B_Kc7AVJjm8_2),.clk(gclk));
	jdff dff_B_QoXqCVU15_2(.din(w_dff_B_Kc7AVJjm8_2),.dout(w_dff_B_QoXqCVU15_2),.clk(gclk));
	jdff dff_B_RkQ1Wc8J6_2(.din(w_dff_B_QoXqCVU15_2),.dout(w_dff_B_RkQ1Wc8J6_2),.clk(gclk));
	jdff dff_B_KsuwzJpz1_2(.din(w_dff_B_RkQ1Wc8J6_2),.dout(w_dff_B_KsuwzJpz1_2),.clk(gclk));
	jdff dff_B_aEWQcq2K0_2(.din(w_dff_B_KsuwzJpz1_2),.dout(w_dff_B_aEWQcq2K0_2),.clk(gclk));
	jdff dff_B_TdSHs97D6_2(.din(w_dff_B_aEWQcq2K0_2),.dout(w_dff_B_TdSHs97D6_2),.clk(gclk));
	jdff dff_B_ojYdJ6xP7_2(.din(w_dff_B_TdSHs97D6_2),.dout(w_dff_B_ojYdJ6xP7_2),.clk(gclk));
	jdff dff_B_2aqGnBmB3_2(.din(w_dff_B_ojYdJ6xP7_2),.dout(w_dff_B_2aqGnBmB3_2),.clk(gclk));
	jdff dff_B_BY9jdHMx3_2(.din(w_dff_B_2aqGnBmB3_2),.dout(w_dff_B_BY9jdHMx3_2),.clk(gclk));
	jdff dff_B_G75FPiZ94_2(.din(w_dff_B_BY9jdHMx3_2),.dout(w_dff_B_G75FPiZ94_2),.clk(gclk));
	jdff dff_B_KH1bkfDM3_2(.din(w_dff_B_G75FPiZ94_2),.dout(w_dff_B_KH1bkfDM3_2),.clk(gclk));
	jdff dff_B_ZCw7RZE63_2(.din(w_dff_B_KH1bkfDM3_2),.dout(w_dff_B_ZCw7RZE63_2),.clk(gclk));
	jdff dff_B_O5R55zZc6_2(.din(w_dff_B_ZCw7RZE63_2),.dout(w_dff_B_O5R55zZc6_2),.clk(gclk));
	jdff dff_B_CltihA214_2(.din(w_dff_B_O5R55zZc6_2),.dout(w_dff_B_CltihA214_2),.clk(gclk));
	jdff dff_B_NFs8nu665_2(.din(w_dff_B_CltihA214_2),.dout(w_dff_B_NFs8nu665_2),.clk(gclk));
	jdff dff_B_dA59S4zW5_2(.din(w_dff_B_NFs8nu665_2),.dout(w_dff_B_dA59S4zW5_2),.clk(gclk));
	jdff dff_B_wZS7RfwH9_2(.din(w_dff_B_dA59S4zW5_2),.dout(w_dff_B_wZS7RfwH9_2),.clk(gclk));
	jdff dff_B_ekZVA6Pp4_2(.din(w_dff_B_wZS7RfwH9_2),.dout(w_dff_B_ekZVA6Pp4_2),.clk(gclk));
	jdff dff_B_qDnt8Nwe4_2(.din(w_dff_B_ekZVA6Pp4_2),.dout(w_dff_B_qDnt8Nwe4_2),.clk(gclk));
	jdff dff_B_5gyJeHCz5_2(.din(w_dff_B_qDnt8Nwe4_2),.dout(w_dff_B_5gyJeHCz5_2),.clk(gclk));
	jdff dff_B_7IOPICYw1_2(.din(w_dff_B_5gyJeHCz5_2),.dout(w_dff_B_7IOPICYw1_2),.clk(gclk));
	jdff dff_B_3b8WpZfL0_2(.din(w_dff_B_7IOPICYw1_2),.dout(w_dff_B_3b8WpZfL0_2),.clk(gclk));
	jdff dff_B_YnabyG0G3_2(.din(w_dff_B_3b8WpZfL0_2),.dout(w_dff_B_YnabyG0G3_2),.clk(gclk));
	jdff dff_B_n77vf1nt9_2(.din(w_dff_B_YnabyG0G3_2),.dout(w_dff_B_n77vf1nt9_2),.clk(gclk));
	jdff dff_B_Vm42VOx80_2(.din(w_dff_B_n77vf1nt9_2),.dout(w_dff_B_Vm42VOx80_2),.clk(gclk));
	jdff dff_B_m0eMMI8i3_2(.din(w_dff_B_Vm42VOx80_2),.dout(w_dff_B_m0eMMI8i3_2),.clk(gclk));
	jdff dff_B_ep9J85lm5_1(.din(n1508),.dout(w_dff_B_ep9J85lm5_1),.clk(gclk));
	jdff dff_B_NITjvwZO1_2(.din(n1436),.dout(w_dff_B_NITjvwZO1_2),.clk(gclk));
	jdff dff_B_pp1IcoEZ3_2(.din(w_dff_B_NITjvwZO1_2),.dout(w_dff_B_pp1IcoEZ3_2),.clk(gclk));
	jdff dff_B_yCg6xIBm2_2(.din(w_dff_B_pp1IcoEZ3_2),.dout(w_dff_B_yCg6xIBm2_2),.clk(gclk));
	jdff dff_B_AXH3ceeX4_2(.din(w_dff_B_yCg6xIBm2_2),.dout(w_dff_B_AXH3ceeX4_2),.clk(gclk));
	jdff dff_B_hBxhxHyA9_2(.din(w_dff_B_AXH3ceeX4_2),.dout(w_dff_B_hBxhxHyA9_2),.clk(gclk));
	jdff dff_B_2VNxjfxP7_2(.din(w_dff_B_hBxhxHyA9_2),.dout(w_dff_B_2VNxjfxP7_2),.clk(gclk));
	jdff dff_B_jUKy0EVc6_2(.din(w_dff_B_2VNxjfxP7_2),.dout(w_dff_B_jUKy0EVc6_2),.clk(gclk));
	jdff dff_B_pVmGhPvx3_2(.din(w_dff_B_jUKy0EVc6_2),.dout(w_dff_B_pVmGhPvx3_2),.clk(gclk));
	jdff dff_B_uKayVfot0_2(.din(w_dff_B_pVmGhPvx3_2),.dout(w_dff_B_uKayVfot0_2),.clk(gclk));
	jdff dff_B_vvfc7eE66_2(.din(w_dff_B_uKayVfot0_2),.dout(w_dff_B_vvfc7eE66_2),.clk(gclk));
	jdff dff_B_5hX1zHPV4_2(.din(w_dff_B_vvfc7eE66_2),.dout(w_dff_B_5hX1zHPV4_2),.clk(gclk));
	jdff dff_B_dcXSkwkr4_2(.din(w_dff_B_5hX1zHPV4_2),.dout(w_dff_B_dcXSkwkr4_2),.clk(gclk));
	jdff dff_B_wirYtMQL7_2(.din(w_dff_B_dcXSkwkr4_2),.dout(w_dff_B_wirYtMQL7_2),.clk(gclk));
	jdff dff_B_o6umcOOP8_2(.din(w_dff_B_wirYtMQL7_2),.dout(w_dff_B_o6umcOOP8_2),.clk(gclk));
	jdff dff_B_d9CUyejE7_2(.din(w_dff_B_o6umcOOP8_2),.dout(w_dff_B_d9CUyejE7_2),.clk(gclk));
	jdff dff_B_L8ISDlfd1_2(.din(w_dff_B_d9CUyejE7_2),.dout(w_dff_B_L8ISDlfd1_2),.clk(gclk));
	jdff dff_B_j1J6srgp4_2(.din(w_dff_B_L8ISDlfd1_2),.dout(w_dff_B_j1J6srgp4_2),.clk(gclk));
	jdff dff_B_VQnKRV0Y2_2(.din(w_dff_B_j1J6srgp4_2),.dout(w_dff_B_VQnKRV0Y2_2),.clk(gclk));
	jdff dff_B_rhduM2fl6_2(.din(w_dff_B_VQnKRV0Y2_2),.dout(w_dff_B_rhduM2fl6_2),.clk(gclk));
	jdff dff_B_lG6L7IyP0_2(.din(w_dff_B_rhduM2fl6_2),.dout(w_dff_B_lG6L7IyP0_2),.clk(gclk));
	jdff dff_B_I4ezPKmf1_2(.din(w_dff_B_lG6L7IyP0_2),.dout(w_dff_B_I4ezPKmf1_2),.clk(gclk));
	jdff dff_B_I5Mn5VT17_2(.din(w_dff_B_I4ezPKmf1_2),.dout(w_dff_B_I5Mn5VT17_2),.clk(gclk));
	jdff dff_B_63fQgczl7_2(.din(w_dff_B_I5Mn5VT17_2),.dout(w_dff_B_63fQgczl7_2),.clk(gclk));
	jdff dff_B_stByCNqY7_2(.din(w_dff_B_63fQgczl7_2),.dout(w_dff_B_stByCNqY7_2),.clk(gclk));
	jdff dff_B_PQDJDI380_2(.din(w_dff_B_stByCNqY7_2),.dout(w_dff_B_PQDJDI380_2),.clk(gclk));
	jdff dff_B_zFRQ0nHT0_2(.din(w_dff_B_PQDJDI380_2),.dout(w_dff_B_zFRQ0nHT0_2),.clk(gclk));
	jdff dff_B_ErKhzT9D7_2(.din(w_dff_B_zFRQ0nHT0_2),.dout(w_dff_B_ErKhzT9D7_2),.clk(gclk));
	jdff dff_B_yXmbOzmP5_2(.din(w_dff_B_ErKhzT9D7_2),.dout(w_dff_B_yXmbOzmP5_2),.clk(gclk));
	jdff dff_B_T5upasdN9_2(.din(w_dff_B_yXmbOzmP5_2),.dout(w_dff_B_T5upasdN9_2),.clk(gclk));
	jdff dff_B_JtUGBNnw2_2(.din(w_dff_B_T5upasdN9_2),.dout(w_dff_B_JtUGBNnw2_2),.clk(gclk));
	jdff dff_B_hI6yFXJz7_2(.din(w_dff_B_JtUGBNnw2_2),.dout(w_dff_B_hI6yFXJz7_2),.clk(gclk));
	jdff dff_B_PNQIdWr74_2(.din(w_dff_B_hI6yFXJz7_2),.dout(w_dff_B_PNQIdWr74_2),.clk(gclk));
	jdff dff_B_wjpq9D6j9_2(.din(w_dff_B_PNQIdWr74_2),.dout(w_dff_B_wjpq9D6j9_2),.clk(gclk));
	jdff dff_B_vRvr2wr26_2(.din(w_dff_B_wjpq9D6j9_2),.dout(w_dff_B_vRvr2wr26_2),.clk(gclk));
	jdff dff_B_Nk3AB6I91_2(.din(w_dff_B_vRvr2wr26_2),.dout(w_dff_B_Nk3AB6I91_2),.clk(gclk));
	jdff dff_B_2ywxSxKj8_2(.din(w_dff_B_Nk3AB6I91_2),.dout(w_dff_B_2ywxSxKj8_2),.clk(gclk));
	jdff dff_B_HISQ8N1N8_2(.din(n1475),.dout(w_dff_B_HISQ8N1N8_2),.clk(gclk));
	jdff dff_B_bc8EOeQJ5_1(.din(n1437),.dout(w_dff_B_bc8EOeQJ5_1),.clk(gclk));
	jdff dff_B_9dobeQkJ7_2(.din(n1358),.dout(w_dff_B_9dobeQkJ7_2),.clk(gclk));
	jdff dff_B_jyVHoDC70_2(.din(w_dff_B_9dobeQkJ7_2),.dout(w_dff_B_jyVHoDC70_2),.clk(gclk));
	jdff dff_B_m7F28Hkb4_2(.din(w_dff_B_jyVHoDC70_2),.dout(w_dff_B_m7F28Hkb4_2),.clk(gclk));
	jdff dff_B_eMQ3XJKt9_2(.din(w_dff_B_m7F28Hkb4_2),.dout(w_dff_B_eMQ3XJKt9_2),.clk(gclk));
	jdff dff_B_fTpM45iT8_2(.din(w_dff_B_eMQ3XJKt9_2),.dout(w_dff_B_fTpM45iT8_2),.clk(gclk));
	jdff dff_B_hhwn8Kaf2_2(.din(w_dff_B_fTpM45iT8_2),.dout(w_dff_B_hhwn8Kaf2_2),.clk(gclk));
	jdff dff_B_1gBks4D78_2(.din(w_dff_B_hhwn8Kaf2_2),.dout(w_dff_B_1gBks4D78_2),.clk(gclk));
	jdff dff_B_EUu8PYPN4_2(.din(w_dff_B_1gBks4D78_2),.dout(w_dff_B_EUu8PYPN4_2),.clk(gclk));
	jdff dff_B_dRIsLWDc5_2(.din(w_dff_B_EUu8PYPN4_2),.dout(w_dff_B_dRIsLWDc5_2),.clk(gclk));
	jdff dff_B_okH6juCc3_2(.din(w_dff_B_dRIsLWDc5_2),.dout(w_dff_B_okH6juCc3_2),.clk(gclk));
	jdff dff_B_HZpdYgyn7_2(.din(w_dff_B_okH6juCc3_2),.dout(w_dff_B_HZpdYgyn7_2),.clk(gclk));
	jdff dff_B_Pj4hLcsP1_2(.din(w_dff_B_HZpdYgyn7_2),.dout(w_dff_B_Pj4hLcsP1_2),.clk(gclk));
	jdff dff_B_NYENvobe8_2(.din(w_dff_B_Pj4hLcsP1_2),.dout(w_dff_B_NYENvobe8_2),.clk(gclk));
	jdff dff_B_wzcWJJa17_2(.din(w_dff_B_NYENvobe8_2),.dout(w_dff_B_wzcWJJa17_2),.clk(gclk));
	jdff dff_B_Y17Tzvel4_2(.din(w_dff_B_wzcWJJa17_2),.dout(w_dff_B_Y17Tzvel4_2),.clk(gclk));
	jdff dff_B_OAL4d9VV7_2(.din(w_dff_B_Y17Tzvel4_2),.dout(w_dff_B_OAL4d9VV7_2),.clk(gclk));
	jdff dff_B_uFMc3xi21_2(.din(w_dff_B_OAL4d9VV7_2),.dout(w_dff_B_uFMc3xi21_2),.clk(gclk));
	jdff dff_B_1CWtZyUO2_2(.din(w_dff_B_uFMc3xi21_2),.dout(w_dff_B_1CWtZyUO2_2),.clk(gclk));
	jdff dff_B_6sOJFOLV6_2(.din(w_dff_B_1CWtZyUO2_2),.dout(w_dff_B_6sOJFOLV6_2),.clk(gclk));
	jdff dff_B_PLWr5jKS6_2(.din(w_dff_B_6sOJFOLV6_2),.dout(w_dff_B_PLWr5jKS6_2),.clk(gclk));
	jdff dff_B_74DTXMSh3_2(.din(w_dff_B_PLWr5jKS6_2),.dout(w_dff_B_74DTXMSh3_2),.clk(gclk));
	jdff dff_B_ajl8NgPG4_2(.din(w_dff_B_74DTXMSh3_2),.dout(w_dff_B_ajl8NgPG4_2),.clk(gclk));
	jdff dff_B_fMU1GJRk7_2(.din(w_dff_B_ajl8NgPG4_2),.dout(w_dff_B_fMU1GJRk7_2),.clk(gclk));
	jdff dff_B_hoNMd5JW0_2(.din(w_dff_B_fMU1GJRk7_2),.dout(w_dff_B_hoNMd5JW0_2),.clk(gclk));
	jdff dff_B_Yn3XMZPW3_2(.din(w_dff_B_hoNMd5JW0_2),.dout(w_dff_B_Yn3XMZPW3_2),.clk(gclk));
	jdff dff_B_muVvpKeL8_2(.din(w_dff_B_Yn3XMZPW3_2),.dout(w_dff_B_muVvpKeL8_2),.clk(gclk));
	jdff dff_B_ownsU5WY6_2(.din(w_dff_B_muVvpKeL8_2),.dout(w_dff_B_ownsU5WY6_2),.clk(gclk));
	jdff dff_B_KaOcZpno8_2(.din(w_dff_B_ownsU5WY6_2),.dout(w_dff_B_KaOcZpno8_2),.clk(gclk));
	jdff dff_B_X3GzVAcQ1_2(.din(w_dff_B_KaOcZpno8_2),.dout(w_dff_B_X3GzVAcQ1_2),.clk(gclk));
	jdff dff_B_0u3Qh3XZ2_2(.din(w_dff_B_X3GzVAcQ1_2),.dout(w_dff_B_0u3Qh3XZ2_2),.clk(gclk));
	jdff dff_B_5S0Pu4gx2_2(.din(w_dff_B_0u3Qh3XZ2_2),.dout(w_dff_B_5S0Pu4gx2_2),.clk(gclk));
	jdff dff_B_gtqgsyJ29_2(.din(w_dff_B_5S0Pu4gx2_2),.dout(w_dff_B_gtqgsyJ29_2),.clk(gclk));
	jdff dff_B_ytPP6zC89_2(.din(w_dff_B_gtqgsyJ29_2),.dout(w_dff_B_ytPP6zC89_2),.clk(gclk));
	jdff dff_B_1JzL5Mq57_2(.din(n1397),.dout(w_dff_B_1JzL5Mq57_2),.clk(gclk));
	jdff dff_B_WVn4gxIs4_1(.din(n1359),.dout(w_dff_B_WVn4gxIs4_1),.clk(gclk));
	jdff dff_B_ip10Dipr1_2(.din(n1273),.dout(w_dff_B_ip10Dipr1_2),.clk(gclk));
	jdff dff_B_F6lJWV9g8_2(.din(w_dff_B_ip10Dipr1_2),.dout(w_dff_B_F6lJWV9g8_2),.clk(gclk));
	jdff dff_B_ZeC5lp6w7_2(.din(w_dff_B_F6lJWV9g8_2),.dout(w_dff_B_ZeC5lp6w7_2),.clk(gclk));
	jdff dff_B_Fe3noJUt0_2(.din(w_dff_B_ZeC5lp6w7_2),.dout(w_dff_B_Fe3noJUt0_2),.clk(gclk));
	jdff dff_B_6rMTpEze6_2(.din(w_dff_B_Fe3noJUt0_2),.dout(w_dff_B_6rMTpEze6_2),.clk(gclk));
	jdff dff_B_iHGDDPCs5_2(.din(w_dff_B_6rMTpEze6_2),.dout(w_dff_B_iHGDDPCs5_2),.clk(gclk));
	jdff dff_B_qAzHfZTW8_2(.din(w_dff_B_iHGDDPCs5_2),.dout(w_dff_B_qAzHfZTW8_2),.clk(gclk));
	jdff dff_B_toU4PPUN8_2(.din(w_dff_B_qAzHfZTW8_2),.dout(w_dff_B_toU4PPUN8_2),.clk(gclk));
	jdff dff_B_ncnBoFdE2_2(.din(w_dff_B_toU4PPUN8_2),.dout(w_dff_B_ncnBoFdE2_2),.clk(gclk));
	jdff dff_B_skqtymb74_2(.din(w_dff_B_ncnBoFdE2_2),.dout(w_dff_B_skqtymb74_2),.clk(gclk));
	jdff dff_B_0VPZXGuf9_2(.din(w_dff_B_skqtymb74_2),.dout(w_dff_B_0VPZXGuf9_2),.clk(gclk));
	jdff dff_B_YBZzA1aF4_2(.din(w_dff_B_0VPZXGuf9_2),.dout(w_dff_B_YBZzA1aF4_2),.clk(gclk));
	jdff dff_B_apHUwt5q6_2(.din(w_dff_B_YBZzA1aF4_2),.dout(w_dff_B_apHUwt5q6_2),.clk(gclk));
	jdff dff_B_9iGDo3O46_2(.din(w_dff_B_apHUwt5q6_2),.dout(w_dff_B_9iGDo3O46_2),.clk(gclk));
	jdff dff_B_iAabzOLN2_2(.din(w_dff_B_9iGDo3O46_2),.dout(w_dff_B_iAabzOLN2_2),.clk(gclk));
	jdff dff_B_64YivDpv3_2(.din(w_dff_B_iAabzOLN2_2),.dout(w_dff_B_64YivDpv3_2),.clk(gclk));
	jdff dff_B_GIcp11qT1_2(.din(w_dff_B_64YivDpv3_2),.dout(w_dff_B_GIcp11qT1_2),.clk(gclk));
	jdff dff_B_Rr24kxsg3_2(.din(w_dff_B_GIcp11qT1_2),.dout(w_dff_B_Rr24kxsg3_2),.clk(gclk));
	jdff dff_B_oxBHb8iV9_2(.din(w_dff_B_Rr24kxsg3_2),.dout(w_dff_B_oxBHb8iV9_2),.clk(gclk));
	jdff dff_B_BEKKcG2v0_2(.din(w_dff_B_oxBHb8iV9_2),.dout(w_dff_B_BEKKcG2v0_2),.clk(gclk));
	jdff dff_B_uM1nMhGN2_2(.din(w_dff_B_BEKKcG2v0_2),.dout(w_dff_B_uM1nMhGN2_2),.clk(gclk));
	jdff dff_B_Z3txKOzB0_2(.din(w_dff_B_uM1nMhGN2_2),.dout(w_dff_B_Z3txKOzB0_2),.clk(gclk));
	jdff dff_B_NsuF8KsE1_2(.din(w_dff_B_Z3txKOzB0_2),.dout(w_dff_B_NsuF8KsE1_2),.clk(gclk));
	jdff dff_B_SAvm11bq7_2(.din(w_dff_B_NsuF8KsE1_2),.dout(w_dff_B_SAvm11bq7_2),.clk(gclk));
	jdff dff_B_L8G6ABRI2_2(.din(w_dff_B_SAvm11bq7_2),.dout(w_dff_B_L8G6ABRI2_2),.clk(gclk));
	jdff dff_B_oFuVGFgH8_2(.din(w_dff_B_L8G6ABRI2_2),.dout(w_dff_B_oFuVGFgH8_2),.clk(gclk));
	jdff dff_B_eFMZsobE9_2(.din(w_dff_B_oFuVGFgH8_2),.dout(w_dff_B_eFMZsobE9_2),.clk(gclk));
	jdff dff_B_2YLg9TQ78_2(.din(w_dff_B_eFMZsobE9_2),.dout(w_dff_B_2YLg9TQ78_2),.clk(gclk));
	jdff dff_B_T1HO2Rd15_2(.din(w_dff_B_2YLg9TQ78_2),.dout(w_dff_B_T1HO2Rd15_2),.clk(gclk));
	jdff dff_B_7zpv10YT7_2(.din(w_dff_B_T1HO2Rd15_2),.dout(w_dff_B_7zpv10YT7_2),.clk(gclk));
	jdff dff_B_mADqmqP18_2(.din(n1312),.dout(w_dff_B_mADqmqP18_2),.clk(gclk));
	jdff dff_B_nwJXkFV64_1(.din(n1274),.dout(w_dff_B_nwJXkFV64_1),.clk(gclk));
	jdff dff_B_LiWGV6py7_2(.din(n1183),.dout(w_dff_B_LiWGV6py7_2),.clk(gclk));
	jdff dff_B_We4PU8jH9_2(.din(w_dff_B_LiWGV6py7_2),.dout(w_dff_B_We4PU8jH9_2),.clk(gclk));
	jdff dff_B_lcrIB0qU5_2(.din(w_dff_B_We4PU8jH9_2),.dout(w_dff_B_lcrIB0qU5_2),.clk(gclk));
	jdff dff_B_cjjx011v3_2(.din(w_dff_B_lcrIB0qU5_2),.dout(w_dff_B_cjjx011v3_2),.clk(gclk));
	jdff dff_B_rrpxWGx76_2(.din(w_dff_B_cjjx011v3_2),.dout(w_dff_B_rrpxWGx76_2),.clk(gclk));
	jdff dff_B_zWgXi6xT9_2(.din(w_dff_B_rrpxWGx76_2),.dout(w_dff_B_zWgXi6xT9_2),.clk(gclk));
	jdff dff_B_eAkQYT9l8_2(.din(w_dff_B_zWgXi6xT9_2),.dout(w_dff_B_eAkQYT9l8_2),.clk(gclk));
	jdff dff_B_K8jmrcin0_2(.din(w_dff_B_eAkQYT9l8_2),.dout(w_dff_B_K8jmrcin0_2),.clk(gclk));
	jdff dff_B_Uqjnyzse5_2(.din(w_dff_B_K8jmrcin0_2),.dout(w_dff_B_Uqjnyzse5_2),.clk(gclk));
	jdff dff_B_2fxMLfWK8_2(.din(w_dff_B_Uqjnyzse5_2),.dout(w_dff_B_2fxMLfWK8_2),.clk(gclk));
	jdff dff_B_jAXTuAWY0_2(.din(w_dff_B_2fxMLfWK8_2),.dout(w_dff_B_jAXTuAWY0_2),.clk(gclk));
	jdff dff_B_WrljdxqX4_2(.din(w_dff_B_jAXTuAWY0_2),.dout(w_dff_B_WrljdxqX4_2),.clk(gclk));
	jdff dff_B_G8Sh7LQa3_2(.din(w_dff_B_WrljdxqX4_2),.dout(w_dff_B_G8Sh7LQa3_2),.clk(gclk));
	jdff dff_B_VyJhSFsX7_2(.din(w_dff_B_G8Sh7LQa3_2),.dout(w_dff_B_VyJhSFsX7_2),.clk(gclk));
	jdff dff_B_n4fjb4Hx4_2(.din(w_dff_B_VyJhSFsX7_2),.dout(w_dff_B_n4fjb4Hx4_2),.clk(gclk));
	jdff dff_B_ctJpDmhB3_2(.din(w_dff_B_n4fjb4Hx4_2),.dout(w_dff_B_ctJpDmhB3_2),.clk(gclk));
	jdff dff_B_dKvI9GS99_2(.din(w_dff_B_ctJpDmhB3_2),.dout(w_dff_B_dKvI9GS99_2),.clk(gclk));
	jdff dff_B_kzUkZZI13_2(.din(w_dff_B_dKvI9GS99_2),.dout(w_dff_B_kzUkZZI13_2),.clk(gclk));
	jdff dff_B_7ZeqhotU4_2(.din(w_dff_B_kzUkZZI13_2),.dout(w_dff_B_7ZeqhotU4_2),.clk(gclk));
	jdff dff_B_FgEaB1x25_2(.din(w_dff_B_7ZeqhotU4_2),.dout(w_dff_B_FgEaB1x25_2),.clk(gclk));
	jdff dff_B_M6ZF9rCk4_2(.din(w_dff_B_FgEaB1x25_2),.dout(w_dff_B_M6ZF9rCk4_2),.clk(gclk));
	jdff dff_B_mRnJoWnI9_2(.din(w_dff_B_M6ZF9rCk4_2),.dout(w_dff_B_mRnJoWnI9_2),.clk(gclk));
	jdff dff_B_uCuvAqPS5_2(.din(w_dff_B_mRnJoWnI9_2),.dout(w_dff_B_uCuvAqPS5_2),.clk(gclk));
	jdff dff_B_aZ27IuzA5_2(.din(w_dff_B_uCuvAqPS5_2),.dout(w_dff_B_aZ27IuzA5_2),.clk(gclk));
	jdff dff_B_x8ueRvEL4_2(.din(w_dff_B_aZ27IuzA5_2),.dout(w_dff_B_x8ueRvEL4_2),.clk(gclk));
	jdff dff_B_V7vgzhww6_2(.din(w_dff_B_x8ueRvEL4_2),.dout(w_dff_B_V7vgzhww6_2),.clk(gclk));
	jdff dff_B_44hlovNk6_2(.din(w_dff_B_V7vgzhww6_2),.dout(w_dff_B_44hlovNk6_2),.clk(gclk));
	jdff dff_B_MsvinaVe8_2(.din(n1221),.dout(w_dff_B_MsvinaVe8_2),.clk(gclk));
	jdff dff_B_k0AmojMX2_1(.din(n1184),.dout(w_dff_B_k0AmojMX2_1),.clk(gclk));
	jdff dff_B_dBxrUPST0_2(.din(n1079),.dout(w_dff_B_dBxrUPST0_2),.clk(gclk));
	jdff dff_B_6FQvDauU0_2(.din(w_dff_B_dBxrUPST0_2),.dout(w_dff_B_6FQvDauU0_2),.clk(gclk));
	jdff dff_B_On3kuz2s7_2(.din(w_dff_B_6FQvDauU0_2),.dout(w_dff_B_On3kuz2s7_2),.clk(gclk));
	jdff dff_B_i4PD0MDB5_2(.din(w_dff_B_On3kuz2s7_2),.dout(w_dff_B_i4PD0MDB5_2),.clk(gclk));
	jdff dff_B_ZAyC6yzB2_2(.din(w_dff_B_i4PD0MDB5_2),.dout(w_dff_B_ZAyC6yzB2_2),.clk(gclk));
	jdff dff_B_ACqCUdJK3_2(.din(w_dff_B_ZAyC6yzB2_2),.dout(w_dff_B_ACqCUdJK3_2),.clk(gclk));
	jdff dff_B_7wAoJzCG3_2(.din(w_dff_B_ACqCUdJK3_2),.dout(w_dff_B_7wAoJzCG3_2),.clk(gclk));
	jdff dff_B_5imdgR868_2(.din(w_dff_B_7wAoJzCG3_2),.dout(w_dff_B_5imdgR868_2),.clk(gclk));
	jdff dff_B_ezW95HMd0_2(.din(w_dff_B_5imdgR868_2),.dout(w_dff_B_ezW95HMd0_2),.clk(gclk));
	jdff dff_B_2hjVwVmF8_2(.din(w_dff_B_ezW95HMd0_2),.dout(w_dff_B_2hjVwVmF8_2),.clk(gclk));
	jdff dff_B_QBlXEqT10_2(.din(w_dff_B_2hjVwVmF8_2),.dout(w_dff_B_QBlXEqT10_2),.clk(gclk));
	jdff dff_B_uAyDHpfw6_2(.din(w_dff_B_QBlXEqT10_2),.dout(w_dff_B_uAyDHpfw6_2),.clk(gclk));
	jdff dff_B_zMbHL9B32_2(.din(w_dff_B_uAyDHpfw6_2),.dout(w_dff_B_zMbHL9B32_2),.clk(gclk));
	jdff dff_B_598SblUx5_2(.din(w_dff_B_zMbHL9B32_2),.dout(w_dff_B_598SblUx5_2),.clk(gclk));
	jdff dff_B_FFHcRYqL3_2(.din(w_dff_B_598SblUx5_2),.dout(w_dff_B_FFHcRYqL3_2),.clk(gclk));
	jdff dff_B_xkdNef0i0_2(.din(w_dff_B_FFHcRYqL3_2),.dout(w_dff_B_xkdNef0i0_2),.clk(gclk));
	jdff dff_B_mKinpzrY2_2(.din(w_dff_B_xkdNef0i0_2),.dout(w_dff_B_mKinpzrY2_2),.clk(gclk));
	jdff dff_B_sVlZZoUM2_2(.din(w_dff_B_mKinpzrY2_2),.dout(w_dff_B_sVlZZoUM2_2),.clk(gclk));
	jdff dff_B_wizdV6E65_2(.din(w_dff_B_sVlZZoUM2_2),.dout(w_dff_B_wizdV6E65_2),.clk(gclk));
	jdff dff_B_WmzQRrq68_2(.din(w_dff_B_wizdV6E65_2),.dout(w_dff_B_WmzQRrq68_2),.clk(gclk));
	jdff dff_B_RfEcLeU20_2(.din(w_dff_B_WmzQRrq68_2),.dout(w_dff_B_RfEcLeU20_2),.clk(gclk));
	jdff dff_B_hpnRPkPl8_2(.din(w_dff_B_RfEcLeU20_2),.dout(w_dff_B_hpnRPkPl8_2),.clk(gclk));
	jdff dff_B_BOHMR4jD0_2(.din(w_dff_B_hpnRPkPl8_2),.dout(w_dff_B_BOHMR4jD0_2),.clk(gclk));
	jdff dff_B_zmFlblHR9_2(.din(w_dff_B_BOHMR4jD0_2),.dout(w_dff_B_zmFlblHR9_2),.clk(gclk));
	jdff dff_B_ArKrp9Jo9_2(.din(n1123),.dout(w_dff_B_ArKrp9Jo9_2),.clk(gclk));
	jdff dff_B_IHPr1Lw29_1(.din(n1080),.dout(w_dff_B_IHPr1Lw29_1),.clk(gclk));
	jdff dff_B_tXrxXVHm9_2(.din(n981),.dout(w_dff_B_tXrxXVHm9_2),.clk(gclk));
	jdff dff_B_MrHLKQ150_2(.din(w_dff_B_tXrxXVHm9_2),.dout(w_dff_B_MrHLKQ150_2),.clk(gclk));
	jdff dff_B_ibuG9Ba73_2(.din(w_dff_B_MrHLKQ150_2),.dout(w_dff_B_ibuG9Ba73_2),.clk(gclk));
	jdff dff_B_naOkVaFF0_2(.din(w_dff_B_ibuG9Ba73_2),.dout(w_dff_B_naOkVaFF0_2),.clk(gclk));
	jdff dff_B_UTSv0xFq2_2(.din(w_dff_B_naOkVaFF0_2),.dout(w_dff_B_UTSv0xFq2_2),.clk(gclk));
	jdff dff_B_H2a9u2ng7_2(.din(w_dff_B_UTSv0xFq2_2),.dout(w_dff_B_H2a9u2ng7_2),.clk(gclk));
	jdff dff_B_ERHndalF5_2(.din(w_dff_B_H2a9u2ng7_2),.dout(w_dff_B_ERHndalF5_2),.clk(gclk));
	jdff dff_B_q2HbTIzh3_2(.din(w_dff_B_ERHndalF5_2),.dout(w_dff_B_q2HbTIzh3_2),.clk(gclk));
	jdff dff_B_wrcCZKqo9_2(.din(w_dff_B_q2HbTIzh3_2),.dout(w_dff_B_wrcCZKqo9_2),.clk(gclk));
	jdff dff_B_ZDwDkWAI9_2(.din(w_dff_B_wrcCZKqo9_2),.dout(w_dff_B_ZDwDkWAI9_2),.clk(gclk));
	jdff dff_B_HWroxUo33_2(.din(w_dff_B_ZDwDkWAI9_2),.dout(w_dff_B_HWroxUo33_2),.clk(gclk));
	jdff dff_B_g1Lf0It04_2(.din(w_dff_B_HWroxUo33_2),.dout(w_dff_B_g1Lf0It04_2),.clk(gclk));
	jdff dff_B_e6WgFQ6R8_2(.din(w_dff_B_g1Lf0It04_2),.dout(w_dff_B_e6WgFQ6R8_2),.clk(gclk));
	jdff dff_B_kpoUAvar0_2(.din(w_dff_B_e6WgFQ6R8_2),.dout(w_dff_B_kpoUAvar0_2),.clk(gclk));
	jdff dff_B_5xcht1sV5_2(.din(w_dff_B_kpoUAvar0_2),.dout(w_dff_B_5xcht1sV5_2),.clk(gclk));
	jdff dff_B_LIuaEXWL2_2(.din(w_dff_B_5xcht1sV5_2),.dout(w_dff_B_LIuaEXWL2_2),.clk(gclk));
	jdff dff_B_JpvsrTgi6_2(.din(w_dff_B_LIuaEXWL2_2),.dout(w_dff_B_JpvsrTgi6_2),.clk(gclk));
	jdff dff_B_j5B9MQpc4_2(.din(w_dff_B_JpvsrTgi6_2),.dout(w_dff_B_j5B9MQpc4_2),.clk(gclk));
	jdff dff_B_0d3qYfrT5_2(.din(w_dff_B_j5B9MQpc4_2),.dout(w_dff_B_0d3qYfrT5_2),.clk(gclk));
	jdff dff_B_NlFy0QL04_2(.din(w_dff_B_0d3qYfrT5_2),.dout(w_dff_B_NlFy0QL04_2),.clk(gclk));
	jdff dff_B_AU6jyrFE3_2(.din(w_dff_B_NlFy0QL04_2),.dout(w_dff_B_AU6jyrFE3_2),.clk(gclk));
	jdff dff_B_hOikBsCD4_2(.din(n1018),.dout(w_dff_B_hOikBsCD4_2),.clk(gclk));
	jdff dff_B_xA5TsFm41_1(.din(n982),.dout(w_dff_B_xA5TsFm41_1),.clk(gclk));
	jdff dff_B_5Xu7gypW2_2(.din(n876),.dout(w_dff_B_5Xu7gypW2_2),.clk(gclk));
	jdff dff_B_VbfjyOeY5_2(.din(w_dff_B_5Xu7gypW2_2),.dout(w_dff_B_VbfjyOeY5_2),.clk(gclk));
	jdff dff_B_rPfXnYEv0_2(.din(w_dff_B_VbfjyOeY5_2),.dout(w_dff_B_rPfXnYEv0_2),.clk(gclk));
	jdff dff_B_Whxa2VIo9_2(.din(w_dff_B_rPfXnYEv0_2),.dout(w_dff_B_Whxa2VIo9_2),.clk(gclk));
	jdff dff_B_JbtUBMFH5_2(.din(w_dff_B_Whxa2VIo9_2),.dout(w_dff_B_JbtUBMFH5_2),.clk(gclk));
	jdff dff_B_eCibOGKe4_2(.din(w_dff_B_JbtUBMFH5_2),.dout(w_dff_B_eCibOGKe4_2),.clk(gclk));
	jdff dff_B_SofNfQdv7_2(.din(w_dff_B_eCibOGKe4_2),.dout(w_dff_B_SofNfQdv7_2),.clk(gclk));
	jdff dff_B_DxpG3HVZ7_2(.din(w_dff_B_SofNfQdv7_2),.dout(w_dff_B_DxpG3HVZ7_2),.clk(gclk));
	jdff dff_B_UMPJEe397_2(.din(w_dff_B_DxpG3HVZ7_2),.dout(w_dff_B_UMPJEe397_2),.clk(gclk));
	jdff dff_B_DEN1JuF13_2(.din(w_dff_B_UMPJEe397_2),.dout(w_dff_B_DEN1JuF13_2),.clk(gclk));
	jdff dff_B_SvVeqdPa7_2(.din(w_dff_B_DEN1JuF13_2),.dout(w_dff_B_SvVeqdPa7_2),.clk(gclk));
	jdff dff_B_jwUptlux1_2(.din(w_dff_B_SvVeqdPa7_2),.dout(w_dff_B_jwUptlux1_2),.clk(gclk));
	jdff dff_B_WFlrYD1e1_2(.din(w_dff_B_jwUptlux1_2),.dout(w_dff_B_WFlrYD1e1_2),.clk(gclk));
	jdff dff_B_jiy5FE7l9_2(.din(w_dff_B_WFlrYD1e1_2),.dout(w_dff_B_jiy5FE7l9_2),.clk(gclk));
	jdff dff_B_BeVZ6VZy0_2(.din(w_dff_B_jiy5FE7l9_2),.dout(w_dff_B_BeVZ6VZy0_2),.clk(gclk));
	jdff dff_B_hipvSVQU7_2(.din(w_dff_B_BeVZ6VZy0_2),.dout(w_dff_B_hipvSVQU7_2),.clk(gclk));
	jdff dff_B_LkHXZCBK7_2(.din(w_dff_B_hipvSVQU7_2),.dout(w_dff_B_LkHXZCBK7_2),.clk(gclk));
	jdff dff_B_pfabGU1z4_2(.din(w_dff_B_LkHXZCBK7_2),.dout(w_dff_B_pfabGU1z4_2),.clk(gclk));
	jdff dff_B_n9EISm401_2(.din(n913),.dout(w_dff_B_n9EISm401_2),.clk(gclk));
	jdff dff_B_HJQyML745_1(.din(n877),.dout(w_dff_B_HJQyML745_1),.clk(gclk));
	jdff dff_B_wQfdFuV10_2(.din(n777),.dout(w_dff_B_wQfdFuV10_2),.clk(gclk));
	jdff dff_B_o73wuKI98_2(.din(w_dff_B_wQfdFuV10_2),.dout(w_dff_B_o73wuKI98_2),.clk(gclk));
	jdff dff_B_wmM4FHRy8_2(.din(w_dff_B_o73wuKI98_2),.dout(w_dff_B_wmM4FHRy8_2),.clk(gclk));
	jdff dff_B_3FrgMzfP3_2(.din(w_dff_B_wmM4FHRy8_2),.dout(w_dff_B_3FrgMzfP3_2),.clk(gclk));
	jdff dff_B_zzCFyGPl5_2(.din(w_dff_B_3FrgMzfP3_2),.dout(w_dff_B_zzCFyGPl5_2),.clk(gclk));
	jdff dff_B_CTrWC2XS6_2(.din(w_dff_B_zzCFyGPl5_2),.dout(w_dff_B_CTrWC2XS6_2),.clk(gclk));
	jdff dff_B_7bFV2QGw0_2(.din(w_dff_B_CTrWC2XS6_2),.dout(w_dff_B_7bFV2QGw0_2),.clk(gclk));
	jdff dff_B_NeFY834T1_2(.din(w_dff_B_7bFV2QGw0_2),.dout(w_dff_B_NeFY834T1_2),.clk(gclk));
	jdff dff_B_7VkI8jLT7_2(.din(w_dff_B_NeFY834T1_2),.dout(w_dff_B_7VkI8jLT7_2),.clk(gclk));
	jdff dff_B_i1IxUYqg2_2(.din(w_dff_B_7VkI8jLT7_2),.dout(w_dff_B_i1IxUYqg2_2),.clk(gclk));
	jdff dff_B_knIISLSD0_2(.din(w_dff_B_i1IxUYqg2_2),.dout(w_dff_B_knIISLSD0_2),.clk(gclk));
	jdff dff_B_lARREP0g7_2(.din(w_dff_B_knIISLSD0_2),.dout(w_dff_B_lARREP0g7_2),.clk(gclk));
	jdff dff_B_g7j7Yk6r6_2(.din(w_dff_B_lARREP0g7_2),.dout(w_dff_B_g7j7Yk6r6_2),.clk(gclk));
	jdff dff_B_XkKe7h4n6_2(.din(w_dff_B_g7j7Yk6r6_2),.dout(w_dff_B_XkKe7h4n6_2),.clk(gclk));
	jdff dff_B_dOQjWle73_2(.din(w_dff_B_XkKe7h4n6_2),.dout(w_dff_B_dOQjWle73_2),.clk(gclk));
	jdff dff_B_yEpiPgRN8_2(.din(n807),.dout(w_dff_B_yEpiPgRN8_2),.clk(gclk));
	jdff dff_B_bSQO3Iix9_1(.din(n778),.dout(w_dff_B_bSQO3Iix9_1),.clk(gclk));
	jdff dff_B_KbwQes492_2(.din(n684),.dout(w_dff_B_KbwQes492_2),.clk(gclk));
	jdff dff_B_IXmf1d398_2(.din(w_dff_B_KbwQes492_2),.dout(w_dff_B_IXmf1d398_2),.clk(gclk));
	jdff dff_B_ix1OoRRr9_2(.din(w_dff_B_IXmf1d398_2),.dout(w_dff_B_ix1OoRRr9_2),.clk(gclk));
	jdff dff_B_uCJoVFSw0_2(.din(w_dff_B_ix1OoRRr9_2),.dout(w_dff_B_uCJoVFSw0_2),.clk(gclk));
	jdff dff_B_5xjfZ3Wp0_2(.din(w_dff_B_uCJoVFSw0_2),.dout(w_dff_B_5xjfZ3Wp0_2),.clk(gclk));
	jdff dff_B_X1viEgLQ7_2(.din(w_dff_B_5xjfZ3Wp0_2),.dout(w_dff_B_X1viEgLQ7_2),.clk(gclk));
	jdff dff_B_YuiNqHBZ8_2(.din(w_dff_B_X1viEgLQ7_2),.dout(w_dff_B_YuiNqHBZ8_2),.clk(gclk));
	jdff dff_B_YOyAP99l4_2(.din(w_dff_B_YuiNqHBZ8_2),.dout(w_dff_B_YOyAP99l4_2),.clk(gclk));
	jdff dff_B_Uk4p2vjt6_2(.din(w_dff_B_YOyAP99l4_2),.dout(w_dff_B_Uk4p2vjt6_2),.clk(gclk));
	jdff dff_B_oQsncDie8_2(.din(w_dff_B_Uk4p2vjt6_2),.dout(w_dff_B_oQsncDie8_2),.clk(gclk));
	jdff dff_B_PqihfLAO8_2(.din(w_dff_B_oQsncDie8_2),.dout(w_dff_B_PqihfLAO8_2),.clk(gclk));
	jdff dff_B_7W6IBFpX8_2(.din(w_dff_B_PqihfLAO8_2),.dout(w_dff_B_7W6IBFpX8_2),.clk(gclk));
	jdff dff_B_Q5STwsBo3_2(.din(n707),.dout(w_dff_B_Q5STwsBo3_2),.clk(gclk));
	jdff dff_B_vavzs6245_1(.din(n685),.dout(w_dff_B_vavzs6245_1),.clk(gclk));
	jdff dff_B_uFybdbnK0_2(.din(n598),.dout(w_dff_B_uFybdbnK0_2),.clk(gclk));
	jdff dff_B_0LVi9f7f4_2(.din(w_dff_B_uFybdbnK0_2),.dout(w_dff_B_0LVi9f7f4_2),.clk(gclk));
	jdff dff_B_ZR15t9k95_2(.din(w_dff_B_0LVi9f7f4_2),.dout(w_dff_B_ZR15t9k95_2),.clk(gclk));
	jdff dff_B_uoKljbTd4_2(.din(w_dff_B_ZR15t9k95_2),.dout(w_dff_B_uoKljbTd4_2),.clk(gclk));
	jdff dff_B_GalnD0kl1_2(.din(w_dff_B_uoKljbTd4_2),.dout(w_dff_B_GalnD0kl1_2),.clk(gclk));
	jdff dff_B_ykNEyVAn8_2(.din(w_dff_B_GalnD0kl1_2),.dout(w_dff_B_ykNEyVAn8_2),.clk(gclk));
	jdff dff_B_WjD1AETW3_2(.din(w_dff_B_ykNEyVAn8_2),.dout(w_dff_B_WjD1AETW3_2),.clk(gclk));
	jdff dff_B_bsuqZ2859_2(.din(w_dff_B_WjD1AETW3_2),.dout(w_dff_B_bsuqZ2859_2),.clk(gclk));
	jdff dff_B_jZe4YHWU3_2(.din(w_dff_B_bsuqZ2859_2),.dout(w_dff_B_jZe4YHWU3_2),.clk(gclk));
	jdff dff_B_OhS1WdKY6_2(.din(n614),.dout(w_dff_B_OhS1WdKY6_2),.clk(gclk));
	jdff dff_B_Y11zjUIr9_2(.din(w_dff_B_OhS1WdKY6_2),.dout(w_dff_B_Y11zjUIr9_2),.clk(gclk));
	jdff dff_B_2NBhPVEo0_1(.din(n599),.dout(w_dff_B_2NBhPVEo0_1),.clk(gclk));
	jdff dff_B_yhRwLhSl0_1(.din(w_dff_B_2NBhPVEo0_1),.dout(w_dff_B_yhRwLhSl0_1),.clk(gclk));
	jdff dff_B_h5csbh3Q4_1(.din(w_dff_B_yhRwLhSl0_1),.dout(w_dff_B_h5csbh3Q4_1),.clk(gclk));
	jdff dff_B_A6id4RZi6_1(.din(w_dff_B_h5csbh3Q4_1),.dout(w_dff_B_A6id4RZi6_1),.clk(gclk));
	jdff dff_B_tz6VrQ7D8_1(.din(w_dff_B_A6id4RZi6_1),.dout(w_dff_B_tz6VrQ7D8_1),.clk(gclk));
	jdff dff_B_CbMh0etk8_1(.din(w_dff_B_tz6VrQ7D8_1),.dout(w_dff_B_CbMh0etk8_1),.clk(gclk));
	jdff dff_B_clarPqnr6_0(.din(n528),.dout(w_dff_B_clarPqnr6_0),.clk(gclk));
	jdff dff_B_5EYqdB1x0_0(.din(w_dff_B_clarPqnr6_0),.dout(w_dff_B_5EYqdB1x0_0),.clk(gclk));
	jdff dff_A_yizNcz2A1_0(.dout(w_n527_0[0]),.din(w_dff_A_yizNcz2A1_0),.clk(gclk));
	jdff dff_A_sFCCDAuD8_0(.dout(w_dff_A_yizNcz2A1_0),.din(w_dff_A_sFCCDAuD8_0),.clk(gclk));
	jdff dff_A_BnbUiBaX3_0(.dout(w_dff_A_sFCCDAuD8_0),.din(w_dff_A_BnbUiBaX3_0),.clk(gclk));
	jdff dff_B_pIrr73m08_1(.din(n521),.dout(w_dff_B_pIrr73m08_1),.clk(gclk));
	jdff dff_A_VEjDMFPq4_0(.dout(w_n446_0[0]),.din(w_dff_A_VEjDMFPq4_0),.clk(gclk));
	jdff dff_A_SAfrAM5U4_1(.dout(w_n446_0[1]),.din(w_dff_A_SAfrAM5U4_1),.clk(gclk));
	jdff dff_A_DzAcwloZ4_1(.dout(w_dff_A_SAfrAM5U4_1),.din(w_dff_A_DzAcwloZ4_1),.clk(gclk));
	jdff dff_A_ajZXznoi4_1(.dout(w_n519_0[1]),.din(w_dff_A_ajZXznoi4_1),.clk(gclk));
	jdff dff_A_2oHCCgGu6_1(.dout(w_dff_A_ajZXznoi4_1),.din(w_dff_A_2oHCCgGu6_1),.clk(gclk));
	jdff dff_A_BK8X57VK0_1(.dout(w_dff_A_2oHCCgGu6_1),.din(w_dff_A_BK8X57VK0_1),.clk(gclk));
	jdff dff_A_PbKr4Kqu4_1(.dout(w_dff_A_BK8X57VK0_1),.din(w_dff_A_PbKr4Kqu4_1),.clk(gclk));
	jdff dff_A_0GWR2Htb6_1(.dout(w_dff_A_PbKr4Kqu4_1),.din(w_dff_A_0GWR2Htb6_1),.clk(gclk));
	jdff dff_A_6STtgGwI6_1(.dout(w_dff_A_0GWR2Htb6_1),.din(w_dff_A_6STtgGwI6_1),.clk(gclk));
	jdff dff_B_TCewL5c97_1(.din(n1760),.dout(w_dff_B_TCewL5c97_1),.clk(gclk));
	jdff dff_A_gs11IcZb5_1(.dout(w_n1728_0[1]),.din(w_dff_A_gs11IcZb5_1),.clk(gclk));
	jdff dff_B_ZNA61zx23_1(.din(n1726),.dout(w_dff_B_ZNA61zx23_1),.clk(gclk));
	jdff dff_B_TkY1yLGK6_2(.din(n1684),.dout(w_dff_B_TkY1yLGK6_2),.clk(gclk));
	jdff dff_B_diW2C7mX8_2(.din(w_dff_B_TkY1yLGK6_2),.dout(w_dff_B_diW2C7mX8_2),.clk(gclk));
	jdff dff_B_rE5T2yVe7_2(.din(w_dff_B_diW2C7mX8_2),.dout(w_dff_B_rE5T2yVe7_2),.clk(gclk));
	jdff dff_B_CS8zggMj5_2(.din(w_dff_B_rE5T2yVe7_2),.dout(w_dff_B_CS8zggMj5_2),.clk(gclk));
	jdff dff_B_b2mo3lKz6_2(.din(w_dff_B_CS8zggMj5_2),.dout(w_dff_B_b2mo3lKz6_2),.clk(gclk));
	jdff dff_B_KLT5Lpxt9_2(.din(w_dff_B_b2mo3lKz6_2),.dout(w_dff_B_KLT5Lpxt9_2),.clk(gclk));
	jdff dff_B_b3FesVu59_2(.din(w_dff_B_KLT5Lpxt9_2),.dout(w_dff_B_b3FesVu59_2),.clk(gclk));
	jdff dff_B_Ph3YzaFY7_2(.din(w_dff_B_b3FesVu59_2),.dout(w_dff_B_Ph3YzaFY7_2),.clk(gclk));
	jdff dff_B_ANayHqti9_2(.din(w_dff_B_Ph3YzaFY7_2),.dout(w_dff_B_ANayHqti9_2),.clk(gclk));
	jdff dff_B_4JXILDJZ6_2(.din(w_dff_B_ANayHqti9_2),.dout(w_dff_B_4JXILDJZ6_2),.clk(gclk));
	jdff dff_B_CfMFsKap0_2(.din(w_dff_B_4JXILDJZ6_2),.dout(w_dff_B_CfMFsKap0_2),.clk(gclk));
	jdff dff_B_RWGSRGPx5_2(.din(w_dff_B_CfMFsKap0_2),.dout(w_dff_B_RWGSRGPx5_2),.clk(gclk));
	jdff dff_B_9K3JBp0j7_2(.din(w_dff_B_RWGSRGPx5_2),.dout(w_dff_B_9K3JBp0j7_2),.clk(gclk));
	jdff dff_B_zJqTLJr99_2(.din(w_dff_B_9K3JBp0j7_2),.dout(w_dff_B_zJqTLJr99_2),.clk(gclk));
	jdff dff_B_99CbURTR4_2(.din(w_dff_B_zJqTLJr99_2),.dout(w_dff_B_99CbURTR4_2),.clk(gclk));
	jdff dff_B_GI3UMVU34_2(.din(w_dff_B_99CbURTR4_2),.dout(w_dff_B_GI3UMVU34_2),.clk(gclk));
	jdff dff_B_5KSbgHdb9_2(.din(w_dff_B_GI3UMVU34_2),.dout(w_dff_B_5KSbgHdb9_2),.clk(gclk));
	jdff dff_B_eGCNUpTC8_2(.din(w_dff_B_5KSbgHdb9_2),.dout(w_dff_B_eGCNUpTC8_2),.clk(gclk));
	jdff dff_B_bu3eTSlq2_2(.din(w_dff_B_eGCNUpTC8_2),.dout(w_dff_B_bu3eTSlq2_2),.clk(gclk));
	jdff dff_B_9otfr0AT1_2(.din(w_dff_B_bu3eTSlq2_2),.dout(w_dff_B_9otfr0AT1_2),.clk(gclk));
	jdff dff_B_eh42FrmY0_2(.din(w_dff_B_9otfr0AT1_2),.dout(w_dff_B_eh42FrmY0_2),.clk(gclk));
	jdff dff_B_rawarsQ76_2(.din(w_dff_B_eh42FrmY0_2),.dout(w_dff_B_rawarsQ76_2),.clk(gclk));
	jdff dff_B_FgThDuMj4_2(.din(w_dff_B_rawarsQ76_2),.dout(w_dff_B_FgThDuMj4_2),.clk(gclk));
	jdff dff_B_vGmS6IKl5_2(.din(w_dff_B_FgThDuMj4_2),.dout(w_dff_B_vGmS6IKl5_2),.clk(gclk));
	jdff dff_B_0C2ytVHC6_2(.din(w_dff_B_vGmS6IKl5_2),.dout(w_dff_B_0C2ytVHC6_2),.clk(gclk));
	jdff dff_B_Jq9SG4xc0_2(.din(w_dff_B_0C2ytVHC6_2),.dout(w_dff_B_Jq9SG4xc0_2),.clk(gclk));
	jdff dff_B_fmhu7x7C5_2(.din(w_dff_B_Jq9SG4xc0_2),.dout(w_dff_B_fmhu7x7C5_2),.clk(gclk));
	jdff dff_B_rWFzzuz68_2(.din(w_dff_B_fmhu7x7C5_2),.dout(w_dff_B_rWFzzuz68_2),.clk(gclk));
	jdff dff_B_F5bXzkmW5_2(.din(w_dff_B_rWFzzuz68_2),.dout(w_dff_B_F5bXzkmW5_2),.clk(gclk));
	jdff dff_B_n9uHyAWm4_2(.din(w_dff_B_F5bXzkmW5_2),.dout(w_dff_B_n9uHyAWm4_2),.clk(gclk));
	jdff dff_B_UWOLfndn8_2(.din(w_dff_B_n9uHyAWm4_2),.dout(w_dff_B_UWOLfndn8_2),.clk(gclk));
	jdff dff_B_oXm7oNef5_2(.din(w_dff_B_UWOLfndn8_2),.dout(w_dff_B_oXm7oNef5_2),.clk(gclk));
	jdff dff_B_CBNzjB7B2_2(.din(w_dff_B_oXm7oNef5_2),.dout(w_dff_B_CBNzjB7B2_2),.clk(gclk));
	jdff dff_B_Syiaelsg1_2(.din(w_dff_B_CBNzjB7B2_2),.dout(w_dff_B_Syiaelsg1_2),.clk(gclk));
	jdff dff_B_3zQJlg3H0_2(.din(w_dff_B_Syiaelsg1_2),.dout(w_dff_B_3zQJlg3H0_2),.clk(gclk));
	jdff dff_B_JI51UZ669_2(.din(w_dff_B_3zQJlg3H0_2),.dout(w_dff_B_JI51UZ669_2),.clk(gclk));
	jdff dff_B_vzn2Bcph8_2(.din(w_dff_B_JI51UZ669_2),.dout(w_dff_B_vzn2Bcph8_2),.clk(gclk));
	jdff dff_B_ppiBzVLm1_2(.din(w_dff_B_vzn2Bcph8_2),.dout(w_dff_B_ppiBzVLm1_2),.clk(gclk));
	jdff dff_B_Mftj1Eta7_2(.din(w_dff_B_ppiBzVLm1_2),.dout(w_dff_B_Mftj1Eta7_2),.clk(gclk));
	jdff dff_B_O4UpiI2e8_2(.din(w_dff_B_Mftj1Eta7_2),.dout(w_dff_B_O4UpiI2e8_2),.clk(gclk));
	jdff dff_B_eRtSiULM4_2(.din(w_dff_B_O4UpiI2e8_2),.dout(w_dff_B_eRtSiULM4_2),.clk(gclk));
	jdff dff_B_aspaOuBq0_2(.din(w_dff_B_eRtSiULM4_2),.dout(w_dff_B_aspaOuBq0_2),.clk(gclk));
	jdff dff_B_9a1SXeoi0_2(.din(w_dff_B_aspaOuBq0_2),.dout(w_dff_B_9a1SXeoi0_2),.clk(gclk));
	jdff dff_B_lWuhQ7km8_2(.din(w_dff_B_9a1SXeoi0_2),.dout(w_dff_B_lWuhQ7km8_2),.clk(gclk));
	jdff dff_B_yP0Jf2nB5_2(.din(w_dff_B_lWuhQ7km8_2),.dout(w_dff_B_yP0Jf2nB5_2),.clk(gclk));
	jdff dff_B_JNbSNTFf9_2(.din(w_dff_B_yP0Jf2nB5_2),.dout(w_dff_B_JNbSNTFf9_2),.clk(gclk));
	jdff dff_B_mAJPjSWK4_2(.din(w_dff_B_JNbSNTFf9_2),.dout(w_dff_B_mAJPjSWK4_2),.clk(gclk));
	jdff dff_B_tcULOzcr5_2(.din(w_dff_B_mAJPjSWK4_2),.dout(w_dff_B_tcULOzcr5_2),.clk(gclk));
	jdff dff_B_1pDKIZ093_2(.din(w_dff_B_tcULOzcr5_2),.dout(w_dff_B_1pDKIZ093_2),.clk(gclk));
	jdff dff_B_N2jdzGk90_2(.din(n1687),.dout(w_dff_B_N2jdzGk90_2),.clk(gclk));
	jdff dff_B_OD8zsOFz3_1(.din(n1685),.dout(w_dff_B_OD8zsOFz3_1),.clk(gclk));
	jdff dff_B_Le2aNLXW1_2(.din(n1633),.dout(w_dff_B_Le2aNLXW1_2),.clk(gclk));
	jdff dff_B_X940kKQk4_2(.din(w_dff_B_Le2aNLXW1_2),.dout(w_dff_B_X940kKQk4_2),.clk(gclk));
	jdff dff_B_WQWOCGvC2_2(.din(w_dff_B_X940kKQk4_2),.dout(w_dff_B_WQWOCGvC2_2),.clk(gclk));
	jdff dff_B_KKy3QRSz1_2(.din(w_dff_B_WQWOCGvC2_2),.dout(w_dff_B_KKy3QRSz1_2),.clk(gclk));
	jdff dff_B_Dbr6G2PZ9_2(.din(w_dff_B_KKy3QRSz1_2),.dout(w_dff_B_Dbr6G2PZ9_2),.clk(gclk));
	jdff dff_B_G0ADHMuC9_2(.din(w_dff_B_Dbr6G2PZ9_2),.dout(w_dff_B_G0ADHMuC9_2),.clk(gclk));
	jdff dff_B_oEcDhbXk8_2(.din(w_dff_B_G0ADHMuC9_2),.dout(w_dff_B_oEcDhbXk8_2),.clk(gclk));
	jdff dff_B_l0jqOEwI9_2(.din(w_dff_B_oEcDhbXk8_2),.dout(w_dff_B_l0jqOEwI9_2),.clk(gclk));
	jdff dff_B_NZYnER997_2(.din(w_dff_B_l0jqOEwI9_2),.dout(w_dff_B_NZYnER997_2),.clk(gclk));
	jdff dff_B_9eFXj9rZ8_2(.din(w_dff_B_NZYnER997_2),.dout(w_dff_B_9eFXj9rZ8_2),.clk(gclk));
	jdff dff_B_lATkhR9x2_2(.din(w_dff_B_9eFXj9rZ8_2),.dout(w_dff_B_lATkhR9x2_2),.clk(gclk));
	jdff dff_B_fjW11Uiw8_2(.din(w_dff_B_lATkhR9x2_2),.dout(w_dff_B_fjW11Uiw8_2),.clk(gclk));
	jdff dff_B_AWWjL4iO7_2(.din(w_dff_B_fjW11Uiw8_2),.dout(w_dff_B_AWWjL4iO7_2),.clk(gclk));
	jdff dff_B_9zkz70Iy8_2(.din(w_dff_B_AWWjL4iO7_2),.dout(w_dff_B_9zkz70Iy8_2),.clk(gclk));
	jdff dff_B_4JdnowO17_2(.din(w_dff_B_9zkz70Iy8_2),.dout(w_dff_B_4JdnowO17_2),.clk(gclk));
	jdff dff_B_PFUZM9UN2_2(.din(w_dff_B_4JdnowO17_2),.dout(w_dff_B_PFUZM9UN2_2),.clk(gclk));
	jdff dff_B_eNZAHqET7_2(.din(w_dff_B_PFUZM9UN2_2),.dout(w_dff_B_eNZAHqET7_2),.clk(gclk));
	jdff dff_B_23GPd94w8_2(.din(w_dff_B_eNZAHqET7_2),.dout(w_dff_B_23GPd94w8_2),.clk(gclk));
	jdff dff_B_U06PEwPw6_2(.din(w_dff_B_23GPd94w8_2),.dout(w_dff_B_U06PEwPw6_2),.clk(gclk));
	jdff dff_B_svnKd5Hb2_2(.din(w_dff_B_U06PEwPw6_2),.dout(w_dff_B_svnKd5Hb2_2),.clk(gclk));
	jdff dff_B_WolfQb4C1_2(.din(w_dff_B_svnKd5Hb2_2),.dout(w_dff_B_WolfQb4C1_2),.clk(gclk));
	jdff dff_B_8sef5ni97_2(.din(w_dff_B_WolfQb4C1_2),.dout(w_dff_B_8sef5ni97_2),.clk(gclk));
	jdff dff_B_COQEwRTS3_2(.din(w_dff_B_8sef5ni97_2),.dout(w_dff_B_COQEwRTS3_2),.clk(gclk));
	jdff dff_B_eNKHHtb45_2(.din(w_dff_B_COQEwRTS3_2),.dout(w_dff_B_eNKHHtb45_2),.clk(gclk));
	jdff dff_B_vZM6LUyC7_2(.din(w_dff_B_eNKHHtb45_2),.dout(w_dff_B_vZM6LUyC7_2),.clk(gclk));
	jdff dff_B_O9ovA19C0_2(.din(w_dff_B_vZM6LUyC7_2),.dout(w_dff_B_O9ovA19C0_2),.clk(gclk));
	jdff dff_B_0ayl8ijC5_2(.din(w_dff_B_O9ovA19C0_2),.dout(w_dff_B_0ayl8ijC5_2),.clk(gclk));
	jdff dff_B_B3NPte5y2_2(.din(w_dff_B_0ayl8ijC5_2),.dout(w_dff_B_B3NPte5y2_2),.clk(gclk));
	jdff dff_B_pkTmhiov8_2(.din(w_dff_B_B3NPte5y2_2),.dout(w_dff_B_pkTmhiov8_2),.clk(gclk));
	jdff dff_B_bU4njUtF6_2(.din(w_dff_B_pkTmhiov8_2),.dout(w_dff_B_bU4njUtF6_2),.clk(gclk));
	jdff dff_B_h9EIukWF0_2(.din(w_dff_B_bU4njUtF6_2),.dout(w_dff_B_h9EIukWF0_2),.clk(gclk));
	jdff dff_B_Qh8KRF7c1_2(.din(w_dff_B_h9EIukWF0_2),.dout(w_dff_B_Qh8KRF7c1_2),.clk(gclk));
	jdff dff_B_MdxlzSYs3_2(.din(w_dff_B_Qh8KRF7c1_2),.dout(w_dff_B_MdxlzSYs3_2),.clk(gclk));
	jdff dff_B_5ocVLUiB6_2(.din(w_dff_B_MdxlzSYs3_2),.dout(w_dff_B_5ocVLUiB6_2),.clk(gclk));
	jdff dff_B_qwmLDYlS5_2(.din(w_dff_B_5ocVLUiB6_2),.dout(w_dff_B_qwmLDYlS5_2),.clk(gclk));
	jdff dff_B_K8LkMMUf4_2(.din(w_dff_B_qwmLDYlS5_2),.dout(w_dff_B_K8LkMMUf4_2),.clk(gclk));
	jdff dff_B_3QpEcBYS5_2(.din(w_dff_B_K8LkMMUf4_2),.dout(w_dff_B_3QpEcBYS5_2),.clk(gclk));
	jdff dff_B_B68IbSmN4_2(.din(w_dff_B_3QpEcBYS5_2),.dout(w_dff_B_B68IbSmN4_2),.clk(gclk));
	jdff dff_B_q2UG8rry9_2(.din(w_dff_B_B68IbSmN4_2),.dout(w_dff_B_q2UG8rry9_2),.clk(gclk));
	jdff dff_B_GWmTiUBi7_2(.din(w_dff_B_q2UG8rry9_2),.dout(w_dff_B_GWmTiUBi7_2),.clk(gclk));
	jdff dff_B_6czhGHEI7_2(.din(w_dff_B_GWmTiUBi7_2),.dout(w_dff_B_6czhGHEI7_2),.clk(gclk));
	jdff dff_B_0dWJxbfB1_2(.din(w_dff_B_6czhGHEI7_2),.dout(w_dff_B_0dWJxbfB1_2),.clk(gclk));
	jdff dff_B_Wiglwtz19_2(.din(w_dff_B_0dWJxbfB1_2),.dout(w_dff_B_Wiglwtz19_2),.clk(gclk));
	jdff dff_B_e4hHRO710_2(.din(w_dff_B_Wiglwtz19_2),.dout(w_dff_B_e4hHRO710_2),.clk(gclk));
	jdff dff_B_t7NTSo022_2(.din(w_dff_B_e4hHRO710_2),.dout(w_dff_B_t7NTSo022_2),.clk(gclk));
	jdff dff_B_gEWZXbi90_2(.din(n1636),.dout(w_dff_B_gEWZXbi90_2),.clk(gclk));
	jdff dff_B_4DM503qx1_1(.din(n1634),.dout(w_dff_B_4DM503qx1_1),.clk(gclk));
	jdff dff_B_XSj0W33P0_2(.din(n1576),.dout(w_dff_B_XSj0W33P0_2),.clk(gclk));
	jdff dff_B_mF69VJTT3_2(.din(w_dff_B_XSj0W33P0_2),.dout(w_dff_B_mF69VJTT3_2),.clk(gclk));
	jdff dff_B_ucASIHuc0_2(.din(w_dff_B_mF69VJTT3_2),.dout(w_dff_B_ucASIHuc0_2),.clk(gclk));
	jdff dff_B_Qftq9QV42_2(.din(w_dff_B_ucASIHuc0_2),.dout(w_dff_B_Qftq9QV42_2),.clk(gclk));
	jdff dff_B_et16hyLE3_2(.din(w_dff_B_Qftq9QV42_2),.dout(w_dff_B_et16hyLE3_2),.clk(gclk));
	jdff dff_B_9Nd1Zc0o6_2(.din(w_dff_B_et16hyLE3_2),.dout(w_dff_B_9Nd1Zc0o6_2),.clk(gclk));
	jdff dff_B_QzZVqoBh7_2(.din(w_dff_B_9Nd1Zc0o6_2),.dout(w_dff_B_QzZVqoBh7_2),.clk(gclk));
	jdff dff_B_IkSMX9aT1_2(.din(w_dff_B_QzZVqoBh7_2),.dout(w_dff_B_IkSMX9aT1_2),.clk(gclk));
	jdff dff_B_vQHBgyYe9_2(.din(w_dff_B_IkSMX9aT1_2),.dout(w_dff_B_vQHBgyYe9_2),.clk(gclk));
	jdff dff_B_vvAv7Okf5_2(.din(w_dff_B_vQHBgyYe9_2),.dout(w_dff_B_vvAv7Okf5_2),.clk(gclk));
	jdff dff_B_5e5HsEMC4_2(.din(w_dff_B_vvAv7Okf5_2),.dout(w_dff_B_5e5HsEMC4_2),.clk(gclk));
	jdff dff_B_pEBgNAwd1_2(.din(w_dff_B_5e5HsEMC4_2),.dout(w_dff_B_pEBgNAwd1_2),.clk(gclk));
	jdff dff_B_Vuefmv1m0_2(.din(w_dff_B_pEBgNAwd1_2),.dout(w_dff_B_Vuefmv1m0_2),.clk(gclk));
	jdff dff_B_COoAiAtz7_2(.din(w_dff_B_Vuefmv1m0_2),.dout(w_dff_B_COoAiAtz7_2),.clk(gclk));
	jdff dff_B_DnnAyAKx2_2(.din(w_dff_B_COoAiAtz7_2),.dout(w_dff_B_DnnAyAKx2_2),.clk(gclk));
	jdff dff_B_muPSitCL1_2(.din(w_dff_B_DnnAyAKx2_2),.dout(w_dff_B_muPSitCL1_2),.clk(gclk));
	jdff dff_B_muLNuAq94_2(.din(w_dff_B_muPSitCL1_2),.dout(w_dff_B_muLNuAq94_2),.clk(gclk));
	jdff dff_B_CAX2kDuR4_2(.din(w_dff_B_muLNuAq94_2),.dout(w_dff_B_CAX2kDuR4_2),.clk(gclk));
	jdff dff_B_TWbd1d8b4_2(.din(w_dff_B_CAX2kDuR4_2),.dout(w_dff_B_TWbd1d8b4_2),.clk(gclk));
	jdff dff_B_JI8RnBij7_2(.din(w_dff_B_TWbd1d8b4_2),.dout(w_dff_B_JI8RnBij7_2),.clk(gclk));
	jdff dff_B_p95ohL3o8_2(.din(w_dff_B_JI8RnBij7_2),.dout(w_dff_B_p95ohL3o8_2),.clk(gclk));
	jdff dff_B_TxH64Jd20_2(.din(w_dff_B_p95ohL3o8_2),.dout(w_dff_B_TxH64Jd20_2),.clk(gclk));
	jdff dff_B_vlsk8rsp8_2(.din(w_dff_B_TxH64Jd20_2),.dout(w_dff_B_vlsk8rsp8_2),.clk(gclk));
	jdff dff_B_HWi3T1sR2_2(.din(w_dff_B_vlsk8rsp8_2),.dout(w_dff_B_HWi3T1sR2_2),.clk(gclk));
	jdff dff_B_syxz5Bew5_2(.din(w_dff_B_HWi3T1sR2_2),.dout(w_dff_B_syxz5Bew5_2),.clk(gclk));
	jdff dff_B_ViomdNKI7_2(.din(w_dff_B_syxz5Bew5_2),.dout(w_dff_B_ViomdNKI7_2),.clk(gclk));
	jdff dff_B_B2IHkcjU0_2(.din(w_dff_B_ViomdNKI7_2),.dout(w_dff_B_B2IHkcjU0_2),.clk(gclk));
	jdff dff_B_JFXiRL2v5_2(.din(w_dff_B_B2IHkcjU0_2),.dout(w_dff_B_JFXiRL2v5_2),.clk(gclk));
	jdff dff_B_qnOSOI3J0_2(.din(w_dff_B_JFXiRL2v5_2),.dout(w_dff_B_qnOSOI3J0_2),.clk(gclk));
	jdff dff_B_o0aGfLs23_2(.din(w_dff_B_qnOSOI3J0_2),.dout(w_dff_B_o0aGfLs23_2),.clk(gclk));
	jdff dff_B_2ZGwtNOI0_2(.din(w_dff_B_o0aGfLs23_2),.dout(w_dff_B_2ZGwtNOI0_2),.clk(gclk));
	jdff dff_B_oYfWgQwj4_2(.din(w_dff_B_2ZGwtNOI0_2),.dout(w_dff_B_oYfWgQwj4_2),.clk(gclk));
	jdff dff_B_vrHRwwY64_2(.din(w_dff_B_oYfWgQwj4_2),.dout(w_dff_B_vrHRwwY64_2),.clk(gclk));
	jdff dff_B_w6MhnlCF4_2(.din(w_dff_B_vrHRwwY64_2),.dout(w_dff_B_w6MhnlCF4_2),.clk(gclk));
	jdff dff_B_dLFBpsyn4_2(.din(w_dff_B_w6MhnlCF4_2),.dout(w_dff_B_dLFBpsyn4_2),.clk(gclk));
	jdff dff_B_lOrcylcN4_2(.din(w_dff_B_dLFBpsyn4_2),.dout(w_dff_B_lOrcylcN4_2),.clk(gclk));
	jdff dff_B_NTf9Cb4h1_2(.din(w_dff_B_lOrcylcN4_2),.dout(w_dff_B_NTf9Cb4h1_2),.clk(gclk));
	jdff dff_B_1xK1Vb336_2(.din(w_dff_B_NTf9Cb4h1_2),.dout(w_dff_B_1xK1Vb336_2),.clk(gclk));
	jdff dff_B_k00PbxRh3_2(.din(w_dff_B_1xK1Vb336_2),.dout(w_dff_B_k00PbxRh3_2),.clk(gclk));
	jdff dff_B_shqddaeU0_2(.din(w_dff_B_k00PbxRh3_2),.dout(w_dff_B_shqddaeU0_2),.clk(gclk));
	jdff dff_B_PlW01fJO6_2(.din(w_dff_B_shqddaeU0_2),.dout(w_dff_B_PlW01fJO6_2),.clk(gclk));
	jdff dff_B_k6Z3dM301_2(.din(n1579),.dout(w_dff_B_k6Z3dM301_2),.clk(gclk));
	jdff dff_B_KWsj1w4I1_1(.din(n1577),.dout(w_dff_B_KWsj1w4I1_1),.clk(gclk));
	jdff dff_B_fnADqmUn2_2(.din(n1512),.dout(w_dff_B_fnADqmUn2_2),.clk(gclk));
	jdff dff_B_HtyjzvXR0_2(.din(w_dff_B_fnADqmUn2_2),.dout(w_dff_B_HtyjzvXR0_2),.clk(gclk));
	jdff dff_B_niEEAyfw3_2(.din(w_dff_B_HtyjzvXR0_2),.dout(w_dff_B_niEEAyfw3_2),.clk(gclk));
	jdff dff_B_nkqB8I3H3_2(.din(w_dff_B_niEEAyfw3_2),.dout(w_dff_B_nkqB8I3H3_2),.clk(gclk));
	jdff dff_B_MBEf3onO7_2(.din(w_dff_B_nkqB8I3H3_2),.dout(w_dff_B_MBEf3onO7_2),.clk(gclk));
	jdff dff_B_xExIR2Qf8_2(.din(w_dff_B_MBEf3onO7_2),.dout(w_dff_B_xExIR2Qf8_2),.clk(gclk));
	jdff dff_B_ZZj8lqqf6_2(.din(w_dff_B_xExIR2Qf8_2),.dout(w_dff_B_ZZj8lqqf6_2),.clk(gclk));
	jdff dff_B_wDnhVLNH7_2(.din(w_dff_B_ZZj8lqqf6_2),.dout(w_dff_B_wDnhVLNH7_2),.clk(gclk));
	jdff dff_B_N5r9Gnzo9_2(.din(w_dff_B_wDnhVLNH7_2),.dout(w_dff_B_N5r9Gnzo9_2),.clk(gclk));
	jdff dff_B_dFgESHhn5_2(.din(w_dff_B_N5r9Gnzo9_2),.dout(w_dff_B_dFgESHhn5_2),.clk(gclk));
	jdff dff_B_I5XpsT1x0_2(.din(w_dff_B_dFgESHhn5_2),.dout(w_dff_B_I5XpsT1x0_2),.clk(gclk));
	jdff dff_B_qxrLQuA97_2(.din(w_dff_B_I5XpsT1x0_2),.dout(w_dff_B_qxrLQuA97_2),.clk(gclk));
	jdff dff_B_TwS7Su2d1_2(.din(w_dff_B_qxrLQuA97_2),.dout(w_dff_B_TwS7Su2d1_2),.clk(gclk));
	jdff dff_B_TI4D2na19_2(.din(w_dff_B_TwS7Su2d1_2),.dout(w_dff_B_TI4D2na19_2),.clk(gclk));
	jdff dff_B_wdtrvRXi8_2(.din(w_dff_B_TI4D2na19_2),.dout(w_dff_B_wdtrvRXi8_2),.clk(gclk));
	jdff dff_B_GE6M4kkh9_2(.din(w_dff_B_wdtrvRXi8_2),.dout(w_dff_B_GE6M4kkh9_2),.clk(gclk));
	jdff dff_B_1v9xkd8r2_2(.din(w_dff_B_GE6M4kkh9_2),.dout(w_dff_B_1v9xkd8r2_2),.clk(gclk));
	jdff dff_B_c8p1SSMr9_2(.din(w_dff_B_1v9xkd8r2_2),.dout(w_dff_B_c8p1SSMr9_2),.clk(gclk));
	jdff dff_B_rG8uYtic6_2(.din(w_dff_B_c8p1SSMr9_2),.dout(w_dff_B_rG8uYtic6_2),.clk(gclk));
	jdff dff_B_G2qFkAGH0_2(.din(w_dff_B_rG8uYtic6_2),.dout(w_dff_B_G2qFkAGH0_2),.clk(gclk));
	jdff dff_B_BmlNWpeI1_2(.din(w_dff_B_G2qFkAGH0_2),.dout(w_dff_B_BmlNWpeI1_2),.clk(gclk));
	jdff dff_B_8s4SRJPV3_2(.din(w_dff_B_BmlNWpeI1_2),.dout(w_dff_B_8s4SRJPV3_2),.clk(gclk));
	jdff dff_B_hxYpHBWI4_2(.din(w_dff_B_8s4SRJPV3_2),.dout(w_dff_B_hxYpHBWI4_2),.clk(gclk));
	jdff dff_B_iqOqpiti7_2(.din(w_dff_B_hxYpHBWI4_2),.dout(w_dff_B_iqOqpiti7_2),.clk(gclk));
	jdff dff_B_1ap5ySk98_2(.din(w_dff_B_iqOqpiti7_2),.dout(w_dff_B_1ap5ySk98_2),.clk(gclk));
	jdff dff_B_ThBV1DCF0_2(.din(w_dff_B_1ap5ySk98_2),.dout(w_dff_B_ThBV1DCF0_2),.clk(gclk));
	jdff dff_B_7iAodSeq2_2(.din(w_dff_B_ThBV1DCF0_2),.dout(w_dff_B_7iAodSeq2_2),.clk(gclk));
	jdff dff_B_wopjOCEN2_2(.din(w_dff_B_7iAodSeq2_2),.dout(w_dff_B_wopjOCEN2_2),.clk(gclk));
	jdff dff_B_1WI3EKo63_2(.din(w_dff_B_wopjOCEN2_2),.dout(w_dff_B_1WI3EKo63_2),.clk(gclk));
	jdff dff_B_NR4hBKQh4_2(.din(w_dff_B_1WI3EKo63_2),.dout(w_dff_B_NR4hBKQh4_2),.clk(gclk));
	jdff dff_B_G5gHnXfc5_2(.din(w_dff_B_NR4hBKQh4_2),.dout(w_dff_B_G5gHnXfc5_2),.clk(gclk));
	jdff dff_B_QN5lWEbu1_2(.din(w_dff_B_G5gHnXfc5_2),.dout(w_dff_B_QN5lWEbu1_2),.clk(gclk));
	jdff dff_B_hL6rvXJP4_2(.din(w_dff_B_QN5lWEbu1_2),.dout(w_dff_B_hL6rvXJP4_2),.clk(gclk));
	jdff dff_B_Xcz8bQt79_2(.din(w_dff_B_hL6rvXJP4_2),.dout(w_dff_B_Xcz8bQt79_2),.clk(gclk));
	jdff dff_B_lrITYiHD2_2(.din(w_dff_B_Xcz8bQt79_2),.dout(w_dff_B_lrITYiHD2_2),.clk(gclk));
	jdff dff_B_BHbMM9XM6_2(.din(w_dff_B_lrITYiHD2_2),.dout(w_dff_B_BHbMM9XM6_2),.clk(gclk));
	jdff dff_B_2q0oM0jv1_2(.din(w_dff_B_BHbMM9XM6_2),.dout(w_dff_B_2q0oM0jv1_2),.clk(gclk));
	jdff dff_B_f4y5ryhm3_2(.din(n1515),.dout(w_dff_B_f4y5ryhm3_2),.clk(gclk));
	jdff dff_B_QlXDA0Gs6_1(.din(n1513),.dout(w_dff_B_QlXDA0Gs6_1),.clk(gclk));
	jdff dff_B_HFuURorS5_2(.din(n1441),.dout(w_dff_B_HFuURorS5_2),.clk(gclk));
	jdff dff_B_HYtwev9K1_2(.din(w_dff_B_HFuURorS5_2),.dout(w_dff_B_HYtwev9K1_2),.clk(gclk));
	jdff dff_B_jsr3QjnB4_2(.din(w_dff_B_HYtwev9K1_2),.dout(w_dff_B_jsr3QjnB4_2),.clk(gclk));
	jdff dff_B_KLGBzTgE6_2(.din(w_dff_B_jsr3QjnB4_2),.dout(w_dff_B_KLGBzTgE6_2),.clk(gclk));
	jdff dff_B_6ChZadHj3_2(.din(w_dff_B_KLGBzTgE6_2),.dout(w_dff_B_6ChZadHj3_2),.clk(gclk));
	jdff dff_B_UbqCyEjC9_2(.din(w_dff_B_6ChZadHj3_2),.dout(w_dff_B_UbqCyEjC9_2),.clk(gclk));
	jdff dff_B_Hhwahzwe4_2(.din(w_dff_B_UbqCyEjC9_2),.dout(w_dff_B_Hhwahzwe4_2),.clk(gclk));
	jdff dff_B_2iJvjgP80_2(.din(w_dff_B_Hhwahzwe4_2),.dout(w_dff_B_2iJvjgP80_2),.clk(gclk));
	jdff dff_B_0rAaLXo55_2(.din(w_dff_B_2iJvjgP80_2),.dout(w_dff_B_0rAaLXo55_2),.clk(gclk));
	jdff dff_B_WKRz6zFz4_2(.din(w_dff_B_0rAaLXo55_2),.dout(w_dff_B_WKRz6zFz4_2),.clk(gclk));
	jdff dff_B_mYj8hEJG2_2(.din(w_dff_B_WKRz6zFz4_2),.dout(w_dff_B_mYj8hEJG2_2),.clk(gclk));
	jdff dff_B_2tDofd421_2(.din(w_dff_B_mYj8hEJG2_2),.dout(w_dff_B_2tDofd421_2),.clk(gclk));
	jdff dff_B_BrDCQca44_2(.din(w_dff_B_2tDofd421_2),.dout(w_dff_B_BrDCQca44_2),.clk(gclk));
	jdff dff_B_ovWFeDIW3_2(.din(w_dff_B_BrDCQca44_2),.dout(w_dff_B_ovWFeDIW3_2),.clk(gclk));
	jdff dff_B_UFvFRXVG7_2(.din(w_dff_B_ovWFeDIW3_2),.dout(w_dff_B_UFvFRXVG7_2),.clk(gclk));
	jdff dff_B_dWjQTx6d2_2(.din(w_dff_B_UFvFRXVG7_2),.dout(w_dff_B_dWjQTx6d2_2),.clk(gclk));
	jdff dff_B_Z1pQawyx2_2(.din(w_dff_B_dWjQTx6d2_2),.dout(w_dff_B_Z1pQawyx2_2),.clk(gclk));
	jdff dff_B_2Mws1gYY1_2(.din(w_dff_B_Z1pQawyx2_2),.dout(w_dff_B_2Mws1gYY1_2),.clk(gclk));
	jdff dff_B_tviATJVO9_2(.din(w_dff_B_2Mws1gYY1_2),.dout(w_dff_B_tviATJVO9_2),.clk(gclk));
	jdff dff_B_GTeB3NYr8_2(.din(w_dff_B_tviATJVO9_2),.dout(w_dff_B_GTeB3NYr8_2),.clk(gclk));
	jdff dff_B_Y6j6lNRV8_2(.din(w_dff_B_GTeB3NYr8_2),.dout(w_dff_B_Y6j6lNRV8_2),.clk(gclk));
	jdff dff_B_unFGG66d8_2(.din(w_dff_B_Y6j6lNRV8_2),.dout(w_dff_B_unFGG66d8_2),.clk(gclk));
	jdff dff_B_7aIpXPD49_2(.din(w_dff_B_unFGG66d8_2),.dout(w_dff_B_7aIpXPD49_2),.clk(gclk));
	jdff dff_B_V2ISwFEN5_2(.din(w_dff_B_7aIpXPD49_2),.dout(w_dff_B_V2ISwFEN5_2),.clk(gclk));
	jdff dff_B_LJw5olb82_2(.din(w_dff_B_V2ISwFEN5_2),.dout(w_dff_B_LJw5olb82_2),.clk(gclk));
	jdff dff_B_Fx76HhxW5_2(.din(w_dff_B_LJw5olb82_2),.dout(w_dff_B_Fx76HhxW5_2),.clk(gclk));
	jdff dff_B_0u5xo9Bq9_2(.din(w_dff_B_Fx76HhxW5_2),.dout(w_dff_B_0u5xo9Bq9_2),.clk(gclk));
	jdff dff_B_GmD0ky7j3_2(.din(w_dff_B_0u5xo9Bq9_2),.dout(w_dff_B_GmD0ky7j3_2),.clk(gclk));
	jdff dff_B_n9K19JA90_2(.din(w_dff_B_GmD0ky7j3_2),.dout(w_dff_B_n9K19JA90_2),.clk(gclk));
	jdff dff_B_fMOdFGYu5_2(.din(w_dff_B_n9K19JA90_2),.dout(w_dff_B_fMOdFGYu5_2),.clk(gclk));
	jdff dff_B_y2k1Dz5Y5_2(.din(w_dff_B_fMOdFGYu5_2),.dout(w_dff_B_y2k1Dz5Y5_2),.clk(gclk));
	jdff dff_B_ogX3M0e88_2(.din(w_dff_B_y2k1Dz5Y5_2),.dout(w_dff_B_ogX3M0e88_2),.clk(gclk));
	jdff dff_B_NIiP5MnK3_2(.din(w_dff_B_ogX3M0e88_2),.dout(w_dff_B_NIiP5MnK3_2),.clk(gclk));
	jdff dff_B_0Ke26RMA9_1(.din(n1442),.dout(w_dff_B_0Ke26RMA9_1),.clk(gclk));
	jdff dff_B_zdur0rHx6_2(.din(n1363),.dout(w_dff_B_zdur0rHx6_2),.clk(gclk));
	jdff dff_B_NHoRZHjM0_2(.din(w_dff_B_zdur0rHx6_2),.dout(w_dff_B_NHoRZHjM0_2),.clk(gclk));
	jdff dff_B_8SYQqcns8_2(.din(w_dff_B_NHoRZHjM0_2),.dout(w_dff_B_8SYQqcns8_2),.clk(gclk));
	jdff dff_B_YBcxg5414_2(.din(w_dff_B_8SYQqcns8_2),.dout(w_dff_B_YBcxg5414_2),.clk(gclk));
	jdff dff_B_erQ4fIHP6_2(.din(w_dff_B_YBcxg5414_2),.dout(w_dff_B_erQ4fIHP6_2),.clk(gclk));
	jdff dff_B_4PuvGxbi5_2(.din(w_dff_B_erQ4fIHP6_2),.dout(w_dff_B_4PuvGxbi5_2),.clk(gclk));
	jdff dff_B_HMFb1ltr6_2(.din(w_dff_B_4PuvGxbi5_2),.dout(w_dff_B_HMFb1ltr6_2),.clk(gclk));
	jdff dff_B_Ife0iku81_2(.din(w_dff_B_HMFb1ltr6_2),.dout(w_dff_B_Ife0iku81_2),.clk(gclk));
	jdff dff_B_f8cjXL9Z2_2(.din(w_dff_B_Ife0iku81_2),.dout(w_dff_B_f8cjXL9Z2_2),.clk(gclk));
	jdff dff_B_UiOIbgrz5_2(.din(w_dff_B_f8cjXL9Z2_2),.dout(w_dff_B_UiOIbgrz5_2),.clk(gclk));
	jdff dff_B_7jUvcbn46_2(.din(w_dff_B_UiOIbgrz5_2),.dout(w_dff_B_7jUvcbn46_2),.clk(gclk));
	jdff dff_B_EVeQGmWW3_2(.din(w_dff_B_7jUvcbn46_2),.dout(w_dff_B_EVeQGmWW3_2),.clk(gclk));
	jdff dff_B_H9Ffuray3_2(.din(w_dff_B_EVeQGmWW3_2),.dout(w_dff_B_H9Ffuray3_2),.clk(gclk));
	jdff dff_B_3akg4uhZ2_2(.din(w_dff_B_H9Ffuray3_2),.dout(w_dff_B_3akg4uhZ2_2),.clk(gclk));
	jdff dff_B_qlAL7DbF5_2(.din(w_dff_B_3akg4uhZ2_2),.dout(w_dff_B_qlAL7DbF5_2),.clk(gclk));
	jdff dff_B_rcyTbpPx5_2(.din(w_dff_B_qlAL7DbF5_2),.dout(w_dff_B_rcyTbpPx5_2),.clk(gclk));
	jdff dff_B_Egp1LORW2_2(.din(w_dff_B_rcyTbpPx5_2),.dout(w_dff_B_Egp1LORW2_2),.clk(gclk));
	jdff dff_B_W59M4nOI8_2(.din(w_dff_B_Egp1LORW2_2),.dout(w_dff_B_W59M4nOI8_2),.clk(gclk));
	jdff dff_B_bxryLyCT7_2(.din(w_dff_B_W59M4nOI8_2),.dout(w_dff_B_bxryLyCT7_2),.clk(gclk));
	jdff dff_B_7WUGfm5W9_2(.din(w_dff_B_bxryLyCT7_2),.dout(w_dff_B_7WUGfm5W9_2),.clk(gclk));
	jdff dff_B_4Lb1V7ce6_2(.din(w_dff_B_7WUGfm5W9_2),.dout(w_dff_B_4Lb1V7ce6_2),.clk(gclk));
	jdff dff_B_VoDIUlxA7_2(.din(w_dff_B_4Lb1V7ce6_2),.dout(w_dff_B_VoDIUlxA7_2),.clk(gclk));
	jdff dff_B_XTgZh5318_2(.din(w_dff_B_VoDIUlxA7_2),.dout(w_dff_B_XTgZh5318_2),.clk(gclk));
	jdff dff_B_CL2iF2yL3_2(.din(w_dff_B_XTgZh5318_2),.dout(w_dff_B_CL2iF2yL3_2),.clk(gclk));
	jdff dff_B_k9owATDD3_2(.din(w_dff_B_CL2iF2yL3_2),.dout(w_dff_B_k9owATDD3_2),.clk(gclk));
	jdff dff_B_iyU4cppo5_2(.din(w_dff_B_k9owATDD3_2),.dout(w_dff_B_iyU4cppo5_2),.clk(gclk));
	jdff dff_B_MsQzurds4_2(.din(w_dff_B_iyU4cppo5_2),.dout(w_dff_B_MsQzurds4_2),.clk(gclk));
	jdff dff_B_TTTi2UUd8_2(.din(w_dff_B_MsQzurds4_2),.dout(w_dff_B_TTTi2UUd8_2),.clk(gclk));
	jdff dff_B_WJEV09jc6_2(.din(w_dff_B_TTTi2UUd8_2),.dout(w_dff_B_WJEV09jc6_2),.clk(gclk));
	jdff dff_B_iqpIQTzU2_2(.din(w_dff_B_WJEV09jc6_2),.dout(w_dff_B_iqpIQTzU2_2),.clk(gclk));
	jdff dff_B_2gb9Bxer1_2(.din(n1395),.dout(w_dff_B_2gb9Bxer1_2),.clk(gclk));
	jdff dff_B_jkB5FMPY5_1(.din(n1364),.dout(w_dff_B_jkB5FMPY5_1),.clk(gclk));
	jdff dff_B_EHNiVPGa5_2(.din(n1278),.dout(w_dff_B_EHNiVPGa5_2),.clk(gclk));
	jdff dff_B_R53KKUYP0_2(.din(w_dff_B_EHNiVPGa5_2),.dout(w_dff_B_R53KKUYP0_2),.clk(gclk));
	jdff dff_B_cZjVBzQE5_2(.din(w_dff_B_R53KKUYP0_2),.dout(w_dff_B_cZjVBzQE5_2),.clk(gclk));
	jdff dff_B_4j4JNBkS9_2(.din(w_dff_B_cZjVBzQE5_2),.dout(w_dff_B_4j4JNBkS9_2),.clk(gclk));
	jdff dff_B_qudDM4mX8_2(.din(w_dff_B_4j4JNBkS9_2),.dout(w_dff_B_qudDM4mX8_2),.clk(gclk));
	jdff dff_B_I2hQy2mV6_2(.din(w_dff_B_qudDM4mX8_2),.dout(w_dff_B_I2hQy2mV6_2),.clk(gclk));
	jdff dff_B_GUVxetKd4_2(.din(w_dff_B_I2hQy2mV6_2),.dout(w_dff_B_GUVxetKd4_2),.clk(gclk));
	jdff dff_B_WlH3N3xI3_2(.din(w_dff_B_GUVxetKd4_2),.dout(w_dff_B_WlH3N3xI3_2),.clk(gclk));
	jdff dff_B_qaD0liny8_2(.din(w_dff_B_WlH3N3xI3_2),.dout(w_dff_B_qaD0liny8_2),.clk(gclk));
	jdff dff_B_pskPLXQP5_2(.din(w_dff_B_qaD0liny8_2),.dout(w_dff_B_pskPLXQP5_2),.clk(gclk));
	jdff dff_B_RY5mHMTT7_2(.din(w_dff_B_pskPLXQP5_2),.dout(w_dff_B_RY5mHMTT7_2),.clk(gclk));
	jdff dff_B_w31ARI7p5_2(.din(w_dff_B_RY5mHMTT7_2),.dout(w_dff_B_w31ARI7p5_2),.clk(gclk));
	jdff dff_B_q0iaNeqA5_2(.din(w_dff_B_w31ARI7p5_2),.dout(w_dff_B_q0iaNeqA5_2),.clk(gclk));
	jdff dff_B_Ktf7kmeC2_2(.din(w_dff_B_q0iaNeqA5_2),.dout(w_dff_B_Ktf7kmeC2_2),.clk(gclk));
	jdff dff_B_DQnPTe6U1_2(.din(w_dff_B_Ktf7kmeC2_2),.dout(w_dff_B_DQnPTe6U1_2),.clk(gclk));
	jdff dff_B_s3baH0L16_2(.din(w_dff_B_DQnPTe6U1_2),.dout(w_dff_B_s3baH0L16_2),.clk(gclk));
	jdff dff_B_smTXGo765_2(.din(w_dff_B_s3baH0L16_2),.dout(w_dff_B_smTXGo765_2),.clk(gclk));
	jdff dff_B_wqyk9ScC3_2(.din(w_dff_B_smTXGo765_2),.dout(w_dff_B_wqyk9ScC3_2),.clk(gclk));
	jdff dff_B_MOC4qZHb7_2(.din(w_dff_B_wqyk9ScC3_2),.dout(w_dff_B_MOC4qZHb7_2),.clk(gclk));
	jdff dff_B_ypz8S9Q79_2(.din(w_dff_B_MOC4qZHb7_2),.dout(w_dff_B_ypz8S9Q79_2),.clk(gclk));
	jdff dff_B_NMepsmpw3_2(.din(w_dff_B_ypz8S9Q79_2),.dout(w_dff_B_NMepsmpw3_2),.clk(gclk));
	jdff dff_B_mbJAJiPN0_2(.din(w_dff_B_NMepsmpw3_2),.dout(w_dff_B_mbJAJiPN0_2),.clk(gclk));
	jdff dff_B_yLgDWa1g2_2(.din(w_dff_B_mbJAJiPN0_2),.dout(w_dff_B_yLgDWa1g2_2),.clk(gclk));
	jdff dff_B_DO6sKrzx2_2(.din(w_dff_B_yLgDWa1g2_2),.dout(w_dff_B_DO6sKrzx2_2),.clk(gclk));
	jdff dff_B_SnAK9J960_2(.din(w_dff_B_DO6sKrzx2_2),.dout(w_dff_B_SnAK9J960_2),.clk(gclk));
	jdff dff_B_EeLLnJ7g4_2(.din(w_dff_B_SnAK9J960_2),.dout(w_dff_B_EeLLnJ7g4_2),.clk(gclk));
	jdff dff_B_1Klk0tMV1_2(.din(w_dff_B_EeLLnJ7g4_2),.dout(w_dff_B_1Klk0tMV1_2),.clk(gclk));
	jdff dff_B_OyczPD237_2(.din(n1310),.dout(w_dff_B_OyczPD237_2),.clk(gclk));
	jdff dff_B_IZsyeWf28_1(.din(n1279),.dout(w_dff_B_IZsyeWf28_1),.clk(gclk));
	jdff dff_B_L1gaHzF19_2(.din(n1188),.dout(w_dff_B_L1gaHzF19_2),.clk(gclk));
	jdff dff_B_cihPYqz81_2(.din(w_dff_B_L1gaHzF19_2),.dout(w_dff_B_cihPYqz81_2),.clk(gclk));
	jdff dff_B_GbGbOR9e9_2(.din(w_dff_B_cihPYqz81_2),.dout(w_dff_B_GbGbOR9e9_2),.clk(gclk));
	jdff dff_B_zOOFACYH8_2(.din(w_dff_B_GbGbOR9e9_2),.dout(w_dff_B_zOOFACYH8_2),.clk(gclk));
	jdff dff_B_NrA7s80c8_2(.din(w_dff_B_zOOFACYH8_2),.dout(w_dff_B_NrA7s80c8_2),.clk(gclk));
	jdff dff_B_HsfuJafL4_2(.din(w_dff_B_NrA7s80c8_2),.dout(w_dff_B_HsfuJafL4_2),.clk(gclk));
	jdff dff_B_z8Spxi6f9_2(.din(w_dff_B_HsfuJafL4_2),.dout(w_dff_B_z8Spxi6f9_2),.clk(gclk));
	jdff dff_B_TMGb5HZq1_2(.din(w_dff_B_z8Spxi6f9_2),.dout(w_dff_B_TMGb5HZq1_2),.clk(gclk));
	jdff dff_B_icSf5HTl1_2(.din(w_dff_B_TMGb5HZq1_2),.dout(w_dff_B_icSf5HTl1_2),.clk(gclk));
	jdff dff_B_EAbTJmvu8_2(.din(w_dff_B_icSf5HTl1_2),.dout(w_dff_B_EAbTJmvu8_2),.clk(gclk));
	jdff dff_B_MqnxQ0SH0_2(.din(w_dff_B_EAbTJmvu8_2),.dout(w_dff_B_MqnxQ0SH0_2),.clk(gclk));
	jdff dff_B_TTRDu9L52_2(.din(w_dff_B_MqnxQ0SH0_2),.dout(w_dff_B_TTRDu9L52_2),.clk(gclk));
	jdff dff_B_UTsSfrOG5_2(.din(w_dff_B_TTRDu9L52_2),.dout(w_dff_B_UTsSfrOG5_2),.clk(gclk));
	jdff dff_B_YY5hh0fQ9_2(.din(w_dff_B_UTsSfrOG5_2),.dout(w_dff_B_YY5hh0fQ9_2),.clk(gclk));
	jdff dff_B_DhV318ib4_2(.din(w_dff_B_YY5hh0fQ9_2),.dout(w_dff_B_DhV318ib4_2),.clk(gclk));
	jdff dff_B_Lf99Nr2G0_2(.din(w_dff_B_DhV318ib4_2),.dout(w_dff_B_Lf99Nr2G0_2),.clk(gclk));
	jdff dff_B_GMR7TjrY2_2(.din(w_dff_B_Lf99Nr2G0_2),.dout(w_dff_B_GMR7TjrY2_2),.clk(gclk));
	jdff dff_B_JLZtvhgW5_2(.din(w_dff_B_GMR7TjrY2_2),.dout(w_dff_B_JLZtvhgW5_2),.clk(gclk));
	jdff dff_B_ih9TGE8T8_2(.din(w_dff_B_JLZtvhgW5_2),.dout(w_dff_B_ih9TGE8T8_2),.clk(gclk));
	jdff dff_B_2WOqcq8D2_2(.din(w_dff_B_ih9TGE8T8_2),.dout(w_dff_B_2WOqcq8D2_2),.clk(gclk));
	jdff dff_B_NxtaKpLL8_2(.din(w_dff_B_2WOqcq8D2_2),.dout(w_dff_B_NxtaKpLL8_2),.clk(gclk));
	jdff dff_B_2FGWKC1H9_2(.din(w_dff_B_NxtaKpLL8_2),.dout(w_dff_B_2FGWKC1H9_2),.clk(gclk));
	jdff dff_B_uomZ3BfG8_2(.din(w_dff_B_2FGWKC1H9_2),.dout(w_dff_B_uomZ3BfG8_2),.clk(gclk));
	jdff dff_B_vuesWQg10_2(.din(w_dff_B_uomZ3BfG8_2),.dout(w_dff_B_vuesWQg10_2),.clk(gclk));
	jdff dff_B_0ln7i3yv3_2(.din(n1219),.dout(w_dff_B_0ln7i3yv3_2),.clk(gclk));
	jdff dff_B_teh9vl1E7_1(.din(n1189),.dout(w_dff_B_teh9vl1E7_1),.clk(gclk));
	jdff dff_B_52OESfC01_2(.din(n1084),.dout(w_dff_B_52OESfC01_2),.clk(gclk));
	jdff dff_B_nySWuDaB3_2(.din(w_dff_B_52OESfC01_2),.dout(w_dff_B_nySWuDaB3_2),.clk(gclk));
	jdff dff_B_0j5IJlxb1_2(.din(w_dff_B_nySWuDaB3_2),.dout(w_dff_B_0j5IJlxb1_2),.clk(gclk));
	jdff dff_B_xUnWSZUa1_2(.din(w_dff_B_0j5IJlxb1_2),.dout(w_dff_B_xUnWSZUa1_2),.clk(gclk));
	jdff dff_B_q6Jh4Fqk1_2(.din(w_dff_B_xUnWSZUa1_2),.dout(w_dff_B_q6Jh4Fqk1_2),.clk(gclk));
	jdff dff_B_VqFUs14A8_2(.din(w_dff_B_q6Jh4Fqk1_2),.dout(w_dff_B_VqFUs14A8_2),.clk(gclk));
	jdff dff_B_PEclydIw9_2(.din(w_dff_B_VqFUs14A8_2),.dout(w_dff_B_PEclydIw9_2),.clk(gclk));
	jdff dff_B_dwJuQe8d3_2(.din(w_dff_B_PEclydIw9_2),.dout(w_dff_B_dwJuQe8d3_2),.clk(gclk));
	jdff dff_B_bEUvZqBd9_2(.din(w_dff_B_dwJuQe8d3_2),.dout(w_dff_B_bEUvZqBd9_2),.clk(gclk));
	jdff dff_B_kn7fbtFZ0_2(.din(w_dff_B_bEUvZqBd9_2),.dout(w_dff_B_kn7fbtFZ0_2),.clk(gclk));
	jdff dff_B_LARXZbmT2_2(.din(w_dff_B_kn7fbtFZ0_2),.dout(w_dff_B_LARXZbmT2_2),.clk(gclk));
	jdff dff_B_6HOxNdgJ9_2(.din(w_dff_B_LARXZbmT2_2),.dout(w_dff_B_6HOxNdgJ9_2),.clk(gclk));
	jdff dff_B_aX6E68Rs5_2(.din(w_dff_B_6HOxNdgJ9_2),.dout(w_dff_B_aX6E68Rs5_2),.clk(gclk));
	jdff dff_B_IfY7yqZW1_2(.din(w_dff_B_aX6E68Rs5_2),.dout(w_dff_B_IfY7yqZW1_2),.clk(gclk));
	jdff dff_B_qxKB7DB39_2(.din(w_dff_B_IfY7yqZW1_2),.dout(w_dff_B_qxKB7DB39_2),.clk(gclk));
	jdff dff_B_KBa7162e0_2(.din(w_dff_B_qxKB7DB39_2),.dout(w_dff_B_KBa7162e0_2),.clk(gclk));
	jdff dff_B_KHTrgNUI6_2(.din(w_dff_B_KBa7162e0_2),.dout(w_dff_B_KHTrgNUI6_2),.clk(gclk));
	jdff dff_B_iNU01zlk3_2(.din(w_dff_B_KHTrgNUI6_2),.dout(w_dff_B_iNU01zlk3_2),.clk(gclk));
	jdff dff_B_Y66iCzaW2_2(.din(w_dff_B_iNU01zlk3_2),.dout(w_dff_B_Y66iCzaW2_2),.clk(gclk));
	jdff dff_B_FIAq9V0Q4_2(.din(w_dff_B_Y66iCzaW2_2),.dout(w_dff_B_FIAq9V0Q4_2),.clk(gclk));
	jdff dff_B_F7lIEWSj0_2(.din(w_dff_B_FIAq9V0Q4_2),.dout(w_dff_B_F7lIEWSj0_2),.clk(gclk));
	jdff dff_B_HKVoNoEe3_2(.din(n1121),.dout(w_dff_B_HKVoNoEe3_2),.clk(gclk));
	jdff dff_B_g9P1r5ym0_1(.din(n1085),.dout(w_dff_B_g9P1r5ym0_1),.clk(gclk));
	jdff dff_B_xiWu0dwT2_2(.din(n986),.dout(w_dff_B_xiWu0dwT2_2),.clk(gclk));
	jdff dff_B_YHrjbzBw9_2(.din(w_dff_B_xiWu0dwT2_2),.dout(w_dff_B_YHrjbzBw9_2),.clk(gclk));
	jdff dff_B_LEWog6le3_2(.din(w_dff_B_YHrjbzBw9_2),.dout(w_dff_B_LEWog6le3_2),.clk(gclk));
	jdff dff_B_gx8vGpJf7_2(.din(w_dff_B_LEWog6le3_2),.dout(w_dff_B_gx8vGpJf7_2),.clk(gclk));
	jdff dff_B_iXjk25ko9_2(.din(w_dff_B_gx8vGpJf7_2),.dout(w_dff_B_iXjk25ko9_2),.clk(gclk));
	jdff dff_B_QmnEWcnm7_2(.din(w_dff_B_iXjk25ko9_2),.dout(w_dff_B_QmnEWcnm7_2),.clk(gclk));
	jdff dff_B_Tk30aquB3_2(.din(w_dff_B_QmnEWcnm7_2),.dout(w_dff_B_Tk30aquB3_2),.clk(gclk));
	jdff dff_B_XUzeh79p2_2(.din(w_dff_B_Tk30aquB3_2),.dout(w_dff_B_XUzeh79p2_2),.clk(gclk));
	jdff dff_B_9RsS1pdi9_2(.din(w_dff_B_XUzeh79p2_2),.dout(w_dff_B_9RsS1pdi9_2),.clk(gclk));
	jdff dff_B_PvucHwYW2_2(.din(w_dff_B_9RsS1pdi9_2),.dout(w_dff_B_PvucHwYW2_2),.clk(gclk));
	jdff dff_B_aHsH2MyB5_2(.din(w_dff_B_PvucHwYW2_2),.dout(w_dff_B_aHsH2MyB5_2),.clk(gclk));
	jdff dff_B_dlJ8ddlK4_2(.din(w_dff_B_aHsH2MyB5_2),.dout(w_dff_B_dlJ8ddlK4_2),.clk(gclk));
	jdff dff_B_xtYAbrtG5_2(.din(w_dff_B_dlJ8ddlK4_2),.dout(w_dff_B_xtYAbrtG5_2),.clk(gclk));
	jdff dff_B_ic7GWx239_2(.din(w_dff_B_xtYAbrtG5_2),.dout(w_dff_B_ic7GWx239_2),.clk(gclk));
	jdff dff_B_ezXa3Q176_2(.din(w_dff_B_ic7GWx239_2),.dout(w_dff_B_ezXa3Q176_2),.clk(gclk));
	jdff dff_B_M7KNXDcu3_2(.din(w_dff_B_ezXa3Q176_2),.dout(w_dff_B_M7KNXDcu3_2),.clk(gclk));
	jdff dff_B_E60SA92c5_2(.din(w_dff_B_M7KNXDcu3_2),.dout(w_dff_B_E60SA92c5_2),.clk(gclk));
	jdff dff_B_A61RqbDr9_2(.din(w_dff_B_E60SA92c5_2),.dout(w_dff_B_A61RqbDr9_2),.clk(gclk));
	jdff dff_B_RcsfpYi26_2(.din(n1016),.dout(w_dff_B_RcsfpYi26_2),.clk(gclk));
	jdff dff_B_nYni0s4q4_1(.din(n987),.dout(w_dff_B_nYni0s4q4_1),.clk(gclk));
	jdff dff_B_16wA4Tok1_2(.din(n881),.dout(w_dff_B_16wA4Tok1_2),.clk(gclk));
	jdff dff_B_HcoFhwj94_2(.din(w_dff_B_16wA4Tok1_2),.dout(w_dff_B_HcoFhwj94_2),.clk(gclk));
	jdff dff_B_ssb5h6nL8_2(.din(w_dff_B_HcoFhwj94_2),.dout(w_dff_B_ssb5h6nL8_2),.clk(gclk));
	jdff dff_B_WhAQoRf68_2(.din(w_dff_B_ssb5h6nL8_2),.dout(w_dff_B_WhAQoRf68_2),.clk(gclk));
	jdff dff_B_1W6cgkrg1_2(.din(w_dff_B_WhAQoRf68_2),.dout(w_dff_B_1W6cgkrg1_2),.clk(gclk));
	jdff dff_B_qcw6OwS11_2(.din(w_dff_B_1W6cgkrg1_2),.dout(w_dff_B_qcw6OwS11_2),.clk(gclk));
	jdff dff_B_eBYhpD1m0_2(.din(w_dff_B_qcw6OwS11_2),.dout(w_dff_B_eBYhpD1m0_2),.clk(gclk));
	jdff dff_B_5Y0gQePj7_2(.din(w_dff_B_eBYhpD1m0_2),.dout(w_dff_B_5Y0gQePj7_2),.clk(gclk));
	jdff dff_B_gqcx2evk1_2(.din(w_dff_B_5Y0gQePj7_2),.dout(w_dff_B_gqcx2evk1_2),.clk(gclk));
	jdff dff_B_rmOU3GDN6_2(.din(w_dff_B_gqcx2evk1_2),.dout(w_dff_B_rmOU3GDN6_2),.clk(gclk));
	jdff dff_B_z7giTpya6_2(.din(w_dff_B_rmOU3GDN6_2),.dout(w_dff_B_z7giTpya6_2),.clk(gclk));
	jdff dff_B_Z3acxj7O5_2(.din(w_dff_B_z7giTpya6_2),.dout(w_dff_B_Z3acxj7O5_2),.clk(gclk));
	jdff dff_B_SG9yeJir4_2(.din(w_dff_B_Z3acxj7O5_2),.dout(w_dff_B_SG9yeJir4_2),.clk(gclk));
	jdff dff_B_f9xz1iH55_2(.din(w_dff_B_SG9yeJir4_2),.dout(w_dff_B_f9xz1iH55_2),.clk(gclk));
	jdff dff_B_JmAnH8nQ3_2(.din(w_dff_B_f9xz1iH55_2),.dout(w_dff_B_JmAnH8nQ3_2),.clk(gclk));
	jdff dff_B_Lcdxw4Xr7_2(.din(n911),.dout(w_dff_B_Lcdxw4Xr7_2),.clk(gclk));
	jdff dff_B_6TftSVYF7_1(.din(n882),.dout(w_dff_B_6TftSVYF7_1),.clk(gclk));
	jdff dff_B_fOZFgnN18_2(.din(n782),.dout(w_dff_B_fOZFgnN18_2),.clk(gclk));
	jdff dff_B_J6dWZeOp2_2(.din(w_dff_B_fOZFgnN18_2),.dout(w_dff_B_J6dWZeOp2_2),.clk(gclk));
	jdff dff_B_NEtTj2Mq9_2(.din(w_dff_B_J6dWZeOp2_2),.dout(w_dff_B_NEtTj2Mq9_2),.clk(gclk));
	jdff dff_B_S3EBGOoQ6_2(.din(w_dff_B_NEtTj2Mq9_2),.dout(w_dff_B_S3EBGOoQ6_2),.clk(gclk));
	jdff dff_B_y1VeWTxt8_2(.din(w_dff_B_S3EBGOoQ6_2),.dout(w_dff_B_y1VeWTxt8_2),.clk(gclk));
	jdff dff_B_jOoHe2UU8_2(.din(w_dff_B_y1VeWTxt8_2),.dout(w_dff_B_jOoHe2UU8_2),.clk(gclk));
	jdff dff_B_gsI5fYDQ3_2(.din(w_dff_B_jOoHe2UU8_2),.dout(w_dff_B_gsI5fYDQ3_2),.clk(gclk));
	jdff dff_B_NBf5rh7b4_2(.din(w_dff_B_gsI5fYDQ3_2),.dout(w_dff_B_NBf5rh7b4_2),.clk(gclk));
	jdff dff_B_OydbojVv2_2(.din(w_dff_B_NBf5rh7b4_2),.dout(w_dff_B_OydbojVv2_2),.clk(gclk));
	jdff dff_B_XepdfhXy6_2(.din(w_dff_B_OydbojVv2_2),.dout(w_dff_B_XepdfhXy6_2),.clk(gclk));
	jdff dff_B_r2F1US2v5_2(.din(w_dff_B_XepdfhXy6_2),.dout(w_dff_B_r2F1US2v5_2),.clk(gclk));
	jdff dff_B_Fx7TQE1T8_2(.din(w_dff_B_r2F1US2v5_2),.dout(w_dff_B_Fx7TQE1T8_2),.clk(gclk));
	jdff dff_B_tWtJj8lm3_2(.din(n805),.dout(w_dff_B_tWtJj8lm3_2),.clk(gclk));
	jdff dff_B_R12el6iH1_1(.din(n783),.dout(w_dff_B_R12el6iH1_1),.clk(gclk));
	jdff dff_B_tdkRVyET1_2(.din(n689),.dout(w_dff_B_tdkRVyET1_2),.clk(gclk));
	jdff dff_B_Dw7Hi8SV3_2(.din(w_dff_B_tdkRVyET1_2),.dout(w_dff_B_Dw7Hi8SV3_2),.clk(gclk));
	jdff dff_B_frbER5xA9_2(.din(w_dff_B_Dw7Hi8SV3_2),.dout(w_dff_B_frbER5xA9_2),.clk(gclk));
	jdff dff_B_rmnmQTaV7_2(.din(w_dff_B_frbER5xA9_2),.dout(w_dff_B_rmnmQTaV7_2),.clk(gclk));
	jdff dff_B_qIGRpHMu2_2(.din(w_dff_B_rmnmQTaV7_2),.dout(w_dff_B_qIGRpHMu2_2),.clk(gclk));
	jdff dff_B_3QBsWR8H1_2(.din(w_dff_B_qIGRpHMu2_2),.dout(w_dff_B_3QBsWR8H1_2),.clk(gclk));
	jdff dff_B_zqHIAowd4_2(.din(w_dff_B_3QBsWR8H1_2),.dout(w_dff_B_zqHIAowd4_2),.clk(gclk));
	jdff dff_B_y05Obsgc0_2(.din(w_dff_B_zqHIAowd4_2),.dout(w_dff_B_y05Obsgc0_2),.clk(gclk));
	jdff dff_B_PumEGzma6_2(.din(w_dff_B_y05Obsgc0_2),.dout(w_dff_B_PumEGzma6_2),.clk(gclk));
	jdff dff_B_yd2VpjQb7_2(.din(n705),.dout(w_dff_B_yd2VpjQb7_2),.clk(gclk));
	jdff dff_B_GTmP2KeA8_2(.din(w_dff_B_yd2VpjQb7_2),.dout(w_dff_B_GTmP2KeA8_2),.clk(gclk));
	jdff dff_B_Y7u0ICTY3_1(.din(n690),.dout(w_dff_B_Y7u0ICTY3_1),.clk(gclk));
	jdff dff_B_vMOoao6P2_1(.din(w_dff_B_Y7u0ICTY3_1),.dout(w_dff_B_vMOoao6P2_1),.clk(gclk));
	jdff dff_B_6wM3bMd49_1(.din(w_dff_B_vMOoao6P2_1),.dout(w_dff_B_6wM3bMd49_1),.clk(gclk));
	jdff dff_B_GKLQP4Ta8_1(.din(w_dff_B_6wM3bMd49_1),.dout(w_dff_B_GKLQP4Ta8_1),.clk(gclk));
	jdff dff_B_pEl37SFF6_1(.din(w_dff_B_GKLQP4Ta8_1),.dout(w_dff_B_pEl37SFF6_1),.clk(gclk));
	jdff dff_B_w4rI4dlB8_1(.din(w_dff_B_pEl37SFF6_1),.dout(w_dff_B_w4rI4dlB8_1),.clk(gclk));
	jdff dff_B_uvHwSihO4_0(.din(n612),.dout(w_dff_B_uvHwSihO4_0),.clk(gclk));
	jdff dff_B_yeWItqQb4_0(.din(w_dff_B_uvHwSihO4_0),.dout(w_dff_B_yeWItqQb4_0),.clk(gclk));
	jdff dff_A_sMSki8O07_0(.dout(w_n611_0[0]),.din(w_dff_A_sMSki8O07_0),.clk(gclk));
	jdff dff_A_mV1ETtr76_0(.dout(w_dff_A_sMSki8O07_0),.din(w_dff_A_mV1ETtr76_0),.clk(gclk));
	jdff dff_A_DwgwG6gr1_0(.dout(w_dff_A_mV1ETtr76_0),.din(w_dff_A_DwgwG6gr1_0),.clk(gclk));
	jdff dff_B_wtlWOni45_1(.din(n605),.dout(w_dff_B_wtlWOni45_1),.clk(gclk));
	jdff dff_A_8UhmKZc75_0(.dout(w_n523_0[0]),.din(w_dff_A_8UhmKZc75_0),.clk(gclk));
	jdff dff_A_TaYnXwFq7_1(.dout(w_n523_0[1]),.din(w_dff_A_TaYnXwFq7_1),.clk(gclk));
	jdff dff_A_NfLo46A38_1(.dout(w_dff_A_TaYnXwFq7_1),.din(w_dff_A_NfLo46A38_1),.clk(gclk));
	jdff dff_A_lD78zEp75_1(.dout(w_n603_0[1]),.din(w_dff_A_lD78zEp75_1),.clk(gclk));
	jdff dff_A_iRN75Ff71_1(.dout(w_dff_A_lD78zEp75_1),.din(w_dff_A_iRN75Ff71_1),.clk(gclk));
	jdff dff_A_U1GsVckW9_1(.dout(w_dff_A_iRN75Ff71_1),.din(w_dff_A_U1GsVckW9_1),.clk(gclk));
	jdff dff_A_kf5tlb256_1(.dout(w_dff_A_U1GsVckW9_1),.din(w_dff_A_kf5tlb256_1),.clk(gclk));
	jdff dff_A_9RwiuLbM9_1(.dout(w_dff_A_kf5tlb256_1),.din(w_dff_A_9RwiuLbM9_1),.clk(gclk));
	jdff dff_A_7lPIcV558_1(.dout(w_dff_A_9RwiuLbM9_1),.din(w_dff_A_7lPIcV558_1),.clk(gclk));
	jdff dff_B_swAYl7xU4_1(.din(n1793),.dout(w_dff_B_swAYl7xU4_1),.clk(gclk));
	jdff dff_A_WItlfLpC4_1(.dout(w_n1768_0[1]),.din(w_dff_A_WItlfLpC4_1),.clk(gclk));
	jdff dff_B_LzPbpWEu3_1(.din(n1766),.dout(w_dff_B_LzPbpWEu3_1),.clk(gclk));
	jdff dff_B_H6mtBv1K6_2(.din(n1730),.dout(w_dff_B_H6mtBv1K6_2),.clk(gclk));
	jdff dff_B_9XvtSTpv6_2(.din(w_dff_B_H6mtBv1K6_2),.dout(w_dff_B_9XvtSTpv6_2),.clk(gclk));
	jdff dff_B_yb1kLai44_2(.din(w_dff_B_9XvtSTpv6_2),.dout(w_dff_B_yb1kLai44_2),.clk(gclk));
	jdff dff_B_9JzcRiYJ3_2(.din(w_dff_B_yb1kLai44_2),.dout(w_dff_B_9JzcRiYJ3_2),.clk(gclk));
	jdff dff_B_kdxV89qc4_2(.din(w_dff_B_9JzcRiYJ3_2),.dout(w_dff_B_kdxV89qc4_2),.clk(gclk));
	jdff dff_B_1nr48IKx1_2(.din(w_dff_B_kdxV89qc4_2),.dout(w_dff_B_1nr48IKx1_2),.clk(gclk));
	jdff dff_B_anXGj3Lk6_2(.din(w_dff_B_1nr48IKx1_2),.dout(w_dff_B_anXGj3Lk6_2),.clk(gclk));
	jdff dff_B_gP6AfZ4R5_2(.din(w_dff_B_anXGj3Lk6_2),.dout(w_dff_B_gP6AfZ4R5_2),.clk(gclk));
	jdff dff_B_l7rqyiSV9_2(.din(w_dff_B_gP6AfZ4R5_2),.dout(w_dff_B_l7rqyiSV9_2),.clk(gclk));
	jdff dff_B_ShfQ0cvR2_2(.din(w_dff_B_l7rqyiSV9_2),.dout(w_dff_B_ShfQ0cvR2_2),.clk(gclk));
	jdff dff_B_svNpG9i57_2(.din(w_dff_B_ShfQ0cvR2_2),.dout(w_dff_B_svNpG9i57_2),.clk(gclk));
	jdff dff_B_xp2N5JwY0_2(.din(w_dff_B_svNpG9i57_2),.dout(w_dff_B_xp2N5JwY0_2),.clk(gclk));
	jdff dff_B_jlivo5LI9_2(.din(w_dff_B_xp2N5JwY0_2),.dout(w_dff_B_jlivo5LI9_2),.clk(gclk));
	jdff dff_B_ej2HIOCH3_2(.din(w_dff_B_jlivo5LI9_2),.dout(w_dff_B_ej2HIOCH3_2),.clk(gclk));
	jdff dff_B_6jU6beEu7_2(.din(w_dff_B_ej2HIOCH3_2),.dout(w_dff_B_6jU6beEu7_2),.clk(gclk));
	jdff dff_B_aEVKyXID7_2(.din(w_dff_B_6jU6beEu7_2),.dout(w_dff_B_aEVKyXID7_2),.clk(gclk));
	jdff dff_B_ZU662TJJ7_2(.din(w_dff_B_aEVKyXID7_2),.dout(w_dff_B_ZU662TJJ7_2),.clk(gclk));
	jdff dff_B_4qnuRD3s8_2(.din(w_dff_B_ZU662TJJ7_2),.dout(w_dff_B_4qnuRD3s8_2),.clk(gclk));
	jdff dff_B_9Gx5wGeG1_2(.din(w_dff_B_4qnuRD3s8_2),.dout(w_dff_B_9Gx5wGeG1_2),.clk(gclk));
	jdff dff_B_Yo0Vf7SH7_2(.din(w_dff_B_9Gx5wGeG1_2),.dout(w_dff_B_Yo0Vf7SH7_2),.clk(gclk));
	jdff dff_B_LbMODvhb2_2(.din(w_dff_B_Yo0Vf7SH7_2),.dout(w_dff_B_LbMODvhb2_2),.clk(gclk));
	jdff dff_B_wrDSOEST9_2(.din(w_dff_B_LbMODvhb2_2),.dout(w_dff_B_wrDSOEST9_2),.clk(gclk));
	jdff dff_B_EIvnxcR78_2(.din(w_dff_B_wrDSOEST9_2),.dout(w_dff_B_EIvnxcR78_2),.clk(gclk));
	jdff dff_B_5v8GyuaA4_2(.din(w_dff_B_EIvnxcR78_2),.dout(w_dff_B_5v8GyuaA4_2),.clk(gclk));
	jdff dff_B_Yhoexs5x1_2(.din(w_dff_B_5v8GyuaA4_2),.dout(w_dff_B_Yhoexs5x1_2),.clk(gclk));
	jdff dff_B_OrtWqyKA3_2(.din(w_dff_B_Yhoexs5x1_2),.dout(w_dff_B_OrtWqyKA3_2),.clk(gclk));
	jdff dff_B_tgn7m4K28_2(.din(w_dff_B_OrtWqyKA3_2),.dout(w_dff_B_tgn7m4K28_2),.clk(gclk));
	jdff dff_B_yJcC1C7Q1_2(.din(w_dff_B_tgn7m4K28_2),.dout(w_dff_B_yJcC1C7Q1_2),.clk(gclk));
	jdff dff_B_UPcYNmSS2_2(.din(w_dff_B_yJcC1C7Q1_2),.dout(w_dff_B_UPcYNmSS2_2),.clk(gclk));
	jdff dff_B_RIwApUQW6_2(.din(w_dff_B_UPcYNmSS2_2),.dout(w_dff_B_RIwApUQW6_2),.clk(gclk));
	jdff dff_B_bQfhKYo91_2(.din(w_dff_B_RIwApUQW6_2),.dout(w_dff_B_bQfhKYo91_2),.clk(gclk));
	jdff dff_B_fMkyXAsr2_2(.din(w_dff_B_bQfhKYo91_2),.dout(w_dff_B_fMkyXAsr2_2),.clk(gclk));
	jdff dff_B_zsGQLSGN9_2(.din(w_dff_B_fMkyXAsr2_2),.dout(w_dff_B_zsGQLSGN9_2),.clk(gclk));
	jdff dff_B_9FlxtoOI5_2(.din(w_dff_B_zsGQLSGN9_2),.dout(w_dff_B_9FlxtoOI5_2),.clk(gclk));
	jdff dff_B_IQdKcivU4_2(.din(w_dff_B_9FlxtoOI5_2),.dout(w_dff_B_IQdKcivU4_2),.clk(gclk));
	jdff dff_B_CUKrA4Cw9_2(.din(w_dff_B_IQdKcivU4_2),.dout(w_dff_B_CUKrA4Cw9_2),.clk(gclk));
	jdff dff_B_Y9PhFo438_2(.din(w_dff_B_CUKrA4Cw9_2),.dout(w_dff_B_Y9PhFo438_2),.clk(gclk));
	jdff dff_B_LzbBETMS3_2(.din(w_dff_B_Y9PhFo438_2),.dout(w_dff_B_LzbBETMS3_2),.clk(gclk));
	jdff dff_B_957WxHNJ7_2(.din(w_dff_B_LzbBETMS3_2),.dout(w_dff_B_957WxHNJ7_2),.clk(gclk));
	jdff dff_B_rqZ2L9jc4_2(.din(w_dff_B_957WxHNJ7_2),.dout(w_dff_B_rqZ2L9jc4_2),.clk(gclk));
	jdff dff_B_tdgePMaP4_2(.din(w_dff_B_rqZ2L9jc4_2),.dout(w_dff_B_tdgePMaP4_2),.clk(gclk));
	jdff dff_B_gUyDHGLI0_2(.din(w_dff_B_tdgePMaP4_2),.dout(w_dff_B_gUyDHGLI0_2),.clk(gclk));
	jdff dff_B_9MgmbgsI1_2(.din(w_dff_B_gUyDHGLI0_2),.dout(w_dff_B_9MgmbgsI1_2),.clk(gclk));
	jdff dff_B_syFGDCgS1_2(.din(w_dff_B_9MgmbgsI1_2),.dout(w_dff_B_syFGDCgS1_2),.clk(gclk));
	jdff dff_B_utdgoEAV1_2(.din(w_dff_B_syFGDCgS1_2),.dout(w_dff_B_utdgoEAV1_2),.clk(gclk));
	jdff dff_B_YSxTucuZ5_2(.din(w_dff_B_utdgoEAV1_2),.dout(w_dff_B_YSxTucuZ5_2),.clk(gclk));
	jdff dff_B_j7cEDYbT1_2(.din(w_dff_B_YSxTucuZ5_2),.dout(w_dff_B_j7cEDYbT1_2),.clk(gclk));
	jdff dff_B_wcq1zbGT0_2(.din(w_dff_B_j7cEDYbT1_2),.dout(w_dff_B_wcq1zbGT0_2),.clk(gclk));
	jdff dff_B_umlEhmbA0_2(.din(w_dff_B_wcq1zbGT0_2),.dout(w_dff_B_umlEhmbA0_2),.clk(gclk));
	jdff dff_B_8T0UyFxb2_2(.din(w_dff_B_umlEhmbA0_2),.dout(w_dff_B_8T0UyFxb2_2),.clk(gclk));
	jdff dff_B_xe0e7oJ50_2(.din(w_dff_B_8T0UyFxb2_2),.dout(w_dff_B_xe0e7oJ50_2),.clk(gclk));
	jdff dff_B_bUQI7BuH1_2(.din(n1733),.dout(w_dff_B_bUQI7BuH1_2),.clk(gclk));
	jdff dff_B_cbqqkSOt3_1(.din(n1731),.dout(w_dff_B_cbqqkSOt3_1),.clk(gclk));
	jdff dff_B_4WuJtOWd5_2(.din(n1689),.dout(w_dff_B_4WuJtOWd5_2),.clk(gclk));
	jdff dff_B_YOyTYtVv5_2(.din(w_dff_B_4WuJtOWd5_2),.dout(w_dff_B_YOyTYtVv5_2),.clk(gclk));
	jdff dff_B_d9tLDOwU8_2(.din(w_dff_B_YOyTYtVv5_2),.dout(w_dff_B_d9tLDOwU8_2),.clk(gclk));
	jdff dff_B_BqLPgxoY5_2(.din(w_dff_B_d9tLDOwU8_2),.dout(w_dff_B_BqLPgxoY5_2),.clk(gclk));
	jdff dff_B_a0WegON35_2(.din(w_dff_B_BqLPgxoY5_2),.dout(w_dff_B_a0WegON35_2),.clk(gclk));
	jdff dff_B_0Z9Q4Un26_2(.din(w_dff_B_a0WegON35_2),.dout(w_dff_B_0Z9Q4Un26_2),.clk(gclk));
	jdff dff_B_N1F4fEdb1_2(.din(w_dff_B_0Z9Q4Un26_2),.dout(w_dff_B_N1F4fEdb1_2),.clk(gclk));
	jdff dff_B_eTMkIJLa1_2(.din(w_dff_B_N1F4fEdb1_2),.dout(w_dff_B_eTMkIJLa1_2),.clk(gclk));
	jdff dff_B_djqRUxpN1_2(.din(w_dff_B_eTMkIJLa1_2),.dout(w_dff_B_djqRUxpN1_2),.clk(gclk));
	jdff dff_B_o3iJ7W9p2_2(.din(w_dff_B_djqRUxpN1_2),.dout(w_dff_B_o3iJ7W9p2_2),.clk(gclk));
	jdff dff_B_QkBUDKmJ9_2(.din(w_dff_B_o3iJ7W9p2_2),.dout(w_dff_B_QkBUDKmJ9_2),.clk(gclk));
	jdff dff_B_HMeZxEat8_2(.din(w_dff_B_QkBUDKmJ9_2),.dout(w_dff_B_HMeZxEat8_2),.clk(gclk));
	jdff dff_B_VgB0xkrC5_2(.din(w_dff_B_HMeZxEat8_2),.dout(w_dff_B_VgB0xkrC5_2),.clk(gclk));
	jdff dff_B_edFqKEm53_2(.din(w_dff_B_VgB0xkrC5_2),.dout(w_dff_B_edFqKEm53_2),.clk(gclk));
	jdff dff_B_fH4Oxttf8_2(.din(w_dff_B_edFqKEm53_2),.dout(w_dff_B_fH4Oxttf8_2),.clk(gclk));
	jdff dff_B_NOTK3CBt7_2(.din(w_dff_B_fH4Oxttf8_2),.dout(w_dff_B_NOTK3CBt7_2),.clk(gclk));
	jdff dff_B_dPVSB4Nc7_2(.din(w_dff_B_NOTK3CBt7_2),.dout(w_dff_B_dPVSB4Nc7_2),.clk(gclk));
	jdff dff_B_aFdUhKba3_2(.din(w_dff_B_dPVSB4Nc7_2),.dout(w_dff_B_aFdUhKba3_2),.clk(gclk));
	jdff dff_B_qMp8mdia4_2(.din(w_dff_B_aFdUhKba3_2),.dout(w_dff_B_qMp8mdia4_2),.clk(gclk));
	jdff dff_B_RoXPRaTS4_2(.din(w_dff_B_qMp8mdia4_2),.dout(w_dff_B_RoXPRaTS4_2),.clk(gclk));
	jdff dff_B_bJhY5KSt2_2(.din(w_dff_B_RoXPRaTS4_2),.dout(w_dff_B_bJhY5KSt2_2),.clk(gclk));
	jdff dff_B_EZ6E0mIH9_2(.din(w_dff_B_bJhY5KSt2_2),.dout(w_dff_B_EZ6E0mIH9_2),.clk(gclk));
	jdff dff_B_LiOHpp0s8_2(.din(w_dff_B_EZ6E0mIH9_2),.dout(w_dff_B_LiOHpp0s8_2),.clk(gclk));
	jdff dff_B_UvNqbsXi3_2(.din(w_dff_B_LiOHpp0s8_2),.dout(w_dff_B_UvNqbsXi3_2),.clk(gclk));
	jdff dff_B_ZYkrU6122_2(.din(w_dff_B_UvNqbsXi3_2),.dout(w_dff_B_ZYkrU6122_2),.clk(gclk));
	jdff dff_B_kyw1KR4g9_2(.din(w_dff_B_ZYkrU6122_2),.dout(w_dff_B_kyw1KR4g9_2),.clk(gclk));
	jdff dff_B_P62hqi5Z4_2(.din(w_dff_B_kyw1KR4g9_2),.dout(w_dff_B_P62hqi5Z4_2),.clk(gclk));
	jdff dff_B_txPKKbPr8_2(.din(w_dff_B_P62hqi5Z4_2),.dout(w_dff_B_txPKKbPr8_2),.clk(gclk));
	jdff dff_B_41AylPxe4_2(.din(w_dff_B_txPKKbPr8_2),.dout(w_dff_B_41AylPxe4_2),.clk(gclk));
	jdff dff_B_mOKvSalK5_2(.din(w_dff_B_41AylPxe4_2),.dout(w_dff_B_mOKvSalK5_2),.clk(gclk));
	jdff dff_B_z47xiuzn1_2(.din(w_dff_B_mOKvSalK5_2),.dout(w_dff_B_z47xiuzn1_2),.clk(gclk));
	jdff dff_B_K2Habuhe4_2(.din(w_dff_B_z47xiuzn1_2),.dout(w_dff_B_K2Habuhe4_2),.clk(gclk));
	jdff dff_B_KRwvONfS6_2(.din(w_dff_B_K2Habuhe4_2),.dout(w_dff_B_KRwvONfS6_2),.clk(gclk));
	jdff dff_B_3NSyxBTa3_2(.din(w_dff_B_KRwvONfS6_2),.dout(w_dff_B_3NSyxBTa3_2),.clk(gclk));
	jdff dff_B_ExW8D8dv7_2(.din(w_dff_B_3NSyxBTa3_2),.dout(w_dff_B_ExW8D8dv7_2),.clk(gclk));
	jdff dff_B_GnmsHfMT3_2(.din(w_dff_B_ExW8D8dv7_2),.dout(w_dff_B_GnmsHfMT3_2),.clk(gclk));
	jdff dff_B_GJ6aRfhb6_2(.din(w_dff_B_GnmsHfMT3_2),.dout(w_dff_B_GJ6aRfhb6_2),.clk(gclk));
	jdff dff_B_yQM7XMqw2_2(.din(w_dff_B_GJ6aRfhb6_2),.dout(w_dff_B_yQM7XMqw2_2),.clk(gclk));
	jdff dff_B_vBvVXIyN1_2(.din(w_dff_B_yQM7XMqw2_2),.dout(w_dff_B_vBvVXIyN1_2),.clk(gclk));
	jdff dff_B_EN9LNgMC8_2(.din(w_dff_B_vBvVXIyN1_2),.dout(w_dff_B_EN9LNgMC8_2),.clk(gclk));
	jdff dff_B_sg1tNUUs7_2(.din(w_dff_B_EN9LNgMC8_2),.dout(w_dff_B_sg1tNUUs7_2),.clk(gclk));
	jdff dff_B_FcxZ8jjA7_2(.din(w_dff_B_sg1tNUUs7_2),.dout(w_dff_B_FcxZ8jjA7_2),.clk(gclk));
	jdff dff_B_Z0iUD3KS2_2(.din(w_dff_B_FcxZ8jjA7_2),.dout(w_dff_B_Z0iUD3KS2_2),.clk(gclk));
	jdff dff_B_GnLQSwgO7_2(.din(w_dff_B_Z0iUD3KS2_2),.dout(w_dff_B_GnLQSwgO7_2),.clk(gclk));
	jdff dff_B_mYHW4hAb0_2(.din(w_dff_B_GnLQSwgO7_2),.dout(w_dff_B_mYHW4hAb0_2),.clk(gclk));
	jdff dff_B_5F8Eq4700_2(.din(w_dff_B_mYHW4hAb0_2),.dout(w_dff_B_5F8Eq4700_2),.clk(gclk));
	jdff dff_B_nj4zgaFg1_2(.din(w_dff_B_5F8Eq4700_2),.dout(w_dff_B_nj4zgaFg1_2),.clk(gclk));
	jdff dff_B_jVVl5q6J8_2(.din(n1692),.dout(w_dff_B_jVVl5q6J8_2),.clk(gclk));
	jdff dff_B_YNu2zp3w3_1(.din(n1690),.dout(w_dff_B_YNu2zp3w3_1),.clk(gclk));
	jdff dff_B_TUQ9DmFl3_2(.din(n1638),.dout(w_dff_B_TUQ9DmFl3_2),.clk(gclk));
	jdff dff_B_2OdILCNc6_2(.din(w_dff_B_TUQ9DmFl3_2),.dout(w_dff_B_2OdILCNc6_2),.clk(gclk));
	jdff dff_B_OjvU5On85_2(.din(w_dff_B_2OdILCNc6_2),.dout(w_dff_B_OjvU5On85_2),.clk(gclk));
	jdff dff_B_mLQhD9fW2_2(.din(w_dff_B_OjvU5On85_2),.dout(w_dff_B_mLQhD9fW2_2),.clk(gclk));
	jdff dff_B_oWwDZk5Y7_2(.din(w_dff_B_mLQhD9fW2_2),.dout(w_dff_B_oWwDZk5Y7_2),.clk(gclk));
	jdff dff_B_GoOhqLBZ2_2(.din(w_dff_B_oWwDZk5Y7_2),.dout(w_dff_B_GoOhqLBZ2_2),.clk(gclk));
	jdff dff_B_eizSrCK38_2(.din(w_dff_B_GoOhqLBZ2_2),.dout(w_dff_B_eizSrCK38_2),.clk(gclk));
	jdff dff_B_bcoynlxS0_2(.din(w_dff_B_eizSrCK38_2),.dout(w_dff_B_bcoynlxS0_2),.clk(gclk));
	jdff dff_B_3A4MX6ls7_2(.din(w_dff_B_bcoynlxS0_2),.dout(w_dff_B_3A4MX6ls7_2),.clk(gclk));
	jdff dff_B_tWhHESrw8_2(.din(w_dff_B_3A4MX6ls7_2),.dout(w_dff_B_tWhHESrw8_2),.clk(gclk));
	jdff dff_B_VIfc0kX26_2(.din(w_dff_B_tWhHESrw8_2),.dout(w_dff_B_VIfc0kX26_2),.clk(gclk));
	jdff dff_B_zEMQBD2f6_2(.din(w_dff_B_VIfc0kX26_2),.dout(w_dff_B_zEMQBD2f6_2),.clk(gclk));
	jdff dff_B_BKvZJwyW9_2(.din(w_dff_B_zEMQBD2f6_2),.dout(w_dff_B_BKvZJwyW9_2),.clk(gclk));
	jdff dff_B_yNQHINSw0_2(.din(w_dff_B_BKvZJwyW9_2),.dout(w_dff_B_yNQHINSw0_2),.clk(gclk));
	jdff dff_B_qfR2ewqZ8_2(.din(w_dff_B_yNQHINSw0_2),.dout(w_dff_B_qfR2ewqZ8_2),.clk(gclk));
	jdff dff_B_K5ZmDyLb1_2(.din(w_dff_B_qfR2ewqZ8_2),.dout(w_dff_B_K5ZmDyLb1_2),.clk(gclk));
	jdff dff_B_0YAJk6Uj1_2(.din(w_dff_B_K5ZmDyLb1_2),.dout(w_dff_B_0YAJk6Uj1_2),.clk(gclk));
	jdff dff_B_z8BhNc4j2_2(.din(w_dff_B_0YAJk6Uj1_2),.dout(w_dff_B_z8BhNc4j2_2),.clk(gclk));
	jdff dff_B_Y3ZIg1M75_2(.din(w_dff_B_z8BhNc4j2_2),.dout(w_dff_B_Y3ZIg1M75_2),.clk(gclk));
	jdff dff_B_YSqnfV811_2(.din(w_dff_B_Y3ZIg1M75_2),.dout(w_dff_B_YSqnfV811_2),.clk(gclk));
	jdff dff_B_ai8j6rzt5_2(.din(w_dff_B_YSqnfV811_2),.dout(w_dff_B_ai8j6rzt5_2),.clk(gclk));
	jdff dff_B_a98vFQd63_2(.din(w_dff_B_ai8j6rzt5_2),.dout(w_dff_B_a98vFQd63_2),.clk(gclk));
	jdff dff_B_CsJ1R2Tr4_2(.din(w_dff_B_a98vFQd63_2),.dout(w_dff_B_CsJ1R2Tr4_2),.clk(gclk));
	jdff dff_B_aDMptzkZ5_2(.din(w_dff_B_CsJ1R2Tr4_2),.dout(w_dff_B_aDMptzkZ5_2),.clk(gclk));
	jdff dff_B_ZLN7o7mO9_2(.din(w_dff_B_aDMptzkZ5_2),.dout(w_dff_B_ZLN7o7mO9_2),.clk(gclk));
	jdff dff_B_W97JhkRO2_2(.din(w_dff_B_ZLN7o7mO9_2),.dout(w_dff_B_W97JhkRO2_2),.clk(gclk));
	jdff dff_B_GUzZIFy88_2(.din(w_dff_B_W97JhkRO2_2),.dout(w_dff_B_GUzZIFy88_2),.clk(gclk));
	jdff dff_B_5vcJ02eG7_2(.din(w_dff_B_GUzZIFy88_2),.dout(w_dff_B_5vcJ02eG7_2),.clk(gclk));
	jdff dff_B_LgymVEUt2_2(.din(w_dff_B_5vcJ02eG7_2),.dout(w_dff_B_LgymVEUt2_2),.clk(gclk));
	jdff dff_B_SrU3J8Tn8_2(.din(w_dff_B_LgymVEUt2_2),.dout(w_dff_B_SrU3J8Tn8_2),.clk(gclk));
	jdff dff_B_90hJe6is0_2(.din(w_dff_B_SrU3J8Tn8_2),.dout(w_dff_B_90hJe6is0_2),.clk(gclk));
	jdff dff_B_An0iTvcV8_2(.din(w_dff_B_90hJe6is0_2),.dout(w_dff_B_An0iTvcV8_2),.clk(gclk));
	jdff dff_B_CV5w5Dn94_2(.din(w_dff_B_An0iTvcV8_2),.dout(w_dff_B_CV5w5Dn94_2),.clk(gclk));
	jdff dff_B_TMIYBPzl7_2(.din(w_dff_B_CV5w5Dn94_2),.dout(w_dff_B_TMIYBPzl7_2),.clk(gclk));
	jdff dff_B_GfeaITEK3_2(.din(w_dff_B_TMIYBPzl7_2),.dout(w_dff_B_GfeaITEK3_2),.clk(gclk));
	jdff dff_B_o6gHOwCh1_2(.din(w_dff_B_GfeaITEK3_2),.dout(w_dff_B_o6gHOwCh1_2),.clk(gclk));
	jdff dff_B_N1nDXXcd8_2(.din(w_dff_B_o6gHOwCh1_2),.dout(w_dff_B_N1nDXXcd8_2),.clk(gclk));
	jdff dff_B_X9SB6rxh9_2(.din(w_dff_B_N1nDXXcd8_2),.dout(w_dff_B_X9SB6rxh9_2),.clk(gclk));
	jdff dff_B_AvYioCkM2_2(.din(w_dff_B_X9SB6rxh9_2),.dout(w_dff_B_AvYioCkM2_2),.clk(gclk));
	jdff dff_B_9ONkPx6P2_2(.din(w_dff_B_AvYioCkM2_2),.dout(w_dff_B_9ONkPx6P2_2),.clk(gclk));
	jdff dff_B_sS0vzrBr8_2(.din(w_dff_B_9ONkPx6P2_2),.dout(w_dff_B_sS0vzrBr8_2),.clk(gclk));
	jdff dff_B_hSEr7CFm3_2(.din(w_dff_B_sS0vzrBr8_2),.dout(w_dff_B_hSEr7CFm3_2),.clk(gclk));
	jdff dff_B_gg96ixUT7_2(.din(w_dff_B_hSEr7CFm3_2),.dout(w_dff_B_gg96ixUT7_2),.clk(gclk));
	jdff dff_B_RlKTCuxy7_2(.din(n1641),.dout(w_dff_B_RlKTCuxy7_2),.clk(gclk));
	jdff dff_B_jPDNsV4f5_1(.din(n1639),.dout(w_dff_B_jPDNsV4f5_1),.clk(gclk));
	jdff dff_B_FWhxwsyp1_2(.din(n1581),.dout(w_dff_B_FWhxwsyp1_2),.clk(gclk));
	jdff dff_B_hN6NoHL09_2(.din(w_dff_B_FWhxwsyp1_2),.dout(w_dff_B_hN6NoHL09_2),.clk(gclk));
	jdff dff_B_LmcKsD8k2_2(.din(w_dff_B_hN6NoHL09_2),.dout(w_dff_B_LmcKsD8k2_2),.clk(gclk));
	jdff dff_B_HEZbZo4H0_2(.din(w_dff_B_LmcKsD8k2_2),.dout(w_dff_B_HEZbZo4H0_2),.clk(gclk));
	jdff dff_B_a5JieUma1_2(.din(w_dff_B_HEZbZo4H0_2),.dout(w_dff_B_a5JieUma1_2),.clk(gclk));
	jdff dff_B_SZllBtwh5_2(.din(w_dff_B_a5JieUma1_2),.dout(w_dff_B_SZllBtwh5_2),.clk(gclk));
	jdff dff_B_CWE7WaOw3_2(.din(w_dff_B_SZllBtwh5_2),.dout(w_dff_B_CWE7WaOw3_2),.clk(gclk));
	jdff dff_B_T5ucWDJP3_2(.din(w_dff_B_CWE7WaOw3_2),.dout(w_dff_B_T5ucWDJP3_2),.clk(gclk));
	jdff dff_B_vUhUwuC36_2(.din(w_dff_B_T5ucWDJP3_2),.dout(w_dff_B_vUhUwuC36_2),.clk(gclk));
	jdff dff_B_qWV9Z5bT0_2(.din(w_dff_B_vUhUwuC36_2),.dout(w_dff_B_qWV9Z5bT0_2),.clk(gclk));
	jdff dff_B_S8Pv2Su02_2(.din(w_dff_B_qWV9Z5bT0_2),.dout(w_dff_B_S8Pv2Su02_2),.clk(gclk));
	jdff dff_B_vTyWXmq13_2(.din(w_dff_B_S8Pv2Su02_2),.dout(w_dff_B_vTyWXmq13_2),.clk(gclk));
	jdff dff_B_bPFVtFv45_2(.din(w_dff_B_vTyWXmq13_2),.dout(w_dff_B_bPFVtFv45_2),.clk(gclk));
	jdff dff_B_N6U4zmN03_2(.din(w_dff_B_bPFVtFv45_2),.dout(w_dff_B_N6U4zmN03_2),.clk(gclk));
	jdff dff_B_SSUob3hE8_2(.din(w_dff_B_N6U4zmN03_2),.dout(w_dff_B_SSUob3hE8_2),.clk(gclk));
	jdff dff_B_NT6MnoK61_2(.din(w_dff_B_SSUob3hE8_2),.dout(w_dff_B_NT6MnoK61_2),.clk(gclk));
	jdff dff_B_5oPMN6Tr6_2(.din(w_dff_B_NT6MnoK61_2),.dout(w_dff_B_5oPMN6Tr6_2),.clk(gclk));
	jdff dff_B_fIFqLAVR8_2(.din(w_dff_B_5oPMN6Tr6_2),.dout(w_dff_B_fIFqLAVR8_2),.clk(gclk));
	jdff dff_B_A35TbZZY1_2(.din(w_dff_B_fIFqLAVR8_2),.dout(w_dff_B_A35TbZZY1_2),.clk(gclk));
	jdff dff_B_TuHtGioY2_2(.din(w_dff_B_A35TbZZY1_2),.dout(w_dff_B_TuHtGioY2_2),.clk(gclk));
	jdff dff_B_EenB9Ik38_2(.din(w_dff_B_TuHtGioY2_2),.dout(w_dff_B_EenB9Ik38_2),.clk(gclk));
	jdff dff_B_zcY1HmAm6_2(.din(w_dff_B_EenB9Ik38_2),.dout(w_dff_B_zcY1HmAm6_2),.clk(gclk));
	jdff dff_B_9DLkRjS03_2(.din(w_dff_B_zcY1HmAm6_2),.dout(w_dff_B_9DLkRjS03_2),.clk(gclk));
	jdff dff_B_vGgx5UOl8_2(.din(w_dff_B_9DLkRjS03_2),.dout(w_dff_B_vGgx5UOl8_2),.clk(gclk));
	jdff dff_B_0ss9W9jf0_2(.din(w_dff_B_vGgx5UOl8_2),.dout(w_dff_B_0ss9W9jf0_2),.clk(gclk));
	jdff dff_B_sQzvEDJH0_2(.din(w_dff_B_0ss9W9jf0_2),.dout(w_dff_B_sQzvEDJH0_2),.clk(gclk));
	jdff dff_B_Hj9Y9dzq5_2(.din(w_dff_B_sQzvEDJH0_2),.dout(w_dff_B_Hj9Y9dzq5_2),.clk(gclk));
	jdff dff_B_RE2q9mKr2_2(.din(w_dff_B_Hj9Y9dzq5_2),.dout(w_dff_B_RE2q9mKr2_2),.clk(gclk));
	jdff dff_B_cgkKqhsh2_2(.din(w_dff_B_RE2q9mKr2_2),.dout(w_dff_B_cgkKqhsh2_2),.clk(gclk));
	jdff dff_B_IllvyTv35_2(.din(w_dff_B_cgkKqhsh2_2),.dout(w_dff_B_IllvyTv35_2),.clk(gclk));
	jdff dff_B_OzYlfES70_2(.din(w_dff_B_IllvyTv35_2),.dout(w_dff_B_OzYlfES70_2),.clk(gclk));
	jdff dff_B_CupDJq5Y7_2(.din(w_dff_B_OzYlfES70_2),.dout(w_dff_B_CupDJq5Y7_2),.clk(gclk));
	jdff dff_B_V3vfjcVw0_2(.din(w_dff_B_CupDJq5Y7_2),.dout(w_dff_B_V3vfjcVw0_2),.clk(gclk));
	jdff dff_B_Cfb4vqSe7_2(.din(w_dff_B_V3vfjcVw0_2),.dout(w_dff_B_Cfb4vqSe7_2),.clk(gclk));
	jdff dff_B_4C0WKNQH4_2(.din(w_dff_B_Cfb4vqSe7_2),.dout(w_dff_B_4C0WKNQH4_2),.clk(gclk));
	jdff dff_B_i96nFEU98_2(.din(w_dff_B_4C0WKNQH4_2),.dout(w_dff_B_i96nFEU98_2),.clk(gclk));
	jdff dff_B_ypZ51DHP7_2(.din(w_dff_B_i96nFEU98_2),.dout(w_dff_B_ypZ51DHP7_2),.clk(gclk));
	jdff dff_B_zk0hrgOT6_2(.din(w_dff_B_ypZ51DHP7_2),.dout(w_dff_B_zk0hrgOT6_2),.clk(gclk));
	jdff dff_B_fmCt4rpQ0_2(.din(w_dff_B_zk0hrgOT6_2),.dout(w_dff_B_fmCt4rpQ0_2),.clk(gclk));
	jdff dff_B_Us3zuZTo6_2(.din(n1584),.dout(w_dff_B_Us3zuZTo6_2),.clk(gclk));
	jdff dff_B_8o2FsipG4_1(.din(n1582),.dout(w_dff_B_8o2FsipG4_1),.clk(gclk));
	jdff dff_B_yvHiPnQw7_2(.din(n1517),.dout(w_dff_B_yvHiPnQw7_2),.clk(gclk));
	jdff dff_B_jUVPFEwC2_2(.din(w_dff_B_yvHiPnQw7_2),.dout(w_dff_B_jUVPFEwC2_2),.clk(gclk));
	jdff dff_B_GJuLF0m44_2(.din(w_dff_B_jUVPFEwC2_2),.dout(w_dff_B_GJuLF0m44_2),.clk(gclk));
	jdff dff_B_b12wuBNb6_2(.din(w_dff_B_GJuLF0m44_2),.dout(w_dff_B_b12wuBNb6_2),.clk(gclk));
	jdff dff_B_qay5OBGx1_2(.din(w_dff_B_b12wuBNb6_2),.dout(w_dff_B_qay5OBGx1_2),.clk(gclk));
	jdff dff_B_lP0gwImO0_2(.din(w_dff_B_qay5OBGx1_2),.dout(w_dff_B_lP0gwImO0_2),.clk(gclk));
	jdff dff_B_k7XucLjP3_2(.din(w_dff_B_lP0gwImO0_2),.dout(w_dff_B_k7XucLjP3_2),.clk(gclk));
	jdff dff_B_NqDDxPS28_2(.din(w_dff_B_k7XucLjP3_2),.dout(w_dff_B_NqDDxPS28_2),.clk(gclk));
	jdff dff_B_0JQlx2xx9_2(.din(w_dff_B_NqDDxPS28_2),.dout(w_dff_B_0JQlx2xx9_2),.clk(gclk));
	jdff dff_B_dDyXOI5Y6_2(.din(w_dff_B_0JQlx2xx9_2),.dout(w_dff_B_dDyXOI5Y6_2),.clk(gclk));
	jdff dff_B_3T4EUipr5_2(.din(w_dff_B_dDyXOI5Y6_2),.dout(w_dff_B_3T4EUipr5_2),.clk(gclk));
	jdff dff_B_EmAbx1th6_2(.din(w_dff_B_3T4EUipr5_2),.dout(w_dff_B_EmAbx1th6_2),.clk(gclk));
	jdff dff_B_zDFDPh4S8_2(.din(w_dff_B_EmAbx1th6_2),.dout(w_dff_B_zDFDPh4S8_2),.clk(gclk));
	jdff dff_B_MmorXoxh8_2(.din(w_dff_B_zDFDPh4S8_2),.dout(w_dff_B_MmorXoxh8_2),.clk(gclk));
	jdff dff_B_7aMezkkc7_2(.din(w_dff_B_MmorXoxh8_2),.dout(w_dff_B_7aMezkkc7_2),.clk(gclk));
	jdff dff_B_PZUNlUiX7_2(.din(w_dff_B_7aMezkkc7_2),.dout(w_dff_B_PZUNlUiX7_2),.clk(gclk));
	jdff dff_B_C1bhB9y15_2(.din(w_dff_B_PZUNlUiX7_2),.dout(w_dff_B_C1bhB9y15_2),.clk(gclk));
	jdff dff_B_wL0SRZO77_2(.din(w_dff_B_C1bhB9y15_2),.dout(w_dff_B_wL0SRZO77_2),.clk(gclk));
	jdff dff_B_PQmflSPZ8_2(.din(w_dff_B_wL0SRZO77_2),.dout(w_dff_B_PQmflSPZ8_2),.clk(gclk));
	jdff dff_B_2bVdqd6s8_2(.din(w_dff_B_PQmflSPZ8_2),.dout(w_dff_B_2bVdqd6s8_2),.clk(gclk));
	jdff dff_B_DQ6r8t1B7_2(.din(w_dff_B_2bVdqd6s8_2),.dout(w_dff_B_DQ6r8t1B7_2),.clk(gclk));
	jdff dff_B_cIbBd5qZ7_2(.din(w_dff_B_DQ6r8t1B7_2),.dout(w_dff_B_cIbBd5qZ7_2),.clk(gclk));
	jdff dff_B_RacqNaBe5_2(.din(w_dff_B_cIbBd5qZ7_2),.dout(w_dff_B_RacqNaBe5_2),.clk(gclk));
	jdff dff_B_nD6vQqlA2_2(.din(w_dff_B_RacqNaBe5_2),.dout(w_dff_B_nD6vQqlA2_2),.clk(gclk));
	jdff dff_B_uNVs8MvF4_2(.din(w_dff_B_nD6vQqlA2_2),.dout(w_dff_B_uNVs8MvF4_2),.clk(gclk));
	jdff dff_B_JQlG46sZ5_2(.din(w_dff_B_uNVs8MvF4_2),.dout(w_dff_B_JQlG46sZ5_2),.clk(gclk));
	jdff dff_B_VGko9RUY8_2(.din(w_dff_B_JQlG46sZ5_2),.dout(w_dff_B_VGko9RUY8_2),.clk(gclk));
	jdff dff_B_HTldysDF6_2(.din(w_dff_B_VGko9RUY8_2),.dout(w_dff_B_HTldysDF6_2),.clk(gclk));
	jdff dff_B_JzVxaj0z2_2(.din(w_dff_B_HTldysDF6_2),.dout(w_dff_B_JzVxaj0z2_2),.clk(gclk));
	jdff dff_B_NyAFTD8h7_2(.din(w_dff_B_JzVxaj0z2_2),.dout(w_dff_B_NyAFTD8h7_2),.clk(gclk));
	jdff dff_B_H3rhAmjQ4_2(.din(w_dff_B_NyAFTD8h7_2),.dout(w_dff_B_H3rhAmjQ4_2),.clk(gclk));
	jdff dff_B_SUOXQVS70_2(.din(w_dff_B_H3rhAmjQ4_2),.dout(w_dff_B_SUOXQVS70_2),.clk(gclk));
	jdff dff_B_9UqHuJWk3_2(.din(w_dff_B_SUOXQVS70_2),.dout(w_dff_B_9UqHuJWk3_2),.clk(gclk));
	jdff dff_B_5af9HRqt5_2(.din(w_dff_B_9UqHuJWk3_2),.dout(w_dff_B_5af9HRqt5_2),.clk(gclk));
	jdff dff_B_68ngA5Vo5_2(.din(w_dff_B_5af9HRqt5_2),.dout(w_dff_B_68ngA5Vo5_2),.clk(gclk));
	jdff dff_B_OMES7jqo9_2(.din(n1520),.dout(w_dff_B_OMES7jqo9_2),.clk(gclk));
	jdff dff_B_u5IVoq2a4_1(.din(n1518),.dout(w_dff_B_u5IVoq2a4_1),.clk(gclk));
	jdff dff_B_YcFCBFPO3_2(.din(n1446),.dout(w_dff_B_YcFCBFPO3_2),.clk(gclk));
	jdff dff_B_w4zDWyvm6_2(.din(w_dff_B_YcFCBFPO3_2),.dout(w_dff_B_w4zDWyvm6_2),.clk(gclk));
	jdff dff_B_2JWSzrzO0_2(.din(w_dff_B_w4zDWyvm6_2),.dout(w_dff_B_2JWSzrzO0_2),.clk(gclk));
	jdff dff_B_oTIs4USt9_2(.din(w_dff_B_2JWSzrzO0_2),.dout(w_dff_B_oTIs4USt9_2),.clk(gclk));
	jdff dff_B_3zipsOJY5_2(.din(w_dff_B_oTIs4USt9_2),.dout(w_dff_B_3zipsOJY5_2),.clk(gclk));
	jdff dff_B_YIFSJtrs0_2(.din(w_dff_B_3zipsOJY5_2),.dout(w_dff_B_YIFSJtrs0_2),.clk(gclk));
	jdff dff_B_N4acTxeA6_2(.din(w_dff_B_YIFSJtrs0_2),.dout(w_dff_B_N4acTxeA6_2),.clk(gclk));
	jdff dff_B_eXEd1Tmq8_2(.din(w_dff_B_N4acTxeA6_2),.dout(w_dff_B_eXEd1Tmq8_2),.clk(gclk));
	jdff dff_B_21cSfqmk9_2(.din(w_dff_B_eXEd1Tmq8_2),.dout(w_dff_B_21cSfqmk9_2),.clk(gclk));
	jdff dff_B_OydAEvk49_2(.din(w_dff_B_21cSfqmk9_2),.dout(w_dff_B_OydAEvk49_2),.clk(gclk));
	jdff dff_B_zLqu2rxX3_2(.din(w_dff_B_OydAEvk49_2),.dout(w_dff_B_zLqu2rxX3_2),.clk(gclk));
	jdff dff_B_zXzp0jIM8_2(.din(w_dff_B_zLqu2rxX3_2),.dout(w_dff_B_zXzp0jIM8_2),.clk(gclk));
	jdff dff_B_anhUD9a27_2(.din(w_dff_B_zXzp0jIM8_2),.dout(w_dff_B_anhUD9a27_2),.clk(gclk));
	jdff dff_B_eE1Wg2bl5_2(.din(w_dff_B_anhUD9a27_2),.dout(w_dff_B_eE1Wg2bl5_2),.clk(gclk));
	jdff dff_B_MDKR1x8E2_2(.din(w_dff_B_eE1Wg2bl5_2),.dout(w_dff_B_MDKR1x8E2_2),.clk(gclk));
	jdff dff_B_2O9MIAMb3_2(.din(w_dff_B_MDKR1x8E2_2),.dout(w_dff_B_2O9MIAMb3_2),.clk(gclk));
	jdff dff_B_iNFgzxZ08_2(.din(w_dff_B_2O9MIAMb3_2),.dout(w_dff_B_iNFgzxZ08_2),.clk(gclk));
	jdff dff_B_U8aDgk9d7_2(.din(w_dff_B_iNFgzxZ08_2),.dout(w_dff_B_U8aDgk9d7_2),.clk(gclk));
	jdff dff_B_ufLv9hl44_2(.din(w_dff_B_U8aDgk9d7_2),.dout(w_dff_B_ufLv9hl44_2),.clk(gclk));
	jdff dff_B_8vwtoFUA6_2(.din(w_dff_B_ufLv9hl44_2),.dout(w_dff_B_8vwtoFUA6_2),.clk(gclk));
	jdff dff_B_n7xiUSD47_2(.din(w_dff_B_8vwtoFUA6_2),.dout(w_dff_B_n7xiUSD47_2),.clk(gclk));
	jdff dff_B_kciiJgb55_2(.din(w_dff_B_n7xiUSD47_2),.dout(w_dff_B_kciiJgb55_2),.clk(gclk));
	jdff dff_B_zEkxCo4z3_2(.din(w_dff_B_kciiJgb55_2),.dout(w_dff_B_zEkxCo4z3_2),.clk(gclk));
	jdff dff_B_pgNjoc4F8_2(.din(w_dff_B_zEkxCo4z3_2),.dout(w_dff_B_pgNjoc4F8_2),.clk(gclk));
	jdff dff_B_u9kmetFt3_2(.din(w_dff_B_pgNjoc4F8_2),.dout(w_dff_B_u9kmetFt3_2),.clk(gclk));
	jdff dff_B_ltVj1MsD6_2(.din(w_dff_B_u9kmetFt3_2),.dout(w_dff_B_ltVj1MsD6_2),.clk(gclk));
	jdff dff_B_W2YPltbM3_2(.din(w_dff_B_ltVj1MsD6_2),.dout(w_dff_B_W2YPltbM3_2),.clk(gclk));
	jdff dff_B_2oCdhB3n3_2(.din(w_dff_B_W2YPltbM3_2),.dout(w_dff_B_2oCdhB3n3_2),.clk(gclk));
	jdff dff_B_ajPvAAUC4_2(.din(w_dff_B_2oCdhB3n3_2),.dout(w_dff_B_ajPvAAUC4_2),.clk(gclk));
	jdff dff_B_jYZV3R8I4_2(.din(w_dff_B_ajPvAAUC4_2),.dout(w_dff_B_jYZV3R8I4_2),.clk(gclk));
	jdff dff_B_jjedWkFG1_2(.din(w_dff_B_jYZV3R8I4_2),.dout(w_dff_B_jjedWkFG1_2),.clk(gclk));
	jdff dff_B_njPQvG9e8_2(.din(n1449),.dout(w_dff_B_njPQvG9e8_2),.clk(gclk));
	jdff dff_B_DeIbx7lP9_1(.din(n1447),.dout(w_dff_B_DeIbx7lP9_1),.clk(gclk));
	jdff dff_B_8e4NqzHw4_2(.din(n1368),.dout(w_dff_B_8e4NqzHw4_2),.clk(gclk));
	jdff dff_B_9Vh8Bn5K4_2(.din(w_dff_B_8e4NqzHw4_2),.dout(w_dff_B_9Vh8Bn5K4_2),.clk(gclk));
	jdff dff_B_yRa6JZ6l7_2(.din(w_dff_B_9Vh8Bn5K4_2),.dout(w_dff_B_yRa6JZ6l7_2),.clk(gclk));
	jdff dff_B_zdwx9JsP5_2(.din(w_dff_B_yRa6JZ6l7_2),.dout(w_dff_B_zdwx9JsP5_2),.clk(gclk));
	jdff dff_B_3RknptOY1_2(.din(w_dff_B_zdwx9JsP5_2),.dout(w_dff_B_3RknptOY1_2),.clk(gclk));
	jdff dff_B_AOVLuSwa7_2(.din(w_dff_B_3RknptOY1_2),.dout(w_dff_B_AOVLuSwa7_2),.clk(gclk));
	jdff dff_B_wrNpn0Rv4_2(.din(w_dff_B_AOVLuSwa7_2),.dout(w_dff_B_wrNpn0Rv4_2),.clk(gclk));
	jdff dff_B_SuxR5NWe6_2(.din(w_dff_B_wrNpn0Rv4_2),.dout(w_dff_B_SuxR5NWe6_2),.clk(gclk));
	jdff dff_B_9Vxltf1N5_2(.din(w_dff_B_SuxR5NWe6_2),.dout(w_dff_B_9Vxltf1N5_2),.clk(gclk));
	jdff dff_B_oSCyB8iY8_2(.din(w_dff_B_9Vxltf1N5_2),.dout(w_dff_B_oSCyB8iY8_2),.clk(gclk));
	jdff dff_B_yrycadkq0_2(.din(w_dff_B_oSCyB8iY8_2),.dout(w_dff_B_yrycadkq0_2),.clk(gclk));
	jdff dff_B_vIIsJsSq8_2(.din(w_dff_B_yrycadkq0_2),.dout(w_dff_B_vIIsJsSq8_2),.clk(gclk));
	jdff dff_B_TgSk8gGZ1_2(.din(w_dff_B_vIIsJsSq8_2),.dout(w_dff_B_TgSk8gGZ1_2),.clk(gclk));
	jdff dff_B_TFTtsks27_2(.din(w_dff_B_TgSk8gGZ1_2),.dout(w_dff_B_TFTtsks27_2),.clk(gclk));
	jdff dff_B_RvZnRIGG5_2(.din(w_dff_B_TFTtsks27_2),.dout(w_dff_B_RvZnRIGG5_2),.clk(gclk));
	jdff dff_B_QD4U42DU1_2(.din(w_dff_B_RvZnRIGG5_2),.dout(w_dff_B_QD4U42DU1_2),.clk(gclk));
	jdff dff_B_0sF7O7788_2(.din(w_dff_B_QD4U42DU1_2),.dout(w_dff_B_0sF7O7788_2),.clk(gclk));
	jdff dff_B_VaE4exiy4_2(.din(w_dff_B_0sF7O7788_2),.dout(w_dff_B_VaE4exiy4_2),.clk(gclk));
	jdff dff_B_xy9r5xCJ6_2(.din(w_dff_B_VaE4exiy4_2),.dout(w_dff_B_xy9r5xCJ6_2),.clk(gclk));
	jdff dff_B_rrP0XZrv6_2(.din(w_dff_B_xy9r5xCJ6_2),.dout(w_dff_B_rrP0XZrv6_2),.clk(gclk));
	jdff dff_B_EjHAvBwx7_2(.din(w_dff_B_rrP0XZrv6_2),.dout(w_dff_B_EjHAvBwx7_2),.clk(gclk));
	jdff dff_B_dbN2Nquh8_2(.din(w_dff_B_EjHAvBwx7_2),.dout(w_dff_B_dbN2Nquh8_2),.clk(gclk));
	jdff dff_B_e34QdL9G8_2(.din(w_dff_B_dbN2Nquh8_2),.dout(w_dff_B_e34QdL9G8_2),.clk(gclk));
	jdff dff_B_8cxraynF3_2(.din(w_dff_B_e34QdL9G8_2),.dout(w_dff_B_8cxraynF3_2),.clk(gclk));
	jdff dff_B_QbmdQVPc6_2(.din(w_dff_B_8cxraynF3_2),.dout(w_dff_B_QbmdQVPc6_2),.clk(gclk));
	jdff dff_B_ouMsuwRl7_2(.din(w_dff_B_QbmdQVPc6_2),.dout(w_dff_B_ouMsuwRl7_2),.clk(gclk));
	jdff dff_B_kHJAgOSm2_2(.din(w_dff_B_ouMsuwRl7_2),.dout(w_dff_B_kHJAgOSm2_2),.clk(gclk));
	jdff dff_B_g4zIW2PC4_1(.din(n1369),.dout(w_dff_B_g4zIW2PC4_1),.clk(gclk));
	jdff dff_B_AYwQZKXF4_2(.din(n1283),.dout(w_dff_B_AYwQZKXF4_2),.clk(gclk));
	jdff dff_B_xaBHkDI30_2(.din(w_dff_B_AYwQZKXF4_2),.dout(w_dff_B_xaBHkDI30_2),.clk(gclk));
	jdff dff_B_jeOGttWN8_2(.din(w_dff_B_xaBHkDI30_2),.dout(w_dff_B_jeOGttWN8_2),.clk(gclk));
	jdff dff_B_dHIOjesb1_2(.din(w_dff_B_jeOGttWN8_2),.dout(w_dff_B_dHIOjesb1_2),.clk(gclk));
	jdff dff_B_ygGQLR5W8_2(.din(w_dff_B_dHIOjesb1_2),.dout(w_dff_B_ygGQLR5W8_2),.clk(gclk));
	jdff dff_B_WynmUHo74_2(.din(w_dff_B_ygGQLR5W8_2),.dout(w_dff_B_WynmUHo74_2),.clk(gclk));
	jdff dff_B_7KpYrw5Z4_2(.din(w_dff_B_WynmUHo74_2),.dout(w_dff_B_7KpYrw5Z4_2),.clk(gclk));
	jdff dff_B_UVypv7lh7_2(.din(w_dff_B_7KpYrw5Z4_2),.dout(w_dff_B_UVypv7lh7_2),.clk(gclk));
	jdff dff_B_Ol5CSGFC4_2(.din(w_dff_B_UVypv7lh7_2),.dout(w_dff_B_Ol5CSGFC4_2),.clk(gclk));
	jdff dff_B_LUr1MXYX4_2(.din(w_dff_B_Ol5CSGFC4_2),.dout(w_dff_B_LUr1MXYX4_2),.clk(gclk));
	jdff dff_B_URSG0eUG4_2(.din(w_dff_B_LUr1MXYX4_2),.dout(w_dff_B_URSG0eUG4_2),.clk(gclk));
	jdff dff_B_7Jq3Nyio3_2(.din(w_dff_B_URSG0eUG4_2),.dout(w_dff_B_7Jq3Nyio3_2),.clk(gclk));
	jdff dff_B_k5Q1N5zD2_2(.din(w_dff_B_7Jq3Nyio3_2),.dout(w_dff_B_k5Q1N5zD2_2),.clk(gclk));
	jdff dff_B_OYPcVGBD1_2(.din(w_dff_B_k5Q1N5zD2_2),.dout(w_dff_B_OYPcVGBD1_2),.clk(gclk));
	jdff dff_B_qXnGpUXg3_2(.din(w_dff_B_OYPcVGBD1_2),.dout(w_dff_B_qXnGpUXg3_2),.clk(gclk));
	jdff dff_B_IPPbY5Lz0_2(.din(w_dff_B_qXnGpUXg3_2),.dout(w_dff_B_IPPbY5Lz0_2),.clk(gclk));
	jdff dff_B_1rwHte9Y5_2(.din(w_dff_B_IPPbY5Lz0_2),.dout(w_dff_B_1rwHte9Y5_2),.clk(gclk));
	jdff dff_B_Np6mHN2u7_2(.din(w_dff_B_1rwHte9Y5_2),.dout(w_dff_B_Np6mHN2u7_2),.clk(gclk));
	jdff dff_B_jslJltsU6_2(.din(w_dff_B_Np6mHN2u7_2),.dout(w_dff_B_jslJltsU6_2),.clk(gclk));
	jdff dff_B_prf6axQ95_2(.din(w_dff_B_jslJltsU6_2),.dout(w_dff_B_prf6axQ95_2),.clk(gclk));
	jdff dff_B_AoafReTF8_2(.din(w_dff_B_prf6axQ95_2),.dout(w_dff_B_AoafReTF8_2),.clk(gclk));
	jdff dff_B_ikuXHfzF8_2(.din(w_dff_B_AoafReTF8_2),.dout(w_dff_B_ikuXHfzF8_2),.clk(gclk));
	jdff dff_B_5rfyVuhh2_2(.din(w_dff_B_ikuXHfzF8_2),.dout(w_dff_B_5rfyVuhh2_2),.clk(gclk));
	jdff dff_B_bpkdk6rt2_2(.din(w_dff_B_5rfyVuhh2_2),.dout(w_dff_B_bpkdk6rt2_2),.clk(gclk));
	jdff dff_B_JJRZtfhZ9_2(.din(n1308),.dout(w_dff_B_JJRZtfhZ9_2),.clk(gclk));
	jdff dff_B_uZ7dF0Vi0_1(.din(n1284),.dout(w_dff_B_uZ7dF0Vi0_1),.clk(gclk));
	jdff dff_B_NOQlrnEz4_2(.din(n1193),.dout(w_dff_B_NOQlrnEz4_2),.clk(gclk));
	jdff dff_B_ivEGhaFx0_2(.din(w_dff_B_NOQlrnEz4_2),.dout(w_dff_B_ivEGhaFx0_2),.clk(gclk));
	jdff dff_B_GRbcs1Zq0_2(.din(w_dff_B_ivEGhaFx0_2),.dout(w_dff_B_GRbcs1Zq0_2),.clk(gclk));
	jdff dff_B_COEcUgMw3_2(.din(w_dff_B_GRbcs1Zq0_2),.dout(w_dff_B_COEcUgMw3_2),.clk(gclk));
	jdff dff_B_gJR63a2E9_2(.din(w_dff_B_COEcUgMw3_2),.dout(w_dff_B_gJR63a2E9_2),.clk(gclk));
	jdff dff_B_GG8SLyLe1_2(.din(w_dff_B_gJR63a2E9_2),.dout(w_dff_B_GG8SLyLe1_2),.clk(gclk));
	jdff dff_B_q7RnC2cO8_2(.din(w_dff_B_GG8SLyLe1_2),.dout(w_dff_B_q7RnC2cO8_2),.clk(gclk));
	jdff dff_B_qG4cZdZk7_2(.din(w_dff_B_q7RnC2cO8_2),.dout(w_dff_B_qG4cZdZk7_2),.clk(gclk));
	jdff dff_B_9R7Dz9iL9_2(.din(w_dff_B_qG4cZdZk7_2),.dout(w_dff_B_9R7Dz9iL9_2),.clk(gclk));
	jdff dff_B_vYsibJJa3_2(.din(w_dff_B_9R7Dz9iL9_2),.dout(w_dff_B_vYsibJJa3_2),.clk(gclk));
	jdff dff_B_eu0eYM0b0_2(.din(w_dff_B_vYsibJJa3_2),.dout(w_dff_B_eu0eYM0b0_2),.clk(gclk));
	jdff dff_B_8myywXnU8_2(.din(w_dff_B_eu0eYM0b0_2),.dout(w_dff_B_8myywXnU8_2),.clk(gclk));
	jdff dff_B_mOsJWtyd9_2(.din(w_dff_B_8myywXnU8_2),.dout(w_dff_B_mOsJWtyd9_2),.clk(gclk));
	jdff dff_B_bH83fHp69_2(.din(w_dff_B_mOsJWtyd9_2),.dout(w_dff_B_bH83fHp69_2),.clk(gclk));
	jdff dff_B_Fzu3Vkti7_2(.din(w_dff_B_bH83fHp69_2),.dout(w_dff_B_Fzu3Vkti7_2),.clk(gclk));
	jdff dff_B_zByCkGqu9_2(.din(w_dff_B_Fzu3Vkti7_2),.dout(w_dff_B_zByCkGqu9_2),.clk(gclk));
	jdff dff_B_Tcx4Y4gi5_2(.din(w_dff_B_zByCkGqu9_2),.dout(w_dff_B_Tcx4Y4gi5_2),.clk(gclk));
	jdff dff_B_JkexPaGh0_2(.din(w_dff_B_Tcx4Y4gi5_2),.dout(w_dff_B_JkexPaGh0_2),.clk(gclk));
	jdff dff_B_o4Lc9StX7_2(.din(w_dff_B_JkexPaGh0_2),.dout(w_dff_B_o4Lc9StX7_2),.clk(gclk));
	jdff dff_B_n4cbJXyH0_2(.din(w_dff_B_o4Lc9StX7_2),.dout(w_dff_B_n4cbJXyH0_2),.clk(gclk));
	jdff dff_B_eXoYxCfj8_2(.din(w_dff_B_n4cbJXyH0_2),.dout(w_dff_B_eXoYxCfj8_2),.clk(gclk));
	jdff dff_B_cMtgVFzy1_2(.din(n1217),.dout(w_dff_B_cMtgVFzy1_2),.clk(gclk));
	jdff dff_B_kK2ESgpI4_1(.din(n1194),.dout(w_dff_B_kK2ESgpI4_1),.clk(gclk));
	jdff dff_B_mHn6A1TG5_2(.din(n1089),.dout(w_dff_B_mHn6A1TG5_2),.clk(gclk));
	jdff dff_B_1vwQrPGr6_2(.din(w_dff_B_mHn6A1TG5_2),.dout(w_dff_B_1vwQrPGr6_2),.clk(gclk));
	jdff dff_B_qlumm9ey3_2(.din(w_dff_B_1vwQrPGr6_2),.dout(w_dff_B_qlumm9ey3_2),.clk(gclk));
	jdff dff_B_buLk5kNv1_2(.din(w_dff_B_qlumm9ey3_2),.dout(w_dff_B_buLk5kNv1_2),.clk(gclk));
	jdff dff_B_brqUSC524_2(.din(w_dff_B_buLk5kNv1_2),.dout(w_dff_B_brqUSC524_2),.clk(gclk));
	jdff dff_B_hmKDX2123_2(.din(w_dff_B_brqUSC524_2),.dout(w_dff_B_hmKDX2123_2),.clk(gclk));
	jdff dff_B_7a6b6YKa7_2(.din(w_dff_B_hmKDX2123_2),.dout(w_dff_B_7a6b6YKa7_2),.clk(gclk));
	jdff dff_B_KfiuQHT62_2(.din(w_dff_B_7a6b6YKa7_2),.dout(w_dff_B_KfiuQHT62_2),.clk(gclk));
	jdff dff_B_UX5K9AA02_2(.din(w_dff_B_KfiuQHT62_2),.dout(w_dff_B_UX5K9AA02_2),.clk(gclk));
	jdff dff_B_5xw0O59C9_2(.din(w_dff_B_UX5K9AA02_2),.dout(w_dff_B_5xw0O59C9_2),.clk(gclk));
	jdff dff_B_XaBd5fvY9_2(.din(w_dff_B_5xw0O59C9_2),.dout(w_dff_B_XaBd5fvY9_2),.clk(gclk));
	jdff dff_B_4Ajmh4Hz1_2(.din(w_dff_B_XaBd5fvY9_2),.dout(w_dff_B_4Ajmh4Hz1_2),.clk(gclk));
	jdff dff_B_GeeD8kzF0_2(.din(w_dff_B_4Ajmh4Hz1_2),.dout(w_dff_B_GeeD8kzF0_2),.clk(gclk));
	jdff dff_B_nEMqyReq9_2(.din(w_dff_B_GeeD8kzF0_2),.dout(w_dff_B_nEMqyReq9_2),.clk(gclk));
	jdff dff_B_jiPdFc5v4_2(.din(w_dff_B_nEMqyReq9_2),.dout(w_dff_B_jiPdFc5v4_2),.clk(gclk));
	jdff dff_B_7nqQFFA68_2(.din(w_dff_B_jiPdFc5v4_2),.dout(w_dff_B_7nqQFFA68_2),.clk(gclk));
	jdff dff_B_KYByy9QX1_2(.din(w_dff_B_7nqQFFA68_2),.dout(w_dff_B_KYByy9QX1_2),.clk(gclk));
	jdff dff_B_9eFiQyfl7_2(.din(w_dff_B_KYByy9QX1_2),.dout(w_dff_B_9eFiQyfl7_2),.clk(gclk));
	jdff dff_B_hZ2lehh50_2(.din(n1119),.dout(w_dff_B_hZ2lehh50_2),.clk(gclk));
	jdff dff_B_yk5YtVJ65_1(.din(n1090),.dout(w_dff_B_yk5YtVJ65_1),.clk(gclk));
	jdff dff_B_iFI0Jw5b8_2(.din(n991),.dout(w_dff_B_iFI0Jw5b8_2),.clk(gclk));
	jdff dff_B_Kv4pRacZ1_2(.din(w_dff_B_iFI0Jw5b8_2),.dout(w_dff_B_Kv4pRacZ1_2),.clk(gclk));
	jdff dff_B_bLaoZtQK9_2(.din(w_dff_B_Kv4pRacZ1_2),.dout(w_dff_B_bLaoZtQK9_2),.clk(gclk));
	jdff dff_B_Tk3tCumm3_2(.din(w_dff_B_bLaoZtQK9_2),.dout(w_dff_B_Tk3tCumm3_2),.clk(gclk));
	jdff dff_B_RIbb9lo81_2(.din(w_dff_B_Tk3tCumm3_2),.dout(w_dff_B_RIbb9lo81_2),.clk(gclk));
	jdff dff_B_fNkKkKfD6_2(.din(w_dff_B_RIbb9lo81_2),.dout(w_dff_B_fNkKkKfD6_2),.clk(gclk));
	jdff dff_B_zRxHkNoV3_2(.din(w_dff_B_fNkKkKfD6_2),.dout(w_dff_B_zRxHkNoV3_2),.clk(gclk));
	jdff dff_B_FNNAJWGs8_2(.din(w_dff_B_zRxHkNoV3_2),.dout(w_dff_B_FNNAJWGs8_2),.clk(gclk));
	jdff dff_B_uVu1qw1Q7_2(.din(w_dff_B_FNNAJWGs8_2),.dout(w_dff_B_uVu1qw1Q7_2),.clk(gclk));
	jdff dff_B_4lKUbKg04_2(.din(w_dff_B_uVu1qw1Q7_2),.dout(w_dff_B_4lKUbKg04_2),.clk(gclk));
	jdff dff_B_Tmmw64Qi2_2(.din(w_dff_B_4lKUbKg04_2),.dout(w_dff_B_Tmmw64Qi2_2),.clk(gclk));
	jdff dff_B_paeWwoNP1_2(.din(w_dff_B_Tmmw64Qi2_2),.dout(w_dff_B_paeWwoNP1_2),.clk(gclk));
	jdff dff_B_vV0WF0t53_2(.din(w_dff_B_paeWwoNP1_2),.dout(w_dff_B_vV0WF0t53_2),.clk(gclk));
	jdff dff_B_blbVkEUT9_2(.din(w_dff_B_vV0WF0t53_2),.dout(w_dff_B_blbVkEUT9_2),.clk(gclk));
	jdff dff_B_bflIGW7s7_2(.din(w_dff_B_blbVkEUT9_2),.dout(w_dff_B_bflIGW7s7_2),.clk(gclk));
	jdff dff_B_i5sM6kEZ8_2(.din(n1014),.dout(w_dff_B_i5sM6kEZ8_2),.clk(gclk));
	jdff dff_B_SB7dlvBc6_1(.din(n992),.dout(w_dff_B_SB7dlvBc6_1),.clk(gclk));
	jdff dff_B_Sklpz0k90_2(.din(n886),.dout(w_dff_B_Sklpz0k90_2),.clk(gclk));
	jdff dff_B_W4v6kaYt6_2(.din(w_dff_B_Sklpz0k90_2),.dout(w_dff_B_W4v6kaYt6_2),.clk(gclk));
	jdff dff_B_E09KK3E12_2(.din(w_dff_B_W4v6kaYt6_2),.dout(w_dff_B_E09KK3E12_2),.clk(gclk));
	jdff dff_B_lPn8Wxfn7_2(.din(w_dff_B_E09KK3E12_2),.dout(w_dff_B_lPn8Wxfn7_2),.clk(gclk));
	jdff dff_B_jxOpEzbY9_2(.din(w_dff_B_lPn8Wxfn7_2),.dout(w_dff_B_jxOpEzbY9_2),.clk(gclk));
	jdff dff_B_aE7bPIxk7_2(.din(w_dff_B_jxOpEzbY9_2),.dout(w_dff_B_aE7bPIxk7_2),.clk(gclk));
	jdff dff_B_kEUTOeIR7_2(.din(w_dff_B_aE7bPIxk7_2),.dout(w_dff_B_kEUTOeIR7_2),.clk(gclk));
	jdff dff_B_v4S3pv8l4_2(.din(w_dff_B_kEUTOeIR7_2),.dout(w_dff_B_v4S3pv8l4_2),.clk(gclk));
	jdff dff_B_EhWVhiBI6_2(.din(w_dff_B_v4S3pv8l4_2),.dout(w_dff_B_EhWVhiBI6_2),.clk(gclk));
	jdff dff_B_LIaiFfNQ6_2(.din(w_dff_B_EhWVhiBI6_2),.dout(w_dff_B_LIaiFfNQ6_2),.clk(gclk));
	jdff dff_B_uKetQiRC1_2(.din(w_dff_B_LIaiFfNQ6_2),.dout(w_dff_B_uKetQiRC1_2),.clk(gclk));
	jdff dff_B_yAr04H9W1_2(.din(w_dff_B_uKetQiRC1_2),.dout(w_dff_B_yAr04H9W1_2),.clk(gclk));
	jdff dff_B_QPpQGM361_2(.din(n909),.dout(w_dff_B_QPpQGM361_2),.clk(gclk));
	jdff dff_B_UNbWXrTi5_1(.din(n887),.dout(w_dff_B_UNbWXrTi5_1),.clk(gclk));
	jdff dff_B_C5q94eMr1_2(.din(n787),.dout(w_dff_B_C5q94eMr1_2),.clk(gclk));
	jdff dff_B_irBegRFQ8_2(.din(w_dff_B_C5q94eMr1_2),.dout(w_dff_B_irBegRFQ8_2),.clk(gclk));
	jdff dff_B_qwRekFJZ8_2(.din(w_dff_B_irBegRFQ8_2),.dout(w_dff_B_qwRekFJZ8_2),.clk(gclk));
	jdff dff_B_eb8W9Ta22_2(.din(w_dff_B_qwRekFJZ8_2),.dout(w_dff_B_eb8W9Ta22_2),.clk(gclk));
	jdff dff_B_l2EDcrU55_2(.din(w_dff_B_eb8W9Ta22_2),.dout(w_dff_B_l2EDcrU55_2),.clk(gclk));
	jdff dff_B_85hhOQCy4_2(.din(w_dff_B_l2EDcrU55_2),.dout(w_dff_B_85hhOQCy4_2),.clk(gclk));
	jdff dff_B_qsBeduna3_2(.din(w_dff_B_85hhOQCy4_2),.dout(w_dff_B_qsBeduna3_2),.clk(gclk));
	jdff dff_B_XGOvkdA66_2(.din(w_dff_B_qsBeduna3_2),.dout(w_dff_B_XGOvkdA66_2),.clk(gclk));
	jdff dff_B_4LFn6EgN7_2(.din(w_dff_B_XGOvkdA66_2),.dout(w_dff_B_4LFn6EgN7_2),.clk(gclk));
	jdff dff_B_6JFRe99A8_2(.din(n803),.dout(w_dff_B_6JFRe99A8_2),.clk(gclk));
	jdff dff_B_nzwKRckY6_2(.din(w_dff_B_6JFRe99A8_2),.dout(w_dff_B_nzwKRckY6_2),.clk(gclk));
	jdff dff_B_F6KKqp0I8_1(.din(n788),.dout(w_dff_B_F6KKqp0I8_1),.clk(gclk));
	jdff dff_B_208H61nz4_1(.din(w_dff_B_F6KKqp0I8_1),.dout(w_dff_B_208H61nz4_1),.clk(gclk));
	jdff dff_B_nfh0Anse2_1(.din(w_dff_B_208H61nz4_1),.dout(w_dff_B_nfh0Anse2_1),.clk(gclk));
	jdff dff_B_aGehSRJq9_1(.din(w_dff_B_nfh0Anse2_1),.dout(w_dff_B_aGehSRJq9_1),.clk(gclk));
	jdff dff_B_pK6cNqnY1_1(.din(w_dff_B_aGehSRJq9_1),.dout(w_dff_B_pK6cNqnY1_1),.clk(gclk));
	jdff dff_B_ycQziHRj5_1(.din(w_dff_B_pK6cNqnY1_1),.dout(w_dff_B_ycQziHRj5_1),.clk(gclk));
	jdff dff_B_ghKvLSbr0_0(.din(n703),.dout(w_dff_B_ghKvLSbr0_0),.clk(gclk));
	jdff dff_B_PYhFfXDa8_0(.din(w_dff_B_ghKvLSbr0_0),.dout(w_dff_B_PYhFfXDa8_0),.clk(gclk));
	jdff dff_A_Iuo8bC7C8_0(.dout(w_n702_0[0]),.din(w_dff_A_Iuo8bC7C8_0),.clk(gclk));
	jdff dff_A_UmkstwiT2_0(.dout(w_dff_A_Iuo8bC7C8_0),.din(w_dff_A_UmkstwiT2_0),.clk(gclk));
	jdff dff_A_LRlOYx2p2_0(.dout(w_dff_A_UmkstwiT2_0),.din(w_dff_A_LRlOYx2p2_0),.clk(gclk));
	jdff dff_B_j6eUikvB2_1(.din(n696),.dout(w_dff_B_j6eUikvB2_1),.clk(gclk));
	jdff dff_A_Ai6ny8Yz9_0(.dout(w_n607_0[0]),.din(w_dff_A_Ai6ny8Yz9_0),.clk(gclk));
	jdff dff_A_sWnJlBNP2_1(.dout(w_n607_0[1]),.din(w_dff_A_sWnJlBNP2_1),.clk(gclk));
	jdff dff_A_MUWNUiji3_1(.dout(w_dff_A_sWnJlBNP2_1),.din(w_dff_A_MUWNUiji3_1),.clk(gclk));
	jdff dff_A_DKGW4iE87_1(.dout(w_n694_0[1]),.din(w_dff_A_DKGW4iE87_1),.clk(gclk));
	jdff dff_A_ZtDRweVm1_1(.dout(w_dff_A_DKGW4iE87_1),.din(w_dff_A_ZtDRweVm1_1),.clk(gclk));
	jdff dff_A_3Pzw6UTd0_1(.dout(w_dff_A_ZtDRweVm1_1),.din(w_dff_A_3Pzw6UTd0_1),.clk(gclk));
	jdff dff_A_1d6TTFCT0_1(.dout(w_dff_A_3Pzw6UTd0_1),.din(w_dff_A_1d6TTFCT0_1),.clk(gclk));
	jdff dff_A_Ophfcl6M1_1(.dout(w_dff_A_1d6TTFCT0_1),.din(w_dff_A_Ophfcl6M1_1),.clk(gclk));
	jdff dff_A_bBP3iweD3_1(.dout(w_dff_A_Ophfcl6M1_1),.din(w_dff_A_bBP3iweD3_1),.clk(gclk));
	jdff dff_B_NiRQ0XUX0_1(.din(n1819),.dout(w_dff_B_NiRQ0XUX0_1),.clk(gclk));
	jdff dff_A_yvPCCEoS2_1(.dout(w_n1801_0[1]),.din(w_dff_A_yvPCCEoS2_1),.clk(gclk));
	jdff dff_B_CTe4bPiS3_1(.din(n1799),.dout(w_dff_B_CTe4bPiS3_1),.clk(gclk));
	jdff dff_B_4nIVDGd25_2(.din(n1770),.dout(w_dff_B_4nIVDGd25_2),.clk(gclk));
	jdff dff_B_QUfPRJAv6_2(.din(w_dff_B_4nIVDGd25_2),.dout(w_dff_B_QUfPRJAv6_2),.clk(gclk));
	jdff dff_B_quiluQjn1_2(.din(w_dff_B_QUfPRJAv6_2),.dout(w_dff_B_quiluQjn1_2),.clk(gclk));
	jdff dff_B_Lwpwq0Rs1_2(.din(w_dff_B_quiluQjn1_2),.dout(w_dff_B_Lwpwq0Rs1_2),.clk(gclk));
	jdff dff_B_go08VVGf3_2(.din(w_dff_B_Lwpwq0Rs1_2),.dout(w_dff_B_go08VVGf3_2),.clk(gclk));
	jdff dff_B_r02VsDN50_2(.din(w_dff_B_go08VVGf3_2),.dout(w_dff_B_r02VsDN50_2),.clk(gclk));
	jdff dff_B_AD3YtUdT3_2(.din(w_dff_B_r02VsDN50_2),.dout(w_dff_B_AD3YtUdT3_2),.clk(gclk));
	jdff dff_B_YidBgOfN1_2(.din(w_dff_B_AD3YtUdT3_2),.dout(w_dff_B_YidBgOfN1_2),.clk(gclk));
	jdff dff_B_Eh6HP9FU7_2(.din(w_dff_B_YidBgOfN1_2),.dout(w_dff_B_Eh6HP9FU7_2),.clk(gclk));
	jdff dff_B_aCqiNgN90_2(.din(w_dff_B_Eh6HP9FU7_2),.dout(w_dff_B_aCqiNgN90_2),.clk(gclk));
	jdff dff_B_O7uZei4a2_2(.din(w_dff_B_aCqiNgN90_2),.dout(w_dff_B_O7uZei4a2_2),.clk(gclk));
	jdff dff_B_KlPistLC0_2(.din(w_dff_B_O7uZei4a2_2),.dout(w_dff_B_KlPistLC0_2),.clk(gclk));
	jdff dff_B_5Uci0xnl4_2(.din(w_dff_B_KlPistLC0_2),.dout(w_dff_B_5Uci0xnl4_2),.clk(gclk));
	jdff dff_B_tsTNUwdT8_2(.din(w_dff_B_5Uci0xnl4_2),.dout(w_dff_B_tsTNUwdT8_2),.clk(gclk));
	jdff dff_B_IhEt0xlD8_2(.din(w_dff_B_tsTNUwdT8_2),.dout(w_dff_B_IhEt0xlD8_2),.clk(gclk));
	jdff dff_B_R5eYr6q44_2(.din(w_dff_B_IhEt0xlD8_2),.dout(w_dff_B_R5eYr6q44_2),.clk(gclk));
	jdff dff_B_HF8XaDwQ5_2(.din(w_dff_B_R5eYr6q44_2),.dout(w_dff_B_HF8XaDwQ5_2),.clk(gclk));
	jdff dff_B_eCZCoMfL5_2(.din(w_dff_B_HF8XaDwQ5_2),.dout(w_dff_B_eCZCoMfL5_2),.clk(gclk));
	jdff dff_B_65c9tFPw6_2(.din(w_dff_B_eCZCoMfL5_2),.dout(w_dff_B_65c9tFPw6_2),.clk(gclk));
	jdff dff_B_c7nY5kDD2_2(.din(w_dff_B_65c9tFPw6_2),.dout(w_dff_B_c7nY5kDD2_2),.clk(gclk));
	jdff dff_B_aUv76SM82_2(.din(w_dff_B_c7nY5kDD2_2),.dout(w_dff_B_aUv76SM82_2),.clk(gclk));
	jdff dff_B_NjvE3s542_2(.din(w_dff_B_aUv76SM82_2),.dout(w_dff_B_NjvE3s542_2),.clk(gclk));
	jdff dff_B_BeEC1Zg71_2(.din(w_dff_B_NjvE3s542_2),.dout(w_dff_B_BeEC1Zg71_2),.clk(gclk));
	jdff dff_B_8o94F5ir9_2(.din(w_dff_B_BeEC1Zg71_2),.dout(w_dff_B_8o94F5ir9_2),.clk(gclk));
	jdff dff_B_6jffrsIL3_2(.din(w_dff_B_8o94F5ir9_2),.dout(w_dff_B_6jffrsIL3_2),.clk(gclk));
	jdff dff_B_obcOtCP87_2(.din(w_dff_B_6jffrsIL3_2),.dout(w_dff_B_obcOtCP87_2),.clk(gclk));
	jdff dff_B_hwvu0FLI9_2(.din(w_dff_B_obcOtCP87_2),.dout(w_dff_B_hwvu0FLI9_2),.clk(gclk));
	jdff dff_B_pbZRBvRS6_2(.din(w_dff_B_hwvu0FLI9_2),.dout(w_dff_B_pbZRBvRS6_2),.clk(gclk));
	jdff dff_B_SPRwxoXi1_2(.din(w_dff_B_pbZRBvRS6_2),.dout(w_dff_B_SPRwxoXi1_2),.clk(gclk));
	jdff dff_B_W5tD9vhU1_2(.din(w_dff_B_SPRwxoXi1_2),.dout(w_dff_B_W5tD9vhU1_2),.clk(gclk));
	jdff dff_B_gKsJZiiL0_2(.din(w_dff_B_W5tD9vhU1_2),.dout(w_dff_B_gKsJZiiL0_2),.clk(gclk));
	jdff dff_B_kiKmBUMo3_2(.din(w_dff_B_gKsJZiiL0_2),.dout(w_dff_B_kiKmBUMo3_2),.clk(gclk));
	jdff dff_B_tROCr7Qy1_2(.din(w_dff_B_kiKmBUMo3_2),.dout(w_dff_B_tROCr7Qy1_2),.clk(gclk));
	jdff dff_B_9DKHQsVB6_2(.din(w_dff_B_tROCr7Qy1_2),.dout(w_dff_B_9DKHQsVB6_2),.clk(gclk));
	jdff dff_B_lvIOlS5B8_2(.din(w_dff_B_9DKHQsVB6_2),.dout(w_dff_B_lvIOlS5B8_2),.clk(gclk));
	jdff dff_B_aULnmtzK4_2(.din(w_dff_B_lvIOlS5B8_2),.dout(w_dff_B_aULnmtzK4_2),.clk(gclk));
	jdff dff_B_gICv0iZF9_2(.din(w_dff_B_aULnmtzK4_2),.dout(w_dff_B_gICv0iZF9_2),.clk(gclk));
	jdff dff_B_qNV9so0P2_2(.din(w_dff_B_gICv0iZF9_2),.dout(w_dff_B_qNV9so0P2_2),.clk(gclk));
	jdff dff_B_ymtchohA0_2(.din(w_dff_B_qNV9so0P2_2),.dout(w_dff_B_ymtchohA0_2),.clk(gclk));
	jdff dff_B_hzjYATWG7_2(.din(w_dff_B_ymtchohA0_2),.dout(w_dff_B_hzjYATWG7_2),.clk(gclk));
	jdff dff_B_mX3K5PLX2_2(.din(w_dff_B_hzjYATWG7_2),.dout(w_dff_B_mX3K5PLX2_2),.clk(gclk));
	jdff dff_B_CxOv5dCV8_2(.din(w_dff_B_mX3K5PLX2_2),.dout(w_dff_B_CxOv5dCV8_2),.clk(gclk));
	jdff dff_B_N9peuzqX8_2(.din(w_dff_B_CxOv5dCV8_2),.dout(w_dff_B_N9peuzqX8_2),.clk(gclk));
	jdff dff_B_ia8C6Jxo2_2(.din(w_dff_B_N9peuzqX8_2),.dout(w_dff_B_ia8C6Jxo2_2),.clk(gclk));
	jdff dff_B_4h1mvUyI5_2(.din(w_dff_B_ia8C6Jxo2_2),.dout(w_dff_B_4h1mvUyI5_2),.clk(gclk));
	jdff dff_B_dFVoXNyH6_2(.din(w_dff_B_4h1mvUyI5_2),.dout(w_dff_B_dFVoXNyH6_2),.clk(gclk));
	jdff dff_B_R2Uyxj707_2(.din(w_dff_B_dFVoXNyH6_2),.dout(w_dff_B_R2Uyxj707_2),.clk(gclk));
	jdff dff_B_t6OTknWa2_2(.din(w_dff_B_R2Uyxj707_2),.dout(w_dff_B_t6OTknWa2_2),.clk(gclk));
	jdff dff_B_KJSXHFsq9_2(.din(w_dff_B_t6OTknWa2_2),.dout(w_dff_B_KJSXHFsq9_2),.clk(gclk));
	jdff dff_B_ZaTVUDFY8_2(.din(w_dff_B_KJSXHFsq9_2),.dout(w_dff_B_ZaTVUDFY8_2),.clk(gclk));
	jdff dff_B_NrKguckG2_2(.din(w_dff_B_ZaTVUDFY8_2),.dout(w_dff_B_NrKguckG2_2),.clk(gclk));
	jdff dff_B_slftNcig9_2(.din(w_dff_B_NrKguckG2_2),.dout(w_dff_B_slftNcig9_2),.clk(gclk));
	jdff dff_B_Yzc9RcZh4_2(.din(w_dff_B_slftNcig9_2),.dout(w_dff_B_Yzc9RcZh4_2),.clk(gclk));
	jdff dff_B_2XG2nvNA2_2(.din(n1773),.dout(w_dff_B_2XG2nvNA2_2),.clk(gclk));
	jdff dff_B_b90Z7vXn8_1(.din(n1771),.dout(w_dff_B_b90Z7vXn8_1),.clk(gclk));
	jdff dff_B_KXCtdLDY9_2(.din(n1735),.dout(w_dff_B_KXCtdLDY9_2),.clk(gclk));
	jdff dff_B_ZPMbSx675_2(.din(w_dff_B_KXCtdLDY9_2),.dout(w_dff_B_ZPMbSx675_2),.clk(gclk));
	jdff dff_B_oabqylBl9_2(.din(w_dff_B_ZPMbSx675_2),.dout(w_dff_B_oabqylBl9_2),.clk(gclk));
	jdff dff_B_A0AcWmW61_2(.din(w_dff_B_oabqylBl9_2),.dout(w_dff_B_A0AcWmW61_2),.clk(gclk));
	jdff dff_B_3pAKkzOx4_2(.din(w_dff_B_A0AcWmW61_2),.dout(w_dff_B_3pAKkzOx4_2),.clk(gclk));
	jdff dff_B_qUoeQIKv6_2(.din(w_dff_B_3pAKkzOx4_2),.dout(w_dff_B_qUoeQIKv6_2),.clk(gclk));
	jdff dff_B_s4PK1PJk0_2(.din(w_dff_B_qUoeQIKv6_2),.dout(w_dff_B_s4PK1PJk0_2),.clk(gclk));
	jdff dff_B_5qVeG1Dk9_2(.din(w_dff_B_s4PK1PJk0_2),.dout(w_dff_B_5qVeG1Dk9_2),.clk(gclk));
	jdff dff_B_ZdHKM6qD3_2(.din(w_dff_B_5qVeG1Dk9_2),.dout(w_dff_B_ZdHKM6qD3_2),.clk(gclk));
	jdff dff_B_i9an8hkh6_2(.din(w_dff_B_ZdHKM6qD3_2),.dout(w_dff_B_i9an8hkh6_2),.clk(gclk));
	jdff dff_B_5sjCzV3N6_2(.din(w_dff_B_i9an8hkh6_2),.dout(w_dff_B_5sjCzV3N6_2),.clk(gclk));
	jdff dff_B_gPof9vDJ0_2(.din(w_dff_B_5sjCzV3N6_2),.dout(w_dff_B_gPof9vDJ0_2),.clk(gclk));
	jdff dff_B_Aq0lgHlt0_2(.din(w_dff_B_gPof9vDJ0_2),.dout(w_dff_B_Aq0lgHlt0_2),.clk(gclk));
	jdff dff_B_Tres6fIH3_2(.din(w_dff_B_Aq0lgHlt0_2),.dout(w_dff_B_Tres6fIH3_2),.clk(gclk));
	jdff dff_B_b7EvgEKd2_2(.din(w_dff_B_Tres6fIH3_2),.dout(w_dff_B_b7EvgEKd2_2),.clk(gclk));
	jdff dff_B_9vI8bOzX1_2(.din(w_dff_B_b7EvgEKd2_2),.dout(w_dff_B_9vI8bOzX1_2),.clk(gclk));
	jdff dff_B_2RDqrGKY7_2(.din(w_dff_B_9vI8bOzX1_2),.dout(w_dff_B_2RDqrGKY7_2),.clk(gclk));
	jdff dff_B_5TwqCLW80_2(.din(w_dff_B_2RDqrGKY7_2),.dout(w_dff_B_5TwqCLW80_2),.clk(gclk));
	jdff dff_B_woQAuOM94_2(.din(w_dff_B_5TwqCLW80_2),.dout(w_dff_B_woQAuOM94_2),.clk(gclk));
	jdff dff_B_f2G8Qthw2_2(.din(w_dff_B_woQAuOM94_2),.dout(w_dff_B_f2G8Qthw2_2),.clk(gclk));
	jdff dff_B_PG6hOt2x3_2(.din(w_dff_B_f2G8Qthw2_2),.dout(w_dff_B_PG6hOt2x3_2),.clk(gclk));
	jdff dff_B_m0ipGKvO8_2(.din(w_dff_B_PG6hOt2x3_2),.dout(w_dff_B_m0ipGKvO8_2),.clk(gclk));
	jdff dff_B_lUtFYRnr3_2(.din(w_dff_B_m0ipGKvO8_2),.dout(w_dff_B_lUtFYRnr3_2),.clk(gclk));
	jdff dff_B_KebbMlSm5_2(.din(w_dff_B_lUtFYRnr3_2),.dout(w_dff_B_KebbMlSm5_2),.clk(gclk));
	jdff dff_B_oNxnqqyu5_2(.din(w_dff_B_KebbMlSm5_2),.dout(w_dff_B_oNxnqqyu5_2),.clk(gclk));
	jdff dff_B_1l8dkLAa2_2(.din(w_dff_B_oNxnqqyu5_2),.dout(w_dff_B_1l8dkLAa2_2),.clk(gclk));
	jdff dff_B_nCz172J18_2(.din(w_dff_B_1l8dkLAa2_2),.dout(w_dff_B_nCz172J18_2),.clk(gclk));
	jdff dff_B_AxL68lvD9_2(.din(w_dff_B_nCz172J18_2),.dout(w_dff_B_AxL68lvD9_2),.clk(gclk));
	jdff dff_B_f5mxh1ET3_2(.din(w_dff_B_AxL68lvD9_2),.dout(w_dff_B_f5mxh1ET3_2),.clk(gclk));
	jdff dff_B_o20zr0du2_2(.din(w_dff_B_f5mxh1ET3_2),.dout(w_dff_B_o20zr0du2_2),.clk(gclk));
	jdff dff_B_ZeIq7Lxt3_2(.din(w_dff_B_o20zr0du2_2),.dout(w_dff_B_ZeIq7Lxt3_2),.clk(gclk));
	jdff dff_B_3OKcia3V4_2(.din(w_dff_B_ZeIq7Lxt3_2),.dout(w_dff_B_3OKcia3V4_2),.clk(gclk));
	jdff dff_B_x1Y6veYi8_2(.din(w_dff_B_3OKcia3V4_2),.dout(w_dff_B_x1Y6veYi8_2),.clk(gclk));
	jdff dff_B_mrBya4Ue2_2(.din(w_dff_B_x1Y6veYi8_2),.dout(w_dff_B_mrBya4Ue2_2),.clk(gclk));
	jdff dff_B_1rR9e1Ob7_2(.din(w_dff_B_mrBya4Ue2_2),.dout(w_dff_B_1rR9e1Ob7_2),.clk(gclk));
	jdff dff_B_VgSSCo7L6_2(.din(w_dff_B_1rR9e1Ob7_2),.dout(w_dff_B_VgSSCo7L6_2),.clk(gclk));
	jdff dff_B_4Inb6VYI6_2(.din(w_dff_B_VgSSCo7L6_2),.dout(w_dff_B_4Inb6VYI6_2),.clk(gclk));
	jdff dff_B_iFlcSjGb2_2(.din(w_dff_B_4Inb6VYI6_2),.dout(w_dff_B_iFlcSjGb2_2),.clk(gclk));
	jdff dff_B_Uc3LKQd95_2(.din(w_dff_B_iFlcSjGb2_2),.dout(w_dff_B_Uc3LKQd95_2),.clk(gclk));
	jdff dff_B_7uSCX6Ej2_2(.din(w_dff_B_Uc3LKQd95_2),.dout(w_dff_B_7uSCX6Ej2_2),.clk(gclk));
	jdff dff_B_VTXlkmTV2_2(.din(w_dff_B_7uSCX6Ej2_2),.dout(w_dff_B_VTXlkmTV2_2),.clk(gclk));
	jdff dff_B_ta4tm3Ee2_2(.din(w_dff_B_VTXlkmTV2_2),.dout(w_dff_B_ta4tm3Ee2_2),.clk(gclk));
	jdff dff_B_ETpWHW4o5_2(.din(w_dff_B_ta4tm3Ee2_2),.dout(w_dff_B_ETpWHW4o5_2),.clk(gclk));
	jdff dff_B_2PiFW1EC3_2(.din(w_dff_B_ETpWHW4o5_2),.dout(w_dff_B_2PiFW1EC3_2),.clk(gclk));
	jdff dff_B_hXelHWkr4_2(.din(w_dff_B_2PiFW1EC3_2),.dout(w_dff_B_hXelHWkr4_2),.clk(gclk));
	jdff dff_B_1YHFoZHD0_2(.din(w_dff_B_hXelHWkr4_2),.dout(w_dff_B_1YHFoZHD0_2),.clk(gclk));
	jdff dff_B_xCbISSsD1_2(.din(w_dff_B_1YHFoZHD0_2),.dout(w_dff_B_xCbISSsD1_2),.clk(gclk));
	jdff dff_B_MIp6UnZx6_2(.din(w_dff_B_xCbISSsD1_2),.dout(w_dff_B_MIp6UnZx6_2),.clk(gclk));
	jdff dff_B_09FlSBNU8_2(.din(w_dff_B_MIp6UnZx6_2),.dout(w_dff_B_09FlSBNU8_2),.clk(gclk));
	jdff dff_B_Hto6pA017_2(.din(n1738),.dout(w_dff_B_Hto6pA017_2),.clk(gclk));
	jdff dff_B_GBFhlqJt1_1(.din(n1736),.dout(w_dff_B_GBFhlqJt1_1),.clk(gclk));
	jdff dff_B_4UDLIoq55_2(.din(n1694),.dout(w_dff_B_4UDLIoq55_2),.clk(gclk));
	jdff dff_B_6W6ZzYxM6_2(.din(w_dff_B_4UDLIoq55_2),.dout(w_dff_B_6W6ZzYxM6_2),.clk(gclk));
	jdff dff_B_XH1xguaG7_2(.din(w_dff_B_6W6ZzYxM6_2),.dout(w_dff_B_XH1xguaG7_2),.clk(gclk));
	jdff dff_B_wEzATMU09_2(.din(w_dff_B_XH1xguaG7_2),.dout(w_dff_B_wEzATMU09_2),.clk(gclk));
	jdff dff_B_nndZOcyO3_2(.din(w_dff_B_wEzATMU09_2),.dout(w_dff_B_nndZOcyO3_2),.clk(gclk));
	jdff dff_B_DFfnGP5J9_2(.din(w_dff_B_nndZOcyO3_2),.dout(w_dff_B_DFfnGP5J9_2),.clk(gclk));
	jdff dff_B_BLdlEHzf0_2(.din(w_dff_B_DFfnGP5J9_2),.dout(w_dff_B_BLdlEHzf0_2),.clk(gclk));
	jdff dff_B_mh1EG16L9_2(.din(w_dff_B_BLdlEHzf0_2),.dout(w_dff_B_mh1EG16L9_2),.clk(gclk));
	jdff dff_B_k5sQI2H94_2(.din(w_dff_B_mh1EG16L9_2),.dout(w_dff_B_k5sQI2H94_2),.clk(gclk));
	jdff dff_B_gIS3kEDz2_2(.din(w_dff_B_k5sQI2H94_2),.dout(w_dff_B_gIS3kEDz2_2),.clk(gclk));
	jdff dff_B_WuTXHVMW8_2(.din(w_dff_B_gIS3kEDz2_2),.dout(w_dff_B_WuTXHVMW8_2),.clk(gclk));
	jdff dff_B_tVhIJKlQ7_2(.din(w_dff_B_WuTXHVMW8_2),.dout(w_dff_B_tVhIJKlQ7_2),.clk(gclk));
	jdff dff_B_cWNrJTbM5_2(.din(w_dff_B_tVhIJKlQ7_2),.dout(w_dff_B_cWNrJTbM5_2),.clk(gclk));
	jdff dff_B_kbAsr9uR3_2(.din(w_dff_B_cWNrJTbM5_2),.dout(w_dff_B_kbAsr9uR3_2),.clk(gclk));
	jdff dff_B_NipPy7uN2_2(.din(w_dff_B_kbAsr9uR3_2),.dout(w_dff_B_NipPy7uN2_2),.clk(gclk));
	jdff dff_B_eiXdaOvx5_2(.din(w_dff_B_NipPy7uN2_2),.dout(w_dff_B_eiXdaOvx5_2),.clk(gclk));
	jdff dff_B_vLi2tK112_2(.din(w_dff_B_eiXdaOvx5_2),.dout(w_dff_B_vLi2tK112_2),.clk(gclk));
	jdff dff_B_ksl1FEt55_2(.din(w_dff_B_vLi2tK112_2),.dout(w_dff_B_ksl1FEt55_2),.clk(gclk));
	jdff dff_B_9juIz4GK3_2(.din(w_dff_B_ksl1FEt55_2),.dout(w_dff_B_9juIz4GK3_2),.clk(gclk));
	jdff dff_B_87lSFLpn4_2(.din(w_dff_B_9juIz4GK3_2),.dout(w_dff_B_87lSFLpn4_2),.clk(gclk));
	jdff dff_B_uX0s9TIR7_2(.din(w_dff_B_87lSFLpn4_2),.dout(w_dff_B_uX0s9TIR7_2),.clk(gclk));
	jdff dff_B_K6W7jNUc1_2(.din(w_dff_B_uX0s9TIR7_2),.dout(w_dff_B_K6W7jNUc1_2),.clk(gclk));
	jdff dff_B_xBMYqHLV8_2(.din(w_dff_B_K6W7jNUc1_2),.dout(w_dff_B_xBMYqHLV8_2),.clk(gclk));
	jdff dff_B_D1VcgLeh7_2(.din(w_dff_B_xBMYqHLV8_2),.dout(w_dff_B_D1VcgLeh7_2),.clk(gclk));
	jdff dff_B_Kc3U1Dgf5_2(.din(w_dff_B_D1VcgLeh7_2),.dout(w_dff_B_Kc3U1Dgf5_2),.clk(gclk));
	jdff dff_B_fS7xFAsa4_2(.din(w_dff_B_Kc3U1Dgf5_2),.dout(w_dff_B_fS7xFAsa4_2),.clk(gclk));
	jdff dff_B_hJgONq219_2(.din(w_dff_B_fS7xFAsa4_2),.dout(w_dff_B_hJgONq219_2),.clk(gclk));
	jdff dff_B_7HZ5Uspp5_2(.din(w_dff_B_hJgONq219_2),.dout(w_dff_B_7HZ5Uspp5_2),.clk(gclk));
	jdff dff_B_lRMMQxUd3_2(.din(w_dff_B_7HZ5Uspp5_2),.dout(w_dff_B_lRMMQxUd3_2),.clk(gclk));
	jdff dff_B_NUYPluOB9_2(.din(w_dff_B_lRMMQxUd3_2),.dout(w_dff_B_NUYPluOB9_2),.clk(gclk));
	jdff dff_B_M4hO2AI63_2(.din(w_dff_B_NUYPluOB9_2),.dout(w_dff_B_M4hO2AI63_2),.clk(gclk));
	jdff dff_B_E38pZlid0_2(.din(w_dff_B_M4hO2AI63_2),.dout(w_dff_B_E38pZlid0_2),.clk(gclk));
	jdff dff_B_v3RGeEgj5_2(.din(w_dff_B_E38pZlid0_2),.dout(w_dff_B_v3RGeEgj5_2),.clk(gclk));
	jdff dff_B_0IskqFG09_2(.din(w_dff_B_v3RGeEgj5_2),.dout(w_dff_B_0IskqFG09_2),.clk(gclk));
	jdff dff_B_s5JImO5R6_2(.din(w_dff_B_0IskqFG09_2),.dout(w_dff_B_s5JImO5R6_2),.clk(gclk));
	jdff dff_B_IFDitTZ19_2(.din(w_dff_B_s5JImO5R6_2),.dout(w_dff_B_IFDitTZ19_2),.clk(gclk));
	jdff dff_B_zqvwS3iM5_2(.din(w_dff_B_IFDitTZ19_2),.dout(w_dff_B_zqvwS3iM5_2),.clk(gclk));
	jdff dff_B_i1aIOw928_2(.din(w_dff_B_zqvwS3iM5_2),.dout(w_dff_B_i1aIOw928_2),.clk(gclk));
	jdff dff_B_Gdc5TsG35_2(.din(w_dff_B_i1aIOw928_2),.dout(w_dff_B_Gdc5TsG35_2),.clk(gclk));
	jdff dff_B_CqHiyiZY7_2(.din(w_dff_B_Gdc5TsG35_2),.dout(w_dff_B_CqHiyiZY7_2),.clk(gclk));
	jdff dff_B_LfEiPaCA7_2(.din(w_dff_B_CqHiyiZY7_2),.dout(w_dff_B_LfEiPaCA7_2),.clk(gclk));
	jdff dff_B_Gpze2ohh9_2(.din(w_dff_B_LfEiPaCA7_2),.dout(w_dff_B_Gpze2ohh9_2),.clk(gclk));
	jdff dff_B_4OrxLSvx8_2(.din(w_dff_B_Gpze2ohh9_2),.dout(w_dff_B_4OrxLSvx8_2),.clk(gclk));
	jdff dff_B_lb9kz3zq0_2(.din(w_dff_B_4OrxLSvx8_2),.dout(w_dff_B_lb9kz3zq0_2),.clk(gclk));
	jdff dff_B_icbpygs14_2(.din(w_dff_B_lb9kz3zq0_2),.dout(w_dff_B_icbpygs14_2),.clk(gclk));
	jdff dff_B_CWjW9Ljq8_2(.din(n1697),.dout(w_dff_B_CWjW9Ljq8_2),.clk(gclk));
	jdff dff_B_IVGV1hWr7_1(.din(n1695),.dout(w_dff_B_IVGV1hWr7_1),.clk(gclk));
	jdff dff_B_273ZWcL18_2(.din(n1643),.dout(w_dff_B_273ZWcL18_2),.clk(gclk));
	jdff dff_B_gLWEgUOH6_2(.din(w_dff_B_273ZWcL18_2),.dout(w_dff_B_gLWEgUOH6_2),.clk(gclk));
	jdff dff_B_oco2Xphf9_2(.din(w_dff_B_gLWEgUOH6_2),.dout(w_dff_B_oco2Xphf9_2),.clk(gclk));
	jdff dff_B_xZiyinH49_2(.din(w_dff_B_oco2Xphf9_2),.dout(w_dff_B_xZiyinH49_2),.clk(gclk));
	jdff dff_B_QtSkH6op7_2(.din(w_dff_B_xZiyinH49_2),.dout(w_dff_B_QtSkH6op7_2),.clk(gclk));
	jdff dff_B_n6Yh4seq7_2(.din(w_dff_B_QtSkH6op7_2),.dout(w_dff_B_n6Yh4seq7_2),.clk(gclk));
	jdff dff_B_7MxdhzbH0_2(.din(w_dff_B_n6Yh4seq7_2),.dout(w_dff_B_7MxdhzbH0_2),.clk(gclk));
	jdff dff_B_g5a79xU07_2(.din(w_dff_B_7MxdhzbH0_2),.dout(w_dff_B_g5a79xU07_2),.clk(gclk));
	jdff dff_B_W0GnBM7v9_2(.din(w_dff_B_g5a79xU07_2),.dout(w_dff_B_W0GnBM7v9_2),.clk(gclk));
	jdff dff_B_ApJ9mZ5m1_2(.din(w_dff_B_W0GnBM7v9_2),.dout(w_dff_B_ApJ9mZ5m1_2),.clk(gclk));
	jdff dff_B_BeobT1ZP5_2(.din(w_dff_B_ApJ9mZ5m1_2),.dout(w_dff_B_BeobT1ZP5_2),.clk(gclk));
	jdff dff_B_vW33an8Q9_2(.din(w_dff_B_BeobT1ZP5_2),.dout(w_dff_B_vW33an8Q9_2),.clk(gclk));
	jdff dff_B_QOIXrkTW8_2(.din(w_dff_B_vW33an8Q9_2),.dout(w_dff_B_QOIXrkTW8_2),.clk(gclk));
	jdff dff_B_NtK0a0m25_2(.din(w_dff_B_QOIXrkTW8_2),.dout(w_dff_B_NtK0a0m25_2),.clk(gclk));
	jdff dff_B_VCgPFZcq9_2(.din(w_dff_B_NtK0a0m25_2),.dout(w_dff_B_VCgPFZcq9_2),.clk(gclk));
	jdff dff_B_g26D1fnS9_2(.din(w_dff_B_VCgPFZcq9_2),.dout(w_dff_B_g26D1fnS9_2),.clk(gclk));
	jdff dff_B_cUQTFXfz3_2(.din(w_dff_B_g26D1fnS9_2),.dout(w_dff_B_cUQTFXfz3_2),.clk(gclk));
	jdff dff_B_fc7bjt8A9_2(.din(w_dff_B_cUQTFXfz3_2),.dout(w_dff_B_fc7bjt8A9_2),.clk(gclk));
	jdff dff_B_QTttfCQz4_2(.din(w_dff_B_fc7bjt8A9_2),.dout(w_dff_B_QTttfCQz4_2),.clk(gclk));
	jdff dff_B_dN2AR35P0_2(.din(w_dff_B_QTttfCQz4_2),.dout(w_dff_B_dN2AR35P0_2),.clk(gclk));
	jdff dff_B_TOHUYWdZ1_2(.din(w_dff_B_dN2AR35P0_2),.dout(w_dff_B_TOHUYWdZ1_2),.clk(gclk));
	jdff dff_B_q6qrVm9B0_2(.din(w_dff_B_TOHUYWdZ1_2),.dout(w_dff_B_q6qrVm9B0_2),.clk(gclk));
	jdff dff_B_OihMuvS32_2(.din(w_dff_B_q6qrVm9B0_2),.dout(w_dff_B_OihMuvS32_2),.clk(gclk));
	jdff dff_B_ndJRK4Ir6_2(.din(w_dff_B_OihMuvS32_2),.dout(w_dff_B_ndJRK4Ir6_2),.clk(gclk));
	jdff dff_B_if7qqmyu3_2(.din(w_dff_B_ndJRK4Ir6_2),.dout(w_dff_B_if7qqmyu3_2),.clk(gclk));
	jdff dff_B_pksl8QHj3_2(.din(w_dff_B_if7qqmyu3_2),.dout(w_dff_B_pksl8QHj3_2),.clk(gclk));
	jdff dff_B_i6IMqcDR0_2(.din(w_dff_B_pksl8QHj3_2),.dout(w_dff_B_i6IMqcDR0_2),.clk(gclk));
	jdff dff_B_k2vqLwNI5_2(.din(w_dff_B_i6IMqcDR0_2),.dout(w_dff_B_k2vqLwNI5_2),.clk(gclk));
	jdff dff_B_JnDYOcxb6_2(.din(w_dff_B_k2vqLwNI5_2),.dout(w_dff_B_JnDYOcxb6_2),.clk(gclk));
	jdff dff_B_u2SVdbn26_2(.din(w_dff_B_JnDYOcxb6_2),.dout(w_dff_B_u2SVdbn26_2),.clk(gclk));
	jdff dff_B_uyYZNR952_2(.din(w_dff_B_u2SVdbn26_2),.dout(w_dff_B_uyYZNR952_2),.clk(gclk));
	jdff dff_B_CaS43xin0_2(.din(w_dff_B_uyYZNR952_2),.dout(w_dff_B_CaS43xin0_2),.clk(gclk));
	jdff dff_B_iTqTfpYg1_2(.din(w_dff_B_CaS43xin0_2),.dout(w_dff_B_iTqTfpYg1_2),.clk(gclk));
	jdff dff_B_JzbMjfsx6_2(.din(w_dff_B_iTqTfpYg1_2),.dout(w_dff_B_JzbMjfsx6_2),.clk(gclk));
	jdff dff_B_Qe7aWXeH0_2(.din(w_dff_B_JzbMjfsx6_2),.dout(w_dff_B_Qe7aWXeH0_2),.clk(gclk));
	jdff dff_B_045T1oLg8_2(.din(w_dff_B_Qe7aWXeH0_2),.dout(w_dff_B_045T1oLg8_2),.clk(gclk));
	jdff dff_B_URcjHMWH7_2(.din(w_dff_B_045T1oLg8_2),.dout(w_dff_B_URcjHMWH7_2),.clk(gclk));
	jdff dff_B_hyrv6va34_2(.din(w_dff_B_URcjHMWH7_2),.dout(w_dff_B_hyrv6va34_2),.clk(gclk));
	jdff dff_B_dnZ792338_2(.din(w_dff_B_hyrv6va34_2),.dout(w_dff_B_dnZ792338_2),.clk(gclk));
	jdff dff_B_mFUXl2Vr0_2(.din(w_dff_B_dnZ792338_2),.dout(w_dff_B_mFUXl2Vr0_2),.clk(gclk));
	jdff dff_B_49g8mCix4_2(.din(w_dff_B_mFUXl2Vr0_2),.dout(w_dff_B_49g8mCix4_2),.clk(gclk));
	jdff dff_B_D0oz23es3_2(.din(n1646),.dout(w_dff_B_D0oz23es3_2),.clk(gclk));
	jdff dff_B_BceJ9HAg2_1(.din(n1644),.dout(w_dff_B_BceJ9HAg2_1),.clk(gclk));
	jdff dff_B_XU1ib5pi4_2(.din(n1586),.dout(w_dff_B_XU1ib5pi4_2),.clk(gclk));
	jdff dff_B_4Hf9CiEg8_2(.din(w_dff_B_XU1ib5pi4_2),.dout(w_dff_B_4Hf9CiEg8_2),.clk(gclk));
	jdff dff_B_PQbTCk5t0_2(.din(w_dff_B_4Hf9CiEg8_2),.dout(w_dff_B_PQbTCk5t0_2),.clk(gclk));
	jdff dff_B_JwZJKHav3_2(.din(w_dff_B_PQbTCk5t0_2),.dout(w_dff_B_JwZJKHav3_2),.clk(gclk));
	jdff dff_B_IU07JJ6l8_2(.din(w_dff_B_JwZJKHav3_2),.dout(w_dff_B_IU07JJ6l8_2),.clk(gclk));
	jdff dff_B_iQyohNPb5_2(.din(w_dff_B_IU07JJ6l8_2),.dout(w_dff_B_iQyohNPb5_2),.clk(gclk));
	jdff dff_B_2syLQrTk8_2(.din(w_dff_B_iQyohNPb5_2),.dout(w_dff_B_2syLQrTk8_2),.clk(gclk));
	jdff dff_B_c6BjeoqK3_2(.din(w_dff_B_2syLQrTk8_2),.dout(w_dff_B_c6BjeoqK3_2),.clk(gclk));
	jdff dff_B_5CWHnyk14_2(.din(w_dff_B_c6BjeoqK3_2),.dout(w_dff_B_5CWHnyk14_2),.clk(gclk));
	jdff dff_B_1ev366XH7_2(.din(w_dff_B_5CWHnyk14_2),.dout(w_dff_B_1ev366XH7_2),.clk(gclk));
	jdff dff_B_kAPCeusT6_2(.din(w_dff_B_1ev366XH7_2),.dout(w_dff_B_kAPCeusT6_2),.clk(gclk));
	jdff dff_B_Ui9tzaJe3_2(.din(w_dff_B_kAPCeusT6_2),.dout(w_dff_B_Ui9tzaJe3_2),.clk(gclk));
	jdff dff_B_8hseRavn4_2(.din(w_dff_B_Ui9tzaJe3_2),.dout(w_dff_B_8hseRavn4_2),.clk(gclk));
	jdff dff_B_1hIBzhWY4_2(.din(w_dff_B_8hseRavn4_2),.dout(w_dff_B_1hIBzhWY4_2),.clk(gclk));
	jdff dff_B_yPUbsZcR6_2(.din(w_dff_B_1hIBzhWY4_2),.dout(w_dff_B_yPUbsZcR6_2),.clk(gclk));
	jdff dff_B_0Yx81Hka1_2(.din(w_dff_B_yPUbsZcR6_2),.dout(w_dff_B_0Yx81Hka1_2),.clk(gclk));
	jdff dff_B_0iY5WYrK6_2(.din(w_dff_B_0Yx81Hka1_2),.dout(w_dff_B_0iY5WYrK6_2),.clk(gclk));
	jdff dff_B_vIluE7Hi3_2(.din(w_dff_B_0iY5WYrK6_2),.dout(w_dff_B_vIluE7Hi3_2),.clk(gclk));
	jdff dff_B_jO7epaEW3_2(.din(w_dff_B_vIluE7Hi3_2),.dout(w_dff_B_jO7epaEW3_2),.clk(gclk));
	jdff dff_B_Qwxy4cgT8_2(.din(w_dff_B_jO7epaEW3_2),.dout(w_dff_B_Qwxy4cgT8_2),.clk(gclk));
	jdff dff_B_6P7mbnmE0_2(.din(w_dff_B_Qwxy4cgT8_2),.dout(w_dff_B_6P7mbnmE0_2),.clk(gclk));
	jdff dff_B_T9lmb8lD4_2(.din(w_dff_B_6P7mbnmE0_2),.dout(w_dff_B_T9lmb8lD4_2),.clk(gclk));
	jdff dff_B_uBmoyWnJ8_2(.din(w_dff_B_T9lmb8lD4_2),.dout(w_dff_B_uBmoyWnJ8_2),.clk(gclk));
	jdff dff_B_aXfjF8iJ7_2(.din(w_dff_B_uBmoyWnJ8_2),.dout(w_dff_B_aXfjF8iJ7_2),.clk(gclk));
	jdff dff_B_L5RnNB3u8_2(.din(w_dff_B_aXfjF8iJ7_2),.dout(w_dff_B_L5RnNB3u8_2),.clk(gclk));
	jdff dff_B_F3I74PE33_2(.din(w_dff_B_L5RnNB3u8_2),.dout(w_dff_B_F3I74PE33_2),.clk(gclk));
	jdff dff_B_OSC9w5fH6_2(.din(w_dff_B_F3I74PE33_2),.dout(w_dff_B_OSC9w5fH6_2),.clk(gclk));
	jdff dff_B_7aV4A1kK0_2(.din(w_dff_B_OSC9w5fH6_2),.dout(w_dff_B_7aV4A1kK0_2),.clk(gclk));
	jdff dff_B_Vqb8uKpm7_2(.din(w_dff_B_7aV4A1kK0_2),.dout(w_dff_B_Vqb8uKpm7_2),.clk(gclk));
	jdff dff_B_VZEGaTD22_2(.din(w_dff_B_Vqb8uKpm7_2),.dout(w_dff_B_VZEGaTD22_2),.clk(gclk));
	jdff dff_B_e2dWQ5mI9_2(.din(w_dff_B_VZEGaTD22_2),.dout(w_dff_B_e2dWQ5mI9_2),.clk(gclk));
	jdff dff_B_eWJ0iAyU8_2(.din(w_dff_B_e2dWQ5mI9_2),.dout(w_dff_B_eWJ0iAyU8_2),.clk(gclk));
	jdff dff_B_yTiDZGKA7_2(.din(w_dff_B_eWJ0iAyU8_2),.dout(w_dff_B_yTiDZGKA7_2),.clk(gclk));
	jdff dff_B_BB7c8lP05_2(.din(w_dff_B_yTiDZGKA7_2),.dout(w_dff_B_BB7c8lP05_2),.clk(gclk));
	jdff dff_B_9VhKkMOn9_2(.din(w_dff_B_BB7c8lP05_2),.dout(w_dff_B_9VhKkMOn9_2),.clk(gclk));
	jdff dff_B_gBhgOVnT1_2(.din(w_dff_B_9VhKkMOn9_2),.dout(w_dff_B_gBhgOVnT1_2),.clk(gclk));
	jdff dff_B_89y1K2Xs8_2(.din(w_dff_B_gBhgOVnT1_2),.dout(w_dff_B_89y1K2Xs8_2),.clk(gclk));
	jdff dff_B_mk4QHZQS7_2(.din(n1589),.dout(w_dff_B_mk4QHZQS7_2),.clk(gclk));
	jdff dff_B_SAOoRhsC9_1(.din(n1587),.dout(w_dff_B_SAOoRhsC9_1),.clk(gclk));
	jdff dff_B_XjefX4721_2(.din(n1522),.dout(w_dff_B_XjefX4721_2),.clk(gclk));
	jdff dff_B_NolhAyI60_2(.din(w_dff_B_XjefX4721_2),.dout(w_dff_B_NolhAyI60_2),.clk(gclk));
	jdff dff_B_5Ux9wGwm5_2(.din(w_dff_B_NolhAyI60_2),.dout(w_dff_B_5Ux9wGwm5_2),.clk(gclk));
	jdff dff_B_LD6nPV3L0_2(.din(w_dff_B_5Ux9wGwm5_2),.dout(w_dff_B_LD6nPV3L0_2),.clk(gclk));
	jdff dff_B_qi2cPUYf2_2(.din(w_dff_B_LD6nPV3L0_2),.dout(w_dff_B_qi2cPUYf2_2),.clk(gclk));
	jdff dff_B_EnY0yLLv9_2(.din(w_dff_B_qi2cPUYf2_2),.dout(w_dff_B_EnY0yLLv9_2),.clk(gclk));
	jdff dff_B_aKQqJcDg9_2(.din(w_dff_B_EnY0yLLv9_2),.dout(w_dff_B_aKQqJcDg9_2),.clk(gclk));
	jdff dff_B_ZClTf7qy1_2(.din(w_dff_B_aKQqJcDg9_2),.dout(w_dff_B_ZClTf7qy1_2),.clk(gclk));
	jdff dff_B_IpAfcqwl0_2(.din(w_dff_B_ZClTf7qy1_2),.dout(w_dff_B_IpAfcqwl0_2),.clk(gclk));
	jdff dff_B_mrKCDw2q9_2(.din(w_dff_B_IpAfcqwl0_2),.dout(w_dff_B_mrKCDw2q9_2),.clk(gclk));
	jdff dff_B_U08s84Q54_2(.din(w_dff_B_mrKCDw2q9_2),.dout(w_dff_B_U08s84Q54_2),.clk(gclk));
	jdff dff_B_YVAuNIrv0_2(.din(w_dff_B_U08s84Q54_2),.dout(w_dff_B_YVAuNIrv0_2),.clk(gclk));
	jdff dff_B_0LxnTeCw2_2(.din(w_dff_B_YVAuNIrv0_2),.dout(w_dff_B_0LxnTeCw2_2),.clk(gclk));
	jdff dff_B_9xHkYdKc0_2(.din(w_dff_B_0LxnTeCw2_2),.dout(w_dff_B_9xHkYdKc0_2),.clk(gclk));
	jdff dff_B_l4Mnnc7U8_2(.din(w_dff_B_9xHkYdKc0_2),.dout(w_dff_B_l4Mnnc7U8_2),.clk(gclk));
	jdff dff_B_W0QLLP3E9_2(.din(w_dff_B_l4Mnnc7U8_2),.dout(w_dff_B_W0QLLP3E9_2),.clk(gclk));
	jdff dff_B_kJ4UVvww1_2(.din(w_dff_B_W0QLLP3E9_2),.dout(w_dff_B_kJ4UVvww1_2),.clk(gclk));
	jdff dff_B_iYxINs7f7_2(.din(w_dff_B_kJ4UVvww1_2),.dout(w_dff_B_iYxINs7f7_2),.clk(gclk));
	jdff dff_B_IS2dR1B27_2(.din(w_dff_B_iYxINs7f7_2),.dout(w_dff_B_IS2dR1B27_2),.clk(gclk));
	jdff dff_B_7k2RvW6g1_2(.din(w_dff_B_IS2dR1B27_2),.dout(w_dff_B_7k2RvW6g1_2),.clk(gclk));
	jdff dff_B_v75OYDqx0_2(.din(w_dff_B_7k2RvW6g1_2),.dout(w_dff_B_v75OYDqx0_2),.clk(gclk));
	jdff dff_B_f3JmymHX2_2(.din(w_dff_B_v75OYDqx0_2),.dout(w_dff_B_f3JmymHX2_2),.clk(gclk));
	jdff dff_B_xnqkOxxm0_2(.din(w_dff_B_f3JmymHX2_2),.dout(w_dff_B_xnqkOxxm0_2),.clk(gclk));
	jdff dff_B_s6uW2cIn2_2(.din(w_dff_B_xnqkOxxm0_2),.dout(w_dff_B_s6uW2cIn2_2),.clk(gclk));
	jdff dff_B_XRBAfsxD8_2(.din(w_dff_B_s6uW2cIn2_2),.dout(w_dff_B_XRBAfsxD8_2),.clk(gclk));
	jdff dff_B_YwwbrA3T6_2(.din(w_dff_B_XRBAfsxD8_2),.dout(w_dff_B_YwwbrA3T6_2),.clk(gclk));
	jdff dff_B_ndj0dHNJ8_2(.din(w_dff_B_YwwbrA3T6_2),.dout(w_dff_B_ndj0dHNJ8_2),.clk(gclk));
	jdff dff_B_6bjCgydK2_2(.din(w_dff_B_ndj0dHNJ8_2),.dout(w_dff_B_6bjCgydK2_2),.clk(gclk));
	jdff dff_B_vpcUPsY24_2(.din(w_dff_B_6bjCgydK2_2),.dout(w_dff_B_vpcUPsY24_2),.clk(gclk));
	jdff dff_B_3eIUFEBL4_2(.din(w_dff_B_vpcUPsY24_2),.dout(w_dff_B_3eIUFEBL4_2),.clk(gclk));
	jdff dff_B_yz6ItiD02_2(.din(w_dff_B_3eIUFEBL4_2),.dout(w_dff_B_yz6ItiD02_2),.clk(gclk));
	jdff dff_B_OYI5TTQ27_2(.din(w_dff_B_yz6ItiD02_2),.dout(w_dff_B_OYI5TTQ27_2),.clk(gclk));
	jdff dff_B_sEVUrz8g0_2(.din(w_dff_B_OYI5TTQ27_2),.dout(w_dff_B_sEVUrz8g0_2),.clk(gclk));
	jdff dff_B_4P5mUltv6_2(.din(n1525),.dout(w_dff_B_4P5mUltv6_2),.clk(gclk));
	jdff dff_B_TCdl79rD8_1(.din(n1523),.dout(w_dff_B_TCdl79rD8_1),.clk(gclk));
	jdff dff_B_edWN1NhW4_2(.din(n1451),.dout(w_dff_B_edWN1NhW4_2),.clk(gclk));
	jdff dff_B_HHx47qXL1_2(.din(w_dff_B_edWN1NhW4_2),.dout(w_dff_B_HHx47qXL1_2),.clk(gclk));
	jdff dff_B_rc7qgt0a3_2(.din(w_dff_B_HHx47qXL1_2),.dout(w_dff_B_rc7qgt0a3_2),.clk(gclk));
	jdff dff_B_dIWe51b91_2(.din(w_dff_B_rc7qgt0a3_2),.dout(w_dff_B_dIWe51b91_2),.clk(gclk));
	jdff dff_B_HHe1uSsr2_2(.din(w_dff_B_dIWe51b91_2),.dout(w_dff_B_HHe1uSsr2_2),.clk(gclk));
	jdff dff_B_UUMlViDm1_2(.din(w_dff_B_HHe1uSsr2_2),.dout(w_dff_B_UUMlViDm1_2),.clk(gclk));
	jdff dff_B_FACeCpGh4_2(.din(w_dff_B_UUMlViDm1_2),.dout(w_dff_B_FACeCpGh4_2),.clk(gclk));
	jdff dff_B_FRwGckXt5_2(.din(w_dff_B_FACeCpGh4_2),.dout(w_dff_B_FRwGckXt5_2),.clk(gclk));
	jdff dff_B_1DapE0cs9_2(.din(w_dff_B_FRwGckXt5_2),.dout(w_dff_B_1DapE0cs9_2),.clk(gclk));
	jdff dff_B_JVZC70tZ0_2(.din(w_dff_B_1DapE0cs9_2),.dout(w_dff_B_JVZC70tZ0_2),.clk(gclk));
	jdff dff_B_ljxaKdkG0_2(.din(w_dff_B_JVZC70tZ0_2),.dout(w_dff_B_ljxaKdkG0_2),.clk(gclk));
	jdff dff_B_VOthYxX98_2(.din(w_dff_B_ljxaKdkG0_2),.dout(w_dff_B_VOthYxX98_2),.clk(gclk));
	jdff dff_B_fdfOxRjd5_2(.din(w_dff_B_VOthYxX98_2),.dout(w_dff_B_fdfOxRjd5_2),.clk(gclk));
	jdff dff_B_XKiqIZ5r4_2(.din(w_dff_B_fdfOxRjd5_2),.dout(w_dff_B_XKiqIZ5r4_2),.clk(gclk));
	jdff dff_B_NeSmKgSE2_2(.din(w_dff_B_XKiqIZ5r4_2),.dout(w_dff_B_NeSmKgSE2_2),.clk(gclk));
	jdff dff_B_F3SclU8R3_2(.din(w_dff_B_NeSmKgSE2_2),.dout(w_dff_B_F3SclU8R3_2),.clk(gclk));
	jdff dff_B_XSyHIbcY0_2(.din(w_dff_B_F3SclU8R3_2),.dout(w_dff_B_XSyHIbcY0_2),.clk(gclk));
	jdff dff_B_4LHxSwYK3_2(.din(w_dff_B_XSyHIbcY0_2),.dout(w_dff_B_4LHxSwYK3_2),.clk(gclk));
	jdff dff_B_P187kyDT4_2(.din(w_dff_B_4LHxSwYK3_2),.dout(w_dff_B_P187kyDT4_2),.clk(gclk));
	jdff dff_B_v0lmHB5I7_2(.din(w_dff_B_P187kyDT4_2),.dout(w_dff_B_v0lmHB5I7_2),.clk(gclk));
	jdff dff_B_wVKtpP5L9_2(.din(w_dff_B_v0lmHB5I7_2),.dout(w_dff_B_wVKtpP5L9_2),.clk(gclk));
	jdff dff_B_vYdEo0Fz2_2(.din(w_dff_B_wVKtpP5L9_2),.dout(w_dff_B_vYdEo0Fz2_2),.clk(gclk));
	jdff dff_B_hz8Uspyn5_2(.din(w_dff_B_vYdEo0Fz2_2),.dout(w_dff_B_hz8Uspyn5_2),.clk(gclk));
	jdff dff_B_zRU4CEaB0_2(.din(w_dff_B_hz8Uspyn5_2),.dout(w_dff_B_zRU4CEaB0_2),.clk(gclk));
	jdff dff_B_5zbn9sFc5_2(.din(w_dff_B_zRU4CEaB0_2),.dout(w_dff_B_5zbn9sFc5_2),.clk(gclk));
	jdff dff_B_7ubZMhHE7_2(.din(w_dff_B_5zbn9sFc5_2),.dout(w_dff_B_7ubZMhHE7_2),.clk(gclk));
	jdff dff_B_7EEoPkXK2_2(.din(w_dff_B_7ubZMhHE7_2),.dout(w_dff_B_7EEoPkXK2_2),.clk(gclk));
	jdff dff_B_VsStI1L86_2(.din(w_dff_B_7EEoPkXK2_2),.dout(w_dff_B_VsStI1L86_2),.clk(gclk));
	jdff dff_B_hT9Ev7Vt9_2(.din(w_dff_B_VsStI1L86_2),.dout(w_dff_B_hT9Ev7Vt9_2),.clk(gclk));
	jdff dff_B_qdYNCKvA2_2(.din(n1454),.dout(w_dff_B_qdYNCKvA2_2),.clk(gclk));
	jdff dff_B_QsPz98oR1_1(.din(n1452),.dout(w_dff_B_QsPz98oR1_1),.clk(gclk));
	jdff dff_B_GrRxEaNu6_2(.din(n1373),.dout(w_dff_B_GrRxEaNu6_2),.clk(gclk));
	jdff dff_B_rEGRSoG71_2(.din(w_dff_B_GrRxEaNu6_2),.dout(w_dff_B_rEGRSoG71_2),.clk(gclk));
	jdff dff_B_tGa8r5Lc4_2(.din(w_dff_B_rEGRSoG71_2),.dout(w_dff_B_tGa8r5Lc4_2),.clk(gclk));
	jdff dff_B_ejkEqu0H3_2(.din(w_dff_B_tGa8r5Lc4_2),.dout(w_dff_B_ejkEqu0H3_2),.clk(gclk));
	jdff dff_B_2NN5B2kf0_2(.din(w_dff_B_ejkEqu0H3_2),.dout(w_dff_B_2NN5B2kf0_2),.clk(gclk));
	jdff dff_B_RHDjHqwB8_2(.din(w_dff_B_2NN5B2kf0_2),.dout(w_dff_B_RHDjHqwB8_2),.clk(gclk));
	jdff dff_B_QEiEL3mN7_2(.din(w_dff_B_RHDjHqwB8_2),.dout(w_dff_B_QEiEL3mN7_2),.clk(gclk));
	jdff dff_B_JJKIdqw52_2(.din(w_dff_B_QEiEL3mN7_2),.dout(w_dff_B_JJKIdqw52_2),.clk(gclk));
	jdff dff_B_OUNeJMVY8_2(.din(w_dff_B_JJKIdqw52_2),.dout(w_dff_B_OUNeJMVY8_2),.clk(gclk));
	jdff dff_B_xkoXLOF85_2(.din(w_dff_B_OUNeJMVY8_2),.dout(w_dff_B_xkoXLOF85_2),.clk(gclk));
	jdff dff_B_Jed5Tjm11_2(.din(w_dff_B_xkoXLOF85_2),.dout(w_dff_B_Jed5Tjm11_2),.clk(gclk));
	jdff dff_B_mp4F1oZH8_2(.din(w_dff_B_Jed5Tjm11_2),.dout(w_dff_B_mp4F1oZH8_2),.clk(gclk));
	jdff dff_B_eEJfo6TG8_2(.din(w_dff_B_mp4F1oZH8_2),.dout(w_dff_B_eEJfo6TG8_2),.clk(gclk));
	jdff dff_B_RO0EvG131_2(.din(w_dff_B_eEJfo6TG8_2),.dout(w_dff_B_RO0EvG131_2),.clk(gclk));
	jdff dff_B_0hbscURz9_2(.din(w_dff_B_RO0EvG131_2),.dout(w_dff_B_0hbscURz9_2),.clk(gclk));
	jdff dff_B_uErcEyIz3_2(.din(w_dff_B_0hbscURz9_2),.dout(w_dff_B_uErcEyIz3_2),.clk(gclk));
	jdff dff_B_8wOoISR05_2(.din(w_dff_B_uErcEyIz3_2),.dout(w_dff_B_8wOoISR05_2),.clk(gclk));
	jdff dff_B_fKU9188e7_2(.din(w_dff_B_8wOoISR05_2),.dout(w_dff_B_fKU9188e7_2),.clk(gclk));
	jdff dff_B_ZbKGSvYT9_2(.din(w_dff_B_fKU9188e7_2),.dout(w_dff_B_ZbKGSvYT9_2),.clk(gclk));
	jdff dff_B_MqbE7NgF3_2(.din(w_dff_B_ZbKGSvYT9_2),.dout(w_dff_B_MqbE7NgF3_2),.clk(gclk));
	jdff dff_B_OoAHvFgV5_2(.din(w_dff_B_MqbE7NgF3_2),.dout(w_dff_B_OoAHvFgV5_2),.clk(gclk));
	jdff dff_B_qf2DMypr4_2(.din(w_dff_B_OoAHvFgV5_2),.dout(w_dff_B_qf2DMypr4_2),.clk(gclk));
	jdff dff_B_pMKCDJvG9_2(.din(w_dff_B_qf2DMypr4_2),.dout(w_dff_B_pMKCDJvG9_2),.clk(gclk));
	jdff dff_B_VrZdiStE9_2(.din(w_dff_B_pMKCDJvG9_2),.dout(w_dff_B_VrZdiStE9_2),.clk(gclk));
	jdff dff_B_7bdxXkSP7_2(.din(w_dff_B_VrZdiStE9_2),.dout(w_dff_B_7bdxXkSP7_2),.clk(gclk));
	jdff dff_B_c1BRs3pm3_2(.din(n1376),.dout(w_dff_B_c1BRs3pm3_2),.clk(gclk));
	jdff dff_B_f3NceXEh7_1(.din(n1374),.dout(w_dff_B_f3NceXEh7_1),.clk(gclk));
	jdff dff_B_lCx35bWy3_2(.din(n1288),.dout(w_dff_B_lCx35bWy3_2),.clk(gclk));
	jdff dff_B_AztIEZv59_2(.din(w_dff_B_lCx35bWy3_2),.dout(w_dff_B_AztIEZv59_2),.clk(gclk));
	jdff dff_B_d7TUXjew0_2(.din(w_dff_B_AztIEZv59_2),.dout(w_dff_B_d7TUXjew0_2),.clk(gclk));
	jdff dff_B_k9Jg1eEh3_2(.din(w_dff_B_d7TUXjew0_2),.dout(w_dff_B_k9Jg1eEh3_2),.clk(gclk));
	jdff dff_B_124TKauY1_2(.din(w_dff_B_k9Jg1eEh3_2),.dout(w_dff_B_124TKauY1_2),.clk(gclk));
	jdff dff_B_mOF0fu9Y5_2(.din(w_dff_B_124TKauY1_2),.dout(w_dff_B_mOF0fu9Y5_2),.clk(gclk));
	jdff dff_B_Kl3R1ejy5_2(.din(w_dff_B_mOF0fu9Y5_2),.dout(w_dff_B_Kl3R1ejy5_2),.clk(gclk));
	jdff dff_B_qfbSuO2U5_2(.din(w_dff_B_Kl3R1ejy5_2),.dout(w_dff_B_qfbSuO2U5_2),.clk(gclk));
	jdff dff_B_iPLNtMfH4_2(.din(w_dff_B_qfbSuO2U5_2),.dout(w_dff_B_iPLNtMfH4_2),.clk(gclk));
	jdff dff_B_LFvrOSLM2_2(.din(w_dff_B_iPLNtMfH4_2),.dout(w_dff_B_LFvrOSLM2_2),.clk(gclk));
	jdff dff_B_y5xnIrsl7_2(.din(w_dff_B_LFvrOSLM2_2),.dout(w_dff_B_y5xnIrsl7_2),.clk(gclk));
	jdff dff_B_KiJengFT6_2(.din(w_dff_B_y5xnIrsl7_2),.dout(w_dff_B_KiJengFT6_2),.clk(gclk));
	jdff dff_B_Ha11kADe9_2(.din(w_dff_B_KiJengFT6_2),.dout(w_dff_B_Ha11kADe9_2),.clk(gclk));
	jdff dff_B_UrtMm4fC2_2(.din(w_dff_B_Ha11kADe9_2),.dout(w_dff_B_UrtMm4fC2_2),.clk(gclk));
	jdff dff_B_n98Zh5Uc4_2(.din(w_dff_B_UrtMm4fC2_2),.dout(w_dff_B_n98Zh5Uc4_2),.clk(gclk));
	jdff dff_B_6BtnarNa7_2(.din(w_dff_B_n98Zh5Uc4_2),.dout(w_dff_B_6BtnarNa7_2),.clk(gclk));
	jdff dff_B_WIL0cb5J4_2(.din(w_dff_B_6BtnarNa7_2),.dout(w_dff_B_WIL0cb5J4_2),.clk(gclk));
	jdff dff_B_NqJgbb3l5_2(.din(w_dff_B_WIL0cb5J4_2),.dout(w_dff_B_NqJgbb3l5_2),.clk(gclk));
	jdff dff_B_bPKMX1LZ2_2(.din(w_dff_B_NqJgbb3l5_2),.dout(w_dff_B_bPKMX1LZ2_2),.clk(gclk));
	jdff dff_B_gOxNeTZb8_2(.din(w_dff_B_bPKMX1LZ2_2),.dout(w_dff_B_gOxNeTZb8_2),.clk(gclk));
	jdff dff_B_3XfacPBE0_2(.din(w_dff_B_gOxNeTZb8_2),.dout(w_dff_B_3XfacPBE0_2),.clk(gclk));
	jdff dff_B_Za8DoiXy7_1(.din(n1289),.dout(w_dff_B_Za8DoiXy7_1),.clk(gclk));
	jdff dff_B_r5fzfAxf9_2(.din(n1198),.dout(w_dff_B_r5fzfAxf9_2),.clk(gclk));
	jdff dff_B_ePE49Jzy5_2(.din(w_dff_B_r5fzfAxf9_2),.dout(w_dff_B_ePE49Jzy5_2),.clk(gclk));
	jdff dff_B_Ve2RcBtt0_2(.din(w_dff_B_ePE49Jzy5_2),.dout(w_dff_B_Ve2RcBtt0_2),.clk(gclk));
	jdff dff_B_Mz06rtE93_2(.din(w_dff_B_Ve2RcBtt0_2),.dout(w_dff_B_Mz06rtE93_2),.clk(gclk));
	jdff dff_B_9CMdKNfD5_2(.din(w_dff_B_Mz06rtE93_2),.dout(w_dff_B_9CMdKNfD5_2),.clk(gclk));
	jdff dff_B_b8GLL0Nk3_2(.din(w_dff_B_9CMdKNfD5_2),.dout(w_dff_B_b8GLL0Nk3_2),.clk(gclk));
	jdff dff_B_h7pYsV878_2(.din(w_dff_B_b8GLL0Nk3_2),.dout(w_dff_B_h7pYsV878_2),.clk(gclk));
	jdff dff_B_lE00m7Z73_2(.din(w_dff_B_h7pYsV878_2),.dout(w_dff_B_lE00m7Z73_2),.clk(gclk));
	jdff dff_B_eRPL2gmp0_2(.din(w_dff_B_lE00m7Z73_2),.dout(w_dff_B_eRPL2gmp0_2),.clk(gclk));
	jdff dff_B_a6kvGCiD9_2(.din(w_dff_B_eRPL2gmp0_2),.dout(w_dff_B_a6kvGCiD9_2),.clk(gclk));
	jdff dff_B_L9TnrSUB8_2(.din(w_dff_B_a6kvGCiD9_2),.dout(w_dff_B_L9TnrSUB8_2),.clk(gclk));
	jdff dff_B_baOIVWVp9_2(.din(w_dff_B_L9TnrSUB8_2),.dout(w_dff_B_baOIVWVp9_2),.clk(gclk));
	jdff dff_B_R8slybch4_2(.din(w_dff_B_baOIVWVp9_2),.dout(w_dff_B_R8slybch4_2),.clk(gclk));
	jdff dff_B_6hbSk1TN9_2(.din(w_dff_B_R8slybch4_2),.dout(w_dff_B_6hbSk1TN9_2),.clk(gclk));
	jdff dff_B_ddo9L6QE0_2(.din(w_dff_B_6hbSk1TN9_2),.dout(w_dff_B_ddo9L6QE0_2),.clk(gclk));
	jdff dff_B_MczcRKuC2_2(.din(w_dff_B_ddo9L6QE0_2),.dout(w_dff_B_MczcRKuC2_2),.clk(gclk));
	jdff dff_B_nvfTUSFu6_2(.din(w_dff_B_MczcRKuC2_2),.dout(w_dff_B_nvfTUSFu6_2),.clk(gclk));
	jdff dff_B_Xiu0xkK29_2(.din(w_dff_B_nvfTUSFu6_2),.dout(w_dff_B_Xiu0xkK29_2),.clk(gclk));
	jdff dff_B_msSltTL19_2(.din(n1215),.dout(w_dff_B_msSltTL19_2),.clk(gclk));
	jdff dff_B_af6URBAC0_1(.din(n1199),.dout(w_dff_B_af6URBAC0_1),.clk(gclk));
	jdff dff_B_oYP1l3rM5_2(.din(n1094),.dout(w_dff_B_oYP1l3rM5_2),.clk(gclk));
	jdff dff_B_gRf78oQM8_2(.din(w_dff_B_oYP1l3rM5_2),.dout(w_dff_B_gRf78oQM8_2),.clk(gclk));
	jdff dff_B_tgN7iGGJ7_2(.din(w_dff_B_gRf78oQM8_2),.dout(w_dff_B_tgN7iGGJ7_2),.clk(gclk));
	jdff dff_B_l7CesZvX9_2(.din(w_dff_B_tgN7iGGJ7_2),.dout(w_dff_B_l7CesZvX9_2),.clk(gclk));
	jdff dff_B_ezaZEJrp5_2(.din(w_dff_B_l7CesZvX9_2),.dout(w_dff_B_ezaZEJrp5_2),.clk(gclk));
	jdff dff_B_RfHQRe791_2(.din(w_dff_B_ezaZEJrp5_2),.dout(w_dff_B_RfHQRe791_2),.clk(gclk));
	jdff dff_B_dsUBNTIy8_2(.din(w_dff_B_RfHQRe791_2),.dout(w_dff_B_dsUBNTIy8_2),.clk(gclk));
	jdff dff_B_nWAzqlwX2_2(.din(w_dff_B_dsUBNTIy8_2),.dout(w_dff_B_nWAzqlwX2_2),.clk(gclk));
	jdff dff_B_RaF2pSzQ5_2(.din(w_dff_B_nWAzqlwX2_2),.dout(w_dff_B_RaF2pSzQ5_2),.clk(gclk));
	jdff dff_B_VZxdJc120_2(.din(w_dff_B_RaF2pSzQ5_2),.dout(w_dff_B_VZxdJc120_2),.clk(gclk));
	jdff dff_B_L5Z5gPi44_2(.din(w_dff_B_VZxdJc120_2),.dout(w_dff_B_L5Z5gPi44_2),.clk(gclk));
	jdff dff_B_Px5rwGni0_2(.din(w_dff_B_L5Z5gPi44_2),.dout(w_dff_B_Px5rwGni0_2),.clk(gclk));
	jdff dff_B_sbDZY1tI2_2(.din(w_dff_B_Px5rwGni0_2),.dout(w_dff_B_sbDZY1tI2_2),.clk(gclk));
	jdff dff_B_WtGIh4183_2(.din(w_dff_B_sbDZY1tI2_2),.dout(w_dff_B_WtGIh4183_2),.clk(gclk));
	jdff dff_B_9P0YEedD2_2(.din(w_dff_B_WtGIh4183_2),.dout(w_dff_B_9P0YEedD2_2),.clk(gclk));
	jdff dff_B_RSnN9Bqc6_2(.din(n1117),.dout(w_dff_B_RSnN9Bqc6_2),.clk(gclk));
	jdff dff_B_GbnFbinF7_2(.din(w_dff_B_RSnN9Bqc6_2),.dout(w_dff_B_GbnFbinF7_2),.clk(gclk));
	jdff dff_B_JdMX0b1g2_1(.din(n1095),.dout(w_dff_B_JdMX0b1g2_1),.clk(gclk));
	jdff dff_B_eeCbMqGg7_2(.din(n996),.dout(w_dff_B_eeCbMqGg7_2),.clk(gclk));
	jdff dff_B_z1LRiTOE0_2(.din(w_dff_B_eeCbMqGg7_2),.dout(w_dff_B_z1LRiTOE0_2),.clk(gclk));
	jdff dff_B_gv3NYn6P6_2(.din(w_dff_B_z1LRiTOE0_2),.dout(w_dff_B_gv3NYn6P6_2),.clk(gclk));
	jdff dff_B_1ENQgEHy7_2(.din(w_dff_B_gv3NYn6P6_2),.dout(w_dff_B_1ENQgEHy7_2),.clk(gclk));
	jdff dff_B_vijbYQq07_2(.din(w_dff_B_1ENQgEHy7_2),.dout(w_dff_B_vijbYQq07_2),.clk(gclk));
	jdff dff_B_BhQpaSSH3_2(.din(w_dff_B_vijbYQq07_2),.dout(w_dff_B_BhQpaSSH3_2),.clk(gclk));
	jdff dff_B_CBo7bbq76_2(.din(w_dff_B_BhQpaSSH3_2),.dout(w_dff_B_CBo7bbq76_2),.clk(gclk));
	jdff dff_B_JYBkCv3n7_2(.din(w_dff_B_CBo7bbq76_2),.dout(w_dff_B_JYBkCv3n7_2),.clk(gclk));
	jdff dff_B_edUcnAT04_2(.din(w_dff_B_JYBkCv3n7_2),.dout(w_dff_B_edUcnAT04_2),.clk(gclk));
	jdff dff_B_yHYHauRk5_2(.din(w_dff_B_edUcnAT04_2),.dout(w_dff_B_yHYHauRk5_2),.clk(gclk));
	jdff dff_B_eCVnUcVL2_2(.din(w_dff_B_yHYHauRk5_2),.dout(w_dff_B_eCVnUcVL2_2),.clk(gclk));
	jdff dff_B_RN7mN8hd4_2(.din(w_dff_B_eCVnUcVL2_2),.dout(w_dff_B_RN7mN8hd4_2),.clk(gclk));
	jdff dff_B_DOAQMQjL2_2(.din(n1012),.dout(w_dff_B_DOAQMQjL2_2),.clk(gclk));
	jdff dff_B_QkUk3v3e1_2(.din(w_dff_B_DOAQMQjL2_2),.dout(w_dff_B_QkUk3v3e1_2),.clk(gclk));
	jdff dff_B_PJf0cWwu9_1(.din(n997),.dout(w_dff_B_PJf0cWwu9_1),.clk(gclk));
	jdff dff_B_h9kLTsBE7_2(.din(n891),.dout(w_dff_B_h9kLTsBE7_2),.clk(gclk));
	jdff dff_B_3IuYWM1f7_2(.din(w_dff_B_h9kLTsBE7_2),.dout(w_dff_B_3IuYWM1f7_2),.clk(gclk));
	jdff dff_B_ZSeLQX9n7_2(.din(w_dff_B_3IuYWM1f7_2),.dout(w_dff_B_ZSeLQX9n7_2),.clk(gclk));
	jdff dff_B_nGXJ12E88_2(.din(w_dff_B_ZSeLQX9n7_2),.dout(w_dff_B_nGXJ12E88_2),.clk(gclk));
	jdff dff_B_HdZ7ZILy2_2(.din(w_dff_B_nGXJ12E88_2),.dout(w_dff_B_HdZ7ZILy2_2),.clk(gclk));
	jdff dff_B_xWtGqVjE0_2(.din(w_dff_B_HdZ7ZILy2_2),.dout(w_dff_B_xWtGqVjE0_2),.clk(gclk));
	jdff dff_B_aTqj50vP2_2(.din(w_dff_B_xWtGqVjE0_2),.dout(w_dff_B_aTqj50vP2_2),.clk(gclk));
	jdff dff_B_FKjZDHFt8_2(.din(w_dff_B_aTqj50vP2_2),.dout(w_dff_B_FKjZDHFt8_2),.clk(gclk));
	jdff dff_B_PJROlhI89_2(.din(w_dff_B_FKjZDHFt8_2),.dout(w_dff_B_PJROlhI89_2),.clk(gclk));
	jdff dff_B_WNF3HEs58_2(.din(n907),.dout(w_dff_B_WNF3HEs58_2),.clk(gclk));
	jdff dff_B_6IN4EJlK2_2(.din(w_dff_B_WNF3HEs58_2),.dout(w_dff_B_6IN4EJlK2_2),.clk(gclk));
	jdff dff_B_sYNSHnuN6_2(.din(w_dff_B_6IN4EJlK2_2),.dout(w_dff_B_sYNSHnuN6_2),.clk(gclk));
	jdff dff_B_yTJ3of4o1_1(.din(n892),.dout(w_dff_B_yTJ3of4o1_1),.clk(gclk));
	jdff dff_B_7Qv96jdo5_1(.din(w_dff_B_yTJ3of4o1_1),.dout(w_dff_B_7Qv96jdo5_1),.clk(gclk));
	jdff dff_B_qojY8BTd6_1(.din(w_dff_B_7Qv96jdo5_1),.dout(w_dff_B_qojY8BTd6_1),.clk(gclk));
	jdff dff_B_3WH9b8qn6_1(.din(w_dff_B_qojY8BTd6_1),.dout(w_dff_B_3WH9b8qn6_1),.clk(gclk));
	jdff dff_B_l0OJj6WW6_1(.din(w_dff_B_3WH9b8qn6_1),.dout(w_dff_B_l0OJj6WW6_1),.clk(gclk));
	jdff dff_B_Q36U5tAt1_1(.din(w_dff_B_l0OJj6WW6_1),.dout(w_dff_B_Q36U5tAt1_1),.clk(gclk));
	jdff dff_B_UmxfwUrb4_0(.din(n801),.dout(w_dff_B_UmxfwUrb4_0),.clk(gclk));
	jdff dff_B_l1FIUshX7_0(.din(w_dff_B_UmxfwUrb4_0),.dout(w_dff_B_l1FIUshX7_0),.clk(gclk));
	jdff dff_A_IZ0xkOZa6_0(.dout(w_n800_0[0]),.din(w_dff_A_IZ0xkOZa6_0),.clk(gclk));
	jdff dff_A_Vp1im4IS8_0(.dout(w_dff_A_IZ0xkOZa6_0),.din(w_dff_A_Vp1im4IS8_0),.clk(gclk));
	jdff dff_A_xxdJDKKt3_0(.dout(w_dff_A_Vp1im4IS8_0),.din(w_dff_A_xxdJDKKt3_0),.clk(gclk));
	jdff dff_B_fexZ1vyZ4_1(.din(n794),.dout(w_dff_B_fexZ1vyZ4_1),.clk(gclk));
	jdff dff_A_PWnxLbLl4_0(.dout(w_n698_0[0]),.din(w_dff_A_PWnxLbLl4_0),.clk(gclk));
	jdff dff_A_sW6BxUtj5_1(.dout(w_n698_0[1]),.din(w_dff_A_sW6BxUtj5_1),.clk(gclk));
	jdff dff_A_j2EXnS4j2_1(.dout(w_dff_A_sW6BxUtj5_1),.din(w_dff_A_j2EXnS4j2_1),.clk(gclk));
	jdff dff_A_Bng07JI51_1(.dout(w_n792_0[1]),.din(w_dff_A_Bng07JI51_1),.clk(gclk));
	jdff dff_A_DMRk3z007_1(.dout(w_dff_A_Bng07JI51_1),.din(w_dff_A_DMRk3z007_1),.clk(gclk));
	jdff dff_A_FPrhdtpG5_1(.dout(w_dff_A_DMRk3z007_1),.din(w_dff_A_FPrhdtpG5_1),.clk(gclk));
	jdff dff_A_kH63j8y58_1(.dout(w_dff_A_FPrhdtpG5_1),.din(w_dff_A_kH63j8y58_1),.clk(gclk));
	jdff dff_A_N3X0YXy17_1(.dout(w_dff_A_kH63j8y58_1),.din(w_dff_A_N3X0YXy17_1),.clk(gclk));
	jdff dff_A_YFE1FYKA7_1(.dout(w_dff_A_N3X0YXy17_1),.din(w_dff_A_YFE1FYKA7_1),.clk(gclk));
	jdff dff_B_G1Be0w1L8_1(.din(n1843),.dout(w_dff_B_G1Be0w1L8_1),.clk(gclk));
	jdff dff_B_BJk9Dbvo7_1(.din(n1830),.dout(w_dff_B_BJk9Dbvo7_1),.clk(gclk));
	jdff dff_B_AxN3HC4J1_1(.din(w_dff_B_BJk9Dbvo7_1),.dout(w_dff_B_AxN3HC4J1_1),.clk(gclk));
	jdff dff_B_9vMD6hbD0_2(.din(n1829),.dout(w_dff_B_9vMD6hbD0_2),.clk(gclk));
	jdff dff_B_iR3Wwocn7_2(.din(w_dff_B_9vMD6hbD0_2),.dout(w_dff_B_iR3Wwocn7_2),.clk(gclk));
	jdff dff_B_y2CLNKJg3_2(.din(w_dff_B_iR3Wwocn7_2),.dout(w_dff_B_y2CLNKJg3_2),.clk(gclk));
	jdff dff_B_thMdE1km3_2(.din(w_dff_B_y2CLNKJg3_2),.dout(w_dff_B_thMdE1km3_2),.clk(gclk));
	jdff dff_B_gqRyL4kK8_2(.din(w_dff_B_thMdE1km3_2),.dout(w_dff_B_gqRyL4kK8_2),.clk(gclk));
	jdff dff_B_2A6sBGJO0_2(.din(w_dff_B_gqRyL4kK8_2),.dout(w_dff_B_2A6sBGJO0_2),.clk(gclk));
	jdff dff_B_1FX43Tc53_2(.din(w_dff_B_2A6sBGJO0_2),.dout(w_dff_B_1FX43Tc53_2),.clk(gclk));
	jdff dff_B_6x2Ex84T7_2(.din(w_dff_B_1FX43Tc53_2),.dout(w_dff_B_6x2Ex84T7_2),.clk(gclk));
	jdff dff_B_LYPyE8tY2_2(.din(w_dff_B_6x2Ex84T7_2),.dout(w_dff_B_LYPyE8tY2_2),.clk(gclk));
	jdff dff_B_zVhitRX36_2(.din(w_dff_B_LYPyE8tY2_2),.dout(w_dff_B_zVhitRX36_2),.clk(gclk));
	jdff dff_B_mtiAUmNd6_2(.din(w_dff_B_zVhitRX36_2),.dout(w_dff_B_mtiAUmNd6_2),.clk(gclk));
	jdff dff_B_7SoSryC90_2(.din(w_dff_B_mtiAUmNd6_2),.dout(w_dff_B_7SoSryC90_2),.clk(gclk));
	jdff dff_B_fP3eqyak0_2(.din(w_dff_B_7SoSryC90_2),.dout(w_dff_B_fP3eqyak0_2),.clk(gclk));
	jdff dff_B_njOaAzGI0_2(.din(w_dff_B_fP3eqyak0_2),.dout(w_dff_B_njOaAzGI0_2),.clk(gclk));
	jdff dff_B_7tPl8Cjy8_2(.din(w_dff_B_njOaAzGI0_2),.dout(w_dff_B_7tPl8Cjy8_2),.clk(gclk));
	jdff dff_B_v8BIbjAg8_2(.din(w_dff_B_7tPl8Cjy8_2),.dout(w_dff_B_v8BIbjAg8_2),.clk(gclk));
	jdff dff_B_StLRGRLP9_2(.din(w_dff_B_v8BIbjAg8_2),.dout(w_dff_B_StLRGRLP9_2),.clk(gclk));
	jdff dff_B_QfVDqDwH8_2(.din(w_dff_B_StLRGRLP9_2),.dout(w_dff_B_QfVDqDwH8_2),.clk(gclk));
	jdff dff_B_B3KWInmO7_2(.din(w_dff_B_QfVDqDwH8_2),.dout(w_dff_B_B3KWInmO7_2),.clk(gclk));
	jdff dff_B_M7DCY9k03_2(.din(w_dff_B_B3KWInmO7_2),.dout(w_dff_B_M7DCY9k03_2),.clk(gclk));
	jdff dff_B_rAUwfWYI2_2(.din(w_dff_B_M7DCY9k03_2),.dout(w_dff_B_rAUwfWYI2_2),.clk(gclk));
	jdff dff_B_52iviQen5_2(.din(w_dff_B_rAUwfWYI2_2),.dout(w_dff_B_52iviQen5_2),.clk(gclk));
	jdff dff_B_nYhK47Pe4_2(.din(w_dff_B_52iviQen5_2),.dout(w_dff_B_nYhK47Pe4_2),.clk(gclk));
	jdff dff_B_ETSoEChk3_2(.din(w_dff_B_nYhK47Pe4_2),.dout(w_dff_B_ETSoEChk3_2),.clk(gclk));
	jdff dff_B_wJZ6jOMz5_2(.din(w_dff_B_ETSoEChk3_2),.dout(w_dff_B_wJZ6jOMz5_2),.clk(gclk));
	jdff dff_B_MnNlc0Ou7_2(.din(w_dff_B_wJZ6jOMz5_2),.dout(w_dff_B_MnNlc0Ou7_2),.clk(gclk));
	jdff dff_B_tEmivrTT0_2(.din(w_dff_B_MnNlc0Ou7_2),.dout(w_dff_B_tEmivrTT0_2),.clk(gclk));
	jdff dff_B_cE7dGaTG7_2(.din(w_dff_B_tEmivrTT0_2),.dout(w_dff_B_cE7dGaTG7_2),.clk(gclk));
	jdff dff_B_eBmY3vh63_2(.din(w_dff_B_cE7dGaTG7_2),.dout(w_dff_B_eBmY3vh63_2),.clk(gclk));
	jdff dff_B_UqrvQW5a4_2(.din(w_dff_B_eBmY3vh63_2),.dout(w_dff_B_UqrvQW5a4_2),.clk(gclk));
	jdff dff_B_9S1WPhc23_2(.din(w_dff_B_UqrvQW5a4_2),.dout(w_dff_B_9S1WPhc23_2),.clk(gclk));
	jdff dff_B_sgCui1Oh6_2(.din(w_dff_B_9S1WPhc23_2),.dout(w_dff_B_sgCui1Oh6_2),.clk(gclk));
	jdff dff_B_dFFw3xfX4_2(.din(w_dff_B_sgCui1Oh6_2),.dout(w_dff_B_dFFw3xfX4_2),.clk(gclk));
	jdff dff_B_KykwPUDp1_2(.din(w_dff_B_dFFw3xfX4_2),.dout(w_dff_B_KykwPUDp1_2),.clk(gclk));
	jdff dff_B_6nFXMZBp9_2(.din(w_dff_B_KykwPUDp1_2),.dout(w_dff_B_6nFXMZBp9_2),.clk(gclk));
	jdff dff_B_Q4CBMmkC9_2(.din(w_dff_B_6nFXMZBp9_2),.dout(w_dff_B_Q4CBMmkC9_2),.clk(gclk));
	jdff dff_B_UC5kuJaV0_2(.din(w_dff_B_Q4CBMmkC9_2),.dout(w_dff_B_UC5kuJaV0_2),.clk(gclk));
	jdff dff_B_1fdUktiK4_2(.din(w_dff_B_UC5kuJaV0_2),.dout(w_dff_B_1fdUktiK4_2),.clk(gclk));
	jdff dff_B_Pmflzgv54_2(.din(w_dff_B_1fdUktiK4_2),.dout(w_dff_B_Pmflzgv54_2),.clk(gclk));
	jdff dff_B_zhUTe2rp2_2(.din(w_dff_B_Pmflzgv54_2),.dout(w_dff_B_zhUTe2rp2_2),.clk(gclk));
	jdff dff_B_D2PBaTFe8_2(.din(w_dff_B_zhUTe2rp2_2),.dout(w_dff_B_D2PBaTFe8_2),.clk(gclk));
	jdff dff_B_sH9z1PyZ3_2(.din(w_dff_B_D2PBaTFe8_2),.dout(w_dff_B_sH9z1PyZ3_2),.clk(gclk));
	jdff dff_B_MvYL5r789_2(.din(w_dff_B_sH9z1PyZ3_2),.dout(w_dff_B_MvYL5r789_2),.clk(gclk));
	jdff dff_B_5BFebvs10_2(.din(w_dff_B_MvYL5r789_2),.dout(w_dff_B_5BFebvs10_2),.clk(gclk));
	jdff dff_B_PULcOqeB0_2(.din(w_dff_B_5BFebvs10_2),.dout(w_dff_B_PULcOqeB0_2),.clk(gclk));
	jdff dff_B_gXqmDAeT8_2(.din(w_dff_B_PULcOqeB0_2),.dout(w_dff_B_gXqmDAeT8_2),.clk(gclk));
	jdff dff_B_xgFFtDeH6_2(.din(w_dff_B_gXqmDAeT8_2),.dout(w_dff_B_xgFFtDeH6_2),.clk(gclk));
	jdff dff_B_3H1iyCRn6_2(.din(w_dff_B_xgFFtDeH6_2),.dout(w_dff_B_3H1iyCRn6_2),.clk(gclk));
	jdff dff_B_06s29llU5_2(.din(w_dff_B_3H1iyCRn6_2),.dout(w_dff_B_06s29llU5_2),.clk(gclk));
	jdff dff_B_NCg4KGXy8_2(.din(w_dff_B_06s29llU5_2),.dout(w_dff_B_NCg4KGXy8_2),.clk(gclk));
	jdff dff_B_aDtcJ0ba2_2(.din(w_dff_B_NCg4KGXy8_2),.dout(w_dff_B_aDtcJ0ba2_2),.clk(gclk));
	jdff dff_B_DBu9MS8x8_2(.din(w_dff_B_aDtcJ0ba2_2),.dout(w_dff_B_DBu9MS8x8_2),.clk(gclk));
	jdff dff_B_WqK2XOQa0_2(.din(w_dff_B_DBu9MS8x8_2),.dout(w_dff_B_WqK2XOQa0_2),.clk(gclk));
	jdff dff_B_K12XMtUH4_2(.din(w_dff_B_WqK2XOQa0_2),.dout(w_dff_B_K12XMtUH4_2),.clk(gclk));
	jdff dff_B_NX47Qo9X3_2(.din(w_dff_B_K12XMtUH4_2),.dout(w_dff_B_NX47Qo9X3_2),.clk(gclk));
	jdff dff_B_1EHsxoj72_2(.din(w_dff_B_NX47Qo9X3_2),.dout(w_dff_B_1EHsxoj72_2),.clk(gclk));
	jdff dff_B_XFzugYOA1_2(.din(n1828),.dout(w_dff_B_XFzugYOA1_2),.clk(gclk));
	jdff dff_B_T28lCIe81_2(.din(w_dff_B_XFzugYOA1_2),.dout(w_dff_B_T28lCIe81_2),.clk(gclk));
	jdff dff_B_wkflulbq7_2(.din(w_dff_B_T28lCIe81_2),.dout(w_dff_B_wkflulbq7_2),.clk(gclk));
	jdff dff_B_U5frjtpA6_2(.din(w_dff_B_wkflulbq7_2),.dout(w_dff_B_U5frjtpA6_2),.clk(gclk));
	jdff dff_B_O6i7BYTM1_2(.din(w_dff_B_U5frjtpA6_2),.dout(w_dff_B_O6i7BYTM1_2),.clk(gclk));
	jdff dff_B_rwByXSln1_2(.din(w_dff_B_O6i7BYTM1_2),.dout(w_dff_B_rwByXSln1_2),.clk(gclk));
	jdff dff_B_rtwrQ7Tv5_2(.din(w_dff_B_rwByXSln1_2),.dout(w_dff_B_rtwrQ7Tv5_2),.clk(gclk));
	jdff dff_B_HDbnImm39_2(.din(w_dff_B_rtwrQ7Tv5_2),.dout(w_dff_B_HDbnImm39_2),.clk(gclk));
	jdff dff_B_AaMS8tfn6_2(.din(w_dff_B_HDbnImm39_2),.dout(w_dff_B_AaMS8tfn6_2),.clk(gclk));
	jdff dff_B_pVk1HtIl5_2(.din(w_dff_B_AaMS8tfn6_2),.dout(w_dff_B_pVk1HtIl5_2),.clk(gclk));
	jdff dff_B_FAc6RLLw4_2(.din(w_dff_B_pVk1HtIl5_2),.dout(w_dff_B_FAc6RLLw4_2),.clk(gclk));
	jdff dff_B_1TFpC6D21_2(.din(w_dff_B_FAc6RLLw4_2),.dout(w_dff_B_1TFpC6D21_2),.clk(gclk));
	jdff dff_B_PfAeb9oB3_2(.din(w_dff_B_1TFpC6D21_2),.dout(w_dff_B_PfAeb9oB3_2),.clk(gclk));
	jdff dff_B_MVQii1Gd8_2(.din(w_dff_B_PfAeb9oB3_2),.dout(w_dff_B_MVQii1Gd8_2),.clk(gclk));
	jdff dff_B_Djsn6kpn7_2(.din(w_dff_B_MVQii1Gd8_2),.dout(w_dff_B_Djsn6kpn7_2),.clk(gclk));
	jdff dff_B_xexikIMK3_2(.din(w_dff_B_Djsn6kpn7_2),.dout(w_dff_B_xexikIMK3_2),.clk(gclk));
	jdff dff_B_ggMbpQ1Y0_2(.din(w_dff_B_xexikIMK3_2),.dout(w_dff_B_ggMbpQ1Y0_2),.clk(gclk));
	jdff dff_B_vCgWseQY3_2(.din(w_dff_B_ggMbpQ1Y0_2),.dout(w_dff_B_vCgWseQY3_2),.clk(gclk));
	jdff dff_B_JdEPa84d2_2(.din(w_dff_B_vCgWseQY3_2),.dout(w_dff_B_JdEPa84d2_2),.clk(gclk));
	jdff dff_B_4BkPHsBH0_2(.din(w_dff_B_JdEPa84d2_2),.dout(w_dff_B_4BkPHsBH0_2),.clk(gclk));
	jdff dff_B_vHAFnp5x2_2(.din(w_dff_B_4BkPHsBH0_2),.dout(w_dff_B_vHAFnp5x2_2),.clk(gclk));
	jdff dff_B_nBcdnM9J5_2(.din(w_dff_B_vHAFnp5x2_2),.dout(w_dff_B_nBcdnM9J5_2),.clk(gclk));
	jdff dff_B_mqHpdWmB4_2(.din(w_dff_B_nBcdnM9J5_2),.dout(w_dff_B_mqHpdWmB4_2),.clk(gclk));
	jdff dff_B_XxhIOBW03_2(.din(w_dff_B_mqHpdWmB4_2),.dout(w_dff_B_XxhIOBW03_2),.clk(gclk));
	jdff dff_B_YerTaQ5M3_2(.din(w_dff_B_XxhIOBW03_2),.dout(w_dff_B_YerTaQ5M3_2),.clk(gclk));
	jdff dff_B_5qeh0qTg4_2(.din(w_dff_B_YerTaQ5M3_2),.dout(w_dff_B_5qeh0qTg4_2),.clk(gclk));
	jdff dff_B_N5mK56Ne9_2(.din(w_dff_B_5qeh0qTg4_2),.dout(w_dff_B_N5mK56Ne9_2),.clk(gclk));
	jdff dff_B_YvHSALV81_2(.din(w_dff_B_N5mK56Ne9_2),.dout(w_dff_B_YvHSALV81_2),.clk(gclk));
	jdff dff_B_SVjep5Kl0_2(.din(w_dff_B_YvHSALV81_2),.dout(w_dff_B_SVjep5Kl0_2),.clk(gclk));
	jdff dff_B_i2mWbpK86_2(.din(w_dff_B_SVjep5Kl0_2),.dout(w_dff_B_i2mWbpK86_2),.clk(gclk));
	jdff dff_B_FxwMyqUs3_2(.din(w_dff_B_i2mWbpK86_2),.dout(w_dff_B_FxwMyqUs3_2),.clk(gclk));
	jdff dff_B_cxmOkPJ61_2(.din(w_dff_B_FxwMyqUs3_2),.dout(w_dff_B_cxmOkPJ61_2),.clk(gclk));
	jdff dff_B_dyIoaoXw8_2(.din(w_dff_B_cxmOkPJ61_2),.dout(w_dff_B_dyIoaoXw8_2),.clk(gclk));
	jdff dff_B_SflPcyWR9_2(.din(w_dff_B_dyIoaoXw8_2),.dout(w_dff_B_SflPcyWR9_2),.clk(gclk));
	jdff dff_B_jrItXETU6_2(.din(w_dff_B_SflPcyWR9_2),.dout(w_dff_B_jrItXETU6_2),.clk(gclk));
	jdff dff_B_WK2EgIWG3_2(.din(w_dff_B_jrItXETU6_2),.dout(w_dff_B_WK2EgIWG3_2),.clk(gclk));
	jdff dff_B_xFAOHMdw9_2(.din(w_dff_B_WK2EgIWG3_2),.dout(w_dff_B_xFAOHMdw9_2),.clk(gclk));
	jdff dff_B_dhnAj0hT9_2(.din(w_dff_B_xFAOHMdw9_2),.dout(w_dff_B_dhnAj0hT9_2),.clk(gclk));
	jdff dff_B_QTDhhjWn0_2(.din(w_dff_B_dhnAj0hT9_2),.dout(w_dff_B_QTDhhjWn0_2),.clk(gclk));
	jdff dff_B_lN3EfoVL0_2(.din(w_dff_B_QTDhhjWn0_2),.dout(w_dff_B_lN3EfoVL0_2),.clk(gclk));
	jdff dff_B_8s5o3v5U4_2(.din(w_dff_B_lN3EfoVL0_2),.dout(w_dff_B_8s5o3v5U4_2),.clk(gclk));
	jdff dff_B_qde6tAky2_2(.din(w_dff_B_8s5o3v5U4_2),.dout(w_dff_B_qde6tAky2_2),.clk(gclk));
	jdff dff_B_In3gVkjm5_2(.din(w_dff_B_qde6tAky2_2),.dout(w_dff_B_In3gVkjm5_2),.clk(gclk));
	jdff dff_B_STu83squ6_2(.din(w_dff_B_In3gVkjm5_2),.dout(w_dff_B_STu83squ6_2),.clk(gclk));
	jdff dff_B_gfdF8Odu5_2(.din(w_dff_B_STu83squ6_2),.dout(w_dff_B_gfdF8Odu5_2),.clk(gclk));
	jdff dff_B_oyiBnt7S7_2(.din(w_dff_B_gfdF8Odu5_2),.dout(w_dff_B_oyiBnt7S7_2),.clk(gclk));
	jdff dff_B_ix5DV3Pj9_2(.din(w_dff_B_oyiBnt7S7_2),.dout(w_dff_B_ix5DV3Pj9_2),.clk(gclk));
	jdff dff_B_DQziWUWh7_2(.din(w_dff_B_ix5DV3Pj9_2),.dout(w_dff_B_DQziWUWh7_2),.clk(gclk));
	jdff dff_B_tKKdVf3h6_2(.din(w_dff_B_DQziWUWh7_2),.dout(w_dff_B_tKKdVf3h6_2),.clk(gclk));
	jdff dff_B_ZnvyxNqF0_2(.din(w_dff_B_tKKdVf3h6_2),.dout(w_dff_B_ZnvyxNqF0_2),.clk(gclk));
	jdff dff_B_bVUR7K3M1_2(.din(w_dff_B_ZnvyxNqF0_2),.dout(w_dff_B_bVUR7K3M1_2),.clk(gclk));
	jdff dff_B_NfQ7qjpF1_2(.din(w_dff_B_bVUR7K3M1_2),.dout(w_dff_B_NfQ7qjpF1_2),.clk(gclk));
	jdff dff_B_KvjGBq3E4_2(.din(w_dff_B_NfQ7qjpF1_2),.dout(w_dff_B_KvjGBq3E4_2),.clk(gclk));
	jdff dff_B_PFWPYXhD6_2(.din(w_dff_B_KvjGBq3E4_2),.dout(w_dff_B_PFWPYXhD6_2),.clk(gclk));
	jdff dff_B_JwSfpbBe7_2(.din(w_dff_B_PFWPYXhD6_2),.dout(w_dff_B_JwSfpbBe7_2),.clk(gclk));
	jdff dff_B_JRF5aHui3_2(.din(w_dff_B_JwSfpbBe7_2),.dout(w_dff_B_JRF5aHui3_2),.clk(gclk));
	jdff dff_B_n6ngT6Yo2_2(.din(w_dff_B_JRF5aHui3_2),.dout(w_dff_B_n6ngT6Yo2_2),.clk(gclk));
	jdff dff_B_eP2sF8fc1_2(.din(w_dff_B_n6ngT6Yo2_2),.dout(w_dff_B_eP2sF8fc1_2),.clk(gclk));
	jdff dff_A_Gl0YM9RQ1_1(.dout(w_n1827_0[1]),.din(w_dff_A_Gl0YM9RQ1_1),.clk(gclk));
	jdff dff_B_mgjKK9GJ3_1(.din(n1825),.dout(w_dff_B_mgjKK9GJ3_1),.clk(gclk));
	jdff dff_B_SCL5FPKf3_2(.din(n1803),.dout(w_dff_B_SCL5FPKf3_2),.clk(gclk));
	jdff dff_B_rzXmh0BJ1_2(.din(w_dff_B_SCL5FPKf3_2),.dout(w_dff_B_rzXmh0BJ1_2),.clk(gclk));
	jdff dff_B_qeZt0Tgx5_2(.din(w_dff_B_rzXmh0BJ1_2),.dout(w_dff_B_qeZt0Tgx5_2),.clk(gclk));
	jdff dff_B_f3WvnnPU4_2(.din(w_dff_B_qeZt0Tgx5_2),.dout(w_dff_B_f3WvnnPU4_2),.clk(gclk));
	jdff dff_B_NyTNzeqe7_2(.din(w_dff_B_f3WvnnPU4_2),.dout(w_dff_B_NyTNzeqe7_2),.clk(gclk));
	jdff dff_B_bu82JbmM1_2(.din(w_dff_B_NyTNzeqe7_2),.dout(w_dff_B_bu82JbmM1_2),.clk(gclk));
	jdff dff_B_PtMZMIJq2_2(.din(w_dff_B_bu82JbmM1_2),.dout(w_dff_B_PtMZMIJq2_2),.clk(gclk));
	jdff dff_B_iAqmL0DB6_2(.din(w_dff_B_PtMZMIJq2_2),.dout(w_dff_B_iAqmL0DB6_2),.clk(gclk));
	jdff dff_B_ljIttL9l9_2(.din(w_dff_B_iAqmL0DB6_2),.dout(w_dff_B_ljIttL9l9_2),.clk(gclk));
	jdff dff_B_nxCSWGlt7_2(.din(w_dff_B_ljIttL9l9_2),.dout(w_dff_B_nxCSWGlt7_2),.clk(gclk));
	jdff dff_B_qwNFtUbC2_2(.din(w_dff_B_nxCSWGlt7_2),.dout(w_dff_B_qwNFtUbC2_2),.clk(gclk));
	jdff dff_B_eX9ZyAfw3_2(.din(w_dff_B_qwNFtUbC2_2),.dout(w_dff_B_eX9ZyAfw3_2),.clk(gclk));
	jdff dff_B_d40C5jOH5_2(.din(w_dff_B_eX9ZyAfw3_2),.dout(w_dff_B_d40C5jOH5_2),.clk(gclk));
	jdff dff_B_QYCke47w0_2(.din(w_dff_B_d40C5jOH5_2),.dout(w_dff_B_QYCke47w0_2),.clk(gclk));
	jdff dff_B_O7ZtqB7H8_2(.din(w_dff_B_QYCke47w0_2),.dout(w_dff_B_O7ZtqB7H8_2),.clk(gclk));
	jdff dff_B_buJwVWIL1_2(.din(w_dff_B_O7ZtqB7H8_2),.dout(w_dff_B_buJwVWIL1_2),.clk(gclk));
	jdff dff_B_4wdRDvXP7_2(.din(w_dff_B_buJwVWIL1_2),.dout(w_dff_B_4wdRDvXP7_2),.clk(gclk));
	jdff dff_B_M027ArTJ2_2(.din(w_dff_B_4wdRDvXP7_2),.dout(w_dff_B_M027ArTJ2_2),.clk(gclk));
	jdff dff_B_IgbOy04R6_2(.din(w_dff_B_M027ArTJ2_2),.dout(w_dff_B_IgbOy04R6_2),.clk(gclk));
	jdff dff_B_JKKOcUY14_2(.din(w_dff_B_IgbOy04R6_2),.dout(w_dff_B_JKKOcUY14_2),.clk(gclk));
	jdff dff_B_uOyyPRu64_2(.din(w_dff_B_JKKOcUY14_2),.dout(w_dff_B_uOyyPRu64_2),.clk(gclk));
	jdff dff_B_Qq5pQ5Py1_2(.din(w_dff_B_uOyyPRu64_2),.dout(w_dff_B_Qq5pQ5Py1_2),.clk(gclk));
	jdff dff_B_RNL4Jt5w8_2(.din(w_dff_B_Qq5pQ5Py1_2),.dout(w_dff_B_RNL4Jt5w8_2),.clk(gclk));
	jdff dff_B_mDVG1MSg6_2(.din(w_dff_B_RNL4Jt5w8_2),.dout(w_dff_B_mDVG1MSg6_2),.clk(gclk));
	jdff dff_B_qPSvWAOh0_2(.din(w_dff_B_mDVG1MSg6_2),.dout(w_dff_B_qPSvWAOh0_2),.clk(gclk));
	jdff dff_B_0OTCxfDP5_2(.din(w_dff_B_qPSvWAOh0_2),.dout(w_dff_B_0OTCxfDP5_2),.clk(gclk));
	jdff dff_B_e3nTQoLs9_2(.din(w_dff_B_0OTCxfDP5_2),.dout(w_dff_B_e3nTQoLs9_2),.clk(gclk));
	jdff dff_B_tpHaKlcI8_2(.din(w_dff_B_e3nTQoLs9_2),.dout(w_dff_B_tpHaKlcI8_2),.clk(gclk));
	jdff dff_B_2ux7tTVC2_2(.din(w_dff_B_tpHaKlcI8_2),.dout(w_dff_B_2ux7tTVC2_2),.clk(gclk));
	jdff dff_B_pVz0MthM3_2(.din(w_dff_B_2ux7tTVC2_2),.dout(w_dff_B_pVz0MthM3_2),.clk(gclk));
	jdff dff_B_xpITjV6J8_2(.din(w_dff_B_pVz0MthM3_2),.dout(w_dff_B_xpITjV6J8_2),.clk(gclk));
	jdff dff_B_zCFukkEW2_2(.din(w_dff_B_xpITjV6J8_2),.dout(w_dff_B_zCFukkEW2_2),.clk(gclk));
	jdff dff_B_6GVByEGo9_2(.din(w_dff_B_zCFukkEW2_2),.dout(w_dff_B_6GVByEGo9_2),.clk(gclk));
	jdff dff_B_PzF4wiI91_2(.din(w_dff_B_6GVByEGo9_2),.dout(w_dff_B_PzF4wiI91_2),.clk(gclk));
	jdff dff_B_PZRbMNPF1_2(.din(w_dff_B_PzF4wiI91_2),.dout(w_dff_B_PZRbMNPF1_2),.clk(gclk));
	jdff dff_B_wE8M9pSE6_2(.din(w_dff_B_PZRbMNPF1_2),.dout(w_dff_B_wE8M9pSE6_2),.clk(gclk));
	jdff dff_B_sxF7Nnto4_2(.din(w_dff_B_wE8M9pSE6_2),.dout(w_dff_B_sxF7Nnto4_2),.clk(gclk));
	jdff dff_B_0s4hG60m4_2(.din(w_dff_B_sxF7Nnto4_2),.dout(w_dff_B_0s4hG60m4_2),.clk(gclk));
	jdff dff_B_5h7NepSj5_2(.din(w_dff_B_0s4hG60m4_2),.dout(w_dff_B_5h7NepSj5_2),.clk(gclk));
	jdff dff_B_pop4QW1h9_2(.din(w_dff_B_5h7NepSj5_2),.dout(w_dff_B_pop4QW1h9_2),.clk(gclk));
	jdff dff_B_upAQuHGD9_2(.din(w_dff_B_pop4QW1h9_2),.dout(w_dff_B_upAQuHGD9_2),.clk(gclk));
	jdff dff_B_vnGnmv5D6_2(.din(w_dff_B_upAQuHGD9_2),.dout(w_dff_B_vnGnmv5D6_2),.clk(gclk));
	jdff dff_B_WsEJNZR41_2(.din(w_dff_B_vnGnmv5D6_2),.dout(w_dff_B_WsEJNZR41_2),.clk(gclk));
	jdff dff_B_t8NUpRFL8_2(.din(w_dff_B_WsEJNZR41_2),.dout(w_dff_B_t8NUpRFL8_2),.clk(gclk));
	jdff dff_B_n4UBlc7K0_2(.din(w_dff_B_t8NUpRFL8_2),.dout(w_dff_B_n4UBlc7K0_2),.clk(gclk));
	jdff dff_B_9QpmV5qC5_2(.din(w_dff_B_n4UBlc7K0_2),.dout(w_dff_B_9QpmV5qC5_2),.clk(gclk));
	jdff dff_B_LTNHYBTm5_2(.din(w_dff_B_9QpmV5qC5_2),.dout(w_dff_B_LTNHYBTm5_2),.clk(gclk));
	jdff dff_B_yZxKMZrc0_2(.din(w_dff_B_LTNHYBTm5_2),.dout(w_dff_B_yZxKMZrc0_2),.clk(gclk));
	jdff dff_B_t5UhvOzR9_2(.din(w_dff_B_yZxKMZrc0_2),.dout(w_dff_B_t5UhvOzR9_2),.clk(gclk));
	jdff dff_B_u4xfTwzc5_2(.din(w_dff_B_t5UhvOzR9_2),.dout(w_dff_B_u4xfTwzc5_2),.clk(gclk));
	jdff dff_B_f5WMARNu2_2(.din(w_dff_B_u4xfTwzc5_2),.dout(w_dff_B_f5WMARNu2_2),.clk(gclk));
	jdff dff_B_kqOINCaK6_2(.din(w_dff_B_f5WMARNu2_2),.dout(w_dff_B_kqOINCaK6_2),.clk(gclk));
	jdff dff_B_pZhfJMe73_2(.din(w_dff_B_kqOINCaK6_2),.dout(w_dff_B_pZhfJMe73_2),.clk(gclk));
	jdff dff_B_DDLXVTVi5_2(.din(w_dff_B_pZhfJMe73_2),.dout(w_dff_B_DDLXVTVi5_2),.clk(gclk));
	jdff dff_B_iy3NUKPE5_2(.din(w_dff_B_DDLXVTVi5_2),.dout(w_dff_B_iy3NUKPE5_2),.clk(gclk));
	jdff dff_B_C5PFZR9b4_1(.din(n1809),.dout(w_dff_B_C5PFZR9b4_1),.clk(gclk));
	jdff dff_B_HF7UIH5v7_1(.din(w_dff_B_C5PFZR9b4_1),.dout(w_dff_B_HF7UIH5v7_1),.clk(gclk));
	jdff dff_B_wHsykZ4H0_2(.din(n1808),.dout(w_dff_B_wHsykZ4H0_2),.clk(gclk));
	jdff dff_B_zhuPOkfj8_2(.din(w_dff_B_wHsykZ4H0_2),.dout(w_dff_B_zhuPOkfj8_2),.clk(gclk));
	jdff dff_B_0XaTQvYi4_2(.din(w_dff_B_zhuPOkfj8_2),.dout(w_dff_B_0XaTQvYi4_2),.clk(gclk));
	jdff dff_B_yDLhR7300_2(.din(w_dff_B_0XaTQvYi4_2),.dout(w_dff_B_yDLhR7300_2),.clk(gclk));
	jdff dff_B_Eex5LyVM5_2(.din(w_dff_B_yDLhR7300_2),.dout(w_dff_B_Eex5LyVM5_2),.clk(gclk));
	jdff dff_B_6ZvvSzvv7_2(.din(w_dff_B_Eex5LyVM5_2),.dout(w_dff_B_6ZvvSzvv7_2),.clk(gclk));
	jdff dff_B_U9JaiPV90_2(.din(w_dff_B_6ZvvSzvv7_2),.dout(w_dff_B_U9JaiPV90_2),.clk(gclk));
	jdff dff_B_3HEWHJvJ7_2(.din(w_dff_B_U9JaiPV90_2),.dout(w_dff_B_3HEWHJvJ7_2),.clk(gclk));
	jdff dff_B_5tC6oTRG6_2(.din(w_dff_B_3HEWHJvJ7_2),.dout(w_dff_B_5tC6oTRG6_2),.clk(gclk));
	jdff dff_B_kaXIRbLv3_2(.din(w_dff_B_5tC6oTRG6_2),.dout(w_dff_B_kaXIRbLv3_2),.clk(gclk));
	jdff dff_B_CP6JXgNu9_2(.din(w_dff_B_kaXIRbLv3_2),.dout(w_dff_B_CP6JXgNu9_2),.clk(gclk));
	jdff dff_B_gzs4q0lq2_2(.din(w_dff_B_CP6JXgNu9_2),.dout(w_dff_B_gzs4q0lq2_2),.clk(gclk));
	jdff dff_B_3esntLel3_2(.din(w_dff_B_gzs4q0lq2_2),.dout(w_dff_B_3esntLel3_2),.clk(gclk));
	jdff dff_B_V4mb45DA0_2(.din(w_dff_B_3esntLel3_2),.dout(w_dff_B_V4mb45DA0_2),.clk(gclk));
	jdff dff_B_BelUqyhy5_2(.din(w_dff_B_V4mb45DA0_2),.dout(w_dff_B_BelUqyhy5_2),.clk(gclk));
	jdff dff_B_6H5KFKj60_2(.din(w_dff_B_BelUqyhy5_2),.dout(w_dff_B_6H5KFKj60_2),.clk(gclk));
	jdff dff_B_s8QpbDgg2_2(.din(w_dff_B_6H5KFKj60_2),.dout(w_dff_B_s8QpbDgg2_2),.clk(gclk));
	jdff dff_B_U7g7E0915_2(.din(w_dff_B_s8QpbDgg2_2),.dout(w_dff_B_U7g7E0915_2),.clk(gclk));
	jdff dff_B_HQwyle1y5_2(.din(w_dff_B_U7g7E0915_2),.dout(w_dff_B_HQwyle1y5_2),.clk(gclk));
	jdff dff_B_0TwLzO5A5_2(.din(w_dff_B_HQwyle1y5_2),.dout(w_dff_B_0TwLzO5A5_2),.clk(gclk));
	jdff dff_B_jmKALU6T0_2(.din(w_dff_B_0TwLzO5A5_2),.dout(w_dff_B_jmKALU6T0_2),.clk(gclk));
	jdff dff_B_eBUFuLKM9_2(.din(w_dff_B_jmKALU6T0_2),.dout(w_dff_B_eBUFuLKM9_2),.clk(gclk));
	jdff dff_B_33O9jhYA3_2(.din(w_dff_B_eBUFuLKM9_2),.dout(w_dff_B_33O9jhYA3_2),.clk(gclk));
	jdff dff_B_YJDYGVz93_2(.din(w_dff_B_33O9jhYA3_2),.dout(w_dff_B_YJDYGVz93_2),.clk(gclk));
	jdff dff_B_pG3Im42M8_2(.din(w_dff_B_YJDYGVz93_2),.dout(w_dff_B_pG3Im42M8_2),.clk(gclk));
	jdff dff_B_IST5TWf49_2(.din(w_dff_B_pG3Im42M8_2),.dout(w_dff_B_IST5TWf49_2),.clk(gclk));
	jdff dff_B_Tl1UPHVz1_2(.din(w_dff_B_IST5TWf49_2),.dout(w_dff_B_Tl1UPHVz1_2),.clk(gclk));
	jdff dff_B_oNE4NWWT9_2(.din(w_dff_B_Tl1UPHVz1_2),.dout(w_dff_B_oNE4NWWT9_2),.clk(gclk));
	jdff dff_B_lyFbzixm0_2(.din(w_dff_B_oNE4NWWT9_2),.dout(w_dff_B_lyFbzixm0_2),.clk(gclk));
	jdff dff_B_TocHg3WY7_2(.din(w_dff_B_lyFbzixm0_2),.dout(w_dff_B_TocHg3WY7_2),.clk(gclk));
	jdff dff_B_3cBaZWW75_2(.din(w_dff_B_TocHg3WY7_2),.dout(w_dff_B_3cBaZWW75_2),.clk(gclk));
	jdff dff_B_SDyoQ5iT4_2(.din(w_dff_B_3cBaZWW75_2),.dout(w_dff_B_SDyoQ5iT4_2),.clk(gclk));
	jdff dff_B_64TKNjo47_2(.din(w_dff_B_SDyoQ5iT4_2),.dout(w_dff_B_64TKNjo47_2),.clk(gclk));
	jdff dff_B_uyHq7NzC1_2(.din(w_dff_B_64TKNjo47_2),.dout(w_dff_B_uyHq7NzC1_2),.clk(gclk));
	jdff dff_B_ZoiUq8a02_2(.din(w_dff_B_uyHq7NzC1_2),.dout(w_dff_B_ZoiUq8a02_2),.clk(gclk));
	jdff dff_B_Ba850tM69_2(.din(w_dff_B_ZoiUq8a02_2),.dout(w_dff_B_Ba850tM69_2),.clk(gclk));
	jdff dff_B_mnXNmXzB8_2(.din(w_dff_B_Ba850tM69_2),.dout(w_dff_B_mnXNmXzB8_2),.clk(gclk));
	jdff dff_B_4gS6xnRA7_2(.din(w_dff_B_mnXNmXzB8_2),.dout(w_dff_B_4gS6xnRA7_2),.clk(gclk));
	jdff dff_B_EbhUxANj2_2(.din(w_dff_B_4gS6xnRA7_2),.dout(w_dff_B_EbhUxANj2_2),.clk(gclk));
	jdff dff_B_vuE5VV8D4_2(.din(w_dff_B_EbhUxANj2_2),.dout(w_dff_B_vuE5VV8D4_2),.clk(gclk));
	jdff dff_B_eT333xhz5_2(.din(w_dff_B_vuE5VV8D4_2),.dout(w_dff_B_eT333xhz5_2),.clk(gclk));
	jdff dff_B_467KL0ma9_2(.din(w_dff_B_eT333xhz5_2),.dout(w_dff_B_467KL0ma9_2),.clk(gclk));
	jdff dff_B_0qy5Wpy23_2(.din(w_dff_B_467KL0ma9_2),.dout(w_dff_B_0qy5Wpy23_2),.clk(gclk));
	jdff dff_B_eFqEJzwg6_2(.din(w_dff_B_0qy5Wpy23_2),.dout(w_dff_B_eFqEJzwg6_2),.clk(gclk));
	jdff dff_B_a8QS7p6D1_2(.din(w_dff_B_eFqEJzwg6_2),.dout(w_dff_B_a8QS7p6D1_2),.clk(gclk));
	jdff dff_B_QPsg3qiV0_2(.din(w_dff_B_a8QS7p6D1_2),.dout(w_dff_B_QPsg3qiV0_2),.clk(gclk));
	jdff dff_B_VjQUnkm02_2(.din(w_dff_B_QPsg3qiV0_2),.dout(w_dff_B_VjQUnkm02_2),.clk(gclk));
	jdff dff_B_Xv7fqjh14_2(.din(w_dff_B_VjQUnkm02_2),.dout(w_dff_B_Xv7fqjh14_2),.clk(gclk));
	jdff dff_B_KY5ozMdg9_2(.din(w_dff_B_Xv7fqjh14_2),.dout(w_dff_B_KY5ozMdg9_2),.clk(gclk));
	jdff dff_B_fD031rCq7_2(.din(w_dff_B_KY5ozMdg9_2),.dout(w_dff_B_fD031rCq7_2),.clk(gclk));
	jdff dff_B_E57eyS4L2_2(.din(w_dff_B_fD031rCq7_2),.dout(w_dff_B_E57eyS4L2_2),.clk(gclk));
	jdff dff_B_qDLH0N856_2(.din(w_dff_B_E57eyS4L2_2),.dout(w_dff_B_qDLH0N856_2),.clk(gclk));
	jdff dff_B_2fPJuVhx8_2(.din(n1807),.dout(w_dff_B_2fPJuVhx8_2),.clk(gclk));
	jdff dff_B_7dzdvXTd5_2(.din(w_dff_B_2fPJuVhx8_2),.dout(w_dff_B_7dzdvXTd5_2),.clk(gclk));
	jdff dff_B_0VyNcSpR3_2(.din(w_dff_B_7dzdvXTd5_2),.dout(w_dff_B_0VyNcSpR3_2),.clk(gclk));
	jdff dff_B_1P0ZU3AO1_2(.din(w_dff_B_0VyNcSpR3_2),.dout(w_dff_B_1P0ZU3AO1_2),.clk(gclk));
	jdff dff_B_9eR9o1238_2(.din(w_dff_B_1P0ZU3AO1_2),.dout(w_dff_B_9eR9o1238_2),.clk(gclk));
	jdff dff_B_Lt9yd9Dk1_2(.din(w_dff_B_9eR9o1238_2),.dout(w_dff_B_Lt9yd9Dk1_2),.clk(gclk));
	jdff dff_B_UuhZQnPW4_2(.din(w_dff_B_Lt9yd9Dk1_2),.dout(w_dff_B_UuhZQnPW4_2),.clk(gclk));
	jdff dff_B_bYhuYC8K5_2(.din(w_dff_B_UuhZQnPW4_2),.dout(w_dff_B_bYhuYC8K5_2),.clk(gclk));
	jdff dff_B_tCOv0GtU3_2(.din(w_dff_B_bYhuYC8K5_2),.dout(w_dff_B_tCOv0GtU3_2),.clk(gclk));
	jdff dff_B_LkK62bDd0_2(.din(w_dff_B_tCOv0GtU3_2),.dout(w_dff_B_LkK62bDd0_2),.clk(gclk));
	jdff dff_B_FdqfFCXn2_2(.din(w_dff_B_LkK62bDd0_2),.dout(w_dff_B_FdqfFCXn2_2),.clk(gclk));
	jdff dff_B_hxVovnc37_2(.din(w_dff_B_FdqfFCXn2_2),.dout(w_dff_B_hxVovnc37_2),.clk(gclk));
	jdff dff_B_tFMXEZ056_2(.din(w_dff_B_hxVovnc37_2),.dout(w_dff_B_tFMXEZ056_2),.clk(gclk));
	jdff dff_B_YG1uLtQO4_2(.din(w_dff_B_tFMXEZ056_2),.dout(w_dff_B_YG1uLtQO4_2),.clk(gclk));
	jdff dff_B_NIhudi1f7_2(.din(w_dff_B_YG1uLtQO4_2),.dout(w_dff_B_NIhudi1f7_2),.clk(gclk));
	jdff dff_B_FBxUjoSz5_2(.din(w_dff_B_NIhudi1f7_2),.dout(w_dff_B_FBxUjoSz5_2),.clk(gclk));
	jdff dff_B_c7fpcYcG8_2(.din(w_dff_B_FBxUjoSz5_2),.dout(w_dff_B_c7fpcYcG8_2),.clk(gclk));
	jdff dff_B_5NAKAHfi0_2(.din(w_dff_B_c7fpcYcG8_2),.dout(w_dff_B_5NAKAHfi0_2),.clk(gclk));
	jdff dff_B_P6j1z3zi3_2(.din(w_dff_B_5NAKAHfi0_2),.dout(w_dff_B_P6j1z3zi3_2),.clk(gclk));
	jdff dff_B_eaU1Od7X3_2(.din(w_dff_B_P6j1z3zi3_2),.dout(w_dff_B_eaU1Od7X3_2),.clk(gclk));
	jdff dff_B_luTLKIV70_2(.din(w_dff_B_eaU1Od7X3_2),.dout(w_dff_B_luTLKIV70_2),.clk(gclk));
	jdff dff_B_czYanEhE8_2(.din(w_dff_B_luTLKIV70_2),.dout(w_dff_B_czYanEhE8_2),.clk(gclk));
	jdff dff_B_X6ighRgX3_2(.din(w_dff_B_czYanEhE8_2),.dout(w_dff_B_X6ighRgX3_2),.clk(gclk));
	jdff dff_B_asnk09Ta4_2(.din(w_dff_B_X6ighRgX3_2),.dout(w_dff_B_asnk09Ta4_2),.clk(gclk));
	jdff dff_B_ijlB5QAU4_2(.din(w_dff_B_asnk09Ta4_2),.dout(w_dff_B_ijlB5QAU4_2),.clk(gclk));
	jdff dff_B_hmkodBnU9_2(.din(w_dff_B_ijlB5QAU4_2),.dout(w_dff_B_hmkodBnU9_2),.clk(gclk));
	jdff dff_B_9m5MlGyv0_2(.din(w_dff_B_hmkodBnU9_2),.dout(w_dff_B_9m5MlGyv0_2),.clk(gclk));
	jdff dff_B_oEHLFViE1_2(.din(w_dff_B_9m5MlGyv0_2),.dout(w_dff_B_oEHLFViE1_2),.clk(gclk));
	jdff dff_B_7IopQFbk8_2(.din(w_dff_B_oEHLFViE1_2),.dout(w_dff_B_7IopQFbk8_2),.clk(gclk));
	jdff dff_B_FJXngTPx4_2(.din(w_dff_B_7IopQFbk8_2),.dout(w_dff_B_FJXngTPx4_2),.clk(gclk));
	jdff dff_B_CcvmYj4K1_2(.din(w_dff_B_FJXngTPx4_2),.dout(w_dff_B_CcvmYj4K1_2),.clk(gclk));
	jdff dff_B_IcljosVj9_2(.din(w_dff_B_CcvmYj4K1_2),.dout(w_dff_B_IcljosVj9_2),.clk(gclk));
	jdff dff_B_D3OS0tOl8_2(.din(w_dff_B_IcljosVj9_2),.dout(w_dff_B_D3OS0tOl8_2),.clk(gclk));
	jdff dff_B_vLq7xXXe6_2(.din(w_dff_B_D3OS0tOl8_2),.dout(w_dff_B_vLq7xXXe6_2),.clk(gclk));
	jdff dff_B_Cxlbn2YH1_2(.din(w_dff_B_vLq7xXXe6_2),.dout(w_dff_B_Cxlbn2YH1_2),.clk(gclk));
	jdff dff_B_bYDkw8ey7_2(.din(w_dff_B_Cxlbn2YH1_2),.dout(w_dff_B_bYDkw8ey7_2),.clk(gclk));
	jdff dff_B_YsVtuTww3_2(.din(w_dff_B_bYDkw8ey7_2),.dout(w_dff_B_YsVtuTww3_2),.clk(gclk));
	jdff dff_B_zeQHvMfS1_2(.din(w_dff_B_YsVtuTww3_2),.dout(w_dff_B_zeQHvMfS1_2),.clk(gclk));
	jdff dff_B_xh3h0ZTH5_2(.din(w_dff_B_zeQHvMfS1_2),.dout(w_dff_B_xh3h0ZTH5_2),.clk(gclk));
	jdff dff_B_Bxbj5GNR9_2(.din(w_dff_B_xh3h0ZTH5_2),.dout(w_dff_B_Bxbj5GNR9_2),.clk(gclk));
	jdff dff_B_DDQoObtD0_2(.din(w_dff_B_Bxbj5GNR9_2),.dout(w_dff_B_DDQoObtD0_2),.clk(gclk));
	jdff dff_B_WPWPEX9p4_2(.din(w_dff_B_DDQoObtD0_2),.dout(w_dff_B_WPWPEX9p4_2),.clk(gclk));
	jdff dff_B_qe5l42G07_2(.din(w_dff_B_WPWPEX9p4_2),.dout(w_dff_B_qe5l42G07_2),.clk(gclk));
	jdff dff_B_5NwC0zyT1_2(.din(w_dff_B_qe5l42G07_2),.dout(w_dff_B_5NwC0zyT1_2),.clk(gclk));
	jdff dff_B_XMJKtRfu1_2(.din(w_dff_B_5NwC0zyT1_2),.dout(w_dff_B_XMJKtRfu1_2),.clk(gclk));
	jdff dff_B_gPYNN6We1_2(.din(w_dff_B_XMJKtRfu1_2),.dout(w_dff_B_gPYNN6We1_2),.clk(gclk));
	jdff dff_B_4X61qpGa9_2(.din(w_dff_B_gPYNN6We1_2),.dout(w_dff_B_4X61qpGa9_2),.clk(gclk));
	jdff dff_B_g88UkIkL3_2(.din(w_dff_B_4X61qpGa9_2),.dout(w_dff_B_g88UkIkL3_2),.clk(gclk));
	jdff dff_B_xm3ajwH93_2(.din(w_dff_B_g88UkIkL3_2),.dout(w_dff_B_xm3ajwH93_2),.clk(gclk));
	jdff dff_B_LgYseWrf1_2(.din(w_dff_B_xm3ajwH93_2),.dout(w_dff_B_LgYseWrf1_2),.clk(gclk));
	jdff dff_B_fwwxPM7b0_2(.din(w_dff_B_LgYseWrf1_2),.dout(w_dff_B_fwwxPM7b0_2),.clk(gclk));
	jdff dff_B_oawvuwEe3_2(.din(w_dff_B_fwwxPM7b0_2),.dout(w_dff_B_oawvuwEe3_2),.clk(gclk));
	jdff dff_B_smj7f7QK1_2(.din(w_dff_B_oawvuwEe3_2),.dout(w_dff_B_smj7f7QK1_2),.clk(gclk));
	jdff dff_B_eAyBbxsi5_2(.din(w_dff_B_smj7f7QK1_2),.dout(w_dff_B_eAyBbxsi5_2),.clk(gclk));
	jdff dff_B_qwcLaNmX5_2(.din(n1806),.dout(w_dff_B_qwcLaNmX5_2),.clk(gclk));
	jdff dff_B_DCVTibQ27_1(.din(n1804),.dout(w_dff_B_DCVTibQ27_1),.clk(gclk));
	jdff dff_B_mBr9zinK6_2(.din(n1775),.dout(w_dff_B_mBr9zinK6_2),.clk(gclk));
	jdff dff_B_LULJaJzn4_2(.din(w_dff_B_mBr9zinK6_2),.dout(w_dff_B_LULJaJzn4_2),.clk(gclk));
	jdff dff_B_sUAEr5C76_2(.din(w_dff_B_LULJaJzn4_2),.dout(w_dff_B_sUAEr5C76_2),.clk(gclk));
	jdff dff_B_7O0dQzBl7_2(.din(w_dff_B_sUAEr5C76_2),.dout(w_dff_B_7O0dQzBl7_2),.clk(gclk));
	jdff dff_B_2bRqSR7K4_2(.din(w_dff_B_7O0dQzBl7_2),.dout(w_dff_B_2bRqSR7K4_2),.clk(gclk));
	jdff dff_B_9oiuXmBM5_2(.din(w_dff_B_2bRqSR7K4_2),.dout(w_dff_B_9oiuXmBM5_2),.clk(gclk));
	jdff dff_B_CWyPJmsp1_2(.din(w_dff_B_9oiuXmBM5_2),.dout(w_dff_B_CWyPJmsp1_2),.clk(gclk));
	jdff dff_B_JQClPjCb6_2(.din(w_dff_B_CWyPJmsp1_2),.dout(w_dff_B_JQClPjCb6_2),.clk(gclk));
	jdff dff_B_vmLGuPmO0_2(.din(w_dff_B_JQClPjCb6_2),.dout(w_dff_B_vmLGuPmO0_2),.clk(gclk));
	jdff dff_B_M3aP8gb95_2(.din(w_dff_B_vmLGuPmO0_2),.dout(w_dff_B_M3aP8gb95_2),.clk(gclk));
	jdff dff_B_wV5zPB190_2(.din(w_dff_B_M3aP8gb95_2),.dout(w_dff_B_wV5zPB190_2),.clk(gclk));
	jdff dff_B_sjcZzzYF5_2(.din(w_dff_B_wV5zPB190_2),.dout(w_dff_B_sjcZzzYF5_2),.clk(gclk));
	jdff dff_B_430T1Hu07_2(.din(w_dff_B_sjcZzzYF5_2),.dout(w_dff_B_430T1Hu07_2),.clk(gclk));
	jdff dff_B_W97Gox2J2_2(.din(w_dff_B_430T1Hu07_2),.dout(w_dff_B_W97Gox2J2_2),.clk(gclk));
	jdff dff_B_y0f3K5dY3_2(.din(w_dff_B_W97Gox2J2_2),.dout(w_dff_B_y0f3K5dY3_2),.clk(gclk));
	jdff dff_B_6msuEzT60_2(.din(w_dff_B_y0f3K5dY3_2),.dout(w_dff_B_6msuEzT60_2),.clk(gclk));
	jdff dff_B_b4ApuG0W5_2(.din(w_dff_B_6msuEzT60_2),.dout(w_dff_B_b4ApuG0W5_2),.clk(gclk));
	jdff dff_B_f0i7id6f0_2(.din(w_dff_B_b4ApuG0W5_2),.dout(w_dff_B_f0i7id6f0_2),.clk(gclk));
	jdff dff_B_fy0ZoZUL7_2(.din(w_dff_B_f0i7id6f0_2),.dout(w_dff_B_fy0ZoZUL7_2),.clk(gclk));
	jdff dff_B_DjY4juBD1_2(.din(w_dff_B_fy0ZoZUL7_2),.dout(w_dff_B_DjY4juBD1_2),.clk(gclk));
	jdff dff_B_NP1GV6ld1_2(.din(w_dff_B_DjY4juBD1_2),.dout(w_dff_B_NP1GV6ld1_2),.clk(gclk));
	jdff dff_B_paD3DpxO7_2(.din(w_dff_B_NP1GV6ld1_2),.dout(w_dff_B_paD3DpxO7_2),.clk(gclk));
	jdff dff_B_sDHHtcpz7_2(.din(w_dff_B_paD3DpxO7_2),.dout(w_dff_B_sDHHtcpz7_2),.clk(gclk));
	jdff dff_B_wjppf0Bc1_2(.din(w_dff_B_sDHHtcpz7_2),.dout(w_dff_B_wjppf0Bc1_2),.clk(gclk));
	jdff dff_B_lbLrs8LF4_2(.din(w_dff_B_wjppf0Bc1_2),.dout(w_dff_B_lbLrs8LF4_2),.clk(gclk));
	jdff dff_B_L0DmwOYo7_2(.din(w_dff_B_lbLrs8LF4_2),.dout(w_dff_B_L0DmwOYo7_2),.clk(gclk));
	jdff dff_B_Ft5TVyL50_2(.din(w_dff_B_L0DmwOYo7_2),.dout(w_dff_B_Ft5TVyL50_2),.clk(gclk));
	jdff dff_B_9aue72Ua0_2(.din(w_dff_B_Ft5TVyL50_2),.dout(w_dff_B_9aue72Ua0_2),.clk(gclk));
	jdff dff_B_cIwxU3zM3_2(.din(w_dff_B_9aue72Ua0_2),.dout(w_dff_B_cIwxU3zM3_2),.clk(gclk));
	jdff dff_B_RHqIKApR7_2(.din(w_dff_B_cIwxU3zM3_2),.dout(w_dff_B_RHqIKApR7_2),.clk(gclk));
	jdff dff_B_ujN89r0g6_2(.din(w_dff_B_RHqIKApR7_2),.dout(w_dff_B_ujN89r0g6_2),.clk(gclk));
	jdff dff_B_wvxQYmri1_2(.din(w_dff_B_ujN89r0g6_2),.dout(w_dff_B_wvxQYmri1_2),.clk(gclk));
	jdff dff_B_ePiEQjG64_2(.din(w_dff_B_wvxQYmri1_2),.dout(w_dff_B_ePiEQjG64_2),.clk(gclk));
	jdff dff_B_GrU9M4Jm8_2(.din(w_dff_B_ePiEQjG64_2),.dout(w_dff_B_GrU9M4Jm8_2),.clk(gclk));
	jdff dff_B_6f4JRWgK8_2(.din(w_dff_B_GrU9M4Jm8_2),.dout(w_dff_B_6f4JRWgK8_2),.clk(gclk));
	jdff dff_B_D5mwCWO32_2(.din(w_dff_B_6f4JRWgK8_2),.dout(w_dff_B_D5mwCWO32_2),.clk(gclk));
	jdff dff_B_xl4p3TSt5_2(.din(w_dff_B_D5mwCWO32_2),.dout(w_dff_B_xl4p3TSt5_2),.clk(gclk));
	jdff dff_B_9GkEsjpZ8_2(.din(w_dff_B_xl4p3TSt5_2),.dout(w_dff_B_9GkEsjpZ8_2),.clk(gclk));
	jdff dff_B_lAUcFlBh4_2(.din(w_dff_B_9GkEsjpZ8_2),.dout(w_dff_B_lAUcFlBh4_2),.clk(gclk));
	jdff dff_B_DOaNXmBB7_2(.din(w_dff_B_lAUcFlBh4_2),.dout(w_dff_B_DOaNXmBB7_2),.clk(gclk));
	jdff dff_B_2MlMu2sh8_2(.din(w_dff_B_DOaNXmBB7_2),.dout(w_dff_B_2MlMu2sh8_2),.clk(gclk));
	jdff dff_B_74oQAdo70_2(.din(w_dff_B_2MlMu2sh8_2),.dout(w_dff_B_74oQAdo70_2),.clk(gclk));
	jdff dff_B_3wHcWuwi0_2(.din(w_dff_B_74oQAdo70_2),.dout(w_dff_B_3wHcWuwi0_2),.clk(gclk));
	jdff dff_B_R67BSxLW1_2(.din(w_dff_B_3wHcWuwi0_2),.dout(w_dff_B_R67BSxLW1_2),.clk(gclk));
	jdff dff_B_Vw8N4D9R7_2(.din(w_dff_B_R67BSxLW1_2),.dout(w_dff_B_Vw8N4D9R7_2),.clk(gclk));
	jdff dff_B_00ZDp0qO0_2(.din(w_dff_B_Vw8N4D9R7_2),.dout(w_dff_B_00ZDp0qO0_2),.clk(gclk));
	jdff dff_B_52nWTJBW9_2(.din(w_dff_B_00ZDp0qO0_2),.dout(w_dff_B_52nWTJBW9_2),.clk(gclk));
	jdff dff_B_gh6p9pkQ1_2(.din(w_dff_B_52nWTJBW9_2),.dout(w_dff_B_gh6p9pkQ1_2),.clk(gclk));
	jdff dff_B_ov1qn2jK9_2(.din(w_dff_B_gh6p9pkQ1_2),.dout(w_dff_B_ov1qn2jK9_2),.clk(gclk));
	jdff dff_B_gKuxhXwY3_2(.din(w_dff_B_ov1qn2jK9_2),.dout(w_dff_B_gKuxhXwY3_2),.clk(gclk));
	jdff dff_B_KRSHZt2L9_2(.din(w_dff_B_gKuxhXwY3_2),.dout(w_dff_B_KRSHZt2L9_2),.clk(gclk));
	jdff dff_B_1pa574RV7_1(.din(n1781),.dout(w_dff_B_1pa574RV7_1),.clk(gclk));
	jdff dff_B_ab685Q2h6_1(.din(w_dff_B_1pa574RV7_1),.dout(w_dff_B_ab685Q2h6_1),.clk(gclk));
	jdff dff_B_ZTQGXS6I4_2(.din(n1780),.dout(w_dff_B_ZTQGXS6I4_2),.clk(gclk));
	jdff dff_B_Lx3mjdSi3_2(.din(w_dff_B_ZTQGXS6I4_2),.dout(w_dff_B_Lx3mjdSi3_2),.clk(gclk));
	jdff dff_B_2yMd3pmf8_2(.din(w_dff_B_Lx3mjdSi3_2),.dout(w_dff_B_2yMd3pmf8_2),.clk(gclk));
	jdff dff_B_GvLXw1Dy4_2(.din(w_dff_B_2yMd3pmf8_2),.dout(w_dff_B_GvLXw1Dy4_2),.clk(gclk));
	jdff dff_B_Y34VWZRz1_2(.din(w_dff_B_GvLXw1Dy4_2),.dout(w_dff_B_Y34VWZRz1_2),.clk(gclk));
	jdff dff_B_ASvUhJ8E6_2(.din(w_dff_B_Y34VWZRz1_2),.dout(w_dff_B_ASvUhJ8E6_2),.clk(gclk));
	jdff dff_B_0DR97vdd7_2(.din(w_dff_B_ASvUhJ8E6_2),.dout(w_dff_B_0DR97vdd7_2),.clk(gclk));
	jdff dff_B_mhEG4gnA9_2(.din(w_dff_B_0DR97vdd7_2),.dout(w_dff_B_mhEG4gnA9_2),.clk(gclk));
	jdff dff_B_NiVKBVR14_2(.din(w_dff_B_mhEG4gnA9_2),.dout(w_dff_B_NiVKBVR14_2),.clk(gclk));
	jdff dff_B_zg14c5Ki7_2(.din(w_dff_B_NiVKBVR14_2),.dout(w_dff_B_zg14c5Ki7_2),.clk(gclk));
	jdff dff_B_KW35wHnr4_2(.din(w_dff_B_zg14c5Ki7_2),.dout(w_dff_B_KW35wHnr4_2),.clk(gclk));
	jdff dff_B_Lr2extkt9_2(.din(w_dff_B_KW35wHnr4_2),.dout(w_dff_B_Lr2extkt9_2),.clk(gclk));
	jdff dff_B_dTuSMScV1_2(.din(w_dff_B_Lr2extkt9_2),.dout(w_dff_B_dTuSMScV1_2),.clk(gclk));
	jdff dff_B_HUyS1SZJ5_2(.din(w_dff_B_dTuSMScV1_2),.dout(w_dff_B_HUyS1SZJ5_2),.clk(gclk));
	jdff dff_B_wi4EoFSo0_2(.din(w_dff_B_HUyS1SZJ5_2),.dout(w_dff_B_wi4EoFSo0_2),.clk(gclk));
	jdff dff_B_JBWjeKvm9_2(.din(w_dff_B_wi4EoFSo0_2),.dout(w_dff_B_JBWjeKvm9_2),.clk(gclk));
	jdff dff_B_nPHj5vVo7_2(.din(w_dff_B_JBWjeKvm9_2),.dout(w_dff_B_nPHj5vVo7_2),.clk(gclk));
	jdff dff_B_zboqbU9m7_2(.din(w_dff_B_nPHj5vVo7_2),.dout(w_dff_B_zboqbU9m7_2),.clk(gclk));
	jdff dff_B_Dpr5pW0F1_2(.din(w_dff_B_zboqbU9m7_2),.dout(w_dff_B_Dpr5pW0F1_2),.clk(gclk));
	jdff dff_B_4Rt9FTG91_2(.din(w_dff_B_Dpr5pW0F1_2),.dout(w_dff_B_4Rt9FTG91_2),.clk(gclk));
	jdff dff_B_poSUiAYG0_2(.din(w_dff_B_4Rt9FTG91_2),.dout(w_dff_B_poSUiAYG0_2),.clk(gclk));
	jdff dff_B_kIyNPvVA4_2(.din(w_dff_B_poSUiAYG0_2),.dout(w_dff_B_kIyNPvVA4_2),.clk(gclk));
	jdff dff_B_jTSwfXPJ8_2(.din(w_dff_B_kIyNPvVA4_2),.dout(w_dff_B_jTSwfXPJ8_2),.clk(gclk));
	jdff dff_B_nOxYfUo26_2(.din(w_dff_B_jTSwfXPJ8_2),.dout(w_dff_B_nOxYfUo26_2),.clk(gclk));
	jdff dff_B_h8cPlX6y5_2(.din(w_dff_B_nOxYfUo26_2),.dout(w_dff_B_h8cPlX6y5_2),.clk(gclk));
	jdff dff_B_WPqMUme29_2(.din(w_dff_B_h8cPlX6y5_2),.dout(w_dff_B_WPqMUme29_2),.clk(gclk));
	jdff dff_B_MI5UAQtl8_2(.din(w_dff_B_WPqMUme29_2),.dout(w_dff_B_MI5UAQtl8_2),.clk(gclk));
	jdff dff_B_WRtTMCzU1_2(.din(w_dff_B_MI5UAQtl8_2),.dout(w_dff_B_WRtTMCzU1_2),.clk(gclk));
	jdff dff_B_5n4V0OA64_2(.din(w_dff_B_WRtTMCzU1_2),.dout(w_dff_B_5n4V0OA64_2),.clk(gclk));
	jdff dff_B_O4WLllGz5_2(.din(w_dff_B_5n4V0OA64_2),.dout(w_dff_B_O4WLllGz5_2),.clk(gclk));
	jdff dff_B_qP2Freca0_2(.din(w_dff_B_O4WLllGz5_2),.dout(w_dff_B_qP2Freca0_2),.clk(gclk));
	jdff dff_B_aYAGfY9R4_2(.din(w_dff_B_qP2Freca0_2),.dout(w_dff_B_aYAGfY9R4_2),.clk(gclk));
	jdff dff_B_HQbZyGRz8_2(.din(w_dff_B_aYAGfY9R4_2),.dout(w_dff_B_HQbZyGRz8_2),.clk(gclk));
	jdff dff_B_6XQUihbW8_2(.din(w_dff_B_HQbZyGRz8_2),.dout(w_dff_B_6XQUihbW8_2),.clk(gclk));
	jdff dff_B_Hn32oo9u0_2(.din(w_dff_B_6XQUihbW8_2),.dout(w_dff_B_Hn32oo9u0_2),.clk(gclk));
	jdff dff_B_aYmWKJlS1_2(.din(w_dff_B_Hn32oo9u0_2),.dout(w_dff_B_aYmWKJlS1_2),.clk(gclk));
	jdff dff_B_RddqjjSj7_2(.din(w_dff_B_aYmWKJlS1_2),.dout(w_dff_B_RddqjjSj7_2),.clk(gclk));
	jdff dff_B_KzTHHdTZ9_2(.din(w_dff_B_RddqjjSj7_2),.dout(w_dff_B_KzTHHdTZ9_2),.clk(gclk));
	jdff dff_B_LQMIU07m6_2(.din(w_dff_B_KzTHHdTZ9_2),.dout(w_dff_B_LQMIU07m6_2),.clk(gclk));
	jdff dff_B_ANxyz6Kb5_2(.din(w_dff_B_LQMIU07m6_2),.dout(w_dff_B_ANxyz6Kb5_2),.clk(gclk));
	jdff dff_B_NCvwvwDQ1_2(.din(w_dff_B_ANxyz6Kb5_2),.dout(w_dff_B_NCvwvwDQ1_2),.clk(gclk));
	jdff dff_B_8ZyEKesh8_2(.din(w_dff_B_NCvwvwDQ1_2),.dout(w_dff_B_8ZyEKesh8_2),.clk(gclk));
	jdff dff_B_12TJV3oR1_2(.din(w_dff_B_8ZyEKesh8_2),.dout(w_dff_B_12TJV3oR1_2),.clk(gclk));
	jdff dff_B_6pviUdXw0_2(.din(w_dff_B_12TJV3oR1_2),.dout(w_dff_B_6pviUdXw0_2),.clk(gclk));
	jdff dff_B_Lgp6UKpm6_2(.din(w_dff_B_6pviUdXw0_2),.dout(w_dff_B_Lgp6UKpm6_2),.clk(gclk));
	jdff dff_B_vPpUmE0L7_2(.din(w_dff_B_Lgp6UKpm6_2),.dout(w_dff_B_vPpUmE0L7_2),.clk(gclk));
	jdff dff_B_JTOL4DZN6_2(.din(w_dff_B_vPpUmE0L7_2),.dout(w_dff_B_JTOL4DZN6_2),.clk(gclk));
	jdff dff_B_T0DnmlcE6_2(.din(w_dff_B_JTOL4DZN6_2),.dout(w_dff_B_T0DnmlcE6_2),.clk(gclk));
	jdff dff_B_UTRszQtn2_2(.din(n1779),.dout(w_dff_B_UTRszQtn2_2),.clk(gclk));
	jdff dff_B_Cr8357xq0_2(.din(w_dff_B_UTRszQtn2_2),.dout(w_dff_B_Cr8357xq0_2),.clk(gclk));
	jdff dff_B_QZf6fSZk6_2(.din(w_dff_B_Cr8357xq0_2),.dout(w_dff_B_QZf6fSZk6_2),.clk(gclk));
	jdff dff_B_KPhStNhc8_2(.din(w_dff_B_QZf6fSZk6_2),.dout(w_dff_B_KPhStNhc8_2),.clk(gclk));
	jdff dff_B_vWPu9wjV8_2(.din(w_dff_B_KPhStNhc8_2),.dout(w_dff_B_vWPu9wjV8_2),.clk(gclk));
	jdff dff_B_YYYBmQsF7_2(.din(w_dff_B_vWPu9wjV8_2),.dout(w_dff_B_YYYBmQsF7_2),.clk(gclk));
	jdff dff_B_ePWIeJ7V6_2(.din(w_dff_B_YYYBmQsF7_2),.dout(w_dff_B_ePWIeJ7V6_2),.clk(gclk));
	jdff dff_B_bzgpolVd7_2(.din(w_dff_B_ePWIeJ7V6_2),.dout(w_dff_B_bzgpolVd7_2),.clk(gclk));
	jdff dff_B_JbbDq3Bd9_2(.din(w_dff_B_bzgpolVd7_2),.dout(w_dff_B_JbbDq3Bd9_2),.clk(gclk));
	jdff dff_B_05NofmFR7_2(.din(w_dff_B_JbbDq3Bd9_2),.dout(w_dff_B_05NofmFR7_2),.clk(gclk));
	jdff dff_B_grb6c2iX6_2(.din(w_dff_B_05NofmFR7_2),.dout(w_dff_B_grb6c2iX6_2),.clk(gclk));
	jdff dff_B_3T42BwSA4_2(.din(w_dff_B_grb6c2iX6_2),.dout(w_dff_B_3T42BwSA4_2),.clk(gclk));
	jdff dff_B_6MX5TUvy2_2(.din(w_dff_B_3T42BwSA4_2),.dout(w_dff_B_6MX5TUvy2_2),.clk(gclk));
	jdff dff_B_vhJlguC05_2(.din(w_dff_B_6MX5TUvy2_2),.dout(w_dff_B_vhJlguC05_2),.clk(gclk));
	jdff dff_B_e7b6DkQD1_2(.din(w_dff_B_vhJlguC05_2),.dout(w_dff_B_e7b6DkQD1_2),.clk(gclk));
	jdff dff_B_Jlhw6XOj4_2(.din(w_dff_B_e7b6DkQD1_2),.dout(w_dff_B_Jlhw6XOj4_2),.clk(gclk));
	jdff dff_B_BztSFJGT6_2(.din(w_dff_B_Jlhw6XOj4_2),.dout(w_dff_B_BztSFJGT6_2),.clk(gclk));
	jdff dff_B_WCvndrbo4_2(.din(w_dff_B_BztSFJGT6_2),.dout(w_dff_B_WCvndrbo4_2),.clk(gclk));
	jdff dff_B_O0eLY8gG7_2(.din(w_dff_B_WCvndrbo4_2),.dout(w_dff_B_O0eLY8gG7_2),.clk(gclk));
	jdff dff_B_XRz4o72X2_2(.din(w_dff_B_O0eLY8gG7_2),.dout(w_dff_B_XRz4o72X2_2),.clk(gclk));
	jdff dff_B_gdE9GhUH5_2(.din(w_dff_B_XRz4o72X2_2),.dout(w_dff_B_gdE9GhUH5_2),.clk(gclk));
	jdff dff_B_owaIawDw8_2(.din(w_dff_B_gdE9GhUH5_2),.dout(w_dff_B_owaIawDw8_2),.clk(gclk));
	jdff dff_B_4DSfg6gF5_2(.din(w_dff_B_owaIawDw8_2),.dout(w_dff_B_4DSfg6gF5_2),.clk(gclk));
	jdff dff_B_2NbcAh0T1_2(.din(w_dff_B_4DSfg6gF5_2),.dout(w_dff_B_2NbcAh0T1_2),.clk(gclk));
	jdff dff_B_gdSaeRLj7_2(.din(w_dff_B_2NbcAh0T1_2),.dout(w_dff_B_gdSaeRLj7_2),.clk(gclk));
	jdff dff_B_9HrCLUZ11_2(.din(w_dff_B_gdSaeRLj7_2),.dout(w_dff_B_9HrCLUZ11_2),.clk(gclk));
	jdff dff_B_pm2HzBRZ3_2(.din(w_dff_B_9HrCLUZ11_2),.dout(w_dff_B_pm2HzBRZ3_2),.clk(gclk));
	jdff dff_B_bGsG0aH45_2(.din(w_dff_B_pm2HzBRZ3_2),.dout(w_dff_B_bGsG0aH45_2),.clk(gclk));
	jdff dff_B_4EO0Me7n0_2(.din(w_dff_B_bGsG0aH45_2),.dout(w_dff_B_4EO0Me7n0_2),.clk(gclk));
	jdff dff_B_xAwSMO3D1_2(.din(w_dff_B_4EO0Me7n0_2),.dout(w_dff_B_xAwSMO3D1_2),.clk(gclk));
	jdff dff_B_z2EjJ4dY6_2(.din(w_dff_B_xAwSMO3D1_2),.dout(w_dff_B_z2EjJ4dY6_2),.clk(gclk));
	jdff dff_B_WsrsDtnA7_2(.din(w_dff_B_z2EjJ4dY6_2),.dout(w_dff_B_WsrsDtnA7_2),.clk(gclk));
	jdff dff_B_Njbn7fqq4_2(.din(w_dff_B_WsrsDtnA7_2),.dout(w_dff_B_Njbn7fqq4_2),.clk(gclk));
	jdff dff_B_5El2Biyu2_2(.din(w_dff_B_Njbn7fqq4_2),.dout(w_dff_B_5El2Biyu2_2),.clk(gclk));
	jdff dff_B_bYCIXVhK1_2(.din(w_dff_B_5El2Biyu2_2),.dout(w_dff_B_bYCIXVhK1_2),.clk(gclk));
	jdff dff_B_Yq0xn5UJ7_2(.din(w_dff_B_bYCIXVhK1_2),.dout(w_dff_B_Yq0xn5UJ7_2),.clk(gclk));
	jdff dff_B_Sxnc3k794_2(.din(w_dff_B_Yq0xn5UJ7_2),.dout(w_dff_B_Sxnc3k794_2),.clk(gclk));
	jdff dff_B_WM4jHbNO0_2(.din(w_dff_B_Sxnc3k794_2),.dout(w_dff_B_WM4jHbNO0_2),.clk(gclk));
	jdff dff_B_8k2UQPcp3_2(.din(w_dff_B_WM4jHbNO0_2),.dout(w_dff_B_8k2UQPcp3_2),.clk(gclk));
	jdff dff_B_CQGVIHtp5_2(.din(w_dff_B_8k2UQPcp3_2),.dout(w_dff_B_CQGVIHtp5_2),.clk(gclk));
	jdff dff_B_WqHq0ZFJ8_2(.din(w_dff_B_CQGVIHtp5_2),.dout(w_dff_B_WqHq0ZFJ8_2),.clk(gclk));
	jdff dff_B_awSFrf515_2(.din(w_dff_B_WqHq0ZFJ8_2),.dout(w_dff_B_awSFrf515_2),.clk(gclk));
	jdff dff_B_rlXqutju2_2(.din(w_dff_B_awSFrf515_2),.dout(w_dff_B_rlXqutju2_2),.clk(gclk));
	jdff dff_B_inKx7PGA4_2(.din(w_dff_B_rlXqutju2_2),.dout(w_dff_B_inKx7PGA4_2),.clk(gclk));
	jdff dff_B_RWuu1e251_2(.din(w_dff_B_inKx7PGA4_2),.dout(w_dff_B_RWuu1e251_2),.clk(gclk));
	jdff dff_B_5rGmhKVO8_2(.din(w_dff_B_RWuu1e251_2),.dout(w_dff_B_5rGmhKVO8_2),.clk(gclk));
	jdff dff_B_dzzTHMoz6_2(.din(w_dff_B_5rGmhKVO8_2),.dout(w_dff_B_dzzTHMoz6_2),.clk(gclk));
	jdff dff_B_eIn0hFC26_2(.din(w_dff_B_dzzTHMoz6_2),.dout(w_dff_B_eIn0hFC26_2),.clk(gclk));
	jdff dff_B_DigdRgnJ2_2(.din(w_dff_B_eIn0hFC26_2),.dout(w_dff_B_DigdRgnJ2_2),.clk(gclk));
	jdff dff_B_qFmd4odf4_2(.din(w_dff_B_DigdRgnJ2_2),.dout(w_dff_B_qFmd4odf4_2),.clk(gclk));
	jdff dff_B_agF8t62T8_2(.din(n1778),.dout(w_dff_B_agF8t62T8_2),.clk(gclk));
	jdff dff_B_3hVnrSk46_1(.din(n1776),.dout(w_dff_B_3hVnrSk46_1),.clk(gclk));
	jdff dff_B_5T2MMC6t4_2(.din(n1740),.dout(w_dff_B_5T2MMC6t4_2),.clk(gclk));
	jdff dff_B_jHJYw1tZ2_2(.din(w_dff_B_5T2MMC6t4_2),.dout(w_dff_B_jHJYw1tZ2_2),.clk(gclk));
	jdff dff_B_ipwt0XsT6_2(.din(w_dff_B_jHJYw1tZ2_2),.dout(w_dff_B_ipwt0XsT6_2),.clk(gclk));
	jdff dff_B_1eZUEalB9_2(.din(w_dff_B_ipwt0XsT6_2),.dout(w_dff_B_1eZUEalB9_2),.clk(gclk));
	jdff dff_B_ZLREOlSh2_2(.din(w_dff_B_1eZUEalB9_2),.dout(w_dff_B_ZLREOlSh2_2),.clk(gclk));
	jdff dff_B_3WHtvTS26_2(.din(w_dff_B_ZLREOlSh2_2),.dout(w_dff_B_3WHtvTS26_2),.clk(gclk));
	jdff dff_B_r3UPrdIk0_2(.din(w_dff_B_3WHtvTS26_2),.dout(w_dff_B_r3UPrdIk0_2),.clk(gclk));
	jdff dff_B_30ZujImX2_2(.din(w_dff_B_r3UPrdIk0_2),.dout(w_dff_B_30ZujImX2_2),.clk(gclk));
	jdff dff_B_LuAgpGXj1_2(.din(w_dff_B_30ZujImX2_2),.dout(w_dff_B_LuAgpGXj1_2),.clk(gclk));
	jdff dff_B_CueCAGRS1_2(.din(w_dff_B_LuAgpGXj1_2),.dout(w_dff_B_CueCAGRS1_2),.clk(gclk));
	jdff dff_B_rR8nMODP8_2(.din(w_dff_B_CueCAGRS1_2),.dout(w_dff_B_rR8nMODP8_2),.clk(gclk));
	jdff dff_B_vlA4WHrT9_2(.din(w_dff_B_rR8nMODP8_2),.dout(w_dff_B_vlA4WHrT9_2),.clk(gclk));
	jdff dff_B_hNPXYkr54_2(.din(w_dff_B_vlA4WHrT9_2),.dout(w_dff_B_hNPXYkr54_2),.clk(gclk));
	jdff dff_B_CbJP7g9z3_2(.din(w_dff_B_hNPXYkr54_2),.dout(w_dff_B_CbJP7g9z3_2),.clk(gclk));
	jdff dff_B_l7GiGpvr5_2(.din(w_dff_B_CbJP7g9z3_2),.dout(w_dff_B_l7GiGpvr5_2),.clk(gclk));
	jdff dff_B_TlmxsKRL8_2(.din(w_dff_B_l7GiGpvr5_2),.dout(w_dff_B_TlmxsKRL8_2),.clk(gclk));
	jdff dff_B_9TkOdnhg8_2(.din(w_dff_B_TlmxsKRL8_2),.dout(w_dff_B_9TkOdnhg8_2),.clk(gclk));
	jdff dff_B_o0H4G08Y3_2(.din(w_dff_B_9TkOdnhg8_2),.dout(w_dff_B_o0H4G08Y3_2),.clk(gclk));
	jdff dff_B_XlcvIfD08_2(.din(w_dff_B_o0H4G08Y3_2),.dout(w_dff_B_XlcvIfD08_2),.clk(gclk));
	jdff dff_B_Rmq9Dlrt6_2(.din(w_dff_B_XlcvIfD08_2),.dout(w_dff_B_Rmq9Dlrt6_2),.clk(gclk));
	jdff dff_B_fu5VFzlx7_2(.din(w_dff_B_Rmq9Dlrt6_2),.dout(w_dff_B_fu5VFzlx7_2),.clk(gclk));
	jdff dff_B_wIA6K3Ev7_2(.din(w_dff_B_fu5VFzlx7_2),.dout(w_dff_B_wIA6K3Ev7_2),.clk(gclk));
	jdff dff_B_ub2kmoWX3_2(.din(w_dff_B_wIA6K3Ev7_2),.dout(w_dff_B_ub2kmoWX3_2),.clk(gclk));
	jdff dff_B_U2zk2YV07_2(.din(w_dff_B_ub2kmoWX3_2),.dout(w_dff_B_U2zk2YV07_2),.clk(gclk));
	jdff dff_B_aYTXs1Rt6_2(.din(w_dff_B_U2zk2YV07_2),.dout(w_dff_B_aYTXs1Rt6_2),.clk(gclk));
	jdff dff_B_4RGwT7B56_2(.din(w_dff_B_aYTXs1Rt6_2),.dout(w_dff_B_4RGwT7B56_2),.clk(gclk));
	jdff dff_B_opA2uA8u9_2(.din(w_dff_B_4RGwT7B56_2),.dout(w_dff_B_opA2uA8u9_2),.clk(gclk));
	jdff dff_B_znimIONV6_2(.din(w_dff_B_opA2uA8u9_2),.dout(w_dff_B_znimIONV6_2),.clk(gclk));
	jdff dff_B_0Is8eCHY6_2(.din(w_dff_B_znimIONV6_2),.dout(w_dff_B_0Is8eCHY6_2),.clk(gclk));
	jdff dff_B_tqvDZqSD6_2(.din(w_dff_B_0Is8eCHY6_2),.dout(w_dff_B_tqvDZqSD6_2),.clk(gclk));
	jdff dff_B_fO3nrgpd7_2(.din(w_dff_B_tqvDZqSD6_2),.dout(w_dff_B_fO3nrgpd7_2),.clk(gclk));
	jdff dff_B_bVnvuLRV5_2(.din(w_dff_B_fO3nrgpd7_2),.dout(w_dff_B_bVnvuLRV5_2),.clk(gclk));
	jdff dff_B_peI1zMN58_2(.din(w_dff_B_bVnvuLRV5_2),.dout(w_dff_B_peI1zMN58_2),.clk(gclk));
	jdff dff_B_uVS5ZH7X4_2(.din(w_dff_B_peI1zMN58_2),.dout(w_dff_B_uVS5ZH7X4_2),.clk(gclk));
	jdff dff_B_m8kkNvOa9_2(.din(w_dff_B_uVS5ZH7X4_2),.dout(w_dff_B_m8kkNvOa9_2),.clk(gclk));
	jdff dff_B_zMTkOWJj4_2(.din(w_dff_B_m8kkNvOa9_2),.dout(w_dff_B_zMTkOWJj4_2),.clk(gclk));
	jdff dff_B_4VO5xxc52_2(.din(w_dff_B_zMTkOWJj4_2),.dout(w_dff_B_4VO5xxc52_2),.clk(gclk));
	jdff dff_B_rsDZjJQp9_2(.din(w_dff_B_4VO5xxc52_2),.dout(w_dff_B_rsDZjJQp9_2),.clk(gclk));
	jdff dff_B_Xx1zgopg7_2(.din(w_dff_B_rsDZjJQp9_2),.dout(w_dff_B_Xx1zgopg7_2),.clk(gclk));
	jdff dff_B_UJiMHZ1T7_2(.din(w_dff_B_Xx1zgopg7_2),.dout(w_dff_B_UJiMHZ1T7_2),.clk(gclk));
	jdff dff_B_CqfMuxuq4_2(.din(w_dff_B_UJiMHZ1T7_2),.dout(w_dff_B_CqfMuxuq4_2),.clk(gclk));
	jdff dff_B_fQriyvUs6_2(.din(w_dff_B_CqfMuxuq4_2),.dout(w_dff_B_fQriyvUs6_2),.clk(gclk));
	jdff dff_B_rbfuiNGA4_2(.din(w_dff_B_fQriyvUs6_2),.dout(w_dff_B_rbfuiNGA4_2),.clk(gclk));
	jdff dff_B_0L2gbH7y8_2(.din(w_dff_B_rbfuiNGA4_2),.dout(w_dff_B_0L2gbH7y8_2),.clk(gclk));
	jdff dff_B_IQenXnjK5_2(.din(w_dff_B_0L2gbH7y8_2),.dout(w_dff_B_IQenXnjK5_2),.clk(gclk));
	jdff dff_B_gVBE3rh19_2(.din(w_dff_B_IQenXnjK5_2),.dout(w_dff_B_gVBE3rh19_2),.clk(gclk));
	jdff dff_B_DyB1IKPC5_2(.din(w_dff_B_gVBE3rh19_2),.dout(w_dff_B_DyB1IKPC5_2),.clk(gclk));
	jdff dff_B_qT5sAETC5_1(.din(n1746),.dout(w_dff_B_qT5sAETC5_1),.clk(gclk));
	jdff dff_B_ITq5ODvv5_1(.din(w_dff_B_qT5sAETC5_1),.dout(w_dff_B_ITq5ODvv5_1),.clk(gclk));
	jdff dff_B_sqPDmQhi6_2(.din(n1745),.dout(w_dff_B_sqPDmQhi6_2),.clk(gclk));
	jdff dff_B_XHC47qVA8_2(.din(w_dff_B_sqPDmQhi6_2),.dout(w_dff_B_XHC47qVA8_2),.clk(gclk));
	jdff dff_B_Lcsrw7ZW2_2(.din(w_dff_B_XHC47qVA8_2),.dout(w_dff_B_Lcsrw7ZW2_2),.clk(gclk));
	jdff dff_B_AghjpGzh2_2(.din(w_dff_B_Lcsrw7ZW2_2),.dout(w_dff_B_AghjpGzh2_2),.clk(gclk));
	jdff dff_B_AsT0YJje5_2(.din(w_dff_B_AghjpGzh2_2),.dout(w_dff_B_AsT0YJje5_2),.clk(gclk));
	jdff dff_B_jMrePLeH8_2(.din(w_dff_B_AsT0YJje5_2),.dout(w_dff_B_jMrePLeH8_2),.clk(gclk));
	jdff dff_B_Ra7XznvX7_2(.din(w_dff_B_jMrePLeH8_2),.dout(w_dff_B_Ra7XznvX7_2),.clk(gclk));
	jdff dff_B_sPrRGCIl5_2(.din(w_dff_B_Ra7XznvX7_2),.dout(w_dff_B_sPrRGCIl5_2),.clk(gclk));
	jdff dff_B_9m5DIBku3_2(.din(w_dff_B_sPrRGCIl5_2),.dout(w_dff_B_9m5DIBku3_2),.clk(gclk));
	jdff dff_B_wd47nu722_2(.din(w_dff_B_9m5DIBku3_2),.dout(w_dff_B_wd47nu722_2),.clk(gclk));
	jdff dff_B_kOheLc7A8_2(.din(w_dff_B_wd47nu722_2),.dout(w_dff_B_kOheLc7A8_2),.clk(gclk));
	jdff dff_B_UBxZJgp13_2(.din(w_dff_B_kOheLc7A8_2),.dout(w_dff_B_UBxZJgp13_2),.clk(gclk));
	jdff dff_B_W3z5arOG0_2(.din(w_dff_B_UBxZJgp13_2),.dout(w_dff_B_W3z5arOG0_2),.clk(gclk));
	jdff dff_B_nEPJvcAE5_2(.din(w_dff_B_W3z5arOG0_2),.dout(w_dff_B_nEPJvcAE5_2),.clk(gclk));
	jdff dff_B_e9AZpvSL1_2(.din(w_dff_B_nEPJvcAE5_2),.dout(w_dff_B_e9AZpvSL1_2),.clk(gclk));
	jdff dff_B_34hCClRC5_2(.din(w_dff_B_e9AZpvSL1_2),.dout(w_dff_B_34hCClRC5_2),.clk(gclk));
	jdff dff_B_QtxlQDeo3_2(.din(w_dff_B_34hCClRC5_2),.dout(w_dff_B_QtxlQDeo3_2),.clk(gclk));
	jdff dff_B_A5G1GQsU1_2(.din(w_dff_B_QtxlQDeo3_2),.dout(w_dff_B_A5G1GQsU1_2),.clk(gclk));
	jdff dff_B_Z6WgYcih9_2(.din(w_dff_B_A5G1GQsU1_2),.dout(w_dff_B_Z6WgYcih9_2),.clk(gclk));
	jdff dff_B_Un0gvM0A3_2(.din(w_dff_B_Z6WgYcih9_2),.dout(w_dff_B_Un0gvM0A3_2),.clk(gclk));
	jdff dff_B_cEG43IBd2_2(.din(w_dff_B_Un0gvM0A3_2),.dout(w_dff_B_cEG43IBd2_2),.clk(gclk));
	jdff dff_B_UmiKB51T9_2(.din(w_dff_B_cEG43IBd2_2),.dout(w_dff_B_UmiKB51T9_2),.clk(gclk));
	jdff dff_B_vmejwXTn7_2(.din(w_dff_B_UmiKB51T9_2),.dout(w_dff_B_vmejwXTn7_2),.clk(gclk));
	jdff dff_B_fBUGWA7r4_2(.din(w_dff_B_vmejwXTn7_2),.dout(w_dff_B_fBUGWA7r4_2),.clk(gclk));
	jdff dff_B_RybLmypm7_2(.din(w_dff_B_fBUGWA7r4_2),.dout(w_dff_B_RybLmypm7_2),.clk(gclk));
	jdff dff_B_TrRCfxIc6_2(.din(w_dff_B_RybLmypm7_2),.dout(w_dff_B_TrRCfxIc6_2),.clk(gclk));
	jdff dff_B_NudGuLI28_2(.din(w_dff_B_TrRCfxIc6_2),.dout(w_dff_B_NudGuLI28_2),.clk(gclk));
	jdff dff_B_Udft1zug1_2(.din(w_dff_B_NudGuLI28_2),.dout(w_dff_B_Udft1zug1_2),.clk(gclk));
	jdff dff_B_bndFKDjV2_2(.din(w_dff_B_Udft1zug1_2),.dout(w_dff_B_bndFKDjV2_2),.clk(gclk));
	jdff dff_B_tRLHHMq32_2(.din(w_dff_B_bndFKDjV2_2),.dout(w_dff_B_tRLHHMq32_2),.clk(gclk));
	jdff dff_B_6oO5qoZ88_2(.din(w_dff_B_tRLHHMq32_2),.dout(w_dff_B_6oO5qoZ88_2),.clk(gclk));
	jdff dff_B_PPkq81yt1_2(.din(w_dff_B_6oO5qoZ88_2),.dout(w_dff_B_PPkq81yt1_2),.clk(gclk));
	jdff dff_B_Up27UF968_2(.din(w_dff_B_PPkq81yt1_2),.dout(w_dff_B_Up27UF968_2),.clk(gclk));
	jdff dff_B_h8i0gn0l5_2(.din(w_dff_B_Up27UF968_2),.dout(w_dff_B_h8i0gn0l5_2),.clk(gclk));
	jdff dff_B_pa97XfOY7_2(.din(w_dff_B_h8i0gn0l5_2),.dout(w_dff_B_pa97XfOY7_2),.clk(gclk));
	jdff dff_B_9G0AjUt00_2(.din(w_dff_B_pa97XfOY7_2),.dout(w_dff_B_9G0AjUt00_2),.clk(gclk));
	jdff dff_B_hDkgm3b39_2(.din(w_dff_B_9G0AjUt00_2),.dout(w_dff_B_hDkgm3b39_2),.clk(gclk));
	jdff dff_B_gRhSfi7Y4_2(.din(w_dff_B_hDkgm3b39_2),.dout(w_dff_B_gRhSfi7Y4_2),.clk(gclk));
	jdff dff_B_kFbdzq0O6_2(.din(w_dff_B_gRhSfi7Y4_2),.dout(w_dff_B_kFbdzq0O6_2),.clk(gclk));
	jdff dff_B_Vk0OT2gT7_2(.din(w_dff_B_kFbdzq0O6_2),.dout(w_dff_B_Vk0OT2gT7_2),.clk(gclk));
	jdff dff_B_0NfvmgbE2_2(.din(w_dff_B_Vk0OT2gT7_2),.dout(w_dff_B_0NfvmgbE2_2),.clk(gclk));
	jdff dff_B_IQFjwthz5_2(.din(w_dff_B_0NfvmgbE2_2),.dout(w_dff_B_IQFjwthz5_2),.clk(gclk));
	jdff dff_B_MgjlpJUQ4_2(.din(w_dff_B_IQFjwthz5_2),.dout(w_dff_B_MgjlpJUQ4_2),.clk(gclk));
	jdff dff_B_XccXmWny7_2(.din(w_dff_B_MgjlpJUQ4_2),.dout(w_dff_B_XccXmWny7_2),.clk(gclk));
	jdff dff_B_bIda4Wl94_2(.din(n1744),.dout(w_dff_B_bIda4Wl94_2),.clk(gclk));
	jdff dff_B_D2cKQdCD6_2(.din(w_dff_B_bIda4Wl94_2),.dout(w_dff_B_D2cKQdCD6_2),.clk(gclk));
	jdff dff_B_WOviowce3_2(.din(w_dff_B_D2cKQdCD6_2),.dout(w_dff_B_WOviowce3_2),.clk(gclk));
	jdff dff_B_RtvW9lIH1_2(.din(w_dff_B_WOviowce3_2),.dout(w_dff_B_RtvW9lIH1_2),.clk(gclk));
	jdff dff_B_ngoc9Dr45_2(.din(w_dff_B_RtvW9lIH1_2),.dout(w_dff_B_ngoc9Dr45_2),.clk(gclk));
	jdff dff_B_yM6Mq15k2_2(.din(w_dff_B_ngoc9Dr45_2),.dout(w_dff_B_yM6Mq15k2_2),.clk(gclk));
	jdff dff_B_YYC0TVfN6_2(.din(w_dff_B_yM6Mq15k2_2),.dout(w_dff_B_YYC0TVfN6_2),.clk(gclk));
	jdff dff_B_LcvQ6Vel9_2(.din(w_dff_B_YYC0TVfN6_2),.dout(w_dff_B_LcvQ6Vel9_2),.clk(gclk));
	jdff dff_B_Gj7zbwEj5_2(.din(w_dff_B_LcvQ6Vel9_2),.dout(w_dff_B_Gj7zbwEj5_2),.clk(gclk));
	jdff dff_B_NIhRWEWa3_2(.din(w_dff_B_Gj7zbwEj5_2),.dout(w_dff_B_NIhRWEWa3_2),.clk(gclk));
	jdff dff_B_6RhbpRHq5_2(.din(w_dff_B_NIhRWEWa3_2),.dout(w_dff_B_6RhbpRHq5_2),.clk(gclk));
	jdff dff_B_xrjWXvYI5_2(.din(w_dff_B_6RhbpRHq5_2),.dout(w_dff_B_xrjWXvYI5_2),.clk(gclk));
	jdff dff_B_nOwczB7i9_2(.din(w_dff_B_xrjWXvYI5_2),.dout(w_dff_B_nOwczB7i9_2),.clk(gclk));
	jdff dff_B_sw9dZln41_2(.din(w_dff_B_nOwczB7i9_2),.dout(w_dff_B_sw9dZln41_2),.clk(gclk));
	jdff dff_B_zBpaf05x4_2(.din(w_dff_B_sw9dZln41_2),.dout(w_dff_B_zBpaf05x4_2),.clk(gclk));
	jdff dff_B_HPBngvMO2_2(.din(w_dff_B_zBpaf05x4_2),.dout(w_dff_B_HPBngvMO2_2),.clk(gclk));
	jdff dff_B_V2xOTHGb5_2(.din(w_dff_B_HPBngvMO2_2),.dout(w_dff_B_V2xOTHGb5_2),.clk(gclk));
	jdff dff_B_M9SZ4K9n7_2(.din(w_dff_B_V2xOTHGb5_2),.dout(w_dff_B_M9SZ4K9n7_2),.clk(gclk));
	jdff dff_B_BVMznqHk9_2(.din(w_dff_B_M9SZ4K9n7_2),.dout(w_dff_B_BVMznqHk9_2),.clk(gclk));
	jdff dff_B_c1B8b2oY8_2(.din(w_dff_B_BVMznqHk9_2),.dout(w_dff_B_c1B8b2oY8_2),.clk(gclk));
	jdff dff_B_idg30Hq10_2(.din(w_dff_B_c1B8b2oY8_2),.dout(w_dff_B_idg30Hq10_2),.clk(gclk));
	jdff dff_B_2RjKTG4C6_2(.din(w_dff_B_idg30Hq10_2),.dout(w_dff_B_2RjKTG4C6_2),.clk(gclk));
	jdff dff_B_ro5LUE5u7_2(.din(w_dff_B_2RjKTG4C6_2),.dout(w_dff_B_ro5LUE5u7_2),.clk(gclk));
	jdff dff_B_COgsj6Jh5_2(.din(w_dff_B_ro5LUE5u7_2),.dout(w_dff_B_COgsj6Jh5_2),.clk(gclk));
	jdff dff_B_IyAuwlPp5_2(.din(w_dff_B_COgsj6Jh5_2),.dout(w_dff_B_IyAuwlPp5_2),.clk(gclk));
	jdff dff_B_Iz5CJ1uM3_2(.din(w_dff_B_IyAuwlPp5_2),.dout(w_dff_B_Iz5CJ1uM3_2),.clk(gclk));
	jdff dff_B_HlG3ISFt2_2(.din(w_dff_B_Iz5CJ1uM3_2),.dout(w_dff_B_HlG3ISFt2_2),.clk(gclk));
	jdff dff_B_Rd4TqUI25_2(.din(w_dff_B_HlG3ISFt2_2),.dout(w_dff_B_Rd4TqUI25_2),.clk(gclk));
	jdff dff_B_cDI7qBXs5_2(.din(w_dff_B_Rd4TqUI25_2),.dout(w_dff_B_cDI7qBXs5_2),.clk(gclk));
	jdff dff_B_EqfTcMKK7_2(.din(w_dff_B_cDI7qBXs5_2),.dout(w_dff_B_EqfTcMKK7_2),.clk(gclk));
	jdff dff_B_dCEUnK2t6_2(.din(w_dff_B_EqfTcMKK7_2),.dout(w_dff_B_dCEUnK2t6_2),.clk(gclk));
	jdff dff_B_8Lpohban6_2(.din(w_dff_B_dCEUnK2t6_2),.dout(w_dff_B_8Lpohban6_2),.clk(gclk));
	jdff dff_B_3mIoPgG90_2(.din(w_dff_B_8Lpohban6_2),.dout(w_dff_B_3mIoPgG90_2),.clk(gclk));
	jdff dff_B_0gNR8ukV1_2(.din(w_dff_B_3mIoPgG90_2),.dout(w_dff_B_0gNR8ukV1_2),.clk(gclk));
	jdff dff_B_ZOUbpQuz2_2(.din(w_dff_B_0gNR8ukV1_2),.dout(w_dff_B_ZOUbpQuz2_2),.clk(gclk));
	jdff dff_B_zi9iEQlJ1_2(.din(w_dff_B_ZOUbpQuz2_2),.dout(w_dff_B_zi9iEQlJ1_2),.clk(gclk));
	jdff dff_B_P4LaNWa51_2(.din(w_dff_B_zi9iEQlJ1_2),.dout(w_dff_B_P4LaNWa51_2),.clk(gclk));
	jdff dff_B_KWCFnulf0_2(.din(w_dff_B_P4LaNWa51_2),.dout(w_dff_B_KWCFnulf0_2),.clk(gclk));
	jdff dff_B_FqOHMpem9_2(.din(w_dff_B_KWCFnulf0_2),.dout(w_dff_B_FqOHMpem9_2),.clk(gclk));
	jdff dff_B_2Xg4DstL1_2(.din(w_dff_B_FqOHMpem9_2),.dout(w_dff_B_2Xg4DstL1_2),.clk(gclk));
	jdff dff_B_1B3fioXq4_2(.din(w_dff_B_2Xg4DstL1_2),.dout(w_dff_B_1B3fioXq4_2),.clk(gclk));
	jdff dff_B_SlOPBWUG4_2(.din(w_dff_B_1B3fioXq4_2),.dout(w_dff_B_SlOPBWUG4_2),.clk(gclk));
	jdff dff_B_ZlrO80Xt4_2(.din(w_dff_B_SlOPBWUG4_2),.dout(w_dff_B_ZlrO80Xt4_2),.clk(gclk));
	jdff dff_B_o2rqvsZX4_2(.din(w_dff_B_ZlrO80Xt4_2),.dout(w_dff_B_o2rqvsZX4_2),.clk(gclk));
	jdff dff_B_DAygf4x11_2(.din(w_dff_B_o2rqvsZX4_2),.dout(w_dff_B_DAygf4x11_2),.clk(gclk));
	jdff dff_B_B7RNIbNT7_2(.din(w_dff_B_DAygf4x11_2),.dout(w_dff_B_B7RNIbNT7_2),.clk(gclk));
	jdff dff_B_0wdXCfdC9_2(.din(n1743),.dout(w_dff_B_0wdXCfdC9_2),.clk(gclk));
	jdff dff_B_UFVwRiwo2_1(.din(n1741),.dout(w_dff_B_UFVwRiwo2_1),.clk(gclk));
	jdff dff_B_4CbQx41F9_2(.din(n1699),.dout(w_dff_B_4CbQx41F9_2),.clk(gclk));
	jdff dff_B_tOzd0Gtu8_2(.din(w_dff_B_4CbQx41F9_2),.dout(w_dff_B_tOzd0Gtu8_2),.clk(gclk));
	jdff dff_B_3RK9jRb23_2(.din(w_dff_B_tOzd0Gtu8_2),.dout(w_dff_B_3RK9jRb23_2),.clk(gclk));
	jdff dff_B_aHLVSmPo4_2(.din(w_dff_B_3RK9jRb23_2),.dout(w_dff_B_aHLVSmPo4_2),.clk(gclk));
	jdff dff_B_njx5V7RV3_2(.din(w_dff_B_aHLVSmPo4_2),.dout(w_dff_B_njx5V7RV3_2),.clk(gclk));
	jdff dff_B_AWLuKZf47_2(.din(w_dff_B_njx5V7RV3_2),.dout(w_dff_B_AWLuKZf47_2),.clk(gclk));
	jdff dff_B_8yo0YQbD7_2(.din(w_dff_B_AWLuKZf47_2),.dout(w_dff_B_8yo0YQbD7_2),.clk(gclk));
	jdff dff_B_R1JKiXfl3_2(.din(w_dff_B_8yo0YQbD7_2),.dout(w_dff_B_R1JKiXfl3_2),.clk(gclk));
	jdff dff_B_hPiNVPYx9_2(.din(w_dff_B_R1JKiXfl3_2),.dout(w_dff_B_hPiNVPYx9_2),.clk(gclk));
	jdff dff_B_xRtlWB7b4_2(.din(w_dff_B_hPiNVPYx9_2),.dout(w_dff_B_xRtlWB7b4_2),.clk(gclk));
	jdff dff_B_7g4ARltO2_2(.din(w_dff_B_xRtlWB7b4_2),.dout(w_dff_B_7g4ARltO2_2),.clk(gclk));
	jdff dff_B_cl3vqZW91_2(.din(w_dff_B_7g4ARltO2_2),.dout(w_dff_B_cl3vqZW91_2),.clk(gclk));
	jdff dff_B_aifoDLxY3_2(.din(w_dff_B_cl3vqZW91_2),.dout(w_dff_B_aifoDLxY3_2),.clk(gclk));
	jdff dff_B_WZ7VcjL10_2(.din(w_dff_B_aifoDLxY3_2),.dout(w_dff_B_WZ7VcjL10_2),.clk(gclk));
	jdff dff_B_6HbPTyBX3_2(.din(w_dff_B_WZ7VcjL10_2),.dout(w_dff_B_6HbPTyBX3_2),.clk(gclk));
	jdff dff_B_UlcXload6_2(.din(w_dff_B_6HbPTyBX3_2),.dout(w_dff_B_UlcXload6_2),.clk(gclk));
	jdff dff_B_DWbaprGE6_2(.din(w_dff_B_UlcXload6_2),.dout(w_dff_B_DWbaprGE6_2),.clk(gclk));
	jdff dff_B_0v5qJSuu3_2(.din(w_dff_B_DWbaprGE6_2),.dout(w_dff_B_0v5qJSuu3_2),.clk(gclk));
	jdff dff_B_rt0SGGiy8_2(.din(w_dff_B_0v5qJSuu3_2),.dout(w_dff_B_rt0SGGiy8_2),.clk(gclk));
	jdff dff_B_uYwP1HhH2_2(.din(w_dff_B_rt0SGGiy8_2),.dout(w_dff_B_uYwP1HhH2_2),.clk(gclk));
	jdff dff_B_8Gn5FTjb7_2(.din(w_dff_B_uYwP1HhH2_2),.dout(w_dff_B_8Gn5FTjb7_2),.clk(gclk));
	jdff dff_B_thXTg66f1_2(.din(w_dff_B_8Gn5FTjb7_2),.dout(w_dff_B_thXTg66f1_2),.clk(gclk));
	jdff dff_B_1C367qgX9_2(.din(w_dff_B_thXTg66f1_2),.dout(w_dff_B_1C367qgX9_2),.clk(gclk));
	jdff dff_B_d8ORhABr8_2(.din(w_dff_B_1C367qgX9_2),.dout(w_dff_B_d8ORhABr8_2),.clk(gclk));
	jdff dff_B_5ixPI9vT5_2(.din(w_dff_B_d8ORhABr8_2),.dout(w_dff_B_5ixPI9vT5_2),.clk(gclk));
	jdff dff_B_s2XpSyNf3_2(.din(w_dff_B_5ixPI9vT5_2),.dout(w_dff_B_s2XpSyNf3_2),.clk(gclk));
	jdff dff_B_FPkc7MQy5_2(.din(w_dff_B_s2XpSyNf3_2),.dout(w_dff_B_FPkc7MQy5_2),.clk(gclk));
	jdff dff_B_Lfo6DpxF6_2(.din(w_dff_B_FPkc7MQy5_2),.dout(w_dff_B_Lfo6DpxF6_2),.clk(gclk));
	jdff dff_B_dgD72bWa6_2(.din(w_dff_B_Lfo6DpxF6_2),.dout(w_dff_B_dgD72bWa6_2),.clk(gclk));
	jdff dff_B_BY1kU5Ct4_2(.din(w_dff_B_dgD72bWa6_2),.dout(w_dff_B_BY1kU5Ct4_2),.clk(gclk));
	jdff dff_B_eFP3B0QO9_2(.din(w_dff_B_BY1kU5Ct4_2),.dout(w_dff_B_eFP3B0QO9_2),.clk(gclk));
	jdff dff_B_HJR4GMn03_2(.din(w_dff_B_eFP3B0QO9_2),.dout(w_dff_B_HJR4GMn03_2),.clk(gclk));
	jdff dff_B_pV2aBFeC8_2(.din(w_dff_B_HJR4GMn03_2),.dout(w_dff_B_pV2aBFeC8_2),.clk(gclk));
	jdff dff_B_UM4RUzm44_2(.din(w_dff_B_pV2aBFeC8_2),.dout(w_dff_B_UM4RUzm44_2),.clk(gclk));
	jdff dff_B_zr5HyVi01_2(.din(w_dff_B_UM4RUzm44_2),.dout(w_dff_B_zr5HyVi01_2),.clk(gclk));
	jdff dff_B_z2ACCUCN5_2(.din(w_dff_B_zr5HyVi01_2),.dout(w_dff_B_z2ACCUCN5_2),.clk(gclk));
	jdff dff_B_szGS4o266_2(.din(w_dff_B_z2ACCUCN5_2),.dout(w_dff_B_szGS4o266_2),.clk(gclk));
	jdff dff_B_gLEu3eWy3_2(.din(w_dff_B_szGS4o266_2),.dout(w_dff_B_gLEu3eWy3_2),.clk(gclk));
	jdff dff_B_BMMSSA753_2(.din(w_dff_B_gLEu3eWy3_2),.dout(w_dff_B_BMMSSA753_2),.clk(gclk));
	jdff dff_B_BBLcp6S29_2(.din(w_dff_B_BMMSSA753_2),.dout(w_dff_B_BBLcp6S29_2),.clk(gclk));
	jdff dff_B_9MIUmrvb4_2(.din(w_dff_B_BBLcp6S29_2),.dout(w_dff_B_9MIUmrvb4_2),.clk(gclk));
	jdff dff_B_WvOsFQZ35_2(.din(w_dff_B_9MIUmrvb4_2),.dout(w_dff_B_WvOsFQZ35_2),.clk(gclk));
	jdff dff_B_YpBZ67h04_2(.din(w_dff_B_WvOsFQZ35_2),.dout(w_dff_B_YpBZ67h04_2),.clk(gclk));
	jdff dff_B_YXZvJO2k0_1(.din(n1705),.dout(w_dff_B_YXZvJO2k0_1),.clk(gclk));
	jdff dff_B_sl9LlNAT0_1(.din(w_dff_B_YXZvJO2k0_1),.dout(w_dff_B_sl9LlNAT0_1),.clk(gclk));
	jdff dff_B_a60FCBK10_2(.din(n1704),.dout(w_dff_B_a60FCBK10_2),.clk(gclk));
	jdff dff_B_s1t0Ne6l1_2(.din(w_dff_B_a60FCBK10_2),.dout(w_dff_B_s1t0Ne6l1_2),.clk(gclk));
	jdff dff_B_8txMS7B40_2(.din(w_dff_B_s1t0Ne6l1_2),.dout(w_dff_B_8txMS7B40_2),.clk(gclk));
	jdff dff_B_DX4hwEel0_2(.din(w_dff_B_8txMS7B40_2),.dout(w_dff_B_DX4hwEel0_2),.clk(gclk));
	jdff dff_B_UALV2Nvv2_2(.din(w_dff_B_DX4hwEel0_2),.dout(w_dff_B_UALV2Nvv2_2),.clk(gclk));
	jdff dff_B_rbZtHZzC4_2(.din(w_dff_B_UALV2Nvv2_2),.dout(w_dff_B_rbZtHZzC4_2),.clk(gclk));
	jdff dff_B_Mckbp9AA5_2(.din(w_dff_B_rbZtHZzC4_2),.dout(w_dff_B_Mckbp9AA5_2),.clk(gclk));
	jdff dff_B_LqIoFn6Q8_2(.din(w_dff_B_Mckbp9AA5_2),.dout(w_dff_B_LqIoFn6Q8_2),.clk(gclk));
	jdff dff_B_f3VAqxAh7_2(.din(w_dff_B_LqIoFn6Q8_2),.dout(w_dff_B_f3VAqxAh7_2),.clk(gclk));
	jdff dff_B_CnYgRNZE5_2(.din(w_dff_B_f3VAqxAh7_2),.dout(w_dff_B_CnYgRNZE5_2),.clk(gclk));
	jdff dff_B_pVWbBQ752_2(.din(w_dff_B_CnYgRNZE5_2),.dout(w_dff_B_pVWbBQ752_2),.clk(gclk));
	jdff dff_B_lQkJtgS43_2(.din(w_dff_B_pVWbBQ752_2),.dout(w_dff_B_lQkJtgS43_2),.clk(gclk));
	jdff dff_B_OoVrgO5r5_2(.din(w_dff_B_lQkJtgS43_2),.dout(w_dff_B_OoVrgO5r5_2),.clk(gclk));
	jdff dff_B_01azvw9k8_2(.din(w_dff_B_OoVrgO5r5_2),.dout(w_dff_B_01azvw9k8_2),.clk(gclk));
	jdff dff_B_vvHpNv2c6_2(.din(w_dff_B_01azvw9k8_2),.dout(w_dff_B_vvHpNv2c6_2),.clk(gclk));
	jdff dff_B_0Nxn7GMb3_2(.din(w_dff_B_vvHpNv2c6_2),.dout(w_dff_B_0Nxn7GMb3_2),.clk(gclk));
	jdff dff_B_oJBPUXTm8_2(.din(w_dff_B_0Nxn7GMb3_2),.dout(w_dff_B_oJBPUXTm8_2),.clk(gclk));
	jdff dff_B_jtkDR4jN2_2(.din(w_dff_B_oJBPUXTm8_2),.dout(w_dff_B_jtkDR4jN2_2),.clk(gclk));
	jdff dff_B_0QZrmuTs4_2(.din(w_dff_B_jtkDR4jN2_2),.dout(w_dff_B_0QZrmuTs4_2),.clk(gclk));
	jdff dff_B_4ONyxXPC6_2(.din(w_dff_B_0QZrmuTs4_2),.dout(w_dff_B_4ONyxXPC6_2),.clk(gclk));
	jdff dff_B_9DXOjNco4_2(.din(w_dff_B_4ONyxXPC6_2),.dout(w_dff_B_9DXOjNco4_2),.clk(gclk));
	jdff dff_B_plsApLue3_2(.din(w_dff_B_9DXOjNco4_2),.dout(w_dff_B_plsApLue3_2),.clk(gclk));
	jdff dff_B_iZ8OwxC19_2(.din(w_dff_B_plsApLue3_2),.dout(w_dff_B_iZ8OwxC19_2),.clk(gclk));
	jdff dff_B_P7ODU0VS2_2(.din(w_dff_B_iZ8OwxC19_2),.dout(w_dff_B_P7ODU0VS2_2),.clk(gclk));
	jdff dff_B_7XkJH0Kl6_2(.din(w_dff_B_P7ODU0VS2_2),.dout(w_dff_B_7XkJH0Kl6_2),.clk(gclk));
	jdff dff_B_J2CyJSVW3_2(.din(w_dff_B_7XkJH0Kl6_2),.dout(w_dff_B_J2CyJSVW3_2),.clk(gclk));
	jdff dff_B_awG32zrH7_2(.din(w_dff_B_J2CyJSVW3_2),.dout(w_dff_B_awG32zrH7_2),.clk(gclk));
	jdff dff_B_G4phLsEV1_2(.din(w_dff_B_awG32zrH7_2),.dout(w_dff_B_G4phLsEV1_2),.clk(gclk));
	jdff dff_B_1sSPCddY0_2(.din(w_dff_B_G4phLsEV1_2),.dout(w_dff_B_1sSPCddY0_2),.clk(gclk));
	jdff dff_B_1KItqeoN9_2(.din(w_dff_B_1sSPCddY0_2),.dout(w_dff_B_1KItqeoN9_2),.clk(gclk));
	jdff dff_B_bjkQGqVN7_2(.din(w_dff_B_1KItqeoN9_2),.dout(w_dff_B_bjkQGqVN7_2),.clk(gclk));
	jdff dff_B_GnKywHke3_2(.din(w_dff_B_bjkQGqVN7_2),.dout(w_dff_B_GnKywHke3_2),.clk(gclk));
	jdff dff_B_hcg06UVb7_2(.din(w_dff_B_GnKywHke3_2),.dout(w_dff_B_hcg06UVb7_2),.clk(gclk));
	jdff dff_B_KMgVGQSX8_2(.din(w_dff_B_hcg06UVb7_2),.dout(w_dff_B_KMgVGQSX8_2),.clk(gclk));
	jdff dff_B_m8TLvjHr8_2(.din(w_dff_B_KMgVGQSX8_2),.dout(w_dff_B_m8TLvjHr8_2),.clk(gclk));
	jdff dff_B_lBGh094G6_2(.din(w_dff_B_m8TLvjHr8_2),.dout(w_dff_B_lBGh094G6_2),.clk(gclk));
	jdff dff_B_A9W44fyG5_2(.din(w_dff_B_lBGh094G6_2),.dout(w_dff_B_A9W44fyG5_2),.clk(gclk));
	jdff dff_B_ITUO9W679_2(.din(w_dff_B_A9W44fyG5_2),.dout(w_dff_B_ITUO9W679_2),.clk(gclk));
	jdff dff_B_jubSsqcg2_2(.din(w_dff_B_ITUO9W679_2),.dout(w_dff_B_jubSsqcg2_2),.clk(gclk));
	jdff dff_B_ftAC1Tv30_2(.din(w_dff_B_jubSsqcg2_2),.dout(w_dff_B_ftAC1Tv30_2),.clk(gclk));
	jdff dff_B_lQcMoh2d5_2(.din(n1703),.dout(w_dff_B_lQcMoh2d5_2),.clk(gclk));
	jdff dff_B_RzhjSOY79_2(.din(w_dff_B_lQcMoh2d5_2),.dout(w_dff_B_RzhjSOY79_2),.clk(gclk));
	jdff dff_B_IVtF71gj1_2(.din(w_dff_B_RzhjSOY79_2),.dout(w_dff_B_IVtF71gj1_2),.clk(gclk));
	jdff dff_B_ne5l9KOw5_2(.din(w_dff_B_IVtF71gj1_2),.dout(w_dff_B_ne5l9KOw5_2),.clk(gclk));
	jdff dff_B_LZv7m9H48_2(.din(w_dff_B_ne5l9KOw5_2),.dout(w_dff_B_LZv7m9H48_2),.clk(gclk));
	jdff dff_B_xLPZGdPs7_2(.din(w_dff_B_LZv7m9H48_2),.dout(w_dff_B_xLPZGdPs7_2),.clk(gclk));
	jdff dff_B_WpcYmYiE8_2(.din(w_dff_B_xLPZGdPs7_2),.dout(w_dff_B_WpcYmYiE8_2),.clk(gclk));
	jdff dff_B_Xe29gkP29_2(.din(w_dff_B_WpcYmYiE8_2),.dout(w_dff_B_Xe29gkP29_2),.clk(gclk));
	jdff dff_B_X8q39fkN9_2(.din(w_dff_B_Xe29gkP29_2),.dout(w_dff_B_X8q39fkN9_2),.clk(gclk));
	jdff dff_B_qEs4RS6u6_2(.din(w_dff_B_X8q39fkN9_2),.dout(w_dff_B_qEs4RS6u6_2),.clk(gclk));
	jdff dff_B_wu1PItlE7_2(.din(w_dff_B_qEs4RS6u6_2),.dout(w_dff_B_wu1PItlE7_2),.clk(gclk));
	jdff dff_B_b7iuyeou2_2(.din(w_dff_B_wu1PItlE7_2),.dout(w_dff_B_b7iuyeou2_2),.clk(gclk));
	jdff dff_B_VMXC3PbE2_2(.din(w_dff_B_b7iuyeou2_2),.dout(w_dff_B_VMXC3PbE2_2),.clk(gclk));
	jdff dff_B_mHuU6GOr7_2(.din(w_dff_B_VMXC3PbE2_2),.dout(w_dff_B_mHuU6GOr7_2),.clk(gclk));
	jdff dff_B_7fl2GvwK8_2(.din(w_dff_B_mHuU6GOr7_2),.dout(w_dff_B_7fl2GvwK8_2),.clk(gclk));
	jdff dff_B_4YiJLsiw6_2(.din(w_dff_B_7fl2GvwK8_2),.dout(w_dff_B_4YiJLsiw6_2),.clk(gclk));
	jdff dff_B_eP5FJVGW1_2(.din(w_dff_B_4YiJLsiw6_2),.dout(w_dff_B_eP5FJVGW1_2),.clk(gclk));
	jdff dff_B_d4gPjic42_2(.din(w_dff_B_eP5FJVGW1_2),.dout(w_dff_B_d4gPjic42_2),.clk(gclk));
	jdff dff_B_JOLA9J4w9_2(.din(w_dff_B_d4gPjic42_2),.dout(w_dff_B_JOLA9J4w9_2),.clk(gclk));
	jdff dff_B_c2lYvNJ78_2(.din(w_dff_B_JOLA9J4w9_2),.dout(w_dff_B_c2lYvNJ78_2),.clk(gclk));
	jdff dff_B_hODBv9zx5_2(.din(w_dff_B_c2lYvNJ78_2),.dout(w_dff_B_hODBv9zx5_2),.clk(gclk));
	jdff dff_B_zNY6mDat2_2(.din(w_dff_B_hODBv9zx5_2),.dout(w_dff_B_zNY6mDat2_2),.clk(gclk));
	jdff dff_B_x8AeANCb1_2(.din(w_dff_B_zNY6mDat2_2),.dout(w_dff_B_x8AeANCb1_2),.clk(gclk));
	jdff dff_B_gqMnlbSj4_2(.din(w_dff_B_x8AeANCb1_2),.dout(w_dff_B_gqMnlbSj4_2),.clk(gclk));
	jdff dff_B_QR4AWM4t6_2(.din(w_dff_B_gqMnlbSj4_2),.dout(w_dff_B_QR4AWM4t6_2),.clk(gclk));
	jdff dff_B_eoTPu0120_2(.din(w_dff_B_QR4AWM4t6_2),.dout(w_dff_B_eoTPu0120_2),.clk(gclk));
	jdff dff_B_KRrr06ro0_2(.din(w_dff_B_eoTPu0120_2),.dout(w_dff_B_KRrr06ro0_2),.clk(gclk));
	jdff dff_B_yPDbsUSp2_2(.din(w_dff_B_KRrr06ro0_2),.dout(w_dff_B_yPDbsUSp2_2),.clk(gclk));
	jdff dff_B_4D4VzV5M7_2(.din(w_dff_B_yPDbsUSp2_2),.dout(w_dff_B_4D4VzV5M7_2),.clk(gclk));
	jdff dff_B_iAMWRmag3_2(.din(w_dff_B_4D4VzV5M7_2),.dout(w_dff_B_iAMWRmag3_2),.clk(gclk));
	jdff dff_B_i7GRGFgO4_2(.din(w_dff_B_iAMWRmag3_2),.dout(w_dff_B_i7GRGFgO4_2),.clk(gclk));
	jdff dff_B_QEukstIO4_2(.din(w_dff_B_i7GRGFgO4_2),.dout(w_dff_B_QEukstIO4_2),.clk(gclk));
	jdff dff_B_Q5QgZt8i7_2(.din(w_dff_B_QEukstIO4_2),.dout(w_dff_B_Q5QgZt8i7_2),.clk(gclk));
	jdff dff_B_89Bz2bgh5_2(.din(w_dff_B_Q5QgZt8i7_2),.dout(w_dff_B_89Bz2bgh5_2),.clk(gclk));
	jdff dff_B_X7fyyJgm1_2(.din(w_dff_B_89Bz2bgh5_2),.dout(w_dff_B_X7fyyJgm1_2),.clk(gclk));
	jdff dff_B_pvEecekj9_2(.din(w_dff_B_X7fyyJgm1_2),.dout(w_dff_B_pvEecekj9_2),.clk(gclk));
	jdff dff_B_epgzQZn99_2(.din(w_dff_B_pvEecekj9_2),.dout(w_dff_B_epgzQZn99_2),.clk(gclk));
	jdff dff_B_WbEVTkPs8_2(.din(w_dff_B_epgzQZn99_2),.dout(w_dff_B_WbEVTkPs8_2),.clk(gclk));
	jdff dff_B_QDa8gHla1_2(.din(w_dff_B_WbEVTkPs8_2),.dout(w_dff_B_QDa8gHla1_2),.clk(gclk));
	jdff dff_B_mEwxybiH7_2(.din(w_dff_B_QDa8gHla1_2),.dout(w_dff_B_mEwxybiH7_2),.clk(gclk));
	jdff dff_B_7lJ4oeRx8_2(.din(w_dff_B_mEwxybiH7_2),.dout(w_dff_B_7lJ4oeRx8_2),.clk(gclk));
	jdff dff_B_kv4gH2Zd2_2(.din(w_dff_B_7lJ4oeRx8_2),.dout(w_dff_B_kv4gH2Zd2_2),.clk(gclk));
	jdff dff_B_hrir7I2z8_2(.din(n1702),.dout(w_dff_B_hrir7I2z8_2),.clk(gclk));
	jdff dff_B_LD9XSOiS3_1(.din(n1700),.dout(w_dff_B_LD9XSOiS3_1),.clk(gclk));
	jdff dff_B_IO8osC6D0_2(.din(n1648),.dout(w_dff_B_IO8osC6D0_2),.clk(gclk));
	jdff dff_B_5YZ5C6Kq6_2(.din(w_dff_B_IO8osC6D0_2),.dout(w_dff_B_5YZ5C6Kq6_2),.clk(gclk));
	jdff dff_B_mt6k1Qos2_2(.din(w_dff_B_5YZ5C6Kq6_2),.dout(w_dff_B_mt6k1Qos2_2),.clk(gclk));
	jdff dff_B_jtmtyrZ36_2(.din(w_dff_B_mt6k1Qos2_2),.dout(w_dff_B_jtmtyrZ36_2),.clk(gclk));
	jdff dff_B_M5YPqomP5_2(.din(w_dff_B_jtmtyrZ36_2),.dout(w_dff_B_M5YPqomP5_2),.clk(gclk));
	jdff dff_B_HgGLTEMa7_2(.din(w_dff_B_M5YPqomP5_2),.dout(w_dff_B_HgGLTEMa7_2),.clk(gclk));
	jdff dff_B_2QcuSjtX7_2(.din(w_dff_B_HgGLTEMa7_2),.dout(w_dff_B_2QcuSjtX7_2),.clk(gclk));
	jdff dff_B_wmwHp6Js4_2(.din(w_dff_B_2QcuSjtX7_2),.dout(w_dff_B_wmwHp6Js4_2),.clk(gclk));
	jdff dff_B_zzYyRr8p3_2(.din(w_dff_B_wmwHp6Js4_2),.dout(w_dff_B_zzYyRr8p3_2),.clk(gclk));
	jdff dff_B_VO1JxMWh7_2(.din(w_dff_B_zzYyRr8p3_2),.dout(w_dff_B_VO1JxMWh7_2),.clk(gclk));
	jdff dff_B_AqsmNwUX4_2(.din(w_dff_B_VO1JxMWh7_2),.dout(w_dff_B_AqsmNwUX4_2),.clk(gclk));
	jdff dff_B_B9KIpRH98_2(.din(w_dff_B_AqsmNwUX4_2),.dout(w_dff_B_B9KIpRH98_2),.clk(gclk));
	jdff dff_B_V2zO15AL1_2(.din(w_dff_B_B9KIpRH98_2),.dout(w_dff_B_V2zO15AL1_2),.clk(gclk));
	jdff dff_B_WGas6kLb8_2(.din(w_dff_B_V2zO15AL1_2),.dout(w_dff_B_WGas6kLb8_2),.clk(gclk));
	jdff dff_B_dxtI1b3L5_2(.din(w_dff_B_WGas6kLb8_2),.dout(w_dff_B_dxtI1b3L5_2),.clk(gclk));
	jdff dff_B_BNkXoz4z2_2(.din(w_dff_B_dxtI1b3L5_2),.dout(w_dff_B_BNkXoz4z2_2),.clk(gclk));
	jdff dff_B_p6AAIeBf7_2(.din(w_dff_B_BNkXoz4z2_2),.dout(w_dff_B_p6AAIeBf7_2),.clk(gclk));
	jdff dff_B_loF9KRgF4_2(.din(w_dff_B_p6AAIeBf7_2),.dout(w_dff_B_loF9KRgF4_2),.clk(gclk));
	jdff dff_B_55OKPuuj6_2(.din(w_dff_B_loF9KRgF4_2),.dout(w_dff_B_55OKPuuj6_2),.clk(gclk));
	jdff dff_B_D5tdWEfJ1_2(.din(w_dff_B_55OKPuuj6_2),.dout(w_dff_B_D5tdWEfJ1_2),.clk(gclk));
	jdff dff_B_uT3CuPGq1_2(.din(w_dff_B_D5tdWEfJ1_2),.dout(w_dff_B_uT3CuPGq1_2),.clk(gclk));
	jdff dff_B_2YkQPLcm9_2(.din(w_dff_B_uT3CuPGq1_2),.dout(w_dff_B_2YkQPLcm9_2),.clk(gclk));
	jdff dff_B_7Ie72Y0Y4_2(.din(w_dff_B_2YkQPLcm9_2),.dout(w_dff_B_7Ie72Y0Y4_2),.clk(gclk));
	jdff dff_B_LQYwPaLL0_2(.din(w_dff_B_7Ie72Y0Y4_2),.dout(w_dff_B_LQYwPaLL0_2),.clk(gclk));
	jdff dff_B_LuE6FoXo9_2(.din(w_dff_B_LQYwPaLL0_2),.dout(w_dff_B_LuE6FoXo9_2),.clk(gclk));
	jdff dff_B_VeGAicis8_2(.din(w_dff_B_LuE6FoXo9_2),.dout(w_dff_B_VeGAicis8_2),.clk(gclk));
	jdff dff_B_OAZR1hcB0_2(.din(w_dff_B_VeGAicis8_2),.dout(w_dff_B_OAZR1hcB0_2),.clk(gclk));
	jdff dff_B_z6tL5lTR1_2(.din(w_dff_B_OAZR1hcB0_2),.dout(w_dff_B_z6tL5lTR1_2),.clk(gclk));
	jdff dff_B_3SOP35U57_2(.din(w_dff_B_z6tL5lTR1_2),.dout(w_dff_B_3SOP35U57_2),.clk(gclk));
	jdff dff_B_4ldaTvvg9_2(.din(w_dff_B_3SOP35U57_2),.dout(w_dff_B_4ldaTvvg9_2),.clk(gclk));
	jdff dff_B_E4V7pNm14_2(.din(w_dff_B_4ldaTvvg9_2),.dout(w_dff_B_E4V7pNm14_2),.clk(gclk));
	jdff dff_B_GjkRbhM33_2(.din(w_dff_B_E4V7pNm14_2),.dout(w_dff_B_GjkRbhM33_2),.clk(gclk));
	jdff dff_B_8RUqxONn7_2(.din(w_dff_B_GjkRbhM33_2),.dout(w_dff_B_8RUqxONn7_2),.clk(gclk));
	jdff dff_B_rjemjsH95_2(.din(w_dff_B_8RUqxONn7_2),.dout(w_dff_B_rjemjsH95_2),.clk(gclk));
	jdff dff_B_pXfP7u089_2(.din(w_dff_B_rjemjsH95_2),.dout(w_dff_B_pXfP7u089_2),.clk(gclk));
	jdff dff_B_6fugebGy4_2(.din(w_dff_B_pXfP7u089_2),.dout(w_dff_B_6fugebGy4_2),.clk(gclk));
	jdff dff_B_SuRv9RT48_2(.din(w_dff_B_6fugebGy4_2),.dout(w_dff_B_SuRv9RT48_2),.clk(gclk));
	jdff dff_B_grxZZwjR0_2(.din(w_dff_B_SuRv9RT48_2),.dout(w_dff_B_grxZZwjR0_2),.clk(gclk));
	jdff dff_B_FH7jW32D5_2(.din(w_dff_B_grxZZwjR0_2),.dout(w_dff_B_FH7jW32D5_2),.clk(gclk));
	jdff dff_B_11h2mnBb6_1(.din(n1654),.dout(w_dff_B_11h2mnBb6_1),.clk(gclk));
	jdff dff_B_QnrhvDJ39_1(.din(w_dff_B_11h2mnBb6_1),.dout(w_dff_B_QnrhvDJ39_1),.clk(gclk));
	jdff dff_B_OjtRWkz85_2(.din(n1653),.dout(w_dff_B_OjtRWkz85_2),.clk(gclk));
	jdff dff_B_H4sLWXAM1_2(.din(w_dff_B_OjtRWkz85_2),.dout(w_dff_B_H4sLWXAM1_2),.clk(gclk));
	jdff dff_B_rhKgKYmg2_2(.din(w_dff_B_H4sLWXAM1_2),.dout(w_dff_B_rhKgKYmg2_2),.clk(gclk));
	jdff dff_B_PrcewLJg3_2(.din(w_dff_B_rhKgKYmg2_2),.dout(w_dff_B_PrcewLJg3_2),.clk(gclk));
	jdff dff_B_ciMQANda1_2(.din(w_dff_B_PrcewLJg3_2),.dout(w_dff_B_ciMQANda1_2),.clk(gclk));
	jdff dff_B_BsoIaXf27_2(.din(w_dff_B_ciMQANda1_2),.dout(w_dff_B_BsoIaXf27_2),.clk(gclk));
	jdff dff_B_oQWgyVv40_2(.din(w_dff_B_BsoIaXf27_2),.dout(w_dff_B_oQWgyVv40_2),.clk(gclk));
	jdff dff_B_yB01E5nB4_2(.din(w_dff_B_oQWgyVv40_2),.dout(w_dff_B_yB01E5nB4_2),.clk(gclk));
	jdff dff_B_7FeFVmGh3_2(.din(w_dff_B_yB01E5nB4_2),.dout(w_dff_B_7FeFVmGh3_2),.clk(gclk));
	jdff dff_B_Tmxh3YeH3_2(.din(w_dff_B_7FeFVmGh3_2),.dout(w_dff_B_Tmxh3YeH3_2),.clk(gclk));
	jdff dff_B_yCsTGjWz8_2(.din(w_dff_B_Tmxh3YeH3_2),.dout(w_dff_B_yCsTGjWz8_2),.clk(gclk));
	jdff dff_B_y9zwp4Az5_2(.din(w_dff_B_yCsTGjWz8_2),.dout(w_dff_B_y9zwp4Az5_2),.clk(gclk));
	jdff dff_B_YFiH6sbf2_2(.din(w_dff_B_y9zwp4Az5_2),.dout(w_dff_B_YFiH6sbf2_2),.clk(gclk));
	jdff dff_B_FnzaljUV9_2(.din(w_dff_B_YFiH6sbf2_2),.dout(w_dff_B_FnzaljUV9_2),.clk(gclk));
	jdff dff_B_ix1L4zjC8_2(.din(w_dff_B_FnzaljUV9_2),.dout(w_dff_B_ix1L4zjC8_2),.clk(gclk));
	jdff dff_B_VVQpPhB32_2(.din(w_dff_B_ix1L4zjC8_2),.dout(w_dff_B_VVQpPhB32_2),.clk(gclk));
	jdff dff_B_sSgwnOrU2_2(.din(w_dff_B_VVQpPhB32_2),.dout(w_dff_B_sSgwnOrU2_2),.clk(gclk));
	jdff dff_B_UJZ3Wht43_2(.din(w_dff_B_sSgwnOrU2_2),.dout(w_dff_B_UJZ3Wht43_2),.clk(gclk));
	jdff dff_B_S6OOM1Kq2_2(.din(w_dff_B_UJZ3Wht43_2),.dout(w_dff_B_S6OOM1Kq2_2),.clk(gclk));
	jdff dff_B_dBV8XEuL1_2(.din(w_dff_B_S6OOM1Kq2_2),.dout(w_dff_B_dBV8XEuL1_2),.clk(gclk));
	jdff dff_B_sxWOfH029_2(.din(w_dff_B_dBV8XEuL1_2),.dout(w_dff_B_sxWOfH029_2),.clk(gclk));
	jdff dff_B_uwtfZuaL3_2(.din(w_dff_B_sxWOfH029_2),.dout(w_dff_B_uwtfZuaL3_2),.clk(gclk));
	jdff dff_B_PRHyGlfj1_2(.din(w_dff_B_uwtfZuaL3_2),.dout(w_dff_B_PRHyGlfj1_2),.clk(gclk));
	jdff dff_B_NwBrKywE1_2(.din(w_dff_B_PRHyGlfj1_2),.dout(w_dff_B_NwBrKywE1_2),.clk(gclk));
	jdff dff_B_mI0wTFno9_2(.din(w_dff_B_NwBrKywE1_2),.dout(w_dff_B_mI0wTFno9_2),.clk(gclk));
	jdff dff_B_hX6AAV445_2(.din(w_dff_B_mI0wTFno9_2),.dout(w_dff_B_hX6AAV445_2),.clk(gclk));
	jdff dff_B_5CvxOZxv5_2(.din(w_dff_B_hX6AAV445_2),.dout(w_dff_B_5CvxOZxv5_2),.clk(gclk));
	jdff dff_B_7c00OjEb2_2(.din(w_dff_B_5CvxOZxv5_2),.dout(w_dff_B_7c00OjEb2_2),.clk(gclk));
	jdff dff_B_MbRKR5KN5_2(.din(w_dff_B_7c00OjEb2_2),.dout(w_dff_B_MbRKR5KN5_2),.clk(gclk));
	jdff dff_B_BkYHmE6V4_2(.din(w_dff_B_MbRKR5KN5_2),.dout(w_dff_B_BkYHmE6V4_2),.clk(gclk));
	jdff dff_B_YE2rx8cE6_2(.din(w_dff_B_BkYHmE6V4_2),.dout(w_dff_B_YE2rx8cE6_2),.clk(gclk));
	jdff dff_B_Q2Bm8MuR8_2(.din(w_dff_B_YE2rx8cE6_2),.dout(w_dff_B_Q2Bm8MuR8_2),.clk(gclk));
	jdff dff_B_5MqNYOMH4_2(.din(w_dff_B_Q2Bm8MuR8_2),.dout(w_dff_B_5MqNYOMH4_2),.clk(gclk));
	jdff dff_B_lnxo9GcD3_2(.din(w_dff_B_5MqNYOMH4_2),.dout(w_dff_B_lnxo9GcD3_2),.clk(gclk));
	jdff dff_B_dOovRSgX9_2(.din(w_dff_B_lnxo9GcD3_2),.dout(w_dff_B_dOovRSgX9_2),.clk(gclk));
	jdff dff_B_gllUR0MF3_2(.din(w_dff_B_dOovRSgX9_2),.dout(w_dff_B_gllUR0MF3_2),.clk(gclk));
	jdff dff_B_XnR8pnxw7_2(.din(n1652),.dout(w_dff_B_XnR8pnxw7_2),.clk(gclk));
	jdff dff_B_GR15E4pp6_2(.din(w_dff_B_XnR8pnxw7_2),.dout(w_dff_B_GR15E4pp6_2),.clk(gclk));
	jdff dff_B_PCIhFuYQ6_2(.din(w_dff_B_GR15E4pp6_2),.dout(w_dff_B_PCIhFuYQ6_2),.clk(gclk));
	jdff dff_B_IKYZ6lqQ6_2(.din(w_dff_B_PCIhFuYQ6_2),.dout(w_dff_B_IKYZ6lqQ6_2),.clk(gclk));
	jdff dff_B_E65ue60G1_2(.din(w_dff_B_IKYZ6lqQ6_2),.dout(w_dff_B_E65ue60G1_2),.clk(gclk));
	jdff dff_B_CuRHdUgE3_2(.din(w_dff_B_E65ue60G1_2),.dout(w_dff_B_CuRHdUgE3_2),.clk(gclk));
	jdff dff_B_vf1kuXxr8_2(.din(w_dff_B_CuRHdUgE3_2),.dout(w_dff_B_vf1kuXxr8_2),.clk(gclk));
	jdff dff_B_jnb87pNR1_2(.din(w_dff_B_vf1kuXxr8_2),.dout(w_dff_B_jnb87pNR1_2),.clk(gclk));
	jdff dff_B_8X9VvcrN1_2(.din(w_dff_B_jnb87pNR1_2),.dout(w_dff_B_8X9VvcrN1_2),.clk(gclk));
	jdff dff_B_nrCLN1p26_2(.din(w_dff_B_8X9VvcrN1_2),.dout(w_dff_B_nrCLN1p26_2),.clk(gclk));
	jdff dff_B_yog6ln8E5_2(.din(w_dff_B_nrCLN1p26_2),.dout(w_dff_B_yog6ln8E5_2),.clk(gclk));
	jdff dff_B_pEmW8hLs0_2(.din(w_dff_B_yog6ln8E5_2),.dout(w_dff_B_pEmW8hLs0_2),.clk(gclk));
	jdff dff_B_TkCdXKA67_2(.din(w_dff_B_pEmW8hLs0_2),.dout(w_dff_B_TkCdXKA67_2),.clk(gclk));
	jdff dff_B_FW6cNoW11_2(.din(w_dff_B_TkCdXKA67_2),.dout(w_dff_B_FW6cNoW11_2),.clk(gclk));
	jdff dff_B_ehuOBwyZ0_2(.din(w_dff_B_FW6cNoW11_2),.dout(w_dff_B_ehuOBwyZ0_2),.clk(gclk));
	jdff dff_B_0ZrObZ2m1_2(.din(w_dff_B_ehuOBwyZ0_2),.dout(w_dff_B_0ZrObZ2m1_2),.clk(gclk));
	jdff dff_B_Eq7tGFbb8_2(.din(w_dff_B_0ZrObZ2m1_2),.dout(w_dff_B_Eq7tGFbb8_2),.clk(gclk));
	jdff dff_B_10mGnbdy4_2(.din(w_dff_B_Eq7tGFbb8_2),.dout(w_dff_B_10mGnbdy4_2),.clk(gclk));
	jdff dff_B_cJiyqwCu8_2(.din(w_dff_B_10mGnbdy4_2),.dout(w_dff_B_cJiyqwCu8_2),.clk(gclk));
	jdff dff_B_CVoOe6WP7_2(.din(w_dff_B_cJiyqwCu8_2),.dout(w_dff_B_CVoOe6WP7_2),.clk(gclk));
	jdff dff_B_868FyOFP4_2(.din(w_dff_B_CVoOe6WP7_2),.dout(w_dff_B_868FyOFP4_2),.clk(gclk));
	jdff dff_B_Q08SRK5p4_2(.din(w_dff_B_868FyOFP4_2),.dout(w_dff_B_Q08SRK5p4_2),.clk(gclk));
	jdff dff_B_alGe5RtK7_2(.din(w_dff_B_Q08SRK5p4_2),.dout(w_dff_B_alGe5RtK7_2),.clk(gclk));
	jdff dff_B_Zp6xdwHW2_2(.din(w_dff_B_alGe5RtK7_2),.dout(w_dff_B_Zp6xdwHW2_2),.clk(gclk));
	jdff dff_B_I8DUJgua2_2(.din(w_dff_B_Zp6xdwHW2_2),.dout(w_dff_B_I8DUJgua2_2),.clk(gclk));
	jdff dff_B_31Sj8Rt25_2(.din(w_dff_B_I8DUJgua2_2),.dout(w_dff_B_31Sj8Rt25_2),.clk(gclk));
	jdff dff_B_JV0yl0MZ1_2(.din(w_dff_B_31Sj8Rt25_2),.dout(w_dff_B_JV0yl0MZ1_2),.clk(gclk));
	jdff dff_B_j9x3Q7nm3_2(.din(w_dff_B_JV0yl0MZ1_2),.dout(w_dff_B_j9x3Q7nm3_2),.clk(gclk));
	jdff dff_B_GnXLaZHG8_2(.din(w_dff_B_j9x3Q7nm3_2),.dout(w_dff_B_GnXLaZHG8_2),.clk(gclk));
	jdff dff_B_Z3pLEOEH0_2(.din(w_dff_B_GnXLaZHG8_2),.dout(w_dff_B_Z3pLEOEH0_2),.clk(gclk));
	jdff dff_B_HbzwnA556_2(.din(w_dff_B_Z3pLEOEH0_2),.dout(w_dff_B_HbzwnA556_2),.clk(gclk));
	jdff dff_B_dv1s7Ykx1_2(.din(w_dff_B_HbzwnA556_2),.dout(w_dff_B_dv1s7Ykx1_2),.clk(gclk));
	jdff dff_B_ObRThRGk1_2(.din(w_dff_B_dv1s7Ykx1_2),.dout(w_dff_B_ObRThRGk1_2),.clk(gclk));
	jdff dff_B_XwJ5JWuj3_2(.din(w_dff_B_ObRThRGk1_2),.dout(w_dff_B_XwJ5JWuj3_2),.clk(gclk));
	jdff dff_B_2q4SW0fe1_2(.din(w_dff_B_XwJ5JWuj3_2),.dout(w_dff_B_2q4SW0fe1_2),.clk(gclk));
	jdff dff_B_ocKxbxSA6_2(.din(w_dff_B_2q4SW0fe1_2),.dout(w_dff_B_ocKxbxSA6_2),.clk(gclk));
	jdff dff_B_9PAd5v7J8_2(.din(w_dff_B_ocKxbxSA6_2),.dout(w_dff_B_9PAd5v7J8_2),.clk(gclk));
	jdff dff_B_NufzxXYp2_2(.din(w_dff_B_9PAd5v7J8_2),.dout(w_dff_B_NufzxXYp2_2),.clk(gclk));
	jdff dff_B_IGBSwx534_2(.din(n1651),.dout(w_dff_B_IGBSwx534_2),.clk(gclk));
	jdff dff_B_PRIZboWh1_1(.din(n1649),.dout(w_dff_B_PRIZboWh1_1),.clk(gclk));
	jdff dff_B_NracL9LR4_2(.din(n1591),.dout(w_dff_B_NracL9LR4_2),.clk(gclk));
	jdff dff_B_0NUeyTxa8_2(.din(w_dff_B_NracL9LR4_2),.dout(w_dff_B_0NUeyTxa8_2),.clk(gclk));
	jdff dff_B_zRK2UE0c0_2(.din(w_dff_B_0NUeyTxa8_2),.dout(w_dff_B_zRK2UE0c0_2),.clk(gclk));
	jdff dff_B_FN3IRPQl4_2(.din(w_dff_B_zRK2UE0c0_2),.dout(w_dff_B_FN3IRPQl4_2),.clk(gclk));
	jdff dff_B_jAv1NIka7_2(.din(w_dff_B_FN3IRPQl4_2),.dout(w_dff_B_jAv1NIka7_2),.clk(gclk));
	jdff dff_B_teeeHzWr1_2(.din(w_dff_B_jAv1NIka7_2),.dout(w_dff_B_teeeHzWr1_2),.clk(gclk));
	jdff dff_B_6fvY58Yc2_2(.din(w_dff_B_teeeHzWr1_2),.dout(w_dff_B_6fvY58Yc2_2),.clk(gclk));
	jdff dff_B_Qwudmptu0_2(.din(w_dff_B_6fvY58Yc2_2),.dout(w_dff_B_Qwudmptu0_2),.clk(gclk));
	jdff dff_B_MCD9BKO21_2(.din(w_dff_B_Qwudmptu0_2),.dout(w_dff_B_MCD9BKO21_2),.clk(gclk));
	jdff dff_B_dgyQrOCl3_2(.din(w_dff_B_MCD9BKO21_2),.dout(w_dff_B_dgyQrOCl3_2),.clk(gclk));
	jdff dff_B_caS2ihKx8_2(.din(w_dff_B_dgyQrOCl3_2),.dout(w_dff_B_caS2ihKx8_2),.clk(gclk));
	jdff dff_B_sERGt8je2_2(.din(w_dff_B_caS2ihKx8_2),.dout(w_dff_B_sERGt8je2_2),.clk(gclk));
	jdff dff_B_wse96MkP4_2(.din(w_dff_B_sERGt8je2_2),.dout(w_dff_B_wse96MkP4_2),.clk(gclk));
	jdff dff_B_YVoBk29T8_2(.din(w_dff_B_wse96MkP4_2),.dout(w_dff_B_YVoBk29T8_2),.clk(gclk));
	jdff dff_B_rNnEPmTd7_2(.din(w_dff_B_YVoBk29T8_2),.dout(w_dff_B_rNnEPmTd7_2),.clk(gclk));
	jdff dff_B_91DkQBZA9_2(.din(w_dff_B_rNnEPmTd7_2),.dout(w_dff_B_91DkQBZA9_2),.clk(gclk));
	jdff dff_B_WzkmCQyW8_2(.din(w_dff_B_91DkQBZA9_2),.dout(w_dff_B_WzkmCQyW8_2),.clk(gclk));
	jdff dff_B_2Mjyl81S8_2(.din(w_dff_B_WzkmCQyW8_2),.dout(w_dff_B_2Mjyl81S8_2),.clk(gclk));
	jdff dff_B_RQRhDMSc3_2(.din(w_dff_B_2Mjyl81S8_2),.dout(w_dff_B_RQRhDMSc3_2),.clk(gclk));
	jdff dff_B_xLWUme7f7_2(.din(w_dff_B_RQRhDMSc3_2),.dout(w_dff_B_xLWUme7f7_2),.clk(gclk));
	jdff dff_B_M4pE5sV05_2(.din(w_dff_B_xLWUme7f7_2),.dout(w_dff_B_M4pE5sV05_2),.clk(gclk));
	jdff dff_B_FiRVVw5h1_2(.din(w_dff_B_M4pE5sV05_2),.dout(w_dff_B_FiRVVw5h1_2),.clk(gclk));
	jdff dff_B_4mzbmJPp6_2(.din(w_dff_B_FiRVVw5h1_2),.dout(w_dff_B_4mzbmJPp6_2),.clk(gclk));
	jdff dff_B_AOlAwuXk7_2(.din(w_dff_B_4mzbmJPp6_2),.dout(w_dff_B_AOlAwuXk7_2),.clk(gclk));
	jdff dff_B_BTHarfsS1_2(.din(w_dff_B_AOlAwuXk7_2),.dout(w_dff_B_BTHarfsS1_2),.clk(gclk));
	jdff dff_B_4UvEFnxN4_2(.din(w_dff_B_BTHarfsS1_2),.dout(w_dff_B_4UvEFnxN4_2),.clk(gclk));
	jdff dff_B_TbSFipsC5_2(.din(w_dff_B_4UvEFnxN4_2),.dout(w_dff_B_TbSFipsC5_2),.clk(gclk));
	jdff dff_B_qCxYuplw6_2(.din(w_dff_B_TbSFipsC5_2),.dout(w_dff_B_qCxYuplw6_2),.clk(gclk));
	jdff dff_B_02PCvWrG3_2(.din(w_dff_B_qCxYuplw6_2),.dout(w_dff_B_02PCvWrG3_2),.clk(gclk));
	jdff dff_B_TwB6wEks6_2(.din(w_dff_B_02PCvWrG3_2),.dout(w_dff_B_TwB6wEks6_2),.clk(gclk));
	jdff dff_B_FDz5upXD3_2(.din(w_dff_B_TwB6wEks6_2),.dout(w_dff_B_FDz5upXD3_2),.clk(gclk));
	jdff dff_B_SiabVybH4_2(.din(w_dff_B_FDz5upXD3_2),.dout(w_dff_B_SiabVybH4_2),.clk(gclk));
	jdff dff_B_VraM9NXu3_2(.din(w_dff_B_SiabVybH4_2),.dout(w_dff_B_VraM9NXu3_2),.clk(gclk));
	jdff dff_B_qJzGZ17T5_2(.din(w_dff_B_VraM9NXu3_2),.dout(w_dff_B_qJzGZ17T5_2),.clk(gclk));
	jdff dff_B_poyiy4tx3_2(.din(w_dff_B_qJzGZ17T5_2),.dout(w_dff_B_poyiy4tx3_2),.clk(gclk));
	jdff dff_B_o269yUIt0_1(.din(n1597),.dout(w_dff_B_o269yUIt0_1),.clk(gclk));
	jdff dff_B_F8seNExg6_1(.din(w_dff_B_o269yUIt0_1),.dout(w_dff_B_F8seNExg6_1),.clk(gclk));
	jdff dff_B_CKhLp4CL1_2(.din(n1596),.dout(w_dff_B_CKhLp4CL1_2),.clk(gclk));
	jdff dff_B_xRDHZbVN6_2(.din(w_dff_B_CKhLp4CL1_2),.dout(w_dff_B_xRDHZbVN6_2),.clk(gclk));
	jdff dff_B_oqi26wSG4_2(.din(w_dff_B_xRDHZbVN6_2),.dout(w_dff_B_oqi26wSG4_2),.clk(gclk));
	jdff dff_B_9tYi3ZoF6_2(.din(w_dff_B_oqi26wSG4_2),.dout(w_dff_B_9tYi3ZoF6_2),.clk(gclk));
	jdff dff_B_wZVMEj6s0_2(.din(w_dff_B_9tYi3ZoF6_2),.dout(w_dff_B_wZVMEj6s0_2),.clk(gclk));
	jdff dff_B_tJibNlXw0_2(.din(w_dff_B_wZVMEj6s0_2),.dout(w_dff_B_tJibNlXw0_2),.clk(gclk));
	jdff dff_B_JbuW4FVZ4_2(.din(w_dff_B_tJibNlXw0_2),.dout(w_dff_B_JbuW4FVZ4_2),.clk(gclk));
	jdff dff_B_JMyUr2pa2_2(.din(w_dff_B_JbuW4FVZ4_2),.dout(w_dff_B_JMyUr2pa2_2),.clk(gclk));
	jdff dff_B_spw74YZt9_2(.din(w_dff_B_JMyUr2pa2_2),.dout(w_dff_B_spw74YZt9_2),.clk(gclk));
	jdff dff_B_68BhCiDL5_2(.din(w_dff_B_spw74YZt9_2),.dout(w_dff_B_68BhCiDL5_2),.clk(gclk));
	jdff dff_B_9pAHtDJY3_2(.din(w_dff_B_68BhCiDL5_2),.dout(w_dff_B_9pAHtDJY3_2),.clk(gclk));
	jdff dff_B_tD8IOVpw4_2(.din(w_dff_B_9pAHtDJY3_2),.dout(w_dff_B_tD8IOVpw4_2),.clk(gclk));
	jdff dff_B_lFHHKp1E1_2(.din(w_dff_B_tD8IOVpw4_2),.dout(w_dff_B_lFHHKp1E1_2),.clk(gclk));
	jdff dff_B_sYNlZP2V8_2(.din(w_dff_B_lFHHKp1E1_2),.dout(w_dff_B_sYNlZP2V8_2),.clk(gclk));
	jdff dff_B_6fJPR5jL1_2(.din(w_dff_B_sYNlZP2V8_2),.dout(w_dff_B_6fJPR5jL1_2),.clk(gclk));
	jdff dff_B_Z1351Jwl1_2(.din(w_dff_B_6fJPR5jL1_2),.dout(w_dff_B_Z1351Jwl1_2),.clk(gclk));
	jdff dff_B_NAhqd4hB7_2(.din(w_dff_B_Z1351Jwl1_2),.dout(w_dff_B_NAhqd4hB7_2),.clk(gclk));
	jdff dff_B_uftwVYDF0_2(.din(w_dff_B_NAhqd4hB7_2),.dout(w_dff_B_uftwVYDF0_2),.clk(gclk));
	jdff dff_B_YTM6FdhP4_2(.din(w_dff_B_uftwVYDF0_2),.dout(w_dff_B_YTM6FdhP4_2),.clk(gclk));
	jdff dff_B_XT5l0IX35_2(.din(w_dff_B_YTM6FdhP4_2),.dout(w_dff_B_XT5l0IX35_2),.clk(gclk));
	jdff dff_B_gfi2GPms9_2(.din(w_dff_B_XT5l0IX35_2),.dout(w_dff_B_gfi2GPms9_2),.clk(gclk));
	jdff dff_B_7LGXwjJU3_2(.din(w_dff_B_gfi2GPms9_2),.dout(w_dff_B_7LGXwjJU3_2),.clk(gclk));
	jdff dff_B_9Bl4KFyY8_2(.din(w_dff_B_7LGXwjJU3_2),.dout(w_dff_B_9Bl4KFyY8_2),.clk(gclk));
	jdff dff_B_P7fVqXY20_2(.din(w_dff_B_9Bl4KFyY8_2),.dout(w_dff_B_P7fVqXY20_2),.clk(gclk));
	jdff dff_B_bcNGexlG7_2(.din(w_dff_B_P7fVqXY20_2),.dout(w_dff_B_bcNGexlG7_2),.clk(gclk));
	jdff dff_B_qkyEtRzg8_2(.din(w_dff_B_bcNGexlG7_2),.dout(w_dff_B_qkyEtRzg8_2),.clk(gclk));
	jdff dff_B_5zXY9Bby4_2(.din(w_dff_B_qkyEtRzg8_2),.dout(w_dff_B_5zXY9Bby4_2),.clk(gclk));
	jdff dff_B_I9nvUdiI9_2(.din(w_dff_B_5zXY9Bby4_2),.dout(w_dff_B_I9nvUdiI9_2),.clk(gclk));
	jdff dff_B_Wzt3jgkN5_2(.din(w_dff_B_I9nvUdiI9_2),.dout(w_dff_B_Wzt3jgkN5_2),.clk(gclk));
	jdff dff_B_qa9CpgJ81_2(.din(w_dff_B_Wzt3jgkN5_2),.dout(w_dff_B_qa9CpgJ81_2),.clk(gclk));
	jdff dff_B_4MP7TjJv7_2(.din(w_dff_B_qa9CpgJ81_2),.dout(w_dff_B_4MP7TjJv7_2),.clk(gclk));
	jdff dff_B_k33KKcJH0_2(.din(w_dff_B_4MP7TjJv7_2),.dout(w_dff_B_k33KKcJH0_2),.clk(gclk));
	jdff dff_B_z5sIHDtl4_2(.din(n1595),.dout(w_dff_B_z5sIHDtl4_2),.clk(gclk));
	jdff dff_B_ceOKQeDm3_2(.din(w_dff_B_z5sIHDtl4_2),.dout(w_dff_B_ceOKQeDm3_2),.clk(gclk));
	jdff dff_B_OIwOBmQ74_2(.din(w_dff_B_ceOKQeDm3_2),.dout(w_dff_B_OIwOBmQ74_2),.clk(gclk));
	jdff dff_B_3VDPHyRE7_2(.din(w_dff_B_OIwOBmQ74_2),.dout(w_dff_B_3VDPHyRE7_2),.clk(gclk));
	jdff dff_B_45xF50ic2_2(.din(w_dff_B_3VDPHyRE7_2),.dout(w_dff_B_45xF50ic2_2),.clk(gclk));
	jdff dff_B_OkN2jMdi2_2(.din(w_dff_B_45xF50ic2_2),.dout(w_dff_B_OkN2jMdi2_2),.clk(gclk));
	jdff dff_B_oH16Peh98_2(.din(w_dff_B_OkN2jMdi2_2),.dout(w_dff_B_oH16Peh98_2),.clk(gclk));
	jdff dff_B_LR98fBSb3_2(.din(w_dff_B_oH16Peh98_2),.dout(w_dff_B_LR98fBSb3_2),.clk(gclk));
	jdff dff_B_m2VBFUQB9_2(.din(w_dff_B_LR98fBSb3_2),.dout(w_dff_B_m2VBFUQB9_2),.clk(gclk));
	jdff dff_B_ofV171bt6_2(.din(w_dff_B_m2VBFUQB9_2),.dout(w_dff_B_ofV171bt6_2),.clk(gclk));
	jdff dff_B_y2q5XDX69_2(.din(w_dff_B_ofV171bt6_2),.dout(w_dff_B_y2q5XDX69_2),.clk(gclk));
	jdff dff_B_XP0fBp7V2_2(.din(w_dff_B_y2q5XDX69_2),.dout(w_dff_B_XP0fBp7V2_2),.clk(gclk));
	jdff dff_B_W8vqF5TY8_2(.din(w_dff_B_XP0fBp7V2_2),.dout(w_dff_B_W8vqF5TY8_2),.clk(gclk));
	jdff dff_B_ieeJvNcR6_2(.din(w_dff_B_W8vqF5TY8_2),.dout(w_dff_B_ieeJvNcR6_2),.clk(gclk));
	jdff dff_B_qfeuUqiQ7_2(.din(w_dff_B_ieeJvNcR6_2),.dout(w_dff_B_qfeuUqiQ7_2),.clk(gclk));
	jdff dff_B_rCIUZCPg8_2(.din(w_dff_B_qfeuUqiQ7_2),.dout(w_dff_B_rCIUZCPg8_2),.clk(gclk));
	jdff dff_B_RJ14PlcM2_2(.din(w_dff_B_rCIUZCPg8_2),.dout(w_dff_B_RJ14PlcM2_2),.clk(gclk));
	jdff dff_B_3ZsxmYPr5_2(.din(w_dff_B_RJ14PlcM2_2),.dout(w_dff_B_3ZsxmYPr5_2),.clk(gclk));
	jdff dff_B_M8SpTF1E4_2(.din(w_dff_B_3ZsxmYPr5_2),.dout(w_dff_B_M8SpTF1E4_2),.clk(gclk));
	jdff dff_B_cXHeC0i30_2(.din(w_dff_B_M8SpTF1E4_2),.dout(w_dff_B_cXHeC0i30_2),.clk(gclk));
	jdff dff_B_3pZV89Ul7_2(.din(w_dff_B_cXHeC0i30_2),.dout(w_dff_B_3pZV89Ul7_2),.clk(gclk));
	jdff dff_B_vKJCAfLp4_2(.din(w_dff_B_3pZV89Ul7_2),.dout(w_dff_B_vKJCAfLp4_2),.clk(gclk));
	jdff dff_B_YlPJwVTa2_2(.din(w_dff_B_vKJCAfLp4_2),.dout(w_dff_B_YlPJwVTa2_2),.clk(gclk));
	jdff dff_B_Ag52ToH48_2(.din(w_dff_B_YlPJwVTa2_2),.dout(w_dff_B_Ag52ToH48_2),.clk(gclk));
	jdff dff_B_In1xradN7_2(.din(w_dff_B_Ag52ToH48_2),.dout(w_dff_B_In1xradN7_2),.clk(gclk));
	jdff dff_B_Ssv5yBim0_2(.din(w_dff_B_In1xradN7_2),.dout(w_dff_B_Ssv5yBim0_2),.clk(gclk));
	jdff dff_B_eW05ITvY5_2(.din(w_dff_B_Ssv5yBim0_2),.dout(w_dff_B_eW05ITvY5_2),.clk(gclk));
	jdff dff_B_VOxdsDCI2_2(.din(w_dff_B_eW05ITvY5_2),.dout(w_dff_B_VOxdsDCI2_2),.clk(gclk));
	jdff dff_B_u4nTYRW40_2(.din(w_dff_B_VOxdsDCI2_2),.dout(w_dff_B_u4nTYRW40_2),.clk(gclk));
	jdff dff_B_3WN5ZGwT8_2(.din(w_dff_B_u4nTYRW40_2),.dout(w_dff_B_3WN5ZGwT8_2),.clk(gclk));
	jdff dff_B_qENnCH9B0_2(.din(w_dff_B_3WN5ZGwT8_2),.dout(w_dff_B_qENnCH9B0_2),.clk(gclk));
	jdff dff_B_KU1oYdmK9_2(.din(w_dff_B_qENnCH9B0_2),.dout(w_dff_B_KU1oYdmK9_2),.clk(gclk));
	jdff dff_B_PCSE2ZYu5_2(.din(w_dff_B_KU1oYdmK9_2),.dout(w_dff_B_PCSE2ZYu5_2),.clk(gclk));
	jdff dff_B_Dk0tMq5b9_2(.din(w_dff_B_PCSE2ZYu5_2),.dout(w_dff_B_Dk0tMq5b9_2),.clk(gclk));
	jdff dff_B_896xBcra0_2(.din(n1594),.dout(w_dff_B_896xBcra0_2),.clk(gclk));
	jdff dff_B_McwKnVtr5_1(.din(n1592),.dout(w_dff_B_McwKnVtr5_1),.clk(gclk));
	jdff dff_B_bZ6WEBNu7_2(.din(n1527),.dout(w_dff_B_bZ6WEBNu7_2),.clk(gclk));
	jdff dff_B_xzEVptqB3_2(.din(w_dff_B_bZ6WEBNu7_2),.dout(w_dff_B_xzEVptqB3_2),.clk(gclk));
	jdff dff_B_ea4bv41s1_2(.din(w_dff_B_xzEVptqB3_2),.dout(w_dff_B_ea4bv41s1_2),.clk(gclk));
	jdff dff_B_EEK7yyOR7_2(.din(w_dff_B_ea4bv41s1_2),.dout(w_dff_B_EEK7yyOR7_2),.clk(gclk));
	jdff dff_B_G5rB0ymr7_2(.din(w_dff_B_EEK7yyOR7_2),.dout(w_dff_B_G5rB0ymr7_2),.clk(gclk));
	jdff dff_B_GLf2xhsH2_2(.din(w_dff_B_G5rB0ymr7_2),.dout(w_dff_B_GLf2xhsH2_2),.clk(gclk));
	jdff dff_B_dXmZjGWX2_2(.din(w_dff_B_GLf2xhsH2_2),.dout(w_dff_B_dXmZjGWX2_2),.clk(gclk));
	jdff dff_B_3muGzQyA3_2(.din(w_dff_B_dXmZjGWX2_2),.dout(w_dff_B_3muGzQyA3_2),.clk(gclk));
	jdff dff_B_2FDjoapF1_2(.din(w_dff_B_3muGzQyA3_2),.dout(w_dff_B_2FDjoapF1_2),.clk(gclk));
	jdff dff_B_KEI8AuKV3_2(.din(w_dff_B_2FDjoapF1_2),.dout(w_dff_B_KEI8AuKV3_2),.clk(gclk));
	jdff dff_B_VDBAvZfu0_2(.din(w_dff_B_KEI8AuKV3_2),.dout(w_dff_B_VDBAvZfu0_2),.clk(gclk));
	jdff dff_B_NgLvRoqM9_2(.din(w_dff_B_VDBAvZfu0_2),.dout(w_dff_B_NgLvRoqM9_2),.clk(gclk));
	jdff dff_B_2ab4lZzW5_2(.din(w_dff_B_NgLvRoqM9_2),.dout(w_dff_B_2ab4lZzW5_2),.clk(gclk));
	jdff dff_B_BrQETskv6_2(.din(w_dff_B_2ab4lZzW5_2),.dout(w_dff_B_BrQETskv6_2),.clk(gclk));
	jdff dff_B_7Y5AYlhf9_2(.din(w_dff_B_BrQETskv6_2),.dout(w_dff_B_7Y5AYlhf9_2),.clk(gclk));
	jdff dff_B_ewG0hSRH3_2(.din(w_dff_B_7Y5AYlhf9_2),.dout(w_dff_B_ewG0hSRH3_2),.clk(gclk));
	jdff dff_B_WPS5zvIH6_2(.din(w_dff_B_ewG0hSRH3_2),.dout(w_dff_B_WPS5zvIH6_2),.clk(gclk));
	jdff dff_B_CBfMUNlC8_2(.din(w_dff_B_WPS5zvIH6_2),.dout(w_dff_B_CBfMUNlC8_2),.clk(gclk));
	jdff dff_B_Q7SK2WP14_2(.din(w_dff_B_CBfMUNlC8_2),.dout(w_dff_B_Q7SK2WP14_2),.clk(gclk));
	jdff dff_B_9RdwN7NJ2_2(.din(w_dff_B_Q7SK2WP14_2),.dout(w_dff_B_9RdwN7NJ2_2),.clk(gclk));
	jdff dff_B_utU1DPPF8_2(.din(w_dff_B_9RdwN7NJ2_2),.dout(w_dff_B_utU1DPPF8_2),.clk(gclk));
	jdff dff_B_dCgsYsmP2_2(.din(w_dff_B_utU1DPPF8_2),.dout(w_dff_B_dCgsYsmP2_2),.clk(gclk));
	jdff dff_B_MD0JMfIu9_2(.din(w_dff_B_dCgsYsmP2_2),.dout(w_dff_B_MD0JMfIu9_2),.clk(gclk));
	jdff dff_B_gBZwyyzt0_2(.din(w_dff_B_MD0JMfIu9_2),.dout(w_dff_B_gBZwyyzt0_2),.clk(gclk));
	jdff dff_B_AhXiICfe0_2(.din(w_dff_B_gBZwyyzt0_2),.dout(w_dff_B_AhXiICfe0_2),.clk(gclk));
	jdff dff_B_v8yKt9CW2_2(.din(w_dff_B_AhXiICfe0_2),.dout(w_dff_B_v8yKt9CW2_2),.clk(gclk));
	jdff dff_B_lMxW56rO1_2(.din(w_dff_B_v8yKt9CW2_2),.dout(w_dff_B_lMxW56rO1_2),.clk(gclk));
	jdff dff_B_M4PoGaBP3_2(.din(w_dff_B_lMxW56rO1_2),.dout(w_dff_B_M4PoGaBP3_2),.clk(gclk));
	jdff dff_B_XT0Pvyyn6_2(.din(w_dff_B_M4PoGaBP3_2),.dout(w_dff_B_XT0Pvyyn6_2),.clk(gclk));
	jdff dff_B_ZOu315Ty6_2(.din(w_dff_B_XT0Pvyyn6_2),.dout(w_dff_B_ZOu315Ty6_2),.clk(gclk));
	jdff dff_B_ugBGSNfa3_2(.din(w_dff_B_ZOu315Ty6_2),.dout(w_dff_B_ugBGSNfa3_2),.clk(gclk));
	jdff dff_B_qoDRJVxL7_1(.din(n1533),.dout(w_dff_B_qoDRJVxL7_1),.clk(gclk));
	jdff dff_B_2ezTw40N3_1(.din(w_dff_B_qoDRJVxL7_1),.dout(w_dff_B_2ezTw40N3_1),.clk(gclk));
	jdff dff_B_58UfveQP3_2(.din(n1532),.dout(w_dff_B_58UfveQP3_2),.clk(gclk));
	jdff dff_B_ADp3j63K0_2(.din(w_dff_B_58UfveQP3_2),.dout(w_dff_B_ADp3j63K0_2),.clk(gclk));
	jdff dff_B_i7itV8O29_2(.din(w_dff_B_ADp3j63K0_2),.dout(w_dff_B_i7itV8O29_2),.clk(gclk));
	jdff dff_B_UAApKXy27_2(.din(w_dff_B_i7itV8O29_2),.dout(w_dff_B_UAApKXy27_2),.clk(gclk));
	jdff dff_B_ualVowA88_2(.din(w_dff_B_UAApKXy27_2),.dout(w_dff_B_ualVowA88_2),.clk(gclk));
	jdff dff_B_QcDY9brj0_2(.din(w_dff_B_ualVowA88_2),.dout(w_dff_B_QcDY9brj0_2),.clk(gclk));
	jdff dff_B_GdyBCVIk3_2(.din(w_dff_B_QcDY9brj0_2),.dout(w_dff_B_GdyBCVIk3_2),.clk(gclk));
	jdff dff_B_TiogwJfi9_2(.din(w_dff_B_GdyBCVIk3_2),.dout(w_dff_B_TiogwJfi9_2),.clk(gclk));
	jdff dff_B_gPw2qPn51_2(.din(w_dff_B_TiogwJfi9_2),.dout(w_dff_B_gPw2qPn51_2),.clk(gclk));
	jdff dff_B_3lSYcOmN9_2(.din(w_dff_B_gPw2qPn51_2),.dout(w_dff_B_3lSYcOmN9_2),.clk(gclk));
	jdff dff_B_RqrDtsIH9_2(.din(w_dff_B_3lSYcOmN9_2),.dout(w_dff_B_RqrDtsIH9_2),.clk(gclk));
	jdff dff_B_nqltyu9W7_2(.din(w_dff_B_RqrDtsIH9_2),.dout(w_dff_B_nqltyu9W7_2),.clk(gclk));
	jdff dff_B_Llt5KdTM8_2(.din(w_dff_B_nqltyu9W7_2),.dout(w_dff_B_Llt5KdTM8_2),.clk(gclk));
	jdff dff_B_Cbi5UaaD9_2(.din(w_dff_B_Llt5KdTM8_2),.dout(w_dff_B_Cbi5UaaD9_2),.clk(gclk));
	jdff dff_B_Y1QeJM9E6_2(.din(w_dff_B_Cbi5UaaD9_2),.dout(w_dff_B_Y1QeJM9E6_2),.clk(gclk));
	jdff dff_B_dPpWhZ6g2_2(.din(w_dff_B_Y1QeJM9E6_2),.dout(w_dff_B_dPpWhZ6g2_2),.clk(gclk));
	jdff dff_B_qwjEigGV2_2(.din(w_dff_B_dPpWhZ6g2_2),.dout(w_dff_B_qwjEigGV2_2),.clk(gclk));
	jdff dff_B_8rUETevF1_2(.din(w_dff_B_qwjEigGV2_2),.dout(w_dff_B_8rUETevF1_2),.clk(gclk));
	jdff dff_B_igXJoIem2_2(.din(w_dff_B_8rUETevF1_2),.dout(w_dff_B_igXJoIem2_2),.clk(gclk));
	jdff dff_B_uZnQPvYp7_2(.din(w_dff_B_igXJoIem2_2),.dout(w_dff_B_uZnQPvYp7_2),.clk(gclk));
	jdff dff_B_y8rwqxq31_2(.din(w_dff_B_uZnQPvYp7_2),.dout(w_dff_B_y8rwqxq31_2),.clk(gclk));
	jdff dff_B_FKTrVXhZ8_2(.din(w_dff_B_y8rwqxq31_2),.dout(w_dff_B_FKTrVXhZ8_2),.clk(gclk));
	jdff dff_B_3nv21eCL6_2(.din(w_dff_B_FKTrVXhZ8_2),.dout(w_dff_B_3nv21eCL6_2),.clk(gclk));
	jdff dff_B_F19CCd8T2_2(.din(w_dff_B_3nv21eCL6_2),.dout(w_dff_B_F19CCd8T2_2),.clk(gclk));
	jdff dff_B_kFLHSc7L3_2(.din(w_dff_B_F19CCd8T2_2),.dout(w_dff_B_kFLHSc7L3_2),.clk(gclk));
	jdff dff_B_VeEQDDQO3_2(.din(w_dff_B_kFLHSc7L3_2),.dout(w_dff_B_VeEQDDQO3_2),.clk(gclk));
	jdff dff_B_vzwqLw0d9_2(.din(w_dff_B_VeEQDDQO3_2),.dout(w_dff_B_vzwqLw0d9_2),.clk(gclk));
	jdff dff_B_7nodYucn0_2(.din(w_dff_B_vzwqLw0d9_2),.dout(w_dff_B_7nodYucn0_2),.clk(gclk));
	jdff dff_B_60a6Xq1l9_2(.din(n1531),.dout(w_dff_B_60a6Xq1l9_2),.clk(gclk));
	jdff dff_B_hodZAB5S2_2(.din(w_dff_B_60a6Xq1l9_2),.dout(w_dff_B_hodZAB5S2_2),.clk(gclk));
	jdff dff_B_KXkbuGap5_2(.din(w_dff_B_hodZAB5S2_2),.dout(w_dff_B_KXkbuGap5_2),.clk(gclk));
	jdff dff_B_q24DgdNX2_2(.din(w_dff_B_KXkbuGap5_2),.dout(w_dff_B_q24DgdNX2_2),.clk(gclk));
	jdff dff_B_lI9Asubr5_2(.din(w_dff_B_q24DgdNX2_2),.dout(w_dff_B_lI9Asubr5_2),.clk(gclk));
	jdff dff_B_C9nG3yxR4_2(.din(w_dff_B_lI9Asubr5_2),.dout(w_dff_B_C9nG3yxR4_2),.clk(gclk));
	jdff dff_B_YcRguUlg1_2(.din(w_dff_B_C9nG3yxR4_2),.dout(w_dff_B_YcRguUlg1_2),.clk(gclk));
	jdff dff_B_3vZBWnPc9_2(.din(w_dff_B_YcRguUlg1_2),.dout(w_dff_B_3vZBWnPc9_2),.clk(gclk));
	jdff dff_B_pbwmV0Pd3_2(.din(w_dff_B_3vZBWnPc9_2),.dout(w_dff_B_pbwmV0Pd3_2),.clk(gclk));
	jdff dff_B_N8ZhIHqc4_2(.din(w_dff_B_pbwmV0Pd3_2),.dout(w_dff_B_N8ZhIHqc4_2),.clk(gclk));
	jdff dff_B_f70K9my72_2(.din(w_dff_B_N8ZhIHqc4_2),.dout(w_dff_B_f70K9my72_2),.clk(gclk));
	jdff dff_B_irg1wuLv2_2(.din(w_dff_B_f70K9my72_2),.dout(w_dff_B_irg1wuLv2_2),.clk(gclk));
	jdff dff_B_z4IAjJXj2_2(.din(w_dff_B_irg1wuLv2_2),.dout(w_dff_B_z4IAjJXj2_2),.clk(gclk));
	jdff dff_B_cbLsPkEf9_2(.din(w_dff_B_z4IAjJXj2_2),.dout(w_dff_B_cbLsPkEf9_2),.clk(gclk));
	jdff dff_B_BRob48bd0_2(.din(w_dff_B_cbLsPkEf9_2),.dout(w_dff_B_BRob48bd0_2),.clk(gclk));
	jdff dff_B_9uiwO0Nl7_2(.din(w_dff_B_BRob48bd0_2),.dout(w_dff_B_9uiwO0Nl7_2),.clk(gclk));
	jdff dff_B_SLiuM5ML4_2(.din(w_dff_B_9uiwO0Nl7_2),.dout(w_dff_B_SLiuM5ML4_2),.clk(gclk));
	jdff dff_B_KYcwbfYM0_2(.din(w_dff_B_SLiuM5ML4_2),.dout(w_dff_B_KYcwbfYM0_2),.clk(gclk));
	jdff dff_B_zRRdla247_2(.din(w_dff_B_KYcwbfYM0_2),.dout(w_dff_B_zRRdla247_2),.clk(gclk));
	jdff dff_B_VYh0AFar9_2(.din(w_dff_B_zRRdla247_2),.dout(w_dff_B_VYh0AFar9_2),.clk(gclk));
	jdff dff_B_BvHwI7er9_2(.din(w_dff_B_VYh0AFar9_2),.dout(w_dff_B_BvHwI7er9_2),.clk(gclk));
	jdff dff_B_SSqH70Pr3_2(.din(w_dff_B_BvHwI7er9_2),.dout(w_dff_B_SSqH70Pr3_2),.clk(gclk));
	jdff dff_B_s0avIIv43_2(.din(w_dff_B_SSqH70Pr3_2),.dout(w_dff_B_s0avIIv43_2),.clk(gclk));
	jdff dff_B_e6Yqgxd20_2(.din(w_dff_B_s0avIIv43_2),.dout(w_dff_B_e6Yqgxd20_2),.clk(gclk));
	jdff dff_B_C41PjQDs7_2(.din(w_dff_B_e6Yqgxd20_2),.dout(w_dff_B_C41PjQDs7_2),.clk(gclk));
	jdff dff_B_voCVrfKC1_2(.din(w_dff_B_C41PjQDs7_2),.dout(w_dff_B_voCVrfKC1_2),.clk(gclk));
	jdff dff_B_Kf2JBVjW1_2(.din(w_dff_B_voCVrfKC1_2),.dout(w_dff_B_Kf2JBVjW1_2),.clk(gclk));
	jdff dff_B_oFa4G7VG1_2(.din(w_dff_B_Kf2JBVjW1_2),.dout(w_dff_B_oFa4G7VG1_2),.clk(gclk));
	jdff dff_B_3CPhrYIH7_2(.din(w_dff_B_oFa4G7VG1_2),.dout(w_dff_B_3CPhrYIH7_2),.clk(gclk));
	jdff dff_B_8YzArT0w9_2(.din(w_dff_B_3CPhrYIH7_2),.dout(w_dff_B_8YzArT0w9_2),.clk(gclk));
	jdff dff_B_jyCedYn23_2(.din(n1530),.dout(w_dff_B_jyCedYn23_2),.clk(gclk));
	jdff dff_B_4ZGyLYI34_1(.din(n1528),.dout(w_dff_B_4ZGyLYI34_1),.clk(gclk));
	jdff dff_B_qFNYwrEz8_2(.din(n1456),.dout(w_dff_B_qFNYwrEz8_2),.clk(gclk));
	jdff dff_B_aPMWol1E1_2(.din(w_dff_B_qFNYwrEz8_2),.dout(w_dff_B_aPMWol1E1_2),.clk(gclk));
	jdff dff_B_YHzQ0G6b9_2(.din(w_dff_B_aPMWol1E1_2),.dout(w_dff_B_YHzQ0G6b9_2),.clk(gclk));
	jdff dff_B_7x82HizO4_2(.din(w_dff_B_YHzQ0G6b9_2),.dout(w_dff_B_7x82HizO4_2),.clk(gclk));
	jdff dff_B_trzPZ1DV9_2(.din(w_dff_B_7x82HizO4_2),.dout(w_dff_B_trzPZ1DV9_2),.clk(gclk));
	jdff dff_B_iTpLJomj2_2(.din(w_dff_B_trzPZ1DV9_2),.dout(w_dff_B_iTpLJomj2_2),.clk(gclk));
	jdff dff_B_Noac6bpN9_2(.din(w_dff_B_iTpLJomj2_2),.dout(w_dff_B_Noac6bpN9_2),.clk(gclk));
	jdff dff_B_ziRsvjyZ2_2(.din(w_dff_B_Noac6bpN9_2),.dout(w_dff_B_ziRsvjyZ2_2),.clk(gclk));
	jdff dff_B_tY7iefEe6_2(.din(w_dff_B_ziRsvjyZ2_2),.dout(w_dff_B_tY7iefEe6_2),.clk(gclk));
	jdff dff_B_sTQAvUcs4_2(.din(w_dff_B_tY7iefEe6_2),.dout(w_dff_B_sTQAvUcs4_2),.clk(gclk));
	jdff dff_B_mXctcUt55_2(.din(w_dff_B_sTQAvUcs4_2),.dout(w_dff_B_mXctcUt55_2),.clk(gclk));
	jdff dff_B_29Y4etSI2_2(.din(w_dff_B_mXctcUt55_2),.dout(w_dff_B_29Y4etSI2_2),.clk(gclk));
	jdff dff_B_WuFtF8pK6_2(.din(w_dff_B_29Y4etSI2_2),.dout(w_dff_B_WuFtF8pK6_2),.clk(gclk));
	jdff dff_B_zO4t1JEV1_2(.din(w_dff_B_WuFtF8pK6_2),.dout(w_dff_B_zO4t1JEV1_2),.clk(gclk));
	jdff dff_B_Hb4tDzjv1_2(.din(w_dff_B_zO4t1JEV1_2),.dout(w_dff_B_Hb4tDzjv1_2),.clk(gclk));
	jdff dff_B_mnmD1hQL7_2(.din(w_dff_B_Hb4tDzjv1_2),.dout(w_dff_B_mnmD1hQL7_2),.clk(gclk));
	jdff dff_B_mMfPWLG28_2(.din(w_dff_B_mnmD1hQL7_2),.dout(w_dff_B_mMfPWLG28_2),.clk(gclk));
	jdff dff_B_F3GEOyI63_2(.din(w_dff_B_mMfPWLG28_2),.dout(w_dff_B_F3GEOyI63_2),.clk(gclk));
	jdff dff_B_QeSoVTIQ9_2(.din(w_dff_B_F3GEOyI63_2),.dout(w_dff_B_QeSoVTIQ9_2),.clk(gclk));
	jdff dff_B_PXKRWx8c6_2(.din(w_dff_B_QeSoVTIQ9_2),.dout(w_dff_B_PXKRWx8c6_2),.clk(gclk));
	jdff dff_B_ofihC0d07_2(.din(w_dff_B_PXKRWx8c6_2),.dout(w_dff_B_ofihC0d07_2),.clk(gclk));
	jdff dff_B_c656eRfT1_2(.din(w_dff_B_ofihC0d07_2),.dout(w_dff_B_c656eRfT1_2),.clk(gclk));
	jdff dff_B_lOISoo5H7_2(.din(w_dff_B_c656eRfT1_2),.dout(w_dff_B_lOISoo5H7_2),.clk(gclk));
	jdff dff_B_rPZS3WR15_2(.din(w_dff_B_lOISoo5H7_2),.dout(w_dff_B_rPZS3WR15_2),.clk(gclk));
	jdff dff_B_t3HreJNU1_2(.din(w_dff_B_rPZS3WR15_2),.dout(w_dff_B_t3HreJNU1_2),.clk(gclk));
	jdff dff_B_gN63ag3Z0_2(.din(w_dff_B_t3HreJNU1_2),.dout(w_dff_B_gN63ag3Z0_2),.clk(gclk));
	jdff dff_B_FDLZUWT77_2(.din(w_dff_B_gN63ag3Z0_2),.dout(w_dff_B_FDLZUWT77_2),.clk(gclk));
	jdff dff_B_VA2S6U9k3_1(.din(n1462),.dout(w_dff_B_VA2S6U9k3_1),.clk(gclk));
	jdff dff_B_RSFFa2ch4_1(.din(w_dff_B_VA2S6U9k3_1),.dout(w_dff_B_RSFFa2ch4_1),.clk(gclk));
	jdff dff_B_qYTGGBHQ4_2(.din(n1461),.dout(w_dff_B_qYTGGBHQ4_2),.clk(gclk));
	jdff dff_B_DnQe1eps2_2(.din(w_dff_B_qYTGGBHQ4_2),.dout(w_dff_B_DnQe1eps2_2),.clk(gclk));
	jdff dff_B_wOc0NqTM3_2(.din(w_dff_B_DnQe1eps2_2),.dout(w_dff_B_wOc0NqTM3_2),.clk(gclk));
	jdff dff_B_l2LCdCB09_2(.din(w_dff_B_wOc0NqTM3_2),.dout(w_dff_B_l2LCdCB09_2),.clk(gclk));
	jdff dff_B_fMjO1sZz7_2(.din(w_dff_B_l2LCdCB09_2),.dout(w_dff_B_fMjO1sZz7_2),.clk(gclk));
	jdff dff_B_D2krJ9sU8_2(.din(w_dff_B_fMjO1sZz7_2),.dout(w_dff_B_D2krJ9sU8_2),.clk(gclk));
	jdff dff_B_V3Tvob7D8_2(.din(w_dff_B_D2krJ9sU8_2),.dout(w_dff_B_V3Tvob7D8_2),.clk(gclk));
	jdff dff_B_aoBNOexl5_2(.din(w_dff_B_V3Tvob7D8_2),.dout(w_dff_B_aoBNOexl5_2),.clk(gclk));
	jdff dff_B_Igy2xp7q7_2(.din(w_dff_B_aoBNOexl5_2),.dout(w_dff_B_Igy2xp7q7_2),.clk(gclk));
	jdff dff_B_fPLs186h5_2(.din(w_dff_B_Igy2xp7q7_2),.dout(w_dff_B_fPLs186h5_2),.clk(gclk));
	jdff dff_B_ooSGm1Wu3_2(.din(w_dff_B_fPLs186h5_2),.dout(w_dff_B_ooSGm1Wu3_2),.clk(gclk));
	jdff dff_B_EPIkemYa6_2(.din(w_dff_B_ooSGm1Wu3_2),.dout(w_dff_B_EPIkemYa6_2),.clk(gclk));
	jdff dff_B_0srqfk369_2(.din(w_dff_B_EPIkemYa6_2),.dout(w_dff_B_0srqfk369_2),.clk(gclk));
	jdff dff_B_mDjfZofs0_2(.din(w_dff_B_0srqfk369_2),.dout(w_dff_B_mDjfZofs0_2),.clk(gclk));
	jdff dff_B_ONRmRIjR0_2(.din(w_dff_B_mDjfZofs0_2),.dout(w_dff_B_ONRmRIjR0_2),.clk(gclk));
	jdff dff_B_Fn0cynub1_2(.din(w_dff_B_ONRmRIjR0_2),.dout(w_dff_B_Fn0cynub1_2),.clk(gclk));
	jdff dff_B_Cy1ke8qC5_2(.din(w_dff_B_Fn0cynub1_2),.dout(w_dff_B_Cy1ke8qC5_2),.clk(gclk));
	jdff dff_B_l3P9r0Z05_2(.din(w_dff_B_Cy1ke8qC5_2),.dout(w_dff_B_l3P9r0Z05_2),.clk(gclk));
	jdff dff_B_tn8Bj7vT3_2(.din(w_dff_B_l3P9r0Z05_2),.dout(w_dff_B_tn8Bj7vT3_2),.clk(gclk));
	jdff dff_B_ZZfgxB8n9_2(.din(w_dff_B_tn8Bj7vT3_2),.dout(w_dff_B_ZZfgxB8n9_2),.clk(gclk));
	jdff dff_B_inr8OxK96_2(.din(w_dff_B_ZZfgxB8n9_2),.dout(w_dff_B_inr8OxK96_2),.clk(gclk));
	jdff dff_B_zqSBWBxZ4_2(.din(w_dff_B_inr8OxK96_2),.dout(w_dff_B_zqSBWBxZ4_2),.clk(gclk));
	jdff dff_B_XdgUDHoV7_2(.din(w_dff_B_zqSBWBxZ4_2),.dout(w_dff_B_XdgUDHoV7_2),.clk(gclk));
	jdff dff_B_qLO6wcXk4_2(.din(w_dff_B_XdgUDHoV7_2),.dout(w_dff_B_qLO6wcXk4_2),.clk(gclk));
	jdff dff_B_2GUUuvJi6_2(.din(n1460),.dout(w_dff_B_2GUUuvJi6_2),.clk(gclk));
	jdff dff_B_BcUnDo3x0_2(.din(w_dff_B_2GUUuvJi6_2),.dout(w_dff_B_BcUnDo3x0_2),.clk(gclk));
	jdff dff_B_ZTUmweih7_2(.din(w_dff_B_BcUnDo3x0_2),.dout(w_dff_B_ZTUmweih7_2),.clk(gclk));
	jdff dff_B_mnxWbeaS7_2(.din(w_dff_B_ZTUmweih7_2),.dout(w_dff_B_mnxWbeaS7_2),.clk(gclk));
	jdff dff_B_mly1ZQ6m9_2(.din(w_dff_B_mnxWbeaS7_2),.dout(w_dff_B_mly1ZQ6m9_2),.clk(gclk));
	jdff dff_B_DsxJIYWN8_2(.din(w_dff_B_mly1ZQ6m9_2),.dout(w_dff_B_DsxJIYWN8_2),.clk(gclk));
	jdff dff_B_cSN5Cmro0_2(.din(w_dff_B_DsxJIYWN8_2),.dout(w_dff_B_cSN5Cmro0_2),.clk(gclk));
	jdff dff_B_CBPklAv78_2(.din(w_dff_B_cSN5Cmro0_2),.dout(w_dff_B_CBPklAv78_2),.clk(gclk));
	jdff dff_B_eYqCWvtK9_2(.din(w_dff_B_CBPklAv78_2),.dout(w_dff_B_eYqCWvtK9_2),.clk(gclk));
	jdff dff_B_JzIh3nX11_2(.din(w_dff_B_eYqCWvtK9_2),.dout(w_dff_B_JzIh3nX11_2),.clk(gclk));
	jdff dff_B_R1tHNeA23_2(.din(w_dff_B_JzIh3nX11_2),.dout(w_dff_B_R1tHNeA23_2),.clk(gclk));
	jdff dff_B_y3sOlxXo1_2(.din(w_dff_B_R1tHNeA23_2),.dout(w_dff_B_y3sOlxXo1_2),.clk(gclk));
	jdff dff_B_FQuTkHes5_2(.din(w_dff_B_y3sOlxXo1_2),.dout(w_dff_B_FQuTkHes5_2),.clk(gclk));
	jdff dff_B_hF9g4pqb5_2(.din(w_dff_B_FQuTkHes5_2),.dout(w_dff_B_hF9g4pqb5_2),.clk(gclk));
	jdff dff_B_hYx4OPiE9_2(.din(w_dff_B_hF9g4pqb5_2),.dout(w_dff_B_hYx4OPiE9_2),.clk(gclk));
	jdff dff_B_wqBGXGS29_2(.din(w_dff_B_hYx4OPiE9_2),.dout(w_dff_B_wqBGXGS29_2),.clk(gclk));
	jdff dff_B_EVUWCY8u1_2(.din(w_dff_B_wqBGXGS29_2),.dout(w_dff_B_EVUWCY8u1_2),.clk(gclk));
	jdff dff_B_AVD8uGbv5_2(.din(w_dff_B_EVUWCY8u1_2),.dout(w_dff_B_AVD8uGbv5_2),.clk(gclk));
	jdff dff_B_LZAS6Ncv7_2(.din(w_dff_B_AVD8uGbv5_2),.dout(w_dff_B_LZAS6Ncv7_2),.clk(gclk));
	jdff dff_B_9Ezn80wH8_2(.din(w_dff_B_LZAS6Ncv7_2),.dout(w_dff_B_9Ezn80wH8_2),.clk(gclk));
	jdff dff_B_drNNHBSY3_2(.din(w_dff_B_9Ezn80wH8_2),.dout(w_dff_B_drNNHBSY3_2),.clk(gclk));
	jdff dff_B_40GxfDLh2_2(.din(w_dff_B_drNNHBSY3_2),.dout(w_dff_B_40GxfDLh2_2),.clk(gclk));
	jdff dff_B_hkNq5KuS4_2(.din(w_dff_B_40GxfDLh2_2),.dout(w_dff_B_hkNq5KuS4_2),.clk(gclk));
	jdff dff_B_0jv3VXap9_2(.din(w_dff_B_hkNq5KuS4_2),.dout(w_dff_B_0jv3VXap9_2),.clk(gclk));
	jdff dff_B_cx3cJiul8_2(.din(w_dff_B_0jv3VXap9_2),.dout(w_dff_B_cx3cJiul8_2),.clk(gclk));
	jdff dff_B_9HjdEJhl7_2(.din(w_dff_B_cx3cJiul8_2),.dout(w_dff_B_9HjdEJhl7_2),.clk(gclk));
	jdff dff_B_jUVca4ae9_2(.din(n1459),.dout(w_dff_B_jUVca4ae9_2),.clk(gclk));
	jdff dff_B_QnmaqLHI3_1(.din(n1457),.dout(w_dff_B_QnmaqLHI3_1),.clk(gclk));
	jdff dff_B_RTYpZfbk8_2(.din(n1378),.dout(w_dff_B_RTYpZfbk8_2),.clk(gclk));
	jdff dff_B_1h5JXzJ86_2(.din(w_dff_B_RTYpZfbk8_2),.dout(w_dff_B_1h5JXzJ86_2),.clk(gclk));
	jdff dff_B_AcHC6nNx6_2(.din(w_dff_B_1h5JXzJ86_2),.dout(w_dff_B_AcHC6nNx6_2),.clk(gclk));
	jdff dff_B_ocXo9ELj4_2(.din(w_dff_B_AcHC6nNx6_2),.dout(w_dff_B_ocXo9ELj4_2),.clk(gclk));
	jdff dff_B_jKH6hJgT0_2(.din(w_dff_B_ocXo9ELj4_2),.dout(w_dff_B_jKH6hJgT0_2),.clk(gclk));
	jdff dff_B_ilvAowbK1_2(.din(w_dff_B_jKH6hJgT0_2),.dout(w_dff_B_ilvAowbK1_2),.clk(gclk));
	jdff dff_B_VLPeSxyM5_2(.din(w_dff_B_ilvAowbK1_2),.dout(w_dff_B_VLPeSxyM5_2),.clk(gclk));
	jdff dff_B_XU5Xcd4s4_2(.din(w_dff_B_VLPeSxyM5_2),.dout(w_dff_B_XU5Xcd4s4_2),.clk(gclk));
	jdff dff_B_B89o1cIh6_2(.din(w_dff_B_XU5Xcd4s4_2),.dout(w_dff_B_B89o1cIh6_2),.clk(gclk));
	jdff dff_B_msrWJA2I1_2(.din(w_dff_B_B89o1cIh6_2),.dout(w_dff_B_msrWJA2I1_2),.clk(gclk));
	jdff dff_B_EzqXSzlB0_2(.din(w_dff_B_msrWJA2I1_2),.dout(w_dff_B_EzqXSzlB0_2),.clk(gclk));
	jdff dff_B_GSA0RLq28_2(.din(w_dff_B_EzqXSzlB0_2),.dout(w_dff_B_GSA0RLq28_2),.clk(gclk));
	jdff dff_B_yF99YuQj5_2(.din(w_dff_B_GSA0RLq28_2),.dout(w_dff_B_yF99YuQj5_2),.clk(gclk));
	jdff dff_B_myVQmF2v8_2(.din(w_dff_B_yF99YuQj5_2),.dout(w_dff_B_myVQmF2v8_2),.clk(gclk));
	jdff dff_B_H9CCqDaM9_2(.din(w_dff_B_myVQmF2v8_2),.dout(w_dff_B_H9CCqDaM9_2),.clk(gclk));
	jdff dff_B_CITYv9zH7_2(.din(w_dff_B_H9CCqDaM9_2),.dout(w_dff_B_CITYv9zH7_2),.clk(gclk));
	jdff dff_B_IqlDVPEu7_2(.din(w_dff_B_CITYv9zH7_2),.dout(w_dff_B_IqlDVPEu7_2),.clk(gclk));
	jdff dff_B_k5spDBxP4_2(.din(w_dff_B_IqlDVPEu7_2),.dout(w_dff_B_k5spDBxP4_2),.clk(gclk));
	jdff dff_B_hGmShCwr1_2(.din(w_dff_B_k5spDBxP4_2),.dout(w_dff_B_hGmShCwr1_2),.clk(gclk));
	jdff dff_B_9OR9JLkl7_2(.din(w_dff_B_hGmShCwr1_2),.dout(w_dff_B_9OR9JLkl7_2),.clk(gclk));
	jdff dff_B_kehTNLxI5_2(.din(w_dff_B_9OR9JLkl7_2),.dout(w_dff_B_kehTNLxI5_2),.clk(gclk));
	jdff dff_B_XzFRErpm5_2(.din(w_dff_B_kehTNLxI5_2),.dout(w_dff_B_XzFRErpm5_2),.clk(gclk));
	jdff dff_B_XOoBHcnR4_2(.din(w_dff_B_XzFRErpm5_2),.dout(w_dff_B_XOoBHcnR4_2),.clk(gclk));
	jdff dff_B_5yASU09a7_1(.din(n1384),.dout(w_dff_B_5yASU09a7_1),.clk(gclk));
	jdff dff_B_OLZWrOjp4_1(.din(w_dff_B_5yASU09a7_1),.dout(w_dff_B_OLZWrOjp4_1),.clk(gclk));
	jdff dff_B_olLFN9c87_2(.din(n1383),.dout(w_dff_B_olLFN9c87_2),.clk(gclk));
	jdff dff_B_Oy1yACP37_2(.din(w_dff_B_olLFN9c87_2),.dout(w_dff_B_Oy1yACP37_2),.clk(gclk));
	jdff dff_B_hILtbE4e4_2(.din(w_dff_B_Oy1yACP37_2),.dout(w_dff_B_hILtbE4e4_2),.clk(gclk));
	jdff dff_B_jAZ0UAPM5_2(.din(w_dff_B_hILtbE4e4_2),.dout(w_dff_B_jAZ0UAPM5_2),.clk(gclk));
	jdff dff_B_tD6kzMRP0_2(.din(w_dff_B_jAZ0UAPM5_2),.dout(w_dff_B_tD6kzMRP0_2),.clk(gclk));
	jdff dff_B_9EfIgV226_2(.din(w_dff_B_tD6kzMRP0_2),.dout(w_dff_B_9EfIgV226_2),.clk(gclk));
	jdff dff_B_2sTwPaFB7_2(.din(w_dff_B_9EfIgV226_2),.dout(w_dff_B_2sTwPaFB7_2),.clk(gclk));
	jdff dff_B_LGlJ9LGR6_2(.din(w_dff_B_2sTwPaFB7_2),.dout(w_dff_B_LGlJ9LGR6_2),.clk(gclk));
	jdff dff_B_Gy1z6sy28_2(.din(w_dff_B_LGlJ9LGR6_2),.dout(w_dff_B_Gy1z6sy28_2),.clk(gclk));
	jdff dff_B_qil5CCJE2_2(.din(w_dff_B_Gy1z6sy28_2),.dout(w_dff_B_qil5CCJE2_2),.clk(gclk));
	jdff dff_B_ugPp0WhU1_2(.din(w_dff_B_qil5CCJE2_2),.dout(w_dff_B_ugPp0WhU1_2),.clk(gclk));
	jdff dff_B_fqUOMK534_2(.din(w_dff_B_ugPp0WhU1_2),.dout(w_dff_B_fqUOMK534_2),.clk(gclk));
	jdff dff_B_mhWh2Hty5_2(.din(w_dff_B_fqUOMK534_2),.dout(w_dff_B_mhWh2Hty5_2),.clk(gclk));
	jdff dff_B_v5OiShYa0_2(.din(w_dff_B_mhWh2Hty5_2),.dout(w_dff_B_v5OiShYa0_2),.clk(gclk));
	jdff dff_B_wVN5XThm4_2(.din(w_dff_B_v5OiShYa0_2),.dout(w_dff_B_wVN5XThm4_2),.clk(gclk));
	jdff dff_B_XR9ue4V19_2(.din(w_dff_B_wVN5XThm4_2),.dout(w_dff_B_XR9ue4V19_2),.clk(gclk));
	jdff dff_B_bKVQjgk65_2(.din(w_dff_B_XR9ue4V19_2),.dout(w_dff_B_bKVQjgk65_2),.clk(gclk));
	jdff dff_B_P6lI9vI11_2(.din(w_dff_B_bKVQjgk65_2),.dout(w_dff_B_P6lI9vI11_2),.clk(gclk));
	jdff dff_B_zQGYo7ns2_2(.din(w_dff_B_P6lI9vI11_2),.dout(w_dff_B_zQGYo7ns2_2),.clk(gclk));
	jdff dff_B_2TsNxkrJ7_2(.din(w_dff_B_zQGYo7ns2_2),.dout(w_dff_B_2TsNxkrJ7_2),.clk(gclk));
	jdff dff_B_u4OSFqmP6_2(.din(n1382),.dout(w_dff_B_u4OSFqmP6_2),.clk(gclk));
	jdff dff_B_nlfaaTG72_2(.din(w_dff_B_u4OSFqmP6_2),.dout(w_dff_B_nlfaaTG72_2),.clk(gclk));
	jdff dff_B_VJVzxNCg7_2(.din(w_dff_B_nlfaaTG72_2),.dout(w_dff_B_VJVzxNCg7_2),.clk(gclk));
	jdff dff_B_30SkPjq55_2(.din(w_dff_B_VJVzxNCg7_2),.dout(w_dff_B_30SkPjq55_2),.clk(gclk));
	jdff dff_B_uSQi8yFR7_2(.din(w_dff_B_30SkPjq55_2),.dout(w_dff_B_uSQi8yFR7_2),.clk(gclk));
	jdff dff_B_3Ahs3CHu0_2(.din(w_dff_B_uSQi8yFR7_2),.dout(w_dff_B_3Ahs3CHu0_2),.clk(gclk));
	jdff dff_B_1jT8OPdh5_2(.din(w_dff_B_3Ahs3CHu0_2),.dout(w_dff_B_1jT8OPdh5_2),.clk(gclk));
	jdff dff_B_5JuWZToz2_2(.din(w_dff_B_1jT8OPdh5_2),.dout(w_dff_B_5JuWZToz2_2),.clk(gclk));
	jdff dff_B_VtPQUMxf3_2(.din(w_dff_B_5JuWZToz2_2),.dout(w_dff_B_VtPQUMxf3_2),.clk(gclk));
	jdff dff_B_YH45DRSu7_2(.din(w_dff_B_VtPQUMxf3_2),.dout(w_dff_B_YH45DRSu7_2),.clk(gclk));
	jdff dff_B_4APZnBpN8_2(.din(w_dff_B_YH45DRSu7_2),.dout(w_dff_B_4APZnBpN8_2),.clk(gclk));
	jdff dff_B_c0tyCitH7_2(.din(w_dff_B_4APZnBpN8_2),.dout(w_dff_B_c0tyCitH7_2),.clk(gclk));
	jdff dff_B_b4kjQ4vj9_2(.din(w_dff_B_c0tyCitH7_2),.dout(w_dff_B_b4kjQ4vj9_2),.clk(gclk));
	jdff dff_B_GtTC14yz3_2(.din(w_dff_B_b4kjQ4vj9_2),.dout(w_dff_B_GtTC14yz3_2),.clk(gclk));
	jdff dff_B_J9YPhhVi8_2(.din(w_dff_B_GtTC14yz3_2),.dout(w_dff_B_J9YPhhVi8_2),.clk(gclk));
	jdff dff_B_ce6ZBtkp1_2(.din(w_dff_B_J9YPhhVi8_2),.dout(w_dff_B_ce6ZBtkp1_2),.clk(gclk));
	jdff dff_B_EagJwI7z3_2(.din(w_dff_B_ce6ZBtkp1_2),.dout(w_dff_B_EagJwI7z3_2),.clk(gclk));
	jdff dff_B_x5wcMjqP2_2(.din(w_dff_B_EagJwI7z3_2),.dout(w_dff_B_x5wcMjqP2_2),.clk(gclk));
	jdff dff_B_dz69GAil1_2(.din(w_dff_B_x5wcMjqP2_2),.dout(w_dff_B_dz69GAil1_2),.clk(gclk));
	jdff dff_B_USR9CEH27_2(.din(w_dff_B_dz69GAil1_2),.dout(w_dff_B_USR9CEH27_2),.clk(gclk));
	jdff dff_B_IVvOEBOt9_2(.din(w_dff_B_USR9CEH27_2),.dout(w_dff_B_IVvOEBOt9_2),.clk(gclk));
	jdff dff_B_IEOErc0A7_2(.din(w_dff_B_IVvOEBOt9_2),.dout(w_dff_B_IEOErc0A7_2),.clk(gclk));
	jdff dff_B_fYYk5f3O9_2(.din(n1381),.dout(w_dff_B_fYYk5f3O9_2),.clk(gclk));
	jdff dff_B_8PWg07E36_1(.din(n1379),.dout(w_dff_B_8PWg07E36_1),.clk(gclk));
	jdff dff_B_OzHhAVOr8_2(.din(n1293),.dout(w_dff_B_OzHhAVOr8_2),.clk(gclk));
	jdff dff_B_VKHez9Q05_2(.din(w_dff_B_OzHhAVOr8_2),.dout(w_dff_B_VKHez9Q05_2),.clk(gclk));
	jdff dff_B_wSxZEkEG6_2(.din(w_dff_B_VKHez9Q05_2),.dout(w_dff_B_wSxZEkEG6_2),.clk(gclk));
	jdff dff_B_bgpXZGrs1_2(.din(w_dff_B_wSxZEkEG6_2),.dout(w_dff_B_bgpXZGrs1_2),.clk(gclk));
	jdff dff_B_TQyk5DZu4_2(.din(w_dff_B_bgpXZGrs1_2),.dout(w_dff_B_TQyk5DZu4_2),.clk(gclk));
	jdff dff_B_iiZ26NXU0_2(.din(w_dff_B_TQyk5DZu4_2),.dout(w_dff_B_iiZ26NXU0_2),.clk(gclk));
	jdff dff_B_u3ZcPFKs5_2(.din(w_dff_B_iiZ26NXU0_2),.dout(w_dff_B_u3ZcPFKs5_2),.clk(gclk));
	jdff dff_B_NH2bHgDY3_2(.din(w_dff_B_u3ZcPFKs5_2),.dout(w_dff_B_NH2bHgDY3_2),.clk(gclk));
	jdff dff_B_KOPAkTZ98_2(.din(w_dff_B_NH2bHgDY3_2),.dout(w_dff_B_KOPAkTZ98_2),.clk(gclk));
	jdff dff_B_GJyHhEcH6_2(.din(w_dff_B_KOPAkTZ98_2),.dout(w_dff_B_GJyHhEcH6_2),.clk(gclk));
	jdff dff_B_H7y5d9bZ3_2(.din(w_dff_B_GJyHhEcH6_2),.dout(w_dff_B_H7y5d9bZ3_2),.clk(gclk));
	jdff dff_B_tslGbXB79_2(.din(w_dff_B_H7y5d9bZ3_2),.dout(w_dff_B_tslGbXB79_2),.clk(gclk));
	jdff dff_B_N1htLnBN3_2(.din(w_dff_B_tslGbXB79_2),.dout(w_dff_B_N1htLnBN3_2),.clk(gclk));
	jdff dff_B_w00JVhEH6_2(.din(w_dff_B_N1htLnBN3_2),.dout(w_dff_B_w00JVhEH6_2),.clk(gclk));
	jdff dff_B_oZbSLAm03_2(.din(w_dff_B_w00JVhEH6_2),.dout(w_dff_B_oZbSLAm03_2),.clk(gclk));
	jdff dff_B_GFeb4tGH0_2(.din(w_dff_B_oZbSLAm03_2),.dout(w_dff_B_GFeb4tGH0_2),.clk(gclk));
	jdff dff_B_2V2Ugc569_2(.din(w_dff_B_GFeb4tGH0_2),.dout(w_dff_B_2V2Ugc569_2),.clk(gclk));
	jdff dff_B_VOrXH5oj5_2(.din(w_dff_B_2V2Ugc569_2),.dout(w_dff_B_VOrXH5oj5_2),.clk(gclk));
	jdff dff_B_EGF4byLT4_2(.din(w_dff_B_VOrXH5oj5_2),.dout(w_dff_B_EGF4byLT4_2),.clk(gclk));
	jdff dff_B_Qv0e2HCL2_1(.din(n1299),.dout(w_dff_B_Qv0e2HCL2_1),.clk(gclk));
	jdff dff_B_e2ET3Y1E7_1(.din(w_dff_B_Qv0e2HCL2_1),.dout(w_dff_B_e2ET3Y1E7_1),.clk(gclk));
	jdff dff_B_Y3Dj646E0_2(.din(n1298),.dout(w_dff_B_Y3Dj646E0_2),.clk(gclk));
	jdff dff_B_7CvXI7ia0_2(.din(w_dff_B_Y3Dj646E0_2),.dout(w_dff_B_7CvXI7ia0_2),.clk(gclk));
	jdff dff_B_9xXQQOur9_2(.din(w_dff_B_7CvXI7ia0_2),.dout(w_dff_B_9xXQQOur9_2),.clk(gclk));
	jdff dff_B_7HO27aZ45_2(.din(w_dff_B_9xXQQOur9_2),.dout(w_dff_B_7HO27aZ45_2),.clk(gclk));
	jdff dff_B_jJNuFAOp9_2(.din(w_dff_B_7HO27aZ45_2),.dout(w_dff_B_jJNuFAOp9_2),.clk(gclk));
	jdff dff_B_cYqN30bH0_2(.din(w_dff_B_jJNuFAOp9_2),.dout(w_dff_B_cYqN30bH0_2),.clk(gclk));
	jdff dff_B_DlhQfQlF8_2(.din(w_dff_B_cYqN30bH0_2),.dout(w_dff_B_DlhQfQlF8_2),.clk(gclk));
	jdff dff_B_exE0wN6I5_2(.din(w_dff_B_DlhQfQlF8_2),.dout(w_dff_B_exE0wN6I5_2),.clk(gclk));
	jdff dff_B_vuCazIXF0_2(.din(w_dff_B_exE0wN6I5_2),.dout(w_dff_B_vuCazIXF0_2),.clk(gclk));
	jdff dff_B_BKjuYlam2_2(.din(w_dff_B_vuCazIXF0_2),.dout(w_dff_B_BKjuYlam2_2),.clk(gclk));
	jdff dff_B_wD24toJc9_2(.din(w_dff_B_BKjuYlam2_2),.dout(w_dff_B_wD24toJc9_2),.clk(gclk));
	jdff dff_B_MQpUhRpQ3_2(.din(w_dff_B_wD24toJc9_2),.dout(w_dff_B_MQpUhRpQ3_2),.clk(gclk));
	jdff dff_B_ziTNQ1Cx2_2(.din(w_dff_B_MQpUhRpQ3_2),.dout(w_dff_B_ziTNQ1Cx2_2),.clk(gclk));
	jdff dff_B_RkkV6wiZ3_2(.din(w_dff_B_ziTNQ1Cx2_2),.dout(w_dff_B_RkkV6wiZ3_2),.clk(gclk));
	jdff dff_B_AxdOm1kF0_2(.din(w_dff_B_RkkV6wiZ3_2),.dout(w_dff_B_AxdOm1kF0_2),.clk(gclk));
	jdff dff_B_7a6jpQSa0_2(.din(w_dff_B_AxdOm1kF0_2),.dout(w_dff_B_7a6jpQSa0_2),.clk(gclk));
	jdff dff_B_LFO4qeg28_2(.din(n1297),.dout(w_dff_B_LFO4qeg28_2),.clk(gclk));
	jdff dff_B_Mw2zSURz3_2(.din(w_dff_B_LFO4qeg28_2),.dout(w_dff_B_Mw2zSURz3_2),.clk(gclk));
	jdff dff_B_BlHRHpQm6_2(.din(w_dff_B_Mw2zSURz3_2),.dout(w_dff_B_BlHRHpQm6_2),.clk(gclk));
	jdff dff_B_g23d2ye54_2(.din(w_dff_B_BlHRHpQm6_2),.dout(w_dff_B_g23d2ye54_2),.clk(gclk));
	jdff dff_B_HslQ4LMC2_2(.din(w_dff_B_g23d2ye54_2),.dout(w_dff_B_HslQ4LMC2_2),.clk(gclk));
	jdff dff_B_qFEL7Ce34_2(.din(w_dff_B_HslQ4LMC2_2),.dout(w_dff_B_qFEL7Ce34_2),.clk(gclk));
	jdff dff_B_NfJh0SOk3_2(.din(w_dff_B_qFEL7Ce34_2),.dout(w_dff_B_NfJh0SOk3_2),.clk(gclk));
	jdff dff_B_0kdqCHKs6_2(.din(w_dff_B_NfJh0SOk3_2),.dout(w_dff_B_0kdqCHKs6_2),.clk(gclk));
	jdff dff_B_RCXf0GSK9_2(.din(w_dff_B_0kdqCHKs6_2),.dout(w_dff_B_RCXf0GSK9_2),.clk(gclk));
	jdff dff_B_SbeIj4EA9_2(.din(w_dff_B_RCXf0GSK9_2),.dout(w_dff_B_SbeIj4EA9_2),.clk(gclk));
	jdff dff_B_oWCisUL88_2(.din(w_dff_B_SbeIj4EA9_2),.dout(w_dff_B_oWCisUL88_2),.clk(gclk));
	jdff dff_B_73KwR9kl1_2(.din(w_dff_B_oWCisUL88_2),.dout(w_dff_B_73KwR9kl1_2),.clk(gclk));
	jdff dff_B_Ws0GHVFN2_2(.din(w_dff_B_73KwR9kl1_2),.dout(w_dff_B_Ws0GHVFN2_2),.clk(gclk));
	jdff dff_B_MSt4HiVG0_2(.din(w_dff_B_Ws0GHVFN2_2),.dout(w_dff_B_MSt4HiVG0_2),.clk(gclk));
	jdff dff_B_yZAGZScQ3_2(.din(w_dff_B_MSt4HiVG0_2),.dout(w_dff_B_yZAGZScQ3_2),.clk(gclk));
	jdff dff_B_pM6Mmx3n7_2(.din(w_dff_B_yZAGZScQ3_2),.dout(w_dff_B_pM6Mmx3n7_2),.clk(gclk));
	jdff dff_B_IjKhdoj22_2(.din(w_dff_B_pM6Mmx3n7_2),.dout(w_dff_B_IjKhdoj22_2),.clk(gclk));
	jdff dff_B_HNwucoHX8_2(.din(w_dff_B_IjKhdoj22_2),.dout(w_dff_B_HNwucoHX8_2),.clk(gclk));
	jdff dff_B_MWaXlhv09_2(.din(n1296),.dout(w_dff_B_MWaXlhv09_2),.clk(gclk));
	jdff dff_B_DZrKGAMs6_1(.din(n1294),.dout(w_dff_B_DZrKGAMs6_1),.clk(gclk));
	jdff dff_B_szCQqSSU2_2(.din(n1203),.dout(w_dff_B_szCQqSSU2_2),.clk(gclk));
	jdff dff_B_lOEFlTU39_2(.din(w_dff_B_szCQqSSU2_2),.dout(w_dff_B_lOEFlTU39_2),.clk(gclk));
	jdff dff_B_Jqv4AdE23_2(.din(w_dff_B_lOEFlTU39_2),.dout(w_dff_B_Jqv4AdE23_2),.clk(gclk));
	jdff dff_B_XiAMtTEU2_2(.din(w_dff_B_Jqv4AdE23_2),.dout(w_dff_B_XiAMtTEU2_2),.clk(gclk));
	jdff dff_B_cbUdpB1v5_2(.din(w_dff_B_XiAMtTEU2_2),.dout(w_dff_B_cbUdpB1v5_2),.clk(gclk));
	jdff dff_B_EZjbtMY64_2(.din(w_dff_B_cbUdpB1v5_2),.dout(w_dff_B_EZjbtMY64_2),.clk(gclk));
	jdff dff_B_kCVwGTK17_2(.din(w_dff_B_EZjbtMY64_2),.dout(w_dff_B_kCVwGTK17_2),.clk(gclk));
	jdff dff_B_IM5IdGkX5_2(.din(w_dff_B_kCVwGTK17_2),.dout(w_dff_B_IM5IdGkX5_2),.clk(gclk));
	jdff dff_B_EWB7lJfj3_2(.din(w_dff_B_IM5IdGkX5_2),.dout(w_dff_B_EWB7lJfj3_2),.clk(gclk));
	jdff dff_B_y4KSNL9q6_2(.din(w_dff_B_EWB7lJfj3_2),.dout(w_dff_B_y4KSNL9q6_2),.clk(gclk));
	jdff dff_B_BruesTkW2_2(.din(w_dff_B_y4KSNL9q6_2),.dout(w_dff_B_BruesTkW2_2),.clk(gclk));
	jdff dff_B_pgFTnIOK6_2(.din(w_dff_B_BruesTkW2_2),.dout(w_dff_B_pgFTnIOK6_2),.clk(gclk));
	jdff dff_B_xVlEOmrX7_2(.din(w_dff_B_pgFTnIOK6_2),.dout(w_dff_B_xVlEOmrX7_2),.clk(gclk));
	jdff dff_B_6J2NyFim8_2(.din(w_dff_B_xVlEOmrX7_2),.dout(w_dff_B_6J2NyFim8_2),.clk(gclk));
	jdff dff_B_B9IrkPD37_2(.din(w_dff_B_6J2NyFim8_2),.dout(w_dff_B_B9IrkPD37_2),.clk(gclk));
	jdff dff_B_RntvHVY90_2(.din(n1208),.dout(w_dff_B_RntvHVY90_2),.clk(gclk));
	jdff dff_B_fG3DPFL78_2(.din(w_dff_B_RntvHVY90_2),.dout(w_dff_B_fG3DPFL78_2),.clk(gclk));
	jdff dff_B_utpFtmHA2_2(.din(w_dff_B_fG3DPFL78_2),.dout(w_dff_B_utpFtmHA2_2),.clk(gclk));
	jdff dff_B_NT2Q9DQR8_2(.din(w_dff_B_utpFtmHA2_2),.dout(w_dff_B_NT2Q9DQR8_2),.clk(gclk));
	jdff dff_B_0q3OCYoI2_2(.din(w_dff_B_NT2Q9DQR8_2),.dout(w_dff_B_0q3OCYoI2_2),.clk(gclk));
	jdff dff_B_v2k9uez14_2(.din(w_dff_B_0q3OCYoI2_2),.dout(w_dff_B_v2k9uez14_2),.clk(gclk));
	jdff dff_B_5AdnHcnK5_2(.din(w_dff_B_v2k9uez14_2),.dout(w_dff_B_5AdnHcnK5_2),.clk(gclk));
	jdff dff_B_QqvYuJ5h8_2(.din(w_dff_B_5AdnHcnK5_2),.dout(w_dff_B_QqvYuJ5h8_2),.clk(gclk));
	jdff dff_B_T2Q7Wbqm2_2(.din(w_dff_B_QqvYuJ5h8_2),.dout(w_dff_B_T2Q7Wbqm2_2),.clk(gclk));
	jdff dff_B_mES2Qmt23_2(.din(w_dff_B_T2Q7Wbqm2_2),.dout(w_dff_B_mES2Qmt23_2),.clk(gclk));
	jdff dff_B_fxYnfF0S9_2(.din(w_dff_B_mES2Qmt23_2),.dout(w_dff_B_fxYnfF0S9_2),.clk(gclk));
	jdff dff_B_RqiMIXOz0_2(.din(w_dff_B_fxYnfF0S9_2),.dout(w_dff_B_RqiMIXOz0_2),.clk(gclk));
	jdff dff_B_wTSyRGBe8_2(.din(n1207),.dout(w_dff_B_wTSyRGBe8_2),.clk(gclk));
	jdff dff_B_R7U1seq15_2(.din(w_dff_B_wTSyRGBe8_2),.dout(w_dff_B_R7U1seq15_2),.clk(gclk));
	jdff dff_B_Cnh3ALpc1_2(.din(w_dff_B_R7U1seq15_2),.dout(w_dff_B_Cnh3ALpc1_2),.clk(gclk));
	jdff dff_B_wAlqMFZK2_2(.din(w_dff_B_Cnh3ALpc1_2),.dout(w_dff_B_wAlqMFZK2_2),.clk(gclk));
	jdff dff_B_YmJ0rA5v8_2(.din(w_dff_B_wAlqMFZK2_2),.dout(w_dff_B_YmJ0rA5v8_2),.clk(gclk));
	jdff dff_B_EqXigxnl2_2(.din(w_dff_B_YmJ0rA5v8_2),.dout(w_dff_B_EqXigxnl2_2),.clk(gclk));
	jdff dff_B_qEd7GUfv1_2(.din(w_dff_B_EqXigxnl2_2),.dout(w_dff_B_qEd7GUfv1_2),.clk(gclk));
	jdff dff_B_USPE4sBL7_2(.din(w_dff_B_qEd7GUfv1_2),.dout(w_dff_B_USPE4sBL7_2),.clk(gclk));
	jdff dff_B_9s7J8j272_2(.din(w_dff_B_USPE4sBL7_2),.dout(w_dff_B_9s7J8j272_2),.clk(gclk));
	jdff dff_B_MW0mOvnW2_2(.din(w_dff_B_9s7J8j272_2),.dout(w_dff_B_MW0mOvnW2_2),.clk(gclk));
	jdff dff_B_uHG8XFyv3_2(.din(w_dff_B_MW0mOvnW2_2),.dout(w_dff_B_uHG8XFyv3_2),.clk(gclk));
	jdff dff_B_VSTZy9ar0_2(.din(w_dff_B_uHG8XFyv3_2),.dout(w_dff_B_VSTZy9ar0_2),.clk(gclk));
	jdff dff_B_5pvmsgAx2_2(.din(w_dff_B_VSTZy9ar0_2),.dout(w_dff_B_5pvmsgAx2_2),.clk(gclk));
	jdff dff_B_y5rNK1No5_2(.din(w_dff_B_5pvmsgAx2_2),.dout(w_dff_B_y5rNK1No5_2),.clk(gclk));
	jdff dff_B_ZnJx9fZ55_2(.din(n1206),.dout(w_dff_B_ZnJx9fZ55_2),.clk(gclk));
	jdff dff_B_ekLgpStc5_1(.din(n1204),.dout(w_dff_B_ekLgpStc5_1),.clk(gclk));
	jdff dff_B_bStYKeD78_2(.din(n1099),.dout(w_dff_B_bStYKeD78_2),.clk(gclk));
	jdff dff_B_tcQEwGcI6_2(.din(w_dff_B_bStYKeD78_2),.dout(w_dff_B_tcQEwGcI6_2),.clk(gclk));
	jdff dff_B_HzGCXw0e3_2(.din(w_dff_B_tcQEwGcI6_2),.dout(w_dff_B_HzGCXw0e3_2),.clk(gclk));
	jdff dff_B_o0zYhiyG4_2(.din(w_dff_B_HzGCXw0e3_2),.dout(w_dff_B_o0zYhiyG4_2),.clk(gclk));
	jdff dff_B_TI8ZuKjZ5_2(.din(w_dff_B_o0zYhiyG4_2),.dout(w_dff_B_TI8ZuKjZ5_2),.clk(gclk));
	jdff dff_B_TpDxDOgf3_2(.din(w_dff_B_TI8ZuKjZ5_2),.dout(w_dff_B_TpDxDOgf3_2),.clk(gclk));
	jdff dff_B_gXurmGlr9_2(.din(w_dff_B_TpDxDOgf3_2),.dout(w_dff_B_gXurmGlr9_2),.clk(gclk));
	jdff dff_B_7IOOwjVc4_2(.din(w_dff_B_gXurmGlr9_2),.dout(w_dff_B_7IOOwjVc4_2),.clk(gclk));
	jdff dff_B_R5OmwPa20_2(.din(w_dff_B_7IOOwjVc4_2),.dout(w_dff_B_R5OmwPa20_2),.clk(gclk));
	jdff dff_B_lIu6VCdA5_2(.din(w_dff_B_R5OmwPa20_2),.dout(w_dff_B_lIu6VCdA5_2),.clk(gclk));
	jdff dff_B_9lWhhvuT2_2(.din(w_dff_B_lIu6VCdA5_2),.dout(w_dff_B_9lWhhvuT2_2),.clk(gclk));
	jdff dff_A_Ajg6pi0s7_0(.dout(w_n1110_0[0]),.din(w_dff_A_Ajg6pi0s7_0),.clk(gclk));
	jdff dff_A_AKZFsUKo0_0(.dout(w_dff_A_Ajg6pi0s7_0),.din(w_dff_A_AKZFsUKo0_0),.clk(gclk));
	jdff dff_A_f2e2Ey2h5_0(.dout(w_dff_A_AKZFsUKo0_0),.din(w_dff_A_f2e2Ey2h5_0),.clk(gclk));
	jdff dff_B_GDoq4Fl55_2(.din(n1110),.dout(w_dff_B_GDoq4Fl55_2),.clk(gclk));
	jdff dff_B_35JBD6cT9_1(.din(n1104),.dout(w_dff_B_35JBD6cT9_1),.clk(gclk));
	jdff dff_B_mznpII4E5_1(.din(w_dff_B_35JBD6cT9_1),.dout(w_dff_B_mznpII4E5_1),.clk(gclk));
	jdff dff_B_vwTQ4LEh0_1(.din(w_dff_B_mznpII4E5_1),.dout(w_dff_B_vwTQ4LEh0_1),.clk(gclk));
	jdff dff_B_tLoMFTzR5_1(.din(w_dff_B_vwTQ4LEh0_1),.dout(w_dff_B_tLoMFTzR5_1),.clk(gclk));
	jdff dff_B_pfb2HwpJ1_1(.din(w_dff_B_tLoMFTzR5_1),.dout(w_dff_B_pfb2HwpJ1_1),.clk(gclk));
	jdff dff_B_B5JNyJST3_1(.din(w_dff_B_pfb2HwpJ1_1),.dout(w_dff_B_B5JNyJST3_1),.clk(gclk));
	jdff dff_B_PQHk8nW76_1(.din(n1105),.dout(w_dff_B_PQHk8nW76_1),.clk(gclk));
	jdff dff_B_IWVdypPc3_1(.din(w_dff_B_PQHk8nW76_1),.dout(w_dff_B_IWVdypPc3_1),.clk(gclk));
	jdff dff_A_TZ6tGNyO8_1(.dout(w_G307gat_2[1]),.din(w_dff_A_TZ6tGNyO8_1),.clk(gclk));
	jdff dff_A_4xiO9KTf8_1(.dout(w_dff_A_TZ6tGNyO8_1),.din(w_dff_A_4xiO9KTf8_1),.clk(gclk));
	jdff dff_A_m2JdDYnS7_1(.dout(w_dff_A_4xiO9KTf8_1),.din(w_dff_A_m2JdDYnS7_1),.clk(gclk));
	jdff dff_A_XdPmzeat0_1(.dout(w_dff_A_m2JdDYnS7_1),.din(w_dff_A_XdPmzeat0_1),.clk(gclk));
	jdff dff_A_vhJuOkKT5_1(.dout(w_dff_A_XdPmzeat0_1),.din(w_dff_A_vhJuOkKT5_1),.clk(gclk));
	jdff dff_A_xXmrnfsi0_1(.dout(w_dff_A_vhJuOkKT5_1),.din(w_dff_A_xXmrnfsi0_1),.clk(gclk));
	jdff dff_A_TGokZRHD9_1(.dout(w_dff_A_xXmrnfsi0_1),.din(w_dff_A_TGokZRHD9_1),.clk(gclk));
	jdff dff_B_RmMAyjat2_2(.din(n1103),.dout(w_dff_B_RmMAyjat2_2),.clk(gclk));
	jdff dff_B_39TboRSy1_2(.din(w_dff_B_RmMAyjat2_2),.dout(w_dff_B_39TboRSy1_2),.clk(gclk));
	jdff dff_B_Ch6Yixrm2_2(.din(w_dff_B_39TboRSy1_2),.dout(w_dff_B_Ch6Yixrm2_2),.clk(gclk));
	jdff dff_B_gZ8hmKrM8_2(.din(w_dff_B_Ch6Yixrm2_2),.dout(w_dff_B_gZ8hmKrM8_2),.clk(gclk));
	jdff dff_B_YNY4Uvzw2_2(.din(w_dff_B_gZ8hmKrM8_2),.dout(w_dff_B_YNY4Uvzw2_2),.clk(gclk));
	jdff dff_B_1yeDeOyg8_2(.din(w_dff_B_YNY4Uvzw2_2),.dout(w_dff_B_1yeDeOyg8_2),.clk(gclk));
	jdff dff_B_dq8Y05WN7_2(.din(w_dff_B_1yeDeOyg8_2),.dout(w_dff_B_dq8Y05WN7_2),.clk(gclk));
	jdff dff_B_UC6AoPgJ6_2(.din(w_dff_B_dq8Y05WN7_2),.dout(w_dff_B_UC6AoPgJ6_2),.clk(gclk));
	jdff dff_B_pKyIMzVa8_2(.din(w_dff_B_UC6AoPgJ6_2),.dout(w_dff_B_pKyIMzVa8_2),.clk(gclk));
	jdff dff_B_cqFfBWP55_2(.din(w_dff_B_pKyIMzVa8_2),.dout(w_dff_B_cqFfBWP55_2),.clk(gclk));
	jdff dff_B_cmfpmCl56_1(.din(n1100),.dout(w_dff_B_cmfpmCl56_1),.clk(gclk));
	jdff dff_B_X1hBfCeL4_2(.din(n1001),.dout(w_dff_B_X1hBfCeL4_2),.clk(gclk));
	jdff dff_B_UfPsd2bc2_2(.din(w_dff_B_X1hBfCeL4_2),.dout(w_dff_B_UfPsd2bc2_2),.clk(gclk));
	jdff dff_B_yV00sn1Q7_2(.din(w_dff_B_UfPsd2bc2_2),.dout(w_dff_B_yV00sn1Q7_2),.clk(gclk));
	jdff dff_B_y9DjVUcg0_2(.din(w_dff_B_yV00sn1Q7_2),.dout(w_dff_B_y9DjVUcg0_2),.clk(gclk));
	jdff dff_B_jWFSNWq73_2(.din(w_dff_B_y9DjVUcg0_2),.dout(w_dff_B_jWFSNWq73_2),.clk(gclk));
	jdff dff_B_JD0A8qP97_2(.din(w_dff_B_jWFSNWq73_2),.dout(w_dff_B_JD0A8qP97_2),.clk(gclk));
	jdff dff_B_snnwlZP56_2(.din(w_dff_B_JD0A8qP97_2),.dout(w_dff_B_snnwlZP56_2),.clk(gclk));
	jdff dff_B_rvbvWtr08_2(.din(w_dff_B_snnwlZP56_2),.dout(w_dff_B_rvbvWtr08_2),.clk(gclk));
	jdff dff_B_aMxbGL8a2_2(.din(n1010),.dout(w_dff_B_aMxbGL8a2_2),.clk(gclk));
	jdff dff_B_WbleH03o3_2(.din(w_dff_B_aMxbGL8a2_2),.dout(w_dff_B_WbleH03o3_2),.clk(gclk));
	jdff dff_B_m1RCkkPH9_2(.din(w_dff_B_WbleH03o3_2),.dout(w_dff_B_m1RCkkPH9_2),.clk(gclk));
	jdff dff_B_Wp4tjeBe1_2(.din(w_dff_B_m1RCkkPH9_2),.dout(w_dff_B_Wp4tjeBe1_2),.clk(gclk));
	jdff dff_B_rbubUt2i7_2(.din(w_dff_B_Wp4tjeBe1_2),.dout(w_dff_B_rbubUt2i7_2),.clk(gclk));
	jdff dff_A_U1HcrelJ0_0(.dout(w_n1008_0[0]),.din(w_dff_A_U1HcrelJ0_0),.clk(gclk));
	jdff dff_A_2ggyHQ8U6_0(.dout(w_dff_A_U1HcrelJ0_0),.din(w_dff_A_2ggyHQ8U6_0),.clk(gclk));
	jdff dff_A_vaNofmMD7_0(.dout(w_dff_A_2ggyHQ8U6_0),.din(w_dff_A_vaNofmMD7_0),.clk(gclk));
	jdff dff_A_uVjBeraU8_0(.dout(w_n793_0[0]),.din(w_dff_A_uVjBeraU8_0),.clk(gclk));
	jdff dff_A_B5pqTIi46_1(.dout(w_n1006_0[1]),.din(w_dff_A_B5pqTIi46_1),.clk(gclk));
	jdff dff_A_DIA0lUDf8_1(.dout(w_dff_A_B5pqTIi46_1),.din(w_dff_A_DIA0lUDf8_1),.clk(gclk));
	jdff dff_B_5oDqQnFC4_1(.din(n1002),.dout(w_dff_B_5oDqQnFC4_1),.clk(gclk));
	jdff dff_B_KZLhzZXj0_1(.din(w_dff_B_5oDqQnFC4_1),.dout(w_dff_B_KZLhzZXj0_1),.clk(gclk));
	jdff dff_B_YmpiVlK80_1(.din(w_dff_B_KZLhzZXj0_1),.dout(w_dff_B_YmpiVlK80_1),.clk(gclk));
	jdff dff_B_bvM5pOaO1_1(.din(w_dff_B_YmpiVlK80_1),.dout(w_dff_B_bvM5pOaO1_1),.clk(gclk));
	jdff dff_B_7ocKJlph9_1(.din(w_dff_B_bvM5pOaO1_1),.dout(w_dff_B_7ocKJlph9_1),.clk(gclk));
	jdff dff_A_3tzYqdid4_0(.dout(w_n903_0[0]),.din(w_dff_A_3tzYqdid4_0),.clk(gclk));
	jdff dff_A_iPbA4AM20_0(.dout(w_dff_A_3tzYqdid4_0),.din(w_dff_A_iPbA4AM20_0),.clk(gclk));
	jdff dff_A_uLByc2El7_0(.dout(w_dff_A_iPbA4AM20_0),.din(w_dff_A_uLByc2El7_0),.clk(gclk));
	jdff dff_A_f2OUeufa5_0(.dout(w_n695_0[0]),.din(w_dff_A_f2OUeufa5_0),.clk(gclk));
	jdff dff_A_0kBr7MwZ8_0(.dout(w_dff_A_f2OUeufa5_0),.din(w_dff_A_0kBr7MwZ8_0),.clk(gclk));
	jdff dff_A_VCHMQp1s7_0(.dout(w_dff_A_0kBr7MwZ8_0),.din(w_dff_A_VCHMQp1s7_0),.clk(gclk));
	jdff dff_B_lLac3uo07_2(.din(n898),.dout(w_dff_B_lLac3uo07_2),.clk(gclk));
	jdff dff_A_HlqjyqD42_1(.dout(w_n896_0[1]),.din(w_dff_A_HlqjyqD42_1),.clk(gclk));
	jdff dff_A_z9GPjSto8_1(.dout(w_dff_A_HlqjyqD42_1),.din(w_dff_A_z9GPjSto8_1),.clk(gclk));
	jdff dff_A_PqR25d2d6_1(.dout(w_dff_A_z9GPjSto8_1),.din(w_dff_A_PqR25d2d6_1),.clk(gclk));
	jdff dff_A_LFZNbteQ8_1(.dout(w_dff_A_PqR25d2d6_1),.din(w_dff_A_LFZNbteQ8_1),.clk(gclk));
	jdff dff_A_AhwbHvEf1_1(.dout(w_dff_A_LFZNbteQ8_1),.din(w_dff_A_AhwbHvEf1_1),.clk(gclk));
	jdff dff_A_rE4qmGgL3_1(.dout(w_dff_A_ZHjSjUI17_0),.din(w_dff_A_rE4qmGgL3_1),.clk(gclk));
	jdff dff_A_ZHjSjUI17_0(.dout(w_dff_A_a5FiIX6v2_0),.din(w_dff_A_ZHjSjUI17_0),.clk(gclk));
	jdff dff_A_a5FiIX6v2_0(.dout(w_dff_A_GjJySaNj3_0),.din(w_dff_A_a5FiIX6v2_0),.clk(gclk));
	jdff dff_A_GjJySaNj3_0(.dout(w_dff_A_qNBEAGXc1_0),.din(w_dff_A_GjJySaNj3_0),.clk(gclk));
	jdff dff_A_qNBEAGXc1_0(.dout(w_dff_A_BU4rTDgm3_0),.din(w_dff_A_qNBEAGXc1_0),.clk(gclk));
	jdff dff_A_BU4rTDgm3_0(.dout(w_dff_A_fGX7JfCv5_0),.din(w_dff_A_BU4rTDgm3_0),.clk(gclk));
	jdff dff_A_fGX7JfCv5_0(.dout(w_dff_A_pr6bOVe40_0),.din(w_dff_A_fGX7JfCv5_0),.clk(gclk));
	jdff dff_A_pr6bOVe40_0(.dout(w_dff_A_fE7kvKyq3_0),.din(w_dff_A_pr6bOVe40_0),.clk(gclk));
	jdff dff_A_fE7kvKyq3_0(.dout(w_dff_A_44kvQYtZ7_0),.din(w_dff_A_fE7kvKyq3_0),.clk(gclk));
	jdff dff_A_44kvQYtZ7_0(.dout(w_dff_A_Qu8OTBtf4_0),.din(w_dff_A_44kvQYtZ7_0),.clk(gclk));
	jdff dff_A_Qu8OTBtf4_0(.dout(w_dff_A_A30gUBkh9_0),.din(w_dff_A_Qu8OTBtf4_0),.clk(gclk));
	jdff dff_A_A30gUBkh9_0(.dout(w_dff_A_sGgHrYJb0_0),.din(w_dff_A_A30gUBkh9_0),.clk(gclk));
	jdff dff_A_sGgHrYJb0_0(.dout(w_dff_A_AlYXZySL1_0),.din(w_dff_A_sGgHrYJb0_0),.clk(gclk));
	jdff dff_A_AlYXZySL1_0(.dout(w_dff_A_7eGlORmV1_0),.din(w_dff_A_AlYXZySL1_0),.clk(gclk));
	jdff dff_A_7eGlORmV1_0(.dout(w_dff_A_4IMo6afp9_0),.din(w_dff_A_7eGlORmV1_0),.clk(gclk));
	jdff dff_A_4IMo6afp9_0(.dout(w_dff_A_9l1niQwx9_0),.din(w_dff_A_4IMo6afp9_0),.clk(gclk));
	jdff dff_A_9l1niQwx9_0(.dout(w_dff_A_77ogvPP86_0),.din(w_dff_A_9l1niQwx9_0),.clk(gclk));
	jdff dff_A_77ogvPP86_0(.dout(w_dff_A_BHSr3EmJ0_0),.din(w_dff_A_77ogvPP86_0),.clk(gclk));
	jdff dff_A_BHSr3EmJ0_0(.dout(w_dff_A_bjAgsrpW0_0),.din(w_dff_A_BHSr3EmJ0_0),.clk(gclk));
	jdff dff_A_bjAgsrpW0_0(.dout(w_dff_A_NrivGG2h2_0),.din(w_dff_A_bjAgsrpW0_0),.clk(gclk));
	jdff dff_A_NrivGG2h2_0(.dout(w_dff_A_XYj3p9UF8_0),.din(w_dff_A_NrivGG2h2_0),.clk(gclk));
	jdff dff_A_XYj3p9UF8_0(.dout(w_dff_A_J9yBLkpz7_0),.din(w_dff_A_XYj3p9UF8_0),.clk(gclk));
	jdff dff_A_J9yBLkpz7_0(.dout(w_dff_A_itn12WyD8_0),.din(w_dff_A_J9yBLkpz7_0),.clk(gclk));
	jdff dff_A_itn12WyD8_0(.dout(w_dff_A_xu7skIGf8_0),.din(w_dff_A_itn12WyD8_0),.clk(gclk));
	jdff dff_A_xu7skIGf8_0(.dout(w_dff_A_JcuAN9sZ9_0),.din(w_dff_A_xu7skIGf8_0),.clk(gclk));
	jdff dff_A_JcuAN9sZ9_0(.dout(w_dff_A_UqtOzkKK3_0),.din(w_dff_A_JcuAN9sZ9_0),.clk(gclk));
	jdff dff_A_UqtOzkKK3_0(.dout(w_dff_A_KdfBZQGv4_0),.din(w_dff_A_UqtOzkKK3_0),.clk(gclk));
	jdff dff_A_KdfBZQGv4_0(.dout(w_dff_A_6YgT5HmA5_0),.din(w_dff_A_KdfBZQGv4_0),.clk(gclk));
	jdff dff_A_6YgT5HmA5_0(.dout(w_dff_A_1TftoEOW8_0),.din(w_dff_A_6YgT5HmA5_0),.clk(gclk));
	jdff dff_A_1TftoEOW8_0(.dout(w_dff_A_USQYQHf75_0),.din(w_dff_A_1TftoEOW8_0),.clk(gclk));
	jdff dff_A_USQYQHf75_0(.dout(w_dff_A_1D1Y6BUd5_0),.din(w_dff_A_USQYQHf75_0),.clk(gclk));
	jdff dff_A_1D1Y6BUd5_0(.dout(w_dff_A_AGJH553l7_0),.din(w_dff_A_1D1Y6BUd5_0),.clk(gclk));
	jdff dff_A_AGJH553l7_0(.dout(w_dff_A_hwq5kgka2_0),.din(w_dff_A_AGJH553l7_0),.clk(gclk));
	jdff dff_A_hwq5kgka2_0(.dout(w_dff_A_YN4nNPtx9_0),.din(w_dff_A_hwq5kgka2_0),.clk(gclk));
	jdff dff_A_YN4nNPtx9_0(.dout(w_dff_A_mtZguglp8_0),.din(w_dff_A_YN4nNPtx9_0),.clk(gclk));
	jdff dff_A_mtZguglp8_0(.dout(w_dff_A_yJGhVhhl3_0),.din(w_dff_A_mtZguglp8_0),.clk(gclk));
	jdff dff_A_yJGhVhhl3_0(.dout(w_dff_A_548WKCsg9_0),.din(w_dff_A_yJGhVhhl3_0),.clk(gclk));
	jdff dff_A_548WKCsg9_0(.dout(w_dff_A_mLPPM5sn6_0),.din(w_dff_A_548WKCsg9_0),.clk(gclk));
	jdff dff_A_mLPPM5sn6_0(.dout(w_dff_A_nrufeGX17_0),.din(w_dff_A_mLPPM5sn6_0),.clk(gclk));
	jdff dff_A_nrufeGX17_0(.dout(w_dff_A_4MqFCvoH0_0),.din(w_dff_A_nrufeGX17_0),.clk(gclk));
	jdff dff_A_4MqFCvoH0_0(.dout(w_dff_A_2zk8f1AU5_0),.din(w_dff_A_4MqFCvoH0_0),.clk(gclk));
	jdff dff_A_2zk8f1AU5_0(.dout(w_dff_A_AguR2ECu4_0),.din(w_dff_A_2zk8f1AU5_0),.clk(gclk));
	jdff dff_A_AguR2ECu4_0(.dout(w_dff_A_ny7PYMA96_0),.din(w_dff_A_AguR2ECu4_0),.clk(gclk));
	jdff dff_A_ny7PYMA96_0(.dout(w_dff_A_98ErYpfl4_0),.din(w_dff_A_ny7PYMA96_0),.clk(gclk));
	jdff dff_A_98ErYpfl4_0(.dout(w_dff_A_qce9Ezw64_0),.din(w_dff_A_98ErYpfl4_0),.clk(gclk));
	jdff dff_A_qce9Ezw64_0(.dout(w_dff_A_LvmED0907_0),.din(w_dff_A_qce9Ezw64_0),.clk(gclk));
	jdff dff_A_LvmED0907_0(.dout(w_dff_A_ZrwPCZx36_0),.din(w_dff_A_LvmED0907_0),.clk(gclk));
	jdff dff_A_ZrwPCZx36_0(.dout(w_dff_A_6Fb6qF1p2_0),.din(w_dff_A_ZrwPCZx36_0),.clk(gclk));
	jdff dff_A_6Fb6qF1p2_0(.dout(w_dff_A_TTH40hc38_0),.din(w_dff_A_6Fb6qF1p2_0),.clk(gclk));
	jdff dff_A_TTH40hc38_0(.dout(w_dff_A_8qhQPsyN2_0),.din(w_dff_A_TTH40hc38_0),.clk(gclk));
	jdff dff_A_8qhQPsyN2_0(.dout(w_dff_A_slabGQfO5_0),.din(w_dff_A_8qhQPsyN2_0),.clk(gclk));
	jdff dff_A_slabGQfO5_0(.dout(w_dff_A_lEDkFNI38_0),.din(w_dff_A_slabGQfO5_0),.clk(gclk));
	jdff dff_A_lEDkFNI38_0(.dout(w_dff_A_iYmAUuzm0_0),.din(w_dff_A_lEDkFNI38_0),.clk(gclk));
	jdff dff_A_iYmAUuzm0_0(.dout(w_dff_A_OlYLz6wX1_0),.din(w_dff_A_iYmAUuzm0_0),.clk(gclk));
	jdff dff_A_OlYLz6wX1_0(.dout(w_dff_A_dALT4q3n8_0),.din(w_dff_A_OlYLz6wX1_0),.clk(gclk));
	jdff dff_A_dALT4q3n8_0(.dout(w_dff_A_CgyGOVCN8_0),.din(w_dff_A_dALT4q3n8_0),.clk(gclk));
	jdff dff_A_CgyGOVCN8_0(.dout(w_dff_A_5gfEFDge0_0),.din(w_dff_A_CgyGOVCN8_0),.clk(gclk));
	jdff dff_A_5gfEFDge0_0(.dout(w_dff_A_s78YTkNL7_0),.din(w_dff_A_5gfEFDge0_0),.clk(gclk));
	jdff dff_A_s78YTkNL7_0(.dout(w_dff_A_kPG8ZVs28_0),.din(w_dff_A_s78YTkNL7_0),.clk(gclk));
	jdff dff_A_kPG8ZVs28_0(.dout(w_dff_A_WAUmUw6U6_0),.din(w_dff_A_kPG8ZVs28_0),.clk(gclk));
	jdff dff_A_WAUmUw6U6_0(.dout(w_dff_A_NPgZlsW65_0),.din(w_dff_A_WAUmUw6U6_0),.clk(gclk));
	jdff dff_A_NPgZlsW65_0(.dout(w_dff_A_jOaAEEDT2_0),.din(w_dff_A_NPgZlsW65_0),.clk(gclk));
	jdff dff_A_jOaAEEDT2_0(.dout(w_dff_A_PWbMRYmD2_0),.din(w_dff_A_jOaAEEDT2_0),.clk(gclk));
	jdff dff_A_PWbMRYmD2_0(.dout(w_dff_A_LM1FenCm6_0),.din(w_dff_A_PWbMRYmD2_0),.clk(gclk));
	jdff dff_A_LM1FenCm6_0(.dout(w_dff_A_qHIUtCQv8_0),.din(w_dff_A_LM1FenCm6_0),.clk(gclk));
	jdff dff_A_qHIUtCQv8_0(.dout(w_dff_A_NTuBIZC16_0),.din(w_dff_A_qHIUtCQv8_0),.clk(gclk));
	jdff dff_A_NTuBIZC16_0(.dout(w_dff_A_irNDFiMt4_0),.din(w_dff_A_NTuBIZC16_0),.clk(gclk));
	jdff dff_A_irNDFiMt4_0(.dout(w_dff_A_P4linBrj6_0),.din(w_dff_A_irNDFiMt4_0),.clk(gclk));
	jdff dff_A_P4linBrj6_0(.dout(w_dff_A_Giinq9195_0),.din(w_dff_A_P4linBrj6_0),.clk(gclk));
	jdff dff_A_Giinq9195_0(.dout(w_dff_A_cYf0crjQ1_0),.din(w_dff_A_Giinq9195_0),.clk(gclk));
	jdff dff_A_cYf0crjQ1_0(.dout(w_dff_A_VBKTxnU93_0),.din(w_dff_A_cYf0crjQ1_0),.clk(gclk));
	jdff dff_A_VBKTxnU93_0(.dout(w_dff_A_aumP3CjT5_0),.din(w_dff_A_VBKTxnU93_0),.clk(gclk));
	jdff dff_A_aumP3CjT5_0(.dout(w_dff_A_98G6dCIX3_0),.din(w_dff_A_aumP3CjT5_0),.clk(gclk));
	jdff dff_A_98G6dCIX3_0(.dout(w_dff_A_P7Rt7lic5_0),.din(w_dff_A_98G6dCIX3_0),.clk(gclk));
	jdff dff_A_P7Rt7lic5_0(.dout(G545gat),.din(w_dff_A_P7Rt7lic5_0),.clk(gclk));
	jdff dff_A_YXiv6Yx23_2(.dout(w_dff_A_p64RLqHA6_0),.din(w_dff_A_YXiv6Yx23_2),.clk(gclk));
	jdff dff_A_p64RLqHA6_0(.dout(w_dff_A_Kc8P7odh1_0),.din(w_dff_A_p64RLqHA6_0),.clk(gclk));
	jdff dff_A_Kc8P7odh1_0(.dout(w_dff_A_SjmfjdMv9_0),.din(w_dff_A_Kc8P7odh1_0),.clk(gclk));
	jdff dff_A_SjmfjdMv9_0(.dout(w_dff_A_5RDbOpvM5_0),.din(w_dff_A_SjmfjdMv9_0),.clk(gclk));
	jdff dff_A_5RDbOpvM5_0(.dout(w_dff_A_peI4Grcg6_0),.din(w_dff_A_5RDbOpvM5_0),.clk(gclk));
	jdff dff_A_peI4Grcg6_0(.dout(w_dff_A_or75KAGO6_0),.din(w_dff_A_peI4Grcg6_0),.clk(gclk));
	jdff dff_A_or75KAGO6_0(.dout(w_dff_A_wGvRFbvr5_0),.din(w_dff_A_or75KAGO6_0),.clk(gclk));
	jdff dff_A_wGvRFbvr5_0(.dout(w_dff_A_8B23OrgM6_0),.din(w_dff_A_wGvRFbvr5_0),.clk(gclk));
	jdff dff_A_8B23OrgM6_0(.dout(w_dff_A_H3ssAJR90_0),.din(w_dff_A_8B23OrgM6_0),.clk(gclk));
	jdff dff_A_H3ssAJR90_0(.dout(w_dff_A_fzAJolga8_0),.din(w_dff_A_H3ssAJR90_0),.clk(gclk));
	jdff dff_A_fzAJolga8_0(.dout(w_dff_A_jDtwgd2i4_0),.din(w_dff_A_fzAJolga8_0),.clk(gclk));
	jdff dff_A_jDtwgd2i4_0(.dout(w_dff_A_W2yE3rvl0_0),.din(w_dff_A_jDtwgd2i4_0),.clk(gclk));
	jdff dff_A_W2yE3rvl0_0(.dout(w_dff_A_PFsb8Yf51_0),.din(w_dff_A_W2yE3rvl0_0),.clk(gclk));
	jdff dff_A_PFsb8Yf51_0(.dout(w_dff_A_p7puu2no7_0),.din(w_dff_A_PFsb8Yf51_0),.clk(gclk));
	jdff dff_A_p7puu2no7_0(.dout(w_dff_A_vfDdvrFO3_0),.din(w_dff_A_p7puu2no7_0),.clk(gclk));
	jdff dff_A_vfDdvrFO3_0(.dout(w_dff_A_TTeC5tV14_0),.din(w_dff_A_vfDdvrFO3_0),.clk(gclk));
	jdff dff_A_TTeC5tV14_0(.dout(w_dff_A_jzfbyS4I7_0),.din(w_dff_A_TTeC5tV14_0),.clk(gclk));
	jdff dff_A_jzfbyS4I7_0(.dout(w_dff_A_i9vzbcfc5_0),.din(w_dff_A_jzfbyS4I7_0),.clk(gclk));
	jdff dff_A_i9vzbcfc5_0(.dout(w_dff_A_ktjbljTE0_0),.din(w_dff_A_i9vzbcfc5_0),.clk(gclk));
	jdff dff_A_ktjbljTE0_0(.dout(w_dff_A_LVV36kZL1_0),.din(w_dff_A_ktjbljTE0_0),.clk(gclk));
	jdff dff_A_LVV36kZL1_0(.dout(w_dff_A_6CjaYoLO1_0),.din(w_dff_A_LVV36kZL1_0),.clk(gclk));
	jdff dff_A_6CjaYoLO1_0(.dout(w_dff_A_HxOUhU9n0_0),.din(w_dff_A_6CjaYoLO1_0),.clk(gclk));
	jdff dff_A_HxOUhU9n0_0(.dout(w_dff_A_By7SmI832_0),.din(w_dff_A_HxOUhU9n0_0),.clk(gclk));
	jdff dff_A_By7SmI832_0(.dout(w_dff_A_zxKvatpL2_0),.din(w_dff_A_By7SmI832_0),.clk(gclk));
	jdff dff_A_zxKvatpL2_0(.dout(w_dff_A_5ameRFIA4_0),.din(w_dff_A_zxKvatpL2_0),.clk(gclk));
	jdff dff_A_5ameRFIA4_0(.dout(w_dff_A_YcFPflsI3_0),.din(w_dff_A_5ameRFIA4_0),.clk(gclk));
	jdff dff_A_YcFPflsI3_0(.dout(w_dff_A_FKECd3dk6_0),.din(w_dff_A_YcFPflsI3_0),.clk(gclk));
	jdff dff_A_FKECd3dk6_0(.dout(w_dff_A_FOjuWzTf0_0),.din(w_dff_A_FKECd3dk6_0),.clk(gclk));
	jdff dff_A_FOjuWzTf0_0(.dout(w_dff_A_OMTNsVM81_0),.din(w_dff_A_FOjuWzTf0_0),.clk(gclk));
	jdff dff_A_OMTNsVM81_0(.dout(w_dff_A_JkSPIyLB4_0),.din(w_dff_A_OMTNsVM81_0),.clk(gclk));
	jdff dff_A_JkSPIyLB4_0(.dout(w_dff_A_merzZsE68_0),.din(w_dff_A_JkSPIyLB4_0),.clk(gclk));
	jdff dff_A_merzZsE68_0(.dout(w_dff_A_cdYbLOH19_0),.din(w_dff_A_merzZsE68_0),.clk(gclk));
	jdff dff_A_cdYbLOH19_0(.dout(w_dff_A_JGeJVqJn3_0),.din(w_dff_A_cdYbLOH19_0),.clk(gclk));
	jdff dff_A_JGeJVqJn3_0(.dout(w_dff_A_S0FYVG1S0_0),.din(w_dff_A_JGeJVqJn3_0),.clk(gclk));
	jdff dff_A_S0FYVG1S0_0(.dout(w_dff_A_xgRwYFbb3_0),.din(w_dff_A_S0FYVG1S0_0),.clk(gclk));
	jdff dff_A_xgRwYFbb3_0(.dout(w_dff_A_8yiAk4tD8_0),.din(w_dff_A_xgRwYFbb3_0),.clk(gclk));
	jdff dff_A_8yiAk4tD8_0(.dout(w_dff_A_kpXii2qt5_0),.din(w_dff_A_8yiAk4tD8_0),.clk(gclk));
	jdff dff_A_kpXii2qt5_0(.dout(w_dff_A_kpY6t2RW1_0),.din(w_dff_A_kpXii2qt5_0),.clk(gclk));
	jdff dff_A_kpY6t2RW1_0(.dout(w_dff_A_LFJqh0xF9_0),.din(w_dff_A_kpY6t2RW1_0),.clk(gclk));
	jdff dff_A_LFJqh0xF9_0(.dout(w_dff_A_Ct3URjSe1_0),.din(w_dff_A_LFJqh0xF9_0),.clk(gclk));
	jdff dff_A_Ct3URjSe1_0(.dout(w_dff_A_LpTzvMRc1_0),.din(w_dff_A_Ct3URjSe1_0),.clk(gclk));
	jdff dff_A_LpTzvMRc1_0(.dout(w_dff_A_agohsC0X8_0),.din(w_dff_A_LpTzvMRc1_0),.clk(gclk));
	jdff dff_A_agohsC0X8_0(.dout(w_dff_A_05f6D0SG2_0),.din(w_dff_A_agohsC0X8_0),.clk(gclk));
	jdff dff_A_05f6D0SG2_0(.dout(w_dff_A_MHH2uqGI2_0),.din(w_dff_A_05f6D0SG2_0),.clk(gclk));
	jdff dff_A_MHH2uqGI2_0(.dout(w_dff_A_M8fUQQ3i5_0),.din(w_dff_A_MHH2uqGI2_0),.clk(gclk));
	jdff dff_A_M8fUQQ3i5_0(.dout(w_dff_A_SF7FExQW6_0),.din(w_dff_A_M8fUQQ3i5_0),.clk(gclk));
	jdff dff_A_SF7FExQW6_0(.dout(w_dff_A_khpJA9Vz3_0),.din(w_dff_A_SF7FExQW6_0),.clk(gclk));
	jdff dff_A_khpJA9Vz3_0(.dout(w_dff_A_N8OZYB3v1_0),.din(w_dff_A_khpJA9Vz3_0),.clk(gclk));
	jdff dff_A_N8OZYB3v1_0(.dout(w_dff_A_7G07MALF0_0),.din(w_dff_A_N8OZYB3v1_0),.clk(gclk));
	jdff dff_A_7G07MALF0_0(.dout(w_dff_A_MXdsDW6I3_0),.din(w_dff_A_7G07MALF0_0),.clk(gclk));
	jdff dff_A_MXdsDW6I3_0(.dout(w_dff_A_1CBWRDSR3_0),.din(w_dff_A_MXdsDW6I3_0),.clk(gclk));
	jdff dff_A_1CBWRDSR3_0(.dout(w_dff_A_YerZPohO3_0),.din(w_dff_A_1CBWRDSR3_0),.clk(gclk));
	jdff dff_A_YerZPohO3_0(.dout(w_dff_A_BhZ3RtV71_0),.din(w_dff_A_YerZPohO3_0),.clk(gclk));
	jdff dff_A_BhZ3RtV71_0(.dout(w_dff_A_rY2wFcGx5_0),.din(w_dff_A_BhZ3RtV71_0),.clk(gclk));
	jdff dff_A_rY2wFcGx5_0(.dout(w_dff_A_NxZsVi9t8_0),.din(w_dff_A_rY2wFcGx5_0),.clk(gclk));
	jdff dff_A_NxZsVi9t8_0(.dout(w_dff_A_7ZVKcPhK8_0),.din(w_dff_A_NxZsVi9t8_0),.clk(gclk));
	jdff dff_A_7ZVKcPhK8_0(.dout(w_dff_A_U4GUl6kQ8_0),.din(w_dff_A_7ZVKcPhK8_0),.clk(gclk));
	jdff dff_A_U4GUl6kQ8_0(.dout(w_dff_A_D1V1DfQ07_0),.din(w_dff_A_U4GUl6kQ8_0),.clk(gclk));
	jdff dff_A_D1V1DfQ07_0(.dout(w_dff_A_35XEmrYb4_0),.din(w_dff_A_D1V1DfQ07_0),.clk(gclk));
	jdff dff_A_35XEmrYb4_0(.dout(w_dff_A_RhiqKDrt0_0),.din(w_dff_A_35XEmrYb4_0),.clk(gclk));
	jdff dff_A_RhiqKDrt0_0(.dout(w_dff_A_Ulr0o6TO5_0),.din(w_dff_A_RhiqKDrt0_0),.clk(gclk));
	jdff dff_A_Ulr0o6TO5_0(.dout(w_dff_A_aligU5lK9_0),.din(w_dff_A_Ulr0o6TO5_0),.clk(gclk));
	jdff dff_A_aligU5lK9_0(.dout(w_dff_A_FAYZJtDj5_0),.din(w_dff_A_aligU5lK9_0),.clk(gclk));
	jdff dff_A_FAYZJtDj5_0(.dout(w_dff_A_JWJAKf7Q0_0),.din(w_dff_A_FAYZJtDj5_0),.clk(gclk));
	jdff dff_A_JWJAKf7Q0_0(.dout(w_dff_A_KseXWj2U4_0),.din(w_dff_A_JWJAKf7Q0_0),.clk(gclk));
	jdff dff_A_KseXWj2U4_0(.dout(w_dff_A_TQU6YDac1_0),.din(w_dff_A_KseXWj2U4_0),.clk(gclk));
	jdff dff_A_TQU6YDac1_0(.dout(w_dff_A_BvEGz6x93_0),.din(w_dff_A_TQU6YDac1_0),.clk(gclk));
	jdff dff_A_BvEGz6x93_0(.dout(w_dff_A_UpFK9dU44_0),.din(w_dff_A_BvEGz6x93_0),.clk(gclk));
	jdff dff_A_UpFK9dU44_0(.dout(w_dff_A_2Yd292y00_0),.din(w_dff_A_UpFK9dU44_0),.clk(gclk));
	jdff dff_A_2Yd292y00_0(.dout(w_dff_A_NoShJDYn0_0),.din(w_dff_A_2Yd292y00_0),.clk(gclk));
	jdff dff_A_NoShJDYn0_0(.dout(w_dff_A_7LlMToQR5_0),.din(w_dff_A_NoShJDYn0_0),.clk(gclk));
	jdff dff_A_7LlMToQR5_0(.dout(G1581gat),.din(w_dff_A_7LlMToQR5_0),.clk(gclk));
	jdff dff_A_bk66JIRc7_2(.dout(w_dff_A_IKCfQeGD9_0),.din(w_dff_A_bk66JIRc7_2),.clk(gclk));
	jdff dff_A_IKCfQeGD9_0(.dout(w_dff_A_lC3t4jek6_0),.din(w_dff_A_IKCfQeGD9_0),.clk(gclk));
	jdff dff_A_lC3t4jek6_0(.dout(w_dff_A_n57bBGQP3_0),.din(w_dff_A_lC3t4jek6_0),.clk(gclk));
	jdff dff_A_n57bBGQP3_0(.dout(w_dff_A_Dpyr2gKH1_0),.din(w_dff_A_n57bBGQP3_0),.clk(gclk));
	jdff dff_A_Dpyr2gKH1_0(.dout(w_dff_A_o8HRGzKQ7_0),.din(w_dff_A_Dpyr2gKH1_0),.clk(gclk));
	jdff dff_A_o8HRGzKQ7_0(.dout(w_dff_A_V99KVqkz2_0),.din(w_dff_A_o8HRGzKQ7_0),.clk(gclk));
	jdff dff_A_V99KVqkz2_0(.dout(w_dff_A_teGtxT7P7_0),.din(w_dff_A_V99KVqkz2_0),.clk(gclk));
	jdff dff_A_teGtxT7P7_0(.dout(w_dff_A_ee17YuJ77_0),.din(w_dff_A_teGtxT7P7_0),.clk(gclk));
	jdff dff_A_ee17YuJ77_0(.dout(w_dff_A_16J9Ltb47_0),.din(w_dff_A_ee17YuJ77_0),.clk(gclk));
	jdff dff_A_16J9Ltb47_0(.dout(w_dff_A_itTsayCO6_0),.din(w_dff_A_16J9Ltb47_0),.clk(gclk));
	jdff dff_A_itTsayCO6_0(.dout(w_dff_A_1ScT891b9_0),.din(w_dff_A_itTsayCO6_0),.clk(gclk));
	jdff dff_A_1ScT891b9_0(.dout(w_dff_A_fiuBGqNA6_0),.din(w_dff_A_1ScT891b9_0),.clk(gclk));
	jdff dff_A_fiuBGqNA6_0(.dout(w_dff_A_J5JYw0Cg9_0),.din(w_dff_A_fiuBGqNA6_0),.clk(gclk));
	jdff dff_A_J5JYw0Cg9_0(.dout(w_dff_A_n6lkNNPd0_0),.din(w_dff_A_J5JYw0Cg9_0),.clk(gclk));
	jdff dff_A_n6lkNNPd0_0(.dout(w_dff_A_GjzVWqgl2_0),.din(w_dff_A_n6lkNNPd0_0),.clk(gclk));
	jdff dff_A_GjzVWqgl2_0(.dout(w_dff_A_OsT9bsmP2_0),.din(w_dff_A_GjzVWqgl2_0),.clk(gclk));
	jdff dff_A_OsT9bsmP2_0(.dout(w_dff_A_IsUssCpU0_0),.din(w_dff_A_OsT9bsmP2_0),.clk(gclk));
	jdff dff_A_IsUssCpU0_0(.dout(w_dff_A_LZmai8il1_0),.din(w_dff_A_IsUssCpU0_0),.clk(gclk));
	jdff dff_A_LZmai8il1_0(.dout(w_dff_A_X0r76xsS0_0),.din(w_dff_A_LZmai8il1_0),.clk(gclk));
	jdff dff_A_X0r76xsS0_0(.dout(w_dff_A_R6ur1G3R4_0),.din(w_dff_A_X0r76xsS0_0),.clk(gclk));
	jdff dff_A_R6ur1G3R4_0(.dout(w_dff_A_WSus9DQn2_0),.din(w_dff_A_R6ur1G3R4_0),.clk(gclk));
	jdff dff_A_WSus9DQn2_0(.dout(w_dff_A_ue27BoMK0_0),.din(w_dff_A_WSus9DQn2_0),.clk(gclk));
	jdff dff_A_ue27BoMK0_0(.dout(w_dff_A_B5EsmqgE8_0),.din(w_dff_A_ue27BoMK0_0),.clk(gclk));
	jdff dff_A_B5EsmqgE8_0(.dout(w_dff_A_tPS7lwTn4_0),.din(w_dff_A_B5EsmqgE8_0),.clk(gclk));
	jdff dff_A_tPS7lwTn4_0(.dout(w_dff_A_sxyqDQwb0_0),.din(w_dff_A_tPS7lwTn4_0),.clk(gclk));
	jdff dff_A_sxyqDQwb0_0(.dout(w_dff_A_fJDhVgOz5_0),.din(w_dff_A_sxyqDQwb0_0),.clk(gclk));
	jdff dff_A_fJDhVgOz5_0(.dout(w_dff_A_Gox6RqJK1_0),.din(w_dff_A_fJDhVgOz5_0),.clk(gclk));
	jdff dff_A_Gox6RqJK1_0(.dout(w_dff_A_yWfJCSsM6_0),.din(w_dff_A_Gox6RqJK1_0),.clk(gclk));
	jdff dff_A_yWfJCSsM6_0(.dout(w_dff_A_npB4fh242_0),.din(w_dff_A_yWfJCSsM6_0),.clk(gclk));
	jdff dff_A_npB4fh242_0(.dout(w_dff_A_ZJOgWIsk0_0),.din(w_dff_A_npB4fh242_0),.clk(gclk));
	jdff dff_A_ZJOgWIsk0_0(.dout(w_dff_A_cdoOIn1i1_0),.din(w_dff_A_ZJOgWIsk0_0),.clk(gclk));
	jdff dff_A_cdoOIn1i1_0(.dout(w_dff_A_cpQj61Q11_0),.din(w_dff_A_cdoOIn1i1_0),.clk(gclk));
	jdff dff_A_cpQj61Q11_0(.dout(w_dff_A_8u57dXdM6_0),.din(w_dff_A_cpQj61Q11_0),.clk(gclk));
	jdff dff_A_8u57dXdM6_0(.dout(w_dff_A_m6TfIlGV0_0),.din(w_dff_A_8u57dXdM6_0),.clk(gclk));
	jdff dff_A_m6TfIlGV0_0(.dout(w_dff_A_YfxDWxVz7_0),.din(w_dff_A_m6TfIlGV0_0),.clk(gclk));
	jdff dff_A_YfxDWxVz7_0(.dout(w_dff_A_0iddeGKK0_0),.din(w_dff_A_YfxDWxVz7_0),.clk(gclk));
	jdff dff_A_0iddeGKK0_0(.dout(w_dff_A_rfogrGqH8_0),.din(w_dff_A_0iddeGKK0_0),.clk(gclk));
	jdff dff_A_rfogrGqH8_0(.dout(w_dff_A_DWnq424u4_0),.din(w_dff_A_rfogrGqH8_0),.clk(gclk));
	jdff dff_A_DWnq424u4_0(.dout(w_dff_A_qLjqvj5B3_0),.din(w_dff_A_DWnq424u4_0),.clk(gclk));
	jdff dff_A_qLjqvj5B3_0(.dout(w_dff_A_RYFMtx8M8_0),.din(w_dff_A_qLjqvj5B3_0),.clk(gclk));
	jdff dff_A_RYFMtx8M8_0(.dout(w_dff_A_9rqH1VZm4_0),.din(w_dff_A_RYFMtx8M8_0),.clk(gclk));
	jdff dff_A_9rqH1VZm4_0(.dout(w_dff_A_wNigYBvw4_0),.din(w_dff_A_9rqH1VZm4_0),.clk(gclk));
	jdff dff_A_wNigYBvw4_0(.dout(w_dff_A_tR05fWiy5_0),.din(w_dff_A_wNigYBvw4_0),.clk(gclk));
	jdff dff_A_tR05fWiy5_0(.dout(w_dff_A_Ia2f72Ci3_0),.din(w_dff_A_tR05fWiy5_0),.clk(gclk));
	jdff dff_A_Ia2f72Ci3_0(.dout(w_dff_A_Yqpxj6UB9_0),.din(w_dff_A_Ia2f72Ci3_0),.clk(gclk));
	jdff dff_A_Yqpxj6UB9_0(.dout(w_dff_A_K11Uetar0_0),.din(w_dff_A_Yqpxj6UB9_0),.clk(gclk));
	jdff dff_A_K11Uetar0_0(.dout(w_dff_A_pIIYnlCH7_0),.din(w_dff_A_K11Uetar0_0),.clk(gclk));
	jdff dff_A_pIIYnlCH7_0(.dout(w_dff_A_P5yrAl677_0),.din(w_dff_A_pIIYnlCH7_0),.clk(gclk));
	jdff dff_A_P5yrAl677_0(.dout(w_dff_A_ATBUR3tj3_0),.din(w_dff_A_P5yrAl677_0),.clk(gclk));
	jdff dff_A_ATBUR3tj3_0(.dout(w_dff_A_nD9hgrCF5_0),.din(w_dff_A_ATBUR3tj3_0),.clk(gclk));
	jdff dff_A_nD9hgrCF5_0(.dout(w_dff_A_NTln6Xsz8_0),.din(w_dff_A_nD9hgrCF5_0),.clk(gclk));
	jdff dff_A_NTln6Xsz8_0(.dout(w_dff_A_G2CKQlSS9_0),.din(w_dff_A_NTln6Xsz8_0),.clk(gclk));
	jdff dff_A_G2CKQlSS9_0(.dout(w_dff_A_qqjCttYu8_0),.din(w_dff_A_G2CKQlSS9_0),.clk(gclk));
	jdff dff_A_qqjCttYu8_0(.dout(w_dff_A_8eNjoxBn4_0),.din(w_dff_A_qqjCttYu8_0),.clk(gclk));
	jdff dff_A_8eNjoxBn4_0(.dout(w_dff_A_JFGtlC5t4_0),.din(w_dff_A_8eNjoxBn4_0),.clk(gclk));
	jdff dff_A_JFGtlC5t4_0(.dout(w_dff_A_KgoDcpQ35_0),.din(w_dff_A_JFGtlC5t4_0),.clk(gclk));
	jdff dff_A_KgoDcpQ35_0(.dout(w_dff_A_zVR9oK5w1_0),.din(w_dff_A_KgoDcpQ35_0),.clk(gclk));
	jdff dff_A_zVR9oK5w1_0(.dout(w_dff_A_mBg5cCz30_0),.din(w_dff_A_zVR9oK5w1_0),.clk(gclk));
	jdff dff_A_mBg5cCz30_0(.dout(w_dff_A_wCUZ1sVW6_0),.din(w_dff_A_mBg5cCz30_0),.clk(gclk));
	jdff dff_A_wCUZ1sVW6_0(.dout(w_dff_A_rYcqg5M32_0),.din(w_dff_A_wCUZ1sVW6_0),.clk(gclk));
	jdff dff_A_rYcqg5M32_0(.dout(w_dff_A_KGNYuGTP1_0),.din(w_dff_A_rYcqg5M32_0),.clk(gclk));
	jdff dff_A_KGNYuGTP1_0(.dout(w_dff_A_1AMb7ab21_0),.din(w_dff_A_KGNYuGTP1_0),.clk(gclk));
	jdff dff_A_1AMb7ab21_0(.dout(w_dff_A_1yl3Tr0K0_0),.din(w_dff_A_1AMb7ab21_0),.clk(gclk));
	jdff dff_A_1yl3Tr0K0_0(.dout(w_dff_A_MYeHyNuP9_0),.din(w_dff_A_1yl3Tr0K0_0),.clk(gclk));
	jdff dff_A_MYeHyNuP9_0(.dout(w_dff_A_dA0i9buk1_0),.din(w_dff_A_MYeHyNuP9_0),.clk(gclk));
	jdff dff_A_dA0i9buk1_0(.dout(w_dff_A_UwY88ub12_0),.din(w_dff_A_dA0i9buk1_0),.clk(gclk));
	jdff dff_A_UwY88ub12_0(.dout(w_dff_A_QOUpQTe75_0),.din(w_dff_A_UwY88ub12_0),.clk(gclk));
	jdff dff_A_QOUpQTe75_0(.dout(w_dff_A_ZO8vVKK11_0),.din(w_dff_A_QOUpQTe75_0),.clk(gclk));
	jdff dff_A_ZO8vVKK11_0(.dout(G1901gat),.din(w_dff_A_ZO8vVKK11_0),.clk(gclk));
	jdff dff_A_ihkYZoXx2_2(.dout(w_dff_A_SC53etb39_0),.din(w_dff_A_ihkYZoXx2_2),.clk(gclk));
	jdff dff_A_SC53etb39_0(.dout(w_dff_A_GTMw07LJ7_0),.din(w_dff_A_SC53etb39_0),.clk(gclk));
	jdff dff_A_GTMw07LJ7_0(.dout(w_dff_A_abpLbixo1_0),.din(w_dff_A_GTMw07LJ7_0),.clk(gclk));
	jdff dff_A_abpLbixo1_0(.dout(w_dff_A_g6MFUHP52_0),.din(w_dff_A_abpLbixo1_0),.clk(gclk));
	jdff dff_A_g6MFUHP52_0(.dout(w_dff_A_dIuFx3vT5_0),.din(w_dff_A_g6MFUHP52_0),.clk(gclk));
	jdff dff_A_dIuFx3vT5_0(.dout(w_dff_A_mwkUC4UP9_0),.din(w_dff_A_dIuFx3vT5_0),.clk(gclk));
	jdff dff_A_mwkUC4UP9_0(.dout(w_dff_A_dVLD3Ro47_0),.din(w_dff_A_mwkUC4UP9_0),.clk(gclk));
	jdff dff_A_dVLD3Ro47_0(.dout(w_dff_A_kWQRDeEs6_0),.din(w_dff_A_dVLD3Ro47_0),.clk(gclk));
	jdff dff_A_kWQRDeEs6_0(.dout(w_dff_A_C5iXU3DY6_0),.din(w_dff_A_kWQRDeEs6_0),.clk(gclk));
	jdff dff_A_C5iXU3DY6_0(.dout(w_dff_A_P9xwoMHP3_0),.din(w_dff_A_C5iXU3DY6_0),.clk(gclk));
	jdff dff_A_P9xwoMHP3_0(.dout(w_dff_A_188WxzeC5_0),.din(w_dff_A_P9xwoMHP3_0),.clk(gclk));
	jdff dff_A_188WxzeC5_0(.dout(w_dff_A_c37TLJfK1_0),.din(w_dff_A_188WxzeC5_0),.clk(gclk));
	jdff dff_A_c37TLJfK1_0(.dout(w_dff_A_l58SNuKq3_0),.din(w_dff_A_c37TLJfK1_0),.clk(gclk));
	jdff dff_A_l58SNuKq3_0(.dout(w_dff_A_guS0juLC7_0),.din(w_dff_A_l58SNuKq3_0),.clk(gclk));
	jdff dff_A_guS0juLC7_0(.dout(w_dff_A_kAcV4oxf0_0),.din(w_dff_A_guS0juLC7_0),.clk(gclk));
	jdff dff_A_kAcV4oxf0_0(.dout(w_dff_A_ZIiaFsVb2_0),.din(w_dff_A_kAcV4oxf0_0),.clk(gclk));
	jdff dff_A_ZIiaFsVb2_0(.dout(w_dff_A_wHt4zteD1_0),.din(w_dff_A_ZIiaFsVb2_0),.clk(gclk));
	jdff dff_A_wHt4zteD1_0(.dout(w_dff_A_DHMaLv0r3_0),.din(w_dff_A_wHt4zteD1_0),.clk(gclk));
	jdff dff_A_DHMaLv0r3_0(.dout(w_dff_A_xzotiHdE6_0),.din(w_dff_A_DHMaLv0r3_0),.clk(gclk));
	jdff dff_A_xzotiHdE6_0(.dout(w_dff_A_OJlLLM5O7_0),.din(w_dff_A_xzotiHdE6_0),.clk(gclk));
	jdff dff_A_OJlLLM5O7_0(.dout(w_dff_A_Yg4WvvCX9_0),.din(w_dff_A_OJlLLM5O7_0),.clk(gclk));
	jdff dff_A_Yg4WvvCX9_0(.dout(w_dff_A_gYj8Sm3I7_0),.din(w_dff_A_Yg4WvvCX9_0),.clk(gclk));
	jdff dff_A_gYj8Sm3I7_0(.dout(w_dff_A_Gi9v8lA62_0),.din(w_dff_A_gYj8Sm3I7_0),.clk(gclk));
	jdff dff_A_Gi9v8lA62_0(.dout(w_dff_A_DSpPYdNM5_0),.din(w_dff_A_Gi9v8lA62_0),.clk(gclk));
	jdff dff_A_DSpPYdNM5_0(.dout(w_dff_A_xly4i3pr4_0),.din(w_dff_A_DSpPYdNM5_0),.clk(gclk));
	jdff dff_A_xly4i3pr4_0(.dout(w_dff_A_lBDkvRUu2_0),.din(w_dff_A_xly4i3pr4_0),.clk(gclk));
	jdff dff_A_lBDkvRUu2_0(.dout(w_dff_A_zQgRC7OG7_0),.din(w_dff_A_lBDkvRUu2_0),.clk(gclk));
	jdff dff_A_zQgRC7OG7_0(.dout(w_dff_A_2QpKr6gk8_0),.din(w_dff_A_zQgRC7OG7_0),.clk(gclk));
	jdff dff_A_2QpKr6gk8_0(.dout(w_dff_A_yZmlUCb06_0),.din(w_dff_A_2QpKr6gk8_0),.clk(gclk));
	jdff dff_A_yZmlUCb06_0(.dout(w_dff_A_ozZXWHbn6_0),.din(w_dff_A_yZmlUCb06_0),.clk(gclk));
	jdff dff_A_ozZXWHbn6_0(.dout(w_dff_A_TglgS7hl8_0),.din(w_dff_A_ozZXWHbn6_0),.clk(gclk));
	jdff dff_A_TglgS7hl8_0(.dout(w_dff_A_E6nEfCKl2_0),.din(w_dff_A_TglgS7hl8_0),.clk(gclk));
	jdff dff_A_E6nEfCKl2_0(.dout(w_dff_A_WvDEKKvF0_0),.din(w_dff_A_E6nEfCKl2_0),.clk(gclk));
	jdff dff_A_WvDEKKvF0_0(.dout(w_dff_A_NhVoXUf70_0),.din(w_dff_A_WvDEKKvF0_0),.clk(gclk));
	jdff dff_A_NhVoXUf70_0(.dout(w_dff_A_Tjw3eYba6_0),.din(w_dff_A_NhVoXUf70_0),.clk(gclk));
	jdff dff_A_Tjw3eYba6_0(.dout(w_dff_A_Df4bkLAL2_0),.din(w_dff_A_Tjw3eYba6_0),.clk(gclk));
	jdff dff_A_Df4bkLAL2_0(.dout(w_dff_A_GwQLWlZ29_0),.din(w_dff_A_Df4bkLAL2_0),.clk(gclk));
	jdff dff_A_GwQLWlZ29_0(.dout(w_dff_A_kJPi2ieZ8_0),.din(w_dff_A_GwQLWlZ29_0),.clk(gclk));
	jdff dff_A_kJPi2ieZ8_0(.dout(w_dff_A_6kIevxMP0_0),.din(w_dff_A_kJPi2ieZ8_0),.clk(gclk));
	jdff dff_A_6kIevxMP0_0(.dout(w_dff_A_yJZO6A449_0),.din(w_dff_A_6kIevxMP0_0),.clk(gclk));
	jdff dff_A_yJZO6A449_0(.dout(w_dff_A_IXbyTuFa5_0),.din(w_dff_A_yJZO6A449_0),.clk(gclk));
	jdff dff_A_IXbyTuFa5_0(.dout(w_dff_A_q8X3NXYg4_0),.din(w_dff_A_IXbyTuFa5_0),.clk(gclk));
	jdff dff_A_q8X3NXYg4_0(.dout(w_dff_A_CuZuBnGt2_0),.din(w_dff_A_q8X3NXYg4_0),.clk(gclk));
	jdff dff_A_CuZuBnGt2_0(.dout(w_dff_A_aUujZGe54_0),.din(w_dff_A_CuZuBnGt2_0),.clk(gclk));
	jdff dff_A_aUujZGe54_0(.dout(w_dff_A_Q9mGDfoZ7_0),.din(w_dff_A_aUujZGe54_0),.clk(gclk));
	jdff dff_A_Q9mGDfoZ7_0(.dout(w_dff_A_EOe5qfW22_0),.din(w_dff_A_Q9mGDfoZ7_0),.clk(gclk));
	jdff dff_A_EOe5qfW22_0(.dout(w_dff_A_FslfGcvR1_0),.din(w_dff_A_EOe5qfW22_0),.clk(gclk));
	jdff dff_A_FslfGcvR1_0(.dout(w_dff_A_fUn8xO5C3_0),.din(w_dff_A_FslfGcvR1_0),.clk(gclk));
	jdff dff_A_fUn8xO5C3_0(.dout(w_dff_A_lJ3FDdwu0_0),.din(w_dff_A_fUn8xO5C3_0),.clk(gclk));
	jdff dff_A_lJ3FDdwu0_0(.dout(w_dff_A_KHvpRFUN1_0),.din(w_dff_A_lJ3FDdwu0_0),.clk(gclk));
	jdff dff_A_KHvpRFUN1_0(.dout(w_dff_A_hVdqspZl2_0),.din(w_dff_A_KHvpRFUN1_0),.clk(gclk));
	jdff dff_A_hVdqspZl2_0(.dout(w_dff_A_u1mu6W740_0),.din(w_dff_A_hVdqspZl2_0),.clk(gclk));
	jdff dff_A_u1mu6W740_0(.dout(w_dff_A_KCMgCse62_0),.din(w_dff_A_u1mu6W740_0),.clk(gclk));
	jdff dff_A_KCMgCse62_0(.dout(w_dff_A_TvsniWpr4_0),.din(w_dff_A_KCMgCse62_0),.clk(gclk));
	jdff dff_A_TvsniWpr4_0(.dout(w_dff_A_K1YnwdvK1_0),.din(w_dff_A_TvsniWpr4_0),.clk(gclk));
	jdff dff_A_K1YnwdvK1_0(.dout(w_dff_A_72m3X7Vd2_0),.din(w_dff_A_K1YnwdvK1_0),.clk(gclk));
	jdff dff_A_72m3X7Vd2_0(.dout(w_dff_A_CrKFiCqf1_0),.din(w_dff_A_72m3X7Vd2_0),.clk(gclk));
	jdff dff_A_CrKFiCqf1_0(.dout(w_dff_A_dahJqzWt9_0),.din(w_dff_A_CrKFiCqf1_0),.clk(gclk));
	jdff dff_A_dahJqzWt9_0(.dout(w_dff_A_HkFVYLsx4_0),.din(w_dff_A_dahJqzWt9_0),.clk(gclk));
	jdff dff_A_HkFVYLsx4_0(.dout(w_dff_A_U61jtEFG5_0),.din(w_dff_A_HkFVYLsx4_0),.clk(gclk));
	jdff dff_A_U61jtEFG5_0(.dout(w_dff_A_G2CYWKhS2_0),.din(w_dff_A_U61jtEFG5_0),.clk(gclk));
	jdff dff_A_G2CYWKhS2_0(.dout(w_dff_A_deKqIOxp6_0),.din(w_dff_A_G2CYWKhS2_0),.clk(gclk));
	jdff dff_A_deKqIOxp6_0(.dout(w_dff_A_jTlifDtK4_0),.din(w_dff_A_deKqIOxp6_0),.clk(gclk));
	jdff dff_A_jTlifDtK4_0(.dout(w_dff_A_7E3bbe5x1_0),.din(w_dff_A_jTlifDtK4_0),.clk(gclk));
	jdff dff_A_7E3bbe5x1_0(.dout(w_dff_A_49Gda4N82_0),.din(w_dff_A_7E3bbe5x1_0),.clk(gclk));
	jdff dff_A_49Gda4N82_0(.dout(G2223gat),.din(w_dff_A_49Gda4N82_0),.clk(gclk));
	jdff dff_A_u59OK6MR6_2(.dout(w_dff_A_AUDRS8GG1_0),.din(w_dff_A_u59OK6MR6_2),.clk(gclk));
	jdff dff_A_AUDRS8GG1_0(.dout(w_dff_A_EdpmgK5y6_0),.din(w_dff_A_AUDRS8GG1_0),.clk(gclk));
	jdff dff_A_EdpmgK5y6_0(.dout(w_dff_A_ZiAS5RSm0_0),.din(w_dff_A_EdpmgK5y6_0),.clk(gclk));
	jdff dff_A_ZiAS5RSm0_0(.dout(w_dff_A_nBUqx7vL4_0),.din(w_dff_A_ZiAS5RSm0_0),.clk(gclk));
	jdff dff_A_nBUqx7vL4_0(.dout(w_dff_A_Tcg6oiJu6_0),.din(w_dff_A_nBUqx7vL4_0),.clk(gclk));
	jdff dff_A_Tcg6oiJu6_0(.dout(w_dff_A_z0wpr7zP6_0),.din(w_dff_A_Tcg6oiJu6_0),.clk(gclk));
	jdff dff_A_z0wpr7zP6_0(.dout(w_dff_A_6gqQAzuL4_0),.din(w_dff_A_z0wpr7zP6_0),.clk(gclk));
	jdff dff_A_6gqQAzuL4_0(.dout(w_dff_A_APpQpcHi8_0),.din(w_dff_A_6gqQAzuL4_0),.clk(gclk));
	jdff dff_A_APpQpcHi8_0(.dout(w_dff_A_nyLnwlWy9_0),.din(w_dff_A_APpQpcHi8_0),.clk(gclk));
	jdff dff_A_nyLnwlWy9_0(.dout(w_dff_A_tbpEb7BY9_0),.din(w_dff_A_nyLnwlWy9_0),.clk(gclk));
	jdff dff_A_tbpEb7BY9_0(.dout(w_dff_A_rOIcZZDu9_0),.din(w_dff_A_tbpEb7BY9_0),.clk(gclk));
	jdff dff_A_rOIcZZDu9_0(.dout(w_dff_A_Ja78ZvCe2_0),.din(w_dff_A_rOIcZZDu9_0),.clk(gclk));
	jdff dff_A_Ja78ZvCe2_0(.dout(w_dff_A_CXGxDzkH2_0),.din(w_dff_A_Ja78ZvCe2_0),.clk(gclk));
	jdff dff_A_CXGxDzkH2_0(.dout(w_dff_A_pnrcnN4J1_0),.din(w_dff_A_CXGxDzkH2_0),.clk(gclk));
	jdff dff_A_pnrcnN4J1_0(.dout(w_dff_A_UGT5LskC9_0),.din(w_dff_A_pnrcnN4J1_0),.clk(gclk));
	jdff dff_A_UGT5LskC9_0(.dout(w_dff_A_AeEhZNnb2_0),.din(w_dff_A_UGT5LskC9_0),.clk(gclk));
	jdff dff_A_AeEhZNnb2_0(.dout(w_dff_A_hJBYENos7_0),.din(w_dff_A_AeEhZNnb2_0),.clk(gclk));
	jdff dff_A_hJBYENos7_0(.dout(w_dff_A_AjK0qOSk1_0),.din(w_dff_A_hJBYENos7_0),.clk(gclk));
	jdff dff_A_AjK0qOSk1_0(.dout(w_dff_A_GBYgOpBd7_0),.din(w_dff_A_AjK0qOSk1_0),.clk(gclk));
	jdff dff_A_GBYgOpBd7_0(.dout(w_dff_A_QnVD2dQL5_0),.din(w_dff_A_GBYgOpBd7_0),.clk(gclk));
	jdff dff_A_QnVD2dQL5_0(.dout(w_dff_A_Fl6TlHCf6_0),.din(w_dff_A_QnVD2dQL5_0),.clk(gclk));
	jdff dff_A_Fl6TlHCf6_0(.dout(w_dff_A_FbLdgRgn8_0),.din(w_dff_A_Fl6TlHCf6_0),.clk(gclk));
	jdff dff_A_FbLdgRgn8_0(.dout(w_dff_A_wZULdw2L9_0),.din(w_dff_A_FbLdgRgn8_0),.clk(gclk));
	jdff dff_A_wZULdw2L9_0(.dout(w_dff_A_QFUs9Ila8_0),.din(w_dff_A_wZULdw2L9_0),.clk(gclk));
	jdff dff_A_QFUs9Ila8_0(.dout(w_dff_A_wJOokmHS5_0),.din(w_dff_A_QFUs9Ila8_0),.clk(gclk));
	jdff dff_A_wJOokmHS5_0(.dout(w_dff_A_dEmfk64u5_0),.din(w_dff_A_wJOokmHS5_0),.clk(gclk));
	jdff dff_A_dEmfk64u5_0(.dout(w_dff_A_FVKsp7M03_0),.din(w_dff_A_dEmfk64u5_0),.clk(gclk));
	jdff dff_A_FVKsp7M03_0(.dout(w_dff_A_MvLXYLxv5_0),.din(w_dff_A_FVKsp7M03_0),.clk(gclk));
	jdff dff_A_MvLXYLxv5_0(.dout(w_dff_A_CFZpnAs40_0),.din(w_dff_A_MvLXYLxv5_0),.clk(gclk));
	jdff dff_A_CFZpnAs40_0(.dout(w_dff_A_LD930DMu4_0),.din(w_dff_A_CFZpnAs40_0),.clk(gclk));
	jdff dff_A_LD930DMu4_0(.dout(w_dff_A_40sP0Bmi0_0),.din(w_dff_A_LD930DMu4_0),.clk(gclk));
	jdff dff_A_40sP0Bmi0_0(.dout(w_dff_A_PY1Wxqvw7_0),.din(w_dff_A_40sP0Bmi0_0),.clk(gclk));
	jdff dff_A_PY1Wxqvw7_0(.dout(w_dff_A_Nk71cV790_0),.din(w_dff_A_PY1Wxqvw7_0),.clk(gclk));
	jdff dff_A_Nk71cV790_0(.dout(w_dff_A_EvxITJEX9_0),.din(w_dff_A_Nk71cV790_0),.clk(gclk));
	jdff dff_A_EvxITJEX9_0(.dout(w_dff_A_Kqrr3aOs4_0),.din(w_dff_A_EvxITJEX9_0),.clk(gclk));
	jdff dff_A_Kqrr3aOs4_0(.dout(w_dff_A_uYbfkqNb0_0),.din(w_dff_A_Kqrr3aOs4_0),.clk(gclk));
	jdff dff_A_uYbfkqNb0_0(.dout(w_dff_A_ysW22CG84_0),.din(w_dff_A_uYbfkqNb0_0),.clk(gclk));
	jdff dff_A_ysW22CG84_0(.dout(w_dff_A_io4ikEzF2_0),.din(w_dff_A_ysW22CG84_0),.clk(gclk));
	jdff dff_A_io4ikEzF2_0(.dout(w_dff_A_R0kt95vW2_0),.din(w_dff_A_io4ikEzF2_0),.clk(gclk));
	jdff dff_A_R0kt95vW2_0(.dout(w_dff_A_3pPmDxCy2_0),.din(w_dff_A_R0kt95vW2_0),.clk(gclk));
	jdff dff_A_3pPmDxCy2_0(.dout(w_dff_A_cS8XrOzc9_0),.din(w_dff_A_3pPmDxCy2_0),.clk(gclk));
	jdff dff_A_cS8XrOzc9_0(.dout(w_dff_A_G4B3b3nI4_0),.din(w_dff_A_cS8XrOzc9_0),.clk(gclk));
	jdff dff_A_G4B3b3nI4_0(.dout(w_dff_A_v8EUxYoE6_0),.din(w_dff_A_G4B3b3nI4_0),.clk(gclk));
	jdff dff_A_v8EUxYoE6_0(.dout(w_dff_A_W1ZfZD3z6_0),.din(w_dff_A_v8EUxYoE6_0),.clk(gclk));
	jdff dff_A_W1ZfZD3z6_0(.dout(w_dff_A_MYsLJGFR8_0),.din(w_dff_A_W1ZfZD3z6_0),.clk(gclk));
	jdff dff_A_MYsLJGFR8_0(.dout(w_dff_A_wR71dWOy1_0),.din(w_dff_A_MYsLJGFR8_0),.clk(gclk));
	jdff dff_A_wR71dWOy1_0(.dout(w_dff_A_xFfKk3BB7_0),.din(w_dff_A_wR71dWOy1_0),.clk(gclk));
	jdff dff_A_xFfKk3BB7_0(.dout(w_dff_A_EPvQzi5F2_0),.din(w_dff_A_xFfKk3BB7_0),.clk(gclk));
	jdff dff_A_EPvQzi5F2_0(.dout(w_dff_A_S1jL8bHB9_0),.din(w_dff_A_EPvQzi5F2_0),.clk(gclk));
	jdff dff_A_S1jL8bHB9_0(.dout(w_dff_A_HnpzXgXD2_0),.din(w_dff_A_S1jL8bHB9_0),.clk(gclk));
	jdff dff_A_HnpzXgXD2_0(.dout(w_dff_A_8AIsEPAw5_0),.din(w_dff_A_HnpzXgXD2_0),.clk(gclk));
	jdff dff_A_8AIsEPAw5_0(.dout(w_dff_A_qpXikVWH1_0),.din(w_dff_A_8AIsEPAw5_0),.clk(gclk));
	jdff dff_A_qpXikVWH1_0(.dout(w_dff_A_09EW2rDW4_0),.din(w_dff_A_qpXikVWH1_0),.clk(gclk));
	jdff dff_A_09EW2rDW4_0(.dout(w_dff_A_fR8LNZsj5_0),.din(w_dff_A_09EW2rDW4_0),.clk(gclk));
	jdff dff_A_fR8LNZsj5_0(.dout(w_dff_A_gArMwLcF2_0),.din(w_dff_A_fR8LNZsj5_0),.clk(gclk));
	jdff dff_A_gArMwLcF2_0(.dout(w_dff_A_csHlvfVS8_0),.din(w_dff_A_gArMwLcF2_0),.clk(gclk));
	jdff dff_A_csHlvfVS8_0(.dout(w_dff_A_qaoRYh0E1_0),.din(w_dff_A_csHlvfVS8_0),.clk(gclk));
	jdff dff_A_qaoRYh0E1_0(.dout(w_dff_A_Ocxo46xu6_0),.din(w_dff_A_qaoRYh0E1_0),.clk(gclk));
	jdff dff_A_Ocxo46xu6_0(.dout(w_dff_A_KGlUjaKO8_0),.din(w_dff_A_Ocxo46xu6_0),.clk(gclk));
	jdff dff_A_KGlUjaKO8_0(.dout(w_dff_A_gkNXnR409_0),.din(w_dff_A_KGlUjaKO8_0),.clk(gclk));
	jdff dff_A_gkNXnR409_0(.dout(w_dff_A_nbpHtQDg8_0),.din(w_dff_A_gkNXnR409_0),.clk(gclk));
	jdff dff_A_nbpHtQDg8_0(.dout(w_dff_A_xu0HXtiL9_0),.din(w_dff_A_nbpHtQDg8_0),.clk(gclk));
	jdff dff_A_xu0HXtiL9_0(.dout(G2548gat),.din(w_dff_A_xu0HXtiL9_0),.clk(gclk));
	jdff dff_A_RUYPQsDY7_2(.dout(w_dff_A_FERBmCp34_0),.din(w_dff_A_RUYPQsDY7_2),.clk(gclk));
	jdff dff_A_FERBmCp34_0(.dout(w_dff_A_lSRreIfz1_0),.din(w_dff_A_FERBmCp34_0),.clk(gclk));
	jdff dff_A_lSRreIfz1_0(.dout(w_dff_A_D8PKPrPK0_0),.din(w_dff_A_lSRreIfz1_0),.clk(gclk));
	jdff dff_A_D8PKPrPK0_0(.dout(w_dff_A_Wgwibnsv3_0),.din(w_dff_A_D8PKPrPK0_0),.clk(gclk));
	jdff dff_A_Wgwibnsv3_0(.dout(w_dff_A_3c7oaCSD7_0),.din(w_dff_A_Wgwibnsv3_0),.clk(gclk));
	jdff dff_A_3c7oaCSD7_0(.dout(w_dff_A_i9vTsd9D9_0),.din(w_dff_A_3c7oaCSD7_0),.clk(gclk));
	jdff dff_A_i9vTsd9D9_0(.dout(w_dff_A_aYXvXpA00_0),.din(w_dff_A_i9vTsd9D9_0),.clk(gclk));
	jdff dff_A_aYXvXpA00_0(.dout(w_dff_A_gqknKMfQ0_0),.din(w_dff_A_aYXvXpA00_0),.clk(gclk));
	jdff dff_A_gqknKMfQ0_0(.dout(w_dff_A_fKVkzAPb6_0),.din(w_dff_A_gqknKMfQ0_0),.clk(gclk));
	jdff dff_A_fKVkzAPb6_0(.dout(w_dff_A_J1woOXAB6_0),.din(w_dff_A_fKVkzAPb6_0),.clk(gclk));
	jdff dff_A_J1woOXAB6_0(.dout(w_dff_A_RDyDpIKL3_0),.din(w_dff_A_J1woOXAB6_0),.clk(gclk));
	jdff dff_A_RDyDpIKL3_0(.dout(w_dff_A_tGrCqxOn3_0),.din(w_dff_A_RDyDpIKL3_0),.clk(gclk));
	jdff dff_A_tGrCqxOn3_0(.dout(w_dff_A_TNghpsKr9_0),.din(w_dff_A_tGrCqxOn3_0),.clk(gclk));
	jdff dff_A_TNghpsKr9_0(.dout(w_dff_A_B9jwKtEi0_0),.din(w_dff_A_TNghpsKr9_0),.clk(gclk));
	jdff dff_A_B9jwKtEi0_0(.dout(w_dff_A_Mh1ZkqB01_0),.din(w_dff_A_B9jwKtEi0_0),.clk(gclk));
	jdff dff_A_Mh1ZkqB01_0(.dout(w_dff_A_zDZVouRh0_0),.din(w_dff_A_Mh1ZkqB01_0),.clk(gclk));
	jdff dff_A_zDZVouRh0_0(.dout(w_dff_A_yUimV0Bh9_0),.din(w_dff_A_zDZVouRh0_0),.clk(gclk));
	jdff dff_A_yUimV0Bh9_0(.dout(w_dff_A_RAueuALN5_0),.din(w_dff_A_yUimV0Bh9_0),.clk(gclk));
	jdff dff_A_RAueuALN5_0(.dout(w_dff_A_AxMvzLU83_0),.din(w_dff_A_RAueuALN5_0),.clk(gclk));
	jdff dff_A_AxMvzLU83_0(.dout(w_dff_A_3gSVC3rH2_0),.din(w_dff_A_AxMvzLU83_0),.clk(gclk));
	jdff dff_A_3gSVC3rH2_0(.dout(w_dff_A_awNIhsVs6_0),.din(w_dff_A_3gSVC3rH2_0),.clk(gclk));
	jdff dff_A_awNIhsVs6_0(.dout(w_dff_A_G3QlGVPr3_0),.din(w_dff_A_awNIhsVs6_0),.clk(gclk));
	jdff dff_A_G3QlGVPr3_0(.dout(w_dff_A_RhKMlQyO5_0),.din(w_dff_A_G3QlGVPr3_0),.clk(gclk));
	jdff dff_A_RhKMlQyO5_0(.dout(w_dff_A_QQyIJLSQ3_0),.din(w_dff_A_RhKMlQyO5_0),.clk(gclk));
	jdff dff_A_QQyIJLSQ3_0(.dout(w_dff_A_O1DAztnV3_0),.din(w_dff_A_QQyIJLSQ3_0),.clk(gclk));
	jdff dff_A_O1DAztnV3_0(.dout(w_dff_A_QxPjcjDw3_0),.din(w_dff_A_O1DAztnV3_0),.clk(gclk));
	jdff dff_A_QxPjcjDw3_0(.dout(w_dff_A_8Uat7pf94_0),.din(w_dff_A_QxPjcjDw3_0),.clk(gclk));
	jdff dff_A_8Uat7pf94_0(.dout(w_dff_A_r8XYs8Hd3_0),.din(w_dff_A_8Uat7pf94_0),.clk(gclk));
	jdff dff_A_r8XYs8Hd3_0(.dout(w_dff_A_BdxTEUHS9_0),.din(w_dff_A_r8XYs8Hd3_0),.clk(gclk));
	jdff dff_A_BdxTEUHS9_0(.dout(w_dff_A_qpsctrvC1_0),.din(w_dff_A_BdxTEUHS9_0),.clk(gclk));
	jdff dff_A_qpsctrvC1_0(.dout(w_dff_A_lpZGXu0y2_0),.din(w_dff_A_qpsctrvC1_0),.clk(gclk));
	jdff dff_A_lpZGXu0y2_0(.dout(w_dff_A_19fCI6Zc0_0),.din(w_dff_A_lpZGXu0y2_0),.clk(gclk));
	jdff dff_A_19fCI6Zc0_0(.dout(w_dff_A_XybjtclJ7_0),.din(w_dff_A_19fCI6Zc0_0),.clk(gclk));
	jdff dff_A_XybjtclJ7_0(.dout(w_dff_A_Czx8K6yD4_0),.din(w_dff_A_XybjtclJ7_0),.clk(gclk));
	jdff dff_A_Czx8K6yD4_0(.dout(w_dff_A_R9sSCIk98_0),.din(w_dff_A_Czx8K6yD4_0),.clk(gclk));
	jdff dff_A_R9sSCIk98_0(.dout(w_dff_A_dn38EZaj9_0),.din(w_dff_A_R9sSCIk98_0),.clk(gclk));
	jdff dff_A_dn38EZaj9_0(.dout(w_dff_A_uQOZSzyv7_0),.din(w_dff_A_dn38EZaj9_0),.clk(gclk));
	jdff dff_A_uQOZSzyv7_0(.dout(w_dff_A_YKdDcgJM5_0),.din(w_dff_A_uQOZSzyv7_0),.clk(gclk));
	jdff dff_A_YKdDcgJM5_0(.dout(w_dff_A_Rj33y8Qg2_0),.din(w_dff_A_YKdDcgJM5_0),.clk(gclk));
	jdff dff_A_Rj33y8Qg2_0(.dout(w_dff_A_H0xHfJn59_0),.din(w_dff_A_Rj33y8Qg2_0),.clk(gclk));
	jdff dff_A_H0xHfJn59_0(.dout(w_dff_A_joOw27Ci1_0),.din(w_dff_A_H0xHfJn59_0),.clk(gclk));
	jdff dff_A_joOw27Ci1_0(.dout(w_dff_A_SH4AX4Fe8_0),.din(w_dff_A_joOw27Ci1_0),.clk(gclk));
	jdff dff_A_SH4AX4Fe8_0(.dout(w_dff_A_YIkkrbas4_0),.din(w_dff_A_SH4AX4Fe8_0),.clk(gclk));
	jdff dff_A_YIkkrbas4_0(.dout(w_dff_A_bnRvhZUK2_0),.din(w_dff_A_YIkkrbas4_0),.clk(gclk));
	jdff dff_A_bnRvhZUK2_0(.dout(w_dff_A_Np5uqXUX6_0),.din(w_dff_A_bnRvhZUK2_0),.clk(gclk));
	jdff dff_A_Np5uqXUX6_0(.dout(w_dff_A_xgSBFmNI2_0),.din(w_dff_A_Np5uqXUX6_0),.clk(gclk));
	jdff dff_A_xgSBFmNI2_0(.dout(w_dff_A_MD9CjD6p0_0),.din(w_dff_A_xgSBFmNI2_0),.clk(gclk));
	jdff dff_A_MD9CjD6p0_0(.dout(w_dff_A_IMUfPG2y2_0),.din(w_dff_A_MD9CjD6p0_0),.clk(gclk));
	jdff dff_A_IMUfPG2y2_0(.dout(w_dff_A_jz5MI4T16_0),.din(w_dff_A_IMUfPG2y2_0),.clk(gclk));
	jdff dff_A_jz5MI4T16_0(.dout(w_dff_A_8MbgAvdt1_0),.din(w_dff_A_jz5MI4T16_0),.clk(gclk));
	jdff dff_A_8MbgAvdt1_0(.dout(w_dff_A_hvHqZMJY9_0),.din(w_dff_A_8MbgAvdt1_0),.clk(gclk));
	jdff dff_A_hvHqZMJY9_0(.dout(w_dff_A_0kYKmnQE1_0),.din(w_dff_A_hvHqZMJY9_0),.clk(gclk));
	jdff dff_A_0kYKmnQE1_0(.dout(w_dff_A_3K3I5SLN9_0),.din(w_dff_A_0kYKmnQE1_0),.clk(gclk));
	jdff dff_A_3K3I5SLN9_0(.dout(w_dff_A_hsBftZC11_0),.din(w_dff_A_3K3I5SLN9_0),.clk(gclk));
	jdff dff_A_hsBftZC11_0(.dout(w_dff_A_fj6EaFpb0_0),.din(w_dff_A_hsBftZC11_0),.clk(gclk));
	jdff dff_A_fj6EaFpb0_0(.dout(w_dff_A_f4420IxB5_0),.din(w_dff_A_fj6EaFpb0_0),.clk(gclk));
	jdff dff_A_f4420IxB5_0(.dout(w_dff_A_wn5HowOg8_0),.din(w_dff_A_f4420IxB5_0),.clk(gclk));
	jdff dff_A_wn5HowOg8_0(.dout(w_dff_A_I9IweMtn6_0),.din(w_dff_A_wn5HowOg8_0),.clk(gclk));
	jdff dff_A_I9IweMtn6_0(.dout(w_dff_A_XQpzOOFe4_0),.din(w_dff_A_I9IweMtn6_0),.clk(gclk));
	jdff dff_A_XQpzOOFe4_0(.dout(G2877gat),.din(w_dff_A_XQpzOOFe4_0),.clk(gclk));
	jdff dff_A_3cNNDt623_2(.dout(w_dff_A_OeD4kmTb0_0),.din(w_dff_A_3cNNDt623_2),.clk(gclk));
	jdff dff_A_OeD4kmTb0_0(.dout(w_dff_A_gbjDoEu50_0),.din(w_dff_A_OeD4kmTb0_0),.clk(gclk));
	jdff dff_A_gbjDoEu50_0(.dout(w_dff_A_sti6URCX3_0),.din(w_dff_A_gbjDoEu50_0),.clk(gclk));
	jdff dff_A_sti6URCX3_0(.dout(w_dff_A_Ixj4wH3s3_0),.din(w_dff_A_sti6URCX3_0),.clk(gclk));
	jdff dff_A_Ixj4wH3s3_0(.dout(w_dff_A_zqHGa9GZ9_0),.din(w_dff_A_Ixj4wH3s3_0),.clk(gclk));
	jdff dff_A_zqHGa9GZ9_0(.dout(w_dff_A_A4V818kf7_0),.din(w_dff_A_zqHGa9GZ9_0),.clk(gclk));
	jdff dff_A_A4V818kf7_0(.dout(w_dff_A_d8LqlvIK9_0),.din(w_dff_A_A4V818kf7_0),.clk(gclk));
	jdff dff_A_d8LqlvIK9_0(.dout(w_dff_A_incpz5RR2_0),.din(w_dff_A_d8LqlvIK9_0),.clk(gclk));
	jdff dff_A_incpz5RR2_0(.dout(w_dff_A_SDcD5pXx9_0),.din(w_dff_A_incpz5RR2_0),.clk(gclk));
	jdff dff_A_SDcD5pXx9_0(.dout(w_dff_A_UIl9BgcD5_0),.din(w_dff_A_SDcD5pXx9_0),.clk(gclk));
	jdff dff_A_UIl9BgcD5_0(.dout(w_dff_A_oZzv7tR73_0),.din(w_dff_A_UIl9BgcD5_0),.clk(gclk));
	jdff dff_A_oZzv7tR73_0(.dout(w_dff_A_RwzAJwkD4_0),.din(w_dff_A_oZzv7tR73_0),.clk(gclk));
	jdff dff_A_RwzAJwkD4_0(.dout(w_dff_A_z4swIlhP5_0),.din(w_dff_A_RwzAJwkD4_0),.clk(gclk));
	jdff dff_A_z4swIlhP5_0(.dout(w_dff_A_ET5BbgDx8_0),.din(w_dff_A_z4swIlhP5_0),.clk(gclk));
	jdff dff_A_ET5BbgDx8_0(.dout(w_dff_A_dLTlhKMU5_0),.din(w_dff_A_ET5BbgDx8_0),.clk(gclk));
	jdff dff_A_dLTlhKMU5_0(.dout(w_dff_A_EIOYCWZT6_0),.din(w_dff_A_dLTlhKMU5_0),.clk(gclk));
	jdff dff_A_EIOYCWZT6_0(.dout(w_dff_A_i55dgTbi1_0),.din(w_dff_A_EIOYCWZT6_0),.clk(gclk));
	jdff dff_A_i55dgTbi1_0(.dout(w_dff_A_lv79t8RY6_0),.din(w_dff_A_i55dgTbi1_0),.clk(gclk));
	jdff dff_A_lv79t8RY6_0(.dout(w_dff_A_m3MsK69G3_0),.din(w_dff_A_lv79t8RY6_0),.clk(gclk));
	jdff dff_A_m3MsK69G3_0(.dout(w_dff_A_wWCHn3aI2_0),.din(w_dff_A_m3MsK69G3_0),.clk(gclk));
	jdff dff_A_wWCHn3aI2_0(.dout(w_dff_A_QYU6znvH3_0),.din(w_dff_A_wWCHn3aI2_0),.clk(gclk));
	jdff dff_A_QYU6znvH3_0(.dout(w_dff_A_Yf2eC9iE3_0),.din(w_dff_A_QYU6znvH3_0),.clk(gclk));
	jdff dff_A_Yf2eC9iE3_0(.dout(w_dff_A_x75KIasX8_0),.din(w_dff_A_Yf2eC9iE3_0),.clk(gclk));
	jdff dff_A_x75KIasX8_0(.dout(w_dff_A_cGlLDSgH2_0),.din(w_dff_A_x75KIasX8_0),.clk(gclk));
	jdff dff_A_cGlLDSgH2_0(.dout(w_dff_A_4BGdnQu19_0),.din(w_dff_A_cGlLDSgH2_0),.clk(gclk));
	jdff dff_A_4BGdnQu19_0(.dout(w_dff_A_aWzaHUEc1_0),.din(w_dff_A_4BGdnQu19_0),.clk(gclk));
	jdff dff_A_aWzaHUEc1_0(.dout(w_dff_A_IMY3fq3d2_0),.din(w_dff_A_aWzaHUEc1_0),.clk(gclk));
	jdff dff_A_IMY3fq3d2_0(.dout(w_dff_A_TfhU36SW1_0),.din(w_dff_A_IMY3fq3d2_0),.clk(gclk));
	jdff dff_A_TfhU36SW1_0(.dout(w_dff_A_8aFoTaVN9_0),.din(w_dff_A_TfhU36SW1_0),.clk(gclk));
	jdff dff_A_8aFoTaVN9_0(.dout(w_dff_A_tZSNMhT42_0),.din(w_dff_A_8aFoTaVN9_0),.clk(gclk));
	jdff dff_A_tZSNMhT42_0(.dout(w_dff_A_P5Laq6MP6_0),.din(w_dff_A_tZSNMhT42_0),.clk(gclk));
	jdff dff_A_P5Laq6MP6_0(.dout(w_dff_A_XhvDV9rF2_0),.din(w_dff_A_P5Laq6MP6_0),.clk(gclk));
	jdff dff_A_XhvDV9rF2_0(.dout(w_dff_A_lcAp889A4_0),.din(w_dff_A_XhvDV9rF2_0),.clk(gclk));
	jdff dff_A_lcAp889A4_0(.dout(w_dff_A_urBqOGvO9_0),.din(w_dff_A_lcAp889A4_0),.clk(gclk));
	jdff dff_A_urBqOGvO9_0(.dout(w_dff_A_h5UpJryP1_0),.din(w_dff_A_urBqOGvO9_0),.clk(gclk));
	jdff dff_A_h5UpJryP1_0(.dout(w_dff_A_V3mBh8Xe1_0),.din(w_dff_A_h5UpJryP1_0),.clk(gclk));
	jdff dff_A_V3mBh8Xe1_0(.dout(w_dff_A_VVRS5WCw3_0),.din(w_dff_A_V3mBh8Xe1_0),.clk(gclk));
	jdff dff_A_VVRS5WCw3_0(.dout(w_dff_A_KQEBDqy60_0),.din(w_dff_A_VVRS5WCw3_0),.clk(gclk));
	jdff dff_A_KQEBDqy60_0(.dout(w_dff_A_mGKEe4Tn7_0),.din(w_dff_A_KQEBDqy60_0),.clk(gclk));
	jdff dff_A_mGKEe4Tn7_0(.dout(w_dff_A_MdjoMgUH1_0),.din(w_dff_A_mGKEe4Tn7_0),.clk(gclk));
	jdff dff_A_MdjoMgUH1_0(.dout(w_dff_A_GD3P4vfF6_0),.din(w_dff_A_MdjoMgUH1_0),.clk(gclk));
	jdff dff_A_GD3P4vfF6_0(.dout(w_dff_A_SPWjq15W3_0),.din(w_dff_A_GD3P4vfF6_0),.clk(gclk));
	jdff dff_A_SPWjq15W3_0(.dout(w_dff_A_SuSjSHB70_0),.din(w_dff_A_SPWjq15W3_0),.clk(gclk));
	jdff dff_A_SuSjSHB70_0(.dout(w_dff_A_KOXpkjoS4_0),.din(w_dff_A_SuSjSHB70_0),.clk(gclk));
	jdff dff_A_KOXpkjoS4_0(.dout(w_dff_A_rPFu5ZpZ8_0),.din(w_dff_A_KOXpkjoS4_0),.clk(gclk));
	jdff dff_A_rPFu5ZpZ8_0(.dout(w_dff_A_Y70DArRS4_0),.din(w_dff_A_rPFu5ZpZ8_0),.clk(gclk));
	jdff dff_A_Y70DArRS4_0(.dout(w_dff_A_nagS59Gw5_0),.din(w_dff_A_Y70DArRS4_0),.clk(gclk));
	jdff dff_A_nagS59Gw5_0(.dout(w_dff_A_DBTLQpSv1_0),.din(w_dff_A_nagS59Gw5_0),.clk(gclk));
	jdff dff_A_DBTLQpSv1_0(.dout(w_dff_A_BWCZocTP7_0),.din(w_dff_A_DBTLQpSv1_0),.clk(gclk));
	jdff dff_A_BWCZocTP7_0(.dout(w_dff_A_qZ22fWx69_0),.din(w_dff_A_BWCZocTP7_0),.clk(gclk));
	jdff dff_A_qZ22fWx69_0(.dout(w_dff_A_XXBn1gv58_0),.din(w_dff_A_qZ22fWx69_0),.clk(gclk));
	jdff dff_A_XXBn1gv58_0(.dout(w_dff_A_z29R41yA9_0),.din(w_dff_A_XXBn1gv58_0),.clk(gclk));
	jdff dff_A_z29R41yA9_0(.dout(w_dff_A_2oBeUSdY0_0),.din(w_dff_A_z29R41yA9_0),.clk(gclk));
	jdff dff_A_2oBeUSdY0_0(.dout(w_dff_A_XdntmXwb6_0),.din(w_dff_A_2oBeUSdY0_0),.clk(gclk));
	jdff dff_A_XdntmXwb6_0(.dout(w_dff_A_1KEcECGy0_0),.din(w_dff_A_XdntmXwb6_0),.clk(gclk));
	jdff dff_A_1KEcECGy0_0(.dout(w_dff_A_yJ4EGLoz5_0),.din(w_dff_A_1KEcECGy0_0),.clk(gclk));
	jdff dff_A_yJ4EGLoz5_0(.dout(G3211gat),.din(w_dff_A_yJ4EGLoz5_0),.clk(gclk));
	jdff dff_A_AWpHub178_2(.dout(w_dff_A_k1paZK0Y2_0),.din(w_dff_A_AWpHub178_2),.clk(gclk));
	jdff dff_A_k1paZK0Y2_0(.dout(w_dff_A_ijtJorKs5_0),.din(w_dff_A_k1paZK0Y2_0),.clk(gclk));
	jdff dff_A_ijtJorKs5_0(.dout(w_dff_A_DQ4C7Sfr2_0),.din(w_dff_A_ijtJorKs5_0),.clk(gclk));
	jdff dff_A_DQ4C7Sfr2_0(.dout(w_dff_A_Xxke3TNk9_0),.din(w_dff_A_DQ4C7Sfr2_0),.clk(gclk));
	jdff dff_A_Xxke3TNk9_0(.dout(w_dff_A_LOY1HQbs4_0),.din(w_dff_A_Xxke3TNk9_0),.clk(gclk));
	jdff dff_A_LOY1HQbs4_0(.dout(w_dff_A_n8Qrp2Vw8_0),.din(w_dff_A_LOY1HQbs4_0),.clk(gclk));
	jdff dff_A_n8Qrp2Vw8_0(.dout(w_dff_A_8teEXTp34_0),.din(w_dff_A_n8Qrp2Vw8_0),.clk(gclk));
	jdff dff_A_8teEXTp34_0(.dout(w_dff_A_iWRwJXu99_0),.din(w_dff_A_8teEXTp34_0),.clk(gclk));
	jdff dff_A_iWRwJXu99_0(.dout(w_dff_A_npqPB1Q28_0),.din(w_dff_A_iWRwJXu99_0),.clk(gclk));
	jdff dff_A_npqPB1Q28_0(.dout(w_dff_A_oijkPitJ0_0),.din(w_dff_A_npqPB1Q28_0),.clk(gclk));
	jdff dff_A_oijkPitJ0_0(.dout(w_dff_A_vZkmqeXs2_0),.din(w_dff_A_oijkPitJ0_0),.clk(gclk));
	jdff dff_A_vZkmqeXs2_0(.dout(w_dff_A_OU5mnSOI7_0),.din(w_dff_A_vZkmqeXs2_0),.clk(gclk));
	jdff dff_A_OU5mnSOI7_0(.dout(w_dff_A_0Ej9uaVS9_0),.din(w_dff_A_OU5mnSOI7_0),.clk(gclk));
	jdff dff_A_0Ej9uaVS9_0(.dout(w_dff_A_hmWynH6E1_0),.din(w_dff_A_0Ej9uaVS9_0),.clk(gclk));
	jdff dff_A_hmWynH6E1_0(.dout(w_dff_A_IAEEHCxV1_0),.din(w_dff_A_hmWynH6E1_0),.clk(gclk));
	jdff dff_A_IAEEHCxV1_0(.dout(w_dff_A_R06KiJGO1_0),.din(w_dff_A_IAEEHCxV1_0),.clk(gclk));
	jdff dff_A_R06KiJGO1_0(.dout(w_dff_A_xgL3MgNv9_0),.din(w_dff_A_R06KiJGO1_0),.clk(gclk));
	jdff dff_A_xgL3MgNv9_0(.dout(w_dff_A_BPh9lray7_0),.din(w_dff_A_xgL3MgNv9_0),.clk(gclk));
	jdff dff_A_BPh9lray7_0(.dout(w_dff_A_AxcYoavu9_0),.din(w_dff_A_BPh9lray7_0),.clk(gclk));
	jdff dff_A_AxcYoavu9_0(.dout(w_dff_A_VHTLPc0a7_0),.din(w_dff_A_AxcYoavu9_0),.clk(gclk));
	jdff dff_A_VHTLPc0a7_0(.dout(w_dff_A_AcMpOlLu9_0),.din(w_dff_A_VHTLPc0a7_0),.clk(gclk));
	jdff dff_A_AcMpOlLu9_0(.dout(w_dff_A_3mqbvP4W1_0),.din(w_dff_A_AcMpOlLu9_0),.clk(gclk));
	jdff dff_A_3mqbvP4W1_0(.dout(w_dff_A_lecah2h29_0),.din(w_dff_A_3mqbvP4W1_0),.clk(gclk));
	jdff dff_A_lecah2h29_0(.dout(w_dff_A_0yWtDODy3_0),.din(w_dff_A_lecah2h29_0),.clk(gclk));
	jdff dff_A_0yWtDODy3_0(.dout(w_dff_A_roPLPGKs4_0),.din(w_dff_A_0yWtDODy3_0),.clk(gclk));
	jdff dff_A_roPLPGKs4_0(.dout(w_dff_A_rfVEkmun7_0),.din(w_dff_A_roPLPGKs4_0),.clk(gclk));
	jdff dff_A_rfVEkmun7_0(.dout(w_dff_A_9nAAV3iw0_0),.din(w_dff_A_rfVEkmun7_0),.clk(gclk));
	jdff dff_A_9nAAV3iw0_0(.dout(w_dff_A_MbeVzEdF9_0),.din(w_dff_A_9nAAV3iw0_0),.clk(gclk));
	jdff dff_A_MbeVzEdF9_0(.dout(w_dff_A_oqXMtO5e1_0),.din(w_dff_A_MbeVzEdF9_0),.clk(gclk));
	jdff dff_A_oqXMtO5e1_0(.dout(w_dff_A_9iXITTRO2_0),.din(w_dff_A_oqXMtO5e1_0),.clk(gclk));
	jdff dff_A_9iXITTRO2_0(.dout(w_dff_A_bW12ClKR0_0),.din(w_dff_A_9iXITTRO2_0),.clk(gclk));
	jdff dff_A_bW12ClKR0_0(.dout(w_dff_A_BglbO1Nb1_0),.din(w_dff_A_bW12ClKR0_0),.clk(gclk));
	jdff dff_A_BglbO1Nb1_0(.dout(w_dff_A_ZKRWuKQ48_0),.din(w_dff_A_BglbO1Nb1_0),.clk(gclk));
	jdff dff_A_ZKRWuKQ48_0(.dout(w_dff_A_gUA9l13G5_0),.din(w_dff_A_ZKRWuKQ48_0),.clk(gclk));
	jdff dff_A_gUA9l13G5_0(.dout(w_dff_A_rYLWwpsi5_0),.din(w_dff_A_gUA9l13G5_0),.clk(gclk));
	jdff dff_A_rYLWwpsi5_0(.dout(w_dff_A_nNAihJVP2_0),.din(w_dff_A_rYLWwpsi5_0),.clk(gclk));
	jdff dff_A_nNAihJVP2_0(.dout(w_dff_A_KpCWsgbB6_0),.din(w_dff_A_nNAihJVP2_0),.clk(gclk));
	jdff dff_A_KpCWsgbB6_0(.dout(w_dff_A_5TP7WeBX6_0),.din(w_dff_A_KpCWsgbB6_0),.clk(gclk));
	jdff dff_A_5TP7WeBX6_0(.dout(w_dff_A_pwjGtfFN2_0),.din(w_dff_A_5TP7WeBX6_0),.clk(gclk));
	jdff dff_A_pwjGtfFN2_0(.dout(w_dff_A_Clh6yr2s4_0),.din(w_dff_A_pwjGtfFN2_0),.clk(gclk));
	jdff dff_A_Clh6yr2s4_0(.dout(w_dff_A_0bmlHtoQ2_0),.din(w_dff_A_Clh6yr2s4_0),.clk(gclk));
	jdff dff_A_0bmlHtoQ2_0(.dout(w_dff_A_NEVy6wJg0_0),.din(w_dff_A_0bmlHtoQ2_0),.clk(gclk));
	jdff dff_A_NEVy6wJg0_0(.dout(w_dff_A_AABDCGJa1_0),.din(w_dff_A_NEVy6wJg0_0),.clk(gclk));
	jdff dff_A_AABDCGJa1_0(.dout(w_dff_A_DyDEiMTR9_0),.din(w_dff_A_AABDCGJa1_0),.clk(gclk));
	jdff dff_A_DyDEiMTR9_0(.dout(w_dff_A_0CHITjur6_0),.din(w_dff_A_DyDEiMTR9_0),.clk(gclk));
	jdff dff_A_0CHITjur6_0(.dout(w_dff_A_NWFLROeL9_0),.din(w_dff_A_0CHITjur6_0),.clk(gclk));
	jdff dff_A_NWFLROeL9_0(.dout(w_dff_A_PrqbpDdw6_0),.din(w_dff_A_NWFLROeL9_0),.clk(gclk));
	jdff dff_A_PrqbpDdw6_0(.dout(w_dff_A_vBxmA6LB5_0),.din(w_dff_A_PrqbpDdw6_0),.clk(gclk));
	jdff dff_A_vBxmA6LB5_0(.dout(w_dff_A_YDg62S291_0),.din(w_dff_A_vBxmA6LB5_0),.clk(gclk));
	jdff dff_A_YDg62S291_0(.dout(w_dff_A_tGZYoIwU7_0),.din(w_dff_A_YDg62S291_0),.clk(gclk));
	jdff dff_A_tGZYoIwU7_0(.dout(w_dff_A_e41qEz0N0_0),.din(w_dff_A_tGZYoIwU7_0),.clk(gclk));
	jdff dff_A_e41qEz0N0_0(.dout(w_dff_A_XFF46Scq2_0),.din(w_dff_A_e41qEz0N0_0),.clk(gclk));
	jdff dff_A_XFF46Scq2_0(.dout(w_dff_A_E6Tczljx8_0),.din(w_dff_A_XFF46Scq2_0),.clk(gclk));
	jdff dff_A_E6Tczljx8_0(.dout(G3552gat),.din(w_dff_A_E6Tczljx8_0),.clk(gclk));
	jdff dff_A_8gCK9mkA1_2(.dout(w_dff_A_gZhCNXNw1_0),.din(w_dff_A_8gCK9mkA1_2),.clk(gclk));
	jdff dff_A_gZhCNXNw1_0(.dout(w_dff_A_JAUFx1H55_0),.din(w_dff_A_gZhCNXNw1_0),.clk(gclk));
	jdff dff_A_JAUFx1H55_0(.dout(w_dff_A_3vcoTw601_0),.din(w_dff_A_JAUFx1H55_0),.clk(gclk));
	jdff dff_A_3vcoTw601_0(.dout(w_dff_A_5YmVidb34_0),.din(w_dff_A_3vcoTw601_0),.clk(gclk));
	jdff dff_A_5YmVidb34_0(.dout(w_dff_A_5J3Q3rFA6_0),.din(w_dff_A_5YmVidb34_0),.clk(gclk));
	jdff dff_A_5J3Q3rFA6_0(.dout(w_dff_A_qAgfKp1R4_0),.din(w_dff_A_5J3Q3rFA6_0),.clk(gclk));
	jdff dff_A_qAgfKp1R4_0(.dout(w_dff_A_d3KWg11b4_0),.din(w_dff_A_qAgfKp1R4_0),.clk(gclk));
	jdff dff_A_d3KWg11b4_0(.dout(w_dff_A_vlL9DLbv4_0),.din(w_dff_A_d3KWg11b4_0),.clk(gclk));
	jdff dff_A_vlL9DLbv4_0(.dout(w_dff_A_mRhjIvPZ4_0),.din(w_dff_A_vlL9DLbv4_0),.clk(gclk));
	jdff dff_A_mRhjIvPZ4_0(.dout(w_dff_A_Bblxg0SQ5_0),.din(w_dff_A_mRhjIvPZ4_0),.clk(gclk));
	jdff dff_A_Bblxg0SQ5_0(.dout(w_dff_A_7wu4IHuK6_0),.din(w_dff_A_Bblxg0SQ5_0),.clk(gclk));
	jdff dff_A_7wu4IHuK6_0(.dout(w_dff_A_rnXu5VpJ8_0),.din(w_dff_A_7wu4IHuK6_0),.clk(gclk));
	jdff dff_A_rnXu5VpJ8_0(.dout(w_dff_A_KWfWl4Vb3_0),.din(w_dff_A_rnXu5VpJ8_0),.clk(gclk));
	jdff dff_A_KWfWl4Vb3_0(.dout(w_dff_A_WIJih7lt7_0),.din(w_dff_A_KWfWl4Vb3_0),.clk(gclk));
	jdff dff_A_WIJih7lt7_0(.dout(w_dff_A_MNG0GSFM8_0),.din(w_dff_A_WIJih7lt7_0),.clk(gclk));
	jdff dff_A_MNG0GSFM8_0(.dout(w_dff_A_Hx307nNz5_0),.din(w_dff_A_MNG0GSFM8_0),.clk(gclk));
	jdff dff_A_Hx307nNz5_0(.dout(w_dff_A_QSNsEGjp8_0),.din(w_dff_A_Hx307nNz5_0),.clk(gclk));
	jdff dff_A_QSNsEGjp8_0(.dout(w_dff_A_IIaFWszV3_0),.din(w_dff_A_QSNsEGjp8_0),.clk(gclk));
	jdff dff_A_IIaFWszV3_0(.dout(w_dff_A_6ljpBP196_0),.din(w_dff_A_IIaFWszV3_0),.clk(gclk));
	jdff dff_A_6ljpBP196_0(.dout(w_dff_A_yzWhyFCM4_0),.din(w_dff_A_6ljpBP196_0),.clk(gclk));
	jdff dff_A_yzWhyFCM4_0(.dout(w_dff_A_79dKQcCA6_0),.din(w_dff_A_yzWhyFCM4_0),.clk(gclk));
	jdff dff_A_79dKQcCA6_0(.dout(w_dff_A_OxNPGvac0_0),.din(w_dff_A_79dKQcCA6_0),.clk(gclk));
	jdff dff_A_OxNPGvac0_0(.dout(w_dff_A_jcMpPvlb7_0),.din(w_dff_A_OxNPGvac0_0),.clk(gclk));
	jdff dff_A_jcMpPvlb7_0(.dout(w_dff_A_FiLwcXha9_0),.din(w_dff_A_jcMpPvlb7_0),.clk(gclk));
	jdff dff_A_FiLwcXha9_0(.dout(w_dff_A_T1zyELv61_0),.din(w_dff_A_FiLwcXha9_0),.clk(gclk));
	jdff dff_A_T1zyELv61_0(.dout(w_dff_A_uwXDEM0t8_0),.din(w_dff_A_T1zyELv61_0),.clk(gclk));
	jdff dff_A_uwXDEM0t8_0(.dout(w_dff_A_WO0q5qOl7_0),.din(w_dff_A_uwXDEM0t8_0),.clk(gclk));
	jdff dff_A_WO0q5qOl7_0(.dout(w_dff_A_fVChj8QF5_0),.din(w_dff_A_WO0q5qOl7_0),.clk(gclk));
	jdff dff_A_fVChj8QF5_0(.dout(w_dff_A_u5lQ2RIG2_0),.din(w_dff_A_fVChj8QF5_0),.clk(gclk));
	jdff dff_A_u5lQ2RIG2_0(.dout(w_dff_A_bMyFap6R8_0),.din(w_dff_A_u5lQ2RIG2_0),.clk(gclk));
	jdff dff_A_bMyFap6R8_0(.dout(w_dff_A_9LJ5SVdU0_0),.din(w_dff_A_bMyFap6R8_0),.clk(gclk));
	jdff dff_A_9LJ5SVdU0_0(.dout(w_dff_A_7SpiseeD3_0),.din(w_dff_A_9LJ5SVdU0_0),.clk(gclk));
	jdff dff_A_7SpiseeD3_0(.dout(w_dff_A_cHyQKoF31_0),.din(w_dff_A_7SpiseeD3_0),.clk(gclk));
	jdff dff_A_cHyQKoF31_0(.dout(w_dff_A_PCqNBvVU8_0),.din(w_dff_A_cHyQKoF31_0),.clk(gclk));
	jdff dff_A_PCqNBvVU8_0(.dout(w_dff_A_UyEANOgG7_0),.din(w_dff_A_PCqNBvVU8_0),.clk(gclk));
	jdff dff_A_UyEANOgG7_0(.dout(w_dff_A_97w0fdhi5_0),.din(w_dff_A_UyEANOgG7_0),.clk(gclk));
	jdff dff_A_97w0fdhi5_0(.dout(w_dff_A_GCTuFQdP2_0),.din(w_dff_A_97w0fdhi5_0),.clk(gclk));
	jdff dff_A_GCTuFQdP2_0(.dout(w_dff_A_8xKbKkRf2_0),.din(w_dff_A_GCTuFQdP2_0),.clk(gclk));
	jdff dff_A_8xKbKkRf2_0(.dout(w_dff_A_GJiTmOg07_0),.din(w_dff_A_8xKbKkRf2_0),.clk(gclk));
	jdff dff_A_GJiTmOg07_0(.dout(w_dff_A_iWyeoXsu8_0),.din(w_dff_A_GJiTmOg07_0),.clk(gclk));
	jdff dff_A_iWyeoXsu8_0(.dout(w_dff_A_vGZPtRr95_0),.din(w_dff_A_iWyeoXsu8_0),.clk(gclk));
	jdff dff_A_vGZPtRr95_0(.dout(w_dff_A_v1wARnUV7_0),.din(w_dff_A_vGZPtRr95_0),.clk(gclk));
	jdff dff_A_v1wARnUV7_0(.dout(w_dff_A_d8ZKm9L55_0),.din(w_dff_A_v1wARnUV7_0),.clk(gclk));
	jdff dff_A_d8ZKm9L55_0(.dout(w_dff_A_uUTRxxwB7_0),.din(w_dff_A_d8ZKm9L55_0),.clk(gclk));
	jdff dff_A_uUTRxxwB7_0(.dout(w_dff_A_1I2yB0dQ3_0),.din(w_dff_A_uUTRxxwB7_0),.clk(gclk));
	jdff dff_A_1I2yB0dQ3_0(.dout(w_dff_A_5tWePsnQ5_0),.din(w_dff_A_1I2yB0dQ3_0),.clk(gclk));
	jdff dff_A_5tWePsnQ5_0(.dout(w_dff_A_QGDy6GMk4_0),.din(w_dff_A_5tWePsnQ5_0),.clk(gclk));
	jdff dff_A_QGDy6GMk4_0(.dout(w_dff_A_WPod74vA5_0),.din(w_dff_A_QGDy6GMk4_0),.clk(gclk));
	jdff dff_A_WPod74vA5_0(.dout(w_dff_A_hZpcWkUB7_0),.din(w_dff_A_WPod74vA5_0),.clk(gclk));
	jdff dff_A_hZpcWkUB7_0(.dout(w_dff_A_G853ioWQ5_0),.din(w_dff_A_hZpcWkUB7_0),.clk(gclk));
	jdff dff_A_G853ioWQ5_0(.dout(G3895gat),.din(w_dff_A_G853ioWQ5_0),.clk(gclk));
	jdff dff_A_mdcJ4ar90_2(.dout(w_dff_A_ucXRuTTy6_0),.din(w_dff_A_mdcJ4ar90_2),.clk(gclk));
	jdff dff_A_ucXRuTTy6_0(.dout(w_dff_A_8wzFp3Rz4_0),.din(w_dff_A_ucXRuTTy6_0),.clk(gclk));
	jdff dff_A_8wzFp3Rz4_0(.dout(w_dff_A_2Q16xPir4_0),.din(w_dff_A_8wzFp3Rz4_0),.clk(gclk));
	jdff dff_A_2Q16xPir4_0(.dout(w_dff_A_RD4HbXrN3_0),.din(w_dff_A_2Q16xPir4_0),.clk(gclk));
	jdff dff_A_RD4HbXrN3_0(.dout(w_dff_A_j0fwaono3_0),.din(w_dff_A_RD4HbXrN3_0),.clk(gclk));
	jdff dff_A_j0fwaono3_0(.dout(w_dff_A_ErXFPDHr2_0),.din(w_dff_A_j0fwaono3_0),.clk(gclk));
	jdff dff_A_ErXFPDHr2_0(.dout(w_dff_A_lNjD4OkO5_0),.din(w_dff_A_ErXFPDHr2_0),.clk(gclk));
	jdff dff_A_lNjD4OkO5_0(.dout(w_dff_A_Ytk9gg1e7_0),.din(w_dff_A_lNjD4OkO5_0),.clk(gclk));
	jdff dff_A_Ytk9gg1e7_0(.dout(w_dff_A_EEAvtlMp8_0),.din(w_dff_A_Ytk9gg1e7_0),.clk(gclk));
	jdff dff_A_EEAvtlMp8_0(.dout(w_dff_A_apc6Yn0R8_0),.din(w_dff_A_EEAvtlMp8_0),.clk(gclk));
	jdff dff_A_apc6Yn0R8_0(.dout(w_dff_A_SDwRpmoh6_0),.din(w_dff_A_apc6Yn0R8_0),.clk(gclk));
	jdff dff_A_SDwRpmoh6_0(.dout(w_dff_A_5rDcnqKM0_0),.din(w_dff_A_SDwRpmoh6_0),.clk(gclk));
	jdff dff_A_5rDcnqKM0_0(.dout(w_dff_A_ewKztJgs5_0),.din(w_dff_A_5rDcnqKM0_0),.clk(gclk));
	jdff dff_A_ewKztJgs5_0(.dout(w_dff_A_TFdvfNZE4_0),.din(w_dff_A_ewKztJgs5_0),.clk(gclk));
	jdff dff_A_TFdvfNZE4_0(.dout(w_dff_A_JMBMXPot0_0),.din(w_dff_A_TFdvfNZE4_0),.clk(gclk));
	jdff dff_A_JMBMXPot0_0(.dout(w_dff_A_FjyxqxJR5_0),.din(w_dff_A_JMBMXPot0_0),.clk(gclk));
	jdff dff_A_FjyxqxJR5_0(.dout(w_dff_A_v1cz1S526_0),.din(w_dff_A_FjyxqxJR5_0),.clk(gclk));
	jdff dff_A_v1cz1S526_0(.dout(w_dff_A_3U3ruLjg7_0),.din(w_dff_A_v1cz1S526_0),.clk(gclk));
	jdff dff_A_3U3ruLjg7_0(.dout(w_dff_A_kdfXz4xG5_0),.din(w_dff_A_3U3ruLjg7_0),.clk(gclk));
	jdff dff_A_kdfXz4xG5_0(.dout(w_dff_A_J6LhkjTI5_0),.din(w_dff_A_kdfXz4xG5_0),.clk(gclk));
	jdff dff_A_J6LhkjTI5_0(.dout(w_dff_A_kkd0xx6G5_0),.din(w_dff_A_J6LhkjTI5_0),.clk(gclk));
	jdff dff_A_kkd0xx6G5_0(.dout(w_dff_A_E2RjHl9D8_0),.din(w_dff_A_kkd0xx6G5_0),.clk(gclk));
	jdff dff_A_E2RjHl9D8_0(.dout(w_dff_A_mPavfK0m8_0),.din(w_dff_A_E2RjHl9D8_0),.clk(gclk));
	jdff dff_A_mPavfK0m8_0(.dout(w_dff_A_C4PI9ZpR7_0),.din(w_dff_A_mPavfK0m8_0),.clk(gclk));
	jdff dff_A_C4PI9ZpR7_0(.dout(w_dff_A_VdZlvEUK6_0),.din(w_dff_A_C4PI9ZpR7_0),.clk(gclk));
	jdff dff_A_VdZlvEUK6_0(.dout(w_dff_A_ZWZPEdqW4_0),.din(w_dff_A_VdZlvEUK6_0),.clk(gclk));
	jdff dff_A_ZWZPEdqW4_0(.dout(w_dff_A_gS7FByvC2_0),.din(w_dff_A_ZWZPEdqW4_0),.clk(gclk));
	jdff dff_A_gS7FByvC2_0(.dout(w_dff_A_EKThDx0b3_0),.din(w_dff_A_gS7FByvC2_0),.clk(gclk));
	jdff dff_A_EKThDx0b3_0(.dout(w_dff_A_zsBQAZrm8_0),.din(w_dff_A_EKThDx0b3_0),.clk(gclk));
	jdff dff_A_zsBQAZrm8_0(.dout(w_dff_A_w6tNTT3C9_0),.din(w_dff_A_zsBQAZrm8_0),.clk(gclk));
	jdff dff_A_w6tNTT3C9_0(.dout(w_dff_A_yfka91WD1_0),.din(w_dff_A_w6tNTT3C9_0),.clk(gclk));
	jdff dff_A_yfka91WD1_0(.dout(w_dff_A_YJElB5c46_0),.din(w_dff_A_yfka91WD1_0),.clk(gclk));
	jdff dff_A_YJElB5c46_0(.dout(w_dff_A_p3iF3YJn8_0),.din(w_dff_A_YJElB5c46_0),.clk(gclk));
	jdff dff_A_p3iF3YJn8_0(.dout(w_dff_A_UFeWtC3S0_0),.din(w_dff_A_p3iF3YJn8_0),.clk(gclk));
	jdff dff_A_UFeWtC3S0_0(.dout(w_dff_A_EsM5A4XG5_0),.din(w_dff_A_UFeWtC3S0_0),.clk(gclk));
	jdff dff_A_EsM5A4XG5_0(.dout(w_dff_A_C06t6JTJ2_0),.din(w_dff_A_EsM5A4XG5_0),.clk(gclk));
	jdff dff_A_C06t6JTJ2_0(.dout(w_dff_A_PAynWK271_0),.din(w_dff_A_C06t6JTJ2_0),.clk(gclk));
	jdff dff_A_PAynWK271_0(.dout(w_dff_A_rIywPZc71_0),.din(w_dff_A_PAynWK271_0),.clk(gclk));
	jdff dff_A_rIywPZc71_0(.dout(w_dff_A_O50fT2260_0),.din(w_dff_A_rIywPZc71_0),.clk(gclk));
	jdff dff_A_O50fT2260_0(.dout(w_dff_A_SjRZRti05_0),.din(w_dff_A_O50fT2260_0),.clk(gclk));
	jdff dff_A_SjRZRti05_0(.dout(w_dff_A_6c2Zg5Hw8_0),.din(w_dff_A_SjRZRti05_0),.clk(gclk));
	jdff dff_A_6c2Zg5Hw8_0(.dout(w_dff_A_qc3faVvK6_0),.din(w_dff_A_6c2Zg5Hw8_0),.clk(gclk));
	jdff dff_A_qc3faVvK6_0(.dout(w_dff_A_d0TPnhfP7_0),.din(w_dff_A_qc3faVvK6_0),.clk(gclk));
	jdff dff_A_d0TPnhfP7_0(.dout(w_dff_A_BCvXb6co5_0),.din(w_dff_A_d0TPnhfP7_0),.clk(gclk));
	jdff dff_A_BCvXb6co5_0(.dout(w_dff_A_kGMURzPc5_0),.din(w_dff_A_BCvXb6co5_0),.clk(gclk));
	jdff dff_A_kGMURzPc5_0(.dout(w_dff_A_TD0rCCw76_0),.din(w_dff_A_kGMURzPc5_0),.clk(gclk));
	jdff dff_A_TD0rCCw76_0(.dout(w_dff_A_UElGlsnx8_0),.din(w_dff_A_TD0rCCw76_0),.clk(gclk));
	jdff dff_A_UElGlsnx8_0(.dout(G4241gat),.din(w_dff_A_UElGlsnx8_0),.clk(gclk));
	jdff dff_A_Phb6U75D9_2(.dout(w_dff_A_mR2Eva228_0),.din(w_dff_A_Phb6U75D9_2),.clk(gclk));
	jdff dff_A_mR2Eva228_0(.dout(w_dff_A_iiBkQspR7_0),.din(w_dff_A_mR2Eva228_0),.clk(gclk));
	jdff dff_A_iiBkQspR7_0(.dout(w_dff_A_q4LRSY5y5_0),.din(w_dff_A_iiBkQspR7_0),.clk(gclk));
	jdff dff_A_q4LRSY5y5_0(.dout(w_dff_A_Y84AA9ZC1_0),.din(w_dff_A_q4LRSY5y5_0),.clk(gclk));
	jdff dff_A_Y84AA9ZC1_0(.dout(w_dff_A_Llfmmfo59_0),.din(w_dff_A_Y84AA9ZC1_0),.clk(gclk));
	jdff dff_A_Llfmmfo59_0(.dout(w_dff_A_DUTLKYQL6_0),.din(w_dff_A_Llfmmfo59_0),.clk(gclk));
	jdff dff_A_DUTLKYQL6_0(.dout(w_dff_A_9aQLkix55_0),.din(w_dff_A_DUTLKYQL6_0),.clk(gclk));
	jdff dff_A_9aQLkix55_0(.dout(w_dff_A_YpfIfAzr6_0),.din(w_dff_A_9aQLkix55_0),.clk(gclk));
	jdff dff_A_YpfIfAzr6_0(.dout(w_dff_A_KNsYc6qM1_0),.din(w_dff_A_YpfIfAzr6_0),.clk(gclk));
	jdff dff_A_KNsYc6qM1_0(.dout(w_dff_A_ngcDbCQN1_0),.din(w_dff_A_KNsYc6qM1_0),.clk(gclk));
	jdff dff_A_ngcDbCQN1_0(.dout(w_dff_A_LUg8UohJ2_0),.din(w_dff_A_ngcDbCQN1_0),.clk(gclk));
	jdff dff_A_LUg8UohJ2_0(.dout(w_dff_A_FB2kpki42_0),.din(w_dff_A_LUg8UohJ2_0),.clk(gclk));
	jdff dff_A_FB2kpki42_0(.dout(w_dff_A_MVtKYeAe9_0),.din(w_dff_A_FB2kpki42_0),.clk(gclk));
	jdff dff_A_MVtKYeAe9_0(.dout(w_dff_A_xEF2irEO8_0),.din(w_dff_A_MVtKYeAe9_0),.clk(gclk));
	jdff dff_A_xEF2irEO8_0(.dout(w_dff_A_nGGdf9zh1_0),.din(w_dff_A_xEF2irEO8_0),.clk(gclk));
	jdff dff_A_nGGdf9zh1_0(.dout(w_dff_A_cTZlejHs1_0),.din(w_dff_A_nGGdf9zh1_0),.clk(gclk));
	jdff dff_A_cTZlejHs1_0(.dout(w_dff_A_0JAzP6X92_0),.din(w_dff_A_cTZlejHs1_0),.clk(gclk));
	jdff dff_A_0JAzP6X92_0(.dout(w_dff_A_TShY5e1Z7_0),.din(w_dff_A_0JAzP6X92_0),.clk(gclk));
	jdff dff_A_TShY5e1Z7_0(.dout(w_dff_A_Vy2WT7NC9_0),.din(w_dff_A_TShY5e1Z7_0),.clk(gclk));
	jdff dff_A_Vy2WT7NC9_0(.dout(w_dff_A_0de3tUVL0_0),.din(w_dff_A_Vy2WT7NC9_0),.clk(gclk));
	jdff dff_A_0de3tUVL0_0(.dout(w_dff_A_GpRypKlf2_0),.din(w_dff_A_0de3tUVL0_0),.clk(gclk));
	jdff dff_A_GpRypKlf2_0(.dout(w_dff_A_iuQwrsgM3_0),.din(w_dff_A_GpRypKlf2_0),.clk(gclk));
	jdff dff_A_iuQwrsgM3_0(.dout(w_dff_A_PZD3Cajo7_0),.din(w_dff_A_iuQwrsgM3_0),.clk(gclk));
	jdff dff_A_PZD3Cajo7_0(.dout(w_dff_A_EPf5hEiT1_0),.din(w_dff_A_PZD3Cajo7_0),.clk(gclk));
	jdff dff_A_EPf5hEiT1_0(.dout(w_dff_A_GoxV6nt89_0),.din(w_dff_A_EPf5hEiT1_0),.clk(gclk));
	jdff dff_A_GoxV6nt89_0(.dout(w_dff_A_hE0m3T3e9_0),.din(w_dff_A_GoxV6nt89_0),.clk(gclk));
	jdff dff_A_hE0m3T3e9_0(.dout(w_dff_A_3tX2e9C44_0),.din(w_dff_A_hE0m3T3e9_0),.clk(gclk));
	jdff dff_A_3tX2e9C44_0(.dout(w_dff_A_jNyxx1wT6_0),.din(w_dff_A_3tX2e9C44_0),.clk(gclk));
	jdff dff_A_jNyxx1wT6_0(.dout(w_dff_A_QJEE8DWm4_0),.din(w_dff_A_jNyxx1wT6_0),.clk(gclk));
	jdff dff_A_QJEE8DWm4_0(.dout(w_dff_A_PuXQpVOz3_0),.din(w_dff_A_QJEE8DWm4_0),.clk(gclk));
	jdff dff_A_PuXQpVOz3_0(.dout(w_dff_A_7XI49bBE6_0),.din(w_dff_A_PuXQpVOz3_0),.clk(gclk));
	jdff dff_A_7XI49bBE6_0(.dout(w_dff_A_6XOZBCHi0_0),.din(w_dff_A_7XI49bBE6_0),.clk(gclk));
	jdff dff_A_6XOZBCHi0_0(.dout(w_dff_A_85U7jzTf1_0),.din(w_dff_A_6XOZBCHi0_0),.clk(gclk));
	jdff dff_A_85U7jzTf1_0(.dout(w_dff_A_MnTObEKb6_0),.din(w_dff_A_85U7jzTf1_0),.clk(gclk));
	jdff dff_A_MnTObEKb6_0(.dout(w_dff_A_o8iwBowI6_0),.din(w_dff_A_MnTObEKb6_0),.clk(gclk));
	jdff dff_A_o8iwBowI6_0(.dout(w_dff_A_nhjQHZwh3_0),.din(w_dff_A_o8iwBowI6_0),.clk(gclk));
	jdff dff_A_nhjQHZwh3_0(.dout(w_dff_A_Oa3dy7Jx0_0),.din(w_dff_A_nhjQHZwh3_0),.clk(gclk));
	jdff dff_A_Oa3dy7Jx0_0(.dout(w_dff_A_moRygh1K1_0),.din(w_dff_A_Oa3dy7Jx0_0),.clk(gclk));
	jdff dff_A_moRygh1K1_0(.dout(w_dff_A_J86AyhRy1_0),.din(w_dff_A_moRygh1K1_0),.clk(gclk));
	jdff dff_A_J86AyhRy1_0(.dout(w_dff_A_zsMZny7A9_0),.din(w_dff_A_J86AyhRy1_0),.clk(gclk));
	jdff dff_A_zsMZny7A9_0(.dout(w_dff_A_9jyakfJn9_0),.din(w_dff_A_zsMZny7A9_0),.clk(gclk));
	jdff dff_A_9jyakfJn9_0(.dout(w_dff_A_YmCBS2ot5_0),.din(w_dff_A_9jyakfJn9_0),.clk(gclk));
	jdff dff_A_YmCBS2ot5_0(.dout(w_dff_A_vsJcTJdJ4_0),.din(w_dff_A_YmCBS2ot5_0),.clk(gclk));
	jdff dff_A_vsJcTJdJ4_0(.dout(w_dff_A_H8sTOo013_0),.din(w_dff_A_vsJcTJdJ4_0),.clk(gclk));
	jdff dff_A_H8sTOo013_0(.dout(G4591gat),.din(w_dff_A_H8sTOo013_0),.clk(gclk));
	jdff dff_A_x2APV6JE4_2(.dout(w_dff_A_4ZUMfstK2_0),.din(w_dff_A_x2APV6JE4_2),.clk(gclk));
	jdff dff_A_4ZUMfstK2_0(.dout(w_dff_A_8isAp7KB2_0),.din(w_dff_A_4ZUMfstK2_0),.clk(gclk));
	jdff dff_A_8isAp7KB2_0(.dout(w_dff_A_4Z7Lme3u0_0),.din(w_dff_A_8isAp7KB2_0),.clk(gclk));
	jdff dff_A_4Z7Lme3u0_0(.dout(w_dff_A_bXFsMF1j7_0),.din(w_dff_A_4Z7Lme3u0_0),.clk(gclk));
	jdff dff_A_bXFsMF1j7_0(.dout(w_dff_A_4IEEwk6D1_0),.din(w_dff_A_bXFsMF1j7_0),.clk(gclk));
	jdff dff_A_4IEEwk6D1_0(.dout(w_dff_A_m8vhnz8X6_0),.din(w_dff_A_4IEEwk6D1_0),.clk(gclk));
	jdff dff_A_m8vhnz8X6_0(.dout(w_dff_A_HYP6mTaq8_0),.din(w_dff_A_m8vhnz8X6_0),.clk(gclk));
	jdff dff_A_HYP6mTaq8_0(.dout(w_dff_A_u2lVkaxh5_0),.din(w_dff_A_HYP6mTaq8_0),.clk(gclk));
	jdff dff_A_u2lVkaxh5_0(.dout(w_dff_A_AdqfIWAB0_0),.din(w_dff_A_u2lVkaxh5_0),.clk(gclk));
	jdff dff_A_AdqfIWAB0_0(.dout(w_dff_A_EWuIz2Yi1_0),.din(w_dff_A_AdqfIWAB0_0),.clk(gclk));
	jdff dff_A_EWuIz2Yi1_0(.dout(w_dff_A_2kzbZG6l7_0),.din(w_dff_A_EWuIz2Yi1_0),.clk(gclk));
	jdff dff_A_2kzbZG6l7_0(.dout(w_dff_A_DeGW5AQc1_0),.din(w_dff_A_2kzbZG6l7_0),.clk(gclk));
	jdff dff_A_DeGW5AQc1_0(.dout(w_dff_A_NiH8YMgt1_0),.din(w_dff_A_DeGW5AQc1_0),.clk(gclk));
	jdff dff_A_NiH8YMgt1_0(.dout(w_dff_A_CnZPTTrA1_0),.din(w_dff_A_NiH8YMgt1_0),.clk(gclk));
	jdff dff_A_CnZPTTrA1_0(.dout(w_dff_A_BNP7UCab2_0),.din(w_dff_A_CnZPTTrA1_0),.clk(gclk));
	jdff dff_A_BNP7UCab2_0(.dout(w_dff_A_KvAm47Gq4_0),.din(w_dff_A_BNP7UCab2_0),.clk(gclk));
	jdff dff_A_KvAm47Gq4_0(.dout(w_dff_A_bMRb5fEI9_0),.din(w_dff_A_KvAm47Gq4_0),.clk(gclk));
	jdff dff_A_bMRb5fEI9_0(.dout(w_dff_A_HBs1nnTQ8_0),.din(w_dff_A_bMRb5fEI9_0),.clk(gclk));
	jdff dff_A_HBs1nnTQ8_0(.dout(w_dff_A_AxWT3cyQ6_0),.din(w_dff_A_HBs1nnTQ8_0),.clk(gclk));
	jdff dff_A_AxWT3cyQ6_0(.dout(w_dff_A_0yEshw0C5_0),.din(w_dff_A_AxWT3cyQ6_0),.clk(gclk));
	jdff dff_A_0yEshw0C5_0(.dout(w_dff_A_hgW0cZ6R3_0),.din(w_dff_A_0yEshw0C5_0),.clk(gclk));
	jdff dff_A_hgW0cZ6R3_0(.dout(w_dff_A_1FU2AFeo8_0),.din(w_dff_A_hgW0cZ6R3_0),.clk(gclk));
	jdff dff_A_1FU2AFeo8_0(.dout(w_dff_A_38nBbQo59_0),.din(w_dff_A_1FU2AFeo8_0),.clk(gclk));
	jdff dff_A_38nBbQo59_0(.dout(w_dff_A_TxihdmPS3_0),.din(w_dff_A_38nBbQo59_0),.clk(gclk));
	jdff dff_A_TxihdmPS3_0(.dout(w_dff_A_PhBFujKQ8_0),.din(w_dff_A_TxihdmPS3_0),.clk(gclk));
	jdff dff_A_PhBFujKQ8_0(.dout(w_dff_A_5R1Urcqo2_0),.din(w_dff_A_PhBFujKQ8_0),.clk(gclk));
	jdff dff_A_5R1Urcqo2_0(.dout(w_dff_A_PlGwnbl21_0),.din(w_dff_A_5R1Urcqo2_0),.clk(gclk));
	jdff dff_A_PlGwnbl21_0(.dout(w_dff_A_9dQXlluI7_0),.din(w_dff_A_PlGwnbl21_0),.clk(gclk));
	jdff dff_A_9dQXlluI7_0(.dout(w_dff_A_2Bc3iSTU2_0),.din(w_dff_A_9dQXlluI7_0),.clk(gclk));
	jdff dff_A_2Bc3iSTU2_0(.dout(w_dff_A_2GQKVBUa4_0),.din(w_dff_A_2Bc3iSTU2_0),.clk(gclk));
	jdff dff_A_2GQKVBUa4_0(.dout(w_dff_A_9BaNkW873_0),.din(w_dff_A_2GQKVBUa4_0),.clk(gclk));
	jdff dff_A_9BaNkW873_0(.dout(w_dff_A_YKM56Nk35_0),.din(w_dff_A_9BaNkW873_0),.clk(gclk));
	jdff dff_A_YKM56Nk35_0(.dout(w_dff_A_iMAxdH4P7_0),.din(w_dff_A_YKM56Nk35_0),.clk(gclk));
	jdff dff_A_iMAxdH4P7_0(.dout(w_dff_A_BMI7anqQ5_0),.din(w_dff_A_iMAxdH4P7_0),.clk(gclk));
	jdff dff_A_BMI7anqQ5_0(.dout(w_dff_A_kVagMUbd2_0),.din(w_dff_A_BMI7anqQ5_0),.clk(gclk));
	jdff dff_A_kVagMUbd2_0(.dout(w_dff_A_bc52apDh2_0),.din(w_dff_A_kVagMUbd2_0),.clk(gclk));
	jdff dff_A_bc52apDh2_0(.dout(w_dff_A_dRqHU3vM2_0),.din(w_dff_A_bc52apDh2_0),.clk(gclk));
	jdff dff_A_dRqHU3vM2_0(.dout(w_dff_A_jBG6z9Zz6_0),.din(w_dff_A_dRqHU3vM2_0),.clk(gclk));
	jdff dff_A_jBG6z9Zz6_0(.dout(w_dff_A_HbMaSnJb1_0),.din(w_dff_A_jBG6z9Zz6_0),.clk(gclk));
	jdff dff_A_HbMaSnJb1_0(.dout(w_dff_A_sGerDx5E0_0),.din(w_dff_A_HbMaSnJb1_0),.clk(gclk));
	jdff dff_A_sGerDx5E0_0(.dout(w_dff_A_xgDN7rc03_0),.din(w_dff_A_sGerDx5E0_0),.clk(gclk));
	jdff dff_A_xgDN7rc03_0(.dout(G4946gat),.din(w_dff_A_xgDN7rc03_0),.clk(gclk));
	jdff dff_A_7vyaZLbT9_2(.dout(w_dff_A_rBGM1luv2_0),.din(w_dff_A_7vyaZLbT9_2),.clk(gclk));
	jdff dff_A_rBGM1luv2_0(.dout(w_dff_A_lSs1vlGz9_0),.din(w_dff_A_rBGM1luv2_0),.clk(gclk));
	jdff dff_A_lSs1vlGz9_0(.dout(w_dff_A_96qz8p685_0),.din(w_dff_A_lSs1vlGz9_0),.clk(gclk));
	jdff dff_A_96qz8p685_0(.dout(w_dff_A_gxl8MQ4C1_0),.din(w_dff_A_96qz8p685_0),.clk(gclk));
	jdff dff_A_gxl8MQ4C1_0(.dout(w_dff_A_6Zc0b0fZ8_0),.din(w_dff_A_gxl8MQ4C1_0),.clk(gclk));
	jdff dff_A_6Zc0b0fZ8_0(.dout(w_dff_A_UKQhSSBv1_0),.din(w_dff_A_6Zc0b0fZ8_0),.clk(gclk));
	jdff dff_A_UKQhSSBv1_0(.dout(w_dff_A_0Uc7yspJ2_0),.din(w_dff_A_UKQhSSBv1_0),.clk(gclk));
	jdff dff_A_0Uc7yspJ2_0(.dout(w_dff_A_p2BWwzJt9_0),.din(w_dff_A_0Uc7yspJ2_0),.clk(gclk));
	jdff dff_A_p2BWwzJt9_0(.dout(w_dff_A_jgqmBM7u3_0),.din(w_dff_A_p2BWwzJt9_0),.clk(gclk));
	jdff dff_A_jgqmBM7u3_0(.dout(w_dff_A_TC6LzhCv1_0),.din(w_dff_A_jgqmBM7u3_0),.clk(gclk));
	jdff dff_A_TC6LzhCv1_0(.dout(w_dff_A_lWMirraW9_0),.din(w_dff_A_TC6LzhCv1_0),.clk(gclk));
	jdff dff_A_lWMirraW9_0(.dout(w_dff_A_2fBCdJA41_0),.din(w_dff_A_lWMirraW9_0),.clk(gclk));
	jdff dff_A_2fBCdJA41_0(.dout(w_dff_A_AgMpUUJg0_0),.din(w_dff_A_2fBCdJA41_0),.clk(gclk));
	jdff dff_A_AgMpUUJg0_0(.dout(w_dff_A_qFMdeTVf4_0),.din(w_dff_A_AgMpUUJg0_0),.clk(gclk));
	jdff dff_A_qFMdeTVf4_0(.dout(w_dff_A_LMHMNP2S0_0),.din(w_dff_A_qFMdeTVf4_0),.clk(gclk));
	jdff dff_A_LMHMNP2S0_0(.dout(w_dff_A_My7pE2MQ1_0),.din(w_dff_A_LMHMNP2S0_0),.clk(gclk));
	jdff dff_A_My7pE2MQ1_0(.dout(w_dff_A_18ITMQEf6_0),.din(w_dff_A_My7pE2MQ1_0),.clk(gclk));
	jdff dff_A_18ITMQEf6_0(.dout(w_dff_A_AUUizrVk3_0),.din(w_dff_A_18ITMQEf6_0),.clk(gclk));
	jdff dff_A_AUUizrVk3_0(.dout(w_dff_A_cEGfUJgl3_0),.din(w_dff_A_AUUizrVk3_0),.clk(gclk));
	jdff dff_A_cEGfUJgl3_0(.dout(w_dff_A_oJXbKlhp9_0),.din(w_dff_A_cEGfUJgl3_0),.clk(gclk));
	jdff dff_A_oJXbKlhp9_0(.dout(w_dff_A_R70apvjg6_0),.din(w_dff_A_oJXbKlhp9_0),.clk(gclk));
	jdff dff_A_R70apvjg6_0(.dout(w_dff_A_hxDU4T4v5_0),.din(w_dff_A_R70apvjg6_0),.clk(gclk));
	jdff dff_A_hxDU4T4v5_0(.dout(w_dff_A_y09MRX6l3_0),.din(w_dff_A_hxDU4T4v5_0),.clk(gclk));
	jdff dff_A_y09MRX6l3_0(.dout(w_dff_A_TUn1Bpxd1_0),.din(w_dff_A_y09MRX6l3_0),.clk(gclk));
	jdff dff_A_TUn1Bpxd1_0(.dout(w_dff_A_xDZBgepc1_0),.din(w_dff_A_TUn1Bpxd1_0),.clk(gclk));
	jdff dff_A_xDZBgepc1_0(.dout(w_dff_A_Avkw0D2G0_0),.din(w_dff_A_xDZBgepc1_0),.clk(gclk));
	jdff dff_A_Avkw0D2G0_0(.dout(w_dff_A_3yAZ8lbo1_0),.din(w_dff_A_Avkw0D2G0_0),.clk(gclk));
	jdff dff_A_3yAZ8lbo1_0(.dout(w_dff_A_Vb4wSG9j9_0),.din(w_dff_A_3yAZ8lbo1_0),.clk(gclk));
	jdff dff_A_Vb4wSG9j9_0(.dout(w_dff_A_Yh73tfam1_0),.din(w_dff_A_Vb4wSG9j9_0),.clk(gclk));
	jdff dff_A_Yh73tfam1_0(.dout(w_dff_A_vROip8wM3_0),.din(w_dff_A_Yh73tfam1_0),.clk(gclk));
	jdff dff_A_vROip8wM3_0(.dout(w_dff_A_u3M4koVj4_0),.din(w_dff_A_vROip8wM3_0),.clk(gclk));
	jdff dff_A_u3M4koVj4_0(.dout(w_dff_A_1OqLBf1z9_0),.din(w_dff_A_u3M4koVj4_0),.clk(gclk));
	jdff dff_A_1OqLBf1z9_0(.dout(w_dff_A_wjoisF5K4_0),.din(w_dff_A_1OqLBf1z9_0),.clk(gclk));
	jdff dff_A_wjoisF5K4_0(.dout(w_dff_A_6Sybiw3c3_0),.din(w_dff_A_wjoisF5K4_0),.clk(gclk));
	jdff dff_A_6Sybiw3c3_0(.dout(w_dff_A_2AMhb9GJ6_0),.din(w_dff_A_6Sybiw3c3_0),.clk(gclk));
	jdff dff_A_2AMhb9GJ6_0(.dout(w_dff_A_xvKm44JZ0_0),.din(w_dff_A_2AMhb9GJ6_0),.clk(gclk));
	jdff dff_A_xvKm44JZ0_0(.dout(w_dff_A_LQ7uLL3z4_0),.din(w_dff_A_xvKm44JZ0_0),.clk(gclk));
	jdff dff_A_LQ7uLL3z4_0(.dout(w_dff_A_SCqH8zVk4_0),.din(w_dff_A_LQ7uLL3z4_0),.clk(gclk));
	jdff dff_A_SCqH8zVk4_0(.dout(G5308gat),.din(w_dff_A_SCqH8zVk4_0),.clk(gclk));
	jdff dff_A_TEKx8qT56_2(.dout(w_dff_A_5mbaOIAJ7_0),.din(w_dff_A_TEKx8qT56_2),.clk(gclk));
	jdff dff_A_5mbaOIAJ7_0(.dout(w_dff_A_EeD76MjA9_0),.din(w_dff_A_5mbaOIAJ7_0),.clk(gclk));
	jdff dff_A_EeD76MjA9_0(.dout(w_dff_A_LEiV6ZbY0_0),.din(w_dff_A_EeD76MjA9_0),.clk(gclk));
	jdff dff_A_LEiV6ZbY0_0(.dout(w_dff_A_k3IAA0DQ1_0),.din(w_dff_A_LEiV6ZbY0_0),.clk(gclk));
	jdff dff_A_k3IAA0DQ1_0(.dout(w_dff_A_hUJ43Mx16_0),.din(w_dff_A_k3IAA0DQ1_0),.clk(gclk));
	jdff dff_A_hUJ43Mx16_0(.dout(w_dff_A_9IUh5jR18_0),.din(w_dff_A_hUJ43Mx16_0),.clk(gclk));
	jdff dff_A_9IUh5jR18_0(.dout(w_dff_A_AhKosuqg5_0),.din(w_dff_A_9IUh5jR18_0),.clk(gclk));
	jdff dff_A_AhKosuqg5_0(.dout(w_dff_A_LPRA2KEJ1_0),.din(w_dff_A_AhKosuqg5_0),.clk(gclk));
	jdff dff_A_LPRA2KEJ1_0(.dout(w_dff_A_2RppvQGd1_0),.din(w_dff_A_LPRA2KEJ1_0),.clk(gclk));
	jdff dff_A_2RppvQGd1_0(.dout(w_dff_A_hhlbElyG8_0),.din(w_dff_A_2RppvQGd1_0),.clk(gclk));
	jdff dff_A_hhlbElyG8_0(.dout(w_dff_A_uzU0o8xR2_0),.din(w_dff_A_hhlbElyG8_0),.clk(gclk));
	jdff dff_A_uzU0o8xR2_0(.dout(w_dff_A_UINZN4gY4_0),.din(w_dff_A_uzU0o8xR2_0),.clk(gclk));
	jdff dff_A_UINZN4gY4_0(.dout(w_dff_A_8cLKzRYr0_0),.din(w_dff_A_UINZN4gY4_0),.clk(gclk));
	jdff dff_A_8cLKzRYr0_0(.dout(w_dff_A_vKxdlqmx2_0),.din(w_dff_A_8cLKzRYr0_0),.clk(gclk));
	jdff dff_A_vKxdlqmx2_0(.dout(w_dff_A_gqh9o9Uh4_0),.din(w_dff_A_vKxdlqmx2_0),.clk(gclk));
	jdff dff_A_gqh9o9Uh4_0(.dout(w_dff_A_24sZSyuT2_0),.din(w_dff_A_gqh9o9Uh4_0),.clk(gclk));
	jdff dff_A_24sZSyuT2_0(.dout(w_dff_A_NqdZPWQn1_0),.din(w_dff_A_24sZSyuT2_0),.clk(gclk));
	jdff dff_A_NqdZPWQn1_0(.dout(w_dff_A_AiBYpJBN9_0),.din(w_dff_A_NqdZPWQn1_0),.clk(gclk));
	jdff dff_A_AiBYpJBN9_0(.dout(w_dff_A_D50d9q789_0),.din(w_dff_A_AiBYpJBN9_0),.clk(gclk));
	jdff dff_A_D50d9q789_0(.dout(w_dff_A_ac4B31Zm5_0),.din(w_dff_A_D50d9q789_0),.clk(gclk));
	jdff dff_A_ac4B31Zm5_0(.dout(w_dff_A_s2yProDA8_0),.din(w_dff_A_ac4B31Zm5_0),.clk(gclk));
	jdff dff_A_s2yProDA8_0(.dout(w_dff_A_brPQUTpK2_0),.din(w_dff_A_s2yProDA8_0),.clk(gclk));
	jdff dff_A_brPQUTpK2_0(.dout(w_dff_A_0XnJtovy0_0),.din(w_dff_A_brPQUTpK2_0),.clk(gclk));
	jdff dff_A_0XnJtovy0_0(.dout(w_dff_A_lsm4iIuD7_0),.din(w_dff_A_0XnJtovy0_0),.clk(gclk));
	jdff dff_A_lsm4iIuD7_0(.dout(w_dff_A_F6jGdstK4_0),.din(w_dff_A_lsm4iIuD7_0),.clk(gclk));
	jdff dff_A_F6jGdstK4_0(.dout(w_dff_A_SVNBHzQj6_0),.din(w_dff_A_F6jGdstK4_0),.clk(gclk));
	jdff dff_A_SVNBHzQj6_0(.dout(w_dff_A_kBXQzIa09_0),.din(w_dff_A_SVNBHzQj6_0),.clk(gclk));
	jdff dff_A_kBXQzIa09_0(.dout(w_dff_A_r43YaIL49_0),.din(w_dff_A_kBXQzIa09_0),.clk(gclk));
	jdff dff_A_r43YaIL49_0(.dout(w_dff_A_Ltom9Con4_0),.din(w_dff_A_r43YaIL49_0),.clk(gclk));
	jdff dff_A_Ltom9Con4_0(.dout(w_dff_A_raTQam683_0),.din(w_dff_A_Ltom9Con4_0),.clk(gclk));
	jdff dff_A_raTQam683_0(.dout(w_dff_A_TiehvIPe1_0),.din(w_dff_A_raTQam683_0),.clk(gclk));
	jdff dff_A_TiehvIPe1_0(.dout(w_dff_A_Vx8PwlVK2_0),.din(w_dff_A_TiehvIPe1_0),.clk(gclk));
	jdff dff_A_Vx8PwlVK2_0(.dout(w_dff_A_lBGpUiJc3_0),.din(w_dff_A_Vx8PwlVK2_0),.clk(gclk));
	jdff dff_A_lBGpUiJc3_0(.dout(w_dff_A_ezVCfewI6_0),.din(w_dff_A_lBGpUiJc3_0),.clk(gclk));
	jdff dff_A_ezVCfewI6_0(.dout(w_dff_A_miMC25NO6_0),.din(w_dff_A_ezVCfewI6_0),.clk(gclk));
	jdff dff_A_miMC25NO6_0(.dout(G5672gat),.din(w_dff_A_miMC25NO6_0),.clk(gclk));
	jdff dff_A_ND5rrPHV5_2(.dout(w_dff_A_rnAfQz647_0),.din(w_dff_A_ND5rrPHV5_2),.clk(gclk));
	jdff dff_A_rnAfQz647_0(.dout(w_dff_A_ZoFID5zg1_0),.din(w_dff_A_rnAfQz647_0),.clk(gclk));
	jdff dff_A_ZoFID5zg1_0(.dout(w_dff_A_noM0juy98_0),.din(w_dff_A_ZoFID5zg1_0),.clk(gclk));
	jdff dff_A_noM0juy98_0(.dout(w_dff_A_UD61nGIn5_0),.din(w_dff_A_noM0juy98_0),.clk(gclk));
	jdff dff_A_UD61nGIn5_0(.dout(w_dff_A_dCcWln6m4_0),.din(w_dff_A_UD61nGIn5_0),.clk(gclk));
	jdff dff_A_dCcWln6m4_0(.dout(w_dff_A_iSE9KQJO4_0),.din(w_dff_A_dCcWln6m4_0),.clk(gclk));
	jdff dff_A_iSE9KQJO4_0(.dout(w_dff_A_6luKBhuP9_0),.din(w_dff_A_iSE9KQJO4_0),.clk(gclk));
	jdff dff_A_6luKBhuP9_0(.dout(w_dff_A_uNvo4nFD0_0),.din(w_dff_A_6luKBhuP9_0),.clk(gclk));
	jdff dff_A_uNvo4nFD0_0(.dout(w_dff_A_64uUHRJo8_0),.din(w_dff_A_uNvo4nFD0_0),.clk(gclk));
	jdff dff_A_64uUHRJo8_0(.dout(w_dff_A_DlEzE1mQ8_0),.din(w_dff_A_64uUHRJo8_0),.clk(gclk));
	jdff dff_A_DlEzE1mQ8_0(.dout(w_dff_A_4oxaVBo92_0),.din(w_dff_A_DlEzE1mQ8_0),.clk(gclk));
	jdff dff_A_4oxaVBo92_0(.dout(w_dff_A_a6yGjMhT8_0),.din(w_dff_A_4oxaVBo92_0),.clk(gclk));
	jdff dff_A_a6yGjMhT8_0(.dout(w_dff_A_3vS5ofQE4_0),.din(w_dff_A_a6yGjMhT8_0),.clk(gclk));
	jdff dff_A_3vS5ofQE4_0(.dout(w_dff_A_uO5GxKNN4_0),.din(w_dff_A_3vS5ofQE4_0),.clk(gclk));
	jdff dff_A_uO5GxKNN4_0(.dout(w_dff_A_QGzY2HHp8_0),.din(w_dff_A_uO5GxKNN4_0),.clk(gclk));
	jdff dff_A_QGzY2HHp8_0(.dout(w_dff_A_ctOe0XbO7_0),.din(w_dff_A_QGzY2HHp8_0),.clk(gclk));
	jdff dff_A_ctOe0XbO7_0(.dout(w_dff_A_seMU5cwB7_0),.din(w_dff_A_ctOe0XbO7_0),.clk(gclk));
	jdff dff_A_seMU5cwB7_0(.dout(w_dff_A_fJ2ksThq7_0),.din(w_dff_A_seMU5cwB7_0),.clk(gclk));
	jdff dff_A_fJ2ksThq7_0(.dout(w_dff_A_kNbLuFPy1_0),.din(w_dff_A_fJ2ksThq7_0),.clk(gclk));
	jdff dff_A_kNbLuFPy1_0(.dout(w_dff_A_tDwSXBuX8_0),.din(w_dff_A_kNbLuFPy1_0),.clk(gclk));
	jdff dff_A_tDwSXBuX8_0(.dout(w_dff_A_TkTttgAE7_0),.din(w_dff_A_tDwSXBuX8_0),.clk(gclk));
	jdff dff_A_TkTttgAE7_0(.dout(w_dff_A_1MceHRts7_0),.din(w_dff_A_TkTttgAE7_0),.clk(gclk));
	jdff dff_A_1MceHRts7_0(.dout(w_dff_A_6ri971VA8_0),.din(w_dff_A_1MceHRts7_0),.clk(gclk));
	jdff dff_A_6ri971VA8_0(.dout(w_dff_A_KIrgp2FT9_0),.din(w_dff_A_6ri971VA8_0),.clk(gclk));
	jdff dff_A_KIrgp2FT9_0(.dout(w_dff_A_FxLDEICg3_0),.din(w_dff_A_KIrgp2FT9_0),.clk(gclk));
	jdff dff_A_FxLDEICg3_0(.dout(w_dff_A_Q7ZELAT24_0),.din(w_dff_A_FxLDEICg3_0),.clk(gclk));
	jdff dff_A_Q7ZELAT24_0(.dout(w_dff_A_49v8goCE1_0),.din(w_dff_A_Q7ZELAT24_0),.clk(gclk));
	jdff dff_A_49v8goCE1_0(.dout(w_dff_A_hBHHZSBk0_0),.din(w_dff_A_49v8goCE1_0),.clk(gclk));
	jdff dff_A_hBHHZSBk0_0(.dout(w_dff_A_yhb5xtMo9_0),.din(w_dff_A_hBHHZSBk0_0),.clk(gclk));
	jdff dff_A_yhb5xtMo9_0(.dout(w_dff_A_fD7qzMXK6_0),.din(w_dff_A_yhb5xtMo9_0),.clk(gclk));
	jdff dff_A_fD7qzMXK6_0(.dout(w_dff_A_BwrTxgv56_0),.din(w_dff_A_fD7qzMXK6_0),.clk(gclk));
	jdff dff_A_BwrTxgv56_0(.dout(w_dff_A_7zApRyyX4_0),.din(w_dff_A_BwrTxgv56_0),.clk(gclk));
	jdff dff_A_7zApRyyX4_0(.dout(G5971gat),.din(w_dff_A_7zApRyyX4_0),.clk(gclk));
	jdff dff_A_NtHJwKOW4_2(.dout(w_dff_A_tTAugpDu8_0),.din(w_dff_A_NtHJwKOW4_2),.clk(gclk));
	jdff dff_A_tTAugpDu8_0(.dout(w_dff_A_YArGBafw5_0),.din(w_dff_A_tTAugpDu8_0),.clk(gclk));
	jdff dff_A_YArGBafw5_0(.dout(w_dff_A_WFPPUgIw0_0),.din(w_dff_A_YArGBafw5_0),.clk(gclk));
	jdff dff_A_WFPPUgIw0_0(.dout(w_dff_A_13jcXOoq3_0),.din(w_dff_A_WFPPUgIw0_0),.clk(gclk));
	jdff dff_A_13jcXOoq3_0(.dout(w_dff_A_CkGOUhHZ3_0),.din(w_dff_A_13jcXOoq3_0),.clk(gclk));
	jdff dff_A_CkGOUhHZ3_0(.dout(w_dff_A_xiSZTgnd1_0),.din(w_dff_A_CkGOUhHZ3_0),.clk(gclk));
	jdff dff_A_xiSZTgnd1_0(.dout(w_dff_A_XaxNQUaZ9_0),.din(w_dff_A_xiSZTgnd1_0),.clk(gclk));
	jdff dff_A_XaxNQUaZ9_0(.dout(w_dff_A_sxEwDzW34_0),.din(w_dff_A_XaxNQUaZ9_0),.clk(gclk));
	jdff dff_A_sxEwDzW34_0(.dout(w_dff_A_aWMd9Avm2_0),.din(w_dff_A_sxEwDzW34_0),.clk(gclk));
	jdff dff_A_aWMd9Avm2_0(.dout(w_dff_A_IjeC78Q92_0),.din(w_dff_A_aWMd9Avm2_0),.clk(gclk));
	jdff dff_A_IjeC78Q92_0(.dout(w_dff_A_ExpXmqPP2_0),.din(w_dff_A_IjeC78Q92_0),.clk(gclk));
	jdff dff_A_ExpXmqPP2_0(.dout(w_dff_A_ChGizsMB3_0),.din(w_dff_A_ExpXmqPP2_0),.clk(gclk));
	jdff dff_A_ChGizsMB3_0(.dout(w_dff_A_jMGqfSc36_0),.din(w_dff_A_ChGizsMB3_0),.clk(gclk));
	jdff dff_A_jMGqfSc36_0(.dout(w_dff_A_4c4B0fIt5_0),.din(w_dff_A_jMGqfSc36_0),.clk(gclk));
	jdff dff_A_4c4B0fIt5_0(.dout(w_dff_A_O2DG3k1q4_0),.din(w_dff_A_4c4B0fIt5_0),.clk(gclk));
	jdff dff_A_O2DG3k1q4_0(.dout(w_dff_A_eUEtAQCo4_0),.din(w_dff_A_O2DG3k1q4_0),.clk(gclk));
	jdff dff_A_eUEtAQCo4_0(.dout(w_dff_A_4bLZjiLN2_0),.din(w_dff_A_eUEtAQCo4_0),.clk(gclk));
	jdff dff_A_4bLZjiLN2_0(.dout(w_dff_A_wBb23zsF9_0),.din(w_dff_A_4bLZjiLN2_0),.clk(gclk));
	jdff dff_A_wBb23zsF9_0(.dout(w_dff_A_Mo48ahrG7_0),.din(w_dff_A_wBb23zsF9_0),.clk(gclk));
	jdff dff_A_Mo48ahrG7_0(.dout(w_dff_A_4uVDk40k9_0),.din(w_dff_A_Mo48ahrG7_0),.clk(gclk));
	jdff dff_A_4uVDk40k9_0(.dout(w_dff_A_QPJq0wl87_0),.din(w_dff_A_4uVDk40k9_0),.clk(gclk));
	jdff dff_A_QPJq0wl87_0(.dout(w_dff_A_RIzwbEFv3_0),.din(w_dff_A_QPJq0wl87_0),.clk(gclk));
	jdff dff_A_RIzwbEFv3_0(.dout(w_dff_A_wW8DdkE31_0),.din(w_dff_A_RIzwbEFv3_0),.clk(gclk));
	jdff dff_A_wW8DdkE31_0(.dout(w_dff_A_G9Hukp1N3_0),.din(w_dff_A_wW8DdkE31_0),.clk(gclk));
	jdff dff_A_G9Hukp1N3_0(.dout(w_dff_A_RqIx8HCk4_0),.din(w_dff_A_G9Hukp1N3_0),.clk(gclk));
	jdff dff_A_RqIx8HCk4_0(.dout(w_dff_A_ALOEaoHQ2_0),.din(w_dff_A_RqIx8HCk4_0),.clk(gclk));
	jdff dff_A_ALOEaoHQ2_0(.dout(w_dff_A_UG3LSBeI9_0),.din(w_dff_A_ALOEaoHQ2_0),.clk(gclk));
	jdff dff_A_UG3LSBeI9_0(.dout(w_dff_A_slTLL1i85_0),.din(w_dff_A_UG3LSBeI9_0),.clk(gclk));
	jdff dff_A_slTLL1i85_0(.dout(w_dff_A_fvjl21Pj0_0),.din(w_dff_A_slTLL1i85_0),.clk(gclk));
	jdff dff_A_fvjl21Pj0_0(.dout(G6123gat),.din(w_dff_A_fvjl21Pj0_0),.clk(gclk));
	jdff dff_A_GkoBMSiy7_2(.dout(w_dff_A_dFa2grTs5_0),.din(w_dff_A_GkoBMSiy7_2),.clk(gclk));
	jdff dff_A_dFa2grTs5_0(.dout(w_dff_A_gJhzoAqT4_0),.din(w_dff_A_dFa2grTs5_0),.clk(gclk));
	jdff dff_A_gJhzoAqT4_0(.dout(w_dff_A_wzQDPlfJ8_0),.din(w_dff_A_gJhzoAqT4_0),.clk(gclk));
	jdff dff_A_wzQDPlfJ8_0(.dout(w_dff_A_79cZBL3i4_0),.din(w_dff_A_wzQDPlfJ8_0),.clk(gclk));
	jdff dff_A_79cZBL3i4_0(.dout(w_dff_A_2pjyHanq4_0),.din(w_dff_A_79cZBL3i4_0),.clk(gclk));
	jdff dff_A_2pjyHanq4_0(.dout(w_dff_A_OSRhVY1y6_0),.din(w_dff_A_2pjyHanq4_0),.clk(gclk));
	jdff dff_A_OSRhVY1y6_0(.dout(w_dff_A_zwZK5P7g3_0),.din(w_dff_A_OSRhVY1y6_0),.clk(gclk));
	jdff dff_A_zwZK5P7g3_0(.dout(w_dff_A_ELBK5l5c3_0),.din(w_dff_A_zwZK5P7g3_0),.clk(gclk));
	jdff dff_A_ELBK5l5c3_0(.dout(w_dff_A_v22zptni0_0),.din(w_dff_A_ELBK5l5c3_0),.clk(gclk));
	jdff dff_A_v22zptni0_0(.dout(w_dff_A_p3wQVyqS2_0),.din(w_dff_A_v22zptni0_0),.clk(gclk));
	jdff dff_A_p3wQVyqS2_0(.dout(w_dff_A_YVwbXvNp5_0),.din(w_dff_A_p3wQVyqS2_0),.clk(gclk));
	jdff dff_A_YVwbXvNp5_0(.dout(w_dff_A_vSa1ery42_0),.din(w_dff_A_YVwbXvNp5_0),.clk(gclk));
	jdff dff_A_vSa1ery42_0(.dout(w_dff_A_gp0tKW2z2_0),.din(w_dff_A_vSa1ery42_0),.clk(gclk));
	jdff dff_A_gp0tKW2z2_0(.dout(w_dff_A_w2Cxhf6o2_0),.din(w_dff_A_gp0tKW2z2_0),.clk(gclk));
	jdff dff_A_w2Cxhf6o2_0(.dout(w_dff_A_q04g2wjQ5_0),.din(w_dff_A_w2Cxhf6o2_0),.clk(gclk));
	jdff dff_A_q04g2wjQ5_0(.dout(w_dff_A_8ywlq8QD5_0),.din(w_dff_A_q04g2wjQ5_0),.clk(gclk));
	jdff dff_A_8ywlq8QD5_0(.dout(w_dff_A_Po2kMWjL0_0),.din(w_dff_A_8ywlq8QD5_0),.clk(gclk));
	jdff dff_A_Po2kMWjL0_0(.dout(w_dff_A_BZaa3w2n4_0),.din(w_dff_A_Po2kMWjL0_0),.clk(gclk));
	jdff dff_A_BZaa3w2n4_0(.dout(w_dff_A_6tTqPnQr9_0),.din(w_dff_A_BZaa3w2n4_0),.clk(gclk));
	jdff dff_A_6tTqPnQr9_0(.dout(w_dff_A_1gZyF6l89_0),.din(w_dff_A_6tTqPnQr9_0),.clk(gclk));
	jdff dff_A_1gZyF6l89_0(.dout(w_dff_A_mjBcYgBA6_0),.din(w_dff_A_1gZyF6l89_0),.clk(gclk));
	jdff dff_A_mjBcYgBA6_0(.dout(w_dff_A_c2YqTHKU9_0),.din(w_dff_A_mjBcYgBA6_0),.clk(gclk));
	jdff dff_A_c2YqTHKU9_0(.dout(w_dff_A_Mig4cTnu4_0),.din(w_dff_A_c2YqTHKU9_0),.clk(gclk));
	jdff dff_A_Mig4cTnu4_0(.dout(w_dff_A_2l8yetws1_0),.din(w_dff_A_Mig4cTnu4_0),.clk(gclk));
	jdff dff_A_2l8yetws1_0(.dout(w_dff_A_Y7CuQ6JA8_0),.din(w_dff_A_2l8yetws1_0),.clk(gclk));
	jdff dff_A_Y7CuQ6JA8_0(.dout(w_dff_A_kQnOLAU39_0),.din(w_dff_A_Y7CuQ6JA8_0),.clk(gclk));
	jdff dff_A_kQnOLAU39_0(.dout(w_dff_A_5SPcpRbO5_0),.din(w_dff_A_kQnOLAU39_0),.clk(gclk));
	jdff dff_A_5SPcpRbO5_0(.dout(G6150gat),.din(w_dff_A_5SPcpRbO5_0),.clk(gclk));
	jdff dff_A_fgq1tWlH0_2(.dout(w_dff_A_FMBJe05O9_0),.din(w_dff_A_fgq1tWlH0_2),.clk(gclk));
	jdff dff_A_FMBJe05O9_0(.dout(w_dff_A_4CLg10dh8_0),.din(w_dff_A_FMBJe05O9_0),.clk(gclk));
	jdff dff_A_4CLg10dh8_0(.dout(w_dff_A_LVL9bFe91_0),.din(w_dff_A_4CLg10dh8_0),.clk(gclk));
	jdff dff_A_LVL9bFe91_0(.dout(w_dff_A_oppvS8j14_0),.din(w_dff_A_LVL9bFe91_0),.clk(gclk));
	jdff dff_A_oppvS8j14_0(.dout(w_dff_A_OSQHFrAg1_0),.din(w_dff_A_oppvS8j14_0),.clk(gclk));
	jdff dff_A_OSQHFrAg1_0(.dout(w_dff_A_ryMO8kaz0_0),.din(w_dff_A_OSQHFrAg1_0),.clk(gclk));
	jdff dff_A_ryMO8kaz0_0(.dout(w_dff_A_rYofgzWO9_0),.din(w_dff_A_ryMO8kaz0_0),.clk(gclk));
	jdff dff_A_rYofgzWO9_0(.dout(w_dff_A_mBkmDaAr7_0),.din(w_dff_A_rYofgzWO9_0),.clk(gclk));
	jdff dff_A_mBkmDaAr7_0(.dout(w_dff_A_oYaKYWwJ3_0),.din(w_dff_A_mBkmDaAr7_0),.clk(gclk));
	jdff dff_A_oYaKYWwJ3_0(.dout(w_dff_A_NEEFFIV93_0),.din(w_dff_A_oYaKYWwJ3_0),.clk(gclk));
	jdff dff_A_NEEFFIV93_0(.dout(w_dff_A_NKLITBXP5_0),.din(w_dff_A_NEEFFIV93_0),.clk(gclk));
	jdff dff_A_NKLITBXP5_0(.dout(w_dff_A_KiciQbBH1_0),.din(w_dff_A_NKLITBXP5_0),.clk(gclk));
	jdff dff_A_KiciQbBH1_0(.dout(w_dff_A_tCRfYsDX5_0),.din(w_dff_A_KiciQbBH1_0),.clk(gclk));
	jdff dff_A_tCRfYsDX5_0(.dout(w_dff_A_XyVUbH8F1_0),.din(w_dff_A_tCRfYsDX5_0),.clk(gclk));
	jdff dff_A_XyVUbH8F1_0(.dout(w_dff_A_diXooZ1c8_0),.din(w_dff_A_XyVUbH8F1_0),.clk(gclk));
	jdff dff_A_diXooZ1c8_0(.dout(w_dff_A_JYl2zW550_0),.din(w_dff_A_diXooZ1c8_0),.clk(gclk));
	jdff dff_A_JYl2zW550_0(.dout(w_dff_A_ChMB0Ynx5_0),.din(w_dff_A_JYl2zW550_0),.clk(gclk));
	jdff dff_A_ChMB0Ynx5_0(.dout(w_dff_A_tLXdZOYV8_0),.din(w_dff_A_ChMB0Ynx5_0),.clk(gclk));
	jdff dff_A_tLXdZOYV8_0(.dout(w_dff_A_aPx83fBB0_0),.din(w_dff_A_tLXdZOYV8_0),.clk(gclk));
	jdff dff_A_aPx83fBB0_0(.dout(w_dff_A_kiSBccT21_0),.din(w_dff_A_aPx83fBB0_0),.clk(gclk));
	jdff dff_A_kiSBccT21_0(.dout(w_dff_A_9aIz1G115_0),.din(w_dff_A_kiSBccT21_0),.clk(gclk));
	jdff dff_A_9aIz1G115_0(.dout(w_dff_A_VrkgbPSv9_0),.din(w_dff_A_9aIz1G115_0),.clk(gclk));
	jdff dff_A_VrkgbPSv9_0(.dout(w_dff_A_VvnvkjsB7_0),.din(w_dff_A_VrkgbPSv9_0),.clk(gclk));
	jdff dff_A_VvnvkjsB7_0(.dout(w_dff_A_bPuLvC5u3_0),.din(w_dff_A_VvnvkjsB7_0),.clk(gclk));
	jdff dff_A_bPuLvC5u3_0(.dout(w_dff_A_K0VMRFxq2_0),.din(w_dff_A_bPuLvC5u3_0),.clk(gclk));
	jdff dff_A_K0VMRFxq2_0(.dout(G6160gat),.din(w_dff_A_K0VMRFxq2_0),.clk(gclk));
	jdff dff_A_obuUdNIl2_2(.dout(w_dff_A_3LVBNeEx3_0),.din(w_dff_A_obuUdNIl2_2),.clk(gclk));
	jdff dff_A_3LVBNeEx3_0(.dout(w_dff_A_Xouw1Ph47_0),.din(w_dff_A_3LVBNeEx3_0),.clk(gclk));
	jdff dff_A_Xouw1Ph47_0(.dout(w_dff_A_wX4PHBXr0_0),.din(w_dff_A_Xouw1Ph47_0),.clk(gclk));
	jdff dff_A_wX4PHBXr0_0(.dout(w_dff_A_uzrl6ITp3_0),.din(w_dff_A_wX4PHBXr0_0),.clk(gclk));
	jdff dff_A_uzrl6ITp3_0(.dout(w_dff_A_RbZnFsIQ5_0),.din(w_dff_A_uzrl6ITp3_0),.clk(gclk));
	jdff dff_A_RbZnFsIQ5_0(.dout(w_dff_A_DggnEZFj7_0),.din(w_dff_A_RbZnFsIQ5_0),.clk(gclk));
	jdff dff_A_DggnEZFj7_0(.dout(w_dff_A_PFmNnG3k8_0),.din(w_dff_A_DggnEZFj7_0),.clk(gclk));
	jdff dff_A_PFmNnG3k8_0(.dout(w_dff_A_K9dQJapv8_0),.din(w_dff_A_PFmNnG3k8_0),.clk(gclk));
	jdff dff_A_K9dQJapv8_0(.dout(w_dff_A_jYnAtpYq3_0),.din(w_dff_A_K9dQJapv8_0),.clk(gclk));
	jdff dff_A_jYnAtpYq3_0(.dout(w_dff_A_ISuhW5kz7_0),.din(w_dff_A_jYnAtpYq3_0),.clk(gclk));
	jdff dff_A_ISuhW5kz7_0(.dout(w_dff_A_j8rDyhVM4_0),.din(w_dff_A_ISuhW5kz7_0),.clk(gclk));
	jdff dff_A_j8rDyhVM4_0(.dout(w_dff_A_ofAzioCB2_0),.din(w_dff_A_j8rDyhVM4_0),.clk(gclk));
	jdff dff_A_ofAzioCB2_0(.dout(w_dff_A_tbZj41kF9_0),.din(w_dff_A_ofAzioCB2_0),.clk(gclk));
	jdff dff_A_tbZj41kF9_0(.dout(w_dff_A_vlDewE9B9_0),.din(w_dff_A_tbZj41kF9_0),.clk(gclk));
	jdff dff_A_vlDewE9B9_0(.dout(w_dff_A_ZPeyBSXX7_0),.din(w_dff_A_vlDewE9B9_0),.clk(gclk));
	jdff dff_A_ZPeyBSXX7_0(.dout(w_dff_A_wK1dcayQ8_0),.din(w_dff_A_ZPeyBSXX7_0),.clk(gclk));
	jdff dff_A_wK1dcayQ8_0(.dout(w_dff_A_WEVIotbk2_0),.din(w_dff_A_wK1dcayQ8_0),.clk(gclk));
	jdff dff_A_WEVIotbk2_0(.dout(w_dff_A_oIOw8cGC7_0),.din(w_dff_A_WEVIotbk2_0),.clk(gclk));
	jdff dff_A_oIOw8cGC7_0(.dout(w_dff_A_HvckR75J2_0),.din(w_dff_A_oIOw8cGC7_0),.clk(gclk));
	jdff dff_A_HvckR75J2_0(.dout(w_dff_A_LwNB3OKs1_0),.din(w_dff_A_HvckR75J2_0),.clk(gclk));
	jdff dff_A_LwNB3OKs1_0(.dout(w_dff_A_kFu9MVUT3_0),.din(w_dff_A_LwNB3OKs1_0),.clk(gclk));
	jdff dff_A_kFu9MVUT3_0(.dout(w_dff_A_gM8cknpP4_0),.din(w_dff_A_kFu9MVUT3_0),.clk(gclk));
	jdff dff_A_gM8cknpP4_0(.dout(w_dff_A_ytUpiMlJ5_0),.din(w_dff_A_gM8cknpP4_0),.clk(gclk));
	jdff dff_A_ytUpiMlJ5_0(.dout(w_dff_A_wJ6PBTgs4_0),.din(w_dff_A_ytUpiMlJ5_0),.clk(gclk));
	jdff dff_A_wJ6PBTgs4_0(.dout(G6170gat),.din(w_dff_A_wJ6PBTgs4_0),.clk(gclk));
	jdff dff_A_XYc3sDAs5_2(.dout(w_dff_A_s8Lz3PP21_0),.din(w_dff_A_XYc3sDAs5_2),.clk(gclk));
	jdff dff_A_s8Lz3PP21_0(.dout(w_dff_A_Vl6XXqKR4_0),.din(w_dff_A_s8Lz3PP21_0),.clk(gclk));
	jdff dff_A_Vl6XXqKR4_0(.dout(w_dff_A_mIRvBGgs2_0),.din(w_dff_A_Vl6XXqKR4_0),.clk(gclk));
	jdff dff_A_mIRvBGgs2_0(.dout(w_dff_A_j61eup6U3_0),.din(w_dff_A_mIRvBGgs2_0),.clk(gclk));
	jdff dff_A_j61eup6U3_0(.dout(w_dff_A_XzSjgAJD4_0),.din(w_dff_A_j61eup6U3_0),.clk(gclk));
	jdff dff_A_XzSjgAJD4_0(.dout(w_dff_A_qN60RfzG1_0),.din(w_dff_A_XzSjgAJD4_0),.clk(gclk));
	jdff dff_A_qN60RfzG1_0(.dout(w_dff_A_gc57QrSY6_0),.din(w_dff_A_qN60RfzG1_0),.clk(gclk));
	jdff dff_A_gc57QrSY6_0(.dout(w_dff_A_l0SLvcbN7_0),.din(w_dff_A_gc57QrSY6_0),.clk(gclk));
	jdff dff_A_l0SLvcbN7_0(.dout(w_dff_A_DrbsFgqW9_0),.din(w_dff_A_l0SLvcbN7_0),.clk(gclk));
	jdff dff_A_DrbsFgqW9_0(.dout(w_dff_A_N4255XaA4_0),.din(w_dff_A_DrbsFgqW9_0),.clk(gclk));
	jdff dff_A_N4255XaA4_0(.dout(w_dff_A_9t9c2ZSL7_0),.din(w_dff_A_N4255XaA4_0),.clk(gclk));
	jdff dff_A_9t9c2ZSL7_0(.dout(w_dff_A_TwcTavwt2_0),.din(w_dff_A_9t9c2ZSL7_0),.clk(gclk));
	jdff dff_A_TwcTavwt2_0(.dout(w_dff_A_gGj8T90x1_0),.din(w_dff_A_TwcTavwt2_0),.clk(gclk));
	jdff dff_A_gGj8T90x1_0(.dout(w_dff_A_gSEeBq5e7_0),.din(w_dff_A_gGj8T90x1_0),.clk(gclk));
	jdff dff_A_gSEeBq5e7_0(.dout(w_dff_A_LYPqDeu10_0),.din(w_dff_A_gSEeBq5e7_0),.clk(gclk));
	jdff dff_A_LYPqDeu10_0(.dout(w_dff_A_Eo0iLPBH0_0),.din(w_dff_A_LYPqDeu10_0),.clk(gclk));
	jdff dff_A_Eo0iLPBH0_0(.dout(w_dff_A_IulUPpmL5_0),.din(w_dff_A_Eo0iLPBH0_0),.clk(gclk));
	jdff dff_A_IulUPpmL5_0(.dout(w_dff_A_qHkWz9bX2_0),.din(w_dff_A_IulUPpmL5_0),.clk(gclk));
	jdff dff_A_qHkWz9bX2_0(.dout(w_dff_A_FdyIXHAm7_0),.din(w_dff_A_qHkWz9bX2_0),.clk(gclk));
	jdff dff_A_FdyIXHAm7_0(.dout(w_dff_A_WwhykUhZ0_0),.din(w_dff_A_FdyIXHAm7_0),.clk(gclk));
	jdff dff_A_WwhykUhZ0_0(.dout(w_dff_A_2s2nWD7l1_0),.din(w_dff_A_WwhykUhZ0_0),.clk(gclk));
	jdff dff_A_2s2nWD7l1_0(.dout(w_dff_A_jIx7cOiV7_0),.din(w_dff_A_2s2nWD7l1_0),.clk(gclk));
	jdff dff_A_jIx7cOiV7_0(.dout(G6180gat),.din(w_dff_A_jIx7cOiV7_0),.clk(gclk));
	jdff dff_A_0iZHqm6h1_2(.dout(w_dff_A_prtqAZc98_0),.din(w_dff_A_0iZHqm6h1_2),.clk(gclk));
	jdff dff_A_prtqAZc98_0(.dout(w_dff_A_YziWlVof8_0),.din(w_dff_A_prtqAZc98_0),.clk(gclk));
	jdff dff_A_YziWlVof8_0(.dout(w_dff_A_UiZcUW5a0_0),.din(w_dff_A_YziWlVof8_0),.clk(gclk));
	jdff dff_A_UiZcUW5a0_0(.dout(w_dff_A_W2hvF0zz0_0),.din(w_dff_A_UiZcUW5a0_0),.clk(gclk));
	jdff dff_A_W2hvF0zz0_0(.dout(w_dff_A_xjdaaH8o2_0),.din(w_dff_A_W2hvF0zz0_0),.clk(gclk));
	jdff dff_A_xjdaaH8o2_0(.dout(w_dff_A_UfmbiT5a1_0),.din(w_dff_A_xjdaaH8o2_0),.clk(gclk));
	jdff dff_A_UfmbiT5a1_0(.dout(w_dff_A_dWzIwmUM7_0),.din(w_dff_A_UfmbiT5a1_0),.clk(gclk));
	jdff dff_A_dWzIwmUM7_0(.dout(w_dff_A_138kPFry8_0),.din(w_dff_A_dWzIwmUM7_0),.clk(gclk));
	jdff dff_A_138kPFry8_0(.dout(w_dff_A_gTtrjauN9_0),.din(w_dff_A_138kPFry8_0),.clk(gclk));
	jdff dff_A_gTtrjauN9_0(.dout(w_dff_A_bLdR2FXj9_0),.din(w_dff_A_gTtrjauN9_0),.clk(gclk));
	jdff dff_A_bLdR2FXj9_0(.dout(w_dff_A_W7qz9fsH8_0),.din(w_dff_A_bLdR2FXj9_0),.clk(gclk));
	jdff dff_A_W7qz9fsH8_0(.dout(w_dff_A_CaEvomZQ3_0),.din(w_dff_A_W7qz9fsH8_0),.clk(gclk));
	jdff dff_A_CaEvomZQ3_0(.dout(w_dff_A_mHVkNbvH7_0),.din(w_dff_A_CaEvomZQ3_0),.clk(gclk));
	jdff dff_A_mHVkNbvH7_0(.dout(w_dff_A_kJMyCwVs3_0),.din(w_dff_A_mHVkNbvH7_0),.clk(gclk));
	jdff dff_A_kJMyCwVs3_0(.dout(w_dff_A_8jUGBtcG2_0),.din(w_dff_A_kJMyCwVs3_0),.clk(gclk));
	jdff dff_A_8jUGBtcG2_0(.dout(w_dff_A_bOQ97r6R4_0),.din(w_dff_A_8jUGBtcG2_0),.clk(gclk));
	jdff dff_A_bOQ97r6R4_0(.dout(w_dff_A_T6qWt4nx7_0),.din(w_dff_A_bOQ97r6R4_0),.clk(gclk));
	jdff dff_A_T6qWt4nx7_0(.dout(w_dff_A_ixdpxXyl9_0),.din(w_dff_A_T6qWt4nx7_0),.clk(gclk));
	jdff dff_A_ixdpxXyl9_0(.dout(w_dff_A_QDexrUex8_0),.din(w_dff_A_ixdpxXyl9_0),.clk(gclk));
	jdff dff_A_QDexrUex8_0(.dout(w_dff_A_4Tot9Ke45_0),.din(w_dff_A_QDexrUex8_0),.clk(gclk));
	jdff dff_A_4Tot9Ke45_0(.dout(G6190gat),.din(w_dff_A_4Tot9Ke45_0),.clk(gclk));
	jdff dff_A_DbIDePej4_2(.dout(w_dff_A_mGau4jRS5_0),.din(w_dff_A_DbIDePej4_2),.clk(gclk));
	jdff dff_A_mGau4jRS5_0(.dout(w_dff_A_aQIhDYMB0_0),.din(w_dff_A_mGau4jRS5_0),.clk(gclk));
	jdff dff_A_aQIhDYMB0_0(.dout(w_dff_A_QVEmwyc12_0),.din(w_dff_A_aQIhDYMB0_0),.clk(gclk));
	jdff dff_A_QVEmwyc12_0(.dout(w_dff_A_1vdIsrcS5_0),.din(w_dff_A_QVEmwyc12_0),.clk(gclk));
	jdff dff_A_1vdIsrcS5_0(.dout(w_dff_A_nUyTD8ts3_0),.din(w_dff_A_1vdIsrcS5_0),.clk(gclk));
	jdff dff_A_nUyTD8ts3_0(.dout(w_dff_A_u2jthr0Z6_0),.din(w_dff_A_nUyTD8ts3_0),.clk(gclk));
	jdff dff_A_u2jthr0Z6_0(.dout(w_dff_A_qQ7jFv5L9_0),.din(w_dff_A_u2jthr0Z6_0),.clk(gclk));
	jdff dff_A_qQ7jFv5L9_0(.dout(w_dff_A_4KyxBQfF9_0),.din(w_dff_A_qQ7jFv5L9_0),.clk(gclk));
	jdff dff_A_4KyxBQfF9_0(.dout(w_dff_A_pzlp7gQm8_0),.din(w_dff_A_4KyxBQfF9_0),.clk(gclk));
	jdff dff_A_pzlp7gQm8_0(.dout(w_dff_A_gQCbsAhm6_0),.din(w_dff_A_pzlp7gQm8_0),.clk(gclk));
	jdff dff_A_gQCbsAhm6_0(.dout(w_dff_A_oTcZHgAl7_0),.din(w_dff_A_gQCbsAhm6_0),.clk(gclk));
	jdff dff_A_oTcZHgAl7_0(.dout(w_dff_A_Tfh6mXU79_0),.din(w_dff_A_oTcZHgAl7_0),.clk(gclk));
	jdff dff_A_Tfh6mXU79_0(.dout(w_dff_A_RiKmipjv3_0),.din(w_dff_A_Tfh6mXU79_0),.clk(gclk));
	jdff dff_A_RiKmipjv3_0(.dout(w_dff_A_JSEHANbP2_0),.din(w_dff_A_RiKmipjv3_0),.clk(gclk));
	jdff dff_A_JSEHANbP2_0(.dout(w_dff_A_OS4F2H9T4_0),.din(w_dff_A_JSEHANbP2_0),.clk(gclk));
	jdff dff_A_OS4F2H9T4_0(.dout(w_dff_A_nNDroKgT3_0),.din(w_dff_A_OS4F2H9T4_0),.clk(gclk));
	jdff dff_A_nNDroKgT3_0(.dout(w_dff_A_ryZ5pVjc1_0),.din(w_dff_A_nNDroKgT3_0),.clk(gclk));
	jdff dff_A_ryZ5pVjc1_0(.dout(w_dff_A_CwF0X3Qt5_0),.din(w_dff_A_ryZ5pVjc1_0),.clk(gclk));
	jdff dff_A_CwF0X3Qt5_0(.dout(G6200gat),.din(w_dff_A_CwF0X3Qt5_0),.clk(gclk));
	jdff dff_A_IUYnNff39_2(.dout(w_dff_A_xQeTjuds5_0),.din(w_dff_A_IUYnNff39_2),.clk(gclk));
	jdff dff_A_xQeTjuds5_0(.dout(w_dff_A_U1EP0ICI1_0),.din(w_dff_A_xQeTjuds5_0),.clk(gclk));
	jdff dff_A_U1EP0ICI1_0(.dout(w_dff_A_XPescyqL8_0),.din(w_dff_A_U1EP0ICI1_0),.clk(gclk));
	jdff dff_A_XPescyqL8_0(.dout(w_dff_A_6lpCmimB2_0),.din(w_dff_A_XPescyqL8_0),.clk(gclk));
	jdff dff_A_6lpCmimB2_0(.dout(w_dff_A_vYYr7qNX5_0),.din(w_dff_A_6lpCmimB2_0),.clk(gclk));
	jdff dff_A_vYYr7qNX5_0(.dout(w_dff_A_taIrpx5f3_0),.din(w_dff_A_vYYr7qNX5_0),.clk(gclk));
	jdff dff_A_taIrpx5f3_0(.dout(w_dff_A_xU2xglG99_0),.din(w_dff_A_taIrpx5f3_0),.clk(gclk));
	jdff dff_A_xU2xglG99_0(.dout(w_dff_A_fr2ZZxGV7_0),.din(w_dff_A_xU2xglG99_0),.clk(gclk));
	jdff dff_A_fr2ZZxGV7_0(.dout(w_dff_A_Yq6pLs3I3_0),.din(w_dff_A_fr2ZZxGV7_0),.clk(gclk));
	jdff dff_A_Yq6pLs3I3_0(.dout(w_dff_A_KxfVw64E6_0),.din(w_dff_A_Yq6pLs3I3_0),.clk(gclk));
	jdff dff_A_KxfVw64E6_0(.dout(w_dff_A_uTlf0yaM5_0),.din(w_dff_A_KxfVw64E6_0),.clk(gclk));
	jdff dff_A_uTlf0yaM5_0(.dout(w_dff_A_b9Imky7T9_0),.din(w_dff_A_uTlf0yaM5_0),.clk(gclk));
	jdff dff_A_b9Imky7T9_0(.dout(w_dff_A_ngYzzIIk4_0),.din(w_dff_A_b9Imky7T9_0),.clk(gclk));
	jdff dff_A_ngYzzIIk4_0(.dout(w_dff_A_LHDF6mO28_0),.din(w_dff_A_ngYzzIIk4_0),.clk(gclk));
	jdff dff_A_LHDF6mO28_0(.dout(w_dff_A_Wqx6ig220_0),.din(w_dff_A_LHDF6mO28_0),.clk(gclk));
	jdff dff_A_Wqx6ig220_0(.dout(w_dff_A_q0ovqedw9_0),.din(w_dff_A_Wqx6ig220_0),.clk(gclk));
	jdff dff_A_q0ovqedw9_0(.dout(G6210gat),.din(w_dff_A_q0ovqedw9_0),.clk(gclk));
	jdff dff_A_bLrqy25k9_2(.dout(w_dff_A_Zvp8zY511_0),.din(w_dff_A_bLrqy25k9_2),.clk(gclk));
	jdff dff_A_Zvp8zY511_0(.dout(w_dff_A_3phXYowu3_0),.din(w_dff_A_Zvp8zY511_0),.clk(gclk));
	jdff dff_A_3phXYowu3_0(.dout(w_dff_A_93feg0hY2_0),.din(w_dff_A_3phXYowu3_0),.clk(gclk));
	jdff dff_A_93feg0hY2_0(.dout(w_dff_A_h9JzAGb39_0),.din(w_dff_A_93feg0hY2_0),.clk(gclk));
	jdff dff_A_h9JzAGb39_0(.dout(w_dff_A_EvwOX0nf7_0),.din(w_dff_A_h9JzAGb39_0),.clk(gclk));
	jdff dff_A_EvwOX0nf7_0(.dout(w_dff_A_csAyt3t46_0),.din(w_dff_A_EvwOX0nf7_0),.clk(gclk));
	jdff dff_A_csAyt3t46_0(.dout(w_dff_A_XiOyo2uX4_0),.din(w_dff_A_csAyt3t46_0),.clk(gclk));
	jdff dff_A_XiOyo2uX4_0(.dout(w_dff_A_p3fTEORF6_0),.din(w_dff_A_XiOyo2uX4_0),.clk(gclk));
	jdff dff_A_p3fTEORF6_0(.dout(w_dff_A_TNemDBlJ5_0),.din(w_dff_A_p3fTEORF6_0),.clk(gclk));
	jdff dff_A_TNemDBlJ5_0(.dout(w_dff_A_AidrJimb7_0),.din(w_dff_A_TNemDBlJ5_0),.clk(gclk));
	jdff dff_A_AidrJimb7_0(.dout(w_dff_A_zvqnxQ0t7_0),.din(w_dff_A_AidrJimb7_0),.clk(gclk));
	jdff dff_A_zvqnxQ0t7_0(.dout(w_dff_A_ReOMoYRg9_0),.din(w_dff_A_zvqnxQ0t7_0),.clk(gclk));
	jdff dff_A_ReOMoYRg9_0(.dout(w_dff_A_FhgJ3KMa0_0),.din(w_dff_A_ReOMoYRg9_0),.clk(gclk));
	jdff dff_A_FhgJ3KMa0_0(.dout(w_dff_A_zFU6cqn04_0),.din(w_dff_A_FhgJ3KMa0_0),.clk(gclk));
	jdff dff_A_zFU6cqn04_0(.dout(G6220gat),.din(w_dff_A_zFU6cqn04_0),.clk(gclk));
	jdff dff_A_LmfDc3mX7_2(.dout(w_dff_A_hboK2Rm15_0),.din(w_dff_A_LmfDc3mX7_2),.clk(gclk));
	jdff dff_A_hboK2Rm15_0(.dout(w_dff_A_At2BKpWp7_0),.din(w_dff_A_hboK2Rm15_0),.clk(gclk));
	jdff dff_A_At2BKpWp7_0(.dout(w_dff_A_QV3e7I3m6_0),.din(w_dff_A_At2BKpWp7_0),.clk(gclk));
	jdff dff_A_QV3e7I3m6_0(.dout(w_dff_A_CltQHqxN1_0),.din(w_dff_A_QV3e7I3m6_0),.clk(gclk));
	jdff dff_A_CltQHqxN1_0(.dout(w_dff_A_EP4Nrif76_0),.din(w_dff_A_CltQHqxN1_0),.clk(gclk));
	jdff dff_A_EP4Nrif76_0(.dout(w_dff_A_EDFDqcWu2_0),.din(w_dff_A_EP4Nrif76_0),.clk(gclk));
	jdff dff_A_EDFDqcWu2_0(.dout(w_dff_A_C9lOJ36M2_0),.din(w_dff_A_EDFDqcWu2_0),.clk(gclk));
	jdff dff_A_C9lOJ36M2_0(.dout(w_dff_A_KMCrbG5i2_0),.din(w_dff_A_C9lOJ36M2_0),.clk(gclk));
	jdff dff_A_KMCrbG5i2_0(.dout(w_dff_A_B1mpiYQK7_0),.din(w_dff_A_KMCrbG5i2_0),.clk(gclk));
	jdff dff_A_B1mpiYQK7_0(.dout(w_dff_A_VxSjdbXL3_0),.din(w_dff_A_B1mpiYQK7_0),.clk(gclk));
	jdff dff_A_VxSjdbXL3_0(.dout(w_dff_A_jemr7PEt7_0),.din(w_dff_A_VxSjdbXL3_0),.clk(gclk));
	jdff dff_A_jemr7PEt7_0(.dout(w_dff_A_tVYZQ0xk2_0),.din(w_dff_A_jemr7PEt7_0),.clk(gclk));
	jdff dff_A_tVYZQ0xk2_0(.dout(G6230gat),.din(w_dff_A_tVYZQ0xk2_0),.clk(gclk));
	jdff dff_A_hXEXHGJP4_2(.dout(w_dff_A_Jd6PsPPu4_0),.din(w_dff_A_hXEXHGJP4_2),.clk(gclk));
	jdff dff_A_Jd6PsPPu4_0(.dout(w_dff_A_JL78wWS26_0),.din(w_dff_A_Jd6PsPPu4_0),.clk(gclk));
	jdff dff_A_JL78wWS26_0(.dout(w_dff_A_BovAFiDd6_0),.din(w_dff_A_JL78wWS26_0),.clk(gclk));
	jdff dff_A_BovAFiDd6_0(.dout(w_dff_A_S33jOICy7_0),.din(w_dff_A_BovAFiDd6_0),.clk(gclk));
	jdff dff_A_S33jOICy7_0(.dout(w_dff_A_LK6wRUxT8_0),.din(w_dff_A_S33jOICy7_0),.clk(gclk));
	jdff dff_A_LK6wRUxT8_0(.dout(w_dff_A_dMe4vE8R8_0),.din(w_dff_A_LK6wRUxT8_0),.clk(gclk));
	jdff dff_A_dMe4vE8R8_0(.dout(w_dff_A_PFx33hNw4_0),.din(w_dff_A_dMe4vE8R8_0),.clk(gclk));
	jdff dff_A_PFx33hNw4_0(.dout(w_dff_A_fwuPYOIa2_0),.din(w_dff_A_PFx33hNw4_0),.clk(gclk));
	jdff dff_A_fwuPYOIa2_0(.dout(w_dff_A_O5HVrv8X7_0),.din(w_dff_A_fwuPYOIa2_0),.clk(gclk));
	jdff dff_A_O5HVrv8X7_0(.dout(w_dff_A_v64lkwQT4_0),.din(w_dff_A_O5HVrv8X7_0),.clk(gclk));
	jdff dff_A_v64lkwQT4_0(.dout(G6240gat),.din(w_dff_A_v64lkwQT4_0),.clk(gclk));
	jdff dff_A_3iLVSEwm9_2(.dout(w_dff_A_4W1dVK516_0),.din(w_dff_A_3iLVSEwm9_2),.clk(gclk));
	jdff dff_A_4W1dVK516_0(.dout(w_dff_A_NaxIzPxG7_0),.din(w_dff_A_4W1dVK516_0),.clk(gclk));
	jdff dff_A_NaxIzPxG7_0(.dout(w_dff_A_EGkVELoi0_0),.din(w_dff_A_NaxIzPxG7_0),.clk(gclk));
	jdff dff_A_EGkVELoi0_0(.dout(w_dff_A_dpmFDk4l4_0),.din(w_dff_A_EGkVELoi0_0),.clk(gclk));
	jdff dff_A_dpmFDk4l4_0(.dout(w_dff_A_zWPEkxoE8_0),.din(w_dff_A_dpmFDk4l4_0),.clk(gclk));
	jdff dff_A_zWPEkxoE8_0(.dout(w_dff_A_S2fxXnOh9_0),.din(w_dff_A_zWPEkxoE8_0),.clk(gclk));
	jdff dff_A_S2fxXnOh9_0(.dout(w_dff_A_pUDoKapv1_0),.din(w_dff_A_S2fxXnOh9_0),.clk(gclk));
	jdff dff_A_pUDoKapv1_0(.dout(w_dff_A_he6AWlgo8_0),.din(w_dff_A_pUDoKapv1_0),.clk(gclk));
	jdff dff_A_he6AWlgo8_0(.dout(G6250gat),.din(w_dff_A_he6AWlgo8_0),.clk(gclk));
	jdff dff_A_ItMjlGlT1_2(.dout(w_dff_A_C1CdSTLN7_0),.din(w_dff_A_ItMjlGlT1_2),.clk(gclk));
	jdff dff_A_C1CdSTLN7_0(.dout(w_dff_A_W6uKVywC5_0),.din(w_dff_A_C1CdSTLN7_0),.clk(gclk));
	jdff dff_A_W6uKVywC5_0(.dout(w_dff_A_GG2KKa2p5_0),.din(w_dff_A_W6uKVywC5_0),.clk(gclk));
	jdff dff_A_GG2KKa2p5_0(.dout(w_dff_A_QFPb4j7j6_0),.din(w_dff_A_GG2KKa2p5_0),.clk(gclk));
	jdff dff_A_QFPb4j7j6_0(.dout(w_dff_A_C1glzCQw2_0),.din(w_dff_A_QFPb4j7j6_0),.clk(gclk));
	jdff dff_A_C1glzCQw2_0(.dout(w_dff_A_VtpZWgPZ6_0),.din(w_dff_A_C1glzCQw2_0),.clk(gclk));
	jdff dff_A_VtpZWgPZ6_0(.dout(G6260gat),.din(w_dff_A_VtpZWgPZ6_0),.clk(gclk));
	jdff dff_A_WJUS03tP8_2(.dout(w_dff_A_4TathcMT6_0),.din(w_dff_A_WJUS03tP8_2),.clk(gclk));
	jdff dff_A_4TathcMT6_0(.dout(w_dff_A_ifSQI7J07_0),.din(w_dff_A_4TathcMT6_0),.clk(gclk));
	jdff dff_A_ifSQI7J07_0(.dout(w_dff_A_6OgvdeOL1_0),.din(w_dff_A_ifSQI7J07_0),.clk(gclk));
	jdff dff_A_6OgvdeOL1_0(.dout(w_dff_A_MHHB6UYJ2_0),.din(w_dff_A_6OgvdeOL1_0),.clk(gclk));
	jdff dff_A_MHHB6UYJ2_0(.dout(G6270gat),.din(w_dff_A_MHHB6UYJ2_0),.clk(gclk));
	jdff dff_A_8IBM46XT7_2(.dout(w_dff_A_PeO9O6Ih5_0),.din(w_dff_A_8IBM46XT7_2),.clk(gclk));
	jdff dff_A_PeO9O6Ih5_0(.dout(w_dff_A_Axb5Z3Rn6_0),.din(w_dff_A_PeO9O6Ih5_0),.clk(gclk));
	jdff dff_A_Axb5Z3Rn6_0(.dout(G6280gat),.din(w_dff_A_Axb5Z3Rn6_0),.clk(gclk));
	jdff dff_A_Sal8trTP1_2(.dout(G6288gat),.din(w_dff_A_Sal8trTP1_2),.clk(gclk));
endmodule

